magic
tech sky130A
magscale 1 2
timestamp 1670026737
<< error_p >>
rect -478 1828 -465 1892
rect -410 1828 -395 1842
rect -376 1830 -363 1892
rect -295 1840 -142 1886
rect -313 1828 -121 1840
rect -42 1828 -29 1893
rect 53 1828 72 1892
rect 87 1828 93 1892
rect 102 1828 115 1892
rect 170 1828 185 1842
rect 204 1830 217 1892
rect 285 1840 438 1886
rect 267 1828 459 1840
rect 538 1828 551 1892
rect 633 1828 652 1892
rect 667 1828 673 1892
rect 682 1828 695 1892
rect 750 1828 765 1842
rect 784 1830 797 1892
rect 865 1840 1018 1886
rect 847 1828 1039 1840
rect 1118 1828 1131 1892
rect 1219 1878 1232 1892
rect 1213 1828 1232 1878
rect 1247 1828 1253 1844
rect 1262 1828 1275 1844
rect 1330 1828 1345 1842
rect 1364 1830 1377 1892
rect 1445 1840 1598 1886
rect 1427 1828 1619 1840
rect 1698 1828 1711 1892
rect 1793 1828 1812 1844
rect 1827 1828 1833 1844
rect 1842 1828 1855 1844
rect 1910 1828 1925 1842
rect 1944 1830 1957 1892
rect 2025 1840 2178 1886
rect 2007 1828 2199 1840
rect 2278 1828 2291 1892
rect 2373 1828 2392 1844
rect 2407 1828 2413 1844
rect 2422 1828 2435 1844
rect -541 1814 2479 1828
rect -478 1744 -465 1814
rect -420 1788 -391 1802
rect -338 1788 -322 1802
rect -284 1798 -278 1800
rect -271 1798 -163 1814
rect -156 1798 -150 1800
rect -142 1798 -127 1814
rect -61 1808 -42 1811
rect -420 1786 -322 1788
rect -295 1786 -127 1798
rect -112 1788 -96 1802
rect -61 1789 -39 1808
rect -29 1795 -13 1803
rect -39 1788 -33 1789
rect -30 1788 -1 1795
rect -112 1787 -1 1788
rect -112 1786 5 1787
rect -436 1778 -385 1786
rect -338 1778 -304 1786
rect -436 1766 -411 1778
rect -404 1766 -385 1778
rect -331 1776 -304 1778
rect -295 1776 -74 1786
rect -39 1783 -33 1786
rect -331 1772 -74 1776
rect -436 1758 -385 1766
rect -338 1758 -74 1772
rect -30 1778 5 1786
rect -484 1710 -465 1744
rect -420 1750 -391 1758
rect -420 1744 -403 1750
rect -420 1742 -386 1744
rect -338 1742 -322 1758
rect -321 1748 -113 1758
rect -112 1748 -96 1758
rect -48 1754 -33 1769
rect -30 1766 -29 1778
rect -22 1766 5 1778
rect -30 1758 5 1766
rect -30 1757 -1 1758
rect -310 1744 -96 1748
rect -295 1742 -96 1744
rect -61 1744 -48 1754
rect -30 1744 -13 1757
rect -61 1742 -13 1744
rect -419 1738 -386 1742
rect -423 1736 -386 1738
rect -423 1735 -356 1736
rect -423 1730 -392 1735
rect -386 1730 -356 1735
rect -423 1726 -356 1730
rect -450 1723 -356 1726
rect -450 1716 -401 1723
rect -450 1710 -420 1716
rect -401 1711 -396 1716
rect -484 1694 -404 1710
rect -392 1702 -356 1723
rect -295 1718 -106 1742
rect -61 1741 -14 1742
rect -48 1736 -14 1741
rect -280 1715 -106 1718
rect -287 1712 -106 1715
rect -78 1735 -14 1736
rect -484 1692 -465 1694
rect -450 1692 -416 1694
rect -484 1676 -404 1692
rect -484 1670 -465 1676
rect -494 1654 -465 1670
rect -450 1660 -420 1676
rect -392 1654 -386 1702
rect -383 1696 -364 1702
rect -349 1696 -319 1704
rect -383 1688 -319 1696
rect -383 1672 -303 1688
rect -287 1681 -225 1712
rect -209 1681 -147 1712
rect -78 1710 -29 1735
rect -14 1710 16 1726
rect -115 1696 -85 1704
rect -78 1702 32 1710
rect -115 1688 -70 1696
rect -383 1670 -364 1672
rect -349 1670 -303 1672
rect -383 1654 -303 1670
rect -276 1668 -241 1681
rect -200 1678 -163 1681
rect -200 1676 -158 1678
rect -271 1665 -241 1668
rect -262 1661 -255 1665
rect -255 1660 -254 1661
rect -296 1654 -286 1660
rect -500 1646 -459 1654
rect -500 1620 -485 1646
rect -478 1620 -459 1646
rect -395 1642 -364 1654
rect -349 1642 -246 1654
rect -234 1644 -208 1670
rect -193 1665 -163 1676
rect -131 1672 -69 1688
rect -131 1670 -85 1672
rect -131 1654 -69 1670
rect -57 1654 -51 1702
rect -48 1694 32 1702
rect -48 1692 -29 1694
rect -14 1692 20 1694
rect -48 1676 32 1692
rect -48 1654 -29 1676
rect -14 1660 16 1676
rect 44 1670 50 1744
rect 53 1670 72 1814
rect 87 1670 93 1814
rect 102 1744 115 1814
rect 160 1788 189 1802
rect 242 1788 258 1802
rect 296 1798 302 1800
rect 309 1798 417 1814
rect 424 1798 430 1800
rect 438 1798 453 1814
rect 519 1808 538 1811
rect 160 1786 258 1788
rect 285 1786 453 1798
rect 468 1788 484 1802
rect 519 1789 541 1808
rect 551 1795 567 1803
rect 541 1788 547 1789
rect 550 1788 579 1795
rect 468 1787 579 1788
rect 468 1786 585 1787
rect 144 1778 195 1786
rect 242 1778 276 1786
rect 144 1766 169 1778
rect 176 1766 195 1778
rect 249 1776 276 1778
rect 285 1776 506 1786
rect 541 1783 547 1786
rect 249 1772 506 1776
rect 144 1758 195 1766
rect 242 1758 506 1772
rect 550 1778 585 1786
rect 96 1710 115 1744
rect 160 1750 189 1758
rect 160 1744 177 1750
rect 160 1742 194 1744
rect 242 1742 258 1758
rect 259 1748 467 1758
rect 468 1748 484 1758
rect 532 1754 547 1769
rect 550 1766 551 1778
rect 558 1766 585 1778
rect 550 1758 585 1766
rect 550 1757 579 1758
rect 270 1744 484 1748
rect 285 1742 484 1744
rect 519 1744 532 1754
rect 550 1744 567 1757
rect 519 1742 567 1744
rect 161 1738 194 1742
rect 157 1736 194 1738
rect 157 1735 224 1736
rect 157 1730 188 1735
rect 194 1730 224 1735
rect 157 1726 224 1730
rect 130 1723 224 1726
rect 130 1716 179 1723
rect 130 1710 160 1716
rect 179 1711 184 1716
rect 96 1694 176 1710
rect 188 1702 224 1723
rect 285 1718 474 1742
rect 519 1741 566 1742
rect 532 1736 566 1741
rect 606 1736 622 1738
rect 300 1715 474 1718
rect 293 1712 474 1715
rect 502 1735 566 1736
rect 96 1692 115 1694
rect 130 1692 164 1694
rect 96 1676 176 1692
rect 96 1670 115 1676
rect -188 1644 -85 1654
rect -234 1642 -85 1644
rect -64 1642 -29 1654
rect -395 1640 -233 1642
rect -383 1620 -364 1640
rect -349 1638 -319 1640
rect -500 1612 -459 1620
rect -377 1616 -364 1620
rect -312 1624 -233 1640
rect -201 1640 -29 1642
rect -201 1624 -122 1640
rect -115 1638 -85 1640
rect -494 1602 -465 1612
rect -450 1602 -420 1616
rect -377 1602 -334 1616
rect -312 1612 -122 1624
rect -57 1620 -51 1640
rect -327 1602 -297 1612
rect -296 1602 -138 1612
rect -134 1602 -104 1612
rect -100 1602 -70 1616
rect -42 1602 -29 1640
rect 43 1654 72 1670
rect 86 1654 115 1670
rect 130 1660 160 1676
rect 188 1654 194 1702
rect 197 1696 216 1702
rect 231 1696 261 1704
rect 197 1688 261 1696
rect 197 1672 277 1688
rect 293 1681 355 1712
rect 371 1681 433 1712
rect 502 1710 551 1735
rect 596 1726 622 1736
rect 566 1710 622 1726
rect 465 1696 495 1704
rect 502 1702 612 1710
rect 465 1688 510 1696
rect 197 1670 216 1672
rect 231 1670 277 1672
rect 197 1654 277 1670
rect 304 1668 339 1681
rect 380 1678 417 1681
rect 380 1676 422 1678
rect 309 1665 339 1668
rect 318 1661 325 1665
rect 325 1660 326 1661
rect 284 1654 294 1660
rect 43 1646 78 1654
rect 43 1620 44 1646
rect 51 1620 78 1646
rect -14 1602 16 1616
rect 43 1612 78 1620
rect 80 1646 121 1654
rect 80 1620 95 1646
rect 102 1620 121 1646
rect 185 1642 216 1654
rect 231 1642 334 1654
rect 346 1644 372 1670
rect 387 1665 417 1676
rect 449 1672 511 1688
rect 449 1670 495 1672
rect 449 1654 511 1670
rect 523 1654 529 1702
rect 532 1694 612 1702
rect 532 1692 551 1694
rect 566 1692 600 1694
rect 532 1676 612 1692
rect 532 1654 551 1676
rect 566 1660 596 1676
rect 624 1670 630 1744
rect 633 1670 652 1814
rect 667 1670 673 1814
rect 682 1744 695 1814
rect 740 1788 769 1802
rect 822 1788 838 1802
rect 876 1798 882 1800
rect 889 1798 997 1814
rect 1004 1798 1010 1800
rect 1018 1798 1033 1814
rect 1099 1808 1118 1811
rect 740 1786 838 1788
rect 865 1786 1033 1798
rect 1048 1788 1064 1802
rect 1099 1789 1121 1808
rect 1131 1795 1147 1803
rect 1121 1788 1127 1789
rect 1130 1788 1159 1795
rect 1048 1787 1159 1788
rect 1048 1786 1165 1787
rect 724 1778 775 1786
rect 822 1778 856 1786
rect 724 1766 749 1778
rect 756 1766 775 1778
rect 829 1776 856 1778
rect 865 1776 1086 1786
rect 1121 1783 1127 1786
rect 829 1772 1086 1776
rect 724 1758 775 1766
rect 822 1758 1086 1772
rect 1130 1778 1165 1786
rect 676 1710 695 1744
rect 740 1750 769 1758
rect 740 1744 757 1750
rect 740 1742 774 1744
rect 822 1742 838 1758
rect 839 1748 1047 1758
rect 1048 1748 1064 1758
rect 1112 1754 1127 1769
rect 1130 1766 1131 1778
rect 1138 1766 1165 1778
rect 1130 1758 1165 1766
rect 1130 1757 1159 1758
rect 850 1744 1064 1748
rect 865 1742 1064 1744
rect 1099 1744 1112 1754
rect 1130 1744 1147 1757
rect 1099 1742 1147 1744
rect 741 1738 774 1742
rect 737 1736 774 1738
rect 737 1735 804 1736
rect 737 1730 768 1735
rect 774 1730 804 1735
rect 737 1726 804 1730
rect 710 1723 804 1726
rect 710 1716 759 1723
rect 710 1710 740 1716
rect 759 1711 764 1716
rect 676 1694 756 1710
rect 768 1702 804 1723
rect 865 1718 1054 1742
rect 1099 1741 1146 1742
rect 1112 1736 1146 1741
rect 880 1715 1054 1718
rect 873 1712 1054 1715
rect 1082 1735 1146 1736
rect 676 1692 695 1694
rect 710 1692 744 1694
rect 676 1676 756 1692
rect 676 1670 695 1676
rect 392 1644 495 1654
rect 346 1642 495 1644
rect 516 1642 551 1654
rect 185 1640 347 1642
rect 197 1620 216 1640
rect 231 1638 261 1640
rect 80 1612 121 1620
rect 203 1616 216 1620
rect 268 1624 347 1640
rect 379 1640 551 1642
rect 379 1624 458 1640
rect 465 1638 495 1640
rect 43 1602 72 1612
rect 86 1602 115 1612
rect 130 1602 160 1616
rect 203 1602 246 1616
rect 268 1612 458 1624
rect 523 1620 529 1640
rect 253 1602 283 1612
rect 284 1602 442 1612
rect 446 1602 476 1612
rect 480 1602 510 1616
rect 538 1602 551 1640
rect 623 1654 652 1670
rect 666 1654 695 1670
rect 710 1660 740 1676
rect 768 1654 774 1702
rect 777 1696 796 1702
rect 811 1696 841 1704
rect 777 1688 841 1696
rect 777 1672 857 1688
rect 873 1681 935 1712
rect 951 1681 1013 1712
rect 1082 1710 1131 1735
rect 1146 1710 1176 1728
rect 1045 1696 1075 1704
rect 1082 1702 1192 1710
rect 1045 1688 1090 1696
rect 777 1670 796 1672
rect 811 1670 857 1672
rect 777 1654 857 1670
rect 884 1668 919 1681
rect 960 1678 997 1681
rect 960 1676 1002 1678
rect 889 1665 919 1668
rect 898 1661 905 1665
rect 905 1660 906 1661
rect 864 1654 874 1660
rect 623 1646 658 1654
rect 623 1620 624 1646
rect 631 1620 658 1646
rect 566 1602 596 1616
rect 623 1612 658 1620
rect 660 1646 701 1654
rect 660 1620 675 1646
rect 682 1620 701 1646
rect 765 1642 796 1654
rect 811 1642 914 1654
rect 926 1644 952 1670
rect 967 1665 997 1676
rect 1029 1672 1091 1688
rect 1029 1670 1075 1672
rect 1029 1654 1091 1670
rect 1103 1654 1109 1702
rect 1112 1694 1192 1702
rect 1112 1692 1131 1694
rect 1146 1692 1180 1694
rect 1112 1677 1192 1692
rect 1112 1676 1198 1677
rect 1112 1654 1131 1676
rect 1146 1660 1176 1676
rect 1204 1670 1210 1744
rect 1213 1670 1232 1814
rect 1247 1670 1253 1814
rect 1262 1744 1275 1814
rect 1320 1788 1349 1802
rect 1402 1788 1418 1802
rect 1456 1798 1462 1800
rect 1469 1798 1577 1814
rect 1584 1798 1590 1800
rect 1598 1798 1613 1814
rect 1679 1808 1698 1811
rect 1320 1786 1418 1788
rect 1445 1786 1613 1798
rect 1628 1788 1644 1802
rect 1679 1789 1701 1808
rect 1711 1795 1727 1803
rect 1701 1788 1707 1789
rect 1710 1788 1739 1795
rect 1628 1787 1739 1788
rect 1628 1786 1745 1787
rect 1304 1778 1355 1786
rect 1402 1778 1436 1786
rect 1304 1766 1329 1778
rect 1336 1766 1355 1778
rect 1409 1776 1436 1778
rect 1445 1776 1666 1786
rect 1701 1783 1707 1786
rect 1409 1772 1666 1776
rect 1304 1758 1355 1766
rect 1402 1758 1666 1772
rect 1710 1778 1745 1786
rect 1256 1710 1275 1744
rect 1320 1750 1349 1758
rect 1320 1744 1337 1750
rect 1320 1742 1354 1744
rect 1402 1742 1418 1758
rect 1419 1748 1627 1758
rect 1628 1748 1644 1758
rect 1692 1754 1707 1769
rect 1710 1766 1711 1778
rect 1718 1766 1745 1778
rect 1710 1758 1745 1766
rect 1710 1757 1739 1758
rect 1430 1744 1644 1748
rect 1445 1742 1644 1744
rect 1679 1744 1692 1754
rect 1710 1744 1727 1757
rect 1679 1742 1727 1744
rect 1321 1738 1354 1742
rect 1317 1736 1354 1738
rect 1317 1735 1384 1736
rect 1317 1730 1348 1735
rect 1354 1730 1384 1735
rect 1317 1726 1384 1730
rect 1290 1723 1384 1726
rect 1290 1716 1339 1723
rect 1290 1710 1320 1716
rect 1339 1711 1344 1716
rect 1256 1694 1336 1710
rect 1348 1702 1384 1723
rect 1445 1718 1634 1742
rect 1679 1741 1726 1742
rect 1692 1736 1726 1741
rect 1766 1736 1782 1738
rect 1460 1715 1634 1718
rect 1453 1712 1634 1715
rect 1662 1735 1726 1736
rect 1256 1692 1275 1694
rect 1290 1692 1324 1694
rect 1256 1676 1336 1692
rect 1256 1670 1275 1676
rect 972 1644 1075 1654
rect 926 1642 1075 1644
rect 1096 1642 1131 1654
rect 765 1640 927 1642
rect 777 1620 796 1640
rect 811 1638 841 1640
rect 660 1612 701 1620
rect 783 1616 796 1620
rect 848 1624 927 1640
rect 959 1640 1131 1642
rect 959 1624 1038 1640
rect 1045 1638 1075 1640
rect 623 1602 652 1612
rect 666 1602 695 1612
rect 710 1602 740 1616
rect 783 1602 826 1616
rect 848 1612 1038 1624
rect 1103 1620 1109 1640
rect 833 1602 863 1612
rect 864 1602 1022 1612
rect 1026 1602 1056 1612
rect 1060 1602 1090 1616
rect 1118 1602 1131 1640
rect 1203 1654 1232 1670
rect 1246 1654 1275 1670
rect 1290 1660 1320 1676
rect 1348 1654 1354 1702
rect 1357 1696 1376 1702
rect 1391 1696 1421 1704
rect 1357 1688 1421 1696
rect 1357 1672 1437 1688
rect 1453 1681 1515 1712
rect 1531 1681 1593 1712
rect 1662 1710 1711 1735
rect 1756 1726 1782 1736
rect 1726 1710 1782 1726
rect 1625 1696 1655 1704
rect 1662 1702 1772 1710
rect 1625 1688 1670 1696
rect 1357 1670 1376 1672
rect 1391 1670 1437 1672
rect 1357 1654 1437 1670
rect 1464 1668 1499 1681
rect 1540 1678 1577 1681
rect 1540 1676 1582 1678
rect 1469 1665 1499 1668
rect 1478 1661 1485 1665
rect 1485 1660 1486 1661
rect 1444 1654 1454 1660
rect 1203 1646 1238 1654
rect 1203 1620 1204 1646
rect 1211 1620 1238 1646
rect 1146 1602 1176 1616
rect 1203 1612 1238 1620
rect 1240 1646 1281 1654
rect 1240 1620 1255 1646
rect 1262 1620 1281 1646
rect 1345 1642 1376 1654
rect 1391 1642 1494 1654
rect 1506 1644 1532 1670
rect 1547 1665 1577 1676
rect 1609 1672 1671 1688
rect 1609 1670 1655 1672
rect 1609 1654 1671 1670
rect 1683 1654 1689 1702
rect 1692 1694 1772 1702
rect 1692 1692 1711 1694
rect 1726 1692 1760 1694
rect 1692 1676 1772 1692
rect 1692 1654 1711 1676
rect 1726 1660 1756 1676
rect 1784 1670 1790 1744
rect 1793 1670 1812 1814
rect 1827 1670 1833 1814
rect 1842 1744 1855 1814
rect 1900 1788 1929 1802
rect 1982 1788 1998 1802
rect 2036 1798 2042 1800
rect 2049 1798 2157 1814
rect 2164 1798 2170 1800
rect 2178 1798 2193 1814
rect 2259 1808 2278 1811
rect 1900 1786 1998 1788
rect 2025 1786 2193 1798
rect 2208 1788 2224 1802
rect 2259 1789 2281 1808
rect 2291 1795 2307 1803
rect 2281 1788 2287 1789
rect 2290 1788 2319 1795
rect 2208 1787 2319 1788
rect 2208 1786 2325 1787
rect 1884 1778 1935 1786
rect 1982 1778 2016 1786
rect 1884 1766 1909 1778
rect 1916 1766 1935 1778
rect 1989 1776 2016 1778
rect 2025 1776 2246 1786
rect 2281 1783 2287 1786
rect 1989 1772 2246 1776
rect 1884 1758 1935 1766
rect 1982 1758 2246 1772
rect 2290 1778 2325 1786
rect 1836 1710 1855 1744
rect 1900 1750 1929 1758
rect 1900 1744 1917 1750
rect 1900 1742 1934 1744
rect 1982 1742 1998 1758
rect 1999 1748 2207 1758
rect 2208 1748 2224 1758
rect 2272 1754 2287 1769
rect 2290 1766 2291 1778
rect 2298 1766 2325 1778
rect 2290 1758 2325 1766
rect 2290 1757 2319 1758
rect 2010 1744 2224 1748
rect 2025 1742 2224 1744
rect 2259 1744 2272 1754
rect 2290 1744 2307 1757
rect 2259 1742 2307 1744
rect 1901 1738 1934 1742
rect 1897 1736 1934 1738
rect 1897 1735 1964 1736
rect 1897 1730 1928 1735
rect 1934 1730 1964 1735
rect 1897 1726 1964 1730
rect 1870 1723 1964 1726
rect 1870 1716 1919 1723
rect 1870 1710 1900 1716
rect 1919 1711 1924 1716
rect 1836 1694 1916 1710
rect 1928 1702 1964 1723
rect 2025 1718 2214 1742
rect 2259 1741 2306 1742
rect 2272 1736 2306 1741
rect 2040 1715 2214 1718
rect 2033 1712 2214 1715
rect 2242 1735 2306 1736
rect 1836 1692 1855 1694
rect 1870 1692 1904 1694
rect 1836 1676 1916 1692
rect 1836 1670 1855 1676
rect 1552 1644 1655 1654
rect 1506 1642 1655 1644
rect 1676 1642 1711 1654
rect 1345 1640 1507 1642
rect 1357 1620 1376 1640
rect 1391 1638 1421 1640
rect 1240 1612 1281 1620
rect 1363 1616 1376 1620
rect 1428 1624 1507 1640
rect 1539 1640 1711 1642
rect 1539 1624 1618 1640
rect 1625 1638 1655 1640
rect 1203 1602 1232 1612
rect 1246 1602 1275 1612
rect 1290 1602 1320 1616
rect 1363 1602 1406 1616
rect 1428 1612 1618 1624
rect 1683 1620 1689 1640
rect 1413 1602 1443 1612
rect 1444 1602 1602 1612
rect 1606 1602 1636 1612
rect 1640 1602 1670 1616
rect 1698 1602 1711 1640
rect 1783 1654 1812 1670
rect 1826 1654 1855 1670
rect 1870 1660 1900 1676
rect 1928 1654 1934 1702
rect 1937 1696 1956 1702
rect 1971 1696 2001 1704
rect 1937 1688 2001 1696
rect 1937 1672 2017 1688
rect 2033 1681 2095 1712
rect 2111 1681 2173 1712
rect 2242 1710 2291 1735
rect 2306 1710 2336 1728
rect 2205 1696 2235 1704
rect 2242 1702 2352 1710
rect 2205 1688 2250 1696
rect 1937 1670 1956 1672
rect 1971 1670 2017 1672
rect 1937 1654 2017 1670
rect 2044 1668 2079 1681
rect 2120 1678 2157 1681
rect 2120 1676 2162 1678
rect 2049 1665 2079 1668
rect 2058 1661 2065 1665
rect 2065 1660 2066 1661
rect 2024 1654 2034 1660
rect 1783 1646 1818 1654
rect 1783 1620 1784 1646
rect 1791 1620 1818 1646
rect 1726 1602 1756 1616
rect 1783 1612 1818 1620
rect 1820 1646 1861 1654
rect 1820 1620 1835 1646
rect 1842 1620 1861 1646
rect 1925 1642 1956 1654
rect 1971 1642 2074 1654
rect 2086 1644 2112 1670
rect 2127 1665 2157 1676
rect 2189 1672 2251 1688
rect 2189 1670 2235 1672
rect 2189 1654 2251 1670
rect 2263 1654 2269 1702
rect 2272 1694 2352 1702
rect 2272 1692 2291 1694
rect 2306 1692 2340 1694
rect 2272 1677 2352 1692
rect 2272 1676 2358 1677
rect 2272 1654 2291 1676
rect 2306 1660 2336 1676
rect 2364 1670 2370 1744
rect 2373 1670 2392 1814
rect 2407 1670 2413 1814
rect 2422 1744 2435 1814
rect 2464 1758 2479 1786
rect 2416 1710 2435 1744
rect 2477 1726 2479 1738
rect 2450 1710 2479 1726
rect 2416 1694 2479 1710
rect 2416 1692 2435 1694
rect 2450 1692 2479 1694
rect 2416 1676 2479 1692
rect 2416 1670 2435 1676
rect 2132 1644 2235 1654
rect 2086 1642 2235 1644
rect 2256 1642 2291 1654
rect 1925 1640 2087 1642
rect 1937 1620 1956 1640
rect 1971 1638 2001 1640
rect 1820 1612 1861 1620
rect 1943 1616 1956 1620
rect 2008 1624 2087 1640
rect 2119 1640 2291 1642
rect 2119 1624 2198 1640
rect 2205 1638 2235 1640
rect 1783 1602 1812 1612
rect 1826 1602 1855 1612
rect 1870 1602 1900 1616
rect 1943 1602 1986 1616
rect 2008 1612 2198 1624
rect 2263 1620 2269 1640
rect 1993 1602 2023 1612
rect 2024 1602 2182 1612
rect 2186 1602 2216 1612
rect 2220 1602 2250 1616
rect 2278 1602 2291 1640
rect 2363 1654 2392 1670
rect 2406 1654 2435 1670
rect 2450 1660 2479 1676
rect 2363 1646 2398 1654
rect 2363 1620 2364 1646
rect 2371 1620 2398 1646
rect 2306 1602 2336 1616
rect 2363 1612 2398 1620
rect 2400 1646 2441 1654
rect 2400 1620 2415 1646
rect 2422 1620 2441 1646
rect 2400 1612 2441 1620
rect 2363 1602 2392 1612
rect 2406 1602 2435 1612
rect 2450 1602 2479 1616
rect -541 1588 2479 1602
rect -478 1558 -465 1588
rect -450 1574 -420 1588
rect -377 1574 -334 1588
rect -327 1574 -107 1588
rect -100 1574 -70 1588
rect -410 1560 -395 1572
rect -376 1560 -363 1574
rect -295 1570 -142 1574
rect -413 1558 -391 1560
rect -313 1558 -121 1570
rect -42 1558 -29 1588
rect -14 1574 16 1588
rect 53 1558 72 1588
rect 87 1558 93 1588
rect 102 1558 115 1588
rect 130 1574 160 1588
rect 203 1574 246 1588
rect 253 1574 473 1588
rect 480 1574 510 1588
rect 170 1560 185 1572
rect 204 1560 217 1574
rect 285 1570 438 1574
rect 167 1558 189 1560
rect 267 1558 459 1570
rect 538 1558 551 1588
rect 566 1574 596 1588
rect 633 1558 652 1588
rect 667 1558 673 1588
rect 682 1558 695 1588
rect 710 1574 740 1588
rect 783 1574 826 1588
rect 833 1574 1053 1588
rect 1060 1574 1090 1588
rect 750 1560 765 1572
rect 784 1560 797 1574
rect 865 1570 1018 1574
rect 747 1558 769 1560
rect 847 1558 1039 1570
rect 1118 1558 1131 1588
rect 1146 1574 1176 1588
rect 1213 1558 1232 1588
rect 1247 1558 1253 1588
rect 1262 1558 1275 1588
rect 1290 1574 1320 1588
rect 1363 1574 1406 1588
rect 1413 1574 1633 1588
rect 1640 1574 1670 1588
rect 1330 1560 1345 1572
rect 1364 1560 1377 1574
rect 1445 1570 1598 1574
rect 1327 1558 1349 1560
rect 1427 1558 1619 1570
rect 1698 1558 1711 1588
rect 1726 1574 1756 1588
rect 1793 1558 1812 1588
rect 1827 1558 1833 1588
rect 1842 1558 1855 1588
rect 1870 1574 1900 1588
rect 1943 1574 1986 1588
rect 1993 1574 2213 1588
rect 2220 1574 2250 1588
rect 1910 1560 1925 1572
rect 1944 1560 1957 1574
rect 2025 1570 2178 1574
rect 1907 1558 1929 1560
rect 2007 1558 2199 1570
rect 2278 1558 2291 1588
rect 2306 1574 2336 1588
rect 2373 1558 2392 1588
rect 2407 1558 2413 1588
rect 2422 1558 2435 1588
rect 2450 1574 2479 1588
rect -541 1544 2479 1558
rect -478 1474 -465 1544
rect -413 1540 -391 1544
rect -420 1518 -391 1532
rect -338 1518 -322 1532
rect -284 1528 -278 1530
rect -271 1528 -163 1544
rect -156 1528 -150 1530
rect -142 1528 -127 1544
rect -61 1538 -42 1541
rect -420 1516 -322 1518
rect -295 1516 -127 1528
rect -112 1518 -96 1532
rect -61 1519 -39 1538
rect -29 1525 -13 1533
rect -39 1518 -33 1519
rect -30 1518 -1 1525
rect -112 1517 -1 1518
rect -112 1516 5 1517
rect -436 1508 -385 1516
rect -338 1508 -304 1516
rect -436 1496 -411 1508
rect -404 1496 -385 1508
rect -331 1506 -304 1508
rect -295 1506 -74 1516
rect -39 1513 -33 1516
rect -331 1502 -74 1506
rect -436 1488 -385 1496
rect -338 1488 -74 1502
rect -30 1508 5 1516
rect -484 1440 -465 1474
rect -420 1480 -391 1488
rect -420 1474 -403 1480
rect -420 1472 -386 1474
rect -338 1472 -322 1488
rect -321 1478 -113 1488
rect -112 1478 -96 1488
rect -48 1484 -33 1499
rect -30 1496 -29 1508
rect -22 1496 5 1508
rect -30 1488 5 1496
rect -30 1487 -1 1488
rect -310 1474 -96 1478
rect -295 1472 -96 1474
rect -61 1474 -48 1484
rect -30 1474 -13 1487
rect -61 1472 -13 1474
rect -419 1468 -386 1472
rect -423 1466 -386 1468
rect -423 1465 -356 1466
rect -423 1460 -392 1465
rect -386 1460 -356 1465
rect -423 1456 -356 1460
rect -450 1453 -356 1456
rect -450 1446 -401 1453
rect -450 1440 -420 1446
rect -401 1441 -396 1446
rect -484 1424 -404 1440
rect -392 1432 -356 1453
rect -295 1448 -106 1472
rect -61 1471 -14 1472
rect -48 1466 -14 1471
rect -280 1445 -106 1448
rect -287 1442 -106 1445
rect -78 1465 -14 1466
rect -484 1422 -465 1424
rect -450 1422 -416 1424
rect -484 1406 -404 1422
rect -484 1400 -465 1406
rect -494 1384 -465 1400
rect -450 1390 -420 1406
rect -392 1384 -386 1432
rect -383 1426 -364 1432
rect -349 1426 -319 1434
rect -383 1418 -319 1426
rect -383 1402 -303 1418
rect -287 1411 -225 1442
rect -209 1411 -147 1442
rect -78 1440 -29 1465
rect -14 1440 16 1458
rect -115 1426 -85 1434
rect -78 1432 32 1440
rect -115 1418 -70 1426
rect -383 1400 -364 1402
rect -349 1400 -303 1402
rect -383 1384 -303 1400
rect -276 1398 -241 1411
rect -200 1408 -163 1411
rect -200 1406 -158 1408
rect -271 1395 -241 1398
rect -262 1391 -255 1395
rect -255 1390 -254 1391
rect -296 1384 -286 1390
rect -500 1376 -459 1384
rect -500 1350 -485 1376
rect -478 1350 -459 1376
rect -395 1372 -364 1384
rect -349 1372 -246 1384
rect -234 1374 -208 1400
rect -193 1395 -163 1406
rect -131 1402 -69 1418
rect -131 1400 -85 1402
rect -131 1384 -69 1400
rect -57 1384 -51 1432
rect -48 1424 32 1432
rect -48 1422 -29 1424
rect -14 1422 20 1424
rect -48 1407 32 1422
rect -48 1406 38 1407
rect -48 1384 -29 1406
rect -14 1390 16 1406
rect 44 1400 50 1474
rect 53 1400 72 1544
rect 87 1400 93 1544
rect 102 1474 115 1544
rect 167 1540 189 1544
rect 160 1518 189 1532
rect 242 1518 258 1532
rect 296 1528 302 1530
rect 309 1528 417 1544
rect 424 1528 430 1530
rect 438 1528 453 1544
rect 519 1538 538 1541
rect 160 1516 258 1518
rect 285 1516 453 1528
rect 468 1518 484 1532
rect 519 1519 541 1538
rect 551 1525 567 1533
rect 541 1518 547 1519
rect 550 1518 579 1525
rect 468 1517 579 1518
rect 468 1516 585 1517
rect 144 1508 195 1516
rect 242 1508 276 1516
rect 144 1496 169 1508
rect 176 1496 195 1508
rect 249 1506 276 1508
rect 285 1506 506 1516
rect 541 1513 547 1516
rect 249 1502 506 1506
rect 144 1488 195 1496
rect 242 1488 506 1502
rect 550 1508 585 1516
rect 96 1440 115 1474
rect 160 1480 189 1488
rect 160 1474 177 1480
rect 160 1472 194 1474
rect 242 1472 258 1488
rect 259 1478 467 1488
rect 468 1478 484 1488
rect 532 1484 547 1499
rect 550 1496 551 1508
rect 558 1496 585 1508
rect 550 1488 585 1496
rect 550 1487 579 1488
rect 270 1474 484 1478
rect 285 1472 484 1474
rect 519 1474 532 1484
rect 550 1474 567 1487
rect 519 1472 567 1474
rect 161 1468 194 1472
rect 157 1466 194 1468
rect 157 1465 224 1466
rect 157 1460 188 1465
rect 194 1460 224 1465
rect 157 1456 224 1460
rect 130 1453 224 1456
rect 130 1446 179 1453
rect 130 1440 160 1446
rect 179 1441 184 1446
rect 96 1424 176 1440
rect 188 1432 224 1453
rect 285 1448 474 1472
rect 519 1471 566 1472
rect 532 1466 566 1471
rect 606 1466 622 1468
rect 300 1445 474 1448
rect 293 1442 474 1445
rect 502 1465 566 1466
rect 96 1422 115 1424
rect 130 1422 164 1424
rect 96 1406 176 1422
rect 96 1400 115 1406
rect -188 1374 -85 1384
rect -234 1372 -85 1374
rect -64 1372 -29 1384
rect -395 1370 -233 1372
rect -383 1352 -364 1370
rect -349 1368 -319 1370
rect -500 1342 -459 1350
rect -376 1346 -364 1352
rect -312 1354 -233 1370
rect -201 1370 -29 1372
rect -201 1354 -122 1370
rect -115 1368 -85 1370
rect -494 1332 -465 1342
rect -450 1332 -420 1346
rect -376 1332 -334 1346
rect -312 1342 -122 1354
rect -57 1350 -51 1370
rect -327 1332 -297 1342
rect -296 1332 -138 1342
rect -134 1332 -104 1342
rect -100 1332 -70 1346
rect -42 1332 -29 1370
rect 43 1384 72 1400
rect 86 1384 115 1400
rect 130 1390 160 1406
rect 188 1384 194 1432
rect 197 1426 216 1432
rect 231 1426 261 1434
rect 197 1418 261 1426
rect 197 1402 277 1418
rect 293 1411 355 1442
rect 371 1411 433 1442
rect 502 1440 551 1465
rect 596 1456 622 1466
rect 566 1440 622 1456
rect 465 1426 495 1434
rect 502 1432 612 1440
rect 465 1418 510 1426
rect 197 1400 216 1402
rect 231 1400 277 1402
rect 197 1384 277 1400
rect 304 1398 339 1411
rect 380 1408 417 1411
rect 380 1406 422 1408
rect 309 1395 339 1398
rect 318 1391 325 1395
rect 325 1390 326 1391
rect 284 1384 294 1390
rect 43 1376 78 1384
rect 43 1350 44 1376
rect 51 1350 78 1376
rect -14 1332 16 1346
rect 43 1342 78 1350
rect 80 1376 121 1384
rect 80 1350 95 1376
rect 102 1350 121 1376
rect 185 1372 216 1384
rect 231 1372 334 1384
rect 346 1374 372 1400
rect 387 1395 417 1406
rect 449 1402 511 1418
rect 449 1400 495 1402
rect 449 1384 511 1400
rect 523 1384 529 1432
rect 532 1424 612 1432
rect 532 1422 551 1424
rect 566 1422 600 1424
rect 532 1406 612 1422
rect 532 1384 551 1406
rect 566 1390 596 1406
rect 624 1400 630 1474
rect 633 1400 652 1544
rect 667 1400 673 1544
rect 682 1474 695 1544
rect 747 1540 769 1544
rect 740 1518 769 1532
rect 822 1518 838 1532
rect 876 1528 882 1530
rect 889 1528 997 1544
rect 1004 1528 1010 1530
rect 1018 1528 1033 1544
rect 1099 1538 1118 1541
rect 740 1516 838 1518
rect 865 1516 1033 1528
rect 1048 1518 1064 1532
rect 1099 1519 1121 1538
rect 1131 1525 1147 1533
rect 1121 1518 1127 1519
rect 1130 1518 1159 1525
rect 1048 1517 1159 1518
rect 1048 1516 1165 1517
rect 724 1508 775 1516
rect 822 1508 856 1516
rect 724 1496 749 1508
rect 756 1496 775 1508
rect 829 1506 856 1508
rect 865 1506 1086 1516
rect 1121 1513 1127 1516
rect 829 1502 1086 1506
rect 724 1488 775 1496
rect 822 1488 1086 1502
rect 1130 1508 1165 1516
rect 676 1440 695 1474
rect 740 1480 769 1488
rect 740 1474 757 1480
rect 740 1472 774 1474
rect 822 1472 838 1488
rect 839 1478 1047 1488
rect 1048 1478 1064 1488
rect 1112 1484 1127 1499
rect 1130 1496 1131 1508
rect 1138 1496 1165 1508
rect 1130 1488 1165 1496
rect 1130 1487 1159 1488
rect 850 1474 1064 1478
rect 865 1472 1064 1474
rect 1099 1474 1112 1484
rect 1130 1474 1147 1487
rect 1099 1472 1147 1474
rect 741 1468 774 1472
rect 737 1466 774 1468
rect 737 1465 804 1466
rect 737 1460 768 1465
rect 774 1460 804 1465
rect 737 1456 804 1460
rect 710 1453 804 1456
rect 710 1446 759 1453
rect 710 1440 740 1446
rect 759 1441 764 1446
rect 676 1424 756 1440
rect 768 1432 804 1453
rect 865 1448 1054 1472
rect 1099 1471 1146 1472
rect 1112 1466 1146 1471
rect 880 1445 1054 1448
rect 873 1442 1054 1445
rect 1082 1465 1146 1466
rect 676 1422 695 1424
rect 710 1422 744 1424
rect 676 1406 756 1422
rect 676 1400 695 1406
rect 392 1374 495 1384
rect 346 1372 495 1374
rect 516 1372 551 1384
rect 185 1370 347 1372
rect 197 1352 216 1370
rect 231 1368 261 1370
rect 80 1342 121 1350
rect 204 1346 216 1352
rect 268 1354 347 1370
rect 379 1370 551 1372
rect 379 1354 458 1370
rect 465 1368 495 1370
rect 43 1332 72 1342
rect 86 1332 115 1342
rect 130 1332 160 1346
rect 204 1332 246 1346
rect 268 1342 458 1354
rect 523 1350 529 1370
rect 253 1332 283 1342
rect 284 1332 442 1342
rect 446 1332 476 1342
rect 480 1332 510 1346
rect 538 1332 551 1370
rect 623 1384 652 1400
rect 666 1384 695 1400
rect 710 1390 740 1406
rect 768 1384 774 1432
rect 777 1426 796 1432
rect 811 1426 841 1434
rect 777 1418 841 1426
rect 777 1402 857 1418
rect 873 1411 935 1442
rect 951 1411 1013 1442
rect 1082 1440 1131 1465
rect 1146 1440 1176 1458
rect 1045 1426 1075 1434
rect 1082 1432 1192 1440
rect 1045 1418 1090 1426
rect 777 1400 796 1402
rect 811 1400 857 1402
rect 777 1384 857 1400
rect 884 1398 919 1411
rect 960 1408 997 1411
rect 960 1406 1002 1408
rect 889 1395 919 1398
rect 898 1391 905 1395
rect 905 1390 906 1391
rect 864 1384 874 1390
rect 623 1376 658 1384
rect 623 1350 624 1376
rect 631 1350 658 1376
rect 566 1332 596 1346
rect 623 1342 658 1350
rect 660 1376 701 1384
rect 660 1350 675 1376
rect 682 1350 701 1376
rect 765 1372 796 1384
rect 811 1372 914 1384
rect 926 1374 952 1400
rect 967 1395 997 1406
rect 1029 1402 1091 1418
rect 1029 1400 1075 1402
rect 1029 1384 1091 1400
rect 1103 1384 1109 1432
rect 1112 1424 1192 1432
rect 1112 1422 1131 1424
rect 1146 1422 1180 1424
rect 1112 1407 1192 1422
rect 1112 1406 1198 1407
rect 1112 1384 1131 1406
rect 1146 1390 1176 1406
rect 1204 1400 1210 1474
rect 1213 1400 1232 1544
rect 1247 1400 1253 1544
rect 1262 1474 1275 1544
rect 1327 1540 1349 1544
rect 1320 1518 1349 1532
rect 1402 1518 1418 1532
rect 1456 1528 1462 1530
rect 1469 1528 1577 1544
rect 1584 1528 1590 1530
rect 1598 1528 1613 1544
rect 1679 1538 1698 1541
rect 1320 1516 1418 1518
rect 1445 1516 1613 1528
rect 1628 1518 1644 1532
rect 1679 1519 1701 1538
rect 1711 1525 1727 1533
rect 1701 1518 1707 1519
rect 1710 1518 1739 1525
rect 1628 1517 1739 1518
rect 1628 1516 1745 1517
rect 1304 1508 1355 1516
rect 1402 1508 1436 1516
rect 1304 1496 1329 1508
rect 1336 1496 1355 1508
rect 1409 1506 1436 1508
rect 1445 1506 1666 1516
rect 1701 1513 1707 1516
rect 1409 1502 1666 1506
rect 1304 1488 1355 1496
rect 1402 1488 1666 1502
rect 1710 1508 1745 1516
rect 1256 1440 1275 1474
rect 1320 1480 1349 1488
rect 1320 1474 1337 1480
rect 1320 1472 1354 1474
rect 1402 1472 1418 1488
rect 1419 1478 1627 1488
rect 1628 1478 1644 1488
rect 1692 1484 1707 1499
rect 1710 1496 1711 1508
rect 1718 1496 1745 1508
rect 1710 1488 1745 1496
rect 1710 1487 1739 1488
rect 1430 1474 1644 1478
rect 1445 1472 1644 1474
rect 1679 1474 1692 1484
rect 1710 1474 1727 1487
rect 1679 1472 1727 1474
rect 1321 1468 1354 1472
rect 1317 1466 1354 1468
rect 1317 1465 1384 1466
rect 1317 1460 1348 1465
rect 1354 1460 1384 1465
rect 1317 1456 1384 1460
rect 1290 1453 1384 1456
rect 1290 1446 1339 1453
rect 1290 1440 1320 1446
rect 1339 1441 1344 1446
rect 1256 1424 1336 1440
rect 1348 1432 1384 1453
rect 1445 1448 1634 1472
rect 1679 1471 1726 1472
rect 1692 1466 1726 1471
rect 1766 1466 1782 1468
rect 1460 1445 1634 1448
rect 1453 1442 1634 1445
rect 1662 1465 1726 1466
rect 1256 1422 1275 1424
rect 1290 1422 1324 1424
rect 1256 1406 1336 1422
rect 1256 1400 1275 1406
rect 972 1374 1075 1384
rect 926 1372 1075 1374
rect 1096 1372 1131 1384
rect 765 1370 927 1372
rect 777 1352 796 1370
rect 811 1368 841 1370
rect 660 1342 701 1350
rect 784 1346 796 1352
rect 848 1354 927 1370
rect 959 1370 1131 1372
rect 959 1354 1038 1370
rect 1045 1368 1075 1370
rect 623 1332 652 1342
rect 666 1332 695 1342
rect 710 1332 740 1346
rect 784 1332 826 1346
rect 848 1342 1038 1354
rect 1103 1350 1109 1370
rect 833 1332 863 1342
rect 864 1332 1022 1342
rect 1026 1332 1056 1342
rect 1060 1332 1090 1346
rect 1118 1332 1131 1370
rect 1203 1384 1232 1400
rect 1246 1384 1275 1400
rect 1290 1390 1320 1406
rect 1348 1384 1354 1432
rect 1357 1426 1376 1432
rect 1391 1426 1421 1434
rect 1357 1418 1421 1426
rect 1357 1402 1437 1418
rect 1453 1411 1515 1442
rect 1531 1411 1593 1442
rect 1662 1440 1711 1465
rect 1756 1456 1782 1466
rect 1726 1440 1782 1456
rect 1625 1426 1655 1434
rect 1662 1432 1772 1440
rect 1625 1418 1670 1426
rect 1357 1400 1376 1402
rect 1391 1400 1437 1402
rect 1357 1384 1437 1400
rect 1464 1398 1499 1411
rect 1540 1408 1577 1411
rect 1540 1406 1582 1408
rect 1469 1395 1499 1398
rect 1478 1391 1485 1395
rect 1485 1390 1486 1391
rect 1444 1384 1454 1390
rect 1203 1376 1238 1384
rect 1203 1350 1204 1376
rect 1211 1350 1238 1376
rect 1146 1332 1176 1346
rect 1203 1342 1238 1350
rect 1240 1376 1281 1384
rect 1240 1350 1255 1376
rect 1262 1350 1281 1376
rect 1345 1372 1376 1384
rect 1391 1372 1494 1384
rect 1506 1374 1532 1400
rect 1547 1395 1577 1406
rect 1609 1402 1671 1418
rect 1609 1400 1655 1402
rect 1609 1384 1671 1400
rect 1683 1384 1689 1432
rect 1692 1424 1772 1432
rect 1692 1422 1711 1424
rect 1726 1422 1760 1424
rect 1692 1406 1772 1422
rect 1692 1384 1711 1406
rect 1726 1390 1756 1406
rect 1784 1400 1790 1474
rect 1793 1400 1812 1544
rect 1827 1400 1833 1544
rect 1842 1474 1855 1544
rect 1907 1540 1929 1544
rect 1900 1518 1929 1532
rect 1982 1518 1998 1532
rect 2036 1528 2042 1530
rect 2049 1528 2157 1544
rect 2164 1528 2170 1530
rect 2178 1528 2193 1544
rect 2259 1538 2278 1541
rect 1900 1516 1998 1518
rect 2025 1516 2193 1528
rect 2208 1518 2224 1532
rect 2259 1519 2281 1538
rect 2291 1525 2307 1533
rect 2281 1518 2287 1519
rect 2290 1518 2319 1525
rect 2208 1517 2319 1518
rect 2208 1516 2325 1517
rect 1884 1508 1935 1516
rect 1982 1508 2016 1516
rect 1884 1496 1909 1508
rect 1916 1496 1935 1508
rect 1989 1506 2016 1508
rect 2025 1506 2246 1516
rect 2281 1513 2287 1516
rect 1989 1502 2246 1506
rect 1884 1488 1935 1496
rect 1982 1488 2246 1502
rect 2290 1508 2325 1516
rect 1836 1440 1855 1474
rect 1900 1480 1929 1488
rect 1900 1474 1917 1480
rect 1900 1472 1934 1474
rect 1982 1472 1998 1488
rect 1999 1478 2207 1488
rect 2208 1478 2224 1488
rect 2272 1484 2287 1499
rect 2290 1496 2291 1508
rect 2298 1496 2325 1508
rect 2290 1488 2325 1496
rect 2290 1487 2319 1488
rect 2010 1474 2224 1478
rect 2025 1472 2224 1474
rect 2259 1474 2272 1484
rect 2290 1474 2307 1487
rect 2259 1472 2307 1474
rect 1901 1468 1934 1472
rect 1897 1466 1934 1468
rect 1897 1465 1964 1466
rect 1897 1460 1928 1465
rect 1934 1460 1964 1465
rect 1897 1456 1964 1460
rect 1870 1453 1964 1456
rect 1870 1446 1919 1453
rect 1870 1440 1900 1446
rect 1919 1441 1924 1446
rect 1836 1424 1916 1440
rect 1928 1432 1964 1453
rect 2025 1448 2214 1472
rect 2259 1471 2306 1472
rect 2272 1466 2306 1471
rect 2040 1445 2214 1448
rect 2033 1442 2214 1445
rect 2242 1465 2306 1466
rect 1836 1422 1855 1424
rect 1870 1422 1904 1424
rect 1836 1406 1916 1422
rect 1836 1400 1855 1406
rect 1552 1374 1655 1384
rect 1506 1372 1655 1374
rect 1676 1372 1711 1384
rect 1345 1370 1507 1372
rect 1357 1352 1376 1370
rect 1391 1368 1421 1370
rect 1240 1342 1281 1350
rect 1364 1346 1376 1352
rect 1428 1354 1507 1370
rect 1539 1370 1711 1372
rect 1539 1354 1618 1370
rect 1625 1368 1655 1370
rect 1203 1332 1232 1342
rect 1246 1332 1275 1342
rect 1290 1332 1320 1346
rect 1364 1332 1406 1346
rect 1428 1342 1618 1354
rect 1683 1350 1689 1370
rect 1413 1332 1443 1342
rect 1444 1332 1602 1342
rect 1606 1332 1636 1342
rect 1640 1332 1670 1346
rect 1698 1332 1711 1370
rect 1783 1384 1812 1400
rect 1826 1384 1855 1400
rect 1870 1390 1900 1406
rect 1928 1384 1934 1432
rect 1937 1426 1956 1432
rect 1971 1426 2001 1434
rect 1937 1418 2001 1426
rect 1937 1402 2017 1418
rect 2033 1411 2095 1442
rect 2111 1411 2173 1442
rect 2242 1440 2291 1465
rect 2306 1440 2336 1458
rect 2205 1426 2235 1434
rect 2242 1432 2352 1440
rect 2205 1418 2250 1426
rect 1937 1400 1956 1402
rect 1971 1400 2017 1402
rect 1937 1384 2017 1400
rect 2044 1398 2079 1411
rect 2120 1408 2157 1411
rect 2120 1406 2162 1408
rect 2049 1395 2079 1398
rect 2058 1391 2065 1395
rect 2065 1390 2066 1391
rect 2024 1384 2034 1390
rect 1783 1376 1818 1384
rect 1783 1350 1784 1376
rect 1791 1350 1818 1376
rect 1726 1332 1756 1346
rect 1783 1342 1818 1350
rect 1820 1376 1861 1384
rect 1820 1350 1835 1376
rect 1842 1350 1861 1376
rect 1925 1372 1956 1384
rect 1971 1372 2074 1384
rect 2086 1374 2112 1400
rect 2127 1395 2157 1406
rect 2189 1402 2251 1418
rect 2189 1400 2235 1402
rect 2189 1384 2251 1400
rect 2263 1384 2269 1432
rect 2272 1424 2352 1432
rect 2272 1422 2291 1424
rect 2306 1422 2340 1424
rect 2272 1407 2352 1422
rect 2272 1406 2358 1407
rect 2272 1384 2291 1406
rect 2306 1390 2336 1406
rect 2364 1400 2370 1474
rect 2373 1400 2392 1544
rect 2407 1400 2413 1544
rect 2422 1474 2435 1544
rect 2464 1488 2479 1516
rect 2416 1440 2435 1474
rect 2477 1456 2479 1468
rect 2450 1440 2479 1456
rect 2416 1424 2479 1440
rect 2416 1422 2435 1424
rect 2450 1422 2479 1424
rect 2416 1406 2479 1422
rect 2416 1400 2435 1406
rect 2132 1374 2235 1384
rect 2086 1372 2235 1374
rect 2256 1372 2291 1384
rect 1925 1370 2087 1372
rect 1937 1352 1956 1370
rect 1971 1368 2001 1370
rect 1820 1342 1861 1350
rect 1944 1346 1956 1352
rect 2008 1354 2087 1370
rect 2119 1370 2291 1372
rect 2119 1354 2198 1370
rect 2205 1368 2235 1370
rect 1783 1332 1812 1342
rect 1826 1332 1855 1342
rect 1870 1332 1900 1346
rect 1944 1332 1986 1346
rect 2008 1342 2198 1354
rect 2263 1350 2269 1370
rect 1993 1332 2023 1342
rect 2024 1332 2182 1342
rect 2186 1332 2216 1342
rect 2220 1332 2250 1346
rect 2278 1332 2291 1370
rect 2363 1384 2392 1400
rect 2406 1384 2435 1400
rect 2450 1390 2479 1406
rect 2363 1376 2398 1384
rect 2363 1350 2364 1376
rect 2371 1350 2398 1376
rect 2306 1332 2336 1346
rect 2363 1342 2398 1350
rect 2400 1376 2441 1384
rect 2400 1350 2415 1376
rect 2422 1350 2441 1376
rect 2400 1342 2441 1350
rect 2363 1332 2392 1342
rect 2406 1332 2435 1342
rect 2450 1332 2479 1346
rect -541 1318 2479 1332
rect -478 1288 -465 1318
rect -450 1304 -420 1318
rect -376 1304 -334 1318
rect -327 1304 -107 1318
rect -100 1304 -70 1318
rect -410 1290 -395 1302
rect -376 1290 -363 1304
rect -295 1300 -142 1304
rect -413 1288 -391 1290
rect -313 1288 -121 1300
rect -42 1288 -29 1318
rect -14 1304 16 1318
rect 53 1288 72 1318
rect 87 1288 93 1318
rect 102 1288 115 1318
rect 130 1304 160 1318
rect 204 1304 246 1318
rect 253 1304 473 1318
rect 480 1304 510 1318
rect 170 1290 185 1302
rect 204 1290 217 1304
rect 285 1300 438 1304
rect 167 1288 189 1290
rect 267 1288 459 1300
rect 538 1288 551 1318
rect 566 1304 596 1318
rect 633 1288 652 1318
rect 667 1288 673 1318
rect 682 1288 695 1318
rect 710 1304 740 1318
rect 784 1304 826 1318
rect 833 1304 1053 1318
rect 1060 1304 1090 1318
rect 750 1290 765 1302
rect 784 1290 797 1304
rect 865 1300 1018 1304
rect 747 1288 769 1290
rect 847 1288 1039 1300
rect 1118 1288 1131 1318
rect 1146 1304 1176 1318
rect 1213 1288 1232 1318
rect 1247 1288 1253 1318
rect 1262 1288 1275 1318
rect 1290 1304 1320 1318
rect 1364 1304 1406 1318
rect 1413 1304 1633 1318
rect 1640 1304 1670 1318
rect 1330 1290 1345 1302
rect 1364 1290 1377 1304
rect 1445 1300 1598 1304
rect 1327 1288 1349 1290
rect 1427 1288 1619 1300
rect 1698 1288 1711 1318
rect 1726 1304 1756 1318
rect 1793 1288 1812 1318
rect 1827 1288 1833 1318
rect 1842 1288 1855 1318
rect 1870 1304 1900 1318
rect 1944 1304 1986 1318
rect 1993 1304 2213 1318
rect 2220 1304 2250 1318
rect 1910 1290 1925 1302
rect 1944 1290 1957 1304
rect 2025 1300 2178 1304
rect 1907 1288 1929 1290
rect 2007 1288 2199 1300
rect 2278 1288 2291 1318
rect 2306 1304 2336 1318
rect 2373 1288 2392 1318
rect 2407 1288 2413 1318
rect 2422 1288 2435 1318
rect 2450 1304 2479 1318
rect -541 1274 2479 1288
rect -478 1204 -465 1274
rect -413 1270 -391 1274
rect -420 1248 -391 1262
rect -338 1248 -322 1262
rect -284 1258 -278 1260
rect -271 1258 -163 1274
rect -156 1258 -150 1260
rect -142 1258 -127 1274
rect -61 1268 -42 1271
rect -420 1246 -322 1248
rect -295 1246 -127 1258
rect -112 1248 -96 1262
rect -61 1249 -39 1268
rect -29 1255 -13 1263
rect -39 1248 -33 1249
rect -30 1248 -1 1255
rect -112 1247 -1 1248
rect -112 1246 5 1247
rect -436 1238 -385 1246
rect -338 1238 -304 1246
rect -436 1226 -411 1238
rect -404 1226 -385 1238
rect -331 1236 -304 1238
rect -295 1236 -74 1246
rect -39 1243 -33 1246
rect -331 1232 -74 1236
rect -436 1218 -385 1226
rect -338 1218 -74 1232
rect -30 1238 5 1246
rect -484 1170 -465 1204
rect -420 1210 -391 1218
rect -420 1204 -403 1210
rect -420 1202 -386 1204
rect -338 1202 -322 1218
rect -321 1208 -113 1218
rect -112 1208 -96 1218
rect -48 1214 -33 1229
rect -30 1226 -29 1238
rect -22 1226 5 1238
rect -30 1218 5 1226
rect -30 1217 -1 1218
rect -310 1204 -96 1208
rect -295 1202 -96 1204
rect -61 1204 -48 1214
rect -30 1204 -13 1217
rect -61 1202 -13 1204
rect -419 1198 -386 1202
rect -423 1196 -386 1198
rect -423 1195 -356 1196
rect -423 1190 -392 1195
rect -386 1190 -356 1195
rect -423 1186 -356 1190
rect -450 1183 -356 1186
rect -450 1176 -401 1183
rect -450 1170 -420 1176
rect -401 1171 -396 1176
rect -484 1154 -404 1170
rect -392 1162 -356 1183
rect -295 1178 -106 1202
rect -61 1201 -14 1202
rect -48 1196 -14 1201
rect -280 1175 -106 1178
rect -287 1172 -106 1175
rect -78 1195 -14 1196
rect -484 1152 -465 1154
rect -450 1152 -416 1154
rect -484 1136 -404 1152
rect -484 1130 -465 1136
rect -494 1114 -465 1130
rect -450 1120 -420 1136
rect -392 1114 -386 1162
rect -383 1156 -364 1162
rect -349 1156 -319 1164
rect -383 1148 -319 1156
rect -383 1132 -303 1148
rect -287 1141 -225 1172
rect -209 1141 -147 1172
rect -78 1170 -29 1195
rect -14 1170 16 1188
rect -115 1156 -85 1164
rect -78 1162 32 1170
rect -115 1148 -70 1156
rect -383 1130 -364 1132
rect -349 1130 -303 1132
rect -383 1114 -303 1130
rect -276 1128 -241 1141
rect -200 1138 -163 1141
rect -200 1136 -158 1138
rect -271 1125 -241 1128
rect -262 1121 -255 1125
rect -255 1120 -254 1121
rect -296 1114 -286 1120
rect -500 1106 -459 1114
rect -500 1080 -485 1106
rect -478 1080 -459 1106
rect -395 1102 -364 1114
rect -349 1102 -246 1114
rect -234 1104 -208 1130
rect -193 1125 -163 1136
rect -131 1132 -69 1148
rect -131 1130 -85 1132
rect -131 1114 -69 1130
rect -57 1114 -51 1162
rect -48 1154 32 1162
rect -48 1152 -29 1154
rect -14 1152 20 1154
rect -48 1137 32 1152
rect -48 1136 38 1137
rect -48 1114 -29 1136
rect -14 1120 16 1136
rect 44 1130 50 1204
rect 53 1130 72 1274
rect 87 1130 93 1274
rect 102 1204 115 1274
rect 167 1270 189 1274
rect 160 1248 189 1262
rect 242 1248 258 1262
rect 296 1258 302 1260
rect 309 1258 417 1274
rect 424 1258 430 1260
rect 438 1258 453 1274
rect 519 1268 538 1271
rect 160 1246 258 1248
rect 285 1246 453 1258
rect 468 1248 484 1262
rect 519 1249 541 1268
rect 551 1255 567 1263
rect 541 1248 547 1249
rect 550 1248 579 1255
rect 468 1247 579 1248
rect 468 1246 585 1247
rect 144 1238 195 1246
rect 242 1238 276 1246
rect 144 1226 169 1238
rect 176 1226 195 1238
rect 249 1236 276 1238
rect 285 1236 506 1246
rect 541 1243 547 1246
rect 249 1232 506 1236
rect 144 1218 195 1226
rect 242 1218 506 1232
rect 550 1238 585 1246
rect 96 1170 115 1204
rect 160 1210 189 1218
rect 160 1204 177 1210
rect 160 1202 194 1204
rect 242 1202 258 1218
rect 259 1208 467 1218
rect 468 1208 484 1218
rect 532 1214 547 1229
rect 550 1226 551 1238
rect 558 1226 585 1238
rect 550 1218 585 1226
rect 550 1217 579 1218
rect 270 1204 484 1208
rect 285 1202 484 1204
rect 519 1204 532 1214
rect 550 1204 567 1217
rect 519 1202 567 1204
rect 161 1198 194 1202
rect 157 1196 194 1198
rect 157 1195 224 1196
rect 157 1190 188 1195
rect 194 1190 224 1195
rect 157 1186 224 1190
rect 130 1183 224 1186
rect 130 1176 179 1183
rect 130 1170 160 1176
rect 179 1171 184 1176
rect 96 1154 176 1170
rect 188 1162 224 1183
rect 285 1178 474 1202
rect 519 1201 566 1202
rect 532 1196 566 1201
rect 606 1196 622 1198
rect 300 1175 474 1178
rect 293 1172 474 1175
rect 502 1195 566 1196
rect 96 1152 115 1154
rect 130 1152 164 1154
rect 96 1136 176 1152
rect 96 1130 115 1136
rect -188 1104 -85 1114
rect -234 1102 -85 1104
rect -64 1102 -29 1114
rect -395 1100 -233 1102
rect -383 1080 -364 1100
rect -349 1098 -319 1100
rect -500 1072 -459 1080
rect -377 1076 -364 1080
rect -312 1084 -233 1100
rect -201 1100 -29 1102
rect -201 1084 -122 1100
rect -115 1098 -85 1100
rect -494 1062 -465 1072
rect -450 1062 -420 1076
rect -377 1062 -334 1076
rect -312 1072 -122 1084
rect -57 1080 -51 1100
rect -327 1062 -297 1072
rect -296 1062 -138 1072
rect -134 1062 -104 1072
rect -100 1062 -70 1076
rect -42 1062 -29 1100
rect 43 1114 72 1130
rect 86 1114 115 1130
rect 130 1120 160 1136
rect 188 1114 194 1162
rect 197 1156 216 1162
rect 231 1156 261 1164
rect 197 1148 261 1156
rect 197 1132 277 1148
rect 293 1141 355 1172
rect 371 1141 433 1172
rect 502 1170 551 1195
rect 596 1186 622 1196
rect 566 1170 622 1186
rect 465 1156 495 1164
rect 502 1162 612 1170
rect 465 1148 510 1156
rect 197 1130 216 1132
rect 231 1130 277 1132
rect 197 1114 277 1130
rect 304 1128 339 1141
rect 380 1138 417 1141
rect 380 1136 422 1138
rect 309 1125 339 1128
rect 318 1121 325 1125
rect 325 1120 326 1121
rect 284 1114 294 1120
rect 43 1106 78 1114
rect 43 1080 44 1106
rect 51 1080 78 1106
rect -14 1062 16 1076
rect 43 1072 78 1080
rect 80 1106 121 1114
rect 80 1080 95 1106
rect 102 1080 121 1106
rect 185 1102 216 1114
rect 231 1102 334 1114
rect 346 1104 372 1130
rect 387 1125 417 1136
rect 449 1132 511 1148
rect 449 1130 495 1132
rect 449 1114 511 1130
rect 523 1114 529 1162
rect 532 1154 612 1162
rect 532 1152 551 1154
rect 566 1152 600 1154
rect 532 1136 612 1152
rect 532 1114 551 1136
rect 566 1120 596 1136
rect 624 1130 630 1204
rect 633 1130 652 1274
rect 667 1130 673 1274
rect 682 1204 695 1274
rect 747 1270 769 1274
rect 740 1248 769 1262
rect 822 1248 838 1262
rect 876 1258 882 1260
rect 889 1258 997 1274
rect 1004 1258 1010 1260
rect 1018 1258 1033 1274
rect 1099 1268 1118 1271
rect 740 1246 838 1248
rect 865 1246 1033 1258
rect 1048 1248 1064 1262
rect 1099 1249 1121 1268
rect 1131 1255 1147 1263
rect 1121 1248 1127 1249
rect 1130 1248 1159 1255
rect 1048 1247 1159 1248
rect 1048 1246 1165 1247
rect 724 1238 775 1246
rect 822 1238 856 1246
rect 724 1226 749 1238
rect 756 1226 775 1238
rect 829 1236 856 1238
rect 865 1236 1086 1246
rect 1121 1243 1127 1246
rect 829 1232 1086 1236
rect 724 1218 775 1226
rect 822 1218 1086 1232
rect 1130 1238 1165 1246
rect 676 1170 695 1204
rect 740 1210 769 1218
rect 740 1204 757 1210
rect 740 1202 774 1204
rect 822 1202 838 1218
rect 839 1208 1047 1218
rect 1048 1208 1064 1218
rect 1112 1214 1127 1229
rect 1130 1226 1131 1238
rect 1138 1226 1165 1238
rect 1130 1218 1165 1226
rect 1130 1217 1159 1218
rect 850 1204 1064 1208
rect 865 1202 1064 1204
rect 1099 1204 1112 1214
rect 1130 1204 1147 1217
rect 1099 1202 1147 1204
rect 741 1198 774 1202
rect 737 1196 774 1198
rect 737 1195 804 1196
rect 737 1190 768 1195
rect 774 1190 804 1195
rect 737 1186 804 1190
rect 710 1183 804 1186
rect 710 1176 759 1183
rect 710 1170 740 1176
rect 759 1171 764 1176
rect 676 1154 756 1170
rect 768 1162 804 1183
rect 865 1178 1054 1202
rect 1099 1201 1146 1202
rect 1112 1196 1146 1201
rect 880 1175 1054 1178
rect 873 1172 1054 1175
rect 1082 1195 1146 1196
rect 676 1152 695 1154
rect 710 1152 744 1154
rect 676 1136 756 1152
rect 676 1130 695 1136
rect 392 1104 495 1114
rect 346 1102 495 1104
rect 516 1102 551 1114
rect 185 1100 347 1102
rect 197 1080 216 1100
rect 231 1098 261 1100
rect 80 1072 121 1080
rect 203 1076 216 1080
rect 268 1084 347 1100
rect 379 1100 551 1102
rect 379 1084 458 1100
rect 465 1098 495 1100
rect 43 1062 72 1072
rect 86 1062 115 1072
rect 130 1062 160 1076
rect 203 1062 246 1076
rect 268 1072 458 1084
rect 523 1080 529 1100
rect 253 1062 283 1072
rect 284 1062 442 1072
rect 446 1062 476 1072
rect 480 1062 510 1076
rect 538 1062 551 1100
rect 623 1114 652 1130
rect 666 1114 695 1130
rect 710 1120 740 1136
rect 768 1114 774 1162
rect 777 1156 796 1162
rect 811 1156 841 1164
rect 777 1148 841 1156
rect 777 1132 857 1148
rect 873 1141 935 1172
rect 951 1141 1013 1172
rect 1082 1170 1131 1195
rect 1146 1170 1176 1188
rect 1045 1156 1075 1164
rect 1082 1162 1192 1170
rect 1045 1148 1090 1156
rect 777 1130 796 1132
rect 811 1130 857 1132
rect 777 1114 857 1130
rect 884 1128 919 1141
rect 960 1138 997 1141
rect 960 1136 1002 1138
rect 889 1125 919 1128
rect 898 1121 905 1125
rect 905 1120 906 1121
rect 864 1114 874 1120
rect 623 1106 658 1114
rect 623 1080 624 1106
rect 631 1080 658 1106
rect 566 1062 596 1076
rect 623 1072 658 1080
rect 660 1106 701 1114
rect 660 1080 675 1106
rect 682 1080 701 1106
rect 765 1102 796 1114
rect 811 1102 914 1114
rect 926 1104 952 1130
rect 967 1125 997 1136
rect 1029 1132 1091 1148
rect 1029 1130 1075 1132
rect 1029 1114 1091 1130
rect 1103 1114 1109 1162
rect 1112 1154 1192 1162
rect 1112 1152 1131 1154
rect 1146 1152 1180 1154
rect 1112 1137 1192 1152
rect 1112 1136 1198 1137
rect 1112 1114 1131 1136
rect 1146 1120 1176 1136
rect 1204 1130 1210 1204
rect 1213 1130 1232 1274
rect 1247 1130 1253 1274
rect 1262 1204 1275 1274
rect 1327 1270 1349 1274
rect 1320 1248 1349 1262
rect 1402 1248 1418 1262
rect 1456 1258 1462 1260
rect 1469 1258 1577 1274
rect 1584 1258 1590 1260
rect 1598 1258 1613 1274
rect 1679 1268 1698 1271
rect 1320 1246 1418 1248
rect 1445 1246 1613 1258
rect 1628 1248 1644 1262
rect 1679 1249 1701 1268
rect 1711 1255 1727 1263
rect 1701 1248 1707 1249
rect 1710 1248 1739 1255
rect 1628 1247 1739 1248
rect 1628 1246 1745 1247
rect 1304 1238 1355 1246
rect 1402 1238 1436 1246
rect 1304 1226 1329 1238
rect 1336 1226 1355 1238
rect 1409 1236 1436 1238
rect 1445 1236 1666 1246
rect 1701 1243 1707 1246
rect 1409 1232 1666 1236
rect 1304 1218 1355 1226
rect 1402 1218 1666 1232
rect 1710 1238 1745 1246
rect 1256 1170 1275 1204
rect 1320 1210 1349 1218
rect 1320 1204 1337 1210
rect 1320 1202 1354 1204
rect 1402 1202 1418 1218
rect 1419 1208 1627 1218
rect 1628 1208 1644 1218
rect 1692 1214 1707 1229
rect 1710 1226 1711 1238
rect 1718 1226 1745 1238
rect 1710 1218 1745 1226
rect 1710 1217 1739 1218
rect 1430 1204 1644 1208
rect 1445 1202 1644 1204
rect 1679 1204 1692 1214
rect 1710 1204 1727 1217
rect 1679 1202 1727 1204
rect 1321 1198 1354 1202
rect 1317 1196 1354 1198
rect 1317 1195 1384 1196
rect 1317 1190 1348 1195
rect 1354 1190 1384 1195
rect 1317 1186 1384 1190
rect 1290 1183 1384 1186
rect 1290 1176 1339 1183
rect 1290 1170 1320 1176
rect 1339 1171 1344 1176
rect 1256 1154 1336 1170
rect 1348 1162 1384 1183
rect 1445 1178 1634 1202
rect 1679 1201 1726 1202
rect 1692 1196 1726 1201
rect 1766 1196 1782 1198
rect 1460 1175 1634 1178
rect 1453 1172 1634 1175
rect 1662 1195 1726 1196
rect 1256 1152 1275 1154
rect 1290 1152 1324 1154
rect 1256 1136 1336 1152
rect 1256 1130 1275 1136
rect 972 1104 1075 1114
rect 926 1102 1075 1104
rect 1096 1102 1131 1114
rect 765 1100 927 1102
rect 777 1080 796 1100
rect 811 1098 841 1100
rect 660 1072 701 1080
rect 783 1076 796 1080
rect 848 1084 927 1100
rect 959 1100 1131 1102
rect 959 1084 1038 1100
rect 1045 1098 1075 1100
rect 623 1062 652 1072
rect 666 1062 695 1072
rect 710 1062 740 1076
rect 783 1062 826 1076
rect 848 1072 1038 1084
rect 1103 1080 1109 1100
rect 833 1062 863 1072
rect 864 1062 1022 1072
rect 1026 1062 1056 1072
rect 1060 1062 1090 1076
rect 1118 1062 1131 1100
rect 1203 1114 1232 1130
rect 1246 1114 1275 1130
rect 1290 1120 1320 1136
rect 1348 1114 1354 1162
rect 1357 1156 1376 1162
rect 1391 1156 1421 1164
rect 1357 1148 1421 1156
rect 1357 1132 1437 1148
rect 1453 1141 1515 1172
rect 1531 1141 1593 1172
rect 1662 1170 1711 1195
rect 1756 1186 1782 1196
rect 1726 1170 1782 1186
rect 1625 1156 1655 1164
rect 1662 1162 1772 1170
rect 1625 1148 1670 1156
rect 1357 1130 1376 1132
rect 1391 1130 1437 1132
rect 1357 1114 1437 1130
rect 1464 1128 1499 1141
rect 1540 1138 1577 1141
rect 1540 1136 1582 1138
rect 1469 1125 1499 1128
rect 1478 1121 1485 1125
rect 1485 1120 1486 1121
rect 1444 1114 1454 1120
rect 1203 1106 1238 1114
rect 1203 1080 1204 1106
rect 1211 1080 1238 1106
rect 1146 1062 1176 1076
rect 1203 1072 1238 1080
rect 1240 1106 1281 1114
rect 1240 1080 1255 1106
rect 1262 1080 1281 1106
rect 1345 1102 1376 1114
rect 1391 1102 1494 1114
rect 1506 1104 1532 1130
rect 1547 1125 1577 1136
rect 1609 1132 1671 1148
rect 1609 1130 1655 1132
rect 1609 1114 1671 1130
rect 1683 1114 1689 1162
rect 1692 1154 1772 1162
rect 1692 1152 1711 1154
rect 1726 1152 1760 1154
rect 1692 1136 1772 1152
rect 1692 1114 1711 1136
rect 1726 1120 1756 1136
rect 1784 1130 1790 1204
rect 1793 1130 1812 1274
rect 1827 1130 1833 1274
rect 1842 1204 1855 1274
rect 1907 1270 1929 1274
rect 1900 1248 1929 1262
rect 1982 1248 1998 1262
rect 2036 1258 2042 1260
rect 2049 1258 2157 1274
rect 2164 1258 2170 1260
rect 2178 1258 2193 1274
rect 2259 1268 2278 1271
rect 1900 1246 1998 1248
rect 2025 1246 2193 1258
rect 2208 1248 2224 1262
rect 2259 1249 2281 1268
rect 2291 1255 2307 1263
rect 2281 1248 2287 1249
rect 2290 1248 2319 1255
rect 2208 1247 2319 1248
rect 2208 1246 2325 1247
rect 1884 1238 1935 1246
rect 1982 1238 2016 1246
rect 1884 1226 1909 1238
rect 1916 1226 1935 1238
rect 1989 1236 2016 1238
rect 2025 1236 2246 1246
rect 2281 1243 2287 1246
rect 1989 1232 2246 1236
rect 1884 1218 1935 1226
rect 1982 1218 2246 1232
rect 2290 1238 2325 1246
rect 1836 1170 1855 1204
rect 1900 1210 1929 1218
rect 1900 1204 1917 1210
rect 1900 1202 1934 1204
rect 1982 1202 1998 1218
rect 1999 1208 2207 1218
rect 2208 1208 2224 1218
rect 2272 1214 2287 1229
rect 2290 1226 2291 1238
rect 2298 1226 2325 1238
rect 2290 1218 2325 1226
rect 2290 1217 2319 1218
rect 2010 1204 2224 1208
rect 2025 1202 2224 1204
rect 2259 1204 2272 1214
rect 2290 1204 2307 1217
rect 2259 1202 2307 1204
rect 1901 1198 1934 1202
rect 1897 1196 1934 1198
rect 1897 1195 1964 1196
rect 1897 1190 1928 1195
rect 1934 1190 1964 1195
rect 1897 1186 1964 1190
rect 1870 1183 1964 1186
rect 1870 1176 1919 1183
rect 1870 1170 1900 1176
rect 1919 1171 1924 1176
rect 1836 1154 1916 1170
rect 1928 1162 1964 1183
rect 2025 1178 2214 1202
rect 2259 1201 2306 1202
rect 2272 1196 2306 1201
rect 2040 1175 2214 1178
rect 2033 1172 2214 1175
rect 2242 1195 2306 1196
rect 1836 1152 1855 1154
rect 1870 1152 1904 1154
rect 1836 1136 1916 1152
rect 1836 1130 1855 1136
rect 1552 1104 1655 1114
rect 1506 1102 1655 1104
rect 1676 1102 1711 1114
rect 1345 1100 1507 1102
rect 1357 1080 1376 1100
rect 1391 1098 1421 1100
rect 1240 1072 1281 1080
rect 1363 1076 1376 1080
rect 1428 1084 1507 1100
rect 1539 1100 1711 1102
rect 1539 1084 1618 1100
rect 1625 1098 1655 1100
rect 1203 1062 1232 1072
rect 1246 1062 1275 1072
rect 1290 1062 1320 1076
rect 1363 1062 1406 1076
rect 1428 1072 1618 1084
rect 1683 1080 1689 1100
rect 1413 1062 1443 1072
rect 1444 1062 1602 1072
rect 1606 1062 1636 1072
rect 1640 1062 1670 1076
rect 1698 1062 1711 1100
rect 1783 1114 1812 1130
rect 1826 1114 1855 1130
rect 1870 1120 1900 1136
rect 1928 1114 1934 1162
rect 1937 1156 1956 1162
rect 1971 1156 2001 1164
rect 1937 1148 2001 1156
rect 1937 1132 2017 1148
rect 2033 1141 2095 1172
rect 2111 1141 2173 1172
rect 2242 1170 2291 1195
rect 2306 1170 2336 1188
rect 2205 1156 2235 1164
rect 2242 1162 2352 1170
rect 2205 1148 2250 1156
rect 1937 1130 1956 1132
rect 1971 1130 2017 1132
rect 1937 1114 2017 1130
rect 2044 1128 2079 1141
rect 2120 1138 2157 1141
rect 2120 1136 2162 1138
rect 2049 1125 2079 1128
rect 2058 1121 2065 1125
rect 2065 1120 2066 1121
rect 2024 1114 2034 1120
rect 1783 1106 1818 1114
rect 1783 1080 1784 1106
rect 1791 1080 1818 1106
rect 1726 1062 1756 1076
rect 1783 1072 1818 1080
rect 1820 1106 1861 1114
rect 1820 1080 1835 1106
rect 1842 1080 1861 1106
rect 1925 1102 1956 1114
rect 1971 1102 2074 1114
rect 2086 1104 2112 1130
rect 2127 1125 2157 1136
rect 2189 1132 2251 1148
rect 2189 1130 2235 1132
rect 2189 1114 2251 1130
rect 2263 1114 2269 1162
rect 2272 1154 2352 1162
rect 2272 1152 2291 1154
rect 2306 1152 2340 1154
rect 2272 1137 2352 1152
rect 2272 1136 2358 1137
rect 2272 1114 2291 1136
rect 2306 1120 2336 1136
rect 2364 1130 2370 1204
rect 2373 1130 2392 1274
rect 2407 1130 2413 1274
rect 2422 1204 2435 1274
rect 2464 1218 2479 1246
rect 2416 1170 2435 1204
rect 2477 1186 2479 1198
rect 2450 1170 2479 1186
rect 2416 1154 2479 1170
rect 2416 1152 2435 1154
rect 2450 1152 2479 1154
rect 2416 1136 2479 1152
rect 2416 1130 2435 1136
rect 2132 1104 2235 1114
rect 2086 1102 2235 1104
rect 2256 1102 2291 1114
rect 1925 1100 2087 1102
rect 1937 1080 1956 1100
rect 1971 1098 2001 1100
rect 1820 1072 1861 1080
rect 1943 1076 1956 1080
rect 2008 1084 2087 1100
rect 2119 1100 2291 1102
rect 2119 1084 2198 1100
rect 2205 1098 2235 1100
rect 1783 1062 1812 1072
rect 1826 1062 1855 1072
rect 1870 1062 1900 1076
rect 1943 1062 1986 1076
rect 2008 1072 2198 1084
rect 2263 1080 2269 1100
rect 1993 1062 2023 1072
rect 2024 1062 2182 1072
rect 2186 1062 2216 1072
rect 2220 1062 2250 1076
rect 2278 1062 2291 1100
rect 2363 1114 2392 1130
rect 2406 1114 2435 1130
rect 2450 1120 2479 1136
rect 2363 1106 2398 1114
rect 2363 1080 2364 1106
rect 2371 1080 2398 1106
rect 2306 1062 2336 1076
rect 2363 1072 2398 1080
rect 2400 1106 2441 1114
rect 2400 1080 2415 1106
rect 2422 1080 2441 1106
rect 2400 1072 2441 1080
rect 2363 1062 2392 1072
rect 2406 1062 2435 1072
rect 2450 1062 2479 1076
rect -541 1048 2479 1062
rect -478 1018 -465 1048
rect -450 1034 -420 1048
rect -377 1034 -334 1048
rect -327 1034 -107 1048
rect -100 1034 -70 1048
rect -410 1020 -395 1032
rect -376 1020 -363 1034
rect -295 1030 -142 1034
rect -413 1018 -391 1020
rect -313 1018 -121 1030
rect -42 1018 -29 1048
rect -14 1034 16 1048
rect 53 1018 72 1048
rect 87 1018 93 1048
rect 102 1018 115 1048
rect 130 1034 160 1048
rect 203 1034 246 1048
rect 253 1034 473 1048
rect 480 1034 510 1048
rect 170 1020 185 1032
rect 204 1020 217 1034
rect 285 1030 438 1034
rect 167 1018 189 1020
rect 267 1018 459 1030
rect 538 1018 551 1048
rect 566 1034 596 1048
rect 633 1018 652 1048
rect 667 1018 673 1048
rect 682 1018 695 1048
rect 710 1034 740 1048
rect 783 1034 826 1048
rect 833 1034 1053 1048
rect 1060 1034 1090 1048
rect 750 1020 765 1032
rect 784 1020 797 1034
rect 865 1030 1018 1034
rect 747 1018 769 1020
rect 847 1018 1039 1030
rect 1118 1018 1131 1048
rect 1146 1034 1176 1048
rect 1213 1018 1232 1048
rect 1247 1018 1253 1048
rect 1262 1018 1275 1048
rect 1290 1034 1320 1048
rect 1363 1034 1406 1048
rect 1413 1034 1633 1048
rect 1640 1034 1670 1048
rect 1330 1020 1345 1032
rect 1364 1020 1377 1034
rect 1445 1030 1598 1034
rect 1327 1018 1349 1020
rect 1427 1018 1619 1030
rect 1698 1018 1711 1048
rect 1726 1034 1756 1048
rect 1793 1018 1812 1048
rect 1827 1018 1833 1048
rect 1842 1018 1855 1048
rect 1870 1034 1900 1048
rect 1943 1034 1986 1048
rect 1993 1034 2213 1048
rect 2220 1034 2250 1048
rect 1910 1020 1925 1032
rect 1944 1020 1957 1034
rect 2025 1030 2178 1034
rect 1907 1018 1929 1020
rect 2007 1018 2199 1030
rect 2278 1018 2291 1048
rect 2306 1034 2336 1048
rect 2373 1018 2392 1048
rect 2407 1018 2413 1048
rect 2422 1018 2435 1048
rect 2450 1034 2479 1048
rect -541 1004 2479 1018
rect -478 934 -465 1004
rect -413 1000 -391 1004
rect -420 978 -391 992
rect -338 978 -322 992
rect -284 988 -278 990
rect -271 988 -163 1004
rect -156 988 -150 990
rect -142 988 -127 1004
rect -61 998 -42 1001
rect -420 976 -322 978
rect -295 976 -127 988
rect -112 978 -96 992
rect -61 979 -39 998
rect -29 985 -13 993
rect -39 978 -33 979
rect -30 978 -1 985
rect -112 977 -1 978
rect -112 976 5 977
rect -436 968 -385 976
rect -338 968 -304 976
rect -436 956 -411 968
rect -404 956 -385 968
rect -331 966 -304 968
rect -295 966 -74 976
rect -39 973 -33 976
rect -331 962 -74 966
rect -436 948 -385 956
rect -338 948 -74 962
rect -30 968 5 976
rect -484 900 -465 934
rect -420 940 -391 948
rect -420 934 -403 940
rect -420 932 -386 934
rect -338 932 -322 948
rect -321 938 -113 948
rect -112 938 -96 948
rect -48 944 -33 959
rect -30 956 -29 968
rect -22 956 5 968
rect -30 948 5 956
rect -30 947 -1 948
rect -310 934 -96 938
rect -295 932 -96 934
rect -61 934 -48 944
rect -30 934 -13 947
rect -61 932 -13 934
rect -419 928 -386 932
rect -423 926 -386 928
rect -423 925 -356 926
rect -423 920 -392 925
rect -386 920 -356 925
rect -423 916 -356 920
rect -450 913 -356 916
rect -450 906 -401 913
rect -450 900 -420 906
rect -401 901 -396 906
rect -484 884 -404 900
rect -392 892 -356 913
rect -295 908 -106 932
rect -61 931 -14 932
rect -48 926 -14 931
rect -280 905 -106 908
rect -287 902 -106 905
rect -78 925 -14 926
rect -484 882 -465 884
rect -450 882 -416 884
rect -484 866 -404 882
rect -484 860 -465 866
rect -494 844 -465 860
rect -450 850 -420 866
rect -392 844 -386 892
rect -383 886 -364 892
rect -349 886 -319 894
rect -383 878 -319 886
rect -383 862 -303 878
rect -287 871 -225 902
rect -209 871 -147 902
rect -78 900 -29 925
rect -14 900 16 918
rect -115 886 -85 894
rect -78 892 32 900
rect -115 878 -70 886
rect -383 860 -364 862
rect -349 860 -303 862
rect -383 844 -303 860
rect -276 858 -241 871
rect -200 868 -163 871
rect -200 866 -158 868
rect -271 855 -241 858
rect -262 851 -255 855
rect -255 850 -254 851
rect -296 844 -286 850
rect -500 836 -459 844
rect -500 810 -485 836
rect -478 810 -459 836
rect -395 832 -364 844
rect -349 832 -246 844
rect -234 834 -208 860
rect -193 855 -163 866
rect -131 862 -69 878
rect -131 860 -85 862
rect -131 844 -69 860
rect -57 844 -51 892
rect -48 884 32 892
rect -48 882 -29 884
rect -14 882 20 884
rect -48 867 32 882
rect -48 866 38 867
rect -48 844 -29 866
rect -14 850 16 866
rect 44 860 50 934
rect 53 860 72 1004
rect 87 860 93 1004
rect 102 934 115 1004
rect 167 1000 189 1004
rect 160 978 189 992
rect 242 978 258 992
rect 296 988 302 990
rect 309 988 417 1004
rect 424 988 430 990
rect 438 988 453 1004
rect 519 998 538 1001
rect 160 976 258 978
rect 285 976 453 988
rect 468 978 484 992
rect 519 979 541 998
rect 551 985 567 993
rect 541 978 547 979
rect 550 978 579 985
rect 468 977 579 978
rect 468 976 585 977
rect 144 968 195 976
rect 242 968 276 976
rect 144 956 169 968
rect 176 956 195 968
rect 249 966 276 968
rect 285 966 506 976
rect 541 973 547 976
rect 249 962 506 966
rect 144 948 195 956
rect 242 948 506 962
rect 550 968 585 976
rect 96 900 115 934
rect 160 940 189 948
rect 160 934 177 940
rect 160 932 194 934
rect 242 932 258 948
rect 259 938 467 948
rect 468 938 484 948
rect 532 944 547 959
rect 550 956 551 968
rect 558 956 585 968
rect 550 948 585 956
rect 550 947 579 948
rect 270 934 484 938
rect 285 932 484 934
rect 519 934 532 944
rect 550 934 567 947
rect 519 932 567 934
rect 161 928 194 932
rect 157 926 194 928
rect 157 925 224 926
rect 157 920 188 925
rect 194 920 224 925
rect 157 916 224 920
rect 130 913 224 916
rect 130 906 179 913
rect 130 900 160 906
rect 179 901 184 906
rect 96 884 176 900
rect 188 892 224 913
rect 285 908 474 932
rect 519 931 566 932
rect 532 926 566 931
rect 606 926 622 928
rect 300 905 474 908
rect 293 902 474 905
rect 502 925 566 926
rect 96 882 115 884
rect 130 882 164 884
rect 96 866 176 882
rect 96 860 115 866
rect -188 834 -85 844
rect -234 832 -85 834
rect -64 832 -29 844
rect -395 830 -233 832
rect -383 812 -364 830
rect -349 828 -319 830
rect -500 802 -459 810
rect -376 806 -364 812
rect -312 814 -233 830
rect -201 830 -29 832
rect -201 814 -122 830
rect -115 828 -85 830
rect -494 792 -465 802
rect -450 792 -420 806
rect -376 792 -334 806
rect -312 802 -122 814
rect -57 810 -51 830
rect -327 792 -297 802
rect -296 792 -138 802
rect -134 792 -104 802
rect -100 792 -70 806
rect -42 792 -29 830
rect 43 844 72 860
rect 86 844 115 860
rect 130 850 160 866
rect 188 844 194 892
rect 197 886 216 892
rect 231 886 261 894
rect 197 878 261 886
rect 197 862 277 878
rect 293 871 355 902
rect 371 871 433 902
rect 502 900 551 925
rect 596 916 622 926
rect 566 900 622 916
rect 465 886 495 894
rect 502 892 612 900
rect 465 878 510 886
rect 197 860 216 862
rect 231 860 277 862
rect 197 844 277 860
rect 304 858 339 871
rect 380 868 417 871
rect 380 866 422 868
rect 309 855 339 858
rect 318 851 325 855
rect 325 850 326 851
rect 284 844 294 850
rect 43 836 78 844
rect 43 810 44 836
rect 51 810 78 836
rect -14 792 16 806
rect 43 802 78 810
rect 80 836 121 844
rect 80 810 95 836
rect 102 810 121 836
rect 185 832 216 844
rect 231 832 334 844
rect 346 834 372 860
rect 387 855 417 866
rect 449 862 511 878
rect 449 860 495 862
rect 449 844 511 860
rect 523 844 529 892
rect 532 884 612 892
rect 532 882 551 884
rect 566 882 600 884
rect 532 866 612 882
rect 532 844 551 866
rect 566 850 596 866
rect 624 860 630 934
rect 633 860 652 1004
rect 667 860 673 1004
rect 682 934 695 1004
rect 747 1000 769 1004
rect 740 978 769 992
rect 822 978 838 992
rect 876 988 882 990
rect 889 988 997 1004
rect 1004 988 1010 990
rect 1018 988 1033 1004
rect 1099 998 1118 1001
rect 740 976 838 978
rect 865 976 1033 988
rect 1048 978 1064 992
rect 1099 979 1121 998
rect 1131 985 1147 993
rect 1121 978 1127 979
rect 1130 978 1159 985
rect 1048 977 1159 978
rect 1048 976 1165 977
rect 724 968 775 976
rect 822 968 856 976
rect 724 956 749 968
rect 756 956 775 968
rect 829 966 856 968
rect 865 966 1086 976
rect 1121 973 1127 976
rect 829 962 1086 966
rect 724 948 775 956
rect 822 948 1086 962
rect 1130 968 1165 976
rect 676 900 695 934
rect 740 940 769 948
rect 740 934 757 940
rect 740 932 774 934
rect 822 932 838 948
rect 839 938 1047 948
rect 1048 938 1064 948
rect 1112 944 1127 959
rect 1130 956 1131 968
rect 1138 956 1165 968
rect 1130 948 1165 956
rect 1130 947 1159 948
rect 850 934 1064 938
rect 865 932 1064 934
rect 1099 934 1112 944
rect 1130 934 1147 947
rect 1099 932 1147 934
rect 741 928 774 932
rect 737 926 774 928
rect 737 925 804 926
rect 737 920 768 925
rect 774 920 804 925
rect 737 916 804 920
rect 710 913 804 916
rect 710 906 759 913
rect 710 900 740 906
rect 759 901 764 906
rect 676 884 756 900
rect 768 892 804 913
rect 865 908 1054 932
rect 1099 931 1146 932
rect 1112 926 1146 931
rect 880 905 1054 908
rect 873 902 1054 905
rect 1082 925 1146 926
rect 676 882 695 884
rect 710 882 744 884
rect 676 866 756 882
rect 676 860 695 866
rect 392 834 495 844
rect 346 832 495 834
rect 516 832 551 844
rect 185 830 347 832
rect 197 812 216 830
rect 231 828 261 830
rect 80 802 121 810
rect 204 806 216 812
rect 268 814 347 830
rect 379 830 551 832
rect 379 814 458 830
rect 465 828 495 830
rect 43 792 72 802
rect 86 792 115 802
rect 130 792 160 806
rect 204 792 246 806
rect 268 802 458 814
rect 523 810 529 830
rect 253 792 283 802
rect 284 792 442 802
rect 446 792 476 802
rect 480 792 510 806
rect 538 792 551 830
rect 623 844 652 860
rect 666 844 695 860
rect 710 850 740 866
rect 768 844 774 892
rect 777 886 796 892
rect 811 886 841 894
rect 777 878 841 886
rect 777 862 857 878
rect 873 871 935 902
rect 951 871 1013 902
rect 1082 900 1131 925
rect 1146 900 1176 918
rect 1045 886 1075 894
rect 1082 892 1192 900
rect 1045 878 1090 886
rect 777 860 796 862
rect 811 860 857 862
rect 777 844 857 860
rect 884 858 919 871
rect 960 868 997 871
rect 960 866 1002 868
rect 889 855 919 858
rect 898 851 905 855
rect 905 850 906 851
rect 864 844 874 850
rect 623 836 658 844
rect 623 810 624 836
rect 631 810 658 836
rect 566 792 596 806
rect 623 802 658 810
rect 660 836 701 844
rect 660 810 675 836
rect 682 810 701 836
rect 765 832 796 844
rect 811 832 914 844
rect 926 834 952 860
rect 967 855 997 866
rect 1029 862 1091 878
rect 1029 860 1075 862
rect 1029 844 1091 860
rect 1103 844 1109 892
rect 1112 884 1192 892
rect 1112 882 1131 884
rect 1146 882 1180 884
rect 1112 867 1192 882
rect 1112 866 1198 867
rect 1112 844 1131 866
rect 1146 850 1176 866
rect 1204 860 1210 934
rect 1213 860 1232 1004
rect 1247 860 1253 1004
rect 1262 934 1275 1004
rect 1327 1000 1349 1004
rect 1320 978 1349 992
rect 1402 978 1418 992
rect 1456 988 1462 990
rect 1469 988 1577 1004
rect 1584 988 1590 990
rect 1598 988 1613 1004
rect 1679 998 1698 1001
rect 1320 976 1418 978
rect 1445 976 1613 988
rect 1628 978 1644 992
rect 1679 979 1701 998
rect 1711 985 1727 993
rect 1701 978 1707 979
rect 1710 978 1739 985
rect 1628 977 1739 978
rect 1628 976 1745 977
rect 1304 968 1355 976
rect 1402 968 1436 976
rect 1304 956 1329 968
rect 1336 956 1355 968
rect 1409 966 1436 968
rect 1445 966 1666 976
rect 1701 973 1707 976
rect 1409 962 1666 966
rect 1304 948 1355 956
rect 1402 948 1666 962
rect 1710 968 1745 976
rect 1256 900 1275 934
rect 1320 940 1349 948
rect 1320 934 1337 940
rect 1320 932 1354 934
rect 1402 932 1418 948
rect 1419 938 1627 948
rect 1628 938 1644 948
rect 1692 944 1707 959
rect 1710 956 1711 968
rect 1718 956 1745 968
rect 1710 948 1745 956
rect 1710 947 1739 948
rect 1430 934 1644 938
rect 1445 932 1644 934
rect 1679 934 1692 944
rect 1710 934 1727 947
rect 1679 932 1727 934
rect 1321 928 1354 932
rect 1317 926 1354 928
rect 1317 925 1384 926
rect 1317 920 1348 925
rect 1354 920 1384 925
rect 1317 916 1384 920
rect 1290 913 1384 916
rect 1290 906 1339 913
rect 1290 900 1320 906
rect 1339 901 1344 906
rect 1256 884 1336 900
rect 1348 892 1384 913
rect 1445 908 1634 932
rect 1679 931 1726 932
rect 1692 926 1726 931
rect 1766 926 1782 928
rect 1460 905 1634 908
rect 1453 902 1634 905
rect 1662 925 1726 926
rect 1256 882 1275 884
rect 1290 882 1324 884
rect 1256 866 1336 882
rect 1256 860 1275 866
rect 972 834 1075 844
rect 926 832 1075 834
rect 1096 832 1131 844
rect 765 830 927 832
rect 777 812 796 830
rect 811 828 841 830
rect 660 802 701 810
rect 784 806 796 812
rect 848 814 927 830
rect 959 830 1131 832
rect 959 814 1038 830
rect 1045 828 1075 830
rect 623 792 652 802
rect 666 792 695 802
rect 710 792 740 806
rect 784 792 826 806
rect 848 802 1038 814
rect 1103 810 1109 830
rect 833 792 863 802
rect 864 792 1022 802
rect 1026 792 1056 802
rect 1060 792 1090 806
rect 1118 792 1131 830
rect 1203 844 1232 860
rect 1246 844 1275 860
rect 1290 850 1320 866
rect 1348 844 1354 892
rect 1357 886 1376 892
rect 1391 886 1421 894
rect 1357 878 1421 886
rect 1357 862 1437 878
rect 1453 871 1515 902
rect 1531 871 1593 902
rect 1662 900 1711 925
rect 1756 916 1782 926
rect 1726 900 1782 916
rect 1625 886 1655 894
rect 1662 892 1772 900
rect 1625 878 1670 886
rect 1357 860 1376 862
rect 1391 860 1437 862
rect 1357 844 1437 860
rect 1464 858 1499 871
rect 1540 868 1577 871
rect 1540 866 1582 868
rect 1469 855 1499 858
rect 1478 851 1485 855
rect 1485 850 1486 851
rect 1444 844 1454 850
rect 1203 836 1238 844
rect 1203 810 1204 836
rect 1211 810 1238 836
rect 1146 792 1176 806
rect 1203 802 1238 810
rect 1240 836 1281 844
rect 1240 810 1255 836
rect 1262 810 1281 836
rect 1345 832 1376 844
rect 1391 832 1494 844
rect 1506 834 1532 860
rect 1547 855 1577 866
rect 1609 862 1671 878
rect 1609 860 1655 862
rect 1609 844 1671 860
rect 1683 844 1689 892
rect 1692 884 1772 892
rect 1692 882 1711 884
rect 1726 882 1760 884
rect 1692 866 1772 882
rect 1692 844 1711 866
rect 1726 850 1756 866
rect 1784 860 1790 934
rect 1793 860 1812 1004
rect 1827 860 1833 1004
rect 1842 934 1855 1004
rect 1907 1000 1929 1004
rect 1900 978 1929 992
rect 1982 978 1998 992
rect 2036 988 2042 990
rect 2049 988 2157 1004
rect 2164 988 2170 990
rect 2178 988 2193 1004
rect 2259 998 2278 1001
rect 1900 976 1998 978
rect 2025 976 2193 988
rect 2208 978 2224 992
rect 2259 979 2281 998
rect 2291 985 2307 993
rect 2281 978 2287 979
rect 2290 978 2319 985
rect 2208 977 2319 978
rect 2208 976 2325 977
rect 1884 968 1935 976
rect 1982 968 2016 976
rect 1884 956 1909 968
rect 1916 956 1935 968
rect 1989 966 2016 968
rect 2025 966 2246 976
rect 2281 973 2287 976
rect 1989 962 2246 966
rect 1884 948 1935 956
rect 1982 948 2246 962
rect 2290 968 2325 976
rect 1836 900 1855 934
rect 1900 940 1929 948
rect 1900 934 1917 940
rect 1900 932 1934 934
rect 1982 932 1998 948
rect 1999 938 2207 948
rect 2208 938 2224 948
rect 2272 944 2287 959
rect 2290 956 2291 968
rect 2298 956 2325 968
rect 2290 948 2325 956
rect 2290 947 2319 948
rect 2010 934 2224 938
rect 2025 932 2224 934
rect 2259 934 2272 944
rect 2290 934 2307 947
rect 2259 932 2307 934
rect 1901 928 1934 932
rect 1897 926 1934 928
rect 1897 925 1964 926
rect 1897 920 1928 925
rect 1934 920 1964 925
rect 1897 916 1964 920
rect 1870 913 1964 916
rect 1870 906 1919 913
rect 1870 900 1900 906
rect 1919 901 1924 906
rect 1836 884 1916 900
rect 1928 892 1964 913
rect 2025 908 2214 932
rect 2259 931 2306 932
rect 2272 926 2306 931
rect 2040 905 2214 908
rect 2033 902 2214 905
rect 2242 925 2306 926
rect 1836 882 1855 884
rect 1870 882 1904 884
rect 1836 866 1916 882
rect 1836 860 1855 866
rect 1552 834 1655 844
rect 1506 832 1655 834
rect 1676 832 1711 844
rect 1345 830 1507 832
rect 1357 812 1376 830
rect 1391 828 1421 830
rect 1240 802 1281 810
rect 1364 806 1376 812
rect 1428 814 1507 830
rect 1539 830 1711 832
rect 1539 814 1618 830
rect 1625 828 1655 830
rect 1203 792 1232 802
rect 1246 792 1275 802
rect 1290 792 1320 806
rect 1364 792 1406 806
rect 1428 802 1618 814
rect 1683 810 1689 830
rect 1413 792 1443 802
rect 1444 792 1602 802
rect 1606 792 1636 802
rect 1640 792 1670 806
rect 1698 792 1711 830
rect 1783 844 1812 860
rect 1826 844 1855 860
rect 1870 850 1900 866
rect 1928 844 1934 892
rect 1937 886 1956 892
rect 1971 886 2001 894
rect 1937 878 2001 886
rect 1937 862 2017 878
rect 2033 871 2095 902
rect 2111 871 2173 902
rect 2242 900 2291 925
rect 2306 900 2336 918
rect 2205 886 2235 894
rect 2242 892 2352 900
rect 2205 878 2250 886
rect 1937 860 1956 862
rect 1971 860 2017 862
rect 1937 844 2017 860
rect 2044 858 2079 871
rect 2120 868 2157 871
rect 2120 866 2162 868
rect 2049 855 2079 858
rect 2058 851 2065 855
rect 2065 850 2066 851
rect 2024 844 2034 850
rect 1783 836 1818 844
rect 1783 810 1784 836
rect 1791 810 1818 836
rect 1726 792 1756 806
rect 1783 802 1818 810
rect 1820 836 1861 844
rect 1820 810 1835 836
rect 1842 810 1861 836
rect 1925 832 1956 844
rect 1971 832 2074 844
rect 2086 834 2112 860
rect 2127 855 2157 866
rect 2189 862 2251 878
rect 2189 860 2235 862
rect 2189 844 2251 860
rect 2263 844 2269 892
rect 2272 884 2352 892
rect 2272 882 2291 884
rect 2306 882 2340 884
rect 2272 867 2352 882
rect 2272 866 2358 867
rect 2272 844 2291 866
rect 2306 850 2336 866
rect 2364 860 2370 934
rect 2373 860 2392 1004
rect 2407 860 2413 1004
rect 2422 934 2435 1004
rect 2464 948 2479 976
rect 2416 900 2435 934
rect 2477 916 2479 928
rect 2450 900 2479 916
rect 2416 884 2479 900
rect 2416 882 2435 884
rect 2450 882 2479 884
rect 2416 866 2479 882
rect 2416 860 2435 866
rect 2132 834 2235 844
rect 2086 832 2235 834
rect 2256 832 2291 844
rect 1925 830 2087 832
rect 1937 812 1956 830
rect 1971 828 2001 830
rect 1820 802 1861 810
rect 1944 806 1956 812
rect 2008 814 2087 830
rect 2119 830 2291 832
rect 2119 814 2198 830
rect 2205 828 2235 830
rect 1783 792 1812 802
rect 1826 792 1855 802
rect 1870 792 1900 806
rect 1944 792 1986 806
rect 2008 802 2198 814
rect 2263 810 2269 830
rect 1993 792 2023 802
rect 2024 792 2182 802
rect 2186 792 2216 802
rect 2220 792 2250 806
rect 2278 792 2291 830
rect 2363 844 2392 860
rect 2406 844 2435 860
rect 2450 850 2479 866
rect 2363 836 2398 844
rect 2363 810 2364 836
rect 2371 810 2398 836
rect 2306 792 2336 806
rect 2363 802 2398 810
rect 2400 836 2441 844
rect 2400 810 2415 836
rect 2422 810 2441 836
rect 2400 802 2441 810
rect 2363 792 2392 802
rect 2406 792 2435 802
rect 2450 792 2479 806
rect -541 778 2479 792
rect -478 748 -465 778
rect -450 764 -420 778
rect -376 764 -334 778
rect -327 764 -107 778
rect -100 764 -70 778
rect -410 750 -395 762
rect -376 750 -363 764
rect -295 760 -142 764
rect -413 748 -391 750
rect -313 748 -121 760
rect -42 748 -29 778
rect -14 764 16 778
rect 53 748 72 778
rect 87 748 93 778
rect 102 748 115 778
rect 130 764 160 778
rect 204 764 246 778
rect 253 764 473 778
rect 480 764 510 778
rect 170 750 185 762
rect 204 750 217 764
rect 285 760 438 764
rect 167 748 189 750
rect 267 748 459 760
rect 538 748 551 778
rect 566 764 596 778
rect 633 748 652 778
rect 667 748 673 778
rect 682 748 695 778
rect 710 764 740 778
rect 784 764 826 778
rect 833 764 1053 778
rect 1060 764 1090 778
rect 750 750 765 762
rect 784 750 797 764
rect 865 760 1018 764
rect 747 748 769 750
rect 847 748 1039 760
rect 1118 748 1131 778
rect 1146 764 1176 778
rect 1213 748 1232 778
rect 1247 748 1253 778
rect 1262 748 1275 778
rect 1290 764 1320 778
rect 1364 764 1406 778
rect 1413 764 1633 778
rect 1640 764 1670 778
rect 1330 750 1345 762
rect 1364 750 1377 764
rect 1445 760 1598 764
rect 1327 748 1349 750
rect 1427 748 1619 760
rect 1698 748 1711 778
rect 1726 764 1756 778
rect 1793 748 1812 778
rect 1827 748 1833 778
rect 1842 748 1855 778
rect 1870 764 1900 778
rect 1944 764 1986 778
rect 1993 764 2213 778
rect 2220 764 2250 778
rect 1910 750 1925 762
rect 1944 750 1957 764
rect 2025 760 2178 764
rect 1907 748 1929 750
rect 2007 748 2199 760
rect 2278 748 2291 778
rect 2306 764 2336 778
rect 2373 748 2392 778
rect 2407 748 2413 778
rect 2422 748 2435 778
rect 2450 764 2479 778
rect -541 734 2479 748
rect -478 664 -465 734
rect -413 730 -391 734
rect -420 708 -391 722
rect -338 708 -322 722
rect -284 718 -278 720
rect -271 718 -163 734
rect -156 718 -150 720
rect -142 718 -127 734
rect -61 728 -42 731
rect -420 706 -322 708
rect -295 706 -127 718
rect -112 708 -96 722
rect -61 709 -39 728
rect -29 715 -13 723
rect -39 708 -33 709
rect -30 708 -1 715
rect -112 707 -1 708
rect -112 706 5 707
rect -436 698 -385 706
rect -338 698 -304 706
rect -436 686 -411 698
rect -404 686 -385 698
rect -331 696 -304 698
rect -295 696 -74 706
rect -39 703 -33 706
rect -331 692 -74 696
rect -436 678 -385 686
rect -338 678 -74 692
rect -30 698 5 706
rect -484 630 -465 664
rect -420 670 -391 678
rect -420 664 -403 670
rect -420 662 -386 664
rect -338 662 -322 678
rect -321 668 -113 678
rect -112 668 -96 678
rect -48 674 -33 689
rect -30 686 -29 698
rect -22 686 5 698
rect -30 678 5 686
rect -30 677 -1 678
rect -310 664 -96 668
rect -295 662 -96 664
rect -61 664 -48 674
rect -30 664 -13 677
rect -61 662 -13 664
rect -419 658 -386 662
rect -423 656 -386 658
rect -423 655 -356 656
rect -423 650 -392 655
rect -386 650 -356 655
rect -423 646 -356 650
rect -450 643 -356 646
rect -450 636 -401 643
rect -450 630 -420 636
rect -401 631 -396 636
rect -484 614 -404 630
rect -392 622 -356 643
rect -295 638 -106 662
rect -61 661 -14 662
rect -48 656 -14 661
rect -280 635 -106 638
rect -287 632 -106 635
rect -78 655 -14 656
rect -484 612 -465 614
rect -450 612 -416 614
rect -484 596 -404 612
rect -484 590 -465 596
rect -494 574 -465 590
rect -450 580 -420 596
rect -392 574 -386 622
rect -383 616 -364 622
rect -349 616 -319 624
rect -383 608 -319 616
rect -383 592 -303 608
rect -287 601 -225 632
rect -209 601 -147 632
rect -78 630 -29 655
rect -14 630 16 648
rect -115 616 -85 624
rect -78 622 32 630
rect -115 608 -70 616
rect -383 590 -364 592
rect -349 590 -303 592
rect -383 574 -303 590
rect -276 588 -241 601
rect -200 598 -163 601
rect -200 596 -158 598
rect -271 585 -241 588
rect -262 581 -255 585
rect -255 580 -254 581
rect -296 574 -286 580
rect -500 566 -459 574
rect -500 540 -485 566
rect -478 540 -459 566
rect -395 562 -364 574
rect -349 562 -246 574
rect -234 564 -208 590
rect -193 585 -163 596
rect -131 592 -69 608
rect -131 590 -85 592
rect -131 574 -69 590
rect -57 574 -51 622
rect -48 614 32 622
rect -48 612 -29 614
rect -14 612 20 614
rect -48 597 32 612
rect -48 596 38 597
rect -48 574 -29 596
rect -14 580 16 596
rect 44 590 50 664
rect 53 590 72 734
rect 87 590 93 734
rect 102 664 115 734
rect 167 730 189 734
rect 160 708 189 722
rect 242 708 258 722
rect 296 718 302 720
rect 309 718 417 734
rect 424 718 430 720
rect 438 718 453 734
rect 519 728 538 731
rect 160 706 258 708
rect 285 706 453 718
rect 468 708 484 722
rect 519 709 541 728
rect 551 715 567 723
rect 541 708 547 709
rect 550 708 579 715
rect 468 707 579 708
rect 468 706 585 707
rect 144 698 195 706
rect 242 698 276 706
rect 144 686 169 698
rect 176 686 195 698
rect 249 696 276 698
rect 285 696 506 706
rect 541 703 547 706
rect 249 692 506 696
rect 144 678 195 686
rect 242 678 506 692
rect 550 698 585 706
rect 96 630 115 664
rect 160 670 189 678
rect 160 664 177 670
rect 160 662 194 664
rect 242 662 258 678
rect 259 668 467 678
rect 468 668 484 678
rect 532 674 547 689
rect 550 686 551 698
rect 558 686 585 698
rect 550 678 585 686
rect 550 677 579 678
rect 270 664 484 668
rect 285 662 484 664
rect 519 664 532 674
rect 550 664 567 677
rect 519 662 567 664
rect 161 658 194 662
rect 157 656 194 658
rect 157 655 224 656
rect 157 650 188 655
rect 194 650 224 655
rect 157 646 224 650
rect 130 643 224 646
rect 130 636 179 643
rect 130 630 160 636
rect 179 631 184 636
rect 96 614 176 630
rect 188 622 224 643
rect 285 638 474 662
rect 519 661 566 662
rect 532 656 566 661
rect 606 656 622 658
rect 300 635 474 638
rect 293 632 474 635
rect 502 655 566 656
rect 96 612 115 614
rect 130 612 164 614
rect 96 596 176 612
rect 96 590 115 596
rect -188 564 -85 574
rect -234 562 -85 564
rect -64 562 -29 574
rect -395 560 -233 562
rect -383 540 -364 560
rect -349 558 -319 560
rect -500 532 -459 540
rect -377 536 -364 540
rect -312 544 -233 560
rect -201 560 -29 562
rect -201 544 -122 560
rect -115 558 -85 560
rect -494 522 -465 532
rect -450 522 -420 536
rect -377 522 -334 536
rect -312 532 -122 544
rect -57 540 -51 560
rect -327 522 -297 532
rect -296 522 -138 532
rect -134 522 -104 532
rect -100 522 -70 536
rect -42 522 -29 560
rect 43 574 72 590
rect 86 574 115 590
rect 130 580 160 596
rect 188 574 194 622
rect 197 616 216 622
rect 231 616 261 624
rect 197 608 261 616
rect 197 592 277 608
rect 293 601 355 632
rect 371 601 433 632
rect 502 630 551 655
rect 596 646 622 656
rect 566 630 622 646
rect 465 616 495 624
rect 502 622 612 630
rect 465 608 510 616
rect 197 590 216 592
rect 231 590 277 592
rect 197 574 277 590
rect 304 588 339 601
rect 380 598 417 601
rect 380 596 422 598
rect 309 585 339 588
rect 318 581 325 585
rect 325 580 326 581
rect 284 574 294 580
rect 43 566 78 574
rect 43 540 44 566
rect 51 540 78 566
rect -14 522 16 536
rect 43 532 78 540
rect 80 566 121 574
rect 80 540 95 566
rect 102 540 121 566
rect 185 562 216 574
rect 231 562 334 574
rect 346 564 372 590
rect 387 585 417 596
rect 449 592 511 608
rect 449 590 495 592
rect 449 574 511 590
rect 523 574 529 622
rect 532 614 612 622
rect 532 612 551 614
rect 566 612 600 614
rect 532 596 612 612
rect 532 574 551 596
rect 566 580 596 596
rect 624 590 630 664
rect 633 590 652 734
rect 667 590 673 734
rect 682 664 695 734
rect 747 730 769 734
rect 740 708 769 722
rect 822 708 838 722
rect 876 718 882 720
rect 889 718 997 734
rect 1004 718 1010 720
rect 1018 718 1033 734
rect 1099 728 1118 731
rect 740 706 838 708
rect 865 706 1033 718
rect 1048 708 1064 722
rect 1099 709 1121 728
rect 1131 715 1147 723
rect 1121 708 1127 709
rect 1130 708 1159 715
rect 1048 707 1159 708
rect 1048 706 1165 707
rect 724 698 775 706
rect 822 698 856 706
rect 724 686 749 698
rect 756 686 775 698
rect 829 696 856 698
rect 865 696 1086 706
rect 1121 703 1127 706
rect 829 692 1086 696
rect 724 678 775 686
rect 822 678 1086 692
rect 1130 698 1165 706
rect 676 630 695 664
rect 740 670 769 678
rect 740 664 757 670
rect 740 662 774 664
rect 822 662 838 678
rect 839 668 1047 678
rect 1048 668 1064 678
rect 1112 674 1127 689
rect 1130 686 1131 698
rect 1138 686 1165 698
rect 1130 678 1165 686
rect 1130 677 1159 678
rect 850 664 1064 668
rect 865 662 1064 664
rect 1099 664 1112 674
rect 1130 664 1147 677
rect 1099 662 1147 664
rect 741 658 774 662
rect 737 656 774 658
rect 737 655 804 656
rect 737 650 768 655
rect 774 650 804 655
rect 737 646 804 650
rect 710 643 804 646
rect 710 636 759 643
rect 710 630 740 636
rect 759 631 764 636
rect 676 614 756 630
rect 768 622 804 643
rect 865 638 1054 662
rect 1099 661 1146 662
rect 1112 656 1146 661
rect 880 635 1054 638
rect 873 632 1054 635
rect 1082 655 1146 656
rect 676 612 695 614
rect 710 612 744 614
rect 676 596 756 612
rect 676 590 695 596
rect 392 564 495 574
rect 346 562 495 564
rect 516 562 551 574
rect 185 560 347 562
rect 197 540 216 560
rect 231 558 261 560
rect 80 532 121 540
rect 203 536 216 540
rect 268 544 347 560
rect 379 560 551 562
rect 379 544 458 560
rect 465 558 495 560
rect 43 522 72 532
rect 86 522 115 532
rect 130 522 160 536
rect 203 522 246 536
rect 268 532 458 544
rect 523 540 529 560
rect 253 522 283 532
rect 284 522 442 532
rect 446 522 476 532
rect 480 522 510 536
rect 538 522 551 560
rect 623 574 652 590
rect 666 574 695 590
rect 710 580 740 596
rect 768 574 774 622
rect 777 616 796 622
rect 811 616 841 624
rect 777 608 841 616
rect 777 592 857 608
rect 873 601 935 632
rect 951 601 1013 632
rect 1082 630 1131 655
rect 1146 630 1176 648
rect 1045 616 1075 624
rect 1082 622 1192 630
rect 1045 608 1090 616
rect 777 590 796 592
rect 811 590 857 592
rect 777 574 857 590
rect 884 588 919 601
rect 960 598 997 601
rect 960 596 1002 598
rect 889 585 919 588
rect 898 581 905 585
rect 905 580 906 581
rect 864 574 874 580
rect 623 566 658 574
rect 623 540 624 566
rect 631 540 658 566
rect 566 522 596 536
rect 623 532 658 540
rect 660 566 701 574
rect 660 540 675 566
rect 682 540 701 566
rect 765 562 796 574
rect 811 562 914 574
rect 926 564 952 590
rect 967 585 997 596
rect 1029 592 1091 608
rect 1029 590 1075 592
rect 1029 574 1091 590
rect 1103 574 1109 622
rect 1112 614 1192 622
rect 1112 612 1131 614
rect 1146 612 1180 614
rect 1112 597 1192 612
rect 1112 596 1198 597
rect 1112 574 1131 596
rect 1146 580 1176 596
rect 1204 590 1210 664
rect 1213 590 1232 734
rect 1247 590 1253 734
rect 1262 664 1275 734
rect 1327 730 1349 734
rect 1320 708 1349 722
rect 1402 708 1418 722
rect 1456 718 1462 720
rect 1469 718 1577 734
rect 1584 718 1590 720
rect 1598 718 1613 734
rect 1679 728 1698 731
rect 1320 706 1418 708
rect 1445 706 1613 718
rect 1628 708 1644 722
rect 1679 709 1701 728
rect 1711 715 1727 723
rect 1701 708 1707 709
rect 1710 708 1739 715
rect 1628 707 1739 708
rect 1628 706 1745 707
rect 1304 698 1355 706
rect 1402 698 1436 706
rect 1304 686 1329 698
rect 1336 686 1355 698
rect 1409 696 1436 698
rect 1445 696 1666 706
rect 1701 703 1707 706
rect 1409 692 1666 696
rect 1304 678 1355 686
rect 1402 678 1666 692
rect 1710 698 1745 706
rect 1256 630 1275 664
rect 1320 670 1349 678
rect 1320 664 1337 670
rect 1320 662 1354 664
rect 1402 662 1418 678
rect 1419 668 1627 678
rect 1628 668 1644 678
rect 1692 674 1707 689
rect 1710 686 1711 698
rect 1718 686 1745 698
rect 1710 678 1745 686
rect 1710 677 1739 678
rect 1430 664 1644 668
rect 1445 662 1644 664
rect 1679 664 1692 674
rect 1710 664 1727 677
rect 1679 662 1727 664
rect 1321 658 1354 662
rect 1317 656 1354 658
rect 1317 655 1384 656
rect 1317 650 1348 655
rect 1354 650 1384 655
rect 1317 646 1384 650
rect 1290 643 1384 646
rect 1290 636 1339 643
rect 1290 630 1320 636
rect 1339 631 1344 636
rect 1256 614 1336 630
rect 1348 622 1384 643
rect 1445 638 1634 662
rect 1679 661 1726 662
rect 1692 656 1726 661
rect 1766 656 1782 658
rect 1460 635 1634 638
rect 1453 632 1634 635
rect 1662 655 1726 656
rect 1256 612 1275 614
rect 1290 612 1324 614
rect 1256 596 1336 612
rect 1256 590 1275 596
rect 972 564 1075 574
rect 926 562 1075 564
rect 1096 562 1131 574
rect 765 560 927 562
rect 777 540 796 560
rect 811 558 841 560
rect 660 532 701 540
rect 783 536 796 540
rect 848 544 927 560
rect 959 560 1131 562
rect 959 544 1038 560
rect 1045 558 1075 560
rect 623 522 652 532
rect 666 522 695 532
rect 710 522 740 536
rect 783 522 826 536
rect 848 532 1038 544
rect 1103 540 1109 560
rect 833 522 863 532
rect 864 522 1022 532
rect 1026 522 1056 532
rect 1060 522 1090 536
rect 1118 522 1131 560
rect 1203 574 1232 590
rect 1246 574 1275 590
rect 1290 584 1320 596
rect 1348 584 1354 622
rect 1357 616 1376 622
rect 1391 616 1421 624
rect 1357 608 1421 616
rect 1357 592 1437 608
rect 1453 601 1515 632
rect 1531 601 1593 632
rect 1662 630 1711 655
rect 1756 646 1782 656
rect 1726 630 1782 646
rect 1625 616 1655 624
rect 1662 622 1772 630
rect 1625 608 1670 616
rect 1357 590 1376 592
rect 1391 590 1437 592
rect 1357 584 1437 590
rect 1464 588 1499 601
rect 1540 598 1577 601
rect 1540 596 1582 598
rect 1469 585 1499 588
rect 1478 584 1485 585
rect 1506 584 1532 590
rect 1547 585 1577 596
rect 1609 592 1671 608
rect 1609 590 1655 592
rect 1609 584 1671 590
rect 1683 584 1689 622
rect 1692 614 1772 622
rect 1692 612 1711 614
rect 1726 612 1760 614
rect 1692 596 1772 612
rect 1692 584 1711 596
rect 1726 584 1756 596
rect 1784 590 1790 664
rect 1793 590 1812 734
rect 1784 584 1812 590
rect 1827 590 1833 734
rect 1842 664 1855 734
rect 1907 730 1929 734
rect 1900 708 1929 722
rect 1982 708 1998 722
rect 2036 718 2042 720
rect 2049 718 2157 734
rect 2164 718 2170 720
rect 2178 718 2193 734
rect 2259 728 2278 731
rect 1900 706 1998 708
rect 2025 706 2193 718
rect 2208 708 2224 722
rect 2259 709 2281 728
rect 2291 715 2307 723
rect 2281 708 2287 709
rect 2290 708 2319 715
rect 2208 707 2319 708
rect 2208 706 2325 707
rect 1884 698 1935 706
rect 1982 698 2016 706
rect 1884 686 1909 698
rect 1916 686 1935 698
rect 1989 696 2016 698
rect 2025 696 2246 706
rect 2281 703 2287 706
rect 1989 692 2246 696
rect 1884 678 1935 686
rect 1982 678 2246 692
rect 2290 698 2325 706
rect 1836 630 1855 664
rect 1900 670 1929 678
rect 1900 664 1917 670
rect 1900 662 1934 664
rect 1982 662 1998 678
rect 1999 668 2207 678
rect 2208 668 2224 678
rect 2272 674 2287 689
rect 2290 686 2291 698
rect 2298 686 2325 698
rect 2290 678 2325 686
rect 2290 677 2319 678
rect 2010 664 2224 668
rect 2025 662 2224 664
rect 2259 664 2272 674
rect 2290 664 2307 677
rect 2259 662 2307 664
rect 1901 658 1934 662
rect 1897 656 1934 658
rect 1897 655 1964 656
rect 1897 650 1928 655
rect 1934 650 1964 655
rect 1897 646 1964 650
rect 1870 643 1964 646
rect 1870 636 1919 643
rect 1870 630 1900 636
rect 1919 631 1924 636
rect 1836 614 1916 630
rect 1928 622 1964 643
rect 2025 638 2214 662
rect 2259 661 2306 662
rect 2272 656 2306 661
rect 2040 635 2214 638
rect 2033 632 2214 635
rect 2242 655 2306 656
rect 1836 612 1855 614
rect 1870 612 1904 614
rect 1836 596 1916 612
rect 1836 590 1855 596
rect 1827 584 1855 590
rect 1870 584 1900 596
rect 1928 584 1934 622
rect 1937 616 1956 622
rect 1971 616 2001 624
rect 1937 608 2001 616
rect 1937 592 2017 608
rect 2033 601 2095 632
rect 2111 601 2173 632
rect 2242 630 2291 655
rect 2306 630 2336 648
rect 2205 616 2235 624
rect 2242 622 2352 630
rect 2205 608 2250 616
rect 1937 590 1956 592
rect 1971 590 2017 592
rect 1937 584 2017 590
rect 2044 588 2079 601
rect 2120 598 2157 601
rect 2120 596 2162 598
rect 2049 585 2079 588
rect 2058 584 2065 585
rect 2086 584 2112 590
rect 2127 585 2157 596
rect 2189 592 2251 608
rect 2189 590 2235 592
rect 2189 584 2251 590
rect 2263 584 2269 622
rect 2272 614 2352 622
rect 2272 612 2291 614
rect 2306 612 2340 614
rect 2272 597 2352 612
rect 2272 596 2358 597
rect 2272 584 2291 596
rect 2306 584 2336 596
rect 2364 590 2370 664
rect 2373 590 2392 734
rect 2364 584 2392 590
rect 2407 590 2413 734
rect 2422 664 2435 734
rect 2464 678 2479 706
rect 2416 630 2435 664
rect 2477 646 2479 658
rect 2450 630 2479 646
rect 2416 614 2479 630
rect 2416 612 2435 614
rect 2450 612 2479 614
rect 2416 596 2479 612
rect 2416 590 2435 596
rect 2407 584 2435 590
rect 2450 584 2479 596
rect 1203 566 1238 574
rect 1203 540 1204 566
rect 1211 540 1238 566
rect 1146 522 1176 536
rect 1203 532 1238 540
rect 1240 566 1276 574
rect 1240 540 1255 566
rect 1262 540 1276 566
rect 1240 532 1276 540
rect 1203 522 1232 532
rect 1246 522 1275 532
rect -541 508 1276 522
rect -478 478 -465 508
rect -450 494 -420 508
rect -377 494 -334 508
rect -327 494 -107 508
rect -100 494 -70 508
rect -410 480 -395 492
rect -376 480 -363 494
rect -295 490 -142 494
rect -413 478 -391 480
rect -313 478 -121 490
rect -42 478 -29 508
rect -14 494 16 508
rect 53 478 72 508
rect 87 478 93 508
rect 102 478 115 508
rect 130 494 160 508
rect 203 494 246 508
rect 253 494 473 508
rect 480 494 510 508
rect 170 480 185 492
rect 204 480 217 494
rect 285 490 438 494
rect 167 478 189 480
rect 267 478 459 490
rect 538 478 551 508
rect 566 494 596 508
rect 633 478 652 508
rect 667 478 673 508
rect 682 478 695 508
rect 710 494 740 508
rect 783 494 826 508
rect 833 494 1053 508
rect 1060 494 1090 508
rect 750 480 765 492
rect 784 480 797 494
rect 865 490 1018 494
rect 747 478 769 480
rect 847 478 1039 490
rect 1118 478 1131 508
rect 1146 494 1176 508
rect 1213 478 1232 508
rect 1247 478 1253 508
rect 1262 478 1275 508
rect -541 464 1276 478
rect -478 413 -465 464
rect -413 460 -391 464
rect -420 438 -391 452
rect -338 438 -322 452
rect -284 448 -278 450
rect -271 448 -163 464
rect -156 448 -150 450
rect -142 448 -127 464
rect -61 458 -42 461
rect -420 436 -322 438
rect -295 436 -127 448
rect -112 438 -96 452
rect -61 439 -39 458
rect -29 445 -13 453
rect -39 438 -33 439
rect -30 438 -1 445
rect -112 437 -1 438
rect -112 436 5 437
rect -436 428 -385 436
rect -338 428 -304 436
rect -436 416 -411 428
rect -404 416 -385 428
rect -331 426 -304 428
rect -295 426 -74 436
rect -39 433 -33 436
rect -331 422 -74 426
rect -436 413 -385 416
rect -338 413 -74 422
rect -30 428 5 436
rect -48 413 -33 419
rect -30 416 -29 428
rect -22 416 5 428
rect -30 413 5 416
rect 53 413 72 464
rect 87 413 93 464
rect 102 413 115 464
rect 167 460 189 464
rect 160 438 189 452
rect 242 438 258 452
rect 296 448 302 450
rect 309 448 417 464
rect 424 448 430 450
rect 438 448 453 464
rect 519 458 538 461
rect 160 436 258 438
rect 285 436 453 448
rect 468 438 484 452
rect 519 439 541 458
rect 551 445 567 453
rect 541 438 547 439
rect 550 438 579 445
rect 468 437 579 438
rect 468 436 585 437
rect 144 428 195 436
rect 242 428 276 436
rect 144 416 169 428
rect 176 416 195 428
rect 249 426 276 428
rect 285 426 506 436
rect 541 433 547 436
rect 249 422 506 426
rect 144 413 195 416
rect 242 413 506 422
rect 550 428 585 436
rect 532 413 547 419
rect 550 416 551 428
rect 558 416 585 428
rect 550 413 585 416
rect 633 413 652 464
rect 667 413 673 464
rect 682 413 695 464
rect 747 460 769 464
rect 740 438 769 452
rect 822 438 838 452
rect 876 448 882 450
rect 889 448 997 464
rect 1004 448 1010 450
rect 1018 448 1033 464
rect 1099 458 1118 461
rect 740 436 838 438
rect 865 436 1033 448
rect 1048 438 1064 452
rect 1099 439 1121 458
rect 1131 445 1147 453
rect 1121 438 1127 439
rect 1130 438 1159 445
rect 1048 437 1159 438
rect 1048 436 1165 437
rect 724 428 775 436
rect 822 428 856 436
rect 724 416 749 428
rect 756 416 775 428
rect 829 426 856 428
rect 865 426 1086 436
rect 1121 433 1127 436
rect 829 422 1086 426
rect 822 416 1086 422
rect 1130 428 1165 436
rect 1112 416 1127 419
rect 1130 416 1131 428
rect 1138 416 1165 428
rect 1213 416 1232 464
rect 1247 416 1253 464
rect 1262 416 1275 464
rect 724 413 757 416
<< nwell >>
rect -295 1718 -142 1814
rect 285 1718 438 1814
rect -295 1448 -142 1544
rect 285 1448 438 1544
rect -295 1178 -142 1274
rect 285 1178 438 1274
rect -295 908 -142 1004
rect 285 908 438 1004
rect -295 638 -142 734
rect 285 638 438 734
rect -295 368 -142 464
rect 285 368 438 464
rect -295 98 -142 194
rect 285 98 438 194
rect -295 -172 -142 -76
rect 285 -172 438 -76
rect -295 -442 -142 -346
rect 285 -442 438 -346
rect -295 -712 -142 -616
rect 285 -712 438 -616
rect -295 -982 -142 -886
rect 285 -982 438 -886
rect -295 -1252 -142 -1156
rect 285 -1252 438 -1156
rect -295 -1522 -142 -1426
rect 285 -1522 438 -1426
rect -295 -1792 -142 -1696
rect 285 -1792 438 -1696
rect -295 -2062 -142 -1966
rect 285 -2062 438 -1966
rect -295 -2332 -142 -2236
rect 285 -2332 438 -2236
rect 865 1718 1018 1814
rect 1445 1718 1598 1814
rect 865 1448 1018 1544
rect 1445 1448 1598 1544
rect 865 1178 1018 1274
rect 1445 1178 1598 1274
rect 865 908 1018 1004
rect 1445 908 1598 1004
rect 865 638 1018 734
rect 1445 638 1598 734
rect 865 368 1018 464
rect 1445 368 1598 464
rect 865 98 1018 194
rect 1445 98 1598 194
rect 865 -172 1018 -76
rect 1445 -172 1598 -76
rect 865 -442 1018 -346
rect 1445 -442 1598 -346
rect 865 -712 1018 -616
rect 1445 -712 1598 -616
rect 865 -982 1018 -886
rect 1445 -982 1598 -886
rect 865 -1252 1018 -1156
rect 1445 -1252 1598 -1156
rect 865 -1522 1018 -1426
rect 1445 -1522 1598 -1426
rect 865 -1792 1018 -1696
rect 1445 -1792 1598 -1696
rect 865 -2062 1018 -1966
rect 1445 -2062 1598 -1966
rect 865 -2332 1018 -2236
rect 1445 -2332 1598 -2236
rect 2025 1718 2178 1814
rect 2605 1718 2758 1814
rect 2025 1448 2178 1544
rect 2605 1448 2758 1544
rect 2025 1178 2178 1274
rect 2605 1178 2758 1274
rect 2025 908 2178 1004
rect 2605 908 2758 1004
rect 2025 638 2178 734
rect 2605 638 2758 734
rect 2025 368 2178 464
rect 2605 368 2758 464
rect 2025 98 2178 194
rect 2605 98 2758 194
rect 2025 -172 2178 -76
rect 2605 -172 2758 -76
rect 2025 -442 2178 -346
rect 2605 -442 2758 -346
rect 2025 -712 2178 -616
rect 2605 -712 2758 -616
rect 2025 -982 2178 -886
rect 2605 -982 2758 -886
rect 2025 -1252 2178 -1156
rect 2605 -1252 2758 -1156
rect 2025 -1522 2178 -1426
rect 2605 -1522 2758 -1426
rect 2025 -1792 2178 -1696
rect 2605 -1792 2758 -1696
rect 2025 -2062 2178 -1966
rect 2605 -2062 2758 -1966
rect 2025 -2332 2178 -2236
rect 2605 -2332 2758 -2236
rect 3185 1718 3338 1814
rect 3765 1718 3918 1814
rect 3185 1448 3338 1544
rect 3765 1448 3918 1544
rect 3185 1178 3338 1274
rect 3765 1178 3918 1274
rect 3185 908 3338 1004
rect 3765 908 3918 1004
rect 3185 638 3338 734
rect 3765 638 3918 734
rect 3185 368 3338 464
rect 3765 368 3918 464
rect 3185 98 3338 194
rect 3765 98 3918 194
rect 3185 -172 3338 -76
rect 3765 -172 3918 -76
rect 3185 -442 3338 -346
rect 3765 -442 3918 -346
rect 3185 -712 3338 -616
rect 3765 -712 3918 -616
rect 3185 -982 3338 -886
rect 3765 -982 3918 -886
rect 3185 -1252 3338 -1156
rect 3765 -1252 3918 -1156
rect 3185 -1522 3338 -1426
rect 3765 -1522 3918 -1426
rect 3185 -1792 3338 -1696
rect 3765 -1792 3918 -1696
rect 3185 -2062 3338 -1966
rect 3765 -2062 3918 -1966
rect 3185 -2332 3338 -2236
rect 3765 -2332 3918 -2236
rect 4345 1718 4498 1814
rect 4925 1718 5078 1814
rect 4345 1448 4498 1544
rect 4925 1448 5078 1544
rect 4345 1178 4498 1274
rect 4925 1178 5078 1274
rect 4345 908 4498 1004
rect 4925 908 5078 1004
rect 4345 638 4498 734
rect 4925 638 5078 734
rect 4345 368 4498 464
rect 4925 368 5078 464
rect 4345 98 4498 194
rect 4925 98 5078 194
rect 4345 -172 4498 -76
rect 4925 -172 5078 -76
rect 4345 -442 4498 -346
rect 4925 -442 5078 -346
rect 4345 -712 4498 -616
rect 4925 -712 5078 -616
rect 4345 -982 4498 -886
rect 4925 -982 5078 -886
rect 4345 -1252 4498 -1156
rect 4925 -1252 5078 -1156
rect 4345 -1522 4498 -1426
rect 4925 -1522 5078 -1426
rect 4345 -1792 4498 -1696
rect 4925 -1792 5078 -1696
rect 4345 -2062 4498 -1966
rect 4925 -2062 5078 -1966
rect 4345 -2332 4498 -2236
rect 4925 -2332 5078 -2236
rect 5505 1718 5658 1814
rect 6085 1718 6238 1814
rect 5505 1448 5658 1544
rect 6085 1448 6238 1544
rect 5505 1178 5658 1274
rect 6085 1178 6238 1274
rect 5505 908 5658 1004
rect 6085 908 6238 1004
rect 5505 638 5658 734
rect 6085 638 6238 734
rect 5505 368 5658 464
rect 6085 368 6238 464
rect 5505 98 5658 194
rect 6085 98 6238 194
rect 5505 -172 5658 -76
rect 6085 -172 6238 -76
rect 5505 -442 5658 -346
rect 6085 -442 6238 -346
rect 5505 -712 5658 -616
rect 6085 -712 6238 -616
rect 5505 -982 5658 -886
rect 6085 -982 6238 -886
rect 5505 -1252 5658 -1156
rect 6085 -1252 6238 -1156
rect 5505 -1522 5658 -1426
rect 6085 -1522 6238 -1426
rect 5505 -1792 5658 -1696
rect 6085 -1792 6238 -1696
rect 5505 -2062 5658 -1966
rect 6085 -2062 6238 -1966
rect 5505 -2332 5658 -2236
rect 6085 -2332 6238 -2236
<< pwell >>
rect -493 1672 -323 1844
rect -111 1672 257 1844
rect 469 1672 639 1844
rect -493 1574 639 1672
rect -493 1402 -323 1574
rect -111 1402 257 1574
rect 469 1402 639 1574
rect -493 1304 639 1402
rect -493 1132 -323 1304
rect -111 1132 257 1304
rect 469 1132 639 1304
rect -493 1034 639 1132
rect -493 862 -323 1034
rect -111 862 257 1034
rect 469 862 639 1034
rect -493 764 639 862
rect -493 592 -323 764
rect -111 592 257 764
rect 469 592 639 764
rect -493 494 639 592
rect -493 322 -323 494
rect -111 322 257 494
rect 469 322 639 494
rect -493 224 639 322
rect -493 52 -323 224
rect -111 52 257 224
rect 469 52 639 224
rect -493 -46 639 52
rect -493 -218 -323 -46
rect -111 -218 257 -46
rect 469 -218 639 -46
rect -493 -316 639 -218
rect -493 -488 -323 -316
rect -111 -488 257 -316
rect 469 -488 639 -316
rect -493 -586 639 -488
rect -493 -758 -323 -586
rect -111 -758 257 -586
rect 469 -758 639 -586
rect -493 -856 639 -758
rect -493 -1028 -323 -856
rect -111 -1028 257 -856
rect 469 -1028 639 -856
rect -493 -1126 639 -1028
rect -493 -1298 -323 -1126
rect -111 -1298 257 -1126
rect 469 -1298 639 -1126
rect -493 -1396 639 -1298
rect -493 -1568 -323 -1396
rect -111 -1568 257 -1396
rect 469 -1568 639 -1396
rect -493 -1666 639 -1568
rect -493 -1838 -323 -1666
rect -111 -1838 257 -1666
rect 469 -1838 639 -1666
rect -493 -1936 639 -1838
rect -493 -2108 -323 -1936
rect -111 -2108 257 -1936
rect 469 -2108 639 -1936
rect -493 -2206 639 -2108
rect -493 -2378 -323 -2206
rect -111 -2378 257 -2206
rect 469 -2378 639 -2206
rect -493 -2476 639 -2378
rect 667 1672 837 1844
rect 1049 1672 1417 1844
rect 1629 1672 1799 1844
rect 667 1574 1799 1672
rect 667 1402 837 1574
rect 1049 1402 1417 1574
rect 1629 1402 1799 1574
rect 667 1304 1799 1402
rect 667 1132 837 1304
rect 1049 1132 1417 1304
rect 1629 1132 1799 1304
rect 667 1034 1799 1132
rect 667 862 837 1034
rect 1049 862 1417 1034
rect 1629 862 1799 1034
rect 667 764 1799 862
rect 667 592 837 764
rect 1049 592 1417 764
rect 1629 592 1799 764
rect 667 494 1799 592
rect 667 322 837 494
rect 1049 322 1417 494
rect 1629 322 1799 494
rect 667 224 1799 322
rect 667 52 837 224
rect 1049 52 1417 224
rect 1629 52 1799 224
rect 667 -46 1799 52
rect 667 -218 837 -46
rect 1049 -218 1417 -46
rect 1629 -218 1799 -46
rect 667 -316 1799 -218
rect 667 -488 837 -316
rect 1049 -488 1417 -316
rect 1629 -488 1799 -316
rect 667 -586 1799 -488
rect 667 -758 837 -586
rect 1049 -758 1417 -586
rect 1629 -758 1799 -586
rect 667 -856 1799 -758
rect 667 -1028 837 -856
rect 1049 -1028 1417 -856
rect 1629 -1028 1799 -856
rect 667 -1126 1799 -1028
rect 667 -1298 837 -1126
rect 1049 -1298 1417 -1126
rect 1629 -1298 1799 -1126
rect 667 -1396 1799 -1298
rect 667 -1568 837 -1396
rect 1049 -1568 1417 -1396
rect 1629 -1568 1799 -1396
rect 667 -1666 1799 -1568
rect 667 -1838 837 -1666
rect 1049 -1838 1417 -1666
rect 1629 -1838 1799 -1666
rect 667 -1936 1799 -1838
rect 667 -2108 837 -1936
rect 1049 -2108 1417 -1936
rect 1629 -2108 1799 -1936
rect 667 -2206 1799 -2108
rect 667 -2378 837 -2206
rect 1049 -2378 1417 -2206
rect 1629 -2378 1799 -2206
rect 667 -2476 1799 -2378
rect 1827 1672 1997 1844
rect 2209 1672 2577 1844
rect 2789 1672 2959 1844
rect 1827 1574 2959 1672
rect 1827 1402 1997 1574
rect 2209 1402 2577 1574
rect 2789 1402 2959 1574
rect 1827 1304 2959 1402
rect 1827 1132 1997 1304
rect 2209 1132 2577 1304
rect 2789 1132 2959 1304
rect 1827 1034 2959 1132
rect 1827 862 1997 1034
rect 2209 862 2577 1034
rect 2789 862 2959 1034
rect 1827 764 2959 862
rect 1827 592 1997 764
rect 2209 592 2577 764
rect 2789 592 2959 764
rect 1827 494 2959 592
rect 1827 322 1997 494
rect 2209 322 2577 494
rect 2789 322 2959 494
rect 1827 224 2959 322
rect 1827 52 1997 224
rect 2209 52 2577 224
rect 2789 52 2959 224
rect 1827 -46 2959 52
rect 1827 -218 1997 -46
rect 2209 -218 2577 -46
rect 2789 -218 2959 -46
rect 1827 -316 2959 -218
rect 1827 -488 1997 -316
rect 2209 -488 2577 -316
rect 2789 -488 2959 -316
rect 1827 -586 2959 -488
rect 1827 -758 1997 -586
rect 2209 -758 2577 -586
rect 2789 -758 2959 -586
rect 1827 -856 2959 -758
rect 1827 -1028 1997 -856
rect 2209 -1028 2577 -856
rect 2789 -1028 2959 -856
rect 1827 -1126 2959 -1028
rect 1827 -1298 1997 -1126
rect 2209 -1298 2577 -1126
rect 2789 -1298 2959 -1126
rect 1827 -1396 2959 -1298
rect 1827 -1568 1997 -1396
rect 2209 -1568 2577 -1396
rect 2789 -1568 2959 -1396
rect 1827 -1666 2959 -1568
rect 1827 -1838 1997 -1666
rect 2209 -1838 2577 -1666
rect 2789 -1838 2959 -1666
rect 1827 -1936 2959 -1838
rect 1827 -2108 1997 -1936
rect 2209 -2108 2577 -1936
rect 2789 -2108 2959 -1936
rect 1827 -2206 2959 -2108
rect 1827 -2378 1997 -2206
rect 2209 -2378 2577 -2206
rect 2789 -2378 2959 -2206
rect 1827 -2476 2959 -2378
rect 2987 1672 3157 1844
rect 3369 1672 3737 1844
rect 3949 1672 4119 1844
rect 2987 1574 4119 1672
rect 2987 1402 3157 1574
rect 3369 1402 3737 1574
rect 3949 1402 4119 1574
rect 2987 1304 4119 1402
rect 2987 1132 3157 1304
rect 3369 1132 3737 1304
rect 3949 1132 4119 1304
rect 2987 1034 4119 1132
rect 2987 862 3157 1034
rect 3369 862 3737 1034
rect 3949 862 4119 1034
rect 2987 764 4119 862
rect 2987 592 3157 764
rect 3369 592 3737 764
rect 3949 592 4119 764
rect 2987 494 4119 592
rect 2987 322 3157 494
rect 3369 322 3737 494
rect 3949 322 4119 494
rect 2987 224 4119 322
rect 2987 52 3157 224
rect 3369 52 3737 224
rect 3949 52 4119 224
rect 2987 -46 4119 52
rect 2987 -218 3157 -46
rect 3369 -218 3737 -46
rect 3949 -218 4119 -46
rect 2987 -316 4119 -218
rect 2987 -488 3157 -316
rect 3369 -488 3737 -316
rect 3949 -488 4119 -316
rect 2987 -586 4119 -488
rect 2987 -758 3157 -586
rect 3369 -758 3737 -586
rect 3949 -758 4119 -586
rect 2987 -856 4119 -758
rect 2987 -1028 3157 -856
rect 3369 -1028 3737 -856
rect 3949 -1028 4119 -856
rect 2987 -1126 4119 -1028
rect 2987 -1298 3157 -1126
rect 3369 -1298 3737 -1126
rect 3949 -1298 4119 -1126
rect 2987 -1396 4119 -1298
rect 2987 -1568 3157 -1396
rect 3369 -1568 3737 -1396
rect 3949 -1568 4119 -1396
rect 2987 -1666 4119 -1568
rect 2987 -1838 3157 -1666
rect 3369 -1838 3737 -1666
rect 3949 -1838 4119 -1666
rect 2987 -1936 4119 -1838
rect 2987 -2108 3157 -1936
rect 3369 -2108 3737 -1936
rect 3949 -2108 4119 -1936
rect 2987 -2206 4119 -2108
rect 2987 -2378 3157 -2206
rect 3369 -2378 3737 -2206
rect 3949 -2378 4119 -2206
rect 2987 -2476 4119 -2378
rect 4147 1672 4317 1844
rect 4529 1672 4897 1844
rect 5109 1672 5279 1844
rect 4147 1574 5279 1672
rect 4147 1402 4317 1574
rect 4529 1402 4897 1574
rect 5109 1402 5279 1574
rect 4147 1304 5279 1402
rect 4147 1132 4317 1304
rect 4529 1132 4897 1304
rect 5109 1132 5279 1304
rect 4147 1034 5279 1132
rect 4147 862 4317 1034
rect 4529 862 4897 1034
rect 5109 862 5279 1034
rect 4147 764 5279 862
rect 4147 592 4317 764
rect 4529 592 4897 764
rect 5109 592 5279 764
rect 4147 494 5279 592
rect 4147 322 4317 494
rect 4529 322 4897 494
rect 5109 322 5279 494
rect 4147 224 5279 322
rect 4147 52 4317 224
rect 4529 52 4897 224
rect 5109 52 5279 224
rect 4147 -46 5279 52
rect 4147 -218 4317 -46
rect 4529 -218 4897 -46
rect 5109 -218 5279 -46
rect 4147 -316 5279 -218
rect 4147 -488 4317 -316
rect 4529 -488 4897 -316
rect 5109 -488 5279 -316
rect 4147 -586 5279 -488
rect 4147 -758 4317 -586
rect 4529 -758 4897 -586
rect 5109 -758 5279 -586
rect 4147 -856 5279 -758
rect 4147 -1028 4317 -856
rect 4529 -1028 4897 -856
rect 5109 -1028 5279 -856
rect 4147 -1126 5279 -1028
rect 4147 -1298 4317 -1126
rect 4529 -1298 4897 -1126
rect 5109 -1298 5279 -1126
rect 4147 -1396 5279 -1298
rect 4147 -1568 4317 -1396
rect 4529 -1568 4897 -1396
rect 5109 -1568 5279 -1396
rect 4147 -1666 5279 -1568
rect 4147 -1838 4317 -1666
rect 4529 -1838 4897 -1666
rect 5109 -1838 5279 -1666
rect 4147 -1936 5279 -1838
rect 4147 -2108 4317 -1936
rect 4529 -2108 4897 -1936
rect 5109 -2108 5279 -1936
rect 4147 -2206 5279 -2108
rect 4147 -2378 4317 -2206
rect 4529 -2378 4897 -2206
rect 5109 -2378 5279 -2206
rect 4147 -2476 5279 -2378
rect 5307 1672 5477 1844
rect 5689 1672 6057 1844
rect 6269 1672 6439 1844
rect 5307 1574 6439 1672
rect 5307 1402 5477 1574
rect 5689 1402 6057 1574
rect 6269 1402 6439 1574
rect 5307 1304 6439 1402
rect 5307 1132 5477 1304
rect 5689 1132 6057 1304
rect 6269 1132 6439 1304
rect 5307 1034 6439 1132
rect 5307 862 5477 1034
rect 5689 862 6057 1034
rect 6269 862 6439 1034
rect 5307 764 6439 862
rect 5307 592 5477 764
rect 5689 592 6057 764
rect 6269 592 6439 764
rect 5307 494 6439 592
rect 5307 322 5477 494
rect 5689 322 6057 494
rect 6269 322 6439 494
rect 5307 224 6439 322
rect 5307 52 5477 224
rect 5689 52 6057 224
rect 6269 52 6439 224
rect 5307 -46 6439 52
rect 5307 -218 5477 -46
rect 5689 -218 6057 -46
rect 6269 -218 6439 -46
rect 5307 -316 6439 -218
rect 5307 -488 5477 -316
rect 5689 -488 6057 -316
rect 6269 -488 6439 -316
rect 5307 -586 6439 -488
rect 5307 -758 5477 -586
rect 5689 -758 6057 -586
rect 6269 -758 6439 -586
rect 5307 -856 6439 -758
rect 5307 -1028 5477 -856
rect 5689 -1028 6057 -856
rect 6269 -1028 6439 -856
rect 5307 -1126 6439 -1028
rect 5307 -1298 5477 -1126
rect 5689 -1298 6057 -1126
rect 6269 -1298 6439 -1126
rect 5307 -1396 6439 -1298
rect 5307 -1568 5477 -1396
rect 5689 -1568 6057 -1396
rect 6269 -1568 6439 -1396
rect 5307 -1666 6439 -1568
rect 5307 -1838 5477 -1666
rect 5689 -1838 6057 -1666
rect 6269 -1838 6439 -1666
rect 5307 -1936 6439 -1838
rect 5307 -2108 5477 -1936
rect 5689 -2108 6057 -1936
rect 6269 -2108 6439 -1936
rect 5307 -2206 6439 -2108
rect 5307 -2378 5477 -2206
rect 5689 -2378 6057 -2206
rect 6269 -2378 6439 -2206
rect 5307 -2476 6439 -2378
<< nmos >>
rect -386 1758 -356 1786
rect -78 1758 -48 1786
rect 194 1758 224 1786
rect 502 1758 532 1786
rect 774 1758 804 1786
rect 1082 1758 1112 1786
rect 1354 1758 1384 1786
rect 1662 1758 1692 1786
rect 1934 1758 1964 1786
rect 2242 1758 2272 1786
rect 2514 1758 2544 1786
rect 2822 1758 2852 1786
rect 3094 1758 3124 1786
rect 3402 1758 3432 1786
rect 3674 1758 3704 1786
rect 3982 1758 4012 1786
rect 4254 1758 4284 1786
rect 4562 1758 4592 1786
rect 4834 1758 4864 1786
rect 5142 1758 5172 1786
rect 5414 1758 5444 1786
rect 5722 1758 5752 1786
rect 5994 1758 6024 1786
rect 6302 1758 6332 1786
rect -450 1612 -420 1654
rect -14 1612 16 1654
rect 130 1612 160 1654
rect 566 1612 596 1654
rect 710 1612 740 1654
rect 1146 1612 1176 1654
rect 1290 1612 1320 1654
rect 1726 1612 1756 1654
rect 1870 1612 1900 1654
rect 2306 1612 2336 1654
rect 2450 1612 2480 1654
rect 2886 1612 2916 1654
rect 3030 1612 3060 1654
rect 3466 1612 3496 1654
rect 3610 1612 3640 1654
rect 4046 1612 4076 1654
rect 4190 1612 4220 1654
rect 4626 1612 4656 1654
rect 4770 1612 4800 1654
rect 5206 1612 5236 1654
rect 5350 1612 5380 1654
rect 5786 1612 5816 1654
rect 5930 1612 5960 1654
rect 6366 1612 6396 1654
rect -386 1488 -356 1516
rect -78 1488 -48 1516
rect 194 1488 224 1516
rect 502 1488 532 1516
rect 774 1488 804 1516
rect 1082 1488 1112 1516
rect 1354 1488 1384 1516
rect 1662 1488 1692 1516
rect 1934 1488 1964 1516
rect 2242 1488 2272 1516
rect 2514 1488 2544 1516
rect 2822 1488 2852 1516
rect 3094 1488 3124 1516
rect 3402 1488 3432 1516
rect 3674 1488 3704 1516
rect 3982 1488 4012 1516
rect 4254 1488 4284 1516
rect 4562 1488 4592 1516
rect 4834 1488 4864 1516
rect 5142 1488 5172 1516
rect 5414 1488 5444 1516
rect 5722 1488 5752 1516
rect 5994 1488 6024 1516
rect 6302 1488 6332 1516
rect -450 1342 -420 1384
rect -14 1342 16 1384
rect 130 1342 160 1384
rect 566 1342 596 1384
rect 710 1342 740 1384
rect 1146 1342 1176 1384
rect 1290 1342 1320 1384
rect 1726 1342 1756 1384
rect 1870 1342 1900 1384
rect 2306 1342 2336 1384
rect 2450 1342 2480 1384
rect 2886 1342 2916 1384
rect 3030 1342 3060 1384
rect 3466 1342 3496 1384
rect 3610 1342 3640 1384
rect 4046 1342 4076 1384
rect 4190 1342 4220 1384
rect 4626 1342 4656 1384
rect 4770 1342 4800 1384
rect 5206 1342 5236 1384
rect 5350 1342 5380 1384
rect 5786 1342 5816 1384
rect 5930 1342 5960 1384
rect 6366 1342 6396 1384
rect -386 1218 -356 1246
rect -78 1218 -48 1246
rect 194 1218 224 1246
rect 502 1218 532 1246
rect 774 1218 804 1246
rect 1082 1218 1112 1246
rect 1354 1218 1384 1246
rect 1662 1218 1692 1246
rect 1934 1218 1964 1246
rect 2242 1218 2272 1246
rect 2514 1218 2544 1246
rect 2822 1218 2852 1246
rect 3094 1218 3124 1246
rect 3402 1218 3432 1246
rect 3674 1218 3704 1246
rect 3982 1218 4012 1246
rect 4254 1218 4284 1246
rect 4562 1218 4592 1246
rect 4834 1218 4864 1246
rect 5142 1218 5172 1246
rect 5414 1218 5444 1246
rect 5722 1218 5752 1246
rect 5994 1218 6024 1246
rect 6302 1218 6332 1246
rect -450 1072 -420 1114
rect -14 1072 16 1114
rect 130 1072 160 1114
rect 566 1072 596 1114
rect 710 1072 740 1114
rect 1146 1072 1176 1114
rect 1290 1072 1320 1114
rect 1726 1072 1756 1114
rect 1870 1072 1900 1114
rect 2306 1072 2336 1114
rect 2450 1072 2480 1114
rect 2886 1072 2916 1114
rect 3030 1072 3060 1114
rect 3466 1072 3496 1114
rect 3610 1072 3640 1114
rect 4046 1072 4076 1114
rect 4190 1072 4220 1114
rect 4626 1072 4656 1114
rect 4770 1072 4800 1114
rect 5206 1072 5236 1114
rect 5350 1072 5380 1114
rect 5786 1072 5816 1114
rect 5930 1072 5960 1114
rect 6366 1072 6396 1114
rect -386 948 -356 976
rect -78 948 -48 976
rect 194 948 224 976
rect 502 948 532 976
rect 774 948 804 976
rect 1082 948 1112 976
rect 1354 948 1384 976
rect 1662 948 1692 976
rect 1934 948 1964 976
rect 2242 948 2272 976
rect 2514 948 2544 976
rect 2822 948 2852 976
rect 3094 948 3124 976
rect 3402 948 3432 976
rect 3674 948 3704 976
rect 3982 948 4012 976
rect 4254 948 4284 976
rect 4562 948 4592 976
rect 4834 948 4864 976
rect 5142 948 5172 976
rect 5414 948 5444 976
rect 5722 948 5752 976
rect 5994 948 6024 976
rect 6302 948 6332 976
rect -450 802 -420 844
rect -14 802 16 844
rect 130 802 160 844
rect 566 802 596 844
rect 710 802 740 844
rect 1146 802 1176 844
rect 1290 802 1320 844
rect 1726 802 1756 844
rect 1870 802 1900 844
rect 2306 802 2336 844
rect 2450 802 2480 844
rect 2886 802 2916 844
rect 3030 802 3060 844
rect 3466 802 3496 844
rect 3610 802 3640 844
rect 4046 802 4076 844
rect 4190 802 4220 844
rect 4626 802 4656 844
rect 4770 802 4800 844
rect 5206 802 5236 844
rect 5350 802 5380 844
rect 5786 802 5816 844
rect 5930 802 5960 844
rect 6366 802 6396 844
rect -386 678 -356 706
rect -78 678 -48 706
rect 194 678 224 706
rect 502 678 532 706
rect 774 678 804 706
rect 1082 678 1112 706
rect 1354 678 1384 706
rect 1662 678 1692 706
rect 1934 678 1964 706
rect 2242 678 2272 706
rect 2514 678 2544 706
rect 2822 678 2852 706
rect 3094 678 3124 706
rect 3402 678 3432 706
rect 3674 678 3704 706
rect 3982 678 4012 706
rect 4254 678 4284 706
rect 4562 678 4592 706
rect 4834 678 4864 706
rect 5142 678 5172 706
rect 5414 678 5444 706
rect 5722 678 5752 706
rect 5994 678 6024 706
rect 6302 678 6332 706
rect -450 532 -420 574
rect -14 532 16 574
rect 130 532 160 574
rect 566 532 596 574
rect 710 532 740 574
rect 1146 532 1176 574
rect 1290 532 1320 574
rect 1726 532 1756 574
rect 1870 532 1900 574
rect 2306 532 2336 574
rect 2450 532 2480 574
rect 2886 532 2916 574
rect 3030 532 3060 574
rect 3466 532 3496 574
rect 3610 532 3640 574
rect 4046 532 4076 574
rect 4190 532 4220 574
rect 4626 532 4656 574
rect 4770 532 4800 574
rect 5206 532 5236 574
rect 5350 532 5380 574
rect 5786 532 5816 574
rect 5930 532 5960 574
rect 6366 532 6396 574
rect -386 408 -356 436
rect -78 408 -48 436
rect 194 408 224 436
rect 502 408 532 436
rect 774 408 804 436
rect 1082 408 1112 436
rect 1354 408 1384 436
rect 1662 408 1692 436
rect 1934 408 1964 436
rect 2242 408 2272 436
rect 2514 408 2544 436
rect 2822 408 2852 436
rect 3094 408 3124 436
rect 3402 408 3432 436
rect 3674 408 3704 436
rect 3982 408 4012 436
rect 4254 408 4284 436
rect 4562 408 4592 436
rect 4834 408 4864 436
rect 5142 408 5172 436
rect 5414 408 5444 436
rect 5722 408 5752 436
rect 5994 408 6024 436
rect 6302 408 6332 436
rect -450 262 -420 304
rect -14 262 16 304
rect 130 262 160 304
rect 566 262 596 304
rect 710 262 740 304
rect 1146 262 1176 304
rect 1290 262 1320 304
rect 1726 262 1756 304
rect 1870 262 1900 304
rect 2306 262 2336 304
rect 2450 262 2480 304
rect 2886 262 2916 304
rect 3030 262 3060 304
rect 3466 262 3496 304
rect 3610 262 3640 304
rect 4046 262 4076 304
rect 4190 262 4220 304
rect 4626 262 4656 304
rect 4770 262 4800 304
rect 5206 262 5236 304
rect 5350 262 5380 304
rect 5786 262 5816 304
rect 5930 262 5960 304
rect 6366 262 6396 304
rect -386 138 -356 166
rect -78 138 -48 166
rect 194 138 224 166
rect 502 138 532 166
rect 774 138 804 166
rect 1082 138 1112 166
rect 1354 138 1384 166
rect 1662 138 1692 166
rect 1934 138 1964 166
rect 2242 138 2272 166
rect 2514 138 2544 166
rect 2822 138 2852 166
rect 3094 138 3124 166
rect 3402 138 3432 166
rect 3674 138 3704 166
rect 3982 138 4012 166
rect 4254 138 4284 166
rect 4562 138 4592 166
rect 4834 138 4864 166
rect 5142 138 5172 166
rect 5414 138 5444 166
rect 5722 138 5752 166
rect 5994 138 6024 166
rect 6302 138 6332 166
rect -450 -8 -420 34
rect -14 -8 16 34
rect 130 -8 160 34
rect 566 -8 596 34
rect 710 -8 740 34
rect 1146 -8 1176 34
rect 1290 -8 1320 34
rect 1726 -8 1756 34
rect 1870 -8 1900 34
rect 2306 -8 2336 34
rect 2450 -8 2480 34
rect 2886 -8 2916 34
rect 3030 -8 3060 34
rect 3466 -8 3496 34
rect 3610 -8 3640 34
rect 4046 -8 4076 34
rect 4190 -8 4220 34
rect 4626 -8 4656 34
rect 4770 -8 4800 34
rect 5206 -8 5236 34
rect 5350 -8 5380 34
rect 5786 -8 5816 34
rect 5930 -8 5960 34
rect 6366 -8 6396 34
rect -386 -132 -356 -104
rect -78 -132 -48 -104
rect 194 -132 224 -104
rect 502 -132 532 -104
rect 774 -132 804 -104
rect 1082 -132 1112 -104
rect 1354 -132 1384 -104
rect 1662 -132 1692 -104
rect 1934 -132 1964 -104
rect 2242 -132 2272 -104
rect 2514 -132 2544 -104
rect 2822 -132 2852 -104
rect 3094 -132 3124 -104
rect 3402 -132 3432 -104
rect 3674 -132 3704 -104
rect 3982 -132 4012 -104
rect 4254 -132 4284 -104
rect 4562 -132 4592 -104
rect 4834 -132 4864 -104
rect 5142 -132 5172 -104
rect 5414 -132 5444 -104
rect 5722 -132 5752 -104
rect 5994 -132 6024 -104
rect 6302 -132 6332 -104
rect -450 -278 -420 -236
rect -14 -278 16 -236
rect 130 -278 160 -236
rect 566 -278 596 -236
rect 710 -278 740 -236
rect 1146 -278 1176 -236
rect 1290 -278 1320 -236
rect 1726 -278 1756 -236
rect 1870 -278 1900 -236
rect 2306 -278 2336 -236
rect 2450 -278 2480 -236
rect 2886 -278 2916 -236
rect 3030 -278 3060 -236
rect 3466 -278 3496 -236
rect 3610 -278 3640 -236
rect 4046 -278 4076 -236
rect 4190 -278 4220 -236
rect 4626 -278 4656 -236
rect 4770 -278 4800 -236
rect 5206 -278 5236 -236
rect 5350 -278 5380 -236
rect 5786 -278 5816 -236
rect 5930 -278 5960 -236
rect 6366 -278 6396 -236
rect -386 -402 -356 -374
rect -78 -402 -48 -374
rect 194 -402 224 -374
rect 502 -402 532 -374
rect 774 -402 804 -374
rect 1082 -402 1112 -374
rect 1354 -402 1384 -374
rect 1662 -402 1692 -374
rect 1934 -402 1964 -374
rect 2242 -402 2272 -374
rect 2514 -402 2544 -374
rect 2822 -402 2852 -374
rect 3094 -402 3124 -374
rect 3402 -402 3432 -374
rect 3674 -402 3704 -374
rect 3982 -402 4012 -374
rect 4254 -402 4284 -374
rect 4562 -402 4592 -374
rect 4834 -402 4864 -374
rect 5142 -402 5172 -374
rect 5414 -402 5444 -374
rect 5722 -402 5752 -374
rect 5994 -402 6024 -374
rect 6302 -402 6332 -374
rect -450 -548 -420 -506
rect -14 -548 16 -506
rect 130 -548 160 -506
rect 566 -548 596 -506
rect 710 -548 740 -506
rect 1146 -548 1176 -506
rect 1290 -548 1320 -506
rect 1726 -548 1756 -506
rect 1870 -548 1900 -506
rect 2306 -548 2336 -506
rect 2450 -548 2480 -506
rect 2886 -548 2916 -506
rect 3030 -548 3060 -506
rect 3466 -548 3496 -506
rect 3610 -548 3640 -506
rect 4046 -548 4076 -506
rect 4190 -548 4220 -506
rect 4626 -548 4656 -506
rect 4770 -548 4800 -506
rect 5206 -548 5236 -506
rect 5350 -548 5380 -506
rect 5786 -548 5816 -506
rect 5930 -548 5960 -506
rect 6366 -548 6396 -506
rect -386 -672 -356 -644
rect -78 -672 -48 -644
rect 194 -672 224 -644
rect 502 -672 532 -644
rect 774 -672 804 -644
rect 1082 -672 1112 -644
rect 1354 -672 1384 -644
rect 1662 -672 1692 -644
rect 1934 -672 1964 -644
rect 2242 -672 2272 -644
rect 2514 -672 2544 -644
rect 2822 -672 2852 -644
rect 3094 -672 3124 -644
rect 3402 -672 3432 -644
rect 3674 -672 3704 -644
rect 3982 -672 4012 -644
rect 4254 -672 4284 -644
rect 4562 -672 4592 -644
rect 4834 -672 4864 -644
rect 5142 -672 5172 -644
rect 5414 -672 5444 -644
rect 5722 -672 5752 -644
rect 5994 -672 6024 -644
rect 6302 -672 6332 -644
rect -450 -818 -420 -776
rect -14 -818 16 -776
rect 130 -818 160 -776
rect 566 -818 596 -776
rect 710 -818 740 -776
rect 1146 -818 1176 -776
rect 1290 -818 1320 -776
rect 1726 -818 1756 -776
rect 1870 -818 1900 -776
rect 2306 -818 2336 -776
rect 2450 -818 2480 -776
rect 2886 -818 2916 -776
rect 3030 -818 3060 -776
rect 3466 -818 3496 -776
rect 3610 -818 3640 -776
rect 4046 -818 4076 -776
rect 4190 -818 4220 -776
rect 4626 -818 4656 -776
rect 4770 -818 4800 -776
rect 5206 -818 5236 -776
rect 5350 -818 5380 -776
rect 5786 -818 5816 -776
rect 5930 -818 5960 -776
rect 6366 -818 6396 -776
rect -386 -942 -356 -914
rect -78 -942 -48 -914
rect 194 -942 224 -914
rect 502 -942 532 -914
rect 774 -942 804 -914
rect 1082 -942 1112 -914
rect 1354 -942 1384 -914
rect 1662 -942 1692 -914
rect 1934 -942 1964 -914
rect 2242 -942 2272 -914
rect 2514 -942 2544 -914
rect 2822 -942 2852 -914
rect 3094 -942 3124 -914
rect 3402 -942 3432 -914
rect 3674 -942 3704 -914
rect 3982 -942 4012 -914
rect 4254 -942 4284 -914
rect 4562 -942 4592 -914
rect 4834 -942 4864 -914
rect 5142 -942 5172 -914
rect 5414 -942 5444 -914
rect 5722 -942 5752 -914
rect 5994 -942 6024 -914
rect 6302 -942 6332 -914
rect -450 -1088 -420 -1046
rect -14 -1088 16 -1046
rect 130 -1088 160 -1046
rect 566 -1088 596 -1046
rect 710 -1088 740 -1046
rect 1146 -1088 1176 -1046
rect 1290 -1088 1320 -1046
rect 1726 -1088 1756 -1046
rect 1870 -1088 1900 -1046
rect 2306 -1088 2336 -1046
rect 2450 -1088 2480 -1046
rect 2886 -1088 2916 -1046
rect 3030 -1088 3060 -1046
rect 3466 -1088 3496 -1046
rect 3610 -1088 3640 -1046
rect 4046 -1088 4076 -1046
rect 4190 -1088 4220 -1046
rect 4626 -1088 4656 -1046
rect 4770 -1088 4800 -1046
rect 5206 -1088 5236 -1046
rect 5350 -1088 5380 -1046
rect 5786 -1088 5816 -1046
rect 5930 -1088 5960 -1046
rect 6366 -1088 6396 -1046
rect -386 -1212 -356 -1184
rect -78 -1212 -48 -1184
rect 194 -1212 224 -1184
rect 502 -1212 532 -1184
rect 774 -1212 804 -1184
rect 1082 -1212 1112 -1184
rect 1354 -1212 1384 -1184
rect 1662 -1212 1692 -1184
rect 1934 -1212 1964 -1184
rect 2242 -1212 2272 -1184
rect 2514 -1212 2544 -1184
rect 2822 -1212 2852 -1184
rect 3094 -1212 3124 -1184
rect 3402 -1212 3432 -1184
rect 3674 -1212 3704 -1184
rect 3982 -1212 4012 -1184
rect 4254 -1212 4284 -1184
rect 4562 -1212 4592 -1184
rect 4834 -1212 4864 -1184
rect 5142 -1212 5172 -1184
rect 5414 -1212 5444 -1184
rect 5722 -1212 5752 -1184
rect 5994 -1212 6024 -1184
rect 6302 -1212 6332 -1184
rect -450 -1358 -420 -1316
rect -14 -1358 16 -1316
rect 130 -1358 160 -1316
rect 566 -1358 596 -1316
rect 710 -1358 740 -1316
rect 1146 -1358 1176 -1316
rect 1290 -1358 1320 -1316
rect 1726 -1358 1756 -1316
rect 1870 -1358 1900 -1316
rect 2306 -1358 2336 -1316
rect 2450 -1358 2480 -1316
rect 2886 -1358 2916 -1316
rect 3030 -1358 3060 -1316
rect 3466 -1358 3496 -1316
rect 3610 -1358 3640 -1316
rect 4046 -1358 4076 -1316
rect 4190 -1358 4220 -1316
rect 4626 -1358 4656 -1316
rect 4770 -1358 4800 -1316
rect 5206 -1358 5236 -1316
rect 5350 -1358 5380 -1316
rect 5786 -1358 5816 -1316
rect 5930 -1358 5960 -1316
rect 6366 -1358 6396 -1316
rect -386 -1482 -356 -1454
rect -78 -1482 -48 -1454
rect 194 -1482 224 -1454
rect 502 -1482 532 -1454
rect 774 -1482 804 -1454
rect 1082 -1482 1112 -1454
rect 1354 -1482 1384 -1454
rect 1662 -1482 1692 -1454
rect 1934 -1482 1964 -1454
rect 2242 -1482 2272 -1454
rect 2514 -1482 2544 -1454
rect 2822 -1482 2852 -1454
rect 3094 -1482 3124 -1454
rect 3402 -1482 3432 -1454
rect 3674 -1482 3704 -1454
rect 3982 -1482 4012 -1454
rect 4254 -1482 4284 -1454
rect 4562 -1482 4592 -1454
rect 4834 -1482 4864 -1454
rect 5142 -1482 5172 -1454
rect 5414 -1482 5444 -1454
rect 5722 -1482 5752 -1454
rect 5994 -1482 6024 -1454
rect 6302 -1482 6332 -1454
rect -450 -1628 -420 -1586
rect -14 -1628 16 -1586
rect 130 -1628 160 -1586
rect 566 -1628 596 -1586
rect 710 -1628 740 -1586
rect 1146 -1628 1176 -1586
rect 1290 -1628 1320 -1586
rect 1726 -1628 1756 -1586
rect 1870 -1628 1900 -1586
rect 2306 -1628 2336 -1586
rect 2450 -1628 2480 -1586
rect 2886 -1628 2916 -1586
rect 3030 -1628 3060 -1586
rect 3466 -1628 3496 -1586
rect 3610 -1628 3640 -1586
rect 4046 -1628 4076 -1586
rect 4190 -1628 4220 -1586
rect 4626 -1628 4656 -1586
rect 4770 -1628 4800 -1586
rect 5206 -1628 5236 -1586
rect 5350 -1628 5380 -1586
rect 5786 -1628 5816 -1586
rect 5930 -1628 5960 -1586
rect 6366 -1628 6396 -1586
rect -386 -1752 -356 -1724
rect -78 -1752 -48 -1724
rect 194 -1752 224 -1724
rect 502 -1752 532 -1724
rect 774 -1752 804 -1724
rect 1082 -1752 1112 -1724
rect 1354 -1752 1384 -1724
rect 1662 -1752 1692 -1724
rect 1934 -1752 1964 -1724
rect 2242 -1752 2272 -1724
rect 2514 -1752 2544 -1724
rect 2822 -1752 2852 -1724
rect 3094 -1752 3124 -1724
rect 3402 -1752 3432 -1724
rect 3674 -1752 3704 -1724
rect 3982 -1752 4012 -1724
rect 4254 -1752 4284 -1724
rect 4562 -1752 4592 -1724
rect 4834 -1752 4864 -1724
rect 5142 -1752 5172 -1724
rect 5414 -1752 5444 -1724
rect 5722 -1752 5752 -1724
rect 5994 -1752 6024 -1724
rect 6302 -1752 6332 -1724
rect -450 -1898 -420 -1856
rect -14 -1898 16 -1856
rect 130 -1898 160 -1856
rect 566 -1898 596 -1856
rect 710 -1898 740 -1856
rect 1146 -1898 1176 -1856
rect 1290 -1898 1320 -1856
rect 1726 -1898 1756 -1856
rect 1870 -1898 1900 -1856
rect 2306 -1898 2336 -1856
rect 2450 -1898 2480 -1856
rect 2886 -1898 2916 -1856
rect 3030 -1898 3060 -1856
rect 3466 -1898 3496 -1856
rect 3610 -1898 3640 -1856
rect 4046 -1898 4076 -1856
rect 4190 -1898 4220 -1856
rect 4626 -1898 4656 -1856
rect 4770 -1898 4800 -1856
rect 5206 -1898 5236 -1856
rect 5350 -1898 5380 -1856
rect 5786 -1898 5816 -1856
rect 5930 -1898 5960 -1856
rect 6366 -1898 6396 -1856
rect -386 -2022 -356 -1994
rect -78 -2022 -48 -1994
rect 194 -2022 224 -1994
rect 502 -2022 532 -1994
rect 774 -2022 804 -1994
rect 1082 -2022 1112 -1994
rect 1354 -2022 1384 -1994
rect 1662 -2022 1692 -1994
rect 1934 -2022 1964 -1994
rect 2242 -2022 2272 -1994
rect 2514 -2022 2544 -1994
rect 2822 -2022 2852 -1994
rect 3094 -2022 3124 -1994
rect 3402 -2022 3432 -1994
rect 3674 -2022 3704 -1994
rect 3982 -2022 4012 -1994
rect 4254 -2022 4284 -1994
rect 4562 -2022 4592 -1994
rect 4834 -2022 4864 -1994
rect 5142 -2022 5172 -1994
rect 5414 -2022 5444 -1994
rect 5722 -2022 5752 -1994
rect 5994 -2022 6024 -1994
rect 6302 -2022 6332 -1994
rect -450 -2168 -420 -2126
rect -14 -2168 16 -2126
rect 130 -2168 160 -2126
rect 566 -2168 596 -2126
rect 710 -2168 740 -2126
rect 1146 -2168 1176 -2126
rect 1290 -2168 1320 -2126
rect 1726 -2168 1756 -2126
rect 1870 -2168 1900 -2126
rect 2306 -2168 2336 -2126
rect 2450 -2168 2480 -2126
rect 2886 -2168 2916 -2126
rect 3030 -2168 3060 -2126
rect 3466 -2168 3496 -2126
rect 3610 -2168 3640 -2126
rect 4046 -2168 4076 -2126
rect 4190 -2168 4220 -2126
rect 4626 -2168 4656 -2126
rect 4770 -2168 4800 -2126
rect 5206 -2168 5236 -2126
rect 5350 -2168 5380 -2126
rect 5786 -2168 5816 -2126
rect 5930 -2168 5960 -2126
rect 6366 -2168 6396 -2126
rect -386 -2292 -356 -2264
rect -78 -2292 -48 -2264
rect 194 -2292 224 -2264
rect 502 -2292 532 -2264
rect 774 -2292 804 -2264
rect 1082 -2292 1112 -2264
rect 1354 -2292 1384 -2264
rect 1662 -2292 1692 -2264
rect 1934 -2292 1964 -2264
rect 2242 -2292 2272 -2264
rect 2514 -2292 2544 -2264
rect 2822 -2292 2852 -2264
rect 3094 -2292 3124 -2264
rect 3402 -2292 3432 -2264
rect 3674 -2292 3704 -2264
rect 3982 -2292 4012 -2264
rect 4254 -2292 4284 -2264
rect 4562 -2292 4592 -2264
rect 4834 -2292 4864 -2264
rect 5142 -2292 5172 -2264
rect 5414 -2292 5444 -2264
rect 5722 -2292 5752 -2264
rect 5994 -2292 6024 -2264
rect 6302 -2292 6332 -2264
rect -450 -2438 -420 -2396
rect -14 -2438 16 -2396
rect 130 -2438 160 -2396
rect 566 -2438 596 -2396
rect 710 -2438 740 -2396
rect 1146 -2438 1176 -2396
rect 1290 -2438 1320 -2396
rect 1726 -2438 1756 -2396
rect 1870 -2438 1900 -2396
rect 2306 -2438 2336 -2396
rect 2450 -2438 2480 -2396
rect 2886 -2438 2916 -2396
rect 3030 -2438 3060 -2396
rect 3466 -2438 3496 -2396
rect 3610 -2438 3640 -2396
rect 4046 -2438 4076 -2396
rect 4190 -2438 4220 -2396
rect 4626 -2438 4656 -2396
rect 4770 -2438 4800 -2396
rect 5206 -2438 5236 -2396
rect 5350 -2438 5380 -2396
rect 5786 -2438 5816 -2396
rect 5930 -2438 5960 -2396
rect 6366 -2438 6396 -2396
<< npd >>
rect -271 1612 -241 1654
rect -193 1612 -163 1654
rect 309 1612 339 1654
rect 387 1612 417 1654
rect 889 1612 919 1654
rect 967 1612 997 1654
rect 1469 1612 1499 1654
rect 1547 1612 1577 1654
rect 2049 1612 2079 1654
rect 2127 1612 2157 1654
rect 2629 1612 2659 1654
rect 2707 1612 2737 1654
rect 3209 1612 3239 1654
rect 3287 1612 3317 1654
rect 3789 1612 3819 1654
rect 3867 1612 3897 1654
rect 4369 1612 4399 1654
rect 4447 1612 4477 1654
rect 4949 1612 4979 1654
rect 5027 1612 5057 1654
rect 5529 1612 5559 1654
rect 5607 1612 5637 1654
rect 6109 1612 6139 1654
rect 6187 1612 6217 1654
rect -271 1342 -241 1384
rect -193 1342 -163 1384
rect 309 1342 339 1384
rect 387 1342 417 1384
rect 889 1342 919 1384
rect 967 1342 997 1384
rect 1469 1342 1499 1384
rect 1547 1342 1577 1384
rect 2049 1342 2079 1384
rect 2127 1342 2157 1384
rect 2629 1342 2659 1384
rect 2707 1342 2737 1384
rect 3209 1342 3239 1384
rect 3287 1342 3317 1384
rect 3789 1342 3819 1384
rect 3867 1342 3897 1384
rect 4369 1342 4399 1384
rect 4447 1342 4477 1384
rect 4949 1342 4979 1384
rect 5027 1342 5057 1384
rect 5529 1342 5559 1384
rect 5607 1342 5637 1384
rect 6109 1342 6139 1384
rect 6187 1342 6217 1384
rect -271 1072 -241 1114
rect -193 1072 -163 1114
rect 309 1072 339 1114
rect 387 1072 417 1114
rect 889 1072 919 1114
rect 967 1072 997 1114
rect 1469 1072 1499 1114
rect 1547 1072 1577 1114
rect 2049 1072 2079 1114
rect 2127 1072 2157 1114
rect 2629 1072 2659 1114
rect 2707 1072 2737 1114
rect 3209 1072 3239 1114
rect 3287 1072 3317 1114
rect 3789 1072 3819 1114
rect 3867 1072 3897 1114
rect 4369 1072 4399 1114
rect 4447 1072 4477 1114
rect 4949 1072 4979 1114
rect 5027 1072 5057 1114
rect 5529 1072 5559 1114
rect 5607 1072 5637 1114
rect 6109 1072 6139 1114
rect 6187 1072 6217 1114
rect -271 802 -241 844
rect -193 802 -163 844
rect 309 802 339 844
rect 387 802 417 844
rect 889 802 919 844
rect 967 802 997 844
rect 1469 802 1499 844
rect 1547 802 1577 844
rect 2049 802 2079 844
rect 2127 802 2157 844
rect 2629 802 2659 844
rect 2707 802 2737 844
rect 3209 802 3239 844
rect 3287 802 3317 844
rect 3789 802 3819 844
rect 3867 802 3897 844
rect 4369 802 4399 844
rect 4447 802 4477 844
rect 4949 802 4979 844
rect 5027 802 5057 844
rect 5529 802 5559 844
rect 5607 802 5637 844
rect 6109 802 6139 844
rect 6187 802 6217 844
rect -271 532 -241 574
rect -193 532 -163 574
rect 309 532 339 574
rect 387 532 417 574
rect 889 532 919 574
rect 967 532 997 574
rect 1469 532 1499 574
rect 1547 532 1577 574
rect 2049 532 2079 574
rect 2127 532 2157 574
rect 2629 532 2659 574
rect 2707 532 2737 574
rect 3209 532 3239 574
rect 3287 532 3317 574
rect 3789 532 3819 574
rect 3867 532 3897 574
rect 4369 532 4399 574
rect 4447 532 4477 574
rect 4949 532 4979 574
rect 5027 532 5057 574
rect 5529 532 5559 574
rect 5607 532 5637 574
rect 6109 532 6139 574
rect 6187 532 6217 574
rect -271 262 -241 304
rect -193 262 -163 304
rect 309 262 339 304
rect 387 262 417 304
rect 889 262 919 304
rect 967 262 997 304
rect 1469 262 1499 304
rect 1547 262 1577 304
rect 2049 262 2079 304
rect 2127 262 2157 304
rect 2629 262 2659 304
rect 2707 262 2737 304
rect 3209 262 3239 304
rect 3287 262 3317 304
rect 3789 262 3819 304
rect 3867 262 3897 304
rect 4369 262 4399 304
rect 4447 262 4477 304
rect 4949 262 4979 304
rect 5027 262 5057 304
rect 5529 262 5559 304
rect 5607 262 5637 304
rect 6109 262 6139 304
rect 6187 262 6217 304
rect -271 -8 -241 34
rect -193 -8 -163 34
rect 309 -8 339 34
rect 387 -8 417 34
rect 889 -8 919 34
rect 967 -8 997 34
rect 1469 -8 1499 34
rect 1547 -8 1577 34
rect 2049 -8 2079 34
rect 2127 -8 2157 34
rect 2629 -8 2659 34
rect 2707 -8 2737 34
rect 3209 -8 3239 34
rect 3287 -8 3317 34
rect 3789 -8 3819 34
rect 3867 -8 3897 34
rect 4369 -8 4399 34
rect 4447 -8 4477 34
rect 4949 -8 4979 34
rect 5027 -8 5057 34
rect 5529 -8 5559 34
rect 5607 -8 5637 34
rect 6109 -8 6139 34
rect 6187 -8 6217 34
rect -271 -278 -241 -236
rect -193 -278 -163 -236
rect 309 -278 339 -236
rect 387 -278 417 -236
rect 889 -278 919 -236
rect 967 -278 997 -236
rect 1469 -278 1499 -236
rect 1547 -278 1577 -236
rect 2049 -278 2079 -236
rect 2127 -278 2157 -236
rect 2629 -278 2659 -236
rect 2707 -278 2737 -236
rect 3209 -278 3239 -236
rect 3287 -278 3317 -236
rect 3789 -278 3819 -236
rect 3867 -278 3897 -236
rect 4369 -278 4399 -236
rect 4447 -278 4477 -236
rect 4949 -278 4979 -236
rect 5027 -278 5057 -236
rect 5529 -278 5559 -236
rect 5607 -278 5637 -236
rect 6109 -278 6139 -236
rect 6187 -278 6217 -236
rect -271 -548 -241 -506
rect -193 -548 -163 -506
rect 309 -548 339 -506
rect 387 -548 417 -506
rect 889 -548 919 -506
rect 967 -548 997 -506
rect 1469 -548 1499 -506
rect 1547 -548 1577 -506
rect 2049 -548 2079 -506
rect 2127 -548 2157 -506
rect 2629 -548 2659 -506
rect 2707 -548 2737 -506
rect 3209 -548 3239 -506
rect 3287 -548 3317 -506
rect 3789 -548 3819 -506
rect 3867 -548 3897 -506
rect 4369 -548 4399 -506
rect 4447 -548 4477 -506
rect 4949 -548 4979 -506
rect 5027 -548 5057 -506
rect 5529 -548 5559 -506
rect 5607 -548 5637 -506
rect 6109 -548 6139 -506
rect 6187 -548 6217 -506
rect -271 -818 -241 -776
rect -193 -818 -163 -776
rect 309 -818 339 -776
rect 387 -818 417 -776
rect 889 -818 919 -776
rect 967 -818 997 -776
rect 1469 -818 1499 -776
rect 1547 -818 1577 -776
rect 2049 -818 2079 -776
rect 2127 -818 2157 -776
rect 2629 -818 2659 -776
rect 2707 -818 2737 -776
rect 3209 -818 3239 -776
rect 3287 -818 3317 -776
rect 3789 -818 3819 -776
rect 3867 -818 3897 -776
rect 4369 -818 4399 -776
rect 4447 -818 4477 -776
rect 4949 -818 4979 -776
rect 5027 -818 5057 -776
rect 5529 -818 5559 -776
rect 5607 -818 5637 -776
rect 6109 -818 6139 -776
rect 6187 -818 6217 -776
rect -271 -1088 -241 -1046
rect -193 -1088 -163 -1046
rect 309 -1088 339 -1046
rect 387 -1088 417 -1046
rect 889 -1088 919 -1046
rect 967 -1088 997 -1046
rect 1469 -1088 1499 -1046
rect 1547 -1088 1577 -1046
rect 2049 -1088 2079 -1046
rect 2127 -1088 2157 -1046
rect 2629 -1088 2659 -1046
rect 2707 -1088 2737 -1046
rect 3209 -1088 3239 -1046
rect 3287 -1088 3317 -1046
rect 3789 -1088 3819 -1046
rect 3867 -1088 3897 -1046
rect 4369 -1088 4399 -1046
rect 4447 -1088 4477 -1046
rect 4949 -1088 4979 -1046
rect 5027 -1088 5057 -1046
rect 5529 -1088 5559 -1046
rect 5607 -1088 5637 -1046
rect 6109 -1088 6139 -1046
rect 6187 -1088 6217 -1046
rect -271 -1358 -241 -1316
rect -193 -1358 -163 -1316
rect 309 -1358 339 -1316
rect 387 -1358 417 -1316
rect 889 -1358 919 -1316
rect 967 -1358 997 -1316
rect 1469 -1358 1499 -1316
rect 1547 -1358 1577 -1316
rect 2049 -1358 2079 -1316
rect 2127 -1358 2157 -1316
rect 2629 -1358 2659 -1316
rect 2707 -1358 2737 -1316
rect 3209 -1358 3239 -1316
rect 3287 -1358 3317 -1316
rect 3789 -1358 3819 -1316
rect 3867 -1358 3897 -1316
rect 4369 -1358 4399 -1316
rect 4447 -1358 4477 -1316
rect 4949 -1358 4979 -1316
rect 5027 -1358 5057 -1316
rect 5529 -1358 5559 -1316
rect 5607 -1358 5637 -1316
rect 6109 -1358 6139 -1316
rect 6187 -1358 6217 -1316
rect -271 -1628 -241 -1586
rect -193 -1628 -163 -1586
rect 309 -1628 339 -1586
rect 387 -1628 417 -1586
rect 889 -1628 919 -1586
rect 967 -1628 997 -1586
rect 1469 -1628 1499 -1586
rect 1547 -1628 1577 -1586
rect 2049 -1628 2079 -1586
rect 2127 -1628 2157 -1586
rect 2629 -1628 2659 -1586
rect 2707 -1628 2737 -1586
rect 3209 -1628 3239 -1586
rect 3287 -1628 3317 -1586
rect 3789 -1628 3819 -1586
rect 3867 -1628 3897 -1586
rect 4369 -1628 4399 -1586
rect 4447 -1628 4477 -1586
rect 4949 -1628 4979 -1586
rect 5027 -1628 5057 -1586
rect 5529 -1628 5559 -1586
rect 5607 -1628 5637 -1586
rect 6109 -1628 6139 -1586
rect 6187 -1628 6217 -1586
rect -271 -1898 -241 -1856
rect -193 -1898 -163 -1856
rect 309 -1898 339 -1856
rect 387 -1898 417 -1856
rect 889 -1898 919 -1856
rect 967 -1898 997 -1856
rect 1469 -1898 1499 -1856
rect 1547 -1898 1577 -1856
rect 2049 -1898 2079 -1856
rect 2127 -1898 2157 -1856
rect 2629 -1898 2659 -1856
rect 2707 -1898 2737 -1856
rect 3209 -1898 3239 -1856
rect 3287 -1898 3317 -1856
rect 3789 -1898 3819 -1856
rect 3867 -1898 3897 -1856
rect 4369 -1898 4399 -1856
rect 4447 -1898 4477 -1856
rect 4949 -1898 4979 -1856
rect 5027 -1898 5057 -1856
rect 5529 -1898 5559 -1856
rect 5607 -1898 5637 -1856
rect 6109 -1898 6139 -1856
rect 6187 -1898 6217 -1856
rect -271 -2168 -241 -2126
rect -193 -2168 -163 -2126
rect 309 -2168 339 -2126
rect 387 -2168 417 -2126
rect 889 -2168 919 -2126
rect 967 -2168 997 -2126
rect 1469 -2168 1499 -2126
rect 1547 -2168 1577 -2126
rect 2049 -2168 2079 -2126
rect 2127 -2168 2157 -2126
rect 2629 -2168 2659 -2126
rect 2707 -2168 2737 -2126
rect 3209 -2168 3239 -2126
rect 3287 -2168 3317 -2126
rect 3789 -2168 3819 -2126
rect 3867 -2168 3897 -2126
rect 4369 -2168 4399 -2126
rect 4447 -2168 4477 -2126
rect 4949 -2168 4979 -2126
rect 5027 -2168 5057 -2126
rect 5529 -2168 5559 -2126
rect 5607 -2168 5637 -2126
rect 6109 -2168 6139 -2126
rect 6187 -2168 6217 -2126
rect -271 -2438 -241 -2396
rect -193 -2438 -163 -2396
rect 309 -2438 339 -2396
rect 387 -2438 417 -2396
rect 889 -2438 919 -2396
rect 967 -2438 997 -2396
rect 1469 -2438 1499 -2396
rect 1547 -2438 1577 -2396
rect 2049 -2438 2079 -2396
rect 2127 -2438 2157 -2396
rect 2629 -2438 2659 -2396
rect 2707 -2438 2737 -2396
rect 3209 -2438 3239 -2396
rect 3287 -2438 3317 -2396
rect 3789 -2438 3819 -2396
rect 3867 -2438 3897 -2396
rect 4369 -2438 4399 -2396
rect 4447 -2438 4477 -2396
rect 4949 -2438 4979 -2396
rect 5027 -2438 5057 -2396
rect 5529 -2438 5559 -2396
rect 5607 -2438 5637 -2396
rect 6109 -2438 6139 -2396
rect 6187 -2438 6217 -2396
<< npass >>
rect -364 1612 -334 1640
rect -100 1612 -70 1640
rect 216 1612 246 1640
rect 480 1612 510 1640
rect 796 1612 826 1640
rect 1060 1612 1090 1640
rect 1376 1612 1406 1640
rect 1640 1612 1670 1640
rect 1956 1612 1986 1640
rect 2220 1612 2250 1640
rect 2536 1612 2566 1640
rect 2800 1612 2830 1640
rect 3116 1612 3146 1640
rect 3380 1612 3410 1640
rect 3696 1612 3726 1640
rect 3960 1612 3990 1640
rect 4276 1612 4306 1640
rect 4540 1612 4570 1640
rect 4856 1612 4886 1640
rect 5120 1612 5150 1640
rect 5436 1612 5466 1640
rect 5700 1612 5730 1640
rect 6016 1612 6046 1640
rect 6280 1612 6310 1640
rect -364 1342 -334 1370
rect -100 1342 -70 1370
rect 216 1342 246 1370
rect 480 1342 510 1370
rect 796 1342 826 1370
rect 1060 1342 1090 1370
rect 1376 1342 1406 1370
rect 1640 1342 1670 1370
rect 1956 1342 1986 1370
rect 2220 1342 2250 1370
rect 2536 1342 2566 1370
rect 2800 1342 2830 1370
rect 3116 1342 3146 1370
rect 3380 1342 3410 1370
rect 3696 1342 3726 1370
rect 3960 1342 3990 1370
rect 4276 1342 4306 1370
rect 4540 1342 4570 1370
rect 4856 1342 4886 1370
rect 5120 1342 5150 1370
rect 5436 1342 5466 1370
rect 5700 1342 5730 1370
rect 6016 1342 6046 1370
rect 6280 1342 6310 1370
rect -364 1072 -334 1100
rect -100 1072 -70 1100
rect 216 1072 246 1100
rect 480 1072 510 1100
rect 796 1072 826 1100
rect 1060 1072 1090 1100
rect 1376 1072 1406 1100
rect 1640 1072 1670 1100
rect 1956 1072 1986 1100
rect 2220 1072 2250 1100
rect 2536 1072 2566 1100
rect 2800 1072 2830 1100
rect 3116 1072 3146 1100
rect 3380 1072 3410 1100
rect 3696 1072 3726 1100
rect 3960 1072 3990 1100
rect 4276 1072 4306 1100
rect 4540 1072 4570 1100
rect 4856 1072 4886 1100
rect 5120 1072 5150 1100
rect 5436 1072 5466 1100
rect 5700 1072 5730 1100
rect 6016 1072 6046 1100
rect 6280 1072 6310 1100
rect -364 802 -334 830
rect -100 802 -70 830
rect 216 802 246 830
rect 480 802 510 830
rect 796 802 826 830
rect 1060 802 1090 830
rect 1376 802 1406 830
rect 1640 802 1670 830
rect 1956 802 1986 830
rect 2220 802 2250 830
rect 2536 802 2566 830
rect 2800 802 2830 830
rect 3116 802 3146 830
rect 3380 802 3410 830
rect 3696 802 3726 830
rect 3960 802 3990 830
rect 4276 802 4306 830
rect 4540 802 4570 830
rect 4856 802 4886 830
rect 5120 802 5150 830
rect 5436 802 5466 830
rect 5700 802 5730 830
rect 6016 802 6046 830
rect 6280 802 6310 830
rect -364 532 -334 560
rect -100 532 -70 560
rect 216 532 246 560
rect 480 532 510 560
rect 796 532 826 560
rect 1060 532 1090 560
rect 1376 532 1406 560
rect 1640 532 1670 560
rect 1956 532 1986 560
rect 2220 532 2250 560
rect 2536 532 2566 560
rect 2800 532 2830 560
rect 3116 532 3146 560
rect 3380 532 3410 560
rect 3696 532 3726 560
rect 3960 532 3990 560
rect 4276 532 4306 560
rect 4540 532 4570 560
rect 4856 532 4886 560
rect 5120 532 5150 560
rect 5436 532 5466 560
rect 5700 532 5730 560
rect 6016 532 6046 560
rect 6280 532 6310 560
rect -364 262 -334 290
rect -100 262 -70 290
rect 216 262 246 290
rect 480 262 510 290
rect 796 262 826 290
rect 1060 262 1090 290
rect 1376 262 1406 290
rect 1640 262 1670 290
rect 1956 262 1986 290
rect 2220 262 2250 290
rect 2536 262 2566 290
rect 2800 262 2830 290
rect 3116 262 3146 290
rect 3380 262 3410 290
rect 3696 262 3726 290
rect 3960 262 3990 290
rect 4276 262 4306 290
rect 4540 262 4570 290
rect 4856 262 4886 290
rect 5120 262 5150 290
rect 5436 262 5466 290
rect 5700 262 5730 290
rect 6016 262 6046 290
rect 6280 262 6310 290
rect -364 -8 -334 20
rect -100 -8 -70 20
rect 216 -8 246 20
rect 480 -8 510 20
rect 796 -8 826 20
rect 1060 -8 1090 20
rect 1376 -8 1406 20
rect 1640 -8 1670 20
rect 1956 -8 1986 20
rect 2220 -8 2250 20
rect 2536 -8 2566 20
rect 2800 -8 2830 20
rect 3116 -8 3146 20
rect 3380 -8 3410 20
rect 3696 -8 3726 20
rect 3960 -8 3990 20
rect 4276 -8 4306 20
rect 4540 -8 4570 20
rect 4856 -8 4886 20
rect 5120 -8 5150 20
rect 5436 -8 5466 20
rect 5700 -8 5730 20
rect 6016 -8 6046 20
rect 6280 -8 6310 20
rect -364 -278 -334 -250
rect -100 -278 -70 -250
rect 216 -278 246 -250
rect 480 -278 510 -250
rect 796 -278 826 -250
rect 1060 -278 1090 -250
rect 1376 -278 1406 -250
rect 1640 -278 1670 -250
rect 1956 -278 1986 -250
rect 2220 -278 2250 -250
rect 2536 -278 2566 -250
rect 2800 -278 2830 -250
rect 3116 -278 3146 -250
rect 3380 -278 3410 -250
rect 3696 -278 3726 -250
rect 3960 -278 3990 -250
rect 4276 -278 4306 -250
rect 4540 -278 4570 -250
rect 4856 -278 4886 -250
rect 5120 -278 5150 -250
rect 5436 -278 5466 -250
rect 5700 -278 5730 -250
rect 6016 -278 6046 -250
rect 6280 -278 6310 -250
rect -364 -548 -334 -520
rect -100 -548 -70 -520
rect 216 -548 246 -520
rect 480 -548 510 -520
rect 796 -548 826 -520
rect 1060 -548 1090 -520
rect 1376 -548 1406 -520
rect 1640 -548 1670 -520
rect 1956 -548 1986 -520
rect 2220 -548 2250 -520
rect 2536 -548 2566 -520
rect 2800 -548 2830 -520
rect 3116 -548 3146 -520
rect 3380 -548 3410 -520
rect 3696 -548 3726 -520
rect 3960 -548 3990 -520
rect 4276 -548 4306 -520
rect 4540 -548 4570 -520
rect 4856 -548 4886 -520
rect 5120 -548 5150 -520
rect 5436 -548 5466 -520
rect 5700 -548 5730 -520
rect 6016 -548 6046 -520
rect 6280 -548 6310 -520
rect -364 -818 -334 -790
rect -100 -818 -70 -790
rect 216 -818 246 -790
rect 480 -818 510 -790
rect 796 -818 826 -790
rect 1060 -818 1090 -790
rect 1376 -818 1406 -790
rect 1640 -818 1670 -790
rect 1956 -818 1986 -790
rect 2220 -818 2250 -790
rect 2536 -818 2566 -790
rect 2800 -818 2830 -790
rect 3116 -818 3146 -790
rect 3380 -818 3410 -790
rect 3696 -818 3726 -790
rect 3960 -818 3990 -790
rect 4276 -818 4306 -790
rect 4540 -818 4570 -790
rect 4856 -818 4886 -790
rect 5120 -818 5150 -790
rect 5436 -818 5466 -790
rect 5700 -818 5730 -790
rect 6016 -818 6046 -790
rect 6280 -818 6310 -790
rect -364 -1088 -334 -1060
rect -100 -1088 -70 -1060
rect 216 -1088 246 -1060
rect 480 -1088 510 -1060
rect 796 -1088 826 -1060
rect 1060 -1088 1090 -1060
rect 1376 -1088 1406 -1060
rect 1640 -1088 1670 -1060
rect 1956 -1088 1986 -1060
rect 2220 -1088 2250 -1060
rect 2536 -1088 2566 -1060
rect 2800 -1088 2830 -1060
rect 3116 -1088 3146 -1060
rect 3380 -1088 3410 -1060
rect 3696 -1088 3726 -1060
rect 3960 -1088 3990 -1060
rect 4276 -1088 4306 -1060
rect 4540 -1088 4570 -1060
rect 4856 -1088 4886 -1060
rect 5120 -1088 5150 -1060
rect 5436 -1088 5466 -1060
rect 5700 -1088 5730 -1060
rect 6016 -1088 6046 -1060
rect 6280 -1088 6310 -1060
rect -364 -1358 -334 -1330
rect -100 -1358 -70 -1330
rect 216 -1358 246 -1330
rect 480 -1358 510 -1330
rect 796 -1358 826 -1330
rect 1060 -1358 1090 -1330
rect 1376 -1358 1406 -1330
rect 1640 -1358 1670 -1330
rect 1956 -1358 1986 -1330
rect 2220 -1358 2250 -1330
rect 2536 -1358 2566 -1330
rect 2800 -1358 2830 -1330
rect 3116 -1358 3146 -1330
rect 3380 -1358 3410 -1330
rect 3696 -1358 3726 -1330
rect 3960 -1358 3990 -1330
rect 4276 -1358 4306 -1330
rect 4540 -1358 4570 -1330
rect 4856 -1358 4886 -1330
rect 5120 -1358 5150 -1330
rect 5436 -1358 5466 -1330
rect 5700 -1358 5730 -1330
rect 6016 -1358 6046 -1330
rect 6280 -1358 6310 -1330
rect -364 -1628 -334 -1600
rect -100 -1628 -70 -1600
rect 216 -1628 246 -1600
rect 480 -1628 510 -1600
rect 796 -1628 826 -1600
rect 1060 -1628 1090 -1600
rect 1376 -1628 1406 -1600
rect 1640 -1628 1670 -1600
rect 1956 -1628 1986 -1600
rect 2220 -1628 2250 -1600
rect 2536 -1628 2566 -1600
rect 2800 -1628 2830 -1600
rect 3116 -1628 3146 -1600
rect 3380 -1628 3410 -1600
rect 3696 -1628 3726 -1600
rect 3960 -1628 3990 -1600
rect 4276 -1628 4306 -1600
rect 4540 -1628 4570 -1600
rect 4856 -1628 4886 -1600
rect 5120 -1628 5150 -1600
rect 5436 -1628 5466 -1600
rect 5700 -1628 5730 -1600
rect 6016 -1628 6046 -1600
rect 6280 -1628 6310 -1600
rect -364 -1898 -334 -1870
rect -100 -1898 -70 -1870
rect 216 -1898 246 -1870
rect 480 -1898 510 -1870
rect 796 -1898 826 -1870
rect 1060 -1898 1090 -1870
rect 1376 -1898 1406 -1870
rect 1640 -1898 1670 -1870
rect 1956 -1898 1986 -1870
rect 2220 -1898 2250 -1870
rect 2536 -1898 2566 -1870
rect 2800 -1898 2830 -1870
rect 3116 -1898 3146 -1870
rect 3380 -1898 3410 -1870
rect 3696 -1898 3726 -1870
rect 3960 -1898 3990 -1870
rect 4276 -1898 4306 -1870
rect 4540 -1898 4570 -1870
rect 4856 -1898 4886 -1870
rect 5120 -1898 5150 -1870
rect 5436 -1898 5466 -1870
rect 5700 -1898 5730 -1870
rect 6016 -1898 6046 -1870
rect 6280 -1898 6310 -1870
rect -364 -2168 -334 -2140
rect -100 -2168 -70 -2140
rect 216 -2168 246 -2140
rect 480 -2168 510 -2140
rect 796 -2168 826 -2140
rect 1060 -2168 1090 -2140
rect 1376 -2168 1406 -2140
rect 1640 -2168 1670 -2140
rect 1956 -2168 1986 -2140
rect 2220 -2168 2250 -2140
rect 2536 -2168 2566 -2140
rect 2800 -2168 2830 -2140
rect 3116 -2168 3146 -2140
rect 3380 -2168 3410 -2140
rect 3696 -2168 3726 -2140
rect 3960 -2168 3990 -2140
rect 4276 -2168 4306 -2140
rect 4540 -2168 4570 -2140
rect 4856 -2168 4886 -2140
rect 5120 -2168 5150 -2140
rect 5436 -2168 5466 -2140
rect 5700 -2168 5730 -2140
rect 6016 -2168 6046 -2140
rect 6280 -2168 6310 -2140
rect -364 -2438 -334 -2410
rect -100 -2438 -70 -2410
rect 216 -2438 246 -2410
rect 480 -2438 510 -2410
rect 796 -2438 826 -2410
rect 1060 -2438 1090 -2410
rect 1376 -2438 1406 -2410
rect 1640 -2438 1670 -2410
rect 1956 -2438 1986 -2410
rect 2220 -2438 2250 -2410
rect 2536 -2438 2566 -2410
rect 2800 -2438 2830 -2410
rect 3116 -2438 3146 -2410
rect 3380 -2438 3410 -2410
rect 3696 -2438 3726 -2410
rect 3960 -2438 3990 -2410
rect 4276 -2438 4306 -2410
rect 4540 -2438 4570 -2410
rect 4856 -2438 4886 -2410
rect 5120 -2438 5150 -2410
rect 5436 -2438 5466 -2410
rect 5700 -2438 5730 -2410
rect 6016 -2438 6046 -2410
rect 6280 -2438 6310 -2410
<< ppu >>
rect -271 1748 -241 1776
rect -193 1748 -163 1776
rect 309 1748 339 1776
rect 387 1748 417 1776
rect 889 1748 919 1776
rect 967 1748 997 1776
rect 1469 1748 1499 1776
rect 1547 1748 1577 1776
rect 2049 1748 2079 1776
rect 2127 1748 2157 1776
rect 2629 1748 2659 1776
rect 2707 1748 2737 1776
rect 3209 1748 3239 1776
rect 3287 1748 3317 1776
rect 3789 1748 3819 1776
rect 3867 1748 3897 1776
rect 4369 1748 4399 1776
rect 4447 1748 4477 1776
rect 4949 1748 4979 1776
rect 5027 1748 5057 1776
rect 5529 1748 5559 1776
rect 5607 1748 5637 1776
rect 6109 1748 6139 1776
rect 6187 1748 6217 1776
rect -271 1478 -241 1506
rect -193 1478 -163 1506
rect 309 1478 339 1506
rect 387 1478 417 1506
rect 889 1478 919 1506
rect 967 1478 997 1506
rect 1469 1478 1499 1506
rect 1547 1478 1577 1506
rect 2049 1478 2079 1506
rect 2127 1478 2157 1506
rect 2629 1478 2659 1506
rect 2707 1478 2737 1506
rect 3209 1478 3239 1506
rect 3287 1478 3317 1506
rect 3789 1478 3819 1506
rect 3867 1478 3897 1506
rect 4369 1478 4399 1506
rect 4447 1478 4477 1506
rect 4949 1478 4979 1506
rect 5027 1478 5057 1506
rect 5529 1478 5559 1506
rect 5607 1478 5637 1506
rect 6109 1478 6139 1506
rect 6187 1478 6217 1506
rect -271 1208 -241 1236
rect -193 1208 -163 1236
rect 309 1208 339 1236
rect 387 1208 417 1236
rect 889 1208 919 1236
rect 967 1208 997 1236
rect 1469 1208 1499 1236
rect 1547 1208 1577 1236
rect 2049 1208 2079 1236
rect 2127 1208 2157 1236
rect 2629 1208 2659 1236
rect 2707 1208 2737 1236
rect 3209 1208 3239 1236
rect 3287 1208 3317 1236
rect 3789 1208 3819 1236
rect 3867 1208 3897 1236
rect 4369 1208 4399 1236
rect 4447 1208 4477 1236
rect 4949 1208 4979 1236
rect 5027 1208 5057 1236
rect 5529 1208 5559 1236
rect 5607 1208 5637 1236
rect 6109 1208 6139 1236
rect 6187 1208 6217 1236
rect -271 938 -241 966
rect -193 938 -163 966
rect 309 938 339 966
rect 387 938 417 966
rect 889 938 919 966
rect 967 938 997 966
rect 1469 938 1499 966
rect 1547 938 1577 966
rect 2049 938 2079 966
rect 2127 938 2157 966
rect 2629 938 2659 966
rect 2707 938 2737 966
rect 3209 938 3239 966
rect 3287 938 3317 966
rect 3789 938 3819 966
rect 3867 938 3897 966
rect 4369 938 4399 966
rect 4447 938 4477 966
rect 4949 938 4979 966
rect 5027 938 5057 966
rect 5529 938 5559 966
rect 5607 938 5637 966
rect 6109 938 6139 966
rect 6187 938 6217 966
rect -271 668 -241 696
rect -193 668 -163 696
rect 309 668 339 696
rect 387 668 417 696
rect 889 668 919 696
rect 967 668 997 696
rect 1469 668 1499 696
rect 1547 668 1577 696
rect 2049 668 2079 696
rect 2127 668 2157 696
rect 2629 668 2659 696
rect 2707 668 2737 696
rect 3209 668 3239 696
rect 3287 668 3317 696
rect 3789 668 3819 696
rect 3867 668 3897 696
rect 4369 668 4399 696
rect 4447 668 4477 696
rect 4949 668 4979 696
rect 5027 668 5057 696
rect 5529 668 5559 696
rect 5607 668 5637 696
rect 6109 668 6139 696
rect 6187 668 6217 696
rect -271 398 -241 426
rect -193 398 -163 426
rect 309 398 339 426
rect 387 398 417 426
rect 889 398 919 426
rect 967 398 997 426
rect 1469 398 1499 426
rect 1547 398 1577 426
rect 2049 398 2079 426
rect 2127 398 2157 426
rect 2629 398 2659 426
rect 2707 398 2737 426
rect 3209 398 3239 426
rect 3287 398 3317 426
rect 3789 398 3819 426
rect 3867 398 3897 426
rect 4369 398 4399 426
rect 4447 398 4477 426
rect 4949 398 4979 426
rect 5027 398 5057 426
rect 5529 398 5559 426
rect 5607 398 5637 426
rect 6109 398 6139 426
rect 6187 398 6217 426
rect -271 128 -241 156
rect -193 128 -163 156
rect 309 128 339 156
rect 387 128 417 156
rect 889 128 919 156
rect 967 128 997 156
rect 1469 128 1499 156
rect 1547 128 1577 156
rect 2049 128 2079 156
rect 2127 128 2157 156
rect 2629 128 2659 156
rect 2707 128 2737 156
rect 3209 128 3239 156
rect 3287 128 3317 156
rect 3789 128 3819 156
rect 3867 128 3897 156
rect 4369 128 4399 156
rect 4447 128 4477 156
rect 4949 128 4979 156
rect 5027 128 5057 156
rect 5529 128 5559 156
rect 5607 128 5637 156
rect 6109 128 6139 156
rect 6187 128 6217 156
rect -271 -142 -241 -114
rect -193 -142 -163 -114
rect 309 -142 339 -114
rect 387 -142 417 -114
rect 889 -142 919 -114
rect 967 -142 997 -114
rect 1469 -142 1499 -114
rect 1547 -142 1577 -114
rect 2049 -142 2079 -114
rect 2127 -142 2157 -114
rect 2629 -142 2659 -114
rect 2707 -142 2737 -114
rect 3209 -142 3239 -114
rect 3287 -142 3317 -114
rect 3789 -142 3819 -114
rect 3867 -142 3897 -114
rect 4369 -142 4399 -114
rect 4447 -142 4477 -114
rect 4949 -142 4979 -114
rect 5027 -142 5057 -114
rect 5529 -142 5559 -114
rect 5607 -142 5637 -114
rect 6109 -142 6139 -114
rect 6187 -142 6217 -114
rect -271 -412 -241 -384
rect -193 -412 -163 -384
rect 309 -412 339 -384
rect 387 -412 417 -384
rect 889 -412 919 -384
rect 967 -412 997 -384
rect 1469 -412 1499 -384
rect 1547 -412 1577 -384
rect 2049 -412 2079 -384
rect 2127 -412 2157 -384
rect 2629 -412 2659 -384
rect 2707 -412 2737 -384
rect 3209 -412 3239 -384
rect 3287 -412 3317 -384
rect 3789 -412 3819 -384
rect 3867 -412 3897 -384
rect 4369 -412 4399 -384
rect 4447 -412 4477 -384
rect 4949 -412 4979 -384
rect 5027 -412 5057 -384
rect 5529 -412 5559 -384
rect 5607 -412 5637 -384
rect 6109 -412 6139 -384
rect 6187 -412 6217 -384
rect -271 -682 -241 -654
rect -193 -682 -163 -654
rect 309 -682 339 -654
rect 387 -682 417 -654
rect 889 -682 919 -654
rect 967 -682 997 -654
rect 1469 -682 1499 -654
rect 1547 -682 1577 -654
rect 2049 -682 2079 -654
rect 2127 -682 2157 -654
rect 2629 -682 2659 -654
rect 2707 -682 2737 -654
rect 3209 -682 3239 -654
rect 3287 -682 3317 -654
rect 3789 -682 3819 -654
rect 3867 -682 3897 -654
rect 4369 -682 4399 -654
rect 4447 -682 4477 -654
rect 4949 -682 4979 -654
rect 5027 -682 5057 -654
rect 5529 -682 5559 -654
rect 5607 -682 5637 -654
rect 6109 -682 6139 -654
rect 6187 -682 6217 -654
rect -271 -952 -241 -924
rect -193 -952 -163 -924
rect 309 -952 339 -924
rect 387 -952 417 -924
rect 889 -952 919 -924
rect 967 -952 997 -924
rect 1469 -952 1499 -924
rect 1547 -952 1577 -924
rect 2049 -952 2079 -924
rect 2127 -952 2157 -924
rect 2629 -952 2659 -924
rect 2707 -952 2737 -924
rect 3209 -952 3239 -924
rect 3287 -952 3317 -924
rect 3789 -952 3819 -924
rect 3867 -952 3897 -924
rect 4369 -952 4399 -924
rect 4447 -952 4477 -924
rect 4949 -952 4979 -924
rect 5027 -952 5057 -924
rect 5529 -952 5559 -924
rect 5607 -952 5637 -924
rect 6109 -952 6139 -924
rect 6187 -952 6217 -924
rect -271 -1222 -241 -1194
rect -193 -1222 -163 -1194
rect 309 -1222 339 -1194
rect 387 -1222 417 -1194
rect 889 -1222 919 -1194
rect 967 -1222 997 -1194
rect 1469 -1222 1499 -1194
rect 1547 -1222 1577 -1194
rect 2049 -1222 2079 -1194
rect 2127 -1222 2157 -1194
rect 2629 -1222 2659 -1194
rect 2707 -1222 2737 -1194
rect 3209 -1222 3239 -1194
rect 3287 -1222 3317 -1194
rect 3789 -1222 3819 -1194
rect 3867 -1222 3897 -1194
rect 4369 -1222 4399 -1194
rect 4447 -1222 4477 -1194
rect 4949 -1222 4979 -1194
rect 5027 -1222 5057 -1194
rect 5529 -1222 5559 -1194
rect 5607 -1222 5637 -1194
rect 6109 -1222 6139 -1194
rect 6187 -1222 6217 -1194
rect -271 -1492 -241 -1464
rect -193 -1492 -163 -1464
rect 309 -1492 339 -1464
rect 387 -1492 417 -1464
rect 889 -1492 919 -1464
rect 967 -1492 997 -1464
rect 1469 -1492 1499 -1464
rect 1547 -1492 1577 -1464
rect 2049 -1492 2079 -1464
rect 2127 -1492 2157 -1464
rect 2629 -1492 2659 -1464
rect 2707 -1492 2737 -1464
rect 3209 -1492 3239 -1464
rect 3287 -1492 3317 -1464
rect 3789 -1492 3819 -1464
rect 3867 -1492 3897 -1464
rect 4369 -1492 4399 -1464
rect 4447 -1492 4477 -1464
rect 4949 -1492 4979 -1464
rect 5027 -1492 5057 -1464
rect 5529 -1492 5559 -1464
rect 5607 -1492 5637 -1464
rect 6109 -1492 6139 -1464
rect 6187 -1492 6217 -1464
rect -271 -1762 -241 -1734
rect -193 -1762 -163 -1734
rect 309 -1762 339 -1734
rect 387 -1762 417 -1734
rect 889 -1762 919 -1734
rect 967 -1762 997 -1734
rect 1469 -1762 1499 -1734
rect 1547 -1762 1577 -1734
rect 2049 -1762 2079 -1734
rect 2127 -1762 2157 -1734
rect 2629 -1762 2659 -1734
rect 2707 -1762 2737 -1734
rect 3209 -1762 3239 -1734
rect 3287 -1762 3317 -1734
rect 3789 -1762 3819 -1734
rect 3867 -1762 3897 -1734
rect 4369 -1762 4399 -1734
rect 4447 -1762 4477 -1734
rect 4949 -1762 4979 -1734
rect 5027 -1762 5057 -1734
rect 5529 -1762 5559 -1734
rect 5607 -1762 5637 -1734
rect 6109 -1762 6139 -1734
rect 6187 -1762 6217 -1734
rect -271 -2032 -241 -2004
rect -193 -2032 -163 -2004
rect 309 -2032 339 -2004
rect 387 -2032 417 -2004
rect 889 -2032 919 -2004
rect 967 -2032 997 -2004
rect 1469 -2032 1499 -2004
rect 1547 -2032 1577 -2004
rect 2049 -2032 2079 -2004
rect 2127 -2032 2157 -2004
rect 2629 -2032 2659 -2004
rect 2707 -2032 2737 -2004
rect 3209 -2032 3239 -2004
rect 3287 -2032 3317 -2004
rect 3789 -2032 3819 -2004
rect 3867 -2032 3897 -2004
rect 4369 -2032 4399 -2004
rect 4447 -2032 4477 -2004
rect 4949 -2032 4979 -2004
rect 5027 -2032 5057 -2004
rect 5529 -2032 5559 -2004
rect 5607 -2032 5637 -2004
rect 6109 -2032 6139 -2004
rect 6187 -2032 6217 -2004
rect -271 -2302 -241 -2274
rect -193 -2302 -163 -2274
rect 309 -2302 339 -2274
rect 387 -2302 417 -2274
rect 889 -2302 919 -2274
rect 967 -2302 997 -2274
rect 1469 -2302 1499 -2274
rect 1547 -2302 1577 -2274
rect 2049 -2302 2079 -2274
rect 2127 -2302 2157 -2274
rect 2629 -2302 2659 -2274
rect 2707 -2302 2737 -2274
rect 3209 -2302 3239 -2274
rect 3287 -2302 3317 -2274
rect 3789 -2302 3819 -2274
rect 3867 -2302 3897 -2274
rect 4369 -2302 4399 -2274
rect 4447 -2302 4477 -2274
rect 4949 -2302 4979 -2274
rect 5027 -2302 5057 -2274
rect 5529 -2302 5559 -2274
rect 5607 -2302 5637 -2274
rect 6109 -2302 6139 -2274
rect 6187 -2302 6217 -2274
<< ndiff >>
rect -404 1758 -386 1786
rect -356 1758 -338 1786
rect -96 1758 -78 1786
rect -48 1758 -29 1786
rect 176 1758 194 1786
rect 224 1758 242 1786
rect 484 1758 502 1786
rect 532 1758 551 1786
rect 756 1758 774 1786
rect 804 1758 822 1786
rect 1064 1758 1082 1786
rect 1112 1758 1131 1786
rect 1336 1758 1354 1786
rect 1384 1758 1402 1786
rect 1644 1758 1662 1786
rect 1692 1758 1711 1786
rect 1916 1758 1934 1786
rect 1964 1758 1982 1786
rect 2224 1758 2242 1786
rect 2272 1758 2291 1786
rect 2496 1758 2514 1786
rect 2544 1758 2562 1786
rect 2804 1758 2822 1786
rect 2852 1758 2871 1786
rect 3076 1758 3094 1786
rect 3124 1758 3142 1786
rect 3384 1758 3402 1786
rect 3432 1758 3451 1786
rect 3656 1758 3674 1786
rect 3704 1758 3722 1786
rect 3964 1758 3982 1786
rect 4012 1758 4031 1786
rect 4236 1758 4254 1786
rect 4284 1758 4302 1786
rect 4544 1758 4562 1786
rect 4592 1758 4611 1786
rect 4816 1758 4834 1786
rect 4864 1758 4882 1786
rect 5124 1758 5142 1786
rect 5172 1758 5191 1786
rect 5396 1758 5414 1786
rect 5444 1758 5462 1786
rect 5704 1758 5722 1786
rect 5752 1758 5771 1786
rect 5976 1758 5994 1786
rect 6024 1758 6042 1786
rect 6284 1758 6302 1786
rect 6332 1758 6351 1786
rect -478 1612 -450 1654
rect -420 1640 -395 1654
rect -296 1644 -271 1654
rect -420 1612 -364 1640
rect -334 1612 -300 1640
tri -286 1637 -279 1644 ne
rect -279 1612 -271 1644
rect -241 1612 -193 1654
rect -163 1644 -138 1654
rect -163 1612 -155 1644
rect -39 1640 -14 1654
rect -134 1612 -100 1640
rect -70 1612 -14 1640
rect 16 1612 44 1654
rect 102 1612 130 1654
rect 160 1640 185 1654
rect 284 1644 309 1654
rect 160 1612 216 1640
rect 246 1612 280 1640
tri 294 1637 301 1644 ne
rect 301 1612 309 1644
rect 339 1612 387 1654
rect 417 1644 442 1654
rect 417 1612 425 1644
rect 541 1640 566 1654
rect 446 1612 480 1640
rect 510 1612 566 1640
rect 596 1612 624 1654
rect 682 1612 710 1654
rect 740 1640 765 1654
rect 864 1644 889 1654
rect 740 1612 796 1640
rect 826 1612 860 1640
tri 874 1637 881 1644 ne
rect 881 1612 889 1644
rect 919 1612 967 1654
rect 997 1644 1022 1654
rect 997 1612 1005 1644
rect 1121 1640 1146 1654
rect 1026 1612 1060 1640
rect 1090 1612 1146 1640
rect 1176 1612 1204 1654
rect 1262 1612 1290 1654
rect 1320 1640 1345 1654
rect 1444 1644 1469 1654
rect 1320 1612 1376 1640
rect 1406 1612 1440 1640
tri 1454 1637 1461 1644 ne
rect 1461 1612 1469 1644
rect 1499 1612 1547 1654
rect 1577 1644 1602 1654
rect 1577 1612 1585 1644
rect 1701 1640 1726 1654
rect 1606 1612 1640 1640
rect 1670 1612 1726 1640
rect 1756 1612 1784 1654
rect 1842 1612 1870 1654
rect 1900 1640 1925 1654
rect 2024 1644 2049 1654
rect 1900 1612 1956 1640
rect 1986 1612 2020 1640
tri 2034 1637 2041 1644 ne
rect 2041 1612 2049 1644
rect 2079 1612 2127 1654
rect 2157 1644 2182 1654
rect 2157 1612 2165 1644
rect 2281 1640 2306 1654
rect 2186 1612 2220 1640
rect 2250 1612 2306 1640
rect 2336 1612 2364 1654
rect 2422 1612 2450 1654
rect 2480 1640 2505 1654
rect 2604 1644 2629 1654
rect 2480 1612 2536 1640
rect 2566 1612 2600 1640
tri 2614 1637 2621 1644 ne
rect 2621 1612 2629 1644
rect 2659 1612 2707 1654
rect 2737 1644 2762 1654
rect 2737 1612 2745 1644
rect 2861 1640 2886 1654
rect 2766 1612 2800 1640
rect 2830 1612 2886 1640
rect 2916 1612 2944 1654
rect 3002 1612 3030 1654
rect 3060 1640 3085 1654
rect 3184 1644 3209 1654
rect 3060 1612 3116 1640
rect 3146 1612 3180 1640
tri 3194 1637 3201 1644 ne
rect 3201 1612 3209 1644
rect 3239 1612 3287 1654
rect 3317 1644 3342 1654
rect 3317 1612 3325 1644
rect 3441 1640 3466 1654
rect 3346 1612 3380 1640
rect 3410 1612 3466 1640
rect 3496 1612 3524 1654
rect 3582 1612 3610 1654
rect 3640 1640 3665 1654
rect 3764 1644 3789 1654
rect 3640 1612 3696 1640
rect 3726 1612 3760 1640
tri 3774 1637 3781 1644 ne
rect 3781 1612 3789 1644
rect 3819 1612 3867 1654
rect 3897 1644 3922 1654
rect 3897 1612 3905 1644
rect 4021 1640 4046 1654
rect 3926 1612 3960 1640
rect 3990 1612 4046 1640
rect 4076 1612 4104 1654
rect 4162 1612 4190 1654
rect 4220 1640 4245 1654
rect 4344 1644 4369 1654
rect 4220 1612 4276 1640
rect 4306 1612 4340 1640
tri 4354 1637 4361 1644 ne
rect 4361 1612 4369 1644
rect 4399 1612 4447 1654
rect 4477 1644 4502 1654
rect 4477 1612 4485 1644
rect 4601 1640 4626 1654
rect 4506 1612 4540 1640
rect 4570 1612 4626 1640
rect 4656 1612 4684 1654
rect 4742 1612 4770 1654
rect 4800 1640 4825 1654
rect 4924 1644 4949 1654
rect 4800 1612 4856 1640
rect 4886 1612 4920 1640
tri 4934 1637 4941 1644 ne
rect 4941 1612 4949 1644
rect 4979 1612 5027 1654
rect 5057 1644 5082 1654
rect 5057 1612 5065 1644
rect 5181 1640 5206 1654
rect 5086 1612 5120 1640
rect 5150 1612 5206 1640
rect 5236 1612 5264 1654
rect 5322 1612 5350 1654
rect 5380 1640 5405 1654
rect 5504 1644 5529 1654
rect 5380 1612 5436 1640
rect 5466 1612 5500 1640
tri 5514 1637 5521 1644 ne
rect 5521 1612 5529 1644
rect 5559 1612 5607 1654
rect 5637 1644 5662 1654
rect 5637 1612 5645 1644
rect 5761 1640 5786 1654
rect 5666 1612 5700 1640
rect 5730 1612 5786 1640
rect 5816 1612 5844 1654
rect 5902 1612 5930 1654
rect 5960 1640 5985 1654
rect 6084 1644 6109 1654
rect 5960 1612 6016 1640
rect 6046 1612 6080 1640
tri 6094 1637 6101 1644 ne
rect 6101 1612 6109 1644
rect 6139 1612 6187 1654
rect 6217 1644 6242 1654
rect 6217 1612 6225 1644
rect 6341 1640 6366 1654
rect 6246 1612 6280 1640
rect 6310 1612 6366 1640
rect 6396 1612 6424 1654
rect -327 1588 -300 1612
rect -233 1590 -201 1612
rect -233 1588 -231 1590
rect -203 1588 -201 1590
rect -134 1588 -107 1612
rect -327 1574 -233 1588
rect -201 1574 -107 1588
rect 253 1588 280 1612
rect 347 1590 379 1612
rect 347 1588 349 1590
rect 377 1588 379 1590
rect 446 1588 473 1612
rect 253 1574 347 1588
rect 379 1574 473 1588
rect 833 1588 860 1612
rect 927 1590 959 1612
rect 927 1588 929 1590
rect 957 1588 959 1590
rect 1026 1588 1053 1612
rect 833 1574 927 1588
rect 959 1574 1053 1588
rect 1413 1588 1440 1612
rect 1507 1590 1539 1612
rect 1507 1588 1509 1590
rect 1537 1588 1539 1590
rect 1606 1588 1633 1612
rect 1413 1574 1507 1588
rect 1539 1574 1633 1588
rect 1993 1588 2020 1612
rect 2087 1590 2119 1612
rect 2087 1588 2089 1590
rect 2117 1588 2119 1590
rect 2186 1588 2213 1612
rect 1993 1574 2087 1588
rect 2119 1574 2213 1588
rect 2573 1588 2600 1612
rect 2667 1590 2699 1612
rect 2667 1588 2669 1590
rect 2697 1588 2699 1590
rect 2766 1588 2793 1612
rect 2573 1574 2667 1588
rect 2699 1574 2793 1588
rect 3153 1588 3180 1612
rect 3247 1590 3279 1612
rect 3247 1588 3249 1590
rect 3277 1588 3279 1590
rect 3346 1588 3373 1612
rect 3153 1574 3247 1588
rect 3279 1574 3373 1588
rect 3733 1588 3760 1612
rect 3827 1590 3859 1612
rect 3827 1588 3829 1590
rect 3857 1588 3859 1590
rect 3926 1588 3953 1612
rect 3733 1574 3827 1588
rect 3859 1574 3953 1588
rect 4313 1588 4340 1612
rect 4407 1590 4439 1612
rect 4407 1588 4409 1590
rect 4437 1588 4439 1590
rect 4506 1588 4533 1612
rect 4313 1574 4407 1588
rect 4439 1574 4533 1588
rect 4893 1588 4920 1612
rect 4987 1590 5019 1612
rect 4987 1588 4989 1590
rect 5017 1588 5019 1590
rect 5086 1588 5113 1612
rect 4893 1574 4987 1588
rect 5019 1574 5113 1588
rect 5473 1588 5500 1612
rect 5567 1590 5599 1612
rect 5567 1588 5569 1590
rect 5597 1588 5599 1590
rect 5666 1588 5693 1612
rect 5473 1574 5567 1588
rect 5599 1574 5693 1588
rect 6053 1588 6080 1612
rect 6147 1590 6179 1612
rect 6147 1588 6149 1590
rect 6177 1588 6179 1590
rect 6246 1588 6273 1612
rect 6053 1574 6147 1588
rect 6179 1574 6273 1588
rect -404 1488 -386 1516
rect -356 1488 -338 1516
rect -96 1488 -78 1516
rect -48 1488 -29 1516
rect 176 1488 194 1516
rect 224 1488 242 1516
rect 484 1488 502 1516
rect 532 1488 551 1516
rect 756 1488 774 1516
rect 804 1488 822 1516
rect 1064 1488 1082 1516
rect 1112 1488 1131 1516
rect 1336 1488 1354 1516
rect 1384 1488 1402 1516
rect 1644 1488 1662 1516
rect 1692 1488 1711 1516
rect 1916 1488 1934 1516
rect 1964 1488 1982 1516
rect 2224 1488 2242 1516
rect 2272 1488 2291 1516
rect 2496 1488 2514 1516
rect 2544 1488 2562 1516
rect 2804 1488 2822 1516
rect 2852 1488 2871 1516
rect 3076 1488 3094 1516
rect 3124 1488 3142 1516
rect 3384 1488 3402 1516
rect 3432 1488 3451 1516
rect 3656 1488 3674 1516
rect 3704 1488 3722 1516
rect 3964 1488 3982 1516
rect 4012 1488 4031 1516
rect 4236 1488 4254 1516
rect 4284 1488 4302 1516
rect 4544 1488 4562 1516
rect 4592 1488 4611 1516
rect 4816 1488 4834 1516
rect 4864 1488 4882 1516
rect 5124 1488 5142 1516
rect 5172 1488 5191 1516
rect 5396 1488 5414 1516
rect 5444 1488 5462 1516
rect 5704 1488 5722 1516
rect 5752 1488 5771 1516
rect 5976 1488 5994 1516
rect 6024 1488 6042 1516
rect 6284 1488 6302 1516
rect 6332 1488 6351 1516
rect -478 1342 -450 1384
rect -420 1370 -395 1384
rect -296 1374 -271 1384
rect -420 1342 -364 1370
rect -334 1342 -300 1370
tri -286 1367 -279 1374 ne
rect -279 1342 -271 1374
rect -241 1342 -193 1384
rect -163 1374 -138 1384
rect -163 1342 -155 1374
rect -39 1370 -14 1384
rect -134 1342 -100 1370
rect -70 1342 -14 1370
rect 16 1342 44 1384
rect 102 1342 130 1384
rect 160 1370 185 1384
rect 284 1374 309 1384
rect 160 1342 216 1370
rect 246 1342 280 1370
tri 294 1367 301 1374 ne
rect 301 1342 309 1374
rect 339 1342 387 1384
rect 417 1374 442 1384
rect 417 1342 425 1374
rect 541 1370 566 1384
rect 446 1342 480 1370
rect 510 1342 566 1370
rect 596 1342 624 1384
rect 682 1342 710 1384
rect 740 1370 765 1384
rect 864 1374 889 1384
rect 740 1342 796 1370
rect 826 1342 860 1370
tri 874 1367 881 1374 ne
rect 881 1342 889 1374
rect 919 1342 967 1384
rect 997 1374 1022 1384
rect 997 1342 1005 1374
rect 1121 1370 1146 1384
rect 1026 1342 1060 1370
rect 1090 1342 1146 1370
rect 1176 1342 1204 1384
rect 1262 1342 1290 1384
rect 1320 1370 1345 1384
rect 1444 1374 1469 1384
rect 1320 1342 1376 1370
rect 1406 1342 1440 1370
tri 1454 1367 1461 1374 ne
rect 1461 1342 1469 1374
rect 1499 1342 1547 1384
rect 1577 1374 1602 1384
rect 1577 1342 1585 1374
rect 1701 1370 1726 1384
rect 1606 1342 1640 1370
rect 1670 1342 1726 1370
rect 1756 1342 1784 1384
rect 1842 1342 1870 1384
rect 1900 1370 1925 1384
rect 2024 1374 2049 1384
rect 1900 1342 1956 1370
rect 1986 1342 2020 1370
tri 2034 1367 2041 1374 ne
rect 2041 1342 2049 1374
rect 2079 1342 2127 1384
rect 2157 1374 2182 1384
rect 2157 1342 2165 1374
rect 2281 1370 2306 1384
rect 2186 1342 2220 1370
rect 2250 1342 2306 1370
rect 2336 1342 2364 1384
rect 2422 1342 2450 1384
rect 2480 1370 2505 1384
rect 2604 1374 2629 1384
rect 2480 1342 2536 1370
rect 2566 1342 2600 1370
tri 2614 1367 2621 1374 ne
rect 2621 1342 2629 1374
rect 2659 1342 2707 1384
rect 2737 1374 2762 1384
rect 2737 1342 2745 1374
rect 2861 1370 2886 1384
rect 2766 1342 2800 1370
rect 2830 1342 2886 1370
rect 2916 1342 2944 1384
rect 3002 1342 3030 1384
rect 3060 1370 3085 1384
rect 3184 1374 3209 1384
rect 3060 1342 3116 1370
rect 3146 1342 3180 1370
tri 3194 1367 3201 1374 ne
rect 3201 1342 3209 1374
rect 3239 1342 3287 1384
rect 3317 1374 3342 1384
rect 3317 1342 3325 1374
rect 3441 1370 3466 1384
rect 3346 1342 3380 1370
rect 3410 1342 3466 1370
rect 3496 1342 3524 1384
rect 3582 1342 3610 1384
rect 3640 1370 3665 1384
rect 3764 1374 3789 1384
rect 3640 1342 3696 1370
rect 3726 1342 3760 1370
tri 3774 1367 3781 1374 ne
rect 3781 1342 3789 1374
rect 3819 1342 3867 1384
rect 3897 1374 3922 1384
rect 3897 1342 3905 1374
rect 4021 1370 4046 1384
rect 3926 1342 3960 1370
rect 3990 1342 4046 1370
rect 4076 1342 4104 1384
rect 4162 1342 4190 1384
rect 4220 1370 4245 1384
rect 4344 1374 4369 1384
rect 4220 1342 4276 1370
rect 4306 1342 4340 1370
tri 4354 1367 4361 1374 ne
rect 4361 1342 4369 1374
rect 4399 1342 4447 1384
rect 4477 1374 4502 1384
rect 4477 1342 4485 1374
rect 4601 1370 4626 1384
rect 4506 1342 4540 1370
rect 4570 1342 4626 1370
rect 4656 1342 4684 1384
rect 4742 1342 4770 1384
rect 4800 1370 4825 1384
rect 4924 1374 4949 1384
rect 4800 1342 4856 1370
rect 4886 1342 4920 1370
tri 4934 1367 4941 1374 ne
rect 4941 1342 4949 1374
rect 4979 1342 5027 1384
rect 5057 1374 5082 1384
rect 5057 1342 5065 1374
rect 5181 1370 5206 1384
rect 5086 1342 5120 1370
rect 5150 1342 5206 1370
rect 5236 1342 5264 1384
rect 5322 1342 5350 1384
rect 5380 1370 5405 1384
rect 5504 1374 5529 1384
rect 5380 1342 5436 1370
rect 5466 1342 5500 1370
tri 5514 1367 5521 1374 ne
rect 5521 1342 5529 1374
rect 5559 1342 5607 1384
rect 5637 1374 5662 1384
rect 5637 1342 5645 1374
rect 5761 1370 5786 1384
rect 5666 1342 5700 1370
rect 5730 1342 5786 1370
rect 5816 1342 5844 1384
rect 5902 1342 5930 1384
rect 5960 1370 5985 1384
rect 6084 1374 6109 1384
rect 5960 1342 6016 1370
rect 6046 1342 6080 1370
tri 6094 1367 6101 1374 ne
rect 6101 1342 6109 1374
rect 6139 1342 6187 1384
rect 6217 1374 6242 1384
rect 6217 1342 6225 1374
rect 6341 1370 6366 1384
rect 6246 1342 6280 1370
rect 6310 1342 6366 1370
rect 6396 1342 6424 1384
rect -327 1318 -300 1342
rect -233 1320 -201 1342
rect -233 1318 -231 1320
rect -203 1318 -201 1320
rect -134 1318 -107 1342
rect -327 1304 -233 1318
rect -201 1304 -107 1318
rect 253 1318 280 1342
rect 347 1320 379 1342
rect 347 1318 349 1320
rect 377 1318 379 1320
rect 446 1318 473 1342
rect 253 1304 347 1318
rect 379 1304 473 1318
rect 833 1318 860 1342
rect 927 1320 959 1342
rect 927 1318 929 1320
rect 957 1318 959 1320
rect 1026 1318 1053 1342
rect 833 1304 927 1318
rect 959 1304 1053 1318
rect 1413 1318 1440 1342
rect 1507 1320 1539 1342
rect 1507 1318 1509 1320
rect 1537 1318 1539 1320
rect 1606 1318 1633 1342
rect 1413 1304 1507 1318
rect 1539 1304 1633 1318
rect 1993 1318 2020 1342
rect 2087 1320 2119 1342
rect 2087 1318 2089 1320
rect 2117 1318 2119 1320
rect 2186 1318 2213 1342
rect 1993 1304 2087 1318
rect 2119 1304 2213 1318
rect 2573 1318 2600 1342
rect 2667 1320 2699 1342
rect 2667 1318 2669 1320
rect 2697 1318 2699 1320
rect 2766 1318 2793 1342
rect 2573 1304 2667 1318
rect 2699 1304 2793 1318
rect 3153 1318 3180 1342
rect 3247 1320 3279 1342
rect 3247 1318 3249 1320
rect 3277 1318 3279 1320
rect 3346 1318 3373 1342
rect 3153 1304 3247 1318
rect 3279 1304 3373 1318
rect 3733 1318 3760 1342
rect 3827 1320 3859 1342
rect 3827 1318 3829 1320
rect 3857 1318 3859 1320
rect 3926 1318 3953 1342
rect 3733 1304 3827 1318
rect 3859 1304 3953 1318
rect 4313 1318 4340 1342
rect 4407 1320 4439 1342
rect 4407 1318 4409 1320
rect 4437 1318 4439 1320
rect 4506 1318 4533 1342
rect 4313 1304 4407 1318
rect 4439 1304 4533 1318
rect 4893 1318 4920 1342
rect 4987 1320 5019 1342
rect 4987 1318 4989 1320
rect 5017 1318 5019 1320
rect 5086 1318 5113 1342
rect 4893 1304 4987 1318
rect 5019 1304 5113 1318
rect 5473 1318 5500 1342
rect 5567 1320 5599 1342
rect 5567 1318 5569 1320
rect 5597 1318 5599 1320
rect 5666 1318 5693 1342
rect 5473 1304 5567 1318
rect 5599 1304 5693 1318
rect 6053 1318 6080 1342
rect 6147 1320 6179 1342
rect 6147 1318 6149 1320
rect 6177 1318 6179 1320
rect 6246 1318 6273 1342
rect 6053 1304 6147 1318
rect 6179 1304 6273 1318
rect -404 1218 -386 1246
rect -356 1218 -338 1246
rect -96 1218 -78 1246
rect -48 1218 -29 1246
rect 176 1218 194 1246
rect 224 1218 242 1246
rect 484 1218 502 1246
rect 532 1218 551 1246
rect 756 1218 774 1246
rect 804 1218 822 1246
rect 1064 1218 1082 1246
rect 1112 1218 1131 1246
rect 1336 1218 1354 1246
rect 1384 1218 1402 1246
rect 1644 1218 1662 1246
rect 1692 1218 1711 1246
rect 1916 1218 1934 1246
rect 1964 1218 1982 1246
rect 2224 1218 2242 1246
rect 2272 1218 2291 1246
rect 2496 1218 2514 1246
rect 2544 1218 2562 1246
rect 2804 1218 2822 1246
rect 2852 1218 2871 1246
rect 3076 1218 3094 1246
rect 3124 1218 3142 1246
rect 3384 1218 3402 1246
rect 3432 1218 3451 1246
rect 3656 1218 3674 1246
rect 3704 1218 3722 1246
rect 3964 1218 3982 1246
rect 4012 1218 4031 1246
rect 4236 1218 4254 1246
rect 4284 1218 4302 1246
rect 4544 1218 4562 1246
rect 4592 1218 4611 1246
rect 4816 1218 4834 1246
rect 4864 1218 4882 1246
rect 5124 1218 5142 1246
rect 5172 1218 5191 1246
rect 5396 1218 5414 1246
rect 5444 1218 5462 1246
rect 5704 1218 5722 1246
rect 5752 1218 5771 1246
rect 5976 1218 5994 1246
rect 6024 1218 6042 1246
rect 6284 1218 6302 1246
rect 6332 1218 6351 1246
rect -478 1072 -450 1114
rect -420 1100 -395 1114
rect -296 1104 -271 1114
rect -420 1072 -364 1100
rect -334 1072 -300 1100
tri -286 1097 -279 1104 ne
rect -279 1072 -271 1104
rect -241 1072 -193 1114
rect -163 1104 -138 1114
rect -163 1072 -155 1104
rect -39 1100 -14 1114
rect -134 1072 -100 1100
rect -70 1072 -14 1100
rect 16 1072 44 1114
rect 102 1072 130 1114
rect 160 1100 185 1114
rect 284 1104 309 1114
rect 160 1072 216 1100
rect 246 1072 280 1100
tri 294 1097 301 1104 ne
rect 301 1072 309 1104
rect 339 1072 387 1114
rect 417 1104 442 1114
rect 417 1072 425 1104
rect 541 1100 566 1114
rect 446 1072 480 1100
rect 510 1072 566 1100
rect 596 1072 624 1114
rect 682 1072 710 1114
rect 740 1100 765 1114
rect 864 1104 889 1114
rect 740 1072 796 1100
rect 826 1072 860 1100
tri 874 1097 881 1104 ne
rect 881 1072 889 1104
rect 919 1072 967 1114
rect 997 1104 1022 1114
rect 997 1072 1005 1104
rect 1121 1100 1146 1114
rect 1026 1072 1060 1100
rect 1090 1072 1146 1100
rect 1176 1072 1204 1114
rect 1262 1072 1290 1114
rect 1320 1100 1345 1114
rect 1444 1104 1469 1114
rect 1320 1072 1376 1100
rect 1406 1072 1440 1100
tri 1454 1097 1461 1104 ne
rect 1461 1072 1469 1104
rect 1499 1072 1547 1114
rect 1577 1104 1602 1114
rect 1577 1072 1585 1104
rect 1701 1100 1726 1114
rect 1606 1072 1640 1100
rect 1670 1072 1726 1100
rect 1756 1072 1784 1114
rect 1842 1072 1870 1114
rect 1900 1100 1925 1114
rect 2024 1104 2049 1114
rect 1900 1072 1956 1100
rect 1986 1072 2020 1100
tri 2034 1097 2041 1104 ne
rect 2041 1072 2049 1104
rect 2079 1072 2127 1114
rect 2157 1104 2182 1114
rect 2157 1072 2165 1104
rect 2281 1100 2306 1114
rect 2186 1072 2220 1100
rect 2250 1072 2306 1100
rect 2336 1072 2364 1114
rect 2422 1072 2450 1114
rect 2480 1100 2505 1114
rect 2604 1104 2629 1114
rect 2480 1072 2536 1100
rect 2566 1072 2600 1100
tri 2614 1097 2621 1104 ne
rect 2621 1072 2629 1104
rect 2659 1072 2707 1114
rect 2737 1104 2762 1114
rect 2737 1072 2745 1104
rect 2861 1100 2886 1114
rect 2766 1072 2800 1100
rect 2830 1072 2886 1100
rect 2916 1072 2944 1114
rect 3002 1072 3030 1114
rect 3060 1100 3085 1114
rect 3184 1104 3209 1114
rect 3060 1072 3116 1100
rect 3146 1072 3180 1100
tri 3194 1097 3201 1104 ne
rect 3201 1072 3209 1104
rect 3239 1072 3287 1114
rect 3317 1104 3342 1114
rect 3317 1072 3325 1104
rect 3441 1100 3466 1114
rect 3346 1072 3380 1100
rect 3410 1072 3466 1100
rect 3496 1072 3524 1114
rect 3582 1072 3610 1114
rect 3640 1100 3665 1114
rect 3764 1104 3789 1114
rect 3640 1072 3696 1100
rect 3726 1072 3760 1100
tri 3774 1097 3781 1104 ne
rect 3781 1072 3789 1104
rect 3819 1072 3867 1114
rect 3897 1104 3922 1114
rect 3897 1072 3905 1104
rect 4021 1100 4046 1114
rect 3926 1072 3960 1100
rect 3990 1072 4046 1100
rect 4076 1072 4104 1114
rect 4162 1072 4190 1114
rect 4220 1100 4245 1114
rect 4344 1104 4369 1114
rect 4220 1072 4276 1100
rect 4306 1072 4340 1100
tri 4354 1097 4361 1104 ne
rect 4361 1072 4369 1104
rect 4399 1072 4447 1114
rect 4477 1104 4502 1114
rect 4477 1072 4485 1104
rect 4601 1100 4626 1114
rect 4506 1072 4540 1100
rect 4570 1072 4626 1100
rect 4656 1072 4684 1114
rect 4742 1072 4770 1114
rect 4800 1100 4825 1114
rect 4924 1104 4949 1114
rect 4800 1072 4856 1100
rect 4886 1072 4920 1100
tri 4934 1097 4941 1104 ne
rect 4941 1072 4949 1104
rect 4979 1072 5027 1114
rect 5057 1104 5082 1114
rect 5057 1072 5065 1104
rect 5181 1100 5206 1114
rect 5086 1072 5120 1100
rect 5150 1072 5206 1100
rect 5236 1072 5264 1114
rect 5322 1072 5350 1114
rect 5380 1100 5405 1114
rect 5504 1104 5529 1114
rect 5380 1072 5436 1100
rect 5466 1072 5500 1100
tri 5514 1097 5521 1104 ne
rect 5521 1072 5529 1104
rect 5559 1072 5607 1114
rect 5637 1104 5662 1114
rect 5637 1072 5645 1104
rect 5761 1100 5786 1114
rect 5666 1072 5700 1100
rect 5730 1072 5786 1100
rect 5816 1072 5844 1114
rect 5902 1072 5930 1114
rect 5960 1100 5985 1114
rect 6084 1104 6109 1114
rect 5960 1072 6016 1100
rect 6046 1072 6080 1100
tri 6094 1097 6101 1104 ne
rect 6101 1072 6109 1104
rect 6139 1072 6187 1114
rect 6217 1104 6242 1114
rect 6217 1072 6225 1104
rect 6341 1100 6366 1114
rect 6246 1072 6280 1100
rect 6310 1072 6366 1100
rect 6396 1072 6424 1114
rect -327 1048 -300 1072
rect -233 1050 -201 1072
rect -233 1048 -231 1050
rect -203 1048 -201 1050
rect -134 1048 -107 1072
rect -327 1034 -233 1048
rect -201 1034 -107 1048
rect 253 1048 280 1072
rect 347 1050 379 1072
rect 347 1048 349 1050
rect 377 1048 379 1050
rect 446 1048 473 1072
rect 253 1034 347 1048
rect 379 1034 473 1048
rect 833 1048 860 1072
rect 927 1050 959 1072
rect 927 1048 929 1050
rect 957 1048 959 1050
rect 1026 1048 1053 1072
rect 833 1034 927 1048
rect 959 1034 1053 1048
rect 1413 1048 1440 1072
rect 1507 1050 1539 1072
rect 1507 1048 1509 1050
rect 1537 1048 1539 1050
rect 1606 1048 1633 1072
rect 1413 1034 1507 1048
rect 1539 1034 1633 1048
rect 1993 1048 2020 1072
rect 2087 1050 2119 1072
rect 2087 1048 2089 1050
rect 2117 1048 2119 1050
rect 2186 1048 2213 1072
rect 1993 1034 2087 1048
rect 2119 1034 2213 1048
rect 2573 1048 2600 1072
rect 2667 1050 2699 1072
rect 2667 1048 2669 1050
rect 2697 1048 2699 1050
rect 2766 1048 2793 1072
rect 2573 1034 2667 1048
rect 2699 1034 2793 1048
rect 3153 1048 3180 1072
rect 3247 1050 3279 1072
rect 3247 1048 3249 1050
rect 3277 1048 3279 1050
rect 3346 1048 3373 1072
rect 3153 1034 3247 1048
rect 3279 1034 3373 1048
rect 3733 1048 3760 1072
rect 3827 1050 3859 1072
rect 3827 1048 3829 1050
rect 3857 1048 3859 1050
rect 3926 1048 3953 1072
rect 3733 1034 3827 1048
rect 3859 1034 3953 1048
rect 4313 1048 4340 1072
rect 4407 1050 4439 1072
rect 4407 1048 4409 1050
rect 4437 1048 4439 1050
rect 4506 1048 4533 1072
rect 4313 1034 4407 1048
rect 4439 1034 4533 1048
rect 4893 1048 4920 1072
rect 4987 1050 5019 1072
rect 4987 1048 4989 1050
rect 5017 1048 5019 1050
rect 5086 1048 5113 1072
rect 4893 1034 4987 1048
rect 5019 1034 5113 1048
rect 5473 1048 5500 1072
rect 5567 1050 5599 1072
rect 5567 1048 5569 1050
rect 5597 1048 5599 1050
rect 5666 1048 5693 1072
rect 5473 1034 5567 1048
rect 5599 1034 5693 1048
rect 6053 1048 6080 1072
rect 6147 1050 6179 1072
rect 6147 1048 6149 1050
rect 6177 1048 6179 1050
rect 6246 1048 6273 1072
rect 6053 1034 6147 1048
rect 6179 1034 6273 1048
rect -404 948 -386 976
rect -356 948 -338 976
rect -96 948 -78 976
rect -48 948 -29 976
rect 176 948 194 976
rect 224 948 242 976
rect 484 948 502 976
rect 532 948 551 976
rect 756 948 774 976
rect 804 948 822 976
rect 1064 948 1082 976
rect 1112 948 1131 976
rect 1336 948 1354 976
rect 1384 948 1402 976
rect 1644 948 1662 976
rect 1692 948 1711 976
rect 1916 948 1934 976
rect 1964 948 1982 976
rect 2224 948 2242 976
rect 2272 948 2291 976
rect 2496 948 2514 976
rect 2544 948 2562 976
rect 2804 948 2822 976
rect 2852 948 2871 976
rect 3076 948 3094 976
rect 3124 948 3142 976
rect 3384 948 3402 976
rect 3432 948 3451 976
rect 3656 948 3674 976
rect 3704 948 3722 976
rect 3964 948 3982 976
rect 4012 948 4031 976
rect 4236 948 4254 976
rect 4284 948 4302 976
rect 4544 948 4562 976
rect 4592 948 4611 976
rect 4816 948 4834 976
rect 4864 948 4882 976
rect 5124 948 5142 976
rect 5172 948 5191 976
rect 5396 948 5414 976
rect 5444 948 5462 976
rect 5704 948 5722 976
rect 5752 948 5771 976
rect 5976 948 5994 976
rect 6024 948 6042 976
rect 6284 948 6302 976
rect 6332 948 6351 976
rect -478 802 -450 844
rect -420 830 -395 844
rect -296 834 -271 844
rect -420 802 -364 830
rect -334 802 -300 830
tri -286 827 -279 834 ne
rect -279 802 -271 834
rect -241 802 -193 844
rect -163 834 -138 844
rect -163 802 -155 834
rect -39 830 -14 844
rect -134 802 -100 830
rect -70 802 -14 830
rect 16 802 44 844
rect 102 802 130 844
rect 160 830 185 844
rect 284 834 309 844
rect 160 802 216 830
rect 246 802 280 830
tri 294 827 301 834 ne
rect 301 802 309 834
rect 339 802 387 844
rect 417 834 442 844
rect 417 802 425 834
rect 541 830 566 844
rect 446 802 480 830
rect 510 802 566 830
rect 596 802 624 844
rect 682 802 710 844
rect 740 830 765 844
rect 864 834 889 844
rect 740 802 796 830
rect 826 802 860 830
tri 874 827 881 834 ne
rect 881 802 889 834
rect 919 802 967 844
rect 997 834 1022 844
rect 997 802 1005 834
rect 1121 830 1146 844
rect 1026 802 1060 830
rect 1090 802 1146 830
rect 1176 802 1204 844
rect 1262 802 1290 844
rect 1320 830 1345 844
rect 1444 834 1469 844
rect 1320 802 1376 830
rect 1406 802 1440 830
tri 1454 827 1461 834 ne
rect 1461 802 1469 834
rect 1499 802 1547 844
rect 1577 834 1602 844
rect 1577 802 1585 834
rect 1701 830 1726 844
rect 1606 802 1640 830
rect 1670 802 1726 830
rect 1756 802 1784 844
rect 1842 802 1870 844
rect 1900 830 1925 844
rect 2024 834 2049 844
rect 1900 802 1956 830
rect 1986 802 2020 830
tri 2034 827 2041 834 ne
rect 2041 802 2049 834
rect 2079 802 2127 844
rect 2157 834 2182 844
rect 2157 802 2165 834
rect 2281 830 2306 844
rect 2186 802 2220 830
rect 2250 802 2306 830
rect 2336 802 2364 844
rect 2422 802 2450 844
rect 2480 830 2505 844
rect 2604 834 2629 844
rect 2480 802 2536 830
rect 2566 802 2600 830
tri 2614 827 2621 834 ne
rect 2621 802 2629 834
rect 2659 802 2707 844
rect 2737 834 2762 844
rect 2737 802 2745 834
rect 2861 830 2886 844
rect 2766 802 2800 830
rect 2830 802 2886 830
rect 2916 802 2944 844
rect 3002 802 3030 844
rect 3060 830 3085 844
rect 3184 834 3209 844
rect 3060 802 3116 830
rect 3146 802 3180 830
tri 3194 827 3201 834 ne
rect 3201 802 3209 834
rect 3239 802 3287 844
rect 3317 834 3342 844
rect 3317 802 3325 834
rect 3441 830 3466 844
rect 3346 802 3380 830
rect 3410 802 3466 830
rect 3496 802 3524 844
rect 3582 802 3610 844
rect 3640 830 3665 844
rect 3764 834 3789 844
rect 3640 802 3696 830
rect 3726 802 3760 830
tri 3774 827 3781 834 ne
rect 3781 802 3789 834
rect 3819 802 3867 844
rect 3897 834 3922 844
rect 3897 802 3905 834
rect 4021 830 4046 844
rect 3926 802 3960 830
rect 3990 802 4046 830
rect 4076 802 4104 844
rect 4162 802 4190 844
rect 4220 830 4245 844
rect 4344 834 4369 844
rect 4220 802 4276 830
rect 4306 802 4340 830
tri 4354 827 4361 834 ne
rect 4361 802 4369 834
rect 4399 802 4447 844
rect 4477 834 4502 844
rect 4477 802 4485 834
rect 4601 830 4626 844
rect 4506 802 4540 830
rect 4570 802 4626 830
rect 4656 802 4684 844
rect 4742 802 4770 844
rect 4800 830 4825 844
rect 4924 834 4949 844
rect 4800 802 4856 830
rect 4886 802 4920 830
tri 4934 827 4941 834 ne
rect 4941 802 4949 834
rect 4979 802 5027 844
rect 5057 834 5082 844
rect 5057 802 5065 834
rect 5181 830 5206 844
rect 5086 802 5120 830
rect 5150 802 5206 830
rect 5236 802 5264 844
rect 5322 802 5350 844
rect 5380 830 5405 844
rect 5504 834 5529 844
rect 5380 802 5436 830
rect 5466 802 5500 830
tri 5514 827 5521 834 ne
rect 5521 802 5529 834
rect 5559 802 5607 844
rect 5637 834 5662 844
rect 5637 802 5645 834
rect 5761 830 5786 844
rect 5666 802 5700 830
rect 5730 802 5786 830
rect 5816 802 5844 844
rect 5902 802 5930 844
rect 5960 830 5985 844
rect 6084 834 6109 844
rect 5960 802 6016 830
rect 6046 802 6080 830
tri 6094 827 6101 834 ne
rect 6101 802 6109 834
rect 6139 802 6187 844
rect 6217 834 6242 844
rect 6217 802 6225 834
rect 6341 830 6366 844
rect 6246 802 6280 830
rect 6310 802 6366 830
rect 6396 802 6424 844
rect -327 778 -300 802
rect -233 780 -201 802
rect -233 778 -231 780
rect -203 778 -201 780
rect -134 778 -107 802
rect -327 764 -233 778
rect -201 764 -107 778
rect 253 778 280 802
rect 347 780 379 802
rect 347 778 349 780
rect 377 778 379 780
rect 446 778 473 802
rect 253 764 347 778
rect 379 764 473 778
rect 833 778 860 802
rect 927 780 959 802
rect 927 778 929 780
rect 957 778 959 780
rect 1026 778 1053 802
rect 833 764 927 778
rect 959 764 1053 778
rect 1413 778 1440 802
rect 1507 780 1539 802
rect 1507 778 1509 780
rect 1537 778 1539 780
rect 1606 778 1633 802
rect 1413 764 1507 778
rect 1539 764 1633 778
rect 1993 778 2020 802
rect 2087 780 2119 802
rect 2087 778 2089 780
rect 2117 778 2119 780
rect 2186 778 2213 802
rect 1993 764 2087 778
rect 2119 764 2213 778
rect 2573 778 2600 802
rect 2667 780 2699 802
rect 2667 778 2669 780
rect 2697 778 2699 780
rect 2766 778 2793 802
rect 2573 764 2667 778
rect 2699 764 2793 778
rect 3153 778 3180 802
rect 3247 780 3279 802
rect 3247 778 3249 780
rect 3277 778 3279 780
rect 3346 778 3373 802
rect 3153 764 3247 778
rect 3279 764 3373 778
rect 3733 778 3760 802
rect 3827 780 3859 802
rect 3827 778 3829 780
rect 3857 778 3859 780
rect 3926 778 3953 802
rect 3733 764 3827 778
rect 3859 764 3953 778
rect 4313 778 4340 802
rect 4407 780 4439 802
rect 4407 778 4409 780
rect 4437 778 4439 780
rect 4506 778 4533 802
rect 4313 764 4407 778
rect 4439 764 4533 778
rect 4893 778 4920 802
rect 4987 780 5019 802
rect 4987 778 4989 780
rect 5017 778 5019 780
rect 5086 778 5113 802
rect 4893 764 4987 778
rect 5019 764 5113 778
rect 5473 778 5500 802
rect 5567 780 5599 802
rect 5567 778 5569 780
rect 5597 778 5599 780
rect 5666 778 5693 802
rect 5473 764 5567 778
rect 5599 764 5693 778
rect 6053 778 6080 802
rect 6147 780 6179 802
rect 6147 778 6149 780
rect 6177 778 6179 780
rect 6246 778 6273 802
rect 6053 764 6147 778
rect 6179 764 6273 778
rect -404 678 -386 706
rect -356 678 -338 706
rect -96 678 -78 706
rect -48 678 -29 706
rect 176 678 194 706
rect 224 678 242 706
rect 484 678 502 706
rect 532 678 551 706
rect 756 678 774 706
rect 804 678 822 706
rect 1064 678 1082 706
rect 1112 678 1131 706
rect 1336 678 1354 706
rect 1384 678 1402 706
rect 1644 678 1662 706
rect 1692 678 1711 706
rect 1916 678 1934 706
rect 1964 678 1982 706
rect 2224 678 2242 706
rect 2272 678 2291 706
rect 2496 678 2514 706
rect 2544 678 2562 706
rect 2804 678 2822 706
rect 2852 678 2871 706
rect 3076 678 3094 706
rect 3124 678 3142 706
rect 3384 678 3402 706
rect 3432 678 3451 706
rect 3656 678 3674 706
rect 3704 678 3722 706
rect 3964 678 3982 706
rect 4012 678 4031 706
rect 4236 678 4254 706
rect 4284 678 4302 706
rect 4544 678 4562 706
rect 4592 678 4611 706
rect 4816 678 4834 706
rect 4864 678 4882 706
rect 5124 678 5142 706
rect 5172 678 5191 706
rect 5396 678 5414 706
rect 5444 678 5462 706
rect 5704 678 5722 706
rect 5752 678 5771 706
rect 5976 678 5994 706
rect 6024 678 6042 706
rect 6284 678 6302 706
rect 6332 678 6351 706
rect -478 532 -450 574
rect -420 560 -395 574
rect -296 564 -271 574
rect -420 532 -364 560
rect -334 532 -300 560
tri -286 557 -279 564 ne
rect -279 532 -271 564
rect -241 532 -193 574
rect -163 564 -138 574
rect -163 532 -155 564
rect -39 560 -14 574
rect -134 532 -100 560
rect -70 532 -14 560
rect 16 532 44 574
rect 102 532 130 574
rect 160 560 185 574
rect 284 564 309 574
rect 160 532 216 560
rect 246 532 280 560
tri 294 557 301 564 ne
rect 301 532 309 564
rect 339 532 387 574
rect 417 564 442 574
rect 417 532 425 564
rect 541 560 566 574
rect 446 532 480 560
rect 510 532 566 560
rect 596 532 624 574
rect 682 532 710 574
rect 740 560 765 574
rect 864 564 889 574
rect 740 532 796 560
rect 826 532 860 560
tri 874 557 881 564 ne
rect 881 532 889 564
rect 919 532 967 574
rect 997 564 1022 574
rect 997 532 1005 564
rect 1121 560 1146 574
rect 1026 532 1060 560
rect 1090 532 1146 560
rect 1176 532 1204 574
rect 1262 532 1290 574
rect 1320 560 1345 574
rect 1444 564 1469 574
rect 1320 532 1376 560
rect 1406 532 1440 560
tri 1454 557 1461 564 ne
rect 1461 532 1469 564
rect 1499 532 1547 574
rect 1577 564 1602 574
rect 1577 532 1585 564
rect 1701 560 1726 574
rect 1606 532 1640 560
rect 1670 532 1726 560
rect 1756 532 1784 574
rect 1842 532 1870 574
rect 1900 560 1925 574
rect 2024 564 2049 574
rect 1900 532 1956 560
rect 1986 532 2020 560
tri 2034 557 2041 564 ne
rect 2041 532 2049 564
rect 2079 532 2127 574
rect 2157 564 2182 574
rect 2157 532 2165 564
rect 2281 560 2306 574
rect 2186 532 2220 560
rect 2250 532 2306 560
rect 2336 532 2364 574
rect 2422 532 2450 574
rect 2480 560 2505 574
rect 2604 564 2629 574
rect 2480 532 2536 560
rect 2566 532 2600 560
tri 2614 557 2621 564 ne
rect 2621 532 2629 564
rect 2659 532 2707 574
rect 2737 564 2762 574
rect 2737 532 2745 564
rect 2861 560 2886 574
rect 2766 532 2800 560
rect 2830 532 2886 560
rect 2916 532 2944 574
rect 3002 532 3030 574
rect 3060 560 3085 574
rect 3184 564 3209 574
rect 3060 532 3116 560
rect 3146 532 3180 560
tri 3194 557 3201 564 ne
rect 3201 532 3209 564
rect 3239 532 3287 574
rect 3317 564 3342 574
rect 3317 532 3325 564
rect 3441 560 3466 574
rect 3346 532 3380 560
rect 3410 532 3466 560
rect 3496 532 3524 574
rect 3582 532 3610 574
rect 3640 560 3665 574
rect 3764 564 3789 574
rect 3640 532 3696 560
rect 3726 532 3760 560
tri 3774 557 3781 564 ne
rect 3781 532 3789 564
rect 3819 532 3867 574
rect 3897 564 3922 574
rect 3897 532 3905 564
rect 4021 560 4046 574
rect 3926 532 3960 560
rect 3990 532 4046 560
rect 4076 532 4104 574
rect 4162 532 4190 574
rect 4220 560 4245 574
rect 4344 564 4369 574
rect 4220 532 4276 560
rect 4306 532 4340 560
tri 4354 557 4361 564 ne
rect 4361 532 4369 564
rect 4399 532 4447 574
rect 4477 564 4502 574
rect 4477 532 4485 564
rect 4601 560 4626 574
rect 4506 532 4540 560
rect 4570 532 4626 560
rect 4656 532 4684 574
rect 4742 532 4770 574
rect 4800 560 4825 574
rect 4924 564 4949 574
rect 4800 532 4856 560
rect 4886 532 4920 560
tri 4934 557 4941 564 ne
rect 4941 532 4949 564
rect 4979 532 5027 574
rect 5057 564 5082 574
rect 5057 532 5065 564
rect 5181 560 5206 574
rect 5086 532 5120 560
rect 5150 532 5206 560
rect 5236 532 5264 574
rect 5322 532 5350 574
rect 5380 560 5405 574
rect 5504 564 5529 574
rect 5380 532 5436 560
rect 5466 532 5500 560
tri 5514 557 5521 564 ne
rect 5521 532 5529 564
rect 5559 532 5607 574
rect 5637 564 5662 574
rect 5637 532 5645 564
rect 5761 560 5786 574
rect 5666 532 5700 560
rect 5730 532 5786 560
rect 5816 532 5844 574
rect 5902 532 5930 574
rect 5960 560 5985 574
rect 6084 564 6109 574
rect 5960 532 6016 560
rect 6046 532 6080 560
tri 6094 557 6101 564 ne
rect 6101 532 6109 564
rect 6139 532 6187 574
rect 6217 564 6242 574
rect 6217 532 6225 564
rect 6341 560 6366 574
rect 6246 532 6280 560
rect 6310 532 6366 560
rect 6396 532 6424 574
rect -327 508 -300 532
rect -233 510 -201 532
rect -233 508 -231 510
rect -203 508 -201 510
rect -134 508 -107 532
rect -327 494 -233 508
rect -201 494 -107 508
rect 253 508 280 532
rect 347 510 379 532
rect 347 508 349 510
rect 377 508 379 510
rect 446 508 473 532
rect 253 494 347 508
rect 379 494 473 508
rect 833 508 860 532
rect 927 510 959 532
rect 927 508 929 510
rect 957 508 959 510
rect 1026 508 1053 532
rect 833 494 927 508
rect 959 494 1053 508
rect 1413 508 1440 532
rect 1507 510 1539 532
rect 1507 508 1509 510
rect 1537 508 1539 510
rect 1606 508 1633 532
rect 1413 494 1507 508
rect 1539 494 1633 508
rect 1993 508 2020 532
rect 2087 510 2119 532
rect 2087 508 2089 510
rect 2117 508 2119 510
rect 2186 508 2213 532
rect 1993 494 2087 508
rect 2119 494 2213 508
rect 2573 508 2600 532
rect 2667 510 2699 532
rect 2667 508 2669 510
rect 2697 508 2699 510
rect 2766 508 2793 532
rect 2573 494 2667 508
rect 2699 494 2793 508
rect 3153 508 3180 532
rect 3247 510 3279 532
rect 3247 508 3249 510
rect 3277 508 3279 510
rect 3346 508 3373 532
rect 3153 494 3247 508
rect 3279 494 3373 508
rect 3733 508 3760 532
rect 3827 510 3859 532
rect 3827 508 3829 510
rect 3857 508 3859 510
rect 3926 508 3953 532
rect 3733 494 3827 508
rect 3859 494 3953 508
rect 4313 508 4340 532
rect 4407 510 4439 532
rect 4407 508 4409 510
rect 4437 508 4439 510
rect 4506 508 4533 532
rect 4313 494 4407 508
rect 4439 494 4533 508
rect 4893 508 4920 532
rect 4987 510 5019 532
rect 4987 508 4989 510
rect 5017 508 5019 510
rect 5086 508 5113 532
rect 4893 494 4987 508
rect 5019 494 5113 508
rect 5473 508 5500 532
rect 5567 510 5599 532
rect 5567 508 5569 510
rect 5597 508 5599 510
rect 5666 508 5693 532
rect 5473 494 5567 508
rect 5599 494 5693 508
rect 6053 508 6080 532
rect 6147 510 6179 532
rect 6147 508 6149 510
rect 6177 508 6179 510
rect 6246 508 6273 532
rect 6053 494 6147 508
rect 6179 494 6273 508
rect -404 408 -386 436
rect -356 408 -338 436
rect -96 408 -78 436
rect -48 408 -29 436
rect 176 408 194 436
rect 224 408 242 436
rect 484 408 502 436
rect 532 408 551 436
rect 756 408 774 436
rect 804 408 822 436
rect 1064 408 1082 436
rect 1112 408 1131 436
rect 1336 408 1354 436
rect 1384 408 1402 436
rect 1644 408 1662 436
rect 1692 408 1711 436
rect 1916 408 1934 436
rect 1964 408 1982 436
rect 2224 408 2242 436
rect 2272 408 2291 436
rect 2496 408 2514 436
rect 2544 408 2562 436
rect 2804 408 2822 436
rect 2852 408 2871 436
rect 3076 408 3094 436
rect 3124 408 3142 436
rect 3384 408 3402 436
rect 3432 408 3451 436
rect 3656 408 3674 436
rect 3704 408 3722 436
rect 3964 408 3982 436
rect 4012 408 4031 436
rect 4236 408 4254 436
rect 4284 408 4302 436
rect 4544 408 4562 436
rect 4592 408 4611 436
rect 4816 408 4834 436
rect 4864 408 4882 436
rect 5124 408 5142 436
rect 5172 408 5191 436
rect 5396 408 5414 436
rect 5444 408 5462 436
rect 5704 408 5722 436
rect 5752 408 5771 436
rect 5976 408 5994 436
rect 6024 408 6042 436
rect 6284 408 6302 436
rect 6332 408 6351 436
rect -478 262 -450 304
rect -420 290 -395 304
rect -296 294 -271 304
rect -420 262 -364 290
rect -334 262 -300 290
tri -286 287 -279 294 ne
rect -279 262 -271 294
rect -241 262 -193 304
rect -163 294 -138 304
rect -163 262 -155 294
rect -39 290 -14 304
rect -134 262 -100 290
rect -70 262 -14 290
rect 16 262 44 304
rect 102 262 130 304
rect 160 290 185 304
rect 284 294 309 304
rect 160 262 216 290
rect 246 262 280 290
tri 294 287 301 294 ne
rect 301 262 309 294
rect 339 262 387 304
rect 417 294 442 304
rect 417 262 425 294
rect 541 290 566 304
rect 446 262 480 290
rect 510 262 566 290
rect 596 262 624 304
rect 682 262 710 304
rect 740 290 765 304
rect 864 294 889 304
rect 740 262 796 290
rect 826 262 860 290
tri 874 287 881 294 ne
rect 881 262 889 294
rect 919 262 967 304
rect 997 294 1022 304
rect 997 262 1005 294
rect 1121 290 1146 304
rect 1026 262 1060 290
rect 1090 262 1146 290
rect 1176 262 1204 304
rect 1262 262 1290 304
rect 1320 290 1345 304
rect 1444 294 1469 304
rect 1320 262 1376 290
rect 1406 262 1440 290
tri 1454 287 1461 294 ne
rect 1461 262 1469 294
rect 1499 262 1547 304
rect 1577 294 1602 304
rect 1577 262 1585 294
rect 1701 290 1726 304
rect 1606 262 1640 290
rect 1670 262 1726 290
rect 1756 262 1784 304
rect 1842 262 1870 304
rect 1900 290 1925 304
rect 2024 294 2049 304
rect 1900 262 1956 290
rect 1986 262 2020 290
tri 2034 287 2041 294 ne
rect 2041 262 2049 294
rect 2079 262 2127 304
rect 2157 294 2182 304
rect 2157 262 2165 294
rect 2281 290 2306 304
rect 2186 262 2220 290
rect 2250 262 2306 290
rect 2336 262 2364 304
rect 2422 262 2450 304
rect 2480 290 2505 304
rect 2604 294 2629 304
rect 2480 262 2536 290
rect 2566 262 2600 290
tri 2614 287 2621 294 ne
rect 2621 262 2629 294
rect 2659 262 2707 304
rect 2737 294 2762 304
rect 2737 262 2745 294
rect 2861 290 2886 304
rect 2766 262 2800 290
rect 2830 262 2886 290
rect 2916 262 2944 304
rect 3002 262 3030 304
rect 3060 290 3085 304
rect 3184 294 3209 304
rect 3060 262 3116 290
rect 3146 262 3180 290
tri 3194 287 3201 294 ne
rect 3201 262 3209 294
rect 3239 262 3287 304
rect 3317 294 3342 304
rect 3317 262 3325 294
rect 3441 290 3466 304
rect 3346 262 3380 290
rect 3410 262 3466 290
rect 3496 262 3524 304
rect 3582 262 3610 304
rect 3640 290 3665 304
rect 3764 294 3789 304
rect 3640 262 3696 290
rect 3726 262 3760 290
tri 3774 287 3781 294 ne
rect 3781 262 3789 294
rect 3819 262 3867 304
rect 3897 294 3922 304
rect 3897 262 3905 294
rect 4021 290 4046 304
rect 3926 262 3960 290
rect 3990 262 4046 290
rect 4076 262 4104 304
rect 4162 262 4190 304
rect 4220 290 4245 304
rect 4344 294 4369 304
rect 4220 262 4276 290
rect 4306 262 4340 290
tri 4354 287 4361 294 ne
rect 4361 262 4369 294
rect 4399 262 4447 304
rect 4477 294 4502 304
rect 4477 262 4485 294
rect 4601 290 4626 304
rect 4506 262 4540 290
rect 4570 262 4626 290
rect 4656 262 4684 304
rect 4742 262 4770 304
rect 4800 290 4825 304
rect 4924 294 4949 304
rect 4800 262 4856 290
rect 4886 262 4920 290
tri 4934 287 4941 294 ne
rect 4941 262 4949 294
rect 4979 262 5027 304
rect 5057 294 5082 304
rect 5057 262 5065 294
rect 5181 290 5206 304
rect 5086 262 5120 290
rect 5150 262 5206 290
rect 5236 262 5264 304
rect 5322 262 5350 304
rect 5380 290 5405 304
rect 5504 294 5529 304
rect 5380 262 5436 290
rect 5466 262 5500 290
tri 5514 287 5521 294 ne
rect 5521 262 5529 294
rect 5559 262 5607 304
rect 5637 294 5662 304
rect 5637 262 5645 294
rect 5761 290 5786 304
rect 5666 262 5700 290
rect 5730 262 5786 290
rect 5816 262 5844 304
rect 5902 262 5930 304
rect 5960 290 5985 304
rect 6084 294 6109 304
rect 5960 262 6016 290
rect 6046 262 6080 290
tri 6094 287 6101 294 ne
rect 6101 262 6109 294
rect 6139 262 6187 304
rect 6217 294 6242 304
rect 6217 262 6225 294
rect 6341 290 6366 304
rect 6246 262 6280 290
rect 6310 262 6366 290
rect 6396 262 6424 304
rect -327 238 -300 262
rect -233 240 -201 262
rect -233 238 -231 240
rect -203 238 -201 240
rect -134 238 -107 262
rect -327 224 -233 238
rect -201 224 -107 238
rect 253 238 280 262
rect 347 240 379 262
rect 347 238 349 240
rect 377 238 379 240
rect 446 238 473 262
rect 253 224 347 238
rect 379 224 473 238
rect 833 238 860 262
rect 927 240 959 262
rect 927 238 929 240
rect 957 238 959 240
rect 1026 238 1053 262
rect 833 224 927 238
rect 959 224 1053 238
rect 1413 238 1440 262
rect 1507 240 1539 262
rect 1507 238 1509 240
rect 1537 238 1539 240
rect 1606 238 1633 262
rect 1413 224 1507 238
rect 1539 224 1633 238
rect 1993 238 2020 262
rect 2087 240 2119 262
rect 2087 238 2089 240
rect 2117 238 2119 240
rect 2186 238 2213 262
rect 1993 224 2087 238
rect 2119 224 2213 238
rect 2573 238 2600 262
rect 2667 240 2699 262
rect 2667 238 2669 240
rect 2697 238 2699 240
rect 2766 238 2793 262
rect 2573 224 2667 238
rect 2699 224 2793 238
rect 3153 238 3180 262
rect 3247 240 3279 262
rect 3247 238 3249 240
rect 3277 238 3279 240
rect 3346 238 3373 262
rect 3153 224 3247 238
rect 3279 224 3373 238
rect 3733 238 3760 262
rect 3827 240 3859 262
rect 3827 238 3829 240
rect 3857 238 3859 240
rect 3926 238 3953 262
rect 3733 224 3827 238
rect 3859 224 3953 238
rect 4313 238 4340 262
rect 4407 240 4439 262
rect 4407 238 4409 240
rect 4437 238 4439 240
rect 4506 238 4533 262
rect 4313 224 4407 238
rect 4439 224 4533 238
rect 4893 238 4920 262
rect 4987 240 5019 262
rect 4987 238 4989 240
rect 5017 238 5019 240
rect 5086 238 5113 262
rect 4893 224 4987 238
rect 5019 224 5113 238
rect 5473 238 5500 262
rect 5567 240 5599 262
rect 5567 238 5569 240
rect 5597 238 5599 240
rect 5666 238 5693 262
rect 5473 224 5567 238
rect 5599 224 5693 238
rect 6053 238 6080 262
rect 6147 240 6179 262
rect 6147 238 6149 240
rect 6177 238 6179 240
rect 6246 238 6273 262
rect 6053 224 6147 238
rect 6179 224 6273 238
rect -404 138 -386 166
rect -356 138 -338 166
rect -96 138 -78 166
rect -48 138 -29 166
rect 176 138 194 166
rect 224 138 242 166
rect 484 138 502 166
rect 532 138 551 166
rect 756 138 774 166
rect 804 138 822 166
rect 1064 138 1082 166
rect 1112 138 1131 166
rect 1336 138 1354 166
rect 1384 138 1402 166
rect 1644 138 1662 166
rect 1692 138 1711 166
rect 1916 138 1934 166
rect 1964 138 1982 166
rect 2224 138 2242 166
rect 2272 138 2291 166
rect 2496 138 2514 166
rect 2544 138 2562 166
rect 2804 138 2822 166
rect 2852 138 2871 166
rect 3076 138 3094 166
rect 3124 138 3142 166
rect 3384 138 3402 166
rect 3432 138 3451 166
rect 3656 138 3674 166
rect 3704 138 3722 166
rect 3964 138 3982 166
rect 4012 138 4031 166
rect 4236 138 4254 166
rect 4284 138 4302 166
rect 4544 138 4562 166
rect 4592 138 4611 166
rect 4816 138 4834 166
rect 4864 138 4882 166
rect 5124 138 5142 166
rect 5172 138 5191 166
rect 5396 138 5414 166
rect 5444 138 5462 166
rect 5704 138 5722 166
rect 5752 138 5771 166
rect 5976 138 5994 166
rect 6024 138 6042 166
rect 6284 138 6302 166
rect 6332 138 6351 166
rect -478 -8 -450 34
rect -420 20 -395 34
rect -296 24 -271 34
rect -420 -8 -364 20
rect -334 -8 -300 20
tri -286 17 -279 24 ne
rect -279 -8 -271 24
rect -241 -8 -193 34
rect -163 24 -138 34
rect -163 -8 -155 24
rect -39 20 -14 34
rect -134 -8 -100 20
rect -70 -8 -14 20
rect 16 -8 44 34
rect 102 -8 130 34
rect 160 20 185 34
rect 284 24 309 34
rect 160 -8 216 20
rect 246 -8 280 20
tri 294 17 301 24 ne
rect 301 -8 309 24
rect 339 -8 387 34
rect 417 24 442 34
rect 417 -8 425 24
rect 541 20 566 34
rect 446 -8 480 20
rect 510 -8 566 20
rect 596 -8 624 34
rect 682 -8 710 34
rect 740 20 765 34
rect 864 24 889 34
rect 740 -8 796 20
rect 826 -8 860 20
tri 874 17 881 24 ne
rect 881 -8 889 24
rect 919 -8 967 34
rect 997 24 1022 34
rect 997 -8 1005 24
rect 1121 20 1146 34
rect 1026 -8 1060 20
rect 1090 -8 1146 20
rect 1176 -8 1204 34
rect 1262 -8 1290 34
rect 1320 20 1345 34
rect 1444 24 1469 34
rect 1320 -8 1376 20
rect 1406 -8 1440 20
tri 1454 17 1461 24 ne
rect 1461 -8 1469 24
rect 1499 -8 1547 34
rect 1577 24 1602 34
rect 1577 -8 1585 24
rect 1701 20 1726 34
rect 1606 -8 1640 20
rect 1670 -8 1726 20
rect 1756 -8 1784 34
rect 1842 -8 1870 34
rect 1900 20 1925 34
rect 2024 24 2049 34
rect 1900 -8 1956 20
rect 1986 -8 2020 20
tri 2034 17 2041 24 ne
rect 2041 -8 2049 24
rect 2079 -8 2127 34
rect 2157 24 2182 34
rect 2157 -8 2165 24
rect 2281 20 2306 34
rect 2186 -8 2220 20
rect 2250 -8 2306 20
rect 2336 -8 2364 34
rect 2422 -8 2450 34
rect 2480 20 2505 34
rect 2604 24 2629 34
rect 2480 -8 2536 20
rect 2566 -8 2600 20
tri 2614 17 2621 24 ne
rect 2621 -8 2629 24
rect 2659 -8 2707 34
rect 2737 24 2762 34
rect 2737 -8 2745 24
rect 2861 20 2886 34
rect 2766 -8 2800 20
rect 2830 -8 2886 20
rect 2916 -8 2944 34
rect 3002 -8 3030 34
rect 3060 20 3085 34
rect 3184 24 3209 34
rect 3060 -8 3116 20
rect 3146 -8 3180 20
tri 3194 17 3201 24 ne
rect 3201 -8 3209 24
rect 3239 -8 3287 34
rect 3317 24 3342 34
rect 3317 -8 3325 24
rect 3441 20 3466 34
rect 3346 -8 3380 20
rect 3410 -8 3466 20
rect 3496 -8 3524 34
rect 3582 -8 3610 34
rect 3640 20 3665 34
rect 3764 24 3789 34
rect 3640 -8 3696 20
rect 3726 -8 3760 20
tri 3774 17 3781 24 ne
rect 3781 -8 3789 24
rect 3819 -8 3867 34
rect 3897 24 3922 34
rect 3897 -8 3905 24
rect 4021 20 4046 34
rect 3926 -8 3960 20
rect 3990 -8 4046 20
rect 4076 -8 4104 34
rect 4162 -8 4190 34
rect 4220 20 4245 34
rect 4344 24 4369 34
rect 4220 -8 4276 20
rect 4306 -8 4340 20
tri 4354 17 4361 24 ne
rect 4361 -8 4369 24
rect 4399 -8 4447 34
rect 4477 24 4502 34
rect 4477 -8 4485 24
rect 4601 20 4626 34
rect 4506 -8 4540 20
rect 4570 -8 4626 20
rect 4656 -8 4684 34
rect 4742 -8 4770 34
rect 4800 20 4825 34
rect 4924 24 4949 34
rect 4800 -8 4856 20
rect 4886 -8 4920 20
tri 4934 17 4941 24 ne
rect 4941 -8 4949 24
rect 4979 -8 5027 34
rect 5057 24 5082 34
rect 5057 -8 5065 24
rect 5181 20 5206 34
rect 5086 -8 5120 20
rect 5150 -8 5206 20
rect 5236 -8 5264 34
rect 5322 -8 5350 34
rect 5380 20 5405 34
rect 5504 24 5529 34
rect 5380 -8 5436 20
rect 5466 -8 5500 20
tri 5514 17 5521 24 ne
rect 5521 -8 5529 24
rect 5559 -8 5607 34
rect 5637 24 5662 34
rect 5637 -8 5645 24
rect 5761 20 5786 34
rect 5666 -8 5700 20
rect 5730 -8 5786 20
rect 5816 -8 5844 34
rect 5902 -8 5930 34
rect 5960 20 5985 34
rect 6084 24 6109 34
rect 5960 -8 6016 20
rect 6046 -8 6080 20
tri 6094 17 6101 24 ne
rect 6101 -8 6109 24
rect 6139 -8 6187 34
rect 6217 24 6242 34
rect 6217 -8 6225 24
rect 6341 20 6366 34
rect 6246 -8 6280 20
rect 6310 -8 6366 20
rect 6396 -8 6424 34
rect -327 -32 -300 -8
rect -233 -30 -201 -8
rect -233 -32 -231 -30
rect -203 -32 -201 -30
rect -134 -32 -107 -8
rect -327 -46 -233 -32
rect -201 -46 -107 -32
rect 253 -32 280 -8
rect 347 -30 379 -8
rect 347 -32 349 -30
rect 377 -32 379 -30
rect 446 -32 473 -8
rect 253 -46 347 -32
rect 379 -46 473 -32
rect 833 -32 860 -8
rect 927 -30 959 -8
rect 927 -32 929 -30
rect 957 -32 959 -30
rect 1026 -32 1053 -8
rect 833 -46 927 -32
rect 959 -46 1053 -32
rect 1413 -32 1440 -8
rect 1507 -30 1539 -8
rect 1507 -32 1509 -30
rect 1537 -32 1539 -30
rect 1606 -32 1633 -8
rect 1413 -46 1507 -32
rect 1539 -46 1633 -32
rect 1993 -32 2020 -8
rect 2087 -30 2119 -8
rect 2087 -32 2089 -30
rect 2117 -32 2119 -30
rect 2186 -32 2213 -8
rect 1993 -46 2087 -32
rect 2119 -46 2213 -32
rect 2573 -32 2600 -8
rect 2667 -30 2699 -8
rect 2667 -32 2669 -30
rect 2697 -32 2699 -30
rect 2766 -32 2793 -8
rect 2573 -46 2667 -32
rect 2699 -46 2793 -32
rect 3153 -32 3180 -8
rect 3247 -30 3279 -8
rect 3247 -32 3249 -30
rect 3277 -32 3279 -30
rect 3346 -32 3373 -8
rect 3153 -46 3247 -32
rect 3279 -46 3373 -32
rect 3733 -32 3760 -8
rect 3827 -30 3859 -8
rect 3827 -32 3829 -30
rect 3857 -32 3859 -30
rect 3926 -32 3953 -8
rect 3733 -46 3827 -32
rect 3859 -46 3953 -32
rect 4313 -32 4340 -8
rect 4407 -30 4439 -8
rect 4407 -32 4409 -30
rect 4437 -32 4439 -30
rect 4506 -32 4533 -8
rect 4313 -46 4407 -32
rect 4439 -46 4533 -32
rect 4893 -32 4920 -8
rect 4987 -30 5019 -8
rect 4987 -32 4989 -30
rect 5017 -32 5019 -30
rect 5086 -32 5113 -8
rect 4893 -46 4987 -32
rect 5019 -46 5113 -32
rect 5473 -32 5500 -8
rect 5567 -30 5599 -8
rect 5567 -32 5569 -30
rect 5597 -32 5599 -30
rect 5666 -32 5693 -8
rect 5473 -46 5567 -32
rect 5599 -46 5693 -32
rect 6053 -32 6080 -8
rect 6147 -30 6179 -8
rect 6147 -32 6149 -30
rect 6177 -32 6179 -30
rect 6246 -32 6273 -8
rect 6053 -46 6147 -32
rect 6179 -46 6273 -32
rect -404 -132 -386 -104
rect -356 -132 -338 -104
rect -96 -132 -78 -104
rect -48 -132 -29 -104
rect 176 -132 194 -104
rect 224 -132 242 -104
rect 484 -132 502 -104
rect 532 -132 551 -104
rect 756 -132 774 -104
rect 804 -132 822 -104
rect 1064 -132 1082 -104
rect 1112 -132 1131 -104
rect 1336 -132 1354 -104
rect 1384 -132 1402 -104
rect 1644 -132 1662 -104
rect 1692 -132 1711 -104
rect 1916 -132 1934 -104
rect 1964 -132 1982 -104
rect 2224 -132 2242 -104
rect 2272 -132 2291 -104
rect 2496 -132 2514 -104
rect 2544 -132 2562 -104
rect 2804 -132 2822 -104
rect 2852 -132 2871 -104
rect 3076 -132 3094 -104
rect 3124 -132 3142 -104
rect 3384 -132 3402 -104
rect 3432 -132 3451 -104
rect 3656 -132 3674 -104
rect 3704 -132 3722 -104
rect 3964 -132 3982 -104
rect 4012 -132 4031 -104
rect 4236 -132 4254 -104
rect 4284 -132 4302 -104
rect 4544 -132 4562 -104
rect 4592 -132 4611 -104
rect 4816 -132 4834 -104
rect 4864 -132 4882 -104
rect 5124 -132 5142 -104
rect 5172 -132 5191 -104
rect 5396 -132 5414 -104
rect 5444 -132 5462 -104
rect 5704 -132 5722 -104
rect 5752 -132 5771 -104
rect 5976 -132 5994 -104
rect 6024 -132 6042 -104
rect 6284 -132 6302 -104
rect 6332 -132 6351 -104
rect -478 -278 -450 -236
rect -420 -250 -395 -236
rect -296 -246 -271 -236
rect -420 -278 -364 -250
rect -334 -278 -300 -250
tri -286 -253 -279 -246 ne
rect -279 -278 -271 -246
rect -241 -278 -193 -236
rect -163 -246 -138 -236
rect -163 -278 -155 -246
rect -39 -250 -14 -236
rect -134 -278 -100 -250
rect -70 -278 -14 -250
rect 16 -278 44 -236
rect 102 -278 130 -236
rect 160 -250 185 -236
rect 284 -246 309 -236
rect 160 -278 216 -250
rect 246 -278 280 -250
tri 294 -253 301 -246 ne
rect 301 -278 309 -246
rect 339 -278 387 -236
rect 417 -246 442 -236
rect 417 -278 425 -246
rect 541 -250 566 -236
rect 446 -278 480 -250
rect 510 -278 566 -250
rect 596 -278 624 -236
rect 682 -278 710 -236
rect 740 -250 765 -236
rect 864 -246 889 -236
rect 740 -278 796 -250
rect 826 -278 860 -250
tri 874 -253 881 -246 ne
rect 881 -278 889 -246
rect 919 -278 967 -236
rect 997 -246 1022 -236
rect 997 -278 1005 -246
rect 1121 -250 1146 -236
rect 1026 -278 1060 -250
rect 1090 -278 1146 -250
rect 1176 -278 1204 -236
rect 1262 -278 1290 -236
rect 1320 -250 1345 -236
rect 1444 -246 1469 -236
rect 1320 -278 1376 -250
rect 1406 -278 1440 -250
tri 1454 -253 1461 -246 ne
rect 1461 -278 1469 -246
rect 1499 -278 1547 -236
rect 1577 -246 1602 -236
rect 1577 -278 1585 -246
rect 1701 -250 1726 -236
rect 1606 -278 1640 -250
rect 1670 -278 1726 -250
rect 1756 -278 1784 -236
rect 1842 -278 1870 -236
rect 1900 -250 1925 -236
rect 2024 -246 2049 -236
rect 1900 -278 1956 -250
rect 1986 -278 2020 -250
tri 2034 -253 2041 -246 ne
rect 2041 -278 2049 -246
rect 2079 -278 2127 -236
rect 2157 -246 2182 -236
rect 2157 -278 2165 -246
rect 2281 -250 2306 -236
rect 2186 -278 2220 -250
rect 2250 -278 2306 -250
rect 2336 -278 2364 -236
rect 2422 -278 2450 -236
rect 2480 -250 2505 -236
rect 2604 -246 2629 -236
rect 2480 -278 2536 -250
rect 2566 -278 2600 -250
tri 2614 -253 2621 -246 ne
rect 2621 -278 2629 -246
rect 2659 -278 2707 -236
rect 2737 -246 2762 -236
rect 2737 -278 2745 -246
rect 2861 -250 2886 -236
rect 2766 -278 2800 -250
rect 2830 -278 2886 -250
rect 2916 -278 2944 -236
rect 3002 -278 3030 -236
rect 3060 -250 3085 -236
rect 3184 -246 3209 -236
rect 3060 -278 3116 -250
rect 3146 -278 3180 -250
tri 3194 -253 3201 -246 ne
rect 3201 -278 3209 -246
rect 3239 -278 3287 -236
rect 3317 -246 3342 -236
rect 3317 -278 3325 -246
rect 3441 -250 3466 -236
rect 3346 -278 3380 -250
rect 3410 -278 3466 -250
rect 3496 -278 3524 -236
rect 3582 -278 3610 -236
rect 3640 -250 3665 -236
rect 3764 -246 3789 -236
rect 3640 -278 3696 -250
rect 3726 -278 3760 -250
tri 3774 -253 3781 -246 ne
rect 3781 -278 3789 -246
rect 3819 -278 3867 -236
rect 3897 -246 3922 -236
rect 3897 -278 3905 -246
rect 4021 -250 4046 -236
rect 3926 -278 3960 -250
rect 3990 -278 4046 -250
rect 4076 -278 4104 -236
rect 4162 -278 4190 -236
rect 4220 -250 4245 -236
rect 4344 -246 4369 -236
rect 4220 -278 4276 -250
rect 4306 -278 4340 -250
tri 4354 -253 4361 -246 ne
rect 4361 -278 4369 -246
rect 4399 -278 4447 -236
rect 4477 -246 4502 -236
rect 4477 -278 4485 -246
rect 4601 -250 4626 -236
rect 4506 -278 4540 -250
rect 4570 -278 4626 -250
rect 4656 -278 4684 -236
rect 4742 -278 4770 -236
rect 4800 -250 4825 -236
rect 4924 -246 4949 -236
rect 4800 -278 4856 -250
rect 4886 -278 4920 -250
tri 4934 -253 4941 -246 ne
rect 4941 -278 4949 -246
rect 4979 -278 5027 -236
rect 5057 -246 5082 -236
rect 5057 -278 5065 -246
rect 5181 -250 5206 -236
rect 5086 -278 5120 -250
rect 5150 -278 5206 -250
rect 5236 -278 5264 -236
rect 5322 -278 5350 -236
rect 5380 -250 5405 -236
rect 5504 -246 5529 -236
rect 5380 -278 5436 -250
rect 5466 -278 5500 -250
tri 5514 -253 5521 -246 ne
rect 5521 -278 5529 -246
rect 5559 -278 5607 -236
rect 5637 -246 5662 -236
rect 5637 -278 5645 -246
rect 5761 -250 5786 -236
rect 5666 -278 5700 -250
rect 5730 -278 5786 -250
rect 5816 -278 5844 -236
rect 5902 -278 5930 -236
rect 5960 -250 5985 -236
rect 6084 -246 6109 -236
rect 5960 -278 6016 -250
rect 6046 -278 6080 -250
tri 6094 -253 6101 -246 ne
rect 6101 -278 6109 -246
rect 6139 -278 6187 -236
rect 6217 -246 6242 -236
rect 6217 -278 6225 -246
rect 6341 -250 6366 -236
rect 6246 -278 6280 -250
rect 6310 -278 6366 -250
rect 6396 -278 6424 -236
rect -327 -302 -300 -278
rect -233 -300 -201 -278
rect -233 -302 -231 -300
rect -203 -302 -201 -300
rect -134 -302 -107 -278
rect -327 -316 -233 -302
rect -201 -316 -107 -302
rect 253 -302 280 -278
rect 347 -300 379 -278
rect 347 -302 349 -300
rect 377 -302 379 -300
rect 446 -302 473 -278
rect 253 -316 347 -302
rect 379 -316 473 -302
rect 833 -302 860 -278
rect 927 -300 959 -278
rect 927 -302 929 -300
rect 957 -302 959 -300
rect 1026 -302 1053 -278
rect 833 -316 927 -302
rect 959 -316 1053 -302
rect 1413 -302 1440 -278
rect 1507 -300 1539 -278
rect 1507 -302 1509 -300
rect 1537 -302 1539 -300
rect 1606 -302 1633 -278
rect 1413 -316 1507 -302
rect 1539 -316 1633 -302
rect 1993 -302 2020 -278
rect 2087 -300 2119 -278
rect 2087 -302 2089 -300
rect 2117 -302 2119 -300
rect 2186 -302 2213 -278
rect 1993 -316 2087 -302
rect 2119 -316 2213 -302
rect 2573 -302 2600 -278
rect 2667 -300 2699 -278
rect 2667 -302 2669 -300
rect 2697 -302 2699 -300
rect 2766 -302 2793 -278
rect 2573 -316 2667 -302
rect 2699 -316 2793 -302
rect 3153 -302 3180 -278
rect 3247 -300 3279 -278
rect 3247 -302 3249 -300
rect 3277 -302 3279 -300
rect 3346 -302 3373 -278
rect 3153 -316 3247 -302
rect 3279 -316 3373 -302
rect 3733 -302 3760 -278
rect 3827 -300 3859 -278
rect 3827 -302 3829 -300
rect 3857 -302 3859 -300
rect 3926 -302 3953 -278
rect 3733 -316 3827 -302
rect 3859 -316 3953 -302
rect 4313 -302 4340 -278
rect 4407 -300 4439 -278
rect 4407 -302 4409 -300
rect 4437 -302 4439 -300
rect 4506 -302 4533 -278
rect 4313 -316 4407 -302
rect 4439 -316 4533 -302
rect 4893 -302 4920 -278
rect 4987 -300 5019 -278
rect 4987 -302 4989 -300
rect 5017 -302 5019 -300
rect 5086 -302 5113 -278
rect 4893 -316 4987 -302
rect 5019 -316 5113 -302
rect 5473 -302 5500 -278
rect 5567 -300 5599 -278
rect 5567 -302 5569 -300
rect 5597 -302 5599 -300
rect 5666 -302 5693 -278
rect 5473 -316 5567 -302
rect 5599 -316 5693 -302
rect 6053 -302 6080 -278
rect 6147 -300 6179 -278
rect 6147 -302 6149 -300
rect 6177 -302 6179 -300
rect 6246 -302 6273 -278
rect 6053 -316 6147 -302
rect 6179 -316 6273 -302
rect -404 -402 -386 -374
rect -356 -402 -338 -374
rect -96 -402 -78 -374
rect -48 -402 -29 -374
rect 176 -402 194 -374
rect 224 -402 242 -374
rect 484 -402 502 -374
rect 532 -402 551 -374
rect 756 -402 774 -374
rect 804 -402 822 -374
rect 1064 -402 1082 -374
rect 1112 -402 1131 -374
rect 1336 -402 1354 -374
rect 1384 -402 1402 -374
rect 1644 -402 1662 -374
rect 1692 -402 1711 -374
rect 1916 -402 1934 -374
rect 1964 -402 1982 -374
rect 2224 -402 2242 -374
rect 2272 -402 2291 -374
rect 2496 -402 2514 -374
rect 2544 -402 2562 -374
rect 2804 -402 2822 -374
rect 2852 -402 2871 -374
rect 3076 -402 3094 -374
rect 3124 -402 3142 -374
rect 3384 -402 3402 -374
rect 3432 -402 3451 -374
rect 3656 -402 3674 -374
rect 3704 -402 3722 -374
rect 3964 -402 3982 -374
rect 4012 -402 4031 -374
rect 4236 -402 4254 -374
rect 4284 -402 4302 -374
rect 4544 -402 4562 -374
rect 4592 -402 4611 -374
rect 4816 -402 4834 -374
rect 4864 -402 4882 -374
rect 5124 -402 5142 -374
rect 5172 -402 5191 -374
rect 5396 -402 5414 -374
rect 5444 -402 5462 -374
rect 5704 -402 5722 -374
rect 5752 -402 5771 -374
rect 5976 -402 5994 -374
rect 6024 -402 6042 -374
rect 6284 -402 6302 -374
rect 6332 -402 6351 -374
rect -478 -548 -450 -506
rect -420 -520 -395 -506
rect -296 -516 -271 -506
rect -420 -548 -364 -520
rect -334 -548 -300 -520
tri -286 -523 -279 -516 ne
rect -279 -548 -271 -516
rect -241 -548 -193 -506
rect -163 -516 -138 -506
rect -163 -548 -155 -516
rect -39 -520 -14 -506
rect -134 -548 -100 -520
rect -70 -548 -14 -520
rect 16 -548 44 -506
rect 102 -548 130 -506
rect 160 -520 185 -506
rect 284 -516 309 -506
rect 160 -548 216 -520
rect 246 -548 280 -520
tri 294 -523 301 -516 ne
rect 301 -548 309 -516
rect 339 -548 387 -506
rect 417 -516 442 -506
rect 417 -548 425 -516
rect 541 -520 566 -506
rect 446 -548 480 -520
rect 510 -548 566 -520
rect 596 -548 624 -506
rect 682 -548 710 -506
rect 740 -520 765 -506
rect 864 -516 889 -506
rect 740 -548 796 -520
rect 826 -548 860 -520
tri 874 -523 881 -516 ne
rect 881 -548 889 -516
rect 919 -548 967 -506
rect 997 -516 1022 -506
rect 997 -548 1005 -516
rect 1121 -520 1146 -506
rect 1026 -548 1060 -520
rect 1090 -548 1146 -520
rect 1176 -548 1204 -506
rect 1262 -548 1290 -506
rect 1320 -520 1345 -506
rect 1444 -516 1469 -506
rect 1320 -548 1376 -520
rect 1406 -548 1440 -520
tri 1454 -523 1461 -516 ne
rect 1461 -548 1469 -516
rect 1499 -548 1547 -506
rect 1577 -516 1602 -506
rect 1577 -548 1585 -516
rect 1701 -520 1726 -506
rect 1606 -548 1640 -520
rect 1670 -548 1726 -520
rect 1756 -548 1784 -506
rect 1842 -548 1870 -506
rect 1900 -520 1925 -506
rect 2024 -516 2049 -506
rect 1900 -548 1956 -520
rect 1986 -548 2020 -520
tri 2034 -523 2041 -516 ne
rect 2041 -548 2049 -516
rect 2079 -548 2127 -506
rect 2157 -516 2182 -506
rect 2157 -548 2165 -516
rect 2281 -520 2306 -506
rect 2186 -548 2220 -520
rect 2250 -548 2306 -520
rect 2336 -548 2364 -506
rect 2422 -548 2450 -506
rect 2480 -520 2505 -506
rect 2604 -516 2629 -506
rect 2480 -548 2536 -520
rect 2566 -548 2600 -520
tri 2614 -523 2621 -516 ne
rect 2621 -548 2629 -516
rect 2659 -548 2707 -506
rect 2737 -516 2762 -506
rect 2737 -548 2745 -516
rect 2861 -520 2886 -506
rect 2766 -548 2800 -520
rect 2830 -548 2886 -520
rect 2916 -548 2944 -506
rect 3002 -548 3030 -506
rect 3060 -520 3085 -506
rect 3184 -516 3209 -506
rect 3060 -548 3116 -520
rect 3146 -548 3180 -520
tri 3194 -523 3201 -516 ne
rect 3201 -548 3209 -516
rect 3239 -548 3287 -506
rect 3317 -516 3342 -506
rect 3317 -548 3325 -516
rect 3441 -520 3466 -506
rect 3346 -548 3380 -520
rect 3410 -548 3466 -520
rect 3496 -548 3524 -506
rect 3582 -548 3610 -506
rect 3640 -520 3665 -506
rect 3764 -516 3789 -506
rect 3640 -548 3696 -520
rect 3726 -548 3760 -520
tri 3774 -523 3781 -516 ne
rect 3781 -548 3789 -516
rect 3819 -548 3867 -506
rect 3897 -516 3922 -506
rect 3897 -548 3905 -516
rect 4021 -520 4046 -506
rect 3926 -548 3960 -520
rect 3990 -548 4046 -520
rect 4076 -548 4104 -506
rect 4162 -548 4190 -506
rect 4220 -520 4245 -506
rect 4344 -516 4369 -506
rect 4220 -548 4276 -520
rect 4306 -548 4340 -520
tri 4354 -523 4361 -516 ne
rect 4361 -548 4369 -516
rect 4399 -548 4447 -506
rect 4477 -516 4502 -506
rect 4477 -548 4485 -516
rect 4601 -520 4626 -506
rect 4506 -548 4540 -520
rect 4570 -548 4626 -520
rect 4656 -548 4684 -506
rect 4742 -548 4770 -506
rect 4800 -520 4825 -506
rect 4924 -516 4949 -506
rect 4800 -548 4856 -520
rect 4886 -548 4920 -520
tri 4934 -523 4941 -516 ne
rect 4941 -548 4949 -516
rect 4979 -548 5027 -506
rect 5057 -516 5082 -506
rect 5057 -548 5065 -516
rect 5181 -520 5206 -506
rect 5086 -548 5120 -520
rect 5150 -548 5206 -520
rect 5236 -548 5264 -506
rect 5322 -548 5350 -506
rect 5380 -520 5405 -506
rect 5504 -516 5529 -506
rect 5380 -548 5436 -520
rect 5466 -548 5500 -520
tri 5514 -523 5521 -516 ne
rect 5521 -548 5529 -516
rect 5559 -548 5607 -506
rect 5637 -516 5662 -506
rect 5637 -548 5645 -516
rect 5761 -520 5786 -506
rect 5666 -548 5700 -520
rect 5730 -548 5786 -520
rect 5816 -548 5844 -506
rect 5902 -548 5930 -506
rect 5960 -520 5985 -506
rect 6084 -516 6109 -506
rect 5960 -548 6016 -520
rect 6046 -548 6080 -520
tri 6094 -523 6101 -516 ne
rect 6101 -548 6109 -516
rect 6139 -548 6187 -506
rect 6217 -516 6242 -506
rect 6217 -548 6225 -516
rect 6341 -520 6366 -506
rect 6246 -548 6280 -520
rect 6310 -548 6366 -520
rect 6396 -548 6424 -506
rect -327 -572 -300 -548
rect -233 -570 -201 -548
rect -233 -572 -231 -570
rect -203 -572 -201 -570
rect -134 -572 -107 -548
rect -327 -586 -233 -572
rect -201 -586 -107 -572
rect 253 -572 280 -548
rect 347 -570 379 -548
rect 347 -572 349 -570
rect 377 -572 379 -570
rect 446 -572 473 -548
rect 253 -586 347 -572
rect 379 -586 473 -572
rect 833 -572 860 -548
rect 927 -570 959 -548
rect 927 -572 929 -570
rect 957 -572 959 -570
rect 1026 -572 1053 -548
rect 833 -586 927 -572
rect 959 -586 1053 -572
rect 1413 -572 1440 -548
rect 1507 -570 1539 -548
rect 1507 -572 1509 -570
rect 1537 -572 1539 -570
rect 1606 -572 1633 -548
rect 1413 -586 1507 -572
rect 1539 -586 1633 -572
rect 1993 -572 2020 -548
rect 2087 -570 2119 -548
rect 2087 -572 2089 -570
rect 2117 -572 2119 -570
rect 2186 -572 2213 -548
rect 1993 -586 2087 -572
rect 2119 -586 2213 -572
rect 2573 -572 2600 -548
rect 2667 -570 2699 -548
rect 2667 -572 2669 -570
rect 2697 -572 2699 -570
rect 2766 -572 2793 -548
rect 2573 -586 2667 -572
rect 2699 -586 2793 -572
rect 3153 -572 3180 -548
rect 3247 -570 3279 -548
rect 3247 -572 3249 -570
rect 3277 -572 3279 -570
rect 3346 -572 3373 -548
rect 3153 -586 3247 -572
rect 3279 -586 3373 -572
rect 3733 -572 3760 -548
rect 3827 -570 3859 -548
rect 3827 -572 3829 -570
rect 3857 -572 3859 -570
rect 3926 -572 3953 -548
rect 3733 -586 3827 -572
rect 3859 -586 3953 -572
rect 4313 -572 4340 -548
rect 4407 -570 4439 -548
rect 4407 -572 4409 -570
rect 4437 -572 4439 -570
rect 4506 -572 4533 -548
rect 4313 -586 4407 -572
rect 4439 -586 4533 -572
rect 4893 -572 4920 -548
rect 4987 -570 5019 -548
rect 4987 -572 4989 -570
rect 5017 -572 5019 -570
rect 5086 -572 5113 -548
rect 4893 -586 4987 -572
rect 5019 -586 5113 -572
rect 5473 -572 5500 -548
rect 5567 -570 5599 -548
rect 5567 -572 5569 -570
rect 5597 -572 5599 -570
rect 5666 -572 5693 -548
rect 5473 -586 5567 -572
rect 5599 -586 5693 -572
rect 6053 -572 6080 -548
rect 6147 -570 6179 -548
rect 6147 -572 6149 -570
rect 6177 -572 6179 -570
rect 6246 -572 6273 -548
rect 6053 -586 6147 -572
rect 6179 -586 6273 -572
rect -404 -672 -386 -644
rect -356 -672 -338 -644
rect -96 -672 -78 -644
rect -48 -672 -29 -644
rect 176 -672 194 -644
rect 224 -672 242 -644
rect 484 -672 502 -644
rect 532 -672 551 -644
rect 756 -672 774 -644
rect 804 -672 822 -644
rect 1064 -672 1082 -644
rect 1112 -672 1131 -644
rect 1336 -672 1354 -644
rect 1384 -672 1402 -644
rect 1644 -672 1662 -644
rect 1692 -672 1711 -644
rect 1916 -672 1934 -644
rect 1964 -672 1982 -644
rect 2224 -672 2242 -644
rect 2272 -672 2291 -644
rect 2496 -672 2514 -644
rect 2544 -672 2562 -644
rect 2804 -672 2822 -644
rect 2852 -672 2871 -644
rect 3076 -672 3094 -644
rect 3124 -672 3142 -644
rect 3384 -672 3402 -644
rect 3432 -672 3451 -644
rect 3656 -672 3674 -644
rect 3704 -672 3722 -644
rect 3964 -672 3982 -644
rect 4012 -672 4031 -644
rect 4236 -672 4254 -644
rect 4284 -672 4302 -644
rect 4544 -672 4562 -644
rect 4592 -672 4611 -644
rect 4816 -672 4834 -644
rect 4864 -672 4882 -644
rect 5124 -672 5142 -644
rect 5172 -672 5191 -644
rect 5396 -672 5414 -644
rect 5444 -672 5462 -644
rect 5704 -672 5722 -644
rect 5752 -672 5771 -644
rect 5976 -672 5994 -644
rect 6024 -672 6042 -644
rect 6284 -672 6302 -644
rect 6332 -672 6351 -644
rect -478 -818 -450 -776
rect -420 -790 -395 -776
rect -296 -786 -271 -776
rect -420 -818 -364 -790
rect -334 -818 -300 -790
tri -286 -793 -279 -786 ne
rect -279 -818 -271 -786
rect -241 -818 -193 -776
rect -163 -786 -138 -776
rect -163 -818 -155 -786
rect -39 -790 -14 -776
rect -134 -818 -100 -790
rect -70 -818 -14 -790
rect 16 -818 44 -776
rect 102 -818 130 -776
rect 160 -790 185 -776
rect 284 -786 309 -776
rect 160 -818 216 -790
rect 246 -818 280 -790
tri 294 -793 301 -786 ne
rect 301 -818 309 -786
rect 339 -818 387 -776
rect 417 -786 442 -776
rect 417 -818 425 -786
rect 541 -790 566 -776
rect 446 -818 480 -790
rect 510 -818 566 -790
rect 596 -818 624 -776
rect 682 -818 710 -776
rect 740 -790 765 -776
rect 864 -786 889 -776
rect 740 -818 796 -790
rect 826 -818 860 -790
tri 874 -793 881 -786 ne
rect 881 -818 889 -786
rect 919 -818 967 -776
rect 997 -786 1022 -776
rect 997 -818 1005 -786
rect 1121 -790 1146 -776
rect 1026 -818 1060 -790
rect 1090 -818 1146 -790
rect 1176 -818 1204 -776
rect 1262 -818 1290 -776
rect 1320 -790 1345 -776
rect 1444 -786 1469 -776
rect 1320 -818 1376 -790
rect 1406 -818 1440 -790
tri 1454 -793 1461 -786 ne
rect 1461 -818 1469 -786
rect 1499 -818 1547 -776
rect 1577 -786 1602 -776
rect 1577 -818 1585 -786
rect 1701 -790 1726 -776
rect 1606 -818 1640 -790
rect 1670 -818 1726 -790
rect 1756 -818 1784 -776
rect 1842 -818 1870 -776
rect 1900 -790 1925 -776
rect 2024 -786 2049 -776
rect 1900 -818 1956 -790
rect 1986 -818 2020 -790
tri 2034 -793 2041 -786 ne
rect 2041 -818 2049 -786
rect 2079 -818 2127 -776
rect 2157 -786 2182 -776
rect 2157 -818 2165 -786
rect 2281 -790 2306 -776
rect 2186 -818 2220 -790
rect 2250 -818 2306 -790
rect 2336 -818 2364 -776
rect 2422 -818 2450 -776
rect 2480 -790 2505 -776
rect 2604 -786 2629 -776
rect 2480 -818 2536 -790
rect 2566 -818 2600 -790
tri 2614 -793 2621 -786 ne
rect 2621 -818 2629 -786
rect 2659 -818 2707 -776
rect 2737 -786 2762 -776
rect 2737 -818 2745 -786
rect 2861 -790 2886 -776
rect 2766 -818 2800 -790
rect 2830 -818 2886 -790
rect 2916 -818 2944 -776
rect 3002 -818 3030 -776
rect 3060 -790 3085 -776
rect 3184 -786 3209 -776
rect 3060 -818 3116 -790
rect 3146 -818 3180 -790
tri 3194 -793 3201 -786 ne
rect 3201 -818 3209 -786
rect 3239 -818 3287 -776
rect 3317 -786 3342 -776
rect 3317 -818 3325 -786
rect 3441 -790 3466 -776
rect 3346 -818 3380 -790
rect 3410 -818 3466 -790
rect 3496 -818 3524 -776
rect 3582 -818 3610 -776
rect 3640 -790 3665 -776
rect 3764 -786 3789 -776
rect 3640 -818 3696 -790
rect 3726 -818 3760 -790
tri 3774 -793 3781 -786 ne
rect 3781 -818 3789 -786
rect 3819 -818 3867 -776
rect 3897 -786 3922 -776
rect 3897 -818 3905 -786
rect 4021 -790 4046 -776
rect 3926 -818 3960 -790
rect 3990 -818 4046 -790
rect 4076 -818 4104 -776
rect 4162 -818 4190 -776
rect 4220 -790 4245 -776
rect 4344 -786 4369 -776
rect 4220 -818 4276 -790
rect 4306 -818 4340 -790
tri 4354 -793 4361 -786 ne
rect 4361 -818 4369 -786
rect 4399 -818 4447 -776
rect 4477 -786 4502 -776
rect 4477 -818 4485 -786
rect 4601 -790 4626 -776
rect 4506 -818 4540 -790
rect 4570 -818 4626 -790
rect 4656 -818 4684 -776
rect 4742 -818 4770 -776
rect 4800 -790 4825 -776
rect 4924 -786 4949 -776
rect 4800 -818 4856 -790
rect 4886 -818 4920 -790
tri 4934 -793 4941 -786 ne
rect 4941 -818 4949 -786
rect 4979 -818 5027 -776
rect 5057 -786 5082 -776
rect 5057 -818 5065 -786
rect 5181 -790 5206 -776
rect 5086 -818 5120 -790
rect 5150 -818 5206 -790
rect 5236 -818 5264 -776
rect 5322 -818 5350 -776
rect 5380 -790 5405 -776
rect 5504 -786 5529 -776
rect 5380 -818 5436 -790
rect 5466 -818 5500 -790
tri 5514 -793 5521 -786 ne
rect 5521 -818 5529 -786
rect 5559 -818 5607 -776
rect 5637 -786 5662 -776
rect 5637 -818 5645 -786
rect 5761 -790 5786 -776
rect 5666 -818 5700 -790
rect 5730 -818 5786 -790
rect 5816 -818 5844 -776
rect 5902 -818 5930 -776
rect 5960 -790 5985 -776
rect 6084 -786 6109 -776
rect 5960 -818 6016 -790
rect 6046 -818 6080 -790
tri 6094 -793 6101 -786 ne
rect 6101 -818 6109 -786
rect 6139 -818 6187 -776
rect 6217 -786 6242 -776
rect 6217 -818 6225 -786
rect 6341 -790 6366 -776
rect 6246 -818 6280 -790
rect 6310 -818 6366 -790
rect 6396 -818 6424 -776
rect -327 -842 -300 -818
rect -233 -840 -201 -818
rect -233 -842 -231 -840
rect -203 -842 -201 -840
rect -134 -842 -107 -818
rect -327 -856 -233 -842
rect -201 -856 -107 -842
rect 253 -842 280 -818
rect 347 -840 379 -818
rect 347 -842 349 -840
rect 377 -842 379 -840
rect 446 -842 473 -818
rect 253 -856 347 -842
rect 379 -856 473 -842
rect 833 -842 860 -818
rect 927 -840 959 -818
rect 927 -842 929 -840
rect 957 -842 959 -840
rect 1026 -842 1053 -818
rect 833 -856 927 -842
rect 959 -856 1053 -842
rect 1413 -842 1440 -818
rect 1507 -840 1539 -818
rect 1507 -842 1509 -840
rect 1537 -842 1539 -840
rect 1606 -842 1633 -818
rect 1413 -856 1507 -842
rect 1539 -856 1633 -842
rect 1993 -842 2020 -818
rect 2087 -840 2119 -818
rect 2087 -842 2089 -840
rect 2117 -842 2119 -840
rect 2186 -842 2213 -818
rect 1993 -856 2087 -842
rect 2119 -856 2213 -842
rect 2573 -842 2600 -818
rect 2667 -840 2699 -818
rect 2667 -842 2669 -840
rect 2697 -842 2699 -840
rect 2766 -842 2793 -818
rect 2573 -856 2667 -842
rect 2699 -856 2793 -842
rect 3153 -842 3180 -818
rect 3247 -840 3279 -818
rect 3247 -842 3249 -840
rect 3277 -842 3279 -840
rect 3346 -842 3373 -818
rect 3153 -856 3247 -842
rect 3279 -856 3373 -842
rect 3733 -842 3760 -818
rect 3827 -840 3859 -818
rect 3827 -842 3829 -840
rect 3857 -842 3859 -840
rect 3926 -842 3953 -818
rect 3733 -856 3827 -842
rect 3859 -856 3953 -842
rect 4313 -842 4340 -818
rect 4407 -840 4439 -818
rect 4407 -842 4409 -840
rect 4437 -842 4439 -840
rect 4506 -842 4533 -818
rect 4313 -856 4407 -842
rect 4439 -856 4533 -842
rect 4893 -842 4920 -818
rect 4987 -840 5019 -818
rect 4987 -842 4989 -840
rect 5017 -842 5019 -840
rect 5086 -842 5113 -818
rect 4893 -856 4987 -842
rect 5019 -856 5113 -842
rect 5473 -842 5500 -818
rect 5567 -840 5599 -818
rect 5567 -842 5569 -840
rect 5597 -842 5599 -840
rect 5666 -842 5693 -818
rect 5473 -856 5567 -842
rect 5599 -856 5693 -842
rect 6053 -842 6080 -818
rect 6147 -840 6179 -818
rect 6147 -842 6149 -840
rect 6177 -842 6179 -840
rect 6246 -842 6273 -818
rect 6053 -856 6147 -842
rect 6179 -856 6273 -842
rect -404 -942 -386 -914
rect -356 -942 -338 -914
rect -96 -942 -78 -914
rect -48 -942 -29 -914
rect 176 -942 194 -914
rect 224 -942 242 -914
rect 484 -942 502 -914
rect 532 -942 551 -914
rect 756 -942 774 -914
rect 804 -942 822 -914
rect 1064 -942 1082 -914
rect 1112 -942 1131 -914
rect 1336 -942 1354 -914
rect 1384 -942 1402 -914
rect 1644 -942 1662 -914
rect 1692 -942 1711 -914
rect 1916 -942 1934 -914
rect 1964 -942 1982 -914
rect 2224 -942 2242 -914
rect 2272 -942 2291 -914
rect 2496 -942 2514 -914
rect 2544 -942 2562 -914
rect 2804 -942 2822 -914
rect 2852 -942 2871 -914
rect 3076 -942 3094 -914
rect 3124 -942 3142 -914
rect 3384 -942 3402 -914
rect 3432 -942 3451 -914
rect 3656 -942 3674 -914
rect 3704 -942 3722 -914
rect 3964 -942 3982 -914
rect 4012 -942 4031 -914
rect 4236 -942 4254 -914
rect 4284 -942 4302 -914
rect 4544 -942 4562 -914
rect 4592 -942 4611 -914
rect 4816 -942 4834 -914
rect 4864 -942 4882 -914
rect 5124 -942 5142 -914
rect 5172 -942 5191 -914
rect 5396 -942 5414 -914
rect 5444 -942 5462 -914
rect 5704 -942 5722 -914
rect 5752 -942 5771 -914
rect 5976 -942 5994 -914
rect 6024 -942 6042 -914
rect 6284 -942 6302 -914
rect 6332 -942 6351 -914
rect -478 -1088 -450 -1046
rect -420 -1060 -395 -1046
rect -296 -1056 -271 -1046
rect -420 -1088 -364 -1060
rect -334 -1088 -300 -1060
tri -286 -1063 -279 -1056 ne
rect -279 -1088 -271 -1056
rect -241 -1088 -193 -1046
rect -163 -1056 -138 -1046
rect -163 -1088 -155 -1056
rect -39 -1060 -14 -1046
rect -134 -1088 -100 -1060
rect -70 -1088 -14 -1060
rect 16 -1088 44 -1046
rect 102 -1088 130 -1046
rect 160 -1060 185 -1046
rect 284 -1056 309 -1046
rect 160 -1088 216 -1060
rect 246 -1088 280 -1060
tri 294 -1063 301 -1056 ne
rect 301 -1088 309 -1056
rect 339 -1088 387 -1046
rect 417 -1056 442 -1046
rect 417 -1088 425 -1056
rect 541 -1060 566 -1046
rect 446 -1088 480 -1060
rect 510 -1088 566 -1060
rect 596 -1088 624 -1046
rect 682 -1088 710 -1046
rect 740 -1060 765 -1046
rect 864 -1056 889 -1046
rect 740 -1088 796 -1060
rect 826 -1088 860 -1060
tri 874 -1063 881 -1056 ne
rect 881 -1088 889 -1056
rect 919 -1088 967 -1046
rect 997 -1056 1022 -1046
rect 997 -1088 1005 -1056
rect 1121 -1060 1146 -1046
rect 1026 -1088 1060 -1060
rect 1090 -1088 1146 -1060
rect 1176 -1088 1204 -1046
rect 1262 -1088 1290 -1046
rect 1320 -1060 1345 -1046
rect 1444 -1056 1469 -1046
rect 1320 -1088 1376 -1060
rect 1406 -1088 1440 -1060
tri 1454 -1063 1461 -1056 ne
rect 1461 -1088 1469 -1056
rect 1499 -1088 1547 -1046
rect 1577 -1056 1602 -1046
rect 1577 -1088 1585 -1056
rect 1701 -1060 1726 -1046
rect 1606 -1088 1640 -1060
rect 1670 -1088 1726 -1060
rect 1756 -1088 1784 -1046
rect 1842 -1088 1870 -1046
rect 1900 -1060 1925 -1046
rect 2024 -1056 2049 -1046
rect 1900 -1088 1956 -1060
rect 1986 -1088 2020 -1060
tri 2034 -1063 2041 -1056 ne
rect 2041 -1088 2049 -1056
rect 2079 -1088 2127 -1046
rect 2157 -1056 2182 -1046
rect 2157 -1088 2165 -1056
rect 2281 -1060 2306 -1046
rect 2186 -1088 2220 -1060
rect 2250 -1088 2306 -1060
rect 2336 -1088 2364 -1046
rect 2422 -1088 2450 -1046
rect 2480 -1060 2505 -1046
rect 2604 -1056 2629 -1046
rect 2480 -1088 2536 -1060
rect 2566 -1088 2600 -1060
tri 2614 -1063 2621 -1056 ne
rect 2621 -1088 2629 -1056
rect 2659 -1088 2707 -1046
rect 2737 -1056 2762 -1046
rect 2737 -1088 2745 -1056
rect 2861 -1060 2886 -1046
rect 2766 -1088 2800 -1060
rect 2830 -1088 2886 -1060
rect 2916 -1088 2944 -1046
rect 3002 -1088 3030 -1046
rect 3060 -1060 3085 -1046
rect 3184 -1056 3209 -1046
rect 3060 -1088 3116 -1060
rect 3146 -1088 3180 -1060
tri 3194 -1063 3201 -1056 ne
rect 3201 -1088 3209 -1056
rect 3239 -1088 3287 -1046
rect 3317 -1056 3342 -1046
rect 3317 -1088 3325 -1056
rect 3441 -1060 3466 -1046
rect 3346 -1088 3380 -1060
rect 3410 -1088 3466 -1060
rect 3496 -1088 3524 -1046
rect 3582 -1088 3610 -1046
rect 3640 -1060 3665 -1046
rect 3764 -1056 3789 -1046
rect 3640 -1088 3696 -1060
rect 3726 -1088 3760 -1060
tri 3774 -1063 3781 -1056 ne
rect 3781 -1088 3789 -1056
rect 3819 -1088 3867 -1046
rect 3897 -1056 3922 -1046
rect 3897 -1088 3905 -1056
rect 4021 -1060 4046 -1046
rect 3926 -1088 3960 -1060
rect 3990 -1088 4046 -1060
rect 4076 -1088 4104 -1046
rect 4162 -1088 4190 -1046
rect 4220 -1060 4245 -1046
rect 4344 -1056 4369 -1046
rect 4220 -1088 4276 -1060
rect 4306 -1088 4340 -1060
tri 4354 -1063 4361 -1056 ne
rect 4361 -1088 4369 -1056
rect 4399 -1088 4447 -1046
rect 4477 -1056 4502 -1046
rect 4477 -1088 4485 -1056
rect 4601 -1060 4626 -1046
rect 4506 -1088 4540 -1060
rect 4570 -1088 4626 -1060
rect 4656 -1088 4684 -1046
rect 4742 -1088 4770 -1046
rect 4800 -1060 4825 -1046
rect 4924 -1056 4949 -1046
rect 4800 -1088 4856 -1060
rect 4886 -1088 4920 -1060
tri 4934 -1063 4941 -1056 ne
rect 4941 -1088 4949 -1056
rect 4979 -1088 5027 -1046
rect 5057 -1056 5082 -1046
rect 5057 -1088 5065 -1056
rect 5181 -1060 5206 -1046
rect 5086 -1088 5120 -1060
rect 5150 -1088 5206 -1060
rect 5236 -1088 5264 -1046
rect 5322 -1088 5350 -1046
rect 5380 -1060 5405 -1046
rect 5504 -1056 5529 -1046
rect 5380 -1088 5436 -1060
rect 5466 -1088 5500 -1060
tri 5514 -1063 5521 -1056 ne
rect 5521 -1088 5529 -1056
rect 5559 -1088 5607 -1046
rect 5637 -1056 5662 -1046
rect 5637 -1088 5645 -1056
rect 5761 -1060 5786 -1046
rect 5666 -1088 5700 -1060
rect 5730 -1088 5786 -1060
rect 5816 -1088 5844 -1046
rect 5902 -1088 5930 -1046
rect 5960 -1060 5985 -1046
rect 6084 -1056 6109 -1046
rect 5960 -1088 6016 -1060
rect 6046 -1088 6080 -1060
tri 6094 -1063 6101 -1056 ne
rect 6101 -1088 6109 -1056
rect 6139 -1088 6187 -1046
rect 6217 -1056 6242 -1046
rect 6217 -1088 6225 -1056
rect 6341 -1060 6366 -1046
rect 6246 -1088 6280 -1060
rect 6310 -1088 6366 -1060
rect 6396 -1088 6424 -1046
rect -327 -1112 -300 -1088
rect -233 -1110 -201 -1088
rect -233 -1112 -231 -1110
rect -203 -1112 -201 -1110
rect -134 -1112 -107 -1088
rect -327 -1126 -233 -1112
rect -201 -1126 -107 -1112
rect 253 -1112 280 -1088
rect 347 -1110 379 -1088
rect 347 -1112 349 -1110
rect 377 -1112 379 -1110
rect 446 -1112 473 -1088
rect 253 -1126 347 -1112
rect 379 -1126 473 -1112
rect 833 -1112 860 -1088
rect 927 -1110 959 -1088
rect 927 -1112 929 -1110
rect 957 -1112 959 -1110
rect 1026 -1112 1053 -1088
rect 833 -1126 927 -1112
rect 959 -1126 1053 -1112
rect 1413 -1112 1440 -1088
rect 1507 -1110 1539 -1088
rect 1507 -1112 1509 -1110
rect 1537 -1112 1539 -1110
rect 1606 -1112 1633 -1088
rect 1413 -1126 1507 -1112
rect 1539 -1126 1633 -1112
rect 1993 -1112 2020 -1088
rect 2087 -1110 2119 -1088
rect 2087 -1112 2089 -1110
rect 2117 -1112 2119 -1110
rect 2186 -1112 2213 -1088
rect 1993 -1126 2087 -1112
rect 2119 -1126 2213 -1112
rect 2573 -1112 2600 -1088
rect 2667 -1110 2699 -1088
rect 2667 -1112 2669 -1110
rect 2697 -1112 2699 -1110
rect 2766 -1112 2793 -1088
rect 2573 -1126 2667 -1112
rect 2699 -1126 2793 -1112
rect 3153 -1112 3180 -1088
rect 3247 -1110 3279 -1088
rect 3247 -1112 3249 -1110
rect 3277 -1112 3279 -1110
rect 3346 -1112 3373 -1088
rect 3153 -1126 3247 -1112
rect 3279 -1126 3373 -1112
rect 3733 -1112 3760 -1088
rect 3827 -1110 3859 -1088
rect 3827 -1112 3829 -1110
rect 3857 -1112 3859 -1110
rect 3926 -1112 3953 -1088
rect 3733 -1126 3827 -1112
rect 3859 -1126 3953 -1112
rect 4313 -1112 4340 -1088
rect 4407 -1110 4439 -1088
rect 4407 -1112 4409 -1110
rect 4437 -1112 4439 -1110
rect 4506 -1112 4533 -1088
rect 4313 -1126 4407 -1112
rect 4439 -1126 4533 -1112
rect 4893 -1112 4920 -1088
rect 4987 -1110 5019 -1088
rect 4987 -1112 4989 -1110
rect 5017 -1112 5019 -1110
rect 5086 -1112 5113 -1088
rect 4893 -1126 4987 -1112
rect 5019 -1126 5113 -1112
rect 5473 -1112 5500 -1088
rect 5567 -1110 5599 -1088
rect 5567 -1112 5569 -1110
rect 5597 -1112 5599 -1110
rect 5666 -1112 5693 -1088
rect 5473 -1126 5567 -1112
rect 5599 -1126 5693 -1112
rect 6053 -1112 6080 -1088
rect 6147 -1110 6179 -1088
rect 6147 -1112 6149 -1110
rect 6177 -1112 6179 -1110
rect 6246 -1112 6273 -1088
rect 6053 -1126 6147 -1112
rect 6179 -1126 6273 -1112
rect -404 -1212 -386 -1184
rect -356 -1212 -338 -1184
rect -96 -1212 -78 -1184
rect -48 -1212 -29 -1184
rect 176 -1212 194 -1184
rect 224 -1212 242 -1184
rect 484 -1212 502 -1184
rect 532 -1212 551 -1184
rect 756 -1212 774 -1184
rect 804 -1212 822 -1184
rect 1064 -1212 1082 -1184
rect 1112 -1212 1131 -1184
rect 1336 -1212 1354 -1184
rect 1384 -1212 1402 -1184
rect 1644 -1212 1662 -1184
rect 1692 -1212 1711 -1184
rect 1916 -1212 1934 -1184
rect 1964 -1212 1982 -1184
rect 2224 -1212 2242 -1184
rect 2272 -1212 2291 -1184
rect 2496 -1212 2514 -1184
rect 2544 -1212 2562 -1184
rect 2804 -1212 2822 -1184
rect 2852 -1212 2871 -1184
rect 3076 -1212 3094 -1184
rect 3124 -1212 3142 -1184
rect 3384 -1212 3402 -1184
rect 3432 -1212 3451 -1184
rect 3656 -1212 3674 -1184
rect 3704 -1212 3722 -1184
rect 3964 -1212 3982 -1184
rect 4012 -1212 4031 -1184
rect 4236 -1212 4254 -1184
rect 4284 -1212 4302 -1184
rect 4544 -1212 4562 -1184
rect 4592 -1212 4611 -1184
rect 4816 -1212 4834 -1184
rect 4864 -1212 4882 -1184
rect 5124 -1212 5142 -1184
rect 5172 -1212 5191 -1184
rect 5396 -1212 5414 -1184
rect 5444 -1212 5462 -1184
rect 5704 -1212 5722 -1184
rect 5752 -1212 5771 -1184
rect 5976 -1212 5994 -1184
rect 6024 -1212 6042 -1184
rect 6284 -1212 6302 -1184
rect 6332 -1212 6351 -1184
rect -478 -1358 -450 -1316
rect -420 -1330 -395 -1316
rect -296 -1326 -271 -1316
rect -420 -1358 -364 -1330
rect -334 -1358 -300 -1330
tri -286 -1333 -279 -1326 ne
rect -279 -1358 -271 -1326
rect -241 -1358 -193 -1316
rect -163 -1326 -138 -1316
rect -163 -1358 -155 -1326
rect -39 -1330 -14 -1316
rect -134 -1358 -100 -1330
rect -70 -1358 -14 -1330
rect 16 -1358 44 -1316
rect 102 -1358 130 -1316
rect 160 -1330 185 -1316
rect 284 -1326 309 -1316
rect 160 -1358 216 -1330
rect 246 -1358 280 -1330
tri 294 -1333 301 -1326 ne
rect 301 -1358 309 -1326
rect 339 -1358 387 -1316
rect 417 -1326 442 -1316
rect 417 -1358 425 -1326
rect 541 -1330 566 -1316
rect 446 -1358 480 -1330
rect 510 -1358 566 -1330
rect 596 -1358 624 -1316
rect 682 -1358 710 -1316
rect 740 -1330 765 -1316
rect 864 -1326 889 -1316
rect 740 -1358 796 -1330
rect 826 -1358 860 -1330
tri 874 -1333 881 -1326 ne
rect 881 -1358 889 -1326
rect 919 -1358 967 -1316
rect 997 -1326 1022 -1316
rect 997 -1358 1005 -1326
rect 1121 -1330 1146 -1316
rect 1026 -1358 1060 -1330
rect 1090 -1358 1146 -1330
rect 1176 -1358 1204 -1316
rect 1262 -1358 1290 -1316
rect 1320 -1330 1345 -1316
rect 1444 -1326 1469 -1316
rect 1320 -1358 1376 -1330
rect 1406 -1358 1440 -1330
tri 1454 -1333 1461 -1326 ne
rect 1461 -1358 1469 -1326
rect 1499 -1358 1547 -1316
rect 1577 -1326 1602 -1316
rect 1577 -1358 1585 -1326
rect 1701 -1330 1726 -1316
rect 1606 -1358 1640 -1330
rect 1670 -1358 1726 -1330
rect 1756 -1358 1784 -1316
rect 1842 -1358 1870 -1316
rect 1900 -1330 1925 -1316
rect 2024 -1326 2049 -1316
rect 1900 -1358 1956 -1330
rect 1986 -1358 2020 -1330
tri 2034 -1333 2041 -1326 ne
rect 2041 -1358 2049 -1326
rect 2079 -1358 2127 -1316
rect 2157 -1326 2182 -1316
rect 2157 -1358 2165 -1326
rect 2281 -1330 2306 -1316
rect 2186 -1358 2220 -1330
rect 2250 -1358 2306 -1330
rect 2336 -1358 2364 -1316
rect 2422 -1358 2450 -1316
rect 2480 -1330 2505 -1316
rect 2604 -1326 2629 -1316
rect 2480 -1358 2536 -1330
rect 2566 -1358 2600 -1330
tri 2614 -1333 2621 -1326 ne
rect 2621 -1358 2629 -1326
rect 2659 -1358 2707 -1316
rect 2737 -1326 2762 -1316
rect 2737 -1358 2745 -1326
rect 2861 -1330 2886 -1316
rect 2766 -1358 2800 -1330
rect 2830 -1358 2886 -1330
rect 2916 -1358 2944 -1316
rect 3002 -1358 3030 -1316
rect 3060 -1330 3085 -1316
rect 3184 -1326 3209 -1316
rect 3060 -1358 3116 -1330
rect 3146 -1358 3180 -1330
tri 3194 -1333 3201 -1326 ne
rect 3201 -1358 3209 -1326
rect 3239 -1358 3287 -1316
rect 3317 -1326 3342 -1316
rect 3317 -1358 3325 -1326
rect 3441 -1330 3466 -1316
rect 3346 -1358 3380 -1330
rect 3410 -1358 3466 -1330
rect 3496 -1358 3524 -1316
rect 3582 -1358 3610 -1316
rect 3640 -1330 3665 -1316
rect 3764 -1326 3789 -1316
rect 3640 -1358 3696 -1330
rect 3726 -1358 3760 -1330
tri 3774 -1333 3781 -1326 ne
rect 3781 -1358 3789 -1326
rect 3819 -1358 3867 -1316
rect 3897 -1326 3922 -1316
rect 3897 -1358 3905 -1326
rect 4021 -1330 4046 -1316
rect 3926 -1358 3960 -1330
rect 3990 -1358 4046 -1330
rect 4076 -1358 4104 -1316
rect 4162 -1358 4190 -1316
rect 4220 -1330 4245 -1316
rect 4344 -1326 4369 -1316
rect 4220 -1358 4276 -1330
rect 4306 -1358 4340 -1330
tri 4354 -1333 4361 -1326 ne
rect 4361 -1358 4369 -1326
rect 4399 -1358 4447 -1316
rect 4477 -1326 4502 -1316
rect 4477 -1358 4485 -1326
rect 4601 -1330 4626 -1316
rect 4506 -1358 4540 -1330
rect 4570 -1358 4626 -1330
rect 4656 -1358 4684 -1316
rect 4742 -1358 4770 -1316
rect 4800 -1330 4825 -1316
rect 4924 -1326 4949 -1316
rect 4800 -1358 4856 -1330
rect 4886 -1358 4920 -1330
tri 4934 -1333 4941 -1326 ne
rect 4941 -1358 4949 -1326
rect 4979 -1358 5027 -1316
rect 5057 -1326 5082 -1316
rect 5057 -1358 5065 -1326
rect 5181 -1330 5206 -1316
rect 5086 -1358 5120 -1330
rect 5150 -1358 5206 -1330
rect 5236 -1358 5264 -1316
rect 5322 -1358 5350 -1316
rect 5380 -1330 5405 -1316
rect 5504 -1326 5529 -1316
rect 5380 -1358 5436 -1330
rect 5466 -1358 5500 -1330
tri 5514 -1333 5521 -1326 ne
rect 5521 -1358 5529 -1326
rect 5559 -1358 5607 -1316
rect 5637 -1326 5662 -1316
rect 5637 -1358 5645 -1326
rect 5761 -1330 5786 -1316
rect 5666 -1358 5700 -1330
rect 5730 -1358 5786 -1330
rect 5816 -1358 5844 -1316
rect 5902 -1358 5930 -1316
rect 5960 -1330 5985 -1316
rect 6084 -1326 6109 -1316
rect 5960 -1358 6016 -1330
rect 6046 -1358 6080 -1330
tri 6094 -1333 6101 -1326 ne
rect 6101 -1358 6109 -1326
rect 6139 -1358 6187 -1316
rect 6217 -1326 6242 -1316
rect 6217 -1358 6225 -1326
rect 6341 -1330 6366 -1316
rect 6246 -1358 6280 -1330
rect 6310 -1358 6366 -1330
rect 6396 -1358 6424 -1316
rect -327 -1382 -300 -1358
rect -233 -1380 -201 -1358
rect -233 -1382 -231 -1380
rect -203 -1382 -201 -1380
rect -134 -1382 -107 -1358
rect -327 -1396 -233 -1382
rect -201 -1396 -107 -1382
rect 253 -1382 280 -1358
rect 347 -1380 379 -1358
rect 347 -1382 349 -1380
rect 377 -1382 379 -1380
rect 446 -1382 473 -1358
rect 253 -1396 347 -1382
rect 379 -1396 473 -1382
rect 833 -1382 860 -1358
rect 927 -1380 959 -1358
rect 927 -1382 929 -1380
rect 957 -1382 959 -1380
rect 1026 -1382 1053 -1358
rect 833 -1396 927 -1382
rect 959 -1396 1053 -1382
rect 1413 -1382 1440 -1358
rect 1507 -1380 1539 -1358
rect 1507 -1382 1509 -1380
rect 1537 -1382 1539 -1380
rect 1606 -1382 1633 -1358
rect 1413 -1396 1507 -1382
rect 1539 -1396 1633 -1382
rect 1993 -1382 2020 -1358
rect 2087 -1380 2119 -1358
rect 2087 -1382 2089 -1380
rect 2117 -1382 2119 -1380
rect 2186 -1382 2213 -1358
rect 1993 -1396 2087 -1382
rect 2119 -1396 2213 -1382
rect 2573 -1382 2600 -1358
rect 2667 -1380 2699 -1358
rect 2667 -1382 2669 -1380
rect 2697 -1382 2699 -1380
rect 2766 -1382 2793 -1358
rect 2573 -1396 2667 -1382
rect 2699 -1396 2793 -1382
rect 3153 -1382 3180 -1358
rect 3247 -1380 3279 -1358
rect 3247 -1382 3249 -1380
rect 3277 -1382 3279 -1380
rect 3346 -1382 3373 -1358
rect 3153 -1396 3247 -1382
rect 3279 -1396 3373 -1382
rect 3733 -1382 3760 -1358
rect 3827 -1380 3859 -1358
rect 3827 -1382 3829 -1380
rect 3857 -1382 3859 -1380
rect 3926 -1382 3953 -1358
rect 3733 -1396 3827 -1382
rect 3859 -1396 3953 -1382
rect 4313 -1382 4340 -1358
rect 4407 -1380 4439 -1358
rect 4407 -1382 4409 -1380
rect 4437 -1382 4439 -1380
rect 4506 -1382 4533 -1358
rect 4313 -1396 4407 -1382
rect 4439 -1396 4533 -1382
rect 4893 -1382 4920 -1358
rect 4987 -1380 5019 -1358
rect 4987 -1382 4989 -1380
rect 5017 -1382 5019 -1380
rect 5086 -1382 5113 -1358
rect 4893 -1396 4987 -1382
rect 5019 -1396 5113 -1382
rect 5473 -1382 5500 -1358
rect 5567 -1380 5599 -1358
rect 5567 -1382 5569 -1380
rect 5597 -1382 5599 -1380
rect 5666 -1382 5693 -1358
rect 5473 -1396 5567 -1382
rect 5599 -1396 5693 -1382
rect 6053 -1382 6080 -1358
rect 6147 -1380 6179 -1358
rect 6147 -1382 6149 -1380
rect 6177 -1382 6179 -1380
rect 6246 -1382 6273 -1358
rect 6053 -1396 6147 -1382
rect 6179 -1396 6273 -1382
rect -404 -1482 -386 -1454
rect -356 -1482 -338 -1454
rect -96 -1482 -78 -1454
rect -48 -1482 -29 -1454
rect 176 -1482 194 -1454
rect 224 -1482 242 -1454
rect 484 -1482 502 -1454
rect 532 -1482 551 -1454
rect 756 -1482 774 -1454
rect 804 -1482 822 -1454
rect 1064 -1482 1082 -1454
rect 1112 -1482 1131 -1454
rect 1336 -1482 1354 -1454
rect 1384 -1482 1402 -1454
rect 1644 -1482 1662 -1454
rect 1692 -1482 1711 -1454
rect 1916 -1482 1934 -1454
rect 1964 -1482 1982 -1454
rect 2224 -1482 2242 -1454
rect 2272 -1482 2291 -1454
rect 2496 -1482 2514 -1454
rect 2544 -1482 2562 -1454
rect 2804 -1482 2822 -1454
rect 2852 -1482 2871 -1454
rect 3076 -1482 3094 -1454
rect 3124 -1482 3142 -1454
rect 3384 -1482 3402 -1454
rect 3432 -1482 3451 -1454
rect 3656 -1482 3674 -1454
rect 3704 -1482 3722 -1454
rect 3964 -1482 3982 -1454
rect 4012 -1482 4031 -1454
rect 4236 -1482 4254 -1454
rect 4284 -1482 4302 -1454
rect 4544 -1482 4562 -1454
rect 4592 -1482 4611 -1454
rect 4816 -1482 4834 -1454
rect 4864 -1482 4882 -1454
rect 5124 -1482 5142 -1454
rect 5172 -1482 5191 -1454
rect 5396 -1482 5414 -1454
rect 5444 -1482 5462 -1454
rect 5704 -1482 5722 -1454
rect 5752 -1482 5771 -1454
rect 5976 -1482 5994 -1454
rect 6024 -1482 6042 -1454
rect 6284 -1482 6302 -1454
rect 6332 -1482 6351 -1454
rect -478 -1628 -450 -1586
rect -420 -1600 -395 -1586
rect -296 -1596 -271 -1586
rect -420 -1628 -364 -1600
rect -334 -1628 -300 -1600
tri -286 -1603 -279 -1596 ne
rect -279 -1628 -271 -1596
rect -241 -1628 -193 -1586
rect -163 -1596 -138 -1586
rect -163 -1628 -155 -1596
rect -39 -1600 -14 -1586
rect -134 -1628 -100 -1600
rect -70 -1628 -14 -1600
rect 16 -1628 44 -1586
rect 102 -1628 130 -1586
rect 160 -1600 185 -1586
rect 284 -1596 309 -1586
rect 160 -1628 216 -1600
rect 246 -1628 280 -1600
tri 294 -1603 301 -1596 ne
rect 301 -1628 309 -1596
rect 339 -1628 387 -1586
rect 417 -1596 442 -1586
rect 417 -1628 425 -1596
rect 541 -1600 566 -1586
rect 446 -1628 480 -1600
rect 510 -1628 566 -1600
rect 596 -1628 624 -1586
rect 682 -1628 710 -1586
rect 740 -1600 765 -1586
rect 864 -1596 889 -1586
rect 740 -1628 796 -1600
rect 826 -1628 860 -1600
tri 874 -1603 881 -1596 ne
rect 881 -1628 889 -1596
rect 919 -1628 967 -1586
rect 997 -1596 1022 -1586
rect 997 -1628 1005 -1596
rect 1121 -1600 1146 -1586
rect 1026 -1628 1060 -1600
rect 1090 -1628 1146 -1600
rect 1176 -1628 1204 -1586
rect 1262 -1628 1290 -1586
rect 1320 -1600 1345 -1586
rect 1444 -1596 1469 -1586
rect 1320 -1628 1376 -1600
rect 1406 -1628 1440 -1600
tri 1454 -1603 1461 -1596 ne
rect 1461 -1628 1469 -1596
rect 1499 -1628 1547 -1586
rect 1577 -1596 1602 -1586
rect 1577 -1628 1585 -1596
rect 1701 -1600 1726 -1586
rect 1606 -1628 1640 -1600
rect 1670 -1628 1726 -1600
rect 1756 -1628 1784 -1586
rect 1842 -1628 1870 -1586
rect 1900 -1600 1925 -1586
rect 2024 -1596 2049 -1586
rect 1900 -1628 1956 -1600
rect 1986 -1628 2020 -1600
tri 2034 -1603 2041 -1596 ne
rect 2041 -1628 2049 -1596
rect 2079 -1628 2127 -1586
rect 2157 -1596 2182 -1586
rect 2157 -1628 2165 -1596
rect 2281 -1600 2306 -1586
rect 2186 -1628 2220 -1600
rect 2250 -1628 2306 -1600
rect 2336 -1628 2364 -1586
rect 2422 -1628 2450 -1586
rect 2480 -1600 2505 -1586
rect 2604 -1596 2629 -1586
rect 2480 -1628 2536 -1600
rect 2566 -1628 2600 -1600
tri 2614 -1603 2621 -1596 ne
rect 2621 -1628 2629 -1596
rect 2659 -1628 2707 -1586
rect 2737 -1596 2762 -1586
rect 2737 -1628 2745 -1596
rect 2861 -1600 2886 -1586
rect 2766 -1628 2800 -1600
rect 2830 -1628 2886 -1600
rect 2916 -1628 2944 -1586
rect 3002 -1628 3030 -1586
rect 3060 -1600 3085 -1586
rect 3184 -1596 3209 -1586
rect 3060 -1628 3116 -1600
rect 3146 -1628 3180 -1600
tri 3194 -1603 3201 -1596 ne
rect 3201 -1628 3209 -1596
rect 3239 -1628 3287 -1586
rect 3317 -1596 3342 -1586
rect 3317 -1628 3325 -1596
rect 3441 -1600 3466 -1586
rect 3346 -1628 3380 -1600
rect 3410 -1628 3466 -1600
rect 3496 -1628 3524 -1586
rect 3582 -1628 3610 -1586
rect 3640 -1600 3665 -1586
rect 3764 -1596 3789 -1586
rect 3640 -1628 3696 -1600
rect 3726 -1628 3760 -1600
tri 3774 -1603 3781 -1596 ne
rect 3781 -1628 3789 -1596
rect 3819 -1628 3867 -1586
rect 3897 -1596 3922 -1586
rect 3897 -1628 3905 -1596
rect 4021 -1600 4046 -1586
rect 3926 -1628 3960 -1600
rect 3990 -1628 4046 -1600
rect 4076 -1628 4104 -1586
rect 4162 -1628 4190 -1586
rect 4220 -1600 4245 -1586
rect 4344 -1596 4369 -1586
rect 4220 -1628 4276 -1600
rect 4306 -1628 4340 -1600
tri 4354 -1603 4361 -1596 ne
rect 4361 -1628 4369 -1596
rect 4399 -1628 4447 -1586
rect 4477 -1596 4502 -1586
rect 4477 -1628 4485 -1596
rect 4601 -1600 4626 -1586
rect 4506 -1628 4540 -1600
rect 4570 -1628 4626 -1600
rect 4656 -1628 4684 -1586
rect 4742 -1628 4770 -1586
rect 4800 -1600 4825 -1586
rect 4924 -1596 4949 -1586
rect 4800 -1628 4856 -1600
rect 4886 -1628 4920 -1600
tri 4934 -1603 4941 -1596 ne
rect 4941 -1628 4949 -1596
rect 4979 -1628 5027 -1586
rect 5057 -1596 5082 -1586
rect 5057 -1628 5065 -1596
rect 5181 -1600 5206 -1586
rect 5086 -1628 5120 -1600
rect 5150 -1628 5206 -1600
rect 5236 -1628 5264 -1586
rect 5322 -1628 5350 -1586
rect 5380 -1600 5405 -1586
rect 5504 -1596 5529 -1586
rect 5380 -1628 5436 -1600
rect 5466 -1628 5500 -1600
tri 5514 -1603 5521 -1596 ne
rect 5521 -1628 5529 -1596
rect 5559 -1628 5607 -1586
rect 5637 -1596 5662 -1586
rect 5637 -1628 5645 -1596
rect 5761 -1600 5786 -1586
rect 5666 -1628 5700 -1600
rect 5730 -1628 5786 -1600
rect 5816 -1628 5844 -1586
rect 5902 -1628 5930 -1586
rect 5960 -1600 5985 -1586
rect 6084 -1596 6109 -1586
rect 5960 -1628 6016 -1600
rect 6046 -1628 6080 -1600
tri 6094 -1603 6101 -1596 ne
rect 6101 -1628 6109 -1596
rect 6139 -1628 6187 -1586
rect 6217 -1596 6242 -1586
rect 6217 -1628 6225 -1596
rect 6341 -1600 6366 -1586
rect 6246 -1628 6280 -1600
rect 6310 -1628 6366 -1600
rect 6396 -1628 6424 -1586
rect -327 -1652 -300 -1628
rect -233 -1650 -201 -1628
rect -233 -1652 -231 -1650
rect -203 -1652 -201 -1650
rect -134 -1652 -107 -1628
rect -327 -1666 -233 -1652
rect -201 -1666 -107 -1652
rect 253 -1652 280 -1628
rect 347 -1650 379 -1628
rect 347 -1652 349 -1650
rect 377 -1652 379 -1650
rect 446 -1652 473 -1628
rect 253 -1666 347 -1652
rect 379 -1666 473 -1652
rect 833 -1652 860 -1628
rect 927 -1650 959 -1628
rect 927 -1652 929 -1650
rect 957 -1652 959 -1650
rect 1026 -1652 1053 -1628
rect 833 -1666 927 -1652
rect 959 -1666 1053 -1652
rect 1413 -1652 1440 -1628
rect 1507 -1650 1539 -1628
rect 1507 -1652 1509 -1650
rect 1537 -1652 1539 -1650
rect 1606 -1652 1633 -1628
rect 1413 -1666 1507 -1652
rect 1539 -1666 1633 -1652
rect 1993 -1652 2020 -1628
rect 2087 -1650 2119 -1628
rect 2087 -1652 2089 -1650
rect 2117 -1652 2119 -1650
rect 2186 -1652 2213 -1628
rect 1993 -1666 2087 -1652
rect 2119 -1666 2213 -1652
rect 2573 -1652 2600 -1628
rect 2667 -1650 2699 -1628
rect 2667 -1652 2669 -1650
rect 2697 -1652 2699 -1650
rect 2766 -1652 2793 -1628
rect 2573 -1666 2667 -1652
rect 2699 -1666 2793 -1652
rect 3153 -1652 3180 -1628
rect 3247 -1650 3279 -1628
rect 3247 -1652 3249 -1650
rect 3277 -1652 3279 -1650
rect 3346 -1652 3373 -1628
rect 3153 -1666 3247 -1652
rect 3279 -1666 3373 -1652
rect 3733 -1652 3760 -1628
rect 3827 -1650 3859 -1628
rect 3827 -1652 3829 -1650
rect 3857 -1652 3859 -1650
rect 3926 -1652 3953 -1628
rect 3733 -1666 3827 -1652
rect 3859 -1666 3953 -1652
rect 4313 -1652 4340 -1628
rect 4407 -1650 4439 -1628
rect 4407 -1652 4409 -1650
rect 4437 -1652 4439 -1650
rect 4506 -1652 4533 -1628
rect 4313 -1666 4407 -1652
rect 4439 -1666 4533 -1652
rect 4893 -1652 4920 -1628
rect 4987 -1650 5019 -1628
rect 4987 -1652 4989 -1650
rect 5017 -1652 5019 -1650
rect 5086 -1652 5113 -1628
rect 4893 -1666 4987 -1652
rect 5019 -1666 5113 -1652
rect 5473 -1652 5500 -1628
rect 5567 -1650 5599 -1628
rect 5567 -1652 5569 -1650
rect 5597 -1652 5599 -1650
rect 5666 -1652 5693 -1628
rect 5473 -1666 5567 -1652
rect 5599 -1666 5693 -1652
rect 6053 -1652 6080 -1628
rect 6147 -1650 6179 -1628
rect 6147 -1652 6149 -1650
rect 6177 -1652 6179 -1650
rect 6246 -1652 6273 -1628
rect 6053 -1666 6147 -1652
rect 6179 -1666 6273 -1652
rect -404 -1752 -386 -1724
rect -356 -1752 -338 -1724
rect -96 -1752 -78 -1724
rect -48 -1752 -29 -1724
rect 176 -1752 194 -1724
rect 224 -1752 242 -1724
rect 484 -1752 502 -1724
rect 532 -1752 551 -1724
rect 756 -1752 774 -1724
rect 804 -1752 822 -1724
rect 1064 -1752 1082 -1724
rect 1112 -1752 1131 -1724
rect 1336 -1752 1354 -1724
rect 1384 -1752 1402 -1724
rect 1644 -1752 1662 -1724
rect 1692 -1752 1711 -1724
rect 1916 -1752 1934 -1724
rect 1964 -1752 1982 -1724
rect 2224 -1752 2242 -1724
rect 2272 -1752 2291 -1724
rect 2496 -1752 2514 -1724
rect 2544 -1752 2562 -1724
rect 2804 -1752 2822 -1724
rect 2852 -1752 2871 -1724
rect 3076 -1752 3094 -1724
rect 3124 -1752 3142 -1724
rect 3384 -1752 3402 -1724
rect 3432 -1752 3451 -1724
rect 3656 -1752 3674 -1724
rect 3704 -1752 3722 -1724
rect 3964 -1752 3982 -1724
rect 4012 -1752 4031 -1724
rect 4236 -1752 4254 -1724
rect 4284 -1752 4302 -1724
rect 4544 -1752 4562 -1724
rect 4592 -1752 4611 -1724
rect 4816 -1752 4834 -1724
rect 4864 -1752 4882 -1724
rect 5124 -1752 5142 -1724
rect 5172 -1752 5191 -1724
rect 5396 -1752 5414 -1724
rect 5444 -1752 5462 -1724
rect 5704 -1752 5722 -1724
rect 5752 -1752 5771 -1724
rect 5976 -1752 5994 -1724
rect 6024 -1752 6042 -1724
rect 6284 -1752 6302 -1724
rect 6332 -1752 6351 -1724
rect -478 -1898 -450 -1856
rect -420 -1870 -395 -1856
rect -296 -1866 -271 -1856
rect -420 -1898 -364 -1870
rect -334 -1898 -300 -1870
tri -286 -1873 -279 -1866 ne
rect -279 -1898 -271 -1866
rect -241 -1898 -193 -1856
rect -163 -1866 -138 -1856
rect -163 -1898 -155 -1866
rect -39 -1870 -14 -1856
rect -134 -1898 -100 -1870
rect -70 -1898 -14 -1870
rect 16 -1898 44 -1856
rect 102 -1898 130 -1856
rect 160 -1870 185 -1856
rect 284 -1866 309 -1856
rect 160 -1898 216 -1870
rect 246 -1898 280 -1870
tri 294 -1873 301 -1866 ne
rect 301 -1898 309 -1866
rect 339 -1898 387 -1856
rect 417 -1866 442 -1856
rect 417 -1898 425 -1866
rect 541 -1870 566 -1856
rect 446 -1898 480 -1870
rect 510 -1898 566 -1870
rect 596 -1898 624 -1856
rect 682 -1898 710 -1856
rect 740 -1870 765 -1856
rect 864 -1866 889 -1856
rect 740 -1898 796 -1870
rect 826 -1898 860 -1870
tri 874 -1873 881 -1866 ne
rect 881 -1898 889 -1866
rect 919 -1898 967 -1856
rect 997 -1866 1022 -1856
rect 997 -1898 1005 -1866
rect 1121 -1870 1146 -1856
rect 1026 -1898 1060 -1870
rect 1090 -1898 1146 -1870
rect 1176 -1898 1204 -1856
rect 1262 -1898 1290 -1856
rect 1320 -1870 1345 -1856
rect 1444 -1866 1469 -1856
rect 1320 -1898 1376 -1870
rect 1406 -1898 1440 -1870
tri 1454 -1873 1461 -1866 ne
rect 1461 -1898 1469 -1866
rect 1499 -1898 1547 -1856
rect 1577 -1866 1602 -1856
rect 1577 -1898 1585 -1866
rect 1701 -1870 1726 -1856
rect 1606 -1898 1640 -1870
rect 1670 -1898 1726 -1870
rect 1756 -1898 1784 -1856
rect 1842 -1898 1870 -1856
rect 1900 -1870 1925 -1856
rect 2024 -1866 2049 -1856
rect 1900 -1898 1956 -1870
rect 1986 -1898 2020 -1870
tri 2034 -1873 2041 -1866 ne
rect 2041 -1898 2049 -1866
rect 2079 -1898 2127 -1856
rect 2157 -1866 2182 -1856
rect 2157 -1898 2165 -1866
rect 2281 -1870 2306 -1856
rect 2186 -1898 2220 -1870
rect 2250 -1898 2306 -1870
rect 2336 -1898 2364 -1856
rect 2422 -1898 2450 -1856
rect 2480 -1870 2505 -1856
rect 2604 -1866 2629 -1856
rect 2480 -1898 2536 -1870
rect 2566 -1898 2600 -1870
tri 2614 -1873 2621 -1866 ne
rect 2621 -1898 2629 -1866
rect 2659 -1898 2707 -1856
rect 2737 -1866 2762 -1856
rect 2737 -1898 2745 -1866
rect 2861 -1870 2886 -1856
rect 2766 -1898 2800 -1870
rect 2830 -1898 2886 -1870
rect 2916 -1898 2944 -1856
rect 3002 -1898 3030 -1856
rect 3060 -1870 3085 -1856
rect 3184 -1866 3209 -1856
rect 3060 -1898 3116 -1870
rect 3146 -1898 3180 -1870
tri 3194 -1873 3201 -1866 ne
rect 3201 -1898 3209 -1866
rect 3239 -1898 3287 -1856
rect 3317 -1866 3342 -1856
rect 3317 -1898 3325 -1866
rect 3441 -1870 3466 -1856
rect 3346 -1898 3380 -1870
rect 3410 -1898 3466 -1870
rect 3496 -1898 3524 -1856
rect 3582 -1898 3610 -1856
rect 3640 -1870 3665 -1856
rect 3764 -1866 3789 -1856
rect 3640 -1898 3696 -1870
rect 3726 -1898 3760 -1870
tri 3774 -1873 3781 -1866 ne
rect 3781 -1898 3789 -1866
rect 3819 -1898 3867 -1856
rect 3897 -1866 3922 -1856
rect 3897 -1898 3905 -1866
rect 4021 -1870 4046 -1856
rect 3926 -1898 3960 -1870
rect 3990 -1898 4046 -1870
rect 4076 -1898 4104 -1856
rect 4162 -1898 4190 -1856
rect 4220 -1870 4245 -1856
rect 4344 -1866 4369 -1856
rect 4220 -1898 4276 -1870
rect 4306 -1898 4340 -1870
tri 4354 -1873 4361 -1866 ne
rect 4361 -1898 4369 -1866
rect 4399 -1898 4447 -1856
rect 4477 -1866 4502 -1856
rect 4477 -1898 4485 -1866
rect 4601 -1870 4626 -1856
rect 4506 -1898 4540 -1870
rect 4570 -1898 4626 -1870
rect 4656 -1898 4684 -1856
rect 4742 -1898 4770 -1856
rect 4800 -1870 4825 -1856
rect 4924 -1866 4949 -1856
rect 4800 -1898 4856 -1870
rect 4886 -1898 4920 -1870
tri 4934 -1873 4941 -1866 ne
rect 4941 -1898 4949 -1866
rect 4979 -1898 5027 -1856
rect 5057 -1866 5082 -1856
rect 5057 -1898 5065 -1866
rect 5181 -1870 5206 -1856
rect 5086 -1898 5120 -1870
rect 5150 -1898 5206 -1870
rect 5236 -1898 5264 -1856
rect 5322 -1898 5350 -1856
rect 5380 -1870 5405 -1856
rect 5504 -1866 5529 -1856
rect 5380 -1898 5436 -1870
rect 5466 -1898 5500 -1870
tri 5514 -1873 5521 -1866 ne
rect 5521 -1898 5529 -1866
rect 5559 -1898 5607 -1856
rect 5637 -1866 5662 -1856
rect 5637 -1898 5645 -1866
rect 5761 -1870 5786 -1856
rect 5666 -1898 5700 -1870
rect 5730 -1898 5786 -1870
rect 5816 -1898 5844 -1856
rect 5902 -1898 5930 -1856
rect 5960 -1870 5985 -1856
rect 6084 -1866 6109 -1856
rect 5960 -1898 6016 -1870
rect 6046 -1898 6080 -1870
tri 6094 -1873 6101 -1866 ne
rect 6101 -1898 6109 -1866
rect 6139 -1898 6187 -1856
rect 6217 -1866 6242 -1856
rect 6217 -1898 6225 -1866
rect 6341 -1870 6366 -1856
rect 6246 -1898 6280 -1870
rect 6310 -1898 6366 -1870
rect 6396 -1898 6424 -1856
rect -327 -1922 -300 -1898
rect -233 -1920 -201 -1898
rect -233 -1922 -231 -1920
rect -203 -1922 -201 -1920
rect -134 -1922 -107 -1898
rect -327 -1936 -233 -1922
rect -201 -1936 -107 -1922
rect 253 -1922 280 -1898
rect 347 -1920 379 -1898
rect 347 -1922 349 -1920
rect 377 -1922 379 -1920
rect 446 -1922 473 -1898
rect 253 -1936 347 -1922
rect 379 -1936 473 -1922
rect 833 -1922 860 -1898
rect 927 -1920 959 -1898
rect 927 -1922 929 -1920
rect 957 -1922 959 -1920
rect 1026 -1922 1053 -1898
rect 833 -1936 927 -1922
rect 959 -1936 1053 -1922
rect 1413 -1922 1440 -1898
rect 1507 -1920 1539 -1898
rect 1507 -1922 1509 -1920
rect 1537 -1922 1539 -1920
rect 1606 -1922 1633 -1898
rect 1413 -1936 1507 -1922
rect 1539 -1936 1633 -1922
rect 1993 -1922 2020 -1898
rect 2087 -1920 2119 -1898
rect 2087 -1922 2089 -1920
rect 2117 -1922 2119 -1920
rect 2186 -1922 2213 -1898
rect 1993 -1936 2087 -1922
rect 2119 -1936 2213 -1922
rect 2573 -1922 2600 -1898
rect 2667 -1920 2699 -1898
rect 2667 -1922 2669 -1920
rect 2697 -1922 2699 -1920
rect 2766 -1922 2793 -1898
rect 2573 -1936 2667 -1922
rect 2699 -1936 2793 -1922
rect 3153 -1922 3180 -1898
rect 3247 -1920 3279 -1898
rect 3247 -1922 3249 -1920
rect 3277 -1922 3279 -1920
rect 3346 -1922 3373 -1898
rect 3153 -1936 3247 -1922
rect 3279 -1936 3373 -1922
rect 3733 -1922 3760 -1898
rect 3827 -1920 3859 -1898
rect 3827 -1922 3829 -1920
rect 3857 -1922 3859 -1920
rect 3926 -1922 3953 -1898
rect 3733 -1936 3827 -1922
rect 3859 -1936 3953 -1922
rect 4313 -1922 4340 -1898
rect 4407 -1920 4439 -1898
rect 4407 -1922 4409 -1920
rect 4437 -1922 4439 -1920
rect 4506 -1922 4533 -1898
rect 4313 -1936 4407 -1922
rect 4439 -1936 4533 -1922
rect 4893 -1922 4920 -1898
rect 4987 -1920 5019 -1898
rect 4987 -1922 4989 -1920
rect 5017 -1922 5019 -1920
rect 5086 -1922 5113 -1898
rect 4893 -1936 4987 -1922
rect 5019 -1936 5113 -1922
rect 5473 -1922 5500 -1898
rect 5567 -1920 5599 -1898
rect 5567 -1922 5569 -1920
rect 5597 -1922 5599 -1920
rect 5666 -1922 5693 -1898
rect 5473 -1936 5567 -1922
rect 5599 -1936 5693 -1922
rect 6053 -1922 6080 -1898
rect 6147 -1920 6179 -1898
rect 6147 -1922 6149 -1920
rect 6177 -1922 6179 -1920
rect 6246 -1922 6273 -1898
rect 6053 -1936 6147 -1922
rect 6179 -1936 6273 -1922
rect -404 -2022 -386 -1994
rect -356 -2022 -338 -1994
rect -96 -2022 -78 -1994
rect -48 -2022 -29 -1994
rect 176 -2022 194 -1994
rect 224 -2022 242 -1994
rect 484 -2022 502 -1994
rect 532 -2022 551 -1994
rect 756 -2022 774 -1994
rect 804 -2022 822 -1994
rect 1064 -2022 1082 -1994
rect 1112 -2022 1131 -1994
rect 1336 -2022 1354 -1994
rect 1384 -2022 1402 -1994
rect 1644 -2022 1662 -1994
rect 1692 -2022 1711 -1994
rect 1916 -2022 1934 -1994
rect 1964 -2022 1982 -1994
rect 2224 -2022 2242 -1994
rect 2272 -2022 2291 -1994
rect 2496 -2022 2514 -1994
rect 2544 -2022 2562 -1994
rect 2804 -2022 2822 -1994
rect 2852 -2022 2871 -1994
rect 3076 -2022 3094 -1994
rect 3124 -2022 3142 -1994
rect 3384 -2022 3402 -1994
rect 3432 -2022 3451 -1994
rect 3656 -2022 3674 -1994
rect 3704 -2022 3722 -1994
rect 3964 -2022 3982 -1994
rect 4012 -2022 4031 -1994
rect 4236 -2022 4254 -1994
rect 4284 -2022 4302 -1994
rect 4544 -2022 4562 -1994
rect 4592 -2022 4611 -1994
rect 4816 -2022 4834 -1994
rect 4864 -2022 4882 -1994
rect 5124 -2022 5142 -1994
rect 5172 -2022 5191 -1994
rect 5396 -2022 5414 -1994
rect 5444 -2022 5462 -1994
rect 5704 -2022 5722 -1994
rect 5752 -2022 5771 -1994
rect 5976 -2022 5994 -1994
rect 6024 -2022 6042 -1994
rect 6284 -2022 6302 -1994
rect 6332 -2022 6351 -1994
rect -478 -2168 -450 -2126
rect -420 -2140 -395 -2126
rect -296 -2136 -271 -2126
rect -420 -2168 -364 -2140
rect -334 -2168 -300 -2140
tri -286 -2143 -279 -2136 ne
rect -279 -2168 -271 -2136
rect -241 -2168 -193 -2126
rect -163 -2136 -138 -2126
rect -163 -2168 -155 -2136
rect -39 -2140 -14 -2126
rect -134 -2168 -100 -2140
rect -70 -2168 -14 -2140
rect 16 -2168 44 -2126
rect 102 -2168 130 -2126
rect 160 -2140 185 -2126
rect 284 -2136 309 -2126
rect 160 -2168 216 -2140
rect 246 -2168 280 -2140
tri 294 -2143 301 -2136 ne
rect 301 -2168 309 -2136
rect 339 -2168 387 -2126
rect 417 -2136 442 -2126
rect 417 -2168 425 -2136
rect 541 -2140 566 -2126
rect 446 -2168 480 -2140
rect 510 -2168 566 -2140
rect 596 -2168 624 -2126
rect 682 -2168 710 -2126
rect 740 -2140 765 -2126
rect 864 -2136 889 -2126
rect 740 -2168 796 -2140
rect 826 -2168 860 -2140
tri 874 -2143 881 -2136 ne
rect 881 -2168 889 -2136
rect 919 -2168 967 -2126
rect 997 -2136 1022 -2126
rect 997 -2168 1005 -2136
rect 1121 -2140 1146 -2126
rect 1026 -2168 1060 -2140
rect 1090 -2168 1146 -2140
rect 1176 -2168 1204 -2126
rect 1262 -2168 1290 -2126
rect 1320 -2140 1345 -2126
rect 1444 -2136 1469 -2126
rect 1320 -2168 1376 -2140
rect 1406 -2168 1440 -2140
tri 1454 -2143 1461 -2136 ne
rect 1461 -2168 1469 -2136
rect 1499 -2168 1547 -2126
rect 1577 -2136 1602 -2126
rect 1577 -2168 1585 -2136
rect 1701 -2140 1726 -2126
rect 1606 -2168 1640 -2140
rect 1670 -2168 1726 -2140
rect 1756 -2168 1784 -2126
rect 1842 -2168 1870 -2126
rect 1900 -2140 1925 -2126
rect 2024 -2136 2049 -2126
rect 1900 -2168 1956 -2140
rect 1986 -2168 2020 -2140
tri 2034 -2143 2041 -2136 ne
rect 2041 -2168 2049 -2136
rect 2079 -2168 2127 -2126
rect 2157 -2136 2182 -2126
rect 2157 -2168 2165 -2136
rect 2281 -2140 2306 -2126
rect 2186 -2168 2220 -2140
rect 2250 -2168 2306 -2140
rect 2336 -2168 2364 -2126
rect 2422 -2168 2450 -2126
rect 2480 -2140 2505 -2126
rect 2604 -2136 2629 -2126
rect 2480 -2168 2536 -2140
rect 2566 -2168 2600 -2140
tri 2614 -2143 2621 -2136 ne
rect 2621 -2168 2629 -2136
rect 2659 -2168 2707 -2126
rect 2737 -2136 2762 -2126
rect 2737 -2168 2745 -2136
rect 2861 -2140 2886 -2126
rect 2766 -2168 2800 -2140
rect 2830 -2168 2886 -2140
rect 2916 -2168 2944 -2126
rect 3002 -2168 3030 -2126
rect 3060 -2140 3085 -2126
rect 3184 -2136 3209 -2126
rect 3060 -2168 3116 -2140
rect 3146 -2168 3180 -2140
tri 3194 -2143 3201 -2136 ne
rect 3201 -2168 3209 -2136
rect 3239 -2168 3287 -2126
rect 3317 -2136 3342 -2126
rect 3317 -2168 3325 -2136
rect 3441 -2140 3466 -2126
rect 3346 -2168 3380 -2140
rect 3410 -2168 3466 -2140
rect 3496 -2168 3524 -2126
rect 3582 -2168 3610 -2126
rect 3640 -2140 3665 -2126
rect 3764 -2136 3789 -2126
rect 3640 -2168 3696 -2140
rect 3726 -2168 3760 -2140
tri 3774 -2143 3781 -2136 ne
rect 3781 -2168 3789 -2136
rect 3819 -2168 3867 -2126
rect 3897 -2136 3922 -2126
rect 3897 -2168 3905 -2136
rect 4021 -2140 4046 -2126
rect 3926 -2168 3960 -2140
rect 3990 -2168 4046 -2140
rect 4076 -2168 4104 -2126
rect 4162 -2168 4190 -2126
rect 4220 -2140 4245 -2126
rect 4344 -2136 4369 -2126
rect 4220 -2168 4276 -2140
rect 4306 -2168 4340 -2140
tri 4354 -2143 4361 -2136 ne
rect 4361 -2168 4369 -2136
rect 4399 -2168 4447 -2126
rect 4477 -2136 4502 -2126
rect 4477 -2168 4485 -2136
rect 4601 -2140 4626 -2126
rect 4506 -2168 4540 -2140
rect 4570 -2168 4626 -2140
rect 4656 -2168 4684 -2126
rect 4742 -2168 4770 -2126
rect 4800 -2140 4825 -2126
rect 4924 -2136 4949 -2126
rect 4800 -2168 4856 -2140
rect 4886 -2168 4920 -2140
tri 4934 -2143 4941 -2136 ne
rect 4941 -2168 4949 -2136
rect 4979 -2168 5027 -2126
rect 5057 -2136 5082 -2126
rect 5057 -2168 5065 -2136
rect 5181 -2140 5206 -2126
rect 5086 -2168 5120 -2140
rect 5150 -2168 5206 -2140
rect 5236 -2168 5264 -2126
rect 5322 -2168 5350 -2126
rect 5380 -2140 5405 -2126
rect 5504 -2136 5529 -2126
rect 5380 -2168 5436 -2140
rect 5466 -2168 5500 -2140
tri 5514 -2143 5521 -2136 ne
rect 5521 -2168 5529 -2136
rect 5559 -2168 5607 -2126
rect 5637 -2136 5662 -2126
rect 5637 -2168 5645 -2136
rect 5761 -2140 5786 -2126
rect 5666 -2168 5700 -2140
rect 5730 -2168 5786 -2140
rect 5816 -2168 5844 -2126
rect 5902 -2168 5930 -2126
rect 5960 -2140 5985 -2126
rect 6084 -2136 6109 -2126
rect 5960 -2168 6016 -2140
rect 6046 -2168 6080 -2140
tri 6094 -2143 6101 -2136 ne
rect 6101 -2168 6109 -2136
rect 6139 -2168 6187 -2126
rect 6217 -2136 6242 -2126
rect 6217 -2168 6225 -2136
rect 6341 -2140 6366 -2126
rect 6246 -2168 6280 -2140
rect 6310 -2168 6366 -2140
rect 6396 -2168 6424 -2126
rect -327 -2192 -300 -2168
rect -233 -2190 -201 -2168
rect -233 -2192 -231 -2190
rect -203 -2192 -201 -2190
rect -134 -2192 -107 -2168
rect -327 -2206 -233 -2192
rect -201 -2206 -107 -2192
rect 253 -2192 280 -2168
rect 347 -2190 379 -2168
rect 347 -2192 349 -2190
rect 377 -2192 379 -2190
rect 446 -2192 473 -2168
rect 253 -2206 347 -2192
rect 379 -2206 473 -2192
rect 833 -2192 860 -2168
rect 927 -2190 959 -2168
rect 927 -2192 929 -2190
rect 957 -2192 959 -2190
rect 1026 -2192 1053 -2168
rect 833 -2206 927 -2192
rect 959 -2206 1053 -2192
rect 1413 -2192 1440 -2168
rect 1507 -2190 1539 -2168
rect 1507 -2192 1509 -2190
rect 1537 -2192 1539 -2190
rect 1606 -2192 1633 -2168
rect 1413 -2206 1507 -2192
rect 1539 -2206 1633 -2192
rect 1993 -2192 2020 -2168
rect 2087 -2190 2119 -2168
rect 2087 -2192 2089 -2190
rect 2117 -2192 2119 -2190
rect 2186 -2192 2213 -2168
rect 1993 -2206 2087 -2192
rect 2119 -2206 2213 -2192
rect 2573 -2192 2600 -2168
rect 2667 -2190 2699 -2168
rect 2667 -2192 2669 -2190
rect 2697 -2192 2699 -2190
rect 2766 -2192 2793 -2168
rect 2573 -2206 2667 -2192
rect 2699 -2206 2793 -2192
rect 3153 -2192 3180 -2168
rect 3247 -2190 3279 -2168
rect 3247 -2192 3249 -2190
rect 3277 -2192 3279 -2190
rect 3346 -2192 3373 -2168
rect 3153 -2206 3247 -2192
rect 3279 -2206 3373 -2192
rect 3733 -2192 3760 -2168
rect 3827 -2190 3859 -2168
rect 3827 -2192 3829 -2190
rect 3857 -2192 3859 -2190
rect 3926 -2192 3953 -2168
rect 3733 -2206 3827 -2192
rect 3859 -2206 3953 -2192
rect 4313 -2192 4340 -2168
rect 4407 -2190 4439 -2168
rect 4407 -2192 4409 -2190
rect 4437 -2192 4439 -2190
rect 4506 -2192 4533 -2168
rect 4313 -2206 4407 -2192
rect 4439 -2206 4533 -2192
rect 4893 -2192 4920 -2168
rect 4987 -2190 5019 -2168
rect 4987 -2192 4989 -2190
rect 5017 -2192 5019 -2190
rect 5086 -2192 5113 -2168
rect 4893 -2206 4987 -2192
rect 5019 -2206 5113 -2192
rect 5473 -2192 5500 -2168
rect 5567 -2190 5599 -2168
rect 5567 -2192 5569 -2190
rect 5597 -2192 5599 -2190
rect 5666 -2192 5693 -2168
rect 5473 -2206 5567 -2192
rect 5599 -2206 5693 -2192
rect 6053 -2192 6080 -2168
rect 6147 -2190 6179 -2168
rect 6147 -2192 6149 -2190
rect 6177 -2192 6179 -2190
rect 6246 -2192 6273 -2168
rect 6053 -2206 6147 -2192
rect 6179 -2206 6273 -2192
rect -404 -2292 -386 -2264
rect -356 -2292 -338 -2264
rect -96 -2292 -78 -2264
rect -48 -2292 -29 -2264
rect 176 -2292 194 -2264
rect 224 -2292 242 -2264
rect 484 -2292 502 -2264
rect 532 -2292 551 -2264
rect 756 -2292 774 -2264
rect 804 -2292 822 -2264
rect 1064 -2292 1082 -2264
rect 1112 -2292 1131 -2264
rect 1336 -2292 1354 -2264
rect 1384 -2292 1402 -2264
rect 1644 -2292 1662 -2264
rect 1692 -2292 1711 -2264
rect 1916 -2292 1934 -2264
rect 1964 -2292 1982 -2264
rect 2224 -2292 2242 -2264
rect 2272 -2292 2291 -2264
rect 2496 -2292 2514 -2264
rect 2544 -2292 2562 -2264
rect 2804 -2292 2822 -2264
rect 2852 -2292 2871 -2264
rect 3076 -2292 3094 -2264
rect 3124 -2292 3142 -2264
rect 3384 -2292 3402 -2264
rect 3432 -2292 3451 -2264
rect 3656 -2292 3674 -2264
rect 3704 -2292 3722 -2264
rect 3964 -2292 3982 -2264
rect 4012 -2292 4031 -2264
rect 4236 -2292 4254 -2264
rect 4284 -2292 4302 -2264
rect 4544 -2292 4562 -2264
rect 4592 -2292 4611 -2264
rect 4816 -2292 4834 -2264
rect 4864 -2292 4882 -2264
rect 5124 -2292 5142 -2264
rect 5172 -2292 5191 -2264
rect 5396 -2292 5414 -2264
rect 5444 -2292 5462 -2264
rect 5704 -2292 5722 -2264
rect 5752 -2292 5771 -2264
rect 5976 -2292 5994 -2264
rect 6024 -2292 6042 -2264
rect 6284 -2292 6302 -2264
rect 6332 -2292 6351 -2264
rect -478 -2438 -450 -2396
rect -420 -2410 -395 -2396
rect -296 -2406 -271 -2396
rect -420 -2438 -364 -2410
rect -334 -2438 -300 -2410
tri -286 -2413 -279 -2406 ne
rect -279 -2438 -271 -2406
rect -241 -2438 -193 -2396
rect -163 -2406 -138 -2396
rect -163 -2438 -155 -2406
rect -39 -2410 -14 -2396
rect -134 -2438 -100 -2410
rect -70 -2438 -14 -2410
rect 16 -2438 44 -2396
rect 102 -2438 130 -2396
rect 160 -2410 185 -2396
rect 284 -2406 309 -2396
rect 160 -2438 216 -2410
rect 246 -2438 280 -2410
tri 294 -2413 301 -2406 ne
rect 301 -2438 309 -2406
rect 339 -2438 387 -2396
rect 417 -2406 442 -2396
rect 417 -2438 425 -2406
rect 541 -2410 566 -2396
rect 446 -2438 480 -2410
rect 510 -2438 566 -2410
rect 596 -2438 624 -2396
rect 682 -2438 710 -2396
rect 740 -2410 765 -2396
rect 864 -2406 889 -2396
rect 740 -2438 796 -2410
rect 826 -2438 860 -2410
tri 874 -2413 881 -2406 ne
rect 881 -2438 889 -2406
rect 919 -2438 967 -2396
rect 997 -2406 1022 -2396
rect 997 -2438 1005 -2406
rect 1121 -2410 1146 -2396
rect 1026 -2438 1060 -2410
rect 1090 -2438 1146 -2410
rect 1176 -2438 1204 -2396
rect 1262 -2438 1290 -2396
rect 1320 -2410 1345 -2396
rect 1444 -2406 1469 -2396
rect 1320 -2438 1376 -2410
rect 1406 -2438 1440 -2410
tri 1454 -2413 1461 -2406 ne
rect 1461 -2438 1469 -2406
rect 1499 -2438 1547 -2396
rect 1577 -2406 1602 -2396
rect 1577 -2438 1585 -2406
rect 1701 -2410 1726 -2396
rect 1606 -2438 1640 -2410
rect 1670 -2438 1726 -2410
rect 1756 -2438 1784 -2396
rect 1842 -2438 1870 -2396
rect 1900 -2410 1925 -2396
rect 2024 -2406 2049 -2396
rect 1900 -2438 1956 -2410
rect 1986 -2438 2020 -2410
tri 2034 -2413 2041 -2406 ne
rect 2041 -2438 2049 -2406
rect 2079 -2438 2127 -2396
rect 2157 -2406 2182 -2396
rect 2157 -2438 2165 -2406
rect 2281 -2410 2306 -2396
rect 2186 -2438 2220 -2410
rect 2250 -2438 2306 -2410
rect 2336 -2438 2364 -2396
rect 2422 -2438 2450 -2396
rect 2480 -2410 2505 -2396
rect 2604 -2406 2629 -2396
rect 2480 -2438 2536 -2410
rect 2566 -2438 2600 -2410
tri 2614 -2413 2621 -2406 ne
rect 2621 -2438 2629 -2406
rect 2659 -2438 2707 -2396
rect 2737 -2406 2762 -2396
rect 2737 -2438 2745 -2406
rect 2861 -2410 2886 -2396
rect 2766 -2438 2800 -2410
rect 2830 -2438 2886 -2410
rect 2916 -2438 2944 -2396
rect 3002 -2438 3030 -2396
rect 3060 -2410 3085 -2396
rect 3184 -2406 3209 -2396
rect 3060 -2438 3116 -2410
rect 3146 -2438 3180 -2410
tri 3194 -2413 3201 -2406 ne
rect 3201 -2438 3209 -2406
rect 3239 -2438 3287 -2396
rect 3317 -2406 3342 -2396
rect 3317 -2438 3325 -2406
rect 3441 -2410 3466 -2396
rect 3346 -2438 3380 -2410
rect 3410 -2438 3466 -2410
rect 3496 -2438 3524 -2396
rect 3582 -2438 3610 -2396
rect 3640 -2410 3665 -2396
rect 3764 -2406 3789 -2396
rect 3640 -2438 3696 -2410
rect 3726 -2438 3760 -2410
tri 3774 -2413 3781 -2406 ne
rect 3781 -2438 3789 -2406
rect 3819 -2438 3867 -2396
rect 3897 -2406 3922 -2396
rect 3897 -2438 3905 -2406
rect 4021 -2410 4046 -2396
rect 3926 -2438 3960 -2410
rect 3990 -2438 4046 -2410
rect 4076 -2438 4104 -2396
rect 4162 -2438 4190 -2396
rect 4220 -2410 4245 -2396
rect 4344 -2406 4369 -2396
rect 4220 -2438 4276 -2410
rect 4306 -2438 4340 -2410
tri 4354 -2413 4361 -2406 ne
rect 4361 -2438 4369 -2406
rect 4399 -2438 4447 -2396
rect 4477 -2406 4502 -2396
rect 4477 -2438 4485 -2406
rect 4601 -2410 4626 -2396
rect 4506 -2438 4540 -2410
rect 4570 -2438 4626 -2410
rect 4656 -2438 4684 -2396
rect 4742 -2438 4770 -2396
rect 4800 -2410 4825 -2396
rect 4924 -2406 4949 -2396
rect 4800 -2438 4856 -2410
rect 4886 -2438 4920 -2410
tri 4934 -2413 4941 -2406 ne
rect 4941 -2438 4949 -2406
rect 4979 -2438 5027 -2396
rect 5057 -2406 5082 -2396
rect 5057 -2438 5065 -2406
rect 5181 -2410 5206 -2396
rect 5086 -2438 5120 -2410
rect 5150 -2438 5206 -2410
rect 5236 -2438 5264 -2396
rect 5322 -2438 5350 -2396
rect 5380 -2410 5405 -2396
rect 5504 -2406 5529 -2396
rect 5380 -2438 5436 -2410
rect 5466 -2438 5500 -2410
tri 5514 -2413 5521 -2406 ne
rect 5521 -2438 5529 -2406
rect 5559 -2438 5607 -2396
rect 5637 -2406 5662 -2396
rect 5637 -2438 5645 -2406
rect 5761 -2410 5786 -2396
rect 5666 -2438 5700 -2410
rect 5730 -2438 5786 -2410
rect 5816 -2438 5844 -2396
rect 5902 -2438 5930 -2396
rect 5960 -2410 5985 -2396
rect 6084 -2406 6109 -2396
rect 5960 -2438 6016 -2410
rect 6046 -2438 6080 -2410
tri 6094 -2413 6101 -2406 ne
rect 6101 -2438 6109 -2406
rect 6139 -2438 6187 -2396
rect 6217 -2406 6242 -2396
rect 6217 -2438 6225 -2406
rect 6341 -2410 6366 -2396
rect 6246 -2438 6280 -2410
rect 6310 -2438 6366 -2410
rect 6396 -2438 6424 -2396
rect -327 -2462 -300 -2438
rect -233 -2460 -201 -2438
rect -233 -2462 -231 -2460
rect -203 -2462 -201 -2460
rect -134 -2462 -107 -2438
rect -327 -2476 -233 -2462
rect -201 -2476 -107 -2462
rect 253 -2462 280 -2438
rect 347 -2460 379 -2438
rect 347 -2462 349 -2460
rect 377 -2462 379 -2460
rect 446 -2462 473 -2438
rect 253 -2476 347 -2462
rect 379 -2476 473 -2462
rect 833 -2462 860 -2438
rect 927 -2460 959 -2438
rect 927 -2462 929 -2460
rect 957 -2462 959 -2460
rect 1026 -2462 1053 -2438
rect 833 -2476 927 -2462
rect 959 -2476 1053 -2462
rect 1413 -2462 1440 -2438
rect 1507 -2460 1539 -2438
rect 1507 -2462 1509 -2460
rect 1537 -2462 1539 -2460
rect 1606 -2462 1633 -2438
rect 1413 -2476 1507 -2462
rect 1539 -2476 1633 -2462
rect 1993 -2462 2020 -2438
rect 2087 -2460 2119 -2438
rect 2087 -2462 2089 -2460
rect 2117 -2462 2119 -2460
rect 2186 -2462 2213 -2438
rect 1993 -2476 2087 -2462
rect 2119 -2476 2213 -2462
rect 2573 -2462 2600 -2438
rect 2667 -2460 2699 -2438
rect 2667 -2462 2669 -2460
rect 2697 -2462 2699 -2460
rect 2766 -2462 2793 -2438
rect 2573 -2476 2667 -2462
rect 2699 -2476 2793 -2462
rect 3153 -2462 3180 -2438
rect 3247 -2460 3279 -2438
rect 3247 -2462 3249 -2460
rect 3277 -2462 3279 -2460
rect 3346 -2462 3373 -2438
rect 3153 -2476 3247 -2462
rect 3279 -2476 3373 -2462
rect 3733 -2462 3760 -2438
rect 3827 -2460 3859 -2438
rect 3827 -2462 3829 -2460
rect 3857 -2462 3859 -2460
rect 3926 -2462 3953 -2438
rect 3733 -2476 3827 -2462
rect 3859 -2476 3953 -2462
rect 4313 -2462 4340 -2438
rect 4407 -2460 4439 -2438
rect 4407 -2462 4409 -2460
rect 4437 -2462 4439 -2460
rect 4506 -2462 4533 -2438
rect 4313 -2476 4407 -2462
rect 4439 -2476 4533 -2462
rect 4893 -2462 4920 -2438
rect 4987 -2460 5019 -2438
rect 4987 -2462 4989 -2460
rect 5017 -2462 5019 -2460
rect 5086 -2462 5113 -2438
rect 4893 -2476 4987 -2462
rect 5019 -2476 5113 -2462
rect 5473 -2462 5500 -2438
rect 5567 -2460 5599 -2438
rect 5567 -2462 5569 -2460
rect 5597 -2462 5599 -2460
rect 5666 -2462 5693 -2438
rect 5473 -2476 5567 -2462
rect 5599 -2476 5693 -2462
rect 6053 -2462 6080 -2438
rect 6147 -2460 6179 -2438
rect 6147 -2462 6149 -2460
rect 6177 -2462 6179 -2460
rect 6246 -2462 6273 -2438
rect 6053 -2476 6147 -2462
rect 6179 -2476 6273 -2462
<< pdiff >>
rect -233 1798 -231 1800
rect -203 1798 -201 1800
rect -233 1776 -201 1798
rect -280 1748 -271 1776
rect -241 1748 -193 1776
rect -163 1748 -154 1776
tri -154 1748 -142 1760 sw
rect 347 1798 349 1800
rect 377 1798 379 1800
rect 347 1776 379 1798
rect 300 1748 309 1776
rect 339 1748 387 1776
rect 417 1748 426 1776
tri 426 1748 438 1760 sw
rect 927 1798 929 1800
rect 957 1798 959 1800
rect 927 1776 959 1798
rect 880 1748 889 1776
rect 919 1748 967 1776
rect 997 1748 1006 1776
tri 1006 1748 1018 1760 sw
rect 1507 1798 1509 1800
rect 1537 1798 1539 1800
rect 1507 1776 1539 1798
rect 1460 1748 1469 1776
rect 1499 1748 1547 1776
rect 1577 1748 1586 1776
tri 1586 1748 1598 1760 sw
rect 2087 1798 2089 1800
rect 2117 1798 2119 1800
rect 2087 1776 2119 1798
rect 2040 1748 2049 1776
rect 2079 1748 2127 1776
rect 2157 1748 2166 1776
tri 2166 1748 2178 1760 sw
rect 2667 1798 2669 1800
rect 2697 1798 2699 1800
rect 2667 1776 2699 1798
rect 2620 1748 2629 1776
rect 2659 1748 2707 1776
rect 2737 1748 2746 1776
tri 2746 1748 2758 1760 sw
rect 3247 1798 3249 1800
rect 3277 1798 3279 1800
rect 3247 1776 3279 1798
rect 3200 1748 3209 1776
rect 3239 1748 3287 1776
rect 3317 1748 3326 1776
tri 3326 1748 3338 1760 sw
rect 3827 1798 3829 1800
rect 3857 1798 3859 1800
rect 3827 1776 3859 1798
rect 3780 1748 3789 1776
rect 3819 1748 3867 1776
rect 3897 1748 3906 1776
tri 3906 1748 3918 1760 sw
rect 4407 1798 4409 1800
rect 4437 1798 4439 1800
rect 4407 1776 4439 1798
rect 4360 1748 4369 1776
rect 4399 1748 4447 1776
rect 4477 1748 4486 1776
tri 4486 1748 4498 1760 sw
rect 4987 1798 4989 1800
rect 5017 1798 5019 1800
rect 4987 1776 5019 1798
rect 4940 1748 4949 1776
rect 4979 1748 5027 1776
rect 5057 1748 5066 1776
tri 5066 1748 5078 1760 sw
rect 5567 1798 5569 1800
rect 5597 1798 5599 1800
rect 5567 1776 5599 1798
rect 5520 1748 5529 1776
rect 5559 1748 5607 1776
rect 5637 1748 5646 1776
tri 5646 1748 5658 1760 sw
rect 6147 1798 6149 1800
rect 6177 1798 6179 1800
rect 6147 1776 6179 1798
rect 6100 1748 6109 1776
rect 6139 1748 6187 1776
rect 6217 1748 6226 1776
tri 6226 1748 6238 1760 sw
rect -233 1528 -231 1530
rect -203 1528 -201 1530
rect -233 1506 -201 1528
rect -280 1478 -271 1506
rect -241 1478 -193 1506
rect -163 1478 -154 1506
tri -154 1478 -142 1490 sw
rect 347 1528 349 1530
rect 377 1528 379 1530
rect 347 1506 379 1528
rect 300 1478 309 1506
rect 339 1478 387 1506
rect 417 1478 426 1506
tri 426 1478 438 1490 sw
rect 927 1528 929 1530
rect 957 1528 959 1530
rect 927 1506 959 1528
rect 880 1478 889 1506
rect 919 1478 967 1506
rect 997 1478 1006 1506
tri 1006 1478 1018 1490 sw
rect 1507 1528 1509 1530
rect 1537 1528 1539 1530
rect 1507 1506 1539 1528
rect 1460 1478 1469 1506
rect 1499 1478 1547 1506
rect 1577 1478 1586 1506
tri 1586 1478 1598 1490 sw
rect 2087 1528 2089 1530
rect 2117 1528 2119 1530
rect 2087 1506 2119 1528
rect 2040 1478 2049 1506
rect 2079 1478 2127 1506
rect 2157 1478 2166 1506
tri 2166 1478 2178 1490 sw
rect 2667 1528 2669 1530
rect 2697 1528 2699 1530
rect 2667 1506 2699 1528
rect 2620 1478 2629 1506
rect 2659 1478 2707 1506
rect 2737 1478 2746 1506
tri 2746 1478 2758 1490 sw
rect 3247 1528 3249 1530
rect 3277 1528 3279 1530
rect 3247 1506 3279 1528
rect 3200 1478 3209 1506
rect 3239 1478 3287 1506
rect 3317 1478 3326 1506
tri 3326 1478 3338 1490 sw
rect 3827 1528 3829 1530
rect 3857 1528 3859 1530
rect 3827 1506 3859 1528
rect 3780 1478 3789 1506
rect 3819 1478 3867 1506
rect 3897 1478 3906 1506
tri 3906 1478 3918 1490 sw
rect 4407 1528 4409 1530
rect 4437 1528 4439 1530
rect 4407 1506 4439 1528
rect 4360 1478 4369 1506
rect 4399 1478 4447 1506
rect 4477 1478 4486 1506
tri 4486 1478 4498 1490 sw
rect 4987 1528 4989 1530
rect 5017 1528 5019 1530
rect 4987 1506 5019 1528
rect 4940 1478 4949 1506
rect 4979 1478 5027 1506
rect 5057 1478 5066 1506
tri 5066 1478 5078 1490 sw
rect 5567 1528 5569 1530
rect 5597 1528 5599 1530
rect 5567 1506 5599 1528
rect 5520 1478 5529 1506
rect 5559 1478 5607 1506
rect 5637 1478 5646 1506
tri 5646 1478 5658 1490 sw
rect 6147 1528 6149 1530
rect 6177 1528 6179 1530
rect 6147 1506 6179 1528
rect 6100 1478 6109 1506
rect 6139 1478 6187 1506
rect 6217 1478 6226 1506
tri 6226 1478 6238 1490 sw
rect -233 1258 -231 1260
rect -203 1258 -201 1260
rect -233 1236 -201 1258
rect -280 1208 -271 1236
rect -241 1208 -193 1236
rect -163 1208 -154 1236
tri -154 1208 -142 1220 sw
rect 347 1258 349 1260
rect 377 1258 379 1260
rect 347 1236 379 1258
rect 300 1208 309 1236
rect 339 1208 387 1236
rect 417 1208 426 1236
tri 426 1208 438 1220 sw
rect 927 1258 929 1260
rect 957 1258 959 1260
rect 927 1236 959 1258
rect 880 1208 889 1236
rect 919 1208 967 1236
rect 997 1208 1006 1236
tri 1006 1208 1018 1220 sw
rect 1507 1258 1509 1260
rect 1537 1258 1539 1260
rect 1507 1236 1539 1258
rect 1460 1208 1469 1236
rect 1499 1208 1547 1236
rect 1577 1208 1586 1236
tri 1586 1208 1598 1220 sw
rect 2087 1258 2089 1260
rect 2117 1258 2119 1260
rect 2087 1236 2119 1258
rect 2040 1208 2049 1236
rect 2079 1208 2127 1236
rect 2157 1208 2166 1236
tri 2166 1208 2178 1220 sw
rect 2667 1258 2669 1260
rect 2697 1258 2699 1260
rect 2667 1236 2699 1258
rect 2620 1208 2629 1236
rect 2659 1208 2707 1236
rect 2737 1208 2746 1236
tri 2746 1208 2758 1220 sw
rect 3247 1258 3249 1260
rect 3277 1258 3279 1260
rect 3247 1236 3279 1258
rect 3200 1208 3209 1236
rect 3239 1208 3287 1236
rect 3317 1208 3326 1236
tri 3326 1208 3338 1220 sw
rect 3827 1258 3829 1260
rect 3857 1258 3859 1260
rect 3827 1236 3859 1258
rect 3780 1208 3789 1236
rect 3819 1208 3867 1236
rect 3897 1208 3906 1236
tri 3906 1208 3918 1220 sw
rect 4407 1258 4409 1260
rect 4437 1258 4439 1260
rect 4407 1236 4439 1258
rect 4360 1208 4369 1236
rect 4399 1208 4447 1236
rect 4477 1208 4486 1236
tri 4486 1208 4498 1220 sw
rect 4987 1258 4989 1260
rect 5017 1258 5019 1260
rect 4987 1236 5019 1258
rect 4940 1208 4949 1236
rect 4979 1208 5027 1236
rect 5057 1208 5066 1236
tri 5066 1208 5078 1220 sw
rect 5567 1258 5569 1260
rect 5597 1258 5599 1260
rect 5567 1236 5599 1258
rect 5520 1208 5529 1236
rect 5559 1208 5607 1236
rect 5637 1208 5646 1236
tri 5646 1208 5658 1220 sw
rect 6147 1258 6149 1260
rect 6177 1258 6179 1260
rect 6147 1236 6179 1258
rect 6100 1208 6109 1236
rect 6139 1208 6187 1236
rect 6217 1208 6226 1236
tri 6226 1208 6238 1220 sw
rect -233 988 -231 990
rect -203 988 -201 990
rect -233 966 -201 988
rect -280 938 -271 966
rect -241 938 -193 966
rect -163 938 -154 966
tri -154 938 -142 950 sw
rect 347 988 349 990
rect 377 988 379 990
rect 347 966 379 988
rect 300 938 309 966
rect 339 938 387 966
rect 417 938 426 966
tri 426 938 438 950 sw
rect 927 988 929 990
rect 957 988 959 990
rect 927 966 959 988
rect 880 938 889 966
rect 919 938 967 966
rect 997 938 1006 966
tri 1006 938 1018 950 sw
rect 1507 988 1509 990
rect 1537 988 1539 990
rect 1507 966 1539 988
rect 1460 938 1469 966
rect 1499 938 1547 966
rect 1577 938 1586 966
tri 1586 938 1598 950 sw
rect 2087 988 2089 990
rect 2117 988 2119 990
rect 2087 966 2119 988
rect 2040 938 2049 966
rect 2079 938 2127 966
rect 2157 938 2166 966
tri 2166 938 2178 950 sw
rect 2667 988 2669 990
rect 2697 988 2699 990
rect 2667 966 2699 988
rect 2620 938 2629 966
rect 2659 938 2707 966
rect 2737 938 2746 966
tri 2746 938 2758 950 sw
rect 3247 988 3249 990
rect 3277 988 3279 990
rect 3247 966 3279 988
rect 3200 938 3209 966
rect 3239 938 3287 966
rect 3317 938 3326 966
tri 3326 938 3338 950 sw
rect 3827 988 3829 990
rect 3857 988 3859 990
rect 3827 966 3859 988
rect 3780 938 3789 966
rect 3819 938 3867 966
rect 3897 938 3906 966
tri 3906 938 3918 950 sw
rect 4407 988 4409 990
rect 4437 988 4439 990
rect 4407 966 4439 988
rect 4360 938 4369 966
rect 4399 938 4447 966
rect 4477 938 4486 966
tri 4486 938 4498 950 sw
rect 4987 988 4989 990
rect 5017 988 5019 990
rect 4987 966 5019 988
rect 4940 938 4949 966
rect 4979 938 5027 966
rect 5057 938 5066 966
tri 5066 938 5078 950 sw
rect 5567 988 5569 990
rect 5597 988 5599 990
rect 5567 966 5599 988
rect 5520 938 5529 966
rect 5559 938 5607 966
rect 5637 938 5646 966
tri 5646 938 5658 950 sw
rect 6147 988 6149 990
rect 6177 988 6179 990
rect 6147 966 6179 988
rect 6100 938 6109 966
rect 6139 938 6187 966
rect 6217 938 6226 966
tri 6226 938 6238 950 sw
rect -233 718 -231 720
rect -203 718 -201 720
rect -233 696 -201 718
rect -280 668 -271 696
rect -241 668 -193 696
rect -163 668 -154 696
tri -154 668 -142 680 sw
rect 347 718 349 720
rect 377 718 379 720
rect 347 696 379 718
rect 300 668 309 696
rect 339 668 387 696
rect 417 668 426 696
tri 426 668 438 680 sw
rect 927 718 929 720
rect 957 718 959 720
rect 927 696 959 718
rect 880 668 889 696
rect 919 668 967 696
rect 997 668 1006 696
tri 1006 668 1018 680 sw
rect 1507 718 1509 720
rect 1537 718 1539 720
rect 1507 696 1539 718
rect 1460 668 1469 696
rect 1499 668 1547 696
rect 1577 668 1586 696
tri 1586 668 1598 680 sw
rect 2087 718 2089 720
rect 2117 718 2119 720
rect 2087 696 2119 718
rect 2040 668 2049 696
rect 2079 668 2127 696
rect 2157 668 2166 696
tri 2166 668 2178 680 sw
rect 2667 718 2669 720
rect 2697 718 2699 720
rect 2667 696 2699 718
rect 2620 668 2629 696
rect 2659 668 2707 696
rect 2737 668 2746 696
tri 2746 668 2758 680 sw
rect 3247 718 3249 720
rect 3277 718 3279 720
rect 3247 696 3279 718
rect 3200 668 3209 696
rect 3239 668 3287 696
rect 3317 668 3326 696
tri 3326 668 3338 680 sw
rect 3827 718 3829 720
rect 3857 718 3859 720
rect 3827 696 3859 718
rect 3780 668 3789 696
rect 3819 668 3867 696
rect 3897 668 3906 696
tri 3906 668 3918 680 sw
rect 4407 718 4409 720
rect 4437 718 4439 720
rect 4407 696 4439 718
rect 4360 668 4369 696
rect 4399 668 4447 696
rect 4477 668 4486 696
tri 4486 668 4498 680 sw
rect 4987 718 4989 720
rect 5017 718 5019 720
rect 4987 696 5019 718
rect 4940 668 4949 696
rect 4979 668 5027 696
rect 5057 668 5066 696
tri 5066 668 5078 680 sw
rect 5567 718 5569 720
rect 5597 718 5599 720
rect 5567 696 5599 718
rect 5520 668 5529 696
rect 5559 668 5607 696
rect 5637 668 5646 696
tri 5646 668 5658 680 sw
rect 6147 718 6149 720
rect 6177 718 6179 720
rect 6147 696 6179 718
rect 6100 668 6109 696
rect 6139 668 6187 696
rect 6217 668 6226 696
tri 6226 668 6238 680 sw
rect -233 448 -231 450
rect -203 448 -201 450
rect -233 426 -201 448
rect -280 398 -271 426
rect -241 398 -193 426
rect -163 398 -154 426
tri -154 398 -142 410 sw
rect 347 448 349 450
rect 377 448 379 450
rect 347 426 379 448
rect 300 398 309 426
rect 339 398 387 426
rect 417 398 426 426
tri 426 398 438 410 sw
rect 927 448 929 450
rect 957 448 959 450
rect 927 426 959 448
rect 880 398 889 426
rect 919 398 967 426
rect 997 398 1006 426
tri 1006 398 1018 410 sw
rect 1507 448 1509 450
rect 1537 448 1539 450
rect 1507 426 1539 448
rect 1460 398 1469 426
rect 1499 398 1547 426
rect 1577 398 1586 426
tri 1586 398 1598 410 sw
rect 2087 448 2089 450
rect 2117 448 2119 450
rect 2087 426 2119 448
rect 2040 398 2049 426
rect 2079 398 2127 426
rect 2157 398 2166 426
tri 2166 398 2178 410 sw
rect 2667 448 2669 450
rect 2697 448 2699 450
rect 2667 426 2699 448
rect 2620 398 2629 426
rect 2659 398 2707 426
rect 2737 398 2746 426
tri 2746 398 2758 410 sw
rect 3247 448 3249 450
rect 3277 448 3279 450
rect 3247 426 3279 448
rect 3200 398 3209 426
rect 3239 398 3287 426
rect 3317 398 3326 426
tri 3326 398 3338 410 sw
rect 3827 448 3829 450
rect 3857 448 3859 450
rect 3827 426 3859 448
rect 3780 398 3789 426
rect 3819 398 3867 426
rect 3897 398 3906 426
tri 3906 398 3918 410 sw
rect 4407 448 4409 450
rect 4437 448 4439 450
rect 4407 426 4439 448
rect 4360 398 4369 426
rect 4399 398 4447 426
rect 4477 398 4486 426
tri 4486 398 4498 410 sw
rect 4987 448 4989 450
rect 5017 448 5019 450
rect 4987 426 5019 448
rect 4940 398 4949 426
rect 4979 398 5027 426
rect 5057 398 5066 426
tri 5066 398 5078 410 sw
rect 5567 448 5569 450
rect 5597 448 5599 450
rect 5567 426 5599 448
rect 5520 398 5529 426
rect 5559 398 5607 426
rect 5637 398 5646 426
tri 5646 398 5658 410 sw
rect 6147 448 6149 450
rect 6177 448 6179 450
rect 6147 426 6179 448
rect 6100 398 6109 426
rect 6139 398 6187 426
rect 6217 398 6226 426
tri 6226 398 6238 410 sw
rect -233 178 -231 180
rect -203 178 -201 180
rect -233 156 -201 178
rect -280 128 -271 156
rect -241 128 -193 156
rect -163 128 -154 156
tri -154 128 -142 140 sw
rect 347 178 349 180
rect 377 178 379 180
rect 347 156 379 178
rect 300 128 309 156
rect 339 128 387 156
rect 417 128 426 156
tri 426 128 438 140 sw
rect 927 178 929 180
rect 957 178 959 180
rect 927 156 959 178
rect 880 128 889 156
rect 919 128 967 156
rect 997 128 1006 156
tri 1006 128 1018 140 sw
rect 1507 178 1509 180
rect 1537 178 1539 180
rect 1507 156 1539 178
rect 1460 128 1469 156
rect 1499 128 1547 156
rect 1577 128 1586 156
tri 1586 128 1598 140 sw
rect 2087 178 2089 180
rect 2117 178 2119 180
rect 2087 156 2119 178
rect 2040 128 2049 156
rect 2079 128 2127 156
rect 2157 128 2166 156
tri 2166 128 2178 140 sw
rect 2667 178 2669 180
rect 2697 178 2699 180
rect 2667 156 2699 178
rect 2620 128 2629 156
rect 2659 128 2707 156
rect 2737 128 2746 156
tri 2746 128 2758 140 sw
rect 3247 178 3249 180
rect 3277 178 3279 180
rect 3247 156 3279 178
rect 3200 128 3209 156
rect 3239 128 3287 156
rect 3317 128 3326 156
tri 3326 128 3338 140 sw
rect 3827 178 3829 180
rect 3857 178 3859 180
rect 3827 156 3859 178
rect 3780 128 3789 156
rect 3819 128 3867 156
rect 3897 128 3906 156
tri 3906 128 3918 140 sw
rect 4407 178 4409 180
rect 4437 178 4439 180
rect 4407 156 4439 178
rect 4360 128 4369 156
rect 4399 128 4447 156
rect 4477 128 4486 156
tri 4486 128 4498 140 sw
rect 4987 178 4989 180
rect 5017 178 5019 180
rect 4987 156 5019 178
rect 4940 128 4949 156
rect 4979 128 5027 156
rect 5057 128 5066 156
tri 5066 128 5078 140 sw
rect 5567 178 5569 180
rect 5597 178 5599 180
rect 5567 156 5599 178
rect 5520 128 5529 156
rect 5559 128 5607 156
rect 5637 128 5646 156
tri 5646 128 5658 140 sw
rect 6147 178 6149 180
rect 6177 178 6179 180
rect 6147 156 6179 178
rect 6100 128 6109 156
rect 6139 128 6187 156
rect 6217 128 6226 156
tri 6226 128 6238 140 sw
rect -233 -92 -231 -90
rect -203 -92 -201 -90
rect -233 -114 -201 -92
rect -280 -142 -271 -114
rect -241 -142 -193 -114
rect -163 -142 -154 -114
tri -154 -142 -142 -130 sw
rect 347 -92 349 -90
rect 377 -92 379 -90
rect 347 -114 379 -92
rect 300 -142 309 -114
rect 339 -142 387 -114
rect 417 -142 426 -114
tri 426 -142 438 -130 sw
rect 927 -92 929 -90
rect 957 -92 959 -90
rect 927 -114 959 -92
rect 880 -142 889 -114
rect 919 -142 967 -114
rect 997 -142 1006 -114
tri 1006 -142 1018 -130 sw
rect 1507 -92 1509 -90
rect 1537 -92 1539 -90
rect 1507 -114 1539 -92
rect 1460 -142 1469 -114
rect 1499 -142 1547 -114
rect 1577 -142 1586 -114
tri 1586 -142 1598 -130 sw
rect 2087 -92 2089 -90
rect 2117 -92 2119 -90
rect 2087 -114 2119 -92
rect 2040 -142 2049 -114
rect 2079 -142 2127 -114
rect 2157 -142 2166 -114
tri 2166 -142 2178 -130 sw
rect 2667 -92 2669 -90
rect 2697 -92 2699 -90
rect 2667 -114 2699 -92
rect 2620 -142 2629 -114
rect 2659 -142 2707 -114
rect 2737 -142 2746 -114
tri 2746 -142 2758 -130 sw
rect 3247 -92 3249 -90
rect 3277 -92 3279 -90
rect 3247 -114 3279 -92
rect 3200 -142 3209 -114
rect 3239 -142 3287 -114
rect 3317 -142 3326 -114
tri 3326 -142 3338 -130 sw
rect 3827 -92 3829 -90
rect 3857 -92 3859 -90
rect 3827 -114 3859 -92
rect 3780 -142 3789 -114
rect 3819 -142 3867 -114
rect 3897 -142 3906 -114
tri 3906 -142 3918 -130 sw
rect 4407 -92 4409 -90
rect 4437 -92 4439 -90
rect 4407 -114 4439 -92
rect 4360 -142 4369 -114
rect 4399 -142 4447 -114
rect 4477 -142 4486 -114
tri 4486 -142 4498 -130 sw
rect 4987 -92 4989 -90
rect 5017 -92 5019 -90
rect 4987 -114 5019 -92
rect 4940 -142 4949 -114
rect 4979 -142 5027 -114
rect 5057 -142 5066 -114
tri 5066 -142 5078 -130 sw
rect 5567 -92 5569 -90
rect 5597 -92 5599 -90
rect 5567 -114 5599 -92
rect 5520 -142 5529 -114
rect 5559 -142 5607 -114
rect 5637 -142 5646 -114
tri 5646 -142 5658 -130 sw
rect 6147 -92 6149 -90
rect 6177 -92 6179 -90
rect 6147 -114 6179 -92
rect 6100 -142 6109 -114
rect 6139 -142 6187 -114
rect 6217 -142 6226 -114
tri 6226 -142 6238 -130 sw
rect -233 -362 -231 -360
rect -203 -362 -201 -360
rect -233 -384 -201 -362
rect -280 -412 -271 -384
rect -241 -412 -193 -384
rect -163 -412 -154 -384
tri -154 -412 -142 -400 sw
rect 347 -362 349 -360
rect 377 -362 379 -360
rect 347 -384 379 -362
rect 300 -412 309 -384
rect 339 -412 387 -384
rect 417 -412 426 -384
tri 426 -412 438 -400 sw
rect 927 -362 929 -360
rect 957 -362 959 -360
rect 927 -384 959 -362
rect 880 -412 889 -384
rect 919 -412 967 -384
rect 997 -412 1006 -384
tri 1006 -412 1018 -400 sw
rect 1507 -362 1509 -360
rect 1537 -362 1539 -360
rect 1507 -384 1539 -362
rect 1460 -412 1469 -384
rect 1499 -412 1547 -384
rect 1577 -412 1586 -384
tri 1586 -412 1598 -400 sw
rect 2087 -362 2089 -360
rect 2117 -362 2119 -360
rect 2087 -384 2119 -362
rect 2040 -412 2049 -384
rect 2079 -412 2127 -384
rect 2157 -412 2166 -384
tri 2166 -412 2178 -400 sw
rect 2667 -362 2669 -360
rect 2697 -362 2699 -360
rect 2667 -384 2699 -362
rect 2620 -412 2629 -384
rect 2659 -412 2707 -384
rect 2737 -412 2746 -384
tri 2746 -412 2758 -400 sw
rect 3247 -362 3249 -360
rect 3277 -362 3279 -360
rect 3247 -384 3279 -362
rect 3200 -412 3209 -384
rect 3239 -412 3287 -384
rect 3317 -412 3326 -384
tri 3326 -412 3338 -400 sw
rect 3827 -362 3829 -360
rect 3857 -362 3859 -360
rect 3827 -384 3859 -362
rect 3780 -412 3789 -384
rect 3819 -412 3867 -384
rect 3897 -412 3906 -384
tri 3906 -412 3918 -400 sw
rect 4407 -362 4409 -360
rect 4437 -362 4439 -360
rect 4407 -384 4439 -362
rect 4360 -412 4369 -384
rect 4399 -412 4447 -384
rect 4477 -412 4486 -384
tri 4486 -412 4498 -400 sw
rect 4987 -362 4989 -360
rect 5017 -362 5019 -360
rect 4987 -384 5019 -362
rect 4940 -412 4949 -384
rect 4979 -412 5027 -384
rect 5057 -412 5066 -384
tri 5066 -412 5078 -400 sw
rect 5567 -362 5569 -360
rect 5597 -362 5599 -360
rect 5567 -384 5599 -362
rect 5520 -412 5529 -384
rect 5559 -412 5607 -384
rect 5637 -412 5646 -384
tri 5646 -412 5658 -400 sw
rect 6147 -362 6149 -360
rect 6177 -362 6179 -360
rect 6147 -384 6179 -362
rect 6100 -412 6109 -384
rect 6139 -412 6187 -384
rect 6217 -412 6226 -384
tri 6226 -412 6238 -400 sw
rect -233 -632 -231 -630
rect -203 -632 -201 -630
rect -233 -654 -201 -632
rect -280 -682 -271 -654
rect -241 -682 -193 -654
rect -163 -682 -154 -654
tri -154 -682 -142 -670 sw
rect 347 -632 349 -630
rect 377 -632 379 -630
rect 347 -654 379 -632
rect 300 -682 309 -654
rect 339 -682 387 -654
rect 417 -682 426 -654
tri 426 -682 438 -670 sw
rect 927 -632 929 -630
rect 957 -632 959 -630
rect 927 -654 959 -632
rect 880 -682 889 -654
rect 919 -682 967 -654
rect 997 -682 1006 -654
tri 1006 -682 1018 -670 sw
rect 1507 -632 1509 -630
rect 1537 -632 1539 -630
rect 1507 -654 1539 -632
rect 1460 -682 1469 -654
rect 1499 -682 1547 -654
rect 1577 -682 1586 -654
tri 1586 -682 1598 -670 sw
rect 2087 -632 2089 -630
rect 2117 -632 2119 -630
rect 2087 -654 2119 -632
rect 2040 -682 2049 -654
rect 2079 -682 2127 -654
rect 2157 -682 2166 -654
tri 2166 -682 2178 -670 sw
rect 2667 -632 2669 -630
rect 2697 -632 2699 -630
rect 2667 -654 2699 -632
rect 2620 -682 2629 -654
rect 2659 -682 2707 -654
rect 2737 -682 2746 -654
tri 2746 -682 2758 -670 sw
rect 3247 -632 3249 -630
rect 3277 -632 3279 -630
rect 3247 -654 3279 -632
rect 3200 -682 3209 -654
rect 3239 -682 3287 -654
rect 3317 -682 3326 -654
tri 3326 -682 3338 -670 sw
rect 3827 -632 3829 -630
rect 3857 -632 3859 -630
rect 3827 -654 3859 -632
rect 3780 -682 3789 -654
rect 3819 -682 3867 -654
rect 3897 -682 3906 -654
tri 3906 -682 3918 -670 sw
rect 4407 -632 4409 -630
rect 4437 -632 4439 -630
rect 4407 -654 4439 -632
rect 4360 -682 4369 -654
rect 4399 -682 4447 -654
rect 4477 -682 4486 -654
tri 4486 -682 4498 -670 sw
rect 4987 -632 4989 -630
rect 5017 -632 5019 -630
rect 4987 -654 5019 -632
rect 4940 -682 4949 -654
rect 4979 -682 5027 -654
rect 5057 -682 5066 -654
tri 5066 -682 5078 -670 sw
rect 5567 -632 5569 -630
rect 5597 -632 5599 -630
rect 5567 -654 5599 -632
rect 5520 -682 5529 -654
rect 5559 -682 5607 -654
rect 5637 -682 5646 -654
tri 5646 -682 5658 -670 sw
rect 6147 -632 6149 -630
rect 6177 -632 6179 -630
rect 6147 -654 6179 -632
rect 6100 -682 6109 -654
rect 6139 -682 6187 -654
rect 6217 -682 6226 -654
tri 6226 -682 6238 -670 sw
rect -233 -902 -231 -900
rect -203 -902 -201 -900
rect -233 -924 -201 -902
rect -280 -952 -271 -924
rect -241 -952 -193 -924
rect -163 -952 -154 -924
tri -154 -952 -142 -940 sw
rect 347 -902 349 -900
rect 377 -902 379 -900
rect 347 -924 379 -902
rect 300 -952 309 -924
rect 339 -952 387 -924
rect 417 -952 426 -924
tri 426 -952 438 -940 sw
rect 927 -902 929 -900
rect 957 -902 959 -900
rect 927 -924 959 -902
rect 880 -952 889 -924
rect 919 -952 967 -924
rect 997 -952 1006 -924
tri 1006 -952 1018 -940 sw
rect 1507 -902 1509 -900
rect 1537 -902 1539 -900
rect 1507 -924 1539 -902
rect 1460 -952 1469 -924
rect 1499 -952 1547 -924
rect 1577 -952 1586 -924
tri 1586 -952 1598 -940 sw
rect 2087 -902 2089 -900
rect 2117 -902 2119 -900
rect 2087 -924 2119 -902
rect 2040 -952 2049 -924
rect 2079 -952 2127 -924
rect 2157 -952 2166 -924
tri 2166 -952 2178 -940 sw
rect 2667 -902 2669 -900
rect 2697 -902 2699 -900
rect 2667 -924 2699 -902
rect 2620 -952 2629 -924
rect 2659 -952 2707 -924
rect 2737 -952 2746 -924
tri 2746 -952 2758 -940 sw
rect 3247 -902 3249 -900
rect 3277 -902 3279 -900
rect 3247 -924 3279 -902
rect 3200 -952 3209 -924
rect 3239 -952 3287 -924
rect 3317 -952 3326 -924
tri 3326 -952 3338 -940 sw
rect 3827 -902 3829 -900
rect 3857 -902 3859 -900
rect 3827 -924 3859 -902
rect 3780 -952 3789 -924
rect 3819 -952 3867 -924
rect 3897 -952 3906 -924
tri 3906 -952 3918 -940 sw
rect 4407 -902 4409 -900
rect 4437 -902 4439 -900
rect 4407 -924 4439 -902
rect 4360 -952 4369 -924
rect 4399 -952 4447 -924
rect 4477 -952 4486 -924
tri 4486 -952 4498 -940 sw
rect 4987 -902 4989 -900
rect 5017 -902 5019 -900
rect 4987 -924 5019 -902
rect 4940 -952 4949 -924
rect 4979 -952 5027 -924
rect 5057 -952 5066 -924
tri 5066 -952 5078 -940 sw
rect 5567 -902 5569 -900
rect 5597 -902 5599 -900
rect 5567 -924 5599 -902
rect 5520 -952 5529 -924
rect 5559 -952 5607 -924
rect 5637 -952 5646 -924
tri 5646 -952 5658 -940 sw
rect 6147 -902 6149 -900
rect 6177 -902 6179 -900
rect 6147 -924 6179 -902
rect 6100 -952 6109 -924
rect 6139 -952 6187 -924
rect 6217 -952 6226 -924
tri 6226 -952 6238 -940 sw
rect -233 -1172 -231 -1170
rect -203 -1172 -201 -1170
rect -233 -1194 -201 -1172
rect -280 -1222 -271 -1194
rect -241 -1222 -193 -1194
rect -163 -1222 -154 -1194
tri -154 -1222 -142 -1210 sw
rect 347 -1172 349 -1170
rect 377 -1172 379 -1170
rect 347 -1194 379 -1172
rect 300 -1222 309 -1194
rect 339 -1222 387 -1194
rect 417 -1222 426 -1194
tri 426 -1222 438 -1210 sw
rect 927 -1172 929 -1170
rect 957 -1172 959 -1170
rect 927 -1194 959 -1172
rect 880 -1222 889 -1194
rect 919 -1222 967 -1194
rect 997 -1222 1006 -1194
tri 1006 -1222 1018 -1210 sw
rect 1507 -1172 1509 -1170
rect 1537 -1172 1539 -1170
rect 1507 -1194 1539 -1172
rect 1460 -1222 1469 -1194
rect 1499 -1222 1547 -1194
rect 1577 -1222 1586 -1194
tri 1586 -1222 1598 -1210 sw
rect 2087 -1172 2089 -1170
rect 2117 -1172 2119 -1170
rect 2087 -1194 2119 -1172
rect 2040 -1222 2049 -1194
rect 2079 -1222 2127 -1194
rect 2157 -1222 2166 -1194
tri 2166 -1222 2178 -1210 sw
rect 2667 -1172 2669 -1170
rect 2697 -1172 2699 -1170
rect 2667 -1194 2699 -1172
rect 2620 -1222 2629 -1194
rect 2659 -1222 2707 -1194
rect 2737 -1222 2746 -1194
tri 2746 -1222 2758 -1210 sw
rect 3247 -1172 3249 -1170
rect 3277 -1172 3279 -1170
rect 3247 -1194 3279 -1172
rect 3200 -1222 3209 -1194
rect 3239 -1222 3287 -1194
rect 3317 -1222 3326 -1194
tri 3326 -1222 3338 -1210 sw
rect 3827 -1172 3829 -1170
rect 3857 -1172 3859 -1170
rect 3827 -1194 3859 -1172
rect 3780 -1222 3789 -1194
rect 3819 -1222 3867 -1194
rect 3897 -1222 3906 -1194
tri 3906 -1222 3918 -1210 sw
rect 4407 -1172 4409 -1170
rect 4437 -1172 4439 -1170
rect 4407 -1194 4439 -1172
rect 4360 -1222 4369 -1194
rect 4399 -1222 4447 -1194
rect 4477 -1222 4486 -1194
tri 4486 -1222 4498 -1210 sw
rect 4987 -1172 4989 -1170
rect 5017 -1172 5019 -1170
rect 4987 -1194 5019 -1172
rect 4940 -1222 4949 -1194
rect 4979 -1222 5027 -1194
rect 5057 -1222 5066 -1194
tri 5066 -1222 5078 -1210 sw
rect 5567 -1172 5569 -1170
rect 5597 -1172 5599 -1170
rect 5567 -1194 5599 -1172
rect 5520 -1222 5529 -1194
rect 5559 -1222 5607 -1194
rect 5637 -1222 5646 -1194
tri 5646 -1222 5658 -1210 sw
rect 6147 -1172 6149 -1170
rect 6177 -1172 6179 -1170
rect 6147 -1194 6179 -1172
rect 6100 -1222 6109 -1194
rect 6139 -1222 6187 -1194
rect 6217 -1222 6226 -1194
tri 6226 -1222 6238 -1210 sw
rect -233 -1442 -231 -1440
rect -203 -1442 -201 -1440
rect -233 -1464 -201 -1442
rect -280 -1492 -271 -1464
rect -241 -1492 -193 -1464
rect -163 -1492 -154 -1464
tri -154 -1492 -142 -1480 sw
rect 347 -1442 349 -1440
rect 377 -1442 379 -1440
rect 347 -1464 379 -1442
rect 300 -1492 309 -1464
rect 339 -1492 387 -1464
rect 417 -1492 426 -1464
tri 426 -1492 438 -1480 sw
rect 927 -1442 929 -1440
rect 957 -1442 959 -1440
rect 927 -1464 959 -1442
rect 880 -1492 889 -1464
rect 919 -1492 967 -1464
rect 997 -1492 1006 -1464
tri 1006 -1492 1018 -1480 sw
rect 1507 -1442 1509 -1440
rect 1537 -1442 1539 -1440
rect 1507 -1464 1539 -1442
rect 1460 -1492 1469 -1464
rect 1499 -1492 1547 -1464
rect 1577 -1492 1586 -1464
tri 1586 -1492 1598 -1480 sw
rect 2087 -1442 2089 -1440
rect 2117 -1442 2119 -1440
rect 2087 -1464 2119 -1442
rect 2040 -1492 2049 -1464
rect 2079 -1492 2127 -1464
rect 2157 -1492 2166 -1464
tri 2166 -1492 2178 -1480 sw
rect 2667 -1442 2669 -1440
rect 2697 -1442 2699 -1440
rect 2667 -1464 2699 -1442
rect 2620 -1492 2629 -1464
rect 2659 -1492 2707 -1464
rect 2737 -1492 2746 -1464
tri 2746 -1492 2758 -1480 sw
rect 3247 -1442 3249 -1440
rect 3277 -1442 3279 -1440
rect 3247 -1464 3279 -1442
rect 3200 -1492 3209 -1464
rect 3239 -1492 3287 -1464
rect 3317 -1492 3326 -1464
tri 3326 -1492 3338 -1480 sw
rect 3827 -1442 3829 -1440
rect 3857 -1442 3859 -1440
rect 3827 -1464 3859 -1442
rect 3780 -1492 3789 -1464
rect 3819 -1492 3867 -1464
rect 3897 -1492 3906 -1464
tri 3906 -1492 3918 -1480 sw
rect 4407 -1442 4409 -1440
rect 4437 -1442 4439 -1440
rect 4407 -1464 4439 -1442
rect 4360 -1492 4369 -1464
rect 4399 -1492 4447 -1464
rect 4477 -1492 4486 -1464
tri 4486 -1492 4498 -1480 sw
rect 4987 -1442 4989 -1440
rect 5017 -1442 5019 -1440
rect 4987 -1464 5019 -1442
rect 4940 -1492 4949 -1464
rect 4979 -1492 5027 -1464
rect 5057 -1492 5066 -1464
tri 5066 -1492 5078 -1480 sw
rect 5567 -1442 5569 -1440
rect 5597 -1442 5599 -1440
rect 5567 -1464 5599 -1442
rect 5520 -1492 5529 -1464
rect 5559 -1492 5607 -1464
rect 5637 -1492 5646 -1464
tri 5646 -1492 5658 -1480 sw
rect 6147 -1442 6149 -1440
rect 6177 -1442 6179 -1440
rect 6147 -1464 6179 -1442
rect 6100 -1492 6109 -1464
rect 6139 -1492 6187 -1464
rect 6217 -1492 6226 -1464
tri 6226 -1492 6238 -1480 sw
rect -233 -1712 -231 -1710
rect -203 -1712 -201 -1710
rect -233 -1734 -201 -1712
rect -280 -1762 -271 -1734
rect -241 -1762 -193 -1734
rect -163 -1762 -154 -1734
tri -154 -1762 -142 -1750 sw
rect 347 -1712 349 -1710
rect 377 -1712 379 -1710
rect 347 -1734 379 -1712
rect 300 -1762 309 -1734
rect 339 -1762 387 -1734
rect 417 -1762 426 -1734
tri 426 -1762 438 -1750 sw
rect 927 -1712 929 -1710
rect 957 -1712 959 -1710
rect 927 -1734 959 -1712
rect 880 -1762 889 -1734
rect 919 -1762 967 -1734
rect 997 -1762 1006 -1734
tri 1006 -1762 1018 -1750 sw
rect 1507 -1712 1509 -1710
rect 1537 -1712 1539 -1710
rect 1507 -1734 1539 -1712
rect 1460 -1762 1469 -1734
rect 1499 -1762 1547 -1734
rect 1577 -1762 1586 -1734
tri 1586 -1762 1598 -1750 sw
rect 2087 -1712 2089 -1710
rect 2117 -1712 2119 -1710
rect 2087 -1734 2119 -1712
rect 2040 -1762 2049 -1734
rect 2079 -1762 2127 -1734
rect 2157 -1762 2166 -1734
tri 2166 -1762 2178 -1750 sw
rect 2667 -1712 2669 -1710
rect 2697 -1712 2699 -1710
rect 2667 -1734 2699 -1712
rect 2620 -1762 2629 -1734
rect 2659 -1762 2707 -1734
rect 2737 -1762 2746 -1734
tri 2746 -1762 2758 -1750 sw
rect 3247 -1712 3249 -1710
rect 3277 -1712 3279 -1710
rect 3247 -1734 3279 -1712
rect 3200 -1762 3209 -1734
rect 3239 -1762 3287 -1734
rect 3317 -1762 3326 -1734
tri 3326 -1762 3338 -1750 sw
rect 3827 -1712 3829 -1710
rect 3857 -1712 3859 -1710
rect 3827 -1734 3859 -1712
rect 3780 -1762 3789 -1734
rect 3819 -1762 3867 -1734
rect 3897 -1762 3906 -1734
tri 3906 -1762 3918 -1750 sw
rect 4407 -1712 4409 -1710
rect 4437 -1712 4439 -1710
rect 4407 -1734 4439 -1712
rect 4360 -1762 4369 -1734
rect 4399 -1762 4447 -1734
rect 4477 -1762 4486 -1734
tri 4486 -1762 4498 -1750 sw
rect 4987 -1712 4989 -1710
rect 5017 -1712 5019 -1710
rect 4987 -1734 5019 -1712
rect 4940 -1762 4949 -1734
rect 4979 -1762 5027 -1734
rect 5057 -1762 5066 -1734
tri 5066 -1762 5078 -1750 sw
rect 5567 -1712 5569 -1710
rect 5597 -1712 5599 -1710
rect 5567 -1734 5599 -1712
rect 5520 -1762 5529 -1734
rect 5559 -1762 5607 -1734
rect 5637 -1762 5646 -1734
tri 5646 -1762 5658 -1750 sw
rect 6147 -1712 6149 -1710
rect 6177 -1712 6179 -1710
rect 6147 -1734 6179 -1712
rect 6100 -1762 6109 -1734
rect 6139 -1762 6187 -1734
rect 6217 -1762 6226 -1734
tri 6226 -1762 6238 -1750 sw
rect -233 -1982 -231 -1980
rect -203 -1982 -201 -1980
rect -233 -2004 -201 -1982
rect -280 -2032 -271 -2004
rect -241 -2032 -193 -2004
rect -163 -2032 -154 -2004
tri -154 -2032 -142 -2020 sw
rect 347 -1982 349 -1980
rect 377 -1982 379 -1980
rect 347 -2004 379 -1982
rect 300 -2032 309 -2004
rect 339 -2032 387 -2004
rect 417 -2032 426 -2004
tri 426 -2032 438 -2020 sw
rect 927 -1982 929 -1980
rect 957 -1982 959 -1980
rect 927 -2004 959 -1982
rect 880 -2032 889 -2004
rect 919 -2032 967 -2004
rect 997 -2032 1006 -2004
tri 1006 -2032 1018 -2020 sw
rect 1507 -1982 1509 -1980
rect 1537 -1982 1539 -1980
rect 1507 -2004 1539 -1982
rect 1460 -2032 1469 -2004
rect 1499 -2032 1547 -2004
rect 1577 -2032 1586 -2004
tri 1586 -2032 1598 -2020 sw
rect 2087 -1982 2089 -1980
rect 2117 -1982 2119 -1980
rect 2087 -2004 2119 -1982
rect 2040 -2032 2049 -2004
rect 2079 -2032 2127 -2004
rect 2157 -2032 2166 -2004
tri 2166 -2032 2178 -2020 sw
rect 2667 -1982 2669 -1980
rect 2697 -1982 2699 -1980
rect 2667 -2004 2699 -1982
rect 2620 -2032 2629 -2004
rect 2659 -2032 2707 -2004
rect 2737 -2032 2746 -2004
tri 2746 -2032 2758 -2020 sw
rect 3247 -1982 3249 -1980
rect 3277 -1982 3279 -1980
rect 3247 -2004 3279 -1982
rect 3200 -2032 3209 -2004
rect 3239 -2032 3287 -2004
rect 3317 -2032 3326 -2004
tri 3326 -2032 3338 -2020 sw
rect 3827 -1982 3829 -1980
rect 3857 -1982 3859 -1980
rect 3827 -2004 3859 -1982
rect 3780 -2032 3789 -2004
rect 3819 -2032 3867 -2004
rect 3897 -2032 3906 -2004
tri 3906 -2032 3918 -2020 sw
rect 4407 -1982 4409 -1980
rect 4437 -1982 4439 -1980
rect 4407 -2004 4439 -1982
rect 4360 -2032 4369 -2004
rect 4399 -2032 4447 -2004
rect 4477 -2032 4486 -2004
tri 4486 -2032 4498 -2020 sw
rect 4987 -1982 4989 -1980
rect 5017 -1982 5019 -1980
rect 4987 -2004 5019 -1982
rect 4940 -2032 4949 -2004
rect 4979 -2032 5027 -2004
rect 5057 -2032 5066 -2004
tri 5066 -2032 5078 -2020 sw
rect 5567 -1982 5569 -1980
rect 5597 -1982 5599 -1980
rect 5567 -2004 5599 -1982
rect 5520 -2032 5529 -2004
rect 5559 -2032 5607 -2004
rect 5637 -2032 5646 -2004
tri 5646 -2032 5658 -2020 sw
rect 6147 -1982 6149 -1980
rect 6177 -1982 6179 -1980
rect 6147 -2004 6179 -1982
rect 6100 -2032 6109 -2004
rect 6139 -2032 6187 -2004
rect 6217 -2032 6226 -2004
tri 6226 -2032 6238 -2020 sw
rect -233 -2252 -231 -2250
rect -203 -2252 -201 -2250
rect -233 -2274 -201 -2252
rect -280 -2302 -271 -2274
rect -241 -2302 -193 -2274
rect -163 -2302 -154 -2274
tri -154 -2302 -142 -2290 sw
rect 347 -2252 349 -2250
rect 377 -2252 379 -2250
rect 347 -2274 379 -2252
rect 300 -2302 309 -2274
rect 339 -2302 387 -2274
rect 417 -2302 426 -2274
tri 426 -2302 438 -2290 sw
rect 927 -2252 929 -2250
rect 957 -2252 959 -2250
rect 927 -2274 959 -2252
rect 880 -2302 889 -2274
rect 919 -2302 967 -2274
rect 997 -2302 1006 -2274
tri 1006 -2302 1018 -2290 sw
rect 1507 -2252 1509 -2250
rect 1537 -2252 1539 -2250
rect 1507 -2274 1539 -2252
rect 1460 -2302 1469 -2274
rect 1499 -2302 1547 -2274
rect 1577 -2302 1586 -2274
tri 1586 -2302 1598 -2290 sw
rect 2087 -2252 2089 -2250
rect 2117 -2252 2119 -2250
rect 2087 -2274 2119 -2252
rect 2040 -2302 2049 -2274
rect 2079 -2302 2127 -2274
rect 2157 -2302 2166 -2274
tri 2166 -2302 2178 -2290 sw
rect 2667 -2252 2669 -2250
rect 2697 -2252 2699 -2250
rect 2667 -2274 2699 -2252
rect 2620 -2302 2629 -2274
rect 2659 -2302 2707 -2274
rect 2737 -2302 2746 -2274
tri 2746 -2302 2758 -2290 sw
rect 3247 -2252 3249 -2250
rect 3277 -2252 3279 -2250
rect 3247 -2274 3279 -2252
rect 3200 -2302 3209 -2274
rect 3239 -2302 3287 -2274
rect 3317 -2302 3326 -2274
tri 3326 -2302 3338 -2290 sw
rect 3827 -2252 3829 -2250
rect 3857 -2252 3859 -2250
rect 3827 -2274 3859 -2252
rect 3780 -2302 3789 -2274
rect 3819 -2302 3867 -2274
rect 3897 -2302 3906 -2274
tri 3906 -2302 3918 -2290 sw
rect 4407 -2252 4409 -2250
rect 4437 -2252 4439 -2250
rect 4407 -2274 4439 -2252
rect 4360 -2302 4369 -2274
rect 4399 -2302 4447 -2274
rect 4477 -2302 4486 -2274
tri 4486 -2302 4498 -2290 sw
rect 4987 -2252 4989 -2250
rect 5017 -2252 5019 -2250
rect 4987 -2274 5019 -2252
rect 4940 -2302 4949 -2274
rect 4979 -2302 5027 -2274
rect 5057 -2302 5066 -2274
tri 5066 -2302 5078 -2290 sw
rect 5567 -2252 5569 -2250
rect 5597 -2252 5599 -2250
rect 5567 -2274 5599 -2252
rect 5520 -2302 5529 -2274
rect 5559 -2302 5607 -2274
rect 5637 -2302 5646 -2274
tri 5646 -2302 5658 -2290 sw
rect 6147 -2252 6149 -2250
rect 6177 -2252 6179 -2250
rect 6147 -2274 6179 -2252
rect 6100 -2302 6109 -2274
rect 6139 -2302 6187 -2274
rect 6217 -2302 6226 -2274
tri 6226 -2302 6238 -2290 sw
<< ndiffc >>
rect -419 1758 -404 1786
rect -338 1758 -323 1786
rect -111 1758 -96 1786
rect -29 1758 -14 1787
rect 161 1758 176 1786
rect 242 1758 257 1786
rect 469 1758 484 1786
rect 551 1758 566 1787
rect 741 1758 756 1786
rect 822 1758 837 1786
rect 1049 1758 1064 1786
rect 1131 1758 1146 1787
rect 1321 1758 1336 1786
rect 1402 1758 1417 1786
rect 1629 1758 1644 1786
rect 1711 1758 1726 1787
rect 1901 1758 1916 1786
rect 1982 1758 1997 1786
rect 2209 1758 2224 1786
rect 2291 1758 2306 1787
rect 2481 1758 2496 1786
rect 2562 1758 2577 1786
rect 2789 1758 2804 1786
rect 2871 1758 2886 1787
rect 3061 1758 3076 1786
rect 3142 1758 3157 1786
rect 3369 1758 3384 1786
rect 3451 1758 3466 1787
rect 3641 1758 3656 1786
rect 3722 1758 3737 1786
rect 3949 1758 3964 1786
rect 4031 1758 4046 1787
rect 4221 1758 4236 1786
rect 4302 1758 4317 1786
rect 4529 1758 4544 1786
rect 4611 1758 4626 1787
rect 4801 1758 4816 1786
rect 4882 1758 4897 1786
rect 5109 1758 5124 1786
rect 5191 1758 5206 1787
rect 5381 1758 5396 1786
rect 5462 1758 5477 1786
rect 5689 1758 5704 1786
rect 5771 1758 5786 1787
rect 5961 1758 5976 1786
rect 6042 1758 6057 1786
rect 6269 1758 6284 1786
rect 6351 1758 6366 1787
rect -493 1612 -478 1654
rect -296 1637 -286 1644
tri -286 1637 -279 1644 sw
rect -296 1612 -279 1637
rect -155 1612 -138 1644
rect 44 1612 59 1654
rect 87 1612 102 1654
rect 284 1637 294 1644
tri 294 1637 301 1644 sw
rect 284 1612 301 1637
rect 425 1612 442 1644
rect 624 1612 639 1654
rect 667 1612 682 1654
rect 864 1637 874 1644
tri 874 1637 881 1644 sw
rect 864 1612 881 1637
rect 1005 1612 1022 1644
rect 1204 1612 1219 1654
rect 1247 1612 1262 1654
rect 1444 1637 1454 1644
tri 1454 1637 1461 1644 sw
rect 1444 1612 1461 1637
rect 1585 1612 1602 1644
rect 1784 1612 1799 1654
rect 1827 1612 1842 1654
rect 2024 1637 2034 1644
tri 2034 1637 2041 1644 sw
rect 2024 1612 2041 1637
rect 2165 1612 2182 1644
rect 2364 1612 2379 1654
rect 2407 1612 2422 1654
rect 2604 1637 2614 1644
tri 2614 1637 2621 1644 sw
rect 2604 1612 2621 1637
rect 2745 1612 2762 1644
rect 2944 1612 2959 1654
rect 2987 1612 3002 1654
rect 3184 1637 3194 1644
tri 3194 1637 3201 1644 sw
rect 3184 1612 3201 1637
rect 3325 1612 3342 1644
rect 3524 1612 3539 1654
rect 3567 1612 3582 1654
rect 3764 1637 3774 1644
tri 3774 1637 3781 1644 sw
rect 3764 1612 3781 1637
rect 3905 1612 3922 1644
rect 4104 1612 4119 1654
rect 4147 1612 4162 1654
rect 4344 1637 4354 1644
tri 4354 1637 4361 1644 sw
rect 4344 1612 4361 1637
rect 4485 1612 4502 1644
rect 4684 1612 4699 1654
rect 4727 1612 4742 1654
rect 4924 1637 4934 1644
tri 4934 1637 4941 1644 sw
rect 4924 1612 4941 1637
rect 5065 1612 5082 1644
rect 5264 1612 5279 1654
rect 5307 1612 5322 1654
rect 5504 1637 5514 1644
tri 5514 1637 5521 1644 sw
rect 5504 1612 5521 1637
rect 5645 1612 5662 1644
rect 5844 1612 5859 1654
rect 5887 1612 5902 1654
rect 6084 1637 6094 1644
tri 6094 1637 6101 1644 sw
rect 6084 1612 6101 1637
rect 6225 1612 6242 1644
rect 6424 1612 6439 1654
rect -233 1574 -201 1588
rect 347 1574 379 1588
rect 927 1574 959 1588
rect 1507 1574 1539 1588
rect 2087 1574 2119 1588
rect 2667 1574 2699 1588
rect 3247 1574 3279 1588
rect 3827 1574 3859 1588
rect 4407 1574 4439 1588
rect 4987 1574 5019 1588
rect 5567 1574 5599 1588
rect 6147 1574 6179 1588
rect -419 1488 -404 1516
rect -338 1488 -323 1516
rect -111 1488 -96 1516
rect -29 1488 -14 1517
rect 161 1488 176 1516
rect 242 1488 257 1516
rect 469 1488 484 1516
rect 551 1488 566 1517
rect 741 1488 756 1516
rect 822 1488 837 1516
rect 1049 1488 1064 1516
rect 1131 1488 1146 1517
rect 1321 1488 1336 1516
rect 1402 1488 1417 1516
rect 1629 1488 1644 1516
rect 1711 1488 1726 1517
rect 1901 1488 1916 1516
rect 1982 1488 1997 1516
rect 2209 1488 2224 1516
rect 2291 1488 2306 1517
rect 2481 1488 2496 1516
rect 2562 1488 2577 1516
rect 2789 1488 2804 1516
rect 2871 1488 2886 1517
rect 3061 1488 3076 1516
rect 3142 1488 3157 1516
rect 3369 1488 3384 1516
rect 3451 1488 3466 1517
rect 3641 1488 3656 1516
rect 3722 1488 3737 1516
rect 3949 1488 3964 1516
rect 4031 1488 4046 1517
rect 4221 1488 4236 1516
rect 4302 1488 4317 1516
rect 4529 1488 4544 1516
rect 4611 1488 4626 1517
rect 4801 1488 4816 1516
rect 4882 1488 4897 1516
rect 5109 1488 5124 1516
rect 5191 1488 5206 1517
rect 5381 1488 5396 1516
rect 5462 1488 5477 1516
rect 5689 1488 5704 1516
rect 5771 1488 5786 1517
rect 5961 1488 5976 1516
rect 6042 1488 6057 1516
rect 6269 1488 6284 1516
rect 6351 1488 6366 1517
rect -493 1342 -478 1384
rect -296 1367 -286 1374
tri -286 1367 -279 1374 sw
rect -296 1342 -279 1367
rect -155 1342 -138 1374
rect 44 1342 59 1384
rect 87 1342 102 1384
rect 284 1367 294 1374
tri 294 1367 301 1374 sw
rect 284 1342 301 1367
rect 425 1342 442 1374
rect 624 1342 639 1384
rect 667 1342 682 1384
rect 864 1367 874 1374
tri 874 1367 881 1374 sw
rect 864 1342 881 1367
rect 1005 1342 1022 1374
rect 1204 1342 1219 1384
rect 1247 1342 1262 1384
rect 1444 1367 1454 1374
tri 1454 1367 1461 1374 sw
rect 1444 1342 1461 1367
rect 1585 1342 1602 1374
rect 1784 1342 1799 1384
rect 1827 1342 1842 1384
rect 2024 1367 2034 1374
tri 2034 1367 2041 1374 sw
rect 2024 1342 2041 1367
rect 2165 1342 2182 1374
rect 2364 1342 2379 1384
rect 2407 1342 2422 1384
rect 2604 1367 2614 1374
tri 2614 1367 2621 1374 sw
rect 2604 1342 2621 1367
rect 2745 1342 2762 1374
rect 2944 1342 2959 1384
rect 2987 1342 3002 1384
rect 3184 1367 3194 1374
tri 3194 1367 3201 1374 sw
rect 3184 1342 3201 1367
rect 3325 1342 3342 1374
rect 3524 1342 3539 1384
rect 3567 1342 3582 1384
rect 3764 1367 3774 1374
tri 3774 1367 3781 1374 sw
rect 3764 1342 3781 1367
rect 3905 1342 3922 1374
rect 4104 1342 4119 1384
rect 4147 1342 4162 1384
rect 4344 1367 4354 1374
tri 4354 1367 4361 1374 sw
rect 4344 1342 4361 1367
rect 4485 1342 4502 1374
rect 4684 1342 4699 1384
rect 4727 1342 4742 1384
rect 4924 1367 4934 1374
tri 4934 1367 4941 1374 sw
rect 4924 1342 4941 1367
rect 5065 1342 5082 1374
rect 5264 1342 5279 1384
rect 5307 1342 5322 1384
rect 5504 1367 5514 1374
tri 5514 1367 5521 1374 sw
rect 5504 1342 5521 1367
rect 5645 1342 5662 1374
rect 5844 1342 5859 1384
rect 5887 1342 5902 1384
rect 6084 1367 6094 1374
tri 6094 1367 6101 1374 sw
rect 6084 1342 6101 1367
rect 6225 1342 6242 1374
rect 6424 1342 6439 1384
rect -233 1304 -201 1318
rect 347 1304 379 1318
rect 927 1304 959 1318
rect 1507 1304 1539 1318
rect 2087 1304 2119 1318
rect 2667 1304 2699 1318
rect 3247 1304 3279 1318
rect 3827 1304 3859 1318
rect 4407 1304 4439 1318
rect 4987 1304 5019 1318
rect 5567 1304 5599 1318
rect 6147 1304 6179 1318
rect -419 1218 -404 1246
rect -338 1218 -323 1246
rect -111 1218 -96 1246
rect -29 1218 -14 1247
rect 161 1218 176 1246
rect 242 1218 257 1246
rect 469 1218 484 1246
rect 551 1218 566 1247
rect 741 1218 756 1246
rect 822 1218 837 1246
rect 1049 1218 1064 1246
rect 1131 1218 1146 1247
rect 1321 1218 1336 1246
rect 1402 1218 1417 1246
rect 1629 1218 1644 1246
rect 1711 1218 1726 1247
rect 1901 1218 1916 1246
rect 1982 1218 1997 1246
rect 2209 1218 2224 1246
rect 2291 1218 2306 1247
rect 2481 1218 2496 1246
rect 2562 1218 2577 1246
rect 2789 1218 2804 1246
rect 2871 1218 2886 1247
rect 3061 1218 3076 1246
rect 3142 1218 3157 1246
rect 3369 1218 3384 1246
rect 3451 1218 3466 1247
rect 3641 1218 3656 1246
rect 3722 1218 3737 1246
rect 3949 1218 3964 1246
rect 4031 1218 4046 1247
rect 4221 1218 4236 1246
rect 4302 1218 4317 1246
rect 4529 1218 4544 1246
rect 4611 1218 4626 1247
rect 4801 1218 4816 1246
rect 4882 1218 4897 1246
rect 5109 1218 5124 1246
rect 5191 1218 5206 1247
rect 5381 1218 5396 1246
rect 5462 1218 5477 1246
rect 5689 1218 5704 1246
rect 5771 1218 5786 1247
rect 5961 1218 5976 1246
rect 6042 1218 6057 1246
rect 6269 1218 6284 1246
rect 6351 1218 6366 1247
rect -493 1072 -478 1114
rect -296 1097 -286 1104
tri -286 1097 -279 1104 sw
rect -296 1072 -279 1097
rect -155 1072 -138 1104
rect 44 1072 59 1114
rect 87 1072 102 1114
rect 284 1097 294 1104
tri 294 1097 301 1104 sw
rect 284 1072 301 1097
rect 425 1072 442 1104
rect 624 1072 639 1114
rect 667 1072 682 1114
rect 864 1097 874 1104
tri 874 1097 881 1104 sw
rect 864 1072 881 1097
rect 1005 1072 1022 1104
rect 1204 1072 1219 1114
rect 1247 1072 1262 1114
rect 1444 1097 1454 1104
tri 1454 1097 1461 1104 sw
rect 1444 1072 1461 1097
rect 1585 1072 1602 1104
rect 1784 1072 1799 1114
rect 1827 1072 1842 1114
rect 2024 1097 2034 1104
tri 2034 1097 2041 1104 sw
rect 2024 1072 2041 1097
rect 2165 1072 2182 1104
rect 2364 1072 2379 1114
rect 2407 1072 2422 1114
rect 2604 1097 2614 1104
tri 2614 1097 2621 1104 sw
rect 2604 1072 2621 1097
rect 2745 1072 2762 1104
rect 2944 1072 2959 1114
rect 2987 1072 3002 1114
rect 3184 1097 3194 1104
tri 3194 1097 3201 1104 sw
rect 3184 1072 3201 1097
rect 3325 1072 3342 1104
rect 3524 1072 3539 1114
rect 3567 1072 3582 1114
rect 3764 1097 3774 1104
tri 3774 1097 3781 1104 sw
rect 3764 1072 3781 1097
rect 3905 1072 3922 1104
rect 4104 1072 4119 1114
rect 4147 1072 4162 1114
rect 4344 1097 4354 1104
tri 4354 1097 4361 1104 sw
rect 4344 1072 4361 1097
rect 4485 1072 4502 1104
rect 4684 1072 4699 1114
rect 4727 1072 4742 1114
rect 4924 1097 4934 1104
tri 4934 1097 4941 1104 sw
rect 4924 1072 4941 1097
rect 5065 1072 5082 1104
rect 5264 1072 5279 1114
rect 5307 1072 5322 1114
rect 5504 1097 5514 1104
tri 5514 1097 5521 1104 sw
rect 5504 1072 5521 1097
rect 5645 1072 5662 1104
rect 5844 1072 5859 1114
rect 5887 1072 5902 1114
rect 6084 1097 6094 1104
tri 6094 1097 6101 1104 sw
rect 6084 1072 6101 1097
rect 6225 1072 6242 1104
rect 6424 1072 6439 1114
rect -233 1034 -201 1048
rect 347 1034 379 1048
rect 927 1034 959 1048
rect 1507 1034 1539 1048
rect 2087 1034 2119 1048
rect 2667 1034 2699 1048
rect 3247 1034 3279 1048
rect 3827 1034 3859 1048
rect 4407 1034 4439 1048
rect 4987 1034 5019 1048
rect 5567 1034 5599 1048
rect 6147 1034 6179 1048
rect -419 948 -404 976
rect -338 948 -323 976
rect -111 948 -96 976
rect -29 948 -14 977
rect 161 948 176 976
rect 242 948 257 976
rect 469 948 484 976
rect 551 948 566 977
rect 741 948 756 976
rect 822 948 837 976
rect 1049 948 1064 976
rect 1131 948 1146 977
rect 1321 948 1336 976
rect 1402 948 1417 976
rect 1629 948 1644 976
rect 1711 948 1726 977
rect 1901 948 1916 976
rect 1982 948 1997 976
rect 2209 948 2224 976
rect 2291 948 2306 977
rect 2481 948 2496 976
rect 2562 948 2577 976
rect 2789 948 2804 976
rect 2871 948 2886 977
rect 3061 948 3076 976
rect 3142 948 3157 976
rect 3369 948 3384 976
rect 3451 948 3466 977
rect 3641 948 3656 976
rect 3722 948 3737 976
rect 3949 948 3964 976
rect 4031 948 4046 977
rect 4221 948 4236 976
rect 4302 948 4317 976
rect 4529 948 4544 976
rect 4611 948 4626 977
rect 4801 948 4816 976
rect 4882 948 4897 976
rect 5109 948 5124 976
rect 5191 948 5206 977
rect 5381 948 5396 976
rect 5462 948 5477 976
rect 5689 948 5704 976
rect 5771 948 5786 977
rect 5961 948 5976 976
rect 6042 948 6057 976
rect 6269 948 6284 976
rect 6351 948 6366 977
rect -493 802 -478 844
rect -296 827 -286 834
tri -286 827 -279 834 sw
rect -296 802 -279 827
rect -155 802 -138 834
rect 44 802 59 844
rect 87 802 102 844
rect 284 827 294 834
tri 294 827 301 834 sw
rect 284 802 301 827
rect 425 802 442 834
rect 624 802 639 844
rect 667 802 682 844
rect 864 827 874 834
tri 874 827 881 834 sw
rect 864 802 881 827
rect 1005 802 1022 834
rect 1204 802 1219 844
rect 1247 802 1262 844
rect 1444 827 1454 834
tri 1454 827 1461 834 sw
rect 1444 802 1461 827
rect 1585 802 1602 834
rect 1784 802 1799 844
rect 1827 802 1842 844
rect 2024 827 2034 834
tri 2034 827 2041 834 sw
rect 2024 802 2041 827
rect 2165 802 2182 834
rect 2364 802 2379 844
rect 2407 802 2422 844
rect 2604 827 2614 834
tri 2614 827 2621 834 sw
rect 2604 802 2621 827
rect 2745 802 2762 834
rect 2944 802 2959 844
rect 2987 802 3002 844
rect 3184 827 3194 834
tri 3194 827 3201 834 sw
rect 3184 802 3201 827
rect 3325 802 3342 834
rect 3524 802 3539 844
rect 3567 802 3582 844
rect 3764 827 3774 834
tri 3774 827 3781 834 sw
rect 3764 802 3781 827
rect 3905 802 3922 834
rect 4104 802 4119 844
rect 4147 802 4162 844
rect 4344 827 4354 834
tri 4354 827 4361 834 sw
rect 4344 802 4361 827
rect 4485 802 4502 834
rect 4684 802 4699 844
rect 4727 802 4742 844
rect 4924 827 4934 834
tri 4934 827 4941 834 sw
rect 4924 802 4941 827
rect 5065 802 5082 834
rect 5264 802 5279 844
rect 5307 802 5322 844
rect 5504 827 5514 834
tri 5514 827 5521 834 sw
rect 5504 802 5521 827
rect 5645 802 5662 834
rect 5844 802 5859 844
rect 5887 802 5902 844
rect 6084 827 6094 834
tri 6094 827 6101 834 sw
rect 6084 802 6101 827
rect 6225 802 6242 834
rect 6424 802 6439 844
rect -233 764 -201 778
rect 347 764 379 778
rect 927 764 959 778
rect 1507 764 1539 778
rect 2087 764 2119 778
rect 2667 764 2699 778
rect 3247 764 3279 778
rect 3827 764 3859 778
rect 4407 764 4439 778
rect 4987 764 5019 778
rect 5567 764 5599 778
rect 6147 764 6179 778
rect -419 678 -404 706
rect -338 678 -323 706
rect -111 678 -96 706
rect -29 678 -14 707
rect 161 678 176 706
rect 242 678 257 706
rect 469 678 484 706
rect 551 678 566 707
rect 741 678 756 706
rect 822 678 837 706
rect 1049 678 1064 706
rect 1131 678 1146 707
rect 1321 678 1336 706
rect 1402 678 1417 706
rect 1629 678 1644 706
rect 1711 678 1726 707
rect 1901 678 1916 706
rect 1982 678 1997 706
rect 2209 678 2224 706
rect 2291 678 2306 707
rect 2481 678 2496 706
rect 2562 678 2577 706
rect 2789 678 2804 706
rect 2871 678 2886 707
rect 3061 678 3076 706
rect 3142 678 3157 706
rect 3369 678 3384 706
rect 3451 678 3466 707
rect 3641 678 3656 706
rect 3722 678 3737 706
rect 3949 678 3964 706
rect 4031 678 4046 707
rect 4221 678 4236 706
rect 4302 678 4317 706
rect 4529 678 4544 706
rect 4611 678 4626 707
rect 4801 678 4816 706
rect 4882 678 4897 706
rect 5109 678 5124 706
rect 5191 678 5206 707
rect 5381 678 5396 706
rect 5462 678 5477 706
rect 5689 678 5704 706
rect 5771 678 5786 707
rect 5961 678 5976 706
rect 6042 678 6057 706
rect 6269 678 6284 706
rect 6351 678 6366 707
rect -493 532 -478 574
rect -296 557 -286 564
tri -286 557 -279 564 sw
rect -296 532 -279 557
rect -155 532 -138 564
rect 44 532 59 574
rect 87 532 102 574
rect 284 557 294 564
tri 294 557 301 564 sw
rect 284 532 301 557
rect 425 532 442 564
rect 624 532 639 574
rect 667 532 682 574
rect 864 557 874 564
tri 874 557 881 564 sw
rect 864 532 881 557
rect 1005 532 1022 564
rect 1204 532 1219 574
rect 1247 532 1262 574
rect 1444 557 1454 564
tri 1454 557 1461 564 sw
rect 1444 532 1461 557
rect 1585 532 1602 564
rect 1784 532 1799 574
rect 1827 532 1842 574
rect 2024 557 2034 564
tri 2034 557 2041 564 sw
rect 2024 532 2041 557
rect 2165 532 2182 564
rect 2364 532 2379 574
rect 2407 532 2422 574
rect 2604 557 2614 564
tri 2614 557 2621 564 sw
rect 2604 532 2621 557
rect 2745 532 2762 564
rect 2944 532 2959 574
rect 2987 532 3002 574
rect 3184 557 3194 564
tri 3194 557 3201 564 sw
rect 3184 532 3201 557
rect 3325 532 3342 564
rect 3524 532 3539 574
rect 3567 532 3582 574
rect 3764 557 3774 564
tri 3774 557 3781 564 sw
rect 3764 532 3781 557
rect 3905 532 3922 564
rect 4104 532 4119 574
rect 4147 532 4162 574
rect 4344 557 4354 564
tri 4354 557 4361 564 sw
rect 4344 532 4361 557
rect 4485 532 4502 564
rect 4684 532 4699 574
rect 4727 532 4742 574
rect 4924 557 4934 564
tri 4934 557 4941 564 sw
rect 4924 532 4941 557
rect 5065 532 5082 564
rect 5264 532 5279 574
rect 5307 532 5322 574
rect 5504 557 5514 564
tri 5514 557 5521 564 sw
rect 5504 532 5521 557
rect 5645 532 5662 564
rect 5844 532 5859 574
rect 5887 532 5902 574
rect 6084 557 6094 564
tri 6094 557 6101 564 sw
rect 6084 532 6101 557
rect 6225 532 6242 564
rect 6424 532 6439 574
rect -233 494 -201 508
rect 347 494 379 508
rect 927 494 959 508
rect 1507 494 1539 508
rect 2087 494 2119 508
rect 2667 494 2699 508
rect 3247 494 3279 508
rect 3827 494 3859 508
rect 4407 494 4439 508
rect 4987 494 5019 508
rect 5567 494 5599 508
rect 6147 494 6179 508
rect -419 408 -404 436
rect -338 408 -323 436
rect -111 408 -96 436
rect -29 408 -14 437
rect 161 408 176 436
rect 242 408 257 436
rect 469 408 484 436
rect 551 408 566 437
rect 741 408 756 436
rect 822 408 837 436
rect 1049 408 1064 436
rect 1131 408 1146 437
rect 1321 408 1336 436
rect 1402 408 1417 436
rect 1629 408 1644 436
rect 1711 408 1726 437
rect 1901 408 1916 436
rect 1982 408 1997 436
rect 2209 408 2224 436
rect 2291 408 2306 437
rect 2481 408 2496 436
rect 2562 408 2577 436
rect 2789 408 2804 436
rect 2871 408 2886 437
rect 3061 408 3076 436
rect 3142 408 3157 436
rect 3369 408 3384 436
rect 3451 408 3466 437
rect 3641 408 3656 436
rect 3722 408 3737 436
rect 3949 408 3964 436
rect 4031 408 4046 437
rect 4221 408 4236 436
rect 4302 408 4317 436
rect 4529 408 4544 436
rect 4611 408 4626 437
rect 4801 408 4816 436
rect 4882 408 4897 436
rect 5109 408 5124 436
rect 5191 408 5206 437
rect 5381 408 5396 436
rect 5462 408 5477 436
rect 5689 408 5704 436
rect 5771 408 5786 437
rect 5961 408 5976 436
rect 6042 408 6057 436
rect 6269 408 6284 436
rect 6351 408 6366 437
rect -493 262 -478 304
rect -296 287 -286 294
tri -286 287 -279 294 sw
rect -296 262 -279 287
rect -155 262 -138 294
rect 44 262 59 304
rect 87 262 102 304
rect 284 287 294 294
tri 294 287 301 294 sw
rect 284 262 301 287
rect 425 262 442 294
rect 624 262 639 304
rect 667 262 682 304
rect 864 287 874 294
tri 874 287 881 294 sw
rect 864 262 881 287
rect 1005 262 1022 294
rect 1204 262 1219 304
rect 1247 262 1262 304
rect 1444 287 1454 294
tri 1454 287 1461 294 sw
rect 1444 262 1461 287
rect 1585 262 1602 294
rect 1784 262 1799 304
rect 1827 262 1842 304
rect 2024 287 2034 294
tri 2034 287 2041 294 sw
rect 2024 262 2041 287
rect 2165 262 2182 294
rect 2364 262 2379 304
rect 2407 262 2422 304
rect 2604 287 2614 294
tri 2614 287 2621 294 sw
rect 2604 262 2621 287
rect 2745 262 2762 294
rect 2944 262 2959 304
rect 2987 262 3002 304
rect 3184 287 3194 294
tri 3194 287 3201 294 sw
rect 3184 262 3201 287
rect 3325 262 3342 294
rect 3524 262 3539 304
rect 3567 262 3582 304
rect 3764 287 3774 294
tri 3774 287 3781 294 sw
rect 3764 262 3781 287
rect 3905 262 3922 294
rect 4104 262 4119 304
rect 4147 262 4162 304
rect 4344 287 4354 294
tri 4354 287 4361 294 sw
rect 4344 262 4361 287
rect 4485 262 4502 294
rect 4684 262 4699 304
rect 4727 262 4742 304
rect 4924 287 4934 294
tri 4934 287 4941 294 sw
rect 4924 262 4941 287
rect 5065 262 5082 294
rect 5264 262 5279 304
rect 5307 262 5322 304
rect 5504 287 5514 294
tri 5514 287 5521 294 sw
rect 5504 262 5521 287
rect 5645 262 5662 294
rect 5844 262 5859 304
rect 5887 262 5902 304
rect 6084 287 6094 294
tri 6094 287 6101 294 sw
rect 6084 262 6101 287
rect 6225 262 6242 294
rect 6424 262 6439 304
rect -233 224 -201 238
rect 347 224 379 238
rect 927 224 959 238
rect 1507 224 1539 238
rect 2087 224 2119 238
rect 2667 224 2699 238
rect 3247 224 3279 238
rect 3827 224 3859 238
rect 4407 224 4439 238
rect 4987 224 5019 238
rect 5567 224 5599 238
rect 6147 224 6179 238
rect -419 138 -404 166
rect -338 138 -323 166
rect -111 138 -96 166
rect -29 138 -14 167
rect 161 138 176 166
rect 242 138 257 166
rect 469 138 484 166
rect 551 138 566 167
rect 741 138 756 166
rect 822 138 837 166
rect 1049 138 1064 166
rect 1131 138 1146 167
rect 1321 138 1336 166
rect 1402 138 1417 166
rect 1629 138 1644 166
rect 1711 138 1726 167
rect 1901 138 1916 166
rect 1982 138 1997 166
rect 2209 138 2224 166
rect 2291 138 2306 167
rect 2481 138 2496 166
rect 2562 138 2577 166
rect 2789 138 2804 166
rect 2871 138 2886 167
rect 3061 138 3076 166
rect 3142 138 3157 166
rect 3369 138 3384 166
rect 3451 138 3466 167
rect 3641 138 3656 166
rect 3722 138 3737 166
rect 3949 138 3964 166
rect 4031 138 4046 167
rect 4221 138 4236 166
rect 4302 138 4317 166
rect 4529 138 4544 166
rect 4611 138 4626 167
rect 4801 138 4816 166
rect 4882 138 4897 166
rect 5109 138 5124 166
rect 5191 138 5206 167
rect 5381 138 5396 166
rect 5462 138 5477 166
rect 5689 138 5704 166
rect 5771 138 5786 167
rect 5961 138 5976 166
rect 6042 138 6057 166
rect 6269 138 6284 166
rect 6351 138 6366 167
rect -493 -8 -478 34
rect -296 17 -286 24
tri -286 17 -279 24 sw
rect -296 -8 -279 17
rect -155 -8 -138 24
rect 44 -8 59 34
rect 87 -8 102 34
rect 284 17 294 24
tri 294 17 301 24 sw
rect 284 -8 301 17
rect 425 -8 442 24
rect 624 -8 639 34
rect 667 -8 682 34
rect 864 17 874 24
tri 874 17 881 24 sw
rect 864 -8 881 17
rect 1005 -8 1022 24
rect 1204 -8 1219 34
rect 1247 -8 1262 34
rect 1444 17 1454 24
tri 1454 17 1461 24 sw
rect 1444 -8 1461 17
rect 1585 -8 1602 24
rect 1784 -8 1799 34
rect 1827 -8 1842 34
rect 2024 17 2034 24
tri 2034 17 2041 24 sw
rect 2024 -8 2041 17
rect 2165 -8 2182 24
rect 2364 -8 2379 34
rect 2407 -8 2422 34
rect 2604 17 2614 24
tri 2614 17 2621 24 sw
rect 2604 -8 2621 17
rect 2745 -8 2762 24
rect 2944 -8 2959 34
rect 2987 -8 3002 34
rect 3184 17 3194 24
tri 3194 17 3201 24 sw
rect 3184 -8 3201 17
rect 3325 -8 3342 24
rect 3524 -8 3539 34
rect 3567 -8 3582 34
rect 3764 17 3774 24
tri 3774 17 3781 24 sw
rect 3764 -8 3781 17
rect 3905 -8 3922 24
rect 4104 -8 4119 34
rect 4147 -8 4162 34
rect 4344 17 4354 24
tri 4354 17 4361 24 sw
rect 4344 -8 4361 17
rect 4485 -8 4502 24
rect 4684 -8 4699 34
rect 4727 -8 4742 34
rect 4924 17 4934 24
tri 4934 17 4941 24 sw
rect 4924 -8 4941 17
rect 5065 -8 5082 24
rect 5264 -8 5279 34
rect 5307 -8 5322 34
rect 5504 17 5514 24
tri 5514 17 5521 24 sw
rect 5504 -8 5521 17
rect 5645 -8 5662 24
rect 5844 -8 5859 34
rect 5887 -8 5902 34
rect 6084 17 6094 24
tri 6094 17 6101 24 sw
rect 6084 -8 6101 17
rect 6225 -8 6242 24
rect 6424 -8 6439 34
rect -233 -46 -201 -32
rect 347 -46 379 -32
rect 927 -46 959 -32
rect 1507 -46 1539 -32
rect 2087 -46 2119 -32
rect 2667 -46 2699 -32
rect 3247 -46 3279 -32
rect 3827 -46 3859 -32
rect 4407 -46 4439 -32
rect 4987 -46 5019 -32
rect 5567 -46 5599 -32
rect 6147 -46 6179 -32
rect -419 -132 -404 -104
rect -338 -132 -323 -104
rect -111 -132 -96 -104
rect -29 -132 -14 -103
rect 161 -132 176 -104
rect 242 -132 257 -104
rect 469 -132 484 -104
rect 551 -132 566 -103
rect 741 -132 756 -104
rect 822 -132 837 -104
rect 1049 -132 1064 -104
rect 1131 -132 1146 -103
rect 1321 -132 1336 -104
rect 1402 -132 1417 -104
rect 1629 -132 1644 -104
rect 1711 -132 1726 -103
rect 1901 -132 1916 -104
rect 1982 -132 1997 -104
rect 2209 -132 2224 -104
rect 2291 -132 2306 -103
rect 2481 -132 2496 -104
rect 2562 -132 2577 -104
rect 2789 -132 2804 -104
rect 2871 -132 2886 -103
rect 3061 -132 3076 -104
rect 3142 -132 3157 -104
rect 3369 -132 3384 -104
rect 3451 -132 3466 -103
rect 3641 -132 3656 -104
rect 3722 -132 3737 -104
rect 3949 -132 3964 -104
rect 4031 -132 4046 -103
rect 4221 -132 4236 -104
rect 4302 -132 4317 -104
rect 4529 -132 4544 -104
rect 4611 -132 4626 -103
rect 4801 -132 4816 -104
rect 4882 -132 4897 -104
rect 5109 -132 5124 -104
rect 5191 -132 5206 -103
rect 5381 -132 5396 -104
rect 5462 -132 5477 -104
rect 5689 -132 5704 -104
rect 5771 -132 5786 -103
rect 5961 -132 5976 -104
rect 6042 -132 6057 -104
rect 6269 -132 6284 -104
rect 6351 -132 6366 -103
rect -493 -278 -478 -236
rect -296 -253 -286 -246
tri -286 -253 -279 -246 sw
rect -296 -278 -279 -253
rect -155 -278 -138 -246
rect 44 -278 59 -236
rect 87 -278 102 -236
rect 284 -253 294 -246
tri 294 -253 301 -246 sw
rect 284 -278 301 -253
rect 425 -278 442 -246
rect 624 -278 639 -236
rect 667 -278 682 -236
rect 864 -253 874 -246
tri 874 -253 881 -246 sw
rect 864 -278 881 -253
rect 1005 -278 1022 -246
rect 1204 -278 1219 -236
rect 1247 -278 1262 -236
rect 1444 -253 1454 -246
tri 1454 -253 1461 -246 sw
rect 1444 -278 1461 -253
rect 1585 -278 1602 -246
rect 1784 -278 1799 -236
rect 1827 -278 1842 -236
rect 2024 -253 2034 -246
tri 2034 -253 2041 -246 sw
rect 2024 -278 2041 -253
rect 2165 -278 2182 -246
rect 2364 -278 2379 -236
rect 2407 -278 2422 -236
rect 2604 -253 2614 -246
tri 2614 -253 2621 -246 sw
rect 2604 -278 2621 -253
rect 2745 -278 2762 -246
rect 2944 -278 2959 -236
rect 2987 -278 3002 -236
rect 3184 -253 3194 -246
tri 3194 -253 3201 -246 sw
rect 3184 -278 3201 -253
rect 3325 -278 3342 -246
rect 3524 -278 3539 -236
rect 3567 -278 3582 -236
rect 3764 -253 3774 -246
tri 3774 -253 3781 -246 sw
rect 3764 -278 3781 -253
rect 3905 -278 3922 -246
rect 4104 -278 4119 -236
rect 4147 -278 4162 -236
rect 4344 -253 4354 -246
tri 4354 -253 4361 -246 sw
rect 4344 -278 4361 -253
rect 4485 -278 4502 -246
rect 4684 -278 4699 -236
rect 4727 -278 4742 -236
rect 4924 -253 4934 -246
tri 4934 -253 4941 -246 sw
rect 4924 -278 4941 -253
rect 5065 -278 5082 -246
rect 5264 -278 5279 -236
rect 5307 -278 5322 -236
rect 5504 -253 5514 -246
tri 5514 -253 5521 -246 sw
rect 5504 -278 5521 -253
rect 5645 -278 5662 -246
rect 5844 -278 5859 -236
rect 5887 -278 5902 -236
rect 6084 -253 6094 -246
tri 6094 -253 6101 -246 sw
rect 6084 -278 6101 -253
rect 6225 -278 6242 -246
rect 6424 -278 6439 -236
rect -233 -316 -201 -302
rect 347 -316 379 -302
rect 927 -316 959 -302
rect 1507 -316 1539 -302
rect 2087 -316 2119 -302
rect 2667 -316 2699 -302
rect 3247 -316 3279 -302
rect 3827 -316 3859 -302
rect 4407 -316 4439 -302
rect 4987 -316 5019 -302
rect 5567 -316 5599 -302
rect 6147 -316 6179 -302
rect -419 -402 -404 -374
rect -338 -402 -323 -374
rect -111 -402 -96 -374
rect -29 -402 -14 -373
rect 161 -402 176 -374
rect 242 -402 257 -374
rect 469 -402 484 -374
rect 551 -402 566 -373
rect 741 -402 756 -374
rect 822 -402 837 -374
rect 1049 -402 1064 -374
rect 1131 -402 1146 -373
rect 1321 -402 1336 -374
rect 1402 -402 1417 -374
rect 1629 -402 1644 -374
rect 1711 -402 1726 -373
rect 1901 -402 1916 -374
rect 1982 -402 1997 -374
rect 2209 -402 2224 -374
rect 2291 -402 2306 -373
rect 2481 -402 2496 -374
rect 2562 -402 2577 -374
rect 2789 -402 2804 -374
rect 2871 -402 2886 -373
rect 3061 -402 3076 -374
rect 3142 -402 3157 -374
rect 3369 -402 3384 -374
rect 3451 -402 3466 -373
rect 3641 -402 3656 -374
rect 3722 -402 3737 -374
rect 3949 -402 3964 -374
rect 4031 -402 4046 -373
rect 4221 -402 4236 -374
rect 4302 -402 4317 -374
rect 4529 -402 4544 -374
rect 4611 -402 4626 -373
rect 4801 -402 4816 -374
rect 4882 -402 4897 -374
rect 5109 -402 5124 -374
rect 5191 -402 5206 -373
rect 5381 -402 5396 -374
rect 5462 -402 5477 -374
rect 5689 -402 5704 -374
rect 5771 -402 5786 -373
rect 5961 -402 5976 -374
rect 6042 -402 6057 -374
rect 6269 -402 6284 -374
rect 6351 -402 6366 -373
rect -493 -548 -478 -506
rect -296 -523 -286 -516
tri -286 -523 -279 -516 sw
rect -296 -548 -279 -523
rect -155 -548 -138 -516
rect 44 -548 59 -506
rect 87 -548 102 -506
rect 284 -523 294 -516
tri 294 -523 301 -516 sw
rect 284 -548 301 -523
rect 425 -548 442 -516
rect 624 -548 639 -506
rect 667 -548 682 -506
rect 864 -523 874 -516
tri 874 -523 881 -516 sw
rect 864 -548 881 -523
rect 1005 -548 1022 -516
rect 1204 -548 1219 -506
rect 1247 -548 1262 -506
rect 1444 -523 1454 -516
tri 1454 -523 1461 -516 sw
rect 1444 -548 1461 -523
rect 1585 -548 1602 -516
rect 1784 -548 1799 -506
rect 1827 -548 1842 -506
rect 2024 -523 2034 -516
tri 2034 -523 2041 -516 sw
rect 2024 -548 2041 -523
rect 2165 -548 2182 -516
rect 2364 -548 2379 -506
rect 2407 -548 2422 -506
rect 2604 -523 2614 -516
tri 2614 -523 2621 -516 sw
rect 2604 -548 2621 -523
rect 2745 -548 2762 -516
rect 2944 -548 2959 -506
rect 2987 -548 3002 -506
rect 3184 -523 3194 -516
tri 3194 -523 3201 -516 sw
rect 3184 -548 3201 -523
rect 3325 -548 3342 -516
rect 3524 -548 3539 -506
rect 3567 -548 3582 -506
rect 3764 -523 3774 -516
tri 3774 -523 3781 -516 sw
rect 3764 -548 3781 -523
rect 3905 -548 3922 -516
rect 4104 -548 4119 -506
rect 4147 -548 4162 -506
rect 4344 -523 4354 -516
tri 4354 -523 4361 -516 sw
rect 4344 -548 4361 -523
rect 4485 -548 4502 -516
rect 4684 -548 4699 -506
rect 4727 -548 4742 -506
rect 4924 -523 4934 -516
tri 4934 -523 4941 -516 sw
rect 4924 -548 4941 -523
rect 5065 -548 5082 -516
rect 5264 -548 5279 -506
rect 5307 -548 5322 -506
rect 5504 -523 5514 -516
tri 5514 -523 5521 -516 sw
rect 5504 -548 5521 -523
rect 5645 -548 5662 -516
rect 5844 -548 5859 -506
rect 5887 -548 5902 -506
rect 6084 -523 6094 -516
tri 6094 -523 6101 -516 sw
rect 6084 -548 6101 -523
rect 6225 -548 6242 -516
rect 6424 -548 6439 -506
rect -233 -586 -201 -572
rect 347 -586 379 -572
rect 927 -586 959 -572
rect 1507 -586 1539 -572
rect 2087 -586 2119 -572
rect 2667 -586 2699 -572
rect 3247 -586 3279 -572
rect 3827 -586 3859 -572
rect 4407 -586 4439 -572
rect 4987 -586 5019 -572
rect 5567 -586 5599 -572
rect 6147 -586 6179 -572
rect -419 -672 -404 -644
rect -338 -672 -323 -644
rect -111 -672 -96 -644
rect -29 -672 -14 -643
rect 161 -672 176 -644
rect 242 -672 257 -644
rect 469 -672 484 -644
rect 551 -672 566 -643
rect 741 -672 756 -644
rect 822 -672 837 -644
rect 1049 -672 1064 -644
rect 1131 -672 1146 -643
rect 1321 -672 1336 -644
rect 1402 -672 1417 -644
rect 1629 -672 1644 -644
rect 1711 -672 1726 -643
rect 1901 -672 1916 -644
rect 1982 -672 1997 -644
rect 2209 -672 2224 -644
rect 2291 -672 2306 -643
rect 2481 -672 2496 -644
rect 2562 -672 2577 -644
rect 2789 -672 2804 -644
rect 2871 -672 2886 -643
rect 3061 -672 3076 -644
rect 3142 -672 3157 -644
rect 3369 -672 3384 -644
rect 3451 -672 3466 -643
rect 3641 -672 3656 -644
rect 3722 -672 3737 -644
rect 3949 -672 3964 -644
rect 4031 -672 4046 -643
rect 4221 -672 4236 -644
rect 4302 -672 4317 -644
rect 4529 -672 4544 -644
rect 4611 -672 4626 -643
rect 4801 -672 4816 -644
rect 4882 -672 4897 -644
rect 5109 -672 5124 -644
rect 5191 -672 5206 -643
rect 5381 -672 5396 -644
rect 5462 -672 5477 -644
rect 5689 -672 5704 -644
rect 5771 -672 5786 -643
rect 5961 -672 5976 -644
rect 6042 -672 6057 -644
rect 6269 -672 6284 -644
rect 6351 -672 6366 -643
rect -493 -818 -478 -776
rect -296 -793 -286 -786
tri -286 -793 -279 -786 sw
rect -296 -818 -279 -793
rect -155 -818 -138 -786
rect 44 -818 59 -776
rect 87 -818 102 -776
rect 284 -793 294 -786
tri 294 -793 301 -786 sw
rect 284 -818 301 -793
rect 425 -818 442 -786
rect 624 -818 639 -776
rect 667 -818 682 -776
rect 864 -793 874 -786
tri 874 -793 881 -786 sw
rect 864 -818 881 -793
rect 1005 -818 1022 -786
rect 1204 -818 1219 -776
rect 1247 -818 1262 -776
rect 1444 -793 1454 -786
tri 1454 -793 1461 -786 sw
rect 1444 -818 1461 -793
rect 1585 -818 1602 -786
rect 1784 -818 1799 -776
rect 1827 -818 1842 -776
rect 2024 -793 2034 -786
tri 2034 -793 2041 -786 sw
rect 2024 -818 2041 -793
rect 2165 -818 2182 -786
rect 2364 -818 2379 -776
rect 2407 -818 2422 -776
rect 2604 -793 2614 -786
tri 2614 -793 2621 -786 sw
rect 2604 -818 2621 -793
rect 2745 -818 2762 -786
rect 2944 -818 2959 -776
rect 2987 -818 3002 -776
rect 3184 -793 3194 -786
tri 3194 -793 3201 -786 sw
rect 3184 -818 3201 -793
rect 3325 -818 3342 -786
rect 3524 -818 3539 -776
rect 3567 -818 3582 -776
rect 3764 -793 3774 -786
tri 3774 -793 3781 -786 sw
rect 3764 -818 3781 -793
rect 3905 -818 3922 -786
rect 4104 -818 4119 -776
rect 4147 -818 4162 -776
rect 4344 -793 4354 -786
tri 4354 -793 4361 -786 sw
rect 4344 -818 4361 -793
rect 4485 -818 4502 -786
rect 4684 -818 4699 -776
rect 4727 -818 4742 -776
rect 4924 -793 4934 -786
tri 4934 -793 4941 -786 sw
rect 4924 -818 4941 -793
rect 5065 -818 5082 -786
rect 5264 -818 5279 -776
rect 5307 -818 5322 -776
rect 5504 -793 5514 -786
tri 5514 -793 5521 -786 sw
rect 5504 -818 5521 -793
rect 5645 -818 5662 -786
rect 5844 -818 5859 -776
rect 5887 -818 5902 -776
rect 6084 -793 6094 -786
tri 6094 -793 6101 -786 sw
rect 6084 -818 6101 -793
rect 6225 -818 6242 -786
rect 6424 -818 6439 -776
rect -233 -856 -201 -842
rect 347 -856 379 -842
rect 927 -856 959 -842
rect 1507 -856 1539 -842
rect 2087 -856 2119 -842
rect 2667 -856 2699 -842
rect 3247 -856 3279 -842
rect 3827 -856 3859 -842
rect 4407 -856 4439 -842
rect 4987 -856 5019 -842
rect 5567 -856 5599 -842
rect 6147 -856 6179 -842
rect -419 -942 -404 -914
rect -338 -942 -323 -914
rect -111 -942 -96 -914
rect -29 -942 -14 -913
rect 161 -942 176 -914
rect 242 -942 257 -914
rect 469 -942 484 -914
rect 551 -942 566 -913
rect 741 -942 756 -914
rect 822 -942 837 -914
rect 1049 -942 1064 -914
rect 1131 -942 1146 -913
rect 1321 -942 1336 -914
rect 1402 -942 1417 -914
rect 1629 -942 1644 -914
rect 1711 -942 1726 -913
rect 1901 -942 1916 -914
rect 1982 -942 1997 -914
rect 2209 -942 2224 -914
rect 2291 -942 2306 -913
rect 2481 -942 2496 -914
rect 2562 -942 2577 -914
rect 2789 -942 2804 -914
rect 2871 -942 2886 -913
rect 3061 -942 3076 -914
rect 3142 -942 3157 -914
rect 3369 -942 3384 -914
rect 3451 -942 3466 -913
rect 3641 -942 3656 -914
rect 3722 -942 3737 -914
rect 3949 -942 3964 -914
rect 4031 -942 4046 -913
rect 4221 -942 4236 -914
rect 4302 -942 4317 -914
rect 4529 -942 4544 -914
rect 4611 -942 4626 -913
rect 4801 -942 4816 -914
rect 4882 -942 4897 -914
rect 5109 -942 5124 -914
rect 5191 -942 5206 -913
rect 5381 -942 5396 -914
rect 5462 -942 5477 -914
rect 5689 -942 5704 -914
rect 5771 -942 5786 -913
rect 5961 -942 5976 -914
rect 6042 -942 6057 -914
rect 6269 -942 6284 -914
rect 6351 -942 6366 -913
rect -493 -1088 -478 -1046
rect -296 -1063 -286 -1056
tri -286 -1063 -279 -1056 sw
rect -296 -1088 -279 -1063
rect -155 -1088 -138 -1056
rect 44 -1088 59 -1046
rect 87 -1088 102 -1046
rect 284 -1063 294 -1056
tri 294 -1063 301 -1056 sw
rect 284 -1088 301 -1063
rect 425 -1088 442 -1056
rect 624 -1088 639 -1046
rect 667 -1088 682 -1046
rect 864 -1063 874 -1056
tri 874 -1063 881 -1056 sw
rect 864 -1088 881 -1063
rect 1005 -1088 1022 -1056
rect 1204 -1088 1219 -1046
rect 1247 -1088 1262 -1046
rect 1444 -1063 1454 -1056
tri 1454 -1063 1461 -1056 sw
rect 1444 -1088 1461 -1063
rect 1585 -1088 1602 -1056
rect 1784 -1088 1799 -1046
rect 1827 -1088 1842 -1046
rect 2024 -1063 2034 -1056
tri 2034 -1063 2041 -1056 sw
rect 2024 -1088 2041 -1063
rect 2165 -1088 2182 -1056
rect 2364 -1088 2379 -1046
rect 2407 -1088 2422 -1046
rect 2604 -1063 2614 -1056
tri 2614 -1063 2621 -1056 sw
rect 2604 -1088 2621 -1063
rect 2745 -1088 2762 -1056
rect 2944 -1088 2959 -1046
rect 2987 -1088 3002 -1046
rect 3184 -1063 3194 -1056
tri 3194 -1063 3201 -1056 sw
rect 3184 -1088 3201 -1063
rect 3325 -1088 3342 -1056
rect 3524 -1088 3539 -1046
rect 3567 -1088 3582 -1046
rect 3764 -1063 3774 -1056
tri 3774 -1063 3781 -1056 sw
rect 3764 -1088 3781 -1063
rect 3905 -1088 3922 -1056
rect 4104 -1088 4119 -1046
rect 4147 -1088 4162 -1046
rect 4344 -1063 4354 -1056
tri 4354 -1063 4361 -1056 sw
rect 4344 -1088 4361 -1063
rect 4485 -1088 4502 -1056
rect 4684 -1088 4699 -1046
rect 4727 -1088 4742 -1046
rect 4924 -1063 4934 -1056
tri 4934 -1063 4941 -1056 sw
rect 4924 -1088 4941 -1063
rect 5065 -1088 5082 -1056
rect 5264 -1088 5279 -1046
rect 5307 -1088 5322 -1046
rect 5504 -1063 5514 -1056
tri 5514 -1063 5521 -1056 sw
rect 5504 -1088 5521 -1063
rect 5645 -1088 5662 -1056
rect 5844 -1088 5859 -1046
rect 5887 -1088 5902 -1046
rect 6084 -1063 6094 -1056
tri 6094 -1063 6101 -1056 sw
rect 6084 -1088 6101 -1063
rect 6225 -1088 6242 -1056
rect 6424 -1088 6439 -1046
rect -233 -1126 -201 -1112
rect 347 -1126 379 -1112
rect 927 -1126 959 -1112
rect 1507 -1126 1539 -1112
rect 2087 -1126 2119 -1112
rect 2667 -1126 2699 -1112
rect 3247 -1126 3279 -1112
rect 3827 -1126 3859 -1112
rect 4407 -1126 4439 -1112
rect 4987 -1126 5019 -1112
rect 5567 -1126 5599 -1112
rect 6147 -1126 6179 -1112
rect -419 -1212 -404 -1184
rect -338 -1212 -323 -1184
rect -111 -1212 -96 -1184
rect -29 -1212 -14 -1183
rect 161 -1212 176 -1184
rect 242 -1212 257 -1184
rect 469 -1212 484 -1184
rect 551 -1212 566 -1183
rect 741 -1212 756 -1184
rect 822 -1212 837 -1184
rect 1049 -1212 1064 -1184
rect 1131 -1212 1146 -1183
rect 1321 -1212 1336 -1184
rect 1402 -1212 1417 -1184
rect 1629 -1212 1644 -1184
rect 1711 -1212 1726 -1183
rect 1901 -1212 1916 -1184
rect 1982 -1212 1997 -1184
rect 2209 -1212 2224 -1184
rect 2291 -1212 2306 -1183
rect 2481 -1212 2496 -1184
rect 2562 -1212 2577 -1184
rect 2789 -1212 2804 -1184
rect 2871 -1212 2886 -1183
rect 3061 -1212 3076 -1184
rect 3142 -1212 3157 -1184
rect 3369 -1212 3384 -1184
rect 3451 -1212 3466 -1183
rect 3641 -1212 3656 -1184
rect 3722 -1212 3737 -1184
rect 3949 -1212 3964 -1184
rect 4031 -1212 4046 -1183
rect 4221 -1212 4236 -1184
rect 4302 -1212 4317 -1184
rect 4529 -1212 4544 -1184
rect 4611 -1212 4626 -1183
rect 4801 -1212 4816 -1184
rect 4882 -1212 4897 -1184
rect 5109 -1212 5124 -1184
rect 5191 -1212 5206 -1183
rect 5381 -1212 5396 -1184
rect 5462 -1212 5477 -1184
rect 5689 -1212 5704 -1184
rect 5771 -1212 5786 -1183
rect 5961 -1212 5976 -1184
rect 6042 -1212 6057 -1184
rect 6269 -1212 6284 -1184
rect 6351 -1212 6366 -1183
rect -493 -1358 -478 -1316
rect -296 -1333 -286 -1326
tri -286 -1333 -279 -1326 sw
rect -296 -1358 -279 -1333
rect -155 -1358 -138 -1326
rect 44 -1358 59 -1316
rect 87 -1358 102 -1316
rect 284 -1333 294 -1326
tri 294 -1333 301 -1326 sw
rect 284 -1358 301 -1333
rect 425 -1358 442 -1326
rect 624 -1358 639 -1316
rect 667 -1358 682 -1316
rect 864 -1333 874 -1326
tri 874 -1333 881 -1326 sw
rect 864 -1358 881 -1333
rect 1005 -1358 1022 -1326
rect 1204 -1358 1219 -1316
rect 1247 -1358 1262 -1316
rect 1444 -1333 1454 -1326
tri 1454 -1333 1461 -1326 sw
rect 1444 -1358 1461 -1333
rect 1585 -1358 1602 -1326
rect 1784 -1358 1799 -1316
rect 1827 -1358 1842 -1316
rect 2024 -1333 2034 -1326
tri 2034 -1333 2041 -1326 sw
rect 2024 -1358 2041 -1333
rect 2165 -1358 2182 -1326
rect 2364 -1358 2379 -1316
rect 2407 -1358 2422 -1316
rect 2604 -1333 2614 -1326
tri 2614 -1333 2621 -1326 sw
rect 2604 -1358 2621 -1333
rect 2745 -1358 2762 -1326
rect 2944 -1358 2959 -1316
rect 2987 -1358 3002 -1316
rect 3184 -1333 3194 -1326
tri 3194 -1333 3201 -1326 sw
rect 3184 -1358 3201 -1333
rect 3325 -1358 3342 -1326
rect 3524 -1358 3539 -1316
rect 3567 -1358 3582 -1316
rect 3764 -1333 3774 -1326
tri 3774 -1333 3781 -1326 sw
rect 3764 -1358 3781 -1333
rect 3905 -1358 3922 -1326
rect 4104 -1358 4119 -1316
rect 4147 -1358 4162 -1316
rect 4344 -1333 4354 -1326
tri 4354 -1333 4361 -1326 sw
rect 4344 -1358 4361 -1333
rect 4485 -1358 4502 -1326
rect 4684 -1358 4699 -1316
rect 4727 -1358 4742 -1316
rect 4924 -1333 4934 -1326
tri 4934 -1333 4941 -1326 sw
rect 4924 -1358 4941 -1333
rect 5065 -1358 5082 -1326
rect 5264 -1358 5279 -1316
rect 5307 -1358 5322 -1316
rect 5504 -1333 5514 -1326
tri 5514 -1333 5521 -1326 sw
rect 5504 -1358 5521 -1333
rect 5645 -1358 5662 -1326
rect 5844 -1358 5859 -1316
rect 5887 -1358 5902 -1316
rect 6084 -1333 6094 -1326
tri 6094 -1333 6101 -1326 sw
rect 6084 -1358 6101 -1333
rect 6225 -1358 6242 -1326
rect 6424 -1358 6439 -1316
rect -233 -1396 -201 -1382
rect 347 -1396 379 -1382
rect 927 -1396 959 -1382
rect 1507 -1396 1539 -1382
rect 2087 -1396 2119 -1382
rect 2667 -1396 2699 -1382
rect 3247 -1396 3279 -1382
rect 3827 -1396 3859 -1382
rect 4407 -1396 4439 -1382
rect 4987 -1396 5019 -1382
rect 5567 -1396 5599 -1382
rect 6147 -1396 6179 -1382
rect -419 -1482 -404 -1454
rect -338 -1482 -323 -1454
rect -111 -1482 -96 -1454
rect -29 -1482 -14 -1453
rect 161 -1482 176 -1454
rect 242 -1482 257 -1454
rect 469 -1482 484 -1454
rect 551 -1482 566 -1453
rect 741 -1482 756 -1454
rect 822 -1482 837 -1454
rect 1049 -1482 1064 -1454
rect 1131 -1482 1146 -1453
rect 1321 -1482 1336 -1454
rect 1402 -1482 1417 -1454
rect 1629 -1482 1644 -1454
rect 1711 -1482 1726 -1453
rect 1901 -1482 1916 -1454
rect 1982 -1482 1997 -1454
rect 2209 -1482 2224 -1454
rect 2291 -1482 2306 -1453
rect 2481 -1482 2496 -1454
rect 2562 -1482 2577 -1454
rect 2789 -1482 2804 -1454
rect 2871 -1482 2886 -1453
rect 3061 -1482 3076 -1454
rect 3142 -1482 3157 -1454
rect 3369 -1482 3384 -1454
rect 3451 -1482 3466 -1453
rect 3641 -1482 3656 -1454
rect 3722 -1482 3737 -1454
rect 3949 -1482 3964 -1454
rect 4031 -1482 4046 -1453
rect 4221 -1482 4236 -1454
rect 4302 -1482 4317 -1454
rect 4529 -1482 4544 -1454
rect 4611 -1482 4626 -1453
rect 4801 -1482 4816 -1454
rect 4882 -1482 4897 -1454
rect 5109 -1482 5124 -1454
rect 5191 -1482 5206 -1453
rect 5381 -1482 5396 -1454
rect 5462 -1482 5477 -1454
rect 5689 -1482 5704 -1454
rect 5771 -1482 5786 -1453
rect 5961 -1482 5976 -1454
rect 6042 -1482 6057 -1454
rect 6269 -1482 6284 -1454
rect 6351 -1482 6366 -1453
rect -493 -1628 -478 -1586
rect -296 -1603 -286 -1596
tri -286 -1603 -279 -1596 sw
rect -296 -1628 -279 -1603
rect -155 -1628 -138 -1596
rect 44 -1628 59 -1586
rect 87 -1628 102 -1586
rect 284 -1603 294 -1596
tri 294 -1603 301 -1596 sw
rect 284 -1628 301 -1603
rect 425 -1628 442 -1596
rect 624 -1628 639 -1586
rect 667 -1628 682 -1586
rect 864 -1603 874 -1596
tri 874 -1603 881 -1596 sw
rect 864 -1628 881 -1603
rect 1005 -1628 1022 -1596
rect 1204 -1628 1219 -1586
rect 1247 -1628 1262 -1586
rect 1444 -1603 1454 -1596
tri 1454 -1603 1461 -1596 sw
rect 1444 -1628 1461 -1603
rect 1585 -1628 1602 -1596
rect 1784 -1628 1799 -1586
rect 1827 -1628 1842 -1586
rect 2024 -1603 2034 -1596
tri 2034 -1603 2041 -1596 sw
rect 2024 -1628 2041 -1603
rect 2165 -1628 2182 -1596
rect 2364 -1628 2379 -1586
rect 2407 -1628 2422 -1586
rect 2604 -1603 2614 -1596
tri 2614 -1603 2621 -1596 sw
rect 2604 -1628 2621 -1603
rect 2745 -1628 2762 -1596
rect 2944 -1628 2959 -1586
rect 2987 -1628 3002 -1586
rect 3184 -1603 3194 -1596
tri 3194 -1603 3201 -1596 sw
rect 3184 -1628 3201 -1603
rect 3325 -1628 3342 -1596
rect 3524 -1628 3539 -1586
rect 3567 -1628 3582 -1586
rect 3764 -1603 3774 -1596
tri 3774 -1603 3781 -1596 sw
rect 3764 -1628 3781 -1603
rect 3905 -1628 3922 -1596
rect 4104 -1628 4119 -1586
rect 4147 -1628 4162 -1586
rect 4344 -1603 4354 -1596
tri 4354 -1603 4361 -1596 sw
rect 4344 -1628 4361 -1603
rect 4485 -1628 4502 -1596
rect 4684 -1628 4699 -1586
rect 4727 -1628 4742 -1586
rect 4924 -1603 4934 -1596
tri 4934 -1603 4941 -1596 sw
rect 4924 -1628 4941 -1603
rect 5065 -1628 5082 -1596
rect 5264 -1628 5279 -1586
rect 5307 -1628 5322 -1586
rect 5504 -1603 5514 -1596
tri 5514 -1603 5521 -1596 sw
rect 5504 -1628 5521 -1603
rect 5645 -1628 5662 -1596
rect 5844 -1628 5859 -1586
rect 5887 -1628 5902 -1586
rect 6084 -1603 6094 -1596
tri 6094 -1603 6101 -1596 sw
rect 6084 -1628 6101 -1603
rect 6225 -1628 6242 -1596
rect 6424 -1628 6439 -1586
rect -233 -1666 -201 -1652
rect 347 -1666 379 -1652
rect 927 -1666 959 -1652
rect 1507 -1666 1539 -1652
rect 2087 -1666 2119 -1652
rect 2667 -1666 2699 -1652
rect 3247 -1666 3279 -1652
rect 3827 -1666 3859 -1652
rect 4407 -1666 4439 -1652
rect 4987 -1666 5019 -1652
rect 5567 -1666 5599 -1652
rect 6147 -1666 6179 -1652
rect -419 -1752 -404 -1724
rect -338 -1752 -323 -1724
rect -111 -1752 -96 -1724
rect -29 -1752 -14 -1723
rect 161 -1752 176 -1724
rect 242 -1752 257 -1724
rect 469 -1752 484 -1724
rect 551 -1752 566 -1723
rect 741 -1752 756 -1724
rect 822 -1752 837 -1724
rect 1049 -1752 1064 -1724
rect 1131 -1752 1146 -1723
rect 1321 -1752 1336 -1724
rect 1402 -1752 1417 -1724
rect 1629 -1752 1644 -1724
rect 1711 -1752 1726 -1723
rect 1901 -1752 1916 -1724
rect 1982 -1752 1997 -1724
rect 2209 -1752 2224 -1724
rect 2291 -1752 2306 -1723
rect 2481 -1752 2496 -1724
rect 2562 -1752 2577 -1724
rect 2789 -1752 2804 -1724
rect 2871 -1752 2886 -1723
rect 3061 -1752 3076 -1724
rect 3142 -1752 3157 -1724
rect 3369 -1752 3384 -1724
rect 3451 -1752 3466 -1723
rect 3641 -1752 3656 -1724
rect 3722 -1752 3737 -1724
rect 3949 -1752 3964 -1724
rect 4031 -1752 4046 -1723
rect 4221 -1752 4236 -1724
rect 4302 -1752 4317 -1724
rect 4529 -1752 4544 -1724
rect 4611 -1752 4626 -1723
rect 4801 -1752 4816 -1724
rect 4882 -1752 4897 -1724
rect 5109 -1752 5124 -1724
rect 5191 -1752 5206 -1723
rect 5381 -1752 5396 -1724
rect 5462 -1752 5477 -1724
rect 5689 -1752 5704 -1724
rect 5771 -1752 5786 -1723
rect 5961 -1752 5976 -1724
rect 6042 -1752 6057 -1724
rect 6269 -1752 6284 -1724
rect 6351 -1752 6366 -1723
rect -493 -1898 -478 -1856
rect -296 -1873 -286 -1866
tri -286 -1873 -279 -1866 sw
rect -296 -1898 -279 -1873
rect -155 -1898 -138 -1866
rect 44 -1898 59 -1856
rect 87 -1898 102 -1856
rect 284 -1873 294 -1866
tri 294 -1873 301 -1866 sw
rect 284 -1898 301 -1873
rect 425 -1898 442 -1866
rect 624 -1898 639 -1856
rect 667 -1898 682 -1856
rect 864 -1873 874 -1866
tri 874 -1873 881 -1866 sw
rect 864 -1898 881 -1873
rect 1005 -1898 1022 -1866
rect 1204 -1898 1219 -1856
rect 1247 -1898 1262 -1856
rect 1444 -1873 1454 -1866
tri 1454 -1873 1461 -1866 sw
rect 1444 -1898 1461 -1873
rect 1585 -1898 1602 -1866
rect 1784 -1898 1799 -1856
rect 1827 -1898 1842 -1856
rect 2024 -1873 2034 -1866
tri 2034 -1873 2041 -1866 sw
rect 2024 -1898 2041 -1873
rect 2165 -1898 2182 -1866
rect 2364 -1898 2379 -1856
rect 2407 -1898 2422 -1856
rect 2604 -1873 2614 -1866
tri 2614 -1873 2621 -1866 sw
rect 2604 -1898 2621 -1873
rect 2745 -1898 2762 -1866
rect 2944 -1898 2959 -1856
rect 2987 -1898 3002 -1856
rect 3184 -1873 3194 -1866
tri 3194 -1873 3201 -1866 sw
rect 3184 -1898 3201 -1873
rect 3325 -1898 3342 -1866
rect 3524 -1898 3539 -1856
rect 3567 -1898 3582 -1856
rect 3764 -1873 3774 -1866
tri 3774 -1873 3781 -1866 sw
rect 3764 -1898 3781 -1873
rect 3905 -1898 3922 -1866
rect 4104 -1898 4119 -1856
rect 4147 -1898 4162 -1856
rect 4344 -1873 4354 -1866
tri 4354 -1873 4361 -1866 sw
rect 4344 -1898 4361 -1873
rect 4485 -1898 4502 -1866
rect 4684 -1898 4699 -1856
rect 4727 -1898 4742 -1856
rect 4924 -1873 4934 -1866
tri 4934 -1873 4941 -1866 sw
rect 4924 -1898 4941 -1873
rect 5065 -1898 5082 -1866
rect 5264 -1898 5279 -1856
rect 5307 -1898 5322 -1856
rect 5504 -1873 5514 -1866
tri 5514 -1873 5521 -1866 sw
rect 5504 -1898 5521 -1873
rect 5645 -1898 5662 -1866
rect 5844 -1898 5859 -1856
rect 5887 -1898 5902 -1856
rect 6084 -1873 6094 -1866
tri 6094 -1873 6101 -1866 sw
rect 6084 -1898 6101 -1873
rect 6225 -1898 6242 -1866
rect 6424 -1898 6439 -1856
rect -233 -1936 -201 -1922
rect 347 -1936 379 -1922
rect 927 -1936 959 -1922
rect 1507 -1936 1539 -1922
rect 2087 -1936 2119 -1922
rect 2667 -1936 2699 -1922
rect 3247 -1936 3279 -1922
rect 3827 -1936 3859 -1922
rect 4407 -1936 4439 -1922
rect 4987 -1936 5019 -1922
rect 5567 -1936 5599 -1922
rect 6147 -1936 6179 -1922
rect -419 -2022 -404 -1994
rect -338 -2022 -323 -1994
rect -111 -2022 -96 -1994
rect -29 -2022 -14 -1993
rect 161 -2022 176 -1994
rect 242 -2022 257 -1994
rect 469 -2022 484 -1994
rect 551 -2022 566 -1993
rect 741 -2022 756 -1994
rect 822 -2022 837 -1994
rect 1049 -2022 1064 -1994
rect 1131 -2022 1146 -1993
rect 1321 -2022 1336 -1994
rect 1402 -2022 1417 -1994
rect 1629 -2022 1644 -1994
rect 1711 -2022 1726 -1993
rect 1901 -2022 1916 -1994
rect 1982 -2022 1997 -1994
rect 2209 -2022 2224 -1994
rect 2291 -2022 2306 -1993
rect 2481 -2022 2496 -1994
rect 2562 -2022 2577 -1994
rect 2789 -2022 2804 -1994
rect 2871 -2022 2886 -1993
rect 3061 -2022 3076 -1994
rect 3142 -2022 3157 -1994
rect 3369 -2022 3384 -1994
rect 3451 -2022 3466 -1993
rect 3641 -2022 3656 -1994
rect 3722 -2022 3737 -1994
rect 3949 -2022 3964 -1994
rect 4031 -2022 4046 -1993
rect 4221 -2022 4236 -1994
rect 4302 -2022 4317 -1994
rect 4529 -2022 4544 -1994
rect 4611 -2022 4626 -1993
rect 4801 -2022 4816 -1994
rect 4882 -2022 4897 -1994
rect 5109 -2022 5124 -1994
rect 5191 -2022 5206 -1993
rect 5381 -2022 5396 -1994
rect 5462 -2022 5477 -1994
rect 5689 -2022 5704 -1994
rect 5771 -2022 5786 -1993
rect 5961 -2022 5976 -1994
rect 6042 -2022 6057 -1994
rect 6269 -2022 6284 -1994
rect 6351 -2022 6366 -1993
rect -493 -2168 -478 -2126
rect -296 -2143 -286 -2136
tri -286 -2143 -279 -2136 sw
rect -296 -2168 -279 -2143
rect -155 -2168 -138 -2136
rect 44 -2168 59 -2126
rect 87 -2168 102 -2126
rect 284 -2143 294 -2136
tri 294 -2143 301 -2136 sw
rect 284 -2168 301 -2143
rect 425 -2168 442 -2136
rect 624 -2168 639 -2126
rect 667 -2168 682 -2126
rect 864 -2143 874 -2136
tri 874 -2143 881 -2136 sw
rect 864 -2168 881 -2143
rect 1005 -2168 1022 -2136
rect 1204 -2168 1219 -2126
rect 1247 -2168 1262 -2126
rect 1444 -2143 1454 -2136
tri 1454 -2143 1461 -2136 sw
rect 1444 -2168 1461 -2143
rect 1585 -2168 1602 -2136
rect 1784 -2168 1799 -2126
rect 1827 -2168 1842 -2126
rect 2024 -2143 2034 -2136
tri 2034 -2143 2041 -2136 sw
rect 2024 -2168 2041 -2143
rect 2165 -2168 2182 -2136
rect 2364 -2168 2379 -2126
rect 2407 -2168 2422 -2126
rect 2604 -2143 2614 -2136
tri 2614 -2143 2621 -2136 sw
rect 2604 -2168 2621 -2143
rect 2745 -2168 2762 -2136
rect 2944 -2168 2959 -2126
rect 2987 -2168 3002 -2126
rect 3184 -2143 3194 -2136
tri 3194 -2143 3201 -2136 sw
rect 3184 -2168 3201 -2143
rect 3325 -2168 3342 -2136
rect 3524 -2168 3539 -2126
rect 3567 -2168 3582 -2126
rect 3764 -2143 3774 -2136
tri 3774 -2143 3781 -2136 sw
rect 3764 -2168 3781 -2143
rect 3905 -2168 3922 -2136
rect 4104 -2168 4119 -2126
rect 4147 -2168 4162 -2126
rect 4344 -2143 4354 -2136
tri 4354 -2143 4361 -2136 sw
rect 4344 -2168 4361 -2143
rect 4485 -2168 4502 -2136
rect 4684 -2168 4699 -2126
rect 4727 -2168 4742 -2126
rect 4924 -2143 4934 -2136
tri 4934 -2143 4941 -2136 sw
rect 4924 -2168 4941 -2143
rect 5065 -2168 5082 -2136
rect 5264 -2168 5279 -2126
rect 5307 -2168 5322 -2126
rect 5504 -2143 5514 -2136
tri 5514 -2143 5521 -2136 sw
rect 5504 -2168 5521 -2143
rect 5645 -2168 5662 -2136
rect 5844 -2168 5859 -2126
rect 5887 -2168 5902 -2126
rect 6084 -2143 6094 -2136
tri 6094 -2143 6101 -2136 sw
rect 6084 -2168 6101 -2143
rect 6225 -2168 6242 -2136
rect 6424 -2168 6439 -2126
rect -233 -2206 -201 -2192
rect 347 -2206 379 -2192
rect 927 -2206 959 -2192
rect 1507 -2206 1539 -2192
rect 2087 -2206 2119 -2192
rect 2667 -2206 2699 -2192
rect 3247 -2206 3279 -2192
rect 3827 -2206 3859 -2192
rect 4407 -2206 4439 -2192
rect 4987 -2206 5019 -2192
rect 5567 -2206 5599 -2192
rect 6147 -2206 6179 -2192
rect -419 -2292 -404 -2264
rect -338 -2292 -323 -2264
rect -111 -2292 -96 -2264
rect -29 -2292 -14 -2263
rect 161 -2292 176 -2264
rect 242 -2292 257 -2264
rect 469 -2292 484 -2264
rect 551 -2292 566 -2263
rect 741 -2292 756 -2264
rect 822 -2292 837 -2264
rect 1049 -2292 1064 -2264
rect 1131 -2292 1146 -2263
rect 1321 -2292 1336 -2264
rect 1402 -2292 1417 -2264
rect 1629 -2292 1644 -2264
rect 1711 -2292 1726 -2263
rect 1901 -2292 1916 -2264
rect 1982 -2292 1997 -2264
rect 2209 -2292 2224 -2264
rect 2291 -2292 2306 -2263
rect 2481 -2292 2496 -2264
rect 2562 -2292 2577 -2264
rect 2789 -2292 2804 -2264
rect 2871 -2292 2886 -2263
rect 3061 -2292 3076 -2264
rect 3142 -2292 3157 -2264
rect 3369 -2292 3384 -2264
rect 3451 -2292 3466 -2263
rect 3641 -2292 3656 -2264
rect 3722 -2292 3737 -2264
rect 3949 -2292 3964 -2264
rect 4031 -2292 4046 -2263
rect 4221 -2292 4236 -2264
rect 4302 -2292 4317 -2264
rect 4529 -2292 4544 -2264
rect 4611 -2292 4626 -2263
rect 4801 -2292 4816 -2264
rect 4882 -2292 4897 -2264
rect 5109 -2292 5124 -2264
rect 5191 -2292 5206 -2263
rect 5381 -2292 5396 -2264
rect 5462 -2292 5477 -2264
rect 5689 -2292 5704 -2264
rect 5771 -2292 5786 -2263
rect 5961 -2292 5976 -2264
rect 6042 -2292 6057 -2264
rect 6269 -2292 6284 -2264
rect 6351 -2292 6366 -2263
rect -493 -2438 -478 -2396
rect -296 -2413 -286 -2406
tri -286 -2413 -279 -2406 sw
rect -296 -2438 -279 -2413
rect -155 -2438 -138 -2406
rect 44 -2438 59 -2396
rect 87 -2438 102 -2396
rect 284 -2413 294 -2406
tri 294 -2413 301 -2406 sw
rect 284 -2438 301 -2413
rect 425 -2438 442 -2406
rect 624 -2438 639 -2396
rect 667 -2438 682 -2396
rect 864 -2413 874 -2406
tri 874 -2413 881 -2406 sw
rect 864 -2438 881 -2413
rect 1005 -2438 1022 -2406
rect 1204 -2438 1219 -2396
rect 1247 -2438 1262 -2396
rect 1444 -2413 1454 -2406
tri 1454 -2413 1461 -2406 sw
rect 1444 -2438 1461 -2413
rect 1585 -2438 1602 -2406
rect 1784 -2438 1799 -2396
rect 1827 -2438 1842 -2396
rect 2024 -2413 2034 -2406
tri 2034 -2413 2041 -2406 sw
rect 2024 -2438 2041 -2413
rect 2165 -2438 2182 -2406
rect 2364 -2438 2379 -2396
rect 2407 -2438 2422 -2396
rect 2604 -2413 2614 -2406
tri 2614 -2413 2621 -2406 sw
rect 2604 -2438 2621 -2413
rect 2745 -2438 2762 -2406
rect 2944 -2438 2959 -2396
rect 2987 -2438 3002 -2396
rect 3184 -2413 3194 -2406
tri 3194 -2413 3201 -2406 sw
rect 3184 -2438 3201 -2413
rect 3325 -2438 3342 -2406
rect 3524 -2438 3539 -2396
rect 3567 -2438 3582 -2396
rect 3764 -2413 3774 -2406
tri 3774 -2413 3781 -2406 sw
rect 3764 -2438 3781 -2413
rect 3905 -2438 3922 -2406
rect 4104 -2438 4119 -2396
rect 4147 -2438 4162 -2396
rect 4344 -2413 4354 -2406
tri 4354 -2413 4361 -2406 sw
rect 4344 -2438 4361 -2413
rect 4485 -2438 4502 -2406
rect 4684 -2438 4699 -2396
rect 4727 -2438 4742 -2396
rect 4924 -2413 4934 -2406
tri 4934 -2413 4941 -2406 sw
rect 4924 -2438 4941 -2413
rect 5065 -2438 5082 -2406
rect 5264 -2438 5279 -2396
rect 5307 -2438 5322 -2396
rect 5504 -2413 5514 -2406
tri 5514 -2413 5521 -2406 sw
rect 5504 -2438 5521 -2413
rect 5645 -2438 5662 -2406
rect 5844 -2438 5859 -2396
rect 5887 -2438 5902 -2396
rect 6084 -2413 6094 -2406
tri 6094 -2413 6101 -2406 sw
rect 6084 -2438 6101 -2413
rect 6225 -2438 6242 -2406
rect 6424 -2438 6439 -2396
rect -233 -2476 -201 -2462
rect 347 -2476 379 -2462
rect 927 -2476 959 -2462
rect 1507 -2476 1539 -2462
rect 2087 -2476 2119 -2462
rect 2667 -2476 2699 -2462
rect 3247 -2476 3279 -2462
rect 3827 -2476 3859 -2462
rect 4407 -2476 4439 -2462
rect 4987 -2476 5019 -2462
rect 5567 -2476 5599 -2462
rect 6147 -2476 6179 -2462
<< pdiffc >>
rect -233 1800 -201 1814
rect -295 1748 -280 1776
rect -154 1760 -142 1776
tri -154 1748 -142 1760 ne
rect 347 1800 379 1814
rect 285 1748 300 1776
rect 426 1760 438 1776
tri 426 1748 438 1760 ne
rect 927 1800 959 1814
rect 865 1748 880 1776
rect 1006 1760 1018 1776
tri 1006 1748 1018 1760 ne
rect 1507 1800 1539 1814
rect 1445 1748 1460 1776
rect 1586 1760 1598 1776
tri 1586 1748 1598 1760 ne
rect 2087 1800 2119 1814
rect 2025 1748 2040 1776
rect 2166 1760 2178 1776
tri 2166 1748 2178 1760 ne
rect 2667 1800 2699 1814
rect 2605 1748 2620 1776
rect 2746 1760 2758 1776
tri 2746 1748 2758 1760 ne
rect 3247 1800 3279 1814
rect 3185 1748 3200 1776
rect 3326 1760 3338 1776
tri 3326 1748 3338 1760 ne
rect 3827 1800 3859 1814
rect 3765 1748 3780 1776
rect 3906 1760 3918 1776
tri 3906 1748 3918 1760 ne
rect 4407 1800 4439 1814
rect 4345 1748 4360 1776
rect 4486 1760 4498 1776
tri 4486 1748 4498 1760 ne
rect 4987 1800 5019 1814
rect 4925 1748 4940 1776
rect 5066 1760 5078 1776
tri 5066 1748 5078 1760 ne
rect 5567 1800 5599 1814
rect 5505 1748 5520 1776
rect 5646 1760 5658 1776
tri 5646 1748 5658 1760 ne
rect 6147 1800 6179 1814
rect 6085 1748 6100 1776
rect 6226 1760 6238 1776
tri 6226 1748 6238 1760 ne
rect -233 1530 -201 1544
rect -295 1478 -280 1506
rect -154 1490 -142 1506
tri -154 1478 -142 1490 ne
rect 347 1530 379 1544
rect 285 1478 300 1506
rect 426 1490 438 1506
tri 426 1478 438 1490 ne
rect 927 1530 959 1544
rect 865 1478 880 1506
rect 1006 1490 1018 1506
tri 1006 1478 1018 1490 ne
rect 1507 1530 1539 1544
rect 1445 1478 1460 1506
rect 1586 1490 1598 1506
tri 1586 1478 1598 1490 ne
rect 2087 1530 2119 1544
rect 2025 1478 2040 1506
rect 2166 1490 2178 1506
tri 2166 1478 2178 1490 ne
rect 2667 1530 2699 1544
rect 2605 1478 2620 1506
rect 2746 1490 2758 1506
tri 2746 1478 2758 1490 ne
rect 3247 1530 3279 1544
rect 3185 1478 3200 1506
rect 3326 1490 3338 1506
tri 3326 1478 3338 1490 ne
rect 3827 1530 3859 1544
rect 3765 1478 3780 1506
rect 3906 1490 3918 1506
tri 3906 1478 3918 1490 ne
rect 4407 1530 4439 1544
rect 4345 1478 4360 1506
rect 4486 1490 4498 1506
tri 4486 1478 4498 1490 ne
rect 4987 1530 5019 1544
rect 4925 1478 4940 1506
rect 5066 1490 5078 1506
tri 5066 1478 5078 1490 ne
rect 5567 1530 5599 1544
rect 5505 1478 5520 1506
rect 5646 1490 5658 1506
tri 5646 1478 5658 1490 ne
rect 6147 1530 6179 1544
rect 6085 1478 6100 1506
rect 6226 1490 6238 1506
tri 6226 1478 6238 1490 ne
rect -233 1260 -201 1274
rect -295 1208 -280 1236
rect -154 1220 -142 1236
tri -154 1208 -142 1220 ne
rect 347 1260 379 1274
rect 285 1208 300 1236
rect 426 1220 438 1236
tri 426 1208 438 1220 ne
rect 927 1260 959 1274
rect 865 1208 880 1236
rect 1006 1220 1018 1236
tri 1006 1208 1018 1220 ne
rect 1507 1260 1539 1274
rect 1445 1208 1460 1236
rect 1586 1220 1598 1236
tri 1586 1208 1598 1220 ne
rect 2087 1260 2119 1274
rect 2025 1208 2040 1236
rect 2166 1220 2178 1236
tri 2166 1208 2178 1220 ne
rect 2667 1260 2699 1274
rect 2605 1208 2620 1236
rect 2746 1220 2758 1236
tri 2746 1208 2758 1220 ne
rect 3247 1260 3279 1274
rect 3185 1208 3200 1236
rect 3326 1220 3338 1236
tri 3326 1208 3338 1220 ne
rect 3827 1260 3859 1274
rect 3765 1208 3780 1236
rect 3906 1220 3918 1236
tri 3906 1208 3918 1220 ne
rect 4407 1260 4439 1274
rect 4345 1208 4360 1236
rect 4486 1220 4498 1236
tri 4486 1208 4498 1220 ne
rect 4987 1260 5019 1274
rect 4925 1208 4940 1236
rect 5066 1220 5078 1236
tri 5066 1208 5078 1220 ne
rect 5567 1260 5599 1274
rect 5505 1208 5520 1236
rect 5646 1220 5658 1236
tri 5646 1208 5658 1220 ne
rect 6147 1260 6179 1274
rect 6085 1208 6100 1236
rect 6226 1220 6238 1236
tri 6226 1208 6238 1220 ne
rect -233 990 -201 1004
rect -295 938 -280 966
rect -154 950 -142 966
tri -154 938 -142 950 ne
rect 347 990 379 1004
rect 285 938 300 966
rect 426 950 438 966
tri 426 938 438 950 ne
rect 927 990 959 1004
rect 865 938 880 966
rect 1006 950 1018 966
tri 1006 938 1018 950 ne
rect 1507 990 1539 1004
rect 1445 938 1460 966
rect 1586 950 1598 966
tri 1586 938 1598 950 ne
rect 2087 990 2119 1004
rect 2025 938 2040 966
rect 2166 950 2178 966
tri 2166 938 2178 950 ne
rect 2667 990 2699 1004
rect 2605 938 2620 966
rect 2746 950 2758 966
tri 2746 938 2758 950 ne
rect 3247 990 3279 1004
rect 3185 938 3200 966
rect 3326 950 3338 966
tri 3326 938 3338 950 ne
rect 3827 990 3859 1004
rect 3765 938 3780 966
rect 3906 950 3918 966
tri 3906 938 3918 950 ne
rect 4407 990 4439 1004
rect 4345 938 4360 966
rect 4486 950 4498 966
tri 4486 938 4498 950 ne
rect 4987 990 5019 1004
rect 4925 938 4940 966
rect 5066 950 5078 966
tri 5066 938 5078 950 ne
rect 5567 990 5599 1004
rect 5505 938 5520 966
rect 5646 950 5658 966
tri 5646 938 5658 950 ne
rect 6147 990 6179 1004
rect 6085 938 6100 966
rect 6226 950 6238 966
tri 6226 938 6238 950 ne
rect -233 720 -201 734
rect -295 668 -280 696
rect -154 680 -142 696
tri -154 668 -142 680 ne
rect 347 720 379 734
rect 285 668 300 696
rect 426 680 438 696
tri 426 668 438 680 ne
rect 927 720 959 734
rect 865 668 880 696
rect 1006 680 1018 696
tri 1006 668 1018 680 ne
rect 1507 720 1539 734
rect 1445 668 1460 696
rect 1586 680 1598 696
tri 1586 668 1598 680 ne
rect 2087 720 2119 734
rect 2025 668 2040 696
rect 2166 680 2178 696
tri 2166 668 2178 680 ne
rect 2667 720 2699 734
rect 2605 668 2620 696
rect 2746 680 2758 696
tri 2746 668 2758 680 ne
rect 3247 720 3279 734
rect 3185 668 3200 696
rect 3326 680 3338 696
tri 3326 668 3338 680 ne
rect 3827 720 3859 734
rect 3765 668 3780 696
rect 3906 680 3918 696
tri 3906 668 3918 680 ne
rect 4407 720 4439 734
rect 4345 668 4360 696
rect 4486 680 4498 696
tri 4486 668 4498 680 ne
rect 4987 720 5019 734
rect 4925 668 4940 696
rect 5066 680 5078 696
tri 5066 668 5078 680 ne
rect 5567 720 5599 734
rect 5505 668 5520 696
rect 5646 680 5658 696
tri 5646 668 5658 680 ne
rect 6147 720 6179 734
rect 6085 668 6100 696
rect 6226 680 6238 696
tri 6226 668 6238 680 ne
rect -233 450 -201 464
rect -295 398 -280 426
rect -154 410 -142 426
tri -154 398 -142 410 ne
rect 347 450 379 464
rect 285 398 300 426
rect 426 410 438 426
tri 426 398 438 410 ne
rect 927 450 959 464
rect 865 398 880 426
rect 1006 410 1018 426
tri 1006 398 1018 410 ne
rect 1507 450 1539 464
rect 1445 398 1460 426
rect 1586 410 1598 426
tri 1586 398 1598 410 ne
rect 2087 450 2119 464
rect 2025 398 2040 426
rect 2166 410 2178 426
tri 2166 398 2178 410 ne
rect 2667 450 2699 464
rect 2605 398 2620 426
rect 2746 410 2758 426
tri 2746 398 2758 410 ne
rect 3247 450 3279 464
rect 3185 398 3200 426
rect 3326 410 3338 426
tri 3326 398 3338 410 ne
rect 3827 450 3859 464
rect 3765 398 3780 426
rect 3906 410 3918 426
tri 3906 398 3918 410 ne
rect 4407 450 4439 464
rect 4345 398 4360 426
rect 4486 410 4498 426
tri 4486 398 4498 410 ne
rect 4987 450 5019 464
rect 4925 398 4940 426
rect 5066 410 5078 426
tri 5066 398 5078 410 ne
rect 5567 450 5599 464
rect 5505 398 5520 426
rect 5646 410 5658 426
tri 5646 398 5658 410 ne
rect 6147 450 6179 464
rect 6085 398 6100 426
rect 6226 410 6238 426
tri 6226 398 6238 410 ne
rect -233 180 -201 194
rect -295 128 -280 156
rect -154 140 -142 156
tri -154 128 -142 140 ne
rect 347 180 379 194
rect 285 128 300 156
rect 426 140 438 156
tri 426 128 438 140 ne
rect 927 180 959 194
rect 865 128 880 156
rect 1006 140 1018 156
tri 1006 128 1018 140 ne
rect 1507 180 1539 194
rect 1445 128 1460 156
rect 1586 140 1598 156
tri 1586 128 1598 140 ne
rect 2087 180 2119 194
rect 2025 128 2040 156
rect 2166 140 2178 156
tri 2166 128 2178 140 ne
rect 2667 180 2699 194
rect 2605 128 2620 156
rect 2746 140 2758 156
tri 2746 128 2758 140 ne
rect 3247 180 3279 194
rect 3185 128 3200 156
rect 3326 140 3338 156
tri 3326 128 3338 140 ne
rect 3827 180 3859 194
rect 3765 128 3780 156
rect 3906 140 3918 156
tri 3906 128 3918 140 ne
rect 4407 180 4439 194
rect 4345 128 4360 156
rect 4486 140 4498 156
tri 4486 128 4498 140 ne
rect 4987 180 5019 194
rect 4925 128 4940 156
rect 5066 140 5078 156
tri 5066 128 5078 140 ne
rect 5567 180 5599 194
rect 5505 128 5520 156
rect 5646 140 5658 156
tri 5646 128 5658 140 ne
rect 6147 180 6179 194
rect 6085 128 6100 156
rect 6226 140 6238 156
tri 6226 128 6238 140 ne
rect -233 -90 -201 -76
rect -295 -142 -280 -114
rect -154 -130 -142 -114
tri -154 -142 -142 -130 ne
rect 347 -90 379 -76
rect 285 -142 300 -114
rect 426 -130 438 -114
tri 426 -142 438 -130 ne
rect 927 -90 959 -76
rect 865 -142 880 -114
rect 1006 -130 1018 -114
tri 1006 -142 1018 -130 ne
rect 1507 -90 1539 -76
rect 1445 -142 1460 -114
rect 1586 -130 1598 -114
tri 1586 -142 1598 -130 ne
rect 2087 -90 2119 -76
rect 2025 -142 2040 -114
rect 2166 -130 2178 -114
tri 2166 -142 2178 -130 ne
rect 2667 -90 2699 -76
rect 2605 -142 2620 -114
rect 2746 -130 2758 -114
tri 2746 -142 2758 -130 ne
rect 3247 -90 3279 -76
rect 3185 -142 3200 -114
rect 3326 -130 3338 -114
tri 3326 -142 3338 -130 ne
rect 3827 -90 3859 -76
rect 3765 -142 3780 -114
rect 3906 -130 3918 -114
tri 3906 -142 3918 -130 ne
rect 4407 -90 4439 -76
rect 4345 -142 4360 -114
rect 4486 -130 4498 -114
tri 4486 -142 4498 -130 ne
rect 4987 -90 5019 -76
rect 4925 -142 4940 -114
rect 5066 -130 5078 -114
tri 5066 -142 5078 -130 ne
rect 5567 -90 5599 -76
rect 5505 -142 5520 -114
rect 5646 -130 5658 -114
tri 5646 -142 5658 -130 ne
rect 6147 -90 6179 -76
rect 6085 -142 6100 -114
rect 6226 -130 6238 -114
tri 6226 -142 6238 -130 ne
rect -233 -360 -201 -346
rect -295 -412 -280 -384
rect -154 -400 -142 -384
tri -154 -412 -142 -400 ne
rect 347 -360 379 -346
rect 285 -412 300 -384
rect 426 -400 438 -384
tri 426 -412 438 -400 ne
rect 927 -360 959 -346
rect 865 -412 880 -384
rect 1006 -400 1018 -384
tri 1006 -412 1018 -400 ne
rect 1507 -360 1539 -346
rect 1445 -412 1460 -384
rect 1586 -400 1598 -384
tri 1586 -412 1598 -400 ne
rect 2087 -360 2119 -346
rect 2025 -412 2040 -384
rect 2166 -400 2178 -384
tri 2166 -412 2178 -400 ne
rect 2667 -360 2699 -346
rect 2605 -412 2620 -384
rect 2746 -400 2758 -384
tri 2746 -412 2758 -400 ne
rect 3247 -360 3279 -346
rect 3185 -412 3200 -384
rect 3326 -400 3338 -384
tri 3326 -412 3338 -400 ne
rect 3827 -360 3859 -346
rect 3765 -412 3780 -384
rect 3906 -400 3918 -384
tri 3906 -412 3918 -400 ne
rect 4407 -360 4439 -346
rect 4345 -412 4360 -384
rect 4486 -400 4498 -384
tri 4486 -412 4498 -400 ne
rect 4987 -360 5019 -346
rect 4925 -412 4940 -384
rect 5066 -400 5078 -384
tri 5066 -412 5078 -400 ne
rect 5567 -360 5599 -346
rect 5505 -412 5520 -384
rect 5646 -400 5658 -384
tri 5646 -412 5658 -400 ne
rect 6147 -360 6179 -346
rect 6085 -412 6100 -384
rect 6226 -400 6238 -384
tri 6226 -412 6238 -400 ne
rect -233 -630 -201 -616
rect -295 -682 -280 -654
rect -154 -670 -142 -654
tri -154 -682 -142 -670 ne
rect 347 -630 379 -616
rect 285 -682 300 -654
rect 426 -670 438 -654
tri 426 -682 438 -670 ne
rect 927 -630 959 -616
rect 865 -682 880 -654
rect 1006 -670 1018 -654
tri 1006 -682 1018 -670 ne
rect 1507 -630 1539 -616
rect 1445 -682 1460 -654
rect 1586 -670 1598 -654
tri 1586 -682 1598 -670 ne
rect 2087 -630 2119 -616
rect 2025 -682 2040 -654
rect 2166 -670 2178 -654
tri 2166 -682 2178 -670 ne
rect 2667 -630 2699 -616
rect 2605 -682 2620 -654
rect 2746 -670 2758 -654
tri 2746 -682 2758 -670 ne
rect 3247 -630 3279 -616
rect 3185 -682 3200 -654
rect 3326 -670 3338 -654
tri 3326 -682 3338 -670 ne
rect 3827 -630 3859 -616
rect 3765 -682 3780 -654
rect 3906 -670 3918 -654
tri 3906 -682 3918 -670 ne
rect 4407 -630 4439 -616
rect 4345 -682 4360 -654
rect 4486 -670 4498 -654
tri 4486 -682 4498 -670 ne
rect 4987 -630 5019 -616
rect 4925 -682 4940 -654
rect 5066 -670 5078 -654
tri 5066 -682 5078 -670 ne
rect 5567 -630 5599 -616
rect 5505 -682 5520 -654
rect 5646 -670 5658 -654
tri 5646 -682 5658 -670 ne
rect 6147 -630 6179 -616
rect 6085 -682 6100 -654
rect 6226 -670 6238 -654
tri 6226 -682 6238 -670 ne
rect -233 -900 -201 -886
rect -295 -952 -280 -924
rect -154 -940 -142 -924
tri -154 -952 -142 -940 ne
rect 347 -900 379 -886
rect 285 -952 300 -924
rect 426 -940 438 -924
tri 426 -952 438 -940 ne
rect 927 -900 959 -886
rect 865 -952 880 -924
rect 1006 -940 1018 -924
tri 1006 -952 1018 -940 ne
rect 1507 -900 1539 -886
rect 1445 -952 1460 -924
rect 1586 -940 1598 -924
tri 1586 -952 1598 -940 ne
rect 2087 -900 2119 -886
rect 2025 -952 2040 -924
rect 2166 -940 2178 -924
tri 2166 -952 2178 -940 ne
rect 2667 -900 2699 -886
rect 2605 -952 2620 -924
rect 2746 -940 2758 -924
tri 2746 -952 2758 -940 ne
rect 3247 -900 3279 -886
rect 3185 -952 3200 -924
rect 3326 -940 3338 -924
tri 3326 -952 3338 -940 ne
rect 3827 -900 3859 -886
rect 3765 -952 3780 -924
rect 3906 -940 3918 -924
tri 3906 -952 3918 -940 ne
rect 4407 -900 4439 -886
rect 4345 -952 4360 -924
rect 4486 -940 4498 -924
tri 4486 -952 4498 -940 ne
rect 4987 -900 5019 -886
rect 4925 -952 4940 -924
rect 5066 -940 5078 -924
tri 5066 -952 5078 -940 ne
rect 5567 -900 5599 -886
rect 5505 -952 5520 -924
rect 5646 -940 5658 -924
tri 5646 -952 5658 -940 ne
rect 6147 -900 6179 -886
rect 6085 -952 6100 -924
rect 6226 -940 6238 -924
tri 6226 -952 6238 -940 ne
rect -233 -1170 -201 -1156
rect -295 -1222 -280 -1194
rect -154 -1210 -142 -1194
tri -154 -1222 -142 -1210 ne
rect 347 -1170 379 -1156
rect 285 -1222 300 -1194
rect 426 -1210 438 -1194
tri 426 -1222 438 -1210 ne
rect 927 -1170 959 -1156
rect 865 -1222 880 -1194
rect 1006 -1210 1018 -1194
tri 1006 -1222 1018 -1210 ne
rect 1507 -1170 1539 -1156
rect 1445 -1222 1460 -1194
rect 1586 -1210 1598 -1194
tri 1586 -1222 1598 -1210 ne
rect 2087 -1170 2119 -1156
rect 2025 -1222 2040 -1194
rect 2166 -1210 2178 -1194
tri 2166 -1222 2178 -1210 ne
rect 2667 -1170 2699 -1156
rect 2605 -1222 2620 -1194
rect 2746 -1210 2758 -1194
tri 2746 -1222 2758 -1210 ne
rect 3247 -1170 3279 -1156
rect 3185 -1222 3200 -1194
rect 3326 -1210 3338 -1194
tri 3326 -1222 3338 -1210 ne
rect 3827 -1170 3859 -1156
rect 3765 -1222 3780 -1194
rect 3906 -1210 3918 -1194
tri 3906 -1222 3918 -1210 ne
rect 4407 -1170 4439 -1156
rect 4345 -1222 4360 -1194
rect 4486 -1210 4498 -1194
tri 4486 -1222 4498 -1210 ne
rect 4987 -1170 5019 -1156
rect 4925 -1222 4940 -1194
rect 5066 -1210 5078 -1194
tri 5066 -1222 5078 -1210 ne
rect 5567 -1170 5599 -1156
rect 5505 -1222 5520 -1194
rect 5646 -1210 5658 -1194
tri 5646 -1222 5658 -1210 ne
rect 6147 -1170 6179 -1156
rect 6085 -1222 6100 -1194
rect 6226 -1210 6238 -1194
tri 6226 -1222 6238 -1210 ne
rect -233 -1440 -201 -1426
rect -295 -1492 -280 -1464
rect -154 -1480 -142 -1464
tri -154 -1492 -142 -1480 ne
rect 347 -1440 379 -1426
rect 285 -1492 300 -1464
rect 426 -1480 438 -1464
tri 426 -1492 438 -1480 ne
rect 927 -1440 959 -1426
rect 865 -1492 880 -1464
rect 1006 -1480 1018 -1464
tri 1006 -1492 1018 -1480 ne
rect 1507 -1440 1539 -1426
rect 1445 -1492 1460 -1464
rect 1586 -1480 1598 -1464
tri 1586 -1492 1598 -1480 ne
rect 2087 -1440 2119 -1426
rect 2025 -1492 2040 -1464
rect 2166 -1480 2178 -1464
tri 2166 -1492 2178 -1480 ne
rect 2667 -1440 2699 -1426
rect 2605 -1492 2620 -1464
rect 2746 -1480 2758 -1464
tri 2746 -1492 2758 -1480 ne
rect 3247 -1440 3279 -1426
rect 3185 -1492 3200 -1464
rect 3326 -1480 3338 -1464
tri 3326 -1492 3338 -1480 ne
rect 3827 -1440 3859 -1426
rect 3765 -1492 3780 -1464
rect 3906 -1480 3918 -1464
tri 3906 -1492 3918 -1480 ne
rect 4407 -1440 4439 -1426
rect 4345 -1492 4360 -1464
rect 4486 -1480 4498 -1464
tri 4486 -1492 4498 -1480 ne
rect 4987 -1440 5019 -1426
rect 4925 -1492 4940 -1464
rect 5066 -1480 5078 -1464
tri 5066 -1492 5078 -1480 ne
rect 5567 -1440 5599 -1426
rect 5505 -1492 5520 -1464
rect 5646 -1480 5658 -1464
tri 5646 -1492 5658 -1480 ne
rect 6147 -1440 6179 -1426
rect 6085 -1492 6100 -1464
rect 6226 -1480 6238 -1464
tri 6226 -1492 6238 -1480 ne
rect -233 -1710 -201 -1696
rect -295 -1762 -280 -1734
rect -154 -1750 -142 -1734
tri -154 -1762 -142 -1750 ne
rect 347 -1710 379 -1696
rect 285 -1762 300 -1734
rect 426 -1750 438 -1734
tri 426 -1762 438 -1750 ne
rect 927 -1710 959 -1696
rect 865 -1762 880 -1734
rect 1006 -1750 1018 -1734
tri 1006 -1762 1018 -1750 ne
rect 1507 -1710 1539 -1696
rect 1445 -1762 1460 -1734
rect 1586 -1750 1598 -1734
tri 1586 -1762 1598 -1750 ne
rect 2087 -1710 2119 -1696
rect 2025 -1762 2040 -1734
rect 2166 -1750 2178 -1734
tri 2166 -1762 2178 -1750 ne
rect 2667 -1710 2699 -1696
rect 2605 -1762 2620 -1734
rect 2746 -1750 2758 -1734
tri 2746 -1762 2758 -1750 ne
rect 3247 -1710 3279 -1696
rect 3185 -1762 3200 -1734
rect 3326 -1750 3338 -1734
tri 3326 -1762 3338 -1750 ne
rect 3827 -1710 3859 -1696
rect 3765 -1762 3780 -1734
rect 3906 -1750 3918 -1734
tri 3906 -1762 3918 -1750 ne
rect 4407 -1710 4439 -1696
rect 4345 -1762 4360 -1734
rect 4486 -1750 4498 -1734
tri 4486 -1762 4498 -1750 ne
rect 4987 -1710 5019 -1696
rect 4925 -1762 4940 -1734
rect 5066 -1750 5078 -1734
tri 5066 -1762 5078 -1750 ne
rect 5567 -1710 5599 -1696
rect 5505 -1762 5520 -1734
rect 5646 -1750 5658 -1734
tri 5646 -1762 5658 -1750 ne
rect 6147 -1710 6179 -1696
rect 6085 -1762 6100 -1734
rect 6226 -1750 6238 -1734
tri 6226 -1762 6238 -1750 ne
rect -233 -1980 -201 -1966
rect -295 -2032 -280 -2004
rect -154 -2020 -142 -2004
tri -154 -2032 -142 -2020 ne
rect 347 -1980 379 -1966
rect 285 -2032 300 -2004
rect 426 -2020 438 -2004
tri 426 -2032 438 -2020 ne
rect 927 -1980 959 -1966
rect 865 -2032 880 -2004
rect 1006 -2020 1018 -2004
tri 1006 -2032 1018 -2020 ne
rect 1507 -1980 1539 -1966
rect 1445 -2032 1460 -2004
rect 1586 -2020 1598 -2004
tri 1586 -2032 1598 -2020 ne
rect 2087 -1980 2119 -1966
rect 2025 -2032 2040 -2004
rect 2166 -2020 2178 -2004
tri 2166 -2032 2178 -2020 ne
rect 2667 -1980 2699 -1966
rect 2605 -2032 2620 -2004
rect 2746 -2020 2758 -2004
tri 2746 -2032 2758 -2020 ne
rect 3247 -1980 3279 -1966
rect 3185 -2032 3200 -2004
rect 3326 -2020 3338 -2004
tri 3326 -2032 3338 -2020 ne
rect 3827 -1980 3859 -1966
rect 3765 -2032 3780 -2004
rect 3906 -2020 3918 -2004
tri 3906 -2032 3918 -2020 ne
rect 4407 -1980 4439 -1966
rect 4345 -2032 4360 -2004
rect 4486 -2020 4498 -2004
tri 4486 -2032 4498 -2020 ne
rect 4987 -1980 5019 -1966
rect 4925 -2032 4940 -2004
rect 5066 -2020 5078 -2004
tri 5066 -2032 5078 -2020 ne
rect 5567 -1980 5599 -1966
rect 5505 -2032 5520 -2004
rect 5646 -2020 5658 -2004
tri 5646 -2032 5658 -2020 ne
rect 6147 -1980 6179 -1966
rect 6085 -2032 6100 -2004
rect 6226 -2020 6238 -2004
tri 6226 -2032 6238 -2020 ne
rect -233 -2250 -201 -2236
rect -295 -2302 -280 -2274
rect -154 -2290 -142 -2274
tri -154 -2302 -142 -2290 ne
rect 347 -2250 379 -2236
rect 285 -2302 300 -2274
rect 426 -2290 438 -2274
tri 426 -2302 438 -2290 ne
rect 927 -2250 959 -2236
rect 865 -2302 880 -2274
rect 1006 -2290 1018 -2274
tri 1006 -2302 1018 -2290 ne
rect 1507 -2250 1539 -2236
rect 1445 -2302 1460 -2274
rect 1586 -2290 1598 -2274
tri 1586 -2302 1598 -2290 ne
rect 2087 -2250 2119 -2236
rect 2025 -2302 2040 -2274
rect 2166 -2290 2178 -2274
tri 2166 -2302 2178 -2290 ne
rect 2667 -2250 2699 -2236
rect 2605 -2302 2620 -2274
rect 2746 -2290 2758 -2274
tri 2746 -2302 2758 -2290 ne
rect 3247 -2250 3279 -2236
rect 3185 -2302 3200 -2274
rect 3326 -2290 3338 -2274
tri 3326 -2302 3338 -2290 ne
rect 3827 -2250 3859 -2236
rect 3765 -2302 3780 -2274
rect 3906 -2290 3918 -2274
tri 3906 -2302 3918 -2290 ne
rect 4407 -2250 4439 -2236
rect 4345 -2302 4360 -2274
rect 4486 -2290 4498 -2274
tri 4486 -2302 4498 -2290 ne
rect 4987 -2250 5019 -2236
rect 4925 -2302 4940 -2274
rect 5066 -2290 5078 -2274
tri 5066 -2302 5078 -2290 ne
rect 5567 -2250 5599 -2236
rect 5505 -2302 5520 -2274
rect 5646 -2290 5658 -2274
tri 5646 -2302 5658 -2290 ne
rect 6147 -2250 6179 -2236
rect 6085 -2302 6100 -2274
rect 6226 -2290 6238 -2274
tri 6226 -2302 6238 -2290 ne
<< psubdiffcont >>
rect -231 1588 -203 1590
rect 349 1588 377 1590
rect 929 1588 957 1590
rect 1509 1588 1537 1590
rect 2089 1588 2117 1590
rect 2669 1588 2697 1590
rect 3249 1588 3277 1590
rect 3829 1588 3857 1590
rect 4409 1588 4437 1590
rect 4989 1588 5017 1590
rect 5569 1588 5597 1590
rect 6149 1588 6177 1590
rect -231 1318 -203 1320
rect 349 1318 377 1320
rect 929 1318 957 1320
rect 1509 1318 1537 1320
rect 2089 1318 2117 1320
rect 2669 1318 2697 1320
rect 3249 1318 3277 1320
rect 3829 1318 3857 1320
rect 4409 1318 4437 1320
rect 4989 1318 5017 1320
rect 5569 1318 5597 1320
rect 6149 1318 6177 1320
rect -231 1048 -203 1050
rect 349 1048 377 1050
rect 929 1048 957 1050
rect 1509 1048 1537 1050
rect 2089 1048 2117 1050
rect 2669 1048 2697 1050
rect 3249 1048 3277 1050
rect 3829 1048 3857 1050
rect 4409 1048 4437 1050
rect 4989 1048 5017 1050
rect 5569 1048 5597 1050
rect 6149 1048 6177 1050
rect -231 778 -203 780
rect 349 778 377 780
rect 929 778 957 780
rect 1509 778 1537 780
rect 2089 778 2117 780
rect 2669 778 2697 780
rect 3249 778 3277 780
rect 3829 778 3857 780
rect 4409 778 4437 780
rect 4989 778 5017 780
rect 5569 778 5597 780
rect 6149 778 6177 780
rect -231 508 -203 510
rect 349 508 377 510
rect 929 508 957 510
rect 1509 508 1537 510
rect 2089 508 2117 510
rect 2669 508 2697 510
rect 3249 508 3277 510
rect 3829 508 3857 510
rect 4409 508 4437 510
rect 4989 508 5017 510
rect 5569 508 5597 510
rect 6149 508 6177 510
rect -231 238 -203 240
rect 349 238 377 240
rect 929 238 957 240
rect 1509 238 1537 240
rect 2089 238 2117 240
rect 2669 238 2697 240
rect 3249 238 3277 240
rect 3829 238 3857 240
rect 4409 238 4437 240
rect 4989 238 5017 240
rect 5569 238 5597 240
rect 6149 238 6177 240
rect -231 -32 -203 -30
rect 349 -32 377 -30
rect 929 -32 957 -30
rect 1509 -32 1537 -30
rect 2089 -32 2117 -30
rect 2669 -32 2697 -30
rect 3249 -32 3277 -30
rect 3829 -32 3857 -30
rect 4409 -32 4437 -30
rect 4989 -32 5017 -30
rect 5569 -32 5597 -30
rect 6149 -32 6177 -30
rect -231 -302 -203 -300
rect 349 -302 377 -300
rect 929 -302 957 -300
rect 1509 -302 1537 -300
rect 2089 -302 2117 -300
rect 2669 -302 2697 -300
rect 3249 -302 3277 -300
rect 3829 -302 3857 -300
rect 4409 -302 4437 -300
rect 4989 -302 5017 -300
rect 5569 -302 5597 -300
rect 6149 -302 6177 -300
rect -231 -572 -203 -570
rect 349 -572 377 -570
rect 929 -572 957 -570
rect 1509 -572 1537 -570
rect 2089 -572 2117 -570
rect 2669 -572 2697 -570
rect 3249 -572 3277 -570
rect 3829 -572 3857 -570
rect 4409 -572 4437 -570
rect 4989 -572 5017 -570
rect 5569 -572 5597 -570
rect 6149 -572 6177 -570
rect -231 -842 -203 -840
rect 349 -842 377 -840
rect 929 -842 957 -840
rect 1509 -842 1537 -840
rect 2089 -842 2117 -840
rect 2669 -842 2697 -840
rect 3249 -842 3277 -840
rect 3829 -842 3857 -840
rect 4409 -842 4437 -840
rect 4989 -842 5017 -840
rect 5569 -842 5597 -840
rect 6149 -842 6177 -840
rect -231 -1112 -203 -1110
rect 349 -1112 377 -1110
rect 929 -1112 957 -1110
rect 1509 -1112 1537 -1110
rect 2089 -1112 2117 -1110
rect 2669 -1112 2697 -1110
rect 3249 -1112 3277 -1110
rect 3829 -1112 3857 -1110
rect 4409 -1112 4437 -1110
rect 4989 -1112 5017 -1110
rect 5569 -1112 5597 -1110
rect 6149 -1112 6177 -1110
rect -231 -1382 -203 -1380
rect 349 -1382 377 -1380
rect 929 -1382 957 -1380
rect 1509 -1382 1537 -1380
rect 2089 -1382 2117 -1380
rect 2669 -1382 2697 -1380
rect 3249 -1382 3277 -1380
rect 3829 -1382 3857 -1380
rect 4409 -1382 4437 -1380
rect 4989 -1382 5017 -1380
rect 5569 -1382 5597 -1380
rect 6149 -1382 6177 -1380
rect -231 -1652 -203 -1650
rect 349 -1652 377 -1650
rect 929 -1652 957 -1650
rect 1509 -1652 1537 -1650
rect 2089 -1652 2117 -1650
rect 2669 -1652 2697 -1650
rect 3249 -1652 3277 -1650
rect 3829 -1652 3857 -1650
rect 4409 -1652 4437 -1650
rect 4989 -1652 5017 -1650
rect 5569 -1652 5597 -1650
rect 6149 -1652 6177 -1650
rect -231 -1922 -203 -1920
rect 349 -1922 377 -1920
rect 929 -1922 957 -1920
rect 1509 -1922 1537 -1920
rect 2089 -1922 2117 -1920
rect 2669 -1922 2697 -1920
rect 3249 -1922 3277 -1920
rect 3829 -1922 3857 -1920
rect 4409 -1922 4437 -1920
rect 4989 -1922 5017 -1920
rect 5569 -1922 5597 -1920
rect 6149 -1922 6177 -1920
rect -231 -2192 -203 -2190
rect 349 -2192 377 -2190
rect 929 -2192 957 -2190
rect 1509 -2192 1537 -2190
rect 2089 -2192 2117 -2190
rect 2669 -2192 2697 -2190
rect 3249 -2192 3277 -2190
rect 3829 -2192 3857 -2190
rect 4409 -2192 4437 -2190
rect 4989 -2192 5017 -2190
rect 5569 -2192 5597 -2190
rect 6149 -2192 6177 -2190
rect -231 -2462 -203 -2460
rect 349 -2462 377 -2460
rect 929 -2462 957 -2460
rect 1509 -2462 1537 -2460
rect 2089 -2462 2117 -2460
rect 2669 -2462 2697 -2460
rect 3249 -2462 3277 -2460
rect 3829 -2462 3857 -2460
rect 4409 -2462 4437 -2460
rect 4989 -2462 5017 -2460
rect 5569 -2462 5597 -2460
rect 6149 -2462 6177 -2460
<< nsubdiffcont >>
rect -231 1798 -203 1800
rect 349 1798 377 1800
rect 929 1798 957 1800
rect 1509 1798 1537 1800
rect 2089 1798 2117 1800
rect 2669 1798 2697 1800
rect 3249 1798 3277 1800
rect 3829 1798 3857 1800
rect 4409 1798 4437 1800
rect 4989 1798 5017 1800
rect 5569 1798 5597 1800
rect 6149 1798 6177 1800
rect -231 1528 -203 1530
rect 349 1528 377 1530
rect 929 1528 957 1530
rect 1509 1528 1537 1530
rect 2089 1528 2117 1530
rect 2669 1528 2697 1530
rect 3249 1528 3277 1530
rect 3829 1528 3857 1530
rect 4409 1528 4437 1530
rect 4989 1528 5017 1530
rect 5569 1528 5597 1530
rect 6149 1528 6177 1530
rect -231 1258 -203 1260
rect 349 1258 377 1260
rect 929 1258 957 1260
rect 1509 1258 1537 1260
rect 2089 1258 2117 1260
rect 2669 1258 2697 1260
rect 3249 1258 3277 1260
rect 3829 1258 3857 1260
rect 4409 1258 4437 1260
rect 4989 1258 5017 1260
rect 5569 1258 5597 1260
rect 6149 1258 6177 1260
rect -231 988 -203 990
rect 349 988 377 990
rect 929 988 957 990
rect 1509 988 1537 990
rect 2089 988 2117 990
rect 2669 988 2697 990
rect 3249 988 3277 990
rect 3829 988 3857 990
rect 4409 988 4437 990
rect 4989 988 5017 990
rect 5569 988 5597 990
rect 6149 988 6177 990
rect -231 718 -203 720
rect 349 718 377 720
rect 929 718 957 720
rect 1509 718 1537 720
rect 2089 718 2117 720
rect 2669 718 2697 720
rect 3249 718 3277 720
rect 3829 718 3857 720
rect 4409 718 4437 720
rect 4989 718 5017 720
rect 5569 718 5597 720
rect 6149 718 6177 720
rect -231 448 -203 450
rect 349 448 377 450
rect 929 448 957 450
rect 1509 448 1537 450
rect 2089 448 2117 450
rect 2669 448 2697 450
rect 3249 448 3277 450
rect 3829 448 3857 450
rect 4409 448 4437 450
rect 4989 448 5017 450
rect 5569 448 5597 450
rect 6149 448 6177 450
rect -231 178 -203 180
rect 349 178 377 180
rect 929 178 957 180
rect 1509 178 1537 180
rect 2089 178 2117 180
rect 2669 178 2697 180
rect 3249 178 3277 180
rect 3829 178 3857 180
rect 4409 178 4437 180
rect 4989 178 5017 180
rect 5569 178 5597 180
rect 6149 178 6177 180
rect -231 -92 -203 -90
rect 349 -92 377 -90
rect 929 -92 957 -90
rect 1509 -92 1537 -90
rect 2089 -92 2117 -90
rect 2669 -92 2697 -90
rect 3249 -92 3277 -90
rect 3829 -92 3857 -90
rect 4409 -92 4437 -90
rect 4989 -92 5017 -90
rect 5569 -92 5597 -90
rect 6149 -92 6177 -90
rect -231 -362 -203 -360
rect 349 -362 377 -360
rect 929 -362 957 -360
rect 1509 -362 1537 -360
rect 2089 -362 2117 -360
rect 2669 -362 2697 -360
rect 3249 -362 3277 -360
rect 3829 -362 3857 -360
rect 4409 -362 4437 -360
rect 4989 -362 5017 -360
rect 5569 -362 5597 -360
rect 6149 -362 6177 -360
rect -231 -632 -203 -630
rect 349 -632 377 -630
rect 929 -632 957 -630
rect 1509 -632 1537 -630
rect 2089 -632 2117 -630
rect 2669 -632 2697 -630
rect 3249 -632 3277 -630
rect 3829 -632 3857 -630
rect 4409 -632 4437 -630
rect 4989 -632 5017 -630
rect 5569 -632 5597 -630
rect 6149 -632 6177 -630
rect -231 -902 -203 -900
rect 349 -902 377 -900
rect 929 -902 957 -900
rect 1509 -902 1537 -900
rect 2089 -902 2117 -900
rect 2669 -902 2697 -900
rect 3249 -902 3277 -900
rect 3829 -902 3857 -900
rect 4409 -902 4437 -900
rect 4989 -902 5017 -900
rect 5569 -902 5597 -900
rect 6149 -902 6177 -900
rect -231 -1172 -203 -1170
rect 349 -1172 377 -1170
rect 929 -1172 957 -1170
rect 1509 -1172 1537 -1170
rect 2089 -1172 2117 -1170
rect 2669 -1172 2697 -1170
rect 3249 -1172 3277 -1170
rect 3829 -1172 3857 -1170
rect 4409 -1172 4437 -1170
rect 4989 -1172 5017 -1170
rect 5569 -1172 5597 -1170
rect 6149 -1172 6177 -1170
rect -231 -1442 -203 -1440
rect 349 -1442 377 -1440
rect 929 -1442 957 -1440
rect 1509 -1442 1537 -1440
rect 2089 -1442 2117 -1440
rect 2669 -1442 2697 -1440
rect 3249 -1442 3277 -1440
rect 3829 -1442 3857 -1440
rect 4409 -1442 4437 -1440
rect 4989 -1442 5017 -1440
rect 5569 -1442 5597 -1440
rect 6149 -1442 6177 -1440
rect -231 -1712 -203 -1710
rect 349 -1712 377 -1710
rect 929 -1712 957 -1710
rect 1509 -1712 1537 -1710
rect 2089 -1712 2117 -1710
rect 2669 -1712 2697 -1710
rect 3249 -1712 3277 -1710
rect 3829 -1712 3857 -1710
rect 4409 -1712 4437 -1710
rect 4989 -1712 5017 -1710
rect 5569 -1712 5597 -1710
rect 6149 -1712 6177 -1710
rect -231 -1982 -203 -1980
rect 349 -1982 377 -1980
rect 929 -1982 957 -1980
rect 1509 -1982 1537 -1980
rect 2089 -1982 2117 -1980
rect 2669 -1982 2697 -1980
rect 3249 -1982 3277 -1980
rect 3829 -1982 3857 -1980
rect 4409 -1982 4437 -1980
rect 4989 -1982 5017 -1980
rect 5569 -1982 5597 -1980
rect 6149 -1982 6177 -1980
rect -231 -2252 -203 -2250
rect 349 -2252 377 -2250
rect 929 -2252 957 -2250
rect 1509 -2252 1537 -2250
rect 2089 -2252 2117 -2250
rect 2669 -2252 2697 -2250
rect 3249 -2252 3277 -2250
rect 3829 -2252 3857 -2250
rect 4409 -2252 4437 -2250
rect 4989 -2252 5017 -2250
rect 5569 -2252 5597 -2250
rect 6149 -2252 6177 -2250
<< poly >>
rect -541 1814 6439 1844
rect -386 1786 -356 1814
rect -271 1776 -241 1798
rect -193 1776 -163 1798
rect -78 1786 -48 1814
rect -386 1736 -356 1758
rect 194 1786 224 1814
rect 309 1776 339 1798
rect 387 1776 417 1798
rect 502 1786 532 1814
rect -271 1715 -241 1748
rect -450 1654 -420 1676
rect -364 1654 -349 1688
rect -271 1654 -241 1681
rect -193 1715 -163 1748
rect -78 1736 -48 1758
rect 194 1736 224 1758
rect 774 1786 804 1814
rect 889 1776 919 1798
rect 967 1776 997 1798
rect 1082 1786 1112 1814
rect 309 1715 339 1748
rect -193 1654 -163 1681
rect -85 1654 -70 1688
rect -14 1654 16 1676
rect 130 1654 160 1676
rect 216 1654 231 1688
rect 309 1654 339 1681
rect 387 1715 417 1748
rect 502 1736 532 1758
rect 774 1736 804 1758
rect 1354 1786 1384 1814
rect 1469 1776 1499 1798
rect 1547 1776 1577 1798
rect 1662 1786 1692 1814
rect 889 1715 919 1748
rect 387 1654 417 1681
rect 495 1654 510 1688
rect 566 1654 596 1676
rect 710 1654 740 1676
rect 796 1654 811 1688
rect 889 1654 919 1681
rect 967 1715 997 1748
rect 1082 1736 1112 1758
rect 1354 1736 1384 1758
rect 1934 1786 1964 1814
rect 2049 1776 2079 1798
rect 2127 1776 2157 1798
rect 2242 1786 2272 1814
rect 1469 1715 1499 1748
rect 967 1654 997 1681
rect 1075 1654 1090 1688
rect 1146 1654 1176 1676
rect 1290 1654 1320 1676
rect 1376 1654 1391 1688
rect 1469 1654 1499 1681
rect 1547 1715 1577 1748
rect 1662 1736 1692 1758
rect 1934 1736 1964 1758
rect 2514 1786 2544 1814
rect 2629 1776 2659 1798
rect 2707 1776 2737 1798
rect 2822 1786 2852 1814
rect 2049 1715 2079 1748
rect 1547 1654 1577 1681
rect 1655 1654 1670 1688
rect 1726 1654 1756 1676
rect 1870 1654 1900 1676
rect 1956 1654 1971 1688
rect 2049 1654 2079 1681
rect 2127 1715 2157 1748
rect 2242 1736 2272 1758
rect 2514 1736 2544 1758
rect 3094 1786 3124 1814
rect 3209 1776 3239 1798
rect 3287 1776 3317 1798
rect 3402 1786 3432 1814
rect 2629 1715 2659 1748
rect 2127 1654 2157 1681
rect 2235 1654 2250 1688
rect 2306 1654 2336 1676
rect 2450 1654 2480 1676
rect 2536 1654 2551 1688
rect 2629 1654 2659 1681
rect 2707 1715 2737 1748
rect 2822 1736 2852 1758
rect 3094 1736 3124 1758
rect 3674 1786 3704 1814
rect 3789 1776 3819 1798
rect 3867 1776 3897 1798
rect 3982 1786 4012 1814
rect 3209 1715 3239 1748
rect 2707 1654 2737 1681
rect 2815 1654 2830 1688
rect 2886 1654 2916 1676
rect 3030 1654 3060 1676
rect 3116 1654 3131 1688
rect 3209 1654 3239 1681
rect 3287 1715 3317 1748
rect 3402 1736 3432 1758
rect 3674 1736 3704 1758
rect 4254 1786 4284 1814
rect 4369 1776 4399 1798
rect 4447 1776 4477 1798
rect 4562 1786 4592 1814
rect 3789 1715 3819 1748
rect 3287 1654 3317 1681
rect 3395 1654 3410 1688
rect 3466 1654 3496 1676
rect 3610 1654 3640 1676
rect 3696 1654 3711 1688
rect 3789 1654 3819 1681
rect 3867 1715 3897 1748
rect 3982 1736 4012 1758
rect 4254 1736 4284 1758
rect 4834 1786 4864 1814
rect 4949 1776 4979 1798
rect 5027 1776 5057 1798
rect 5142 1786 5172 1814
rect 4369 1715 4399 1748
rect 3867 1654 3897 1681
rect 3975 1654 3990 1688
rect 4046 1654 4076 1676
rect 4190 1654 4220 1676
rect 4276 1654 4291 1688
rect 4369 1654 4399 1681
rect 4447 1715 4477 1748
rect 4562 1736 4592 1758
rect 4834 1736 4864 1758
rect 5414 1786 5444 1814
rect 5529 1776 5559 1798
rect 5607 1776 5637 1798
rect 5722 1786 5752 1814
rect 4949 1715 4979 1748
rect 4447 1654 4477 1681
rect 4555 1654 4570 1688
rect 4626 1654 4656 1676
rect 4770 1654 4800 1676
rect 4856 1654 4871 1688
rect 4949 1654 4979 1681
rect 5027 1715 5057 1748
rect 5142 1736 5172 1758
rect 5414 1736 5444 1758
rect 5994 1786 6024 1814
rect 6109 1776 6139 1798
rect 6187 1776 6217 1798
rect 6302 1786 6332 1814
rect 5529 1715 5559 1748
rect 5027 1654 5057 1681
rect 5135 1654 5150 1688
rect 5206 1654 5236 1676
rect 5350 1654 5380 1676
rect 5436 1654 5451 1688
rect 5529 1654 5559 1681
rect 5607 1715 5637 1748
rect 5722 1736 5752 1758
rect 5994 1736 6024 1758
rect 6109 1715 6139 1748
rect 5607 1654 5637 1681
rect 5715 1654 5730 1688
rect 5786 1654 5816 1676
rect 5930 1654 5960 1676
rect 6016 1654 6031 1688
rect 6109 1654 6139 1681
rect 6187 1715 6217 1748
rect 6302 1736 6332 1758
rect 6187 1654 6217 1681
rect 6295 1654 6310 1688
rect 6366 1654 6396 1676
rect -364 1640 -334 1654
rect -100 1640 -70 1654
rect 216 1640 246 1654
rect 480 1640 510 1654
rect 796 1640 826 1654
rect 1060 1640 1090 1654
rect 1376 1640 1406 1654
rect 1640 1640 1670 1654
rect 1956 1640 1986 1654
rect 2220 1640 2250 1654
rect 2536 1640 2566 1654
rect 2800 1640 2830 1654
rect 3116 1640 3146 1654
rect 3380 1640 3410 1654
rect 3696 1640 3726 1654
rect 3960 1640 3990 1654
rect 4276 1640 4306 1654
rect 4540 1640 4570 1654
rect 4856 1640 4886 1654
rect 5120 1640 5150 1654
rect 5436 1640 5466 1654
rect 5700 1640 5730 1654
rect 6016 1640 6046 1654
rect 6280 1640 6310 1654
rect -450 1590 -420 1612
rect -364 1590 -334 1612
rect -271 1590 -241 1612
rect -193 1590 -163 1612
rect -100 1590 -70 1612
rect -14 1590 16 1612
rect 130 1590 160 1612
rect 216 1590 246 1612
rect 309 1590 339 1612
rect 387 1590 417 1612
rect 480 1590 510 1612
rect 566 1590 596 1612
rect 710 1590 740 1612
rect 796 1590 826 1612
rect 889 1590 919 1612
rect 967 1590 997 1612
rect 1060 1590 1090 1612
rect 1146 1590 1176 1612
rect 1290 1590 1320 1612
rect 1376 1590 1406 1612
rect 1469 1590 1499 1612
rect 1547 1590 1577 1612
rect 1640 1590 1670 1612
rect 1726 1590 1756 1612
rect 1870 1590 1900 1612
rect 1956 1590 1986 1612
rect 2049 1590 2079 1612
rect 2127 1590 2157 1612
rect 2220 1590 2250 1612
rect 2306 1590 2336 1612
rect 2450 1590 2480 1612
rect 2536 1590 2566 1612
rect 2629 1590 2659 1612
rect 2707 1590 2737 1612
rect 2800 1590 2830 1612
rect 2886 1590 2916 1612
rect 3030 1590 3060 1612
rect 3116 1590 3146 1612
rect 3209 1590 3239 1612
rect 3287 1590 3317 1612
rect 3380 1590 3410 1612
rect 3466 1590 3496 1612
rect 3610 1590 3640 1612
rect 3696 1590 3726 1612
rect 3789 1590 3819 1612
rect 3867 1590 3897 1612
rect 3960 1590 3990 1612
rect 4046 1590 4076 1612
rect 4190 1590 4220 1612
rect 4276 1590 4306 1612
rect 4369 1590 4399 1612
rect 4447 1590 4477 1612
rect 4540 1590 4570 1612
rect 4626 1590 4656 1612
rect 4770 1590 4800 1612
rect 4856 1590 4886 1612
rect 4949 1590 4979 1612
rect 5027 1590 5057 1612
rect 5120 1590 5150 1612
rect 5206 1590 5236 1612
rect 5350 1590 5380 1612
rect 5436 1590 5466 1612
rect 5529 1590 5559 1612
rect 5607 1590 5637 1612
rect 5700 1590 5730 1612
rect 5786 1590 5816 1612
rect 5930 1590 5960 1612
rect 6016 1590 6046 1612
rect 6109 1590 6139 1612
rect 6187 1590 6217 1612
rect 6280 1590 6310 1612
rect 6366 1590 6396 1612
rect -541 1544 6439 1574
rect -386 1516 -356 1544
rect -271 1506 -241 1528
rect -193 1506 -163 1528
rect -78 1516 -48 1544
rect -386 1466 -356 1488
rect 194 1516 224 1544
rect 309 1506 339 1528
rect 387 1506 417 1528
rect 502 1516 532 1544
rect -271 1445 -241 1478
rect -450 1384 -420 1406
rect -364 1384 -349 1418
rect -271 1384 -241 1411
rect -193 1445 -163 1478
rect -78 1466 -48 1488
rect 194 1466 224 1488
rect 774 1516 804 1544
rect 889 1506 919 1528
rect 967 1506 997 1528
rect 1082 1516 1112 1544
rect 309 1445 339 1478
rect -193 1384 -163 1411
rect -85 1384 -70 1418
rect -14 1384 16 1406
rect 130 1384 160 1406
rect 216 1384 231 1418
rect 309 1384 339 1411
rect 387 1445 417 1478
rect 502 1466 532 1488
rect 774 1466 804 1488
rect 1354 1516 1384 1544
rect 1469 1506 1499 1528
rect 1547 1506 1577 1528
rect 1662 1516 1692 1544
rect 889 1445 919 1478
rect 387 1384 417 1411
rect 495 1384 510 1418
rect 566 1384 596 1406
rect 710 1384 740 1406
rect 796 1384 811 1418
rect 889 1384 919 1411
rect 967 1445 997 1478
rect 1082 1466 1112 1488
rect 1354 1466 1384 1488
rect 1934 1516 1964 1544
rect 2049 1506 2079 1528
rect 2127 1506 2157 1528
rect 2242 1516 2272 1544
rect 1469 1445 1499 1478
rect 967 1384 997 1411
rect 1075 1384 1090 1418
rect 1146 1384 1176 1406
rect 1290 1384 1320 1406
rect 1376 1384 1391 1418
rect 1469 1384 1499 1411
rect 1547 1445 1577 1478
rect 1662 1466 1692 1488
rect 1934 1466 1964 1488
rect 2514 1516 2544 1544
rect 2629 1506 2659 1528
rect 2707 1506 2737 1528
rect 2822 1516 2852 1544
rect 2049 1445 2079 1478
rect 1547 1384 1577 1411
rect 1655 1384 1670 1418
rect 1726 1384 1756 1406
rect 1870 1384 1900 1406
rect 1956 1384 1971 1418
rect 2049 1384 2079 1411
rect 2127 1445 2157 1478
rect 2242 1466 2272 1488
rect 2514 1466 2544 1488
rect 3094 1516 3124 1544
rect 3209 1506 3239 1528
rect 3287 1506 3317 1528
rect 3402 1516 3432 1544
rect 2629 1445 2659 1478
rect 2127 1384 2157 1411
rect 2235 1384 2250 1418
rect 2306 1384 2336 1406
rect 2450 1384 2480 1406
rect 2536 1384 2551 1418
rect 2629 1384 2659 1411
rect 2707 1445 2737 1478
rect 2822 1466 2852 1488
rect 3094 1466 3124 1488
rect 3674 1516 3704 1544
rect 3789 1506 3819 1528
rect 3867 1506 3897 1528
rect 3982 1516 4012 1544
rect 3209 1445 3239 1478
rect 2707 1384 2737 1411
rect 2815 1384 2830 1418
rect 2886 1384 2916 1406
rect 3030 1384 3060 1406
rect 3116 1384 3131 1418
rect 3209 1384 3239 1411
rect 3287 1445 3317 1478
rect 3402 1466 3432 1488
rect 3674 1466 3704 1488
rect 4254 1516 4284 1544
rect 4369 1506 4399 1528
rect 4447 1506 4477 1528
rect 4562 1516 4592 1544
rect 3789 1445 3819 1478
rect 3287 1384 3317 1411
rect 3395 1384 3410 1418
rect 3466 1384 3496 1406
rect 3610 1384 3640 1406
rect 3696 1384 3711 1418
rect 3789 1384 3819 1411
rect 3867 1445 3897 1478
rect 3982 1466 4012 1488
rect 4254 1466 4284 1488
rect 4834 1516 4864 1544
rect 4949 1506 4979 1528
rect 5027 1506 5057 1528
rect 5142 1516 5172 1544
rect 4369 1445 4399 1478
rect 3867 1384 3897 1411
rect 3975 1384 3990 1418
rect 4046 1384 4076 1406
rect 4190 1384 4220 1406
rect 4276 1384 4291 1418
rect 4369 1384 4399 1411
rect 4447 1445 4477 1478
rect 4562 1466 4592 1488
rect 4834 1466 4864 1488
rect 5414 1516 5444 1544
rect 5529 1506 5559 1528
rect 5607 1506 5637 1528
rect 5722 1516 5752 1544
rect 4949 1445 4979 1478
rect 4447 1384 4477 1411
rect 4555 1384 4570 1418
rect 4626 1384 4656 1406
rect 4770 1384 4800 1406
rect 4856 1384 4871 1418
rect 4949 1384 4979 1411
rect 5027 1445 5057 1478
rect 5142 1466 5172 1488
rect 5414 1466 5444 1488
rect 5994 1516 6024 1544
rect 6109 1506 6139 1528
rect 6187 1506 6217 1528
rect 6302 1516 6332 1544
rect 5529 1445 5559 1478
rect 5027 1384 5057 1411
rect 5135 1384 5150 1418
rect 5206 1384 5236 1406
rect 5350 1384 5380 1406
rect 5436 1384 5451 1418
rect 5529 1384 5559 1411
rect 5607 1445 5637 1478
rect 5722 1466 5752 1488
rect 5994 1466 6024 1488
rect 6109 1445 6139 1478
rect 5607 1384 5637 1411
rect 5715 1384 5730 1418
rect 5786 1384 5816 1406
rect 5930 1384 5960 1406
rect 6016 1384 6031 1418
rect 6109 1384 6139 1411
rect 6187 1445 6217 1478
rect 6302 1466 6332 1488
rect 6187 1384 6217 1411
rect 6295 1384 6310 1418
rect 6366 1384 6396 1406
rect -364 1370 -334 1384
rect -100 1370 -70 1384
rect 216 1370 246 1384
rect 480 1370 510 1384
rect 796 1370 826 1384
rect 1060 1370 1090 1384
rect 1376 1370 1406 1384
rect 1640 1370 1670 1384
rect 1956 1370 1986 1384
rect 2220 1370 2250 1384
rect 2536 1370 2566 1384
rect 2800 1370 2830 1384
rect 3116 1370 3146 1384
rect 3380 1370 3410 1384
rect 3696 1370 3726 1384
rect 3960 1370 3990 1384
rect 4276 1370 4306 1384
rect 4540 1370 4570 1384
rect 4856 1370 4886 1384
rect 5120 1370 5150 1384
rect 5436 1370 5466 1384
rect 5700 1370 5730 1384
rect 6016 1370 6046 1384
rect 6280 1370 6310 1384
rect -450 1320 -420 1342
rect -364 1320 -334 1342
rect -271 1320 -241 1342
rect -193 1320 -163 1342
rect -100 1320 -70 1342
rect -14 1320 16 1342
rect 130 1320 160 1342
rect 216 1320 246 1342
rect 309 1320 339 1342
rect 387 1320 417 1342
rect 480 1320 510 1342
rect 566 1320 596 1342
rect 710 1320 740 1342
rect 796 1320 826 1342
rect 889 1320 919 1342
rect 967 1320 997 1342
rect 1060 1320 1090 1342
rect 1146 1320 1176 1342
rect 1290 1320 1320 1342
rect 1376 1320 1406 1342
rect 1469 1320 1499 1342
rect 1547 1320 1577 1342
rect 1640 1320 1670 1342
rect 1726 1320 1756 1342
rect 1870 1320 1900 1342
rect 1956 1320 1986 1342
rect 2049 1320 2079 1342
rect 2127 1320 2157 1342
rect 2220 1320 2250 1342
rect 2306 1320 2336 1342
rect 2450 1320 2480 1342
rect 2536 1320 2566 1342
rect 2629 1320 2659 1342
rect 2707 1320 2737 1342
rect 2800 1320 2830 1342
rect 2886 1320 2916 1342
rect 3030 1320 3060 1342
rect 3116 1320 3146 1342
rect 3209 1320 3239 1342
rect 3287 1320 3317 1342
rect 3380 1320 3410 1342
rect 3466 1320 3496 1342
rect 3610 1320 3640 1342
rect 3696 1320 3726 1342
rect 3789 1320 3819 1342
rect 3867 1320 3897 1342
rect 3960 1320 3990 1342
rect 4046 1320 4076 1342
rect 4190 1320 4220 1342
rect 4276 1320 4306 1342
rect 4369 1320 4399 1342
rect 4447 1320 4477 1342
rect 4540 1320 4570 1342
rect 4626 1320 4656 1342
rect 4770 1320 4800 1342
rect 4856 1320 4886 1342
rect 4949 1320 4979 1342
rect 5027 1320 5057 1342
rect 5120 1320 5150 1342
rect 5206 1320 5236 1342
rect 5350 1320 5380 1342
rect 5436 1320 5466 1342
rect 5529 1320 5559 1342
rect 5607 1320 5637 1342
rect 5700 1320 5730 1342
rect 5786 1320 5816 1342
rect 5930 1320 5960 1342
rect 6016 1320 6046 1342
rect 6109 1320 6139 1342
rect 6187 1320 6217 1342
rect 6280 1320 6310 1342
rect 6366 1320 6396 1342
rect -541 1274 6439 1304
rect -386 1246 -356 1274
rect -271 1236 -241 1258
rect -193 1236 -163 1258
rect -78 1246 -48 1274
rect -386 1196 -356 1218
rect 194 1246 224 1274
rect 309 1236 339 1258
rect 387 1236 417 1258
rect 502 1246 532 1274
rect -271 1175 -241 1208
rect -450 1114 -420 1136
rect -364 1114 -349 1148
rect -271 1114 -241 1141
rect -193 1175 -163 1208
rect -78 1196 -48 1218
rect 194 1196 224 1218
rect 774 1246 804 1274
rect 889 1236 919 1258
rect 967 1236 997 1258
rect 1082 1246 1112 1274
rect 309 1175 339 1208
rect -193 1114 -163 1141
rect -85 1114 -70 1148
rect -14 1114 16 1136
rect 130 1114 160 1136
rect 216 1114 231 1148
rect 309 1114 339 1141
rect 387 1175 417 1208
rect 502 1196 532 1218
rect 774 1196 804 1218
rect 1354 1246 1384 1274
rect 1469 1236 1499 1258
rect 1547 1236 1577 1258
rect 1662 1246 1692 1274
rect 889 1175 919 1208
rect 387 1114 417 1141
rect 495 1114 510 1148
rect 566 1114 596 1136
rect 710 1114 740 1136
rect 796 1114 811 1148
rect 889 1114 919 1141
rect 967 1175 997 1208
rect 1082 1196 1112 1218
rect 1354 1196 1384 1218
rect 1934 1246 1964 1274
rect 2049 1236 2079 1258
rect 2127 1236 2157 1258
rect 2242 1246 2272 1274
rect 1469 1175 1499 1208
rect 967 1114 997 1141
rect 1075 1114 1090 1148
rect 1146 1114 1176 1136
rect 1290 1114 1320 1136
rect 1376 1114 1391 1148
rect 1469 1114 1499 1141
rect 1547 1175 1577 1208
rect 1662 1196 1692 1218
rect 1934 1196 1964 1218
rect 2514 1246 2544 1274
rect 2629 1236 2659 1258
rect 2707 1236 2737 1258
rect 2822 1246 2852 1274
rect 2049 1175 2079 1208
rect 1547 1114 1577 1141
rect 1655 1114 1670 1148
rect 1726 1114 1756 1136
rect 1870 1114 1900 1136
rect 1956 1114 1971 1148
rect 2049 1114 2079 1141
rect 2127 1175 2157 1208
rect 2242 1196 2272 1218
rect 2514 1196 2544 1218
rect 3094 1246 3124 1274
rect 3209 1236 3239 1258
rect 3287 1236 3317 1258
rect 3402 1246 3432 1274
rect 2629 1175 2659 1208
rect 2127 1114 2157 1141
rect 2235 1114 2250 1148
rect 2306 1114 2336 1136
rect 2450 1114 2480 1136
rect 2536 1114 2551 1148
rect 2629 1114 2659 1141
rect 2707 1175 2737 1208
rect 2822 1196 2852 1218
rect 3094 1196 3124 1218
rect 3674 1246 3704 1274
rect 3789 1236 3819 1258
rect 3867 1236 3897 1258
rect 3982 1246 4012 1274
rect 3209 1175 3239 1208
rect 2707 1114 2737 1141
rect 2815 1114 2830 1148
rect 2886 1114 2916 1136
rect 3030 1114 3060 1136
rect 3116 1114 3131 1148
rect 3209 1114 3239 1141
rect 3287 1175 3317 1208
rect 3402 1196 3432 1218
rect 3674 1196 3704 1218
rect 4254 1246 4284 1274
rect 4369 1236 4399 1258
rect 4447 1236 4477 1258
rect 4562 1246 4592 1274
rect 3789 1175 3819 1208
rect 3287 1114 3317 1141
rect 3395 1114 3410 1148
rect 3466 1114 3496 1136
rect 3610 1114 3640 1136
rect 3696 1114 3711 1148
rect 3789 1114 3819 1141
rect 3867 1175 3897 1208
rect 3982 1196 4012 1218
rect 4254 1196 4284 1218
rect 4834 1246 4864 1274
rect 4949 1236 4979 1258
rect 5027 1236 5057 1258
rect 5142 1246 5172 1274
rect 4369 1175 4399 1208
rect 3867 1114 3897 1141
rect 3975 1114 3990 1148
rect 4046 1114 4076 1136
rect 4190 1114 4220 1136
rect 4276 1114 4291 1148
rect 4369 1114 4399 1141
rect 4447 1175 4477 1208
rect 4562 1196 4592 1218
rect 4834 1196 4864 1218
rect 5414 1246 5444 1274
rect 5529 1236 5559 1258
rect 5607 1236 5637 1258
rect 5722 1246 5752 1274
rect 4949 1175 4979 1208
rect 4447 1114 4477 1141
rect 4555 1114 4570 1148
rect 4626 1114 4656 1136
rect 4770 1114 4800 1136
rect 4856 1114 4871 1148
rect 4949 1114 4979 1141
rect 5027 1175 5057 1208
rect 5142 1196 5172 1218
rect 5414 1196 5444 1218
rect 5994 1246 6024 1274
rect 6109 1236 6139 1258
rect 6187 1236 6217 1258
rect 6302 1246 6332 1274
rect 5529 1175 5559 1208
rect 5027 1114 5057 1141
rect 5135 1114 5150 1148
rect 5206 1114 5236 1136
rect 5350 1114 5380 1136
rect 5436 1114 5451 1148
rect 5529 1114 5559 1141
rect 5607 1175 5637 1208
rect 5722 1196 5752 1218
rect 5994 1196 6024 1218
rect 6109 1175 6139 1208
rect 5607 1114 5637 1141
rect 5715 1114 5730 1148
rect 5786 1114 5816 1136
rect 5930 1114 5960 1136
rect 6016 1114 6031 1148
rect 6109 1114 6139 1141
rect 6187 1175 6217 1208
rect 6302 1196 6332 1218
rect 6187 1114 6217 1141
rect 6295 1114 6310 1148
rect 6366 1114 6396 1136
rect -364 1100 -334 1114
rect -100 1100 -70 1114
rect 216 1100 246 1114
rect 480 1100 510 1114
rect 796 1100 826 1114
rect 1060 1100 1090 1114
rect 1376 1100 1406 1114
rect 1640 1100 1670 1114
rect 1956 1100 1986 1114
rect 2220 1100 2250 1114
rect 2536 1100 2566 1114
rect 2800 1100 2830 1114
rect 3116 1100 3146 1114
rect 3380 1100 3410 1114
rect 3696 1100 3726 1114
rect 3960 1100 3990 1114
rect 4276 1100 4306 1114
rect 4540 1100 4570 1114
rect 4856 1100 4886 1114
rect 5120 1100 5150 1114
rect 5436 1100 5466 1114
rect 5700 1100 5730 1114
rect 6016 1100 6046 1114
rect 6280 1100 6310 1114
rect -450 1050 -420 1072
rect -364 1050 -334 1072
rect -271 1050 -241 1072
rect -193 1050 -163 1072
rect -100 1050 -70 1072
rect -14 1050 16 1072
rect 130 1050 160 1072
rect 216 1050 246 1072
rect 309 1050 339 1072
rect 387 1050 417 1072
rect 480 1050 510 1072
rect 566 1050 596 1072
rect 710 1050 740 1072
rect 796 1050 826 1072
rect 889 1050 919 1072
rect 967 1050 997 1072
rect 1060 1050 1090 1072
rect 1146 1050 1176 1072
rect 1290 1050 1320 1072
rect 1376 1050 1406 1072
rect 1469 1050 1499 1072
rect 1547 1050 1577 1072
rect 1640 1050 1670 1072
rect 1726 1050 1756 1072
rect 1870 1050 1900 1072
rect 1956 1050 1986 1072
rect 2049 1050 2079 1072
rect 2127 1050 2157 1072
rect 2220 1050 2250 1072
rect 2306 1050 2336 1072
rect 2450 1050 2480 1072
rect 2536 1050 2566 1072
rect 2629 1050 2659 1072
rect 2707 1050 2737 1072
rect 2800 1050 2830 1072
rect 2886 1050 2916 1072
rect 3030 1050 3060 1072
rect 3116 1050 3146 1072
rect 3209 1050 3239 1072
rect 3287 1050 3317 1072
rect 3380 1050 3410 1072
rect 3466 1050 3496 1072
rect 3610 1050 3640 1072
rect 3696 1050 3726 1072
rect 3789 1050 3819 1072
rect 3867 1050 3897 1072
rect 3960 1050 3990 1072
rect 4046 1050 4076 1072
rect 4190 1050 4220 1072
rect 4276 1050 4306 1072
rect 4369 1050 4399 1072
rect 4447 1050 4477 1072
rect 4540 1050 4570 1072
rect 4626 1050 4656 1072
rect 4770 1050 4800 1072
rect 4856 1050 4886 1072
rect 4949 1050 4979 1072
rect 5027 1050 5057 1072
rect 5120 1050 5150 1072
rect 5206 1050 5236 1072
rect 5350 1050 5380 1072
rect 5436 1050 5466 1072
rect 5529 1050 5559 1072
rect 5607 1050 5637 1072
rect 5700 1050 5730 1072
rect 5786 1050 5816 1072
rect 5930 1050 5960 1072
rect 6016 1050 6046 1072
rect 6109 1050 6139 1072
rect 6187 1050 6217 1072
rect 6280 1050 6310 1072
rect 6366 1050 6396 1072
rect -541 1004 6439 1034
rect -386 976 -356 1004
rect -271 966 -241 988
rect -193 966 -163 988
rect -78 976 -48 1004
rect -386 926 -356 948
rect 194 976 224 1004
rect 309 966 339 988
rect 387 966 417 988
rect 502 976 532 1004
rect -271 905 -241 938
rect -450 844 -420 866
rect -364 844 -349 878
rect -271 844 -241 871
rect -193 905 -163 938
rect -78 926 -48 948
rect 194 926 224 948
rect 774 976 804 1004
rect 889 966 919 988
rect 967 966 997 988
rect 1082 976 1112 1004
rect 309 905 339 938
rect -193 844 -163 871
rect -85 844 -70 878
rect -14 844 16 866
rect 130 844 160 866
rect 216 844 231 878
rect 309 844 339 871
rect 387 905 417 938
rect 502 926 532 948
rect 774 926 804 948
rect 1354 976 1384 1004
rect 1469 966 1499 988
rect 1547 966 1577 988
rect 1662 976 1692 1004
rect 889 905 919 938
rect 387 844 417 871
rect 495 844 510 878
rect 566 844 596 866
rect 710 844 740 866
rect 796 844 811 878
rect 889 844 919 871
rect 967 905 997 938
rect 1082 926 1112 948
rect 1354 926 1384 948
rect 1934 976 1964 1004
rect 2049 966 2079 988
rect 2127 966 2157 988
rect 2242 976 2272 1004
rect 1469 905 1499 938
rect 967 844 997 871
rect 1075 844 1090 878
rect 1146 844 1176 866
rect 1290 844 1320 866
rect 1376 844 1391 878
rect 1469 844 1499 871
rect 1547 905 1577 938
rect 1662 926 1692 948
rect 1934 926 1964 948
rect 2514 976 2544 1004
rect 2629 966 2659 988
rect 2707 966 2737 988
rect 2822 976 2852 1004
rect 2049 905 2079 938
rect 1547 844 1577 871
rect 1655 844 1670 878
rect 1726 844 1756 866
rect 1870 844 1900 866
rect 1956 844 1971 878
rect 2049 844 2079 871
rect 2127 905 2157 938
rect 2242 926 2272 948
rect 2514 926 2544 948
rect 3094 976 3124 1004
rect 3209 966 3239 988
rect 3287 966 3317 988
rect 3402 976 3432 1004
rect 2629 905 2659 938
rect 2127 844 2157 871
rect 2235 844 2250 878
rect 2306 844 2336 866
rect 2450 844 2480 866
rect 2536 844 2551 878
rect 2629 844 2659 871
rect 2707 905 2737 938
rect 2822 926 2852 948
rect 3094 926 3124 948
rect 3674 976 3704 1004
rect 3789 966 3819 988
rect 3867 966 3897 988
rect 3982 976 4012 1004
rect 3209 905 3239 938
rect 2707 844 2737 871
rect 2815 844 2830 878
rect 2886 844 2916 866
rect 3030 844 3060 866
rect 3116 844 3131 878
rect 3209 844 3239 871
rect 3287 905 3317 938
rect 3402 926 3432 948
rect 3674 926 3704 948
rect 4254 976 4284 1004
rect 4369 966 4399 988
rect 4447 966 4477 988
rect 4562 976 4592 1004
rect 3789 905 3819 938
rect 3287 844 3317 871
rect 3395 844 3410 878
rect 3466 844 3496 866
rect 3610 844 3640 866
rect 3696 844 3711 878
rect 3789 844 3819 871
rect 3867 905 3897 938
rect 3982 926 4012 948
rect 4254 926 4284 948
rect 4834 976 4864 1004
rect 4949 966 4979 988
rect 5027 966 5057 988
rect 5142 976 5172 1004
rect 4369 905 4399 938
rect 3867 844 3897 871
rect 3975 844 3990 878
rect 4046 844 4076 866
rect 4190 844 4220 866
rect 4276 844 4291 878
rect 4369 844 4399 871
rect 4447 905 4477 938
rect 4562 926 4592 948
rect 4834 926 4864 948
rect 5414 976 5444 1004
rect 5529 966 5559 988
rect 5607 966 5637 988
rect 5722 976 5752 1004
rect 4949 905 4979 938
rect 4447 844 4477 871
rect 4555 844 4570 878
rect 4626 844 4656 866
rect 4770 844 4800 866
rect 4856 844 4871 878
rect 4949 844 4979 871
rect 5027 905 5057 938
rect 5142 926 5172 948
rect 5414 926 5444 948
rect 5994 976 6024 1004
rect 6109 966 6139 988
rect 6187 966 6217 988
rect 6302 976 6332 1004
rect 5529 905 5559 938
rect 5027 844 5057 871
rect 5135 844 5150 878
rect 5206 844 5236 866
rect 5350 844 5380 866
rect 5436 844 5451 878
rect 5529 844 5559 871
rect 5607 905 5637 938
rect 5722 926 5752 948
rect 5994 926 6024 948
rect 6109 905 6139 938
rect 5607 844 5637 871
rect 5715 844 5730 878
rect 5786 844 5816 866
rect 5930 844 5960 866
rect 6016 844 6031 878
rect 6109 844 6139 871
rect 6187 905 6217 938
rect 6302 926 6332 948
rect 6187 844 6217 871
rect 6295 844 6310 878
rect 6366 844 6396 866
rect -364 830 -334 844
rect -100 830 -70 844
rect 216 830 246 844
rect 480 830 510 844
rect 796 830 826 844
rect 1060 830 1090 844
rect 1376 830 1406 844
rect 1640 830 1670 844
rect 1956 830 1986 844
rect 2220 830 2250 844
rect 2536 830 2566 844
rect 2800 830 2830 844
rect 3116 830 3146 844
rect 3380 830 3410 844
rect 3696 830 3726 844
rect 3960 830 3990 844
rect 4276 830 4306 844
rect 4540 830 4570 844
rect 4856 830 4886 844
rect 5120 830 5150 844
rect 5436 830 5466 844
rect 5700 830 5730 844
rect 6016 830 6046 844
rect 6280 830 6310 844
rect -450 780 -420 802
rect -364 780 -334 802
rect -271 780 -241 802
rect -193 780 -163 802
rect -100 780 -70 802
rect -14 780 16 802
rect 130 780 160 802
rect 216 780 246 802
rect 309 780 339 802
rect 387 780 417 802
rect 480 780 510 802
rect 566 780 596 802
rect 710 780 740 802
rect 796 780 826 802
rect 889 780 919 802
rect 967 780 997 802
rect 1060 780 1090 802
rect 1146 780 1176 802
rect 1290 780 1320 802
rect 1376 780 1406 802
rect 1469 780 1499 802
rect 1547 780 1577 802
rect 1640 780 1670 802
rect 1726 780 1756 802
rect 1870 780 1900 802
rect 1956 780 1986 802
rect 2049 780 2079 802
rect 2127 780 2157 802
rect 2220 780 2250 802
rect 2306 780 2336 802
rect 2450 780 2480 802
rect 2536 780 2566 802
rect 2629 780 2659 802
rect 2707 780 2737 802
rect 2800 780 2830 802
rect 2886 780 2916 802
rect 3030 780 3060 802
rect 3116 780 3146 802
rect 3209 780 3239 802
rect 3287 780 3317 802
rect 3380 780 3410 802
rect 3466 780 3496 802
rect 3610 780 3640 802
rect 3696 780 3726 802
rect 3789 780 3819 802
rect 3867 780 3897 802
rect 3960 780 3990 802
rect 4046 780 4076 802
rect 4190 780 4220 802
rect 4276 780 4306 802
rect 4369 780 4399 802
rect 4447 780 4477 802
rect 4540 780 4570 802
rect 4626 780 4656 802
rect 4770 780 4800 802
rect 4856 780 4886 802
rect 4949 780 4979 802
rect 5027 780 5057 802
rect 5120 780 5150 802
rect 5206 780 5236 802
rect 5350 780 5380 802
rect 5436 780 5466 802
rect 5529 780 5559 802
rect 5607 780 5637 802
rect 5700 780 5730 802
rect 5786 780 5816 802
rect 5930 780 5960 802
rect 6016 780 6046 802
rect 6109 780 6139 802
rect 6187 780 6217 802
rect 6280 780 6310 802
rect 6366 780 6396 802
rect -541 734 6439 764
rect -386 706 -356 734
rect -271 696 -241 718
rect -193 696 -163 718
rect -78 706 -48 734
rect -386 656 -356 678
rect 194 706 224 734
rect 309 696 339 718
rect 387 696 417 718
rect 502 706 532 734
rect -271 635 -241 668
rect -450 574 -420 596
rect -364 574 -349 608
rect -271 574 -241 601
rect -193 635 -163 668
rect -78 656 -48 678
rect 194 656 224 678
rect 774 706 804 734
rect 889 696 919 718
rect 967 696 997 718
rect 1082 706 1112 734
rect 309 635 339 668
rect -193 574 -163 601
rect -85 574 -70 608
rect -14 574 16 596
rect 130 574 160 596
rect 216 574 231 608
rect 309 574 339 601
rect 387 635 417 668
rect 502 656 532 678
rect 774 656 804 678
rect 1354 706 1384 734
rect 1469 696 1499 718
rect 1547 696 1577 718
rect 1662 706 1692 734
rect 889 635 919 668
rect 387 574 417 601
rect 495 574 510 608
rect 566 574 596 596
rect 710 574 740 596
rect 796 574 811 608
rect 889 574 919 601
rect 967 635 997 668
rect 1082 656 1112 678
rect 1354 656 1384 678
rect 1934 706 1964 734
rect 2049 696 2079 718
rect 2127 696 2157 718
rect 2242 706 2272 734
rect 1469 635 1499 668
rect 967 574 997 601
rect 1075 574 1090 608
rect 1146 574 1176 596
rect 1290 574 1320 596
rect 1376 574 1391 608
rect 1469 574 1499 601
rect 1547 635 1577 668
rect 1662 656 1692 678
rect 1934 656 1964 678
rect 2514 706 2544 734
rect 2629 696 2659 718
rect 2707 696 2737 718
rect 2822 706 2852 734
rect 2049 635 2079 668
rect 1547 574 1577 601
rect 1655 574 1670 608
rect 1726 574 1756 596
rect 1870 574 1900 596
rect 1956 574 1971 608
rect 2049 574 2079 601
rect 2127 635 2157 668
rect 2242 656 2272 678
rect 2514 656 2544 678
rect 3094 706 3124 734
rect 3209 696 3239 718
rect 3287 696 3317 718
rect 3402 706 3432 734
rect 2629 635 2659 668
rect 2127 574 2157 601
rect 2235 574 2250 608
rect 2306 574 2336 596
rect 2450 574 2480 596
rect 2536 574 2551 608
rect 2629 574 2659 601
rect 2707 635 2737 668
rect 2822 656 2852 678
rect 3094 656 3124 678
rect 3674 706 3704 734
rect 3789 696 3819 718
rect 3867 696 3897 718
rect 3982 706 4012 734
rect 3209 635 3239 668
rect 2707 574 2737 601
rect 2815 574 2830 608
rect 2886 574 2916 596
rect 3030 574 3060 596
rect 3116 574 3131 608
rect 3209 574 3239 601
rect 3287 635 3317 668
rect 3402 656 3432 678
rect 3674 656 3704 678
rect 4254 706 4284 734
rect 4369 696 4399 718
rect 4447 696 4477 718
rect 4562 706 4592 734
rect 3789 635 3819 668
rect 3287 574 3317 601
rect 3395 574 3410 608
rect 3466 574 3496 596
rect 3610 574 3640 596
rect 3696 574 3711 608
rect 3789 574 3819 601
rect 3867 635 3897 668
rect 3982 656 4012 678
rect 4254 656 4284 678
rect 4834 706 4864 734
rect 4949 696 4979 718
rect 5027 696 5057 718
rect 5142 706 5172 734
rect 4369 635 4399 668
rect 3867 574 3897 601
rect 3975 574 3990 608
rect 4046 574 4076 596
rect 4190 574 4220 596
rect 4276 574 4291 608
rect 4369 574 4399 601
rect 4447 635 4477 668
rect 4562 656 4592 678
rect 4834 656 4864 678
rect 5414 706 5444 734
rect 5529 696 5559 718
rect 5607 696 5637 718
rect 5722 706 5752 734
rect 4949 635 4979 668
rect 4447 574 4477 601
rect 4555 574 4570 608
rect 4626 574 4656 596
rect 4770 574 4800 596
rect 4856 574 4871 608
rect 4949 574 4979 601
rect 5027 635 5057 668
rect 5142 656 5172 678
rect 5414 656 5444 678
rect 5994 706 6024 734
rect 6109 696 6139 718
rect 6187 696 6217 718
rect 6302 706 6332 734
rect 5529 635 5559 668
rect 5027 574 5057 601
rect 5135 574 5150 608
rect 5206 574 5236 596
rect 5350 574 5380 596
rect 5436 574 5451 608
rect 5529 574 5559 601
rect 5607 635 5637 668
rect 5722 656 5752 678
rect 5994 656 6024 678
rect 6109 635 6139 668
rect 5607 574 5637 601
rect 5715 574 5730 608
rect 5786 574 5816 596
rect 5930 574 5960 596
rect 6016 574 6031 608
rect 6109 574 6139 601
rect 6187 635 6217 668
rect 6302 656 6332 678
rect 6187 574 6217 601
rect 6295 574 6310 608
rect 6366 574 6396 596
rect -364 560 -334 574
rect -100 560 -70 574
rect 216 560 246 574
rect 480 560 510 574
rect 796 560 826 574
rect 1060 560 1090 574
rect 1376 560 1406 574
rect 1640 560 1670 574
rect 1956 560 1986 574
rect 2220 560 2250 574
rect 2536 560 2566 574
rect 2800 560 2830 574
rect 3116 560 3146 574
rect 3380 560 3410 574
rect 3696 560 3726 574
rect 3960 560 3990 574
rect 4276 560 4306 574
rect 4540 560 4570 574
rect 4856 560 4886 574
rect 5120 560 5150 574
rect 5436 560 5466 574
rect 5700 560 5730 574
rect 6016 560 6046 574
rect 6280 560 6310 574
rect -450 510 -420 532
rect -364 510 -334 532
rect -271 510 -241 532
rect -193 510 -163 532
rect -100 510 -70 532
rect -14 510 16 532
rect 130 510 160 532
rect 216 510 246 532
rect 309 510 339 532
rect 387 510 417 532
rect 480 510 510 532
rect 566 510 596 532
rect 710 510 740 532
rect 796 510 826 532
rect 889 510 919 532
rect 967 510 997 532
rect 1060 510 1090 532
rect 1146 510 1176 532
rect 1290 510 1320 532
rect 1376 510 1406 532
rect 1469 510 1499 532
rect 1547 510 1577 532
rect 1640 510 1670 532
rect 1726 510 1756 532
rect 1870 510 1900 532
rect 1956 510 1986 532
rect 2049 510 2079 532
rect 2127 510 2157 532
rect 2220 510 2250 532
rect 2306 510 2336 532
rect 2450 510 2480 532
rect 2536 510 2566 532
rect 2629 510 2659 532
rect 2707 510 2737 532
rect 2800 510 2830 532
rect 2886 510 2916 532
rect 3030 510 3060 532
rect 3116 510 3146 532
rect 3209 510 3239 532
rect 3287 510 3317 532
rect 3380 510 3410 532
rect 3466 510 3496 532
rect 3610 510 3640 532
rect 3696 510 3726 532
rect 3789 510 3819 532
rect 3867 510 3897 532
rect 3960 510 3990 532
rect 4046 510 4076 532
rect 4190 510 4220 532
rect 4276 510 4306 532
rect 4369 510 4399 532
rect 4447 510 4477 532
rect 4540 510 4570 532
rect 4626 510 4656 532
rect 4770 510 4800 532
rect 4856 510 4886 532
rect 4949 510 4979 532
rect 5027 510 5057 532
rect 5120 510 5150 532
rect 5206 510 5236 532
rect 5350 510 5380 532
rect 5436 510 5466 532
rect 5529 510 5559 532
rect 5607 510 5637 532
rect 5700 510 5730 532
rect 5786 510 5816 532
rect 5930 510 5960 532
rect 6016 510 6046 532
rect 6109 510 6139 532
rect 6187 510 6217 532
rect 6280 510 6310 532
rect 6366 510 6396 532
rect -541 464 6439 494
rect -386 436 -356 464
rect -271 426 -241 448
rect -193 426 -163 448
rect -78 436 -48 464
rect -386 386 -356 408
rect 194 436 224 464
rect 309 426 339 448
rect 387 426 417 448
rect 502 436 532 464
rect -271 365 -241 398
rect -450 304 -420 326
rect -364 304 -349 338
rect -271 304 -241 331
rect -193 365 -163 398
rect -78 386 -48 408
rect 194 386 224 408
rect 774 436 804 464
rect 889 426 919 448
rect 967 426 997 448
rect 1082 436 1112 464
rect 309 365 339 398
rect -193 304 -163 331
rect -85 304 -70 338
rect -14 304 16 326
rect 130 304 160 326
rect 216 304 231 338
rect 309 304 339 331
rect 387 365 417 398
rect 502 386 532 408
rect 774 386 804 408
rect 1354 436 1384 464
rect 1469 426 1499 448
rect 1547 426 1577 448
rect 1662 436 1692 464
rect 889 365 919 398
rect 387 304 417 331
rect 495 304 510 338
rect 566 304 596 326
rect 710 304 740 326
rect 796 304 811 338
rect 889 304 919 331
rect 967 365 997 398
rect 1082 386 1112 408
rect 1354 386 1384 408
rect 1934 436 1964 464
rect 2049 426 2079 448
rect 2127 426 2157 448
rect 2242 436 2272 464
rect 1469 365 1499 398
rect 967 304 997 331
rect 1075 304 1090 338
rect 1146 304 1176 326
rect 1290 304 1320 326
rect 1376 304 1391 338
rect 1469 304 1499 331
rect 1547 365 1577 398
rect 1662 386 1692 408
rect 1934 386 1964 408
rect 2514 436 2544 464
rect 2629 426 2659 448
rect 2707 426 2737 448
rect 2822 436 2852 464
rect 2049 365 2079 398
rect 1547 304 1577 331
rect 1655 304 1670 338
rect 1726 304 1756 326
rect 1870 304 1900 326
rect 1956 304 1971 338
rect 2049 304 2079 331
rect 2127 365 2157 398
rect 2242 386 2272 408
rect 2514 386 2544 408
rect 3094 436 3124 464
rect 3209 426 3239 448
rect 3287 426 3317 448
rect 3402 436 3432 464
rect 2629 365 2659 398
rect 2127 304 2157 331
rect 2235 304 2250 338
rect 2306 304 2336 326
rect 2450 304 2480 326
rect 2536 304 2551 338
rect 2629 304 2659 331
rect 2707 365 2737 398
rect 2822 386 2852 408
rect 3094 386 3124 408
rect 3674 436 3704 464
rect 3789 426 3819 448
rect 3867 426 3897 448
rect 3982 436 4012 464
rect 3209 365 3239 398
rect 2707 304 2737 331
rect 2815 304 2830 338
rect 2886 304 2916 326
rect 3030 304 3060 326
rect 3116 304 3131 338
rect 3209 304 3239 331
rect 3287 365 3317 398
rect 3402 386 3432 408
rect 3674 386 3704 408
rect 4254 436 4284 464
rect 4369 426 4399 448
rect 4447 426 4477 448
rect 4562 436 4592 464
rect 3789 365 3819 398
rect 3287 304 3317 331
rect 3395 304 3410 338
rect 3466 304 3496 326
rect 3610 304 3640 326
rect 3696 304 3711 338
rect 3789 304 3819 331
rect 3867 365 3897 398
rect 3982 386 4012 408
rect 4254 386 4284 408
rect 4834 436 4864 464
rect 4949 426 4979 448
rect 5027 426 5057 448
rect 5142 436 5172 464
rect 4369 365 4399 398
rect 3867 304 3897 331
rect 3975 304 3990 338
rect 4046 304 4076 326
rect 4190 304 4220 326
rect 4276 304 4291 338
rect 4369 304 4399 331
rect 4447 365 4477 398
rect 4562 386 4592 408
rect 4834 386 4864 408
rect 5414 436 5444 464
rect 5529 426 5559 448
rect 5607 426 5637 448
rect 5722 436 5752 464
rect 4949 365 4979 398
rect 4447 304 4477 331
rect 4555 304 4570 338
rect 4626 304 4656 326
rect 4770 304 4800 326
rect 4856 304 4871 338
rect 4949 304 4979 331
rect 5027 365 5057 398
rect 5142 386 5172 408
rect 5414 386 5444 408
rect 5994 436 6024 464
rect 6109 426 6139 448
rect 6187 426 6217 448
rect 6302 436 6332 464
rect 5529 365 5559 398
rect 5027 304 5057 331
rect 5135 304 5150 338
rect 5206 304 5236 326
rect 5350 304 5380 326
rect 5436 304 5451 338
rect 5529 304 5559 331
rect 5607 365 5637 398
rect 5722 386 5752 408
rect 5994 386 6024 408
rect 6109 365 6139 398
rect 5607 304 5637 331
rect 5715 304 5730 338
rect 5786 304 5816 326
rect 5930 304 5960 326
rect 6016 304 6031 338
rect 6109 304 6139 331
rect 6187 365 6217 398
rect 6302 386 6332 408
rect 6187 304 6217 331
rect 6295 304 6310 338
rect 6366 304 6396 326
rect -364 290 -334 304
rect -100 290 -70 304
rect 216 290 246 304
rect 480 290 510 304
rect 796 290 826 304
rect 1060 290 1090 304
rect 1376 290 1406 304
rect 1640 290 1670 304
rect 1956 290 1986 304
rect 2220 290 2250 304
rect 2536 290 2566 304
rect 2800 290 2830 304
rect 3116 290 3146 304
rect 3380 290 3410 304
rect 3696 290 3726 304
rect 3960 290 3990 304
rect 4276 290 4306 304
rect 4540 290 4570 304
rect 4856 290 4886 304
rect 5120 290 5150 304
rect 5436 290 5466 304
rect 5700 290 5730 304
rect 6016 290 6046 304
rect 6280 290 6310 304
rect -450 240 -420 262
rect -364 240 -334 262
rect -271 240 -241 262
rect -193 240 -163 262
rect -100 240 -70 262
rect -14 240 16 262
rect 130 240 160 262
rect 216 240 246 262
rect 309 240 339 262
rect 387 240 417 262
rect 480 240 510 262
rect 566 240 596 262
rect 710 240 740 262
rect 796 240 826 262
rect 889 240 919 262
rect 967 240 997 262
rect 1060 240 1090 262
rect 1146 240 1176 262
rect 1290 240 1320 262
rect 1376 240 1406 262
rect 1469 240 1499 262
rect 1547 240 1577 262
rect 1640 240 1670 262
rect 1726 240 1756 262
rect 1870 240 1900 262
rect 1956 240 1986 262
rect 2049 240 2079 262
rect 2127 240 2157 262
rect 2220 240 2250 262
rect 2306 240 2336 262
rect 2450 240 2480 262
rect 2536 240 2566 262
rect 2629 240 2659 262
rect 2707 240 2737 262
rect 2800 240 2830 262
rect 2886 240 2916 262
rect 3030 240 3060 262
rect 3116 240 3146 262
rect 3209 240 3239 262
rect 3287 240 3317 262
rect 3380 240 3410 262
rect 3466 240 3496 262
rect 3610 240 3640 262
rect 3696 240 3726 262
rect 3789 240 3819 262
rect 3867 240 3897 262
rect 3960 240 3990 262
rect 4046 240 4076 262
rect 4190 240 4220 262
rect 4276 240 4306 262
rect 4369 240 4399 262
rect 4447 240 4477 262
rect 4540 240 4570 262
rect 4626 240 4656 262
rect 4770 240 4800 262
rect 4856 240 4886 262
rect 4949 240 4979 262
rect 5027 240 5057 262
rect 5120 240 5150 262
rect 5206 240 5236 262
rect 5350 240 5380 262
rect 5436 240 5466 262
rect 5529 240 5559 262
rect 5607 240 5637 262
rect 5700 240 5730 262
rect 5786 240 5816 262
rect 5930 240 5960 262
rect 6016 240 6046 262
rect 6109 240 6139 262
rect 6187 240 6217 262
rect 6280 240 6310 262
rect 6366 240 6396 262
rect -541 194 6439 224
rect -386 166 -356 194
rect -271 156 -241 178
rect -193 156 -163 178
rect -78 166 -48 194
rect -386 116 -356 138
rect 194 166 224 194
rect 309 156 339 178
rect 387 156 417 178
rect 502 166 532 194
rect -271 95 -241 128
rect -450 34 -420 56
rect -364 34 -349 68
rect -271 34 -241 61
rect -193 95 -163 128
rect -78 116 -48 138
rect 194 116 224 138
rect 774 166 804 194
rect 889 156 919 178
rect 967 156 997 178
rect 1082 166 1112 194
rect 309 95 339 128
rect -193 34 -163 61
rect -85 34 -70 68
rect -14 34 16 56
rect 130 34 160 56
rect 216 34 231 68
rect 309 34 339 61
rect 387 95 417 128
rect 502 116 532 138
rect 774 116 804 138
rect 1354 166 1384 194
rect 1469 156 1499 178
rect 1547 156 1577 178
rect 1662 166 1692 194
rect 889 95 919 128
rect 387 34 417 61
rect 495 34 510 68
rect 566 34 596 56
rect 710 34 740 56
rect 796 34 811 68
rect 889 34 919 61
rect 967 95 997 128
rect 1082 116 1112 138
rect 1354 116 1384 138
rect 1934 166 1964 194
rect 2049 156 2079 178
rect 2127 156 2157 178
rect 2242 166 2272 194
rect 1469 95 1499 128
rect 967 34 997 61
rect 1075 34 1090 68
rect 1146 34 1176 56
rect 1290 34 1320 56
rect 1376 34 1391 68
rect 1469 34 1499 61
rect 1547 95 1577 128
rect 1662 116 1692 138
rect 1934 116 1964 138
rect 2514 166 2544 194
rect 2629 156 2659 178
rect 2707 156 2737 178
rect 2822 166 2852 194
rect 2049 95 2079 128
rect 1547 34 1577 61
rect 1655 34 1670 68
rect 1726 34 1756 56
rect 1870 34 1900 56
rect 1956 34 1971 68
rect 2049 34 2079 61
rect 2127 95 2157 128
rect 2242 116 2272 138
rect 2514 116 2544 138
rect 3094 166 3124 194
rect 3209 156 3239 178
rect 3287 156 3317 178
rect 3402 166 3432 194
rect 2629 95 2659 128
rect 2127 34 2157 61
rect 2235 34 2250 68
rect 2306 34 2336 56
rect 2450 34 2480 56
rect 2536 34 2551 68
rect 2629 34 2659 61
rect 2707 95 2737 128
rect 2822 116 2852 138
rect 3094 116 3124 138
rect 3674 166 3704 194
rect 3789 156 3819 178
rect 3867 156 3897 178
rect 3982 166 4012 194
rect 3209 95 3239 128
rect 2707 34 2737 61
rect 2815 34 2830 68
rect 2886 34 2916 56
rect 3030 34 3060 56
rect 3116 34 3131 68
rect 3209 34 3239 61
rect 3287 95 3317 128
rect 3402 116 3432 138
rect 3674 116 3704 138
rect 4254 166 4284 194
rect 4369 156 4399 178
rect 4447 156 4477 178
rect 4562 166 4592 194
rect 3789 95 3819 128
rect 3287 34 3317 61
rect 3395 34 3410 68
rect 3466 34 3496 56
rect 3610 34 3640 56
rect 3696 34 3711 68
rect 3789 34 3819 61
rect 3867 95 3897 128
rect 3982 116 4012 138
rect 4254 116 4284 138
rect 4834 166 4864 194
rect 4949 156 4979 178
rect 5027 156 5057 178
rect 5142 166 5172 194
rect 4369 95 4399 128
rect 3867 34 3897 61
rect 3975 34 3990 68
rect 4046 34 4076 56
rect 4190 34 4220 56
rect 4276 34 4291 68
rect 4369 34 4399 61
rect 4447 95 4477 128
rect 4562 116 4592 138
rect 4834 116 4864 138
rect 5414 166 5444 194
rect 5529 156 5559 178
rect 5607 156 5637 178
rect 5722 166 5752 194
rect 4949 95 4979 128
rect 4447 34 4477 61
rect 4555 34 4570 68
rect 4626 34 4656 56
rect 4770 34 4800 56
rect 4856 34 4871 68
rect 4949 34 4979 61
rect 5027 95 5057 128
rect 5142 116 5172 138
rect 5414 116 5444 138
rect 5994 166 6024 194
rect 6109 156 6139 178
rect 6187 156 6217 178
rect 6302 166 6332 194
rect 5529 95 5559 128
rect 5027 34 5057 61
rect 5135 34 5150 68
rect 5206 34 5236 56
rect 5350 34 5380 56
rect 5436 34 5451 68
rect 5529 34 5559 61
rect 5607 95 5637 128
rect 5722 116 5752 138
rect 5994 116 6024 138
rect 6109 95 6139 128
rect 5607 34 5637 61
rect 5715 34 5730 68
rect 5786 34 5816 56
rect 5930 34 5960 56
rect 6016 34 6031 68
rect 6109 34 6139 61
rect 6187 95 6217 128
rect 6302 116 6332 138
rect 6187 34 6217 61
rect 6295 34 6310 68
rect 6366 34 6396 56
rect -364 20 -334 34
rect -100 20 -70 34
rect 216 20 246 34
rect 480 20 510 34
rect 796 20 826 34
rect 1060 20 1090 34
rect 1376 20 1406 34
rect 1640 20 1670 34
rect 1956 20 1986 34
rect 2220 20 2250 34
rect 2536 20 2566 34
rect 2800 20 2830 34
rect 3116 20 3146 34
rect 3380 20 3410 34
rect 3696 20 3726 34
rect 3960 20 3990 34
rect 4276 20 4306 34
rect 4540 20 4570 34
rect 4856 20 4886 34
rect 5120 20 5150 34
rect 5436 20 5466 34
rect 5700 20 5730 34
rect 6016 20 6046 34
rect 6280 20 6310 34
rect -450 -30 -420 -8
rect -364 -30 -334 -8
rect -271 -30 -241 -8
rect -193 -30 -163 -8
rect -100 -30 -70 -8
rect -14 -30 16 -8
rect 130 -30 160 -8
rect 216 -30 246 -8
rect 309 -30 339 -8
rect 387 -30 417 -8
rect 480 -30 510 -8
rect 566 -30 596 -8
rect 710 -30 740 -8
rect 796 -30 826 -8
rect 889 -30 919 -8
rect 967 -30 997 -8
rect 1060 -30 1090 -8
rect 1146 -30 1176 -8
rect 1290 -30 1320 -8
rect 1376 -30 1406 -8
rect 1469 -30 1499 -8
rect 1547 -30 1577 -8
rect 1640 -30 1670 -8
rect 1726 -30 1756 -8
rect 1870 -30 1900 -8
rect 1956 -30 1986 -8
rect 2049 -30 2079 -8
rect 2127 -30 2157 -8
rect 2220 -30 2250 -8
rect 2306 -30 2336 -8
rect 2450 -30 2480 -8
rect 2536 -30 2566 -8
rect 2629 -30 2659 -8
rect 2707 -30 2737 -8
rect 2800 -30 2830 -8
rect 2886 -30 2916 -8
rect 3030 -30 3060 -8
rect 3116 -30 3146 -8
rect 3209 -30 3239 -8
rect 3287 -30 3317 -8
rect 3380 -30 3410 -8
rect 3466 -30 3496 -8
rect 3610 -30 3640 -8
rect 3696 -30 3726 -8
rect 3789 -30 3819 -8
rect 3867 -30 3897 -8
rect 3960 -30 3990 -8
rect 4046 -30 4076 -8
rect 4190 -30 4220 -8
rect 4276 -30 4306 -8
rect 4369 -30 4399 -8
rect 4447 -30 4477 -8
rect 4540 -30 4570 -8
rect 4626 -30 4656 -8
rect 4770 -30 4800 -8
rect 4856 -30 4886 -8
rect 4949 -30 4979 -8
rect 5027 -30 5057 -8
rect 5120 -30 5150 -8
rect 5206 -30 5236 -8
rect 5350 -30 5380 -8
rect 5436 -30 5466 -8
rect 5529 -30 5559 -8
rect 5607 -30 5637 -8
rect 5700 -30 5730 -8
rect 5786 -30 5816 -8
rect 5930 -30 5960 -8
rect 6016 -30 6046 -8
rect 6109 -30 6139 -8
rect 6187 -30 6217 -8
rect 6280 -30 6310 -8
rect 6366 -30 6396 -8
rect -541 -76 6439 -46
rect -386 -104 -356 -76
rect -271 -114 -241 -92
rect -193 -114 -163 -92
rect -78 -104 -48 -76
rect -386 -154 -356 -132
rect 194 -104 224 -76
rect 309 -114 339 -92
rect 387 -114 417 -92
rect 502 -104 532 -76
rect -271 -175 -241 -142
rect -450 -236 -420 -214
rect -364 -236 -349 -202
rect -271 -236 -241 -209
rect -193 -175 -163 -142
rect -78 -154 -48 -132
rect 194 -154 224 -132
rect 774 -104 804 -76
rect 889 -114 919 -92
rect 967 -114 997 -92
rect 1082 -104 1112 -76
rect 309 -175 339 -142
rect -193 -236 -163 -209
rect -85 -236 -70 -202
rect -14 -236 16 -214
rect 130 -236 160 -214
rect 216 -236 231 -202
rect 309 -236 339 -209
rect 387 -175 417 -142
rect 502 -154 532 -132
rect 774 -154 804 -132
rect 1354 -104 1384 -76
rect 1469 -114 1499 -92
rect 1547 -114 1577 -92
rect 1662 -104 1692 -76
rect 889 -175 919 -142
rect 387 -236 417 -209
rect 495 -236 510 -202
rect 566 -236 596 -214
rect 710 -236 740 -214
rect 796 -236 811 -202
rect 889 -236 919 -209
rect 967 -175 997 -142
rect 1082 -154 1112 -132
rect 1354 -154 1384 -132
rect 1934 -104 1964 -76
rect 2049 -114 2079 -92
rect 2127 -114 2157 -92
rect 2242 -104 2272 -76
rect 1469 -175 1499 -142
rect 967 -236 997 -209
rect 1075 -236 1090 -202
rect 1146 -236 1176 -214
rect 1290 -236 1320 -214
rect 1376 -236 1391 -202
rect 1469 -236 1499 -209
rect 1547 -175 1577 -142
rect 1662 -154 1692 -132
rect 1934 -154 1964 -132
rect 2514 -104 2544 -76
rect 2629 -114 2659 -92
rect 2707 -114 2737 -92
rect 2822 -104 2852 -76
rect 2049 -175 2079 -142
rect 1547 -236 1577 -209
rect 1655 -236 1670 -202
rect 1726 -236 1756 -214
rect 1870 -236 1900 -214
rect 1956 -236 1971 -202
rect 2049 -236 2079 -209
rect 2127 -175 2157 -142
rect 2242 -154 2272 -132
rect 2514 -154 2544 -132
rect 3094 -104 3124 -76
rect 3209 -114 3239 -92
rect 3287 -114 3317 -92
rect 3402 -104 3432 -76
rect 2629 -175 2659 -142
rect 2127 -236 2157 -209
rect 2235 -236 2250 -202
rect 2306 -236 2336 -214
rect 2450 -236 2480 -214
rect 2536 -236 2551 -202
rect 2629 -236 2659 -209
rect 2707 -175 2737 -142
rect 2822 -154 2852 -132
rect 3094 -154 3124 -132
rect 3674 -104 3704 -76
rect 3789 -114 3819 -92
rect 3867 -114 3897 -92
rect 3982 -104 4012 -76
rect 3209 -175 3239 -142
rect 2707 -236 2737 -209
rect 2815 -236 2830 -202
rect 2886 -236 2916 -214
rect 3030 -236 3060 -214
rect 3116 -236 3131 -202
rect 3209 -236 3239 -209
rect 3287 -175 3317 -142
rect 3402 -154 3432 -132
rect 3674 -154 3704 -132
rect 4254 -104 4284 -76
rect 4369 -114 4399 -92
rect 4447 -114 4477 -92
rect 4562 -104 4592 -76
rect 3789 -175 3819 -142
rect 3287 -236 3317 -209
rect 3395 -236 3410 -202
rect 3466 -236 3496 -214
rect 3610 -236 3640 -214
rect 3696 -236 3711 -202
rect 3789 -236 3819 -209
rect 3867 -175 3897 -142
rect 3982 -154 4012 -132
rect 4254 -154 4284 -132
rect 4834 -104 4864 -76
rect 4949 -114 4979 -92
rect 5027 -114 5057 -92
rect 5142 -104 5172 -76
rect 4369 -175 4399 -142
rect 3867 -236 3897 -209
rect 3975 -236 3990 -202
rect 4046 -236 4076 -214
rect 4190 -236 4220 -214
rect 4276 -236 4291 -202
rect 4369 -236 4399 -209
rect 4447 -175 4477 -142
rect 4562 -154 4592 -132
rect 4834 -154 4864 -132
rect 5414 -104 5444 -76
rect 5529 -114 5559 -92
rect 5607 -114 5637 -92
rect 5722 -104 5752 -76
rect 4949 -175 4979 -142
rect 4447 -236 4477 -209
rect 4555 -236 4570 -202
rect 4626 -236 4656 -214
rect 4770 -236 4800 -214
rect 4856 -236 4871 -202
rect 4949 -236 4979 -209
rect 5027 -175 5057 -142
rect 5142 -154 5172 -132
rect 5414 -154 5444 -132
rect 5994 -104 6024 -76
rect 6109 -114 6139 -92
rect 6187 -114 6217 -92
rect 6302 -104 6332 -76
rect 5529 -175 5559 -142
rect 5027 -236 5057 -209
rect 5135 -236 5150 -202
rect 5206 -236 5236 -214
rect 5350 -236 5380 -214
rect 5436 -236 5451 -202
rect 5529 -236 5559 -209
rect 5607 -175 5637 -142
rect 5722 -154 5752 -132
rect 5994 -154 6024 -132
rect 6109 -175 6139 -142
rect 5607 -236 5637 -209
rect 5715 -236 5730 -202
rect 5786 -236 5816 -214
rect 5930 -236 5960 -214
rect 6016 -236 6031 -202
rect 6109 -236 6139 -209
rect 6187 -175 6217 -142
rect 6302 -154 6332 -132
rect 6187 -236 6217 -209
rect 6295 -236 6310 -202
rect 6366 -236 6396 -214
rect -364 -250 -334 -236
rect -100 -250 -70 -236
rect 216 -250 246 -236
rect 480 -250 510 -236
rect 796 -250 826 -236
rect 1060 -250 1090 -236
rect 1376 -250 1406 -236
rect 1640 -250 1670 -236
rect 1956 -250 1986 -236
rect 2220 -250 2250 -236
rect 2536 -250 2566 -236
rect 2800 -250 2830 -236
rect 3116 -250 3146 -236
rect 3380 -250 3410 -236
rect 3696 -250 3726 -236
rect 3960 -250 3990 -236
rect 4276 -250 4306 -236
rect 4540 -250 4570 -236
rect 4856 -250 4886 -236
rect 5120 -250 5150 -236
rect 5436 -250 5466 -236
rect 5700 -250 5730 -236
rect 6016 -250 6046 -236
rect 6280 -250 6310 -236
rect -450 -300 -420 -278
rect -364 -300 -334 -278
rect -271 -300 -241 -278
rect -193 -300 -163 -278
rect -100 -300 -70 -278
rect -14 -300 16 -278
rect 130 -300 160 -278
rect 216 -300 246 -278
rect 309 -300 339 -278
rect 387 -300 417 -278
rect 480 -300 510 -278
rect 566 -300 596 -278
rect 710 -300 740 -278
rect 796 -300 826 -278
rect 889 -300 919 -278
rect 967 -300 997 -278
rect 1060 -300 1090 -278
rect 1146 -300 1176 -278
rect 1290 -300 1320 -278
rect 1376 -300 1406 -278
rect 1469 -300 1499 -278
rect 1547 -300 1577 -278
rect 1640 -300 1670 -278
rect 1726 -300 1756 -278
rect 1870 -300 1900 -278
rect 1956 -300 1986 -278
rect 2049 -300 2079 -278
rect 2127 -300 2157 -278
rect 2220 -300 2250 -278
rect 2306 -300 2336 -278
rect 2450 -300 2480 -278
rect 2536 -300 2566 -278
rect 2629 -300 2659 -278
rect 2707 -300 2737 -278
rect 2800 -300 2830 -278
rect 2886 -300 2916 -278
rect 3030 -300 3060 -278
rect 3116 -300 3146 -278
rect 3209 -300 3239 -278
rect 3287 -300 3317 -278
rect 3380 -300 3410 -278
rect 3466 -300 3496 -278
rect 3610 -300 3640 -278
rect 3696 -300 3726 -278
rect 3789 -300 3819 -278
rect 3867 -300 3897 -278
rect 3960 -300 3990 -278
rect 4046 -300 4076 -278
rect 4190 -300 4220 -278
rect 4276 -300 4306 -278
rect 4369 -300 4399 -278
rect 4447 -300 4477 -278
rect 4540 -300 4570 -278
rect 4626 -300 4656 -278
rect 4770 -300 4800 -278
rect 4856 -300 4886 -278
rect 4949 -300 4979 -278
rect 5027 -300 5057 -278
rect 5120 -300 5150 -278
rect 5206 -300 5236 -278
rect 5350 -300 5380 -278
rect 5436 -300 5466 -278
rect 5529 -300 5559 -278
rect 5607 -300 5637 -278
rect 5700 -300 5730 -278
rect 5786 -300 5816 -278
rect 5930 -300 5960 -278
rect 6016 -300 6046 -278
rect 6109 -300 6139 -278
rect 6187 -300 6217 -278
rect 6280 -300 6310 -278
rect 6366 -300 6396 -278
rect -541 -346 6439 -316
rect -386 -374 -356 -346
rect -271 -384 -241 -362
rect -193 -384 -163 -362
rect -78 -374 -48 -346
rect -386 -424 -356 -402
rect 194 -374 224 -346
rect 309 -384 339 -362
rect 387 -384 417 -362
rect 502 -374 532 -346
rect -271 -445 -241 -412
rect -450 -506 -420 -484
rect -364 -506 -349 -472
rect -271 -506 -241 -479
rect -193 -445 -163 -412
rect -78 -424 -48 -402
rect 194 -424 224 -402
rect 774 -374 804 -346
rect 889 -384 919 -362
rect 967 -384 997 -362
rect 1082 -374 1112 -346
rect 309 -445 339 -412
rect -193 -506 -163 -479
rect -85 -506 -70 -472
rect -14 -506 16 -484
rect 130 -506 160 -484
rect 216 -506 231 -472
rect 309 -506 339 -479
rect 387 -445 417 -412
rect 502 -424 532 -402
rect 774 -424 804 -402
rect 1354 -374 1384 -346
rect 1469 -384 1499 -362
rect 1547 -384 1577 -362
rect 1662 -374 1692 -346
rect 889 -445 919 -412
rect 387 -506 417 -479
rect 495 -506 510 -472
rect 566 -506 596 -484
rect 710 -506 740 -484
rect 796 -506 811 -472
rect 889 -506 919 -479
rect 967 -445 997 -412
rect 1082 -424 1112 -402
rect 1354 -424 1384 -402
rect 1934 -374 1964 -346
rect 2049 -384 2079 -362
rect 2127 -384 2157 -362
rect 2242 -374 2272 -346
rect 1469 -445 1499 -412
rect 967 -506 997 -479
rect 1075 -506 1090 -472
rect 1146 -506 1176 -484
rect 1290 -506 1320 -484
rect 1376 -506 1391 -472
rect 1469 -506 1499 -479
rect 1547 -445 1577 -412
rect 1662 -424 1692 -402
rect 1934 -424 1964 -402
rect 2514 -374 2544 -346
rect 2629 -384 2659 -362
rect 2707 -384 2737 -362
rect 2822 -374 2852 -346
rect 2049 -445 2079 -412
rect 1547 -506 1577 -479
rect 1655 -506 1670 -472
rect 1726 -506 1756 -484
rect 1870 -506 1900 -484
rect 1956 -506 1971 -472
rect 2049 -506 2079 -479
rect 2127 -445 2157 -412
rect 2242 -424 2272 -402
rect 2514 -424 2544 -402
rect 3094 -374 3124 -346
rect 3209 -384 3239 -362
rect 3287 -384 3317 -362
rect 3402 -374 3432 -346
rect 2629 -445 2659 -412
rect 2127 -506 2157 -479
rect 2235 -506 2250 -472
rect 2306 -506 2336 -484
rect 2450 -506 2480 -484
rect 2536 -506 2551 -472
rect 2629 -506 2659 -479
rect 2707 -445 2737 -412
rect 2822 -424 2852 -402
rect 3094 -424 3124 -402
rect 3674 -374 3704 -346
rect 3789 -384 3819 -362
rect 3867 -384 3897 -362
rect 3982 -374 4012 -346
rect 3209 -445 3239 -412
rect 2707 -506 2737 -479
rect 2815 -506 2830 -472
rect 2886 -506 2916 -484
rect 3030 -506 3060 -484
rect 3116 -506 3131 -472
rect 3209 -506 3239 -479
rect 3287 -445 3317 -412
rect 3402 -424 3432 -402
rect 3674 -424 3704 -402
rect 4254 -374 4284 -346
rect 4369 -384 4399 -362
rect 4447 -384 4477 -362
rect 4562 -374 4592 -346
rect 3789 -445 3819 -412
rect 3287 -506 3317 -479
rect 3395 -506 3410 -472
rect 3466 -506 3496 -484
rect 3610 -506 3640 -484
rect 3696 -506 3711 -472
rect 3789 -506 3819 -479
rect 3867 -445 3897 -412
rect 3982 -424 4012 -402
rect 4254 -424 4284 -402
rect 4834 -374 4864 -346
rect 4949 -384 4979 -362
rect 5027 -384 5057 -362
rect 5142 -374 5172 -346
rect 4369 -445 4399 -412
rect 3867 -506 3897 -479
rect 3975 -506 3990 -472
rect 4046 -506 4076 -484
rect 4190 -506 4220 -484
rect 4276 -506 4291 -472
rect 4369 -506 4399 -479
rect 4447 -445 4477 -412
rect 4562 -424 4592 -402
rect 4834 -424 4864 -402
rect 5414 -374 5444 -346
rect 5529 -384 5559 -362
rect 5607 -384 5637 -362
rect 5722 -374 5752 -346
rect 4949 -445 4979 -412
rect 4447 -506 4477 -479
rect 4555 -506 4570 -472
rect 4626 -506 4656 -484
rect 4770 -506 4800 -484
rect 4856 -506 4871 -472
rect 4949 -506 4979 -479
rect 5027 -445 5057 -412
rect 5142 -424 5172 -402
rect 5414 -424 5444 -402
rect 5994 -374 6024 -346
rect 6109 -384 6139 -362
rect 6187 -384 6217 -362
rect 6302 -374 6332 -346
rect 5529 -445 5559 -412
rect 5027 -506 5057 -479
rect 5135 -506 5150 -472
rect 5206 -506 5236 -484
rect 5350 -506 5380 -484
rect 5436 -506 5451 -472
rect 5529 -506 5559 -479
rect 5607 -445 5637 -412
rect 5722 -424 5752 -402
rect 5994 -424 6024 -402
rect 6109 -445 6139 -412
rect 5607 -506 5637 -479
rect 5715 -506 5730 -472
rect 5786 -506 5816 -484
rect 5930 -506 5960 -484
rect 6016 -506 6031 -472
rect 6109 -506 6139 -479
rect 6187 -445 6217 -412
rect 6302 -424 6332 -402
rect 6187 -506 6217 -479
rect 6295 -506 6310 -472
rect 6366 -506 6396 -484
rect -364 -520 -334 -506
rect -100 -520 -70 -506
rect 216 -520 246 -506
rect 480 -520 510 -506
rect 796 -520 826 -506
rect 1060 -520 1090 -506
rect 1376 -520 1406 -506
rect 1640 -520 1670 -506
rect 1956 -520 1986 -506
rect 2220 -520 2250 -506
rect 2536 -520 2566 -506
rect 2800 -520 2830 -506
rect 3116 -520 3146 -506
rect 3380 -520 3410 -506
rect 3696 -520 3726 -506
rect 3960 -520 3990 -506
rect 4276 -520 4306 -506
rect 4540 -520 4570 -506
rect 4856 -520 4886 -506
rect 5120 -520 5150 -506
rect 5436 -520 5466 -506
rect 5700 -520 5730 -506
rect 6016 -520 6046 -506
rect 6280 -520 6310 -506
rect -450 -570 -420 -548
rect -364 -570 -334 -548
rect -271 -570 -241 -548
rect -193 -570 -163 -548
rect -100 -570 -70 -548
rect -14 -570 16 -548
rect 130 -570 160 -548
rect 216 -570 246 -548
rect 309 -570 339 -548
rect 387 -570 417 -548
rect 480 -570 510 -548
rect 566 -570 596 -548
rect 710 -570 740 -548
rect 796 -570 826 -548
rect 889 -570 919 -548
rect 967 -570 997 -548
rect 1060 -570 1090 -548
rect 1146 -570 1176 -548
rect 1290 -570 1320 -548
rect 1376 -570 1406 -548
rect 1469 -570 1499 -548
rect 1547 -570 1577 -548
rect 1640 -570 1670 -548
rect 1726 -570 1756 -548
rect 1870 -570 1900 -548
rect 1956 -570 1986 -548
rect 2049 -570 2079 -548
rect 2127 -570 2157 -548
rect 2220 -570 2250 -548
rect 2306 -570 2336 -548
rect 2450 -570 2480 -548
rect 2536 -570 2566 -548
rect 2629 -570 2659 -548
rect 2707 -570 2737 -548
rect 2800 -570 2830 -548
rect 2886 -570 2916 -548
rect 3030 -570 3060 -548
rect 3116 -570 3146 -548
rect 3209 -570 3239 -548
rect 3287 -570 3317 -548
rect 3380 -570 3410 -548
rect 3466 -570 3496 -548
rect 3610 -570 3640 -548
rect 3696 -570 3726 -548
rect 3789 -570 3819 -548
rect 3867 -570 3897 -548
rect 3960 -570 3990 -548
rect 4046 -570 4076 -548
rect 4190 -570 4220 -548
rect 4276 -570 4306 -548
rect 4369 -570 4399 -548
rect 4447 -570 4477 -548
rect 4540 -570 4570 -548
rect 4626 -570 4656 -548
rect 4770 -570 4800 -548
rect 4856 -570 4886 -548
rect 4949 -570 4979 -548
rect 5027 -570 5057 -548
rect 5120 -570 5150 -548
rect 5206 -570 5236 -548
rect 5350 -570 5380 -548
rect 5436 -570 5466 -548
rect 5529 -570 5559 -548
rect 5607 -570 5637 -548
rect 5700 -570 5730 -548
rect 5786 -570 5816 -548
rect 5930 -570 5960 -548
rect 6016 -570 6046 -548
rect 6109 -570 6139 -548
rect 6187 -570 6217 -548
rect 6280 -570 6310 -548
rect 6366 -570 6396 -548
rect -541 -616 6439 -586
rect -386 -644 -356 -616
rect -271 -654 -241 -632
rect -193 -654 -163 -632
rect -78 -644 -48 -616
rect -386 -694 -356 -672
rect 194 -644 224 -616
rect 309 -654 339 -632
rect 387 -654 417 -632
rect 502 -644 532 -616
rect -271 -715 -241 -682
rect -450 -776 -420 -754
rect -364 -776 -349 -742
rect -271 -776 -241 -749
rect -193 -715 -163 -682
rect -78 -694 -48 -672
rect 194 -694 224 -672
rect 774 -644 804 -616
rect 889 -654 919 -632
rect 967 -654 997 -632
rect 1082 -644 1112 -616
rect 309 -715 339 -682
rect -193 -776 -163 -749
rect -85 -776 -70 -742
rect -14 -776 16 -754
rect 130 -776 160 -754
rect 216 -776 231 -742
rect 309 -776 339 -749
rect 387 -715 417 -682
rect 502 -694 532 -672
rect 774 -694 804 -672
rect 1354 -644 1384 -616
rect 1469 -654 1499 -632
rect 1547 -654 1577 -632
rect 1662 -644 1692 -616
rect 889 -715 919 -682
rect 387 -776 417 -749
rect 495 -776 510 -742
rect 566 -776 596 -754
rect 710 -776 740 -754
rect 796 -776 811 -742
rect 889 -776 919 -749
rect 967 -715 997 -682
rect 1082 -694 1112 -672
rect 1354 -694 1384 -672
rect 1934 -644 1964 -616
rect 2049 -654 2079 -632
rect 2127 -654 2157 -632
rect 2242 -644 2272 -616
rect 1469 -715 1499 -682
rect 967 -776 997 -749
rect 1075 -776 1090 -742
rect 1146 -776 1176 -754
rect 1290 -776 1320 -754
rect 1376 -776 1391 -742
rect 1469 -776 1499 -749
rect 1547 -715 1577 -682
rect 1662 -694 1692 -672
rect 1934 -694 1964 -672
rect 2514 -644 2544 -616
rect 2629 -654 2659 -632
rect 2707 -654 2737 -632
rect 2822 -644 2852 -616
rect 2049 -715 2079 -682
rect 1547 -776 1577 -749
rect 1655 -776 1670 -742
rect 1726 -776 1756 -754
rect 1870 -776 1900 -754
rect 1956 -776 1971 -742
rect 2049 -776 2079 -749
rect 2127 -715 2157 -682
rect 2242 -694 2272 -672
rect 2514 -694 2544 -672
rect 3094 -644 3124 -616
rect 3209 -654 3239 -632
rect 3287 -654 3317 -632
rect 3402 -644 3432 -616
rect 2629 -715 2659 -682
rect 2127 -776 2157 -749
rect 2235 -776 2250 -742
rect 2306 -776 2336 -754
rect 2450 -776 2480 -754
rect 2536 -776 2551 -742
rect 2629 -776 2659 -749
rect 2707 -715 2737 -682
rect 2822 -694 2852 -672
rect 3094 -694 3124 -672
rect 3674 -644 3704 -616
rect 3789 -654 3819 -632
rect 3867 -654 3897 -632
rect 3982 -644 4012 -616
rect 3209 -715 3239 -682
rect 2707 -776 2737 -749
rect 2815 -776 2830 -742
rect 2886 -776 2916 -754
rect 3030 -776 3060 -754
rect 3116 -776 3131 -742
rect 3209 -776 3239 -749
rect 3287 -715 3317 -682
rect 3402 -694 3432 -672
rect 3674 -694 3704 -672
rect 4254 -644 4284 -616
rect 4369 -654 4399 -632
rect 4447 -654 4477 -632
rect 4562 -644 4592 -616
rect 3789 -715 3819 -682
rect 3287 -776 3317 -749
rect 3395 -776 3410 -742
rect 3466 -776 3496 -754
rect 3610 -776 3640 -754
rect 3696 -776 3711 -742
rect 3789 -776 3819 -749
rect 3867 -715 3897 -682
rect 3982 -694 4012 -672
rect 4254 -694 4284 -672
rect 4834 -644 4864 -616
rect 4949 -654 4979 -632
rect 5027 -654 5057 -632
rect 5142 -644 5172 -616
rect 4369 -715 4399 -682
rect 3867 -776 3897 -749
rect 3975 -776 3990 -742
rect 4046 -776 4076 -754
rect 4190 -776 4220 -754
rect 4276 -776 4291 -742
rect 4369 -776 4399 -749
rect 4447 -715 4477 -682
rect 4562 -694 4592 -672
rect 4834 -694 4864 -672
rect 5414 -644 5444 -616
rect 5529 -654 5559 -632
rect 5607 -654 5637 -632
rect 5722 -644 5752 -616
rect 4949 -715 4979 -682
rect 4447 -776 4477 -749
rect 4555 -776 4570 -742
rect 4626 -776 4656 -754
rect 4770 -776 4800 -754
rect 4856 -776 4871 -742
rect 4949 -776 4979 -749
rect 5027 -715 5057 -682
rect 5142 -694 5172 -672
rect 5414 -694 5444 -672
rect 5994 -644 6024 -616
rect 6109 -654 6139 -632
rect 6187 -654 6217 -632
rect 6302 -644 6332 -616
rect 5529 -715 5559 -682
rect 5027 -776 5057 -749
rect 5135 -776 5150 -742
rect 5206 -776 5236 -754
rect 5350 -776 5380 -754
rect 5436 -776 5451 -742
rect 5529 -776 5559 -749
rect 5607 -715 5637 -682
rect 5722 -694 5752 -672
rect 5994 -694 6024 -672
rect 6109 -715 6139 -682
rect 5607 -776 5637 -749
rect 5715 -776 5730 -742
rect 5786 -776 5816 -754
rect 5930 -776 5960 -754
rect 6016 -776 6031 -742
rect 6109 -776 6139 -749
rect 6187 -715 6217 -682
rect 6302 -694 6332 -672
rect 6187 -776 6217 -749
rect 6295 -776 6310 -742
rect 6366 -776 6396 -754
rect -364 -790 -334 -776
rect -100 -790 -70 -776
rect 216 -790 246 -776
rect 480 -790 510 -776
rect 796 -790 826 -776
rect 1060 -790 1090 -776
rect 1376 -790 1406 -776
rect 1640 -790 1670 -776
rect 1956 -790 1986 -776
rect 2220 -790 2250 -776
rect 2536 -790 2566 -776
rect 2800 -790 2830 -776
rect 3116 -790 3146 -776
rect 3380 -790 3410 -776
rect 3696 -790 3726 -776
rect 3960 -790 3990 -776
rect 4276 -790 4306 -776
rect 4540 -790 4570 -776
rect 4856 -790 4886 -776
rect 5120 -790 5150 -776
rect 5436 -790 5466 -776
rect 5700 -790 5730 -776
rect 6016 -790 6046 -776
rect 6280 -790 6310 -776
rect -450 -840 -420 -818
rect -364 -840 -334 -818
rect -271 -840 -241 -818
rect -193 -840 -163 -818
rect -100 -840 -70 -818
rect -14 -840 16 -818
rect 130 -840 160 -818
rect 216 -840 246 -818
rect 309 -840 339 -818
rect 387 -840 417 -818
rect 480 -840 510 -818
rect 566 -840 596 -818
rect 710 -840 740 -818
rect 796 -840 826 -818
rect 889 -840 919 -818
rect 967 -840 997 -818
rect 1060 -840 1090 -818
rect 1146 -840 1176 -818
rect 1290 -840 1320 -818
rect 1376 -840 1406 -818
rect 1469 -840 1499 -818
rect 1547 -840 1577 -818
rect 1640 -840 1670 -818
rect 1726 -840 1756 -818
rect 1870 -840 1900 -818
rect 1956 -840 1986 -818
rect 2049 -840 2079 -818
rect 2127 -840 2157 -818
rect 2220 -840 2250 -818
rect 2306 -840 2336 -818
rect 2450 -840 2480 -818
rect 2536 -840 2566 -818
rect 2629 -840 2659 -818
rect 2707 -840 2737 -818
rect 2800 -840 2830 -818
rect 2886 -840 2916 -818
rect 3030 -840 3060 -818
rect 3116 -840 3146 -818
rect 3209 -840 3239 -818
rect 3287 -840 3317 -818
rect 3380 -840 3410 -818
rect 3466 -840 3496 -818
rect 3610 -840 3640 -818
rect 3696 -840 3726 -818
rect 3789 -840 3819 -818
rect 3867 -840 3897 -818
rect 3960 -840 3990 -818
rect 4046 -840 4076 -818
rect 4190 -840 4220 -818
rect 4276 -840 4306 -818
rect 4369 -840 4399 -818
rect 4447 -840 4477 -818
rect 4540 -840 4570 -818
rect 4626 -840 4656 -818
rect 4770 -840 4800 -818
rect 4856 -840 4886 -818
rect 4949 -840 4979 -818
rect 5027 -840 5057 -818
rect 5120 -840 5150 -818
rect 5206 -840 5236 -818
rect 5350 -840 5380 -818
rect 5436 -840 5466 -818
rect 5529 -840 5559 -818
rect 5607 -840 5637 -818
rect 5700 -840 5730 -818
rect 5786 -840 5816 -818
rect 5930 -840 5960 -818
rect 6016 -840 6046 -818
rect 6109 -840 6139 -818
rect 6187 -840 6217 -818
rect 6280 -840 6310 -818
rect 6366 -840 6396 -818
rect -541 -886 6439 -856
rect -386 -914 -356 -886
rect -271 -924 -241 -902
rect -193 -924 -163 -902
rect -78 -914 -48 -886
rect -386 -964 -356 -942
rect 194 -914 224 -886
rect 309 -924 339 -902
rect 387 -924 417 -902
rect 502 -914 532 -886
rect -271 -985 -241 -952
rect -450 -1046 -420 -1024
rect -364 -1046 -349 -1012
rect -271 -1046 -241 -1019
rect -193 -985 -163 -952
rect -78 -964 -48 -942
rect 194 -964 224 -942
rect 774 -914 804 -886
rect 889 -924 919 -902
rect 967 -924 997 -902
rect 1082 -914 1112 -886
rect 309 -985 339 -952
rect -193 -1046 -163 -1019
rect -85 -1046 -70 -1012
rect -14 -1046 16 -1024
rect 130 -1046 160 -1024
rect 216 -1046 231 -1012
rect 309 -1046 339 -1019
rect 387 -985 417 -952
rect 502 -964 532 -942
rect 774 -964 804 -942
rect 1354 -914 1384 -886
rect 1469 -924 1499 -902
rect 1547 -924 1577 -902
rect 1662 -914 1692 -886
rect 889 -985 919 -952
rect 387 -1046 417 -1019
rect 495 -1046 510 -1012
rect 566 -1046 596 -1024
rect 710 -1046 740 -1024
rect 796 -1046 811 -1012
rect 889 -1046 919 -1019
rect 967 -985 997 -952
rect 1082 -964 1112 -942
rect 1354 -964 1384 -942
rect 1934 -914 1964 -886
rect 2049 -924 2079 -902
rect 2127 -924 2157 -902
rect 2242 -914 2272 -886
rect 1469 -985 1499 -952
rect 967 -1046 997 -1019
rect 1075 -1046 1090 -1012
rect 1146 -1046 1176 -1024
rect 1290 -1046 1320 -1024
rect 1376 -1046 1391 -1012
rect 1469 -1046 1499 -1019
rect 1547 -985 1577 -952
rect 1662 -964 1692 -942
rect 1934 -964 1964 -942
rect 2514 -914 2544 -886
rect 2629 -924 2659 -902
rect 2707 -924 2737 -902
rect 2822 -914 2852 -886
rect 2049 -985 2079 -952
rect 1547 -1046 1577 -1019
rect 1655 -1046 1670 -1012
rect 1726 -1046 1756 -1024
rect 1870 -1046 1900 -1024
rect 1956 -1046 1971 -1012
rect 2049 -1046 2079 -1019
rect 2127 -985 2157 -952
rect 2242 -964 2272 -942
rect 2514 -964 2544 -942
rect 3094 -914 3124 -886
rect 3209 -924 3239 -902
rect 3287 -924 3317 -902
rect 3402 -914 3432 -886
rect 2629 -985 2659 -952
rect 2127 -1046 2157 -1019
rect 2235 -1046 2250 -1012
rect 2306 -1046 2336 -1024
rect 2450 -1046 2480 -1024
rect 2536 -1046 2551 -1012
rect 2629 -1046 2659 -1019
rect 2707 -985 2737 -952
rect 2822 -964 2852 -942
rect 3094 -964 3124 -942
rect 3674 -914 3704 -886
rect 3789 -924 3819 -902
rect 3867 -924 3897 -902
rect 3982 -914 4012 -886
rect 3209 -985 3239 -952
rect 2707 -1046 2737 -1019
rect 2815 -1046 2830 -1012
rect 2886 -1046 2916 -1024
rect 3030 -1046 3060 -1024
rect 3116 -1046 3131 -1012
rect 3209 -1046 3239 -1019
rect 3287 -985 3317 -952
rect 3402 -964 3432 -942
rect 3674 -964 3704 -942
rect 4254 -914 4284 -886
rect 4369 -924 4399 -902
rect 4447 -924 4477 -902
rect 4562 -914 4592 -886
rect 3789 -985 3819 -952
rect 3287 -1046 3317 -1019
rect 3395 -1046 3410 -1012
rect 3466 -1046 3496 -1024
rect 3610 -1046 3640 -1024
rect 3696 -1046 3711 -1012
rect 3789 -1046 3819 -1019
rect 3867 -985 3897 -952
rect 3982 -964 4012 -942
rect 4254 -964 4284 -942
rect 4834 -914 4864 -886
rect 4949 -924 4979 -902
rect 5027 -924 5057 -902
rect 5142 -914 5172 -886
rect 4369 -985 4399 -952
rect 3867 -1046 3897 -1019
rect 3975 -1046 3990 -1012
rect 4046 -1046 4076 -1024
rect 4190 -1046 4220 -1024
rect 4276 -1046 4291 -1012
rect 4369 -1046 4399 -1019
rect 4447 -985 4477 -952
rect 4562 -964 4592 -942
rect 4834 -964 4864 -942
rect 5414 -914 5444 -886
rect 5529 -924 5559 -902
rect 5607 -924 5637 -902
rect 5722 -914 5752 -886
rect 4949 -985 4979 -952
rect 4447 -1046 4477 -1019
rect 4555 -1046 4570 -1012
rect 4626 -1046 4656 -1024
rect 4770 -1046 4800 -1024
rect 4856 -1046 4871 -1012
rect 4949 -1046 4979 -1019
rect 5027 -985 5057 -952
rect 5142 -964 5172 -942
rect 5414 -964 5444 -942
rect 5994 -914 6024 -886
rect 6109 -924 6139 -902
rect 6187 -924 6217 -902
rect 6302 -914 6332 -886
rect 5529 -985 5559 -952
rect 5027 -1046 5057 -1019
rect 5135 -1046 5150 -1012
rect 5206 -1046 5236 -1024
rect 5350 -1046 5380 -1024
rect 5436 -1046 5451 -1012
rect 5529 -1046 5559 -1019
rect 5607 -985 5637 -952
rect 5722 -964 5752 -942
rect 5994 -964 6024 -942
rect 6109 -985 6139 -952
rect 5607 -1046 5637 -1019
rect 5715 -1046 5730 -1012
rect 5786 -1046 5816 -1024
rect 5930 -1046 5960 -1024
rect 6016 -1046 6031 -1012
rect 6109 -1046 6139 -1019
rect 6187 -985 6217 -952
rect 6302 -964 6332 -942
rect 6187 -1046 6217 -1019
rect 6295 -1046 6310 -1012
rect 6366 -1046 6396 -1024
rect -364 -1060 -334 -1046
rect -100 -1060 -70 -1046
rect 216 -1060 246 -1046
rect 480 -1060 510 -1046
rect 796 -1060 826 -1046
rect 1060 -1060 1090 -1046
rect 1376 -1060 1406 -1046
rect 1640 -1060 1670 -1046
rect 1956 -1060 1986 -1046
rect 2220 -1060 2250 -1046
rect 2536 -1060 2566 -1046
rect 2800 -1060 2830 -1046
rect 3116 -1060 3146 -1046
rect 3380 -1060 3410 -1046
rect 3696 -1060 3726 -1046
rect 3960 -1060 3990 -1046
rect 4276 -1060 4306 -1046
rect 4540 -1060 4570 -1046
rect 4856 -1060 4886 -1046
rect 5120 -1060 5150 -1046
rect 5436 -1060 5466 -1046
rect 5700 -1060 5730 -1046
rect 6016 -1060 6046 -1046
rect 6280 -1060 6310 -1046
rect -450 -1110 -420 -1088
rect -364 -1110 -334 -1088
rect -271 -1110 -241 -1088
rect -193 -1110 -163 -1088
rect -100 -1110 -70 -1088
rect -14 -1110 16 -1088
rect 130 -1110 160 -1088
rect 216 -1110 246 -1088
rect 309 -1110 339 -1088
rect 387 -1110 417 -1088
rect 480 -1110 510 -1088
rect 566 -1110 596 -1088
rect 710 -1110 740 -1088
rect 796 -1110 826 -1088
rect 889 -1110 919 -1088
rect 967 -1110 997 -1088
rect 1060 -1110 1090 -1088
rect 1146 -1110 1176 -1088
rect 1290 -1110 1320 -1088
rect 1376 -1110 1406 -1088
rect 1469 -1110 1499 -1088
rect 1547 -1110 1577 -1088
rect 1640 -1110 1670 -1088
rect 1726 -1110 1756 -1088
rect 1870 -1110 1900 -1088
rect 1956 -1110 1986 -1088
rect 2049 -1110 2079 -1088
rect 2127 -1110 2157 -1088
rect 2220 -1110 2250 -1088
rect 2306 -1110 2336 -1088
rect 2450 -1110 2480 -1088
rect 2536 -1110 2566 -1088
rect 2629 -1110 2659 -1088
rect 2707 -1110 2737 -1088
rect 2800 -1110 2830 -1088
rect 2886 -1110 2916 -1088
rect 3030 -1110 3060 -1088
rect 3116 -1110 3146 -1088
rect 3209 -1110 3239 -1088
rect 3287 -1110 3317 -1088
rect 3380 -1110 3410 -1088
rect 3466 -1110 3496 -1088
rect 3610 -1110 3640 -1088
rect 3696 -1110 3726 -1088
rect 3789 -1110 3819 -1088
rect 3867 -1110 3897 -1088
rect 3960 -1110 3990 -1088
rect 4046 -1110 4076 -1088
rect 4190 -1110 4220 -1088
rect 4276 -1110 4306 -1088
rect 4369 -1110 4399 -1088
rect 4447 -1110 4477 -1088
rect 4540 -1110 4570 -1088
rect 4626 -1110 4656 -1088
rect 4770 -1110 4800 -1088
rect 4856 -1110 4886 -1088
rect 4949 -1110 4979 -1088
rect 5027 -1110 5057 -1088
rect 5120 -1110 5150 -1088
rect 5206 -1110 5236 -1088
rect 5350 -1110 5380 -1088
rect 5436 -1110 5466 -1088
rect 5529 -1110 5559 -1088
rect 5607 -1110 5637 -1088
rect 5700 -1110 5730 -1088
rect 5786 -1110 5816 -1088
rect 5930 -1110 5960 -1088
rect 6016 -1110 6046 -1088
rect 6109 -1110 6139 -1088
rect 6187 -1110 6217 -1088
rect 6280 -1110 6310 -1088
rect 6366 -1110 6396 -1088
rect -541 -1156 6439 -1126
rect -386 -1184 -356 -1156
rect -271 -1194 -241 -1172
rect -193 -1194 -163 -1172
rect -78 -1184 -48 -1156
rect -386 -1234 -356 -1212
rect 194 -1184 224 -1156
rect 309 -1194 339 -1172
rect 387 -1194 417 -1172
rect 502 -1184 532 -1156
rect -271 -1255 -241 -1222
rect -450 -1316 -420 -1294
rect -364 -1316 -349 -1282
rect -271 -1316 -241 -1289
rect -193 -1255 -163 -1222
rect -78 -1234 -48 -1212
rect 194 -1234 224 -1212
rect 774 -1184 804 -1156
rect 889 -1194 919 -1172
rect 967 -1194 997 -1172
rect 1082 -1184 1112 -1156
rect 309 -1255 339 -1222
rect -193 -1316 -163 -1289
rect -85 -1316 -70 -1282
rect -14 -1316 16 -1294
rect 130 -1316 160 -1294
rect 216 -1316 231 -1282
rect 309 -1316 339 -1289
rect 387 -1255 417 -1222
rect 502 -1234 532 -1212
rect 774 -1234 804 -1212
rect 1354 -1184 1384 -1156
rect 1469 -1194 1499 -1172
rect 1547 -1194 1577 -1172
rect 1662 -1184 1692 -1156
rect 889 -1255 919 -1222
rect 387 -1316 417 -1289
rect 495 -1316 510 -1282
rect 566 -1316 596 -1294
rect 710 -1316 740 -1294
rect 796 -1316 811 -1282
rect 889 -1316 919 -1289
rect 967 -1255 997 -1222
rect 1082 -1234 1112 -1212
rect 1354 -1234 1384 -1212
rect 1934 -1184 1964 -1156
rect 2049 -1194 2079 -1172
rect 2127 -1194 2157 -1172
rect 2242 -1184 2272 -1156
rect 1469 -1255 1499 -1222
rect 967 -1316 997 -1289
rect 1075 -1316 1090 -1282
rect 1146 -1316 1176 -1294
rect 1290 -1316 1320 -1294
rect 1376 -1316 1391 -1282
rect 1469 -1316 1499 -1289
rect 1547 -1255 1577 -1222
rect 1662 -1234 1692 -1212
rect 1934 -1234 1964 -1212
rect 2514 -1184 2544 -1156
rect 2629 -1194 2659 -1172
rect 2707 -1194 2737 -1172
rect 2822 -1184 2852 -1156
rect 2049 -1255 2079 -1222
rect 1547 -1316 1577 -1289
rect 1655 -1316 1670 -1282
rect 1726 -1316 1756 -1294
rect 1870 -1316 1900 -1294
rect 1956 -1316 1971 -1282
rect 2049 -1316 2079 -1289
rect 2127 -1255 2157 -1222
rect 2242 -1234 2272 -1212
rect 2514 -1234 2544 -1212
rect 3094 -1184 3124 -1156
rect 3209 -1194 3239 -1172
rect 3287 -1194 3317 -1172
rect 3402 -1184 3432 -1156
rect 2629 -1255 2659 -1222
rect 2127 -1316 2157 -1289
rect 2235 -1316 2250 -1282
rect 2306 -1316 2336 -1294
rect 2450 -1316 2480 -1294
rect 2536 -1316 2551 -1282
rect 2629 -1316 2659 -1289
rect 2707 -1255 2737 -1222
rect 2822 -1234 2852 -1212
rect 3094 -1234 3124 -1212
rect 3674 -1184 3704 -1156
rect 3789 -1194 3819 -1172
rect 3867 -1194 3897 -1172
rect 3982 -1184 4012 -1156
rect 3209 -1255 3239 -1222
rect 2707 -1316 2737 -1289
rect 2815 -1316 2830 -1282
rect 2886 -1316 2916 -1294
rect 3030 -1316 3060 -1294
rect 3116 -1316 3131 -1282
rect 3209 -1316 3239 -1289
rect 3287 -1255 3317 -1222
rect 3402 -1234 3432 -1212
rect 3674 -1234 3704 -1212
rect 4254 -1184 4284 -1156
rect 4369 -1194 4399 -1172
rect 4447 -1194 4477 -1172
rect 4562 -1184 4592 -1156
rect 3789 -1255 3819 -1222
rect 3287 -1316 3317 -1289
rect 3395 -1316 3410 -1282
rect 3466 -1316 3496 -1294
rect 3610 -1316 3640 -1294
rect 3696 -1316 3711 -1282
rect 3789 -1316 3819 -1289
rect 3867 -1255 3897 -1222
rect 3982 -1234 4012 -1212
rect 4254 -1234 4284 -1212
rect 4834 -1184 4864 -1156
rect 4949 -1194 4979 -1172
rect 5027 -1194 5057 -1172
rect 5142 -1184 5172 -1156
rect 4369 -1255 4399 -1222
rect 3867 -1316 3897 -1289
rect 3975 -1316 3990 -1282
rect 4046 -1316 4076 -1294
rect 4190 -1316 4220 -1294
rect 4276 -1316 4291 -1282
rect 4369 -1316 4399 -1289
rect 4447 -1255 4477 -1222
rect 4562 -1234 4592 -1212
rect 4834 -1234 4864 -1212
rect 5414 -1184 5444 -1156
rect 5529 -1194 5559 -1172
rect 5607 -1194 5637 -1172
rect 5722 -1184 5752 -1156
rect 4949 -1255 4979 -1222
rect 4447 -1316 4477 -1289
rect 4555 -1316 4570 -1282
rect 4626 -1316 4656 -1294
rect 4770 -1316 4800 -1294
rect 4856 -1316 4871 -1282
rect 4949 -1316 4979 -1289
rect 5027 -1255 5057 -1222
rect 5142 -1234 5172 -1212
rect 5414 -1234 5444 -1212
rect 5994 -1184 6024 -1156
rect 6109 -1194 6139 -1172
rect 6187 -1194 6217 -1172
rect 6302 -1184 6332 -1156
rect 5529 -1255 5559 -1222
rect 5027 -1316 5057 -1289
rect 5135 -1316 5150 -1282
rect 5206 -1316 5236 -1294
rect 5350 -1316 5380 -1294
rect 5436 -1316 5451 -1282
rect 5529 -1316 5559 -1289
rect 5607 -1255 5637 -1222
rect 5722 -1234 5752 -1212
rect 5994 -1234 6024 -1212
rect 6109 -1255 6139 -1222
rect 5607 -1316 5637 -1289
rect 5715 -1316 5730 -1282
rect 5786 -1316 5816 -1294
rect 5930 -1316 5960 -1294
rect 6016 -1316 6031 -1282
rect 6109 -1316 6139 -1289
rect 6187 -1255 6217 -1222
rect 6302 -1234 6332 -1212
rect 6187 -1316 6217 -1289
rect 6295 -1316 6310 -1282
rect 6366 -1316 6396 -1294
rect -364 -1330 -334 -1316
rect -100 -1330 -70 -1316
rect 216 -1330 246 -1316
rect 480 -1330 510 -1316
rect 796 -1330 826 -1316
rect 1060 -1330 1090 -1316
rect 1376 -1330 1406 -1316
rect 1640 -1330 1670 -1316
rect 1956 -1330 1986 -1316
rect 2220 -1330 2250 -1316
rect 2536 -1330 2566 -1316
rect 2800 -1330 2830 -1316
rect 3116 -1330 3146 -1316
rect 3380 -1330 3410 -1316
rect 3696 -1330 3726 -1316
rect 3960 -1330 3990 -1316
rect 4276 -1330 4306 -1316
rect 4540 -1330 4570 -1316
rect 4856 -1330 4886 -1316
rect 5120 -1330 5150 -1316
rect 5436 -1330 5466 -1316
rect 5700 -1330 5730 -1316
rect 6016 -1330 6046 -1316
rect 6280 -1330 6310 -1316
rect -450 -1380 -420 -1358
rect -364 -1380 -334 -1358
rect -271 -1380 -241 -1358
rect -193 -1380 -163 -1358
rect -100 -1380 -70 -1358
rect -14 -1380 16 -1358
rect 130 -1380 160 -1358
rect 216 -1380 246 -1358
rect 309 -1380 339 -1358
rect 387 -1380 417 -1358
rect 480 -1380 510 -1358
rect 566 -1380 596 -1358
rect 710 -1380 740 -1358
rect 796 -1380 826 -1358
rect 889 -1380 919 -1358
rect 967 -1380 997 -1358
rect 1060 -1380 1090 -1358
rect 1146 -1380 1176 -1358
rect 1290 -1380 1320 -1358
rect 1376 -1380 1406 -1358
rect 1469 -1380 1499 -1358
rect 1547 -1380 1577 -1358
rect 1640 -1380 1670 -1358
rect 1726 -1380 1756 -1358
rect 1870 -1380 1900 -1358
rect 1956 -1380 1986 -1358
rect 2049 -1380 2079 -1358
rect 2127 -1380 2157 -1358
rect 2220 -1380 2250 -1358
rect 2306 -1380 2336 -1358
rect 2450 -1380 2480 -1358
rect 2536 -1380 2566 -1358
rect 2629 -1380 2659 -1358
rect 2707 -1380 2737 -1358
rect 2800 -1380 2830 -1358
rect 2886 -1380 2916 -1358
rect 3030 -1380 3060 -1358
rect 3116 -1380 3146 -1358
rect 3209 -1380 3239 -1358
rect 3287 -1380 3317 -1358
rect 3380 -1380 3410 -1358
rect 3466 -1380 3496 -1358
rect 3610 -1380 3640 -1358
rect 3696 -1380 3726 -1358
rect 3789 -1380 3819 -1358
rect 3867 -1380 3897 -1358
rect 3960 -1380 3990 -1358
rect 4046 -1380 4076 -1358
rect 4190 -1380 4220 -1358
rect 4276 -1380 4306 -1358
rect 4369 -1380 4399 -1358
rect 4447 -1380 4477 -1358
rect 4540 -1380 4570 -1358
rect 4626 -1380 4656 -1358
rect 4770 -1380 4800 -1358
rect 4856 -1380 4886 -1358
rect 4949 -1380 4979 -1358
rect 5027 -1380 5057 -1358
rect 5120 -1380 5150 -1358
rect 5206 -1380 5236 -1358
rect 5350 -1380 5380 -1358
rect 5436 -1380 5466 -1358
rect 5529 -1380 5559 -1358
rect 5607 -1380 5637 -1358
rect 5700 -1380 5730 -1358
rect 5786 -1380 5816 -1358
rect 5930 -1380 5960 -1358
rect 6016 -1380 6046 -1358
rect 6109 -1380 6139 -1358
rect 6187 -1380 6217 -1358
rect 6280 -1380 6310 -1358
rect 6366 -1380 6396 -1358
rect -541 -1426 6439 -1396
rect -386 -1454 -356 -1426
rect -271 -1464 -241 -1442
rect -193 -1464 -163 -1442
rect -78 -1454 -48 -1426
rect -386 -1504 -356 -1482
rect 194 -1454 224 -1426
rect 309 -1464 339 -1442
rect 387 -1464 417 -1442
rect 502 -1454 532 -1426
rect -271 -1525 -241 -1492
rect -450 -1586 -420 -1564
rect -364 -1586 -349 -1552
rect -271 -1586 -241 -1559
rect -193 -1525 -163 -1492
rect -78 -1504 -48 -1482
rect 194 -1504 224 -1482
rect 774 -1454 804 -1426
rect 889 -1464 919 -1442
rect 967 -1464 997 -1442
rect 1082 -1454 1112 -1426
rect 309 -1525 339 -1492
rect -193 -1586 -163 -1559
rect -85 -1586 -70 -1552
rect -14 -1586 16 -1564
rect 130 -1586 160 -1564
rect 216 -1586 231 -1552
rect 309 -1586 339 -1559
rect 387 -1525 417 -1492
rect 502 -1504 532 -1482
rect 774 -1504 804 -1482
rect 1354 -1454 1384 -1426
rect 1469 -1464 1499 -1442
rect 1547 -1464 1577 -1442
rect 1662 -1454 1692 -1426
rect 889 -1525 919 -1492
rect 387 -1586 417 -1559
rect 495 -1586 510 -1552
rect 566 -1586 596 -1564
rect 710 -1586 740 -1564
rect 796 -1586 811 -1552
rect 889 -1586 919 -1559
rect 967 -1525 997 -1492
rect 1082 -1504 1112 -1482
rect 1354 -1504 1384 -1482
rect 1934 -1454 1964 -1426
rect 2049 -1464 2079 -1442
rect 2127 -1464 2157 -1442
rect 2242 -1454 2272 -1426
rect 1469 -1525 1499 -1492
rect 967 -1586 997 -1559
rect 1075 -1586 1090 -1552
rect 1146 -1586 1176 -1564
rect 1290 -1586 1320 -1564
rect 1376 -1586 1391 -1552
rect 1469 -1586 1499 -1559
rect 1547 -1525 1577 -1492
rect 1662 -1504 1692 -1482
rect 1934 -1504 1964 -1482
rect 2514 -1454 2544 -1426
rect 2629 -1464 2659 -1442
rect 2707 -1464 2737 -1442
rect 2822 -1454 2852 -1426
rect 2049 -1525 2079 -1492
rect 1547 -1586 1577 -1559
rect 1655 -1586 1670 -1552
rect 1726 -1586 1756 -1564
rect 1870 -1586 1900 -1564
rect 1956 -1586 1971 -1552
rect 2049 -1586 2079 -1559
rect 2127 -1525 2157 -1492
rect 2242 -1504 2272 -1482
rect 2514 -1504 2544 -1482
rect 3094 -1454 3124 -1426
rect 3209 -1464 3239 -1442
rect 3287 -1464 3317 -1442
rect 3402 -1454 3432 -1426
rect 2629 -1525 2659 -1492
rect 2127 -1586 2157 -1559
rect 2235 -1586 2250 -1552
rect 2306 -1586 2336 -1564
rect 2450 -1586 2480 -1564
rect 2536 -1586 2551 -1552
rect 2629 -1586 2659 -1559
rect 2707 -1525 2737 -1492
rect 2822 -1504 2852 -1482
rect 3094 -1504 3124 -1482
rect 3674 -1454 3704 -1426
rect 3789 -1464 3819 -1442
rect 3867 -1464 3897 -1442
rect 3982 -1454 4012 -1426
rect 3209 -1525 3239 -1492
rect 2707 -1586 2737 -1559
rect 2815 -1586 2830 -1552
rect 2886 -1586 2916 -1564
rect 3030 -1586 3060 -1564
rect 3116 -1586 3131 -1552
rect 3209 -1586 3239 -1559
rect 3287 -1525 3317 -1492
rect 3402 -1504 3432 -1482
rect 3674 -1504 3704 -1482
rect 4254 -1454 4284 -1426
rect 4369 -1464 4399 -1442
rect 4447 -1464 4477 -1442
rect 4562 -1454 4592 -1426
rect 3789 -1525 3819 -1492
rect 3287 -1586 3317 -1559
rect 3395 -1586 3410 -1552
rect 3466 -1586 3496 -1564
rect 3610 -1586 3640 -1564
rect 3696 -1586 3711 -1552
rect 3789 -1586 3819 -1559
rect 3867 -1525 3897 -1492
rect 3982 -1504 4012 -1482
rect 4254 -1504 4284 -1482
rect 4834 -1454 4864 -1426
rect 4949 -1464 4979 -1442
rect 5027 -1464 5057 -1442
rect 5142 -1454 5172 -1426
rect 4369 -1525 4399 -1492
rect 3867 -1586 3897 -1559
rect 3975 -1586 3990 -1552
rect 4046 -1586 4076 -1564
rect 4190 -1586 4220 -1564
rect 4276 -1586 4291 -1552
rect 4369 -1586 4399 -1559
rect 4447 -1525 4477 -1492
rect 4562 -1504 4592 -1482
rect 4834 -1504 4864 -1482
rect 5414 -1454 5444 -1426
rect 5529 -1464 5559 -1442
rect 5607 -1464 5637 -1442
rect 5722 -1454 5752 -1426
rect 4949 -1525 4979 -1492
rect 4447 -1586 4477 -1559
rect 4555 -1586 4570 -1552
rect 4626 -1586 4656 -1564
rect 4770 -1586 4800 -1564
rect 4856 -1586 4871 -1552
rect 4949 -1586 4979 -1559
rect 5027 -1525 5057 -1492
rect 5142 -1504 5172 -1482
rect 5414 -1504 5444 -1482
rect 5994 -1454 6024 -1426
rect 6109 -1464 6139 -1442
rect 6187 -1464 6217 -1442
rect 6302 -1454 6332 -1426
rect 5529 -1525 5559 -1492
rect 5027 -1586 5057 -1559
rect 5135 -1586 5150 -1552
rect 5206 -1586 5236 -1564
rect 5350 -1586 5380 -1564
rect 5436 -1586 5451 -1552
rect 5529 -1586 5559 -1559
rect 5607 -1525 5637 -1492
rect 5722 -1504 5752 -1482
rect 5994 -1504 6024 -1482
rect 6109 -1525 6139 -1492
rect 5607 -1586 5637 -1559
rect 5715 -1586 5730 -1552
rect 5786 -1586 5816 -1564
rect 5930 -1586 5960 -1564
rect 6016 -1586 6031 -1552
rect 6109 -1586 6139 -1559
rect 6187 -1525 6217 -1492
rect 6302 -1504 6332 -1482
rect 6187 -1586 6217 -1559
rect 6295 -1586 6310 -1552
rect 6366 -1586 6396 -1564
rect -364 -1600 -334 -1586
rect -100 -1600 -70 -1586
rect 216 -1600 246 -1586
rect 480 -1600 510 -1586
rect 796 -1600 826 -1586
rect 1060 -1600 1090 -1586
rect 1376 -1600 1406 -1586
rect 1640 -1600 1670 -1586
rect 1956 -1600 1986 -1586
rect 2220 -1600 2250 -1586
rect 2536 -1600 2566 -1586
rect 2800 -1600 2830 -1586
rect 3116 -1600 3146 -1586
rect 3380 -1600 3410 -1586
rect 3696 -1600 3726 -1586
rect 3960 -1600 3990 -1586
rect 4276 -1600 4306 -1586
rect 4540 -1600 4570 -1586
rect 4856 -1600 4886 -1586
rect 5120 -1600 5150 -1586
rect 5436 -1600 5466 -1586
rect 5700 -1600 5730 -1586
rect 6016 -1600 6046 -1586
rect 6280 -1600 6310 -1586
rect -450 -1650 -420 -1628
rect -364 -1650 -334 -1628
rect -271 -1650 -241 -1628
rect -193 -1650 -163 -1628
rect -100 -1650 -70 -1628
rect -14 -1650 16 -1628
rect 130 -1650 160 -1628
rect 216 -1650 246 -1628
rect 309 -1650 339 -1628
rect 387 -1650 417 -1628
rect 480 -1650 510 -1628
rect 566 -1650 596 -1628
rect 710 -1650 740 -1628
rect 796 -1650 826 -1628
rect 889 -1650 919 -1628
rect 967 -1650 997 -1628
rect 1060 -1650 1090 -1628
rect 1146 -1650 1176 -1628
rect 1290 -1650 1320 -1628
rect 1376 -1650 1406 -1628
rect 1469 -1650 1499 -1628
rect 1547 -1650 1577 -1628
rect 1640 -1650 1670 -1628
rect 1726 -1650 1756 -1628
rect 1870 -1650 1900 -1628
rect 1956 -1650 1986 -1628
rect 2049 -1650 2079 -1628
rect 2127 -1650 2157 -1628
rect 2220 -1650 2250 -1628
rect 2306 -1650 2336 -1628
rect 2450 -1650 2480 -1628
rect 2536 -1650 2566 -1628
rect 2629 -1650 2659 -1628
rect 2707 -1650 2737 -1628
rect 2800 -1650 2830 -1628
rect 2886 -1650 2916 -1628
rect 3030 -1650 3060 -1628
rect 3116 -1650 3146 -1628
rect 3209 -1650 3239 -1628
rect 3287 -1650 3317 -1628
rect 3380 -1650 3410 -1628
rect 3466 -1650 3496 -1628
rect 3610 -1650 3640 -1628
rect 3696 -1650 3726 -1628
rect 3789 -1650 3819 -1628
rect 3867 -1650 3897 -1628
rect 3960 -1650 3990 -1628
rect 4046 -1650 4076 -1628
rect 4190 -1650 4220 -1628
rect 4276 -1650 4306 -1628
rect 4369 -1650 4399 -1628
rect 4447 -1650 4477 -1628
rect 4540 -1650 4570 -1628
rect 4626 -1650 4656 -1628
rect 4770 -1650 4800 -1628
rect 4856 -1650 4886 -1628
rect 4949 -1650 4979 -1628
rect 5027 -1650 5057 -1628
rect 5120 -1650 5150 -1628
rect 5206 -1650 5236 -1628
rect 5350 -1650 5380 -1628
rect 5436 -1650 5466 -1628
rect 5529 -1650 5559 -1628
rect 5607 -1650 5637 -1628
rect 5700 -1650 5730 -1628
rect 5786 -1650 5816 -1628
rect 5930 -1650 5960 -1628
rect 6016 -1650 6046 -1628
rect 6109 -1650 6139 -1628
rect 6187 -1650 6217 -1628
rect 6280 -1650 6310 -1628
rect 6366 -1650 6396 -1628
rect -541 -1696 6439 -1666
rect -386 -1724 -356 -1696
rect -271 -1734 -241 -1712
rect -193 -1734 -163 -1712
rect -78 -1724 -48 -1696
rect -386 -1774 -356 -1752
rect 194 -1724 224 -1696
rect 309 -1734 339 -1712
rect 387 -1734 417 -1712
rect 502 -1724 532 -1696
rect -271 -1795 -241 -1762
rect -450 -1856 -420 -1834
rect -364 -1856 -349 -1822
rect -271 -1856 -241 -1829
rect -193 -1795 -163 -1762
rect -78 -1774 -48 -1752
rect 194 -1774 224 -1752
rect 774 -1724 804 -1696
rect 889 -1734 919 -1712
rect 967 -1734 997 -1712
rect 1082 -1724 1112 -1696
rect 309 -1795 339 -1762
rect -193 -1856 -163 -1829
rect -85 -1856 -70 -1822
rect -14 -1856 16 -1834
rect 130 -1856 160 -1834
rect 216 -1856 231 -1822
rect 309 -1856 339 -1829
rect 387 -1795 417 -1762
rect 502 -1774 532 -1752
rect 774 -1774 804 -1752
rect 1354 -1724 1384 -1696
rect 1469 -1734 1499 -1712
rect 1547 -1734 1577 -1712
rect 1662 -1724 1692 -1696
rect 889 -1795 919 -1762
rect 387 -1856 417 -1829
rect 495 -1856 510 -1822
rect 566 -1856 596 -1834
rect 710 -1856 740 -1834
rect 796 -1856 811 -1822
rect 889 -1856 919 -1829
rect 967 -1795 997 -1762
rect 1082 -1774 1112 -1752
rect 1354 -1774 1384 -1752
rect 1934 -1724 1964 -1696
rect 2049 -1734 2079 -1712
rect 2127 -1734 2157 -1712
rect 2242 -1724 2272 -1696
rect 1469 -1795 1499 -1762
rect 967 -1856 997 -1829
rect 1075 -1856 1090 -1822
rect 1146 -1856 1176 -1834
rect 1290 -1856 1320 -1834
rect 1376 -1856 1391 -1822
rect 1469 -1856 1499 -1829
rect 1547 -1795 1577 -1762
rect 1662 -1774 1692 -1752
rect 1934 -1774 1964 -1752
rect 2514 -1724 2544 -1696
rect 2629 -1734 2659 -1712
rect 2707 -1734 2737 -1712
rect 2822 -1724 2852 -1696
rect 2049 -1795 2079 -1762
rect 1547 -1856 1577 -1829
rect 1655 -1856 1670 -1822
rect 1726 -1856 1756 -1834
rect 1870 -1856 1900 -1834
rect 1956 -1856 1971 -1822
rect 2049 -1856 2079 -1829
rect 2127 -1795 2157 -1762
rect 2242 -1774 2272 -1752
rect 2514 -1774 2544 -1752
rect 3094 -1724 3124 -1696
rect 3209 -1734 3239 -1712
rect 3287 -1734 3317 -1712
rect 3402 -1724 3432 -1696
rect 2629 -1795 2659 -1762
rect 2127 -1856 2157 -1829
rect 2235 -1856 2250 -1822
rect 2306 -1856 2336 -1834
rect 2450 -1856 2480 -1834
rect 2536 -1856 2551 -1822
rect 2629 -1856 2659 -1829
rect 2707 -1795 2737 -1762
rect 2822 -1774 2852 -1752
rect 3094 -1774 3124 -1752
rect 3674 -1724 3704 -1696
rect 3789 -1734 3819 -1712
rect 3867 -1734 3897 -1712
rect 3982 -1724 4012 -1696
rect 3209 -1795 3239 -1762
rect 2707 -1856 2737 -1829
rect 2815 -1856 2830 -1822
rect 2886 -1856 2916 -1834
rect 3030 -1856 3060 -1834
rect 3116 -1856 3131 -1822
rect 3209 -1856 3239 -1829
rect 3287 -1795 3317 -1762
rect 3402 -1774 3432 -1752
rect 3674 -1774 3704 -1752
rect 4254 -1724 4284 -1696
rect 4369 -1734 4399 -1712
rect 4447 -1734 4477 -1712
rect 4562 -1724 4592 -1696
rect 3789 -1795 3819 -1762
rect 3287 -1856 3317 -1829
rect 3395 -1856 3410 -1822
rect 3466 -1856 3496 -1834
rect 3610 -1856 3640 -1834
rect 3696 -1856 3711 -1822
rect 3789 -1856 3819 -1829
rect 3867 -1795 3897 -1762
rect 3982 -1774 4012 -1752
rect 4254 -1774 4284 -1752
rect 4834 -1724 4864 -1696
rect 4949 -1734 4979 -1712
rect 5027 -1734 5057 -1712
rect 5142 -1724 5172 -1696
rect 4369 -1795 4399 -1762
rect 3867 -1856 3897 -1829
rect 3975 -1856 3990 -1822
rect 4046 -1856 4076 -1834
rect 4190 -1856 4220 -1834
rect 4276 -1856 4291 -1822
rect 4369 -1856 4399 -1829
rect 4447 -1795 4477 -1762
rect 4562 -1774 4592 -1752
rect 4834 -1774 4864 -1752
rect 5414 -1724 5444 -1696
rect 5529 -1734 5559 -1712
rect 5607 -1734 5637 -1712
rect 5722 -1724 5752 -1696
rect 4949 -1795 4979 -1762
rect 4447 -1856 4477 -1829
rect 4555 -1856 4570 -1822
rect 4626 -1856 4656 -1834
rect 4770 -1856 4800 -1834
rect 4856 -1856 4871 -1822
rect 4949 -1856 4979 -1829
rect 5027 -1795 5057 -1762
rect 5142 -1774 5172 -1752
rect 5414 -1774 5444 -1752
rect 5994 -1724 6024 -1696
rect 6109 -1734 6139 -1712
rect 6187 -1734 6217 -1712
rect 6302 -1724 6332 -1696
rect 5529 -1795 5559 -1762
rect 5027 -1856 5057 -1829
rect 5135 -1856 5150 -1822
rect 5206 -1856 5236 -1834
rect 5350 -1856 5380 -1834
rect 5436 -1856 5451 -1822
rect 5529 -1856 5559 -1829
rect 5607 -1795 5637 -1762
rect 5722 -1774 5752 -1752
rect 5994 -1774 6024 -1752
rect 6109 -1795 6139 -1762
rect 5607 -1856 5637 -1829
rect 5715 -1856 5730 -1822
rect 5786 -1856 5816 -1834
rect 5930 -1856 5960 -1834
rect 6016 -1856 6031 -1822
rect 6109 -1856 6139 -1829
rect 6187 -1795 6217 -1762
rect 6302 -1774 6332 -1752
rect 6187 -1856 6217 -1829
rect 6295 -1856 6310 -1822
rect 6366 -1856 6396 -1834
rect -364 -1870 -334 -1856
rect -100 -1870 -70 -1856
rect 216 -1870 246 -1856
rect 480 -1870 510 -1856
rect 796 -1870 826 -1856
rect 1060 -1870 1090 -1856
rect 1376 -1870 1406 -1856
rect 1640 -1870 1670 -1856
rect 1956 -1870 1986 -1856
rect 2220 -1870 2250 -1856
rect 2536 -1870 2566 -1856
rect 2800 -1870 2830 -1856
rect 3116 -1870 3146 -1856
rect 3380 -1870 3410 -1856
rect 3696 -1870 3726 -1856
rect 3960 -1870 3990 -1856
rect 4276 -1870 4306 -1856
rect 4540 -1870 4570 -1856
rect 4856 -1870 4886 -1856
rect 5120 -1870 5150 -1856
rect 5436 -1870 5466 -1856
rect 5700 -1870 5730 -1856
rect 6016 -1870 6046 -1856
rect 6280 -1870 6310 -1856
rect -450 -1920 -420 -1898
rect -364 -1920 -334 -1898
rect -271 -1920 -241 -1898
rect -193 -1920 -163 -1898
rect -100 -1920 -70 -1898
rect -14 -1920 16 -1898
rect 130 -1920 160 -1898
rect 216 -1920 246 -1898
rect 309 -1920 339 -1898
rect 387 -1920 417 -1898
rect 480 -1920 510 -1898
rect 566 -1920 596 -1898
rect 710 -1920 740 -1898
rect 796 -1920 826 -1898
rect 889 -1920 919 -1898
rect 967 -1920 997 -1898
rect 1060 -1920 1090 -1898
rect 1146 -1920 1176 -1898
rect 1290 -1920 1320 -1898
rect 1376 -1920 1406 -1898
rect 1469 -1920 1499 -1898
rect 1547 -1920 1577 -1898
rect 1640 -1920 1670 -1898
rect 1726 -1920 1756 -1898
rect 1870 -1920 1900 -1898
rect 1956 -1920 1986 -1898
rect 2049 -1920 2079 -1898
rect 2127 -1920 2157 -1898
rect 2220 -1920 2250 -1898
rect 2306 -1920 2336 -1898
rect 2450 -1920 2480 -1898
rect 2536 -1920 2566 -1898
rect 2629 -1920 2659 -1898
rect 2707 -1920 2737 -1898
rect 2800 -1920 2830 -1898
rect 2886 -1920 2916 -1898
rect 3030 -1920 3060 -1898
rect 3116 -1920 3146 -1898
rect 3209 -1920 3239 -1898
rect 3287 -1920 3317 -1898
rect 3380 -1920 3410 -1898
rect 3466 -1920 3496 -1898
rect 3610 -1920 3640 -1898
rect 3696 -1920 3726 -1898
rect 3789 -1920 3819 -1898
rect 3867 -1920 3897 -1898
rect 3960 -1920 3990 -1898
rect 4046 -1920 4076 -1898
rect 4190 -1920 4220 -1898
rect 4276 -1920 4306 -1898
rect 4369 -1920 4399 -1898
rect 4447 -1920 4477 -1898
rect 4540 -1920 4570 -1898
rect 4626 -1920 4656 -1898
rect 4770 -1920 4800 -1898
rect 4856 -1920 4886 -1898
rect 4949 -1920 4979 -1898
rect 5027 -1920 5057 -1898
rect 5120 -1920 5150 -1898
rect 5206 -1920 5236 -1898
rect 5350 -1920 5380 -1898
rect 5436 -1920 5466 -1898
rect 5529 -1920 5559 -1898
rect 5607 -1920 5637 -1898
rect 5700 -1920 5730 -1898
rect 5786 -1920 5816 -1898
rect 5930 -1920 5960 -1898
rect 6016 -1920 6046 -1898
rect 6109 -1920 6139 -1898
rect 6187 -1920 6217 -1898
rect 6280 -1920 6310 -1898
rect 6366 -1920 6396 -1898
rect -541 -1966 6439 -1936
rect -386 -1994 -356 -1966
rect -271 -2004 -241 -1982
rect -193 -2004 -163 -1982
rect -78 -1994 -48 -1966
rect -386 -2044 -356 -2022
rect 194 -1994 224 -1966
rect 309 -2004 339 -1982
rect 387 -2004 417 -1982
rect 502 -1994 532 -1966
rect -271 -2065 -241 -2032
rect -450 -2126 -420 -2104
rect -364 -2126 -349 -2092
rect -271 -2126 -241 -2099
rect -193 -2065 -163 -2032
rect -78 -2044 -48 -2022
rect 194 -2044 224 -2022
rect 774 -1994 804 -1966
rect 889 -2004 919 -1982
rect 967 -2004 997 -1982
rect 1082 -1994 1112 -1966
rect 309 -2065 339 -2032
rect -193 -2126 -163 -2099
rect -85 -2126 -70 -2092
rect -14 -2126 16 -2104
rect 130 -2126 160 -2104
rect 216 -2126 231 -2092
rect 309 -2126 339 -2099
rect 387 -2065 417 -2032
rect 502 -2044 532 -2022
rect 774 -2044 804 -2022
rect 1354 -1994 1384 -1966
rect 1469 -2004 1499 -1982
rect 1547 -2004 1577 -1982
rect 1662 -1994 1692 -1966
rect 889 -2065 919 -2032
rect 387 -2126 417 -2099
rect 495 -2126 510 -2092
rect 566 -2126 596 -2104
rect 710 -2126 740 -2104
rect 796 -2126 811 -2092
rect 889 -2126 919 -2099
rect 967 -2065 997 -2032
rect 1082 -2044 1112 -2022
rect 1354 -2044 1384 -2022
rect 1934 -1994 1964 -1966
rect 2049 -2004 2079 -1982
rect 2127 -2004 2157 -1982
rect 2242 -1994 2272 -1966
rect 1469 -2065 1499 -2032
rect 967 -2126 997 -2099
rect 1075 -2126 1090 -2092
rect 1146 -2126 1176 -2104
rect 1290 -2126 1320 -2104
rect 1376 -2126 1391 -2092
rect 1469 -2126 1499 -2099
rect 1547 -2065 1577 -2032
rect 1662 -2044 1692 -2022
rect 1934 -2044 1964 -2022
rect 2514 -1994 2544 -1966
rect 2629 -2004 2659 -1982
rect 2707 -2004 2737 -1982
rect 2822 -1994 2852 -1966
rect 2049 -2065 2079 -2032
rect 1547 -2126 1577 -2099
rect 1655 -2126 1670 -2092
rect 1726 -2126 1756 -2104
rect 1870 -2126 1900 -2104
rect 1956 -2126 1971 -2092
rect 2049 -2126 2079 -2099
rect 2127 -2065 2157 -2032
rect 2242 -2044 2272 -2022
rect 2514 -2044 2544 -2022
rect 3094 -1994 3124 -1966
rect 3209 -2004 3239 -1982
rect 3287 -2004 3317 -1982
rect 3402 -1994 3432 -1966
rect 2629 -2065 2659 -2032
rect 2127 -2126 2157 -2099
rect 2235 -2126 2250 -2092
rect 2306 -2126 2336 -2104
rect 2450 -2126 2480 -2104
rect 2536 -2126 2551 -2092
rect 2629 -2126 2659 -2099
rect 2707 -2065 2737 -2032
rect 2822 -2044 2852 -2022
rect 3094 -2044 3124 -2022
rect 3674 -1994 3704 -1966
rect 3789 -2004 3819 -1982
rect 3867 -2004 3897 -1982
rect 3982 -1994 4012 -1966
rect 3209 -2065 3239 -2032
rect 2707 -2126 2737 -2099
rect 2815 -2126 2830 -2092
rect 2886 -2126 2916 -2104
rect 3030 -2126 3060 -2104
rect 3116 -2126 3131 -2092
rect 3209 -2126 3239 -2099
rect 3287 -2065 3317 -2032
rect 3402 -2044 3432 -2022
rect 3674 -2044 3704 -2022
rect 4254 -1994 4284 -1966
rect 4369 -2004 4399 -1982
rect 4447 -2004 4477 -1982
rect 4562 -1994 4592 -1966
rect 3789 -2065 3819 -2032
rect 3287 -2126 3317 -2099
rect 3395 -2126 3410 -2092
rect 3466 -2126 3496 -2104
rect 3610 -2126 3640 -2104
rect 3696 -2126 3711 -2092
rect 3789 -2126 3819 -2099
rect 3867 -2065 3897 -2032
rect 3982 -2044 4012 -2022
rect 4254 -2044 4284 -2022
rect 4834 -1994 4864 -1966
rect 4949 -2004 4979 -1982
rect 5027 -2004 5057 -1982
rect 5142 -1994 5172 -1966
rect 4369 -2065 4399 -2032
rect 3867 -2126 3897 -2099
rect 3975 -2126 3990 -2092
rect 4046 -2126 4076 -2104
rect 4190 -2126 4220 -2104
rect 4276 -2126 4291 -2092
rect 4369 -2126 4399 -2099
rect 4447 -2065 4477 -2032
rect 4562 -2044 4592 -2022
rect 4834 -2044 4864 -2022
rect 5414 -1994 5444 -1966
rect 5529 -2004 5559 -1982
rect 5607 -2004 5637 -1982
rect 5722 -1994 5752 -1966
rect 4949 -2065 4979 -2032
rect 4447 -2126 4477 -2099
rect 4555 -2126 4570 -2092
rect 4626 -2126 4656 -2104
rect 4770 -2126 4800 -2104
rect 4856 -2126 4871 -2092
rect 4949 -2126 4979 -2099
rect 5027 -2065 5057 -2032
rect 5142 -2044 5172 -2022
rect 5414 -2044 5444 -2022
rect 5994 -1994 6024 -1966
rect 6109 -2004 6139 -1982
rect 6187 -2004 6217 -1982
rect 6302 -1994 6332 -1966
rect 5529 -2065 5559 -2032
rect 5027 -2126 5057 -2099
rect 5135 -2126 5150 -2092
rect 5206 -2126 5236 -2104
rect 5350 -2126 5380 -2104
rect 5436 -2126 5451 -2092
rect 5529 -2126 5559 -2099
rect 5607 -2065 5637 -2032
rect 5722 -2044 5752 -2022
rect 5994 -2044 6024 -2022
rect 6109 -2065 6139 -2032
rect 5607 -2126 5637 -2099
rect 5715 -2126 5730 -2092
rect 5786 -2126 5816 -2104
rect 5930 -2126 5960 -2104
rect 6016 -2126 6031 -2092
rect 6109 -2126 6139 -2099
rect 6187 -2065 6217 -2032
rect 6302 -2044 6332 -2022
rect 6187 -2126 6217 -2099
rect 6295 -2126 6310 -2092
rect 6366 -2126 6396 -2104
rect -364 -2140 -334 -2126
rect -100 -2140 -70 -2126
rect 216 -2140 246 -2126
rect 480 -2140 510 -2126
rect 796 -2140 826 -2126
rect 1060 -2140 1090 -2126
rect 1376 -2140 1406 -2126
rect 1640 -2140 1670 -2126
rect 1956 -2140 1986 -2126
rect 2220 -2140 2250 -2126
rect 2536 -2140 2566 -2126
rect 2800 -2140 2830 -2126
rect 3116 -2140 3146 -2126
rect 3380 -2140 3410 -2126
rect 3696 -2140 3726 -2126
rect 3960 -2140 3990 -2126
rect 4276 -2140 4306 -2126
rect 4540 -2140 4570 -2126
rect 4856 -2140 4886 -2126
rect 5120 -2140 5150 -2126
rect 5436 -2140 5466 -2126
rect 5700 -2140 5730 -2126
rect 6016 -2140 6046 -2126
rect 6280 -2140 6310 -2126
rect -450 -2190 -420 -2168
rect -364 -2190 -334 -2168
rect -271 -2190 -241 -2168
rect -193 -2190 -163 -2168
rect -100 -2190 -70 -2168
rect -14 -2190 16 -2168
rect 130 -2190 160 -2168
rect 216 -2190 246 -2168
rect 309 -2190 339 -2168
rect 387 -2190 417 -2168
rect 480 -2190 510 -2168
rect 566 -2190 596 -2168
rect 710 -2190 740 -2168
rect 796 -2190 826 -2168
rect 889 -2190 919 -2168
rect 967 -2190 997 -2168
rect 1060 -2190 1090 -2168
rect 1146 -2190 1176 -2168
rect 1290 -2190 1320 -2168
rect 1376 -2190 1406 -2168
rect 1469 -2190 1499 -2168
rect 1547 -2190 1577 -2168
rect 1640 -2190 1670 -2168
rect 1726 -2190 1756 -2168
rect 1870 -2190 1900 -2168
rect 1956 -2190 1986 -2168
rect 2049 -2190 2079 -2168
rect 2127 -2190 2157 -2168
rect 2220 -2190 2250 -2168
rect 2306 -2190 2336 -2168
rect 2450 -2190 2480 -2168
rect 2536 -2190 2566 -2168
rect 2629 -2190 2659 -2168
rect 2707 -2190 2737 -2168
rect 2800 -2190 2830 -2168
rect 2886 -2190 2916 -2168
rect 3030 -2190 3060 -2168
rect 3116 -2190 3146 -2168
rect 3209 -2190 3239 -2168
rect 3287 -2190 3317 -2168
rect 3380 -2190 3410 -2168
rect 3466 -2190 3496 -2168
rect 3610 -2190 3640 -2168
rect 3696 -2190 3726 -2168
rect 3789 -2190 3819 -2168
rect 3867 -2190 3897 -2168
rect 3960 -2190 3990 -2168
rect 4046 -2190 4076 -2168
rect 4190 -2190 4220 -2168
rect 4276 -2190 4306 -2168
rect 4369 -2190 4399 -2168
rect 4447 -2190 4477 -2168
rect 4540 -2190 4570 -2168
rect 4626 -2190 4656 -2168
rect 4770 -2190 4800 -2168
rect 4856 -2190 4886 -2168
rect 4949 -2190 4979 -2168
rect 5027 -2190 5057 -2168
rect 5120 -2190 5150 -2168
rect 5206 -2190 5236 -2168
rect 5350 -2190 5380 -2168
rect 5436 -2190 5466 -2168
rect 5529 -2190 5559 -2168
rect 5607 -2190 5637 -2168
rect 5700 -2190 5730 -2168
rect 5786 -2190 5816 -2168
rect 5930 -2190 5960 -2168
rect 6016 -2190 6046 -2168
rect 6109 -2190 6139 -2168
rect 6187 -2190 6217 -2168
rect 6280 -2190 6310 -2168
rect 6366 -2190 6396 -2168
rect -541 -2236 6439 -2206
rect -386 -2264 -356 -2236
rect -271 -2274 -241 -2252
rect -193 -2274 -163 -2252
rect -78 -2264 -48 -2236
rect -386 -2314 -356 -2292
rect 194 -2264 224 -2236
rect 309 -2274 339 -2252
rect 387 -2274 417 -2252
rect 502 -2264 532 -2236
rect -271 -2335 -241 -2302
rect -450 -2396 -420 -2374
rect -364 -2396 -349 -2362
rect -271 -2396 -241 -2369
rect -193 -2335 -163 -2302
rect -78 -2314 -48 -2292
rect 194 -2314 224 -2292
rect 774 -2264 804 -2236
rect 889 -2274 919 -2252
rect 967 -2274 997 -2252
rect 1082 -2264 1112 -2236
rect 309 -2335 339 -2302
rect -193 -2396 -163 -2369
rect -85 -2396 -70 -2362
rect -14 -2396 16 -2374
rect 130 -2396 160 -2374
rect 216 -2396 231 -2362
rect 309 -2396 339 -2369
rect 387 -2335 417 -2302
rect 502 -2314 532 -2292
rect 774 -2314 804 -2292
rect 1354 -2264 1384 -2236
rect 1469 -2274 1499 -2252
rect 1547 -2274 1577 -2252
rect 1662 -2264 1692 -2236
rect 889 -2335 919 -2302
rect 387 -2396 417 -2369
rect 495 -2396 510 -2362
rect 566 -2396 596 -2374
rect 710 -2396 740 -2374
rect 796 -2396 811 -2362
rect 889 -2396 919 -2369
rect 967 -2335 997 -2302
rect 1082 -2314 1112 -2292
rect 1354 -2314 1384 -2292
rect 1934 -2264 1964 -2236
rect 2049 -2274 2079 -2252
rect 2127 -2274 2157 -2252
rect 2242 -2264 2272 -2236
rect 1469 -2335 1499 -2302
rect 967 -2396 997 -2369
rect 1075 -2396 1090 -2362
rect 1146 -2396 1176 -2374
rect 1290 -2396 1320 -2374
rect 1376 -2396 1391 -2362
rect 1469 -2396 1499 -2369
rect 1547 -2335 1577 -2302
rect 1662 -2314 1692 -2292
rect 1934 -2314 1964 -2292
rect 2514 -2264 2544 -2236
rect 2629 -2274 2659 -2252
rect 2707 -2274 2737 -2252
rect 2822 -2264 2852 -2236
rect 2049 -2335 2079 -2302
rect 1547 -2396 1577 -2369
rect 1655 -2396 1670 -2362
rect 1726 -2396 1756 -2374
rect 1870 -2396 1900 -2374
rect 1956 -2396 1971 -2362
rect 2049 -2396 2079 -2369
rect 2127 -2335 2157 -2302
rect 2242 -2314 2272 -2292
rect 2514 -2314 2544 -2292
rect 3094 -2264 3124 -2236
rect 3209 -2274 3239 -2252
rect 3287 -2274 3317 -2252
rect 3402 -2264 3432 -2236
rect 2629 -2335 2659 -2302
rect 2127 -2396 2157 -2369
rect 2235 -2396 2250 -2362
rect 2306 -2396 2336 -2374
rect 2450 -2396 2480 -2374
rect 2536 -2396 2551 -2362
rect 2629 -2396 2659 -2369
rect 2707 -2335 2737 -2302
rect 2822 -2314 2852 -2292
rect 3094 -2314 3124 -2292
rect 3674 -2264 3704 -2236
rect 3789 -2274 3819 -2252
rect 3867 -2274 3897 -2252
rect 3982 -2264 4012 -2236
rect 3209 -2335 3239 -2302
rect 2707 -2396 2737 -2369
rect 2815 -2396 2830 -2362
rect 2886 -2396 2916 -2374
rect 3030 -2396 3060 -2374
rect 3116 -2396 3131 -2362
rect 3209 -2396 3239 -2369
rect 3287 -2335 3317 -2302
rect 3402 -2314 3432 -2292
rect 3674 -2314 3704 -2292
rect 4254 -2264 4284 -2236
rect 4369 -2274 4399 -2252
rect 4447 -2274 4477 -2252
rect 4562 -2264 4592 -2236
rect 3789 -2335 3819 -2302
rect 3287 -2396 3317 -2369
rect 3395 -2396 3410 -2362
rect 3466 -2396 3496 -2374
rect 3610 -2396 3640 -2374
rect 3696 -2396 3711 -2362
rect 3789 -2396 3819 -2369
rect 3867 -2335 3897 -2302
rect 3982 -2314 4012 -2292
rect 4254 -2314 4284 -2292
rect 4834 -2264 4864 -2236
rect 4949 -2274 4979 -2252
rect 5027 -2274 5057 -2252
rect 5142 -2264 5172 -2236
rect 4369 -2335 4399 -2302
rect 3867 -2396 3897 -2369
rect 3975 -2396 3990 -2362
rect 4046 -2396 4076 -2374
rect 4190 -2396 4220 -2374
rect 4276 -2396 4291 -2362
rect 4369 -2396 4399 -2369
rect 4447 -2335 4477 -2302
rect 4562 -2314 4592 -2292
rect 4834 -2314 4864 -2292
rect 5414 -2264 5444 -2236
rect 5529 -2274 5559 -2252
rect 5607 -2274 5637 -2252
rect 5722 -2264 5752 -2236
rect 4949 -2335 4979 -2302
rect 4447 -2396 4477 -2369
rect 4555 -2396 4570 -2362
rect 4626 -2396 4656 -2374
rect 4770 -2396 4800 -2374
rect 4856 -2396 4871 -2362
rect 4949 -2396 4979 -2369
rect 5027 -2335 5057 -2302
rect 5142 -2314 5172 -2292
rect 5414 -2314 5444 -2292
rect 5994 -2264 6024 -2236
rect 6109 -2274 6139 -2252
rect 6187 -2274 6217 -2252
rect 6302 -2264 6332 -2236
rect 5529 -2335 5559 -2302
rect 5027 -2396 5057 -2369
rect 5135 -2396 5150 -2362
rect 5206 -2396 5236 -2374
rect 5350 -2396 5380 -2374
rect 5436 -2396 5451 -2362
rect 5529 -2396 5559 -2369
rect 5607 -2335 5637 -2302
rect 5722 -2314 5752 -2292
rect 5994 -2314 6024 -2292
rect 6109 -2335 6139 -2302
rect 5607 -2396 5637 -2369
rect 5715 -2396 5730 -2362
rect 5786 -2396 5816 -2374
rect 5930 -2396 5960 -2374
rect 6016 -2396 6031 -2362
rect 6109 -2396 6139 -2369
rect 6187 -2335 6217 -2302
rect 6302 -2314 6332 -2292
rect 6187 -2396 6217 -2369
rect 6295 -2396 6310 -2362
rect 6366 -2396 6396 -2374
rect -364 -2410 -334 -2396
rect -100 -2410 -70 -2396
rect 216 -2410 246 -2396
rect 480 -2410 510 -2396
rect 796 -2410 826 -2396
rect 1060 -2410 1090 -2396
rect 1376 -2410 1406 -2396
rect 1640 -2410 1670 -2396
rect 1956 -2410 1986 -2396
rect 2220 -2410 2250 -2396
rect 2536 -2410 2566 -2396
rect 2800 -2410 2830 -2396
rect 3116 -2410 3146 -2396
rect 3380 -2410 3410 -2396
rect 3696 -2410 3726 -2396
rect 3960 -2410 3990 -2396
rect 4276 -2410 4306 -2396
rect 4540 -2410 4570 -2396
rect 4856 -2410 4886 -2396
rect 5120 -2410 5150 -2396
rect 5436 -2410 5466 -2396
rect 5700 -2410 5730 -2396
rect 6016 -2410 6046 -2396
rect 6280 -2410 6310 -2396
rect -450 -2460 -420 -2438
rect -364 -2460 -334 -2438
rect -271 -2460 -241 -2438
rect -193 -2460 -163 -2438
rect -100 -2460 -70 -2438
rect -14 -2460 16 -2438
rect 130 -2460 160 -2438
rect 216 -2460 246 -2438
rect 309 -2460 339 -2438
rect 387 -2460 417 -2438
rect 480 -2460 510 -2438
rect 566 -2460 596 -2438
rect 710 -2460 740 -2438
rect 796 -2460 826 -2438
rect 889 -2460 919 -2438
rect 967 -2460 997 -2438
rect 1060 -2460 1090 -2438
rect 1146 -2460 1176 -2438
rect 1290 -2460 1320 -2438
rect 1376 -2460 1406 -2438
rect 1469 -2460 1499 -2438
rect 1547 -2460 1577 -2438
rect 1640 -2460 1670 -2438
rect 1726 -2460 1756 -2438
rect 1870 -2460 1900 -2438
rect 1956 -2460 1986 -2438
rect 2049 -2460 2079 -2438
rect 2127 -2460 2157 -2438
rect 2220 -2460 2250 -2438
rect 2306 -2460 2336 -2438
rect 2450 -2460 2480 -2438
rect 2536 -2460 2566 -2438
rect 2629 -2460 2659 -2438
rect 2707 -2460 2737 -2438
rect 2800 -2460 2830 -2438
rect 2886 -2460 2916 -2438
rect 3030 -2460 3060 -2438
rect 3116 -2460 3146 -2438
rect 3209 -2460 3239 -2438
rect 3287 -2460 3317 -2438
rect 3380 -2460 3410 -2438
rect 3466 -2460 3496 -2438
rect 3610 -2460 3640 -2438
rect 3696 -2460 3726 -2438
rect 3789 -2460 3819 -2438
rect 3867 -2460 3897 -2438
rect 3960 -2460 3990 -2438
rect 4046 -2460 4076 -2438
rect 4190 -2460 4220 -2438
rect 4276 -2460 4306 -2438
rect 4369 -2460 4399 -2438
rect 4447 -2460 4477 -2438
rect 4540 -2460 4570 -2438
rect 4626 -2460 4656 -2438
rect 4770 -2460 4800 -2438
rect 4856 -2460 4886 -2438
rect 4949 -2460 4979 -2438
rect 5027 -2460 5057 -2438
rect 5120 -2460 5150 -2438
rect 5206 -2460 5236 -2438
rect 5350 -2460 5380 -2438
rect 5436 -2460 5466 -2438
rect 5529 -2460 5559 -2438
rect 5607 -2460 5637 -2438
rect 5700 -2460 5730 -2438
rect 5786 -2460 5816 -2438
rect 5930 -2460 5960 -2438
rect 6016 -2460 6046 -2438
rect 6109 -2460 6139 -2438
rect 6187 -2460 6217 -2438
rect 6280 -2460 6310 -2438
rect 6366 -2460 6396 -2438
<< polycont >>
rect -450 1676 -420 1710
rect -349 1654 -319 1688
rect -271 1681 -241 1715
rect -193 1681 -163 1715
rect -115 1654 -85 1688
rect -14 1676 16 1710
rect 130 1676 160 1710
rect 231 1654 261 1688
rect 309 1681 339 1715
rect 387 1681 417 1715
rect 465 1654 495 1688
rect 566 1676 596 1710
rect 710 1676 740 1710
rect 811 1654 841 1688
rect 889 1681 919 1715
rect 967 1681 997 1715
rect 1045 1654 1075 1688
rect 1146 1676 1176 1710
rect 1290 1676 1320 1710
rect 1391 1654 1421 1688
rect 1469 1681 1499 1715
rect 1547 1681 1577 1715
rect 1625 1654 1655 1688
rect 1726 1676 1756 1710
rect 1870 1676 1900 1710
rect 1971 1654 2001 1688
rect 2049 1681 2079 1715
rect 2127 1681 2157 1715
rect 2205 1654 2235 1688
rect 2306 1676 2336 1710
rect 2450 1676 2480 1710
rect 2551 1654 2581 1688
rect 2629 1681 2659 1715
rect 2707 1681 2737 1715
rect 2785 1654 2815 1688
rect 2886 1676 2916 1710
rect 3030 1676 3060 1710
rect 3131 1654 3161 1688
rect 3209 1681 3239 1715
rect 3287 1681 3317 1715
rect 3365 1654 3395 1688
rect 3466 1676 3496 1710
rect 3610 1676 3640 1710
rect 3711 1654 3741 1688
rect 3789 1681 3819 1715
rect 3867 1681 3897 1715
rect 3945 1654 3975 1688
rect 4046 1676 4076 1710
rect 4190 1676 4220 1710
rect 4291 1654 4321 1688
rect 4369 1681 4399 1715
rect 4447 1681 4477 1715
rect 4525 1654 4555 1688
rect 4626 1676 4656 1710
rect 4770 1676 4800 1710
rect 4871 1654 4901 1688
rect 4949 1681 4979 1715
rect 5027 1681 5057 1715
rect 5105 1654 5135 1688
rect 5206 1676 5236 1710
rect 5350 1676 5380 1710
rect 5451 1654 5481 1688
rect 5529 1681 5559 1715
rect 5607 1681 5637 1715
rect 5685 1654 5715 1688
rect 5786 1676 5816 1710
rect 5930 1676 5960 1710
rect 6031 1654 6061 1688
rect 6109 1681 6139 1715
rect 6187 1681 6217 1715
rect 6265 1654 6295 1688
rect 6366 1676 6396 1710
rect -450 1406 -420 1440
rect -349 1384 -319 1418
rect -271 1411 -241 1445
rect -193 1411 -163 1445
rect -115 1384 -85 1418
rect -14 1406 16 1440
rect 130 1406 160 1440
rect 231 1384 261 1418
rect 309 1411 339 1445
rect 387 1411 417 1445
rect 465 1384 495 1418
rect 566 1406 596 1440
rect 710 1406 740 1440
rect 811 1384 841 1418
rect 889 1411 919 1445
rect 967 1411 997 1445
rect 1045 1384 1075 1418
rect 1146 1406 1176 1440
rect 1290 1406 1320 1440
rect 1391 1384 1421 1418
rect 1469 1411 1499 1445
rect 1547 1411 1577 1445
rect 1625 1384 1655 1418
rect 1726 1406 1756 1440
rect 1870 1406 1900 1440
rect 1971 1384 2001 1418
rect 2049 1411 2079 1445
rect 2127 1411 2157 1445
rect 2205 1384 2235 1418
rect 2306 1406 2336 1440
rect 2450 1406 2480 1440
rect 2551 1384 2581 1418
rect 2629 1411 2659 1445
rect 2707 1411 2737 1445
rect 2785 1384 2815 1418
rect 2886 1406 2916 1440
rect 3030 1406 3060 1440
rect 3131 1384 3161 1418
rect 3209 1411 3239 1445
rect 3287 1411 3317 1445
rect 3365 1384 3395 1418
rect 3466 1406 3496 1440
rect 3610 1406 3640 1440
rect 3711 1384 3741 1418
rect 3789 1411 3819 1445
rect 3867 1411 3897 1445
rect 3945 1384 3975 1418
rect 4046 1406 4076 1440
rect 4190 1406 4220 1440
rect 4291 1384 4321 1418
rect 4369 1411 4399 1445
rect 4447 1411 4477 1445
rect 4525 1384 4555 1418
rect 4626 1406 4656 1440
rect 4770 1406 4800 1440
rect 4871 1384 4901 1418
rect 4949 1411 4979 1445
rect 5027 1411 5057 1445
rect 5105 1384 5135 1418
rect 5206 1406 5236 1440
rect 5350 1406 5380 1440
rect 5451 1384 5481 1418
rect 5529 1411 5559 1445
rect 5607 1411 5637 1445
rect 5685 1384 5715 1418
rect 5786 1406 5816 1440
rect 5930 1406 5960 1440
rect 6031 1384 6061 1418
rect 6109 1411 6139 1445
rect 6187 1411 6217 1445
rect 6265 1384 6295 1418
rect 6366 1406 6396 1440
rect -450 1136 -420 1170
rect -349 1114 -319 1148
rect -271 1141 -241 1175
rect -193 1141 -163 1175
rect -115 1114 -85 1148
rect -14 1136 16 1170
rect 130 1136 160 1170
rect 231 1114 261 1148
rect 309 1141 339 1175
rect 387 1141 417 1175
rect 465 1114 495 1148
rect 566 1136 596 1170
rect 710 1136 740 1170
rect 811 1114 841 1148
rect 889 1141 919 1175
rect 967 1141 997 1175
rect 1045 1114 1075 1148
rect 1146 1136 1176 1170
rect 1290 1136 1320 1170
rect 1391 1114 1421 1148
rect 1469 1141 1499 1175
rect 1547 1141 1577 1175
rect 1625 1114 1655 1148
rect 1726 1136 1756 1170
rect 1870 1136 1900 1170
rect 1971 1114 2001 1148
rect 2049 1141 2079 1175
rect 2127 1141 2157 1175
rect 2205 1114 2235 1148
rect 2306 1136 2336 1170
rect 2450 1136 2480 1170
rect 2551 1114 2581 1148
rect 2629 1141 2659 1175
rect 2707 1141 2737 1175
rect 2785 1114 2815 1148
rect 2886 1136 2916 1170
rect 3030 1136 3060 1170
rect 3131 1114 3161 1148
rect 3209 1141 3239 1175
rect 3287 1141 3317 1175
rect 3365 1114 3395 1148
rect 3466 1136 3496 1170
rect 3610 1136 3640 1170
rect 3711 1114 3741 1148
rect 3789 1141 3819 1175
rect 3867 1141 3897 1175
rect 3945 1114 3975 1148
rect 4046 1136 4076 1170
rect 4190 1136 4220 1170
rect 4291 1114 4321 1148
rect 4369 1141 4399 1175
rect 4447 1141 4477 1175
rect 4525 1114 4555 1148
rect 4626 1136 4656 1170
rect 4770 1136 4800 1170
rect 4871 1114 4901 1148
rect 4949 1141 4979 1175
rect 5027 1141 5057 1175
rect 5105 1114 5135 1148
rect 5206 1136 5236 1170
rect 5350 1136 5380 1170
rect 5451 1114 5481 1148
rect 5529 1141 5559 1175
rect 5607 1141 5637 1175
rect 5685 1114 5715 1148
rect 5786 1136 5816 1170
rect 5930 1136 5960 1170
rect 6031 1114 6061 1148
rect 6109 1141 6139 1175
rect 6187 1141 6217 1175
rect 6265 1114 6295 1148
rect 6366 1136 6396 1170
rect -450 866 -420 900
rect -349 844 -319 878
rect -271 871 -241 905
rect -193 871 -163 905
rect -115 844 -85 878
rect -14 866 16 900
rect 130 866 160 900
rect 231 844 261 878
rect 309 871 339 905
rect 387 871 417 905
rect 465 844 495 878
rect 566 866 596 900
rect 710 866 740 900
rect 811 844 841 878
rect 889 871 919 905
rect 967 871 997 905
rect 1045 844 1075 878
rect 1146 866 1176 900
rect 1290 866 1320 900
rect 1391 844 1421 878
rect 1469 871 1499 905
rect 1547 871 1577 905
rect 1625 844 1655 878
rect 1726 866 1756 900
rect 1870 866 1900 900
rect 1971 844 2001 878
rect 2049 871 2079 905
rect 2127 871 2157 905
rect 2205 844 2235 878
rect 2306 866 2336 900
rect 2450 866 2480 900
rect 2551 844 2581 878
rect 2629 871 2659 905
rect 2707 871 2737 905
rect 2785 844 2815 878
rect 2886 866 2916 900
rect 3030 866 3060 900
rect 3131 844 3161 878
rect 3209 871 3239 905
rect 3287 871 3317 905
rect 3365 844 3395 878
rect 3466 866 3496 900
rect 3610 866 3640 900
rect 3711 844 3741 878
rect 3789 871 3819 905
rect 3867 871 3897 905
rect 3945 844 3975 878
rect 4046 866 4076 900
rect 4190 866 4220 900
rect 4291 844 4321 878
rect 4369 871 4399 905
rect 4447 871 4477 905
rect 4525 844 4555 878
rect 4626 866 4656 900
rect 4770 866 4800 900
rect 4871 844 4901 878
rect 4949 871 4979 905
rect 5027 871 5057 905
rect 5105 844 5135 878
rect 5206 866 5236 900
rect 5350 866 5380 900
rect 5451 844 5481 878
rect 5529 871 5559 905
rect 5607 871 5637 905
rect 5685 844 5715 878
rect 5786 866 5816 900
rect 5930 866 5960 900
rect 6031 844 6061 878
rect 6109 871 6139 905
rect 6187 871 6217 905
rect 6265 844 6295 878
rect 6366 866 6396 900
rect -450 596 -420 630
rect -349 574 -319 608
rect -271 601 -241 635
rect -193 601 -163 635
rect -115 574 -85 608
rect -14 596 16 630
rect 130 596 160 630
rect 231 574 261 608
rect 309 601 339 635
rect 387 601 417 635
rect 465 574 495 608
rect 566 596 596 630
rect 710 596 740 630
rect 811 574 841 608
rect 889 601 919 635
rect 967 601 997 635
rect 1045 574 1075 608
rect 1146 596 1176 630
rect 1290 596 1320 630
rect 1391 574 1421 608
rect 1469 601 1499 635
rect 1547 601 1577 635
rect 1625 574 1655 608
rect 1726 596 1756 630
rect 1870 596 1900 630
rect 1971 574 2001 608
rect 2049 601 2079 635
rect 2127 601 2157 635
rect 2205 574 2235 608
rect 2306 596 2336 630
rect 2450 596 2480 630
rect 2551 574 2581 608
rect 2629 601 2659 635
rect 2707 601 2737 635
rect 2785 574 2815 608
rect 2886 596 2916 630
rect 3030 596 3060 630
rect 3131 574 3161 608
rect 3209 601 3239 635
rect 3287 601 3317 635
rect 3365 574 3395 608
rect 3466 596 3496 630
rect 3610 596 3640 630
rect 3711 574 3741 608
rect 3789 601 3819 635
rect 3867 601 3897 635
rect 3945 574 3975 608
rect 4046 596 4076 630
rect 4190 596 4220 630
rect 4291 574 4321 608
rect 4369 601 4399 635
rect 4447 601 4477 635
rect 4525 574 4555 608
rect 4626 596 4656 630
rect 4770 596 4800 630
rect 4871 574 4901 608
rect 4949 601 4979 635
rect 5027 601 5057 635
rect 5105 574 5135 608
rect 5206 596 5236 630
rect 5350 596 5380 630
rect 5451 574 5481 608
rect 5529 601 5559 635
rect 5607 601 5637 635
rect 5685 574 5715 608
rect 5786 596 5816 630
rect 5930 596 5960 630
rect 6031 574 6061 608
rect 6109 601 6139 635
rect 6187 601 6217 635
rect 6265 574 6295 608
rect 6366 596 6396 630
rect -450 326 -420 360
rect -349 304 -319 338
rect -271 331 -241 365
rect -193 331 -163 365
rect -115 304 -85 338
rect -14 326 16 360
rect 130 326 160 360
rect 231 304 261 338
rect 309 331 339 365
rect 387 331 417 365
rect 465 304 495 338
rect 566 326 596 360
rect 710 326 740 360
rect 811 304 841 338
rect 889 331 919 365
rect 967 331 997 365
rect 1045 304 1075 338
rect 1146 326 1176 360
rect 1290 326 1320 360
rect 1391 304 1421 338
rect 1469 331 1499 365
rect 1547 331 1577 365
rect 1625 304 1655 338
rect 1726 326 1756 360
rect 1870 326 1900 360
rect 1971 304 2001 338
rect 2049 331 2079 365
rect 2127 331 2157 365
rect 2205 304 2235 338
rect 2306 326 2336 360
rect 2450 326 2480 360
rect 2551 304 2581 338
rect 2629 331 2659 365
rect 2707 331 2737 365
rect 2785 304 2815 338
rect 2886 326 2916 360
rect 3030 326 3060 360
rect 3131 304 3161 338
rect 3209 331 3239 365
rect 3287 331 3317 365
rect 3365 304 3395 338
rect 3466 326 3496 360
rect 3610 326 3640 360
rect 3711 304 3741 338
rect 3789 331 3819 365
rect 3867 331 3897 365
rect 3945 304 3975 338
rect 4046 326 4076 360
rect 4190 326 4220 360
rect 4291 304 4321 338
rect 4369 331 4399 365
rect 4447 331 4477 365
rect 4525 304 4555 338
rect 4626 326 4656 360
rect 4770 326 4800 360
rect 4871 304 4901 338
rect 4949 331 4979 365
rect 5027 331 5057 365
rect 5105 304 5135 338
rect 5206 326 5236 360
rect 5350 326 5380 360
rect 5451 304 5481 338
rect 5529 331 5559 365
rect 5607 331 5637 365
rect 5685 304 5715 338
rect 5786 326 5816 360
rect 5930 326 5960 360
rect 6031 304 6061 338
rect 6109 331 6139 365
rect 6187 331 6217 365
rect 6265 304 6295 338
rect 6366 326 6396 360
rect -450 56 -420 90
rect -349 34 -319 68
rect -271 61 -241 95
rect -193 61 -163 95
rect -115 34 -85 68
rect -14 56 16 90
rect 130 56 160 90
rect 231 34 261 68
rect 309 61 339 95
rect 387 61 417 95
rect 465 34 495 68
rect 566 56 596 90
rect 710 56 740 90
rect 811 34 841 68
rect 889 61 919 95
rect 967 61 997 95
rect 1045 34 1075 68
rect 1146 56 1176 90
rect 1290 56 1320 90
rect 1391 34 1421 68
rect 1469 61 1499 95
rect 1547 61 1577 95
rect 1625 34 1655 68
rect 1726 56 1756 90
rect 1870 56 1900 90
rect 1971 34 2001 68
rect 2049 61 2079 95
rect 2127 61 2157 95
rect 2205 34 2235 68
rect 2306 56 2336 90
rect 2450 56 2480 90
rect 2551 34 2581 68
rect 2629 61 2659 95
rect 2707 61 2737 95
rect 2785 34 2815 68
rect 2886 56 2916 90
rect 3030 56 3060 90
rect 3131 34 3161 68
rect 3209 61 3239 95
rect 3287 61 3317 95
rect 3365 34 3395 68
rect 3466 56 3496 90
rect 3610 56 3640 90
rect 3711 34 3741 68
rect 3789 61 3819 95
rect 3867 61 3897 95
rect 3945 34 3975 68
rect 4046 56 4076 90
rect 4190 56 4220 90
rect 4291 34 4321 68
rect 4369 61 4399 95
rect 4447 61 4477 95
rect 4525 34 4555 68
rect 4626 56 4656 90
rect 4770 56 4800 90
rect 4871 34 4901 68
rect 4949 61 4979 95
rect 5027 61 5057 95
rect 5105 34 5135 68
rect 5206 56 5236 90
rect 5350 56 5380 90
rect 5451 34 5481 68
rect 5529 61 5559 95
rect 5607 61 5637 95
rect 5685 34 5715 68
rect 5786 56 5816 90
rect 5930 56 5960 90
rect 6031 34 6061 68
rect 6109 61 6139 95
rect 6187 61 6217 95
rect 6265 34 6295 68
rect 6366 56 6396 90
rect -450 -214 -420 -180
rect -349 -236 -319 -202
rect -271 -209 -241 -175
rect -193 -209 -163 -175
rect -115 -236 -85 -202
rect -14 -214 16 -180
rect 130 -214 160 -180
rect 231 -236 261 -202
rect 309 -209 339 -175
rect 387 -209 417 -175
rect 465 -236 495 -202
rect 566 -214 596 -180
rect 710 -214 740 -180
rect 811 -236 841 -202
rect 889 -209 919 -175
rect 967 -209 997 -175
rect 1045 -236 1075 -202
rect 1146 -214 1176 -180
rect 1290 -214 1320 -180
rect 1391 -236 1421 -202
rect 1469 -209 1499 -175
rect 1547 -209 1577 -175
rect 1625 -236 1655 -202
rect 1726 -214 1756 -180
rect 1870 -214 1900 -180
rect 1971 -236 2001 -202
rect 2049 -209 2079 -175
rect 2127 -209 2157 -175
rect 2205 -236 2235 -202
rect 2306 -214 2336 -180
rect 2450 -214 2480 -180
rect 2551 -236 2581 -202
rect 2629 -209 2659 -175
rect 2707 -209 2737 -175
rect 2785 -236 2815 -202
rect 2886 -214 2916 -180
rect 3030 -214 3060 -180
rect 3131 -236 3161 -202
rect 3209 -209 3239 -175
rect 3287 -209 3317 -175
rect 3365 -236 3395 -202
rect 3466 -214 3496 -180
rect 3610 -214 3640 -180
rect 3711 -236 3741 -202
rect 3789 -209 3819 -175
rect 3867 -209 3897 -175
rect 3945 -236 3975 -202
rect 4046 -214 4076 -180
rect 4190 -214 4220 -180
rect 4291 -236 4321 -202
rect 4369 -209 4399 -175
rect 4447 -209 4477 -175
rect 4525 -236 4555 -202
rect 4626 -214 4656 -180
rect 4770 -214 4800 -180
rect 4871 -236 4901 -202
rect 4949 -209 4979 -175
rect 5027 -209 5057 -175
rect 5105 -236 5135 -202
rect 5206 -214 5236 -180
rect 5350 -214 5380 -180
rect 5451 -236 5481 -202
rect 5529 -209 5559 -175
rect 5607 -209 5637 -175
rect 5685 -236 5715 -202
rect 5786 -214 5816 -180
rect 5930 -214 5960 -180
rect 6031 -236 6061 -202
rect 6109 -209 6139 -175
rect 6187 -209 6217 -175
rect 6265 -236 6295 -202
rect 6366 -214 6396 -180
rect -450 -484 -420 -450
rect -349 -506 -319 -472
rect -271 -479 -241 -445
rect -193 -479 -163 -445
rect -115 -506 -85 -472
rect -14 -484 16 -450
rect 130 -484 160 -450
rect 231 -506 261 -472
rect 309 -479 339 -445
rect 387 -479 417 -445
rect 465 -506 495 -472
rect 566 -484 596 -450
rect 710 -484 740 -450
rect 811 -506 841 -472
rect 889 -479 919 -445
rect 967 -479 997 -445
rect 1045 -506 1075 -472
rect 1146 -484 1176 -450
rect 1290 -484 1320 -450
rect 1391 -506 1421 -472
rect 1469 -479 1499 -445
rect 1547 -479 1577 -445
rect 1625 -506 1655 -472
rect 1726 -484 1756 -450
rect 1870 -484 1900 -450
rect 1971 -506 2001 -472
rect 2049 -479 2079 -445
rect 2127 -479 2157 -445
rect 2205 -506 2235 -472
rect 2306 -484 2336 -450
rect 2450 -484 2480 -450
rect 2551 -506 2581 -472
rect 2629 -479 2659 -445
rect 2707 -479 2737 -445
rect 2785 -506 2815 -472
rect 2886 -484 2916 -450
rect 3030 -484 3060 -450
rect 3131 -506 3161 -472
rect 3209 -479 3239 -445
rect 3287 -479 3317 -445
rect 3365 -506 3395 -472
rect 3466 -484 3496 -450
rect 3610 -484 3640 -450
rect 3711 -506 3741 -472
rect 3789 -479 3819 -445
rect 3867 -479 3897 -445
rect 3945 -506 3975 -472
rect 4046 -484 4076 -450
rect 4190 -484 4220 -450
rect 4291 -506 4321 -472
rect 4369 -479 4399 -445
rect 4447 -479 4477 -445
rect 4525 -506 4555 -472
rect 4626 -484 4656 -450
rect 4770 -484 4800 -450
rect 4871 -506 4901 -472
rect 4949 -479 4979 -445
rect 5027 -479 5057 -445
rect 5105 -506 5135 -472
rect 5206 -484 5236 -450
rect 5350 -484 5380 -450
rect 5451 -506 5481 -472
rect 5529 -479 5559 -445
rect 5607 -479 5637 -445
rect 5685 -506 5715 -472
rect 5786 -484 5816 -450
rect 5930 -484 5960 -450
rect 6031 -506 6061 -472
rect 6109 -479 6139 -445
rect 6187 -479 6217 -445
rect 6265 -506 6295 -472
rect 6366 -484 6396 -450
rect -450 -754 -420 -720
rect -349 -776 -319 -742
rect -271 -749 -241 -715
rect -193 -749 -163 -715
rect -115 -776 -85 -742
rect -14 -754 16 -720
rect 130 -754 160 -720
rect 231 -776 261 -742
rect 309 -749 339 -715
rect 387 -749 417 -715
rect 465 -776 495 -742
rect 566 -754 596 -720
rect 710 -754 740 -720
rect 811 -776 841 -742
rect 889 -749 919 -715
rect 967 -749 997 -715
rect 1045 -776 1075 -742
rect 1146 -754 1176 -720
rect 1290 -754 1320 -720
rect 1391 -776 1421 -742
rect 1469 -749 1499 -715
rect 1547 -749 1577 -715
rect 1625 -776 1655 -742
rect 1726 -754 1756 -720
rect 1870 -754 1900 -720
rect 1971 -776 2001 -742
rect 2049 -749 2079 -715
rect 2127 -749 2157 -715
rect 2205 -776 2235 -742
rect 2306 -754 2336 -720
rect 2450 -754 2480 -720
rect 2551 -776 2581 -742
rect 2629 -749 2659 -715
rect 2707 -749 2737 -715
rect 2785 -776 2815 -742
rect 2886 -754 2916 -720
rect 3030 -754 3060 -720
rect 3131 -776 3161 -742
rect 3209 -749 3239 -715
rect 3287 -749 3317 -715
rect 3365 -776 3395 -742
rect 3466 -754 3496 -720
rect 3610 -754 3640 -720
rect 3711 -776 3741 -742
rect 3789 -749 3819 -715
rect 3867 -749 3897 -715
rect 3945 -776 3975 -742
rect 4046 -754 4076 -720
rect 4190 -754 4220 -720
rect 4291 -776 4321 -742
rect 4369 -749 4399 -715
rect 4447 -749 4477 -715
rect 4525 -776 4555 -742
rect 4626 -754 4656 -720
rect 4770 -754 4800 -720
rect 4871 -776 4901 -742
rect 4949 -749 4979 -715
rect 5027 -749 5057 -715
rect 5105 -776 5135 -742
rect 5206 -754 5236 -720
rect 5350 -754 5380 -720
rect 5451 -776 5481 -742
rect 5529 -749 5559 -715
rect 5607 -749 5637 -715
rect 5685 -776 5715 -742
rect 5786 -754 5816 -720
rect 5930 -754 5960 -720
rect 6031 -776 6061 -742
rect 6109 -749 6139 -715
rect 6187 -749 6217 -715
rect 6265 -776 6295 -742
rect 6366 -754 6396 -720
rect -450 -1024 -420 -990
rect -349 -1046 -319 -1012
rect -271 -1019 -241 -985
rect -193 -1019 -163 -985
rect -115 -1046 -85 -1012
rect -14 -1024 16 -990
rect 130 -1024 160 -990
rect 231 -1046 261 -1012
rect 309 -1019 339 -985
rect 387 -1019 417 -985
rect 465 -1046 495 -1012
rect 566 -1024 596 -990
rect 710 -1024 740 -990
rect 811 -1046 841 -1012
rect 889 -1019 919 -985
rect 967 -1019 997 -985
rect 1045 -1046 1075 -1012
rect 1146 -1024 1176 -990
rect 1290 -1024 1320 -990
rect 1391 -1046 1421 -1012
rect 1469 -1019 1499 -985
rect 1547 -1019 1577 -985
rect 1625 -1046 1655 -1012
rect 1726 -1024 1756 -990
rect 1870 -1024 1900 -990
rect 1971 -1046 2001 -1012
rect 2049 -1019 2079 -985
rect 2127 -1019 2157 -985
rect 2205 -1046 2235 -1012
rect 2306 -1024 2336 -990
rect 2450 -1024 2480 -990
rect 2551 -1046 2581 -1012
rect 2629 -1019 2659 -985
rect 2707 -1019 2737 -985
rect 2785 -1046 2815 -1012
rect 2886 -1024 2916 -990
rect 3030 -1024 3060 -990
rect 3131 -1046 3161 -1012
rect 3209 -1019 3239 -985
rect 3287 -1019 3317 -985
rect 3365 -1046 3395 -1012
rect 3466 -1024 3496 -990
rect 3610 -1024 3640 -990
rect 3711 -1046 3741 -1012
rect 3789 -1019 3819 -985
rect 3867 -1019 3897 -985
rect 3945 -1046 3975 -1012
rect 4046 -1024 4076 -990
rect 4190 -1024 4220 -990
rect 4291 -1046 4321 -1012
rect 4369 -1019 4399 -985
rect 4447 -1019 4477 -985
rect 4525 -1046 4555 -1012
rect 4626 -1024 4656 -990
rect 4770 -1024 4800 -990
rect 4871 -1046 4901 -1012
rect 4949 -1019 4979 -985
rect 5027 -1019 5057 -985
rect 5105 -1046 5135 -1012
rect 5206 -1024 5236 -990
rect 5350 -1024 5380 -990
rect 5451 -1046 5481 -1012
rect 5529 -1019 5559 -985
rect 5607 -1019 5637 -985
rect 5685 -1046 5715 -1012
rect 5786 -1024 5816 -990
rect 5930 -1024 5960 -990
rect 6031 -1046 6061 -1012
rect 6109 -1019 6139 -985
rect 6187 -1019 6217 -985
rect 6265 -1046 6295 -1012
rect 6366 -1024 6396 -990
rect -450 -1294 -420 -1260
rect -349 -1316 -319 -1282
rect -271 -1289 -241 -1255
rect -193 -1289 -163 -1255
rect -115 -1316 -85 -1282
rect -14 -1294 16 -1260
rect 130 -1294 160 -1260
rect 231 -1316 261 -1282
rect 309 -1289 339 -1255
rect 387 -1289 417 -1255
rect 465 -1316 495 -1282
rect 566 -1294 596 -1260
rect 710 -1294 740 -1260
rect 811 -1316 841 -1282
rect 889 -1289 919 -1255
rect 967 -1289 997 -1255
rect 1045 -1316 1075 -1282
rect 1146 -1294 1176 -1260
rect 1290 -1294 1320 -1260
rect 1391 -1316 1421 -1282
rect 1469 -1289 1499 -1255
rect 1547 -1289 1577 -1255
rect 1625 -1316 1655 -1282
rect 1726 -1294 1756 -1260
rect 1870 -1294 1900 -1260
rect 1971 -1316 2001 -1282
rect 2049 -1289 2079 -1255
rect 2127 -1289 2157 -1255
rect 2205 -1316 2235 -1282
rect 2306 -1294 2336 -1260
rect 2450 -1294 2480 -1260
rect 2551 -1316 2581 -1282
rect 2629 -1289 2659 -1255
rect 2707 -1289 2737 -1255
rect 2785 -1316 2815 -1282
rect 2886 -1294 2916 -1260
rect 3030 -1294 3060 -1260
rect 3131 -1316 3161 -1282
rect 3209 -1289 3239 -1255
rect 3287 -1289 3317 -1255
rect 3365 -1316 3395 -1282
rect 3466 -1294 3496 -1260
rect 3610 -1294 3640 -1260
rect 3711 -1316 3741 -1282
rect 3789 -1289 3819 -1255
rect 3867 -1289 3897 -1255
rect 3945 -1316 3975 -1282
rect 4046 -1294 4076 -1260
rect 4190 -1294 4220 -1260
rect 4291 -1316 4321 -1282
rect 4369 -1289 4399 -1255
rect 4447 -1289 4477 -1255
rect 4525 -1316 4555 -1282
rect 4626 -1294 4656 -1260
rect 4770 -1294 4800 -1260
rect 4871 -1316 4901 -1282
rect 4949 -1289 4979 -1255
rect 5027 -1289 5057 -1255
rect 5105 -1316 5135 -1282
rect 5206 -1294 5236 -1260
rect 5350 -1294 5380 -1260
rect 5451 -1316 5481 -1282
rect 5529 -1289 5559 -1255
rect 5607 -1289 5637 -1255
rect 5685 -1316 5715 -1282
rect 5786 -1294 5816 -1260
rect 5930 -1294 5960 -1260
rect 6031 -1316 6061 -1282
rect 6109 -1289 6139 -1255
rect 6187 -1289 6217 -1255
rect 6265 -1316 6295 -1282
rect 6366 -1294 6396 -1260
rect -450 -1564 -420 -1530
rect -349 -1586 -319 -1552
rect -271 -1559 -241 -1525
rect -193 -1559 -163 -1525
rect -115 -1586 -85 -1552
rect -14 -1564 16 -1530
rect 130 -1564 160 -1530
rect 231 -1586 261 -1552
rect 309 -1559 339 -1525
rect 387 -1559 417 -1525
rect 465 -1586 495 -1552
rect 566 -1564 596 -1530
rect 710 -1564 740 -1530
rect 811 -1586 841 -1552
rect 889 -1559 919 -1525
rect 967 -1559 997 -1525
rect 1045 -1586 1075 -1552
rect 1146 -1564 1176 -1530
rect 1290 -1564 1320 -1530
rect 1391 -1586 1421 -1552
rect 1469 -1559 1499 -1525
rect 1547 -1559 1577 -1525
rect 1625 -1586 1655 -1552
rect 1726 -1564 1756 -1530
rect 1870 -1564 1900 -1530
rect 1971 -1586 2001 -1552
rect 2049 -1559 2079 -1525
rect 2127 -1559 2157 -1525
rect 2205 -1586 2235 -1552
rect 2306 -1564 2336 -1530
rect 2450 -1564 2480 -1530
rect 2551 -1586 2581 -1552
rect 2629 -1559 2659 -1525
rect 2707 -1559 2737 -1525
rect 2785 -1586 2815 -1552
rect 2886 -1564 2916 -1530
rect 3030 -1564 3060 -1530
rect 3131 -1586 3161 -1552
rect 3209 -1559 3239 -1525
rect 3287 -1559 3317 -1525
rect 3365 -1586 3395 -1552
rect 3466 -1564 3496 -1530
rect 3610 -1564 3640 -1530
rect 3711 -1586 3741 -1552
rect 3789 -1559 3819 -1525
rect 3867 -1559 3897 -1525
rect 3945 -1586 3975 -1552
rect 4046 -1564 4076 -1530
rect 4190 -1564 4220 -1530
rect 4291 -1586 4321 -1552
rect 4369 -1559 4399 -1525
rect 4447 -1559 4477 -1525
rect 4525 -1586 4555 -1552
rect 4626 -1564 4656 -1530
rect 4770 -1564 4800 -1530
rect 4871 -1586 4901 -1552
rect 4949 -1559 4979 -1525
rect 5027 -1559 5057 -1525
rect 5105 -1586 5135 -1552
rect 5206 -1564 5236 -1530
rect 5350 -1564 5380 -1530
rect 5451 -1586 5481 -1552
rect 5529 -1559 5559 -1525
rect 5607 -1559 5637 -1525
rect 5685 -1586 5715 -1552
rect 5786 -1564 5816 -1530
rect 5930 -1564 5960 -1530
rect 6031 -1586 6061 -1552
rect 6109 -1559 6139 -1525
rect 6187 -1559 6217 -1525
rect 6265 -1586 6295 -1552
rect 6366 -1564 6396 -1530
rect -450 -1834 -420 -1800
rect -349 -1856 -319 -1822
rect -271 -1829 -241 -1795
rect -193 -1829 -163 -1795
rect -115 -1856 -85 -1822
rect -14 -1834 16 -1800
rect 130 -1834 160 -1800
rect 231 -1856 261 -1822
rect 309 -1829 339 -1795
rect 387 -1829 417 -1795
rect 465 -1856 495 -1822
rect 566 -1834 596 -1800
rect 710 -1834 740 -1800
rect 811 -1856 841 -1822
rect 889 -1829 919 -1795
rect 967 -1829 997 -1795
rect 1045 -1856 1075 -1822
rect 1146 -1834 1176 -1800
rect 1290 -1834 1320 -1800
rect 1391 -1856 1421 -1822
rect 1469 -1829 1499 -1795
rect 1547 -1829 1577 -1795
rect 1625 -1856 1655 -1822
rect 1726 -1834 1756 -1800
rect 1870 -1834 1900 -1800
rect 1971 -1856 2001 -1822
rect 2049 -1829 2079 -1795
rect 2127 -1829 2157 -1795
rect 2205 -1856 2235 -1822
rect 2306 -1834 2336 -1800
rect 2450 -1834 2480 -1800
rect 2551 -1856 2581 -1822
rect 2629 -1829 2659 -1795
rect 2707 -1829 2737 -1795
rect 2785 -1856 2815 -1822
rect 2886 -1834 2916 -1800
rect 3030 -1834 3060 -1800
rect 3131 -1856 3161 -1822
rect 3209 -1829 3239 -1795
rect 3287 -1829 3317 -1795
rect 3365 -1856 3395 -1822
rect 3466 -1834 3496 -1800
rect 3610 -1834 3640 -1800
rect 3711 -1856 3741 -1822
rect 3789 -1829 3819 -1795
rect 3867 -1829 3897 -1795
rect 3945 -1856 3975 -1822
rect 4046 -1834 4076 -1800
rect 4190 -1834 4220 -1800
rect 4291 -1856 4321 -1822
rect 4369 -1829 4399 -1795
rect 4447 -1829 4477 -1795
rect 4525 -1856 4555 -1822
rect 4626 -1834 4656 -1800
rect 4770 -1834 4800 -1800
rect 4871 -1856 4901 -1822
rect 4949 -1829 4979 -1795
rect 5027 -1829 5057 -1795
rect 5105 -1856 5135 -1822
rect 5206 -1834 5236 -1800
rect 5350 -1834 5380 -1800
rect 5451 -1856 5481 -1822
rect 5529 -1829 5559 -1795
rect 5607 -1829 5637 -1795
rect 5685 -1856 5715 -1822
rect 5786 -1834 5816 -1800
rect 5930 -1834 5960 -1800
rect 6031 -1856 6061 -1822
rect 6109 -1829 6139 -1795
rect 6187 -1829 6217 -1795
rect 6265 -1856 6295 -1822
rect 6366 -1834 6396 -1800
rect -450 -2104 -420 -2070
rect -349 -2126 -319 -2092
rect -271 -2099 -241 -2065
rect -193 -2099 -163 -2065
rect -115 -2126 -85 -2092
rect -14 -2104 16 -2070
rect 130 -2104 160 -2070
rect 231 -2126 261 -2092
rect 309 -2099 339 -2065
rect 387 -2099 417 -2065
rect 465 -2126 495 -2092
rect 566 -2104 596 -2070
rect 710 -2104 740 -2070
rect 811 -2126 841 -2092
rect 889 -2099 919 -2065
rect 967 -2099 997 -2065
rect 1045 -2126 1075 -2092
rect 1146 -2104 1176 -2070
rect 1290 -2104 1320 -2070
rect 1391 -2126 1421 -2092
rect 1469 -2099 1499 -2065
rect 1547 -2099 1577 -2065
rect 1625 -2126 1655 -2092
rect 1726 -2104 1756 -2070
rect 1870 -2104 1900 -2070
rect 1971 -2126 2001 -2092
rect 2049 -2099 2079 -2065
rect 2127 -2099 2157 -2065
rect 2205 -2126 2235 -2092
rect 2306 -2104 2336 -2070
rect 2450 -2104 2480 -2070
rect 2551 -2126 2581 -2092
rect 2629 -2099 2659 -2065
rect 2707 -2099 2737 -2065
rect 2785 -2126 2815 -2092
rect 2886 -2104 2916 -2070
rect 3030 -2104 3060 -2070
rect 3131 -2126 3161 -2092
rect 3209 -2099 3239 -2065
rect 3287 -2099 3317 -2065
rect 3365 -2126 3395 -2092
rect 3466 -2104 3496 -2070
rect 3610 -2104 3640 -2070
rect 3711 -2126 3741 -2092
rect 3789 -2099 3819 -2065
rect 3867 -2099 3897 -2065
rect 3945 -2126 3975 -2092
rect 4046 -2104 4076 -2070
rect 4190 -2104 4220 -2070
rect 4291 -2126 4321 -2092
rect 4369 -2099 4399 -2065
rect 4447 -2099 4477 -2065
rect 4525 -2126 4555 -2092
rect 4626 -2104 4656 -2070
rect 4770 -2104 4800 -2070
rect 4871 -2126 4901 -2092
rect 4949 -2099 4979 -2065
rect 5027 -2099 5057 -2065
rect 5105 -2126 5135 -2092
rect 5206 -2104 5236 -2070
rect 5350 -2104 5380 -2070
rect 5451 -2126 5481 -2092
rect 5529 -2099 5559 -2065
rect 5607 -2099 5637 -2065
rect 5685 -2126 5715 -2092
rect 5786 -2104 5816 -2070
rect 5930 -2104 5960 -2070
rect 6031 -2126 6061 -2092
rect 6109 -2099 6139 -2065
rect 6187 -2099 6217 -2065
rect 6265 -2126 6295 -2092
rect 6366 -2104 6396 -2070
rect -450 -2374 -420 -2340
rect -349 -2396 -319 -2362
rect -271 -2369 -241 -2335
rect -193 -2369 -163 -2335
rect -115 -2396 -85 -2362
rect -14 -2374 16 -2340
rect 130 -2374 160 -2340
rect 231 -2396 261 -2362
rect 309 -2369 339 -2335
rect 387 -2369 417 -2335
rect 465 -2396 495 -2362
rect 566 -2374 596 -2340
rect 710 -2374 740 -2340
rect 811 -2396 841 -2362
rect 889 -2369 919 -2335
rect 967 -2369 997 -2335
rect 1045 -2396 1075 -2362
rect 1146 -2374 1176 -2340
rect 1290 -2374 1320 -2340
rect 1391 -2396 1421 -2362
rect 1469 -2369 1499 -2335
rect 1547 -2369 1577 -2335
rect 1625 -2396 1655 -2362
rect 1726 -2374 1756 -2340
rect 1870 -2374 1900 -2340
rect 1971 -2396 2001 -2362
rect 2049 -2369 2079 -2335
rect 2127 -2369 2157 -2335
rect 2205 -2396 2235 -2362
rect 2306 -2374 2336 -2340
rect 2450 -2374 2480 -2340
rect 2551 -2396 2581 -2362
rect 2629 -2369 2659 -2335
rect 2707 -2369 2737 -2335
rect 2785 -2396 2815 -2362
rect 2886 -2374 2916 -2340
rect 3030 -2374 3060 -2340
rect 3131 -2396 3161 -2362
rect 3209 -2369 3239 -2335
rect 3287 -2369 3317 -2335
rect 3365 -2396 3395 -2362
rect 3466 -2374 3496 -2340
rect 3610 -2374 3640 -2340
rect 3711 -2396 3741 -2362
rect 3789 -2369 3819 -2335
rect 3867 -2369 3897 -2335
rect 3945 -2396 3975 -2362
rect 4046 -2374 4076 -2340
rect 4190 -2374 4220 -2340
rect 4291 -2396 4321 -2362
rect 4369 -2369 4399 -2335
rect 4447 -2369 4477 -2335
rect 4525 -2396 4555 -2362
rect 4626 -2374 4656 -2340
rect 4770 -2374 4800 -2340
rect 4871 -2396 4901 -2362
rect 4949 -2369 4979 -2335
rect 5027 -2369 5057 -2335
rect 5105 -2396 5135 -2362
rect 5206 -2374 5236 -2340
rect 5350 -2374 5380 -2340
rect 5451 -2396 5481 -2362
rect 5529 -2369 5559 -2335
rect 5607 -2369 5637 -2335
rect 5685 -2396 5715 -2362
rect 5786 -2374 5816 -2340
rect 5930 -2374 5960 -2340
rect 6031 -2396 6061 -2362
rect 6109 -2369 6139 -2335
rect 6187 -2369 6217 -2335
rect 6265 -2396 6295 -2362
rect 6366 -2374 6396 -2340
<< corelocali >>
rect -493 1654 -478 1892
tri -413 1808 -391 1830 se
rect -391 1823 -376 1892
tri -391 1808 -376 1823 nw
rect -57 1823 -42 1893
tri -419 1802 -413 1808 se
rect -413 1802 -404 1808
rect -419 1786 -404 1802
tri -404 1795 -391 1808 nw
rect -250 1800 -233 1814
rect -201 1800 -184 1814
tri -57 1808 -42 1823 ne
tri -42 1808 -20 1830 sw
rect -419 1750 -404 1758
rect -338 1786 -278 1800
rect -323 1776 -278 1786
rect -323 1758 -295 1776
tri -419 1735 -404 1750 ne
tri -404 1735 -382 1757 sw
rect -338 1748 -295 1758
rect -280 1772 -278 1776
rect -156 1786 -96 1800
tri -42 1795 -29 1808 ne
rect -29 1802 -20 1808
tri -20 1802 -14 1808 sw
rect -156 1776 -111 1786
rect -280 1748 -206 1772
rect -338 1744 -206 1748
tri -206 1744 -178 1772 sw
rect -156 1762 -154 1776
tri -156 1760 -154 1762 ne
rect -142 1758 -111 1776
rect -142 1748 -96 1758
rect -29 1787 -14 1802
tri -404 1723 -392 1735 ne
rect -392 1730 -382 1735
tri -382 1730 -377 1735 sw
rect -493 1384 -478 1612
rect -392 1574 -377 1730
rect -338 1688 -310 1744
tri -218 1726 -200 1744 ne
rect -200 1724 -178 1744
tri -178 1724 -158 1744 sw
tri -142 1730 -124 1748 ne
rect -319 1654 -310 1688
rect -276 1715 -234 1716
rect -276 1681 -271 1715
rect -241 1681 -234 1715
rect -276 1672 -234 1681
rect -200 1715 -158 1724
rect -200 1681 -193 1715
rect -163 1681 -158 1715
rect -200 1676 -158 1681
rect -124 1688 -96 1748
tri -51 1735 -29 1757 se
rect -29 1750 -14 1758
tri -29 1735 -14 1750 nw
tri -57 1729 -51 1735 se
rect -51 1729 -42 1735
rect -338 1644 -310 1654
tri -310 1644 -286 1668 sw
rect -338 1612 -296 1644
tri -279 1636 -278 1637 sw
rect -279 1612 -278 1636
tri -276 1635 -239 1672 ne
rect -239 1644 -234 1672
tri -234 1644 -208 1670 sw
rect -124 1654 -115 1688
rect -124 1644 -96 1654
rect -239 1635 -155 1644
tri -239 1616 -220 1635 ne
rect -220 1616 -155 1635
rect -338 1590 -278 1612
rect -156 1612 -155 1616
rect -138 1612 -96 1644
rect -156 1590 -96 1612
rect -250 1574 -233 1588
rect -201 1574 -184 1588
tri -413 1538 -391 1560 se
rect -391 1553 -376 1574
tri -391 1538 -376 1553 nw
rect -57 1553 -42 1729
tri -42 1722 -29 1735 nw
rect 44 1654 59 1892
tri -419 1532 -413 1538 se
rect -413 1532 -404 1538
rect -419 1516 -404 1532
tri -404 1525 -391 1538 nw
rect -250 1530 -233 1544
rect -201 1530 -184 1544
tri -57 1538 -42 1553 ne
tri -42 1538 -20 1560 sw
rect -419 1480 -404 1488
rect -338 1516 -278 1530
rect -323 1506 -278 1516
rect -323 1488 -295 1506
tri -419 1465 -404 1480 ne
tri -404 1465 -382 1487 sw
rect -338 1478 -295 1488
rect -280 1502 -278 1506
rect -156 1516 -96 1530
tri -42 1525 -29 1538 ne
rect -29 1532 -20 1538
tri -20 1532 -14 1538 sw
rect -156 1506 -111 1516
rect -280 1478 -206 1502
rect -338 1474 -206 1478
tri -206 1474 -178 1502 sw
rect -156 1492 -154 1506
tri -156 1490 -154 1492 ne
rect -142 1488 -111 1506
rect -142 1478 -96 1488
rect -29 1517 -14 1532
tri -404 1453 -392 1465 ne
rect -392 1460 -382 1465
tri -382 1460 -377 1465 sw
rect -493 1114 -478 1342
rect -392 1352 -377 1460
rect -338 1418 -310 1474
tri -218 1456 -200 1474 ne
rect -200 1454 -178 1474
tri -178 1454 -158 1474 sw
tri -142 1460 -124 1478 ne
rect -319 1384 -310 1418
rect -276 1445 -234 1446
rect -276 1411 -271 1445
rect -241 1411 -234 1445
rect -276 1402 -234 1411
rect -200 1445 -158 1454
rect -200 1411 -193 1445
rect -163 1411 -158 1445
rect -200 1406 -158 1411
rect -124 1418 -96 1478
tri -51 1465 -29 1487 se
rect -29 1480 -14 1488
tri -29 1465 -14 1480 nw
tri -57 1459 -51 1465 se
rect -51 1459 -42 1465
rect -338 1374 -310 1384
tri -310 1374 -286 1398 sw
rect -392 1304 -376 1352
rect -338 1342 -296 1374
tri -279 1366 -278 1367 sw
rect -279 1342 -278 1366
tri -276 1365 -239 1402 ne
rect -239 1374 -234 1402
tri -234 1374 -208 1400 sw
rect -124 1384 -115 1418
rect -124 1374 -96 1384
rect -239 1365 -155 1374
tri -239 1346 -220 1365 ne
rect -220 1346 -155 1365
rect -338 1320 -278 1342
rect -156 1342 -155 1346
rect -138 1342 -96 1374
rect -156 1320 -96 1342
rect -250 1304 -233 1318
rect -201 1304 -184 1318
tri -413 1268 -391 1290 se
rect -391 1283 -376 1304
tri -391 1268 -376 1283 nw
rect -57 1283 -42 1459
tri -42 1452 -29 1465 nw
rect 44 1384 59 1612
tri -419 1262 -413 1268 se
rect -413 1262 -404 1268
rect -419 1246 -404 1262
tri -404 1255 -391 1268 nw
rect -250 1260 -233 1274
rect -201 1260 -184 1274
tri -57 1268 -42 1283 ne
tri -42 1268 -20 1290 sw
rect -419 1210 -404 1218
rect -338 1246 -278 1260
rect -323 1236 -278 1246
rect -323 1218 -295 1236
tri -419 1195 -404 1210 ne
tri -404 1195 -382 1217 sw
rect -338 1208 -295 1218
rect -280 1232 -278 1236
rect -156 1246 -96 1260
tri -42 1255 -29 1268 ne
rect -29 1262 -20 1268
tri -20 1262 -14 1268 sw
rect -156 1236 -111 1246
rect -280 1208 -206 1232
rect -338 1204 -206 1208
tri -206 1204 -178 1232 sw
rect -156 1222 -154 1236
tri -156 1220 -154 1222 ne
rect -142 1218 -111 1236
rect -142 1208 -96 1218
rect -29 1247 -14 1262
tri -404 1183 -392 1195 ne
rect -392 1190 -382 1195
tri -382 1190 -377 1195 sw
rect -493 844 -478 1072
rect -392 1034 -377 1190
rect -338 1148 -310 1204
tri -218 1186 -200 1204 ne
rect -200 1184 -178 1204
tri -178 1184 -158 1204 sw
tri -142 1190 -124 1208 ne
rect -319 1114 -310 1148
rect -276 1175 -234 1176
rect -276 1141 -271 1175
rect -241 1141 -234 1175
rect -276 1132 -234 1141
rect -200 1175 -158 1184
rect -200 1141 -193 1175
rect -163 1141 -158 1175
rect -200 1136 -158 1141
rect -124 1148 -96 1208
tri -51 1195 -29 1217 se
rect -29 1210 -14 1218
tri -29 1195 -14 1210 nw
tri -57 1189 -51 1195 se
rect -51 1189 -42 1195
rect -338 1104 -310 1114
tri -310 1104 -286 1128 sw
rect -338 1072 -296 1104
tri -279 1096 -278 1097 sw
rect -279 1072 -278 1096
tri -276 1095 -239 1132 ne
rect -239 1104 -234 1132
tri -234 1104 -208 1130 sw
rect -124 1114 -115 1148
rect -124 1104 -96 1114
rect -239 1095 -155 1104
tri -239 1076 -220 1095 ne
rect -220 1076 -155 1095
rect -338 1050 -278 1072
rect -156 1072 -155 1076
rect -138 1072 -96 1104
rect -156 1050 -96 1072
rect -250 1034 -233 1048
rect -201 1034 -184 1048
tri -413 998 -391 1020 se
rect -391 1013 -376 1034
tri -391 998 -376 1013 nw
rect -57 1013 -42 1189
tri -42 1182 -29 1195 nw
rect 44 1114 59 1342
tri -419 992 -413 998 se
rect -413 992 -404 998
rect -419 976 -404 992
tri -404 985 -391 998 nw
rect -250 990 -233 1004
rect -201 990 -184 1004
tri -57 998 -42 1013 ne
tri -42 998 -20 1020 sw
rect -419 940 -404 948
rect -338 976 -278 990
rect -323 966 -278 976
rect -323 948 -295 966
tri -419 925 -404 940 ne
tri -404 925 -382 947 sw
rect -338 938 -295 948
rect -280 962 -278 966
rect -156 976 -96 990
tri -42 985 -29 998 ne
rect -29 992 -20 998
tri -20 992 -14 998 sw
rect -156 966 -111 976
rect -280 938 -206 962
rect -338 934 -206 938
tri -206 934 -178 962 sw
rect -156 952 -154 966
tri -156 950 -154 952 ne
rect -142 948 -111 966
rect -142 938 -96 948
rect -29 977 -14 992
tri -404 913 -392 925 ne
rect -392 920 -382 925
tri -382 920 -377 925 sw
rect -493 574 -478 802
rect -392 812 -377 920
rect -338 878 -310 934
tri -218 916 -200 934 ne
rect -200 914 -178 934
tri -178 914 -158 934 sw
tri -142 920 -124 938 ne
rect -319 844 -310 878
rect -276 905 -234 906
rect -276 871 -271 905
rect -241 871 -234 905
rect -276 862 -234 871
rect -200 905 -158 914
rect -200 871 -193 905
rect -163 871 -158 905
rect -200 866 -158 871
rect -124 878 -96 938
tri -51 925 -29 947 se
rect -29 940 -14 948
tri -29 925 -14 940 nw
tri -57 919 -51 925 se
rect -51 919 -42 925
rect -338 834 -310 844
tri -310 834 -286 858 sw
rect -392 764 -376 812
rect -338 802 -296 834
tri -279 826 -278 827 sw
rect -279 802 -278 826
tri -276 825 -239 862 ne
rect -239 834 -234 862
tri -234 834 -208 860 sw
rect -124 844 -115 878
rect -124 834 -96 844
rect -239 825 -155 834
tri -239 806 -220 825 ne
rect -220 806 -155 825
rect -338 780 -278 802
rect -156 802 -155 806
rect -138 802 -96 834
rect -156 780 -96 802
rect -250 764 -233 778
rect -201 764 -184 778
tri -413 728 -391 750 se
rect -391 743 -376 764
tri -391 728 -376 743 nw
rect -57 743 -42 919
tri -42 912 -29 925 nw
rect 44 844 59 1072
tri -419 722 -413 728 se
rect -413 722 -404 728
rect -419 706 -404 722
tri -404 715 -391 728 nw
rect -250 720 -233 734
rect -201 720 -184 734
tri -57 728 -42 743 ne
tri -42 728 -20 750 sw
rect -419 670 -404 678
rect -338 706 -278 720
rect -323 696 -278 706
rect -323 678 -295 696
tri -419 655 -404 670 ne
tri -404 655 -382 677 sw
rect -338 668 -295 678
rect -280 692 -278 696
rect -156 706 -96 720
tri -42 715 -29 728 ne
rect -29 722 -20 728
tri -20 722 -14 728 sw
rect -156 696 -111 706
rect -280 668 -206 692
rect -338 664 -206 668
tri -206 664 -178 692 sw
rect -156 682 -154 696
tri -156 680 -154 682 ne
rect -142 678 -111 696
rect -142 668 -96 678
rect -29 707 -14 722
tri -404 643 -392 655 ne
rect -392 650 -382 655
tri -382 650 -377 655 sw
rect -493 304 -478 532
rect -392 494 -377 650
rect -338 608 -310 664
tri -218 646 -200 664 ne
rect -200 644 -178 664
tri -178 644 -158 664 sw
tri -142 650 -124 668 ne
rect -319 574 -310 608
rect -276 635 -234 636
rect -276 601 -271 635
rect -241 601 -234 635
rect -276 592 -234 601
rect -200 635 -158 644
rect -200 601 -193 635
rect -163 601 -158 635
rect -200 596 -158 601
rect -124 608 -96 668
tri -51 655 -29 677 se
rect -29 670 -14 678
tri -29 655 -14 670 nw
tri -57 649 -51 655 se
rect -51 649 -42 655
rect -338 564 -310 574
tri -310 564 -286 588 sw
rect -338 532 -296 564
tri -279 556 -278 557 sw
rect -279 532 -278 556
tri -276 555 -239 592 ne
rect -239 564 -234 592
tri -234 564 -208 590 sw
rect -124 574 -115 608
rect -124 564 -96 574
rect -239 555 -155 564
tri -239 536 -220 555 ne
rect -220 536 -155 555
rect -338 510 -278 532
rect -156 532 -155 536
rect -138 532 -96 564
rect -156 510 -96 532
rect -250 494 -233 508
rect -201 494 -184 508
tri -413 458 -391 480 se
rect -391 473 -376 494
tri -391 458 -376 473 nw
rect -57 473 -42 649
tri -42 642 -29 655 nw
rect 44 574 59 802
tri -419 452 -413 458 se
rect -413 452 -404 458
rect -419 436 -404 452
tri -404 445 -391 458 nw
rect -250 450 -233 464
rect -201 450 -184 464
tri -57 458 -42 473 ne
tri -42 458 -20 480 sw
rect -419 400 -404 408
rect -338 436 -278 450
rect -323 426 -278 436
rect -323 408 -295 426
tri -419 385 -404 400 ne
tri -404 385 -382 407 sw
rect -338 398 -295 408
rect -280 422 -278 426
rect -156 436 -96 450
tri -42 445 -29 458 ne
rect -29 452 -20 458
tri -20 452 -14 458 sw
rect -156 426 -111 436
rect -280 398 -206 422
rect -338 394 -206 398
tri -206 394 -178 422 sw
rect -156 412 -154 426
tri -156 410 -154 412 ne
rect -142 408 -111 426
rect -142 398 -96 408
rect -29 437 -14 452
tri -404 373 -392 385 ne
rect -392 380 -382 385
tri -382 380 -377 385 sw
rect -493 34 -478 262
rect -392 272 -377 380
rect -338 338 -310 394
tri -218 376 -200 394 ne
rect -200 374 -178 394
tri -178 374 -158 394 sw
tri -142 380 -124 398 ne
rect -319 304 -310 338
rect -276 365 -234 366
rect -276 331 -271 365
rect -241 331 -234 365
rect -276 322 -234 331
rect -200 365 -158 374
rect -200 331 -193 365
rect -163 331 -158 365
rect -200 326 -158 331
rect -124 338 -96 398
tri -51 385 -29 407 se
rect -29 400 -14 408
tri -29 385 -14 400 nw
tri -57 379 -51 385 se
rect -51 379 -42 385
rect -338 294 -310 304
tri -310 294 -286 318 sw
rect -392 224 -376 272
rect -338 262 -296 294
tri -279 286 -278 287 sw
rect -279 262 -278 286
tri -276 285 -239 322 ne
rect -239 294 -234 322
tri -234 294 -208 320 sw
rect -124 304 -115 338
rect -124 294 -96 304
rect -239 285 -155 294
tri -239 266 -220 285 ne
rect -220 266 -155 285
rect -338 240 -278 262
rect -156 262 -155 266
rect -138 262 -96 294
rect -156 240 -96 262
rect -250 224 -233 238
rect -201 224 -184 238
tri -413 188 -391 210 se
rect -391 203 -376 224
tri -391 188 -376 203 nw
rect -57 203 -42 379
tri -42 372 -29 385 nw
rect 44 304 59 532
tri -419 182 -413 188 se
rect -413 182 -404 188
rect -419 166 -404 182
tri -404 175 -391 188 nw
rect -250 180 -233 194
rect -201 180 -184 194
tri -57 188 -42 203 ne
tri -42 188 -20 210 sw
rect -419 130 -404 138
rect -338 166 -278 180
rect -323 156 -278 166
rect -323 138 -295 156
tri -419 115 -404 130 ne
tri -404 115 -382 137 sw
rect -338 128 -295 138
rect -280 152 -278 156
rect -156 166 -96 180
tri -42 175 -29 188 ne
rect -29 182 -20 188
tri -20 182 -14 188 sw
rect -156 156 -111 166
rect -280 128 -206 152
rect -338 124 -206 128
tri -206 124 -178 152 sw
rect -156 142 -154 156
tri -156 140 -154 142 ne
rect -142 138 -111 156
rect -142 128 -96 138
rect -29 167 -14 182
tri -404 103 -392 115 ne
rect -392 110 -382 115
tri -382 110 -377 115 sw
rect -493 -236 -478 -8
rect -392 -46 -377 110
rect -338 68 -310 124
tri -218 106 -200 124 ne
rect -200 104 -178 124
tri -178 104 -158 124 sw
tri -142 110 -124 128 ne
rect -319 34 -310 68
rect -276 95 -234 96
rect -276 61 -271 95
rect -241 61 -234 95
rect -276 52 -234 61
rect -200 95 -158 104
rect -200 61 -193 95
rect -163 61 -158 95
rect -200 56 -158 61
rect -124 68 -96 128
tri -51 115 -29 137 se
rect -29 130 -14 138
tri -29 115 -14 130 nw
tri -57 109 -51 115 se
rect -51 109 -42 115
rect -338 24 -310 34
tri -310 24 -286 48 sw
rect -338 -8 -296 24
tri -279 16 -278 17 sw
rect -279 -8 -278 16
tri -276 15 -239 52 ne
rect -239 24 -234 52
tri -234 24 -208 50 sw
rect -124 34 -115 68
rect -124 24 -96 34
rect -239 15 -155 24
tri -239 -4 -220 15 ne
rect -220 -4 -155 15
rect -338 -30 -278 -8
rect -156 -8 -155 -4
rect -138 -8 -96 24
rect -156 -30 -96 -8
rect -250 -46 -233 -32
rect -201 -46 -184 -32
tri -413 -82 -391 -60 se
rect -391 -67 -376 -46
tri -391 -82 -376 -67 nw
rect -57 -67 -42 109
tri -42 102 -29 115 nw
rect 44 34 59 262
tri -419 -88 -413 -82 se
rect -413 -88 -404 -82
rect -419 -104 -404 -88
tri -404 -95 -391 -82 nw
rect -250 -90 -233 -76
rect -201 -90 -184 -76
tri -57 -82 -42 -67 ne
tri -42 -82 -20 -60 sw
rect -419 -140 -404 -132
rect -338 -104 -278 -90
rect -323 -114 -278 -104
rect -323 -132 -295 -114
tri -419 -155 -404 -140 ne
tri -404 -155 -382 -133 sw
rect -338 -142 -295 -132
rect -280 -118 -278 -114
rect -156 -104 -96 -90
tri -42 -95 -29 -82 ne
rect -29 -88 -20 -82
tri -20 -88 -14 -82 sw
rect -156 -114 -111 -104
rect -280 -142 -206 -118
rect -338 -146 -206 -142
tri -206 -146 -178 -118 sw
rect -156 -128 -154 -114
tri -156 -130 -154 -128 ne
rect -142 -132 -111 -114
rect -142 -142 -96 -132
rect -29 -103 -14 -88
tri -404 -167 -392 -155 ne
rect -392 -160 -382 -155
tri -382 -160 -377 -155 sw
rect -493 -506 -478 -278
rect -392 -268 -377 -160
rect -338 -202 -310 -146
tri -218 -164 -200 -146 ne
rect -200 -166 -178 -146
tri -178 -166 -158 -146 sw
tri -142 -160 -124 -142 ne
rect -319 -236 -310 -202
rect -276 -175 -234 -174
rect -276 -209 -271 -175
rect -241 -209 -234 -175
rect -276 -218 -234 -209
rect -200 -175 -158 -166
rect -200 -209 -193 -175
rect -163 -209 -158 -175
rect -200 -214 -158 -209
rect -124 -202 -96 -142
tri -51 -155 -29 -133 se
rect -29 -140 -14 -132
tri -29 -155 -14 -140 nw
tri -57 -161 -51 -155 se
rect -51 -161 -42 -155
rect -338 -246 -310 -236
tri -310 -246 -286 -222 sw
rect -392 -316 -376 -268
rect -338 -278 -296 -246
tri -279 -254 -278 -253 sw
rect -279 -278 -278 -254
tri -276 -255 -239 -218 ne
rect -239 -246 -234 -218
tri -234 -246 -208 -220 sw
rect -124 -236 -115 -202
rect -124 -246 -96 -236
rect -239 -255 -155 -246
tri -239 -274 -220 -255 ne
rect -220 -274 -155 -255
rect -338 -300 -278 -278
rect -156 -278 -155 -274
rect -138 -278 -96 -246
rect -156 -300 -96 -278
rect -250 -316 -233 -302
rect -201 -316 -184 -302
tri -413 -352 -391 -330 se
rect -391 -337 -376 -316
tri -391 -352 -376 -337 nw
rect -57 -337 -42 -161
tri -42 -168 -29 -155 nw
rect 44 -236 59 -8
tri -419 -358 -413 -352 se
rect -413 -358 -404 -352
rect -419 -374 -404 -358
tri -404 -365 -391 -352 nw
rect -250 -360 -233 -346
rect -201 -360 -184 -346
tri -57 -352 -42 -337 ne
tri -42 -352 -20 -330 sw
rect -419 -410 -404 -402
rect -338 -374 -278 -360
rect -323 -384 -278 -374
rect -323 -402 -295 -384
tri -419 -425 -404 -410 ne
tri -404 -425 -382 -403 sw
rect -338 -412 -295 -402
rect -280 -388 -278 -384
rect -156 -374 -96 -360
tri -42 -365 -29 -352 ne
rect -29 -358 -20 -352
tri -20 -358 -14 -352 sw
rect -156 -384 -111 -374
rect -280 -412 -206 -388
rect -338 -416 -206 -412
tri -206 -416 -178 -388 sw
rect -156 -398 -154 -384
tri -156 -400 -154 -398 ne
rect -142 -402 -111 -384
rect -142 -412 -96 -402
rect -29 -373 -14 -358
tri -404 -437 -392 -425 ne
rect -392 -430 -382 -425
tri -382 -430 -377 -425 sw
rect -493 -776 -478 -548
rect -392 -586 -377 -430
rect -338 -472 -310 -416
tri -218 -434 -200 -416 ne
rect -200 -436 -178 -416
tri -178 -436 -158 -416 sw
tri -142 -430 -124 -412 ne
rect -319 -506 -310 -472
rect -276 -445 -234 -444
rect -276 -479 -271 -445
rect -241 -479 -234 -445
rect -276 -488 -234 -479
rect -200 -445 -158 -436
rect -200 -479 -193 -445
rect -163 -479 -158 -445
rect -200 -484 -158 -479
rect -124 -472 -96 -412
tri -51 -425 -29 -403 se
rect -29 -410 -14 -402
tri -29 -425 -14 -410 nw
tri -57 -431 -51 -425 se
rect -51 -431 -42 -425
rect -338 -516 -310 -506
tri -310 -516 -286 -492 sw
rect -338 -548 -296 -516
tri -279 -524 -278 -523 sw
rect -279 -548 -278 -524
tri -276 -525 -239 -488 ne
rect -239 -516 -234 -488
tri -234 -516 -208 -490 sw
rect -124 -506 -115 -472
rect -124 -516 -96 -506
rect -239 -525 -155 -516
tri -239 -544 -220 -525 ne
rect -220 -544 -155 -525
rect -338 -570 -278 -548
rect -156 -548 -155 -544
rect -138 -548 -96 -516
rect -156 -570 -96 -548
rect -250 -586 -233 -572
rect -201 -586 -184 -572
tri -413 -622 -391 -600 se
rect -391 -607 -376 -586
tri -391 -622 -376 -607 nw
rect -57 -607 -42 -431
tri -42 -438 -29 -425 nw
rect 44 -506 59 -278
tri -419 -628 -413 -622 se
rect -413 -628 -404 -622
rect -419 -644 -404 -628
tri -404 -635 -391 -622 nw
rect -250 -630 -233 -616
rect -201 -630 -184 -616
tri -57 -622 -42 -607 ne
tri -42 -622 -20 -600 sw
rect -419 -680 -404 -672
rect -338 -644 -278 -630
rect -323 -654 -278 -644
rect -323 -672 -295 -654
tri -419 -695 -404 -680 ne
tri -404 -695 -382 -673 sw
rect -338 -682 -295 -672
rect -280 -658 -278 -654
rect -156 -644 -96 -630
tri -42 -635 -29 -622 ne
rect -29 -628 -20 -622
tri -20 -628 -14 -622 sw
rect -156 -654 -111 -644
rect -280 -682 -206 -658
rect -338 -686 -206 -682
tri -206 -686 -178 -658 sw
rect -156 -668 -154 -654
tri -156 -670 -154 -668 ne
rect -142 -672 -111 -654
rect -142 -682 -96 -672
rect -29 -643 -14 -628
tri -404 -707 -392 -695 ne
rect -392 -700 -382 -695
tri -382 -700 -377 -695 sw
rect -493 -1046 -478 -818
rect -392 -808 -377 -700
rect -338 -742 -310 -686
tri -218 -704 -200 -686 ne
rect -200 -706 -178 -686
tri -178 -706 -158 -686 sw
tri -142 -700 -124 -682 ne
rect -319 -776 -310 -742
rect -276 -715 -234 -714
rect -276 -749 -271 -715
rect -241 -749 -234 -715
rect -276 -758 -234 -749
rect -200 -715 -158 -706
rect -200 -749 -193 -715
rect -163 -749 -158 -715
rect -200 -754 -158 -749
rect -124 -742 -96 -682
tri -51 -695 -29 -673 se
rect -29 -680 -14 -672
tri -29 -695 -14 -680 nw
tri -57 -701 -51 -695 se
rect -51 -701 -42 -695
rect -338 -786 -310 -776
tri -310 -786 -286 -762 sw
rect -392 -856 -376 -808
rect -338 -818 -296 -786
tri -279 -794 -278 -793 sw
rect -279 -818 -278 -794
tri -276 -795 -239 -758 ne
rect -239 -786 -234 -758
tri -234 -786 -208 -760 sw
rect -124 -776 -115 -742
rect -124 -786 -96 -776
rect -239 -795 -155 -786
tri -239 -814 -220 -795 ne
rect -220 -814 -155 -795
rect -338 -840 -278 -818
rect -156 -818 -155 -814
rect -138 -818 -96 -786
rect -156 -840 -96 -818
rect -250 -856 -233 -842
rect -201 -856 -184 -842
tri -413 -892 -391 -870 se
rect -391 -877 -376 -856
tri -391 -892 -376 -877 nw
rect -57 -877 -42 -701
tri -42 -708 -29 -695 nw
rect 44 -776 59 -548
tri -419 -898 -413 -892 se
rect -413 -898 -404 -892
rect -419 -914 -404 -898
tri -404 -905 -391 -892 nw
rect -250 -900 -233 -886
rect -201 -900 -184 -886
tri -57 -892 -42 -877 ne
tri -42 -892 -20 -870 sw
rect -419 -950 -404 -942
rect -338 -914 -278 -900
rect -323 -924 -278 -914
rect -323 -942 -295 -924
tri -419 -965 -404 -950 ne
tri -404 -965 -382 -943 sw
rect -338 -952 -295 -942
rect -280 -928 -278 -924
rect -156 -914 -96 -900
tri -42 -905 -29 -892 ne
rect -29 -898 -20 -892
tri -20 -898 -14 -892 sw
rect -156 -924 -111 -914
rect -280 -952 -206 -928
rect -338 -956 -206 -952
tri -206 -956 -178 -928 sw
rect -156 -938 -154 -924
tri -156 -940 -154 -938 ne
rect -142 -942 -111 -924
rect -142 -952 -96 -942
rect -29 -913 -14 -898
tri -404 -977 -392 -965 ne
rect -392 -970 -382 -965
tri -382 -970 -377 -965 sw
rect -493 -1316 -478 -1088
rect -392 -1126 -377 -970
rect -338 -1012 -310 -956
tri -218 -974 -200 -956 ne
rect -200 -976 -178 -956
tri -178 -976 -158 -956 sw
tri -142 -970 -124 -952 ne
rect -319 -1046 -310 -1012
rect -276 -985 -234 -984
rect -276 -1019 -271 -985
rect -241 -1019 -234 -985
rect -276 -1028 -234 -1019
rect -200 -985 -158 -976
rect -200 -1019 -193 -985
rect -163 -1019 -158 -985
rect -200 -1024 -158 -1019
rect -124 -1012 -96 -952
tri -51 -965 -29 -943 se
rect -29 -950 -14 -942
tri -29 -965 -14 -950 nw
tri -57 -971 -51 -965 se
rect -51 -971 -42 -965
rect -338 -1056 -310 -1046
tri -310 -1056 -286 -1032 sw
rect -338 -1088 -296 -1056
tri -279 -1064 -278 -1063 sw
rect -279 -1088 -278 -1064
tri -276 -1065 -239 -1028 ne
rect -239 -1056 -234 -1028
tri -234 -1056 -208 -1030 sw
rect -124 -1046 -115 -1012
rect -124 -1056 -96 -1046
rect -239 -1065 -155 -1056
tri -239 -1084 -220 -1065 ne
rect -220 -1084 -155 -1065
rect -338 -1110 -278 -1088
rect -156 -1088 -155 -1084
rect -138 -1088 -96 -1056
rect -156 -1110 -96 -1088
rect -250 -1126 -233 -1112
rect -201 -1126 -184 -1112
tri -413 -1162 -391 -1140 se
rect -391 -1147 -376 -1126
tri -391 -1162 -376 -1147 nw
rect -57 -1147 -42 -971
tri -42 -978 -29 -965 nw
rect 44 -1046 59 -818
tri -419 -1168 -413 -1162 se
rect -413 -1168 -404 -1162
rect -419 -1184 -404 -1168
tri -404 -1175 -391 -1162 nw
rect -250 -1170 -233 -1156
rect -201 -1170 -184 -1156
tri -57 -1162 -42 -1147 ne
tri -42 -1162 -20 -1140 sw
rect -419 -1220 -404 -1212
rect -338 -1184 -278 -1170
rect -323 -1194 -278 -1184
rect -323 -1212 -295 -1194
tri -419 -1235 -404 -1220 ne
tri -404 -1235 -382 -1213 sw
rect -338 -1222 -295 -1212
rect -280 -1198 -278 -1194
rect -156 -1184 -96 -1170
tri -42 -1175 -29 -1162 ne
rect -29 -1168 -20 -1162
tri -20 -1168 -14 -1162 sw
rect -156 -1194 -111 -1184
rect -280 -1222 -206 -1198
rect -338 -1226 -206 -1222
tri -206 -1226 -178 -1198 sw
rect -156 -1208 -154 -1194
tri -156 -1210 -154 -1208 ne
rect -142 -1212 -111 -1194
rect -142 -1222 -96 -1212
rect -29 -1183 -14 -1168
tri -404 -1247 -392 -1235 ne
rect -392 -1240 -382 -1235
tri -382 -1240 -377 -1235 sw
rect -493 -1586 -478 -1358
rect -392 -1348 -377 -1240
rect -338 -1282 -310 -1226
tri -218 -1244 -200 -1226 ne
rect -200 -1246 -178 -1226
tri -178 -1246 -158 -1226 sw
tri -142 -1240 -124 -1222 ne
rect -319 -1316 -310 -1282
rect -276 -1255 -234 -1254
rect -276 -1289 -271 -1255
rect -241 -1289 -234 -1255
rect -276 -1298 -234 -1289
rect -200 -1255 -158 -1246
rect -200 -1289 -193 -1255
rect -163 -1289 -158 -1255
rect -200 -1294 -158 -1289
rect -124 -1282 -96 -1222
tri -51 -1235 -29 -1213 se
rect -29 -1220 -14 -1212
tri -29 -1235 -14 -1220 nw
tri -57 -1241 -51 -1235 se
rect -51 -1241 -42 -1235
rect -338 -1326 -310 -1316
tri -310 -1326 -286 -1302 sw
rect -392 -1396 -376 -1348
rect -338 -1358 -296 -1326
tri -279 -1334 -278 -1333 sw
rect -279 -1358 -278 -1334
tri -276 -1335 -239 -1298 ne
rect -239 -1326 -234 -1298
tri -234 -1326 -208 -1300 sw
rect -124 -1316 -115 -1282
rect -124 -1326 -96 -1316
rect -239 -1335 -155 -1326
tri -239 -1354 -220 -1335 ne
rect -220 -1354 -155 -1335
rect -338 -1380 -278 -1358
rect -156 -1358 -155 -1354
rect -138 -1358 -96 -1326
rect -156 -1380 -96 -1358
rect -250 -1396 -233 -1382
rect -201 -1396 -184 -1382
tri -413 -1432 -391 -1410 se
rect -391 -1417 -376 -1396
tri -391 -1432 -376 -1417 nw
rect -57 -1417 -42 -1241
tri -42 -1248 -29 -1235 nw
rect 44 -1316 59 -1088
tri -419 -1438 -413 -1432 se
rect -413 -1438 -404 -1432
rect -419 -1454 -404 -1438
tri -404 -1445 -391 -1432 nw
rect -250 -1440 -233 -1426
rect -201 -1440 -184 -1426
tri -57 -1432 -42 -1417 ne
tri -42 -1432 -20 -1410 sw
rect -419 -1490 -404 -1482
rect -338 -1454 -278 -1440
rect -323 -1464 -278 -1454
rect -323 -1482 -295 -1464
tri -419 -1505 -404 -1490 ne
tri -404 -1505 -382 -1483 sw
rect -338 -1492 -295 -1482
rect -280 -1468 -278 -1464
rect -156 -1454 -96 -1440
tri -42 -1445 -29 -1432 ne
rect -29 -1438 -20 -1432
tri -20 -1438 -14 -1432 sw
rect -156 -1464 -111 -1454
rect -280 -1492 -206 -1468
rect -338 -1496 -206 -1492
tri -206 -1496 -178 -1468 sw
rect -156 -1478 -154 -1464
tri -156 -1480 -154 -1478 ne
rect -142 -1482 -111 -1464
rect -142 -1492 -96 -1482
rect -29 -1453 -14 -1438
tri -404 -1517 -392 -1505 ne
rect -392 -1510 -382 -1505
tri -382 -1510 -377 -1505 sw
rect -493 -1856 -478 -1628
rect -392 -1666 -377 -1510
rect -338 -1552 -310 -1496
tri -218 -1514 -200 -1496 ne
rect -200 -1516 -178 -1496
tri -178 -1516 -158 -1496 sw
tri -142 -1510 -124 -1492 ne
rect -319 -1586 -310 -1552
rect -276 -1525 -234 -1524
rect -276 -1559 -271 -1525
rect -241 -1559 -234 -1525
rect -276 -1568 -234 -1559
rect -200 -1525 -158 -1516
rect -200 -1559 -193 -1525
rect -163 -1559 -158 -1525
rect -200 -1564 -158 -1559
rect -124 -1552 -96 -1492
tri -51 -1505 -29 -1483 se
rect -29 -1490 -14 -1482
tri -29 -1505 -14 -1490 nw
tri -57 -1511 -51 -1505 se
rect -51 -1511 -42 -1505
rect -338 -1596 -310 -1586
tri -310 -1596 -286 -1572 sw
rect -338 -1628 -296 -1596
tri -279 -1604 -278 -1603 sw
rect -279 -1628 -278 -1604
tri -276 -1605 -239 -1568 ne
rect -239 -1596 -234 -1568
tri -234 -1596 -208 -1570 sw
rect -124 -1586 -115 -1552
rect -124 -1596 -96 -1586
rect -239 -1605 -155 -1596
tri -239 -1624 -220 -1605 ne
rect -220 -1624 -155 -1605
rect -338 -1650 -278 -1628
rect -156 -1628 -155 -1624
rect -138 -1628 -96 -1596
rect -156 -1650 -96 -1628
rect -250 -1666 -233 -1652
rect -201 -1666 -184 -1652
tri -413 -1702 -391 -1680 se
rect -391 -1687 -376 -1666
tri -391 -1702 -376 -1687 nw
rect -57 -1687 -42 -1511
tri -42 -1518 -29 -1505 nw
rect 44 -1586 59 -1358
tri -419 -1708 -413 -1702 se
rect -413 -1708 -404 -1702
rect -419 -1724 -404 -1708
tri -404 -1715 -391 -1702 nw
rect -250 -1710 -233 -1696
rect -201 -1710 -184 -1696
tri -57 -1702 -42 -1687 ne
tri -42 -1702 -20 -1680 sw
rect -419 -1760 -404 -1752
rect -338 -1724 -278 -1710
rect -323 -1734 -278 -1724
rect -323 -1752 -295 -1734
tri -419 -1775 -404 -1760 ne
tri -404 -1775 -382 -1753 sw
rect -338 -1762 -295 -1752
rect -280 -1738 -278 -1734
rect -156 -1724 -96 -1710
tri -42 -1715 -29 -1702 ne
rect -29 -1708 -20 -1702
tri -20 -1708 -14 -1702 sw
rect -156 -1734 -111 -1724
rect -280 -1762 -206 -1738
rect -338 -1766 -206 -1762
tri -206 -1766 -178 -1738 sw
rect -156 -1748 -154 -1734
tri -156 -1750 -154 -1748 ne
rect -142 -1752 -111 -1734
rect -142 -1762 -96 -1752
rect -29 -1723 -14 -1708
tri -404 -1787 -392 -1775 ne
rect -392 -1780 -382 -1775
tri -382 -1780 -377 -1775 sw
rect -493 -2126 -478 -1898
rect -392 -1888 -377 -1780
rect -338 -1822 -310 -1766
tri -218 -1784 -200 -1766 ne
rect -200 -1786 -178 -1766
tri -178 -1786 -158 -1766 sw
tri -142 -1780 -124 -1762 ne
rect -319 -1856 -310 -1822
rect -276 -1795 -234 -1794
rect -276 -1829 -271 -1795
rect -241 -1829 -234 -1795
rect -276 -1838 -234 -1829
rect -200 -1795 -158 -1786
rect -200 -1829 -193 -1795
rect -163 -1829 -158 -1795
rect -200 -1834 -158 -1829
rect -124 -1822 -96 -1762
tri -51 -1775 -29 -1753 se
rect -29 -1760 -14 -1752
tri -29 -1775 -14 -1760 nw
tri -57 -1781 -51 -1775 se
rect -51 -1781 -42 -1775
rect -338 -1866 -310 -1856
tri -310 -1866 -286 -1842 sw
rect -392 -1936 -376 -1888
rect -338 -1898 -296 -1866
tri -279 -1874 -278 -1873 sw
rect -279 -1898 -278 -1874
tri -276 -1875 -239 -1838 ne
rect -239 -1866 -234 -1838
tri -234 -1866 -208 -1840 sw
rect -124 -1856 -115 -1822
rect -124 -1866 -96 -1856
rect -239 -1875 -155 -1866
tri -239 -1894 -220 -1875 ne
rect -220 -1894 -155 -1875
rect -338 -1920 -278 -1898
rect -156 -1898 -155 -1894
rect -138 -1898 -96 -1866
rect -156 -1920 -96 -1898
rect -250 -1936 -233 -1922
rect -201 -1936 -184 -1922
tri -413 -1972 -391 -1950 se
rect -391 -1957 -376 -1936
tri -391 -1972 -376 -1957 nw
rect -57 -1957 -42 -1781
tri -42 -1788 -29 -1775 nw
rect 44 -1856 59 -1628
tri -419 -1978 -413 -1972 se
rect -413 -1978 -404 -1972
rect -419 -1994 -404 -1978
tri -404 -1985 -391 -1972 nw
rect -250 -1980 -233 -1966
rect -201 -1980 -184 -1966
tri -57 -1972 -42 -1957 ne
tri -42 -1972 -20 -1950 sw
rect -419 -2030 -404 -2022
rect -338 -1994 -278 -1980
rect -323 -2004 -278 -1994
rect -323 -2022 -295 -2004
tri -419 -2045 -404 -2030 ne
tri -404 -2045 -382 -2023 sw
rect -338 -2032 -295 -2022
rect -280 -2008 -278 -2004
rect -156 -1994 -96 -1980
tri -42 -1985 -29 -1972 ne
rect -29 -1978 -20 -1972
tri -20 -1978 -14 -1972 sw
rect -156 -2004 -111 -1994
rect -280 -2032 -206 -2008
rect -338 -2036 -206 -2032
tri -206 -2036 -178 -2008 sw
rect -156 -2018 -154 -2004
tri -156 -2020 -154 -2018 ne
rect -142 -2022 -111 -2004
rect -142 -2032 -96 -2022
rect -29 -1993 -14 -1978
tri -404 -2057 -392 -2045 ne
rect -392 -2050 -382 -2045
tri -382 -2050 -377 -2045 sw
rect -493 -2396 -478 -2168
rect -392 -2206 -377 -2050
rect -338 -2092 -310 -2036
tri -218 -2054 -200 -2036 ne
rect -200 -2056 -178 -2036
tri -178 -2056 -158 -2036 sw
tri -142 -2050 -124 -2032 ne
rect -319 -2126 -310 -2092
rect -276 -2065 -234 -2064
rect -276 -2099 -271 -2065
rect -241 -2099 -234 -2065
rect -276 -2108 -234 -2099
rect -200 -2065 -158 -2056
rect -200 -2099 -193 -2065
rect -163 -2099 -158 -2065
rect -200 -2104 -158 -2099
rect -124 -2092 -96 -2032
tri -51 -2045 -29 -2023 se
rect -29 -2030 -14 -2022
tri -29 -2045 -14 -2030 nw
tri -57 -2051 -51 -2045 se
rect -51 -2051 -42 -2045
rect -338 -2136 -310 -2126
tri -310 -2136 -286 -2112 sw
rect -338 -2168 -296 -2136
tri -279 -2144 -278 -2143 sw
rect -279 -2168 -278 -2144
tri -276 -2145 -239 -2108 ne
rect -239 -2136 -234 -2108
tri -234 -2136 -208 -2110 sw
rect -124 -2126 -115 -2092
rect -124 -2136 -96 -2126
rect -239 -2145 -155 -2136
tri -239 -2164 -220 -2145 ne
rect -220 -2164 -155 -2145
rect -338 -2190 -278 -2168
rect -156 -2168 -155 -2164
rect -138 -2168 -96 -2136
rect -156 -2190 -96 -2168
rect -250 -2206 -233 -2192
rect -201 -2206 -184 -2192
tri -413 -2242 -391 -2220 se
rect -391 -2227 -376 -2206
tri -391 -2242 -376 -2227 nw
rect -57 -2227 -42 -2051
tri -42 -2058 -29 -2045 nw
rect 44 -2126 59 -1898
tri -419 -2248 -413 -2242 se
rect -413 -2248 -404 -2242
rect -419 -2264 -404 -2248
tri -404 -2255 -391 -2242 nw
rect -250 -2250 -233 -2236
rect -201 -2250 -184 -2236
tri -57 -2242 -42 -2227 ne
tri -42 -2242 -20 -2220 sw
rect -419 -2300 -404 -2292
rect -338 -2264 -278 -2250
rect -323 -2274 -278 -2264
rect -323 -2292 -295 -2274
tri -419 -2315 -404 -2300 ne
tri -404 -2315 -382 -2293 sw
rect -338 -2302 -295 -2292
rect -280 -2278 -278 -2274
rect -156 -2264 -96 -2250
tri -42 -2255 -29 -2242 ne
rect -29 -2248 -20 -2242
tri -20 -2248 -14 -2242 sw
rect -156 -2274 -111 -2264
rect -280 -2302 -206 -2278
rect -338 -2306 -206 -2302
tri -206 -2306 -178 -2278 sw
rect -156 -2288 -154 -2274
tri -156 -2290 -154 -2288 ne
rect -142 -2292 -111 -2274
rect -142 -2302 -96 -2292
rect -29 -2263 -14 -2248
tri -404 -2327 -392 -2315 ne
rect -392 -2320 -382 -2315
tri -382 -2320 -377 -2315 sw
rect -493 -2524 -478 -2438
rect -392 -2476 -377 -2320
rect -338 -2362 -310 -2306
tri -218 -2324 -200 -2306 ne
rect -200 -2326 -178 -2306
tri -178 -2326 -158 -2306 sw
tri -142 -2320 -124 -2302 ne
rect -319 -2396 -310 -2362
rect -276 -2335 -234 -2334
rect -276 -2369 -271 -2335
rect -241 -2369 -234 -2335
rect -276 -2378 -234 -2369
rect -200 -2335 -158 -2326
rect -200 -2369 -193 -2335
rect -163 -2369 -158 -2335
rect -200 -2374 -158 -2369
rect -124 -2362 -96 -2302
tri -51 -2315 -29 -2293 se
rect -29 -2300 -14 -2292
tri -29 -2315 -14 -2300 nw
tri -57 -2321 -51 -2315 se
rect -51 -2321 -42 -2315
rect -338 -2406 -310 -2396
tri -310 -2406 -286 -2382 sw
rect -338 -2438 -296 -2406
tri -279 -2414 -278 -2413 sw
rect -279 -2438 -278 -2414
tri -276 -2415 -239 -2378 ne
rect -239 -2406 -234 -2378
tri -234 -2406 -208 -2380 sw
rect -124 -2396 -115 -2362
rect -124 -2406 -96 -2396
rect -239 -2415 -155 -2406
tri -239 -2434 -220 -2415 ne
rect -220 -2434 -155 -2415
rect -338 -2460 -278 -2438
rect -156 -2438 -155 -2434
rect -138 -2438 -96 -2406
rect -156 -2460 -96 -2438
rect -250 -2476 -233 -2462
rect -201 -2476 -184 -2462
rect -57 -2476 -42 -2321
tri -42 -2328 -29 -2315 nw
rect 44 -2396 59 -2168
rect 44 -2524 59 -2438
rect 87 1654 102 1892
tri 167 1808 189 1830 se
rect 189 1823 204 1892
tri 189 1808 204 1823 nw
rect 523 1823 538 1892
tri 161 1802 167 1808 se
rect 167 1802 176 1808
rect 161 1786 176 1802
tri 176 1795 189 1808 nw
rect 330 1800 347 1814
rect 379 1800 396 1814
tri 523 1808 538 1823 ne
tri 538 1808 560 1830 sw
rect 161 1750 176 1758
rect 242 1786 302 1800
rect 257 1776 302 1786
rect 257 1758 285 1776
tri 161 1735 176 1750 ne
tri 176 1735 198 1757 sw
rect 242 1748 285 1758
rect 300 1772 302 1776
rect 424 1786 484 1800
tri 538 1795 551 1808 ne
rect 551 1802 560 1808
tri 560 1802 566 1808 sw
rect 424 1776 469 1786
rect 300 1748 374 1772
rect 242 1744 374 1748
tri 374 1744 402 1772 sw
rect 424 1762 426 1776
tri 424 1760 426 1762 ne
rect 438 1758 469 1776
rect 438 1748 484 1758
rect 551 1787 566 1802
tri 176 1723 188 1735 ne
rect 188 1730 198 1735
tri 198 1730 203 1735 sw
rect 87 1384 102 1612
rect 188 1574 203 1730
rect 242 1688 270 1744
tri 362 1726 380 1744 ne
rect 380 1724 402 1744
tri 402 1724 422 1744 sw
tri 438 1730 456 1748 ne
rect 261 1654 270 1688
rect 304 1715 346 1716
rect 304 1681 309 1715
rect 339 1681 346 1715
rect 304 1672 346 1681
rect 380 1715 422 1724
rect 380 1681 387 1715
rect 417 1681 422 1715
rect 380 1676 422 1681
rect 456 1688 484 1748
tri 529 1735 551 1757 se
rect 551 1750 566 1758
tri 551 1735 566 1750 nw
tri 523 1729 529 1735 se
rect 529 1729 538 1735
rect 242 1644 270 1654
tri 270 1644 294 1668 sw
rect 242 1612 284 1644
tri 301 1636 302 1637 sw
rect 301 1612 302 1636
tri 304 1635 341 1672 ne
rect 341 1644 346 1672
tri 346 1644 372 1670 sw
rect 456 1654 465 1688
rect 456 1644 484 1654
rect 341 1635 425 1644
tri 341 1616 360 1635 ne
rect 360 1616 425 1635
rect 242 1590 302 1612
rect 424 1612 425 1616
rect 442 1612 484 1644
rect 424 1590 484 1612
rect 330 1574 347 1588
rect 379 1574 396 1588
tri 167 1538 189 1560 se
rect 189 1553 204 1574
tri 189 1538 204 1553 nw
rect 523 1553 538 1729
tri 538 1722 551 1735 nw
rect 624 1654 639 1892
tri 161 1532 167 1538 se
rect 167 1532 176 1538
rect 161 1516 176 1532
tri 176 1525 189 1538 nw
rect 330 1530 347 1544
rect 379 1530 396 1544
tri 523 1538 538 1553 ne
tri 538 1538 560 1560 sw
rect 161 1480 176 1488
rect 242 1516 302 1530
rect 257 1506 302 1516
rect 257 1488 285 1506
tri 161 1465 176 1480 ne
tri 176 1465 198 1487 sw
rect 242 1478 285 1488
rect 300 1502 302 1506
rect 424 1516 484 1530
tri 538 1525 551 1538 ne
rect 551 1532 560 1538
tri 560 1532 566 1538 sw
rect 424 1506 469 1516
rect 300 1478 374 1502
rect 242 1474 374 1478
tri 374 1474 402 1502 sw
rect 424 1492 426 1506
tri 424 1490 426 1492 ne
rect 438 1488 469 1506
rect 438 1478 484 1488
rect 551 1517 566 1532
tri 176 1453 188 1465 ne
rect 188 1460 198 1465
tri 198 1460 203 1465 sw
rect 87 1114 102 1342
rect 188 1352 203 1460
rect 242 1418 270 1474
tri 362 1456 380 1474 ne
rect 380 1454 402 1474
tri 402 1454 422 1474 sw
tri 438 1460 456 1478 ne
rect 261 1384 270 1418
rect 304 1445 346 1446
rect 304 1411 309 1445
rect 339 1411 346 1445
rect 304 1402 346 1411
rect 380 1445 422 1454
rect 380 1411 387 1445
rect 417 1411 422 1445
rect 380 1406 422 1411
rect 456 1418 484 1478
tri 529 1465 551 1487 se
rect 551 1480 566 1488
tri 551 1465 566 1480 nw
tri 523 1459 529 1465 se
rect 529 1459 538 1465
rect 242 1374 270 1384
tri 270 1374 294 1398 sw
rect 188 1304 204 1352
rect 242 1342 284 1374
tri 301 1366 302 1367 sw
rect 301 1342 302 1366
tri 304 1365 341 1402 ne
rect 341 1374 346 1402
tri 346 1374 372 1400 sw
rect 456 1384 465 1418
rect 456 1374 484 1384
rect 341 1365 425 1374
tri 341 1346 360 1365 ne
rect 360 1346 425 1365
rect 242 1320 302 1342
rect 424 1342 425 1346
rect 442 1342 484 1374
rect 424 1320 484 1342
rect 330 1304 347 1318
rect 379 1304 396 1318
tri 167 1268 189 1290 se
rect 189 1283 204 1304
tri 189 1268 204 1283 nw
rect 523 1283 538 1459
tri 538 1452 551 1465 nw
rect 624 1384 639 1612
tri 161 1262 167 1268 se
rect 167 1262 176 1268
rect 161 1246 176 1262
tri 176 1255 189 1268 nw
rect 330 1260 347 1274
rect 379 1260 396 1274
tri 523 1268 538 1283 ne
tri 538 1268 560 1290 sw
rect 161 1210 176 1218
rect 242 1246 302 1260
rect 257 1236 302 1246
rect 257 1218 285 1236
tri 161 1195 176 1210 ne
tri 176 1195 198 1217 sw
rect 242 1208 285 1218
rect 300 1232 302 1236
rect 424 1246 484 1260
tri 538 1255 551 1268 ne
rect 551 1262 560 1268
tri 560 1262 566 1268 sw
rect 424 1236 469 1246
rect 300 1208 374 1232
rect 242 1204 374 1208
tri 374 1204 402 1232 sw
rect 424 1222 426 1236
tri 424 1220 426 1222 ne
rect 438 1218 469 1236
rect 438 1208 484 1218
rect 551 1247 566 1262
tri 176 1183 188 1195 ne
rect 188 1190 198 1195
tri 198 1190 203 1195 sw
rect 87 844 102 1072
rect 188 1034 203 1190
rect 242 1148 270 1204
tri 362 1186 380 1204 ne
rect 380 1184 402 1204
tri 402 1184 422 1204 sw
tri 438 1190 456 1208 ne
rect 261 1114 270 1148
rect 304 1175 346 1176
rect 304 1141 309 1175
rect 339 1141 346 1175
rect 304 1132 346 1141
rect 380 1175 422 1184
rect 380 1141 387 1175
rect 417 1141 422 1175
rect 380 1136 422 1141
rect 456 1148 484 1208
tri 529 1195 551 1217 se
rect 551 1210 566 1218
tri 551 1195 566 1210 nw
tri 523 1189 529 1195 se
rect 529 1189 538 1195
rect 242 1104 270 1114
tri 270 1104 294 1128 sw
rect 242 1072 284 1104
tri 301 1096 302 1097 sw
rect 301 1072 302 1096
tri 304 1095 341 1132 ne
rect 341 1104 346 1132
tri 346 1104 372 1130 sw
rect 456 1114 465 1148
rect 456 1104 484 1114
rect 341 1095 425 1104
tri 341 1076 360 1095 ne
rect 360 1076 425 1095
rect 242 1050 302 1072
rect 424 1072 425 1076
rect 442 1072 484 1104
rect 424 1050 484 1072
rect 330 1034 347 1048
rect 379 1034 396 1048
tri 167 998 189 1020 se
rect 189 1013 204 1034
tri 189 998 204 1013 nw
rect 523 1013 538 1189
tri 538 1182 551 1195 nw
rect 624 1114 639 1342
tri 161 992 167 998 se
rect 167 992 176 998
rect 161 976 176 992
tri 176 985 189 998 nw
rect 330 990 347 1004
rect 379 990 396 1004
tri 523 998 538 1013 ne
tri 538 998 560 1020 sw
rect 161 940 176 948
rect 242 976 302 990
rect 257 966 302 976
rect 257 948 285 966
tri 161 925 176 940 ne
tri 176 925 198 947 sw
rect 242 938 285 948
rect 300 962 302 966
rect 424 976 484 990
tri 538 985 551 998 ne
rect 551 992 560 998
tri 560 992 566 998 sw
rect 424 966 469 976
rect 300 938 374 962
rect 242 934 374 938
tri 374 934 402 962 sw
rect 424 952 426 966
tri 424 950 426 952 ne
rect 438 948 469 966
rect 438 938 484 948
rect 551 977 566 992
tri 176 913 188 925 ne
rect 188 920 198 925
tri 198 920 203 925 sw
rect 87 574 102 802
rect 188 812 203 920
rect 242 878 270 934
tri 362 916 380 934 ne
rect 380 914 402 934
tri 402 914 422 934 sw
tri 438 920 456 938 ne
rect 261 844 270 878
rect 304 905 346 906
rect 304 871 309 905
rect 339 871 346 905
rect 304 862 346 871
rect 380 905 422 914
rect 380 871 387 905
rect 417 871 422 905
rect 380 866 422 871
rect 456 878 484 938
tri 529 925 551 947 se
rect 551 940 566 948
tri 551 925 566 940 nw
tri 523 919 529 925 se
rect 529 919 538 925
rect 242 834 270 844
tri 270 834 294 858 sw
rect 188 764 204 812
rect 242 802 284 834
tri 301 826 302 827 sw
rect 301 802 302 826
tri 304 825 341 862 ne
rect 341 834 346 862
tri 346 834 372 860 sw
rect 456 844 465 878
rect 456 834 484 844
rect 341 825 425 834
tri 341 806 360 825 ne
rect 360 806 425 825
rect 242 780 302 802
rect 424 802 425 806
rect 442 802 484 834
rect 424 780 484 802
rect 330 764 347 778
rect 379 764 396 778
tri 167 728 189 750 se
rect 189 743 204 764
tri 189 728 204 743 nw
rect 523 743 538 919
tri 538 912 551 925 nw
rect 624 844 639 1072
tri 161 722 167 728 se
rect 167 722 176 728
rect 161 706 176 722
tri 176 715 189 728 nw
rect 330 720 347 734
rect 379 720 396 734
tri 523 728 538 743 ne
tri 538 728 560 750 sw
rect 161 670 176 678
rect 242 706 302 720
rect 257 696 302 706
rect 257 678 285 696
tri 161 655 176 670 ne
tri 176 655 198 677 sw
rect 242 668 285 678
rect 300 692 302 696
rect 424 706 484 720
tri 538 715 551 728 ne
rect 551 722 560 728
tri 560 722 566 728 sw
rect 424 696 469 706
rect 300 668 374 692
rect 242 664 374 668
tri 374 664 402 692 sw
rect 424 682 426 696
tri 424 680 426 682 ne
rect 438 678 469 696
rect 438 668 484 678
rect 551 707 566 722
tri 176 643 188 655 ne
rect 188 650 198 655
tri 198 650 203 655 sw
rect 87 304 102 532
rect 188 494 203 650
rect 242 608 270 664
tri 362 646 380 664 ne
rect 380 644 402 664
tri 402 644 422 664 sw
tri 438 650 456 668 ne
rect 261 574 270 608
rect 304 635 346 636
rect 304 601 309 635
rect 339 601 346 635
rect 304 592 346 601
rect 380 635 422 644
rect 380 601 387 635
rect 417 601 422 635
rect 380 596 422 601
rect 456 608 484 668
tri 529 655 551 677 se
rect 551 670 566 678
tri 551 655 566 670 nw
tri 523 649 529 655 se
rect 529 649 538 655
rect 242 564 270 574
tri 270 564 294 588 sw
rect 242 532 284 564
tri 301 556 302 557 sw
rect 301 532 302 556
tri 304 555 341 592 ne
rect 341 564 346 592
tri 346 564 372 590 sw
rect 456 574 465 608
rect 456 564 484 574
rect 341 555 425 564
tri 341 536 360 555 ne
rect 360 536 425 555
rect 242 510 302 532
rect 424 532 425 536
rect 442 532 484 564
rect 424 510 484 532
rect 330 494 347 508
rect 379 494 396 508
tri 167 458 189 480 se
rect 189 473 204 494
tri 189 458 204 473 nw
rect 523 473 538 649
tri 538 642 551 655 nw
rect 624 574 639 802
tri 161 452 167 458 se
rect 167 452 176 458
rect 161 436 176 452
tri 176 445 189 458 nw
rect 330 450 347 464
rect 379 450 396 464
tri 523 458 538 473 ne
tri 538 458 560 480 sw
rect 161 400 176 408
rect 242 436 302 450
rect 257 426 302 436
rect 257 408 285 426
tri 161 385 176 400 ne
tri 176 385 198 407 sw
rect 242 398 285 408
rect 300 422 302 426
rect 424 436 484 450
tri 538 445 551 458 ne
rect 551 452 560 458
tri 560 452 566 458 sw
rect 424 426 469 436
rect 300 398 374 422
rect 242 394 374 398
tri 374 394 402 422 sw
rect 424 412 426 426
tri 424 410 426 412 ne
rect 438 408 469 426
rect 438 398 484 408
rect 551 437 566 452
tri 176 373 188 385 ne
rect 188 380 198 385
tri 198 380 203 385 sw
rect 87 34 102 262
rect 188 272 203 380
rect 242 338 270 394
tri 362 376 380 394 ne
rect 380 374 402 394
tri 402 374 422 394 sw
tri 438 380 456 398 ne
rect 261 304 270 338
rect 304 365 346 366
rect 304 331 309 365
rect 339 331 346 365
rect 304 322 346 331
rect 380 365 422 374
rect 380 331 387 365
rect 417 331 422 365
rect 380 326 422 331
rect 456 338 484 398
tri 529 385 551 407 se
rect 551 400 566 408
tri 551 385 566 400 nw
tri 523 379 529 385 se
rect 529 379 538 385
rect 242 294 270 304
tri 270 294 294 318 sw
rect 188 224 204 272
rect 242 262 284 294
tri 301 286 302 287 sw
rect 301 262 302 286
tri 304 285 341 322 ne
rect 341 294 346 322
tri 346 294 372 320 sw
rect 456 304 465 338
rect 456 294 484 304
rect 341 285 425 294
tri 341 266 360 285 ne
rect 360 266 425 285
rect 242 240 302 262
rect 424 262 425 266
rect 442 262 484 294
rect 424 240 484 262
rect 330 224 347 238
rect 379 224 396 238
tri 167 188 189 210 se
rect 189 203 204 224
tri 189 188 204 203 nw
rect 523 203 538 379
tri 538 372 551 385 nw
rect 624 304 639 532
tri 161 182 167 188 se
rect 167 182 176 188
rect 161 166 176 182
tri 176 175 189 188 nw
rect 330 180 347 194
rect 379 180 396 194
tri 523 188 538 203 ne
tri 538 188 560 210 sw
rect 161 130 176 138
rect 242 166 302 180
rect 257 156 302 166
rect 257 138 285 156
tri 161 115 176 130 ne
tri 176 115 198 137 sw
rect 242 128 285 138
rect 300 152 302 156
rect 424 166 484 180
tri 538 175 551 188 ne
rect 551 182 560 188
tri 560 182 566 188 sw
rect 424 156 469 166
rect 300 128 374 152
rect 242 124 374 128
tri 374 124 402 152 sw
rect 424 142 426 156
tri 424 140 426 142 ne
rect 438 138 469 156
rect 438 128 484 138
rect 551 167 566 182
tri 176 103 188 115 ne
rect 188 110 198 115
tri 198 110 203 115 sw
rect 87 -236 102 -8
rect 188 -46 203 110
rect 242 68 270 124
tri 362 106 380 124 ne
rect 380 104 402 124
tri 402 104 422 124 sw
tri 438 110 456 128 ne
rect 261 34 270 68
rect 304 95 346 96
rect 304 61 309 95
rect 339 61 346 95
rect 304 52 346 61
rect 380 95 422 104
rect 380 61 387 95
rect 417 61 422 95
rect 380 56 422 61
rect 456 68 484 128
tri 529 115 551 137 se
rect 551 130 566 138
tri 551 115 566 130 nw
tri 523 109 529 115 se
rect 529 109 538 115
rect 242 24 270 34
tri 270 24 294 48 sw
rect 242 -8 284 24
tri 301 16 302 17 sw
rect 301 -8 302 16
tri 304 15 341 52 ne
rect 341 24 346 52
tri 346 24 372 50 sw
rect 456 34 465 68
rect 456 24 484 34
rect 341 15 425 24
tri 341 -4 360 15 ne
rect 360 -4 425 15
rect 242 -30 302 -8
rect 424 -8 425 -4
rect 442 -8 484 24
rect 424 -30 484 -8
rect 330 -46 347 -32
rect 379 -46 396 -32
tri 167 -82 189 -60 se
rect 189 -67 204 -46
tri 189 -82 204 -67 nw
rect 523 -67 538 109
tri 538 102 551 115 nw
rect 624 34 639 262
tri 161 -88 167 -82 se
rect 167 -88 176 -82
rect 161 -104 176 -88
tri 176 -95 189 -82 nw
rect 330 -90 347 -76
rect 379 -90 396 -76
tri 523 -82 538 -67 ne
tri 538 -82 560 -60 sw
rect 161 -140 176 -132
rect 242 -104 302 -90
rect 257 -114 302 -104
rect 257 -132 285 -114
tri 161 -155 176 -140 ne
tri 176 -155 198 -133 sw
rect 242 -142 285 -132
rect 300 -118 302 -114
rect 424 -104 484 -90
tri 538 -95 551 -82 ne
rect 551 -88 560 -82
tri 560 -88 566 -82 sw
rect 424 -114 469 -104
rect 300 -142 374 -118
rect 242 -146 374 -142
tri 374 -146 402 -118 sw
rect 424 -128 426 -114
tri 424 -130 426 -128 ne
rect 438 -132 469 -114
rect 438 -142 484 -132
rect 551 -103 566 -88
tri 176 -167 188 -155 ne
rect 188 -160 198 -155
tri 198 -160 203 -155 sw
rect 87 -506 102 -278
rect 188 -268 203 -160
rect 242 -202 270 -146
tri 362 -164 380 -146 ne
rect 380 -166 402 -146
tri 402 -166 422 -146 sw
tri 438 -160 456 -142 ne
rect 261 -236 270 -202
rect 304 -175 346 -174
rect 304 -209 309 -175
rect 339 -209 346 -175
rect 304 -218 346 -209
rect 380 -175 422 -166
rect 380 -209 387 -175
rect 417 -209 422 -175
rect 380 -214 422 -209
rect 456 -202 484 -142
tri 529 -155 551 -133 se
rect 551 -140 566 -132
tri 551 -155 566 -140 nw
tri 523 -161 529 -155 se
rect 529 -161 538 -155
rect 242 -246 270 -236
tri 270 -246 294 -222 sw
rect 188 -316 204 -268
rect 242 -278 284 -246
tri 301 -254 302 -253 sw
rect 301 -278 302 -254
tri 304 -255 341 -218 ne
rect 341 -246 346 -218
tri 346 -246 372 -220 sw
rect 456 -236 465 -202
rect 456 -246 484 -236
rect 341 -255 425 -246
tri 341 -274 360 -255 ne
rect 360 -274 425 -255
rect 242 -300 302 -278
rect 424 -278 425 -274
rect 442 -278 484 -246
rect 424 -300 484 -278
rect 330 -316 347 -302
rect 379 -316 396 -302
tri 167 -352 189 -330 se
rect 189 -337 204 -316
tri 189 -352 204 -337 nw
rect 523 -337 538 -161
tri 538 -168 551 -155 nw
rect 624 -236 639 -8
tri 161 -358 167 -352 se
rect 167 -358 176 -352
rect 161 -374 176 -358
tri 176 -365 189 -352 nw
rect 330 -360 347 -346
rect 379 -360 396 -346
tri 523 -352 538 -337 ne
tri 538 -352 560 -330 sw
rect 161 -410 176 -402
rect 242 -374 302 -360
rect 257 -384 302 -374
rect 257 -402 285 -384
tri 161 -425 176 -410 ne
tri 176 -425 198 -403 sw
rect 242 -412 285 -402
rect 300 -388 302 -384
rect 424 -374 484 -360
tri 538 -365 551 -352 ne
rect 551 -358 560 -352
tri 560 -358 566 -352 sw
rect 424 -384 469 -374
rect 300 -412 374 -388
rect 242 -416 374 -412
tri 374 -416 402 -388 sw
rect 424 -398 426 -384
tri 424 -400 426 -398 ne
rect 438 -402 469 -384
rect 438 -412 484 -402
rect 551 -373 566 -358
tri 176 -437 188 -425 ne
rect 188 -430 198 -425
tri 198 -430 203 -425 sw
rect 87 -776 102 -548
rect 188 -586 203 -430
rect 242 -472 270 -416
tri 362 -434 380 -416 ne
rect 380 -436 402 -416
tri 402 -436 422 -416 sw
tri 438 -430 456 -412 ne
rect 261 -506 270 -472
rect 304 -445 346 -444
rect 304 -479 309 -445
rect 339 -479 346 -445
rect 304 -488 346 -479
rect 380 -445 422 -436
rect 380 -479 387 -445
rect 417 -479 422 -445
rect 380 -484 422 -479
rect 456 -472 484 -412
tri 529 -425 551 -403 se
rect 551 -410 566 -402
tri 551 -425 566 -410 nw
tri 523 -431 529 -425 se
rect 529 -431 538 -425
rect 242 -516 270 -506
tri 270 -516 294 -492 sw
rect 242 -548 284 -516
tri 301 -524 302 -523 sw
rect 301 -548 302 -524
tri 304 -525 341 -488 ne
rect 341 -516 346 -488
tri 346 -516 372 -490 sw
rect 456 -506 465 -472
rect 456 -516 484 -506
rect 341 -525 425 -516
tri 341 -544 360 -525 ne
rect 360 -544 425 -525
rect 242 -570 302 -548
rect 424 -548 425 -544
rect 442 -548 484 -516
rect 424 -570 484 -548
rect 330 -586 347 -572
rect 379 -586 396 -572
tri 167 -622 189 -600 se
rect 189 -607 204 -586
tri 189 -622 204 -607 nw
rect 523 -607 538 -431
tri 538 -438 551 -425 nw
rect 624 -506 639 -278
tri 161 -628 167 -622 se
rect 167 -628 176 -622
rect 161 -644 176 -628
tri 176 -635 189 -622 nw
rect 330 -630 347 -616
rect 379 -630 396 -616
tri 523 -622 538 -607 ne
tri 538 -622 560 -600 sw
rect 161 -680 176 -672
rect 242 -644 302 -630
rect 257 -654 302 -644
rect 257 -672 285 -654
tri 161 -695 176 -680 ne
tri 176 -695 198 -673 sw
rect 242 -682 285 -672
rect 300 -658 302 -654
rect 424 -644 484 -630
tri 538 -635 551 -622 ne
rect 551 -628 560 -622
tri 560 -628 566 -622 sw
rect 424 -654 469 -644
rect 300 -682 374 -658
rect 242 -686 374 -682
tri 374 -686 402 -658 sw
rect 424 -668 426 -654
tri 424 -670 426 -668 ne
rect 438 -672 469 -654
rect 438 -682 484 -672
rect 551 -643 566 -628
tri 176 -707 188 -695 ne
rect 188 -700 198 -695
tri 198 -700 203 -695 sw
rect 87 -1046 102 -818
rect 188 -808 203 -700
rect 242 -742 270 -686
tri 362 -704 380 -686 ne
rect 380 -706 402 -686
tri 402 -706 422 -686 sw
tri 438 -700 456 -682 ne
rect 261 -776 270 -742
rect 304 -715 346 -714
rect 304 -749 309 -715
rect 339 -749 346 -715
rect 304 -758 346 -749
rect 380 -715 422 -706
rect 380 -749 387 -715
rect 417 -749 422 -715
rect 380 -754 422 -749
rect 456 -742 484 -682
tri 529 -695 551 -673 se
rect 551 -680 566 -672
tri 551 -695 566 -680 nw
tri 523 -701 529 -695 se
rect 529 -701 538 -695
rect 242 -786 270 -776
tri 270 -786 294 -762 sw
rect 188 -856 204 -808
rect 242 -818 284 -786
tri 301 -794 302 -793 sw
rect 301 -818 302 -794
tri 304 -795 341 -758 ne
rect 341 -786 346 -758
tri 346 -786 372 -760 sw
rect 456 -776 465 -742
rect 456 -786 484 -776
rect 341 -795 425 -786
tri 341 -814 360 -795 ne
rect 360 -814 425 -795
rect 242 -840 302 -818
rect 424 -818 425 -814
rect 442 -818 484 -786
rect 424 -840 484 -818
rect 330 -856 347 -842
rect 379 -856 396 -842
tri 167 -892 189 -870 se
rect 189 -877 204 -856
tri 189 -892 204 -877 nw
rect 523 -877 538 -701
tri 538 -708 551 -695 nw
rect 624 -776 639 -548
tri 161 -898 167 -892 se
rect 167 -898 176 -892
rect 161 -914 176 -898
tri 176 -905 189 -892 nw
rect 330 -900 347 -886
rect 379 -900 396 -886
tri 523 -892 538 -877 ne
tri 538 -892 560 -870 sw
rect 161 -950 176 -942
rect 242 -914 302 -900
rect 257 -924 302 -914
rect 257 -942 285 -924
tri 161 -965 176 -950 ne
tri 176 -965 198 -943 sw
rect 242 -952 285 -942
rect 300 -928 302 -924
rect 424 -914 484 -900
tri 538 -905 551 -892 ne
rect 551 -898 560 -892
tri 560 -898 566 -892 sw
rect 424 -924 469 -914
rect 300 -952 374 -928
rect 242 -956 374 -952
tri 374 -956 402 -928 sw
rect 424 -938 426 -924
tri 424 -940 426 -938 ne
rect 438 -942 469 -924
rect 438 -952 484 -942
rect 551 -913 566 -898
tri 176 -977 188 -965 ne
rect 188 -970 198 -965
tri 198 -970 203 -965 sw
rect 87 -1316 102 -1088
rect 188 -1126 203 -970
rect 242 -1012 270 -956
tri 362 -974 380 -956 ne
rect 380 -976 402 -956
tri 402 -976 422 -956 sw
tri 438 -970 456 -952 ne
rect 261 -1046 270 -1012
rect 304 -985 346 -984
rect 304 -1019 309 -985
rect 339 -1019 346 -985
rect 304 -1028 346 -1019
rect 380 -985 422 -976
rect 380 -1019 387 -985
rect 417 -1019 422 -985
rect 380 -1024 422 -1019
rect 456 -1012 484 -952
tri 529 -965 551 -943 se
rect 551 -950 566 -942
tri 551 -965 566 -950 nw
tri 523 -971 529 -965 se
rect 529 -971 538 -965
rect 242 -1056 270 -1046
tri 270 -1056 294 -1032 sw
rect 242 -1088 284 -1056
tri 301 -1064 302 -1063 sw
rect 301 -1088 302 -1064
tri 304 -1065 341 -1028 ne
rect 341 -1056 346 -1028
tri 346 -1056 372 -1030 sw
rect 456 -1046 465 -1012
rect 456 -1056 484 -1046
rect 341 -1065 425 -1056
tri 341 -1084 360 -1065 ne
rect 360 -1084 425 -1065
rect 242 -1110 302 -1088
rect 424 -1088 425 -1084
rect 442 -1088 484 -1056
rect 424 -1110 484 -1088
rect 330 -1126 347 -1112
rect 379 -1126 396 -1112
tri 167 -1162 189 -1140 se
rect 189 -1147 204 -1126
tri 189 -1162 204 -1147 nw
rect 523 -1147 538 -971
tri 538 -978 551 -965 nw
rect 624 -1046 639 -818
tri 161 -1168 167 -1162 se
rect 167 -1168 176 -1162
rect 161 -1184 176 -1168
tri 176 -1175 189 -1162 nw
rect 330 -1170 347 -1156
rect 379 -1170 396 -1156
tri 523 -1162 538 -1147 ne
tri 538 -1162 560 -1140 sw
rect 161 -1220 176 -1212
rect 242 -1184 302 -1170
rect 257 -1194 302 -1184
rect 257 -1212 285 -1194
tri 161 -1235 176 -1220 ne
tri 176 -1235 198 -1213 sw
rect 242 -1222 285 -1212
rect 300 -1198 302 -1194
rect 424 -1184 484 -1170
tri 538 -1175 551 -1162 ne
rect 551 -1168 560 -1162
tri 560 -1168 566 -1162 sw
rect 424 -1194 469 -1184
rect 300 -1222 374 -1198
rect 242 -1226 374 -1222
tri 374 -1226 402 -1198 sw
rect 424 -1208 426 -1194
tri 424 -1210 426 -1208 ne
rect 438 -1212 469 -1194
rect 438 -1222 484 -1212
rect 551 -1183 566 -1168
tri 176 -1247 188 -1235 ne
rect 188 -1240 198 -1235
tri 198 -1240 203 -1235 sw
rect 87 -1586 102 -1358
rect 188 -1348 203 -1240
rect 242 -1282 270 -1226
tri 362 -1244 380 -1226 ne
rect 380 -1246 402 -1226
tri 402 -1246 422 -1226 sw
tri 438 -1240 456 -1222 ne
rect 261 -1316 270 -1282
rect 304 -1255 346 -1254
rect 304 -1289 309 -1255
rect 339 -1289 346 -1255
rect 304 -1298 346 -1289
rect 380 -1255 422 -1246
rect 380 -1289 387 -1255
rect 417 -1289 422 -1255
rect 380 -1294 422 -1289
rect 456 -1282 484 -1222
tri 529 -1235 551 -1213 se
rect 551 -1220 566 -1212
tri 551 -1235 566 -1220 nw
tri 523 -1241 529 -1235 se
rect 529 -1241 538 -1235
rect 242 -1326 270 -1316
tri 270 -1326 294 -1302 sw
rect 188 -1396 204 -1348
rect 242 -1358 284 -1326
tri 301 -1334 302 -1333 sw
rect 301 -1358 302 -1334
tri 304 -1335 341 -1298 ne
rect 341 -1326 346 -1298
tri 346 -1326 372 -1300 sw
rect 456 -1316 465 -1282
rect 456 -1326 484 -1316
rect 341 -1335 425 -1326
tri 341 -1354 360 -1335 ne
rect 360 -1354 425 -1335
rect 242 -1380 302 -1358
rect 424 -1358 425 -1354
rect 442 -1358 484 -1326
rect 424 -1380 484 -1358
rect 330 -1396 347 -1382
rect 379 -1396 396 -1382
tri 167 -1432 189 -1410 se
rect 189 -1417 204 -1396
tri 189 -1432 204 -1417 nw
rect 523 -1417 538 -1241
tri 538 -1248 551 -1235 nw
rect 624 -1316 639 -1088
tri 161 -1438 167 -1432 se
rect 167 -1438 176 -1432
rect 161 -1454 176 -1438
tri 176 -1445 189 -1432 nw
rect 330 -1440 347 -1426
rect 379 -1440 396 -1426
tri 523 -1432 538 -1417 ne
tri 538 -1432 560 -1410 sw
rect 161 -1490 176 -1482
rect 242 -1454 302 -1440
rect 257 -1464 302 -1454
rect 257 -1482 285 -1464
tri 161 -1505 176 -1490 ne
tri 176 -1505 198 -1483 sw
rect 242 -1492 285 -1482
rect 300 -1468 302 -1464
rect 424 -1454 484 -1440
tri 538 -1445 551 -1432 ne
rect 551 -1438 560 -1432
tri 560 -1438 566 -1432 sw
rect 424 -1464 469 -1454
rect 300 -1492 374 -1468
rect 242 -1496 374 -1492
tri 374 -1496 402 -1468 sw
rect 424 -1478 426 -1464
tri 424 -1480 426 -1478 ne
rect 438 -1482 469 -1464
rect 438 -1492 484 -1482
rect 551 -1453 566 -1438
tri 176 -1517 188 -1505 ne
rect 188 -1510 198 -1505
tri 198 -1510 203 -1505 sw
rect 87 -1856 102 -1628
rect 188 -1666 203 -1510
rect 242 -1552 270 -1496
tri 362 -1514 380 -1496 ne
rect 380 -1516 402 -1496
tri 402 -1516 422 -1496 sw
tri 438 -1510 456 -1492 ne
rect 261 -1586 270 -1552
rect 304 -1525 346 -1524
rect 304 -1559 309 -1525
rect 339 -1559 346 -1525
rect 304 -1568 346 -1559
rect 380 -1525 422 -1516
rect 380 -1559 387 -1525
rect 417 -1559 422 -1525
rect 380 -1564 422 -1559
rect 456 -1552 484 -1492
tri 529 -1505 551 -1483 se
rect 551 -1490 566 -1482
tri 551 -1505 566 -1490 nw
tri 523 -1511 529 -1505 se
rect 529 -1511 538 -1505
rect 242 -1596 270 -1586
tri 270 -1596 294 -1572 sw
rect 242 -1628 284 -1596
tri 301 -1604 302 -1603 sw
rect 301 -1628 302 -1604
tri 304 -1605 341 -1568 ne
rect 341 -1596 346 -1568
tri 346 -1596 372 -1570 sw
rect 456 -1586 465 -1552
rect 456 -1596 484 -1586
rect 341 -1605 425 -1596
tri 341 -1624 360 -1605 ne
rect 360 -1624 425 -1605
rect 242 -1650 302 -1628
rect 424 -1628 425 -1624
rect 442 -1628 484 -1596
rect 424 -1650 484 -1628
rect 330 -1666 347 -1652
rect 379 -1666 396 -1652
tri 167 -1702 189 -1680 se
rect 189 -1687 204 -1666
tri 189 -1702 204 -1687 nw
rect 523 -1687 538 -1511
tri 538 -1518 551 -1505 nw
rect 624 -1586 639 -1358
tri 161 -1708 167 -1702 se
rect 167 -1708 176 -1702
rect 161 -1724 176 -1708
tri 176 -1715 189 -1702 nw
rect 330 -1710 347 -1696
rect 379 -1710 396 -1696
tri 523 -1702 538 -1687 ne
tri 538 -1702 560 -1680 sw
rect 161 -1760 176 -1752
rect 242 -1724 302 -1710
rect 257 -1734 302 -1724
rect 257 -1752 285 -1734
tri 161 -1775 176 -1760 ne
tri 176 -1775 198 -1753 sw
rect 242 -1762 285 -1752
rect 300 -1738 302 -1734
rect 424 -1724 484 -1710
tri 538 -1715 551 -1702 ne
rect 551 -1708 560 -1702
tri 560 -1708 566 -1702 sw
rect 424 -1734 469 -1724
rect 300 -1762 374 -1738
rect 242 -1766 374 -1762
tri 374 -1766 402 -1738 sw
rect 424 -1748 426 -1734
tri 424 -1750 426 -1748 ne
rect 438 -1752 469 -1734
rect 438 -1762 484 -1752
rect 551 -1723 566 -1708
tri 176 -1787 188 -1775 ne
rect 188 -1780 198 -1775
tri 198 -1780 203 -1775 sw
rect 87 -2126 102 -1898
rect 188 -1888 203 -1780
rect 242 -1822 270 -1766
tri 362 -1784 380 -1766 ne
rect 380 -1786 402 -1766
tri 402 -1786 422 -1766 sw
tri 438 -1780 456 -1762 ne
rect 261 -1856 270 -1822
rect 304 -1795 346 -1794
rect 304 -1829 309 -1795
rect 339 -1829 346 -1795
rect 304 -1838 346 -1829
rect 380 -1795 422 -1786
rect 380 -1829 387 -1795
rect 417 -1829 422 -1795
rect 380 -1834 422 -1829
rect 456 -1822 484 -1762
tri 529 -1775 551 -1753 se
rect 551 -1760 566 -1752
tri 551 -1775 566 -1760 nw
tri 523 -1781 529 -1775 se
rect 529 -1781 538 -1775
rect 242 -1866 270 -1856
tri 270 -1866 294 -1842 sw
rect 188 -1936 204 -1888
rect 242 -1898 284 -1866
tri 301 -1874 302 -1873 sw
rect 301 -1898 302 -1874
tri 304 -1875 341 -1838 ne
rect 341 -1866 346 -1838
tri 346 -1866 372 -1840 sw
rect 456 -1856 465 -1822
rect 456 -1866 484 -1856
rect 341 -1875 425 -1866
tri 341 -1894 360 -1875 ne
rect 360 -1894 425 -1875
rect 242 -1920 302 -1898
rect 424 -1898 425 -1894
rect 442 -1898 484 -1866
rect 424 -1920 484 -1898
rect 330 -1936 347 -1922
rect 379 -1936 396 -1922
tri 167 -1972 189 -1950 se
rect 189 -1957 204 -1936
tri 189 -1972 204 -1957 nw
rect 523 -1957 538 -1781
tri 538 -1788 551 -1775 nw
rect 624 -1856 639 -1628
tri 161 -1978 167 -1972 se
rect 167 -1978 176 -1972
rect 161 -1994 176 -1978
tri 176 -1985 189 -1972 nw
rect 330 -1980 347 -1966
rect 379 -1980 396 -1966
tri 523 -1972 538 -1957 ne
tri 538 -1972 560 -1950 sw
rect 161 -2030 176 -2022
rect 242 -1994 302 -1980
rect 257 -2004 302 -1994
rect 257 -2022 285 -2004
tri 161 -2045 176 -2030 ne
tri 176 -2045 198 -2023 sw
rect 242 -2032 285 -2022
rect 300 -2008 302 -2004
rect 424 -1994 484 -1980
tri 538 -1985 551 -1972 ne
rect 551 -1978 560 -1972
tri 560 -1978 566 -1972 sw
rect 424 -2004 469 -1994
rect 300 -2032 374 -2008
rect 242 -2036 374 -2032
tri 374 -2036 402 -2008 sw
rect 424 -2018 426 -2004
tri 424 -2020 426 -2018 ne
rect 438 -2022 469 -2004
rect 438 -2032 484 -2022
rect 551 -1993 566 -1978
tri 176 -2057 188 -2045 ne
rect 188 -2050 198 -2045
tri 198 -2050 203 -2045 sw
rect 87 -2396 102 -2168
rect 188 -2206 203 -2050
rect 242 -2092 270 -2036
tri 362 -2054 380 -2036 ne
rect 380 -2056 402 -2036
tri 402 -2056 422 -2036 sw
tri 438 -2050 456 -2032 ne
rect 261 -2126 270 -2092
rect 304 -2065 346 -2064
rect 304 -2099 309 -2065
rect 339 -2099 346 -2065
rect 304 -2108 346 -2099
rect 380 -2065 422 -2056
rect 380 -2099 387 -2065
rect 417 -2099 422 -2065
rect 380 -2104 422 -2099
rect 456 -2092 484 -2032
tri 529 -2045 551 -2023 se
rect 551 -2030 566 -2022
tri 551 -2045 566 -2030 nw
tri 523 -2051 529 -2045 se
rect 529 -2051 538 -2045
rect 242 -2136 270 -2126
tri 270 -2136 294 -2112 sw
rect 242 -2168 284 -2136
tri 301 -2144 302 -2143 sw
rect 301 -2168 302 -2144
tri 304 -2145 341 -2108 ne
rect 341 -2136 346 -2108
tri 346 -2136 372 -2110 sw
rect 456 -2126 465 -2092
rect 456 -2136 484 -2126
rect 341 -2145 425 -2136
tri 341 -2164 360 -2145 ne
rect 360 -2164 425 -2145
rect 242 -2190 302 -2168
rect 424 -2168 425 -2164
rect 442 -2168 484 -2136
rect 424 -2190 484 -2168
rect 330 -2206 347 -2192
rect 379 -2206 396 -2192
tri 167 -2242 189 -2220 se
rect 189 -2227 204 -2206
tri 189 -2242 204 -2227 nw
rect 523 -2227 538 -2051
tri 538 -2058 551 -2045 nw
rect 624 -2126 639 -1898
tri 161 -2248 167 -2242 se
rect 167 -2248 176 -2242
rect 161 -2264 176 -2248
tri 176 -2255 189 -2242 nw
rect 330 -2250 347 -2236
rect 379 -2250 396 -2236
tri 523 -2242 538 -2227 ne
tri 538 -2242 560 -2220 sw
rect 161 -2300 176 -2292
rect 242 -2264 302 -2250
rect 257 -2274 302 -2264
rect 257 -2292 285 -2274
tri 161 -2315 176 -2300 ne
tri 176 -2315 198 -2293 sw
rect 242 -2302 285 -2292
rect 300 -2278 302 -2274
rect 424 -2264 484 -2250
tri 538 -2255 551 -2242 ne
rect 551 -2248 560 -2242
tri 560 -2248 566 -2242 sw
rect 424 -2274 469 -2264
rect 300 -2302 374 -2278
rect 242 -2306 374 -2302
tri 374 -2306 402 -2278 sw
rect 424 -2288 426 -2274
tri 424 -2290 426 -2288 ne
rect 438 -2292 469 -2274
rect 438 -2302 484 -2292
rect 551 -2263 566 -2248
tri 176 -2327 188 -2315 ne
rect 188 -2320 198 -2315
tri 198 -2320 203 -2315 sw
rect 87 -2524 102 -2438
rect 188 -2476 203 -2320
rect 242 -2362 270 -2306
tri 362 -2324 380 -2306 ne
rect 380 -2326 402 -2306
tri 402 -2326 422 -2306 sw
tri 438 -2320 456 -2302 ne
rect 261 -2396 270 -2362
rect 304 -2335 346 -2334
rect 304 -2369 309 -2335
rect 339 -2369 346 -2335
rect 304 -2378 346 -2369
rect 380 -2335 422 -2326
rect 380 -2369 387 -2335
rect 417 -2369 422 -2335
rect 380 -2374 422 -2369
rect 456 -2362 484 -2302
tri 529 -2315 551 -2293 se
rect 551 -2300 566 -2292
tri 551 -2315 566 -2300 nw
tri 523 -2321 529 -2315 se
rect 529 -2321 538 -2315
rect 242 -2406 270 -2396
tri 270 -2406 294 -2382 sw
rect 242 -2438 284 -2406
tri 301 -2414 302 -2413 sw
rect 301 -2438 302 -2414
tri 304 -2415 341 -2378 ne
rect 341 -2406 346 -2378
tri 346 -2406 372 -2380 sw
rect 456 -2396 465 -2362
rect 456 -2406 484 -2396
rect 341 -2415 425 -2406
tri 341 -2434 360 -2415 ne
rect 360 -2434 425 -2415
rect 242 -2460 302 -2438
rect 424 -2438 425 -2434
rect 442 -2438 484 -2406
rect 424 -2460 484 -2438
rect 330 -2476 347 -2462
rect 379 -2476 396 -2462
rect 523 -2476 538 -2321
tri 538 -2328 551 -2315 nw
rect 624 -2396 639 -2168
rect 624 -2524 639 -2438
rect 667 1654 682 1892
tri 747 1808 769 1830 se
rect 769 1823 784 1892
tri 769 1808 784 1823 nw
rect 1103 1823 1118 1892
tri 741 1802 747 1808 se
rect 747 1802 756 1808
rect 741 1786 756 1802
tri 756 1795 769 1808 nw
rect 910 1800 927 1814
rect 959 1800 976 1814
tri 1103 1808 1118 1823 ne
tri 1118 1808 1140 1830 sw
rect 741 1750 756 1758
rect 822 1786 882 1800
rect 837 1776 882 1786
rect 837 1758 865 1776
tri 741 1735 756 1750 ne
tri 756 1735 778 1757 sw
rect 822 1748 865 1758
rect 880 1772 882 1776
rect 1004 1786 1064 1800
tri 1118 1795 1131 1808 ne
rect 1131 1802 1140 1808
tri 1140 1802 1146 1808 sw
rect 1004 1776 1049 1786
rect 880 1748 954 1772
rect 822 1744 954 1748
tri 954 1744 982 1772 sw
rect 1004 1762 1006 1776
tri 1004 1760 1006 1762 ne
rect 1018 1758 1049 1776
rect 1018 1748 1064 1758
rect 1131 1787 1146 1802
tri 756 1723 768 1735 ne
rect 768 1730 778 1735
tri 778 1730 783 1735 sw
rect 667 1384 682 1612
rect 768 1574 783 1730
rect 822 1688 850 1744
tri 942 1726 960 1744 ne
rect 960 1724 982 1744
tri 982 1724 1002 1744 sw
tri 1018 1730 1036 1748 ne
rect 841 1654 850 1688
rect 884 1715 926 1716
rect 884 1681 889 1715
rect 919 1681 926 1715
rect 884 1672 926 1681
rect 960 1715 1002 1724
rect 960 1681 967 1715
rect 997 1681 1002 1715
rect 960 1676 1002 1681
rect 1036 1688 1064 1748
tri 1109 1735 1131 1757 se
rect 1131 1750 1146 1758
tri 1131 1735 1146 1750 nw
tri 1103 1729 1109 1735 se
rect 1109 1729 1118 1735
rect 822 1644 850 1654
tri 850 1644 874 1668 sw
rect 822 1612 864 1644
tri 881 1636 882 1637 sw
rect 881 1612 882 1636
tri 884 1635 921 1672 ne
rect 921 1644 926 1672
tri 926 1644 952 1670 sw
rect 1036 1654 1045 1688
rect 1036 1644 1064 1654
rect 921 1635 1005 1644
tri 921 1616 940 1635 ne
rect 940 1616 1005 1635
rect 822 1590 882 1612
rect 1004 1612 1005 1616
rect 1022 1612 1064 1644
rect 1004 1590 1064 1612
rect 910 1574 927 1588
rect 959 1574 976 1588
tri 747 1538 769 1560 se
rect 769 1553 784 1574
tri 769 1538 784 1553 nw
rect 1103 1553 1118 1729
tri 1118 1722 1131 1735 nw
rect 1204 1654 1219 1892
tri 741 1532 747 1538 se
rect 747 1532 756 1538
rect 741 1516 756 1532
tri 756 1525 769 1538 nw
rect 910 1530 927 1544
rect 959 1530 976 1544
tri 1103 1538 1118 1553 ne
tri 1118 1538 1140 1560 sw
rect 741 1480 756 1488
rect 822 1516 882 1530
rect 837 1506 882 1516
rect 837 1488 865 1506
tri 741 1465 756 1480 ne
tri 756 1465 778 1487 sw
rect 822 1478 865 1488
rect 880 1502 882 1506
rect 1004 1516 1064 1530
tri 1118 1525 1131 1538 ne
rect 1131 1532 1140 1538
tri 1140 1532 1146 1538 sw
rect 1004 1506 1049 1516
rect 880 1478 954 1502
rect 822 1474 954 1478
tri 954 1474 982 1502 sw
rect 1004 1492 1006 1506
tri 1004 1490 1006 1492 ne
rect 1018 1488 1049 1506
rect 1018 1478 1064 1488
rect 1131 1517 1146 1532
tri 756 1453 768 1465 ne
rect 768 1460 778 1465
tri 778 1460 783 1465 sw
rect 667 1114 682 1342
rect 768 1352 783 1460
rect 822 1418 850 1474
tri 942 1456 960 1474 ne
rect 960 1454 982 1474
tri 982 1454 1002 1474 sw
tri 1018 1460 1036 1478 ne
rect 841 1384 850 1418
rect 884 1445 926 1446
rect 884 1411 889 1445
rect 919 1411 926 1445
rect 884 1402 926 1411
rect 960 1445 1002 1454
rect 960 1411 967 1445
rect 997 1411 1002 1445
rect 960 1406 1002 1411
rect 1036 1418 1064 1478
tri 1109 1465 1131 1487 se
rect 1131 1480 1146 1488
tri 1131 1465 1146 1480 nw
tri 1103 1459 1109 1465 se
rect 1109 1459 1118 1465
rect 822 1374 850 1384
tri 850 1374 874 1398 sw
rect 768 1304 784 1352
rect 822 1342 864 1374
tri 881 1366 882 1367 sw
rect 881 1342 882 1366
tri 884 1365 921 1402 ne
rect 921 1374 926 1402
tri 926 1374 952 1400 sw
rect 1036 1384 1045 1418
rect 1036 1374 1064 1384
rect 921 1365 1005 1374
tri 921 1346 940 1365 ne
rect 940 1346 1005 1365
rect 822 1320 882 1342
rect 1004 1342 1005 1346
rect 1022 1342 1064 1374
rect 1004 1320 1064 1342
rect 910 1304 927 1318
rect 959 1304 976 1318
tri 747 1268 769 1290 se
rect 769 1283 784 1304
tri 769 1268 784 1283 nw
rect 1103 1283 1118 1459
tri 1118 1452 1131 1465 nw
rect 1204 1384 1219 1612
tri 741 1262 747 1268 se
rect 747 1262 756 1268
rect 741 1246 756 1262
tri 756 1255 769 1268 nw
rect 910 1260 927 1274
rect 959 1260 976 1274
tri 1103 1268 1118 1283 ne
tri 1118 1268 1140 1290 sw
rect 741 1210 756 1218
rect 822 1246 882 1260
rect 837 1236 882 1246
rect 837 1218 865 1236
tri 741 1195 756 1210 ne
tri 756 1195 778 1217 sw
rect 822 1208 865 1218
rect 880 1232 882 1236
rect 1004 1246 1064 1260
tri 1118 1255 1131 1268 ne
rect 1131 1262 1140 1268
tri 1140 1262 1146 1268 sw
rect 1004 1236 1049 1246
rect 880 1208 954 1232
rect 822 1204 954 1208
tri 954 1204 982 1232 sw
rect 1004 1222 1006 1236
tri 1004 1220 1006 1222 ne
rect 1018 1218 1049 1236
rect 1018 1208 1064 1218
rect 1131 1247 1146 1262
tri 756 1183 768 1195 ne
rect 768 1190 778 1195
tri 778 1190 783 1195 sw
rect 667 844 682 1072
rect 768 1034 783 1190
rect 822 1148 850 1204
tri 942 1186 960 1204 ne
rect 960 1184 982 1204
tri 982 1184 1002 1204 sw
tri 1018 1190 1036 1208 ne
rect 841 1114 850 1148
rect 884 1175 926 1176
rect 884 1141 889 1175
rect 919 1141 926 1175
rect 884 1132 926 1141
rect 960 1175 1002 1184
rect 960 1141 967 1175
rect 997 1141 1002 1175
rect 960 1136 1002 1141
rect 1036 1148 1064 1208
tri 1109 1195 1131 1217 se
rect 1131 1210 1146 1218
tri 1131 1195 1146 1210 nw
tri 1103 1189 1109 1195 se
rect 1109 1189 1118 1195
rect 822 1104 850 1114
tri 850 1104 874 1128 sw
rect 822 1072 864 1104
tri 881 1096 882 1097 sw
rect 881 1072 882 1096
tri 884 1095 921 1132 ne
rect 921 1104 926 1132
tri 926 1104 952 1130 sw
rect 1036 1114 1045 1148
rect 1036 1104 1064 1114
rect 921 1095 1005 1104
tri 921 1076 940 1095 ne
rect 940 1076 1005 1095
rect 822 1050 882 1072
rect 1004 1072 1005 1076
rect 1022 1072 1064 1104
rect 1004 1050 1064 1072
rect 910 1034 927 1048
rect 959 1034 976 1048
tri 747 998 769 1020 se
rect 769 1013 784 1034
tri 769 998 784 1013 nw
rect 1103 1013 1118 1189
tri 1118 1182 1131 1195 nw
rect 1204 1114 1219 1342
tri 741 992 747 998 se
rect 747 992 756 998
rect 741 976 756 992
tri 756 985 769 998 nw
rect 910 990 927 1004
rect 959 990 976 1004
tri 1103 998 1118 1013 ne
tri 1118 998 1140 1020 sw
rect 741 940 756 948
rect 822 976 882 990
rect 837 966 882 976
rect 837 948 865 966
tri 741 925 756 940 ne
tri 756 925 778 947 sw
rect 822 938 865 948
rect 880 962 882 966
rect 1004 976 1064 990
tri 1118 985 1131 998 ne
rect 1131 992 1140 998
tri 1140 992 1146 998 sw
rect 1004 966 1049 976
rect 880 938 954 962
rect 822 934 954 938
tri 954 934 982 962 sw
rect 1004 952 1006 966
tri 1004 950 1006 952 ne
rect 1018 948 1049 966
rect 1018 938 1064 948
rect 1131 977 1146 992
tri 756 913 768 925 ne
rect 768 920 778 925
tri 778 920 783 925 sw
rect 667 574 682 802
rect 768 812 783 920
rect 822 878 850 934
tri 942 916 960 934 ne
rect 960 914 982 934
tri 982 914 1002 934 sw
tri 1018 920 1036 938 ne
rect 841 844 850 878
rect 884 905 926 906
rect 884 871 889 905
rect 919 871 926 905
rect 884 862 926 871
rect 960 905 1002 914
rect 960 871 967 905
rect 997 871 1002 905
rect 960 866 1002 871
rect 1036 878 1064 938
tri 1109 925 1131 947 se
rect 1131 940 1146 948
tri 1131 925 1146 940 nw
tri 1103 919 1109 925 se
rect 1109 919 1118 925
rect 822 834 850 844
tri 850 834 874 858 sw
rect 768 764 784 812
rect 822 802 864 834
tri 881 826 882 827 sw
rect 881 802 882 826
tri 884 825 921 862 ne
rect 921 834 926 862
tri 926 834 952 860 sw
rect 1036 844 1045 878
rect 1036 834 1064 844
rect 921 825 1005 834
tri 921 806 940 825 ne
rect 940 806 1005 825
rect 822 780 882 802
rect 1004 802 1005 806
rect 1022 802 1064 834
rect 1004 780 1064 802
rect 910 764 927 778
rect 959 764 976 778
tri 747 728 769 750 se
rect 769 743 784 764
tri 769 728 784 743 nw
rect 1103 743 1118 919
tri 1118 912 1131 925 nw
rect 1204 844 1219 1072
tri 741 722 747 728 se
rect 747 722 756 728
rect 741 706 756 722
tri 756 715 769 728 nw
rect 910 720 927 734
rect 959 720 976 734
tri 1103 728 1118 743 ne
tri 1118 728 1140 750 sw
rect 741 670 756 678
rect 822 706 882 720
rect 837 696 882 706
rect 837 678 865 696
tri 741 655 756 670 ne
tri 756 655 778 677 sw
rect 822 668 865 678
rect 880 692 882 696
rect 1004 706 1064 720
tri 1118 715 1131 728 ne
rect 1131 722 1140 728
tri 1140 722 1146 728 sw
rect 1004 696 1049 706
rect 880 668 954 692
rect 822 664 954 668
tri 954 664 982 692 sw
rect 1004 682 1006 696
tri 1004 680 1006 682 ne
rect 1018 678 1049 696
rect 1018 668 1064 678
rect 1131 707 1146 722
tri 756 643 768 655 ne
rect 768 650 778 655
tri 778 650 783 655 sw
rect 667 304 682 532
rect 768 494 783 650
rect 822 608 850 664
tri 942 646 960 664 ne
rect 960 644 982 664
tri 982 644 1002 664 sw
tri 1018 650 1036 668 ne
rect 841 574 850 608
rect 884 635 926 636
rect 884 601 889 635
rect 919 601 926 635
rect 884 592 926 601
rect 960 635 1002 644
rect 960 601 967 635
rect 997 601 1002 635
rect 960 596 1002 601
rect 1036 608 1064 668
tri 1109 655 1131 677 se
rect 1131 670 1146 678
tri 1131 655 1146 670 nw
tri 1103 649 1109 655 se
rect 1109 649 1118 655
rect 822 564 850 574
tri 850 564 874 588 sw
rect 822 532 864 564
tri 881 556 882 557 sw
rect 881 532 882 556
tri 884 555 921 592 ne
rect 921 564 926 592
tri 926 564 952 590 sw
rect 1036 574 1045 608
rect 1036 564 1064 574
rect 921 555 1005 564
tri 921 536 940 555 ne
rect 940 536 1005 555
rect 822 510 882 532
rect 1004 532 1005 536
rect 1022 532 1064 564
rect 1004 510 1064 532
rect 910 494 927 508
rect 959 494 976 508
tri 747 458 769 480 se
rect 769 473 784 494
tri 769 458 784 473 nw
rect 1103 473 1118 649
tri 1118 642 1131 655 nw
rect 1204 574 1219 802
tri 741 452 747 458 se
rect 747 452 756 458
rect 741 436 756 452
tri 756 445 769 458 nw
rect 910 450 927 464
rect 959 450 976 464
tri 1103 458 1118 473 ne
tri 1118 458 1140 480 sw
rect 741 400 756 408
rect 822 436 882 450
rect 837 426 882 436
rect 837 408 865 426
tri 741 385 756 400 ne
tri 756 385 778 407 sw
rect 822 398 865 408
rect 880 422 882 426
rect 1004 436 1064 450
tri 1118 445 1131 458 ne
rect 1131 452 1140 458
tri 1140 452 1146 458 sw
rect 1004 426 1049 436
rect 880 398 954 422
rect 822 394 954 398
tri 954 394 982 422 sw
rect 1004 412 1006 426
tri 1004 410 1006 412 ne
rect 1018 408 1049 426
rect 1018 398 1064 408
rect 1131 437 1146 452
tri 756 373 768 385 ne
rect 768 380 778 385
tri 778 380 783 385 sw
rect 667 34 682 262
rect 768 272 783 380
rect 822 338 850 394
tri 942 376 960 394 ne
rect 960 374 982 394
tri 982 374 1002 394 sw
tri 1018 380 1036 398 ne
rect 841 304 850 338
rect 884 365 926 366
rect 884 331 889 365
rect 919 331 926 365
rect 884 322 926 331
rect 960 365 1002 374
rect 960 331 967 365
rect 997 331 1002 365
rect 960 326 1002 331
rect 1036 338 1064 398
tri 1109 385 1131 407 se
rect 1131 400 1146 408
tri 1131 385 1146 400 nw
tri 1103 379 1109 385 se
rect 1109 379 1118 385
rect 822 294 850 304
tri 850 294 874 318 sw
rect 768 224 784 272
rect 822 262 864 294
tri 881 286 882 287 sw
rect 881 262 882 286
tri 884 285 921 322 ne
rect 921 294 926 322
tri 926 294 952 320 sw
rect 1036 304 1045 338
rect 1036 294 1064 304
rect 921 285 1005 294
tri 921 266 940 285 ne
rect 940 266 1005 285
rect 822 240 882 262
rect 1004 262 1005 266
rect 1022 262 1064 294
rect 1004 240 1064 262
rect 910 224 927 238
rect 959 224 976 238
tri 747 188 769 210 se
rect 769 203 784 224
tri 769 188 784 203 nw
rect 1103 203 1118 379
tri 1118 372 1131 385 nw
rect 1204 304 1219 532
tri 741 182 747 188 se
rect 747 182 756 188
rect 741 166 756 182
tri 756 175 769 188 nw
rect 910 180 927 194
rect 959 180 976 194
tri 1103 188 1118 203 ne
tri 1118 188 1140 210 sw
rect 741 130 756 138
rect 822 166 882 180
rect 837 156 882 166
rect 837 138 865 156
tri 741 115 756 130 ne
tri 756 115 778 137 sw
rect 822 128 865 138
rect 880 152 882 156
rect 1004 166 1064 180
tri 1118 175 1131 188 ne
rect 1131 182 1140 188
tri 1140 182 1146 188 sw
rect 1004 156 1049 166
rect 880 128 954 152
rect 822 124 954 128
tri 954 124 982 152 sw
rect 1004 142 1006 156
tri 1004 140 1006 142 ne
rect 1018 138 1049 156
rect 1018 128 1064 138
rect 1131 167 1146 182
tri 756 103 768 115 ne
rect 768 110 778 115
tri 778 110 783 115 sw
rect 667 -236 682 -8
rect 768 -46 783 110
rect 822 68 850 124
tri 942 106 960 124 ne
rect 960 104 982 124
tri 982 104 1002 124 sw
tri 1018 110 1036 128 ne
rect 841 34 850 68
rect 884 95 926 96
rect 884 61 889 95
rect 919 61 926 95
rect 884 52 926 61
rect 960 95 1002 104
rect 960 61 967 95
rect 997 61 1002 95
rect 960 56 1002 61
rect 1036 68 1064 128
tri 1109 115 1131 137 se
rect 1131 130 1146 138
tri 1131 115 1146 130 nw
tri 1103 109 1109 115 se
rect 1109 109 1118 115
rect 822 24 850 34
tri 850 24 874 48 sw
rect 822 -8 864 24
tri 881 16 882 17 sw
rect 881 -8 882 16
tri 884 15 921 52 ne
rect 921 24 926 52
tri 926 24 952 50 sw
rect 1036 34 1045 68
rect 1036 24 1064 34
rect 921 15 1005 24
tri 921 -4 940 15 ne
rect 940 -4 1005 15
rect 822 -30 882 -8
rect 1004 -8 1005 -4
rect 1022 -8 1064 24
rect 1004 -30 1064 -8
rect 910 -46 927 -32
rect 959 -46 976 -32
tri 747 -82 769 -60 se
rect 769 -67 784 -46
tri 769 -82 784 -67 nw
rect 1103 -67 1118 109
tri 1118 102 1131 115 nw
rect 1204 34 1219 262
tri 741 -88 747 -82 se
rect 747 -88 756 -82
rect 741 -104 756 -88
tri 756 -95 769 -82 nw
rect 910 -90 927 -76
rect 959 -90 976 -76
tri 1103 -82 1118 -67 ne
tri 1118 -82 1140 -60 sw
rect 741 -140 756 -132
rect 822 -104 882 -90
rect 837 -114 882 -104
rect 837 -132 865 -114
tri 741 -155 756 -140 ne
tri 756 -155 778 -133 sw
rect 822 -142 865 -132
rect 880 -118 882 -114
rect 1004 -104 1064 -90
tri 1118 -95 1131 -82 ne
rect 1131 -88 1140 -82
tri 1140 -88 1146 -82 sw
rect 1004 -114 1049 -104
rect 880 -142 954 -118
rect 822 -146 954 -142
tri 954 -146 982 -118 sw
rect 1004 -128 1006 -114
tri 1004 -130 1006 -128 ne
rect 1018 -132 1049 -114
rect 1018 -142 1064 -132
rect 1131 -103 1146 -88
tri 756 -167 768 -155 ne
rect 768 -160 778 -155
tri 778 -160 783 -155 sw
rect 667 -506 682 -278
rect 768 -268 783 -160
rect 822 -202 850 -146
tri 942 -164 960 -146 ne
rect 960 -166 982 -146
tri 982 -166 1002 -146 sw
tri 1018 -160 1036 -142 ne
rect 841 -236 850 -202
rect 884 -175 926 -174
rect 884 -209 889 -175
rect 919 -209 926 -175
rect 884 -218 926 -209
rect 960 -175 1002 -166
rect 960 -209 967 -175
rect 997 -209 1002 -175
rect 960 -214 1002 -209
rect 1036 -202 1064 -142
tri 1109 -155 1131 -133 se
rect 1131 -140 1146 -132
tri 1131 -155 1146 -140 nw
tri 1103 -161 1109 -155 se
rect 1109 -161 1118 -155
rect 822 -246 850 -236
tri 850 -246 874 -222 sw
rect 768 -316 784 -268
rect 822 -278 864 -246
tri 881 -254 882 -253 sw
rect 881 -278 882 -254
tri 884 -255 921 -218 ne
rect 921 -246 926 -218
tri 926 -246 952 -220 sw
rect 1036 -236 1045 -202
rect 1036 -246 1064 -236
rect 921 -255 1005 -246
tri 921 -274 940 -255 ne
rect 940 -274 1005 -255
rect 822 -300 882 -278
rect 1004 -278 1005 -274
rect 1022 -278 1064 -246
rect 1004 -300 1064 -278
rect 910 -316 927 -302
rect 959 -316 976 -302
tri 747 -352 769 -330 se
rect 769 -337 784 -316
tri 769 -352 784 -337 nw
rect 1103 -337 1118 -161
tri 1118 -168 1131 -155 nw
rect 1204 -236 1219 -8
tri 741 -358 747 -352 se
rect 747 -358 756 -352
rect 741 -374 756 -358
tri 756 -365 769 -352 nw
rect 910 -360 927 -346
rect 959 -360 976 -346
tri 1103 -352 1118 -337 ne
tri 1118 -352 1140 -330 sw
rect 741 -410 756 -402
rect 822 -374 882 -360
rect 837 -384 882 -374
rect 837 -402 865 -384
tri 741 -425 756 -410 ne
tri 756 -425 778 -403 sw
rect 822 -412 865 -402
rect 880 -388 882 -384
rect 1004 -374 1064 -360
tri 1118 -365 1131 -352 ne
rect 1131 -358 1140 -352
tri 1140 -358 1146 -352 sw
rect 1004 -384 1049 -374
rect 880 -412 954 -388
rect 822 -416 954 -412
tri 954 -416 982 -388 sw
rect 1004 -398 1006 -384
tri 1004 -400 1006 -398 ne
rect 1018 -402 1049 -384
rect 1018 -412 1064 -402
rect 1131 -373 1146 -358
tri 756 -437 768 -425 ne
rect 768 -430 778 -425
tri 778 -430 783 -425 sw
rect 667 -776 682 -548
rect 768 -586 783 -430
rect 822 -472 850 -416
tri 942 -434 960 -416 ne
rect 960 -436 982 -416
tri 982 -436 1002 -416 sw
tri 1018 -430 1036 -412 ne
rect 841 -506 850 -472
rect 884 -445 926 -444
rect 884 -479 889 -445
rect 919 -479 926 -445
rect 884 -488 926 -479
rect 960 -445 1002 -436
rect 960 -479 967 -445
rect 997 -479 1002 -445
rect 960 -484 1002 -479
rect 1036 -472 1064 -412
tri 1109 -425 1131 -403 se
rect 1131 -410 1146 -402
tri 1131 -425 1146 -410 nw
tri 1103 -431 1109 -425 se
rect 1109 -431 1118 -425
rect 822 -516 850 -506
tri 850 -516 874 -492 sw
rect 822 -548 864 -516
tri 881 -524 882 -523 sw
rect 881 -548 882 -524
tri 884 -525 921 -488 ne
rect 921 -516 926 -488
tri 926 -516 952 -490 sw
rect 1036 -506 1045 -472
rect 1036 -516 1064 -506
rect 921 -525 1005 -516
tri 921 -544 940 -525 ne
rect 940 -544 1005 -525
rect 822 -570 882 -548
rect 1004 -548 1005 -544
rect 1022 -548 1064 -516
rect 1004 -570 1064 -548
rect 910 -586 927 -572
rect 959 -586 976 -572
tri 747 -622 769 -600 se
rect 769 -607 784 -586
tri 769 -622 784 -607 nw
rect 1103 -607 1118 -431
tri 1118 -438 1131 -425 nw
rect 1204 -506 1219 -278
tri 741 -628 747 -622 se
rect 747 -628 756 -622
rect 741 -644 756 -628
tri 756 -635 769 -622 nw
rect 910 -630 927 -616
rect 959 -630 976 -616
tri 1103 -622 1118 -607 ne
tri 1118 -622 1140 -600 sw
rect 741 -680 756 -672
rect 822 -644 882 -630
rect 837 -654 882 -644
rect 837 -672 865 -654
tri 741 -695 756 -680 ne
tri 756 -695 778 -673 sw
rect 822 -682 865 -672
rect 880 -658 882 -654
rect 1004 -644 1064 -630
tri 1118 -635 1131 -622 ne
rect 1131 -628 1140 -622
tri 1140 -628 1146 -622 sw
rect 1004 -654 1049 -644
rect 880 -682 954 -658
rect 822 -686 954 -682
tri 954 -686 982 -658 sw
rect 1004 -668 1006 -654
tri 1004 -670 1006 -668 ne
rect 1018 -672 1049 -654
rect 1018 -682 1064 -672
rect 1131 -643 1146 -628
tri 756 -707 768 -695 ne
rect 768 -700 778 -695
tri 778 -700 783 -695 sw
rect 667 -1046 682 -818
rect 768 -808 783 -700
rect 822 -742 850 -686
tri 942 -704 960 -686 ne
rect 960 -706 982 -686
tri 982 -706 1002 -686 sw
tri 1018 -700 1036 -682 ne
rect 841 -776 850 -742
rect 884 -715 926 -714
rect 884 -749 889 -715
rect 919 -749 926 -715
rect 884 -758 926 -749
rect 960 -715 1002 -706
rect 960 -749 967 -715
rect 997 -749 1002 -715
rect 960 -754 1002 -749
rect 1036 -742 1064 -682
tri 1109 -695 1131 -673 se
rect 1131 -680 1146 -672
tri 1131 -695 1146 -680 nw
tri 1103 -701 1109 -695 se
rect 1109 -701 1118 -695
rect 822 -786 850 -776
tri 850 -786 874 -762 sw
rect 768 -856 784 -808
rect 822 -818 864 -786
tri 881 -794 882 -793 sw
rect 881 -818 882 -794
tri 884 -795 921 -758 ne
rect 921 -786 926 -758
tri 926 -786 952 -760 sw
rect 1036 -776 1045 -742
rect 1036 -786 1064 -776
rect 921 -795 1005 -786
tri 921 -814 940 -795 ne
rect 940 -814 1005 -795
rect 822 -840 882 -818
rect 1004 -818 1005 -814
rect 1022 -818 1064 -786
rect 1004 -840 1064 -818
rect 910 -856 927 -842
rect 959 -856 976 -842
tri 747 -892 769 -870 se
rect 769 -877 784 -856
tri 769 -892 784 -877 nw
rect 1103 -877 1118 -701
tri 1118 -708 1131 -695 nw
rect 1204 -776 1219 -548
tri 741 -898 747 -892 se
rect 747 -898 756 -892
rect 741 -914 756 -898
tri 756 -905 769 -892 nw
rect 910 -900 927 -886
rect 959 -900 976 -886
tri 1103 -892 1118 -877 ne
tri 1118 -892 1140 -870 sw
rect 741 -950 756 -942
rect 822 -914 882 -900
rect 837 -924 882 -914
rect 837 -942 865 -924
tri 741 -965 756 -950 ne
tri 756 -965 778 -943 sw
rect 822 -952 865 -942
rect 880 -928 882 -924
rect 1004 -914 1064 -900
tri 1118 -905 1131 -892 ne
rect 1131 -898 1140 -892
tri 1140 -898 1146 -892 sw
rect 1004 -924 1049 -914
rect 880 -952 954 -928
rect 822 -956 954 -952
tri 954 -956 982 -928 sw
rect 1004 -938 1006 -924
tri 1004 -940 1006 -938 ne
rect 1018 -942 1049 -924
rect 1018 -952 1064 -942
rect 1131 -913 1146 -898
tri 756 -977 768 -965 ne
rect 768 -970 778 -965
tri 778 -970 783 -965 sw
rect 667 -1316 682 -1088
rect 768 -1126 783 -970
rect 822 -1012 850 -956
tri 942 -974 960 -956 ne
rect 960 -976 982 -956
tri 982 -976 1002 -956 sw
tri 1018 -970 1036 -952 ne
rect 841 -1046 850 -1012
rect 884 -985 926 -984
rect 884 -1019 889 -985
rect 919 -1019 926 -985
rect 884 -1028 926 -1019
rect 960 -985 1002 -976
rect 960 -1019 967 -985
rect 997 -1019 1002 -985
rect 960 -1024 1002 -1019
rect 1036 -1012 1064 -952
tri 1109 -965 1131 -943 se
rect 1131 -950 1146 -942
tri 1131 -965 1146 -950 nw
tri 1103 -971 1109 -965 se
rect 1109 -971 1118 -965
rect 822 -1056 850 -1046
tri 850 -1056 874 -1032 sw
rect 822 -1088 864 -1056
tri 881 -1064 882 -1063 sw
rect 881 -1088 882 -1064
tri 884 -1065 921 -1028 ne
rect 921 -1056 926 -1028
tri 926 -1056 952 -1030 sw
rect 1036 -1046 1045 -1012
rect 1036 -1056 1064 -1046
rect 921 -1065 1005 -1056
tri 921 -1084 940 -1065 ne
rect 940 -1084 1005 -1065
rect 822 -1110 882 -1088
rect 1004 -1088 1005 -1084
rect 1022 -1088 1064 -1056
rect 1004 -1110 1064 -1088
rect 910 -1126 927 -1112
rect 959 -1126 976 -1112
tri 747 -1162 769 -1140 se
rect 769 -1147 784 -1126
tri 769 -1162 784 -1147 nw
rect 1103 -1147 1118 -971
tri 1118 -978 1131 -965 nw
rect 1204 -1046 1219 -818
tri 741 -1168 747 -1162 se
rect 747 -1168 756 -1162
rect 741 -1184 756 -1168
tri 756 -1175 769 -1162 nw
rect 910 -1170 927 -1156
rect 959 -1170 976 -1156
tri 1103 -1162 1118 -1147 ne
tri 1118 -1162 1140 -1140 sw
rect 741 -1220 756 -1212
rect 822 -1184 882 -1170
rect 837 -1194 882 -1184
rect 837 -1212 865 -1194
tri 741 -1235 756 -1220 ne
tri 756 -1235 778 -1213 sw
rect 822 -1222 865 -1212
rect 880 -1198 882 -1194
rect 1004 -1184 1064 -1170
tri 1118 -1175 1131 -1162 ne
rect 1131 -1168 1140 -1162
tri 1140 -1168 1146 -1162 sw
rect 1004 -1194 1049 -1184
rect 880 -1222 954 -1198
rect 822 -1226 954 -1222
tri 954 -1226 982 -1198 sw
rect 1004 -1208 1006 -1194
tri 1004 -1210 1006 -1208 ne
rect 1018 -1212 1049 -1194
rect 1018 -1222 1064 -1212
rect 1131 -1183 1146 -1168
tri 756 -1247 768 -1235 ne
rect 768 -1240 778 -1235
tri 778 -1240 783 -1235 sw
rect 667 -1586 682 -1358
rect 768 -1348 783 -1240
rect 822 -1282 850 -1226
tri 942 -1244 960 -1226 ne
rect 960 -1246 982 -1226
tri 982 -1246 1002 -1226 sw
tri 1018 -1240 1036 -1222 ne
rect 841 -1316 850 -1282
rect 884 -1255 926 -1254
rect 884 -1289 889 -1255
rect 919 -1289 926 -1255
rect 884 -1298 926 -1289
rect 960 -1255 1002 -1246
rect 960 -1289 967 -1255
rect 997 -1289 1002 -1255
rect 960 -1294 1002 -1289
rect 1036 -1282 1064 -1222
tri 1109 -1235 1131 -1213 se
rect 1131 -1220 1146 -1212
tri 1131 -1235 1146 -1220 nw
tri 1103 -1241 1109 -1235 se
rect 1109 -1241 1118 -1235
rect 822 -1326 850 -1316
tri 850 -1326 874 -1302 sw
rect 768 -1396 784 -1348
rect 822 -1358 864 -1326
tri 881 -1334 882 -1333 sw
rect 881 -1358 882 -1334
tri 884 -1335 921 -1298 ne
rect 921 -1326 926 -1298
tri 926 -1326 952 -1300 sw
rect 1036 -1316 1045 -1282
rect 1036 -1326 1064 -1316
rect 921 -1335 1005 -1326
tri 921 -1354 940 -1335 ne
rect 940 -1354 1005 -1335
rect 822 -1380 882 -1358
rect 1004 -1358 1005 -1354
rect 1022 -1358 1064 -1326
rect 1004 -1380 1064 -1358
rect 910 -1396 927 -1382
rect 959 -1396 976 -1382
tri 747 -1432 769 -1410 se
rect 769 -1417 784 -1396
tri 769 -1432 784 -1417 nw
rect 1103 -1417 1118 -1241
tri 1118 -1248 1131 -1235 nw
rect 1204 -1316 1219 -1088
tri 741 -1438 747 -1432 se
rect 747 -1438 756 -1432
rect 741 -1454 756 -1438
tri 756 -1445 769 -1432 nw
rect 910 -1440 927 -1426
rect 959 -1440 976 -1426
tri 1103 -1432 1118 -1417 ne
tri 1118 -1432 1140 -1410 sw
rect 741 -1490 756 -1482
rect 822 -1454 882 -1440
rect 837 -1464 882 -1454
rect 837 -1482 865 -1464
tri 741 -1505 756 -1490 ne
tri 756 -1505 778 -1483 sw
rect 822 -1492 865 -1482
rect 880 -1468 882 -1464
rect 1004 -1454 1064 -1440
tri 1118 -1445 1131 -1432 ne
rect 1131 -1438 1140 -1432
tri 1140 -1438 1146 -1432 sw
rect 1004 -1464 1049 -1454
rect 880 -1492 954 -1468
rect 822 -1496 954 -1492
tri 954 -1496 982 -1468 sw
rect 1004 -1478 1006 -1464
tri 1004 -1480 1006 -1478 ne
rect 1018 -1482 1049 -1464
rect 1018 -1492 1064 -1482
rect 1131 -1453 1146 -1438
tri 756 -1517 768 -1505 ne
rect 768 -1510 778 -1505
tri 778 -1510 783 -1505 sw
rect 667 -1856 682 -1628
rect 768 -1666 783 -1510
rect 822 -1552 850 -1496
tri 942 -1514 960 -1496 ne
rect 960 -1516 982 -1496
tri 982 -1516 1002 -1496 sw
tri 1018 -1510 1036 -1492 ne
rect 841 -1586 850 -1552
rect 884 -1525 926 -1524
rect 884 -1559 889 -1525
rect 919 -1559 926 -1525
rect 884 -1568 926 -1559
rect 960 -1525 1002 -1516
rect 960 -1559 967 -1525
rect 997 -1559 1002 -1525
rect 960 -1564 1002 -1559
rect 1036 -1552 1064 -1492
tri 1109 -1505 1131 -1483 se
rect 1131 -1490 1146 -1482
tri 1131 -1505 1146 -1490 nw
tri 1103 -1511 1109 -1505 se
rect 1109 -1511 1118 -1505
rect 822 -1596 850 -1586
tri 850 -1596 874 -1572 sw
rect 822 -1628 864 -1596
tri 881 -1604 882 -1603 sw
rect 881 -1628 882 -1604
tri 884 -1605 921 -1568 ne
rect 921 -1596 926 -1568
tri 926 -1596 952 -1570 sw
rect 1036 -1586 1045 -1552
rect 1036 -1596 1064 -1586
rect 921 -1605 1005 -1596
tri 921 -1624 940 -1605 ne
rect 940 -1624 1005 -1605
rect 822 -1650 882 -1628
rect 1004 -1628 1005 -1624
rect 1022 -1628 1064 -1596
rect 1004 -1650 1064 -1628
rect 910 -1666 927 -1652
rect 959 -1666 976 -1652
tri 747 -1702 769 -1680 se
rect 769 -1687 784 -1666
tri 769 -1702 784 -1687 nw
rect 1103 -1687 1118 -1511
tri 1118 -1518 1131 -1505 nw
rect 1204 -1586 1219 -1358
tri 741 -1708 747 -1702 se
rect 747 -1708 756 -1702
rect 741 -1724 756 -1708
tri 756 -1715 769 -1702 nw
rect 910 -1710 927 -1696
rect 959 -1710 976 -1696
tri 1103 -1702 1118 -1687 ne
tri 1118 -1702 1140 -1680 sw
rect 741 -1760 756 -1752
rect 822 -1724 882 -1710
rect 837 -1734 882 -1724
rect 837 -1752 865 -1734
tri 741 -1775 756 -1760 ne
tri 756 -1775 778 -1753 sw
rect 822 -1762 865 -1752
rect 880 -1738 882 -1734
rect 1004 -1724 1064 -1710
tri 1118 -1715 1131 -1702 ne
rect 1131 -1708 1140 -1702
tri 1140 -1708 1146 -1702 sw
rect 1004 -1734 1049 -1724
rect 880 -1762 954 -1738
rect 822 -1766 954 -1762
tri 954 -1766 982 -1738 sw
rect 1004 -1748 1006 -1734
tri 1004 -1750 1006 -1748 ne
rect 1018 -1752 1049 -1734
rect 1018 -1762 1064 -1752
rect 1131 -1723 1146 -1708
tri 756 -1787 768 -1775 ne
rect 768 -1780 778 -1775
tri 778 -1780 783 -1775 sw
rect 667 -2126 682 -1898
rect 768 -1888 783 -1780
rect 822 -1822 850 -1766
tri 942 -1784 960 -1766 ne
rect 960 -1786 982 -1766
tri 982 -1786 1002 -1766 sw
tri 1018 -1780 1036 -1762 ne
rect 841 -1856 850 -1822
rect 884 -1795 926 -1794
rect 884 -1829 889 -1795
rect 919 -1829 926 -1795
rect 884 -1838 926 -1829
rect 960 -1795 1002 -1786
rect 960 -1829 967 -1795
rect 997 -1829 1002 -1795
rect 960 -1834 1002 -1829
rect 1036 -1822 1064 -1762
tri 1109 -1775 1131 -1753 se
rect 1131 -1760 1146 -1752
tri 1131 -1775 1146 -1760 nw
tri 1103 -1781 1109 -1775 se
rect 1109 -1781 1118 -1775
rect 822 -1866 850 -1856
tri 850 -1866 874 -1842 sw
rect 768 -1936 784 -1888
rect 822 -1898 864 -1866
tri 881 -1874 882 -1873 sw
rect 881 -1898 882 -1874
tri 884 -1875 921 -1838 ne
rect 921 -1866 926 -1838
tri 926 -1866 952 -1840 sw
rect 1036 -1856 1045 -1822
rect 1036 -1866 1064 -1856
rect 921 -1875 1005 -1866
tri 921 -1894 940 -1875 ne
rect 940 -1894 1005 -1875
rect 822 -1920 882 -1898
rect 1004 -1898 1005 -1894
rect 1022 -1898 1064 -1866
rect 1004 -1920 1064 -1898
rect 910 -1936 927 -1922
rect 959 -1936 976 -1922
tri 747 -1972 769 -1950 se
rect 769 -1957 784 -1936
tri 769 -1972 784 -1957 nw
rect 1103 -1957 1118 -1781
tri 1118 -1788 1131 -1775 nw
rect 1204 -1856 1219 -1628
tri 741 -1978 747 -1972 se
rect 747 -1978 756 -1972
rect 741 -1994 756 -1978
tri 756 -1985 769 -1972 nw
rect 910 -1980 927 -1966
rect 959 -1980 976 -1966
tri 1103 -1972 1118 -1957 ne
tri 1118 -1972 1140 -1950 sw
rect 741 -2030 756 -2022
rect 822 -1994 882 -1980
rect 837 -2004 882 -1994
rect 837 -2022 865 -2004
tri 741 -2045 756 -2030 ne
tri 756 -2045 778 -2023 sw
rect 822 -2032 865 -2022
rect 880 -2008 882 -2004
rect 1004 -1994 1064 -1980
tri 1118 -1985 1131 -1972 ne
rect 1131 -1978 1140 -1972
tri 1140 -1978 1146 -1972 sw
rect 1004 -2004 1049 -1994
rect 880 -2032 954 -2008
rect 822 -2036 954 -2032
tri 954 -2036 982 -2008 sw
rect 1004 -2018 1006 -2004
tri 1004 -2020 1006 -2018 ne
rect 1018 -2022 1049 -2004
rect 1018 -2032 1064 -2022
rect 1131 -1993 1146 -1978
tri 756 -2057 768 -2045 ne
rect 768 -2050 778 -2045
tri 778 -2050 783 -2045 sw
rect 667 -2396 682 -2168
rect 768 -2206 783 -2050
rect 822 -2092 850 -2036
tri 942 -2054 960 -2036 ne
rect 960 -2056 982 -2036
tri 982 -2056 1002 -2036 sw
tri 1018 -2050 1036 -2032 ne
rect 841 -2126 850 -2092
rect 884 -2065 926 -2064
rect 884 -2099 889 -2065
rect 919 -2099 926 -2065
rect 884 -2108 926 -2099
rect 960 -2065 1002 -2056
rect 960 -2099 967 -2065
rect 997 -2099 1002 -2065
rect 960 -2104 1002 -2099
rect 1036 -2092 1064 -2032
tri 1109 -2045 1131 -2023 se
rect 1131 -2030 1146 -2022
tri 1131 -2045 1146 -2030 nw
tri 1103 -2051 1109 -2045 se
rect 1109 -2051 1118 -2045
rect 822 -2136 850 -2126
tri 850 -2136 874 -2112 sw
rect 822 -2168 864 -2136
tri 881 -2144 882 -2143 sw
rect 881 -2168 882 -2144
tri 884 -2145 921 -2108 ne
rect 921 -2136 926 -2108
tri 926 -2136 952 -2110 sw
rect 1036 -2126 1045 -2092
rect 1036 -2136 1064 -2126
rect 921 -2145 1005 -2136
tri 921 -2164 940 -2145 ne
rect 940 -2164 1005 -2145
rect 822 -2190 882 -2168
rect 1004 -2168 1005 -2164
rect 1022 -2168 1064 -2136
rect 1004 -2190 1064 -2168
rect 910 -2206 927 -2192
rect 959 -2206 976 -2192
tri 747 -2242 769 -2220 se
rect 769 -2227 784 -2206
tri 769 -2242 784 -2227 nw
rect 1103 -2227 1118 -2051
tri 1118 -2058 1131 -2045 nw
rect 1204 -2126 1219 -1898
tri 741 -2248 747 -2242 se
rect 747 -2248 756 -2242
rect 741 -2264 756 -2248
tri 756 -2255 769 -2242 nw
rect 910 -2250 927 -2236
rect 959 -2250 976 -2236
tri 1103 -2242 1118 -2227 ne
tri 1118 -2242 1140 -2220 sw
rect 741 -2300 756 -2292
rect 822 -2264 882 -2250
rect 837 -2274 882 -2264
rect 837 -2292 865 -2274
tri 741 -2315 756 -2300 ne
tri 756 -2315 778 -2293 sw
rect 822 -2302 865 -2292
rect 880 -2278 882 -2274
rect 1004 -2264 1064 -2250
tri 1118 -2255 1131 -2242 ne
rect 1131 -2248 1140 -2242
tri 1140 -2248 1146 -2242 sw
rect 1004 -2274 1049 -2264
rect 880 -2302 954 -2278
rect 822 -2306 954 -2302
tri 954 -2306 982 -2278 sw
rect 1004 -2288 1006 -2274
tri 1004 -2290 1006 -2288 ne
rect 1018 -2292 1049 -2274
rect 1018 -2302 1064 -2292
rect 1131 -2263 1146 -2248
tri 756 -2327 768 -2315 ne
rect 768 -2320 778 -2315
tri 778 -2320 783 -2315 sw
rect 667 -2524 682 -2438
rect 768 -2476 783 -2320
rect 822 -2362 850 -2306
tri 942 -2324 960 -2306 ne
rect 960 -2326 982 -2306
tri 982 -2326 1002 -2306 sw
tri 1018 -2320 1036 -2302 ne
rect 841 -2396 850 -2362
rect 884 -2335 926 -2334
rect 884 -2369 889 -2335
rect 919 -2369 926 -2335
rect 884 -2378 926 -2369
rect 960 -2335 1002 -2326
rect 960 -2369 967 -2335
rect 997 -2369 1002 -2335
rect 960 -2374 1002 -2369
rect 1036 -2362 1064 -2302
tri 1109 -2315 1131 -2293 se
rect 1131 -2300 1146 -2292
tri 1131 -2315 1146 -2300 nw
tri 1103 -2321 1109 -2315 se
rect 1109 -2321 1118 -2315
rect 822 -2406 850 -2396
tri 850 -2406 874 -2382 sw
rect 822 -2438 864 -2406
tri 881 -2414 882 -2413 sw
rect 881 -2438 882 -2414
tri 884 -2415 921 -2378 ne
rect 921 -2406 926 -2378
tri 926 -2406 952 -2380 sw
rect 1036 -2396 1045 -2362
rect 1036 -2406 1064 -2396
rect 921 -2415 1005 -2406
tri 921 -2434 940 -2415 ne
rect 940 -2434 1005 -2415
rect 822 -2460 882 -2438
rect 1004 -2438 1005 -2434
rect 1022 -2438 1064 -2406
rect 1004 -2460 1064 -2438
rect 910 -2476 927 -2462
rect 959 -2476 976 -2462
rect 1103 -2476 1118 -2321
tri 1118 -2328 1131 -2315 nw
rect 1204 -2396 1219 -2168
rect 1204 -2524 1219 -2438
rect 1247 1654 1262 1844
tri 1327 1808 1349 1830 se
rect 1349 1823 1364 1892
tri 1349 1808 1364 1823 nw
rect 1683 1823 1698 1892
tri 1321 1802 1327 1808 se
rect 1327 1802 1336 1808
rect 1321 1786 1336 1802
tri 1336 1795 1349 1808 nw
rect 1490 1800 1507 1814
rect 1539 1800 1556 1814
tri 1683 1808 1698 1823 ne
tri 1698 1808 1720 1830 sw
rect 1321 1750 1336 1758
rect 1402 1786 1462 1800
rect 1417 1776 1462 1786
rect 1417 1758 1445 1776
tri 1321 1735 1336 1750 ne
tri 1336 1735 1358 1757 sw
rect 1402 1748 1445 1758
rect 1460 1772 1462 1776
rect 1584 1786 1644 1800
tri 1698 1795 1711 1808 ne
rect 1711 1802 1720 1808
tri 1720 1802 1726 1808 sw
rect 1584 1776 1629 1786
rect 1460 1748 1534 1772
rect 1402 1744 1534 1748
tri 1534 1744 1562 1772 sw
rect 1584 1762 1586 1776
tri 1584 1760 1586 1762 ne
rect 1598 1758 1629 1776
rect 1598 1748 1644 1758
rect 1711 1787 1726 1802
tri 1336 1723 1348 1735 ne
rect 1348 1730 1358 1735
tri 1358 1730 1363 1735 sw
rect 1247 1384 1262 1612
rect 1348 1574 1363 1730
rect 1402 1688 1430 1744
tri 1522 1726 1540 1744 ne
rect 1540 1724 1562 1744
tri 1562 1724 1582 1744 sw
tri 1598 1730 1616 1748 ne
rect 1421 1654 1430 1688
rect 1464 1715 1506 1716
rect 1464 1681 1469 1715
rect 1499 1681 1506 1715
rect 1464 1672 1506 1681
rect 1540 1715 1582 1724
rect 1540 1681 1547 1715
rect 1577 1681 1582 1715
rect 1540 1676 1582 1681
rect 1616 1688 1644 1748
tri 1689 1735 1711 1757 se
rect 1711 1750 1726 1758
tri 1711 1735 1726 1750 nw
tri 1683 1729 1689 1735 se
rect 1689 1729 1698 1735
rect 1402 1644 1430 1654
tri 1430 1644 1454 1668 sw
rect 1402 1612 1444 1644
tri 1461 1636 1462 1637 sw
rect 1461 1612 1462 1636
tri 1464 1635 1501 1672 ne
rect 1501 1644 1506 1672
tri 1506 1644 1532 1670 sw
rect 1616 1654 1625 1688
rect 1616 1644 1644 1654
rect 1501 1635 1585 1644
tri 1501 1616 1520 1635 ne
rect 1520 1616 1585 1635
rect 1402 1590 1462 1612
rect 1584 1612 1585 1616
rect 1602 1612 1644 1644
rect 1584 1590 1644 1612
rect 1490 1574 1507 1588
rect 1539 1574 1556 1588
tri 1327 1538 1349 1560 se
rect 1349 1553 1364 1574
tri 1349 1538 1364 1553 nw
rect 1683 1553 1698 1729
tri 1698 1722 1711 1735 nw
rect 1784 1654 1799 1844
tri 1321 1532 1327 1538 se
rect 1327 1532 1336 1538
rect 1321 1516 1336 1532
tri 1336 1525 1349 1538 nw
rect 1490 1530 1507 1544
rect 1539 1530 1556 1544
tri 1683 1538 1698 1553 ne
tri 1698 1538 1720 1560 sw
rect 1321 1480 1336 1488
rect 1402 1516 1462 1530
rect 1417 1506 1462 1516
rect 1417 1488 1445 1506
tri 1321 1465 1336 1480 ne
tri 1336 1465 1358 1487 sw
rect 1402 1478 1445 1488
rect 1460 1502 1462 1506
rect 1584 1516 1644 1530
tri 1698 1525 1711 1538 ne
rect 1711 1532 1720 1538
tri 1720 1532 1726 1538 sw
rect 1584 1506 1629 1516
rect 1460 1478 1534 1502
rect 1402 1474 1534 1478
tri 1534 1474 1562 1502 sw
rect 1584 1492 1586 1506
tri 1584 1490 1586 1492 ne
rect 1598 1488 1629 1506
rect 1598 1478 1644 1488
rect 1711 1517 1726 1532
tri 1336 1453 1348 1465 ne
rect 1348 1460 1358 1465
tri 1358 1460 1363 1465 sw
rect 1247 1114 1262 1342
rect 1348 1352 1363 1460
rect 1402 1418 1430 1474
tri 1522 1456 1540 1474 ne
rect 1540 1454 1562 1474
tri 1562 1454 1582 1474 sw
tri 1598 1460 1616 1478 ne
rect 1421 1384 1430 1418
rect 1464 1445 1506 1446
rect 1464 1411 1469 1445
rect 1499 1411 1506 1445
rect 1464 1402 1506 1411
rect 1540 1445 1582 1454
rect 1540 1411 1547 1445
rect 1577 1411 1582 1445
rect 1540 1406 1582 1411
rect 1616 1418 1644 1478
tri 1689 1465 1711 1487 se
rect 1711 1480 1726 1488
tri 1711 1465 1726 1480 nw
tri 1683 1459 1689 1465 se
rect 1689 1459 1698 1465
rect 1402 1374 1430 1384
tri 1430 1374 1454 1398 sw
rect 1348 1304 1364 1352
rect 1402 1342 1444 1374
tri 1461 1366 1462 1367 sw
rect 1461 1342 1462 1366
tri 1464 1365 1501 1402 ne
rect 1501 1374 1506 1402
tri 1506 1374 1532 1400 sw
rect 1616 1384 1625 1418
rect 1616 1374 1644 1384
rect 1501 1365 1585 1374
tri 1501 1346 1520 1365 ne
rect 1520 1346 1585 1365
rect 1402 1320 1462 1342
rect 1584 1342 1585 1346
rect 1602 1342 1644 1374
rect 1584 1320 1644 1342
rect 1490 1304 1507 1318
rect 1539 1304 1556 1318
tri 1327 1268 1349 1290 se
rect 1349 1283 1364 1304
tri 1349 1268 1364 1283 nw
rect 1683 1283 1698 1459
tri 1698 1452 1711 1465 nw
rect 1784 1384 1799 1612
tri 1321 1262 1327 1268 se
rect 1327 1262 1336 1268
rect 1321 1246 1336 1262
tri 1336 1255 1349 1268 nw
rect 1490 1260 1507 1274
rect 1539 1260 1556 1274
tri 1683 1268 1698 1283 ne
tri 1698 1268 1720 1290 sw
rect 1321 1210 1336 1218
rect 1402 1246 1462 1260
rect 1417 1236 1462 1246
rect 1417 1218 1445 1236
tri 1321 1195 1336 1210 ne
tri 1336 1195 1358 1217 sw
rect 1402 1208 1445 1218
rect 1460 1232 1462 1236
rect 1584 1246 1644 1260
tri 1698 1255 1711 1268 ne
rect 1711 1262 1720 1268
tri 1720 1262 1726 1268 sw
rect 1584 1236 1629 1246
rect 1460 1208 1534 1232
rect 1402 1204 1534 1208
tri 1534 1204 1562 1232 sw
rect 1584 1222 1586 1236
tri 1584 1220 1586 1222 ne
rect 1598 1218 1629 1236
rect 1598 1208 1644 1218
rect 1711 1247 1726 1262
tri 1336 1183 1348 1195 ne
rect 1348 1190 1358 1195
tri 1358 1190 1363 1195 sw
rect 1247 844 1262 1072
rect 1348 1034 1363 1190
rect 1402 1148 1430 1204
tri 1522 1186 1540 1204 ne
rect 1540 1184 1562 1204
tri 1562 1184 1582 1204 sw
tri 1598 1190 1616 1208 ne
rect 1421 1114 1430 1148
rect 1464 1175 1506 1176
rect 1464 1141 1469 1175
rect 1499 1141 1506 1175
rect 1464 1132 1506 1141
rect 1540 1175 1582 1184
rect 1540 1141 1547 1175
rect 1577 1141 1582 1175
rect 1540 1136 1582 1141
rect 1616 1148 1644 1208
tri 1689 1195 1711 1217 se
rect 1711 1210 1726 1218
tri 1711 1195 1726 1210 nw
tri 1683 1189 1689 1195 se
rect 1689 1189 1698 1195
rect 1402 1104 1430 1114
tri 1430 1104 1454 1128 sw
rect 1402 1072 1444 1104
tri 1461 1096 1462 1097 sw
rect 1461 1072 1462 1096
tri 1464 1095 1501 1132 ne
rect 1501 1104 1506 1132
tri 1506 1104 1532 1130 sw
rect 1616 1114 1625 1148
rect 1616 1104 1644 1114
rect 1501 1095 1585 1104
tri 1501 1076 1520 1095 ne
rect 1520 1076 1585 1095
rect 1402 1050 1462 1072
rect 1584 1072 1585 1076
rect 1602 1072 1644 1104
rect 1584 1050 1644 1072
rect 1490 1034 1507 1048
rect 1539 1034 1556 1048
tri 1327 998 1349 1020 se
rect 1349 1013 1364 1034
tri 1349 998 1364 1013 nw
rect 1683 1013 1698 1189
tri 1698 1182 1711 1195 nw
rect 1784 1114 1799 1342
tri 1321 992 1327 998 se
rect 1327 992 1336 998
rect 1321 976 1336 992
tri 1336 985 1349 998 nw
rect 1490 990 1507 1004
rect 1539 990 1556 1004
tri 1683 998 1698 1013 ne
tri 1698 998 1720 1020 sw
rect 1321 940 1336 948
rect 1402 976 1462 990
rect 1417 966 1462 976
rect 1417 948 1445 966
tri 1321 925 1336 940 ne
tri 1336 925 1358 947 sw
rect 1402 938 1445 948
rect 1460 962 1462 966
rect 1584 976 1644 990
tri 1698 985 1711 998 ne
rect 1711 992 1720 998
tri 1720 992 1726 998 sw
rect 1584 966 1629 976
rect 1460 938 1534 962
rect 1402 934 1534 938
tri 1534 934 1562 962 sw
rect 1584 952 1586 966
tri 1584 950 1586 952 ne
rect 1598 948 1629 966
rect 1598 938 1644 948
rect 1711 977 1726 992
tri 1336 913 1348 925 ne
rect 1348 920 1358 925
tri 1358 920 1363 925 sw
rect 1247 574 1262 802
rect 1348 812 1363 920
rect 1402 878 1430 934
tri 1522 916 1540 934 ne
rect 1540 914 1562 934
tri 1562 914 1582 934 sw
tri 1598 920 1616 938 ne
rect 1421 844 1430 878
rect 1464 905 1506 906
rect 1464 871 1469 905
rect 1499 871 1506 905
rect 1464 862 1506 871
rect 1540 905 1582 914
rect 1540 871 1547 905
rect 1577 871 1582 905
rect 1540 866 1582 871
rect 1616 878 1644 938
tri 1689 925 1711 947 se
rect 1711 940 1726 948
tri 1711 925 1726 940 nw
tri 1683 919 1689 925 se
rect 1689 919 1698 925
rect 1402 834 1430 844
tri 1430 834 1454 858 sw
rect 1348 764 1364 812
rect 1402 802 1444 834
tri 1461 826 1462 827 sw
rect 1461 802 1462 826
tri 1464 825 1501 862 ne
rect 1501 834 1506 862
tri 1506 834 1532 860 sw
rect 1616 844 1625 878
rect 1616 834 1644 844
rect 1501 825 1585 834
tri 1501 806 1520 825 ne
rect 1520 806 1585 825
rect 1402 780 1462 802
rect 1584 802 1585 806
rect 1602 802 1644 834
rect 1584 780 1644 802
rect 1490 764 1507 778
rect 1539 764 1556 778
tri 1327 728 1349 750 se
rect 1349 743 1364 764
tri 1349 728 1364 743 nw
rect 1683 743 1698 919
tri 1698 912 1711 925 nw
rect 1784 844 1799 1072
tri 1321 722 1327 728 se
rect 1327 722 1336 728
rect 1321 706 1336 722
tri 1336 715 1349 728 nw
rect 1490 720 1507 734
rect 1539 720 1556 734
tri 1683 728 1698 743 ne
tri 1698 728 1720 750 sw
rect 1321 670 1336 678
rect 1402 706 1462 720
rect 1417 696 1462 706
rect 1417 678 1445 696
tri 1321 655 1336 670 ne
tri 1336 655 1358 677 sw
rect 1402 668 1445 678
rect 1460 692 1462 696
rect 1584 706 1644 720
tri 1698 715 1711 728 ne
rect 1711 722 1720 728
tri 1720 722 1726 728 sw
rect 1584 696 1629 706
rect 1460 668 1534 692
rect 1402 664 1534 668
tri 1534 664 1562 692 sw
rect 1584 682 1586 696
tri 1584 680 1586 682 ne
rect 1598 678 1629 696
rect 1598 668 1644 678
rect 1711 707 1726 722
tri 1336 643 1348 655 ne
rect 1348 650 1358 655
tri 1358 650 1363 655 sw
rect 1247 304 1262 532
rect 1348 494 1363 650
rect 1402 608 1430 664
tri 1522 646 1540 664 ne
rect 1540 644 1562 664
tri 1562 644 1582 664 sw
tri 1598 650 1616 668 ne
rect 1421 574 1430 608
rect 1464 635 1506 636
rect 1464 601 1469 635
rect 1499 601 1506 635
rect 1464 592 1506 601
rect 1540 635 1582 644
rect 1540 601 1547 635
rect 1577 601 1582 635
rect 1540 596 1582 601
rect 1616 608 1644 668
tri 1689 655 1711 677 se
rect 1711 670 1726 678
tri 1711 655 1726 670 nw
tri 1683 649 1689 655 se
rect 1689 649 1698 655
rect 1402 564 1430 574
tri 1430 564 1454 588 sw
rect 1402 532 1444 564
tri 1461 556 1462 557 sw
rect 1461 532 1462 556
tri 1464 555 1501 592 ne
rect 1501 564 1506 592
tri 1506 564 1532 590 sw
rect 1616 574 1625 608
rect 1616 564 1644 574
rect 1501 555 1585 564
tri 1501 536 1520 555 ne
rect 1520 536 1585 555
rect 1402 510 1462 532
rect 1584 532 1585 536
rect 1602 532 1644 564
rect 1584 510 1644 532
rect 1490 494 1507 508
rect 1539 494 1556 508
tri 1327 458 1349 480 se
rect 1349 473 1364 494
tri 1349 458 1364 473 nw
rect 1683 473 1698 649
tri 1698 642 1711 655 nw
rect 1784 574 1799 802
tri 1321 452 1327 458 se
rect 1327 452 1336 458
rect 1321 436 1336 452
tri 1336 445 1349 458 nw
rect 1490 450 1507 464
rect 1539 450 1556 464
tri 1683 458 1698 473 ne
tri 1698 458 1720 480 sw
rect 1321 400 1336 408
rect 1402 436 1462 450
rect 1417 426 1462 436
rect 1417 408 1445 426
tri 1321 385 1336 400 ne
tri 1336 385 1358 407 sw
rect 1402 398 1445 408
rect 1460 422 1462 426
rect 1584 436 1644 450
tri 1698 445 1711 458 ne
rect 1711 452 1720 458
tri 1720 452 1726 458 sw
rect 1584 426 1629 436
rect 1460 398 1534 422
rect 1402 394 1534 398
tri 1534 394 1562 422 sw
rect 1584 412 1586 426
tri 1584 410 1586 412 ne
rect 1598 408 1629 426
rect 1598 398 1644 408
rect 1711 437 1726 452
tri 1336 373 1348 385 ne
rect 1348 380 1358 385
tri 1358 380 1363 385 sw
rect 1247 34 1262 262
rect 1348 272 1363 380
rect 1402 338 1430 394
tri 1522 376 1540 394 ne
rect 1540 374 1562 394
tri 1562 374 1582 394 sw
tri 1598 380 1616 398 ne
rect 1421 304 1430 338
rect 1464 365 1506 366
rect 1464 331 1469 365
rect 1499 331 1506 365
rect 1464 322 1506 331
rect 1540 365 1582 374
rect 1540 331 1547 365
rect 1577 331 1582 365
rect 1540 326 1582 331
rect 1616 338 1644 398
tri 1689 385 1711 407 se
rect 1711 400 1726 408
tri 1711 385 1726 400 nw
tri 1683 379 1689 385 se
rect 1689 379 1698 385
rect 1402 294 1430 304
tri 1430 294 1454 318 sw
rect 1348 224 1364 272
rect 1402 262 1444 294
tri 1461 286 1462 287 sw
rect 1461 262 1462 286
tri 1464 285 1501 322 ne
rect 1501 294 1506 322
tri 1506 294 1532 320 sw
rect 1616 304 1625 338
rect 1616 294 1644 304
rect 1501 285 1585 294
tri 1501 266 1520 285 ne
rect 1520 266 1585 285
rect 1402 240 1462 262
rect 1584 262 1585 266
rect 1602 262 1644 294
rect 1584 240 1644 262
rect 1490 224 1507 238
rect 1539 224 1556 238
tri 1327 188 1349 210 se
rect 1349 203 1364 224
tri 1349 188 1364 203 nw
rect 1683 203 1698 379
tri 1698 372 1711 385 nw
rect 1784 304 1799 532
tri 1321 182 1327 188 se
rect 1327 182 1336 188
rect 1321 166 1336 182
tri 1336 175 1349 188 nw
rect 1490 180 1507 194
rect 1539 180 1556 194
tri 1683 188 1698 203 ne
tri 1698 188 1720 210 sw
rect 1321 130 1336 138
rect 1402 166 1462 180
rect 1417 156 1462 166
rect 1417 138 1445 156
tri 1321 115 1336 130 ne
tri 1336 115 1358 137 sw
rect 1402 128 1445 138
rect 1460 152 1462 156
rect 1584 166 1644 180
tri 1698 175 1711 188 ne
rect 1711 182 1720 188
tri 1720 182 1726 188 sw
rect 1584 156 1629 166
rect 1460 128 1534 152
rect 1402 124 1534 128
tri 1534 124 1562 152 sw
rect 1584 142 1586 156
tri 1584 140 1586 142 ne
rect 1598 138 1629 156
rect 1598 128 1644 138
rect 1711 167 1726 182
tri 1336 103 1348 115 ne
rect 1348 110 1358 115
tri 1358 110 1363 115 sw
rect 1247 -236 1262 -8
rect 1348 -46 1363 110
rect 1402 68 1430 124
tri 1522 106 1540 124 ne
rect 1540 104 1562 124
tri 1562 104 1582 124 sw
tri 1598 110 1616 128 ne
rect 1421 34 1430 68
rect 1464 95 1506 96
rect 1464 61 1469 95
rect 1499 61 1506 95
rect 1464 52 1506 61
rect 1540 95 1582 104
rect 1540 61 1547 95
rect 1577 61 1582 95
rect 1540 56 1582 61
rect 1616 68 1644 128
tri 1689 115 1711 137 se
rect 1711 130 1726 138
tri 1711 115 1726 130 nw
tri 1683 109 1689 115 se
rect 1689 109 1698 115
rect 1402 24 1430 34
tri 1430 24 1454 48 sw
rect 1402 -8 1444 24
tri 1461 16 1462 17 sw
rect 1461 -8 1462 16
tri 1464 15 1501 52 ne
rect 1501 24 1506 52
tri 1506 24 1532 50 sw
rect 1616 34 1625 68
rect 1616 24 1644 34
rect 1501 15 1585 24
tri 1501 -4 1520 15 ne
rect 1520 -4 1585 15
rect 1402 -30 1462 -8
rect 1584 -8 1585 -4
rect 1602 -8 1644 24
rect 1584 -30 1644 -8
rect 1490 -46 1507 -32
rect 1539 -46 1556 -32
tri 1327 -82 1349 -60 se
rect 1349 -67 1364 -46
tri 1349 -82 1364 -67 nw
rect 1683 -67 1698 109
tri 1698 102 1711 115 nw
rect 1784 34 1799 262
tri 1321 -88 1327 -82 se
rect 1327 -88 1336 -82
rect 1321 -104 1336 -88
tri 1336 -95 1349 -82 nw
rect 1490 -90 1507 -76
rect 1539 -90 1556 -76
tri 1683 -82 1698 -67 ne
tri 1698 -82 1720 -60 sw
rect 1321 -140 1336 -132
rect 1402 -104 1462 -90
rect 1417 -114 1462 -104
rect 1417 -132 1445 -114
tri 1321 -155 1336 -140 ne
tri 1336 -155 1358 -133 sw
rect 1402 -142 1445 -132
rect 1460 -118 1462 -114
rect 1584 -104 1644 -90
tri 1698 -95 1711 -82 ne
rect 1711 -88 1720 -82
tri 1720 -88 1726 -82 sw
rect 1584 -114 1629 -104
rect 1460 -142 1534 -118
rect 1402 -146 1534 -142
tri 1534 -146 1562 -118 sw
rect 1584 -128 1586 -114
tri 1584 -130 1586 -128 ne
rect 1598 -132 1629 -114
rect 1598 -142 1644 -132
rect 1711 -103 1726 -88
tri 1336 -167 1348 -155 ne
rect 1348 -160 1358 -155
tri 1358 -160 1363 -155 sw
rect 1247 -506 1262 -278
rect 1348 -268 1363 -160
rect 1402 -202 1430 -146
tri 1522 -164 1540 -146 ne
rect 1540 -166 1562 -146
tri 1562 -166 1582 -146 sw
tri 1598 -160 1616 -142 ne
rect 1421 -236 1430 -202
rect 1464 -175 1506 -174
rect 1464 -209 1469 -175
rect 1499 -209 1506 -175
rect 1464 -218 1506 -209
rect 1540 -175 1582 -166
rect 1540 -209 1547 -175
rect 1577 -209 1582 -175
rect 1540 -214 1582 -209
rect 1616 -202 1644 -142
tri 1689 -155 1711 -133 se
rect 1711 -140 1726 -132
tri 1711 -155 1726 -140 nw
tri 1683 -161 1689 -155 se
rect 1689 -161 1698 -155
rect 1402 -246 1430 -236
tri 1430 -246 1454 -222 sw
rect 1348 -316 1364 -268
rect 1402 -278 1444 -246
tri 1461 -254 1462 -253 sw
rect 1461 -278 1462 -254
tri 1464 -255 1501 -218 ne
rect 1501 -246 1506 -218
tri 1506 -246 1532 -220 sw
rect 1616 -236 1625 -202
rect 1616 -246 1644 -236
rect 1501 -255 1585 -246
tri 1501 -274 1520 -255 ne
rect 1520 -274 1585 -255
rect 1402 -300 1462 -278
rect 1584 -278 1585 -274
rect 1602 -278 1644 -246
rect 1584 -300 1644 -278
rect 1490 -316 1507 -302
rect 1539 -316 1556 -302
tri 1327 -352 1349 -330 se
rect 1349 -337 1364 -316
tri 1349 -352 1364 -337 nw
rect 1683 -337 1698 -161
tri 1698 -168 1711 -155 nw
rect 1784 -236 1799 -8
tri 1321 -358 1327 -352 se
rect 1327 -358 1336 -352
rect 1321 -374 1336 -358
tri 1336 -365 1349 -352 nw
rect 1490 -360 1507 -346
rect 1539 -360 1556 -346
tri 1683 -352 1698 -337 ne
tri 1698 -352 1720 -330 sw
rect 1321 -410 1336 -402
rect 1402 -374 1462 -360
rect 1417 -384 1462 -374
rect 1417 -402 1445 -384
tri 1321 -425 1336 -410 ne
tri 1336 -425 1358 -403 sw
rect 1402 -412 1445 -402
rect 1460 -388 1462 -384
rect 1584 -374 1644 -360
tri 1698 -365 1711 -352 ne
rect 1711 -358 1720 -352
tri 1720 -358 1726 -352 sw
rect 1584 -384 1629 -374
rect 1460 -412 1534 -388
rect 1402 -416 1534 -412
tri 1534 -416 1562 -388 sw
rect 1584 -398 1586 -384
tri 1584 -400 1586 -398 ne
rect 1598 -402 1629 -384
rect 1598 -412 1644 -402
rect 1711 -373 1726 -358
tri 1336 -437 1348 -425 ne
rect 1348 -430 1358 -425
tri 1358 -430 1363 -425 sw
rect 1247 -776 1262 -548
rect 1348 -586 1363 -430
rect 1402 -472 1430 -416
tri 1522 -434 1540 -416 ne
rect 1540 -436 1562 -416
tri 1562 -436 1582 -416 sw
tri 1598 -430 1616 -412 ne
rect 1421 -506 1430 -472
rect 1464 -445 1506 -444
rect 1464 -479 1469 -445
rect 1499 -479 1506 -445
rect 1464 -488 1506 -479
rect 1540 -445 1582 -436
rect 1540 -479 1547 -445
rect 1577 -479 1582 -445
rect 1540 -484 1582 -479
rect 1616 -472 1644 -412
tri 1689 -425 1711 -403 se
rect 1711 -410 1726 -402
tri 1711 -425 1726 -410 nw
tri 1683 -431 1689 -425 se
rect 1689 -431 1698 -425
rect 1402 -516 1430 -506
tri 1430 -516 1454 -492 sw
rect 1402 -548 1444 -516
tri 1461 -524 1462 -523 sw
rect 1461 -548 1462 -524
tri 1464 -525 1501 -488 ne
rect 1501 -516 1506 -488
tri 1506 -516 1532 -490 sw
rect 1616 -506 1625 -472
rect 1616 -516 1644 -506
rect 1501 -525 1585 -516
tri 1501 -544 1520 -525 ne
rect 1520 -544 1585 -525
rect 1402 -570 1462 -548
rect 1584 -548 1585 -544
rect 1602 -548 1644 -516
rect 1584 -570 1644 -548
rect 1490 -586 1507 -572
rect 1539 -586 1556 -572
tri 1327 -622 1349 -600 se
rect 1349 -607 1364 -586
tri 1349 -622 1364 -607 nw
rect 1683 -607 1698 -431
tri 1698 -438 1711 -425 nw
rect 1784 -506 1799 -278
tri 1321 -628 1327 -622 se
rect 1327 -628 1336 -622
rect 1321 -644 1336 -628
tri 1336 -635 1349 -622 nw
rect 1490 -630 1507 -616
rect 1539 -630 1556 -616
tri 1683 -622 1698 -607 ne
tri 1698 -622 1720 -600 sw
rect 1321 -680 1336 -672
rect 1402 -644 1462 -630
rect 1417 -654 1462 -644
rect 1417 -672 1445 -654
tri 1321 -695 1336 -680 ne
tri 1336 -695 1358 -673 sw
rect 1402 -682 1445 -672
rect 1460 -658 1462 -654
rect 1584 -644 1644 -630
tri 1698 -635 1711 -622 ne
rect 1711 -628 1720 -622
tri 1720 -628 1726 -622 sw
rect 1584 -654 1629 -644
rect 1460 -682 1534 -658
rect 1402 -686 1534 -682
tri 1534 -686 1562 -658 sw
rect 1584 -668 1586 -654
tri 1584 -670 1586 -668 ne
rect 1598 -672 1629 -654
rect 1598 -682 1644 -672
rect 1711 -643 1726 -628
tri 1336 -707 1348 -695 ne
rect 1348 -700 1358 -695
tri 1358 -700 1363 -695 sw
rect 1247 -1046 1262 -818
rect 1348 -808 1363 -700
rect 1402 -742 1430 -686
tri 1522 -704 1540 -686 ne
rect 1540 -706 1562 -686
tri 1562 -706 1582 -686 sw
tri 1598 -700 1616 -682 ne
rect 1421 -776 1430 -742
rect 1464 -715 1506 -714
rect 1464 -749 1469 -715
rect 1499 -749 1506 -715
rect 1464 -758 1506 -749
rect 1540 -715 1582 -706
rect 1540 -749 1547 -715
rect 1577 -749 1582 -715
rect 1540 -754 1582 -749
rect 1616 -742 1644 -682
tri 1689 -695 1711 -673 se
rect 1711 -680 1726 -672
tri 1711 -695 1726 -680 nw
tri 1683 -701 1689 -695 se
rect 1689 -701 1698 -695
rect 1402 -786 1430 -776
tri 1430 -786 1454 -762 sw
rect 1348 -856 1364 -808
rect 1402 -818 1444 -786
tri 1461 -794 1462 -793 sw
rect 1461 -818 1462 -794
tri 1464 -795 1501 -758 ne
rect 1501 -786 1506 -758
tri 1506 -786 1532 -760 sw
rect 1616 -776 1625 -742
rect 1616 -786 1644 -776
rect 1501 -795 1585 -786
tri 1501 -814 1520 -795 ne
rect 1520 -814 1585 -795
rect 1402 -840 1462 -818
rect 1584 -818 1585 -814
rect 1602 -818 1644 -786
rect 1584 -840 1644 -818
rect 1490 -856 1507 -842
rect 1539 -856 1556 -842
tri 1327 -892 1349 -870 se
rect 1349 -877 1364 -856
tri 1349 -892 1364 -877 nw
rect 1683 -877 1698 -701
tri 1698 -708 1711 -695 nw
rect 1784 -776 1799 -548
tri 1321 -898 1327 -892 se
rect 1327 -898 1336 -892
rect 1321 -914 1336 -898
tri 1336 -905 1349 -892 nw
rect 1490 -900 1507 -886
rect 1539 -900 1556 -886
tri 1683 -892 1698 -877 ne
tri 1698 -892 1720 -870 sw
rect 1321 -950 1336 -942
rect 1402 -914 1462 -900
rect 1417 -924 1462 -914
rect 1417 -942 1445 -924
tri 1321 -965 1336 -950 ne
tri 1336 -965 1358 -943 sw
rect 1402 -952 1445 -942
rect 1460 -928 1462 -924
rect 1584 -914 1644 -900
tri 1698 -905 1711 -892 ne
rect 1711 -898 1720 -892
tri 1720 -898 1726 -892 sw
rect 1584 -924 1629 -914
rect 1460 -952 1534 -928
rect 1402 -956 1534 -952
tri 1534 -956 1562 -928 sw
rect 1584 -938 1586 -924
tri 1584 -940 1586 -938 ne
rect 1598 -942 1629 -924
rect 1598 -952 1644 -942
rect 1711 -913 1726 -898
tri 1336 -977 1348 -965 ne
rect 1348 -970 1358 -965
tri 1358 -970 1363 -965 sw
rect 1247 -1316 1262 -1088
rect 1348 -1126 1363 -970
rect 1402 -1012 1430 -956
tri 1522 -974 1540 -956 ne
rect 1540 -976 1562 -956
tri 1562 -976 1582 -956 sw
tri 1598 -970 1616 -952 ne
rect 1421 -1046 1430 -1012
rect 1464 -985 1506 -984
rect 1464 -1019 1469 -985
rect 1499 -1019 1506 -985
rect 1464 -1028 1506 -1019
rect 1540 -985 1582 -976
rect 1540 -1019 1547 -985
rect 1577 -1019 1582 -985
rect 1540 -1024 1582 -1019
rect 1616 -1012 1644 -952
tri 1689 -965 1711 -943 se
rect 1711 -950 1726 -942
tri 1711 -965 1726 -950 nw
tri 1683 -971 1689 -965 se
rect 1689 -971 1698 -965
rect 1402 -1056 1430 -1046
tri 1430 -1056 1454 -1032 sw
rect 1402 -1088 1444 -1056
tri 1461 -1064 1462 -1063 sw
rect 1461 -1088 1462 -1064
tri 1464 -1065 1501 -1028 ne
rect 1501 -1056 1506 -1028
tri 1506 -1056 1532 -1030 sw
rect 1616 -1046 1625 -1012
rect 1616 -1056 1644 -1046
rect 1501 -1065 1585 -1056
tri 1501 -1084 1520 -1065 ne
rect 1520 -1084 1585 -1065
rect 1402 -1110 1462 -1088
rect 1584 -1088 1585 -1084
rect 1602 -1088 1644 -1056
rect 1584 -1110 1644 -1088
rect 1490 -1126 1507 -1112
rect 1539 -1126 1556 -1112
tri 1327 -1162 1349 -1140 se
rect 1349 -1147 1364 -1126
tri 1349 -1162 1364 -1147 nw
rect 1683 -1147 1698 -971
tri 1698 -978 1711 -965 nw
rect 1784 -1046 1799 -818
tri 1321 -1168 1327 -1162 se
rect 1327 -1168 1336 -1162
rect 1321 -1184 1336 -1168
tri 1336 -1175 1349 -1162 nw
rect 1490 -1170 1507 -1156
rect 1539 -1170 1556 -1156
tri 1683 -1162 1698 -1147 ne
tri 1698 -1162 1720 -1140 sw
rect 1321 -1220 1336 -1212
rect 1402 -1184 1462 -1170
rect 1417 -1194 1462 -1184
rect 1417 -1212 1445 -1194
tri 1321 -1235 1336 -1220 ne
tri 1336 -1235 1358 -1213 sw
rect 1402 -1222 1445 -1212
rect 1460 -1198 1462 -1194
rect 1584 -1184 1644 -1170
tri 1698 -1175 1711 -1162 ne
rect 1711 -1168 1720 -1162
tri 1720 -1168 1726 -1162 sw
rect 1584 -1194 1629 -1184
rect 1460 -1222 1534 -1198
rect 1402 -1226 1534 -1222
tri 1534 -1226 1562 -1198 sw
rect 1584 -1208 1586 -1194
tri 1584 -1210 1586 -1208 ne
rect 1598 -1212 1629 -1194
rect 1598 -1222 1644 -1212
rect 1711 -1183 1726 -1168
tri 1336 -1247 1348 -1235 ne
rect 1348 -1240 1358 -1235
tri 1358 -1240 1363 -1235 sw
rect 1247 -1586 1262 -1358
rect 1348 -1348 1363 -1240
rect 1402 -1282 1430 -1226
tri 1522 -1244 1540 -1226 ne
rect 1540 -1246 1562 -1226
tri 1562 -1246 1582 -1226 sw
tri 1598 -1240 1616 -1222 ne
rect 1421 -1316 1430 -1282
rect 1464 -1255 1506 -1254
rect 1464 -1289 1469 -1255
rect 1499 -1289 1506 -1255
rect 1464 -1298 1506 -1289
rect 1540 -1255 1582 -1246
rect 1540 -1289 1547 -1255
rect 1577 -1289 1582 -1255
rect 1540 -1294 1582 -1289
rect 1616 -1282 1644 -1222
tri 1689 -1235 1711 -1213 se
rect 1711 -1220 1726 -1212
tri 1711 -1235 1726 -1220 nw
tri 1683 -1241 1689 -1235 se
rect 1689 -1241 1698 -1235
rect 1402 -1326 1430 -1316
tri 1430 -1326 1454 -1302 sw
rect 1348 -1396 1364 -1348
rect 1402 -1358 1444 -1326
tri 1461 -1334 1462 -1333 sw
rect 1461 -1358 1462 -1334
tri 1464 -1335 1501 -1298 ne
rect 1501 -1326 1506 -1298
tri 1506 -1326 1532 -1300 sw
rect 1616 -1316 1625 -1282
rect 1616 -1326 1644 -1316
rect 1501 -1335 1585 -1326
tri 1501 -1354 1520 -1335 ne
rect 1520 -1354 1585 -1335
rect 1402 -1380 1462 -1358
rect 1584 -1358 1585 -1354
rect 1602 -1358 1644 -1326
rect 1584 -1380 1644 -1358
rect 1490 -1396 1507 -1382
rect 1539 -1396 1556 -1382
tri 1327 -1432 1349 -1410 se
rect 1349 -1417 1364 -1396
tri 1349 -1432 1364 -1417 nw
rect 1683 -1417 1698 -1241
tri 1698 -1248 1711 -1235 nw
rect 1784 -1316 1799 -1088
tri 1321 -1438 1327 -1432 se
rect 1327 -1438 1336 -1432
rect 1321 -1454 1336 -1438
tri 1336 -1445 1349 -1432 nw
rect 1490 -1440 1507 -1426
rect 1539 -1440 1556 -1426
tri 1683 -1432 1698 -1417 ne
tri 1698 -1432 1720 -1410 sw
rect 1321 -1490 1336 -1482
rect 1402 -1454 1462 -1440
rect 1417 -1464 1462 -1454
rect 1417 -1482 1445 -1464
tri 1321 -1505 1336 -1490 ne
tri 1336 -1505 1358 -1483 sw
rect 1402 -1492 1445 -1482
rect 1460 -1468 1462 -1464
rect 1584 -1454 1644 -1440
tri 1698 -1445 1711 -1432 ne
rect 1711 -1438 1720 -1432
tri 1720 -1438 1726 -1432 sw
rect 1584 -1464 1629 -1454
rect 1460 -1492 1534 -1468
rect 1402 -1496 1534 -1492
tri 1534 -1496 1562 -1468 sw
rect 1584 -1478 1586 -1464
tri 1584 -1480 1586 -1478 ne
rect 1598 -1482 1629 -1464
rect 1598 -1492 1644 -1482
rect 1711 -1453 1726 -1438
tri 1336 -1517 1348 -1505 ne
rect 1348 -1510 1358 -1505
tri 1358 -1510 1363 -1505 sw
rect 1247 -1856 1262 -1628
rect 1348 -1666 1363 -1510
rect 1402 -1552 1430 -1496
tri 1522 -1514 1540 -1496 ne
rect 1540 -1516 1562 -1496
tri 1562 -1516 1582 -1496 sw
tri 1598 -1510 1616 -1492 ne
rect 1421 -1586 1430 -1552
rect 1464 -1525 1506 -1524
rect 1464 -1559 1469 -1525
rect 1499 -1559 1506 -1525
rect 1464 -1568 1506 -1559
rect 1540 -1525 1582 -1516
rect 1540 -1559 1547 -1525
rect 1577 -1559 1582 -1525
rect 1540 -1564 1582 -1559
rect 1616 -1552 1644 -1492
tri 1689 -1505 1711 -1483 se
rect 1711 -1490 1726 -1482
tri 1711 -1505 1726 -1490 nw
tri 1683 -1511 1689 -1505 se
rect 1689 -1511 1698 -1505
rect 1402 -1596 1430 -1586
tri 1430 -1596 1454 -1572 sw
rect 1402 -1628 1444 -1596
tri 1461 -1604 1462 -1603 sw
rect 1461 -1628 1462 -1604
tri 1464 -1605 1501 -1568 ne
rect 1501 -1596 1506 -1568
tri 1506 -1596 1532 -1570 sw
rect 1616 -1586 1625 -1552
rect 1616 -1596 1644 -1586
rect 1501 -1605 1585 -1596
tri 1501 -1624 1520 -1605 ne
rect 1520 -1624 1585 -1605
rect 1402 -1650 1462 -1628
rect 1584 -1628 1585 -1624
rect 1602 -1628 1644 -1596
rect 1584 -1650 1644 -1628
rect 1490 -1666 1507 -1652
rect 1539 -1666 1556 -1652
tri 1327 -1702 1349 -1680 se
rect 1349 -1687 1364 -1666
tri 1349 -1702 1364 -1687 nw
rect 1683 -1687 1698 -1511
tri 1698 -1518 1711 -1505 nw
rect 1784 -1586 1799 -1358
tri 1321 -1708 1327 -1702 se
rect 1327 -1708 1336 -1702
rect 1321 -1724 1336 -1708
tri 1336 -1715 1349 -1702 nw
rect 1490 -1710 1507 -1696
rect 1539 -1710 1556 -1696
tri 1683 -1702 1698 -1687 ne
tri 1698 -1702 1720 -1680 sw
rect 1321 -1760 1336 -1752
rect 1402 -1724 1462 -1710
rect 1417 -1734 1462 -1724
rect 1417 -1752 1445 -1734
tri 1321 -1775 1336 -1760 ne
tri 1336 -1775 1358 -1753 sw
rect 1402 -1762 1445 -1752
rect 1460 -1738 1462 -1734
rect 1584 -1724 1644 -1710
tri 1698 -1715 1711 -1702 ne
rect 1711 -1708 1720 -1702
tri 1720 -1708 1726 -1702 sw
rect 1584 -1734 1629 -1724
rect 1460 -1762 1534 -1738
rect 1402 -1766 1534 -1762
tri 1534 -1766 1562 -1738 sw
rect 1584 -1748 1586 -1734
tri 1584 -1750 1586 -1748 ne
rect 1598 -1752 1629 -1734
rect 1598 -1762 1644 -1752
rect 1711 -1723 1726 -1708
tri 1336 -1787 1348 -1775 ne
rect 1348 -1780 1358 -1775
tri 1358 -1780 1363 -1775 sw
rect 1247 -2126 1262 -1898
rect 1348 -1888 1363 -1780
rect 1402 -1822 1430 -1766
tri 1522 -1784 1540 -1766 ne
rect 1540 -1786 1562 -1766
tri 1562 -1786 1582 -1766 sw
tri 1598 -1780 1616 -1762 ne
rect 1421 -1856 1430 -1822
rect 1464 -1795 1506 -1794
rect 1464 -1829 1469 -1795
rect 1499 -1829 1506 -1795
rect 1464 -1838 1506 -1829
rect 1540 -1795 1582 -1786
rect 1540 -1829 1547 -1795
rect 1577 -1829 1582 -1795
rect 1540 -1834 1582 -1829
rect 1616 -1822 1644 -1762
tri 1689 -1775 1711 -1753 se
rect 1711 -1760 1726 -1752
tri 1711 -1775 1726 -1760 nw
tri 1683 -1781 1689 -1775 se
rect 1689 -1781 1698 -1775
rect 1402 -1866 1430 -1856
tri 1430 -1866 1454 -1842 sw
rect 1348 -1936 1364 -1888
rect 1402 -1898 1444 -1866
tri 1461 -1874 1462 -1873 sw
rect 1461 -1898 1462 -1874
tri 1464 -1875 1501 -1838 ne
rect 1501 -1866 1506 -1838
tri 1506 -1866 1532 -1840 sw
rect 1616 -1856 1625 -1822
rect 1616 -1866 1644 -1856
rect 1501 -1875 1585 -1866
tri 1501 -1894 1520 -1875 ne
rect 1520 -1894 1585 -1875
rect 1402 -1920 1462 -1898
rect 1584 -1898 1585 -1894
rect 1602 -1898 1644 -1866
rect 1584 -1920 1644 -1898
rect 1490 -1936 1507 -1922
rect 1539 -1936 1556 -1922
tri 1327 -1972 1349 -1950 se
rect 1349 -1957 1364 -1936
tri 1349 -1972 1364 -1957 nw
rect 1683 -1957 1698 -1781
tri 1698 -1788 1711 -1775 nw
rect 1784 -1856 1799 -1628
tri 1321 -1978 1327 -1972 se
rect 1327 -1978 1336 -1972
rect 1321 -1994 1336 -1978
tri 1336 -1985 1349 -1972 nw
rect 1490 -1980 1507 -1966
rect 1539 -1980 1556 -1966
tri 1683 -1972 1698 -1957 ne
tri 1698 -1972 1720 -1950 sw
rect 1321 -2030 1336 -2022
rect 1402 -1994 1462 -1980
rect 1417 -2004 1462 -1994
rect 1417 -2022 1445 -2004
tri 1321 -2045 1336 -2030 ne
tri 1336 -2045 1358 -2023 sw
rect 1402 -2032 1445 -2022
rect 1460 -2008 1462 -2004
rect 1584 -1994 1644 -1980
tri 1698 -1985 1711 -1972 ne
rect 1711 -1978 1720 -1972
tri 1720 -1978 1726 -1972 sw
rect 1584 -2004 1629 -1994
rect 1460 -2032 1534 -2008
rect 1402 -2036 1534 -2032
tri 1534 -2036 1562 -2008 sw
rect 1584 -2018 1586 -2004
tri 1584 -2020 1586 -2018 ne
rect 1598 -2022 1629 -2004
rect 1598 -2032 1644 -2022
rect 1711 -1993 1726 -1978
tri 1336 -2057 1348 -2045 ne
rect 1348 -2050 1358 -2045
tri 1358 -2050 1363 -2045 sw
rect 1247 -2396 1262 -2168
rect 1348 -2206 1363 -2050
rect 1402 -2092 1430 -2036
tri 1522 -2054 1540 -2036 ne
rect 1540 -2056 1562 -2036
tri 1562 -2056 1582 -2036 sw
tri 1598 -2050 1616 -2032 ne
rect 1421 -2126 1430 -2092
rect 1464 -2065 1506 -2064
rect 1464 -2099 1469 -2065
rect 1499 -2099 1506 -2065
rect 1464 -2108 1506 -2099
rect 1540 -2065 1582 -2056
rect 1540 -2099 1547 -2065
rect 1577 -2099 1582 -2065
rect 1540 -2104 1582 -2099
rect 1616 -2092 1644 -2032
tri 1689 -2045 1711 -2023 se
rect 1711 -2030 1726 -2022
tri 1711 -2045 1726 -2030 nw
tri 1683 -2051 1689 -2045 se
rect 1689 -2051 1698 -2045
rect 1402 -2136 1430 -2126
tri 1430 -2136 1454 -2112 sw
rect 1402 -2168 1444 -2136
tri 1461 -2144 1462 -2143 sw
rect 1461 -2168 1462 -2144
tri 1464 -2145 1501 -2108 ne
rect 1501 -2136 1506 -2108
tri 1506 -2136 1532 -2110 sw
rect 1616 -2126 1625 -2092
rect 1616 -2136 1644 -2126
rect 1501 -2145 1585 -2136
tri 1501 -2164 1520 -2145 ne
rect 1520 -2164 1585 -2145
rect 1402 -2190 1462 -2168
rect 1584 -2168 1585 -2164
rect 1602 -2168 1644 -2136
rect 1584 -2190 1644 -2168
rect 1490 -2206 1507 -2192
rect 1539 -2206 1556 -2192
tri 1327 -2242 1349 -2220 se
rect 1349 -2227 1364 -2206
tri 1349 -2242 1364 -2227 nw
rect 1683 -2227 1698 -2051
tri 1698 -2058 1711 -2045 nw
rect 1784 -2126 1799 -1898
tri 1321 -2248 1327 -2242 se
rect 1327 -2248 1336 -2242
rect 1321 -2264 1336 -2248
tri 1336 -2255 1349 -2242 nw
rect 1490 -2250 1507 -2236
rect 1539 -2250 1556 -2236
tri 1683 -2242 1698 -2227 ne
tri 1698 -2242 1720 -2220 sw
rect 1321 -2300 1336 -2292
rect 1402 -2264 1462 -2250
rect 1417 -2274 1462 -2264
rect 1417 -2292 1445 -2274
tri 1321 -2315 1336 -2300 ne
tri 1336 -2315 1358 -2293 sw
rect 1402 -2302 1445 -2292
rect 1460 -2278 1462 -2274
rect 1584 -2264 1644 -2250
tri 1698 -2255 1711 -2242 ne
rect 1711 -2248 1720 -2242
tri 1720 -2248 1726 -2242 sw
rect 1584 -2274 1629 -2264
rect 1460 -2302 1534 -2278
rect 1402 -2306 1534 -2302
tri 1534 -2306 1562 -2278 sw
rect 1584 -2288 1586 -2274
tri 1584 -2290 1586 -2288 ne
rect 1598 -2292 1629 -2274
rect 1598 -2302 1644 -2292
rect 1711 -2263 1726 -2248
tri 1336 -2327 1348 -2315 ne
rect 1348 -2320 1358 -2315
tri 1358 -2320 1363 -2315 sw
rect 1247 -2524 1262 -2438
rect 1348 -2476 1363 -2320
rect 1402 -2362 1430 -2306
tri 1522 -2324 1540 -2306 ne
rect 1540 -2326 1562 -2306
tri 1562 -2326 1582 -2306 sw
tri 1598 -2320 1616 -2302 ne
rect 1421 -2396 1430 -2362
rect 1464 -2335 1506 -2334
rect 1464 -2369 1469 -2335
rect 1499 -2369 1506 -2335
rect 1464 -2378 1506 -2369
rect 1540 -2335 1582 -2326
rect 1540 -2369 1547 -2335
rect 1577 -2369 1582 -2335
rect 1540 -2374 1582 -2369
rect 1616 -2362 1644 -2302
tri 1689 -2315 1711 -2293 se
rect 1711 -2300 1726 -2292
tri 1711 -2315 1726 -2300 nw
tri 1683 -2321 1689 -2315 se
rect 1689 -2321 1698 -2315
rect 1402 -2406 1430 -2396
tri 1430 -2406 1454 -2382 sw
rect 1402 -2438 1444 -2406
tri 1461 -2414 1462 -2413 sw
rect 1461 -2438 1462 -2414
tri 1464 -2415 1501 -2378 ne
rect 1501 -2406 1506 -2378
tri 1506 -2406 1532 -2380 sw
rect 1616 -2396 1625 -2362
rect 1616 -2406 1644 -2396
rect 1501 -2415 1585 -2406
tri 1501 -2434 1520 -2415 ne
rect 1520 -2434 1585 -2415
rect 1402 -2460 1462 -2438
rect 1584 -2438 1585 -2434
rect 1602 -2438 1644 -2406
rect 1584 -2460 1644 -2438
rect 1490 -2476 1507 -2462
rect 1539 -2476 1556 -2462
rect 1683 -2476 1698 -2321
tri 1698 -2328 1711 -2315 nw
rect 1784 -2396 1799 -2168
rect 1784 -2524 1799 -2438
rect 1827 1654 1842 1844
tri 1907 1808 1929 1830 se
rect 1929 1823 1944 1892
tri 1929 1808 1944 1823 nw
rect 2263 1823 2278 1892
tri 1901 1802 1907 1808 se
rect 1907 1802 1916 1808
rect 1901 1786 1916 1802
tri 1916 1795 1929 1808 nw
rect 2070 1800 2087 1814
rect 2119 1800 2136 1814
tri 2263 1808 2278 1823 ne
tri 2278 1808 2300 1830 sw
rect 1901 1750 1916 1758
rect 1982 1786 2042 1800
rect 1997 1776 2042 1786
rect 1997 1758 2025 1776
tri 1901 1735 1916 1750 ne
tri 1916 1735 1938 1757 sw
rect 1982 1748 2025 1758
rect 2040 1772 2042 1776
rect 2164 1786 2224 1800
tri 2278 1795 2291 1808 ne
rect 2291 1802 2300 1808
tri 2300 1802 2306 1808 sw
rect 2164 1776 2209 1786
rect 2040 1748 2114 1772
rect 1982 1744 2114 1748
tri 2114 1744 2142 1772 sw
rect 2164 1762 2166 1776
tri 2164 1760 2166 1762 ne
rect 2178 1758 2209 1776
rect 2178 1748 2224 1758
rect 2291 1787 2306 1802
tri 1916 1723 1928 1735 ne
rect 1928 1730 1938 1735
tri 1938 1730 1943 1735 sw
rect 1827 1384 1842 1612
rect 1928 1574 1943 1730
rect 1982 1688 2010 1744
tri 2102 1726 2120 1744 ne
rect 2120 1724 2142 1744
tri 2142 1724 2162 1744 sw
tri 2178 1730 2196 1748 ne
rect 2001 1654 2010 1688
rect 2044 1715 2086 1716
rect 2044 1681 2049 1715
rect 2079 1681 2086 1715
rect 2044 1672 2086 1681
rect 2120 1715 2162 1724
rect 2120 1681 2127 1715
rect 2157 1681 2162 1715
rect 2120 1676 2162 1681
rect 2196 1688 2224 1748
tri 2269 1735 2291 1757 se
rect 2291 1750 2306 1758
tri 2291 1735 2306 1750 nw
tri 2263 1729 2269 1735 se
rect 2269 1729 2278 1735
rect 1982 1644 2010 1654
tri 2010 1644 2034 1668 sw
rect 1982 1612 2024 1644
tri 2041 1636 2042 1637 sw
rect 2041 1612 2042 1636
tri 2044 1635 2081 1672 ne
rect 2081 1644 2086 1672
tri 2086 1644 2112 1670 sw
rect 2196 1654 2205 1688
rect 2196 1644 2224 1654
rect 2081 1635 2165 1644
tri 2081 1616 2100 1635 ne
rect 2100 1616 2165 1635
rect 1982 1590 2042 1612
rect 2164 1612 2165 1616
rect 2182 1612 2224 1644
rect 2164 1590 2224 1612
rect 2070 1574 2087 1588
rect 2119 1574 2136 1588
tri 1907 1538 1929 1560 se
rect 1929 1553 1944 1574
tri 1929 1538 1944 1553 nw
rect 2263 1553 2278 1729
tri 2278 1722 2291 1735 nw
rect 2364 1654 2379 1844
tri 1901 1532 1907 1538 se
rect 1907 1532 1916 1538
rect 1901 1516 1916 1532
tri 1916 1525 1929 1538 nw
rect 2070 1530 2087 1544
rect 2119 1530 2136 1544
tri 2263 1538 2278 1553 ne
tri 2278 1538 2300 1560 sw
rect 1901 1480 1916 1488
rect 1982 1516 2042 1530
rect 1997 1506 2042 1516
rect 1997 1488 2025 1506
tri 1901 1465 1916 1480 ne
tri 1916 1465 1938 1487 sw
rect 1982 1478 2025 1488
rect 2040 1502 2042 1506
rect 2164 1516 2224 1530
tri 2278 1525 2291 1538 ne
rect 2291 1532 2300 1538
tri 2300 1532 2306 1538 sw
rect 2164 1506 2209 1516
rect 2040 1478 2114 1502
rect 1982 1474 2114 1478
tri 2114 1474 2142 1502 sw
rect 2164 1492 2166 1506
tri 2164 1490 2166 1492 ne
rect 2178 1488 2209 1506
rect 2178 1478 2224 1488
rect 2291 1517 2306 1532
tri 1916 1453 1928 1465 ne
rect 1928 1460 1938 1465
tri 1938 1460 1943 1465 sw
rect 1827 1114 1842 1342
rect 1928 1352 1943 1460
rect 1982 1418 2010 1474
tri 2102 1456 2120 1474 ne
rect 2120 1454 2142 1474
tri 2142 1454 2162 1474 sw
tri 2178 1460 2196 1478 ne
rect 2001 1384 2010 1418
rect 2044 1445 2086 1446
rect 2044 1411 2049 1445
rect 2079 1411 2086 1445
rect 2044 1402 2086 1411
rect 2120 1445 2162 1454
rect 2120 1411 2127 1445
rect 2157 1411 2162 1445
rect 2120 1406 2162 1411
rect 2196 1418 2224 1478
tri 2269 1465 2291 1487 se
rect 2291 1480 2306 1488
tri 2291 1465 2306 1480 nw
tri 2263 1459 2269 1465 se
rect 2269 1459 2278 1465
rect 1982 1374 2010 1384
tri 2010 1374 2034 1398 sw
rect 1928 1304 1944 1352
rect 1982 1342 2024 1374
tri 2041 1366 2042 1367 sw
rect 2041 1342 2042 1366
tri 2044 1365 2081 1402 ne
rect 2081 1374 2086 1402
tri 2086 1374 2112 1400 sw
rect 2196 1384 2205 1418
rect 2196 1374 2224 1384
rect 2081 1365 2165 1374
tri 2081 1346 2100 1365 ne
rect 2100 1346 2165 1365
rect 1982 1320 2042 1342
rect 2164 1342 2165 1346
rect 2182 1342 2224 1374
rect 2164 1320 2224 1342
rect 2070 1304 2087 1318
rect 2119 1304 2136 1318
tri 1907 1268 1929 1290 se
rect 1929 1283 1944 1304
tri 1929 1268 1944 1283 nw
rect 2263 1283 2278 1459
tri 2278 1452 2291 1465 nw
rect 2364 1384 2379 1612
tri 1901 1262 1907 1268 se
rect 1907 1262 1916 1268
rect 1901 1246 1916 1262
tri 1916 1255 1929 1268 nw
rect 2070 1260 2087 1274
rect 2119 1260 2136 1274
tri 2263 1268 2278 1283 ne
tri 2278 1268 2300 1290 sw
rect 1901 1210 1916 1218
rect 1982 1246 2042 1260
rect 1997 1236 2042 1246
rect 1997 1218 2025 1236
tri 1901 1195 1916 1210 ne
tri 1916 1195 1938 1217 sw
rect 1982 1208 2025 1218
rect 2040 1232 2042 1236
rect 2164 1246 2224 1260
tri 2278 1255 2291 1268 ne
rect 2291 1262 2300 1268
tri 2300 1262 2306 1268 sw
rect 2164 1236 2209 1246
rect 2040 1208 2114 1232
rect 1982 1204 2114 1208
tri 2114 1204 2142 1232 sw
rect 2164 1222 2166 1236
tri 2164 1220 2166 1222 ne
rect 2178 1218 2209 1236
rect 2178 1208 2224 1218
rect 2291 1247 2306 1262
tri 1916 1183 1928 1195 ne
rect 1928 1190 1938 1195
tri 1938 1190 1943 1195 sw
rect 1827 844 1842 1072
rect 1928 1034 1943 1190
rect 1982 1148 2010 1204
tri 2102 1186 2120 1204 ne
rect 2120 1184 2142 1204
tri 2142 1184 2162 1204 sw
tri 2178 1190 2196 1208 ne
rect 2001 1114 2010 1148
rect 2044 1175 2086 1176
rect 2044 1141 2049 1175
rect 2079 1141 2086 1175
rect 2044 1132 2086 1141
rect 2120 1175 2162 1184
rect 2120 1141 2127 1175
rect 2157 1141 2162 1175
rect 2120 1136 2162 1141
rect 2196 1148 2224 1208
tri 2269 1195 2291 1217 se
rect 2291 1210 2306 1218
tri 2291 1195 2306 1210 nw
tri 2263 1189 2269 1195 se
rect 2269 1189 2278 1195
rect 1982 1104 2010 1114
tri 2010 1104 2034 1128 sw
rect 1982 1072 2024 1104
tri 2041 1096 2042 1097 sw
rect 2041 1072 2042 1096
tri 2044 1095 2081 1132 ne
rect 2081 1104 2086 1132
tri 2086 1104 2112 1130 sw
rect 2196 1114 2205 1148
rect 2196 1104 2224 1114
rect 2081 1095 2165 1104
tri 2081 1076 2100 1095 ne
rect 2100 1076 2165 1095
rect 1982 1050 2042 1072
rect 2164 1072 2165 1076
rect 2182 1072 2224 1104
rect 2164 1050 2224 1072
rect 2070 1034 2087 1048
rect 2119 1034 2136 1048
tri 1907 998 1929 1020 se
rect 1929 1013 1944 1034
tri 1929 998 1944 1013 nw
rect 2263 1013 2278 1189
tri 2278 1182 2291 1195 nw
rect 2364 1114 2379 1342
tri 1901 992 1907 998 se
rect 1907 992 1916 998
rect 1901 976 1916 992
tri 1916 985 1929 998 nw
rect 2070 990 2087 1004
rect 2119 990 2136 1004
tri 2263 998 2278 1013 ne
tri 2278 998 2300 1020 sw
rect 1901 940 1916 948
rect 1982 976 2042 990
rect 1997 966 2042 976
rect 1997 948 2025 966
tri 1901 925 1916 940 ne
tri 1916 925 1938 947 sw
rect 1982 938 2025 948
rect 2040 962 2042 966
rect 2164 976 2224 990
tri 2278 985 2291 998 ne
rect 2291 992 2300 998
tri 2300 992 2306 998 sw
rect 2164 966 2209 976
rect 2040 938 2114 962
rect 1982 934 2114 938
tri 2114 934 2142 962 sw
rect 2164 952 2166 966
tri 2164 950 2166 952 ne
rect 2178 948 2209 966
rect 2178 938 2224 948
rect 2291 977 2306 992
tri 1916 913 1928 925 ne
rect 1928 920 1938 925
tri 1938 920 1943 925 sw
rect 1827 574 1842 802
rect 1928 812 1943 920
rect 1982 878 2010 934
tri 2102 916 2120 934 ne
rect 2120 914 2142 934
tri 2142 914 2162 934 sw
tri 2178 920 2196 938 ne
rect 2001 844 2010 878
rect 2044 905 2086 906
rect 2044 871 2049 905
rect 2079 871 2086 905
rect 2044 862 2086 871
rect 2120 905 2162 914
rect 2120 871 2127 905
rect 2157 871 2162 905
rect 2120 866 2162 871
rect 2196 878 2224 938
tri 2269 925 2291 947 se
rect 2291 940 2306 948
tri 2291 925 2306 940 nw
tri 2263 919 2269 925 se
rect 2269 919 2278 925
rect 1982 834 2010 844
tri 2010 834 2034 858 sw
rect 1928 764 1944 812
rect 1982 802 2024 834
tri 2041 826 2042 827 sw
rect 2041 802 2042 826
tri 2044 825 2081 862 ne
rect 2081 834 2086 862
tri 2086 834 2112 860 sw
rect 2196 844 2205 878
rect 2196 834 2224 844
rect 2081 825 2165 834
tri 2081 806 2100 825 ne
rect 2100 806 2165 825
rect 1982 780 2042 802
rect 2164 802 2165 806
rect 2182 802 2224 834
rect 2164 780 2224 802
rect 2070 764 2087 778
rect 2119 764 2136 778
tri 1907 728 1929 750 se
rect 1929 743 1944 764
tri 1929 728 1944 743 nw
rect 2263 743 2278 919
tri 2278 912 2291 925 nw
rect 2364 844 2379 1072
tri 1901 722 1907 728 se
rect 1907 722 1916 728
rect 1901 706 1916 722
tri 1916 715 1929 728 nw
rect 2070 720 2087 734
rect 2119 720 2136 734
tri 2263 728 2278 743 ne
tri 2278 728 2300 750 sw
rect 1901 670 1916 678
rect 1982 706 2042 720
rect 1997 696 2042 706
rect 1997 678 2025 696
tri 1901 655 1916 670 ne
tri 1916 655 1938 677 sw
rect 1982 668 2025 678
rect 2040 692 2042 696
rect 2164 706 2224 720
tri 2278 715 2291 728 ne
rect 2291 722 2300 728
tri 2300 722 2306 728 sw
rect 2164 696 2209 706
rect 2040 668 2114 692
rect 1982 664 2114 668
tri 2114 664 2142 692 sw
rect 2164 682 2166 696
tri 2164 680 2166 682 ne
rect 2178 678 2209 696
rect 2178 668 2224 678
rect 2291 707 2306 722
tri 1916 643 1928 655 ne
rect 1928 650 1938 655
tri 1938 650 1943 655 sw
rect 1827 304 1842 532
rect 1928 494 1943 650
rect 1982 608 2010 664
tri 2102 646 2120 664 ne
rect 2120 644 2142 664
tri 2142 644 2162 664 sw
tri 2178 650 2196 668 ne
rect 2001 574 2010 608
rect 2044 635 2086 636
rect 2044 601 2049 635
rect 2079 601 2086 635
rect 2044 592 2086 601
rect 2120 635 2162 644
rect 2120 601 2127 635
rect 2157 601 2162 635
rect 2120 596 2162 601
rect 2196 608 2224 668
tri 2269 655 2291 677 se
rect 2291 670 2306 678
tri 2291 655 2306 670 nw
tri 2263 649 2269 655 se
rect 2269 649 2278 655
rect 1982 564 2010 574
tri 2010 564 2034 588 sw
rect 1982 532 2024 564
tri 2041 556 2042 557 sw
rect 2041 532 2042 556
tri 2044 555 2081 592 ne
rect 2081 564 2086 592
tri 2086 564 2112 590 sw
rect 2196 574 2205 608
rect 2196 564 2224 574
rect 2081 555 2165 564
tri 2081 536 2100 555 ne
rect 2100 536 2165 555
rect 1982 510 2042 532
rect 2164 532 2165 536
rect 2182 532 2224 564
rect 2164 510 2224 532
rect 2070 494 2087 508
rect 2119 494 2136 508
tri 1907 458 1929 480 se
rect 1929 473 1944 494
tri 1929 458 1944 473 nw
rect 2263 473 2278 649
tri 2278 642 2291 655 nw
rect 2364 574 2379 802
tri 1901 452 1907 458 se
rect 1907 452 1916 458
rect 1901 436 1916 452
tri 1916 445 1929 458 nw
rect 2070 450 2087 464
rect 2119 450 2136 464
tri 2263 458 2278 473 ne
tri 2278 458 2300 480 sw
rect 1901 400 1916 408
rect 1982 436 2042 450
rect 1997 426 2042 436
rect 1997 408 2025 426
tri 1901 385 1916 400 ne
tri 1916 385 1938 407 sw
rect 1982 398 2025 408
rect 2040 422 2042 426
rect 2164 436 2224 450
tri 2278 445 2291 458 ne
rect 2291 452 2300 458
tri 2300 452 2306 458 sw
rect 2164 426 2209 436
rect 2040 398 2114 422
rect 1982 394 2114 398
tri 2114 394 2142 422 sw
rect 2164 412 2166 426
tri 2164 410 2166 412 ne
rect 2178 408 2209 426
rect 2178 398 2224 408
rect 2291 437 2306 452
tri 1916 373 1928 385 ne
rect 1928 380 1938 385
tri 1938 380 1943 385 sw
rect 1827 34 1842 262
rect 1928 272 1943 380
rect 1982 338 2010 394
tri 2102 376 2120 394 ne
rect 2120 374 2142 394
tri 2142 374 2162 394 sw
tri 2178 380 2196 398 ne
rect 2001 304 2010 338
rect 2044 365 2086 366
rect 2044 331 2049 365
rect 2079 331 2086 365
rect 2044 322 2086 331
rect 2120 365 2162 374
rect 2120 331 2127 365
rect 2157 331 2162 365
rect 2120 326 2162 331
rect 2196 338 2224 398
tri 2269 385 2291 407 se
rect 2291 400 2306 408
tri 2291 385 2306 400 nw
tri 2263 379 2269 385 se
rect 2269 379 2278 385
rect 1982 294 2010 304
tri 2010 294 2034 318 sw
rect 1928 224 1944 272
rect 1982 262 2024 294
tri 2041 286 2042 287 sw
rect 2041 262 2042 286
tri 2044 285 2081 322 ne
rect 2081 294 2086 322
tri 2086 294 2112 320 sw
rect 2196 304 2205 338
rect 2196 294 2224 304
rect 2081 285 2165 294
tri 2081 266 2100 285 ne
rect 2100 266 2165 285
rect 1982 240 2042 262
rect 2164 262 2165 266
rect 2182 262 2224 294
rect 2164 240 2224 262
rect 2070 224 2087 238
rect 2119 224 2136 238
tri 1907 188 1929 210 se
rect 1929 203 1944 224
tri 1929 188 1944 203 nw
rect 2263 203 2278 379
tri 2278 372 2291 385 nw
rect 2364 304 2379 532
tri 1901 182 1907 188 se
rect 1907 182 1916 188
rect 1901 166 1916 182
tri 1916 175 1929 188 nw
rect 2070 180 2087 194
rect 2119 180 2136 194
tri 2263 188 2278 203 ne
tri 2278 188 2300 210 sw
rect 1901 130 1916 138
rect 1982 166 2042 180
rect 1997 156 2042 166
rect 1997 138 2025 156
tri 1901 115 1916 130 ne
tri 1916 115 1938 137 sw
rect 1982 128 2025 138
rect 2040 152 2042 156
rect 2164 166 2224 180
tri 2278 175 2291 188 ne
rect 2291 182 2300 188
tri 2300 182 2306 188 sw
rect 2164 156 2209 166
rect 2040 128 2114 152
rect 1982 124 2114 128
tri 2114 124 2142 152 sw
rect 2164 142 2166 156
tri 2164 140 2166 142 ne
rect 2178 138 2209 156
rect 2178 128 2224 138
rect 2291 167 2306 182
tri 1916 103 1928 115 ne
rect 1928 110 1938 115
tri 1938 110 1943 115 sw
rect 1827 -236 1842 -8
rect 1928 -46 1943 110
rect 1982 68 2010 124
tri 2102 106 2120 124 ne
rect 2120 104 2142 124
tri 2142 104 2162 124 sw
tri 2178 110 2196 128 ne
rect 2001 34 2010 68
rect 2044 95 2086 96
rect 2044 61 2049 95
rect 2079 61 2086 95
rect 2044 52 2086 61
rect 2120 95 2162 104
rect 2120 61 2127 95
rect 2157 61 2162 95
rect 2120 56 2162 61
rect 2196 68 2224 128
tri 2269 115 2291 137 se
rect 2291 130 2306 138
tri 2291 115 2306 130 nw
tri 2263 109 2269 115 se
rect 2269 109 2278 115
rect 1982 24 2010 34
tri 2010 24 2034 48 sw
rect 1982 -8 2024 24
tri 2041 16 2042 17 sw
rect 2041 -8 2042 16
tri 2044 15 2081 52 ne
rect 2081 24 2086 52
tri 2086 24 2112 50 sw
rect 2196 34 2205 68
rect 2196 24 2224 34
rect 2081 15 2165 24
tri 2081 -4 2100 15 ne
rect 2100 -4 2165 15
rect 1982 -30 2042 -8
rect 2164 -8 2165 -4
rect 2182 -8 2224 24
rect 2164 -30 2224 -8
rect 2070 -46 2087 -32
rect 2119 -46 2136 -32
tri 1907 -82 1929 -60 se
rect 1929 -67 1944 -46
tri 1929 -82 1944 -67 nw
rect 2263 -67 2278 109
tri 2278 102 2291 115 nw
rect 2364 34 2379 262
tri 1901 -88 1907 -82 se
rect 1907 -88 1916 -82
rect 1901 -104 1916 -88
tri 1916 -95 1929 -82 nw
rect 2070 -90 2087 -76
rect 2119 -90 2136 -76
tri 2263 -82 2278 -67 ne
tri 2278 -82 2300 -60 sw
rect 1901 -140 1916 -132
rect 1982 -104 2042 -90
rect 1997 -114 2042 -104
rect 1997 -132 2025 -114
tri 1901 -155 1916 -140 ne
tri 1916 -155 1938 -133 sw
rect 1982 -142 2025 -132
rect 2040 -118 2042 -114
rect 2164 -104 2224 -90
tri 2278 -95 2291 -82 ne
rect 2291 -88 2300 -82
tri 2300 -88 2306 -82 sw
rect 2164 -114 2209 -104
rect 2040 -142 2114 -118
rect 1982 -146 2114 -142
tri 2114 -146 2142 -118 sw
rect 2164 -128 2166 -114
tri 2164 -130 2166 -128 ne
rect 2178 -132 2209 -114
rect 2178 -142 2224 -132
rect 2291 -103 2306 -88
tri 1916 -167 1928 -155 ne
rect 1928 -160 1938 -155
tri 1938 -160 1943 -155 sw
rect 1827 -506 1842 -278
rect 1928 -268 1943 -160
rect 1982 -202 2010 -146
tri 2102 -164 2120 -146 ne
rect 2120 -166 2142 -146
tri 2142 -166 2162 -146 sw
tri 2178 -160 2196 -142 ne
rect 2001 -236 2010 -202
rect 2044 -175 2086 -174
rect 2044 -209 2049 -175
rect 2079 -209 2086 -175
rect 2044 -218 2086 -209
rect 2120 -175 2162 -166
rect 2120 -209 2127 -175
rect 2157 -209 2162 -175
rect 2120 -214 2162 -209
rect 2196 -202 2224 -142
tri 2269 -155 2291 -133 se
rect 2291 -140 2306 -132
tri 2291 -155 2306 -140 nw
tri 2263 -161 2269 -155 se
rect 2269 -161 2278 -155
rect 1982 -246 2010 -236
tri 2010 -246 2034 -222 sw
rect 1928 -316 1944 -268
rect 1982 -278 2024 -246
tri 2041 -254 2042 -253 sw
rect 2041 -278 2042 -254
tri 2044 -255 2081 -218 ne
rect 2081 -246 2086 -218
tri 2086 -246 2112 -220 sw
rect 2196 -236 2205 -202
rect 2196 -246 2224 -236
rect 2081 -255 2165 -246
tri 2081 -274 2100 -255 ne
rect 2100 -274 2165 -255
rect 1982 -300 2042 -278
rect 2164 -278 2165 -274
rect 2182 -278 2224 -246
rect 2164 -300 2224 -278
rect 2070 -316 2087 -302
rect 2119 -316 2136 -302
tri 1907 -352 1929 -330 se
rect 1929 -337 1944 -316
tri 1929 -352 1944 -337 nw
rect 2263 -337 2278 -161
tri 2278 -168 2291 -155 nw
rect 2364 -236 2379 -8
tri 1901 -358 1907 -352 se
rect 1907 -358 1916 -352
rect 1901 -374 1916 -358
tri 1916 -365 1929 -352 nw
rect 2070 -360 2087 -346
rect 2119 -360 2136 -346
tri 2263 -352 2278 -337 ne
tri 2278 -352 2300 -330 sw
rect 1901 -410 1916 -402
rect 1982 -374 2042 -360
rect 1997 -384 2042 -374
rect 1997 -402 2025 -384
tri 1901 -425 1916 -410 ne
tri 1916 -425 1938 -403 sw
rect 1982 -412 2025 -402
rect 2040 -388 2042 -384
rect 2164 -374 2224 -360
tri 2278 -365 2291 -352 ne
rect 2291 -358 2300 -352
tri 2300 -358 2306 -352 sw
rect 2164 -384 2209 -374
rect 2040 -412 2114 -388
rect 1982 -416 2114 -412
tri 2114 -416 2142 -388 sw
rect 2164 -398 2166 -384
tri 2164 -400 2166 -398 ne
rect 2178 -402 2209 -384
rect 2178 -412 2224 -402
rect 2291 -373 2306 -358
tri 1916 -437 1928 -425 ne
rect 1928 -430 1938 -425
tri 1938 -430 1943 -425 sw
rect 1827 -776 1842 -548
rect 1928 -586 1943 -430
rect 1982 -472 2010 -416
tri 2102 -434 2120 -416 ne
rect 2120 -436 2142 -416
tri 2142 -436 2162 -416 sw
tri 2178 -430 2196 -412 ne
rect 2001 -506 2010 -472
rect 2044 -445 2086 -444
rect 2044 -479 2049 -445
rect 2079 -479 2086 -445
rect 2044 -488 2086 -479
rect 2120 -445 2162 -436
rect 2120 -479 2127 -445
rect 2157 -479 2162 -445
rect 2120 -484 2162 -479
rect 2196 -472 2224 -412
tri 2269 -425 2291 -403 se
rect 2291 -410 2306 -402
tri 2291 -425 2306 -410 nw
tri 2263 -431 2269 -425 se
rect 2269 -431 2278 -425
rect 1982 -516 2010 -506
tri 2010 -516 2034 -492 sw
rect 1982 -548 2024 -516
tri 2041 -524 2042 -523 sw
rect 2041 -548 2042 -524
tri 2044 -525 2081 -488 ne
rect 2081 -516 2086 -488
tri 2086 -516 2112 -490 sw
rect 2196 -506 2205 -472
rect 2196 -516 2224 -506
rect 2081 -525 2165 -516
tri 2081 -544 2100 -525 ne
rect 2100 -544 2165 -525
rect 1982 -570 2042 -548
rect 2164 -548 2165 -544
rect 2182 -548 2224 -516
rect 2164 -570 2224 -548
rect 2070 -586 2087 -572
rect 2119 -586 2136 -572
tri 1907 -622 1929 -600 se
rect 1929 -607 1944 -586
tri 1929 -622 1944 -607 nw
rect 2263 -607 2278 -431
tri 2278 -438 2291 -425 nw
rect 2364 -506 2379 -278
tri 1901 -628 1907 -622 se
rect 1907 -628 1916 -622
rect 1901 -644 1916 -628
tri 1916 -635 1929 -622 nw
rect 2070 -630 2087 -616
rect 2119 -630 2136 -616
tri 2263 -622 2278 -607 ne
tri 2278 -622 2300 -600 sw
rect 1901 -680 1916 -672
rect 1982 -644 2042 -630
rect 1997 -654 2042 -644
rect 1997 -672 2025 -654
tri 1901 -695 1916 -680 ne
tri 1916 -695 1938 -673 sw
rect 1982 -682 2025 -672
rect 2040 -658 2042 -654
rect 2164 -644 2224 -630
tri 2278 -635 2291 -622 ne
rect 2291 -628 2300 -622
tri 2300 -628 2306 -622 sw
rect 2164 -654 2209 -644
rect 2040 -682 2114 -658
rect 1982 -686 2114 -682
tri 2114 -686 2142 -658 sw
rect 2164 -668 2166 -654
tri 2164 -670 2166 -668 ne
rect 2178 -672 2209 -654
rect 2178 -682 2224 -672
rect 2291 -643 2306 -628
tri 1916 -707 1928 -695 ne
rect 1928 -700 1938 -695
tri 1938 -700 1943 -695 sw
rect 1827 -1046 1842 -818
rect 1928 -808 1943 -700
rect 1982 -742 2010 -686
tri 2102 -704 2120 -686 ne
rect 2120 -706 2142 -686
tri 2142 -706 2162 -686 sw
tri 2178 -700 2196 -682 ne
rect 2001 -776 2010 -742
rect 2044 -715 2086 -714
rect 2044 -749 2049 -715
rect 2079 -749 2086 -715
rect 2044 -758 2086 -749
rect 2120 -715 2162 -706
rect 2120 -749 2127 -715
rect 2157 -749 2162 -715
rect 2120 -754 2162 -749
rect 2196 -742 2224 -682
tri 2269 -695 2291 -673 se
rect 2291 -680 2306 -672
tri 2291 -695 2306 -680 nw
tri 2263 -701 2269 -695 se
rect 2269 -701 2278 -695
rect 1982 -786 2010 -776
tri 2010 -786 2034 -762 sw
rect 1928 -856 1944 -808
rect 1982 -818 2024 -786
tri 2041 -794 2042 -793 sw
rect 2041 -818 2042 -794
tri 2044 -795 2081 -758 ne
rect 2081 -786 2086 -758
tri 2086 -786 2112 -760 sw
rect 2196 -776 2205 -742
rect 2196 -786 2224 -776
rect 2081 -795 2165 -786
tri 2081 -814 2100 -795 ne
rect 2100 -814 2165 -795
rect 1982 -840 2042 -818
rect 2164 -818 2165 -814
rect 2182 -818 2224 -786
rect 2164 -840 2224 -818
rect 2070 -856 2087 -842
rect 2119 -856 2136 -842
tri 1907 -892 1929 -870 se
rect 1929 -877 1944 -856
tri 1929 -892 1944 -877 nw
rect 2263 -877 2278 -701
tri 2278 -708 2291 -695 nw
rect 2364 -776 2379 -548
tri 1901 -898 1907 -892 se
rect 1907 -898 1916 -892
rect 1901 -914 1916 -898
tri 1916 -905 1929 -892 nw
rect 2070 -900 2087 -886
rect 2119 -900 2136 -886
tri 2263 -892 2278 -877 ne
tri 2278 -892 2300 -870 sw
rect 1901 -950 1916 -942
rect 1982 -914 2042 -900
rect 1997 -924 2042 -914
rect 1997 -942 2025 -924
tri 1901 -965 1916 -950 ne
tri 1916 -965 1938 -943 sw
rect 1982 -952 2025 -942
rect 2040 -928 2042 -924
rect 2164 -914 2224 -900
tri 2278 -905 2291 -892 ne
rect 2291 -898 2300 -892
tri 2300 -898 2306 -892 sw
rect 2164 -924 2209 -914
rect 2040 -952 2114 -928
rect 1982 -956 2114 -952
tri 2114 -956 2142 -928 sw
rect 2164 -938 2166 -924
tri 2164 -940 2166 -938 ne
rect 2178 -942 2209 -924
rect 2178 -952 2224 -942
rect 2291 -913 2306 -898
tri 1916 -977 1928 -965 ne
rect 1928 -970 1938 -965
tri 1938 -970 1943 -965 sw
rect 1827 -1316 1842 -1088
rect 1928 -1126 1943 -970
rect 1982 -1012 2010 -956
tri 2102 -974 2120 -956 ne
rect 2120 -976 2142 -956
tri 2142 -976 2162 -956 sw
tri 2178 -970 2196 -952 ne
rect 2001 -1046 2010 -1012
rect 2044 -985 2086 -984
rect 2044 -1019 2049 -985
rect 2079 -1019 2086 -985
rect 2044 -1028 2086 -1019
rect 2120 -985 2162 -976
rect 2120 -1019 2127 -985
rect 2157 -1019 2162 -985
rect 2120 -1024 2162 -1019
rect 2196 -1012 2224 -952
tri 2269 -965 2291 -943 se
rect 2291 -950 2306 -942
tri 2291 -965 2306 -950 nw
tri 2263 -971 2269 -965 se
rect 2269 -971 2278 -965
rect 1982 -1056 2010 -1046
tri 2010 -1056 2034 -1032 sw
rect 1982 -1088 2024 -1056
tri 2041 -1064 2042 -1063 sw
rect 2041 -1088 2042 -1064
tri 2044 -1065 2081 -1028 ne
rect 2081 -1056 2086 -1028
tri 2086 -1056 2112 -1030 sw
rect 2196 -1046 2205 -1012
rect 2196 -1056 2224 -1046
rect 2081 -1065 2165 -1056
tri 2081 -1084 2100 -1065 ne
rect 2100 -1084 2165 -1065
rect 1982 -1110 2042 -1088
rect 2164 -1088 2165 -1084
rect 2182 -1088 2224 -1056
rect 2164 -1110 2224 -1088
rect 2070 -1126 2087 -1112
rect 2119 -1126 2136 -1112
tri 1907 -1162 1929 -1140 se
rect 1929 -1147 1944 -1126
tri 1929 -1162 1944 -1147 nw
rect 2263 -1147 2278 -971
tri 2278 -978 2291 -965 nw
rect 2364 -1046 2379 -818
tri 1901 -1168 1907 -1162 se
rect 1907 -1168 1916 -1162
rect 1901 -1184 1916 -1168
tri 1916 -1175 1929 -1162 nw
rect 2070 -1170 2087 -1156
rect 2119 -1170 2136 -1156
tri 2263 -1162 2278 -1147 ne
tri 2278 -1162 2300 -1140 sw
rect 1901 -1220 1916 -1212
rect 1982 -1184 2042 -1170
rect 1997 -1194 2042 -1184
rect 1997 -1212 2025 -1194
tri 1901 -1235 1916 -1220 ne
tri 1916 -1235 1938 -1213 sw
rect 1982 -1222 2025 -1212
rect 2040 -1198 2042 -1194
rect 2164 -1184 2224 -1170
tri 2278 -1175 2291 -1162 ne
rect 2291 -1168 2300 -1162
tri 2300 -1168 2306 -1162 sw
rect 2164 -1194 2209 -1184
rect 2040 -1222 2114 -1198
rect 1982 -1226 2114 -1222
tri 2114 -1226 2142 -1198 sw
rect 2164 -1208 2166 -1194
tri 2164 -1210 2166 -1208 ne
rect 2178 -1212 2209 -1194
rect 2178 -1222 2224 -1212
rect 2291 -1183 2306 -1168
tri 1916 -1247 1928 -1235 ne
rect 1928 -1240 1938 -1235
tri 1938 -1240 1943 -1235 sw
rect 1827 -1586 1842 -1358
rect 1928 -1348 1943 -1240
rect 1982 -1282 2010 -1226
tri 2102 -1244 2120 -1226 ne
rect 2120 -1246 2142 -1226
tri 2142 -1246 2162 -1226 sw
tri 2178 -1240 2196 -1222 ne
rect 2001 -1316 2010 -1282
rect 2044 -1255 2086 -1254
rect 2044 -1289 2049 -1255
rect 2079 -1289 2086 -1255
rect 2044 -1298 2086 -1289
rect 2120 -1255 2162 -1246
rect 2120 -1289 2127 -1255
rect 2157 -1289 2162 -1255
rect 2120 -1294 2162 -1289
rect 2196 -1282 2224 -1222
tri 2269 -1235 2291 -1213 se
rect 2291 -1220 2306 -1212
tri 2291 -1235 2306 -1220 nw
tri 2263 -1241 2269 -1235 se
rect 2269 -1241 2278 -1235
rect 1982 -1326 2010 -1316
tri 2010 -1326 2034 -1302 sw
rect 1928 -1396 1944 -1348
rect 1982 -1358 2024 -1326
tri 2041 -1334 2042 -1333 sw
rect 2041 -1358 2042 -1334
tri 2044 -1335 2081 -1298 ne
rect 2081 -1326 2086 -1298
tri 2086 -1326 2112 -1300 sw
rect 2196 -1316 2205 -1282
rect 2196 -1326 2224 -1316
rect 2081 -1335 2165 -1326
tri 2081 -1354 2100 -1335 ne
rect 2100 -1354 2165 -1335
rect 1982 -1380 2042 -1358
rect 2164 -1358 2165 -1354
rect 2182 -1358 2224 -1326
rect 2164 -1380 2224 -1358
rect 2070 -1396 2087 -1382
rect 2119 -1396 2136 -1382
tri 1907 -1432 1929 -1410 se
rect 1929 -1417 1944 -1396
tri 1929 -1432 1944 -1417 nw
rect 2263 -1417 2278 -1241
tri 2278 -1248 2291 -1235 nw
rect 2364 -1316 2379 -1088
tri 1901 -1438 1907 -1432 se
rect 1907 -1438 1916 -1432
rect 1901 -1454 1916 -1438
tri 1916 -1445 1929 -1432 nw
rect 2070 -1440 2087 -1426
rect 2119 -1440 2136 -1426
tri 2263 -1432 2278 -1417 ne
tri 2278 -1432 2300 -1410 sw
rect 1901 -1490 1916 -1482
rect 1982 -1454 2042 -1440
rect 1997 -1464 2042 -1454
rect 1997 -1482 2025 -1464
tri 1901 -1505 1916 -1490 ne
tri 1916 -1505 1938 -1483 sw
rect 1982 -1492 2025 -1482
rect 2040 -1468 2042 -1464
rect 2164 -1454 2224 -1440
tri 2278 -1445 2291 -1432 ne
rect 2291 -1438 2300 -1432
tri 2300 -1438 2306 -1432 sw
rect 2164 -1464 2209 -1454
rect 2040 -1492 2114 -1468
rect 1982 -1496 2114 -1492
tri 2114 -1496 2142 -1468 sw
rect 2164 -1478 2166 -1464
tri 2164 -1480 2166 -1478 ne
rect 2178 -1482 2209 -1464
rect 2178 -1492 2224 -1482
rect 2291 -1453 2306 -1438
tri 1916 -1517 1928 -1505 ne
rect 1928 -1510 1938 -1505
tri 1938 -1510 1943 -1505 sw
rect 1827 -1856 1842 -1628
rect 1928 -1666 1943 -1510
rect 1982 -1552 2010 -1496
tri 2102 -1514 2120 -1496 ne
rect 2120 -1516 2142 -1496
tri 2142 -1516 2162 -1496 sw
tri 2178 -1510 2196 -1492 ne
rect 2001 -1586 2010 -1552
rect 2044 -1525 2086 -1524
rect 2044 -1559 2049 -1525
rect 2079 -1559 2086 -1525
rect 2044 -1568 2086 -1559
rect 2120 -1525 2162 -1516
rect 2120 -1559 2127 -1525
rect 2157 -1559 2162 -1525
rect 2120 -1564 2162 -1559
rect 2196 -1552 2224 -1492
tri 2269 -1505 2291 -1483 se
rect 2291 -1490 2306 -1482
tri 2291 -1505 2306 -1490 nw
tri 2263 -1511 2269 -1505 se
rect 2269 -1511 2278 -1505
rect 1982 -1596 2010 -1586
tri 2010 -1596 2034 -1572 sw
rect 1982 -1628 2024 -1596
tri 2041 -1604 2042 -1603 sw
rect 2041 -1628 2042 -1604
tri 2044 -1605 2081 -1568 ne
rect 2081 -1596 2086 -1568
tri 2086 -1596 2112 -1570 sw
rect 2196 -1586 2205 -1552
rect 2196 -1596 2224 -1586
rect 2081 -1605 2165 -1596
tri 2081 -1624 2100 -1605 ne
rect 2100 -1624 2165 -1605
rect 1982 -1650 2042 -1628
rect 2164 -1628 2165 -1624
rect 2182 -1628 2224 -1596
rect 2164 -1650 2224 -1628
rect 2070 -1666 2087 -1652
rect 2119 -1666 2136 -1652
tri 1907 -1702 1929 -1680 se
rect 1929 -1687 1944 -1666
tri 1929 -1702 1944 -1687 nw
rect 2263 -1687 2278 -1511
tri 2278 -1518 2291 -1505 nw
rect 2364 -1586 2379 -1358
tri 1901 -1708 1907 -1702 se
rect 1907 -1708 1916 -1702
rect 1901 -1724 1916 -1708
tri 1916 -1715 1929 -1702 nw
rect 2070 -1710 2087 -1696
rect 2119 -1710 2136 -1696
tri 2263 -1702 2278 -1687 ne
tri 2278 -1702 2300 -1680 sw
rect 1901 -1760 1916 -1752
rect 1982 -1724 2042 -1710
rect 1997 -1734 2042 -1724
rect 1997 -1752 2025 -1734
tri 1901 -1775 1916 -1760 ne
tri 1916 -1775 1938 -1753 sw
rect 1982 -1762 2025 -1752
rect 2040 -1738 2042 -1734
rect 2164 -1724 2224 -1710
tri 2278 -1715 2291 -1702 ne
rect 2291 -1708 2300 -1702
tri 2300 -1708 2306 -1702 sw
rect 2164 -1734 2209 -1724
rect 2040 -1762 2114 -1738
rect 1982 -1766 2114 -1762
tri 2114 -1766 2142 -1738 sw
rect 2164 -1748 2166 -1734
tri 2164 -1750 2166 -1748 ne
rect 2178 -1752 2209 -1734
rect 2178 -1762 2224 -1752
rect 2291 -1723 2306 -1708
tri 1916 -1787 1928 -1775 ne
rect 1928 -1780 1938 -1775
tri 1938 -1780 1943 -1775 sw
rect 1827 -2126 1842 -1898
rect 1928 -1888 1943 -1780
rect 1982 -1822 2010 -1766
tri 2102 -1784 2120 -1766 ne
rect 2120 -1786 2142 -1766
tri 2142 -1786 2162 -1766 sw
tri 2178 -1780 2196 -1762 ne
rect 2001 -1856 2010 -1822
rect 2044 -1795 2086 -1794
rect 2044 -1829 2049 -1795
rect 2079 -1829 2086 -1795
rect 2044 -1838 2086 -1829
rect 2120 -1795 2162 -1786
rect 2120 -1829 2127 -1795
rect 2157 -1829 2162 -1795
rect 2120 -1834 2162 -1829
rect 2196 -1822 2224 -1762
tri 2269 -1775 2291 -1753 se
rect 2291 -1760 2306 -1752
tri 2291 -1775 2306 -1760 nw
tri 2263 -1781 2269 -1775 se
rect 2269 -1781 2278 -1775
rect 1982 -1866 2010 -1856
tri 2010 -1866 2034 -1842 sw
rect 1928 -1936 1944 -1888
rect 1982 -1898 2024 -1866
tri 2041 -1874 2042 -1873 sw
rect 2041 -1898 2042 -1874
tri 2044 -1875 2081 -1838 ne
rect 2081 -1866 2086 -1838
tri 2086 -1866 2112 -1840 sw
rect 2196 -1856 2205 -1822
rect 2196 -1866 2224 -1856
rect 2081 -1875 2165 -1866
tri 2081 -1894 2100 -1875 ne
rect 2100 -1894 2165 -1875
rect 1982 -1920 2042 -1898
rect 2164 -1898 2165 -1894
rect 2182 -1898 2224 -1866
rect 2164 -1920 2224 -1898
rect 2070 -1936 2087 -1922
rect 2119 -1936 2136 -1922
tri 1907 -1972 1929 -1950 se
rect 1929 -1957 1944 -1936
tri 1929 -1972 1944 -1957 nw
rect 2263 -1957 2278 -1781
tri 2278 -1788 2291 -1775 nw
rect 2364 -1856 2379 -1628
tri 1901 -1978 1907 -1972 se
rect 1907 -1978 1916 -1972
rect 1901 -1994 1916 -1978
tri 1916 -1985 1929 -1972 nw
rect 2070 -1980 2087 -1966
rect 2119 -1980 2136 -1966
tri 2263 -1972 2278 -1957 ne
tri 2278 -1972 2300 -1950 sw
rect 1901 -2030 1916 -2022
rect 1982 -1994 2042 -1980
rect 1997 -2004 2042 -1994
rect 1997 -2022 2025 -2004
tri 1901 -2045 1916 -2030 ne
tri 1916 -2045 1938 -2023 sw
rect 1982 -2032 2025 -2022
rect 2040 -2008 2042 -2004
rect 2164 -1994 2224 -1980
tri 2278 -1985 2291 -1972 ne
rect 2291 -1978 2300 -1972
tri 2300 -1978 2306 -1972 sw
rect 2164 -2004 2209 -1994
rect 2040 -2032 2114 -2008
rect 1982 -2036 2114 -2032
tri 2114 -2036 2142 -2008 sw
rect 2164 -2018 2166 -2004
tri 2164 -2020 2166 -2018 ne
rect 2178 -2022 2209 -2004
rect 2178 -2032 2224 -2022
rect 2291 -1993 2306 -1978
tri 1916 -2057 1928 -2045 ne
rect 1928 -2050 1938 -2045
tri 1938 -2050 1943 -2045 sw
rect 1827 -2396 1842 -2168
rect 1928 -2206 1943 -2050
rect 1982 -2092 2010 -2036
tri 2102 -2054 2120 -2036 ne
rect 2120 -2056 2142 -2036
tri 2142 -2056 2162 -2036 sw
tri 2178 -2050 2196 -2032 ne
rect 2001 -2126 2010 -2092
rect 2044 -2065 2086 -2064
rect 2044 -2099 2049 -2065
rect 2079 -2099 2086 -2065
rect 2044 -2108 2086 -2099
rect 2120 -2065 2162 -2056
rect 2120 -2099 2127 -2065
rect 2157 -2099 2162 -2065
rect 2120 -2104 2162 -2099
rect 2196 -2092 2224 -2032
tri 2269 -2045 2291 -2023 se
rect 2291 -2030 2306 -2022
tri 2291 -2045 2306 -2030 nw
tri 2263 -2051 2269 -2045 se
rect 2269 -2051 2278 -2045
rect 1982 -2136 2010 -2126
tri 2010 -2136 2034 -2112 sw
rect 1982 -2168 2024 -2136
tri 2041 -2144 2042 -2143 sw
rect 2041 -2168 2042 -2144
tri 2044 -2145 2081 -2108 ne
rect 2081 -2136 2086 -2108
tri 2086 -2136 2112 -2110 sw
rect 2196 -2126 2205 -2092
rect 2196 -2136 2224 -2126
rect 2081 -2145 2165 -2136
tri 2081 -2164 2100 -2145 ne
rect 2100 -2164 2165 -2145
rect 1982 -2190 2042 -2168
rect 2164 -2168 2165 -2164
rect 2182 -2168 2224 -2136
rect 2164 -2190 2224 -2168
rect 2070 -2206 2087 -2192
rect 2119 -2206 2136 -2192
tri 1907 -2242 1929 -2220 se
rect 1929 -2227 1944 -2206
tri 1929 -2242 1944 -2227 nw
rect 2263 -2227 2278 -2051
tri 2278 -2058 2291 -2045 nw
rect 2364 -2126 2379 -1898
tri 1901 -2248 1907 -2242 se
rect 1907 -2248 1916 -2242
rect 1901 -2264 1916 -2248
tri 1916 -2255 1929 -2242 nw
rect 2070 -2250 2087 -2236
rect 2119 -2250 2136 -2236
tri 2263 -2242 2278 -2227 ne
tri 2278 -2242 2300 -2220 sw
rect 1901 -2300 1916 -2292
rect 1982 -2264 2042 -2250
rect 1997 -2274 2042 -2264
rect 1997 -2292 2025 -2274
tri 1901 -2315 1916 -2300 ne
tri 1916 -2315 1938 -2293 sw
rect 1982 -2302 2025 -2292
rect 2040 -2278 2042 -2274
rect 2164 -2264 2224 -2250
tri 2278 -2255 2291 -2242 ne
rect 2291 -2248 2300 -2242
tri 2300 -2248 2306 -2242 sw
rect 2164 -2274 2209 -2264
rect 2040 -2302 2114 -2278
rect 1982 -2306 2114 -2302
tri 2114 -2306 2142 -2278 sw
rect 2164 -2288 2166 -2274
tri 2164 -2290 2166 -2288 ne
rect 2178 -2292 2209 -2274
rect 2178 -2302 2224 -2292
rect 2291 -2263 2306 -2248
tri 1916 -2327 1928 -2315 ne
rect 1928 -2320 1938 -2315
tri 1938 -2320 1943 -2315 sw
rect 1827 -2524 1842 -2438
rect 1928 -2476 1943 -2320
rect 1982 -2362 2010 -2306
tri 2102 -2324 2120 -2306 ne
rect 2120 -2326 2142 -2306
tri 2142 -2326 2162 -2306 sw
tri 2178 -2320 2196 -2302 ne
rect 2001 -2396 2010 -2362
rect 2044 -2335 2086 -2334
rect 2044 -2369 2049 -2335
rect 2079 -2369 2086 -2335
rect 2044 -2378 2086 -2369
rect 2120 -2335 2162 -2326
rect 2120 -2369 2127 -2335
rect 2157 -2369 2162 -2335
rect 2120 -2374 2162 -2369
rect 2196 -2362 2224 -2302
tri 2269 -2315 2291 -2293 se
rect 2291 -2300 2306 -2292
tri 2291 -2315 2306 -2300 nw
tri 2263 -2321 2269 -2315 se
rect 2269 -2321 2278 -2315
rect 1982 -2406 2010 -2396
tri 2010 -2406 2034 -2382 sw
rect 1982 -2438 2024 -2406
tri 2041 -2414 2042 -2413 sw
rect 2041 -2438 2042 -2414
tri 2044 -2415 2081 -2378 ne
rect 2081 -2406 2086 -2378
tri 2086 -2406 2112 -2380 sw
rect 2196 -2396 2205 -2362
rect 2196 -2406 2224 -2396
rect 2081 -2415 2165 -2406
tri 2081 -2434 2100 -2415 ne
rect 2100 -2434 2165 -2415
rect 1982 -2460 2042 -2438
rect 2164 -2438 2165 -2434
rect 2182 -2438 2224 -2406
rect 2164 -2460 2224 -2438
rect 2070 -2476 2087 -2462
rect 2119 -2476 2136 -2462
rect 2263 -2476 2278 -2321
tri 2278 -2328 2291 -2315 nw
rect 2364 -2396 2379 -2168
rect 2364 -2524 2379 -2438
rect 2407 1654 2422 1844
tri 2487 1808 2509 1830 se
rect 2509 1823 2524 1892
tri 2509 1808 2524 1823 nw
rect 2843 1823 2858 1892
tri 2481 1802 2487 1808 se
rect 2487 1802 2496 1808
rect 2481 1786 2496 1802
tri 2496 1795 2509 1808 nw
rect 2650 1800 2667 1814
rect 2699 1800 2716 1814
tri 2843 1808 2858 1823 ne
tri 2858 1808 2880 1830 sw
rect 2481 1750 2496 1758
rect 2562 1786 2622 1800
rect 2577 1776 2622 1786
rect 2577 1758 2605 1776
tri 2481 1735 2496 1750 ne
tri 2496 1735 2518 1757 sw
rect 2562 1748 2605 1758
rect 2620 1772 2622 1776
rect 2744 1786 2804 1800
tri 2858 1795 2871 1808 ne
rect 2871 1802 2880 1808
tri 2880 1802 2886 1808 sw
rect 2744 1776 2789 1786
rect 2620 1748 2694 1772
rect 2562 1744 2694 1748
tri 2694 1744 2722 1772 sw
rect 2744 1762 2746 1776
tri 2744 1760 2746 1762 ne
rect 2758 1758 2789 1776
rect 2758 1748 2804 1758
rect 2871 1787 2886 1802
tri 2496 1723 2508 1735 ne
rect 2508 1730 2518 1735
tri 2518 1730 2523 1735 sw
rect 2407 1384 2422 1612
rect 2508 1574 2523 1730
rect 2562 1688 2590 1744
tri 2682 1726 2700 1744 ne
rect 2700 1724 2722 1744
tri 2722 1724 2742 1744 sw
tri 2758 1730 2776 1748 ne
rect 2581 1654 2590 1688
rect 2624 1715 2666 1716
rect 2624 1681 2629 1715
rect 2659 1681 2666 1715
rect 2624 1672 2666 1681
rect 2700 1715 2742 1724
rect 2700 1681 2707 1715
rect 2737 1681 2742 1715
rect 2700 1676 2742 1681
rect 2776 1688 2804 1748
tri 2849 1735 2871 1757 se
rect 2871 1750 2886 1758
tri 2871 1735 2886 1750 nw
tri 2843 1729 2849 1735 se
rect 2849 1729 2858 1735
rect 2562 1644 2590 1654
tri 2590 1644 2614 1668 sw
rect 2562 1612 2604 1644
tri 2621 1636 2622 1637 sw
rect 2621 1612 2622 1636
tri 2624 1635 2661 1672 ne
rect 2661 1644 2666 1672
tri 2666 1644 2692 1670 sw
rect 2776 1654 2785 1688
rect 2776 1644 2804 1654
rect 2661 1635 2745 1644
tri 2661 1616 2680 1635 ne
rect 2680 1616 2745 1635
rect 2562 1590 2622 1612
rect 2744 1612 2745 1616
rect 2762 1612 2804 1644
rect 2744 1590 2804 1612
rect 2650 1574 2667 1588
rect 2699 1574 2716 1588
tri 2487 1538 2509 1560 se
rect 2509 1553 2524 1574
tri 2509 1538 2524 1553 nw
rect 2843 1553 2858 1729
tri 2858 1722 2871 1735 nw
rect 2944 1654 2959 1844
tri 2481 1532 2487 1538 se
rect 2487 1532 2496 1538
rect 2481 1516 2496 1532
tri 2496 1525 2509 1538 nw
rect 2650 1530 2667 1544
rect 2699 1530 2716 1544
tri 2843 1538 2858 1553 ne
tri 2858 1538 2880 1560 sw
rect 2481 1480 2496 1488
rect 2562 1516 2622 1530
rect 2577 1506 2622 1516
rect 2577 1488 2605 1506
tri 2481 1465 2496 1480 ne
tri 2496 1465 2518 1487 sw
rect 2562 1478 2605 1488
rect 2620 1502 2622 1506
rect 2744 1516 2804 1530
tri 2858 1525 2871 1538 ne
rect 2871 1532 2880 1538
tri 2880 1532 2886 1538 sw
rect 2744 1506 2789 1516
rect 2620 1478 2694 1502
rect 2562 1474 2694 1478
tri 2694 1474 2722 1502 sw
rect 2744 1492 2746 1506
tri 2744 1490 2746 1492 ne
rect 2758 1488 2789 1506
rect 2758 1478 2804 1488
rect 2871 1517 2886 1532
tri 2496 1453 2508 1465 ne
rect 2508 1460 2518 1465
tri 2518 1460 2523 1465 sw
rect 2407 1114 2422 1342
rect 2508 1352 2523 1460
rect 2562 1418 2590 1474
tri 2682 1456 2700 1474 ne
rect 2700 1454 2722 1474
tri 2722 1454 2742 1474 sw
tri 2758 1460 2776 1478 ne
rect 2581 1384 2590 1418
rect 2624 1445 2666 1446
rect 2624 1411 2629 1445
rect 2659 1411 2666 1445
rect 2624 1402 2666 1411
rect 2700 1445 2742 1454
rect 2700 1411 2707 1445
rect 2737 1411 2742 1445
rect 2700 1406 2742 1411
rect 2776 1418 2804 1478
tri 2849 1465 2871 1487 se
rect 2871 1480 2886 1488
tri 2871 1465 2886 1480 nw
tri 2843 1459 2849 1465 se
rect 2849 1459 2858 1465
rect 2562 1374 2590 1384
tri 2590 1374 2614 1398 sw
rect 2508 1304 2524 1352
rect 2562 1342 2604 1374
tri 2621 1366 2622 1367 sw
rect 2621 1342 2622 1366
tri 2624 1365 2661 1402 ne
rect 2661 1374 2666 1402
tri 2666 1374 2692 1400 sw
rect 2776 1384 2785 1418
rect 2776 1374 2804 1384
rect 2661 1365 2745 1374
tri 2661 1346 2680 1365 ne
rect 2680 1346 2745 1365
rect 2562 1320 2622 1342
rect 2744 1342 2745 1346
rect 2762 1342 2804 1374
rect 2744 1320 2804 1342
rect 2650 1304 2667 1318
rect 2699 1304 2716 1318
tri 2487 1268 2509 1290 se
rect 2509 1283 2524 1304
tri 2509 1268 2524 1283 nw
rect 2843 1283 2858 1459
tri 2858 1452 2871 1465 nw
rect 2944 1384 2959 1612
tri 2481 1262 2487 1268 se
rect 2487 1262 2496 1268
rect 2481 1246 2496 1262
tri 2496 1255 2509 1268 nw
rect 2650 1260 2667 1274
rect 2699 1260 2716 1274
tri 2843 1268 2858 1283 ne
tri 2858 1268 2880 1290 sw
rect 2481 1210 2496 1218
rect 2562 1246 2622 1260
rect 2577 1236 2622 1246
rect 2577 1218 2605 1236
tri 2481 1195 2496 1210 ne
tri 2496 1195 2518 1217 sw
rect 2562 1208 2605 1218
rect 2620 1232 2622 1236
rect 2744 1246 2804 1260
tri 2858 1255 2871 1268 ne
rect 2871 1262 2880 1268
tri 2880 1262 2886 1268 sw
rect 2744 1236 2789 1246
rect 2620 1208 2694 1232
rect 2562 1204 2694 1208
tri 2694 1204 2722 1232 sw
rect 2744 1222 2746 1236
tri 2744 1220 2746 1222 ne
rect 2758 1218 2789 1236
rect 2758 1208 2804 1218
rect 2871 1247 2886 1262
tri 2496 1183 2508 1195 ne
rect 2508 1190 2518 1195
tri 2518 1190 2523 1195 sw
rect 2407 844 2422 1072
rect 2508 1034 2523 1190
rect 2562 1148 2590 1204
tri 2682 1186 2700 1204 ne
rect 2700 1184 2722 1204
tri 2722 1184 2742 1204 sw
tri 2758 1190 2776 1208 ne
rect 2581 1114 2590 1148
rect 2624 1175 2666 1176
rect 2624 1141 2629 1175
rect 2659 1141 2666 1175
rect 2624 1132 2666 1141
rect 2700 1175 2742 1184
rect 2700 1141 2707 1175
rect 2737 1141 2742 1175
rect 2700 1136 2742 1141
rect 2776 1148 2804 1208
tri 2849 1195 2871 1217 se
rect 2871 1210 2886 1218
tri 2871 1195 2886 1210 nw
tri 2843 1189 2849 1195 se
rect 2849 1189 2858 1195
rect 2562 1104 2590 1114
tri 2590 1104 2614 1128 sw
rect 2562 1072 2604 1104
tri 2621 1096 2622 1097 sw
rect 2621 1072 2622 1096
tri 2624 1095 2661 1132 ne
rect 2661 1104 2666 1132
tri 2666 1104 2692 1130 sw
rect 2776 1114 2785 1148
rect 2776 1104 2804 1114
rect 2661 1095 2745 1104
tri 2661 1076 2680 1095 ne
rect 2680 1076 2745 1095
rect 2562 1050 2622 1072
rect 2744 1072 2745 1076
rect 2762 1072 2804 1104
rect 2744 1050 2804 1072
rect 2650 1034 2667 1048
rect 2699 1034 2716 1048
tri 2487 998 2509 1020 se
rect 2509 1013 2524 1034
tri 2509 998 2524 1013 nw
rect 2843 1013 2858 1189
tri 2858 1182 2871 1195 nw
rect 2944 1114 2959 1342
tri 2481 992 2487 998 se
rect 2487 992 2496 998
rect 2481 976 2496 992
tri 2496 985 2509 998 nw
rect 2650 990 2667 1004
rect 2699 990 2716 1004
tri 2843 998 2858 1013 ne
tri 2858 998 2880 1020 sw
rect 2481 940 2496 948
rect 2562 976 2622 990
rect 2577 966 2622 976
rect 2577 948 2605 966
tri 2481 925 2496 940 ne
tri 2496 925 2518 947 sw
rect 2562 938 2605 948
rect 2620 962 2622 966
rect 2744 976 2804 990
tri 2858 985 2871 998 ne
rect 2871 992 2880 998
tri 2880 992 2886 998 sw
rect 2744 966 2789 976
rect 2620 938 2694 962
rect 2562 934 2694 938
tri 2694 934 2722 962 sw
rect 2744 952 2746 966
tri 2744 950 2746 952 ne
rect 2758 948 2789 966
rect 2758 938 2804 948
rect 2871 977 2886 992
tri 2496 913 2508 925 ne
rect 2508 920 2518 925
tri 2518 920 2523 925 sw
rect 2407 574 2422 802
rect 2508 812 2523 920
rect 2562 878 2590 934
tri 2682 916 2700 934 ne
rect 2700 914 2722 934
tri 2722 914 2742 934 sw
tri 2758 920 2776 938 ne
rect 2581 844 2590 878
rect 2624 905 2666 906
rect 2624 871 2629 905
rect 2659 871 2666 905
rect 2624 862 2666 871
rect 2700 905 2742 914
rect 2700 871 2707 905
rect 2737 871 2742 905
rect 2700 866 2742 871
rect 2776 878 2804 938
tri 2849 925 2871 947 se
rect 2871 940 2886 948
tri 2871 925 2886 940 nw
tri 2843 919 2849 925 se
rect 2849 919 2858 925
rect 2562 834 2590 844
tri 2590 834 2614 858 sw
rect 2508 764 2524 812
rect 2562 802 2604 834
tri 2621 826 2622 827 sw
rect 2621 802 2622 826
tri 2624 825 2661 862 ne
rect 2661 834 2666 862
tri 2666 834 2692 860 sw
rect 2776 844 2785 878
rect 2776 834 2804 844
rect 2661 825 2745 834
tri 2661 806 2680 825 ne
rect 2680 806 2745 825
rect 2562 780 2622 802
rect 2744 802 2745 806
rect 2762 802 2804 834
rect 2744 780 2804 802
rect 2650 764 2667 778
rect 2699 764 2716 778
tri 2487 728 2509 750 se
rect 2509 743 2524 764
tri 2509 728 2524 743 nw
rect 2843 743 2858 919
tri 2858 912 2871 925 nw
rect 2944 844 2959 1072
tri 2481 722 2487 728 se
rect 2487 722 2496 728
rect 2481 706 2496 722
tri 2496 715 2509 728 nw
rect 2650 720 2667 734
rect 2699 720 2716 734
tri 2843 728 2858 743 ne
tri 2858 728 2880 750 sw
rect 2481 670 2496 678
rect 2562 706 2622 720
rect 2577 696 2622 706
rect 2577 678 2605 696
tri 2481 655 2496 670 ne
tri 2496 655 2518 677 sw
rect 2562 668 2605 678
rect 2620 692 2622 696
rect 2744 706 2804 720
tri 2858 715 2871 728 ne
rect 2871 722 2880 728
tri 2880 722 2886 728 sw
rect 2744 696 2789 706
rect 2620 668 2694 692
rect 2562 664 2694 668
tri 2694 664 2722 692 sw
rect 2744 682 2746 696
tri 2744 680 2746 682 ne
rect 2758 678 2789 696
rect 2758 668 2804 678
rect 2871 707 2886 722
tri 2496 643 2508 655 ne
rect 2508 650 2518 655
tri 2518 650 2523 655 sw
rect 2407 304 2422 532
rect 2508 494 2523 650
rect 2562 608 2590 664
tri 2682 646 2700 664 ne
rect 2700 644 2722 664
tri 2722 644 2742 664 sw
tri 2758 650 2776 668 ne
rect 2581 574 2590 608
rect 2624 635 2666 636
rect 2624 601 2629 635
rect 2659 601 2666 635
rect 2624 592 2666 601
rect 2700 635 2742 644
rect 2700 601 2707 635
rect 2737 601 2742 635
rect 2700 596 2742 601
rect 2776 608 2804 668
tri 2849 655 2871 677 se
rect 2871 670 2886 678
tri 2871 655 2886 670 nw
tri 2843 649 2849 655 se
rect 2849 649 2858 655
rect 2562 564 2590 574
tri 2590 564 2614 588 sw
rect 2562 532 2604 564
tri 2621 556 2622 557 sw
rect 2621 532 2622 556
tri 2624 555 2661 592 ne
rect 2661 564 2666 592
tri 2666 564 2692 590 sw
rect 2776 574 2785 608
rect 2776 564 2804 574
rect 2661 555 2745 564
tri 2661 536 2680 555 ne
rect 2680 536 2745 555
rect 2562 510 2622 532
rect 2744 532 2745 536
rect 2762 532 2804 564
rect 2744 510 2804 532
rect 2650 494 2667 508
rect 2699 494 2716 508
tri 2487 458 2509 480 se
rect 2509 473 2524 494
tri 2509 458 2524 473 nw
rect 2843 473 2858 649
tri 2858 642 2871 655 nw
rect 2944 574 2959 802
tri 2481 452 2487 458 se
rect 2487 452 2496 458
rect 2481 436 2496 452
tri 2496 445 2509 458 nw
rect 2650 450 2667 464
rect 2699 450 2716 464
tri 2843 458 2858 473 ne
tri 2858 458 2880 480 sw
rect 2481 400 2496 408
rect 2562 436 2622 450
rect 2577 426 2622 436
rect 2577 408 2605 426
tri 2481 385 2496 400 ne
tri 2496 385 2518 407 sw
rect 2562 398 2605 408
rect 2620 422 2622 426
rect 2744 436 2804 450
tri 2858 445 2871 458 ne
rect 2871 452 2880 458
tri 2880 452 2886 458 sw
rect 2744 426 2789 436
rect 2620 398 2694 422
rect 2562 394 2694 398
tri 2694 394 2722 422 sw
rect 2744 412 2746 426
tri 2744 410 2746 412 ne
rect 2758 408 2789 426
rect 2758 398 2804 408
rect 2871 437 2886 452
tri 2496 373 2508 385 ne
rect 2508 380 2518 385
tri 2518 380 2523 385 sw
rect 2407 34 2422 262
rect 2508 272 2523 380
rect 2562 338 2590 394
tri 2682 376 2700 394 ne
rect 2700 374 2722 394
tri 2722 374 2742 394 sw
tri 2758 380 2776 398 ne
rect 2581 304 2590 338
rect 2624 365 2666 366
rect 2624 331 2629 365
rect 2659 331 2666 365
rect 2624 322 2666 331
rect 2700 365 2742 374
rect 2700 331 2707 365
rect 2737 331 2742 365
rect 2700 326 2742 331
rect 2776 338 2804 398
tri 2849 385 2871 407 se
rect 2871 400 2886 408
tri 2871 385 2886 400 nw
tri 2843 379 2849 385 se
rect 2849 379 2858 385
rect 2562 294 2590 304
tri 2590 294 2614 318 sw
rect 2508 224 2524 272
rect 2562 262 2604 294
tri 2621 286 2622 287 sw
rect 2621 262 2622 286
tri 2624 285 2661 322 ne
rect 2661 294 2666 322
tri 2666 294 2692 320 sw
rect 2776 304 2785 338
rect 2776 294 2804 304
rect 2661 285 2745 294
tri 2661 266 2680 285 ne
rect 2680 266 2745 285
rect 2562 240 2622 262
rect 2744 262 2745 266
rect 2762 262 2804 294
rect 2744 240 2804 262
rect 2650 224 2667 238
rect 2699 224 2716 238
tri 2487 188 2509 210 se
rect 2509 203 2524 224
tri 2509 188 2524 203 nw
rect 2843 203 2858 379
tri 2858 372 2871 385 nw
rect 2944 304 2959 532
tri 2481 182 2487 188 se
rect 2487 182 2496 188
rect 2481 166 2496 182
tri 2496 175 2509 188 nw
rect 2650 180 2667 194
rect 2699 180 2716 194
tri 2843 188 2858 203 ne
tri 2858 188 2880 210 sw
rect 2481 130 2496 138
rect 2562 166 2622 180
rect 2577 156 2622 166
rect 2577 138 2605 156
tri 2481 115 2496 130 ne
tri 2496 115 2518 137 sw
rect 2562 128 2605 138
rect 2620 152 2622 156
rect 2744 166 2804 180
tri 2858 175 2871 188 ne
rect 2871 182 2880 188
tri 2880 182 2886 188 sw
rect 2744 156 2789 166
rect 2620 128 2694 152
rect 2562 124 2694 128
tri 2694 124 2722 152 sw
rect 2744 142 2746 156
tri 2744 140 2746 142 ne
rect 2758 138 2789 156
rect 2758 128 2804 138
rect 2871 167 2886 182
tri 2496 103 2508 115 ne
rect 2508 110 2518 115
tri 2518 110 2523 115 sw
rect 2407 -236 2422 -8
rect 2508 -46 2523 110
rect 2562 68 2590 124
tri 2682 106 2700 124 ne
rect 2700 104 2722 124
tri 2722 104 2742 124 sw
tri 2758 110 2776 128 ne
rect 2581 34 2590 68
rect 2624 95 2666 96
rect 2624 61 2629 95
rect 2659 61 2666 95
rect 2624 52 2666 61
rect 2700 95 2742 104
rect 2700 61 2707 95
rect 2737 61 2742 95
rect 2700 56 2742 61
rect 2776 68 2804 128
tri 2849 115 2871 137 se
rect 2871 130 2886 138
tri 2871 115 2886 130 nw
tri 2843 109 2849 115 se
rect 2849 109 2858 115
rect 2562 24 2590 34
tri 2590 24 2614 48 sw
rect 2562 -8 2604 24
tri 2621 16 2622 17 sw
rect 2621 -8 2622 16
tri 2624 15 2661 52 ne
rect 2661 24 2666 52
tri 2666 24 2692 50 sw
rect 2776 34 2785 68
rect 2776 24 2804 34
rect 2661 15 2745 24
tri 2661 -4 2680 15 ne
rect 2680 -4 2745 15
rect 2562 -30 2622 -8
rect 2744 -8 2745 -4
rect 2762 -8 2804 24
rect 2744 -30 2804 -8
rect 2650 -46 2667 -32
rect 2699 -46 2716 -32
tri 2487 -82 2509 -60 se
rect 2509 -67 2524 -46
tri 2509 -82 2524 -67 nw
rect 2843 -67 2858 109
tri 2858 102 2871 115 nw
rect 2944 34 2959 262
tri 2481 -88 2487 -82 se
rect 2487 -88 2496 -82
rect 2481 -104 2496 -88
tri 2496 -95 2509 -82 nw
rect 2650 -90 2667 -76
rect 2699 -90 2716 -76
tri 2843 -82 2858 -67 ne
tri 2858 -82 2880 -60 sw
rect 2481 -140 2496 -132
rect 2562 -104 2622 -90
rect 2577 -114 2622 -104
rect 2577 -132 2605 -114
tri 2481 -155 2496 -140 ne
tri 2496 -155 2518 -133 sw
rect 2562 -142 2605 -132
rect 2620 -118 2622 -114
rect 2744 -104 2804 -90
tri 2858 -95 2871 -82 ne
rect 2871 -88 2880 -82
tri 2880 -88 2886 -82 sw
rect 2744 -114 2789 -104
rect 2620 -142 2694 -118
rect 2562 -146 2694 -142
tri 2694 -146 2722 -118 sw
rect 2744 -128 2746 -114
tri 2744 -130 2746 -128 ne
rect 2758 -132 2789 -114
rect 2758 -142 2804 -132
rect 2871 -103 2886 -88
tri 2496 -167 2508 -155 ne
rect 2508 -160 2518 -155
tri 2518 -160 2523 -155 sw
rect 2407 -506 2422 -278
rect 2508 -268 2523 -160
rect 2562 -202 2590 -146
tri 2682 -164 2700 -146 ne
rect 2700 -166 2722 -146
tri 2722 -166 2742 -146 sw
tri 2758 -160 2776 -142 ne
rect 2581 -236 2590 -202
rect 2624 -175 2666 -174
rect 2624 -209 2629 -175
rect 2659 -209 2666 -175
rect 2624 -218 2666 -209
rect 2700 -175 2742 -166
rect 2700 -209 2707 -175
rect 2737 -209 2742 -175
rect 2700 -214 2742 -209
rect 2776 -202 2804 -142
tri 2849 -155 2871 -133 se
rect 2871 -140 2886 -132
tri 2871 -155 2886 -140 nw
tri 2843 -161 2849 -155 se
rect 2849 -161 2858 -155
rect 2562 -246 2590 -236
tri 2590 -246 2614 -222 sw
rect 2508 -316 2524 -268
rect 2562 -278 2604 -246
tri 2621 -254 2622 -253 sw
rect 2621 -278 2622 -254
tri 2624 -255 2661 -218 ne
rect 2661 -246 2666 -218
tri 2666 -246 2692 -220 sw
rect 2776 -236 2785 -202
rect 2776 -246 2804 -236
rect 2661 -255 2745 -246
tri 2661 -274 2680 -255 ne
rect 2680 -274 2745 -255
rect 2562 -300 2622 -278
rect 2744 -278 2745 -274
rect 2762 -278 2804 -246
rect 2744 -300 2804 -278
rect 2650 -316 2667 -302
rect 2699 -316 2716 -302
tri 2487 -352 2509 -330 se
rect 2509 -337 2524 -316
tri 2509 -352 2524 -337 nw
rect 2843 -337 2858 -161
tri 2858 -168 2871 -155 nw
rect 2944 -236 2959 -8
tri 2481 -358 2487 -352 se
rect 2487 -358 2496 -352
rect 2481 -374 2496 -358
tri 2496 -365 2509 -352 nw
rect 2650 -360 2667 -346
rect 2699 -360 2716 -346
tri 2843 -352 2858 -337 ne
tri 2858 -352 2880 -330 sw
rect 2481 -410 2496 -402
rect 2562 -374 2622 -360
rect 2577 -384 2622 -374
rect 2577 -402 2605 -384
tri 2481 -425 2496 -410 ne
tri 2496 -425 2518 -403 sw
rect 2562 -412 2605 -402
rect 2620 -388 2622 -384
rect 2744 -374 2804 -360
tri 2858 -365 2871 -352 ne
rect 2871 -358 2880 -352
tri 2880 -358 2886 -352 sw
rect 2744 -384 2789 -374
rect 2620 -412 2694 -388
rect 2562 -416 2694 -412
tri 2694 -416 2722 -388 sw
rect 2744 -398 2746 -384
tri 2744 -400 2746 -398 ne
rect 2758 -402 2789 -384
rect 2758 -412 2804 -402
rect 2871 -373 2886 -358
tri 2496 -437 2508 -425 ne
rect 2508 -430 2518 -425
tri 2518 -430 2523 -425 sw
rect 2407 -776 2422 -548
rect 2508 -586 2523 -430
rect 2562 -472 2590 -416
tri 2682 -434 2700 -416 ne
rect 2700 -436 2722 -416
tri 2722 -436 2742 -416 sw
tri 2758 -430 2776 -412 ne
rect 2581 -506 2590 -472
rect 2624 -445 2666 -444
rect 2624 -479 2629 -445
rect 2659 -479 2666 -445
rect 2624 -488 2666 -479
rect 2700 -445 2742 -436
rect 2700 -479 2707 -445
rect 2737 -479 2742 -445
rect 2700 -484 2742 -479
rect 2776 -472 2804 -412
tri 2849 -425 2871 -403 se
rect 2871 -410 2886 -402
tri 2871 -425 2886 -410 nw
tri 2843 -431 2849 -425 se
rect 2849 -431 2858 -425
rect 2562 -516 2590 -506
tri 2590 -516 2614 -492 sw
rect 2562 -548 2604 -516
tri 2621 -524 2622 -523 sw
rect 2621 -548 2622 -524
tri 2624 -525 2661 -488 ne
rect 2661 -516 2666 -488
tri 2666 -516 2692 -490 sw
rect 2776 -506 2785 -472
rect 2776 -516 2804 -506
rect 2661 -525 2745 -516
tri 2661 -544 2680 -525 ne
rect 2680 -544 2745 -525
rect 2562 -570 2622 -548
rect 2744 -548 2745 -544
rect 2762 -548 2804 -516
rect 2744 -570 2804 -548
rect 2650 -586 2667 -572
rect 2699 -586 2716 -572
tri 2487 -622 2509 -600 se
rect 2509 -607 2524 -586
tri 2509 -622 2524 -607 nw
rect 2843 -607 2858 -431
tri 2858 -438 2871 -425 nw
rect 2944 -506 2959 -278
tri 2481 -628 2487 -622 se
rect 2487 -628 2496 -622
rect 2481 -644 2496 -628
tri 2496 -635 2509 -622 nw
rect 2650 -630 2667 -616
rect 2699 -630 2716 -616
tri 2843 -622 2858 -607 ne
tri 2858 -622 2880 -600 sw
rect 2481 -680 2496 -672
rect 2562 -644 2622 -630
rect 2577 -654 2622 -644
rect 2577 -672 2605 -654
tri 2481 -695 2496 -680 ne
tri 2496 -695 2518 -673 sw
rect 2562 -682 2605 -672
rect 2620 -658 2622 -654
rect 2744 -644 2804 -630
tri 2858 -635 2871 -622 ne
rect 2871 -628 2880 -622
tri 2880 -628 2886 -622 sw
rect 2744 -654 2789 -644
rect 2620 -682 2694 -658
rect 2562 -686 2694 -682
tri 2694 -686 2722 -658 sw
rect 2744 -668 2746 -654
tri 2744 -670 2746 -668 ne
rect 2758 -672 2789 -654
rect 2758 -682 2804 -672
rect 2871 -643 2886 -628
tri 2496 -707 2508 -695 ne
rect 2508 -700 2518 -695
tri 2518 -700 2523 -695 sw
rect 2407 -1046 2422 -818
rect 2508 -808 2523 -700
rect 2562 -742 2590 -686
tri 2682 -704 2700 -686 ne
rect 2700 -706 2722 -686
tri 2722 -706 2742 -686 sw
tri 2758 -700 2776 -682 ne
rect 2581 -776 2590 -742
rect 2624 -715 2666 -714
rect 2624 -749 2629 -715
rect 2659 -749 2666 -715
rect 2624 -758 2666 -749
rect 2700 -715 2742 -706
rect 2700 -749 2707 -715
rect 2737 -749 2742 -715
rect 2700 -754 2742 -749
rect 2776 -742 2804 -682
tri 2849 -695 2871 -673 se
rect 2871 -680 2886 -672
tri 2871 -695 2886 -680 nw
tri 2843 -701 2849 -695 se
rect 2849 -701 2858 -695
rect 2562 -786 2590 -776
tri 2590 -786 2614 -762 sw
rect 2508 -856 2524 -808
rect 2562 -818 2604 -786
tri 2621 -794 2622 -793 sw
rect 2621 -818 2622 -794
tri 2624 -795 2661 -758 ne
rect 2661 -786 2666 -758
tri 2666 -786 2692 -760 sw
rect 2776 -776 2785 -742
rect 2776 -786 2804 -776
rect 2661 -795 2745 -786
tri 2661 -814 2680 -795 ne
rect 2680 -814 2745 -795
rect 2562 -840 2622 -818
rect 2744 -818 2745 -814
rect 2762 -818 2804 -786
rect 2744 -840 2804 -818
rect 2650 -856 2667 -842
rect 2699 -856 2716 -842
tri 2487 -892 2509 -870 se
rect 2509 -877 2524 -856
tri 2509 -892 2524 -877 nw
rect 2843 -877 2858 -701
tri 2858 -708 2871 -695 nw
rect 2944 -776 2959 -548
tri 2481 -898 2487 -892 se
rect 2487 -898 2496 -892
rect 2481 -914 2496 -898
tri 2496 -905 2509 -892 nw
rect 2650 -900 2667 -886
rect 2699 -900 2716 -886
tri 2843 -892 2858 -877 ne
tri 2858 -892 2880 -870 sw
rect 2481 -950 2496 -942
rect 2562 -914 2622 -900
rect 2577 -924 2622 -914
rect 2577 -942 2605 -924
tri 2481 -965 2496 -950 ne
tri 2496 -965 2518 -943 sw
rect 2562 -952 2605 -942
rect 2620 -928 2622 -924
rect 2744 -914 2804 -900
tri 2858 -905 2871 -892 ne
rect 2871 -898 2880 -892
tri 2880 -898 2886 -892 sw
rect 2744 -924 2789 -914
rect 2620 -952 2694 -928
rect 2562 -956 2694 -952
tri 2694 -956 2722 -928 sw
rect 2744 -938 2746 -924
tri 2744 -940 2746 -938 ne
rect 2758 -942 2789 -924
rect 2758 -952 2804 -942
rect 2871 -913 2886 -898
tri 2496 -977 2508 -965 ne
rect 2508 -970 2518 -965
tri 2518 -970 2523 -965 sw
rect 2407 -1316 2422 -1088
rect 2508 -1126 2523 -970
rect 2562 -1012 2590 -956
tri 2682 -974 2700 -956 ne
rect 2700 -976 2722 -956
tri 2722 -976 2742 -956 sw
tri 2758 -970 2776 -952 ne
rect 2581 -1046 2590 -1012
rect 2624 -985 2666 -984
rect 2624 -1019 2629 -985
rect 2659 -1019 2666 -985
rect 2624 -1028 2666 -1019
rect 2700 -985 2742 -976
rect 2700 -1019 2707 -985
rect 2737 -1019 2742 -985
rect 2700 -1024 2742 -1019
rect 2776 -1012 2804 -952
tri 2849 -965 2871 -943 se
rect 2871 -950 2886 -942
tri 2871 -965 2886 -950 nw
tri 2843 -971 2849 -965 se
rect 2849 -971 2858 -965
rect 2562 -1056 2590 -1046
tri 2590 -1056 2614 -1032 sw
rect 2562 -1088 2604 -1056
tri 2621 -1064 2622 -1063 sw
rect 2621 -1088 2622 -1064
tri 2624 -1065 2661 -1028 ne
rect 2661 -1056 2666 -1028
tri 2666 -1056 2692 -1030 sw
rect 2776 -1046 2785 -1012
rect 2776 -1056 2804 -1046
rect 2661 -1065 2745 -1056
tri 2661 -1084 2680 -1065 ne
rect 2680 -1084 2745 -1065
rect 2562 -1110 2622 -1088
rect 2744 -1088 2745 -1084
rect 2762 -1088 2804 -1056
rect 2744 -1110 2804 -1088
rect 2650 -1126 2667 -1112
rect 2699 -1126 2716 -1112
tri 2487 -1162 2509 -1140 se
rect 2509 -1147 2524 -1126
tri 2509 -1162 2524 -1147 nw
rect 2843 -1147 2858 -971
tri 2858 -978 2871 -965 nw
rect 2944 -1046 2959 -818
tri 2481 -1168 2487 -1162 se
rect 2487 -1168 2496 -1162
rect 2481 -1184 2496 -1168
tri 2496 -1175 2509 -1162 nw
rect 2650 -1170 2667 -1156
rect 2699 -1170 2716 -1156
tri 2843 -1162 2858 -1147 ne
tri 2858 -1162 2880 -1140 sw
rect 2481 -1220 2496 -1212
rect 2562 -1184 2622 -1170
rect 2577 -1194 2622 -1184
rect 2577 -1212 2605 -1194
tri 2481 -1235 2496 -1220 ne
tri 2496 -1235 2518 -1213 sw
rect 2562 -1222 2605 -1212
rect 2620 -1198 2622 -1194
rect 2744 -1184 2804 -1170
tri 2858 -1175 2871 -1162 ne
rect 2871 -1168 2880 -1162
tri 2880 -1168 2886 -1162 sw
rect 2744 -1194 2789 -1184
rect 2620 -1222 2694 -1198
rect 2562 -1226 2694 -1222
tri 2694 -1226 2722 -1198 sw
rect 2744 -1208 2746 -1194
tri 2744 -1210 2746 -1208 ne
rect 2758 -1212 2789 -1194
rect 2758 -1222 2804 -1212
rect 2871 -1183 2886 -1168
tri 2496 -1247 2508 -1235 ne
rect 2508 -1240 2518 -1235
tri 2518 -1240 2523 -1235 sw
rect 2407 -1586 2422 -1358
rect 2508 -1348 2523 -1240
rect 2562 -1282 2590 -1226
tri 2682 -1244 2700 -1226 ne
rect 2700 -1246 2722 -1226
tri 2722 -1246 2742 -1226 sw
tri 2758 -1240 2776 -1222 ne
rect 2581 -1316 2590 -1282
rect 2624 -1255 2666 -1254
rect 2624 -1289 2629 -1255
rect 2659 -1289 2666 -1255
rect 2624 -1298 2666 -1289
rect 2700 -1255 2742 -1246
rect 2700 -1289 2707 -1255
rect 2737 -1289 2742 -1255
rect 2700 -1294 2742 -1289
rect 2776 -1282 2804 -1222
tri 2849 -1235 2871 -1213 se
rect 2871 -1220 2886 -1212
tri 2871 -1235 2886 -1220 nw
tri 2843 -1241 2849 -1235 se
rect 2849 -1241 2858 -1235
rect 2562 -1326 2590 -1316
tri 2590 -1326 2614 -1302 sw
rect 2508 -1396 2524 -1348
rect 2562 -1358 2604 -1326
tri 2621 -1334 2622 -1333 sw
rect 2621 -1358 2622 -1334
tri 2624 -1335 2661 -1298 ne
rect 2661 -1326 2666 -1298
tri 2666 -1326 2692 -1300 sw
rect 2776 -1316 2785 -1282
rect 2776 -1326 2804 -1316
rect 2661 -1335 2745 -1326
tri 2661 -1354 2680 -1335 ne
rect 2680 -1354 2745 -1335
rect 2562 -1380 2622 -1358
rect 2744 -1358 2745 -1354
rect 2762 -1358 2804 -1326
rect 2744 -1380 2804 -1358
rect 2650 -1396 2667 -1382
rect 2699 -1396 2716 -1382
tri 2487 -1432 2509 -1410 se
rect 2509 -1417 2524 -1396
tri 2509 -1432 2524 -1417 nw
rect 2843 -1417 2858 -1241
tri 2858 -1248 2871 -1235 nw
rect 2944 -1316 2959 -1088
tri 2481 -1438 2487 -1432 se
rect 2487 -1438 2496 -1432
rect 2481 -1454 2496 -1438
tri 2496 -1445 2509 -1432 nw
rect 2650 -1440 2667 -1426
rect 2699 -1440 2716 -1426
tri 2843 -1432 2858 -1417 ne
tri 2858 -1432 2880 -1410 sw
rect 2481 -1490 2496 -1482
rect 2562 -1454 2622 -1440
rect 2577 -1464 2622 -1454
rect 2577 -1482 2605 -1464
tri 2481 -1505 2496 -1490 ne
tri 2496 -1505 2518 -1483 sw
rect 2562 -1492 2605 -1482
rect 2620 -1468 2622 -1464
rect 2744 -1454 2804 -1440
tri 2858 -1445 2871 -1432 ne
rect 2871 -1438 2880 -1432
tri 2880 -1438 2886 -1432 sw
rect 2744 -1464 2789 -1454
rect 2620 -1492 2694 -1468
rect 2562 -1496 2694 -1492
tri 2694 -1496 2722 -1468 sw
rect 2744 -1478 2746 -1464
tri 2744 -1480 2746 -1478 ne
rect 2758 -1482 2789 -1464
rect 2758 -1492 2804 -1482
rect 2871 -1453 2886 -1438
tri 2496 -1517 2508 -1505 ne
rect 2508 -1510 2518 -1505
tri 2518 -1510 2523 -1505 sw
rect 2407 -1856 2422 -1628
rect 2508 -1666 2523 -1510
rect 2562 -1552 2590 -1496
tri 2682 -1514 2700 -1496 ne
rect 2700 -1516 2722 -1496
tri 2722 -1516 2742 -1496 sw
tri 2758 -1510 2776 -1492 ne
rect 2581 -1586 2590 -1552
rect 2624 -1525 2666 -1524
rect 2624 -1559 2629 -1525
rect 2659 -1559 2666 -1525
rect 2624 -1568 2666 -1559
rect 2700 -1525 2742 -1516
rect 2700 -1559 2707 -1525
rect 2737 -1559 2742 -1525
rect 2700 -1564 2742 -1559
rect 2776 -1552 2804 -1492
tri 2849 -1505 2871 -1483 se
rect 2871 -1490 2886 -1482
tri 2871 -1505 2886 -1490 nw
tri 2843 -1511 2849 -1505 se
rect 2849 -1511 2858 -1505
rect 2562 -1596 2590 -1586
tri 2590 -1596 2614 -1572 sw
rect 2562 -1628 2604 -1596
tri 2621 -1604 2622 -1603 sw
rect 2621 -1628 2622 -1604
tri 2624 -1605 2661 -1568 ne
rect 2661 -1596 2666 -1568
tri 2666 -1596 2692 -1570 sw
rect 2776 -1586 2785 -1552
rect 2776 -1596 2804 -1586
rect 2661 -1605 2745 -1596
tri 2661 -1624 2680 -1605 ne
rect 2680 -1624 2745 -1605
rect 2562 -1650 2622 -1628
rect 2744 -1628 2745 -1624
rect 2762 -1628 2804 -1596
rect 2744 -1650 2804 -1628
rect 2650 -1666 2667 -1652
rect 2699 -1666 2716 -1652
tri 2487 -1702 2509 -1680 se
rect 2509 -1687 2524 -1666
tri 2509 -1702 2524 -1687 nw
rect 2843 -1687 2858 -1511
tri 2858 -1518 2871 -1505 nw
rect 2944 -1586 2959 -1358
tri 2481 -1708 2487 -1702 se
rect 2487 -1708 2496 -1702
rect 2481 -1724 2496 -1708
tri 2496 -1715 2509 -1702 nw
rect 2650 -1710 2667 -1696
rect 2699 -1710 2716 -1696
tri 2843 -1702 2858 -1687 ne
tri 2858 -1702 2880 -1680 sw
rect 2481 -1760 2496 -1752
rect 2562 -1724 2622 -1710
rect 2577 -1734 2622 -1724
rect 2577 -1752 2605 -1734
tri 2481 -1775 2496 -1760 ne
tri 2496 -1775 2518 -1753 sw
rect 2562 -1762 2605 -1752
rect 2620 -1738 2622 -1734
rect 2744 -1724 2804 -1710
tri 2858 -1715 2871 -1702 ne
rect 2871 -1708 2880 -1702
tri 2880 -1708 2886 -1702 sw
rect 2744 -1734 2789 -1724
rect 2620 -1762 2694 -1738
rect 2562 -1766 2694 -1762
tri 2694 -1766 2722 -1738 sw
rect 2744 -1748 2746 -1734
tri 2744 -1750 2746 -1748 ne
rect 2758 -1752 2789 -1734
rect 2758 -1762 2804 -1752
rect 2871 -1723 2886 -1708
tri 2496 -1787 2508 -1775 ne
rect 2508 -1780 2518 -1775
tri 2518 -1780 2523 -1775 sw
rect 2407 -2126 2422 -1898
rect 2508 -1888 2523 -1780
rect 2562 -1822 2590 -1766
tri 2682 -1784 2700 -1766 ne
rect 2700 -1786 2722 -1766
tri 2722 -1786 2742 -1766 sw
tri 2758 -1780 2776 -1762 ne
rect 2581 -1856 2590 -1822
rect 2624 -1795 2666 -1794
rect 2624 -1829 2629 -1795
rect 2659 -1829 2666 -1795
rect 2624 -1838 2666 -1829
rect 2700 -1795 2742 -1786
rect 2700 -1829 2707 -1795
rect 2737 -1829 2742 -1795
rect 2700 -1834 2742 -1829
rect 2776 -1822 2804 -1762
tri 2849 -1775 2871 -1753 se
rect 2871 -1760 2886 -1752
tri 2871 -1775 2886 -1760 nw
tri 2843 -1781 2849 -1775 se
rect 2849 -1781 2858 -1775
rect 2562 -1866 2590 -1856
tri 2590 -1866 2614 -1842 sw
rect 2508 -1936 2524 -1888
rect 2562 -1898 2604 -1866
tri 2621 -1874 2622 -1873 sw
rect 2621 -1898 2622 -1874
tri 2624 -1875 2661 -1838 ne
rect 2661 -1866 2666 -1838
tri 2666 -1866 2692 -1840 sw
rect 2776 -1856 2785 -1822
rect 2776 -1866 2804 -1856
rect 2661 -1875 2745 -1866
tri 2661 -1894 2680 -1875 ne
rect 2680 -1894 2745 -1875
rect 2562 -1920 2622 -1898
rect 2744 -1898 2745 -1894
rect 2762 -1898 2804 -1866
rect 2744 -1920 2804 -1898
rect 2650 -1936 2667 -1922
rect 2699 -1936 2716 -1922
tri 2487 -1972 2509 -1950 se
rect 2509 -1957 2524 -1936
tri 2509 -1972 2524 -1957 nw
rect 2843 -1957 2858 -1781
tri 2858 -1788 2871 -1775 nw
rect 2944 -1856 2959 -1628
tri 2481 -1978 2487 -1972 se
rect 2487 -1978 2496 -1972
rect 2481 -1994 2496 -1978
tri 2496 -1985 2509 -1972 nw
rect 2650 -1980 2667 -1966
rect 2699 -1980 2716 -1966
tri 2843 -1972 2858 -1957 ne
tri 2858 -1972 2880 -1950 sw
rect 2481 -2030 2496 -2022
rect 2562 -1994 2622 -1980
rect 2577 -2004 2622 -1994
rect 2577 -2022 2605 -2004
tri 2481 -2045 2496 -2030 ne
tri 2496 -2045 2518 -2023 sw
rect 2562 -2032 2605 -2022
rect 2620 -2008 2622 -2004
rect 2744 -1994 2804 -1980
tri 2858 -1985 2871 -1972 ne
rect 2871 -1978 2880 -1972
tri 2880 -1978 2886 -1972 sw
rect 2744 -2004 2789 -1994
rect 2620 -2032 2694 -2008
rect 2562 -2036 2694 -2032
tri 2694 -2036 2722 -2008 sw
rect 2744 -2018 2746 -2004
tri 2744 -2020 2746 -2018 ne
rect 2758 -2022 2789 -2004
rect 2758 -2032 2804 -2022
rect 2871 -1993 2886 -1978
tri 2496 -2057 2508 -2045 ne
rect 2508 -2050 2518 -2045
tri 2518 -2050 2523 -2045 sw
rect 2407 -2396 2422 -2168
rect 2508 -2206 2523 -2050
rect 2562 -2092 2590 -2036
tri 2682 -2054 2700 -2036 ne
rect 2700 -2056 2722 -2036
tri 2722 -2056 2742 -2036 sw
tri 2758 -2050 2776 -2032 ne
rect 2581 -2126 2590 -2092
rect 2624 -2065 2666 -2064
rect 2624 -2099 2629 -2065
rect 2659 -2099 2666 -2065
rect 2624 -2108 2666 -2099
rect 2700 -2065 2742 -2056
rect 2700 -2099 2707 -2065
rect 2737 -2099 2742 -2065
rect 2700 -2104 2742 -2099
rect 2776 -2092 2804 -2032
tri 2849 -2045 2871 -2023 se
rect 2871 -2030 2886 -2022
tri 2871 -2045 2886 -2030 nw
tri 2843 -2051 2849 -2045 se
rect 2849 -2051 2858 -2045
rect 2562 -2136 2590 -2126
tri 2590 -2136 2614 -2112 sw
rect 2562 -2168 2604 -2136
tri 2621 -2144 2622 -2143 sw
rect 2621 -2168 2622 -2144
tri 2624 -2145 2661 -2108 ne
rect 2661 -2136 2666 -2108
tri 2666 -2136 2692 -2110 sw
rect 2776 -2126 2785 -2092
rect 2776 -2136 2804 -2126
rect 2661 -2145 2745 -2136
tri 2661 -2164 2680 -2145 ne
rect 2680 -2164 2745 -2145
rect 2562 -2190 2622 -2168
rect 2744 -2168 2745 -2164
rect 2762 -2168 2804 -2136
rect 2744 -2190 2804 -2168
rect 2650 -2206 2667 -2192
rect 2699 -2206 2716 -2192
tri 2487 -2242 2509 -2220 se
rect 2509 -2227 2524 -2206
tri 2509 -2242 2524 -2227 nw
rect 2843 -2227 2858 -2051
tri 2858 -2058 2871 -2045 nw
rect 2944 -2126 2959 -1898
tri 2481 -2248 2487 -2242 se
rect 2487 -2248 2496 -2242
rect 2481 -2264 2496 -2248
tri 2496 -2255 2509 -2242 nw
rect 2650 -2250 2667 -2236
rect 2699 -2250 2716 -2236
tri 2843 -2242 2858 -2227 ne
tri 2858 -2242 2880 -2220 sw
rect 2481 -2300 2496 -2292
rect 2562 -2264 2622 -2250
rect 2577 -2274 2622 -2264
rect 2577 -2292 2605 -2274
tri 2481 -2315 2496 -2300 ne
tri 2496 -2315 2518 -2293 sw
rect 2562 -2302 2605 -2292
rect 2620 -2278 2622 -2274
rect 2744 -2264 2804 -2250
tri 2858 -2255 2871 -2242 ne
rect 2871 -2248 2880 -2242
tri 2880 -2248 2886 -2242 sw
rect 2744 -2274 2789 -2264
rect 2620 -2302 2694 -2278
rect 2562 -2306 2694 -2302
tri 2694 -2306 2722 -2278 sw
rect 2744 -2288 2746 -2274
tri 2744 -2290 2746 -2288 ne
rect 2758 -2292 2789 -2274
rect 2758 -2302 2804 -2292
rect 2871 -2263 2886 -2248
tri 2496 -2327 2508 -2315 ne
rect 2508 -2320 2518 -2315
tri 2518 -2320 2523 -2315 sw
rect 2407 -2524 2422 -2438
rect 2508 -2476 2523 -2320
rect 2562 -2362 2590 -2306
tri 2682 -2324 2700 -2306 ne
rect 2700 -2326 2722 -2306
tri 2722 -2326 2742 -2306 sw
tri 2758 -2320 2776 -2302 ne
rect 2581 -2396 2590 -2362
rect 2624 -2335 2666 -2334
rect 2624 -2369 2629 -2335
rect 2659 -2369 2666 -2335
rect 2624 -2378 2666 -2369
rect 2700 -2335 2742 -2326
rect 2700 -2369 2707 -2335
rect 2737 -2369 2742 -2335
rect 2700 -2374 2742 -2369
rect 2776 -2362 2804 -2302
tri 2849 -2315 2871 -2293 se
rect 2871 -2300 2886 -2292
tri 2871 -2315 2886 -2300 nw
tri 2843 -2321 2849 -2315 se
rect 2849 -2321 2858 -2315
rect 2562 -2406 2590 -2396
tri 2590 -2406 2614 -2382 sw
rect 2562 -2438 2604 -2406
tri 2621 -2414 2622 -2413 sw
rect 2621 -2438 2622 -2414
tri 2624 -2415 2661 -2378 ne
rect 2661 -2406 2666 -2378
tri 2666 -2406 2692 -2380 sw
rect 2776 -2396 2785 -2362
rect 2776 -2406 2804 -2396
rect 2661 -2415 2745 -2406
tri 2661 -2434 2680 -2415 ne
rect 2680 -2434 2745 -2415
rect 2562 -2460 2622 -2438
rect 2744 -2438 2745 -2434
rect 2762 -2438 2804 -2406
rect 2744 -2460 2804 -2438
rect 2650 -2476 2667 -2462
rect 2699 -2476 2716 -2462
rect 2843 -2476 2858 -2321
tri 2858 -2328 2871 -2315 nw
rect 2944 -2396 2959 -2168
rect 2944 -2524 2959 -2438
rect 2987 1654 3002 1844
tri 3067 1808 3089 1830 se
rect 3089 1823 3104 1892
tri 3089 1808 3104 1823 nw
rect 3423 1823 3438 1892
tri 3061 1802 3067 1808 se
rect 3067 1802 3076 1808
rect 3061 1786 3076 1802
tri 3076 1795 3089 1808 nw
rect 3230 1800 3247 1814
rect 3279 1800 3296 1814
tri 3423 1808 3438 1823 ne
tri 3438 1808 3460 1830 sw
rect 3061 1750 3076 1758
rect 3142 1786 3202 1800
rect 3157 1776 3202 1786
rect 3157 1758 3185 1776
tri 3061 1735 3076 1750 ne
tri 3076 1735 3098 1757 sw
rect 3142 1748 3185 1758
rect 3200 1772 3202 1776
rect 3324 1786 3384 1800
tri 3438 1795 3451 1808 ne
rect 3451 1802 3460 1808
tri 3460 1802 3466 1808 sw
rect 3324 1776 3369 1786
rect 3200 1748 3274 1772
rect 3142 1744 3274 1748
tri 3274 1744 3302 1772 sw
rect 3324 1762 3326 1776
tri 3324 1760 3326 1762 ne
rect 3338 1758 3369 1776
rect 3338 1748 3384 1758
rect 3451 1787 3466 1802
tri 3076 1723 3088 1735 ne
rect 3088 1730 3098 1735
tri 3098 1730 3103 1735 sw
rect 2987 1384 3002 1612
rect 3088 1574 3103 1730
rect 3142 1688 3170 1744
tri 3262 1726 3280 1744 ne
rect 3280 1724 3302 1744
tri 3302 1724 3322 1744 sw
tri 3338 1730 3356 1748 ne
rect 3161 1654 3170 1688
rect 3204 1715 3246 1716
rect 3204 1681 3209 1715
rect 3239 1681 3246 1715
rect 3204 1672 3246 1681
rect 3280 1715 3322 1724
rect 3280 1681 3287 1715
rect 3317 1681 3322 1715
rect 3280 1676 3322 1681
rect 3356 1688 3384 1748
tri 3429 1735 3451 1757 se
rect 3451 1750 3466 1758
tri 3451 1735 3466 1750 nw
tri 3423 1729 3429 1735 se
rect 3429 1729 3438 1735
rect 3142 1644 3170 1654
tri 3170 1644 3194 1668 sw
rect 3142 1612 3184 1644
tri 3201 1636 3202 1637 sw
rect 3201 1612 3202 1636
tri 3204 1635 3241 1672 ne
rect 3241 1644 3246 1672
tri 3246 1644 3272 1670 sw
rect 3356 1654 3365 1688
rect 3356 1644 3384 1654
rect 3241 1635 3325 1644
tri 3241 1616 3260 1635 ne
rect 3260 1616 3325 1635
rect 3142 1590 3202 1612
rect 3324 1612 3325 1616
rect 3342 1612 3384 1644
rect 3324 1590 3384 1612
rect 3230 1574 3247 1588
rect 3279 1574 3296 1588
tri 3067 1538 3089 1560 se
rect 3089 1553 3104 1574
tri 3089 1538 3104 1553 nw
rect 3423 1553 3438 1729
tri 3438 1722 3451 1735 nw
rect 3524 1654 3539 1844
tri 3061 1532 3067 1538 se
rect 3067 1532 3076 1538
rect 3061 1516 3076 1532
tri 3076 1525 3089 1538 nw
rect 3230 1530 3247 1544
rect 3279 1530 3296 1544
tri 3423 1538 3438 1553 ne
tri 3438 1538 3460 1560 sw
rect 3061 1480 3076 1488
rect 3142 1516 3202 1530
rect 3157 1506 3202 1516
rect 3157 1488 3185 1506
tri 3061 1465 3076 1480 ne
tri 3076 1465 3098 1487 sw
rect 3142 1478 3185 1488
rect 3200 1502 3202 1506
rect 3324 1516 3384 1530
tri 3438 1525 3451 1538 ne
rect 3451 1532 3460 1538
tri 3460 1532 3466 1538 sw
rect 3324 1506 3369 1516
rect 3200 1478 3274 1502
rect 3142 1474 3274 1478
tri 3274 1474 3302 1502 sw
rect 3324 1492 3326 1506
tri 3324 1490 3326 1492 ne
rect 3338 1488 3369 1506
rect 3338 1478 3384 1488
rect 3451 1517 3466 1532
tri 3076 1453 3088 1465 ne
rect 3088 1460 3098 1465
tri 3098 1460 3103 1465 sw
rect 2987 1114 3002 1342
rect 3088 1352 3103 1460
rect 3142 1418 3170 1474
tri 3262 1456 3280 1474 ne
rect 3280 1454 3302 1474
tri 3302 1454 3322 1474 sw
tri 3338 1460 3356 1478 ne
rect 3161 1384 3170 1418
rect 3204 1445 3246 1446
rect 3204 1411 3209 1445
rect 3239 1411 3246 1445
rect 3204 1402 3246 1411
rect 3280 1445 3322 1454
rect 3280 1411 3287 1445
rect 3317 1411 3322 1445
rect 3280 1406 3322 1411
rect 3356 1418 3384 1478
tri 3429 1465 3451 1487 se
rect 3451 1480 3466 1488
tri 3451 1465 3466 1480 nw
tri 3423 1459 3429 1465 se
rect 3429 1459 3438 1465
rect 3142 1374 3170 1384
tri 3170 1374 3194 1398 sw
rect 3088 1304 3104 1352
rect 3142 1342 3184 1374
tri 3201 1366 3202 1367 sw
rect 3201 1342 3202 1366
tri 3204 1365 3241 1402 ne
rect 3241 1374 3246 1402
tri 3246 1374 3272 1400 sw
rect 3356 1384 3365 1418
rect 3356 1374 3384 1384
rect 3241 1365 3325 1374
tri 3241 1346 3260 1365 ne
rect 3260 1346 3325 1365
rect 3142 1320 3202 1342
rect 3324 1342 3325 1346
rect 3342 1342 3384 1374
rect 3324 1320 3384 1342
rect 3230 1304 3247 1318
rect 3279 1304 3296 1318
tri 3067 1268 3089 1290 se
rect 3089 1283 3104 1304
tri 3089 1268 3104 1283 nw
rect 3423 1283 3438 1459
tri 3438 1452 3451 1465 nw
rect 3524 1384 3539 1612
tri 3061 1262 3067 1268 se
rect 3067 1262 3076 1268
rect 3061 1246 3076 1262
tri 3076 1255 3089 1268 nw
rect 3230 1260 3247 1274
rect 3279 1260 3296 1274
tri 3423 1268 3438 1283 ne
tri 3438 1268 3460 1290 sw
rect 3061 1210 3076 1218
rect 3142 1246 3202 1260
rect 3157 1236 3202 1246
rect 3157 1218 3185 1236
tri 3061 1195 3076 1210 ne
tri 3076 1195 3098 1217 sw
rect 3142 1208 3185 1218
rect 3200 1232 3202 1236
rect 3324 1246 3384 1260
tri 3438 1255 3451 1268 ne
rect 3451 1262 3460 1268
tri 3460 1262 3466 1268 sw
rect 3324 1236 3369 1246
rect 3200 1208 3274 1232
rect 3142 1204 3274 1208
tri 3274 1204 3302 1232 sw
rect 3324 1222 3326 1236
tri 3324 1220 3326 1222 ne
rect 3338 1218 3369 1236
rect 3338 1208 3384 1218
rect 3451 1247 3466 1262
tri 3076 1183 3088 1195 ne
rect 3088 1190 3098 1195
tri 3098 1190 3103 1195 sw
rect 2987 844 3002 1072
rect 3088 1034 3103 1190
rect 3142 1148 3170 1204
tri 3262 1186 3280 1204 ne
rect 3280 1184 3302 1204
tri 3302 1184 3322 1204 sw
tri 3338 1190 3356 1208 ne
rect 3161 1114 3170 1148
rect 3204 1175 3246 1176
rect 3204 1141 3209 1175
rect 3239 1141 3246 1175
rect 3204 1132 3246 1141
rect 3280 1175 3322 1184
rect 3280 1141 3287 1175
rect 3317 1141 3322 1175
rect 3280 1136 3322 1141
rect 3356 1148 3384 1208
tri 3429 1195 3451 1217 se
rect 3451 1210 3466 1218
tri 3451 1195 3466 1210 nw
tri 3423 1189 3429 1195 se
rect 3429 1189 3438 1195
rect 3142 1104 3170 1114
tri 3170 1104 3194 1128 sw
rect 3142 1072 3184 1104
tri 3201 1096 3202 1097 sw
rect 3201 1072 3202 1096
tri 3204 1095 3241 1132 ne
rect 3241 1104 3246 1132
tri 3246 1104 3272 1130 sw
rect 3356 1114 3365 1148
rect 3356 1104 3384 1114
rect 3241 1095 3325 1104
tri 3241 1076 3260 1095 ne
rect 3260 1076 3325 1095
rect 3142 1050 3202 1072
rect 3324 1072 3325 1076
rect 3342 1072 3384 1104
rect 3324 1050 3384 1072
rect 3230 1034 3247 1048
rect 3279 1034 3296 1048
tri 3067 998 3089 1020 se
rect 3089 1013 3104 1034
tri 3089 998 3104 1013 nw
rect 3423 1013 3438 1189
tri 3438 1182 3451 1195 nw
rect 3524 1114 3539 1342
tri 3061 992 3067 998 se
rect 3067 992 3076 998
rect 3061 976 3076 992
tri 3076 985 3089 998 nw
rect 3230 990 3247 1004
rect 3279 990 3296 1004
tri 3423 998 3438 1013 ne
tri 3438 998 3460 1020 sw
rect 3061 940 3076 948
rect 3142 976 3202 990
rect 3157 966 3202 976
rect 3157 948 3185 966
tri 3061 925 3076 940 ne
tri 3076 925 3098 947 sw
rect 3142 938 3185 948
rect 3200 962 3202 966
rect 3324 976 3384 990
tri 3438 985 3451 998 ne
rect 3451 992 3460 998
tri 3460 992 3466 998 sw
rect 3324 966 3369 976
rect 3200 938 3274 962
rect 3142 934 3274 938
tri 3274 934 3302 962 sw
rect 3324 952 3326 966
tri 3324 950 3326 952 ne
rect 3338 948 3369 966
rect 3338 938 3384 948
rect 3451 977 3466 992
tri 3076 913 3088 925 ne
rect 3088 920 3098 925
tri 3098 920 3103 925 sw
rect 2987 574 3002 802
rect 3088 812 3103 920
rect 3142 878 3170 934
tri 3262 916 3280 934 ne
rect 3280 914 3302 934
tri 3302 914 3322 934 sw
tri 3338 920 3356 938 ne
rect 3161 844 3170 878
rect 3204 905 3246 906
rect 3204 871 3209 905
rect 3239 871 3246 905
rect 3204 862 3246 871
rect 3280 905 3322 914
rect 3280 871 3287 905
rect 3317 871 3322 905
rect 3280 866 3322 871
rect 3356 878 3384 938
tri 3429 925 3451 947 se
rect 3451 940 3466 948
tri 3451 925 3466 940 nw
tri 3423 919 3429 925 se
rect 3429 919 3438 925
rect 3142 834 3170 844
tri 3170 834 3194 858 sw
rect 3088 764 3104 812
rect 3142 802 3184 834
tri 3201 826 3202 827 sw
rect 3201 802 3202 826
tri 3204 825 3241 862 ne
rect 3241 834 3246 862
tri 3246 834 3272 860 sw
rect 3356 844 3365 878
rect 3356 834 3384 844
rect 3241 825 3325 834
tri 3241 806 3260 825 ne
rect 3260 806 3325 825
rect 3142 780 3202 802
rect 3324 802 3325 806
rect 3342 802 3384 834
rect 3324 780 3384 802
rect 3230 764 3247 778
rect 3279 764 3296 778
tri 3067 728 3089 750 se
rect 3089 743 3104 764
tri 3089 728 3104 743 nw
rect 3423 743 3438 919
tri 3438 912 3451 925 nw
rect 3524 844 3539 1072
tri 3061 722 3067 728 se
rect 3067 722 3076 728
rect 3061 706 3076 722
tri 3076 715 3089 728 nw
rect 3230 720 3247 734
rect 3279 720 3296 734
tri 3423 728 3438 743 ne
tri 3438 728 3460 750 sw
rect 3061 670 3076 678
rect 3142 706 3202 720
rect 3157 696 3202 706
rect 3157 678 3185 696
tri 3061 655 3076 670 ne
tri 3076 655 3098 677 sw
rect 3142 668 3185 678
rect 3200 692 3202 696
rect 3324 706 3384 720
tri 3438 715 3451 728 ne
rect 3451 722 3460 728
tri 3460 722 3466 728 sw
rect 3324 696 3369 706
rect 3200 668 3274 692
rect 3142 664 3274 668
tri 3274 664 3302 692 sw
rect 3324 682 3326 696
tri 3324 680 3326 682 ne
rect 3338 678 3369 696
rect 3338 668 3384 678
rect 3451 707 3466 722
tri 3076 643 3088 655 ne
rect 3088 650 3098 655
tri 3098 650 3103 655 sw
rect 2987 304 3002 532
rect 3088 494 3103 650
rect 3142 608 3170 664
tri 3262 646 3280 664 ne
rect 3280 644 3302 664
tri 3302 644 3322 664 sw
tri 3338 650 3356 668 ne
rect 3161 574 3170 608
rect 3204 635 3246 636
rect 3204 601 3209 635
rect 3239 601 3246 635
rect 3204 592 3246 601
rect 3280 635 3322 644
rect 3280 601 3287 635
rect 3317 601 3322 635
rect 3280 596 3322 601
rect 3356 608 3384 668
tri 3429 655 3451 677 se
rect 3451 670 3466 678
tri 3451 655 3466 670 nw
tri 3423 649 3429 655 se
rect 3429 649 3438 655
rect 3142 564 3170 574
tri 3170 564 3194 588 sw
rect 3142 532 3184 564
tri 3201 556 3202 557 sw
rect 3201 532 3202 556
tri 3204 555 3241 592 ne
rect 3241 564 3246 592
tri 3246 564 3272 590 sw
rect 3356 574 3365 608
rect 3356 564 3384 574
rect 3241 555 3325 564
tri 3241 536 3260 555 ne
rect 3260 536 3325 555
rect 3142 510 3202 532
rect 3324 532 3325 536
rect 3342 532 3384 564
rect 3324 510 3384 532
rect 3230 494 3247 508
rect 3279 494 3296 508
tri 3067 458 3089 480 se
rect 3089 473 3104 494
tri 3089 458 3104 473 nw
rect 3423 473 3438 649
tri 3438 642 3451 655 nw
rect 3524 574 3539 802
tri 3061 452 3067 458 se
rect 3067 452 3076 458
rect 3061 436 3076 452
tri 3076 445 3089 458 nw
rect 3230 450 3247 464
rect 3279 450 3296 464
tri 3423 458 3438 473 ne
tri 3438 458 3460 480 sw
rect 3061 400 3076 408
rect 3142 436 3202 450
rect 3157 426 3202 436
rect 3157 408 3185 426
tri 3061 385 3076 400 ne
tri 3076 385 3098 407 sw
rect 3142 398 3185 408
rect 3200 422 3202 426
rect 3324 436 3384 450
tri 3438 445 3451 458 ne
rect 3451 452 3460 458
tri 3460 452 3466 458 sw
rect 3324 426 3369 436
rect 3200 398 3274 422
rect 3142 394 3274 398
tri 3274 394 3302 422 sw
rect 3324 412 3326 426
tri 3324 410 3326 412 ne
rect 3338 408 3369 426
rect 3338 398 3384 408
rect 3451 437 3466 452
tri 3076 373 3088 385 ne
rect 3088 380 3098 385
tri 3098 380 3103 385 sw
rect 2987 34 3002 262
rect 3088 272 3103 380
rect 3142 338 3170 394
tri 3262 376 3280 394 ne
rect 3280 374 3302 394
tri 3302 374 3322 394 sw
tri 3338 380 3356 398 ne
rect 3161 304 3170 338
rect 3204 365 3246 366
rect 3204 331 3209 365
rect 3239 331 3246 365
rect 3204 322 3246 331
rect 3280 365 3322 374
rect 3280 331 3287 365
rect 3317 331 3322 365
rect 3280 326 3322 331
rect 3356 338 3384 398
tri 3429 385 3451 407 se
rect 3451 400 3466 408
tri 3451 385 3466 400 nw
tri 3423 379 3429 385 se
rect 3429 379 3438 385
rect 3142 294 3170 304
tri 3170 294 3194 318 sw
rect 3088 224 3104 272
rect 3142 262 3184 294
tri 3201 286 3202 287 sw
rect 3201 262 3202 286
tri 3204 285 3241 322 ne
rect 3241 294 3246 322
tri 3246 294 3272 320 sw
rect 3356 304 3365 338
rect 3356 294 3384 304
rect 3241 285 3325 294
tri 3241 266 3260 285 ne
rect 3260 266 3325 285
rect 3142 240 3202 262
rect 3324 262 3325 266
rect 3342 262 3384 294
rect 3324 240 3384 262
rect 3230 224 3247 238
rect 3279 224 3296 238
tri 3067 188 3089 210 se
rect 3089 203 3104 224
tri 3089 188 3104 203 nw
rect 3423 203 3438 379
tri 3438 372 3451 385 nw
rect 3524 304 3539 532
tri 3061 182 3067 188 se
rect 3067 182 3076 188
rect 3061 166 3076 182
tri 3076 175 3089 188 nw
rect 3230 180 3247 194
rect 3279 180 3296 194
tri 3423 188 3438 203 ne
tri 3438 188 3460 210 sw
rect 3061 130 3076 138
rect 3142 166 3202 180
rect 3157 156 3202 166
rect 3157 138 3185 156
tri 3061 115 3076 130 ne
tri 3076 115 3098 137 sw
rect 3142 128 3185 138
rect 3200 152 3202 156
rect 3324 166 3384 180
tri 3438 175 3451 188 ne
rect 3451 182 3460 188
tri 3460 182 3466 188 sw
rect 3324 156 3369 166
rect 3200 128 3274 152
rect 3142 124 3274 128
tri 3274 124 3302 152 sw
rect 3324 142 3326 156
tri 3324 140 3326 142 ne
rect 3338 138 3369 156
rect 3338 128 3384 138
rect 3451 167 3466 182
tri 3076 103 3088 115 ne
rect 3088 110 3098 115
tri 3098 110 3103 115 sw
rect 2987 -236 3002 -8
rect 3088 -46 3103 110
rect 3142 68 3170 124
tri 3262 106 3280 124 ne
rect 3280 104 3302 124
tri 3302 104 3322 124 sw
tri 3338 110 3356 128 ne
rect 3161 34 3170 68
rect 3204 95 3246 96
rect 3204 61 3209 95
rect 3239 61 3246 95
rect 3204 52 3246 61
rect 3280 95 3322 104
rect 3280 61 3287 95
rect 3317 61 3322 95
rect 3280 56 3322 61
rect 3356 68 3384 128
tri 3429 115 3451 137 se
rect 3451 130 3466 138
tri 3451 115 3466 130 nw
tri 3423 109 3429 115 se
rect 3429 109 3438 115
rect 3142 24 3170 34
tri 3170 24 3194 48 sw
rect 3142 -8 3184 24
tri 3201 16 3202 17 sw
rect 3201 -8 3202 16
tri 3204 15 3241 52 ne
rect 3241 24 3246 52
tri 3246 24 3272 50 sw
rect 3356 34 3365 68
rect 3356 24 3384 34
rect 3241 15 3325 24
tri 3241 -4 3260 15 ne
rect 3260 -4 3325 15
rect 3142 -30 3202 -8
rect 3324 -8 3325 -4
rect 3342 -8 3384 24
rect 3324 -30 3384 -8
rect 3230 -46 3247 -32
rect 3279 -46 3296 -32
tri 3067 -82 3089 -60 se
rect 3089 -67 3104 -46
tri 3089 -82 3104 -67 nw
rect 3423 -67 3438 109
tri 3438 102 3451 115 nw
rect 3524 34 3539 262
tri 3061 -88 3067 -82 se
rect 3067 -88 3076 -82
rect 3061 -104 3076 -88
tri 3076 -95 3089 -82 nw
rect 3230 -90 3247 -76
rect 3279 -90 3296 -76
tri 3423 -82 3438 -67 ne
tri 3438 -82 3460 -60 sw
rect 3061 -140 3076 -132
rect 3142 -104 3202 -90
rect 3157 -114 3202 -104
rect 3157 -132 3185 -114
tri 3061 -155 3076 -140 ne
tri 3076 -155 3098 -133 sw
rect 3142 -142 3185 -132
rect 3200 -118 3202 -114
rect 3324 -104 3384 -90
tri 3438 -95 3451 -82 ne
rect 3451 -88 3460 -82
tri 3460 -88 3466 -82 sw
rect 3324 -114 3369 -104
rect 3200 -142 3274 -118
rect 3142 -146 3274 -142
tri 3274 -146 3302 -118 sw
rect 3324 -128 3326 -114
tri 3324 -130 3326 -128 ne
rect 3338 -132 3369 -114
rect 3338 -142 3384 -132
rect 3451 -103 3466 -88
tri 3076 -167 3088 -155 ne
rect 3088 -160 3098 -155
tri 3098 -160 3103 -155 sw
rect 2987 -506 3002 -278
rect 3088 -268 3103 -160
rect 3142 -202 3170 -146
tri 3262 -164 3280 -146 ne
rect 3280 -166 3302 -146
tri 3302 -166 3322 -146 sw
tri 3338 -160 3356 -142 ne
rect 3161 -236 3170 -202
rect 3204 -175 3246 -174
rect 3204 -209 3209 -175
rect 3239 -209 3246 -175
rect 3204 -218 3246 -209
rect 3280 -175 3322 -166
rect 3280 -209 3287 -175
rect 3317 -209 3322 -175
rect 3280 -214 3322 -209
rect 3356 -202 3384 -142
tri 3429 -155 3451 -133 se
rect 3451 -140 3466 -132
tri 3451 -155 3466 -140 nw
tri 3423 -161 3429 -155 se
rect 3429 -161 3438 -155
rect 3142 -246 3170 -236
tri 3170 -246 3194 -222 sw
rect 3088 -316 3104 -268
rect 3142 -278 3184 -246
tri 3201 -254 3202 -253 sw
rect 3201 -278 3202 -254
tri 3204 -255 3241 -218 ne
rect 3241 -246 3246 -218
tri 3246 -246 3272 -220 sw
rect 3356 -236 3365 -202
rect 3356 -246 3384 -236
rect 3241 -255 3325 -246
tri 3241 -274 3260 -255 ne
rect 3260 -274 3325 -255
rect 3142 -300 3202 -278
rect 3324 -278 3325 -274
rect 3342 -278 3384 -246
rect 3324 -300 3384 -278
rect 3230 -316 3247 -302
rect 3279 -316 3296 -302
tri 3067 -352 3089 -330 se
rect 3089 -337 3104 -316
tri 3089 -352 3104 -337 nw
rect 3423 -337 3438 -161
tri 3438 -168 3451 -155 nw
rect 3524 -236 3539 -8
tri 3061 -358 3067 -352 se
rect 3067 -358 3076 -352
rect 3061 -374 3076 -358
tri 3076 -365 3089 -352 nw
rect 3230 -360 3247 -346
rect 3279 -360 3296 -346
tri 3423 -352 3438 -337 ne
tri 3438 -352 3460 -330 sw
rect 3061 -410 3076 -402
rect 3142 -374 3202 -360
rect 3157 -384 3202 -374
rect 3157 -402 3185 -384
tri 3061 -425 3076 -410 ne
tri 3076 -425 3098 -403 sw
rect 3142 -412 3185 -402
rect 3200 -388 3202 -384
rect 3324 -374 3384 -360
tri 3438 -365 3451 -352 ne
rect 3451 -358 3460 -352
tri 3460 -358 3466 -352 sw
rect 3324 -384 3369 -374
rect 3200 -412 3274 -388
rect 3142 -416 3274 -412
tri 3274 -416 3302 -388 sw
rect 3324 -398 3326 -384
tri 3324 -400 3326 -398 ne
rect 3338 -402 3369 -384
rect 3338 -412 3384 -402
rect 3451 -373 3466 -358
tri 3076 -437 3088 -425 ne
rect 3088 -430 3098 -425
tri 3098 -430 3103 -425 sw
rect 2987 -776 3002 -548
rect 3088 -586 3103 -430
rect 3142 -472 3170 -416
tri 3262 -434 3280 -416 ne
rect 3280 -436 3302 -416
tri 3302 -436 3322 -416 sw
tri 3338 -430 3356 -412 ne
rect 3161 -506 3170 -472
rect 3204 -445 3246 -444
rect 3204 -479 3209 -445
rect 3239 -479 3246 -445
rect 3204 -488 3246 -479
rect 3280 -445 3322 -436
rect 3280 -479 3287 -445
rect 3317 -479 3322 -445
rect 3280 -484 3322 -479
rect 3356 -472 3384 -412
tri 3429 -425 3451 -403 se
rect 3451 -410 3466 -402
tri 3451 -425 3466 -410 nw
tri 3423 -431 3429 -425 se
rect 3429 -431 3438 -425
rect 3142 -516 3170 -506
tri 3170 -516 3194 -492 sw
rect 3142 -548 3184 -516
tri 3201 -524 3202 -523 sw
rect 3201 -548 3202 -524
tri 3204 -525 3241 -488 ne
rect 3241 -516 3246 -488
tri 3246 -516 3272 -490 sw
rect 3356 -506 3365 -472
rect 3356 -516 3384 -506
rect 3241 -525 3325 -516
tri 3241 -544 3260 -525 ne
rect 3260 -544 3325 -525
rect 3142 -570 3202 -548
rect 3324 -548 3325 -544
rect 3342 -548 3384 -516
rect 3324 -570 3384 -548
rect 3230 -586 3247 -572
rect 3279 -586 3296 -572
tri 3067 -622 3089 -600 se
rect 3089 -607 3104 -586
tri 3089 -622 3104 -607 nw
rect 3423 -607 3438 -431
tri 3438 -438 3451 -425 nw
rect 3524 -506 3539 -278
tri 3061 -628 3067 -622 se
rect 3067 -628 3076 -622
rect 3061 -644 3076 -628
tri 3076 -635 3089 -622 nw
rect 3230 -630 3247 -616
rect 3279 -630 3296 -616
tri 3423 -622 3438 -607 ne
tri 3438 -622 3460 -600 sw
rect 3061 -680 3076 -672
rect 3142 -644 3202 -630
rect 3157 -654 3202 -644
rect 3157 -672 3185 -654
tri 3061 -695 3076 -680 ne
tri 3076 -695 3098 -673 sw
rect 3142 -682 3185 -672
rect 3200 -658 3202 -654
rect 3324 -644 3384 -630
tri 3438 -635 3451 -622 ne
rect 3451 -628 3460 -622
tri 3460 -628 3466 -622 sw
rect 3324 -654 3369 -644
rect 3200 -682 3274 -658
rect 3142 -686 3274 -682
tri 3274 -686 3302 -658 sw
rect 3324 -668 3326 -654
tri 3324 -670 3326 -668 ne
rect 3338 -672 3369 -654
rect 3338 -682 3384 -672
rect 3451 -643 3466 -628
tri 3076 -707 3088 -695 ne
rect 3088 -700 3098 -695
tri 3098 -700 3103 -695 sw
rect 2987 -1046 3002 -818
rect 3088 -808 3103 -700
rect 3142 -742 3170 -686
tri 3262 -704 3280 -686 ne
rect 3280 -706 3302 -686
tri 3302 -706 3322 -686 sw
tri 3338 -700 3356 -682 ne
rect 3161 -776 3170 -742
rect 3204 -715 3246 -714
rect 3204 -749 3209 -715
rect 3239 -749 3246 -715
rect 3204 -758 3246 -749
rect 3280 -715 3322 -706
rect 3280 -749 3287 -715
rect 3317 -749 3322 -715
rect 3280 -754 3322 -749
rect 3356 -742 3384 -682
tri 3429 -695 3451 -673 se
rect 3451 -680 3466 -672
tri 3451 -695 3466 -680 nw
tri 3423 -701 3429 -695 se
rect 3429 -701 3438 -695
rect 3142 -786 3170 -776
tri 3170 -786 3194 -762 sw
rect 3088 -856 3104 -808
rect 3142 -818 3184 -786
tri 3201 -794 3202 -793 sw
rect 3201 -818 3202 -794
tri 3204 -795 3241 -758 ne
rect 3241 -786 3246 -758
tri 3246 -786 3272 -760 sw
rect 3356 -776 3365 -742
rect 3356 -786 3384 -776
rect 3241 -795 3325 -786
tri 3241 -814 3260 -795 ne
rect 3260 -814 3325 -795
rect 3142 -840 3202 -818
rect 3324 -818 3325 -814
rect 3342 -818 3384 -786
rect 3324 -840 3384 -818
rect 3230 -856 3247 -842
rect 3279 -856 3296 -842
tri 3067 -892 3089 -870 se
rect 3089 -877 3104 -856
tri 3089 -892 3104 -877 nw
rect 3423 -877 3438 -701
tri 3438 -708 3451 -695 nw
rect 3524 -776 3539 -548
tri 3061 -898 3067 -892 se
rect 3067 -898 3076 -892
rect 3061 -914 3076 -898
tri 3076 -905 3089 -892 nw
rect 3230 -900 3247 -886
rect 3279 -900 3296 -886
tri 3423 -892 3438 -877 ne
tri 3438 -892 3460 -870 sw
rect 3061 -950 3076 -942
rect 3142 -914 3202 -900
rect 3157 -924 3202 -914
rect 3157 -942 3185 -924
tri 3061 -965 3076 -950 ne
tri 3076 -965 3098 -943 sw
rect 3142 -952 3185 -942
rect 3200 -928 3202 -924
rect 3324 -914 3384 -900
tri 3438 -905 3451 -892 ne
rect 3451 -898 3460 -892
tri 3460 -898 3466 -892 sw
rect 3324 -924 3369 -914
rect 3200 -952 3274 -928
rect 3142 -956 3274 -952
tri 3274 -956 3302 -928 sw
rect 3324 -938 3326 -924
tri 3324 -940 3326 -938 ne
rect 3338 -942 3369 -924
rect 3338 -952 3384 -942
rect 3451 -913 3466 -898
tri 3076 -977 3088 -965 ne
rect 3088 -970 3098 -965
tri 3098 -970 3103 -965 sw
rect 2987 -1316 3002 -1088
rect 3088 -1126 3103 -970
rect 3142 -1012 3170 -956
tri 3262 -974 3280 -956 ne
rect 3280 -976 3302 -956
tri 3302 -976 3322 -956 sw
tri 3338 -970 3356 -952 ne
rect 3161 -1046 3170 -1012
rect 3204 -985 3246 -984
rect 3204 -1019 3209 -985
rect 3239 -1019 3246 -985
rect 3204 -1028 3246 -1019
rect 3280 -985 3322 -976
rect 3280 -1019 3287 -985
rect 3317 -1019 3322 -985
rect 3280 -1024 3322 -1019
rect 3356 -1012 3384 -952
tri 3429 -965 3451 -943 se
rect 3451 -950 3466 -942
tri 3451 -965 3466 -950 nw
tri 3423 -971 3429 -965 se
rect 3429 -971 3438 -965
rect 3142 -1056 3170 -1046
tri 3170 -1056 3194 -1032 sw
rect 3142 -1088 3184 -1056
tri 3201 -1064 3202 -1063 sw
rect 3201 -1088 3202 -1064
tri 3204 -1065 3241 -1028 ne
rect 3241 -1056 3246 -1028
tri 3246 -1056 3272 -1030 sw
rect 3356 -1046 3365 -1012
rect 3356 -1056 3384 -1046
rect 3241 -1065 3325 -1056
tri 3241 -1084 3260 -1065 ne
rect 3260 -1084 3325 -1065
rect 3142 -1110 3202 -1088
rect 3324 -1088 3325 -1084
rect 3342 -1088 3384 -1056
rect 3324 -1110 3384 -1088
rect 3230 -1126 3247 -1112
rect 3279 -1126 3296 -1112
tri 3067 -1162 3089 -1140 se
rect 3089 -1147 3104 -1126
tri 3089 -1162 3104 -1147 nw
rect 3423 -1147 3438 -971
tri 3438 -978 3451 -965 nw
rect 3524 -1046 3539 -818
tri 3061 -1168 3067 -1162 se
rect 3067 -1168 3076 -1162
rect 3061 -1184 3076 -1168
tri 3076 -1175 3089 -1162 nw
rect 3230 -1170 3247 -1156
rect 3279 -1170 3296 -1156
tri 3423 -1162 3438 -1147 ne
tri 3438 -1162 3460 -1140 sw
rect 3061 -1220 3076 -1212
rect 3142 -1184 3202 -1170
rect 3157 -1194 3202 -1184
rect 3157 -1212 3185 -1194
tri 3061 -1235 3076 -1220 ne
tri 3076 -1235 3098 -1213 sw
rect 3142 -1222 3185 -1212
rect 3200 -1198 3202 -1194
rect 3324 -1184 3384 -1170
tri 3438 -1175 3451 -1162 ne
rect 3451 -1168 3460 -1162
tri 3460 -1168 3466 -1162 sw
rect 3324 -1194 3369 -1184
rect 3200 -1222 3274 -1198
rect 3142 -1226 3274 -1222
tri 3274 -1226 3302 -1198 sw
rect 3324 -1208 3326 -1194
tri 3324 -1210 3326 -1208 ne
rect 3338 -1212 3369 -1194
rect 3338 -1222 3384 -1212
rect 3451 -1183 3466 -1168
tri 3076 -1247 3088 -1235 ne
rect 3088 -1240 3098 -1235
tri 3098 -1240 3103 -1235 sw
rect 2987 -1586 3002 -1358
rect 3088 -1348 3103 -1240
rect 3142 -1282 3170 -1226
tri 3262 -1244 3280 -1226 ne
rect 3280 -1246 3302 -1226
tri 3302 -1246 3322 -1226 sw
tri 3338 -1240 3356 -1222 ne
rect 3161 -1316 3170 -1282
rect 3204 -1255 3246 -1254
rect 3204 -1289 3209 -1255
rect 3239 -1289 3246 -1255
rect 3204 -1298 3246 -1289
rect 3280 -1255 3322 -1246
rect 3280 -1289 3287 -1255
rect 3317 -1289 3322 -1255
rect 3280 -1294 3322 -1289
rect 3356 -1282 3384 -1222
tri 3429 -1235 3451 -1213 se
rect 3451 -1220 3466 -1212
tri 3451 -1235 3466 -1220 nw
tri 3423 -1241 3429 -1235 se
rect 3429 -1241 3438 -1235
rect 3142 -1326 3170 -1316
tri 3170 -1326 3194 -1302 sw
rect 3088 -1396 3104 -1348
rect 3142 -1358 3184 -1326
tri 3201 -1334 3202 -1333 sw
rect 3201 -1358 3202 -1334
tri 3204 -1335 3241 -1298 ne
rect 3241 -1326 3246 -1298
tri 3246 -1326 3272 -1300 sw
rect 3356 -1316 3365 -1282
rect 3356 -1326 3384 -1316
rect 3241 -1335 3325 -1326
tri 3241 -1354 3260 -1335 ne
rect 3260 -1354 3325 -1335
rect 3142 -1380 3202 -1358
rect 3324 -1358 3325 -1354
rect 3342 -1358 3384 -1326
rect 3324 -1380 3384 -1358
rect 3230 -1396 3247 -1382
rect 3279 -1396 3296 -1382
tri 3067 -1432 3089 -1410 se
rect 3089 -1417 3104 -1396
tri 3089 -1432 3104 -1417 nw
rect 3423 -1417 3438 -1241
tri 3438 -1248 3451 -1235 nw
rect 3524 -1316 3539 -1088
tri 3061 -1438 3067 -1432 se
rect 3067 -1438 3076 -1432
rect 3061 -1454 3076 -1438
tri 3076 -1445 3089 -1432 nw
rect 3230 -1440 3247 -1426
rect 3279 -1440 3296 -1426
tri 3423 -1432 3438 -1417 ne
tri 3438 -1432 3460 -1410 sw
rect 3061 -1490 3076 -1482
rect 3142 -1454 3202 -1440
rect 3157 -1464 3202 -1454
rect 3157 -1482 3185 -1464
tri 3061 -1505 3076 -1490 ne
tri 3076 -1505 3098 -1483 sw
rect 3142 -1492 3185 -1482
rect 3200 -1468 3202 -1464
rect 3324 -1454 3384 -1440
tri 3438 -1445 3451 -1432 ne
rect 3451 -1438 3460 -1432
tri 3460 -1438 3466 -1432 sw
rect 3324 -1464 3369 -1454
rect 3200 -1492 3274 -1468
rect 3142 -1496 3274 -1492
tri 3274 -1496 3302 -1468 sw
rect 3324 -1478 3326 -1464
tri 3324 -1480 3326 -1478 ne
rect 3338 -1482 3369 -1464
rect 3338 -1492 3384 -1482
rect 3451 -1453 3466 -1438
tri 3076 -1517 3088 -1505 ne
rect 3088 -1510 3098 -1505
tri 3098 -1510 3103 -1505 sw
rect 2987 -1856 3002 -1628
rect 3088 -1666 3103 -1510
rect 3142 -1552 3170 -1496
tri 3262 -1514 3280 -1496 ne
rect 3280 -1516 3302 -1496
tri 3302 -1516 3322 -1496 sw
tri 3338 -1510 3356 -1492 ne
rect 3161 -1586 3170 -1552
rect 3204 -1525 3246 -1524
rect 3204 -1559 3209 -1525
rect 3239 -1559 3246 -1525
rect 3204 -1568 3246 -1559
rect 3280 -1525 3322 -1516
rect 3280 -1559 3287 -1525
rect 3317 -1559 3322 -1525
rect 3280 -1564 3322 -1559
rect 3356 -1552 3384 -1492
tri 3429 -1505 3451 -1483 se
rect 3451 -1490 3466 -1482
tri 3451 -1505 3466 -1490 nw
tri 3423 -1511 3429 -1505 se
rect 3429 -1511 3438 -1505
rect 3142 -1596 3170 -1586
tri 3170 -1596 3194 -1572 sw
rect 3142 -1628 3184 -1596
tri 3201 -1604 3202 -1603 sw
rect 3201 -1628 3202 -1604
tri 3204 -1605 3241 -1568 ne
rect 3241 -1596 3246 -1568
tri 3246 -1596 3272 -1570 sw
rect 3356 -1586 3365 -1552
rect 3356 -1596 3384 -1586
rect 3241 -1605 3325 -1596
tri 3241 -1624 3260 -1605 ne
rect 3260 -1624 3325 -1605
rect 3142 -1650 3202 -1628
rect 3324 -1628 3325 -1624
rect 3342 -1628 3384 -1596
rect 3324 -1650 3384 -1628
rect 3230 -1666 3247 -1652
rect 3279 -1666 3296 -1652
tri 3067 -1702 3089 -1680 se
rect 3089 -1687 3104 -1666
tri 3089 -1702 3104 -1687 nw
rect 3423 -1687 3438 -1511
tri 3438 -1518 3451 -1505 nw
rect 3524 -1586 3539 -1358
tri 3061 -1708 3067 -1702 se
rect 3067 -1708 3076 -1702
rect 3061 -1724 3076 -1708
tri 3076 -1715 3089 -1702 nw
rect 3230 -1710 3247 -1696
rect 3279 -1710 3296 -1696
tri 3423 -1702 3438 -1687 ne
tri 3438 -1702 3460 -1680 sw
rect 3061 -1760 3076 -1752
rect 3142 -1724 3202 -1710
rect 3157 -1734 3202 -1724
rect 3157 -1752 3185 -1734
tri 3061 -1775 3076 -1760 ne
tri 3076 -1775 3098 -1753 sw
rect 3142 -1762 3185 -1752
rect 3200 -1738 3202 -1734
rect 3324 -1724 3384 -1710
tri 3438 -1715 3451 -1702 ne
rect 3451 -1708 3460 -1702
tri 3460 -1708 3466 -1702 sw
rect 3324 -1734 3369 -1724
rect 3200 -1762 3274 -1738
rect 3142 -1766 3274 -1762
tri 3274 -1766 3302 -1738 sw
rect 3324 -1748 3326 -1734
tri 3324 -1750 3326 -1748 ne
rect 3338 -1752 3369 -1734
rect 3338 -1762 3384 -1752
rect 3451 -1723 3466 -1708
tri 3076 -1787 3088 -1775 ne
rect 3088 -1780 3098 -1775
tri 3098 -1780 3103 -1775 sw
rect 2987 -2126 3002 -1898
rect 3088 -1888 3103 -1780
rect 3142 -1822 3170 -1766
tri 3262 -1784 3280 -1766 ne
rect 3280 -1786 3302 -1766
tri 3302 -1786 3322 -1766 sw
tri 3338 -1780 3356 -1762 ne
rect 3161 -1856 3170 -1822
rect 3204 -1795 3246 -1794
rect 3204 -1829 3209 -1795
rect 3239 -1829 3246 -1795
rect 3204 -1838 3246 -1829
rect 3280 -1795 3322 -1786
rect 3280 -1829 3287 -1795
rect 3317 -1829 3322 -1795
rect 3280 -1834 3322 -1829
rect 3356 -1822 3384 -1762
tri 3429 -1775 3451 -1753 se
rect 3451 -1760 3466 -1752
tri 3451 -1775 3466 -1760 nw
tri 3423 -1781 3429 -1775 se
rect 3429 -1781 3438 -1775
rect 3142 -1866 3170 -1856
tri 3170 -1866 3194 -1842 sw
rect 3088 -1936 3104 -1888
rect 3142 -1898 3184 -1866
tri 3201 -1874 3202 -1873 sw
rect 3201 -1898 3202 -1874
tri 3204 -1875 3241 -1838 ne
rect 3241 -1866 3246 -1838
tri 3246 -1866 3272 -1840 sw
rect 3356 -1856 3365 -1822
rect 3356 -1866 3384 -1856
rect 3241 -1875 3325 -1866
tri 3241 -1894 3260 -1875 ne
rect 3260 -1894 3325 -1875
rect 3142 -1920 3202 -1898
rect 3324 -1898 3325 -1894
rect 3342 -1898 3384 -1866
rect 3324 -1920 3384 -1898
rect 3230 -1936 3247 -1922
rect 3279 -1936 3296 -1922
tri 3067 -1972 3089 -1950 se
rect 3089 -1957 3104 -1936
tri 3089 -1972 3104 -1957 nw
rect 3423 -1957 3438 -1781
tri 3438 -1788 3451 -1775 nw
rect 3524 -1856 3539 -1628
tri 3061 -1978 3067 -1972 se
rect 3067 -1978 3076 -1972
rect 3061 -1994 3076 -1978
tri 3076 -1985 3089 -1972 nw
rect 3230 -1980 3247 -1966
rect 3279 -1980 3296 -1966
tri 3423 -1972 3438 -1957 ne
tri 3438 -1972 3460 -1950 sw
rect 3061 -2030 3076 -2022
rect 3142 -1994 3202 -1980
rect 3157 -2004 3202 -1994
rect 3157 -2022 3185 -2004
tri 3061 -2045 3076 -2030 ne
tri 3076 -2045 3098 -2023 sw
rect 3142 -2032 3185 -2022
rect 3200 -2008 3202 -2004
rect 3324 -1994 3384 -1980
tri 3438 -1985 3451 -1972 ne
rect 3451 -1978 3460 -1972
tri 3460 -1978 3466 -1972 sw
rect 3324 -2004 3369 -1994
rect 3200 -2032 3274 -2008
rect 3142 -2036 3274 -2032
tri 3274 -2036 3302 -2008 sw
rect 3324 -2018 3326 -2004
tri 3324 -2020 3326 -2018 ne
rect 3338 -2022 3369 -2004
rect 3338 -2032 3384 -2022
rect 3451 -1993 3466 -1978
tri 3076 -2057 3088 -2045 ne
rect 3088 -2050 3098 -2045
tri 3098 -2050 3103 -2045 sw
rect 2987 -2396 3002 -2168
rect 3088 -2206 3103 -2050
rect 3142 -2092 3170 -2036
tri 3262 -2054 3280 -2036 ne
rect 3280 -2056 3302 -2036
tri 3302 -2056 3322 -2036 sw
tri 3338 -2050 3356 -2032 ne
rect 3161 -2126 3170 -2092
rect 3204 -2065 3246 -2064
rect 3204 -2099 3209 -2065
rect 3239 -2099 3246 -2065
rect 3204 -2108 3246 -2099
rect 3280 -2065 3322 -2056
rect 3280 -2099 3287 -2065
rect 3317 -2099 3322 -2065
rect 3280 -2104 3322 -2099
rect 3356 -2092 3384 -2032
tri 3429 -2045 3451 -2023 se
rect 3451 -2030 3466 -2022
tri 3451 -2045 3466 -2030 nw
tri 3423 -2051 3429 -2045 se
rect 3429 -2051 3438 -2045
rect 3142 -2136 3170 -2126
tri 3170 -2136 3194 -2112 sw
rect 3142 -2168 3184 -2136
tri 3201 -2144 3202 -2143 sw
rect 3201 -2168 3202 -2144
tri 3204 -2145 3241 -2108 ne
rect 3241 -2136 3246 -2108
tri 3246 -2136 3272 -2110 sw
rect 3356 -2126 3365 -2092
rect 3356 -2136 3384 -2126
rect 3241 -2145 3325 -2136
tri 3241 -2164 3260 -2145 ne
rect 3260 -2164 3325 -2145
rect 3142 -2190 3202 -2168
rect 3324 -2168 3325 -2164
rect 3342 -2168 3384 -2136
rect 3324 -2190 3384 -2168
rect 3230 -2206 3247 -2192
rect 3279 -2206 3296 -2192
tri 3067 -2242 3089 -2220 se
rect 3089 -2227 3104 -2206
tri 3089 -2242 3104 -2227 nw
rect 3423 -2227 3438 -2051
tri 3438 -2058 3451 -2045 nw
rect 3524 -2126 3539 -1898
tri 3061 -2248 3067 -2242 se
rect 3067 -2248 3076 -2242
rect 3061 -2264 3076 -2248
tri 3076 -2255 3089 -2242 nw
rect 3230 -2250 3247 -2236
rect 3279 -2250 3296 -2236
tri 3423 -2242 3438 -2227 ne
tri 3438 -2242 3460 -2220 sw
rect 3061 -2300 3076 -2292
rect 3142 -2264 3202 -2250
rect 3157 -2274 3202 -2264
rect 3157 -2292 3185 -2274
tri 3061 -2315 3076 -2300 ne
tri 3076 -2315 3098 -2293 sw
rect 3142 -2302 3185 -2292
rect 3200 -2278 3202 -2274
rect 3324 -2264 3384 -2250
tri 3438 -2255 3451 -2242 ne
rect 3451 -2248 3460 -2242
tri 3460 -2248 3466 -2242 sw
rect 3324 -2274 3369 -2264
rect 3200 -2302 3274 -2278
rect 3142 -2306 3274 -2302
tri 3274 -2306 3302 -2278 sw
rect 3324 -2288 3326 -2274
tri 3324 -2290 3326 -2288 ne
rect 3338 -2292 3369 -2274
rect 3338 -2302 3384 -2292
rect 3451 -2263 3466 -2248
tri 3076 -2327 3088 -2315 ne
rect 3088 -2320 3098 -2315
tri 3098 -2320 3103 -2315 sw
rect 2987 -2524 3002 -2438
rect 3088 -2476 3103 -2320
rect 3142 -2362 3170 -2306
tri 3262 -2324 3280 -2306 ne
rect 3280 -2326 3302 -2306
tri 3302 -2326 3322 -2306 sw
tri 3338 -2320 3356 -2302 ne
rect 3161 -2396 3170 -2362
rect 3204 -2335 3246 -2334
rect 3204 -2369 3209 -2335
rect 3239 -2369 3246 -2335
rect 3204 -2378 3246 -2369
rect 3280 -2335 3322 -2326
rect 3280 -2369 3287 -2335
rect 3317 -2369 3322 -2335
rect 3280 -2374 3322 -2369
rect 3356 -2362 3384 -2302
tri 3429 -2315 3451 -2293 se
rect 3451 -2300 3466 -2292
tri 3451 -2315 3466 -2300 nw
tri 3423 -2321 3429 -2315 se
rect 3429 -2321 3438 -2315
rect 3142 -2406 3170 -2396
tri 3170 -2406 3194 -2382 sw
rect 3142 -2438 3184 -2406
tri 3201 -2414 3202 -2413 sw
rect 3201 -2438 3202 -2414
tri 3204 -2415 3241 -2378 ne
rect 3241 -2406 3246 -2378
tri 3246 -2406 3272 -2380 sw
rect 3356 -2396 3365 -2362
rect 3356 -2406 3384 -2396
rect 3241 -2415 3325 -2406
tri 3241 -2434 3260 -2415 ne
rect 3260 -2434 3325 -2415
rect 3142 -2460 3202 -2438
rect 3324 -2438 3325 -2434
rect 3342 -2438 3384 -2406
rect 3324 -2460 3384 -2438
rect 3230 -2476 3247 -2462
rect 3279 -2476 3296 -2462
rect 3423 -2476 3438 -2321
tri 3438 -2328 3451 -2315 nw
rect 3524 -2396 3539 -2168
rect 3524 -2524 3539 -2438
rect 3567 1654 3582 1844
tri 3647 1808 3669 1830 se
rect 3669 1823 3684 1892
tri 3669 1808 3684 1823 nw
rect 4003 1823 4018 1892
tri 3641 1802 3647 1808 se
rect 3647 1802 3656 1808
rect 3641 1786 3656 1802
tri 3656 1795 3669 1808 nw
rect 3810 1800 3827 1814
rect 3859 1800 3876 1814
tri 4003 1808 4018 1823 ne
tri 4018 1808 4040 1830 sw
rect 3641 1750 3656 1758
rect 3722 1786 3782 1800
rect 3737 1776 3782 1786
rect 3737 1758 3765 1776
tri 3641 1735 3656 1750 ne
tri 3656 1735 3678 1757 sw
rect 3722 1748 3765 1758
rect 3780 1772 3782 1776
rect 3904 1786 3964 1800
tri 4018 1795 4031 1808 ne
rect 4031 1802 4040 1808
tri 4040 1802 4046 1808 sw
rect 3904 1776 3949 1786
rect 3780 1748 3854 1772
rect 3722 1744 3854 1748
tri 3854 1744 3882 1772 sw
rect 3904 1762 3906 1776
tri 3904 1760 3906 1762 ne
rect 3918 1758 3949 1776
rect 3918 1748 3964 1758
rect 4031 1787 4046 1802
tri 3656 1723 3668 1735 ne
rect 3668 1730 3678 1735
tri 3678 1730 3683 1735 sw
rect 3567 1384 3582 1612
rect 3668 1574 3683 1730
rect 3722 1688 3750 1744
tri 3842 1726 3860 1744 ne
rect 3860 1724 3882 1744
tri 3882 1724 3902 1744 sw
tri 3918 1730 3936 1748 ne
rect 3741 1654 3750 1688
rect 3784 1715 3826 1716
rect 3784 1681 3789 1715
rect 3819 1681 3826 1715
rect 3784 1672 3826 1681
rect 3860 1715 3902 1724
rect 3860 1681 3867 1715
rect 3897 1681 3902 1715
rect 3860 1676 3902 1681
rect 3936 1688 3964 1748
tri 4009 1735 4031 1757 se
rect 4031 1750 4046 1758
tri 4031 1735 4046 1750 nw
tri 4003 1729 4009 1735 se
rect 4009 1729 4018 1735
rect 3722 1644 3750 1654
tri 3750 1644 3774 1668 sw
rect 3722 1612 3764 1644
tri 3781 1636 3782 1637 sw
rect 3781 1612 3782 1636
tri 3784 1635 3821 1672 ne
rect 3821 1644 3826 1672
tri 3826 1644 3852 1670 sw
rect 3936 1654 3945 1688
rect 3936 1644 3964 1654
rect 3821 1635 3905 1644
tri 3821 1616 3840 1635 ne
rect 3840 1616 3905 1635
rect 3722 1590 3782 1612
rect 3904 1612 3905 1616
rect 3922 1612 3964 1644
rect 3904 1590 3964 1612
rect 3810 1574 3827 1588
rect 3859 1574 3876 1588
tri 3647 1538 3669 1560 se
rect 3669 1553 3684 1574
tri 3669 1538 3684 1553 nw
rect 4003 1553 4018 1729
tri 4018 1722 4031 1735 nw
rect 4104 1654 4119 1844
tri 3641 1532 3647 1538 se
rect 3647 1532 3656 1538
rect 3641 1516 3656 1532
tri 3656 1525 3669 1538 nw
rect 3810 1530 3827 1544
rect 3859 1530 3876 1544
tri 4003 1538 4018 1553 ne
tri 4018 1538 4040 1560 sw
rect 3641 1480 3656 1488
rect 3722 1516 3782 1530
rect 3737 1506 3782 1516
rect 3737 1488 3765 1506
tri 3641 1465 3656 1480 ne
tri 3656 1465 3678 1487 sw
rect 3722 1478 3765 1488
rect 3780 1502 3782 1506
rect 3904 1516 3964 1530
tri 4018 1525 4031 1538 ne
rect 4031 1532 4040 1538
tri 4040 1532 4046 1538 sw
rect 3904 1506 3949 1516
rect 3780 1478 3854 1502
rect 3722 1474 3854 1478
tri 3854 1474 3882 1502 sw
rect 3904 1492 3906 1506
tri 3904 1490 3906 1492 ne
rect 3918 1488 3949 1506
rect 3918 1478 3964 1488
rect 4031 1517 4046 1532
tri 3656 1453 3668 1465 ne
rect 3668 1460 3678 1465
tri 3678 1460 3683 1465 sw
rect 3567 1114 3582 1342
rect 3668 1352 3683 1460
rect 3722 1418 3750 1474
tri 3842 1456 3860 1474 ne
rect 3860 1454 3882 1474
tri 3882 1454 3902 1474 sw
tri 3918 1460 3936 1478 ne
rect 3741 1384 3750 1418
rect 3784 1445 3826 1446
rect 3784 1411 3789 1445
rect 3819 1411 3826 1445
rect 3784 1402 3826 1411
rect 3860 1445 3902 1454
rect 3860 1411 3867 1445
rect 3897 1411 3902 1445
rect 3860 1406 3902 1411
rect 3936 1418 3964 1478
tri 4009 1465 4031 1487 se
rect 4031 1480 4046 1488
tri 4031 1465 4046 1480 nw
tri 4003 1459 4009 1465 se
rect 4009 1459 4018 1465
rect 3722 1374 3750 1384
tri 3750 1374 3774 1398 sw
rect 3668 1304 3684 1352
rect 3722 1342 3764 1374
tri 3781 1366 3782 1367 sw
rect 3781 1342 3782 1366
tri 3784 1365 3821 1402 ne
rect 3821 1374 3826 1402
tri 3826 1374 3852 1400 sw
rect 3936 1384 3945 1418
rect 3936 1374 3964 1384
rect 3821 1365 3905 1374
tri 3821 1346 3840 1365 ne
rect 3840 1346 3905 1365
rect 3722 1320 3782 1342
rect 3904 1342 3905 1346
rect 3922 1342 3964 1374
rect 3904 1320 3964 1342
rect 3810 1304 3827 1318
rect 3859 1304 3876 1318
tri 3647 1268 3669 1290 se
rect 3669 1283 3684 1304
tri 3669 1268 3684 1283 nw
rect 4003 1283 4018 1459
tri 4018 1452 4031 1465 nw
rect 4104 1384 4119 1612
tri 3641 1262 3647 1268 se
rect 3647 1262 3656 1268
rect 3641 1246 3656 1262
tri 3656 1255 3669 1268 nw
rect 3810 1260 3827 1274
rect 3859 1260 3876 1274
tri 4003 1268 4018 1283 ne
tri 4018 1268 4040 1290 sw
rect 3641 1210 3656 1218
rect 3722 1246 3782 1260
rect 3737 1236 3782 1246
rect 3737 1218 3765 1236
tri 3641 1195 3656 1210 ne
tri 3656 1195 3678 1217 sw
rect 3722 1208 3765 1218
rect 3780 1232 3782 1236
rect 3904 1246 3964 1260
tri 4018 1255 4031 1268 ne
rect 4031 1262 4040 1268
tri 4040 1262 4046 1268 sw
rect 3904 1236 3949 1246
rect 3780 1208 3854 1232
rect 3722 1204 3854 1208
tri 3854 1204 3882 1232 sw
rect 3904 1222 3906 1236
tri 3904 1220 3906 1222 ne
rect 3918 1218 3949 1236
rect 3918 1208 3964 1218
rect 4031 1247 4046 1262
tri 3656 1183 3668 1195 ne
rect 3668 1190 3678 1195
tri 3678 1190 3683 1195 sw
rect 3567 844 3582 1072
rect 3668 1034 3683 1190
rect 3722 1148 3750 1204
tri 3842 1186 3860 1204 ne
rect 3860 1184 3882 1204
tri 3882 1184 3902 1204 sw
tri 3918 1190 3936 1208 ne
rect 3741 1114 3750 1148
rect 3784 1175 3826 1176
rect 3784 1141 3789 1175
rect 3819 1141 3826 1175
rect 3784 1132 3826 1141
rect 3860 1175 3902 1184
rect 3860 1141 3867 1175
rect 3897 1141 3902 1175
rect 3860 1136 3902 1141
rect 3936 1148 3964 1208
tri 4009 1195 4031 1217 se
rect 4031 1210 4046 1218
tri 4031 1195 4046 1210 nw
tri 4003 1189 4009 1195 se
rect 4009 1189 4018 1195
rect 3722 1104 3750 1114
tri 3750 1104 3774 1128 sw
rect 3722 1072 3764 1104
tri 3781 1096 3782 1097 sw
rect 3781 1072 3782 1096
tri 3784 1095 3821 1132 ne
rect 3821 1104 3826 1132
tri 3826 1104 3852 1130 sw
rect 3936 1114 3945 1148
rect 3936 1104 3964 1114
rect 3821 1095 3905 1104
tri 3821 1076 3840 1095 ne
rect 3840 1076 3905 1095
rect 3722 1050 3782 1072
rect 3904 1072 3905 1076
rect 3922 1072 3964 1104
rect 3904 1050 3964 1072
rect 3810 1034 3827 1048
rect 3859 1034 3876 1048
tri 3647 998 3669 1020 se
rect 3669 1013 3684 1034
tri 3669 998 3684 1013 nw
rect 4003 1013 4018 1189
tri 4018 1182 4031 1195 nw
rect 4104 1114 4119 1342
tri 3641 992 3647 998 se
rect 3647 992 3656 998
rect 3641 976 3656 992
tri 3656 985 3669 998 nw
rect 3810 990 3827 1004
rect 3859 990 3876 1004
tri 4003 998 4018 1013 ne
tri 4018 998 4040 1020 sw
rect 3641 940 3656 948
rect 3722 976 3782 990
rect 3737 966 3782 976
rect 3737 948 3765 966
tri 3641 925 3656 940 ne
tri 3656 925 3678 947 sw
rect 3722 938 3765 948
rect 3780 962 3782 966
rect 3904 976 3964 990
tri 4018 985 4031 998 ne
rect 4031 992 4040 998
tri 4040 992 4046 998 sw
rect 3904 966 3949 976
rect 3780 938 3854 962
rect 3722 934 3854 938
tri 3854 934 3882 962 sw
rect 3904 952 3906 966
tri 3904 950 3906 952 ne
rect 3918 948 3949 966
rect 3918 938 3964 948
rect 4031 977 4046 992
tri 3656 913 3668 925 ne
rect 3668 920 3678 925
tri 3678 920 3683 925 sw
rect 3567 574 3582 802
rect 3668 812 3683 920
rect 3722 878 3750 934
tri 3842 916 3860 934 ne
rect 3860 914 3882 934
tri 3882 914 3902 934 sw
tri 3918 920 3936 938 ne
rect 3741 844 3750 878
rect 3784 905 3826 906
rect 3784 871 3789 905
rect 3819 871 3826 905
rect 3784 862 3826 871
rect 3860 905 3902 914
rect 3860 871 3867 905
rect 3897 871 3902 905
rect 3860 866 3902 871
rect 3936 878 3964 938
tri 4009 925 4031 947 se
rect 4031 940 4046 948
tri 4031 925 4046 940 nw
tri 4003 919 4009 925 se
rect 4009 919 4018 925
rect 3722 834 3750 844
tri 3750 834 3774 858 sw
rect 3668 764 3684 812
rect 3722 802 3764 834
tri 3781 826 3782 827 sw
rect 3781 802 3782 826
tri 3784 825 3821 862 ne
rect 3821 834 3826 862
tri 3826 834 3852 860 sw
rect 3936 844 3945 878
rect 3936 834 3964 844
rect 3821 825 3905 834
tri 3821 806 3840 825 ne
rect 3840 806 3905 825
rect 3722 780 3782 802
rect 3904 802 3905 806
rect 3922 802 3964 834
rect 3904 780 3964 802
rect 3810 764 3827 778
rect 3859 764 3876 778
tri 3647 728 3669 750 se
rect 3669 743 3684 764
tri 3669 728 3684 743 nw
rect 4003 743 4018 919
tri 4018 912 4031 925 nw
rect 4104 844 4119 1072
tri 3641 722 3647 728 se
rect 3647 722 3656 728
rect 3641 706 3656 722
tri 3656 715 3669 728 nw
rect 3810 720 3827 734
rect 3859 720 3876 734
tri 4003 728 4018 743 ne
tri 4018 728 4040 750 sw
rect 3641 670 3656 678
rect 3722 706 3782 720
rect 3737 696 3782 706
rect 3737 678 3765 696
tri 3641 655 3656 670 ne
tri 3656 655 3678 677 sw
rect 3722 668 3765 678
rect 3780 692 3782 696
rect 3904 706 3964 720
tri 4018 715 4031 728 ne
rect 4031 722 4040 728
tri 4040 722 4046 728 sw
rect 3904 696 3949 706
rect 3780 668 3854 692
rect 3722 664 3854 668
tri 3854 664 3882 692 sw
rect 3904 682 3906 696
tri 3904 680 3906 682 ne
rect 3918 678 3949 696
rect 3918 668 3964 678
rect 4031 707 4046 722
tri 3656 643 3668 655 ne
rect 3668 650 3678 655
tri 3678 650 3683 655 sw
rect 3567 304 3582 532
rect 3668 494 3683 650
rect 3722 608 3750 664
tri 3842 646 3860 664 ne
rect 3860 644 3882 664
tri 3882 644 3902 664 sw
tri 3918 650 3936 668 ne
rect 3741 574 3750 608
rect 3784 635 3826 636
rect 3784 601 3789 635
rect 3819 601 3826 635
rect 3784 592 3826 601
rect 3860 635 3902 644
rect 3860 601 3867 635
rect 3897 601 3902 635
rect 3860 596 3902 601
rect 3936 608 3964 668
tri 4009 655 4031 677 se
rect 4031 670 4046 678
tri 4031 655 4046 670 nw
tri 4003 649 4009 655 se
rect 4009 649 4018 655
rect 3722 564 3750 574
tri 3750 564 3774 588 sw
rect 3722 532 3764 564
tri 3781 556 3782 557 sw
rect 3781 532 3782 556
tri 3784 555 3821 592 ne
rect 3821 564 3826 592
tri 3826 564 3852 590 sw
rect 3936 574 3945 608
rect 3936 564 3964 574
rect 3821 555 3905 564
tri 3821 536 3840 555 ne
rect 3840 536 3905 555
rect 3722 510 3782 532
rect 3904 532 3905 536
rect 3922 532 3964 564
rect 3904 510 3964 532
rect 3810 494 3827 508
rect 3859 494 3876 508
tri 3647 458 3669 480 se
rect 3669 473 3684 494
tri 3669 458 3684 473 nw
rect 4003 473 4018 649
tri 4018 642 4031 655 nw
rect 4104 574 4119 802
tri 3641 452 3647 458 se
rect 3647 452 3656 458
rect 3641 436 3656 452
tri 3656 445 3669 458 nw
rect 3810 450 3827 464
rect 3859 450 3876 464
tri 4003 458 4018 473 ne
tri 4018 458 4040 480 sw
rect 3641 400 3656 408
rect 3722 436 3782 450
rect 3737 426 3782 436
rect 3737 408 3765 426
tri 3641 385 3656 400 ne
tri 3656 385 3678 407 sw
rect 3722 398 3765 408
rect 3780 422 3782 426
rect 3904 436 3964 450
tri 4018 445 4031 458 ne
rect 4031 452 4040 458
tri 4040 452 4046 458 sw
rect 3904 426 3949 436
rect 3780 398 3854 422
rect 3722 394 3854 398
tri 3854 394 3882 422 sw
rect 3904 412 3906 426
tri 3904 410 3906 412 ne
rect 3918 408 3949 426
rect 3918 398 3964 408
rect 4031 437 4046 452
tri 3656 373 3668 385 ne
rect 3668 380 3678 385
tri 3678 380 3683 385 sw
rect 3567 34 3582 262
rect 3668 272 3683 380
rect 3722 338 3750 394
tri 3842 376 3860 394 ne
rect 3860 374 3882 394
tri 3882 374 3902 394 sw
tri 3918 380 3936 398 ne
rect 3741 304 3750 338
rect 3784 365 3826 366
rect 3784 331 3789 365
rect 3819 331 3826 365
rect 3784 322 3826 331
rect 3860 365 3902 374
rect 3860 331 3867 365
rect 3897 331 3902 365
rect 3860 326 3902 331
rect 3936 338 3964 398
tri 4009 385 4031 407 se
rect 4031 400 4046 408
tri 4031 385 4046 400 nw
tri 4003 379 4009 385 se
rect 4009 379 4018 385
rect 3722 294 3750 304
tri 3750 294 3774 318 sw
rect 3668 224 3684 272
rect 3722 262 3764 294
tri 3781 286 3782 287 sw
rect 3781 262 3782 286
tri 3784 285 3821 322 ne
rect 3821 294 3826 322
tri 3826 294 3852 320 sw
rect 3936 304 3945 338
rect 3936 294 3964 304
rect 3821 285 3905 294
tri 3821 266 3840 285 ne
rect 3840 266 3905 285
rect 3722 240 3782 262
rect 3904 262 3905 266
rect 3922 262 3964 294
rect 3904 240 3964 262
rect 3810 224 3827 238
rect 3859 224 3876 238
tri 3647 188 3669 210 se
rect 3669 203 3684 224
tri 3669 188 3684 203 nw
rect 4003 203 4018 379
tri 4018 372 4031 385 nw
rect 4104 304 4119 532
tri 3641 182 3647 188 se
rect 3647 182 3656 188
rect 3641 166 3656 182
tri 3656 175 3669 188 nw
rect 3810 180 3827 194
rect 3859 180 3876 194
tri 4003 188 4018 203 ne
tri 4018 188 4040 210 sw
rect 3641 130 3656 138
rect 3722 166 3782 180
rect 3737 156 3782 166
rect 3737 138 3765 156
tri 3641 115 3656 130 ne
tri 3656 115 3678 137 sw
rect 3722 128 3765 138
rect 3780 152 3782 156
rect 3904 166 3964 180
tri 4018 175 4031 188 ne
rect 4031 182 4040 188
tri 4040 182 4046 188 sw
rect 3904 156 3949 166
rect 3780 128 3854 152
rect 3722 124 3854 128
tri 3854 124 3882 152 sw
rect 3904 142 3906 156
tri 3904 140 3906 142 ne
rect 3918 138 3949 156
rect 3918 128 3964 138
rect 4031 167 4046 182
tri 3656 103 3668 115 ne
rect 3668 110 3678 115
tri 3678 110 3683 115 sw
rect 3567 -236 3582 -8
rect 3668 -46 3683 110
rect 3722 68 3750 124
tri 3842 106 3860 124 ne
rect 3860 104 3882 124
tri 3882 104 3902 124 sw
tri 3918 110 3936 128 ne
rect 3741 34 3750 68
rect 3784 95 3826 96
rect 3784 61 3789 95
rect 3819 61 3826 95
rect 3784 52 3826 61
rect 3860 95 3902 104
rect 3860 61 3867 95
rect 3897 61 3902 95
rect 3860 56 3902 61
rect 3936 68 3964 128
tri 4009 115 4031 137 se
rect 4031 130 4046 138
tri 4031 115 4046 130 nw
tri 4003 109 4009 115 se
rect 4009 109 4018 115
rect 3722 24 3750 34
tri 3750 24 3774 48 sw
rect 3722 -8 3764 24
tri 3781 16 3782 17 sw
rect 3781 -8 3782 16
tri 3784 15 3821 52 ne
rect 3821 24 3826 52
tri 3826 24 3852 50 sw
rect 3936 34 3945 68
rect 3936 24 3964 34
rect 3821 15 3905 24
tri 3821 -4 3840 15 ne
rect 3840 -4 3905 15
rect 3722 -30 3782 -8
rect 3904 -8 3905 -4
rect 3922 -8 3964 24
rect 3904 -30 3964 -8
rect 3810 -46 3827 -32
rect 3859 -46 3876 -32
tri 3647 -82 3669 -60 se
rect 3669 -67 3684 -46
tri 3669 -82 3684 -67 nw
rect 4003 -67 4018 109
tri 4018 102 4031 115 nw
rect 4104 34 4119 262
tri 3641 -88 3647 -82 se
rect 3647 -88 3656 -82
rect 3641 -104 3656 -88
tri 3656 -95 3669 -82 nw
rect 3810 -90 3827 -76
rect 3859 -90 3876 -76
tri 4003 -82 4018 -67 ne
tri 4018 -82 4040 -60 sw
rect 3641 -140 3656 -132
rect 3722 -104 3782 -90
rect 3737 -114 3782 -104
rect 3737 -132 3765 -114
tri 3641 -155 3656 -140 ne
tri 3656 -155 3678 -133 sw
rect 3722 -142 3765 -132
rect 3780 -118 3782 -114
rect 3904 -104 3964 -90
tri 4018 -95 4031 -82 ne
rect 4031 -88 4040 -82
tri 4040 -88 4046 -82 sw
rect 3904 -114 3949 -104
rect 3780 -142 3854 -118
rect 3722 -146 3854 -142
tri 3854 -146 3882 -118 sw
rect 3904 -128 3906 -114
tri 3904 -130 3906 -128 ne
rect 3918 -132 3949 -114
rect 3918 -142 3964 -132
rect 4031 -103 4046 -88
tri 3656 -167 3668 -155 ne
rect 3668 -160 3678 -155
tri 3678 -160 3683 -155 sw
rect 3567 -506 3582 -278
rect 3668 -268 3683 -160
rect 3722 -202 3750 -146
tri 3842 -164 3860 -146 ne
rect 3860 -166 3882 -146
tri 3882 -166 3902 -146 sw
tri 3918 -160 3936 -142 ne
rect 3741 -236 3750 -202
rect 3784 -175 3826 -174
rect 3784 -209 3789 -175
rect 3819 -209 3826 -175
rect 3784 -218 3826 -209
rect 3860 -175 3902 -166
rect 3860 -209 3867 -175
rect 3897 -209 3902 -175
rect 3860 -214 3902 -209
rect 3936 -202 3964 -142
tri 4009 -155 4031 -133 se
rect 4031 -140 4046 -132
tri 4031 -155 4046 -140 nw
tri 4003 -161 4009 -155 se
rect 4009 -161 4018 -155
rect 3722 -246 3750 -236
tri 3750 -246 3774 -222 sw
rect 3668 -316 3684 -268
rect 3722 -278 3764 -246
tri 3781 -254 3782 -253 sw
rect 3781 -278 3782 -254
tri 3784 -255 3821 -218 ne
rect 3821 -246 3826 -218
tri 3826 -246 3852 -220 sw
rect 3936 -236 3945 -202
rect 3936 -246 3964 -236
rect 3821 -255 3905 -246
tri 3821 -274 3840 -255 ne
rect 3840 -274 3905 -255
rect 3722 -300 3782 -278
rect 3904 -278 3905 -274
rect 3922 -278 3964 -246
rect 3904 -300 3964 -278
rect 3810 -316 3827 -302
rect 3859 -316 3876 -302
tri 3647 -352 3669 -330 se
rect 3669 -337 3684 -316
tri 3669 -352 3684 -337 nw
rect 4003 -337 4018 -161
tri 4018 -168 4031 -155 nw
rect 4104 -236 4119 -8
tri 3641 -358 3647 -352 se
rect 3647 -358 3656 -352
rect 3641 -374 3656 -358
tri 3656 -365 3669 -352 nw
rect 3810 -360 3827 -346
rect 3859 -360 3876 -346
tri 4003 -352 4018 -337 ne
tri 4018 -352 4040 -330 sw
rect 3641 -410 3656 -402
rect 3722 -374 3782 -360
rect 3737 -384 3782 -374
rect 3737 -402 3765 -384
tri 3641 -425 3656 -410 ne
tri 3656 -425 3678 -403 sw
rect 3722 -412 3765 -402
rect 3780 -388 3782 -384
rect 3904 -374 3964 -360
tri 4018 -365 4031 -352 ne
rect 4031 -358 4040 -352
tri 4040 -358 4046 -352 sw
rect 3904 -384 3949 -374
rect 3780 -412 3854 -388
rect 3722 -416 3854 -412
tri 3854 -416 3882 -388 sw
rect 3904 -398 3906 -384
tri 3904 -400 3906 -398 ne
rect 3918 -402 3949 -384
rect 3918 -412 3964 -402
rect 4031 -373 4046 -358
tri 3656 -437 3668 -425 ne
rect 3668 -430 3678 -425
tri 3678 -430 3683 -425 sw
rect 3567 -776 3582 -548
rect 3668 -586 3683 -430
rect 3722 -472 3750 -416
tri 3842 -434 3860 -416 ne
rect 3860 -436 3882 -416
tri 3882 -436 3902 -416 sw
tri 3918 -430 3936 -412 ne
rect 3741 -506 3750 -472
rect 3784 -445 3826 -444
rect 3784 -479 3789 -445
rect 3819 -479 3826 -445
rect 3784 -488 3826 -479
rect 3860 -445 3902 -436
rect 3860 -479 3867 -445
rect 3897 -479 3902 -445
rect 3860 -484 3902 -479
rect 3936 -472 3964 -412
tri 4009 -425 4031 -403 se
rect 4031 -410 4046 -402
tri 4031 -425 4046 -410 nw
tri 4003 -431 4009 -425 se
rect 4009 -431 4018 -425
rect 3722 -516 3750 -506
tri 3750 -516 3774 -492 sw
rect 3722 -548 3764 -516
tri 3781 -524 3782 -523 sw
rect 3781 -548 3782 -524
tri 3784 -525 3821 -488 ne
rect 3821 -516 3826 -488
tri 3826 -516 3852 -490 sw
rect 3936 -506 3945 -472
rect 3936 -516 3964 -506
rect 3821 -525 3905 -516
tri 3821 -544 3840 -525 ne
rect 3840 -544 3905 -525
rect 3722 -570 3782 -548
rect 3904 -548 3905 -544
rect 3922 -548 3964 -516
rect 3904 -570 3964 -548
rect 3810 -586 3827 -572
rect 3859 -586 3876 -572
tri 3647 -622 3669 -600 se
rect 3669 -607 3684 -586
tri 3669 -622 3684 -607 nw
rect 4003 -607 4018 -431
tri 4018 -438 4031 -425 nw
rect 4104 -506 4119 -278
tri 3641 -628 3647 -622 se
rect 3647 -628 3656 -622
rect 3641 -644 3656 -628
tri 3656 -635 3669 -622 nw
rect 3810 -630 3827 -616
rect 3859 -630 3876 -616
tri 4003 -622 4018 -607 ne
tri 4018 -622 4040 -600 sw
rect 3641 -680 3656 -672
rect 3722 -644 3782 -630
rect 3737 -654 3782 -644
rect 3737 -672 3765 -654
tri 3641 -695 3656 -680 ne
tri 3656 -695 3678 -673 sw
rect 3722 -682 3765 -672
rect 3780 -658 3782 -654
rect 3904 -644 3964 -630
tri 4018 -635 4031 -622 ne
rect 4031 -628 4040 -622
tri 4040 -628 4046 -622 sw
rect 3904 -654 3949 -644
rect 3780 -682 3854 -658
rect 3722 -686 3854 -682
tri 3854 -686 3882 -658 sw
rect 3904 -668 3906 -654
tri 3904 -670 3906 -668 ne
rect 3918 -672 3949 -654
rect 3918 -682 3964 -672
rect 4031 -643 4046 -628
tri 3656 -707 3668 -695 ne
rect 3668 -700 3678 -695
tri 3678 -700 3683 -695 sw
rect 3567 -1046 3582 -818
rect 3668 -808 3683 -700
rect 3722 -742 3750 -686
tri 3842 -704 3860 -686 ne
rect 3860 -706 3882 -686
tri 3882 -706 3902 -686 sw
tri 3918 -700 3936 -682 ne
rect 3741 -776 3750 -742
rect 3784 -715 3826 -714
rect 3784 -749 3789 -715
rect 3819 -749 3826 -715
rect 3784 -758 3826 -749
rect 3860 -715 3902 -706
rect 3860 -749 3867 -715
rect 3897 -749 3902 -715
rect 3860 -754 3902 -749
rect 3936 -742 3964 -682
tri 4009 -695 4031 -673 se
rect 4031 -680 4046 -672
tri 4031 -695 4046 -680 nw
tri 4003 -701 4009 -695 se
rect 4009 -701 4018 -695
rect 3722 -786 3750 -776
tri 3750 -786 3774 -762 sw
rect 3668 -856 3684 -808
rect 3722 -818 3764 -786
tri 3781 -794 3782 -793 sw
rect 3781 -818 3782 -794
tri 3784 -795 3821 -758 ne
rect 3821 -786 3826 -758
tri 3826 -786 3852 -760 sw
rect 3936 -776 3945 -742
rect 3936 -786 3964 -776
rect 3821 -795 3905 -786
tri 3821 -814 3840 -795 ne
rect 3840 -814 3905 -795
rect 3722 -840 3782 -818
rect 3904 -818 3905 -814
rect 3922 -818 3964 -786
rect 3904 -840 3964 -818
rect 3810 -856 3827 -842
rect 3859 -856 3876 -842
tri 3647 -892 3669 -870 se
rect 3669 -877 3684 -856
tri 3669 -892 3684 -877 nw
rect 4003 -877 4018 -701
tri 4018 -708 4031 -695 nw
rect 4104 -776 4119 -548
tri 3641 -898 3647 -892 se
rect 3647 -898 3656 -892
rect 3641 -914 3656 -898
tri 3656 -905 3669 -892 nw
rect 3810 -900 3827 -886
rect 3859 -900 3876 -886
tri 4003 -892 4018 -877 ne
tri 4018 -892 4040 -870 sw
rect 3641 -950 3656 -942
rect 3722 -914 3782 -900
rect 3737 -924 3782 -914
rect 3737 -942 3765 -924
tri 3641 -965 3656 -950 ne
tri 3656 -965 3678 -943 sw
rect 3722 -952 3765 -942
rect 3780 -928 3782 -924
rect 3904 -914 3964 -900
tri 4018 -905 4031 -892 ne
rect 4031 -898 4040 -892
tri 4040 -898 4046 -892 sw
rect 3904 -924 3949 -914
rect 3780 -952 3854 -928
rect 3722 -956 3854 -952
tri 3854 -956 3882 -928 sw
rect 3904 -938 3906 -924
tri 3904 -940 3906 -938 ne
rect 3918 -942 3949 -924
rect 3918 -952 3964 -942
rect 4031 -913 4046 -898
tri 3656 -977 3668 -965 ne
rect 3668 -970 3678 -965
tri 3678 -970 3683 -965 sw
rect 3567 -1316 3582 -1088
rect 3668 -1126 3683 -970
rect 3722 -1012 3750 -956
tri 3842 -974 3860 -956 ne
rect 3860 -976 3882 -956
tri 3882 -976 3902 -956 sw
tri 3918 -970 3936 -952 ne
rect 3741 -1046 3750 -1012
rect 3784 -985 3826 -984
rect 3784 -1019 3789 -985
rect 3819 -1019 3826 -985
rect 3784 -1028 3826 -1019
rect 3860 -985 3902 -976
rect 3860 -1019 3867 -985
rect 3897 -1019 3902 -985
rect 3860 -1024 3902 -1019
rect 3936 -1012 3964 -952
tri 4009 -965 4031 -943 se
rect 4031 -950 4046 -942
tri 4031 -965 4046 -950 nw
tri 4003 -971 4009 -965 se
rect 4009 -971 4018 -965
rect 3722 -1056 3750 -1046
tri 3750 -1056 3774 -1032 sw
rect 3722 -1088 3764 -1056
tri 3781 -1064 3782 -1063 sw
rect 3781 -1088 3782 -1064
tri 3784 -1065 3821 -1028 ne
rect 3821 -1056 3826 -1028
tri 3826 -1056 3852 -1030 sw
rect 3936 -1046 3945 -1012
rect 3936 -1056 3964 -1046
rect 3821 -1065 3905 -1056
tri 3821 -1084 3840 -1065 ne
rect 3840 -1084 3905 -1065
rect 3722 -1110 3782 -1088
rect 3904 -1088 3905 -1084
rect 3922 -1088 3964 -1056
rect 3904 -1110 3964 -1088
rect 3810 -1126 3827 -1112
rect 3859 -1126 3876 -1112
tri 3647 -1162 3669 -1140 se
rect 3669 -1147 3684 -1126
tri 3669 -1162 3684 -1147 nw
rect 4003 -1147 4018 -971
tri 4018 -978 4031 -965 nw
rect 4104 -1046 4119 -818
tri 3641 -1168 3647 -1162 se
rect 3647 -1168 3656 -1162
rect 3641 -1184 3656 -1168
tri 3656 -1175 3669 -1162 nw
rect 3810 -1170 3827 -1156
rect 3859 -1170 3876 -1156
tri 4003 -1162 4018 -1147 ne
tri 4018 -1162 4040 -1140 sw
rect 3641 -1220 3656 -1212
rect 3722 -1184 3782 -1170
rect 3737 -1194 3782 -1184
rect 3737 -1212 3765 -1194
tri 3641 -1235 3656 -1220 ne
tri 3656 -1235 3678 -1213 sw
rect 3722 -1222 3765 -1212
rect 3780 -1198 3782 -1194
rect 3904 -1184 3964 -1170
tri 4018 -1175 4031 -1162 ne
rect 4031 -1168 4040 -1162
tri 4040 -1168 4046 -1162 sw
rect 3904 -1194 3949 -1184
rect 3780 -1222 3854 -1198
rect 3722 -1226 3854 -1222
tri 3854 -1226 3882 -1198 sw
rect 3904 -1208 3906 -1194
tri 3904 -1210 3906 -1208 ne
rect 3918 -1212 3949 -1194
rect 3918 -1222 3964 -1212
rect 4031 -1183 4046 -1168
tri 3656 -1247 3668 -1235 ne
rect 3668 -1240 3678 -1235
tri 3678 -1240 3683 -1235 sw
rect 3567 -1586 3582 -1358
rect 3668 -1348 3683 -1240
rect 3722 -1282 3750 -1226
tri 3842 -1244 3860 -1226 ne
rect 3860 -1246 3882 -1226
tri 3882 -1246 3902 -1226 sw
tri 3918 -1240 3936 -1222 ne
rect 3741 -1316 3750 -1282
rect 3784 -1255 3826 -1254
rect 3784 -1289 3789 -1255
rect 3819 -1289 3826 -1255
rect 3784 -1298 3826 -1289
rect 3860 -1255 3902 -1246
rect 3860 -1289 3867 -1255
rect 3897 -1289 3902 -1255
rect 3860 -1294 3902 -1289
rect 3936 -1282 3964 -1222
tri 4009 -1235 4031 -1213 se
rect 4031 -1220 4046 -1212
tri 4031 -1235 4046 -1220 nw
tri 4003 -1241 4009 -1235 se
rect 4009 -1241 4018 -1235
rect 3722 -1326 3750 -1316
tri 3750 -1326 3774 -1302 sw
rect 3668 -1396 3684 -1348
rect 3722 -1358 3764 -1326
tri 3781 -1334 3782 -1333 sw
rect 3781 -1358 3782 -1334
tri 3784 -1335 3821 -1298 ne
rect 3821 -1326 3826 -1298
tri 3826 -1326 3852 -1300 sw
rect 3936 -1316 3945 -1282
rect 3936 -1326 3964 -1316
rect 3821 -1335 3905 -1326
tri 3821 -1354 3840 -1335 ne
rect 3840 -1354 3905 -1335
rect 3722 -1380 3782 -1358
rect 3904 -1358 3905 -1354
rect 3922 -1358 3964 -1326
rect 3904 -1380 3964 -1358
rect 3810 -1396 3827 -1382
rect 3859 -1396 3876 -1382
tri 3647 -1432 3669 -1410 se
rect 3669 -1417 3684 -1396
tri 3669 -1432 3684 -1417 nw
rect 4003 -1417 4018 -1241
tri 4018 -1248 4031 -1235 nw
rect 4104 -1316 4119 -1088
tri 3641 -1438 3647 -1432 se
rect 3647 -1438 3656 -1432
rect 3641 -1454 3656 -1438
tri 3656 -1445 3669 -1432 nw
rect 3810 -1440 3827 -1426
rect 3859 -1440 3876 -1426
tri 4003 -1432 4018 -1417 ne
tri 4018 -1432 4040 -1410 sw
rect 3641 -1490 3656 -1482
rect 3722 -1454 3782 -1440
rect 3737 -1464 3782 -1454
rect 3737 -1482 3765 -1464
tri 3641 -1505 3656 -1490 ne
tri 3656 -1505 3678 -1483 sw
rect 3722 -1492 3765 -1482
rect 3780 -1468 3782 -1464
rect 3904 -1454 3964 -1440
tri 4018 -1445 4031 -1432 ne
rect 4031 -1438 4040 -1432
tri 4040 -1438 4046 -1432 sw
rect 3904 -1464 3949 -1454
rect 3780 -1492 3854 -1468
rect 3722 -1496 3854 -1492
tri 3854 -1496 3882 -1468 sw
rect 3904 -1478 3906 -1464
tri 3904 -1480 3906 -1478 ne
rect 3918 -1482 3949 -1464
rect 3918 -1492 3964 -1482
rect 4031 -1453 4046 -1438
tri 3656 -1517 3668 -1505 ne
rect 3668 -1510 3678 -1505
tri 3678 -1510 3683 -1505 sw
rect 3567 -1856 3582 -1628
rect 3668 -1666 3683 -1510
rect 3722 -1552 3750 -1496
tri 3842 -1514 3860 -1496 ne
rect 3860 -1516 3882 -1496
tri 3882 -1516 3902 -1496 sw
tri 3918 -1510 3936 -1492 ne
rect 3741 -1586 3750 -1552
rect 3784 -1525 3826 -1524
rect 3784 -1559 3789 -1525
rect 3819 -1559 3826 -1525
rect 3784 -1568 3826 -1559
rect 3860 -1525 3902 -1516
rect 3860 -1559 3867 -1525
rect 3897 -1559 3902 -1525
rect 3860 -1564 3902 -1559
rect 3936 -1552 3964 -1492
tri 4009 -1505 4031 -1483 se
rect 4031 -1490 4046 -1482
tri 4031 -1505 4046 -1490 nw
tri 4003 -1511 4009 -1505 se
rect 4009 -1511 4018 -1505
rect 3722 -1596 3750 -1586
tri 3750 -1596 3774 -1572 sw
rect 3722 -1628 3764 -1596
tri 3781 -1604 3782 -1603 sw
rect 3781 -1628 3782 -1604
tri 3784 -1605 3821 -1568 ne
rect 3821 -1596 3826 -1568
tri 3826 -1596 3852 -1570 sw
rect 3936 -1586 3945 -1552
rect 3936 -1596 3964 -1586
rect 3821 -1605 3905 -1596
tri 3821 -1624 3840 -1605 ne
rect 3840 -1624 3905 -1605
rect 3722 -1650 3782 -1628
rect 3904 -1628 3905 -1624
rect 3922 -1628 3964 -1596
rect 3904 -1650 3964 -1628
rect 3810 -1666 3827 -1652
rect 3859 -1666 3876 -1652
tri 3647 -1702 3669 -1680 se
rect 3669 -1687 3684 -1666
tri 3669 -1702 3684 -1687 nw
rect 4003 -1687 4018 -1511
tri 4018 -1518 4031 -1505 nw
rect 4104 -1586 4119 -1358
tri 3641 -1708 3647 -1702 se
rect 3647 -1708 3656 -1702
rect 3641 -1724 3656 -1708
tri 3656 -1715 3669 -1702 nw
rect 3810 -1710 3827 -1696
rect 3859 -1710 3876 -1696
tri 4003 -1702 4018 -1687 ne
tri 4018 -1702 4040 -1680 sw
rect 3641 -1760 3656 -1752
rect 3722 -1724 3782 -1710
rect 3737 -1734 3782 -1724
rect 3737 -1752 3765 -1734
tri 3641 -1775 3656 -1760 ne
tri 3656 -1775 3678 -1753 sw
rect 3722 -1762 3765 -1752
rect 3780 -1738 3782 -1734
rect 3904 -1724 3964 -1710
tri 4018 -1715 4031 -1702 ne
rect 4031 -1708 4040 -1702
tri 4040 -1708 4046 -1702 sw
rect 3904 -1734 3949 -1724
rect 3780 -1762 3854 -1738
rect 3722 -1766 3854 -1762
tri 3854 -1766 3882 -1738 sw
rect 3904 -1748 3906 -1734
tri 3904 -1750 3906 -1748 ne
rect 3918 -1752 3949 -1734
rect 3918 -1762 3964 -1752
rect 4031 -1723 4046 -1708
tri 3656 -1787 3668 -1775 ne
rect 3668 -1780 3678 -1775
tri 3678 -1780 3683 -1775 sw
rect 3567 -2126 3582 -1898
rect 3668 -1888 3683 -1780
rect 3722 -1822 3750 -1766
tri 3842 -1784 3860 -1766 ne
rect 3860 -1786 3882 -1766
tri 3882 -1786 3902 -1766 sw
tri 3918 -1780 3936 -1762 ne
rect 3741 -1856 3750 -1822
rect 3784 -1795 3826 -1794
rect 3784 -1829 3789 -1795
rect 3819 -1829 3826 -1795
rect 3784 -1838 3826 -1829
rect 3860 -1795 3902 -1786
rect 3860 -1829 3867 -1795
rect 3897 -1829 3902 -1795
rect 3860 -1834 3902 -1829
rect 3936 -1822 3964 -1762
tri 4009 -1775 4031 -1753 se
rect 4031 -1760 4046 -1752
tri 4031 -1775 4046 -1760 nw
tri 4003 -1781 4009 -1775 se
rect 4009 -1781 4018 -1775
rect 3722 -1866 3750 -1856
tri 3750 -1866 3774 -1842 sw
rect 3668 -1936 3684 -1888
rect 3722 -1898 3764 -1866
tri 3781 -1874 3782 -1873 sw
rect 3781 -1898 3782 -1874
tri 3784 -1875 3821 -1838 ne
rect 3821 -1866 3826 -1838
tri 3826 -1866 3852 -1840 sw
rect 3936 -1856 3945 -1822
rect 3936 -1866 3964 -1856
rect 3821 -1875 3905 -1866
tri 3821 -1894 3840 -1875 ne
rect 3840 -1894 3905 -1875
rect 3722 -1920 3782 -1898
rect 3904 -1898 3905 -1894
rect 3922 -1898 3964 -1866
rect 3904 -1920 3964 -1898
rect 3810 -1936 3827 -1922
rect 3859 -1936 3876 -1922
tri 3647 -1972 3669 -1950 se
rect 3669 -1957 3684 -1936
tri 3669 -1972 3684 -1957 nw
rect 4003 -1957 4018 -1781
tri 4018 -1788 4031 -1775 nw
rect 4104 -1856 4119 -1628
tri 3641 -1978 3647 -1972 se
rect 3647 -1978 3656 -1972
rect 3641 -1994 3656 -1978
tri 3656 -1985 3669 -1972 nw
rect 3810 -1980 3827 -1966
rect 3859 -1980 3876 -1966
tri 4003 -1972 4018 -1957 ne
tri 4018 -1972 4040 -1950 sw
rect 3641 -2030 3656 -2022
rect 3722 -1994 3782 -1980
rect 3737 -2004 3782 -1994
rect 3737 -2022 3765 -2004
tri 3641 -2045 3656 -2030 ne
tri 3656 -2045 3678 -2023 sw
rect 3722 -2032 3765 -2022
rect 3780 -2008 3782 -2004
rect 3904 -1994 3964 -1980
tri 4018 -1985 4031 -1972 ne
rect 4031 -1978 4040 -1972
tri 4040 -1978 4046 -1972 sw
rect 3904 -2004 3949 -1994
rect 3780 -2032 3854 -2008
rect 3722 -2036 3854 -2032
tri 3854 -2036 3882 -2008 sw
rect 3904 -2018 3906 -2004
tri 3904 -2020 3906 -2018 ne
rect 3918 -2022 3949 -2004
rect 3918 -2032 3964 -2022
rect 4031 -1993 4046 -1978
tri 3656 -2057 3668 -2045 ne
rect 3668 -2050 3678 -2045
tri 3678 -2050 3683 -2045 sw
rect 3567 -2396 3582 -2168
rect 3668 -2206 3683 -2050
rect 3722 -2092 3750 -2036
tri 3842 -2054 3860 -2036 ne
rect 3860 -2056 3882 -2036
tri 3882 -2056 3902 -2036 sw
tri 3918 -2050 3936 -2032 ne
rect 3741 -2126 3750 -2092
rect 3784 -2065 3826 -2064
rect 3784 -2099 3789 -2065
rect 3819 -2099 3826 -2065
rect 3784 -2108 3826 -2099
rect 3860 -2065 3902 -2056
rect 3860 -2099 3867 -2065
rect 3897 -2099 3902 -2065
rect 3860 -2104 3902 -2099
rect 3936 -2092 3964 -2032
tri 4009 -2045 4031 -2023 se
rect 4031 -2030 4046 -2022
tri 4031 -2045 4046 -2030 nw
tri 4003 -2051 4009 -2045 se
rect 4009 -2051 4018 -2045
rect 3722 -2136 3750 -2126
tri 3750 -2136 3774 -2112 sw
rect 3722 -2168 3764 -2136
tri 3781 -2144 3782 -2143 sw
rect 3781 -2168 3782 -2144
tri 3784 -2145 3821 -2108 ne
rect 3821 -2136 3826 -2108
tri 3826 -2136 3852 -2110 sw
rect 3936 -2126 3945 -2092
rect 3936 -2136 3964 -2126
rect 3821 -2145 3905 -2136
tri 3821 -2164 3840 -2145 ne
rect 3840 -2164 3905 -2145
rect 3722 -2190 3782 -2168
rect 3904 -2168 3905 -2164
rect 3922 -2168 3964 -2136
rect 3904 -2190 3964 -2168
rect 3810 -2206 3827 -2192
rect 3859 -2206 3876 -2192
tri 3647 -2242 3669 -2220 se
rect 3669 -2227 3684 -2206
tri 3669 -2242 3684 -2227 nw
rect 4003 -2227 4018 -2051
tri 4018 -2058 4031 -2045 nw
rect 4104 -2126 4119 -1898
tri 3641 -2248 3647 -2242 se
rect 3647 -2248 3656 -2242
rect 3641 -2264 3656 -2248
tri 3656 -2255 3669 -2242 nw
rect 3810 -2250 3827 -2236
rect 3859 -2250 3876 -2236
tri 4003 -2242 4018 -2227 ne
tri 4018 -2242 4040 -2220 sw
rect 3641 -2300 3656 -2292
rect 3722 -2264 3782 -2250
rect 3737 -2274 3782 -2264
rect 3737 -2292 3765 -2274
tri 3641 -2315 3656 -2300 ne
tri 3656 -2315 3678 -2293 sw
rect 3722 -2302 3765 -2292
rect 3780 -2278 3782 -2274
rect 3904 -2264 3964 -2250
tri 4018 -2255 4031 -2242 ne
rect 4031 -2248 4040 -2242
tri 4040 -2248 4046 -2242 sw
rect 3904 -2274 3949 -2264
rect 3780 -2302 3854 -2278
rect 3722 -2306 3854 -2302
tri 3854 -2306 3882 -2278 sw
rect 3904 -2288 3906 -2274
tri 3904 -2290 3906 -2288 ne
rect 3918 -2292 3949 -2274
rect 3918 -2302 3964 -2292
rect 4031 -2263 4046 -2248
tri 3656 -2327 3668 -2315 ne
rect 3668 -2320 3678 -2315
tri 3678 -2320 3683 -2315 sw
rect 3567 -2524 3582 -2438
rect 3668 -2476 3683 -2320
rect 3722 -2362 3750 -2306
tri 3842 -2324 3860 -2306 ne
rect 3860 -2326 3882 -2306
tri 3882 -2326 3902 -2306 sw
tri 3918 -2320 3936 -2302 ne
rect 3741 -2396 3750 -2362
rect 3784 -2335 3826 -2334
rect 3784 -2369 3789 -2335
rect 3819 -2369 3826 -2335
rect 3784 -2378 3826 -2369
rect 3860 -2335 3902 -2326
rect 3860 -2369 3867 -2335
rect 3897 -2369 3902 -2335
rect 3860 -2374 3902 -2369
rect 3936 -2362 3964 -2302
tri 4009 -2315 4031 -2293 se
rect 4031 -2300 4046 -2292
tri 4031 -2315 4046 -2300 nw
tri 4003 -2321 4009 -2315 se
rect 4009 -2321 4018 -2315
rect 3722 -2406 3750 -2396
tri 3750 -2406 3774 -2382 sw
rect 3722 -2438 3764 -2406
tri 3781 -2414 3782 -2413 sw
rect 3781 -2438 3782 -2414
tri 3784 -2415 3821 -2378 ne
rect 3821 -2406 3826 -2378
tri 3826 -2406 3852 -2380 sw
rect 3936 -2396 3945 -2362
rect 3936 -2406 3964 -2396
rect 3821 -2415 3905 -2406
tri 3821 -2434 3840 -2415 ne
rect 3840 -2434 3905 -2415
rect 3722 -2460 3782 -2438
rect 3904 -2438 3905 -2434
rect 3922 -2438 3964 -2406
rect 3904 -2460 3964 -2438
rect 3810 -2476 3827 -2462
rect 3859 -2476 3876 -2462
rect 4003 -2476 4018 -2321
tri 4018 -2328 4031 -2315 nw
rect 4104 -2396 4119 -2168
rect 4104 -2524 4119 -2438
rect 4147 1654 4162 1844
tri 4227 1808 4249 1830 se
rect 4249 1823 4264 1892
tri 4249 1808 4264 1823 nw
rect 4583 1823 4598 1892
tri 4221 1802 4227 1808 se
rect 4227 1802 4236 1808
rect 4221 1786 4236 1802
tri 4236 1795 4249 1808 nw
rect 4390 1800 4407 1814
rect 4439 1800 4456 1814
tri 4583 1808 4598 1823 ne
tri 4598 1808 4620 1830 sw
rect 4221 1750 4236 1758
rect 4302 1786 4362 1800
rect 4317 1776 4362 1786
rect 4317 1758 4345 1776
tri 4221 1735 4236 1750 ne
tri 4236 1735 4258 1757 sw
rect 4302 1748 4345 1758
rect 4360 1772 4362 1776
rect 4484 1786 4544 1800
tri 4598 1795 4611 1808 ne
rect 4611 1802 4620 1808
tri 4620 1802 4626 1808 sw
rect 4484 1776 4529 1786
rect 4360 1748 4434 1772
rect 4302 1744 4434 1748
tri 4434 1744 4462 1772 sw
rect 4484 1762 4486 1776
tri 4484 1760 4486 1762 ne
rect 4498 1758 4529 1776
rect 4498 1748 4544 1758
rect 4611 1787 4626 1802
tri 4236 1723 4248 1735 ne
rect 4248 1730 4258 1735
tri 4258 1730 4263 1735 sw
rect 4147 1384 4162 1612
rect 4248 1574 4263 1730
rect 4302 1688 4330 1744
tri 4422 1726 4440 1744 ne
rect 4440 1724 4462 1744
tri 4462 1724 4482 1744 sw
tri 4498 1730 4516 1748 ne
rect 4321 1654 4330 1688
rect 4364 1715 4406 1716
rect 4364 1681 4369 1715
rect 4399 1681 4406 1715
rect 4364 1672 4406 1681
rect 4440 1715 4482 1724
rect 4440 1681 4447 1715
rect 4477 1681 4482 1715
rect 4440 1676 4482 1681
rect 4516 1688 4544 1748
tri 4589 1735 4611 1757 se
rect 4611 1750 4626 1758
tri 4611 1735 4626 1750 nw
tri 4583 1729 4589 1735 se
rect 4589 1729 4598 1735
rect 4302 1644 4330 1654
tri 4330 1644 4354 1668 sw
rect 4302 1612 4344 1644
tri 4361 1636 4362 1637 sw
rect 4361 1612 4362 1636
tri 4364 1635 4401 1672 ne
rect 4401 1644 4406 1672
tri 4406 1644 4432 1670 sw
rect 4516 1654 4525 1688
rect 4516 1644 4544 1654
rect 4401 1635 4485 1644
tri 4401 1616 4420 1635 ne
rect 4420 1616 4485 1635
rect 4302 1590 4362 1612
rect 4484 1612 4485 1616
rect 4502 1612 4544 1644
rect 4484 1590 4544 1612
rect 4390 1574 4407 1588
rect 4439 1574 4456 1588
tri 4227 1538 4249 1560 se
rect 4249 1553 4264 1574
tri 4249 1538 4264 1553 nw
rect 4583 1553 4598 1729
tri 4598 1722 4611 1735 nw
rect 4684 1654 4699 1844
tri 4221 1532 4227 1538 se
rect 4227 1532 4236 1538
rect 4221 1516 4236 1532
tri 4236 1525 4249 1538 nw
rect 4390 1530 4407 1544
rect 4439 1530 4456 1544
tri 4583 1538 4598 1553 ne
tri 4598 1538 4620 1560 sw
rect 4221 1480 4236 1488
rect 4302 1516 4362 1530
rect 4317 1506 4362 1516
rect 4317 1488 4345 1506
tri 4221 1465 4236 1480 ne
tri 4236 1465 4258 1487 sw
rect 4302 1478 4345 1488
rect 4360 1502 4362 1506
rect 4484 1516 4544 1530
tri 4598 1525 4611 1538 ne
rect 4611 1532 4620 1538
tri 4620 1532 4626 1538 sw
rect 4484 1506 4529 1516
rect 4360 1478 4434 1502
rect 4302 1474 4434 1478
tri 4434 1474 4462 1502 sw
rect 4484 1492 4486 1506
tri 4484 1490 4486 1492 ne
rect 4498 1488 4529 1506
rect 4498 1478 4544 1488
rect 4611 1517 4626 1532
tri 4236 1453 4248 1465 ne
rect 4248 1460 4258 1465
tri 4258 1460 4263 1465 sw
rect 4147 1114 4162 1342
rect 4248 1352 4263 1460
rect 4302 1418 4330 1474
tri 4422 1456 4440 1474 ne
rect 4440 1454 4462 1474
tri 4462 1454 4482 1474 sw
tri 4498 1460 4516 1478 ne
rect 4321 1384 4330 1418
rect 4364 1445 4406 1446
rect 4364 1411 4369 1445
rect 4399 1411 4406 1445
rect 4364 1402 4406 1411
rect 4440 1445 4482 1454
rect 4440 1411 4447 1445
rect 4477 1411 4482 1445
rect 4440 1406 4482 1411
rect 4516 1418 4544 1478
tri 4589 1465 4611 1487 se
rect 4611 1480 4626 1488
tri 4611 1465 4626 1480 nw
tri 4583 1459 4589 1465 se
rect 4589 1459 4598 1465
rect 4302 1374 4330 1384
tri 4330 1374 4354 1398 sw
rect 4248 1304 4264 1352
rect 4302 1342 4344 1374
tri 4361 1366 4362 1367 sw
rect 4361 1342 4362 1366
tri 4364 1365 4401 1402 ne
rect 4401 1374 4406 1402
tri 4406 1374 4432 1400 sw
rect 4516 1384 4525 1418
rect 4516 1374 4544 1384
rect 4401 1365 4485 1374
tri 4401 1346 4420 1365 ne
rect 4420 1346 4485 1365
rect 4302 1320 4362 1342
rect 4484 1342 4485 1346
rect 4502 1342 4544 1374
rect 4484 1320 4544 1342
rect 4390 1304 4407 1318
rect 4439 1304 4456 1318
tri 4227 1268 4249 1290 se
rect 4249 1283 4264 1304
tri 4249 1268 4264 1283 nw
rect 4583 1283 4598 1459
tri 4598 1452 4611 1465 nw
rect 4684 1384 4699 1612
tri 4221 1262 4227 1268 se
rect 4227 1262 4236 1268
rect 4221 1246 4236 1262
tri 4236 1255 4249 1268 nw
rect 4390 1260 4407 1274
rect 4439 1260 4456 1274
tri 4583 1268 4598 1283 ne
tri 4598 1268 4620 1290 sw
rect 4221 1210 4236 1218
rect 4302 1246 4362 1260
rect 4317 1236 4362 1246
rect 4317 1218 4345 1236
tri 4221 1195 4236 1210 ne
tri 4236 1195 4258 1217 sw
rect 4302 1208 4345 1218
rect 4360 1232 4362 1236
rect 4484 1246 4544 1260
tri 4598 1255 4611 1268 ne
rect 4611 1262 4620 1268
tri 4620 1262 4626 1268 sw
rect 4484 1236 4529 1246
rect 4360 1208 4434 1232
rect 4302 1204 4434 1208
tri 4434 1204 4462 1232 sw
rect 4484 1222 4486 1236
tri 4484 1220 4486 1222 ne
rect 4498 1218 4529 1236
rect 4498 1208 4544 1218
rect 4611 1247 4626 1262
tri 4236 1183 4248 1195 ne
rect 4248 1190 4258 1195
tri 4258 1190 4263 1195 sw
rect 4147 844 4162 1072
rect 4248 1034 4263 1190
rect 4302 1148 4330 1204
tri 4422 1186 4440 1204 ne
rect 4440 1184 4462 1204
tri 4462 1184 4482 1204 sw
tri 4498 1190 4516 1208 ne
rect 4321 1114 4330 1148
rect 4364 1175 4406 1176
rect 4364 1141 4369 1175
rect 4399 1141 4406 1175
rect 4364 1132 4406 1141
rect 4440 1175 4482 1184
rect 4440 1141 4447 1175
rect 4477 1141 4482 1175
rect 4440 1136 4482 1141
rect 4516 1148 4544 1208
tri 4589 1195 4611 1217 se
rect 4611 1210 4626 1218
tri 4611 1195 4626 1210 nw
tri 4583 1189 4589 1195 se
rect 4589 1189 4598 1195
rect 4302 1104 4330 1114
tri 4330 1104 4354 1128 sw
rect 4302 1072 4344 1104
tri 4361 1096 4362 1097 sw
rect 4361 1072 4362 1096
tri 4364 1095 4401 1132 ne
rect 4401 1104 4406 1132
tri 4406 1104 4432 1130 sw
rect 4516 1114 4525 1148
rect 4516 1104 4544 1114
rect 4401 1095 4485 1104
tri 4401 1076 4420 1095 ne
rect 4420 1076 4485 1095
rect 4302 1050 4362 1072
rect 4484 1072 4485 1076
rect 4502 1072 4544 1104
rect 4484 1050 4544 1072
rect 4390 1034 4407 1048
rect 4439 1034 4456 1048
tri 4227 998 4249 1020 se
rect 4249 1013 4264 1034
tri 4249 998 4264 1013 nw
rect 4583 1013 4598 1189
tri 4598 1182 4611 1195 nw
rect 4684 1114 4699 1342
tri 4221 992 4227 998 se
rect 4227 992 4236 998
rect 4221 976 4236 992
tri 4236 985 4249 998 nw
rect 4390 990 4407 1004
rect 4439 990 4456 1004
tri 4583 998 4598 1013 ne
tri 4598 998 4620 1020 sw
rect 4221 940 4236 948
rect 4302 976 4362 990
rect 4317 966 4362 976
rect 4317 948 4345 966
tri 4221 925 4236 940 ne
tri 4236 925 4258 947 sw
rect 4302 938 4345 948
rect 4360 962 4362 966
rect 4484 976 4544 990
tri 4598 985 4611 998 ne
rect 4611 992 4620 998
tri 4620 992 4626 998 sw
rect 4484 966 4529 976
rect 4360 938 4434 962
rect 4302 934 4434 938
tri 4434 934 4462 962 sw
rect 4484 952 4486 966
tri 4484 950 4486 952 ne
rect 4498 948 4529 966
rect 4498 938 4544 948
rect 4611 977 4626 992
tri 4236 913 4248 925 ne
rect 4248 920 4258 925
tri 4258 920 4263 925 sw
rect 4147 574 4162 802
rect 4248 812 4263 920
rect 4302 878 4330 934
tri 4422 916 4440 934 ne
rect 4440 914 4462 934
tri 4462 914 4482 934 sw
tri 4498 920 4516 938 ne
rect 4321 844 4330 878
rect 4364 905 4406 906
rect 4364 871 4369 905
rect 4399 871 4406 905
rect 4364 862 4406 871
rect 4440 905 4482 914
rect 4440 871 4447 905
rect 4477 871 4482 905
rect 4440 866 4482 871
rect 4516 878 4544 938
tri 4589 925 4611 947 se
rect 4611 940 4626 948
tri 4611 925 4626 940 nw
tri 4583 919 4589 925 se
rect 4589 919 4598 925
rect 4302 834 4330 844
tri 4330 834 4354 858 sw
rect 4248 764 4264 812
rect 4302 802 4344 834
tri 4361 826 4362 827 sw
rect 4361 802 4362 826
tri 4364 825 4401 862 ne
rect 4401 834 4406 862
tri 4406 834 4432 860 sw
rect 4516 844 4525 878
rect 4516 834 4544 844
rect 4401 825 4485 834
tri 4401 806 4420 825 ne
rect 4420 806 4485 825
rect 4302 780 4362 802
rect 4484 802 4485 806
rect 4502 802 4544 834
rect 4484 780 4544 802
rect 4390 764 4407 778
rect 4439 764 4456 778
tri 4227 728 4249 750 se
rect 4249 743 4264 764
tri 4249 728 4264 743 nw
rect 4583 743 4598 919
tri 4598 912 4611 925 nw
rect 4684 844 4699 1072
tri 4221 722 4227 728 se
rect 4227 722 4236 728
rect 4221 706 4236 722
tri 4236 715 4249 728 nw
rect 4390 720 4407 734
rect 4439 720 4456 734
tri 4583 728 4598 743 ne
tri 4598 728 4620 750 sw
rect 4221 670 4236 678
rect 4302 706 4362 720
rect 4317 696 4362 706
rect 4317 678 4345 696
tri 4221 655 4236 670 ne
tri 4236 655 4258 677 sw
rect 4302 668 4345 678
rect 4360 692 4362 696
rect 4484 706 4544 720
tri 4598 715 4611 728 ne
rect 4611 722 4620 728
tri 4620 722 4626 728 sw
rect 4484 696 4529 706
rect 4360 668 4434 692
rect 4302 664 4434 668
tri 4434 664 4462 692 sw
rect 4484 682 4486 696
tri 4484 680 4486 682 ne
rect 4498 678 4529 696
rect 4498 668 4544 678
rect 4611 707 4626 722
tri 4236 643 4248 655 ne
rect 4248 650 4258 655
tri 4258 650 4263 655 sw
rect 4147 304 4162 532
rect 4248 494 4263 650
rect 4302 608 4330 664
tri 4422 646 4440 664 ne
rect 4440 644 4462 664
tri 4462 644 4482 664 sw
tri 4498 650 4516 668 ne
rect 4321 574 4330 608
rect 4364 635 4406 636
rect 4364 601 4369 635
rect 4399 601 4406 635
rect 4364 592 4406 601
rect 4440 635 4482 644
rect 4440 601 4447 635
rect 4477 601 4482 635
rect 4440 596 4482 601
rect 4516 608 4544 668
tri 4589 655 4611 677 se
rect 4611 670 4626 678
tri 4611 655 4626 670 nw
tri 4583 649 4589 655 se
rect 4589 649 4598 655
rect 4302 564 4330 574
tri 4330 564 4354 588 sw
rect 4302 532 4344 564
tri 4361 556 4362 557 sw
rect 4361 532 4362 556
tri 4364 555 4401 592 ne
rect 4401 564 4406 592
tri 4406 564 4432 590 sw
rect 4516 574 4525 608
rect 4516 564 4544 574
rect 4401 555 4485 564
tri 4401 536 4420 555 ne
rect 4420 536 4485 555
rect 4302 510 4362 532
rect 4484 532 4485 536
rect 4502 532 4544 564
rect 4484 510 4544 532
rect 4390 494 4407 508
rect 4439 494 4456 508
tri 4227 458 4249 480 se
rect 4249 473 4264 494
tri 4249 458 4264 473 nw
rect 4583 473 4598 649
tri 4598 642 4611 655 nw
rect 4684 574 4699 802
tri 4221 452 4227 458 se
rect 4227 452 4236 458
rect 4221 436 4236 452
tri 4236 445 4249 458 nw
rect 4390 450 4407 464
rect 4439 450 4456 464
tri 4583 458 4598 473 ne
tri 4598 458 4620 480 sw
rect 4221 400 4236 408
rect 4302 436 4362 450
rect 4317 426 4362 436
rect 4317 408 4345 426
tri 4221 385 4236 400 ne
tri 4236 385 4258 407 sw
rect 4302 398 4345 408
rect 4360 422 4362 426
rect 4484 436 4544 450
tri 4598 445 4611 458 ne
rect 4611 452 4620 458
tri 4620 452 4626 458 sw
rect 4484 426 4529 436
rect 4360 398 4434 422
rect 4302 394 4434 398
tri 4434 394 4462 422 sw
rect 4484 412 4486 426
tri 4484 410 4486 412 ne
rect 4498 408 4529 426
rect 4498 398 4544 408
rect 4611 437 4626 452
tri 4236 373 4248 385 ne
rect 4248 380 4258 385
tri 4258 380 4263 385 sw
rect 4147 34 4162 262
rect 4248 272 4263 380
rect 4302 338 4330 394
tri 4422 376 4440 394 ne
rect 4440 374 4462 394
tri 4462 374 4482 394 sw
tri 4498 380 4516 398 ne
rect 4321 304 4330 338
rect 4364 365 4406 366
rect 4364 331 4369 365
rect 4399 331 4406 365
rect 4364 322 4406 331
rect 4440 365 4482 374
rect 4440 331 4447 365
rect 4477 331 4482 365
rect 4440 326 4482 331
rect 4516 338 4544 398
tri 4589 385 4611 407 se
rect 4611 400 4626 408
tri 4611 385 4626 400 nw
tri 4583 379 4589 385 se
rect 4589 379 4598 385
rect 4302 294 4330 304
tri 4330 294 4354 318 sw
rect 4248 224 4264 272
rect 4302 262 4344 294
tri 4361 286 4362 287 sw
rect 4361 262 4362 286
tri 4364 285 4401 322 ne
rect 4401 294 4406 322
tri 4406 294 4432 320 sw
rect 4516 304 4525 338
rect 4516 294 4544 304
rect 4401 285 4485 294
tri 4401 266 4420 285 ne
rect 4420 266 4485 285
rect 4302 240 4362 262
rect 4484 262 4485 266
rect 4502 262 4544 294
rect 4484 240 4544 262
rect 4390 224 4407 238
rect 4439 224 4456 238
tri 4227 188 4249 210 se
rect 4249 203 4264 224
tri 4249 188 4264 203 nw
rect 4583 203 4598 379
tri 4598 372 4611 385 nw
rect 4684 304 4699 532
tri 4221 182 4227 188 se
rect 4227 182 4236 188
rect 4221 166 4236 182
tri 4236 175 4249 188 nw
rect 4390 180 4407 194
rect 4439 180 4456 194
tri 4583 188 4598 203 ne
tri 4598 188 4620 210 sw
rect 4221 130 4236 138
rect 4302 166 4362 180
rect 4317 156 4362 166
rect 4317 138 4345 156
tri 4221 115 4236 130 ne
tri 4236 115 4258 137 sw
rect 4302 128 4345 138
rect 4360 152 4362 156
rect 4484 166 4544 180
tri 4598 175 4611 188 ne
rect 4611 182 4620 188
tri 4620 182 4626 188 sw
rect 4484 156 4529 166
rect 4360 128 4434 152
rect 4302 124 4434 128
tri 4434 124 4462 152 sw
rect 4484 142 4486 156
tri 4484 140 4486 142 ne
rect 4498 138 4529 156
rect 4498 128 4544 138
rect 4611 167 4626 182
tri 4236 103 4248 115 ne
rect 4248 110 4258 115
tri 4258 110 4263 115 sw
rect 4147 -236 4162 -8
rect 4248 -46 4263 110
rect 4302 68 4330 124
tri 4422 106 4440 124 ne
rect 4440 104 4462 124
tri 4462 104 4482 124 sw
tri 4498 110 4516 128 ne
rect 4321 34 4330 68
rect 4364 95 4406 96
rect 4364 61 4369 95
rect 4399 61 4406 95
rect 4364 52 4406 61
rect 4440 95 4482 104
rect 4440 61 4447 95
rect 4477 61 4482 95
rect 4440 56 4482 61
rect 4516 68 4544 128
tri 4589 115 4611 137 se
rect 4611 130 4626 138
tri 4611 115 4626 130 nw
tri 4583 109 4589 115 se
rect 4589 109 4598 115
rect 4302 24 4330 34
tri 4330 24 4354 48 sw
rect 4302 -8 4344 24
tri 4361 16 4362 17 sw
rect 4361 -8 4362 16
tri 4364 15 4401 52 ne
rect 4401 24 4406 52
tri 4406 24 4432 50 sw
rect 4516 34 4525 68
rect 4516 24 4544 34
rect 4401 15 4485 24
tri 4401 -4 4420 15 ne
rect 4420 -4 4485 15
rect 4302 -30 4362 -8
rect 4484 -8 4485 -4
rect 4502 -8 4544 24
rect 4484 -30 4544 -8
rect 4390 -46 4407 -32
rect 4439 -46 4456 -32
tri 4227 -82 4249 -60 se
rect 4249 -67 4264 -46
tri 4249 -82 4264 -67 nw
rect 4583 -67 4598 109
tri 4598 102 4611 115 nw
rect 4684 34 4699 262
tri 4221 -88 4227 -82 se
rect 4227 -88 4236 -82
rect 4221 -104 4236 -88
tri 4236 -95 4249 -82 nw
rect 4390 -90 4407 -76
rect 4439 -90 4456 -76
tri 4583 -82 4598 -67 ne
tri 4598 -82 4620 -60 sw
rect 4221 -140 4236 -132
rect 4302 -104 4362 -90
rect 4317 -114 4362 -104
rect 4317 -132 4345 -114
tri 4221 -155 4236 -140 ne
tri 4236 -155 4258 -133 sw
rect 4302 -142 4345 -132
rect 4360 -118 4362 -114
rect 4484 -104 4544 -90
tri 4598 -95 4611 -82 ne
rect 4611 -88 4620 -82
tri 4620 -88 4626 -82 sw
rect 4484 -114 4529 -104
rect 4360 -142 4434 -118
rect 4302 -146 4434 -142
tri 4434 -146 4462 -118 sw
rect 4484 -128 4486 -114
tri 4484 -130 4486 -128 ne
rect 4498 -132 4529 -114
rect 4498 -142 4544 -132
rect 4611 -103 4626 -88
tri 4236 -167 4248 -155 ne
rect 4248 -160 4258 -155
tri 4258 -160 4263 -155 sw
rect 4147 -506 4162 -278
rect 4248 -268 4263 -160
rect 4302 -202 4330 -146
tri 4422 -164 4440 -146 ne
rect 4440 -166 4462 -146
tri 4462 -166 4482 -146 sw
tri 4498 -160 4516 -142 ne
rect 4321 -236 4330 -202
rect 4364 -175 4406 -174
rect 4364 -209 4369 -175
rect 4399 -209 4406 -175
rect 4364 -218 4406 -209
rect 4440 -175 4482 -166
rect 4440 -209 4447 -175
rect 4477 -209 4482 -175
rect 4440 -214 4482 -209
rect 4516 -202 4544 -142
tri 4589 -155 4611 -133 se
rect 4611 -140 4626 -132
tri 4611 -155 4626 -140 nw
tri 4583 -161 4589 -155 se
rect 4589 -161 4598 -155
rect 4302 -246 4330 -236
tri 4330 -246 4354 -222 sw
rect 4248 -316 4264 -268
rect 4302 -278 4344 -246
tri 4361 -254 4362 -253 sw
rect 4361 -278 4362 -254
tri 4364 -255 4401 -218 ne
rect 4401 -246 4406 -218
tri 4406 -246 4432 -220 sw
rect 4516 -236 4525 -202
rect 4516 -246 4544 -236
rect 4401 -255 4485 -246
tri 4401 -274 4420 -255 ne
rect 4420 -274 4485 -255
rect 4302 -300 4362 -278
rect 4484 -278 4485 -274
rect 4502 -278 4544 -246
rect 4484 -300 4544 -278
rect 4390 -316 4407 -302
rect 4439 -316 4456 -302
tri 4227 -352 4249 -330 se
rect 4249 -337 4264 -316
tri 4249 -352 4264 -337 nw
rect 4583 -337 4598 -161
tri 4598 -168 4611 -155 nw
rect 4684 -236 4699 -8
tri 4221 -358 4227 -352 se
rect 4227 -358 4236 -352
rect 4221 -374 4236 -358
tri 4236 -365 4249 -352 nw
rect 4390 -360 4407 -346
rect 4439 -360 4456 -346
tri 4583 -352 4598 -337 ne
tri 4598 -352 4620 -330 sw
rect 4221 -410 4236 -402
rect 4302 -374 4362 -360
rect 4317 -384 4362 -374
rect 4317 -402 4345 -384
tri 4221 -425 4236 -410 ne
tri 4236 -425 4258 -403 sw
rect 4302 -412 4345 -402
rect 4360 -388 4362 -384
rect 4484 -374 4544 -360
tri 4598 -365 4611 -352 ne
rect 4611 -358 4620 -352
tri 4620 -358 4626 -352 sw
rect 4484 -384 4529 -374
rect 4360 -412 4434 -388
rect 4302 -416 4434 -412
tri 4434 -416 4462 -388 sw
rect 4484 -398 4486 -384
tri 4484 -400 4486 -398 ne
rect 4498 -402 4529 -384
rect 4498 -412 4544 -402
rect 4611 -373 4626 -358
tri 4236 -437 4248 -425 ne
rect 4248 -430 4258 -425
tri 4258 -430 4263 -425 sw
rect 4147 -776 4162 -548
rect 4248 -586 4263 -430
rect 4302 -472 4330 -416
tri 4422 -434 4440 -416 ne
rect 4440 -436 4462 -416
tri 4462 -436 4482 -416 sw
tri 4498 -430 4516 -412 ne
rect 4321 -506 4330 -472
rect 4364 -445 4406 -444
rect 4364 -479 4369 -445
rect 4399 -479 4406 -445
rect 4364 -488 4406 -479
rect 4440 -445 4482 -436
rect 4440 -479 4447 -445
rect 4477 -479 4482 -445
rect 4440 -484 4482 -479
rect 4516 -472 4544 -412
tri 4589 -425 4611 -403 se
rect 4611 -410 4626 -402
tri 4611 -425 4626 -410 nw
tri 4583 -431 4589 -425 se
rect 4589 -431 4598 -425
rect 4302 -516 4330 -506
tri 4330 -516 4354 -492 sw
rect 4302 -548 4344 -516
tri 4361 -524 4362 -523 sw
rect 4361 -548 4362 -524
tri 4364 -525 4401 -488 ne
rect 4401 -516 4406 -488
tri 4406 -516 4432 -490 sw
rect 4516 -506 4525 -472
rect 4516 -516 4544 -506
rect 4401 -525 4485 -516
tri 4401 -544 4420 -525 ne
rect 4420 -544 4485 -525
rect 4302 -570 4362 -548
rect 4484 -548 4485 -544
rect 4502 -548 4544 -516
rect 4484 -570 4544 -548
rect 4390 -586 4407 -572
rect 4439 -586 4456 -572
tri 4227 -622 4249 -600 se
rect 4249 -607 4264 -586
tri 4249 -622 4264 -607 nw
rect 4583 -607 4598 -431
tri 4598 -438 4611 -425 nw
rect 4684 -506 4699 -278
tri 4221 -628 4227 -622 se
rect 4227 -628 4236 -622
rect 4221 -644 4236 -628
tri 4236 -635 4249 -622 nw
rect 4390 -630 4407 -616
rect 4439 -630 4456 -616
tri 4583 -622 4598 -607 ne
tri 4598 -622 4620 -600 sw
rect 4221 -680 4236 -672
rect 4302 -644 4362 -630
rect 4317 -654 4362 -644
rect 4317 -672 4345 -654
tri 4221 -695 4236 -680 ne
tri 4236 -695 4258 -673 sw
rect 4302 -682 4345 -672
rect 4360 -658 4362 -654
rect 4484 -644 4544 -630
tri 4598 -635 4611 -622 ne
rect 4611 -628 4620 -622
tri 4620 -628 4626 -622 sw
rect 4484 -654 4529 -644
rect 4360 -682 4434 -658
rect 4302 -686 4434 -682
tri 4434 -686 4462 -658 sw
rect 4484 -668 4486 -654
tri 4484 -670 4486 -668 ne
rect 4498 -672 4529 -654
rect 4498 -682 4544 -672
rect 4611 -643 4626 -628
tri 4236 -707 4248 -695 ne
rect 4248 -700 4258 -695
tri 4258 -700 4263 -695 sw
rect 4147 -1046 4162 -818
rect 4248 -808 4263 -700
rect 4302 -742 4330 -686
tri 4422 -704 4440 -686 ne
rect 4440 -706 4462 -686
tri 4462 -706 4482 -686 sw
tri 4498 -700 4516 -682 ne
rect 4321 -776 4330 -742
rect 4364 -715 4406 -714
rect 4364 -749 4369 -715
rect 4399 -749 4406 -715
rect 4364 -758 4406 -749
rect 4440 -715 4482 -706
rect 4440 -749 4447 -715
rect 4477 -749 4482 -715
rect 4440 -754 4482 -749
rect 4516 -742 4544 -682
tri 4589 -695 4611 -673 se
rect 4611 -680 4626 -672
tri 4611 -695 4626 -680 nw
tri 4583 -701 4589 -695 se
rect 4589 -701 4598 -695
rect 4302 -786 4330 -776
tri 4330 -786 4354 -762 sw
rect 4248 -856 4264 -808
rect 4302 -818 4344 -786
tri 4361 -794 4362 -793 sw
rect 4361 -818 4362 -794
tri 4364 -795 4401 -758 ne
rect 4401 -786 4406 -758
tri 4406 -786 4432 -760 sw
rect 4516 -776 4525 -742
rect 4516 -786 4544 -776
rect 4401 -795 4485 -786
tri 4401 -814 4420 -795 ne
rect 4420 -814 4485 -795
rect 4302 -840 4362 -818
rect 4484 -818 4485 -814
rect 4502 -818 4544 -786
rect 4484 -840 4544 -818
rect 4390 -856 4407 -842
rect 4439 -856 4456 -842
tri 4227 -892 4249 -870 se
rect 4249 -877 4264 -856
tri 4249 -892 4264 -877 nw
rect 4583 -877 4598 -701
tri 4598 -708 4611 -695 nw
rect 4684 -776 4699 -548
tri 4221 -898 4227 -892 se
rect 4227 -898 4236 -892
rect 4221 -914 4236 -898
tri 4236 -905 4249 -892 nw
rect 4390 -900 4407 -886
rect 4439 -900 4456 -886
tri 4583 -892 4598 -877 ne
tri 4598 -892 4620 -870 sw
rect 4221 -950 4236 -942
rect 4302 -914 4362 -900
rect 4317 -924 4362 -914
rect 4317 -942 4345 -924
tri 4221 -965 4236 -950 ne
tri 4236 -965 4258 -943 sw
rect 4302 -952 4345 -942
rect 4360 -928 4362 -924
rect 4484 -914 4544 -900
tri 4598 -905 4611 -892 ne
rect 4611 -898 4620 -892
tri 4620 -898 4626 -892 sw
rect 4484 -924 4529 -914
rect 4360 -952 4434 -928
rect 4302 -956 4434 -952
tri 4434 -956 4462 -928 sw
rect 4484 -938 4486 -924
tri 4484 -940 4486 -938 ne
rect 4498 -942 4529 -924
rect 4498 -952 4544 -942
rect 4611 -913 4626 -898
tri 4236 -977 4248 -965 ne
rect 4248 -970 4258 -965
tri 4258 -970 4263 -965 sw
rect 4147 -1316 4162 -1088
rect 4248 -1126 4263 -970
rect 4302 -1012 4330 -956
tri 4422 -974 4440 -956 ne
rect 4440 -976 4462 -956
tri 4462 -976 4482 -956 sw
tri 4498 -970 4516 -952 ne
rect 4321 -1046 4330 -1012
rect 4364 -985 4406 -984
rect 4364 -1019 4369 -985
rect 4399 -1019 4406 -985
rect 4364 -1028 4406 -1019
rect 4440 -985 4482 -976
rect 4440 -1019 4447 -985
rect 4477 -1019 4482 -985
rect 4440 -1024 4482 -1019
rect 4516 -1012 4544 -952
tri 4589 -965 4611 -943 se
rect 4611 -950 4626 -942
tri 4611 -965 4626 -950 nw
tri 4583 -971 4589 -965 se
rect 4589 -971 4598 -965
rect 4302 -1056 4330 -1046
tri 4330 -1056 4354 -1032 sw
rect 4302 -1088 4344 -1056
tri 4361 -1064 4362 -1063 sw
rect 4361 -1088 4362 -1064
tri 4364 -1065 4401 -1028 ne
rect 4401 -1056 4406 -1028
tri 4406 -1056 4432 -1030 sw
rect 4516 -1046 4525 -1012
rect 4516 -1056 4544 -1046
rect 4401 -1065 4485 -1056
tri 4401 -1084 4420 -1065 ne
rect 4420 -1084 4485 -1065
rect 4302 -1110 4362 -1088
rect 4484 -1088 4485 -1084
rect 4502 -1088 4544 -1056
rect 4484 -1110 4544 -1088
rect 4390 -1126 4407 -1112
rect 4439 -1126 4456 -1112
tri 4227 -1162 4249 -1140 se
rect 4249 -1147 4264 -1126
tri 4249 -1162 4264 -1147 nw
rect 4583 -1147 4598 -971
tri 4598 -978 4611 -965 nw
rect 4684 -1046 4699 -818
tri 4221 -1168 4227 -1162 se
rect 4227 -1168 4236 -1162
rect 4221 -1184 4236 -1168
tri 4236 -1175 4249 -1162 nw
rect 4390 -1170 4407 -1156
rect 4439 -1170 4456 -1156
tri 4583 -1162 4598 -1147 ne
tri 4598 -1162 4620 -1140 sw
rect 4221 -1220 4236 -1212
rect 4302 -1184 4362 -1170
rect 4317 -1194 4362 -1184
rect 4317 -1212 4345 -1194
tri 4221 -1235 4236 -1220 ne
tri 4236 -1235 4258 -1213 sw
rect 4302 -1222 4345 -1212
rect 4360 -1198 4362 -1194
rect 4484 -1184 4544 -1170
tri 4598 -1175 4611 -1162 ne
rect 4611 -1168 4620 -1162
tri 4620 -1168 4626 -1162 sw
rect 4484 -1194 4529 -1184
rect 4360 -1222 4434 -1198
rect 4302 -1226 4434 -1222
tri 4434 -1226 4462 -1198 sw
rect 4484 -1208 4486 -1194
tri 4484 -1210 4486 -1208 ne
rect 4498 -1212 4529 -1194
rect 4498 -1222 4544 -1212
rect 4611 -1183 4626 -1168
tri 4236 -1247 4248 -1235 ne
rect 4248 -1240 4258 -1235
tri 4258 -1240 4263 -1235 sw
rect 4147 -1586 4162 -1358
rect 4248 -1348 4263 -1240
rect 4302 -1282 4330 -1226
tri 4422 -1244 4440 -1226 ne
rect 4440 -1246 4462 -1226
tri 4462 -1246 4482 -1226 sw
tri 4498 -1240 4516 -1222 ne
rect 4321 -1316 4330 -1282
rect 4364 -1255 4406 -1254
rect 4364 -1289 4369 -1255
rect 4399 -1289 4406 -1255
rect 4364 -1298 4406 -1289
rect 4440 -1255 4482 -1246
rect 4440 -1289 4447 -1255
rect 4477 -1289 4482 -1255
rect 4440 -1294 4482 -1289
rect 4516 -1282 4544 -1222
tri 4589 -1235 4611 -1213 se
rect 4611 -1220 4626 -1212
tri 4611 -1235 4626 -1220 nw
tri 4583 -1241 4589 -1235 se
rect 4589 -1241 4598 -1235
rect 4302 -1326 4330 -1316
tri 4330 -1326 4354 -1302 sw
rect 4248 -1396 4264 -1348
rect 4302 -1358 4344 -1326
tri 4361 -1334 4362 -1333 sw
rect 4361 -1358 4362 -1334
tri 4364 -1335 4401 -1298 ne
rect 4401 -1326 4406 -1298
tri 4406 -1326 4432 -1300 sw
rect 4516 -1316 4525 -1282
rect 4516 -1326 4544 -1316
rect 4401 -1335 4485 -1326
tri 4401 -1354 4420 -1335 ne
rect 4420 -1354 4485 -1335
rect 4302 -1380 4362 -1358
rect 4484 -1358 4485 -1354
rect 4502 -1358 4544 -1326
rect 4484 -1380 4544 -1358
rect 4390 -1396 4407 -1382
rect 4439 -1396 4456 -1382
tri 4227 -1432 4249 -1410 se
rect 4249 -1417 4264 -1396
tri 4249 -1432 4264 -1417 nw
rect 4583 -1417 4598 -1241
tri 4598 -1248 4611 -1235 nw
rect 4684 -1316 4699 -1088
tri 4221 -1438 4227 -1432 se
rect 4227 -1438 4236 -1432
rect 4221 -1454 4236 -1438
tri 4236 -1445 4249 -1432 nw
rect 4390 -1440 4407 -1426
rect 4439 -1440 4456 -1426
tri 4583 -1432 4598 -1417 ne
tri 4598 -1432 4620 -1410 sw
rect 4221 -1490 4236 -1482
rect 4302 -1454 4362 -1440
rect 4317 -1464 4362 -1454
rect 4317 -1482 4345 -1464
tri 4221 -1505 4236 -1490 ne
tri 4236 -1505 4258 -1483 sw
rect 4302 -1492 4345 -1482
rect 4360 -1468 4362 -1464
rect 4484 -1454 4544 -1440
tri 4598 -1445 4611 -1432 ne
rect 4611 -1438 4620 -1432
tri 4620 -1438 4626 -1432 sw
rect 4484 -1464 4529 -1454
rect 4360 -1492 4434 -1468
rect 4302 -1496 4434 -1492
tri 4434 -1496 4462 -1468 sw
rect 4484 -1478 4486 -1464
tri 4484 -1480 4486 -1478 ne
rect 4498 -1482 4529 -1464
rect 4498 -1492 4544 -1482
rect 4611 -1453 4626 -1438
tri 4236 -1517 4248 -1505 ne
rect 4248 -1510 4258 -1505
tri 4258 -1510 4263 -1505 sw
rect 4147 -1856 4162 -1628
rect 4248 -1666 4263 -1510
rect 4302 -1552 4330 -1496
tri 4422 -1514 4440 -1496 ne
rect 4440 -1516 4462 -1496
tri 4462 -1516 4482 -1496 sw
tri 4498 -1510 4516 -1492 ne
rect 4321 -1586 4330 -1552
rect 4364 -1525 4406 -1524
rect 4364 -1559 4369 -1525
rect 4399 -1559 4406 -1525
rect 4364 -1568 4406 -1559
rect 4440 -1525 4482 -1516
rect 4440 -1559 4447 -1525
rect 4477 -1559 4482 -1525
rect 4440 -1564 4482 -1559
rect 4516 -1552 4544 -1492
tri 4589 -1505 4611 -1483 se
rect 4611 -1490 4626 -1482
tri 4611 -1505 4626 -1490 nw
tri 4583 -1511 4589 -1505 se
rect 4589 -1511 4598 -1505
rect 4302 -1596 4330 -1586
tri 4330 -1596 4354 -1572 sw
rect 4302 -1628 4344 -1596
tri 4361 -1604 4362 -1603 sw
rect 4361 -1628 4362 -1604
tri 4364 -1605 4401 -1568 ne
rect 4401 -1596 4406 -1568
tri 4406 -1596 4432 -1570 sw
rect 4516 -1586 4525 -1552
rect 4516 -1596 4544 -1586
rect 4401 -1605 4485 -1596
tri 4401 -1624 4420 -1605 ne
rect 4420 -1624 4485 -1605
rect 4302 -1650 4362 -1628
rect 4484 -1628 4485 -1624
rect 4502 -1628 4544 -1596
rect 4484 -1650 4544 -1628
rect 4390 -1666 4407 -1652
rect 4439 -1666 4456 -1652
tri 4227 -1702 4249 -1680 se
rect 4249 -1687 4264 -1666
tri 4249 -1702 4264 -1687 nw
rect 4583 -1687 4598 -1511
tri 4598 -1518 4611 -1505 nw
rect 4684 -1586 4699 -1358
tri 4221 -1708 4227 -1702 se
rect 4227 -1708 4236 -1702
rect 4221 -1724 4236 -1708
tri 4236 -1715 4249 -1702 nw
rect 4390 -1710 4407 -1696
rect 4439 -1710 4456 -1696
tri 4583 -1702 4598 -1687 ne
tri 4598 -1702 4620 -1680 sw
rect 4221 -1760 4236 -1752
rect 4302 -1724 4362 -1710
rect 4317 -1734 4362 -1724
rect 4317 -1752 4345 -1734
tri 4221 -1775 4236 -1760 ne
tri 4236 -1775 4258 -1753 sw
rect 4302 -1762 4345 -1752
rect 4360 -1738 4362 -1734
rect 4484 -1724 4544 -1710
tri 4598 -1715 4611 -1702 ne
rect 4611 -1708 4620 -1702
tri 4620 -1708 4626 -1702 sw
rect 4484 -1734 4529 -1724
rect 4360 -1762 4434 -1738
rect 4302 -1766 4434 -1762
tri 4434 -1766 4462 -1738 sw
rect 4484 -1748 4486 -1734
tri 4484 -1750 4486 -1748 ne
rect 4498 -1752 4529 -1734
rect 4498 -1762 4544 -1752
rect 4611 -1723 4626 -1708
tri 4236 -1787 4248 -1775 ne
rect 4248 -1780 4258 -1775
tri 4258 -1780 4263 -1775 sw
rect 4147 -2126 4162 -1898
rect 4248 -1888 4263 -1780
rect 4302 -1822 4330 -1766
tri 4422 -1784 4440 -1766 ne
rect 4440 -1786 4462 -1766
tri 4462 -1786 4482 -1766 sw
tri 4498 -1780 4516 -1762 ne
rect 4321 -1856 4330 -1822
rect 4364 -1795 4406 -1794
rect 4364 -1829 4369 -1795
rect 4399 -1829 4406 -1795
rect 4364 -1838 4406 -1829
rect 4440 -1795 4482 -1786
rect 4440 -1829 4447 -1795
rect 4477 -1829 4482 -1795
rect 4440 -1834 4482 -1829
rect 4516 -1822 4544 -1762
tri 4589 -1775 4611 -1753 se
rect 4611 -1760 4626 -1752
tri 4611 -1775 4626 -1760 nw
tri 4583 -1781 4589 -1775 se
rect 4589 -1781 4598 -1775
rect 4302 -1866 4330 -1856
tri 4330 -1866 4354 -1842 sw
rect 4248 -1936 4264 -1888
rect 4302 -1898 4344 -1866
tri 4361 -1874 4362 -1873 sw
rect 4361 -1898 4362 -1874
tri 4364 -1875 4401 -1838 ne
rect 4401 -1866 4406 -1838
tri 4406 -1866 4432 -1840 sw
rect 4516 -1856 4525 -1822
rect 4516 -1866 4544 -1856
rect 4401 -1875 4485 -1866
tri 4401 -1894 4420 -1875 ne
rect 4420 -1894 4485 -1875
rect 4302 -1920 4362 -1898
rect 4484 -1898 4485 -1894
rect 4502 -1898 4544 -1866
rect 4484 -1920 4544 -1898
rect 4390 -1936 4407 -1922
rect 4439 -1936 4456 -1922
tri 4227 -1972 4249 -1950 se
rect 4249 -1957 4264 -1936
tri 4249 -1972 4264 -1957 nw
rect 4583 -1957 4598 -1781
tri 4598 -1788 4611 -1775 nw
rect 4684 -1856 4699 -1628
tri 4221 -1978 4227 -1972 se
rect 4227 -1978 4236 -1972
rect 4221 -1994 4236 -1978
tri 4236 -1985 4249 -1972 nw
rect 4390 -1980 4407 -1966
rect 4439 -1980 4456 -1966
tri 4583 -1972 4598 -1957 ne
tri 4598 -1972 4620 -1950 sw
rect 4221 -2030 4236 -2022
rect 4302 -1994 4362 -1980
rect 4317 -2004 4362 -1994
rect 4317 -2022 4345 -2004
tri 4221 -2045 4236 -2030 ne
tri 4236 -2045 4258 -2023 sw
rect 4302 -2032 4345 -2022
rect 4360 -2008 4362 -2004
rect 4484 -1994 4544 -1980
tri 4598 -1985 4611 -1972 ne
rect 4611 -1978 4620 -1972
tri 4620 -1978 4626 -1972 sw
rect 4484 -2004 4529 -1994
rect 4360 -2032 4434 -2008
rect 4302 -2036 4434 -2032
tri 4434 -2036 4462 -2008 sw
rect 4484 -2018 4486 -2004
tri 4484 -2020 4486 -2018 ne
rect 4498 -2022 4529 -2004
rect 4498 -2032 4544 -2022
rect 4611 -1993 4626 -1978
tri 4236 -2057 4248 -2045 ne
rect 4248 -2050 4258 -2045
tri 4258 -2050 4263 -2045 sw
rect 4147 -2396 4162 -2168
rect 4248 -2206 4263 -2050
rect 4302 -2092 4330 -2036
tri 4422 -2054 4440 -2036 ne
rect 4440 -2056 4462 -2036
tri 4462 -2056 4482 -2036 sw
tri 4498 -2050 4516 -2032 ne
rect 4321 -2126 4330 -2092
rect 4364 -2065 4406 -2064
rect 4364 -2099 4369 -2065
rect 4399 -2099 4406 -2065
rect 4364 -2108 4406 -2099
rect 4440 -2065 4482 -2056
rect 4440 -2099 4447 -2065
rect 4477 -2099 4482 -2065
rect 4440 -2104 4482 -2099
rect 4516 -2092 4544 -2032
tri 4589 -2045 4611 -2023 se
rect 4611 -2030 4626 -2022
tri 4611 -2045 4626 -2030 nw
tri 4583 -2051 4589 -2045 se
rect 4589 -2051 4598 -2045
rect 4302 -2136 4330 -2126
tri 4330 -2136 4354 -2112 sw
rect 4302 -2168 4344 -2136
tri 4361 -2144 4362 -2143 sw
rect 4361 -2168 4362 -2144
tri 4364 -2145 4401 -2108 ne
rect 4401 -2136 4406 -2108
tri 4406 -2136 4432 -2110 sw
rect 4516 -2126 4525 -2092
rect 4516 -2136 4544 -2126
rect 4401 -2145 4485 -2136
tri 4401 -2164 4420 -2145 ne
rect 4420 -2164 4485 -2145
rect 4302 -2190 4362 -2168
rect 4484 -2168 4485 -2164
rect 4502 -2168 4544 -2136
rect 4484 -2190 4544 -2168
rect 4390 -2206 4407 -2192
rect 4439 -2206 4456 -2192
tri 4227 -2242 4249 -2220 se
rect 4249 -2227 4264 -2206
tri 4249 -2242 4264 -2227 nw
rect 4583 -2227 4598 -2051
tri 4598 -2058 4611 -2045 nw
rect 4684 -2126 4699 -1898
tri 4221 -2248 4227 -2242 se
rect 4227 -2248 4236 -2242
rect 4221 -2264 4236 -2248
tri 4236 -2255 4249 -2242 nw
rect 4390 -2250 4407 -2236
rect 4439 -2250 4456 -2236
tri 4583 -2242 4598 -2227 ne
tri 4598 -2242 4620 -2220 sw
rect 4221 -2300 4236 -2292
rect 4302 -2264 4362 -2250
rect 4317 -2274 4362 -2264
rect 4317 -2292 4345 -2274
tri 4221 -2315 4236 -2300 ne
tri 4236 -2315 4258 -2293 sw
rect 4302 -2302 4345 -2292
rect 4360 -2278 4362 -2274
rect 4484 -2264 4544 -2250
tri 4598 -2255 4611 -2242 ne
rect 4611 -2248 4620 -2242
tri 4620 -2248 4626 -2242 sw
rect 4484 -2274 4529 -2264
rect 4360 -2302 4434 -2278
rect 4302 -2306 4434 -2302
tri 4434 -2306 4462 -2278 sw
rect 4484 -2288 4486 -2274
tri 4484 -2290 4486 -2288 ne
rect 4498 -2292 4529 -2274
rect 4498 -2302 4544 -2292
rect 4611 -2263 4626 -2248
tri 4236 -2327 4248 -2315 ne
rect 4248 -2320 4258 -2315
tri 4258 -2320 4263 -2315 sw
rect 4147 -2524 4162 -2438
rect 4248 -2476 4263 -2320
rect 4302 -2362 4330 -2306
tri 4422 -2324 4440 -2306 ne
rect 4440 -2326 4462 -2306
tri 4462 -2326 4482 -2306 sw
tri 4498 -2320 4516 -2302 ne
rect 4321 -2396 4330 -2362
rect 4364 -2335 4406 -2334
rect 4364 -2369 4369 -2335
rect 4399 -2369 4406 -2335
rect 4364 -2378 4406 -2369
rect 4440 -2335 4482 -2326
rect 4440 -2369 4447 -2335
rect 4477 -2369 4482 -2335
rect 4440 -2374 4482 -2369
rect 4516 -2362 4544 -2302
tri 4589 -2315 4611 -2293 se
rect 4611 -2300 4626 -2292
tri 4611 -2315 4626 -2300 nw
tri 4583 -2321 4589 -2315 se
rect 4589 -2321 4598 -2315
rect 4302 -2406 4330 -2396
tri 4330 -2406 4354 -2382 sw
rect 4302 -2438 4344 -2406
tri 4361 -2414 4362 -2413 sw
rect 4361 -2438 4362 -2414
tri 4364 -2415 4401 -2378 ne
rect 4401 -2406 4406 -2378
tri 4406 -2406 4432 -2380 sw
rect 4516 -2396 4525 -2362
rect 4516 -2406 4544 -2396
rect 4401 -2415 4485 -2406
tri 4401 -2434 4420 -2415 ne
rect 4420 -2434 4485 -2415
rect 4302 -2460 4362 -2438
rect 4484 -2438 4485 -2434
rect 4502 -2438 4544 -2406
rect 4484 -2460 4544 -2438
rect 4390 -2476 4407 -2462
rect 4439 -2476 4456 -2462
rect 4583 -2476 4598 -2321
tri 4598 -2328 4611 -2315 nw
rect 4684 -2396 4699 -2168
rect 4684 -2524 4699 -2438
rect 4727 1654 4742 1844
tri 4807 1808 4829 1830 se
rect 4829 1823 4844 1892
tri 4829 1808 4844 1823 nw
rect 5163 1823 5178 1892
tri 4801 1802 4807 1808 se
rect 4807 1802 4816 1808
rect 4801 1786 4816 1802
tri 4816 1795 4829 1808 nw
rect 4970 1800 4987 1814
rect 5019 1800 5036 1814
tri 5163 1808 5178 1823 ne
tri 5178 1808 5200 1830 sw
rect 4801 1750 4816 1758
rect 4882 1786 4942 1800
rect 4897 1776 4942 1786
rect 4897 1758 4925 1776
tri 4801 1735 4816 1750 ne
tri 4816 1735 4838 1757 sw
rect 4882 1748 4925 1758
rect 4940 1772 4942 1776
rect 5064 1786 5124 1800
tri 5178 1795 5191 1808 ne
rect 5191 1802 5200 1808
tri 5200 1802 5206 1808 sw
rect 5064 1776 5109 1786
rect 4940 1748 5014 1772
rect 4882 1744 5014 1748
tri 5014 1744 5042 1772 sw
rect 5064 1762 5066 1776
tri 5064 1760 5066 1762 ne
rect 5078 1758 5109 1776
rect 5078 1748 5124 1758
rect 5191 1787 5206 1802
tri 4816 1723 4828 1735 ne
rect 4828 1730 4838 1735
tri 4838 1730 4843 1735 sw
rect 4727 1384 4742 1612
rect 4828 1574 4843 1730
rect 4882 1688 4910 1744
tri 5002 1726 5020 1744 ne
rect 5020 1724 5042 1744
tri 5042 1724 5062 1744 sw
tri 5078 1730 5096 1748 ne
rect 4901 1654 4910 1688
rect 4944 1715 4986 1716
rect 4944 1681 4949 1715
rect 4979 1681 4986 1715
rect 4944 1672 4986 1681
rect 5020 1715 5062 1724
rect 5020 1681 5027 1715
rect 5057 1681 5062 1715
rect 5020 1676 5062 1681
rect 5096 1688 5124 1748
tri 5169 1735 5191 1757 se
rect 5191 1750 5206 1758
tri 5191 1735 5206 1750 nw
tri 5163 1729 5169 1735 se
rect 5169 1729 5178 1735
rect 4882 1644 4910 1654
tri 4910 1644 4934 1668 sw
rect 4882 1612 4924 1644
tri 4941 1636 4942 1637 sw
rect 4941 1612 4942 1636
tri 4944 1635 4981 1672 ne
rect 4981 1644 4986 1672
tri 4986 1644 5012 1670 sw
rect 5096 1654 5105 1688
rect 5096 1644 5124 1654
rect 4981 1635 5065 1644
tri 4981 1616 5000 1635 ne
rect 5000 1616 5065 1635
rect 4882 1590 4942 1612
rect 5064 1612 5065 1616
rect 5082 1612 5124 1644
rect 5064 1590 5124 1612
rect 4970 1574 4987 1588
rect 5019 1574 5036 1588
tri 4807 1538 4829 1560 se
rect 4829 1553 4844 1574
tri 4829 1538 4844 1553 nw
rect 5163 1553 5178 1729
tri 5178 1722 5191 1735 nw
rect 5264 1654 5279 1844
tri 4801 1532 4807 1538 se
rect 4807 1532 4816 1538
rect 4801 1516 4816 1532
tri 4816 1525 4829 1538 nw
rect 4970 1530 4987 1544
rect 5019 1530 5036 1544
tri 5163 1538 5178 1553 ne
tri 5178 1538 5200 1560 sw
rect 4801 1480 4816 1488
rect 4882 1516 4942 1530
rect 4897 1506 4942 1516
rect 4897 1488 4925 1506
tri 4801 1465 4816 1480 ne
tri 4816 1465 4838 1487 sw
rect 4882 1478 4925 1488
rect 4940 1502 4942 1506
rect 5064 1516 5124 1530
tri 5178 1525 5191 1538 ne
rect 5191 1532 5200 1538
tri 5200 1532 5206 1538 sw
rect 5064 1506 5109 1516
rect 4940 1478 5014 1502
rect 4882 1474 5014 1478
tri 5014 1474 5042 1502 sw
rect 5064 1492 5066 1506
tri 5064 1490 5066 1492 ne
rect 5078 1488 5109 1506
rect 5078 1478 5124 1488
rect 5191 1517 5206 1532
tri 4816 1453 4828 1465 ne
rect 4828 1460 4838 1465
tri 4838 1460 4843 1465 sw
rect 4727 1114 4742 1342
rect 4828 1352 4843 1460
rect 4882 1418 4910 1474
tri 5002 1456 5020 1474 ne
rect 5020 1454 5042 1474
tri 5042 1454 5062 1474 sw
tri 5078 1460 5096 1478 ne
rect 4901 1384 4910 1418
rect 4944 1445 4986 1446
rect 4944 1411 4949 1445
rect 4979 1411 4986 1445
rect 4944 1402 4986 1411
rect 5020 1445 5062 1454
rect 5020 1411 5027 1445
rect 5057 1411 5062 1445
rect 5020 1406 5062 1411
rect 5096 1418 5124 1478
tri 5169 1465 5191 1487 se
rect 5191 1480 5206 1488
tri 5191 1465 5206 1480 nw
tri 5163 1459 5169 1465 se
rect 5169 1459 5178 1465
rect 4882 1374 4910 1384
tri 4910 1374 4934 1398 sw
rect 4828 1304 4844 1352
rect 4882 1342 4924 1374
tri 4941 1366 4942 1367 sw
rect 4941 1342 4942 1366
tri 4944 1365 4981 1402 ne
rect 4981 1374 4986 1402
tri 4986 1374 5012 1400 sw
rect 5096 1384 5105 1418
rect 5096 1374 5124 1384
rect 4981 1365 5065 1374
tri 4981 1346 5000 1365 ne
rect 5000 1346 5065 1365
rect 4882 1320 4942 1342
rect 5064 1342 5065 1346
rect 5082 1342 5124 1374
rect 5064 1320 5124 1342
rect 4970 1304 4987 1318
rect 5019 1304 5036 1318
tri 4807 1268 4829 1290 se
rect 4829 1283 4844 1304
tri 4829 1268 4844 1283 nw
rect 5163 1283 5178 1459
tri 5178 1452 5191 1465 nw
rect 5264 1384 5279 1612
tri 4801 1262 4807 1268 se
rect 4807 1262 4816 1268
rect 4801 1246 4816 1262
tri 4816 1255 4829 1268 nw
rect 4970 1260 4987 1274
rect 5019 1260 5036 1274
tri 5163 1268 5178 1283 ne
tri 5178 1268 5200 1290 sw
rect 4801 1210 4816 1218
rect 4882 1246 4942 1260
rect 4897 1236 4942 1246
rect 4897 1218 4925 1236
tri 4801 1195 4816 1210 ne
tri 4816 1195 4838 1217 sw
rect 4882 1208 4925 1218
rect 4940 1232 4942 1236
rect 5064 1246 5124 1260
tri 5178 1255 5191 1268 ne
rect 5191 1262 5200 1268
tri 5200 1262 5206 1268 sw
rect 5064 1236 5109 1246
rect 4940 1208 5014 1232
rect 4882 1204 5014 1208
tri 5014 1204 5042 1232 sw
rect 5064 1222 5066 1236
tri 5064 1220 5066 1222 ne
rect 5078 1218 5109 1236
rect 5078 1208 5124 1218
rect 5191 1247 5206 1262
tri 4816 1183 4828 1195 ne
rect 4828 1190 4838 1195
tri 4838 1190 4843 1195 sw
rect 4727 844 4742 1072
rect 4828 1034 4843 1190
rect 4882 1148 4910 1204
tri 5002 1186 5020 1204 ne
rect 5020 1184 5042 1204
tri 5042 1184 5062 1204 sw
tri 5078 1190 5096 1208 ne
rect 4901 1114 4910 1148
rect 4944 1175 4986 1176
rect 4944 1141 4949 1175
rect 4979 1141 4986 1175
rect 4944 1132 4986 1141
rect 5020 1175 5062 1184
rect 5020 1141 5027 1175
rect 5057 1141 5062 1175
rect 5020 1136 5062 1141
rect 5096 1148 5124 1208
tri 5169 1195 5191 1217 se
rect 5191 1210 5206 1218
tri 5191 1195 5206 1210 nw
tri 5163 1189 5169 1195 se
rect 5169 1189 5178 1195
rect 4882 1104 4910 1114
tri 4910 1104 4934 1128 sw
rect 4882 1072 4924 1104
tri 4941 1096 4942 1097 sw
rect 4941 1072 4942 1096
tri 4944 1095 4981 1132 ne
rect 4981 1104 4986 1132
tri 4986 1104 5012 1130 sw
rect 5096 1114 5105 1148
rect 5096 1104 5124 1114
rect 4981 1095 5065 1104
tri 4981 1076 5000 1095 ne
rect 5000 1076 5065 1095
rect 4882 1050 4942 1072
rect 5064 1072 5065 1076
rect 5082 1072 5124 1104
rect 5064 1050 5124 1072
rect 4970 1034 4987 1048
rect 5019 1034 5036 1048
tri 4807 998 4829 1020 se
rect 4829 1013 4844 1034
tri 4829 998 4844 1013 nw
rect 5163 1013 5178 1189
tri 5178 1182 5191 1195 nw
rect 5264 1114 5279 1342
tri 4801 992 4807 998 se
rect 4807 992 4816 998
rect 4801 976 4816 992
tri 4816 985 4829 998 nw
rect 4970 990 4987 1004
rect 5019 990 5036 1004
tri 5163 998 5178 1013 ne
tri 5178 998 5200 1020 sw
rect 4801 940 4816 948
rect 4882 976 4942 990
rect 4897 966 4942 976
rect 4897 948 4925 966
tri 4801 925 4816 940 ne
tri 4816 925 4838 947 sw
rect 4882 938 4925 948
rect 4940 962 4942 966
rect 5064 976 5124 990
tri 5178 985 5191 998 ne
rect 5191 992 5200 998
tri 5200 992 5206 998 sw
rect 5064 966 5109 976
rect 4940 938 5014 962
rect 4882 934 5014 938
tri 5014 934 5042 962 sw
rect 5064 952 5066 966
tri 5064 950 5066 952 ne
rect 5078 948 5109 966
rect 5078 938 5124 948
rect 5191 977 5206 992
tri 4816 913 4828 925 ne
rect 4828 920 4838 925
tri 4838 920 4843 925 sw
rect 4727 574 4742 802
rect 4828 812 4843 920
rect 4882 878 4910 934
tri 5002 916 5020 934 ne
rect 5020 914 5042 934
tri 5042 914 5062 934 sw
tri 5078 920 5096 938 ne
rect 4901 844 4910 878
rect 4944 905 4986 906
rect 4944 871 4949 905
rect 4979 871 4986 905
rect 4944 862 4986 871
rect 5020 905 5062 914
rect 5020 871 5027 905
rect 5057 871 5062 905
rect 5020 866 5062 871
rect 5096 878 5124 938
tri 5169 925 5191 947 se
rect 5191 940 5206 948
tri 5191 925 5206 940 nw
tri 5163 919 5169 925 se
rect 5169 919 5178 925
rect 4882 834 4910 844
tri 4910 834 4934 858 sw
rect 4828 764 4844 812
rect 4882 802 4924 834
tri 4941 826 4942 827 sw
rect 4941 802 4942 826
tri 4944 825 4981 862 ne
rect 4981 834 4986 862
tri 4986 834 5012 860 sw
rect 5096 844 5105 878
rect 5096 834 5124 844
rect 4981 825 5065 834
tri 4981 806 5000 825 ne
rect 5000 806 5065 825
rect 4882 780 4942 802
rect 5064 802 5065 806
rect 5082 802 5124 834
rect 5064 780 5124 802
rect 4970 764 4987 778
rect 5019 764 5036 778
tri 4807 728 4829 750 se
rect 4829 743 4844 764
tri 4829 728 4844 743 nw
rect 5163 743 5178 919
tri 5178 912 5191 925 nw
rect 5264 844 5279 1072
tri 4801 722 4807 728 se
rect 4807 722 4816 728
rect 4801 706 4816 722
tri 4816 715 4829 728 nw
rect 4970 720 4987 734
rect 5019 720 5036 734
tri 5163 728 5178 743 ne
tri 5178 728 5200 750 sw
rect 4801 670 4816 678
rect 4882 706 4942 720
rect 4897 696 4942 706
rect 4897 678 4925 696
tri 4801 655 4816 670 ne
tri 4816 655 4838 677 sw
rect 4882 668 4925 678
rect 4940 692 4942 696
rect 5064 706 5124 720
tri 5178 715 5191 728 ne
rect 5191 722 5200 728
tri 5200 722 5206 728 sw
rect 5064 696 5109 706
rect 4940 668 5014 692
rect 4882 664 5014 668
tri 5014 664 5042 692 sw
rect 5064 682 5066 696
tri 5064 680 5066 682 ne
rect 5078 678 5109 696
rect 5078 668 5124 678
rect 5191 707 5206 722
tri 4816 643 4828 655 ne
rect 4828 650 4838 655
tri 4838 650 4843 655 sw
rect 4727 304 4742 532
rect 4828 494 4843 650
rect 4882 608 4910 664
tri 5002 646 5020 664 ne
rect 5020 644 5042 664
tri 5042 644 5062 664 sw
tri 5078 650 5096 668 ne
rect 4901 574 4910 608
rect 4944 635 4986 636
rect 4944 601 4949 635
rect 4979 601 4986 635
rect 4944 592 4986 601
rect 5020 635 5062 644
rect 5020 601 5027 635
rect 5057 601 5062 635
rect 5020 596 5062 601
rect 5096 608 5124 668
tri 5169 655 5191 677 se
rect 5191 670 5206 678
tri 5191 655 5206 670 nw
tri 5163 649 5169 655 se
rect 5169 649 5178 655
rect 4882 564 4910 574
tri 4910 564 4934 588 sw
rect 4882 532 4924 564
tri 4941 556 4942 557 sw
rect 4941 532 4942 556
tri 4944 555 4981 592 ne
rect 4981 564 4986 592
tri 4986 564 5012 590 sw
rect 5096 574 5105 608
rect 5096 564 5124 574
rect 4981 555 5065 564
tri 4981 536 5000 555 ne
rect 5000 536 5065 555
rect 4882 510 4942 532
rect 5064 532 5065 536
rect 5082 532 5124 564
rect 5064 510 5124 532
rect 4970 494 4987 508
rect 5019 494 5036 508
tri 4807 458 4829 480 se
rect 4829 473 4844 494
tri 4829 458 4844 473 nw
rect 5163 473 5178 649
tri 5178 642 5191 655 nw
rect 5264 574 5279 802
tri 4801 452 4807 458 se
rect 4807 452 4816 458
rect 4801 436 4816 452
tri 4816 445 4829 458 nw
rect 4970 450 4987 464
rect 5019 450 5036 464
tri 5163 458 5178 473 ne
tri 5178 458 5200 480 sw
rect 4801 400 4816 408
rect 4882 436 4942 450
rect 4897 426 4942 436
rect 4897 408 4925 426
tri 4801 385 4816 400 ne
tri 4816 385 4838 407 sw
rect 4882 398 4925 408
rect 4940 422 4942 426
rect 5064 436 5124 450
tri 5178 445 5191 458 ne
rect 5191 452 5200 458
tri 5200 452 5206 458 sw
rect 5064 426 5109 436
rect 4940 398 5014 422
rect 4882 394 5014 398
tri 5014 394 5042 422 sw
rect 5064 412 5066 426
tri 5064 410 5066 412 ne
rect 5078 408 5109 426
rect 5078 398 5124 408
rect 5191 437 5206 452
tri 4816 373 4828 385 ne
rect 4828 380 4838 385
tri 4838 380 4843 385 sw
rect 4727 34 4742 262
rect 4828 272 4843 380
rect 4882 338 4910 394
tri 5002 376 5020 394 ne
rect 5020 374 5042 394
tri 5042 374 5062 394 sw
tri 5078 380 5096 398 ne
rect 4901 304 4910 338
rect 4944 365 4986 366
rect 4944 331 4949 365
rect 4979 331 4986 365
rect 4944 322 4986 331
rect 5020 365 5062 374
rect 5020 331 5027 365
rect 5057 331 5062 365
rect 5020 326 5062 331
rect 5096 338 5124 398
tri 5169 385 5191 407 se
rect 5191 400 5206 408
tri 5191 385 5206 400 nw
tri 5163 379 5169 385 se
rect 5169 379 5178 385
rect 4882 294 4910 304
tri 4910 294 4934 318 sw
rect 4828 224 4844 272
rect 4882 262 4924 294
tri 4941 286 4942 287 sw
rect 4941 262 4942 286
tri 4944 285 4981 322 ne
rect 4981 294 4986 322
tri 4986 294 5012 320 sw
rect 5096 304 5105 338
rect 5096 294 5124 304
rect 4981 285 5065 294
tri 4981 266 5000 285 ne
rect 5000 266 5065 285
rect 4882 240 4942 262
rect 5064 262 5065 266
rect 5082 262 5124 294
rect 5064 240 5124 262
rect 4970 224 4987 238
rect 5019 224 5036 238
tri 4807 188 4829 210 se
rect 4829 203 4844 224
tri 4829 188 4844 203 nw
rect 5163 203 5178 379
tri 5178 372 5191 385 nw
rect 5264 304 5279 532
tri 4801 182 4807 188 se
rect 4807 182 4816 188
rect 4801 166 4816 182
tri 4816 175 4829 188 nw
rect 4970 180 4987 194
rect 5019 180 5036 194
tri 5163 188 5178 203 ne
tri 5178 188 5200 210 sw
rect 4801 130 4816 138
rect 4882 166 4942 180
rect 4897 156 4942 166
rect 4897 138 4925 156
tri 4801 115 4816 130 ne
tri 4816 115 4838 137 sw
rect 4882 128 4925 138
rect 4940 152 4942 156
rect 5064 166 5124 180
tri 5178 175 5191 188 ne
rect 5191 182 5200 188
tri 5200 182 5206 188 sw
rect 5064 156 5109 166
rect 4940 128 5014 152
rect 4882 124 5014 128
tri 5014 124 5042 152 sw
rect 5064 142 5066 156
tri 5064 140 5066 142 ne
rect 5078 138 5109 156
rect 5078 128 5124 138
rect 5191 167 5206 182
tri 4816 103 4828 115 ne
rect 4828 110 4838 115
tri 4838 110 4843 115 sw
rect 4727 -236 4742 -8
rect 4828 -46 4843 110
rect 4882 68 4910 124
tri 5002 106 5020 124 ne
rect 5020 104 5042 124
tri 5042 104 5062 124 sw
tri 5078 110 5096 128 ne
rect 4901 34 4910 68
rect 4944 95 4986 96
rect 4944 61 4949 95
rect 4979 61 4986 95
rect 4944 52 4986 61
rect 5020 95 5062 104
rect 5020 61 5027 95
rect 5057 61 5062 95
rect 5020 56 5062 61
rect 5096 68 5124 128
tri 5169 115 5191 137 se
rect 5191 130 5206 138
tri 5191 115 5206 130 nw
tri 5163 109 5169 115 se
rect 5169 109 5178 115
rect 4882 24 4910 34
tri 4910 24 4934 48 sw
rect 4882 -8 4924 24
tri 4941 16 4942 17 sw
rect 4941 -8 4942 16
tri 4944 15 4981 52 ne
rect 4981 24 4986 52
tri 4986 24 5012 50 sw
rect 5096 34 5105 68
rect 5096 24 5124 34
rect 4981 15 5065 24
tri 4981 -4 5000 15 ne
rect 5000 -4 5065 15
rect 4882 -30 4942 -8
rect 5064 -8 5065 -4
rect 5082 -8 5124 24
rect 5064 -30 5124 -8
rect 4970 -46 4987 -32
rect 5019 -46 5036 -32
tri 4807 -82 4829 -60 se
rect 4829 -67 4844 -46
tri 4829 -82 4844 -67 nw
rect 5163 -67 5178 109
tri 5178 102 5191 115 nw
rect 5264 34 5279 262
tri 4801 -88 4807 -82 se
rect 4807 -88 4816 -82
rect 4801 -104 4816 -88
tri 4816 -95 4829 -82 nw
rect 4970 -90 4987 -76
rect 5019 -90 5036 -76
tri 5163 -82 5178 -67 ne
tri 5178 -82 5200 -60 sw
rect 4801 -140 4816 -132
rect 4882 -104 4942 -90
rect 4897 -114 4942 -104
rect 4897 -132 4925 -114
tri 4801 -155 4816 -140 ne
tri 4816 -155 4838 -133 sw
rect 4882 -142 4925 -132
rect 4940 -118 4942 -114
rect 5064 -104 5124 -90
tri 5178 -95 5191 -82 ne
rect 5191 -88 5200 -82
tri 5200 -88 5206 -82 sw
rect 5064 -114 5109 -104
rect 4940 -142 5014 -118
rect 4882 -146 5014 -142
tri 5014 -146 5042 -118 sw
rect 5064 -128 5066 -114
tri 5064 -130 5066 -128 ne
rect 5078 -132 5109 -114
rect 5078 -142 5124 -132
rect 5191 -103 5206 -88
tri 4816 -167 4828 -155 ne
rect 4828 -160 4838 -155
tri 4838 -160 4843 -155 sw
rect 4727 -506 4742 -278
rect 4828 -268 4843 -160
rect 4882 -202 4910 -146
tri 5002 -164 5020 -146 ne
rect 5020 -166 5042 -146
tri 5042 -166 5062 -146 sw
tri 5078 -160 5096 -142 ne
rect 4901 -236 4910 -202
rect 4944 -175 4986 -174
rect 4944 -209 4949 -175
rect 4979 -209 4986 -175
rect 4944 -218 4986 -209
rect 5020 -175 5062 -166
rect 5020 -209 5027 -175
rect 5057 -209 5062 -175
rect 5020 -214 5062 -209
rect 5096 -202 5124 -142
tri 5169 -155 5191 -133 se
rect 5191 -140 5206 -132
tri 5191 -155 5206 -140 nw
tri 5163 -161 5169 -155 se
rect 5169 -161 5178 -155
rect 4882 -246 4910 -236
tri 4910 -246 4934 -222 sw
rect 4828 -316 4844 -268
rect 4882 -278 4924 -246
tri 4941 -254 4942 -253 sw
rect 4941 -278 4942 -254
tri 4944 -255 4981 -218 ne
rect 4981 -246 4986 -218
tri 4986 -246 5012 -220 sw
rect 5096 -236 5105 -202
rect 5096 -246 5124 -236
rect 4981 -255 5065 -246
tri 4981 -274 5000 -255 ne
rect 5000 -274 5065 -255
rect 4882 -300 4942 -278
rect 5064 -278 5065 -274
rect 5082 -278 5124 -246
rect 5064 -300 5124 -278
rect 4970 -316 4987 -302
rect 5019 -316 5036 -302
tri 4807 -352 4829 -330 se
rect 4829 -337 4844 -316
tri 4829 -352 4844 -337 nw
rect 5163 -337 5178 -161
tri 5178 -168 5191 -155 nw
rect 5264 -236 5279 -8
tri 4801 -358 4807 -352 se
rect 4807 -358 4816 -352
rect 4801 -374 4816 -358
tri 4816 -365 4829 -352 nw
rect 4970 -360 4987 -346
rect 5019 -360 5036 -346
tri 5163 -352 5178 -337 ne
tri 5178 -352 5200 -330 sw
rect 4801 -410 4816 -402
rect 4882 -374 4942 -360
rect 4897 -384 4942 -374
rect 4897 -402 4925 -384
tri 4801 -425 4816 -410 ne
tri 4816 -425 4838 -403 sw
rect 4882 -412 4925 -402
rect 4940 -388 4942 -384
rect 5064 -374 5124 -360
tri 5178 -365 5191 -352 ne
rect 5191 -358 5200 -352
tri 5200 -358 5206 -352 sw
rect 5064 -384 5109 -374
rect 4940 -412 5014 -388
rect 4882 -416 5014 -412
tri 5014 -416 5042 -388 sw
rect 5064 -398 5066 -384
tri 5064 -400 5066 -398 ne
rect 5078 -402 5109 -384
rect 5078 -412 5124 -402
rect 5191 -373 5206 -358
tri 4816 -437 4828 -425 ne
rect 4828 -430 4838 -425
tri 4838 -430 4843 -425 sw
rect 4727 -776 4742 -548
rect 4828 -586 4843 -430
rect 4882 -472 4910 -416
tri 5002 -434 5020 -416 ne
rect 5020 -436 5042 -416
tri 5042 -436 5062 -416 sw
tri 5078 -430 5096 -412 ne
rect 4901 -506 4910 -472
rect 4944 -445 4986 -444
rect 4944 -479 4949 -445
rect 4979 -479 4986 -445
rect 4944 -488 4986 -479
rect 5020 -445 5062 -436
rect 5020 -479 5027 -445
rect 5057 -479 5062 -445
rect 5020 -484 5062 -479
rect 5096 -472 5124 -412
tri 5169 -425 5191 -403 se
rect 5191 -410 5206 -402
tri 5191 -425 5206 -410 nw
tri 5163 -431 5169 -425 se
rect 5169 -431 5178 -425
rect 4882 -516 4910 -506
tri 4910 -516 4934 -492 sw
rect 4882 -548 4924 -516
tri 4941 -524 4942 -523 sw
rect 4941 -548 4942 -524
tri 4944 -525 4981 -488 ne
rect 4981 -516 4986 -488
tri 4986 -516 5012 -490 sw
rect 5096 -506 5105 -472
rect 5096 -516 5124 -506
rect 4981 -525 5065 -516
tri 4981 -544 5000 -525 ne
rect 5000 -544 5065 -525
rect 4882 -570 4942 -548
rect 5064 -548 5065 -544
rect 5082 -548 5124 -516
rect 5064 -570 5124 -548
rect 4970 -586 4987 -572
rect 5019 -586 5036 -572
tri 4807 -622 4829 -600 se
rect 4829 -607 4844 -586
tri 4829 -622 4844 -607 nw
rect 5163 -607 5178 -431
tri 5178 -438 5191 -425 nw
rect 5264 -506 5279 -278
tri 4801 -628 4807 -622 se
rect 4807 -628 4816 -622
rect 4801 -644 4816 -628
tri 4816 -635 4829 -622 nw
rect 4970 -630 4987 -616
rect 5019 -630 5036 -616
tri 5163 -622 5178 -607 ne
tri 5178 -622 5200 -600 sw
rect 4801 -680 4816 -672
rect 4882 -644 4942 -630
rect 4897 -654 4942 -644
rect 4897 -672 4925 -654
tri 4801 -695 4816 -680 ne
tri 4816 -695 4838 -673 sw
rect 4882 -682 4925 -672
rect 4940 -658 4942 -654
rect 5064 -644 5124 -630
tri 5178 -635 5191 -622 ne
rect 5191 -628 5200 -622
tri 5200 -628 5206 -622 sw
rect 5064 -654 5109 -644
rect 4940 -682 5014 -658
rect 4882 -686 5014 -682
tri 5014 -686 5042 -658 sw
rect 5064 -668 5066 -654
tri 5064 -670 5066 -668 ne
rect 5078 -672 5109 -654
rect 5078 -682 5124 -672
rect 5191 -643 5206 -628
tri 4816 -707 4828 -695 ne
rect 4828 -700 4838 -695
tri 4838 -700 4843 -695 sw
rect 4727 -1046 4742 -818
rect 4828 -808 4843 -700
rect 4882 -742 4910 -686
tri 5002 -704 5020 -686 ne
rect 5020 -706 5042 -686
tri 5042 -706 5062 -686 sw
tri 5078 -700 5096 -682 ne
rect 4901 -776 4910 -742
rect 4944 -715 4986 -714
rect 4944 -749 4949 -715
rect 4979 -749 4986 -715
rect 4944 -758 4986 -749
rect 5020 -715 5062 -706
rect 5020 -749 5027 -715
rect 5057 -749 5062 -715
rect 5020 -754 5062 -749
rect 5096 -742 5124 -682
tri 5169 -695 5191 -673 se
rect 5191 -680 5206 -672
tri 5191 -695 5206 -680 nw
tri 5163 -701 5169 -695 se
rect 5169 -701 5178 -695
rect 4882 -786 4910 -776
tri 4910 -786 4934 -762 sw
rect 4828 -856 4844 -808
rect 4882 -818 4924 -786
tri 4941 -794 4942 -793 sw
rect 4941 -818 4942 -794
tri 4944 -795 4981 -758 ne
rect 4981 -786 4986 -758
tri 4986 -786 5012 -760 sw
rect 5096 -776 5105 -742
rect 5096 -786 5124 -776
rect 4981 -795 5065 -786
tri 4981 -814 5000 -795 ne
rect 5000 -814 5065 -795
rect 4882 -840 4942 -818
rect 5064 -818 5065 -814
rect 5082 -818 5124 -786
rect 5064 -840 5124 -818
rect 4970 -856 4987 -842
rect 5019 -856 5036 -842
tri 4807 -892 4829 -870 se
rect 4829 -877 4844 -856
tri 4829 -892 4844 -877 nw
rect 5163 -877 5178 -701
tri 5178 -708 5191 -695 nw
rect 5264 -776 5279 -548
tri 4801 -898 4807 -892 se
rect 4807 -898 4816 -892
rect 4801 -914 4816 -898
tri 4816 -905 4829 -892 nw
rect 4970 -900 4987 -886
rect 5019 -900 5036 -886
tri 5163 -892 5178 -877 ne
tri 5178 -892 5200 -870 sw
rect 4801 -950 4816 -942
rect 4882 -914 4942 -900
rect 4897 -924 4942 -914
rect 4897 -942 4925 -924
tri 4801 -965 4816 -950 ne
tri 4816 -965 4838 -943 sw
rect 4882 -952 4925 -942
rect 4940 -928 4942 -924
rect 5064 -914 5124 -900
tri 5178 -905 5191 -892 ne
rect 5191 -898 5200 -892
tri 5200 -898 5206 -892 sw
rect 5064 -924 5109 -914
rect 4940 -952 5014 -928
rect 4882 -956 5014 -952
tri 5014 -956 5042 -928 sw
rect 5064 -938 5066 -924
tri 5064 -940 5066 -938 ne
rect 5078 -942 5109 -924
rect 5078 -952 5124 -942
rect 5191 -913 5206 -898
tri 4816 -977 4828 -965 ne
rect 4828 -970 4838 -965
tri 4838 -970 4843 -965 sw
rect 4727 -1316 4742 -1088
rect 4828 -1126 4843 -970
rect 4882 -1012 4910 -956
tri 5002 -974 5020 -956 ne
rect 5020 -976 5042 -956
tri 5042 -976 5062 -956 sw
tri 5078 -970 5096 -952 ne
rect 4901 -1046 4910 -1012
rect 4944 -985 4986 -984
rect 4944 -1019 4949 -985
rect 4979 -1019 4986 -985
rect 4944 -1028 4986 -1019
rect 5020 -985 5062 -976
rect 5020 -1019 5027 -985
rect 5057 -1019 5062 -985
rect 5020 -1024 5062 -1019
rect 5096 -1012 5124 -952
tri 5169 -965 5191 -943 se
rect 5191 -950 5206 -942
tri 5191 -965 5206 -950 nw
tri 5163 -971 5169 -965 se
rect 5169 -971 5178 -965
rect 4882 -1056 4910 -1046
tri 4910 -1056 4934 -1032 sw
rect 4882 -1088 4924 -1056
tri 4941 -1064 4942 -1063 sw
rect 4941 -1088 4942 -1064
tri 4944 -1065 4981 -1028 ne
rect 4981 -1056 4986 -1028
tri 4986 -1056 5012 -1030 sw
rect 5096 -1046 5105 -1012
rect 5096 -1056 5124 -1046
rect 4981 -1065 5065 -1056
tri 4981 -1084 5000 -1065 ne
rect 5000 -1084 5065 -1065
rect 4882 -1110 4942 -1088
rect 5064 -1088 5065 -1084
rect 5082 -1088 5124 -1056
rect 5064 -1110 5124 -1088
rect 4970 -1126 4987 -1112
rect 5019 -1126 5036 -1112
tri 4807 -1162 4829 -1140 se
rect 4829 -1147 4844 -1126
tri 4829 -1162 4844 -1147 nw
rect 5163 -1147 5178 -971
tri 5178 -978 5191 -965 nw
rect 5264 -1046 5279 -818
tri 4801 -1168 4807 -1162 se
rect 4807 -1168 4816 -1162
rect 4801 -1184 4816 -1168
tri 4816 -1175 4829 -1162 nw
rect 4970 -1170 4987 -1156
rect 5019 -1170 5036 -1156
tri 5163 -1162 5178 -1147 ne
tri 5178 -1162 5200 -1140 sw
rect 4801 -1220 4816 -1212
rect 4882 -1184 4942 -1170
rect 4897 -1194 4942 -1184
rect 4897 -1212 4925 -1194
tri 4801 -1235 4816 -1220 ne
tri 4816 -1235 4838 -1213 sw
rect 4882 -1222 4925 -1212
rect 4940 -1198 4942 -1194
rect 5064 -1184 5124 -1170
tri 5178 -1175 5191 -1162 ne
rect 5191 -1168 5200 -1162
tri 5200 -1168 5206 -1162 sw
rect 5064 -1194 5109 -1184
rect 4940 -1222 5014 -1198
rect 4882 -1226 5014 -1222
tri 5014 -1226 5042 -1198 sw
rect 5064 -1208 5066 -1194
tri 5064 -1210 5066 -1208 ne
rect 5078 -1212 5109 -1194
rect 5078 -1222 5124 -1212
rect 5191 -1183 5206 -1168
tri 4816 -1247 4828 -1235 ne
rect 4828 -1240 4838 -1235
tri 4838 -1240 4843 -1235 sw
rect 4727 -1586 4742 -1358
rect 4828 -1348 4843 -1240
rect 4882 -1282 4910 -1226
tri 5002 -1244 5020 -1226 ne
rect 5020 -1246 5042 -1226
tri 5042 -1246 5062 -1226 sw
tri 5078 -1240 5096 -1222 ne
rect 4901 -1316 4910 -1282
rect 4944 -1255 4986 -1254
rect 4944 -1289 4949 -1255
rect 4979 -1289 4986 -1255
rect 4944 -1298 4986 -1289
rect 5020 -1255 5062 -1246
rect 5020 -1289 5027 -1255
rect 5057 -1289 5062 -1255
rect 5020 -1294 5062 -1289
rect 5096 -1282 5124 -1222
tri 5169 -1235 5191 -1213 se
rect 5191 -1220 5206 -1212
tri 5191 -1235 5206 -1220 nw
tri 5163 -1241 5169 -1235 se
rect 5169 -1241 5178 -1235
rect 4882 -1326 4910 -1316
tri 4910 -1326 4934 -1302 sw
rect 4828 -1396 4844 -1348
rect 4882 -1358 4924 -1326
tri 4941 -1334 4942 -1333 sw
rect 4941 -1358 4942 -1334
tri 4944 -1335 4981 -1298 ne
rect 4981 -1326 4986 -1298
tri 4986 -1326 5012 -1300 sw
rect 5096 -1316 5105 -1282
rect 5096 -1326 5124 -1316
rect 4981 -1335 5065 -1326
tri 4981 -1354 5000 -1335 ne
rect 5000 -1354 5065 -1335
rect 4882 -1380 4942 -1358
rect 5064 -1358 5065 -1354
rect 5082 -1358 5124 -1326
rect 5064 -1380 5124 -1358
rect 4970 -1396 4987 -1382
rect 5019 -1396 5036 -1382
tri 4807 -1432 4829 -1410 se
rect 4829 -1417 4844 -1396
tri 4829 -1432 4844 -1417 nw
rect 5163 -1417 5178 -1241
tri 5178 -1248 5191 -1235 nw
rect 5264 -1316 5279 -1088
tri 4801 -1438 4807 -1432 se
rect 4807 -1438 4816 -1432
rect 4801 -1454 4816 -1438
tri 4816 -1445 4829 -1432 nw
rect 4970 -1440 4987 -1426
rect 5019 -1440 5036 -1426
tri 5163 -1432 5178 -1417 ne
tri 5178 -1432 5200 -1410 sw
rect 4801 -1490 4816 -1482
rect 4882 -1454 4942 -1440
rect 4897 -1464 4942 -1454
rect 4897 -1482 4925 -1464
tri 4801 -1505 4816 -1490 ne
tri 4816 -1505 4838 -1483 sw
rect 4882 -1492 4925 -1482
rect 4940 -1468 4942 -1464
rect 5064 -1454 5124 -1440
tri 5178 -1445 5191 -1432 ne
rect 5191 -1438 5200 -1432
tri 5200 -1438 5206 -1432 sw
rect 5064 -1464 5109 -1454
rect 4940 -1492 5014 -1468
rect 4882 -1496 5014 -1492
tri 5014 -1496 5042 -1468 sw
rect 5064 -1478 5066 -1464
tri 5064 -1480 5066 -1478 ne
rect 5078 -1482 5109 -1464
rect 5078 -1492 5124 -1482
rect 5191 -1453 5206 -1438
tri 4816 -1517 4828 -1505 ne
rect 4828 -1510 4838 -1505
tri 4838 -1510 4843 -1505 sw
rect 4727 -1856 4742 -1628
rect 4828 -1666 4843 -1510
rect 4882 -1552 4910 -1496
tri 5002 -1514 5020 -1496 ne
rect 5020 -1516 5042 -1496
tri 5042 -1516 5062 -1496 sw
tri 5078 -1510 5096 -1492 ne
rect 4901 -1586 4910 -1552
rect 4944 -1525 4986 -1524
rect 4944 -1559 4949 -1525
rect 4979 -1559 4986 -1525
rect 4944 -1568 4986 -1559
rect 5020 -1525 5062 -1516
rect 5020 -1559 5027 -1525
rect 5057 -1559 5062 -1525
rect 5020 -1564 5062 -1559
rect 5096 -1552 5124 -1492
tri 5169 -1505 5191 -1483 se
rect 5191 -1490 5206 -1482
tri 5191 -1505 5206 -1490 nw
tri 5163 -1511 5169 -1505 se
rect 5169 -1511 5178 -1505
rect 4882 -1596 4910 -1586
tri 4910 -1596 4934 -1572 sw
rect 4882 -1628 4924 -1596
tri 4941 -1604 4942 -1603 sw
rect 4941 -1628 4942 -1604
tri 4944 -1605 4981 -1568 ne
rect 4981 -1596 4986 -1568
tri 4986 -1596 5012 -1570 sw
rect 5096 -1586 5105 -1552
rect 5096 -1596 5124 -1586
rect 4981 -1605 5065 -1596
tri 4981 -1624 5000 -1605 ne
rect 5000 -1624 5065 -1605
rect 4882 -1650 4942 -1628
rect 5064 -1628 5065 -1624
rect 5082 -1628 5124 -1596
rect 5064 -1650 5124 -1628
rect 4970 -1666 4987 -1652
rect 5019 -1666 5036 -1652
tri 4807 -1702 4829 -1680 se
rect 4829 -1687 4844 -1666
tri 4829 -1702 4844 -1687 nw
rect 5163 -1687 5178 -1511
tri 5178 -1518 5191 -1505 nw
rect 5264 -1586 5279 -1358
tri 4801 -1708 4807 -1702 se
rect 4807 -1708 4816 -1702
rect 4801 -1724 4816 -1708
tri 4816 -1715 4829 -1702 nw
rect 4970 -1710 4987 -1696
rect 5019 -1710 5036 -1696
tri 5163 -1702 5178 -1687 ne
tri 5178 -1702 5200 -1680 sw
rect 4801 -1760 4816 -1752
rect 4882 -1724 4942 -1710
rect 4897 -1734 4942 -1724
rect 4897 -1752 4925 -1734
tri 4801 -1775 4816 -1760 ne
tri 4816 -1775 4838 -1753 sw
rect 4882 -1762 4925 -1752
rect 4940 -1738 4942 -1734
rect 5064 -1724 5124 -1710
tri 5178 -1715 5191 -1702 ne
rect 5191 -1708 5200 -1702
tri 5200 -1708 5206 -1702 sw
rect 5064 -1734 5109 -1724
rect 4940 -1762 5014 -1738
rect 4882 -1766 5014 -1762
tri 5014 -1766 5042 -1738 sw
rect 5064 -1748 5066 -1734
tri 5064 -1750 5066 -1748 ne
rect 5078 -1752 5109 -1734
rect 5078 -1762 5124 -1752
rect 5191 -1723 5206 -1708
tri 4816 -1787 4828 -1775 ne
rect 4828 -1780 4838 -1775
tri 4838 -1780 4843 -1775 sw
rect 4727 -2126 4742 -1898
rect 4828 -1888 4843 -1780
rect 4882 -1822 4910 -1766
tri 5002 -1784 5020 -1766 ne
rect 5020 -1786 5042 -1766
tri 5042 -1786 5062 -1766 sw
tri 5078 -1780 5096 -1762 ne
rect 4901 -1856 4910 -1822
rect 4944 -1795 4986 -1794
rect 4944 -1829 4949 -1795
rect 4979 -1829 4986 -1795
rect 4944 -1838 4986 -1829
rect 5020 -1795 5062 -1786
rect 5020 -1829 5027 -1795
rect 5057 -1829 5062 -1795
rect 5020 -1834 5062 -1829
rect 5096 -1822 5124 -1762
tri 5169 -1775 5191 -1753 se
rect 5191 -1760 5206 -1752
tri 5191 -1775 5206 -1760 nw
tri 5163 -1781 5169 -1775 se
rect 5169 -1781 5178 -1775
rect 4882 -1866 4910 -1856
tri 4910 -1866 4934 -1842 sw
rect 4828 -1936 4844 -1888
rect 4882 -1898 4924 -1866
tri 4941 -1874 4942 -1873 sw
rect 4941 -1898 4942 -1874
tri 4944 -1875 4981 -1838 ne
rect 4981 -1866 4986 -1838
tri 4986 -1866 5012 -1840 sw
rect 5096 -1856 5105 -1822
rect 5096 -1866 5124 -1856
rect 4981 -1875 5065 -1866
tri 4981 -1894 5000 -1875 ne
rect 5000 -1894 5065 -1875
rect 4882 -1920 4942 -1898
rect 5064 -1898 5065 -1894
rect 5082 -1898 5124 -1866
rect 5064 -1920 5124 -1898
rect 4970 -1936 4987 -1922
rect 5019 -1936 5036 -1922
tri 4807 -1972 4829 -1950 se
rect 4829 -1957 4844 -1936
tri 4829 -1972 4844 -1957 nw
rect 5163 -1957 5178 -1781
tri 5178 -1788 5191 -1775 nw
rect 5264 -1856 5279 -1628
tri 4801 -1978 4807 -1972 se
rect 4807 -1978 4816 -1972
rect 4801 -1994 4816 -1978
tri 4816 -1985 4829 -1972 nw
rect 4970 -1980 4987 -1966
rect 5019 -1980 5036 -1966
tri 5163 -1972 5178 -1957 ne
tri 5178 -1972 5200 -1950 sw
rect 4801 -2030 4816 -2022
rect 4882 -1994 4942 -1980
rect 4897 -2004 4942 -1994
rect 4897 -2022 4925 -2004
tri 4801 -2045 4816 -2030 ne
tri 4816 -2045 4838 -2023 sw
rect 4882 -2032 4925 -2022
rect 4940 -2008 4942 -2004
rect 5064 -1994 5124 -1980
tri 5178 -1985 5191 -1972 ne
rect 5191 -1978 5200 -1972
tri 5200 -1978 5206 -1972 sw
rect 5064 -2004 5109 -1994
rect 4940 -2032 5014 -2008
rect 4882 -2036 5014 -2032
tri 5014 -2036 5042 -2008 sw
rect 5064 -2018 5066 -2004
tri 5064 -2020 5066 -2018 ne
rect 5078 -2022 5109 -2004
rect 5078 -2032 5124 -2022
rect 5191 -1993 5206 -1978
tri 4816 -2057 4828 -2045 ne
rect 4828 -2050 4838 -2045
tri 4838 -2050 4843 -2045 sw
rect 4727 -2396 4742 -2168
rect 4828 -2206 4843 -2050
rect 4882 -2092 4910 -2036
tri 5002 -2054 5020 -2036 ne
rect 5020 -2056 5042 -2036
tri 5042 -2056 5062 -2036 sw
tri 5078 -2050 5096 -2032 ne
rect 4901 -2126 4910 -2092
rect 4944 -2065 4986 -2064
rect 4944 -2099 4949 -2065
rect 4979 -2099 4986 -2065
rect 4944 -2108 4986 -2099
rect 5020 -2065 5062 -2056
rect 5020 -2099 5027 -2065
rect 5057 -2099 5062 -2065
rect 5020 -2104 5062 -2099
rect 5096 -2092 5124 -2032
tri 5169 -2045 5191 -2023 se
rect 5191 -2030 5206 -2022
tri 5191 -2045 5206 -2030 nw
tri 5163 -2051 5169 -2045 se
rect 5169 -2051 5178 -2045
rect 4882 -2136 4910 -2126
tri 4910 -2136 4934 -2112 sw
rect 4882 -2168 4924 -2136
tri 4941 -2144 4942 -2143 sw
rect 4941 -2168 4942 -2144
tri 4944 -2145 4981 -2108 ne
rect 4981 -2136 4986 -2108
tri 4986 -2136 5012 -2110 sw
rect 5096 -2126 5105 -2092
rect 5096 -2136 5124 -2126
rect 4981 -2145 5065 -2136
tri 4981 -2164 5000 -2145 ne
rect 5000 -2164 5065 -2145
rect 4882 -2190 4942 -2168
rect 5064 -2168 5065 -2164
rect 5082 -2168 5124 -2136
rect 5064 -2190 5124 -2168
rect 4970 -2206 4987 -2192
rect 5019 -2206 5036 -2192
tri 4807 -2242 4829 -2220 se
rect 4829 -2227 4844 -2206
tri 4829 -2242 4844 -2227 nw
rect 5163 -2227 5178 -2051
tri 5178 -2058 5191 -2045 nw
rect 5264 -2126 5279 -1898
tri 4801 -2248 4807 -2242 se
rect 4807 -2248 4816 -2242
rect 4801 -2264 4816 -2248
tri 4816 -2255 4829 -2242 nw
rect 4970 -2250 4987 -2236
rect 5019 -2250 5036 -2236
tri 5163 -2242 5178 -2227 ne
tri 5178 -2242 5200 -2220 sw
rect 4801 -2300 4816 -2292
rect 4882 -2264 4942 -2250
rect 4897 -2274 4942 -2264
rect 4897 -2292 4925 -2274
tri 4801 -2315 4816 -2300 ne
tri 4816 -2315 4838 -2293 sw
rect 4882 -2302 4925 -2292
rect 4940 -2278 4942 -2274
rect 5064 -2264 5124 -2250
tri 5178 -2255 5191 -2242 ne
rect 5191 -2248 5200 -2242
tri 5200 -2248 5206 -2242 sw
rect 5064 -2274 5109 -2264
rect 4940 -2302 5014 -2278
rect 4882 -2306 5014 -2302
tri 5014 -2306 5042 -2278 sw
rect 5064 -2288 5066 -2274
tri 5064 -2290 5066 -2288 ne
rect 5078 -2292 5109 -2274
rect 5078 -2302 5124 -2292
rect 5191 -2263 5206 -2248
tri 4816 -2327 4828 -2315 ne
rect 4828 -2320 4838 -2315
tri 4838 -2320 4843 -2315 sw
rect 4727 -2524 4742 -2438
rect 4828 -2476 4843 -2320
rect 4882 -2362 4910 -2306
tri 5002 -2324 5020 -2306 ne
rect 5020 -2326 5042 -2306
tri 5042 -2326 5062 -2306 sw
tri 5078 -2320 5096 -2302 ne
rect 4901 -2396 4910 -2362
rect 4944 -2335 4986 -2334
rect 4944 -2369 4949 -2335
rect 4979 -2369 4986 -2335
rect 4944 -2378 4986 -2369
rect 5020 -2335 5062 -2326
rect 5020 -2369 5027 -2335
rect 5057 -2369 5062 -2335
rect 5020 -2374 5062 -2369
rect 5096 -2362 5124 -2302
tri 5169 -2315 5191 -2293 se
rect 5191 -2300 5206 -2292
tri 5191 -2315 5206 -2300 nw
tri 5163 -2321 5169 -2315 se
rect 5169 -2321 5178 -2315
rect 4882 -2406 4910 -2396
tri 4910 -2406 4934 -2382 sw
rect 4882 -2438 4924 -2406
tri 4941 -2414 4942 -2413 sw
rect 4941 -2438 4942 -2414
tri 4944 -2415 4981 -2378 ne
rect 4981 -2406 4986 -2378
tri 4986 -2406 5012 -2380 sw
rect 5096 -2396 5105 -2362
rect 5096 -2406 5124 -2396
rect 4981 -2415 5065 -2406
tri 4981 -2434 5000 -2415 ne
rect 5000 -2434 5065 -2415
rect 4882 -2460 4942 -2438
rect 5064 -2438 5065 -2434
rect 5082 -2438 5124 -2406
rect 5064 -2460 5124 -2438
rect 4970 -2476 4987 -2462
rect 5019 -2476 5036 -2462
rect 5163 -2476 5178 -2321
tri 5178 -2328 5191 -2315 nw
rect 5264 -2396 5279 -2168
rect 5264 -2524 5279 -2438
rect 5307 1654 5322 1844
tri 5387 1808 5409 1830 se
rect 5409 1823 5424 1892
tri 5409 1808 5424 1823 nw
rect 5743 1823 5758 1892
tri 5381 1802 5387 1808 se
rect 5387 1802 5396 1808
rect 5381 1786 5396 1802
tri 5396 1795 5409 1808 nw
rect 5550 1800 5567 1814
rect 5599 1800 5616 1814
tri 5743 1808 5758 1823 ne
tri 5758 1808 5780 1830 sw
rect 5381 1750 5396 1758
rect 5462 1786 5522 1800
rect 5477 1776 5522 1786
rect 5477 1758 5505 1776
tri 5381 1735 5396 1750 ne
tri 5396 1735 5418 1757 sw
rect 5462 1748 5505 1758
rect 5520 1772 5522 1776
rect 5644 1786 5704 1800
tri 5758 1795 5771 1808 ne
rect 5771 1802 5780 1808
tri 5780 1802 5786 1808 sw
rect 5644 1776 5689 1786
rect 5520 1748 5594 1772
rect 5462 1744 5594 1748
tri 5594 1744 5622 1772 sw
rect 5644 1762 5646 1776
tri 5644 1760 5646 1762 ne
rect 5658 1758 5689 1776
rect 5658 1748 5704 1758
rect 5771 1787 5786 1802
tri 5396 1723 5408 1735 ne
rect 5408 1730 5418 1735
tri 5418 1730 5423 1735 sw
rect 5307 1384 5322 1612
rect 5408 1574 5423 1730
rect 5462 1688 5490 1744
tri 5582 1726 5600 1744 ne
rect 5600 1724 5622 1744
tri 5622 1724 5642 1744 sw
tri 5658 1730 5676 1748 ne
rect 5481 1654 5490 1688
rect 5524 1715 5566 1716
rect 5524 1681 5529 1715
rect 5559 1681 5566 1715
rect 5524 1672 5566 1681
rect 5600 1715 5642 1724
rect 5600 1681 5607 1715
rect 5637 1681 5642 1715
rect 5600 1676 5642 1681
rect 5676 1688 5704 1748
tri 5749 1735 5771 1757 se
rect 5771 1750 5786 1758
tri 5771 1735 5786 1750 nw
tri 5743 1729 5749 1735 se
rect 5749 1729 5758 1735
rect 5462 1644 5490 1654
tri 5490 1644 5514 1668 sw
rect 5462 1612 5504 1644
tri 5521 1636 5522 1637 sw
rect 5521 1612 5522 1636
tri 5524 1635 5561 1672 ne
rect 5561 1644 5566 1672
tri 5566 1644 5592 1670 sw
rect 5676 1654 5685 1688
rect 5676 1644 5704 1654
rect 5561 1635 5645 1644
tri 5561 1616 5580 1635 ne
rect 5580 1616 5645 1635
rect 5462 1590 5522 1612
rect 5644 1612 5645 1616
rect 5662 1612 5704 1644
rect 5644 1590 5704 1612
rect 5550 1574 5567 1588
rect 5599 1574 5616 1588
tri 5387 1538 5409 1560 se
rect 5409 1553 5424 1574
tri 5409 1538 5424 1553 nw
rect 5743 1553 5758 1729
tri 5758 1722 5771 1735 nw
rect 5844 1654 5859 1844
tri 5381 1532 5387 1538 se
rect 5387 1532 5396 1538
rect 5381 1516 5396 1532
tri 5396 1525 5409 1538 nw
rect 5550 1530 5567 1544
rect 5599 1530 5616 1544
tri 5743 1538 5758 1553 ne
tri 5758 1538 5780 1560 sw
rect 5381 1480 5396 1488
rect 5462 1516 5522 1530
rect 5477 1506 5522 1516
rect 5477 1488 5505 1506
tri 5381 1465 5396 1480 ne
tri 5396 1465 5418 1487 sw
rect 5462 1478 5505 1488
rect 5520 1502 5522 1506
rect 5644 1516 5704 1530
tri 5758 1525 5771 1538 ne
rect 5771 1532 5780 1538
tri 5780 1532 5786 1538 sw
rect 5644 1506 5689 1516
rect 5520 1478 5594 1502
rect 5462 1474 5594 1478
tri 5594 1474 5622 1502 sw
rect 5644 1492 5646 1506
tri 5644 1490 5646 1492 ne
rect 5658 1488 5689 1506
rect 5658 1478 5704 1488
rect 5771 1517 5786 1532
tri 5396 1453 5408 1465 ne
rect 5408 1460 5418 1465
tri 5418 1460 5423 1465 sw
rect 5307 1114 5322 1342
rect 5408 1352 5423 1460
rect 5462 1418 5490 1474
tri 5582 1456 5600 1474 ne
rect 5600 1454 5622 1474
tri 5622 1454 5642 1474 sw
tri 5658 1460 5676 1478 ne
rect 5481 1384 5490 1418
rect 5524 1445 5566 1446
rect 5524 1411 5529 1445
rect 5559 1411 5566 1445
rect 5524 1402 5566 1411
rect 5600 1445 5642 1454
rect 5600 1411 5607 1445
rect 5637 1411 5642 1445
rect 5600 1406 5642 1411
rect 5676 1418 5704 1478
tri 5749 1465 5771 1487 se
rect 5771 1480 5786 1488
tri 5771 1465 5786 1480 nw
tri 5743 1459 5749 1465 se
rect 5749 1459 5758 1465
rect 5462 1374 5490 1384
tri 5490 1374 5514 1398 sw
rect 5408 1304 5424 1352
rect 5462 1342 5504 1374
tri 5521 1366 5522 1367 sw
rect 5521 1342 5522 1366
tri 5524 1365 5561 1402 ne
rect 5561 1374 5566 1402
tri 5566 1374 5592 1400 sw
rect 5676 1384 5685 1418
rect 5676 1374 5704 1384
rect 5561 1365 5645 1374
tri 5561 1346 5580 1365 ne
rect 5580 1346 5645 1365
rect 5462 1320 5522 1342
rect 5644 1342 5645 1346
rect 5662 1342 5704 1374
rect 5644 1320 5704 1342
rect 5550 1304 5567 1318
rect 5599 1304 5616 1318
tri 5387 1268 5409 1290 se
rect 5409 1283 5424 1304
tri 5409 1268 5424 1283 nw
rect 5743 1283 5758 1459
tri 5758 1452 5771 1465 nw
rect 5844 1384 5859 1612
tri 5381 1262 5387 1268 se
rect 5387 1262 5396 1268
rect 5381 1246 5396 1262
tri 5396 1255 5409 1268 nw
rect 5550 1260 5567 1274
rect 5599 1260 5616 1274
tri 5743 1268 5758 1283 ne
tri 5758 1268 5780 1290 sw
rect 5381 1210 5396 1218
rect 5462 1246 5522 1260
rect 5477 1236 5522 1246
rect 5477 1218 5505 1236
tri 5381 1195 5396 1210 ne
tri 5396 1195 5418 1217 sw
rect 5462 1208 5505 1218
rect 5520 1232 5522 1236
rect 5644 1246 5704 1260
tri 5758 1255 5771 1268 ne
rect 5771 1262 5780 1268
tri 5780 1262 5786 1268 sw
rect 5644 1236 5689 1246
rect 5520 1208 5594 1232
rect 5462 1204 5594 1208
tri 5594 1204 5622 1232 sw
rect 5644 1222 5646 1236
tri 5644 1220 5646 1222 ne
rect 5658 1218 5689 1236
rect 5658 1208 5704 1218
rect 5771 1247 5786 1262
tri 5396 1183 5408 1195 ne
rect 5408 1190 5418 1195
tri 5418 1190 5423 1195 sw
rect 5307 844 5322 1072
rect 5408 1034 5423 1190
rect 5462 1148 5490 1204
tri 5582 1186 5600 1204 ne
rect 5600 1184 5622 1204
tri 5622 1184 5642 1204 sw
tri 5658 1190 5676 1208 ne
rect 5481 1114 5490 1148
rect 5524 1175 5566 1176
rect 5524 1141 5529 1175
rect 5559 1141 5566 1175
rect 5524 1132 5566 1141
rect 5600 1175 5642 1184
rect 5600 1141 5607 1175
rect 5637 1141 5642 1175
rect 5600 1136 5642 1141
rect 5676 1148 5704 1208
tri 5749 1195 5771 1217 se
rect 5771 1210 5786 1218
tri 5771 1195 5786 1210 nw
tri 5743 1189 5749 1195 se
rect 5749 1189 5758 1195
rect 5462 1104 5490 1114
tri 5490 1104 5514 1128 sw
rect 5462 1072 5504 1104
tri 5521 1096 5522 1097 sw
rect 5521 1072 5522 1096
tri 5524 1095 5561 1132 ne
rect 5561 1104 5566 1132
tri 5566 1104 5592 1130 sw
rect 5676 1114 5685 1148
rect 5676 1104 5704 1114
rect 5561 1095 5645 1104
tri 5561 1076 5580 1095 ne
rect 5580 1076 5645 1095
rect 5462 1050 5522 1072
rect 5644 1072 5645 1076
rect 5662 1072 5704 1104
rect 5644 1050 5704 1072
rect 5550 1034 5567 1048
rect 5599 1034 5616 1048
tri 5387 998 5409 1020 se
rect 5409 1013 5424 1034
tri 5409 998 5424 1013 nw
rect 5743 1013 5758 1189
tri 5758 1182 5771 1195 nw
rect 5844 1114 5859 1342
tri 5381 992 5387 998 se
rect 5387 992 5396 998
rect 5381 976 5396 992
tri 5396 985 5409 998 nw
rect 5550 990 5567 1004
rect 5599 990 5616 1004
tri 5743 998 5758 1013 ne
tri 5758 998 5780 1020 sw
rect 5381 940 5396 948
rect 5462 976 5522 990
rect 5477 966 5522 976
rect 5477 948 5505 966
tri 5381 925 5396 940 ne
tri 5396 925 5418 947 sw
rect 5462 938 5505 948
rect 5520 962 5522 966
rect 5644 976 5704 990
tri 5758 985 5771 998 ne
rect 5771 992 5780 998
tri 5780 992 5786 998 sw
rect 5644 966 5689 976
rect 5520 938 5594 962
rect 5462 934 5594 938
tri 5594 934 5622 962 sw
rect 5644 952 5646 966
tri 5644 950 5646 952 ne
rect 5658 948 5689 966
rect 5658 938 5704 948
rect 5771 977 5786 992
tri 5396 913 5408 925 ne
rect 5408 920 5418 925
tri 5418 920 5423 925 sw
rect 5307 574 5322 802
rect 5408 812 5423 920
rect 5462 878 5490 934
tri 5582 916 5600 934 ne
rect 5600 914 5622 934
tri 5622 914 5642 934 sw
tri 5658 920 5676 938 ne
rect 5481 844 5490 878
rect 5524 905 5566 906
rect 5524 871 5529 905
rect 5559 871 5566 905
rect 5524 862 5566 871
rect 5600 905 5642 914
rect 5600 871 5607 905
rect 5637 871 5642 905
rect 5600 866 5642 871
rect 5676 878 5704 938
tri 5749 925 5771 947 se
rect 5771 940 5786 948
tri 5771 925 5786 940 nw
tri 5743 919 5749 925 se
rect 5749 919 5758 925
rect 5462 834 5490 844
tri 5490 834 5514 858 sw
rect 5408 764 5424 812
rect 5462 802 5504 834
tri 5521 826 5522 827 sw
rect 5521 802 5522 826
tri 5524 825 5561 862 ne
rect 5561 834 5566 862
tri 5566 834 5592 860 sw
rect 5676 844 5685 878
rect 5676 834 5704 844
rect 5561 825 5645 834
tri 5561 806 5580 825 ne
rect 5580 806 5645 825
rect 5462 780 5522 802
rect 5644 802 5645 806
rect 5662 802 5704 834
rect 5644 780 5704 802
rect 5550 764 5567 778
rect 5599 764 5616 778
tri 5387 728 5409 750 se
rect 5409 743 5424 764
tri 5409 728 5424 743 nw
rect 5743 743 5758 919
tri 5758 912 5771 925 nw
rect 5844 844 5859 1072
tri 5381 722 5387 728 se
rect 5387 722 5396 728
rect 5381 706 5396 722
tri 5396 715 5409 728 nw
rect 5550 720 5567 734
rect 5599 720 5616 734
tri 5743 728 5758 743 ne
tri 5758 728 5780 750 sw
rect 5381 670 5396 678
rect 5462 706 5522 720
rect 5477 696 5522 706
rect 5477 678 5505 696
tri 5381 655 5396 670 ne
tri 5396 655 5418 677 sw
rect 5462 668 5505 678
rect 5520 692 5522 696
rect 5644 706 5704 720
tri 5758 715 5771 728 ne
rect 5771 722 5780 728
tri 5780 722 5786 728 sw
rect 5644 696 5689 706
rect 5520 668 5594 692
rect 5462 664 5594 668
tri 5594 664 5622 692 sw
rect 5644 682 5646 696
tri 5644 680 5646 682 ne
rect 5658 678 5689 696
rect 5658 668 5704 678
rect 5771 707 5786 722
tri 5396 643 5408 655 ne
rect 5408 650 5418 655
tri 5418 650 5423 655 sw
rect 5307 304 5322 532
rect 5408 494 5423 650
rect 5462 608 5490 664
tri 5582 646 5600 664 ne
rect 5600 644 5622 664
tri 5622 644 5642 664 sw
tri 5658 650 5676 668 ne
rect 5481 574 5490 608
rect 5524 635 5566 636
rect 5524 601 5529 635
rect 5559 601 5566 635
rect 5524 592 5566 601
rect 5600 635 5642 644
rect 5600 601 5607 635
rect 5637 601 5642 635
rect 5600 596 5642 601
rect 5676 608 5704 668
tri 5749 655 5771 677 se
rect 5771 670 5786 678
tri 5771 655 5786 670 nw
tri 5743 649 5749 655 se
rect 5749 649 5758 655
rect 5462 564 5490 574
tri 5490 564 5514 588 sw
rect 5462 532 5504 564
tri 5521 556 5522 557 sw
rect 5521 532 5522 556
tri 5524 555 5561 592 ne
rect 5561 564 5566 592
tri 5566 564 5592 590 sw
rect 5676 574 5685 608
rect 5676 564 5704 574
rect 5561 555 5645 564
tri 5561 536 5580 555 ne
rect 5580 536 5645 555
rect 5462 510 5522 532
rect 5644 532 5645 536
rect 5662 532 5704 564
rect 5644 510 5704 532
rect 5550 494 5567 508
rect 5599 494 5616 508
tri 5387 458 5409 480 se
rect 5409 473 5424 494
tri 5409 458 5424 473 nw
rect 5743 473 5758 649
tri 5758 642 5771 655 nw
rect 5844 574 5859 802
tri 5381 452 5387 458 se
rect 5387 452 5396 458
rect 5381 436 5396 452
tri 5396 445 5409 458 nw
rect 5550 450 5567 464
rect 5599 450 5616 464
tri 5743 458 5758 473 ne
tri 5758 458 5780 480 sw
rect 5381 400 5396 408
rect 5462 436 5522 450
rect 5477 426 5522 436
rect 5477 408 5505 426
tri 5381 385 5396 400 ne
tri 5396 385 5418 407 sw
rect 5462 398 5505 408
rect 5520 422 5522 426
rect 5644 436 5704 450
tri 5758 445 5771 458 ne
rect 5771 452 5780 458
tri 5780 452 5786 458 sw
rect 5644 426 5689 436
rect 5520 398 5594 422
rect 5462 394 5594 398
tri 5594 394 5622 422 sw
rect 5644 412 5646 426
tri 5644 410 5646 412 ne
rect 5658 408 5689 426
rect 5658 398 5704 408
rect 5771 437 5786 452
tri 5396 373 5408 385 ne
rect 5408 380 5418 385
tri 5418 380 5423 385 sw
rect 5307 34 5322 262
rect 5408 272 5423 380
rect 5462 338 5490 394
tri 5582 376 5600 394 ne
rect 5600 374 5622 394
tri 5622 374 5642 394 sw
tri 5658 380 5676 398 ne
rect 5481 304 5490 338
rect 5524 365 5566 366
rect 5524 331 5529 365
rect 5559 331 5566 365
rect 5524 322 5566 331
rect 5600 365 5642 374
rect 5600 331 5607 365
rect 5637 331 5642 365
rect 5600 326 5642 331
rect 5676 338 5704 398
tri 5749 385 5771 407 se
rect 5771 400 5786 408
tri 5771 385 5786 400 nw
tri 5743 379 5749 385 se
rect 5749 379 5758 385
rect 5462 294 5490 304
tri 5490 294 5514 318 sw
rect 5408 224 5424 272
rect 5462 262 5504 294
tri 5521 286 5522 287 sw
rect 5521 262 5522 286
tri 5524 285 5561 322 ne
rect 5561 294 5566 322
tri 5566 294 5592 320 sw
rect 5676 304 5685 338
rect 5676 294 5704 304
rect 5561 285 5645 294
tri 5561 266 5580 285 ne
rect 5580 266 5645 285
rect 5462 240 5522 262
rect 5644 262 5645 266
rect 5662 262 5704 294
rect 5644 240 5704 262
rect 5550 224 5567 238
rect 5599 224 5616 238
tri 5387 188 5409 210 se
rect 5409 203 5424 224
tri 5409 188 5424 203 nw
rect 5743 203 5758 379
tri 5758 372 5771 385 nw
rect 5844 304 5859 532
tri 5381 182 5387 188 se
rect 5387 182 5396 188
rect 5381 166 5396 182
tri 5396 175 5409 188 nw
rect 5550 180 5567 194
rect 5599 180 5616 194
tri 5743 188 5758 203 ne
tri 5758 188 5780 210 sw
rect 5381 130 5396 138
rect 5462 166 5522 180
rect 5477 156 5522 166
rect 5477 138 5505 156
tri 5381 115 5396 130 ne
tri 5396 115 5418 137 sw
rect 5462 128 5505 138
rect 5520 152 5522 156
rect 5644 166 5704 180
tri 5758 175 5771 188 ne
rect 5771 182 5780 188
tri 5780 182 5786 188 sw
rect 5644 156 5689 166
rect 5520 128 5594 152
rect 5462 124 5594 128
tri 5594 124 5622 152 sw
rect 5644 142 5646 156
tri 5644 140 5646 142 ne
rect 5658 138 5689 156
rect 5658 128 5704 138
rect 5771 167 5786 182
tri 5396 103 5408 115 ne
rect 5408 110 5418 115
tri 5418 110 5423 115 sw
rect 5307 -236 5322 -8
rect 5408 -46 5423 110
rect 5462 68 5490 124
tri 5582 106 5600 124 ne
rect 5600 104 5622 124
tri 5622 104 5642 124 sw
tri 5658 110 5676 128 ne
rect 5481 34 5490 68
rect 5524 95 5566 96
rect 5524 61 5529 95
rect 5559 61 5566 95
rect 5524 52 5566 61
rect 5600 95 5642 104
rect 5600 61 5607 95
rect 5637 61 5642 95
rect 5600 56 5642 61
rect 5676 68 5704 128
tri 5749 115 5771 137 se
rect 5771 130 5786 138
tri 5771 115 5786 130 nw
tri 5743 109 5749 115 se
rect 5749 109 5758 115
rect 5462 24 5490 34
tri 5490 24 5514 48 sw
rect 5462 -8 5504 24
tri 5521 16 5522 17 sw
rect 5521 -8 5522 16
tri 5524 15 5561 52 ne
rect 5561 24 5566 52
tri 5566 24 5592 50 sw
rect 5676 34 5685 68
rect 5676 24 5704 34
rect 5561 15 5645 24
tri 5561 -4 5580 15 ne
rect 5580 -4 5645 15
rect 5462 -30 5522 -8
rect 5644 -8 5645 -4
rect 5662 -8 5704 24
rect 5644 -30 5704 -8
rect 5550 -46 5567 -32
rect 5599 -46 5616 -32
tri 5387 -82 5409 -60 se
rect 5409 -67 5424 -46
tri 5409 -82 5424 -67 nw
rect 5743 -67 5758 109
tri 5758 102 5771 115 nw
rect 5844 34 5859 262
tri 5381 -88 5387 -82 se
rect 5387 -88 5396 -82
rect 5381 -104 5396 -88
tri 5396 -95 5409 -82 nw
rect 5550 -90 5567 -76
rect 5599 -90 5616 -76
tri 5743 -82 5758 -67 ne
tri 5758 -82 5780 -60 sw
rect 5381 -140 5396 -132
rect 5462 -104 5522 -90
rect 5477 -114 5522 -104
rect 5477 -132 5505 -114
tri 5381 -155 5396 -140 ne
tri 5396 -155 5418 -133 sw
rect 5462 -142 5505 -132
rect 5520 -118 5522 -114
rect 5644 -104 5704 -90
tri 5758 -95 5771 -82 ne
rect 5771 -88 5780 -82
tri 5780 -88 5786 -82 sw
rect 5644 -114 5689 -104
rect 5520 -142 5594 -118
rect 5462 -146 5594 -142
tri 5594 -146 5622 -118 sw
rect 5644 -128 5646 -114
tri 5644 -130 5646 -128 ne
rect 5658 -132 5689 -114
rect 5658 -142 5704 -132
rect 5771 -103 5786 -88
tri 5396 -167 5408 -155 ne
rect 5408 -160 5418 -155
tri 5418 -160 5423 -155 sw
rect 5307 -506 5322 -278
rect 5408 -268 5423 -160
rect 5462 -202 5490 -146
tri 5582 -164 5600 -146 ne
rect 5600 -166 5622 -146
tri 5622 -166 5642 -146 sw
tri 5658 -160 5676 -142 ne
rect 5481 -236 5490 -202
rect 5524 -175 5566 -174
rect 5524 -209 5529 -175
rect 5559 -209 5566 -175
rect 5524 -218 5566 -209
rect 5600 -175 5642 -166
rect 5600 -209 5607 -175
rect 5637 -209 5642 -175
rect 5600 -214 5642 -209
rect 5676 -202 5704 -142
tri 5749 -155 5771 -133 se
rect 5771 -140 5786 -132
tri 5771 -155 5786 -140 nw
tri 5743 -161 5749 -155 se
rect 5749 -161 5758 -155
rect 5462 -246 5490 -236
tri 5490 -246 5514 -222 sw
rect 5408 -316 5424 -268
rect 5462 -278 5504 -246
tri 5521 -254 5522 -253 sw
rect 5521 -278 5522 -254
tri 5524 -255 5561 -218 ne
rect 5561 -246 5566 -218
tri 5566 -246 5592 -220 sw
rect 5676 -236 5685 -202
rect 5676 -246 5704 -236
rect 5561 -255 5645 -246
tri 5561 -274 5580 -255 ne
rect 5580 -274 5645 -255
rect 5462 -300 5522 -278
rect 5644 -278 5645 -274
rect 5662 -278 5704 -246
rect 5644 -300 5704 -278
rect 5550 -316 5567 -302
rect 5599 -316 5616 -302
tri 5387 -352 5409 -330 se
rect 5409 -337 5424 -316
tri 5409 -352 5424 -337 nw
rect 5743 -337 5758 -161
tri 5758 -168 5771 -155 nw
rect 5844 -236 5859 -8
tri 5381 -358 5387 -352 se
rect 5387 -358 5396 -352
rect 5381 -374 5396 -358
tri 5396 -365 5409 -352 nw
rect 5550 -360 5567 -346
rect 5599 -360 5616 -346
tri 5743 -352 5758 -337 ne
tri 5758 -352 5780 -330 sw
rect 5381 -410 5396 -402
rect 5462 -374 5522 -360
rect 5477 -384 5522 -374
rect 5477 -402 5505 -384
tri 5381 -425 5396 -410 ne
tri 5396 -425 5418 -403 sw
rect 5462 -412 5505 -402
rect 5520 -388 5522 -384
rect 5644 -374 5704 -360
tri 5758 -365 5771 -352 ne
rect 5771 -358 5780 -352
tri 5780 -358 5786 -352 sw
rect 5644 -384 5689 -374
rect 5520 -412 5594 -388
rect 5462 -416 5594 -412
tri 5594 -416 5622 -388 sw
rect 5644 -398 5646 -384
tri 5644 -400 5646 -398 ne
rect 5658 -402 5689 -384
rect 5658 -412 5704 -402
rect 5771 -373 5786 -358
tri 5396 -437 5408 -425 ne
rect 5408 -430 5418 -425
tri 5418 -430 5423 -425 sw
rect 5307 -776 5322 -548
rect 5408 -586 5423 -430
rect 5462 -472 5490 -416
tri 5582 -434 5600 -416 ne
rect 5600 -436 5622 -416
tri 5622 -436 5642 -416 sw
tri 5658 -430 5676 -412 ne
rect 5481 -506 5490 -472
rect 5524 -445 5566 -444
rect 5524 -479 5529 -445
rect 5559 -479 5566 -445
rect 5524 -488 5566 -479
rect 5600 -445 5642 -436
rect 5600 -479 5607 -445
rect 5637 -479 5642 -445
rect 5600 -484 5642 -479
rect 5676 -472 5704 -412
tri 5749 -425 5771 -403 se
rect 5771 -410 5786 -402
tri 5771 -425 5786 -410 nw
tri 5743 -431 5749 -425 se
rect 5749 -431 5758 -425
rect 5462 -516 5490 -506
tri 5490 -516 5514 -492 sw
rect 5462 -548 5504 -516
tri 5521 -524 5522 -523 sw
rect 5521 -548 5522 -524
tri 5524 -525 5561 -488 ne
rect 5561 -516 5566 -488
tri 5566 -516 5592 -490 sw
rect 5676 -506 5685 -472
rect 5676 -516 5704 -506
rect 5561 -525 5645 -516
tri 5561 -544 5580 -525 ne
rect 5580 -544 5645 -525
rect 5462 -570 5522 -548
rect 5644 -548 5645 -544
rect 5662 -548 5704 -516
rect 5644 -570 5704 -548
rect 5550 -586 5567 -572
rect 5599 -586 5616 -572
tri 5387 -622 5409 -600 se
rect 5409 -607 5424 -586
tri 5409 -622 5424 -607 nw
rect 5743 -607 5758 -431
tri 5758 -438 5771 -425 nw
rect 5844 -506 5859 -278
tri 5381 -628 5387 -622 se
rect 5387 -628 5396 -622
rect 5381 -644 5396 -628
tri 5396 -635 5409 -622 nw
rect 5550 -630 5567 -616
rect 5599 -630 5616 -616
tri 5743 -622 5758 -607 ne
tri 5758 -622 5780 -600 sw
rect 5381 -680 5396 -672
rect 5462 -644 5522 -630
rect 5477 -654 5522 -644
rect 5477 -672 5505 -654
tri 5381 -695 5396 -680 ne
tri 5396 -695 5418 -673 sw
rect 5462 -682 5505 -672
rect 5520 -658 5522 -654
rect 5644 -644 5704 -630
tri 5758 -635 5771 -622 ne
rect 5771 -628 5780 -622
tri 5780 -628 5786 -622 sw
rect 5644 -654 5689 -644
rect 5520 -682 5594 -658
rect 5462 -686 5594 -682
tri 5594 -686 5622 -658 sw
rect 5644 -668 5646 -654
tri 5644 -670 5646 -668 ne
rect 5658 -672 5689 -654
rect 5658 -682 5704 -672
rect 5771 -643 5786 -628
tri 5396 -707 5408 -695 ne
rect 5408 -700 5418 -695
tri 5418 -700 5423 -695 sw
rect 5307 -1046 5322 -818
rect 5408 -808 5423 -700
rect 5462 -742 5490 -686
tri 5582 -704 5600 -686 ne
rect 5600 -706 5622 -686
tri 5622 -706 5642 -686 sw
tri 5658 -700 5676 -682 ne
rect 5481 -776 5490 -742
rect 5524 -715 5566 -714
rect 5524 -749 5529 -715
rect 5559 -749 5566 -715
rect 5524 -758 5566 -749
rect 5600 -715 5642 -706
rect 5600 -749 5607 -715
rect 5637 -749 5642 -715
rect 5600 -754 5642 -749
rect 5676 -742 5704 -682
tri 5749 -695 5771 -673 se
rect 5771 -680 5786 -672
tri 5771 -695 5786 -680 nw
tri 5743 -701 5749 -695 se
rect 5749 -701 5758 -695
rect 5462 -786 5490 -776
tri 5490 -786 5514 -762 sw
rect 5408 -856 5424 -808
rect 5462 -818 5504 -786
tri 5521 -794 5522 -793 sw
rect 5521 -818 5522 -794
tri 5524 -795 5561 -758 ne
rect 5561 -786 5566 -758
tri 5566 -786 5592 -760 sw
rect 5676 -776 5685 -742
rect 5676 -786 5704 -776
rect 5561 -795 5645 -786
tri 5561 -814 5580 -795 ne
rect 5580 -814 5645 -795
rect 5462 -840 5522 -818
rect 5644 -818 5645 -814
rect 5662 -818 5704 -786
rect 5644 -840 5704 -818
rect 5550 -856 5567 -842
rect 5599 -856 5616 -842
tri 5387 -892 5409 -870 se
rect 5409 -877 5424 -856
tri 5409 -892 5424 -877 nw
rect 5743 -877 5758 -701
tri 5758 -708 5771 -695 nw
rect 5844 -776 5859 -548
tri 5381 -898 5387 -892 se
rect 5387 -898 5396 -892
rect 5381 -914 5396 -898
tri 5396 -905 5409 -892 nw
rect 5550 -900 5567 -886
rect 5599 -900 5616 -886
tri 5743 -892 5758 -877 ne
tri 5758 -892 5780 -870 sw
rect 5381 -950 5396 -942
rect 5462 -914 5522 -900
rect 5477 -924 5522 -914
rect 5477 -942 5505 -924
tri 5381 -965 5396 -950 ne
tri 5396 -965 5418 -943 sw
rect 5462 -952 5505 -942
rect 5520 -928 5522 -924
rect 5644 -914 5704 -900
tri 5758 -905 5771 -892 ne
rect 5771 -898 5780 -892
tri 5780 -898 5786 -892 sw
rect 5644 -924 5689 -914
rect 5520 -952 5594 -928
rect 5462 -956 5594 -952
tri 5594 -956 5622 -928 sw
rect 5644 -938 5646 -924
tri 5644 -940 5646 -938 ne
rect 5658 -942 5689 -924
rect 5658 -952 5704 -942
rect 5771 -913 5786 -898
tri 5396 -977 5408 -965 ne
rect 5408 -970 5418 -965
tri 5418 -970 5423 -965 sw
rect 5307 -1316 5322 -1088
rect 5408 -1126 5423 -970
rect 5462 -1012 5490 -956
tri 5582 -974 5600 -956 ne
rect 5600 -976 5622 -956
tri 5622 -976 5642 -956 sw
tri 5658 -970 5676 -952 ne
rect 5481 -1046 5490 -1012
rect 5524 -985 5566 -984
rect 5524 -1019 5529 -985
rect 5559 -1019 5566 -985
rect 5524 -1028 5566 -1019
rect 5600 -985 5642 -976
rect 5600 -1019 5607 -985
rect 5637 -1019 5642 -985
rect 5600 -1024 5642 -1019
rect 5676 -1012 5704 -952
tri 5749 -965 5771 -943 se
rect 5771 -950 5786 -942
tri 5771 -965 5786 -950 nw
tri 5743 -971 5749 -965 se
rect 5749 -971 5758 -965
rect 5462 -1056 5490 -1046
tri 5490 -1056 5514 -1032 sw
rect 5462 -1088 5504 -1056
tri 5521 -1064 5522 -1063 sw
rect 5521 -1088 5522 -1064
tri 5524 -1065 5561 -1028 ne
rect 5561 -1056 5566 -1028
tri 5566 -1056 5592 -1030 sw
rect 5676 -1046 5685 -1012
rect 5676 -1056 5704 -1046
rect 5561 -1065 5645 -1056
tri 5561 -1084 5580 -1065 ne
rect 5580 -1084 5645 -1065
rect 5462 -1110 5522 -1088
rect 5644 -1088 5645 -1084
rect 5662 -1088 5704 -1056
rect 5644 -1110 5704 -1088
rect 5550 -1126 5567 -1112
rect 5599 -1126 5616 -1112
tri 5387 -1162 5409 -1140 se
rect 5409 -1147 5424 -1126
tri 5409 -1162 5424 -1147 nw
rect 5743 -1147 5758 -971
tri 5758 -978 5771 -965 nw
rect 5844 -1046 5859 -818
tri 5381 -1168 5387 -1162 se
rect 5387 -1168 5396 -1162
rect 5381 -1184 5396 -1168
tri 5396 -1175 5409 -1162 nw
rect 5550 -1170 5567 -1156
rect 5599 -1170 5616 -1156
tri 5743 -1162 5758 -1147 ne
tri 5758 -1162 5780 -1140 sw
rect 5381 -1220 5396 -1212
rect 5462 -1184 5522 -1170
rect 5477 -1194 5522 -1184
rect 5477 -1212 5505 -1194
tri 5381 -1235 5396 -1220 ne
tri 5396 -1235 5418 -1213 sw
rect 5462 -1222 5505 -1212
rect 5520 -1198 5522 -1194
rect 5644 -1184 5704 -1170
tri 5758 -1175 5771 -1162 ne
rect 5771 -1168 5780 -1162
tri 5780 -1168 5786 -1162 sw
rect 5644 -1194 5689 -1184
rect 5520 -1222 5594 -1198
rect 5462 -1226 5594 -1222
tri 5594 -1226 5622 -1198 sw
rect 5644 -1208 5646 -1194
tri 5644 -1210 5646 -1208 ne
rect 5658 -1212 5689 -1194
rect 5658 -1222 5704 -1212
rect 5771 -1183 5786 -1168
tri 5396 -1247 5408 -1235 ne
rect 5408 -1240 5418 -1235
tri 5418 -1240 5423 -1235 sw
rect 5307 -1586 5322 -1358
rect 5408 -1348 5423 -1240
rect 5462 -1282 5490 -1226
tri 5582 -1244 5600 -1226 ne
rect 5600 -1246 5622 -1226
tri 5622 -1246 5642 -1226 sw
tri 5658 -1240 5676 -1222 ne
rect 5481 -1316 5490 -1282
rect 5524 -1255 5566 -1254
rect 5524 -1289 5529 -1255
rect 5559 -1289 5566 -1255
rect 5524 -1298 5566 -1289
rect 5600 -1255 5642 -1246
rect 5600 -1289 5607 -1255
rect 5637 -1289 5642 -1255
rect 5600 -1294 5642 -1289
rect 5676 -1282 5704 -1222
tri 5749 -1235 5771 -1213 se
rect 5771 -1220 5786 -1212
tri 5771 -1235 5786 -1220 nw
tri 5743 -1241 5749 -1235 se
rect 5749 -1241 5758 -1235
rect 5462 -1326 5490 -1316
tri 5490 -1326 5514 -1302 sw
rect 5408 -1396 5424 -1348
rect 5462 -1358 5504 -1326
tri 5521 -1334 5522 -1333 sw
rect 5521 -1358 5522 -1334
tri 5524 -1335 5561 -1298 ne
rect 5561 -1326 5566 -1298
tri 5566 -1326 5592 -1300 sw
rect 5676 -1316 5685 -1282
rect 5676 -1326 5704 -1316
rect 5561 -1335 5645 -1326
tri 5561 -1354 5580 -1335 ne
rect 5580 -1354 5645 -1335
rect 5462 -1380 5522 -1358
rect 5644 -1358 5645 -1354
rect 5662 -1358 5704 -1326
rect 5644 -1380 5704 -1358
rect 5550 -1396 5567 -1382
rect 5599 -1396 5616 -1382
tri 5387 -1432 5409 -1410 se
rect 5409 -1417 5424 -1396
tri 5409 -1432 5424 -1417 nw
rect 5743 -1417 5758 -1241
tri 5758 -1248 5771 -1235 nw
rect 5844 -1316 5859 -1088
tri 5381 -1438 5387 -1432 se
rect 5387 -1438 5396 -1432
rect 5381 -1454 5396 -1438
tri 5396 -1445 5409 -1432 nw
rect 5550 -1440 5567 -1426
rect 5599 -1440 5616 -1426
tri 5743 -1432 5758 -1417 ne
tri 5758 -1432 5780 -1410 sw
rect 5381 -1490 5396 -1482
rect 5462 -1454 5522 -1440
rect 5477 -1464 5522 -1454
rect 5477 -1482 5505 -1464
tri 5381 -1505 5396 -1490 ne
tri 5396 -1505 5418 -1483 sw
rect 5462 -1492 5505 -1482
rect 5520 -1468 5522 -1464
rect 5644 -1454 5704 -1440
tri 5758 -1445 5771 -1432 ne
rect 5771 -1438 5780 -1432
tri 5780 -1438 5786 -1432 sw
rect 5644 -1464 5689 -1454
rect 5520 -1492 5594 -1468
rect 5462 -1496 5594 -1492
tri 5594 -1496 5622 -1468 sw
rect 5644 -1478 5646 -1464
tri 5644 -1480 5646 -1478 ne
rect 5658 -1482 5689 -1464
rect 5658 -1492 5704 -1482
rect 5771 -1453 5786 -1438
tri 5396 -1517 5408 -1505 ne
rect 5408 -1510 5418 -1505
tri 5418 -1510 5423 -1505 sw
rect 5307 -1856 5322 -1628
rect 5408 -1666 5423 -1510
rect 5462 -1552 5490 -1496
tri 5582 -1514 5600 -1496 ne
rect 5600 -1516 5622 -1496
tri 5622 -1516 5642 -1496 sw
tri 5658 -1510 5676 -1492 ne
rect 5481 -1586 5490 -1552
rect 5524 -1525 5566 -1524
rect 5524 -1559 5529 -1525
rect 5559 -1559 5566 -1525
rect 5524 -1568 5566 -1559
rect 5600 -1525 5642 -1516
rect 5600 -1559 5607 -1525
rect 5637 -1559 5642 -1525
rect 5600 -1564 5642 -1559
rect 5676 -1552 5704 -1492
tri 5749 -1505 5771 -1483 se
rect 5771 -1490 5786 -1482
tri 5771 -1505 5786 -1490 nw
tri 5743 -1511 5749 -1505 se
rect 5749 -1511 5758 -1505
rect 5462 -1596 5490 -1586
tri 5490 -1596 5514 -1572 sw
rect 5462 -1628 5504 -1596
tri 5521 -1604 5522 -1603 sw
rect 5521 -1628 5522 -1604
tri 5524 -1605 5561 -1568 ne
rect 5561 -1596 5566 -1568
tri 5566 -1596 5592 -1570 sw
rect 5676 -1586 5685 -1552
rect 5676 -1596 5704 -1586
rect 5561 -1605 5645 -1596
tri 5561 -1624 5580 -1605 ne
rect 5580 -1624 5645 -1605
rect 5462 -1650 5522 -1628
rect 5644 -1628 5645 -1624
rect 5662 -1628 5704 -1596
rect 5644 -1650 5704 -1628
rect 5550 -1666 5567 -1652
rect 5599 -1666 5616 -1652
tri 5387 -1702 5409 -1680 se
rect 5409 -1687 5424 -1666
tri 5409 -1702 5424 -1687 nw
rect 5743 -1687 5758 -1511
tri 5758 -1518 5771 -1505 nw
rect 5844 -1586 5859 -1358
tri 5381 -1708 5387 -1702 se
rect 5387 -1708 5396 -1702
rect 5381 -1724 5396 -1708
tri 5396 -1715 5409 -1702 nw
rect 5550 -1710 5567 -1696
rect 5599 -1710 5616 -1696
tri 5743 -1702 5758 -1687 ne
tri 5758 -1702 5780 -1680 sw
rect 5381 -1760 5396 -1752
rect 5462 -1724 5522 -1710
rect 5477 -1734 5522 -1724
rect 5477 -1752 5505 -1734
tri 5381 -1775 5396 -1760 ne
tri 5396 -1775 5418 -1753 sw
rect 5462 -1762 5505 -1752
rect 5520 -1738 5522 -1734
rect 5644 -1724 5704 -1710
tri 5758 -1715 5771 -1702 ne
rect 5771 -1708 5780 -1702
tri 5780 -1708 5786 -1702 sw
rect 5644 -1734 5689 -1724
rect 5520 -1762 5594 -1738
rect 5462 -1766 5594 -1762
tri 5594 -1766 5622 -1738 sw
rect 5644 -1748 5646 -1734
tri 5644 -1750 5646 -1748 ne
rect 5658 -1752 5689 -1734
rect 5658 -1762 5704 -1752
rect 5771 -1723 5786 -1708
tri 5396 -1787 5408 -1775 ne
rect 5408 -1780 5418 -1775
tri 5418 -1780 5423 -1775 sw
rect 5307 -2126 5322 -1898
rect 5408 -1888 5423 -1780
rect 5462 -1822 5490 -1766
tri 5582 -1784 5600 -1766 ne
rect 5600 -1786 5622 -1766
tri 5622 -1786 5642 -1766 sw
tri 5658 -1780 5676 -1762 ne
rect 5481 -1856 5490 -1822
rect 5524 -1795 5566 -1794
rect 5524 -1829 5529 -1795
rect 5559 -1829 5566 -1795
rect 5524 -1838 5566 -1829
rect 5600 -1795 5642 -1786
rect 5600 -1829 5607 -1795
rect 5637 -1829 5642 -1795
rect 5600 -1834 5642 -1829
rect 5676 -1822 5704 -1762
tri 5749 -1775 5771 -1753 se
rect 5771 -1760 5786 -1752
tri 5771 -1775 5786 -1760 nw
tri 5743 -1781 5749 -1775 se
rect 5749 -1781 5758 -1775
rect 5462 -1866 5490 -1856
tri 5490 -1866 5514 -1842 sw
rect 5408 -1936 5424 -1888
rect 5462 -1898 5504 -1866
tri 5521 -1874 5522 -1873 sw
rect 5521 -1898 5522 -1874
tri 5524 -1875 5561 -1838 ne
rect 5561 -1866 5566 -1838
tri 5566 -1866 5592 -1840 sw
rect 5676 -1856 5685 -1822
rect 5676 -1866 5704 -1856
rect 5561 -1875 5645 -1866
tri 5561 -1894 5580 -1875 ne
rect 5580 -1894 5645 -1875
rect 5462 -1920 5522 -1898
rect 5644 -1898 5645 -1894
rect 5662 -1898 5704 -1866
rect 5644 -1920 5704 -1898
rect 5550 -1936 5567 -1922
rect 5599 -1936 5616 -1922
tri 5387 -1972 5409 -1950 se
rect 5409 -1957 5424 -1936
tri 5409 -1972 5424 -1957 nw
rect 5743 -1957 5758 -1781
tri 5758 -1788 5771 -1775 nw
rect 5844 -1856 5859 -1628
tri 5381 -1978 5387 -1972 se
rect 5387 -1978 5396 -1972
rect 5381 -1994 5396 -1978
tri 5396 -1985 5409 -1972 nw
rect 5550 -1980 5567 -1966
rect 5599 -1980 5616 -1966
tri 5743 -1972 5758 -1957 ne
tri 5758 -1972 5780 -1950 sw
rect 5381 -2030 5396 -2022
rect 5462 -1994 5522 -1980
rect 5477 -2004 5522 -1994
rect 5477 -2022 5505 -2004
tri 5381 -2045 5396 -2030 ne
tri 5396 -2045 5418 -2023 sw
rect 5462 -2032 5505 -2022
rect 5520 -2008 5522 -2004
rect 5644 -1994 5704 -1980
tri 5758 -1985 5771 -1972 ne
rect 5771 -1978 5780 -1972
tri 5780 -1978 5786 -1972 sw
rect 5644 -2004 5689 -1994
rect 5520 -2032 5594 -2008
rect 5462 -2036 5594 -2032
tri 5594 -2036 5622 -2008 sw
rect 5644 -2018 5646 -2004
tri 5644 -2020 5646 -2018 ne
rect 5658 -2022 5689 -2004
rect 5658 -2032 5704 -2022
rect 5771 -1993 5786 -1978
tri 5396 -2057 5408 -2045 ne
rect 5408 -2050 5418 -2045
tri 5418 -2050 5423 -2045 sw
rect 5307 -2396 5322 -2168
rect 5408 -2206 5423 -2050
rect 5462 -2092 5490 -2036
tri 5582 -2054 5600 -2036 ne
rect 5600 -2056 5622 -2036
tri 5622 -2056 5642 -2036 sw
tri 5658 -2050 5676 -2032 ne
rect 5481 -2126 5490 -2092
rect 5524 -2065 5566 -2064
rect 5524 -2099 5529 -2065
rect 5559 -2099 5566 -2065
rect 5524 -2108 5566 -2099
rect 5600 -2065 5642 -2056
rect 5600 -2099 5607 -2065
rect 5637 -2099 5642 -2065
rect 5600 -2104 5642 -2099
rect 5676 -2092 5704 -2032
tri 5749 -2045 5771 -2023 se
rect 5771 -2030 5786 -2022
tri 5771 -2045 5786 -2030 nw
tri 5743 -2051 5749 -2045 se
rect 5749 -2051 5758 -2045
rect 5462 -2136 5490 -2126
tri 5490 -2136 5514 -2112 sw
rect 5462 -2168 5504 -2136
tri 5521 -2144 5522 -2143 sw
rect 5521 -2168 5522 -2144
tri 5524 -2145 5561 -2108 ne
rect 5561 -2136 5566 -2108
tri 5566 -2136 5592 -2110 sw
rect 5676 -2126 5685 -2092
rect 5676 -2136 5704 -2126
rect 5561 -2145 5645 -2136
tri 5561 -2164 5580 -2145 ne
rect 5580 -2164 5645 -2145
rect 5462 -2190 5522 -2168
rect 5644 -2168 5645 -2164
rect 5662 -2168 5704 -2136
rect 5644 -2190 5704 -2168
rect 5550 -2206 5567 -2192
rect 5599 -2206 5616 -2192
tri 5387 -2242 5409 -2220 se
rect 5409 -2227 5424 -2206
tri 5409 -2242 5424 -2227 nw
rect 5743 -2227 5758 -2051
tri 5758 -2058 5771 -2045 nw
rect 5844 -2126 5859 -1898
tri 5381 -2248 5387 -2242 se
rect 5387 -2248 5396 -2242
rect 5381 -2264 5396 -2248
tri 5396 -2255 5409 -2242 nw
rect 5550 -2250 5567 -2236
rect 5599 -2250 5616 -2236
tri 5743 -2242 5758 -2227 ne
tri 5758 -2242 5780 -2220 sw
rect 5381 -2300 5396 -2292
rect 5462 -2264 5522 -2250
rect 5477 -2274 5522 -2264
rect 5477 -2292 5505 -2274
tri 5381 -2315 5396 -2300 ne
tri 5396 -2315 5418 -2293 sw
rect 5462 -2302 5505 -2292
rect 5520 -2278 5522 -2274
rect 5644 -2264 5704 -2250
tri 5758 -2255 5771 -2242 ne
rect 5771 -2248 5780 -2242
tri 5780 -2248 5786 -2242 sw
rect 5644 -2274 5689 -2264
rect 5520 -2302 5594 -2278
rect 5462 -2306 5594 -2302
tri 5594 -2306 5622 -2278 sw
rect 5644 -2288 5646 -2274
tri 5644 -2290 5646 -2288 ne
rect 5658 -2292 5689 -2274
rect 5658 -2302 5704 -2292
rect 5771 -2263 5786 -2248
tri 5396 -2327 5408 -2315 ne
rect 5408 -2320 5418 -2315
tri 5418 -2320 5423 -2315 sw
rect 5307 -2524 5322 -2438
rect 5408 -2476 5423 -2320
rect 5462 -2362 5490 -2306
tri 5582 -2324 5600 -2306 ne
rect 5600 -2326 5622 -2306
tri 5622 -2326 5642 -2306 sw
tri 5658 -2320 5676 -2302 ne
rect 5481 -2396 5490 -2362
rect 5524 -2335 5566 -2334
rect 5524 -2369 5529 -2335
rect 5559 -2369 5566 -2335
rect 5524 -2378 5566 -2369
rect 5600 -2335 5642 -2326
rect 5600 -2369 5607 -2335
rect 5637 -2369 5642 -2335
rect 5600 -2374 5642 -2369
rect 5676 -2362 5704 -2302
tri 5749 -2315 5771 -2293 se
rect 5771 -2300 5786 -2292
tri 5771 -2315 5786 -2300 nw
tri 5743 -2321 5749 -2315 se
rect 5749 -2321 5758 -2315
rect 5462 -2406 5490 -2396
tri 5490 -2406 5514 -2382 sw
rect 5462 -2438 5504 -2406
tri 5521 -2414 5522 -2413 sw
rect 5521 -2438 5522 -2414
tri 5524 -2415 5561 -2378 ne
rect 5561 -2406 5566 -2378
tri 5566 -2406 5592 -2380 sw
rect 5676 -2396 5685 -2362
rect 5676 -2406 5704 -2396
rect 5561 -2415 5645 -2406
tri 5561 -2434 5580 -2415 ne
rect 5580 -2434 5645 -2415
rect 5462 -2460 5522 -2438
rect 5644 -2438 5645 -2434
rect 5662 -2438 5704 -2406
rect 5644 -2460 5704 -2438
rect 5550 -2476 5567 -2462
rect 5599 -2476 5616 -2462
rect 5743 -2476 5758 -2321
tri 5758 -2328 5771 -2315 nw
rect 5844 -2396 5859 -2168
rect 5844 -2524 5859 -2438
rect 5887 1654 5902 1844
tri 5967 1808 5989 1830 se
rect 5989 1823 6004 1892
tri 5989 1808 6004 1823 nw
rect 6323 1823 6338 1892
tri 5961 1802 5967 1808 se
rect 5967 1802 5976 1808
rect 5961 1786 5976 1802
tri 5976 1795 5989 1808 nw
rect 6130 1800 6147 1814
rect 6179 1800 6196 1814
tri 6323 1808 6338 1823 ne
tri 6338 1808 6360 1830 sw
rect 5961 1750 5976 1758
rect 6042 1786 6102 1800
rect 6057 1776 6102 1786
rect 6057 1758 6085 1776
tri 5961 1735 5976 1750 ne
tri 5976 1735 5998 1757 sw
rect 6042 1748 6085 1758
rect 6100 1772 6102 1776
rect 6224 1786 6284 1800
tri 6338 1795 6351 1808 ne
rect 6351 1802 6360 1808
tri 6360 1802 6366 1808 sw
rect 6224 1776 6269 1786
rect 6100 1748 6174 1772
rect 6042 1744 6174 1748
tri 6174 1744 6202 1772 sw
rect 6224 1762 6226 1776
tri 6224 1760 6226 1762 ne
rect 6238 1758 6269 1776
rect 6238 1748 6284 1758
rect 6351 1787 6366 1802
tri 5976 1723 5988 1735 ne
rect 5988 1730 5998 1735
tri 5998 1730 6003 1735 sw
rect 5887 1384 5902 1612
rect 5988 1574 6003 1730
rect 6042 1688 6070 1744
tri 6162 1726 6180 1744 ne
rect 6180 1724 6202 1744
tri 6202 1724 6222 1744 sw
tri 6238 1730 6256 1748 ne
rect 6061 1654 6070 1688
rect 6104 1715 6146 1716
rect 6104 1681 6109 1715
rect 6139 1681 6146 1715
rect 6104 1672 6146 1681
rect 6180 1715 6222 1724
rect 6180 1681 6187 1715
rect 6217 1681 6222 1715
rect 6180 1676 6222 1681
rect 6256 1688 6284 1748
tri 6329 1735 6351 1757 se
rect 6351 1750 6366 1758
tri 6351 1735 6366 1750 nw
tri 6323 1729 6329 1735 se
rect 6329 1729 6338 1735
rect 6042 1644 6070 1654
tri 6070 1644 6094 1668 sw
rect 6042 1612 6084 1644
tri 6101 1636 6102 1637 sw
rect 6101 1612 6102 1636
tri 6104 1635 6141 1672 ne
rect 6141 1644 6146 1672
tri 6146 1644 6172 1670 sw
rect 6256 1654 6265 1688
rect 6256 1644 6284 1654
rect 6141 1635 6225 1644
tri 6141 1616 6160 1635 ne
rect 6160 1616 6225 1635
rect 6042 1590 6102 1612
rect 6224 1612 6225 1616
rect 6242 1612 6284 1644
rect 6224 1590 6284 1612
rect 6130 1574 6147 1588
rect 6179 1574 6196 1588
tri 5967 1538 5989 1560 se
rect 5989 1553 6004 1574
tri 5989 1538 6004 1553 nw
rect 6323 1553 6338 1729
tri 6338 1722 6351 1735 nw
rect 6424 1654 6439 1844
tri 5961 1532 5967 1538 se
rect 5967 1532 5976 1538
rect 5961 1516 5976 1532
tri 5976 1525 5989 1538 nw
rect 6130 1530 6147 1544
rect 6179 1530 6196 1544
tri 6323 1538 6338 1553 ne
tri 6338 1538 6360 1560 sw
rect 5961 1480 5976 1488
rect 6042 1516 6102 1530
rect 6057 1506 6102 1516
rect 6057 1488 6085 1506
tri 5961 1465 5976 1480 ne
tri 5976 1465 5998 1487 sw
rect 6042 1478 6085 1488
rect 6100 1502 6102 1506
rect 6224 1516 6284 1530
tri 6338 1525 6351 1538 ne
rect 6351 1532 6360 1538
tri 6360 1532 6366 1538 sw
rect 6224 1506 6269 1516
rect 6100 1478 6174 1502
rect 6042 1474 6174 1478
tri 6174 1474 6202 1502 sw
rect 6224 1492 6226 1506
tri 6224 1490 6226 1492 ne
rect 6238 1488 6269 1506
rect 6238 1478 6284 1488
rect 6351 1517 6366 1532
tri 5976 1453 5988 1465 ne
rect 5988 1460 5998 1465
tri 5998 1460 6003 1465 sw
rect 5887 1114 5902 1342
rect 5988 1352 6003 1460
rect 6042 1418 6070 1474
tri 6162 1456 6180 1474 ne
rect 6180 1454 6202 1474
tri 6202 1454 6222 1474 sw
tri 6238 1460 6256 1478 ne
rect 6061 1384 6070 1418
rect 6104 1445 6146 1446
rect 6104 1411 6109 1445
rect 6139 1411 6146 1445
rect 6104 1402 6146 1411
rect 6180 1445 6222 1454
rect 6180 1411 6187 1445
rect 6217 1411 6222 1445
rect 6180 1406 6222 1411
rect 6256 1418 6284 1478
tri 6329 1465 6351 1487 se
rect 6351 1480 6366 1488
tri 6351 1465 6366 1480 nw
tri 6323 1459 6329 1465 se
rect 6329 1459 6338 1465
rect 6042 1374 6070 1384
tri 6070 1374 6094 1398 sw
rect 5988 1304 6004 1352
rect 6042 1342 6084 1374
tri 6101 1366 6102 1367 sw
rect 6101 1342 6102 1366
tri 6104 1365 6141 1402 ne
rect 6141 1374 6146 1402
tri 6146 1374 6172 1400 sw
rect 6256 1384 6265 1418
rect 6256 1374 6284 1384
rect 6141 1365 6225 1374
tri 6141 1346 6160 1365 ne
rect 6160 1346 6225 1365
rect 6042 1320 6102 1342
rect 6224 1342 6225 1346
rect 6242 1342 6284 1374
rect 6224 1320 6284 1342
rect 6130 1304 6147 1318
rect 6179 1304 6196 1318
tri 5967 1268 5989 1290 se
rect 5989 1283 6004 1304
tri 5989 1268 6004 1283 nw
rect 6323 1283 6338 1459
tri 6338 1452 6351 1465 nw
rect 6424 1384 6439 1612
tri 5961 1262 5967 1268 se
rect 5967 1262 5976 1268
rect 5961 1246 5976 1262
tri 5976 1255 5989 1268 nw
rect 6130 1260 6147 1274
rect 6179 1260 6196 1274
tri 6323 1268 6338 1283 ne
tri 6338 1268 6360 1290 sw
rect 5961 1210 5976 1218
rect 6042 1246 6102 1260
rect 6057 1236 6102 1246
rect 6057 1218 6085 1236
tri 5961 1195 5976 1210 ne
tri 5976 1195 5998 1217 sw
rect 6042 1208 6085 1218
rect 6100 1232 6102 1236
rect 6224 1246 6284 1260
tri 6338 1255 6351 1268 ne
rect 6351 1262 6360 1268
tri 6360 1262 6366 1268 sw
rect 6224 1236 6269 1246
rect 6100 1208 6174 1232
rect 6042 1204 6174 1208
tri 6174 1204 6202 1232 sw
rect 6224 1222 6226 1236
tri 6224 1220 6226 1222 ne
rect 6238 1218 6269 1236
rect 6238 1208 6284 1218
rect 6351 1247 6366 1262
tri 5976 1183 5988 1195 ne
rect 5988 1190 5998 1195
tri 5998 1190 6003 1195 sw
rect 5887 844 5902 1072
rect 5988 1034 6003 1190
rect 6042 1148 6070 1204
tri 6162 1186 6180 1204 ne
rect 6180 1184 6202 1204
tri 6202 1184 6222 1204 sw
tri 6238 1190 6256 1208 ne
rect 6061 1114 6070 1148
rect 6104 1175 6146 1176
rect 6104 1141 6109 1175
rect 6139 1141 6146 1175
rect 6104 1132 6146 1141
rect 6180 1175 6222 1184
rect 6180 1141 6187 1175
rect 6217 1141 6222 1175
rect 6180 1136 6222 1141
rect 6256 1148 6284 1208
tri 6329 1195 6351 1217 se
rect 6351 1210 6366 1218
tri 6351 1195 6366 1210 nw
tri 6323 1189 6329 1195 se
rect 6329 1189 6338 1195
rect 6042 1104 6070 1114
tri 6070 1104 6094 1128 sw
rect 6042 1072 6084 1104
tri 6101 1096 6102 1097 sw
rect 6101 1072 6102 1096
tri 6104 1095 6141 1132 ne
rect 6141 1104 6146 1132
tri 6146 1104 6172 1130 sw
rect 6256 1114 6265 1148
rect 6256 1104 6284 1114
rect 6141 1095 6225 1104
tri 6141 1076 6160 1095 ne
rect 6160 1076 6225 1095
rect 6042 1050 6102 1072
rect 6224 1072 6225 1076
rect 6242 1072 6284 1104
rect 6224 1050 6284 1072
rect 6130 1034 6147 1048
rect 6179 1034 6196 1048
tri 5967 998 5989 1020 se
rect 5989 1013 6004 1034
tri 5989 998 6004 1013 nw
rect 6323 1013 6338 1189
tri 6338 1182 6351 1195 nw
rect 6424 1114 6439 1342
tri 5961 992 5967 998 se
rect 5967 992 5976 998
rect 5961 976 5976 992
tri 5976 985 5989 998 nw
rect 6130 990 6147 1004
rect 6179 990 6196 1004
tri 6323 998 6338 1013 ne
tri 6338 998 6360 1020 sw
rect 5961 940 5976 948
rect 6042 976 6102 990
rect 6057 966 6102 976
rect 6057 948 6085 966
tri 5961 925 5976 940 ne
tri 5976 925 5998 947 sw
rect 6042 938 6085 948
rect 6100 962 6102 966
rect 6224 976 6284 990
tri 6338 985 6351 998 ne
rect 6351 992 6360 998
tri 6360 992 6366 998 sw
rect 6224 966 6269 976
rect 6100 938 6174 962
rect 6042 934 6174 938
tri 6174 934 6202 962 sw
rect 6224 952 6226 966
tri 6224 950 6226 952 ne
rect 6238 948 6269 966
rect 6238 938 6284 948
rect 6351 977 6366 992
tri 5976 913 5988 925 ne
rect 5988 920 5998 925
tri 5998 920 6003 925 sw
rect 5887 574 5902 802
rect 5988 812 6003 920
rect 6042 878 6070 934
tri 6162 916 6180 934 ne
rect 6180 914 6202 934
tri 6202 914 6222 934 sw
tri 6238 920 6256 938 ne
rect 6061 844 6070 878
rect 6104 905 6146 906
rect 6104 871 6109 905
rect 6139 871 6146 905
rect 6104 862 6146 871
rect 6180 905 6222 914
rect 6180 871 6187 905
rect 6217 871 6222 905
rect 6180 866 6222 871
rect 6256 878 6284 938
tri 6329 925 6351 947 se
rect 6351 940 6366 948
tri 6351 925 6366 940 nw
tri 6323 919 6329 925 se
rect 6329 919 6338 925
rect 6042 834 6070 844
tri 6070 834 6094 858 sw
rect 5988 764 6004 812
rect 6042 802 6084 834
tri 6101 826 6102 827 sw
rect 6101 802 6102 826
tri 6104 825 6141 862 ne
rect 6141 834 6146 862
tri 6146 834 6172 860 sw
rect 6256 844 6265 878
rect 6256 834 6284 844
rect 6141 825 6225 834
tri 6141 806 6160 825 ne
rect 6160 806 6225 825
rect 6042 780 6102 802
rect 6224 802 6225 806
rect 6242 802 6284 834
rect 6224 780 6284 802
rect 6130 764 6147 778
rect 6179 764 6196 778
tri 5967 728 5989 750 se
rect 5989 743 6004 764
tri 5989 728 6004 743 nw
rect 6323 743 6338 919
tri 6338 912 6351 925 nw
rect 6424 844 6439 1072
tri 5961 722 5967 728 se
rect 5967 722 5976 728
rect 5961 706 5976 722
tri 5976 715 5989 728 nw
rect 6130 720 6147 734
rect 6179 720 6196 734
tri 6323 728 6338 743 ne
tri 6338 728 6360 750 sw
rect 5961 670 5976 678
rect 6042 706 6102 720
rect 6057 696 6102 706
rect 6057 678 6085 696
tri 5961 655 5976 670 ne
tri 5976 655 5998 677 sw
rect 6042 668 6085 678
rect 6100 692 6102 696
rect 6224 706 6284 720
tri 6338 715 6351 728 ne
rect 6351 722 6360 728
tri 6360 722 6366 728 sw
rect 6224 696 6269 706
rect 6100 668 6174 692
rect 6042 664 6174 668
tri 6174 664 6202 692 sw
rect 6224 682 6226 696
tri 6224 680 6226 682 ne
rect 6238 678 6269 696
rect 6238 668 6284 678
rect 6351 707 6366 722
tri 5976 643 5988 655 ne
rect 5988 650 5998 655
tri 5998 650 6003 655 sw
rect 5887 304 5902 532
rect 5988 494 6003 650
rect 6042 608 6070 664
tri 6162 646 6180 664 ne
rect 6180 644 6202 664
tri 6202 644 6222 664 sw
tri 6238 650 6256 668 ne
rect 6061 574 6070 608
rect 6104 635 6146 636
rect 6104 601 6109 635
rect 6139 601 6146 635
rect 6104 592 6146 601
rect 6180 635 6222 644
rect 6180 601 6187 635
rect 6217 601 6222 635
rect 6180 596 6222 601
rect 6256 608 6284 668
tri 6329 655 6351 677 se
rect 6351 670 6366 678
tri 6351 655 6366 670 nw
tri 6323 649 6329 655 se
rect 6329 649 6338 655
rect 6042 564 6070 574
tri 6070 564 6094 588 sw
rect 6042 532 6084 564
tri 6101 556 6102 557 sw
rect 6101 532 6102 556
tri 6104 555 6141 592 ne
rect 6141 564 6146 592
tri 6146 564 6172 590 sw
rect 6256 574 6265 608
rect 6256 564 6284 574
rect 6141 555 6225 564
tri 6141 536 6160 555 ne
rect 6160 536 6225 555
rect 6042 510 6102 532
rect 6224 532 6225 536
rect 6242 532 6284 564
rect 6224 510 6284 532
rect 6130 494 6147 508
rect 6179 494 6196 508
tri 5967 458 5989 480 se
rect 5989 473 6004 494
tri 5989 458 6004 473 nw
rect 6323 473 6338 649
tri 6338 642 6351 655 nw
rect 6424 574 6439 802
tri 5961 452 5967 458 se
rect 5967 452 5976 458
rect 5961 436 5976 452
tri 5976 445 5989 458 nw
rect 6130 450 6147 464
rect 6179 450 6196 464
tri 6323 458 6338 473 ne
tri 6338 458 6360 480 sw
rect 5961 400 5976 408
rect 6042 436 6102 450
rect 6057 426 6102 436
rect 6057 408 6085 426
tri 5961 385 5976 400 ne
tri 5976 385 5998 407 sw
rect 6042 398 6085 408
rect 6100 422 6102 426
rect 6224 436 6284 450
tri 6338 445 6351 458 ne
rect 6351 452 6360 458
tri 6360 452 6366 458 sw
rect 6224 426 6269 436
rect 6100 398 6174 422
rect 6042 394 6174 398
tri 6174 394 6202 422 sw
rect 6224 412 6226 426
tri 6224 410 6226 412 ne
rect 6238 408 6269 426
rect 6238 398 6284 408
rect 6351 437 6366 452
tri 5976 373 5988 385 ne
rect 5988 380 5998 385
tri 5998 380 6003 385 sw
rect 5887 34 5902 262
rect 5988 272 6003 380
rect 6042 338 6070 394
tri 6162 376 6180 394 ne
rect 6180 374 6202 394
tri 6202 374 6222 394 sw
tri 6238 380 6256 398 ne
rect 6061 304 6070 338
rect 6104 365 6146 366
rect 6104 331 6109 365
rect 6139 331 6146 365
rect 6104 322 6146 331
rect 6180 365 6222 374
rect 6180 331 6187 365
rect 6217 331 6222 365
rect 6180 326 6222 331
rect 6256 338 6284 398
tri 6329 385 6351 407 se
rect 6351 400 6366 408
tri 6351 385 6366 400 nw
tri 6323 379 6329 385 se
rect 6329 379 6338 385
rect 6042 294 6070 304
tri 6070 294 6094 318 sw
rect 5988 224 6004 272
rect 6042 262 6084 294
tri 6101 286 6102 287 sw
rect 6101 262 6102 286
tri 6104 285 6141 322 ne
rect 6141 294 6146 322
tri 6146 294 6172 320 sw
rect 6256 304 6265 338
rect 6256 294 6284 304
rect 6141 285 6225 294
tri 6141 266 6160 285 ne
rect 6160 266 6225 285
rect 6042 240 6102 262
rect 6224 262 6225 266
rect 6242 262 6284 294
rect 6224 240 6284 262
rect 6130 224 6147 238
rect 6179 224 6196 238
tri 5967 188 5989 210 se
rect 5989 203 6004 224
tri 5989 188 6004 203 nw
rect 6323 203 6338 379
tri 6338 372 6351 385 nw
rect 6424 304 6439 532
tri 5961 182 5967 188 se
rect 5967 182 5976 188
rect 5961 166 5976 182
tri 5976 175 5989 188 nw
rect 6130 180 6147 194
rect 6179 180 6196 194
tri 6323 188 6338 203 ne
tri 6338 188 6360 210 sw
rect 5961 130 5976 138
rect 6042 166 6102 180
rect 6057 156 6102 166
rect 6057 138 6085 156
tri 5961 115 5976 130 ne
tri 5976 115 5998 137 sw
rect 6042 128 6085 138
rect 6100 152 6102 156
rect 6224 166 6284 180
tri 6338 175 6351 188 ne
rect 6351 182 6360 188
tri 6360 182 6366 188 sw
rect 6224 156 6269 166
rect 6100 128 6174 152
rect 6042 124 6174 128
tri 6174 124 6202 152 sw
rect 6224 142 6226 156
tri 6224 140 6226 142 ne
rect 6238 138 6269 156
rect 6238 128 6284 138
rect 6351 167 6366 182
tri 5976 103 5988 115 ne
rect 5988 110 5998 115
tri 5998 110 6003 115 sw
rect 5887 -236 5902 -8
rect 5988 -46 6003 110
rect 6042 68 6070 124
tri 6162 106 6180 124 ne
rect 6180 104 6202 124
tri 6202 104 6222 124 sw
tri 6238 110 6256 128 ne
rect 6061 34 6070 68
rect 6104 95 6146 96
rect 6104 61 6109 95
rect 6139 61 6146 95
rect 6104 52 6146 61
rect 6180 95 6222 104
rect 6180 61 6187 95
rect 6217 61 6222 95
rect 6180 56 6222 61
rect 6256 68 6284 128
tri 6329 115 6351 137 se
rect 6351 130 6366 138
tri 6351 115 6366 130 nw
tri 6323 109 6329 115 se
rect 6329 109 6338 115
rect 6042 24 6070 34
tri 6070 24 6094 48 sw
rect 6042 -8 6084 24
tri 6101 16 6102 17 sw
rect 6101 -8 6102 16
tri 6104 15 6141 52 ne
rect 6141 24 6146 52
tri 6146 24 6172 50 sw
rect 6256 34 6265 68
rect 6256 24 6284 34
rect 6141 15 6225 24
tri 6141 -4 6160 15 ne
rect 6160 -4 6225 15
rect 6042 -30 6102 -8
rect 6224 -8 6225 -4
rect 6242 -8 6284 24
rect 6224 -30 6284 -8
rect 6130 -46 6147 -32
rect 6179 -46 6196 -32
tri 5967 -82 5989 -60 se
rect 5989 -67 6004 -46
tri 5989 -82 6004 -67 nw
rect 6323 -67 6338 109
tri 6338 102 6351 115 nw
rect 6424 34 6439 262
tri 5961 -88 5967 -82 se
rect 5967 -88 5976 -82
rect 5961 -104 5976 -88
tri 5976 -95 5989 -82 nw
rect 6130 -90 6147 -76
rect 6179 -90 6196 -76
tri 6323 -82 6338 -67 ne
tri 6338 -82 6360 -60 sw
rect 5961 -140 5976 -132
rect 6042 -104 6102 -90
rect 6057 -114 6102 -104
rect 6057 -132 6085 -114
tri 5961 -155 5976 -140 ne
tri 5976 -155 5998 -133 sw
rect 6042 -142 6085 -132
rect 6100 -118 6102 -114
rect 6224 -104 6284 -90
tri 6338 -95 6351 -82 ne
rect 6351 -88 6360 -82
tri 6360 -88 6366 -82 sw
rect 6224 -114 6269 -104
rect 6100 -142 6174 -118
rect 6042 -146 6174 -142
tri 6174 -146 6202 -118 sw
rect 6224 -128 6226 -114
tri 6224 -130 6226 -128 ne
rect 6238 -132 6269 -114
rect 6238 -142 6284 -132
rect 6351 -103 6366 -88
tri 5976 -167 5988 -155 ne
rect 5988 -160 5998 -155
tri 5998 -160 6003 -155 sw
rect 5887 -506 5902 -278
rect 5988 -268 6003 -160
rect 6042 -202 6070 -146
tri 6162 -164 6180 -146 ne
rect 6180 -166 6202 -146
tri 6202 -166 6222 -146 sw
tri 6238 -160 6256 -142 ne
rect 6061 -236 6070 -202
rect 6104 -175 6146 -174
rect 6104 -209 6109 -175
rect 6139 -209 6146 -175
rect 6104 -218 6146 -209
rect 6180 -175 6222 -166
rect 6180 -209 6187 -175
rect 6217 -209 6222 -175
rect 6180 -214 6222 -209
rect 6256 -202 6284 -142
tri 6329 -155 6351 -133 se
rect 6351 -140 6366 -132
tri 6351 -155 6366 -140 nw
tri 6323 -161 6329 -155 se
rect 6329 -161 6338 -155
rect 6042 -246 6070 -236
tri 6070 -246 6094 -222 sw
rect 5988 -316 6004 -268
rect 6042 -278 6084 -246
tri 6101 -254 6102 -253 sw
rect 6101 -278 6102 -254
tri 6104 -255 6141 -218 ne
rect 6141 -246 6146 -218
tri 6146 -246 6172 -220 sw
rect 6256 -236 6265 -202
rect 6256 -246 6284 -236
rect 6141 -255 6225 -246
tri 6141 -274 6160 -255 ne
rect 6160 -274 6225 -255
rect 6042 -300 6102 -278
rect 6224 -278 6225 -274
rect 6242 -278 6284 -246
rect 6224 -300 6284 -278
rect 6130 -316 6147 -302
rect 6179 -316 6196 -302
tri 5967 -352 5989 -330 se
rect 5989 -337 6004 -316
tri 5989 -352 6004 -337 nw
rect 6323 -337 6338 -161
tri 6338 -168 6351 -155 nw
rect 6424 -236 6439 -8
tri 5961 -358 5967 -352 se
rect 5967 -358 5976 -352
rect 5961 -374 5976 -358
tri 5976 -365 5989 -352 nw
rect 6130 -360 6147 -346
rect 6179 -360 6196 -346
tri 6323 -352 6338 -337 ne
tri 6338 -352 6360 -330 sw
rect 5961 -410 5976 -402
rect 6042 -374 6102 -360
rect 6057 -384 6102 -374
rect 6057 -402 6085 -384
tri 5961 -425 5976 -410 ne
tri 5976 -425 5998 -403 sw
rect 6042 -412 6085 -402
rect 6100 -388 6102 -384
rect 6224 -374 6284 -360
tri 6338 -365 6351 -352 ne
rect 6351 -358 6360 -352
tri 6360 -358 6366 -352 sw
rect 6224 -384 6269 -374
rect 6100 -412 6174 -388
rect 6042 -416 6174 -412
tri 6174 -416 6202 -388 sw
rect 6224 -398 6226 -384
tri 6224 -400 6226 -398 ne
rect 6238 -402 6269 -384
rect 6238 -412 6284 -402
rect 6351 -373 6366 -358
tri 5976 -437 5988 -425 ne
rect 5988 -430 5998 -425
tri 5998 -430 6003 -425 sw
rect 5887 -776 5902 -548
rect 5988 -586 6003 -430
rect 6042 -472 6070 -416
tri 6162 -434 6180 -416 ne
rect 6180 -436 6202 -416
tri 6202 -436 6222 -416 sw
tri 6238 -430 6256 -412 ne
rect 6061 -506 6070 -472
rect 6104 -445 6146 -444
rect 6104 -479 6109 -445
rect 6139 -479 6146 -445
rect 6104 -488 6146 -479
rect 6180 -445 6222 -436
rect 6180 -479 6187 -445
rect 6217 -479 6222 -445
rect 6180 -484 6222 -479
rect 6256 -472 6284 -412
tri 6329 -425 6351 -403 se
rect 6351 -410 6366 -402
tri 6351 -425 6366 -410 nw
tri 6323 -431 6329 -425 se
rect 6329 -431 6338 -425
rect 6042 -516 6070 -506
tri 6070 -516 6094 -492 sw
rect 6042 -548 6084 -516
tri 6101 -524 6102 -523 sw
rect 6101 -548 6102 -524
tri 6104 -525 6141 -488 ne
rect 6141 -516 6146 -488
tri 6146 -516 6172 -490 sw
rect 6256 -506 6265 -472
rect 6256 -516 6284 -506
rect 6141 -525 6225 -516
tri 6141 -544 6160 -525 ne
rect 6160 -544 6225 -525
rect 6042 -570 6102 -548
rect 6224 -548 6225 -544
rect 6242 -548 6284 -516
rect 6224 -570 6284 -548
rect 6130 -586 6147 -572
rect 6179 -586 6196 -572
tri 5967 -622 5989 -600 se
rect 5989 -607 6004 -586
tri 5989 -622 6004 -607 nw
rect 6323 -607 6338 -431
tri 6338 -438 6351 -425 nw
rect 6424 -506 6439 -278
tri 5961 -628 5967 -622 se
rect 5967 -628 5976 -622
rect 5961 -644 5976 -628
tri 5976 -635 5989 -622 nw
rect 6130 -630 6147 -616
rect 6179 -630 6196 -616
tri 6323 -622 6338 -607 ne
tri 6338 -622 6360 -600 sw
rect 5961 -680 5976 -672
rect 6042 -644 6102 -630
rect 6057 -654 6102 -644
rect 6057 -672 6085 -654
tri 5961 -695 5976 -680 ne
tri 5976 -695 5998 -673 sw
rect 6042 -682 6085 -672
rect 6100 -658 6102 -654
rect 6224 -644 6284 -630
tri 6338 -635 6351 -622 ne
rect 6351 -628 6360 -622
tri 6360 -628 6366 -622 sw
rect 6224 -654 6269 -644
rect 6100 -682 6174 -658
rect 6042 -686 6174 -682
tri 6174 -686 6202 -658 sw
rect 6224 -668 6226 -654
tri 6224 -670 6226 -668 ne
rect 6238 -672 6269 -654
rect 6238 -682 6284 -672
rect 6351 -643 6366 -628
tri 5976 -707 5988 -695 ne
rect 5988 -700 5998 -695
tri 5998 -700 6003 -695 sw
rect 5887 -1046 5902 -818
rect 5988 -808 6003 -700
rect 6042 -742 6070 -686
tri 6162 -704 6180 -686 ne
rect 6180 -706 6202 -686
tri 6202 -706 6222 -686 sw
tri 6238 -700 6256 -682 ne
rect 6061 -776 6070 -742
rect 6104 -715 6146 -714
rect 6104 -749 6109 -715
rect 6139 -749 6146 -715
rect 6104 -758 6146 -749
rect 6180 -715 6222 -706
rect 6180 -749 6187 -715
rect 6217 -749 6222 -715
rect 6180 -754 6222 -749
rect 6256 -742 6284 -682
tri 6329 -695 6351 -673 se
rect 6351 -680 6366 -672
tri 6351 -695 6366 -680 nw
tri 6323 -701 6329 -695 se
rect 6329 -701 6338 -695
rect 6042 -786 6070 -776
tri 6070 -786 6094 -762 sw
rect 5988 -856 6004 -808
rect 6042 -818 6084 -786
tri 6101 -794 6102 -793 sw
rect 6101 -818 6102 -794
tri 6104 -795 6141 -758 ne
rect 6141 -786 6146 -758
tri 6146 -786 6172 -760 sw
rect 6256 -776 6265 -742
rect 6256 -786 6284 -776
rect 6141 -795 6225 -786
tri 6141 -814 6160 -795 ne
rect 6160 -814 6225 -795
rect 6042 -840 6102 -818
rect 6224 -818 6225 -814
rect 6242 -818 6284 -786
rect 6224 -840 6284 -818
rect 6130 -856 6147 -842
rect 6179 -856 6196 -842
tri 5967 -892 5989 -870 se
rect 5989 -877 6004 -856
tri 5989 -892 6004 -877 nw
rect 6323 -877 6338 -701
tri 6338 -708 6351 -695 nw
rect 6424 -776 6439 -548
tri 5961 -898 5967 -892 se
rect 5967 -898 5976 -892
rect 5961 -914 5976 -898
tri 5976 -905 5989 -892 nw
rect 6130 -900 6147 -886
rect 6179 -900 6196 -886
tri 6323 -892 6338 -877 ne
tri 6338 -892 6360 -870 sw
rect 5961 -950 5976 -942
rect 6042 -914 6102 -900
rect 6057 -924 6102 -914
rect 6057 -942 6085 -924
tri 5961 -965 5976 -950 ne
tri 5976 -965 5998 -943 sw
rect 6042 -952 6085 -942
rect 6100 -928 6102 -924
rect 6224 -914 6284 -900
tri 6338 -905 6351 -892 ne
rect 6351 -898 6360 -892
tri 6360 -898 6366 -892 sw
rect 6224 -924 6269 -914
rect 6100 -952 6174 -928
rect 6042 -956 6174 -952
tri 6174 -956 6202 -928 sw
rect 6224 -938 6226 -924
tri 6224 -940 6226 -938 ne
rect 6238 -942 6269 -924
rect 6238 -952 6284 -942
rect 6351 -913 6366 -898
tri 5976 -977 5988 -965 ne
rect 5988 -970 5998 -965
tri 5998 -970 6003 -965 sw
rect 5887 -1316 5902 -1088
rect 5988 -1126 6003 -970
rect 6042 -1012 6070 -956
tri 6162 -974 6180 -956 ne
rect 6180 -976 6202 -956
tri 6202 -976 6222 -956 sw
tri 6238 -970 6256 -952 ne
rect 6061 -1046 6070 -1012
rect 6104 -985 6146 -984
rect 6104 -1019 6109 -985
rect 6139 -1019 6146 -985
rect 6104 -1028 6146 -1019
rect 6180 -985 6222 -976
rect 6180 -1019 6187 -985
rect 6217 -1019 6222 -985
rect 6180 -1024 6222 -1019
rect 6256 -1012 6284 -952
tri 6329 -965 6351 -943 se
rect 6351 -950 6366 -942
tri 6351 -965 6366 -950 nw
tri 6323 -971 6329 -965 se
rect 6329 -971 6338 -965
rect 6042 -1056 6070 -1046
tri 6070 -1056 6094 -1032 sw
rect 6042 -1088 6084 -1056
tri 6101 -1064 6102 -1063 sw
rect 6101 -1088 6102 -1064
tri 6104 -1065 6141 -1028 ne
rect 6141 -1056 6146 -1028
tri 6146 -1056 6172 -1030 sw
rect 6256 -1046 6265 -1012
rect 6256 -1056 6284 -1046
rect 6141 -1065 6225 -1056
tri 6141 -1084 6160 -1065 ne
rect 6160 -1084 6225 -1065
rect 6042 -1110 6102 -1088
rect 6224 -1088 6225 -1084
rect 6242 -1088 6284 -1056
rect 6224 -1110 6284 -1088
rect 6130 -1126 6147 -1112
rect 6179 -1126 6196 -1112
tri 5967 -1162 5989 -1140 se
rect 5989 -1147 6004 -1126
tri 5989 -1162 6004 -1147 nw
rect 6323 -1147 6338 -971
tri 6338 -978 6351 -965 nw
rect 6424 -1046 6439 -818
tri 5961 -1168 5967 -1162 se
rect 5967 -1168 5976 -1162
rect 5961 -1184 5976 -1168
tri 5976 -1175 5989 -1162 nw
rect 6130 -1170 6147 -1156
rect 6179 -1170 6196 -1156
tri 6323 -1162 6338 -1147 ne
tri 6338 -1162 6360 -1140 sw
rect 5961 -1220 5976 -1212
rect 6042 -1184 6102 -1170
rect 6057 -1194 6102 -1184
rect 6057 -1212 6085 -1194
tri 5961 -1235 5976 -1220 ne
tri 5976 -1235 5998 -1213 sw
rect 6042 -1222 6085 -1212
rect 6100 -1198 6102 -1194
rect 6224 -1184 6284 -1170
tri 6338 -1175 6351 -1162 ne
rect 6351 -1168 6360 -1162
tri 6360 -1168 6366 -1162 sw
rect 6224 -1194 6269 -1184
rect 6100 -1222 6174 -1198
rect 6042 -1226 6174 -1222
tri 6174 -1226 6202 -1198 sw
rect 6224 -1208 6226 -1194
tri 6224 -1210 6226 -1208 ne
rect 6238 -1212 6269 -1194
rect 6238 -1222 6284 -1212
rect 6351 -1183 6366 -1168
tri 5976 -1247 5988 -1235 ne
rect 5988 -1240 5998 -1235
tri 5998 -1240 6003 -1235 sw
rect 5887 -1586 5902 -1358
rect 5988 -1348 6003 -1240
rect 6042 -1282 6070 -1226
tri 6162 -1244 6180 -1226 ne
rect 6180 -1246 6202 -1226
tri 6202 -1246 6222 -1226 sw
tri 6238 -1240 6256 -1222 ne
rect 6061 -1316 6070 -1282
rect 6104 -1255 6146 -1254
rect 6104 -1289 6109 -1255
rect 6139 -1289 6146 -1255
rect 6104 -1298 6146 -1289
rect 6180 -1255 6222 -1246
rect 6180 -1289 6187 -1255
rect 6217 -1289 6222 -1255
rect 6180 -1294 6222 -1289
rect 6256 -1282 6284 -1222
tri 6329 -1235 6351 -1213 se
rect 6351 -1220 6366 -1212
tri 6351 -1235 6366 -1220 nw
tri 6323 -1241 6329 -1235 se
rect 6329 -1241 6338 -1235
rect 6042 -1326 6070 -1316
tri 6070 -1326 6094 -1302 sw
rect 5988 -1396 6004 -1348
rect 6042 -1358 6084 -1326
tri 6101 -1334 6102 -1333 sw
rect 6101 -1358 6102 -1334
tri 6104 -1335 6141 -1298 ne
rect 6141 -1326 6146 -1298
tri 6146 -1326 6172 -1300 sw
rect 6256 -1316 6265 -1282
rect 6256 -1326 6284 -1316
rect 6141 -1335 6225 -1326
tri 6141 -1354 6160 -1335 ne
rect 6160 -1354 6225 -1335
rect 6042 -1380 6102 -1358
rect 6224 -1358 6225 -1354
rect 6242 -1358 6284 -1326
rect 6224 -1380 6284 -1358
rect 6130 -1396 6147 -1382
rect 6179 -1396 6196 -1382
tri 5967 -1432 5989 -1410 se
rect 5989 -1417 6004 -1396
tri 5989 -1432 6004 -1417 nw
rect 6323 -1417 6338 -1241
tri 6338 -1248 6351 -1235 nw
rect 6424 -1316 6439 -1088
tri 5961 -1438 5967 -1432 se
rect 5967 -1438 5976 -1432
rect 5961 -1454 5976 -1438
tri 5976 -1445 5989 -1432 nw
rect 6130 -1440 6147 -1426
rect 6179 -1440 6196 -1426
tri 6323 -1432 6338 -1417 ne
tri 6338 -1432 6360 -1410 sw
rect 5961 -1490 5976 -1482
rect 6042 -1454 6102 -1440
rect 6057 -1464 6102 -1454
rect 6057 -1482 6085 -1464
tri 5961 -1505 5976 -1490 ne
tri 5976 -1505 5998 -1483 sw
rect 6042 -1492 6085 -1482
rect 6100 -1468 6102 -1464
rect 6224 -1454 6284 -1440
tri 6338 -1445 6351 -1432 ne
rect 6351 -1438 6360 -1432
tri 6360 -1438 6366 -1432 sw
rect 6224 -1464 6269 -1454
rect 6100 -1492 6174 -1468
rect 6042 -1496 6174 -1492
tri 6174 -1496 6202 -1468 sw
rect 6224 -1478 6226 -1464
tri 6224 -1480 6226 -1478 ne
rect 6238 -1482 6269 -1464
rect 6238 -1492 6284 -1482
rect 6351 -1453 6366 -1438
tri 5976 -1517 5988 -1505 ne
rect 5988 -1510 5998 -1505
tri 5998 -1510 6003 -1505 sw
rect 5887 -1856 5902 -1628
rect 5988 -1666 6003 -1510
rect 6042 -1552 6070 -1496
tri 6162 -1514 6180 -1496 ne
rect 6180 -1516 6202 -1496
tri 6202 -1516 6222 -1496 sw
tri 6238 -1510 6256 -1492 ne
rect 6061 -1586 6070 -1552
rect 6104 -1525 6146 -1524
rect 6104 -1559 6109 -1525
rect 6139 -1559 6146 -1525
rect 6104 -1568 6146 -1559
rect 6180 -1525 6222 -1516
rect 6180 -1559 6187 -1525
rect 6217 -1559 6222 -1525
rect 6180 -1564 6222 -1559
rect 6256 -1552 6284 -1492
tri 6329 -1505 6351 -1483 se
rect 6351 -1490 6366 -1482
tri 6351 -1505 6366 -1490 nw
tri 6323 -1511 6329 -1505 se
rect 6329 -1511 6338 -1505
rect 6042 -1596 6070 -1586
tri 6070 -1596 6094 -1572 sw
rect 6042 -1628 6084 -1596
tri 6101 -1604 6102 -1603 sw
rect 6101 -1628 6102 -1604
tri 6104 -1605 6141 -1568 ne
rect 6141 -1596 6146 -1568
tri 6146 -1596 6172 -1570 sw
rect 6256 -1586 6265 -1552
rect 6256 -1596 6284 -1586
rect 6141 -1605 6225 -1596
tri 6141 -1624 6160 -1605 ne
rect 6160 -1624 6225 -1605
rect 6042 -1650 6102 -1628
rect 6224 -1628 6225 -1624
rect 6242 -1628 6284 -1596
rect 6224 -1650 6284 -1628
rect 6130 -1666 6147 -1652
rect 6179 -1666 6196 -1652
tri 5967 -1702 5989 -1680 se
rect 5989 -1687 6004 -1666
tri 5989 -1702 6004 -1687 nw
rect 6323 -1687 6338 -1511
tri 6338 -1518 6351 -1505 nw
rect 6424 -1586 6439 -1358
tri 5961 -1708 5967 -1702 se
rect 5967 -1708 5976 -1702
rect 5961 -1724 5976 -1708
tri 5976 -1715 5989 -1702 nw
rect 6130 -1710 6147 -1696
rect 6179 -1710 6196 -1696
tri 6323 -1702 6338 -1687 ne
tri 6338 -1702 6360 -1680 sw
rect 5961 -1760 5976 -1752
rect 6042 -1724 6102 -1710
rect 6057 -1734 6102 -1724
rect 6057 -1752 6085 -1734
tri 5961 -1775 5976 -1760 ne
tri 5976 -1775 5998 -1753 sw
rect 6042 -1762 6085 -1752
rect 6100 -1738 6102 -1734
rect 6224 -1724 6284 -1710
tri 6338 -1715 6351 -1702 ne
rect 6351 -1708 6360 -1702
tri 6360 -1708 6366 -1702 sw
rect 6224 -1734 6269 -1724
rect 6100 -1762 6174 -1738
rect 6042 -1766 6174 -1762
tri 6174 -1766 6202 -1738 sw
rect 6224 -1748 6226 -1734
tri 6224 -1750 6226 -1748 ne
rect 6238 -1752 6269 -1734
rect 6238 -1762 6284 -1752
rect 6351 -1723 6366 -1708
tri 5976 -1787 5988 -1775 ne
rect 5988 -1780 5998 -1775
tri 5998 -1780 6003 -1775 sw
rect 5887 -2126 5902 -1898
rect 5988 -1888 6003 -1780
rect 6042 -1822 6070 -1766
tri 6162 -1784 6180 -1766 ne
rect 6180 -1786 6202 -1766
tri 6202 -1786 6222 -1766 sw
tri 6238 -1780 6256 -1762 ne
rect 6061 -1856 6070 -1822
rect 6104 -1795 6146 -1794
rect 6104 -1829 6109 -1795
rect 6139 -1829 6146 -1795
rect 6104 -1838 6146 -1829
rect 6180 -1795 6222 -1786
rect 6180 -1829 6187 -1795
rect 6217 -1829 6222 -1795
rect 6180 -1834 6222 -1829
rect 6256 -1822 6284 -1762
tri 6329 -1775 6351 -1753 se
rect 6351 -1760 6366 -1752
tri 6351 -1775 6366 -1760 nw
tri 6323 -1781 6329 -1775 se
rect 6329 -1781 6338 -1775
rect 6042 -1866 6070 -1856
tri 6070 -1866 6094 -1842 sw
rect 5988 -1936 6004 -1888
rect 6042 -1898 6084 -1866
tri 6101 -1874 6102 -1873 sw
rect 6101 -1898 6102 -1874
tri 6104 -1875 6141 -1838 ne
rect 6141 -1866 6146 -1838
tri 6146 -1866 6172 -1840 sw
rect 6256 -1856 6265 -1822
rect 6256 -1866 6284 -1856
rect 6141 -1875 6225 -1866
tri 6141 -1894 6160 -1875 ne
rect 6160 -1894 6225 -1875
rect 6042 -1920 6102 -1898
rect 6224 -1898 6225 -1894
rect 6242 -1898 6284 -1866
rect 6224 -1920 6284 -1898
rect 6130 -1936 6147 -1922
rect 6179 -1936 6196 -1922
tri 5967 -1972 5989 -1950 se
rect 5989 -1957 6004 -1936
tri 5989 -1972 6004 -1957 nw
rect 6323 -1957 6338 -1781
tri 6338 -1788 6351 -1775 nw
rect 6424 -1856 6439 -1628
tri 5961 -1978 5967 -1972 se
rect 5967 -1978 5976 -1972
rect 5961 -1994 5976 -1978
tri 5976 -1985 5989 -1972 nw
rect 6130 -1980 6147 -1966
rect 6179 -1980 6196 -1966
tri 6323 -1972 6338 -1957 ne
tri 6338 -1972 6360 -1950 sw
rect 5961 -2030 5976 -2022
rect 6042 -1994 6102 -1980
rect 6057 -2004 6102 -1994
rect 6057 -2022 6085 -2004
tri 5961 -2045 5976 -2030 ne
tri 5976 -2045 5998 -2023 sw
rect 6042 -2032 6085 -2022
rect 6100 -2008 6102 -2004
rect 6224 -1994 6284 -1980
tri 6338 -1985 6351 -1972 ne
rect 6351 -1978 6360 -1972
tri 6360 -1978 6366 -1972 sw
rect 6224 -2004 6269 -1994
rect 6100 -2032 6174 -2008
rect 6042 -2036 6174 -2032
tri 6174 -2036 6202 -2008 sw
rect 6224 -2018 6226 -2004
tri 6224 -2020 6226 -2018 ne
rect 6238 -2022 6269 -2004
rect 6238 -2032 6284 -2022
rect 6351 -1993 6366 -1978
tri 5976 -2057 5988 -2045 ne
rect 5988 -2050 5998 -2045
tri 5998 -2050 6003 -2045 sw
rect 5887 -2396 5902 -2168
rect 5988 -2206 6003 -2050
rect 6042 -2092 6070 -2036
tri 6162 -2054 6180 -2036 ne
rect 6180 -2056 6202 -2036
tri 6202 -2056 6222 -2036 sw
tri 6238 -2050 6256 -2032 ne
rect 6061 -2126 6070 -2092
rect 6104 -2065 6146 -2064
rect 6104 -2099 6109 -2065
rect 6139 -2099 6146 -2065
rect 6104 -2108 6146 -2099
rect 6180 -2065 6222 -2056
rect 6180 -2099 6187 -2065
rect 6217 -2099 6222 -2065
rect 6180 -2104 6222 -2099
rect 6256 -2092 6284 -2032
tri 6329 -2045 6351 -2023 se
rect 6351 -2030 6366 -2022
tri 6351 -2045 6366 -2030 nw
tri 6323 -2051 6329 -2045 se
rect 6329 -2051 6338 -2045
rect 6042 -2136 6070 -2126
tri 6070 -2136 6094 -2112 sw
rect 6042 -2168 6084 -2136
tri 6101 -2144 6102 -2143 sw
rect 6101 -2168 6102 -2144
tri 6104 -2145 6141 -2108 ne
rect 6141 -2136 6146 -2108
tri 6146 -2136 6172 -2110 sw
rect 6256 -2126 6265 -2092
rect 6256 -2136 6284 -2126
rect 6141 -2145 6225 -2136
tri 6141 -2164 6160 -2145 ne
rect 6160 -2164 6225 -2145
rect 6042 -2190 6102 -2168
rect 6224 -2168 6225 -2164
rect 6242 -2168 6284 -2136
rect 6224 -2190 6284 -2168
rect 6130 -2206 6147 -2192
rect 6179 -2206 6196 -2192
tri 5967 -2242 5989 -2220 se
rect 5989 -2227 6004 -2206
tri 5989 -2242 6004 -2227 nw
rect 6323 -2227 6338 -2051
tri 6338 -2058 6351 -2045 nw
rect 6424 -2126 6439 -1898
tri 5961 -2248 5967 -2242 se
rect 5967 -2248 5976 -2242
rect 5961 -2264 5976 -2248
tri 5976 -2255 5989 -2242 nw
rect 6130 -2250 6147 -2236
rect 6179 -2250 6196 -2236
tri 6323 -2242 6338 -2227 ne
tri 6338 -2242 6360 -2220 sw
rect 5961 -2300 5976 -2292
rect 6042 -2264 6102 -2250
rect 6057 -2274 6102 -2264
rect 6057 -2292 6085 -2274
tri 5961 -2315 5976 -2300 ne
tri 5976 -2315 5998 -2293 sw
rect 6042 -2302 6085 -2292
rect 6100 -2278 6102 -2274
rect 6224 -2264 6284 -2250
tri 6338 -2255 6351 -2242 ne
rect 6351 -2248 6360 -2242
tri 6360 -2248 6366 -2242 sw
rect 6224 -2274 6269 -2264
rect 6100 -2302 6174 -2278
rect 6042 -2306 6174 -2302
tri 6174 -2306 6202 -2278 sw
rect 6224 -2288 6226 -2274
tri 6224 -2290 6226 -2288 ne
rect 6238 -2292 6269 -2274
rect 6238 -2302 6284 -2292
rect 6351 -2263 6366 -2248
tri 5976 -2327 5988 -2315 ne
rect 5988 -2320 5998 -2315
tri 5998 -2320 6003 -2315 sw
rect 5887 -2524 5902 -2438
rect 5988 -2476 6003 -2320
rect 6042 -2362 6070 -2306
tri 6162 -2324 6180 -2306 ne
rect 6180 -2326 6202 -2306
tri 6202 -2326 6222 -2306 sw
tri 6238 -2320 6256 -2302 ne
rect 6061 -2396 6070 -2362
rect 6104 -2335 6146 -2334
rect 6104 -2369 6109 -2335
rect 6139 -2369 6146 -2335
rect 6104 -2378 6146 -2369
rect 6180 -2335 6222 -2326
rect 6180 -2369 6187 -2335
rect 6217 -2369 6222 -2335
rect 6180 -2374 6222 -2369
rect 6256 -2362 6284 -2302
tri 6329 -2315 6351 -2293 se
rect 6351 -2300 6366 -2292
tri 6351 -2315 6366 -2300 nw
tri 6323 -2321 6329 -2315 se
rect 6329 -2321 6338 -2315
rect 6042 -2406 6070 -2396
tri 6070 -2406 6094 -2382 sw
rect 6042 -2438 6084 -2406
tri 6101 -2414 6102 -2413 sw
rect 6101 -2438 6102 -2414
tri 6104 -2415 6141 -2378 ne
rect 6141 -2406 6146 -2378
tri 6146 -2406 6172 -2380 sw
rect 6256 -2396 6265 -2362
rect 6256 -2406 6284 -2396
rect 6141 -2415 6225 -2406
tri 6141 -2434 6160 -2415 ne
rect 6160 -2434 6225 -2415
rect 6042 -2460 6102 -2438
rect 6224 -2438 6225 -2434
rect 6242 -2438 6284 -2406
rect 6224 -2460 6284 -2438
rect 6130 -2476 6147 -2462
rect 6179 -2476 6196 -2462
rect 6323 -2476 6338 -2321
tri 6338 -2328 6351 -2315 nw
rect 6424 -2396 6439 -2168
rect 6424 -2524 6439 -2438
<< viali >>
rect -233 1800 -201 1814
rect -450 1676 -420 1710
rect -233 1574 -201 1588
rect -14 1676 16 1710
rect -233 1530 -201 1544
rect -450 1406 -420 1440
rect -233 1304 -201 1318
rect -14 1407 16 1440
rect -233 1260 -201 1274
rect -450 1136 -420 1170
rect -233 1034 -201 1048
rect -14 1137 16 1170
rect -233 990 -201 1004
rect -450 866 -420 900
rect -233 764 -201 778
rect -14 867 16 900
rect -233 720 -201 734
rect -450 596 -420 630
rect -233 494 -201 508
rect -14 597 16 630
rect -233 450 -201 464
rect -450 326 -420 360
rect -233 224 -201 238
rect -14 327 16 360
rect -233 180 -201 194
rect -450 56 -420 90
rect -233 -46 -201 -32
rect -14 57 16 90
rect -233 -90 -201 -76
rect -450 -214 -420 -180
rect -233 -316 -201 -302
rect -14 -213 16 -180
rect -233 -360 -201 -346
rect -450 -484 -420 -450
rect -233 -586 -201 -572
rect -14 -483 16 -450
rect -233 -630 -201 -616
rect -450 -754 -420 -720
rect -233 -856 -201 -842
rect -14 -753 16 -720
rect -233 -900 -201 -886
rect -450 -1024 -420 -990
rect -233 -1126 -201 -1112
rect -14 -1023 16 -990
rect -233 -1170 -201 -1156
rect -450 -1294 -420 -1260
rect -233 -1396 -201 -1382
rect -14 -1293 16 -1260
rect -233 -1440 -201 -1426
rect -450 -1564 -420 -1530
rect -233 -1666 -201 -1652
rect -14 -1563 16 -1530
rect -233 -1710 -201 -1696
rect -450 -1834 -420 -1800
rect -233 -1936 -201 -1922
rect -14 -1833 16 -1800
rect -233 -1980 -201 -1966
rect -450 -2104 -420 -2070
rect -233 -2206 -201 -2192
rect -14 -2103 16 -2070
rect -233 -2250 -201 -2236
rect -450 -2374 -420 -2340
rect -233 -2476 -201 -2462
rect -14 -2373 16 -2340
rect 347 1800 379 1814
rect 130 1676 160 1710
rect 347 1574 379 1588
rect 566 1676 596 1710
rect 347 1530 379 1544
rect 130 1406 160 1440
rect 347 1304 379 1318
rect 566 1406 596 1440
rect 347 1260 379 1274
rect 130 1136 160 1170
rect 347 1034 379 1048
rect 566 1136 596 1170
rect 347 990 379 1004
rect 130 866 160 900
rect 347 764 379 778
rect 566 866 596 900
rect 347 720 379 734
rect 130 596 160 630
rect 347 494 379 508
rect 566 596 596 630
rect 347 450 379 464
rect 130 326 160 360
rect 347 224 379 238
rect 566 326 596 360
rect 347 180 379 194
rect 130 56 160 90
rect 347 -46 379 -32
rect 566 56 596 90
rect 347 -90 379 -76
rect 130 -214 160 -180
rect 347 -316 379 -302
rect 566 -214 596 -180
rect 347 -360 379 -346
rect 130 -484 160 -450
rect 347 -586 379 -572
rect 566 -484 596 -450
rect 347 -630 379 -616
rect 130 -754 160 -720
rect 347 -856 379 -842
rect 566 -754 596 -720
rect 347 -900 379 -886
rect 130 -1024 160 -990
rect 347 -1126 379 -1112
rect 566 -1024 596 -990
rect 347 -1170 379 -1156
rect 130 -1294 160 -1260
rect 347 -1396 379 -1382
rect 566 -1294 596 -1260
rect 347 -1440 379 -1426
rect 130 -1564 160 -1530
rect 347 -1666 379 -1652
rect 566 -1564 596 -1530
rect 347 -1710 379 -1696
rect 130 -1834 160 -1800
rect 347 -1936 379 -1922
rect 566 -1834 596 -1800
rect 347 -1980 379 -1966
rect 130 -2104 160 -2070
rect 347 -2206 379 -2192
rect 566 -2104 596 -2070
rect 347 -2250 379 -2236
rect 130 -2374 160 -2340
rect 347 -2476 379 -2462
rect 566 -2374 596 -2340
rect 927 1800 959 1814
rect 710 1676 740 1710
rect 927 1574 959 1588
rect 1146 1677 1176 1710
rect 927 1530 959 1544
rect 710 1406 740 1440
rect 927 1304 959 1318
rect 1146 1407 1176 1440
rect 927 1260 959 1274
rect 710 1136 740 1170
rect 927 1034 959 1048
rect 1146 1137 1176 1170
rect 927 990 959 1004
rect 710 866 740 900
rect 927 764 959 778
rect 1146 867 1176 900
rect 927 720 959 734
rect 710 596 740 630
rect 927 494 959 508
rect 1146 597 1176 630
rect 927 450 959 464
rect 710 326 740 360
rect 927 224 959 238
rect 1146 327 1176 360
rect 927 180 959 194
rect 710 56 740 90
rect 927 -46 959 -32
rect 1146 57 1176 90
rect 927 -90 959 -76
rect 710 -214 740 -180
rect 927 -316 959 -302
rect 1146 -213 1176 -180
rect 927 -360 959 -346
rect 710 -484 740 -450
rect 927 -586 959 -572
rect 1146 -483 1176 -450
rect 927 -630 959 -616
rect 710 -754 740 -720
rect 927 -856 959 -842
rect 1146 -753 1176 -720
rect 927 -900 959 -886
rect 710 -1024 740 -990
rect 927 -1126 959 -1112
rect 1146 -1023 1176 -990
rect 927 -1170 959 -1156
rect 710 -1294 740 -1260
rect 927 -1396 959 -1382
rect 1146 -1293 1176 -1260
rect 927 -1440 959 -1426
rect 710 -1564 740 -1530
rect 927 -1666 959 -1652
rect 1146 -1563 1176 -1530
rect 927 -1710 959 -1696
rect 710 -1834 740 -1800
rect 927 -1936 959 -1922
rect 1146 -1833 1176 -1800
rect 927 -1980 959 -1966
rect 710 -2104 740 -2070
rect 927 -2206 959 -2192
rect 1146 -2103 1176 -2070
rect 927 -2250 959 -2236
rect 710 -2374 740 -2340
rect 927 -2476 959 -2462
rect 1146 -2373 1176 -2340
rect 1507 1800 1539 1814
rect 1290 1676 1320 1710
rect 1507 1574 1539 1588
rect 1726 1676 1756 1710
rect 1507 1530 1539 1544
rect 1290 1406 1320 1440
rect 1507 1304 1539 1318
rect 1726 1406 1756 1440
rect 1507 1260 1539 1274
rect 1290 1136 1320 1170
rect 1507 1034 1539 1048
rect 1726 1136 1756 1170
rect 1507 990 1539 1004
rect 1290 866 1320 900
rect 1507 764 1539 778
rect 1726 866 1756 900
rect 1507 720 1539 734
rect 1290 596 1320 630
rect 1507 494 1539 508
rect 1726 596 1756 630
rect 1507 450 1539 464
rect 1290 326 1320 360
rect 1507 224 1539 238
rect 1726 326 1756 360
rect 1507 180 1539 194
rect 1290 56 1320 90
rect 1507 -46 1539 -32
rect 1726 56 1756 90
rect 1507 -90 1539 -76
rect 1290 -214 1320 -180
rect 1507 -316 1539 -302
rect 1726 -214 1756 -180
rect 1507 -360 1539 -346
rect 1290 -484 1320 -450
rect 1507 -586 1539 -572
rect 1726 -484 1756 -450
rect 1507 -630 1539 -616
rect 1290 -754 1320 -720
rect 1507 -856 1539 -842
rect 1726 -754 1756 -720
rect 1507 -900 1539 -886
rect 1290 -1024 1320 -990
rect 1507 -1126 1539 -1112
rect 1726 -1024 1756 -990
rect 1507 -1170 1539 -1156
rect 1290 -1294 1320 -1260
rect 1507 -1396 1539 -1382
rect 1726 -1294 1756 -1260
rect 1507 -1440 1539 -1426
rect 1290 -1564 1320 -1530
rect 1507 -1666 1539 -1652
rect 1726 -1564 1756 -1530
rect 1507 -1710 1539 -1696
rect 1290 -1834 1320 -1800
rect 1507 -1936 1539 -1922
rect 1726 -1834 1756 -1800
rect 1507 -1980 1539 -1966
rect 1290 -2104 1320 -2070
rect 1507 -2206 1539 -2192
rect 1726 -2104 1756 -2070
rect 1507 -2250 1539 -2236
rect 1290 -2374 1320 -2340
rect 1507 -2476 1539 -2462
rect 1726 -2374 1756 -2340
rect 2087 1800 2119 1814
rect 1870 1676 1900 1710
rect 2087 1574 2119 1588
rect 2306 1677 2336 1710
rect 2087 1530 2119 1544
rect 1870 1406 1900 1440
rect 2087 1304 2119 1318
rect 2306 1407 2336 1440
rect 2087 1260 2119 1274
rect 1870 1136 1900 1170
rect 2087 1034 2119 1048
rect 2306 1137 2336 1170
rect 2087 990 2119 1004
rect 1870 866 1900 900
rect 2087 764 2119 778
rect 2306 867 2336 900
rect 2087 720 2119 734
rect 1870 596 1900 630
rect 2087 494 2119 508
rect 2306 597 2336 630
rect 2087 450 2119 464
rect 1870 326 1900 360
rect 2087 224 2119 238
rect 2306 327 2336 360
rect 2087 180 2119 194
rect 1870 56 1900 90
rect 2087 -46 2119 -32
rect 2306 57 2336 90
rect 2087 -90 2119 -76
rect 1870 -214 1900 -180
rect 2087 -316 2119 -302
rect 2306 -213 2336 -180
rect 2087 -360 2119 -346
rect 1870 -484 1900 -450
rect 2087 -586 2119 -572
rect 2306 -483 2336 -450
rect 2087 -630 2119 -616
rect 1870 -754 1900 -720
rect 2087 -856 2119 -842
rect 2306 -753 2336 -720
rect 2087 -900 2119 -886
rect 1870 -1024 1900 -990
rect 2087 -1126 2119 -1112
rect 2306 -1023 2336 -990
rect 2087 -1170 2119 -1156
rect 1870 -1294 1900 -1260
rect 2087 -1396 2119 -1382
rect 2306 -1293 2336 -1260
rect 2087 -1440 2119 -1426
rect 1870 -1564 1900 -1530
rect 2087 -1666 2119 -1652
rect 2306 -1563 2336 -1530
rect 2087 -1710 2119 -1696
rect 1870 -1834 1900 -1800
rect 2087 -1936 2119 -1922
rect 2306 -1833 2336 -1800
rect 2087 -1980 2119 -1966
rect 1870 -2104 1900 -2070
rect 2087 -2206 2119 -2192
rect 2306 -2103 2336 -2070
rect 2087 -2250 2119 -2236
rect 1870 -2374 1900 -2340
rect 2087 -2476 2119 -2462
rect 2306 -2373 2336 -2340
rect 2667 1800 2699 1814
rect 2450 1676 2480 1710
rect 2667 1574 2699 1588
rect 2886 1676 2916 1710
rect 2667 1530 2699 1544
rect 2450 1406 2480 1440
rect 2667 1304 2699 1318
rect 2886 1406 2916 1440
rect 2667 1260 2699 1274
rect 2450 1136 2480 1170
rect 2667 1034 2699 1048
rect 2886 1136 2916 1170
rect 2667 990 2699 1004
rect 2450 866 2480 900
rect 2667 764 2699 778
rect 2886 866 2916 900
rect 2667 720 2699 734
rect 2450 596 2480 630
rect 2667 494 2699 508
rect 2886 596 2916 630
rect 2667 450 2699 464
rect 2450 326 2480 360
rect 2667 224 2699 238
rect 2886 326 2916 360
rect 2667 180 2699 194
rect 2450 56 2480 90
rect 2667 -46 2699 -32
rect 2886 56 2916 90
rect 2667 -90 2699 -76
rect 2450 -214 2480 -180
rect 2667 -316 2699 -302
rect 2886 -214 2916 -180
rect 2667 -360 2699 -346
rect 2450 -484 2480 -450
rect 2667 -586 2699 -572
rect 2886 -484 2916 -450
rect 2667 -630 2699 -616
rect 2450 -754 2480 -720
rect 2667 -856 2699 -842
rect 2886 -754 2916 -720
rect 2667 -900 2699 -886
rect 2450 -1024 2480 -990
rect 2667 -1126 2699 -1112
rect 2886 -1024 2916 -990
rect 2667 -1170 2699 -1156
rect 2450 -1294 2480 -1260
rect 2667 -1396 2699 -1382
rect 2886 -1294 2916 -1260
rect 2667 -1440 2699 -1426
rect 2450 -1564 2480 -1530
rect 2667 -1666 2699 -1652
rect 2886 -1564 2916 -1530
rect 2667 -1710 2699 -1696
rect 2450 -1834 2480 -1800
rect 2667 -1936 2699 -1922
rect 2886 -1834 2916 -1800
rect 2667 -1980 2699 -1966
rect 2450 -2104 2480 -2070
rect 2667 -2206 2699 -2192
rect 2886 -2104 2916 -2070
rect 2667 -2250 2699 -2236
rect 2450 -2374 2480 -2340
rect 2667 -2476 2699 -2462
rect 2886 -2374 2916 -2340
rect 3247 1800 3279 1814
rect 3030 1676 3060 1710
rect 3247 1574 3279 1588
rect 3466 1677 3496 1710
rect 3247 1530 3279 1544
rect 3030 1406 3060 1440
rect 3247 1304 3279 1318
rect 3466 1407 3496 1440
rect 3247 1260 3279 1274
rect 3030 1136 3060 1170
rect 3247 1034 3279 1048
rect 3466 1137 3496 1170
rect 3247 990 3279 1004
rect 3030 866 3060 900
rect 3247 764 3279 778
rect 3466 867 3496 900
rect 3247 720 3279 734
rect 3030 596 3060 630
rect 3247 494 3279 508
rect 3466 597 3496 630
rect 3247 450 3279 464
rect 3030 326 3060 360
rect 3247 224 3279 238
rect 3466 327 3496 360
rect 3247 180 3279 194
rect 3030 56 3060 90
rect 3247 -46 3279 -32
rect 3466 57 3496 90
rect 3247 -90 3279 -76
rect 3030 -214 3060 -180
rect 3247 -316 3279 -302
rect 3466 -213 3496 -180
rect 3247 -360 3279 -346
rect 3030 -484 3060 -450
rect 3247 -586 3279 -572
rect 3466 -483 3496 -450
rect 3247 -630 3279 -616
rect 3030 -754 3060 -720
rect 3247 -856 3279 -842
rect 3466 -753 3496 -720
rect 3247 -900 3279 -886
rect 3030 -1024 3060 -990
rect 3247 -1126 3279 -1112
rect 3466 -1023 3496 -990
rect 3247 -1170 3279 -1156
rect 3030 -1294 3060 -1260
rect 3247 -1396 3279 -1382
rect 3466 -1293 3496 -1260
rect 3247 -1440 3279 -1426
rect 3030 -1564 3060 -1530
rect 3247 -1666 3279 -1652
rect 3466 -1563 3496 -1530
rect 3247 -1710 3279 -1696
rect 3030 -1834 3060 -1800
rect 3247 -1936 3279 -1922
rect 3466 -1833 3496 -1800
rect 3247 -1980 3279 -1966
rect 3030 -2104 3060 -2070
rect 3247 -2206 3279 -2192
rect 3466 -2103 3496 -2070
rect 3247 -2250 3279 -2236
rect 3030 -2374 3060 -2340
rect 3247 -2476 3279 -2462
rect 3466 -2373 3496 -2340
rect 3827 1800 3859 1814
rect 3610 1676 3640 1710
rect 3827 1574 3859 1588
rect 4046 1676 4076 1710
rect 3827 1530 3859 1544
rect 3610 1406 3640 1440
rect 3827 1304 3859 1318
rect 4046 1406 4076 1440
rect 3827 1260 3859 1274
rect 3610 1136 3640 1170
rect 3827 1034 3859 1048
rect 4046 1136 4076 1170
rect 3827 990 3859 1004
rect 3610 866 3640 900
rect 3827 764 3859 778
rect 4046 866 4076 900
rect 3827 720 3859 734
rect 3610 596 3640 630
rect 3827 494 3859 508
rect 4046 596 4076 630
rect 3827 450 3859 464
rect 3610 326 3640 360
rect 3827 224 3859 238
rect 4046 326 4076 360
rect 3827 180 3859 194
rect 3610 56 3640 90
rect 3827 -46 3859 -32
rect 4046 56 4076 90
rect 3827 -90 3859 -76
rect 3610 -214 3640 -180
rect 3827 -316 3859 -302
rect 4046 -214 4076 -180
rect 3827 -360 3859 -346
rect 3610 -484 3640 -450
rect 3827 -586 3859 -572
rect 4046 -484 4076 -450
rect 3827 -630 3859 -616
rect 3610 -754 3640 -720
rect 3827 -856 3859 -842
rect 4046 -754 4076 -720
rect 3827 -900 3859 -886
rect 3610 -1024 3640 -990
rect 3827 -1126 3859 -1112
rect 4046 -1024 4076 -990
rect 3827 -1170 3859 -1156
rect 3610 -1294 3640 -1260
rect 3827 -1396 3859 -1382
rect 4046 -1294 4076 -1260
rect 3827 -1440 3859 -1426
rect 3610 -1564 3640 -1530
rect 3827 -1666 3859 -1652
rect 4046 -1564 4076 -1530
rect 3827 -1710 3859 -1696
rect 3610 -1834 3640 -1800
rect 3827 -1936 3859 -1922
rect 4046 -1834 4076 -1800
rect 3827 -1980 3859 -1966
rect 3610 -2104 3640 -2070
rect 3827 -2206 3859 -2192
rect 4046 -2104 4076 -2070
rect 3827 -2250 3859 -2236
rect 3610 -2374 3640 -2340
rect 3827 -2476 3859 -2462
rect 4046 -2374 4076 -2340
rect 4407 1800 4439 1814
rect 4190 1676 4220 1710
rect 4407 1574 4439 1588
rect 4626 1677 4656 1710
rect 4407 1530 4439 1544
rect 4190 1406 4220 1440
rect 4407 1304 4439 1318
rect 4626 1407 4656 1440
rect 4407 1260 4439 1274
rect 4190 1136 4220 1170
rect 4407 1034 4439 1048
rect 4626 1137 4656 1170
rect 4407 990 4439 1004
rect 4190 866 4220 900
rect 4407 764 4439 778
rect 4626 867 4656 900
rect 4407 720 4439 734
rect 4190 596 4220 630
rect 4407 494 4439 508
rect 4626 597 4656 630
rect 4407 450 4439 464
rect 4190 326 4220 360
rect 4407 224 4439 238
rect 4626 327 4656 360
rect 4407 180 4439 194
rect 4190 56 4220 90
rect 4407 -46 4439 -32
rect 4626 57 4656 90
rect 4407 -90 4439 -76
rect 4190 -214 4220 -180
rect 4407 -316 4439 -302
rect 4626 -213 4656 -180
rect 4407 -360 4439 -346
rect 4190 -484 4220 -450
rect 4407 -586 4439 -572
rect 4626 -483 4656 -450
rect 4407 -630 4439 -616
rect 4190 -754 4220 -720
rect 4407 -856 4439 -842
rect 4626 -753 4656 -720
rect 4407 -900 4439 -886
rect 4190 -1024 4220 -990
rect 4407 -1126 4439 -1112
rect 4626 -1023 4656 -990
rect 4407 -1170 4439 -1156
rect 4190 -1294 4220 -1260
rect 4407 -1396 4439 -1382
rect 4626 -1293 4656 -1260
rect 4407 -1440 4439 -1426
rect 4190 -1564 4220 -1530
rect 4407 -1666 4439 -1652
rect 4626 -1563 4656 -1530
rect 4407 -1710 4439 -1696
rect 4190 -1834 4220 -1800
rect 4407 -1936 4439 -1922
rect 4626 -1833 4656 -1800
rect 4407 -1980 4439 -1966
rect 4190 -2104 4220 -2070
rect 4407 -2206 4439 -2192
rect 4626 -2103 4656 -2070
rect 4407 -2250 4439 -2236
rect 4190 -2374 4220 -2340
rect 4407 -2476 4439 -2462
rect 4626 -2373 4656 -2340
rect 4987 1800 5019 1814
rect 4770 1676 4800 1710
rect 4987 1574 5019 1588
rect 5206 1676 5236 1710
rect 4987 1530 5019 1544
rect 4770 1406 4800 1440
rect 4987 1304 5019 1318
rect 5206 1406 5236 1440
rect 4987 1260 5019 1274
rect 4770 1136 4800 1170
rect 4987 1034 5019 1048
rect 5206 1136 5236 1170
rect 4987 990 5019 1004
rect 4770 866 4800 900
rect 4987 764 5019 778
rect 5206 866 5236 900
rect 4987 720 5019 734
rect 4770 596 4800 630
rect 4987 494 5019 508
rect 5206 596 5236 630
rect 4987 450 5019 464
rect 4770 326 4800 360
rect 4987 224 5019 238
rect 5206 326 5236 360
rect 4987 180 5019 194
rect 4770 56 4800 90
rect 4987 -46 5019 -32
rect 5206 56 5236 90
rect 4987 -90 5019 -76
rect 4770 -214 4800 -180
rect 4987 -316 5019 -302
rect 5206 -214 5236 -180
rect 4987 -360 5019 -346
rect 4770 -484 4800 -450
rect 4987 -586 5019 -572
rect 5206 -484 5236 -450
rect 4987 -630 5019 -616
rect 4770 -754 4800 -720
rect 4987 -856 5019 -842
rect 5206 -754 5236 -720
rect 4987 -900 5019 -886
rect 4770 -1024 4800 -990
rect 4987 -1126 5019 -1112
rect 5206 -1024 5236 -990
rect 4987 -1170 5019 -1156
rect 4770 -1294 4800 -1260
rect 4987 -1396 5019 -1382
rect 5206 -1294 5236 -1260
rect 4987 -1440 5019 -1426
rect 4770 -1564 4800 -1530
rect 4987 -1666 5019 -1652
rect 5206 -1564 5236 -1530
rect 4987 -1710 5019 -1696
rect 4770 -1834 4800 -1800
rect 4987 -1936 5019 -1922
rect 5206 -1834 5236 -1800
rect 4987 -1980 5019 -1966
rect 4770 -2104 4800 -2070
rect 4987 -2206 5019 -2192
rect 5206 -2104 5236 -2070
rect 4987 -2250 5019 -2236
rect 4770 -2374 4800 -2340
rect 4987 -2476 5019 -2462
rect 5206 -2374 5236 -2340
rect 5567 1800 5599 1814
rect 5350 1676 5380 1710
rect 5567 1574 5599 1588
rect 5786 1677 5816 1710
rect 5567 1530 5599 1544
rect 5350 1406 5380 1440
rect 5567 1304 5599 1318
rect 5786 1407 5816 1440
rect 5567 1260 5599 1274
rect 5350 1136 5380 1170
rect 5567 1034 5599 1048
rect 5786 1137 5816 1170
rect 5567 990 5599 1004
rect 5350 866 5380 900
rect 5567 764 5599 778
rect 5786 867 5816 900
rect 5567 720 5599 734
rect 5350 596 5380 630
rect 5567 494 5599 508
rect 5786 597 5816 630
rect 5567 450 5599 464
rect 5350 326 5380 360
rect 5567 224 5599 238
rect 5786 327 5816 360
rect 5567 180 5599 194
rect 5350 56 5380 90
rect 5567 -46 5599 -32
rect 5786 57 5816 90
rect 5567 -90 5599 -76
rect 5350 -214 5380 -180
rect 5567 -316 5599 -302
rect 5786 -213 5816 -180
rect 5567 -360 5599 -346
rect 5350 -484 5380 -450
rect 5567 -586 5599 -572
rect 5786 -483 5816 -450
rect 5567 -630 5599 -616
rect 5350 -754 5380 -720
rect 5567 -856 5599 -842
rect 5786 -753 5816 -720
rect 5567 -900 5599 -886
rect 5350 -1024 5380 -990
rect 5567 -1126 5599 -1112
rect 5786 -1023 5816 -990
rect 5567 -1170 5599 -1156
rect 5350 -1294 5380 -1260
rect 5567 -1396 5599 -1382
rect 5786 -1293 5816 -1260
rect 5567 -1440 5599 -1426
rect 5350 -1564 5380 -1530
rect 5567 -1666 5599 -1652
rect 5786 -1563 5816 -1530
rect 5567 -1710 5599 -1696
rect 5350 -1834 5380 -1800
rect 5567 -1936 5599 -1922
rect 5786 -1833 5816 -1800
rect 5567 -1980 5599 -1966
rect 5350 -2104 5380 -2070
rect 5567 -2206 5599 -2192
rect 5786 -2103 5816 -2070
rect 5567 -2250 5599 -2236
rect 5350 -2374 5380 -2340
rect 5567 -2476 5599 -2462
rect 5786 -2373 5816 -2340
rect 6147 1800 6179 1814
rect 5930 1676 5960 1710
rect 6147 1574 6179 1588
rect 6366 1676 6396 1710
rect 6147 1530 6179 1544
rect 5930 1406 5960 1440
rect 6147 1304 6179 1318
rect 6366 1406 6396 1440
rect 6147 1260 6179 1274
rect 5930 1136 5960 1170
rect 6147 1034 6179 1048
rect 6366 1136 6396 1170
rect 6147 990 6179 1004
rect 5930 866 5960 900
rect 6147 764 6179 778
rect 6366 866 6396 900
rect 6147 720 6179 734
rect 5930 596 5960 630
rect 6147 494 6179 508
rect 6366 596 6396 630
rect 6147 450 6179 464
rect 5930 326 5960 360
rect 6147 224 6179 238
rect 6366 326 6396 360
rect 6147 180 6179 194
rect 5930 56 5960 90
rect 6147 -46 6179 -32
rect 6366 56 6396 90
rect 6147 -90 6179 -76
rect 5930 -214 5960 -180
rect 6147 -316 6179 -302
rect 6366 -214 6396 -180
rect 6147 -360 6179 -346
rect 5930 -484 5960 -450
rect 6147 -586 6179 -572
rect 6366 -484 6396 -450
rect 6147 -630 6179 -616
rect 5930 -754 5960 -720
rect 6147 -856 6179 -842
rect 6366 -754 6396 -720
rect 6147 -900 6179 -886
rect 5930 -1024 5960 -990
rect 6147 -1126 6179 -1112
rect 6366 -1024 6396 -990
rect 6147 -1170 6179 -1156
rect 5930 -1294 5960 -1260
rect 6147 -1396 6179 -1382
rect 6366 -1294 6396 -1260
rect 6147 -1440 6179 -1426
rect 5930 -1564 5960 -1530
rect 6147 -1666 6179 -1652
rect 6366 -1564 6396 -1530
rect 6147 -1710 6179 -1696
rect 5930 -1834 5960 -1800
rect 6147 -1936 6179 -1922
rect 6366 -1834 6396 -1800
rect 6147 -1980 6179 -1966
rect 5930 -2104 5960 -2070
rect 6147 -2206 6179 -2192
rect 6366 -2104 6396 -2070
rect 6147 -2250 6179 -2236
rect 5930 -2374 5960 -2340
rect 6147 -2476 6179 -2462
rect 6366 -2374 6396 -2340
<< metal1 >>
rect -541 1800 -233 1814
rect -201 1800 347 1814
rect 379 1800 927 1814
rect 959 1800 1507 1814
rect 1539 1800 2087 1814
rect 2119 1800 2667 1814
rect 2699 1800 3247 1814
rect 3279 1800 3827 1814
rect 3859 1800 4407 1814
rect 4439 1800 4987 1814
rect 5019 1800 5567 1814
rect 5599 1800 6147 1814
rect 6179 1800 6439 1814
tri -58 1736 -24 1770 se
rect -24 1736 26 1770
tri 26 1736 60 1770 sw
tri 522 1736 556 1770 se
rect 556 1736 606 1770
tri 606 1736 640 1770 sw
tri 1102 1736 1136 1770 se
rect 1136 1736 1186 1770
tri 1186 1736 1220 1770 sw
tri 1682 1736 1716 1770 se
rect 1716 1736 1766 1770
tri 1766 1736 1800 1770 sw
tri 2262 1736 2296 1770 se
rect 2296 1736 2346 1770
tri 2346 1736 2380 1770 sw
tri 2842 1736 2876 1770 se
rect 2876 1736 2926 1770
tri 2926 1736 2960 1770 sw
tri 3422 1736 3456 1770 se
rect 3456 1736 3506 1770
tri 3506 1736 3540 1770 sw
tri 4002 1736 4036 1770 se
rect 4036 1736 4086 1770
tri 4086 1736 4120 1770 sw
tri 4582 1736 4616 1770 se
rect 4616 1736 4666 1770
tri 4666 1736 4700 1770 sw
tri 5162 1736 5196 1770 se
rect 5196 1736 5246 1770
tri 5246 1736 5280 1770 sw
tri 5742 1736 5776 1770 se
rect 5776 1736 5826 1770
tri 5826 1736 5860 1770 sw
tri 6322 1736 6356 1770 se
rect 6356 1736 6406 1770
tri 6406 1736 6440 1770 sw
tri -84 1710 -58 1736 se
rect -58 1710 -40 1736
tri -40 1710 -14 1736 nw
tri 16 1710 42 1736 ne
rect 42 1710 60 1736
tri 60 1710 86 1736 sw
tri 496 1710 522 1736 se
rect 522 1710 540 1736
tri 540 1710 566 1736 nw
tri 596 1710 622 1736 ne
rect 622 1710 640 1736
tri 640 1710 666 1736 sw
tri 1076 1710 1102 1736 se
rect 1102 1710 1120 1736
tri 1120 1710 1146 1736 nw
tri 1176 1710 1202 1736 ne
rect 1202 1710 1220 1736
tri 1220 1710 1246 1736 sw
tri 1656 1710 1682 1736 se
rect 1682 1710 1700 1736
tri 1700 1710 1726 1736 nw
tri 1756 1710 1782 1736 ne
rect 1782 1710 1800 1736
tri 1800 1710 1826 1736 sw
tri 2236 1710 2262 1736 se
rect 2262 1710 2280 1736
tri 2280 1710 2306 1736 nw
tri 2336 1710 2362 1736 ne
rect 2362 1710 2380 1736
tri 2380 1710 2406 1736 sw
tri 2816 1710 2842 1736 se
rect 2842 1710 2860 1736
tri 2860 1710 2886 1736 nw
tri 2916 1710 2942 1736 ne
rect 2942 1710 2960 1736
tri 2960 1710 2986 1736 sw
tri 3396 1710 3422 1736 se
rect 3422 1710 3440 1736
tri 3440 1710 3466 1736 nw
tri 3496 1710 3522 1736 ne
rect 3522 1710 3540 1736
tri 3540 1710 3566 1736 sw
tri 3976 1710 4002 1736 se
rect 4002 1710 4020 1736
tri 4020 1710 4046 1736 nw
tri 4076 1710 4102 1736 ne
rect 4102 1710 4120 1736
tri 4120 1710 4146 1736 sw
tri 4556 1710 4582 1736 se
rect 4582 1710 4600 1736
tri 4600 1710 4626 1736 nw
tri 4656 1710 4682 1736 ne
rect 4682 1710 4700 1736
tri 4700 1710 4726 1736 sw
tri 5136 1710 5162 1736 se
rect 5162 1710 5180 1736
tri 5180 1710 5206 1736 nw
tri 5236 1710 5262 1736 ne
rect 5262 1710 5280 1736
tri 5280 1710 5306 1736 sw
tri 5716 1710 5742 1736 se
rect 5742 1710 5760 1736
tri 5760 1710 5786 1736 nw
tri 5816 1710 5842 1736 ne
rect 5842 1710 5860 1736
tri 5860 1710 5886 1736 sw
tri 6296 1710 6322 1736 se
rect 6322 1710 6340 1736
tri 6340 1710 6366 1736 nw
tri 6396 1710 6422 1736 ne
rect 6422 1710 6440 1736
tri 6440 1710 6466 1736 sw
rect -541 1676 -450 1710
rect -420 1676 -74 1710
tri -74 1676 -40 1710 nw
tri 42 1676 76 1710 ne
rect 76 1676 130 1710
rect 160 1676 506 1710
tri 506 1676 540 1710 nw
rect 619 1676 710 1710
rect 740 1676 1086 1710
tri 1086 1676 1120 1710 nw
tri 1202 1676 1236 1710 ne
rect 1236 1676 1290 1710
rect 1320 1676 1666 1710
tri 1666 1676 1700 1710 nw
rect 1779 1676 1870 1710
rect 1900 1676 2246 1710
tri 2246 1676 2280 1710 nw
tri 2362 1676 2396 1710 ne
rect 2396 1676 2450 1710
rect 2480 1676 2826 1710
tri 2826 1676 2860 1710 nw
rect 2939 1676 3030 1710
rect 3060 1676 3406 1710
tri 3406 1676 3440 1710 nw
tri 3522 1676 3556 1710 ne
rect 3556 1676 3610 1710
rect 3640 1676 3986 1710
tri 3986 1676 4020 1710 nw
rect 4099 1676 4190 1710
rect 4220 1676 4566 1710
tri 4566 1676 4600 1710 nw
tri 4682 1676 4716 1710 ne
rect 4716 1676 4770 1710
rect 4800 1676 5146 1710
tri 5146 1676 5180 1710 nw
rect 5259 1676 5350 1710
rect 5380 1676 5726 1710
tri 5726 1676 5760 1710 nw
tri 5842 1676 5876 1710 ne
rect 5876 1676 5930 1710
rect 5960 1676 6306 1710
tri 6306 1676 6340 1710 nw
tri 6422 1676 6456 1710 ne
rect 6456 1676 6466 1710
rect -541 1574 -233 1588
rect -201 1574 347 1588
rect 379 1574 927 1588
rect 959 1574 1507 1588
rect 1539 1574 2087 1588
rect 2119 1574 2667 1588
rect 2699 1574 3247 1588
rect 3279 1574 3827 1588
rect 3859 1574 4407 1588
rect 4439 1574 4987 1588
rect 5019 1574 5567 1588
rect 5599 1574 6147 1588
rect 6179 1574 6439 1588
rect -541 1530 -233 1544
rect -201 1530 347 1544
rect 379 1530 927 1544
rect 959 1530 1507 1544
rect 1539 1530 2087 1544
rect 2119 1530 2667 1544
rect 2699 1530 3247 1544
rect 3279 1530 3827 1544
rect 3859 1530 4407 1544
rect 4439 1530 4987 1544
rect 5019 1530 5567 1544
rect 5599 1530 6147 1544
rect 6179 1530 6439 1544
tri -58 1466 -24 1500 se
rect -24 1466 26 1500
tri 26 1466 60 1500 sw
tri 522 1466 556 1500 se
rect 556 1466 606 1500
tri 606 1466 640 1500 sw
tri 1102 1466 1136 1500 se
rect 1136 1466 1186 1500
tri 1186 1466 1220 1500 sw
tri 1682 1466 1716 1500 se
rect 1716 1466 1766 1500
tri 1766 1466 1800 1500 sw
tri 2262 1466 2296 1500 se
rect 2296 1466 2346 1500
tri 2346 1466 2380 1500 sw
tri 2842 1466 2876 1500 se
rect 2876 1466 2926 1500
tri 2926 1466 2960 1500 sw
tri 3422 1466 3456 1500 se
rect 3456 1466 3506 1500
tri 3506 1466 3540 1500 sw
tri 4002 1466 4036 1500 se
rect 4036 1466 4086 1500
tri 4086 1466 4120 1500 sw
tri 4582 1466 4616 1500 se
rect 4616 1466 4666 1500
tri 4666 1466 4700 1500 sw
tri 5162 1466 5196 1500 se
rect 5196 1466 5246 1500
tri 5246 1466 5280 1500 sw
tri 5742 1466 5776 1500 se
rect 5776 1466 5826 1500
tri 5826 1466 5860 1500 sw
tri 6322 1466 6356 1500 se
rect 6356 1466 6406 1500
tri 6406 1466 6440 1500 sw
tri -84 1440 -58 1466 se
rect -58 1440 -40 1466
tri -40 1440 -14 1466 nw
tri 16 1440 42 1466 ne
rect 42 1440 60 1466
tri 60 1440 86 1466 sw
tri 496 1440 522 1466 se
rect 522 1440 540 1466
tri 540 1440 566 1466 nw
tri 596 1440 622 1466 ne
rect 622 1440 640 1466
tri 640 1440 666 1466 sw
tri 1076 1440 1102 1466 se
rect 1102 1440 1120 1466
tri 1120 1440 1146 1466 nw
tri 1176 1440 1202 1466 ne
rect 1202 1440 1220 1466
tri 1220 1440 1246 1466 sw
tri 1656 1440 1682 1466 se
rect 1682 1440 1700 1466
tri 1700 1440 1726 1466 nw
tri 1756 1440 1782 1466 ne
rect 1782 1440 1800 1466
tri 1800 1440 1826 1466 sw
tri 2236 1440 2262 1466 se
rect 2262 1440 2280 1466
tri 2280 1440 2306 1466 nw
tri 2336 1440 2362 1466 ne
rect 2362 1440 2380 1466
tri 2380 1440 2406 1466 sw
tri 2816 1440 2842 1466 se
rect 2842 1440 2860 1466
tri 2860 1440 2886 1466 nw
tri 2916 1440 2942 1466 ne
rect 2942 1440 2960 1466
tri 2960 1440 2986 1466 sw
tri 3396 1440 3422 1466 se
rect 3422 1440 3440 1466
tri 3440 1440 3466 1466 nw
tri 3496 1440 3522 1466 ne
rect 3522 1440 3540 1466
tri 3540 1440 3566 1466 sw
tri 3976 1440 4002 1466 se
rect 4002 1440 4020 1466
tri 4020 1440 4046 1466 nw
tri 4076 1440 4102 1466 ne
rect 4102 1440 4120 1466
tri 4120 1440 4146 1466 sw
tri 4556 1440 4582 1466 se
rect 4582 1440 4600 1466
tri 4600 1440 4626 1466 nw
tri 4656 1440 4682 1466 ne
rect 4682 1440 4700 1466
tri 4700 1440 4726 1466 sw
tri 5136 1440 5162 1466 se
rect 5162 1440 5180 1466
tri 5180 1440 5206 1466 nw
tri 5236 1440 5262 1466 ne
rect 5262 1440 5280 1466
tri 5280 1440 5306 1466 sw
tri 5716 1440 5742 1466 se
rect 5742 1440 5760 1466
tri 5760 1440 5786 1466 nw
tri 5816 1440 5842 1466 ne
rect 5842 1440 5860 1466
tri 5860 1440 5886 1466 sw
tri 6296 1440 6322 1466 se
rect 6322 1440 6340 1466
tri 6340 1440 6366 1466 nw
tri 6396 1440 6422 1466 ne
rect 6422 1440 6440 1466
tri 6440 1440 6466 1466 sw
rect -541 1406 -450 1440
rect -420 1406 -74 1440
tri -74 1406 -40 1440 nw
tri 42 1406 76 1440 ne
rect 76 1406 130 1440
rect 160 1406 506 1440
tri 506 1406 540 1440 nw
rect 619 1406 710 1440
rect 740 1406 1086 1440
tri 1086 1406 1120 1440 nw
tri 1202 1406 1236 1440 ne
rect 1236 1406 1290 1440
rect 1320 1406 1666 1440
tri 1666 1406 1700 1440 nw
rect 1779 1406 1870 1440
rect 1900 1406 2246 1440
tri 2246 1406 2280 1440 nw
tri 2362 1406 2396 1440 ne
rect 2396 1406 2450 1440
rect 2480 1406 2826 1440
tri 2826 1406 2860 1440 nw
rect 2939 1406 3030 1440
rect 3060 1406 3406 1440
tri 3406 1406 3440 1440 nw
tri 3522 1406 3556 1440 ne
rect 3556 1406 3610 1440
rect 3640 1406 3986 1440
tri 3986 1406 4020 1440 nw
rect 4099 1406 4190 1440
rect 4220 1406 4566 1440
tri 4566 1406 4600 1440 nw
tri 4682 1406 4716 1440 ne
rect 4716 1406 4770 1440
rect 4800 1406 5146 1440
tri 5146 1406 5180 1440 nw
rect 5259 1406 5350 1440
rect 5380 1406 5726 1440
tri 5726 1406 5760 1440 nw
tri 5842 1406 5876 1440 ne
rect 5876 1406 5930 1440
rect 5960 1406 6306 1440
tri 6306 1406 6340 1440 nw
tri 6422 1406 6456 1440 ne
rect 6456 1406 6466 1440
rect -541 1304 -233 1318
rect -201 1304 347 1318
rect 379 1304 927 1318
rect 959 1304 1507 1318
rect 1539 1304 2087 1318
rect 2119 1304 2667 1318
rect 2699 1304 3247 1318
rect 3279 1304 3827 1318
rect 3859 1304 4407 1318
rect 4439 1304 4987 1318
rect 5019 1304 5567 1318
rect 5599 1304 6147 1318
rect 6179 1304 6439 1318
rect -541 1260 -233 1274
rect -201 1260 347 1274
rect 379 1260 927 1274
rect 959 1260 1507 1274
rect 1539 1260 2087 1274
rect 2119 1260 2667 1274
rect 2699 1260 3247 1274
rect 3279 1260 3827 1274
rect 3859 1260 4407 1274
rect 4439 1260 4987 1274
rect 5019 1260 5567 1274
rect 5599 1260 6147 1274
rect 6179 1260 6439 1274
tri -58 1196 -24 1230 se
rect -24 1196 26 1230
tri 26 1196 60 1230 sw
tri 522 1196 556 1230 se
rect 556 1196 606 1230
tri 606 1196 640 1230 sw
tri 1102 1196 1136 1230 se
rect 1136 1196 1186 1230
tri 1186 1196 1220 1230 sw
tri 1682 1196 1716 1230 se
rect 1716 1196 1766 1230
tri 1766 1196 1800 1230 sw
tri 2262 1196 2296 1230 se
rect 2296 1196 2346 1230
tri 2346 1196 2380 1230 sw
tri 2842 1196 2876 1230 se
rect 2876 1196 2926 1230
tri 2926 1196 2960 1230 sw
tri 3422 1196 3456 1230 se
rect 3456 1196 3506 1230
tri 3506 1196 3540 1230 sw
tri 4002 1196 4036 1230 se
rect 4036 1196 4086 1230
tri 4086 1196 4120 1230 sw
tri 4582 1196 4616 1230 se
rect 4616 1196 4666 1230
tri 4666 1196 4700 1230 sw
tri 5162 1196 5196 1230 se
rect 5196 1196 5246 1230
tri 5246 1196 5280 1230 sw
tri 5742 1196 5776 1230 se
rect 5776 1196 5826 1230
tri 5826 1196 5860 1230 sw
tri 6322 1196 6356 1230 se
rect 6356 1196 6406 1230
tri 6406 1196 6440 1230 sw
tri -84 1170 -58 1196 se
rect -58 1170 -40 1196
tri -40 1170 -14 1196 nw
tri 16 1170 42 1196 ne
rect 42 1170 60 1196
tri 60 1170 86 1196 sw
tri 496 1170 522 1196 se
rect 522 1170 540 1196
tri 540 1170 566 1196 nw
tri 596 1170 622 1196 ne
rect 622 1170 640 1196
tri 640 1170 666 1196 sw
tri 1076 1170 1102 1196 se
rect 1102 1170 1120 1196
tri 1120 1170 1146 1196 nw
tri 1176 1170 1202 1196 ne
rect 1202 1170 1220 1196
tri 1220 1170 1246 1196 sw
tri 1656 1170 1682 1196 se
rect 1682 1170 1700 1196
tri 1700 1170 1726 1196 nw
tri 1756 1170 1782 1196 ne
rect 1782 1170 1800 1196
tri 1800 1170 1826 1196 sw
tri 2236 1170 2262 1196 se
rect 2262 1170 2280 1196
tri 2280 1170 2306 1196 nw
tri 2336 1170 2362 1196 ne
rect 2362 1170 2380 1196
tri 2380 1170 2406 1196 sw
tri 2816 1170 2842 1196 se
rect 2842 1170 2860 1196
tri 2860 1170 2886 1196 nw
tri 2916 1170 2942 1196 ne
rect 2942 1170 2960 1196
tri 2960 1170 2986 1196 sw
tri 3396 1170 3422 1196 se
rect 3422 1170 3440 1196
tri 3440 1170 3466 1196 nw
tri 3496 1170 3522 1196 ne
rect 3522 1170 3540 1196
tri 3540 1170 3566 1196 sw
tri 3976 1170 4002 1196 se
rect 4002 1170 4020 1196
tri 4020 1170 4046 1196 nw
tri 4076 1170 4102 1196 ne
rect 4102 1170 4120 1196
tri 4120 1170 4146 1196 sw
tri 4556 1170 4582 1196 se
rect 4582 1170 4600 1196
tri 4600 1170 4626 1196 nw
tri 4656 1170 4682 1196 ne
rect 4682 1170 4700 1196
tri 4700 1170 4726 1196 sw
tri 5136 1170 5162 1196 se
rect 5162 1170 5180 1196
tri 5180 1170 5206 1196 nw
tri 5236 1170 5262 1196 ne
rect 5262 1170 5280 1196
tri 5280 1170 5306 1196 sw
tri 5716 1170 5742 1196 se
rect 5742 1170 5760 1196
tri 5760 1170 5786 1196 nw
tri 5816 1170 5842 1196 ne
rect 5842 1170 5860 1196
tri 5860 1170 5886 1196 sw
tri 6296 1170 6322 1196 se
rect 6322 1170 6340 1196
tri 6340 1170 6366 1196 nw
tri 6396 1170 6422 1196 ne
rect 6422 1170 6440 1196
tri 6440 1170 6466 1196 sw
rect -541 1136 -450 1170
rect -420 1136 -74 1170
tri -74 1136 -40 1170 nw
tri 42 1136 76 1170 ne
rect 76 1136 130 1170
rect 160 1136 506 1170
tri 506 1136 540 1170 nw
rect 619 1136 710 1170
rect 740 1136 1086 1170
tri 1086 1136 1120 1170 nw
tri 1202 1136 1236 1170 ne
rect 1236 1136 1290 1170
rect 1320 1136 1666 1170
tri 1666 1136 1700 1170 nw
rect 1779 1136 1870 1170
rect 1900 1136 2246 1170
tri 2246 1136 2280 1170 nw
tri 2362 1136 2396 1170 ne
rect 2396 1136 2450 1170
rect 2480 1136 2826 1170
tri 2826 1136 2860 1170 nw
rect 2939 1136 3030 1170
rect 3060 1136 3406 1170
tri 3406 1136 3440 1170 nw
tri 3522 1136 3556 1170 ne
rect 3556 1136 3610 1170
rect 3640 1136 3986 1170
tri 3986 1136 4020 1170 nw
rect 4099 1136 4190 1170
rect 4220 1136 4566 1170
tri 4566 1136 4600 1170 nw
tri 4682 1136 4716 1170 ne
rect 4716 1136 4770 1170
rect 4800 1136 5146 1170
tri 5146 1136 5180 1170 nw
rect 5259 1136 5350 1170
rect 5380 1136 5726 1170
tri 5726 1136 5760 1170 nw
tri 5842 1136 5876 1170 ne
rect 5876 1136 5930 1170
rect 5960 1136 6306 1170
tri 6306 1136 6340 1170 nw
tri 6422 1136 6456 1170 ne
rect 6456 1136 6466 1170
rect -541 1034 -233 1048
rect -201 1034 347 1048
rect 379 1034 927 1048
rect 959 1034 1507 1048
rect 1539 1034 2087 1048
rect 2119 1034 2667 1048
rect 2699 1034 3247 1048
rect 3279 1034 3827 1048
rect 3859 1034 4407 1048
rect 4439 1034 4987 1048
rect 5019 1034 5567 1048
rect 5599 1034 6147 1048
rect 6179 1034 6439 1048
rect -541 990 -233 1004
rect -201 990 347 1004
rect 379 990 927 1004
rect 959 990 1507 1004
rect 1539 990 2087 1004
rect 2119 990 2667 1004
rect 2699 990 3247 1004
rect 3279 990 3827 1004
rect 3859 990 4407 1004
rect 4439 990 4987 1004
rect 5019 990 5567 1004
rect 5599 990 6147 1004
rect 6179 990 6439 1004
tri -58 926 -24 960 se
rect -24 926 26 960
tri 26 926 60 960 sw
tri 522 926 556 960 se
rect 556 926 606 960
tri 606 926 640 960 sw
tri 1102 926 1136 960 se
rect 1136 926 1186 960
tri 1186 926 1220 960 sw
tri 1682 926 1716 960 se
rect 1716 926 1766 960
tri 1766 926 1800 960 sw
tri 2262 926 2296 960 se
rect 2296 926 2346 960
tri 2346 926 2380 960 sw
tri 2842 926 2876 960 se
rect 2876 926 2926 960
tri 2926 926 2960 960 sw
tri 3422 926 3456 960 se
rect 3456 926 3506 960
tri 3506 926 3540 960 sw
tri 4002 926 4036 960 se
rect 4036 926 4086 960
tri 4086 926 4120 960 sw
tri 4582 926 4616 960 se
rect 4616 926 4666 960
tri 4666 926 4700 960 sw
tri 5162 926 5196 960 se
rect 5196 926 5246 960
tri 5246 926 5280 960 sw
tri 5742 926 5776 960 se
rect 5776 926 5826 960
tri 5826 926 5860 960 sw
tri 6322 926 6356 960 se
rect 6356 926 6406 960
tri 6406 926 6440 960 sw
tri -84 900 -58 926 se
rect -58 900 -40 926
tri -40 900 -14 926 nw
tri 16 900 42 926 ne
rect 42 900 60 926
tri 60 900 86 926 sw
tri 496 900 522 926 se
rect 522 900 540 926
tri 540 900 566 926 nw
tri 596 900 622 926 ne
rect 622 900 640 926
tri 640 900 666 926 sw
tri 1076 900 1102 926 se
rect 1102 900 1120 926
tri 1120 900 1146 926 nw
tri 1176 900 1202 926 ne
rect 1202 900 1220 926
tri 1220 900 1246 926 sw
tri 1656 900 1682 926 se
rect 1682 900 1700 926
tri 1700 900 1726 926 nw
tri 1756 900 1782 926 ne
rect 1782 900 1800 926
tri 1800 900 1826 926 sw
tri 2236 900 2262 926 se
rect 2262 900 2280 926
tri 2280 900 2306 926 nw
tri 2336 900 2362 926 ne
rect 2362 900 2380 926
tri 2380 900 2406 926 sw
tri 2816 900 2842 926 se
rect 2842 900 2860 926
tri 2860 900 2886 926 nw
tri 2916 900 2942 926 ne
rect 2942 900 2960 926
tri 2960 900 2986 926 sw
tri 3396 900 3422 926 se
rect 3422 900 3440 926
tri 3440 900 3466 926 nw
tri 3496 900 3522 926 ne
rect 3522 900 3540 926
tri 3540 900 3566 926 sw
tri 3976 900 4002 926 se
rect 4002 900 4020 926
tri 4020 900 4046 926 nw
tri 4076 900 4102 926 ne
rect 4102 900 4120 926
tri 4120 900 4146 926 sw
tri 4556 900 4582 926 se
rect 4582 900 4600 926
tri 4600 900 4626 926 nw
tri 4656 900 4682 926 ne
rect 4682 900 4700 926
tri 4700 900 4726 926 sw
tri 5136 900 5162 926 se
rect 5162 900 5180 926
tri 5180 900 5206 926 nw
tri 5236 900 5262 926 ne
rect 5262 900 5280 926
tri 5280 900 5306 926 sw
tri 5716 900 5742 926 se
rect 5742 900 5760 926
tri 5760 900 5786 926 nw
tri 5816 900 5842 926 ne
rect 5842 900 5860 926
tri 5860 900 5886 926 sw
tri 6296 900 6322 926 se
rect 6322 900 6340 926
tri 6340 900 6366 926 nw
tri 6396 900 6422 926 ne
rect 6422 900 6440 926
tri 6440 900 6466 926 sw
rect -541 866 -450 900
rect -420 866 -74 900
tri -74 866 -40 900 nw
tri 42 866 76 900 ne
rect 76 866 130 900
rect 160 866 506 900
tri 506 866 540 900 nw
rect 619 866 710 900
rect 740 866 1086 900
tri 1086 866 1120 900 nw
tri 1202 866 1236 900 ne
rect 1236 866 1290 900
rect 1320 866 1666 900
tri 1666 866 1700 900 nw
rect 1779 866 1870 900
rect 1900 866 2246 900
tri 2246 866 2280 900 nw
tri 2362 866 2396 900 ne
rect 2396 866 2450 900
rect 2480 866 2826 900
tri 2826 866 2860 900 nw
rect 2939 866 3030 900
rect 3060 866 3406 900
tri 3406 866 3440 900 nw
tri 3522 866 3556 900 ne
rect 3556 866 3610 900
rect 3640 866 3986 900
tri 3986 866 4020 900 nw
rect 4099 866 4190 900
rect 4220 866 4566 900
tri 4566 866 4600 900 nw
tri 4682 866 4716 900 ne
rect 4716 866 4770 900
rect 4800 866 5146 900
tri 5146 866 5180 900 nw
rect 5259 866 5350 900
rect 5380 866 5726 900
tri 5726 866 5760 900 nw
tri 5842 866 5876 900 ne
rect 5876 866 5930 900
rect 5960 866 6306 900
tri 6306 866 6340 900 nw
tri 6422 866 6456 900 ne
rect 6456 866 6466 900
rect -541 764 -233 778
rect -201 764 347 778
rect 379 764 927 778
rect 959 764 1507 778
rect 1539 764 2087 778
rect 2119 764 2667 778
rect 2699 764 3247 778
rect 3279 764 3827 778
rect 3859 764 4407 778
rect 4439 764 4987 778
rect 5019 764 5567 778
rect 5599 764 6147 778
rect 6179 764 6439 778
rect -541 720 -233 734
rect -201 720 347 734
rect 379 720 927 734
rect 959 720 1507 734
rect 1539 720 2087 734
rect 2119 720 2667 734
rect 2699 720 3247 734
rect 3279 720 3827 734
rect 3859 720 4407 734
rect 4439 720 4987 734
rect 5019 720 5567 734
rect 5599 720 6147 734
rect 6179 720 6439 734
tri -58 656 -24 690 se
rect -24 656 26 690
tri 26 656 60 690 sw
tri 522 656 556 690 se
rect 556 656 606 690
tri 606 656 640 690 sw
tri 1102 656 1136 690 se
rect 1136 656 1186 690
tri 1186 656 1220 690 sw
tri 1682 656 1716 690 se
rect 1716 656 1766 690
tri 1766 656 1800 690 sw
tri 2262 656 2296 690 se
rect 2296 656 2346 690
tri 2346 656 2380 690 sw
tri 2842 656 2876 690 se
rect 2876 656 2926 690
tri 2926 656 2960 690 sw
tri 3422 656 3456 690 se
rect 3456 656 3506 690
tri 3506 656 3540 690 sw
tri 4002 656 4036 690 se
rect 4036 656 4086 690
tri 4086 656 4120 690 sw
tri 4582 656 4616 690 se
rect 4616 656 4666 690
tri 4666 656 4700 690 sw
tri 5162 656 5196 690 se
rect 5196 656 5246 690
tri 5246 656 5280 690 sw
tri 5742 656 5776 690 se
rect 5776 656 5826 690
tri 5826 656 5860 690 sw
tri 6322 656 6356 690 se
rect 6356 656 6406 690
tri 6406 656 6440 690 sw
tri -84 630 -58 656 se
rect -58 630 -40 656
tri -40 630 -14 656 nw
tri 16 630 42 656 ne
rect 42 630 60 656
tri 60 630 86 656 sw
tri 496 630 522 656 se
rect 522 630 540 656
tri 540 630 566 656 nw
tri 596 630 622 656 ne
rect 622 630 640 656
tri 640 630 666 656 sw
tri 1076 630 1102 656 se
rect 1102 630 1120 656
tri 1120 630 1146 656 nw
tri 1176 630 1202 656 ne
rect 1202 630 1220 656
tri 1220 630 1246 656 sw
tri 1656 630 1682 656 se
rect 1682 630 1700 656
tri 1700 630 1726 656 nw
tri 1756 630 1782 656 ne
rect 1782 630 1800 656
tri 1800 630 1826 656 sw
tri 2236 630 2262 656 se
rect 2262 630 2280 656
tri 2280 630 2306 656 nw
tri 2336 630 2362 656 ne
rect 2362 630 2380 656
tri 2380 630 2406 656 sw
tri 2816 630 2842 656 se
rect 2842 630 2860 656
tri 2860 630 2886 656 nw
tri 2916 630 2942 656 ne
rect 2942 630 2960 656
tri 2960 630 2986 656 sw
tri 3396 630 3422 656 se
rect 3422 630 3440 656
tri 3440 630 3466 656 nw
tri 3496 630 3522 656 ne
rect 3522 630 3540 656
tri 3540 630 3566 656 sw
tri 3976 630 4002 656 se
rect 4002 630 4020 656
tri 4020 630 4046 656 nw
tri 4076 630 4102 656 ne
rect 4102 630 4120 656
tri 4120 630 4146 656 sw
tri 4556 630 4582 656 se
rect 4582 630 4600 656
tri 4600 630 4626 656 nw
tri 4656 630 4682 656 ne
rect 4682 630 4700 656
tri 4700 630 4726 656 sw
tri 5136 630 5162 656 se
rect 5162 630 5180 656
tri 5180 630 5206 656 nw
tri 5236 630 5262 656 ne
rect 5262 630 5280 656
tri 5280 630 5306 656 sw
tri 5716 630 5742 656 se
rect 5742 630 5760 656
tri 5760 630 5786 656 nw
tri 5816 630 5842 656 ne
rect 5842 630 5860 656
tri 5860 630 5886 656 sw
tri 6296 630 6322 656 se
rect 6322 630 6340 656
tri 6340 630 6366 656 nw
tri 6396 630 6422 656 ne
rect 6422 630 6440 656
tri 6440 630 6466 656 sw
rect -541 596 -450 630
rect -420 596 -74 630
tri -74 596 -40 630 nw
tri 42 596 76 630 ne
rect 76 596 130 630
rect 160 596 506 630
tri 506 596 540 630 nw
rect 619 596 710 630
rect 740 596 1086 630
tri 1086 596 1120 630 nw
tri 1202 596 1236 630 ne
rect 1236 596 1290 630
rect 1320 596 1666 630
tri 1666 596 1700 630 nw
rect 1779 596 1870 630
rect 1900 596 2246 630
tri 2246 596 2280 630 nw
tri 2362 596 2396 630 ne
rect 2396 596 2450 630
rect 2480 596 2826 630
tri 2826 596 2860 630 nw
rect 2939 596 3030 630
rect 3060 596 3406 630
tri 3406 596 3440 630 nw
tri 3522 596 3556 630 ne
rect 3556 596 3610 630
rect 3640 596 3986 630
tri 3986 596 4020 630 nw
rect 4099 596 4190 630
rect 4220 596 4566 630
tri 4566 596 4600 630 nw
tri 4682 596 4716 630 ne
rect 4716 596 4770 630
rect 4800 596 5146 630
tri 5146 596 5180 630 nw
rect 5259 596 5350 630
rect 5380 596 5726 630
tri 5726 596 5760 630 nw
tri 5842 596 5876 630 ne
rect 5876 596 5930 630
rect 5960 596 6306 630
tri 6306 596 6340 630 nw
tri 6422 596 6456 630 ne
rect 6456 596 6466 630
rect -541 494 -233 508
rect -201 494 347 508
rect 379 494 927 508
rect 959 494 1507 508
rect 1539 494 2087 508
rect 2119 494 2667 508
rect 2699 494 3247 508
rect 3279 494 3827 508
rect 3859 494 4407 508
rect 4439 494 4987 508
rect 5019 494 5567 508
rect 5599 494 6147 508
rect 6179 494 6439 508
rect -541 450 -233 464
rect -201 450 347 464
rect 379 450 927 464
rect 959 450 1507 464
rect 1539 450 2087 464
rect 2119 450 2667 464
rect 2699 450 3247 464
rect 3279 450 3827 464
rect 3859 450 4407 464
rect 4439 450 4987 464
rect 5019 450 5567 464
rect 5599 450 6147 464
rect 6179 450 6439 464
tri -58 386 -24 420 se
rect -24 386 26 420
tri 26 386 60 420 sw
tri 522 386 556 420 se
rect 556 386 606 420
tri 606 386 640 420 sw
tri 1102 386 1136 420 se
rect 1136 386 1186 420
tri 1186 386 1220 420 sw
tri 1682 386 1716 420 se
rect 1716 386 1766 420
tri 1766 386 1800 420 sw
tri 2262 386 2296 420 se
rect 2296 386 2346 420
tri 2346 386 2380 420 sw
tri 2842 386 2876 420 se
rect 2876 386 2926 420
tri 2926 386 2960 420 sw
tri 3422 386 3456 420 se
rect 3456 386 3506 420
tri 3506 386 3540 420 sw
tri 4002 386 4036 420 se
rect 4036 386 4086 420
tri 4086 386 4120 420 sw
tri 4582 386 4616 420 se
rect 4616 386 4666 420
tri 4666 386 4700 420 sw
tri 5162 386 5196 420 se
rect 5196 386 5246 420
tri 5246 386 5280 420 sw
tri 5742 386 5776 420 se
rect 5776 386 5826 420
tri 5826 386 5860 420 sw
tri 6322 386 6356 420 se
rect 6356 386 6406 420
tri 6406 386 6440 420 sw
tri -84 360 -58 386 se
rect -58 360 -40 386
tri -40 360 -14 386 nw
tri 16 360 42 386 ne
rect 42 360 60 386
tri 60 360 86 386 sw
tri 496 360 522 386 se
rect 522 360 540 386
tri 540 360 566 386 nw
tri 596 360 622 386 ne
rect 622 360 640 386
tri 640 360 666 386 sw
tri 1076 360 1102 386 se
rect 1102 360 1120 386
tri 1120 360 1146 386 nw
tri 1176 360 1202 386 ne
rect 1202 360 1220 386
tri 1220 360 1246 386 sw
tri 1656 360 1682 386 se
rect 1682 360 1700 386
tri 1700 360 1726 386 nw
tri 1756 360 1782 386 ne
rect 1782 360 1800 386
tri 1800 360 1826 386 sw
tri 2236 360 2262 386 se
rect 2262 360 2280 386
tri 2280 360 2306 386 nw
tri 2336 360 2362 386 ne
rect 2362 360 2380 386
tri 2380 360 2406 386 sw
tri 2816 360 2842 386 se
rect 2842 360 2860 386
tri 2860 360 2886 386 nw
tri 2916 360 2942 386 ne
rect 2942 360 2960 386
tri 2960 360 2986 386 sw
tri 3396 360 3422 386 se
rect 3422 360 3440 386
tri 3440 360 3466 386 nw
tri 3496 360 3522 386 ne
rect 3522 360 3540 386
tri 3540 360 3566 386 sw
tri 3976 360 4002 386 se
rect 4002 360 4020 386
tri 4020 360 4046 386 nw
tri 4076 360 4102 386 ne
rect 4102 360 4120 386
tri 4120 360 4146 386 sw
tri 4556 360 4582 386 se
rect 4582 360 4600 386
tri 4600 360 4626 386 nw
tri 4656 360 4682 386 ne
rect 4682 360 4700 386
tri 4700 360 4726 386 sw
tri 5136 360 5162 386 se
rect 5162 360 5180 386
tri 5180 360 5206 386 nw
tri 5236 360 5262 386 ne
rect 5262 360 5280 386
tri 5280 360 5306 386 sw
tri 5716 360 5742 386 se
rect 5742 360 5760 386
tri 5760 360 5786 386 nw
tri 5816 360 5842 386 ne
rect 5842 360 5860 386
tri 5860 360 5886 386 sw
tri 6296 360 6322 386 se
rect 6322 360 6340 386
tri 6340 360 6366 386 nw
tri 6396 360 6422 386 ne
rect 6422 360 6440 386
tri 6440 360 6466 386 sw
rect -541 326 -450 360
rect -420 326 -74 360
tri -74 326 -40 360 nw
tri 42 326 76 360 ne
rect 76 326 130 360
rect 160 326 506 360
tri 506 326 540 360 nw
rect 619 326 710 360
rect 740 326 1086 360
tri 1086 326 1120 360 nw
tri 1202 326 1236 360 ne
rect 1236 326 1290 360
rect 1320 326 1666 360
tri 1666 326 1700 360 nw
rect 1779 326 1870 360
rect 1900 326 2246 360
tri 2246 326 2280 360 nw
tri 2362 326 2396 360 ne
rect 2396 326 2450 360
rect 2480 326 2826 360
tri 2826 326 2860 360 nw
rect 2939 326 3030 360
rect 3060 326 3406 360
tri 3406 326 3440 360 nw
tri 3522 326 3556 360 ne
rect 3556 326 3610 360
rect 3640 326 3986 360
tri 3986 326 4020 360 nw
rect 4099 326 4190 360
rect 4220 326 4566 360
tri 4566 326 4600 360 nw
tri 4682 326 4716 360 ne
rect 4716 326 4770 360
rect 4800 326 5146 360
tri 5146 326 5180 360 nw
rect 5259 326 5350 360
rect 5380 326 5726 360
tri 5726 326 5760 360 nw
tri 5842 326 5876 360 ne
rect 5876 326 5930 360
rect 5960 326 6306 360
tri 6306 326 6340 360 nw
tri 6422 326 6456 360 ne
rect 6456 326 6466 360
rect -541 224 -233 238
rect -201 224 347 238
rect 379 224 927 238
rect 959 224 1507 238
rect 1539 224 2087 238
rect 2119 224 2667 238
rect 2699 224 3247 238
rect 3279 224 3827 238
rect 3859 224 4407 238
rect 4439 224 4987 238
rect 5019 224 5567 238
rect 5599 224 6147 238
rect 6179 224 6439 238
rect -541 180 -233 194
rect -201 180 347 194
rect 379 180 927 194
rect 959 180 1507 194
rect 1539 180 2087 194
rect 2119 180 2667 194
rect 2699 180 3247 194
rect 3279 180 3827 194
rect 3859 180 4407 194
rect 4439 180 4987 194
rect 5019 180 5567 194
rect 5599 180 6147 194
rect 6179 180 6439 194
tri -58 116 -24 150 se
rect -24 116 26 150
tri 26 116 60 150 sw
tri 522 116 556 150 se
rect 556 116 606 150
tri 606 116 640 150 sw
tri 1102 116 1136 150 se
rect 1136 116 1186 150
tri 1186 116 1220 150 sw
tri 1682 116 1716 150 se
rect 1716 116 1766 150
tri 1766 116 1800 150 sw
tri 2262 116 2296 150 se
rect 2296 116 2346 150
tri 2346 116 2380 150 sw
tri 2842 116 2876 150 se
rect 2876 116 2926 150
tri 2926 116 2960 150 sw
tri 3422 116 3456 150 se
rect 3456 116 3506 150
tri 3506 116 3540 150 sw
tri 4002 116 4036 150 se
rect 4036 116 4086 150
tri 4086 116 4120 150 sw
tri 4582 116 4616 150 se
rect 4616 116 4666 150
tri 4666 116 4700 150 sw
tri 5162 116 5196 150 se
rect 5196 116 5246 150
tri 5246 116 5280 150 sw
tri 5742 116 5776 150 se
rect 5776 116 5826 150
tri 5826 116 5860 150 sw
tri 6322 116 6356 150 se
rect 6356 116 6406 150
tri 6406 116 6440 150 sw
tri -84 90 -58 116 se
rect -58 90 -40 116
tri -40 90 -14 116 nw
tri 16 90 42 116 ne
rect 42 90 60 116
tri 60 90 86 116 sw
tri 496 90 522 116 se
rect 522 90 540 116
tri 540 90 566 116 nw
tri 596 90 622 116 ne
rect 622 90 640 116
tri 640 90 666 116 sw
tri 1076 90 1102 116 se
rect 1102 90 1120 116
tri 1120 90 1146 116 nw
tri 1176 90 1202 116 ne
rect 1202 90 1220 116
tri 1220 90 1246 116 sw
tri 1656 90 1682 116 se
rect 1682 90 1700 116
tri 1700 90 1726 116 nw
tri 1756 90 1782 116 ne
rect 1782 90 1800 116
tri 1800 90 1826 116 sw
tri 2236 90 2262 116 se
rect 2262 90 2280 116
tri 2280 90 2306 116 nw
tri 2336 90 2362 116 ne
rect 2362 90 2380 116
tri 2380 90 2406 116 sw
tri 2816 90 2842 116 se
rect 2842 90 2860 116
tri 2860 90 2886 116 nw
tri 2916 90 2942 116 ne
rect 2942 90 2960 116
tri 2960 90 2986 116 sw
tri 3396 90 3422 116 se
rect 3422 90 3440 116
tri 3440 90 3466 116 nw
tri 3496 90 3522 116 ne
rect 3522 90 3540 116
tri 3540 90 3566 116 sw
tri 3976 90 4002 116 se
rect 4002 90 4020 116
tri 4020 90 4046 116 nw
tri 4076 90 4102 116 ne
rect 4102 90 4120 116
tri 4120 90 4146 116 sw
tri 4556 90 4582 116 se
rect 4582 90 4600 116
tri 4600 90 4626 116 nw
tri 4656 90 4682 116 ne
rect 4682 90 4700 116
tri 4700 90 4726 116 sw
tri 5136 90 5162 116 se
rect 5162 90 5180 116
tri 5180 90 5206 116 nw
tri 5236 90 5262 116 ne
rect 5262 90 5280 116
tri 5280 90 5306 116 sw
tri 5716 90 5742 116 se
rect 5742 90 5760 116
tri 5760 90 5786 116 nw
tri 5816 90 5842 116 ne
rect 5842 90 5860 116
tri 5860 90 5886 116 sw
tri 6296 90 6322 116 se
rect 6322 90 6340 116
tri 6340 90 6366 116 nw
tri 6396 90 6422 116 ne
rect 6422 90 6440 116
tri 6440 90 6466 116 sw
rect -541 56 -450 90
rect -420 56 -74 90
tri -74 56 -40 90 nw
tri 42 56 76 90 ne
rect 76 56 130 90
rect 160 56 506 90
tri 506 56 540 90 nw
rect 619 56 710 90
rect 740 56 1086 90
tri 1086 56 1120 90 nw
tri 1202 56 1236 90 ne
rect 1236 56 1290 90
rect 1320 56 1666 90
tri 1666 56 1700 90 nw
rect 1779 56 1870 90
rect 1900 56 2246 90
tri 2246 56 2280 90 nw
tri 2362 56 2396 90 ne
rect 2396 56 2450 90
rect 2480 56 2826 90
tri 2826 56 2860 90 nw
rect 2939 56 3030 90
rect 3060 56 3406 90
tri 3406 56 3440 90 nw
tri 3522 56 3556 90 ne
rect 3556 56 3610 90
rect 3640 56 3986 90
tri 3986 56 4020 90 nw
rect 4099 56 4190 90
rect 4220 56 4566 90
tri 4566 56 4600 90 nw
tri 4682 56 4716 90 ne
rect 4716 56 4770 90
rect 4800 56 5146 90
tri 5146 56 5180 90 nw
rect 5259 56 5350 90
rect 5380 56 5726 90
tri 5726 56 5760 90 nw
tri 5842 56 5876 90 ne
rect 5876 56 5930 90
rect 5960 56 6306 90
tri 6306 56 6340 90 nw
tri 6422 56 6456 90 ne
rect 6456 56 6466 90
rect -541 -46 -233 -32
rect -201 -46 347 -32
rect 379 -46 927 -32
rect 959 -46 1507 -32
rect 1539 -46 2087 -32
rect 2119 -46 2667 -32
rect 2699 -46 3247 -32
rect 3279 -46 3827 -32
rect 3859 -46 4407 -32
rect 4439 -46 4987 -32
rect 5019 -46 5567 -32
rect 5599 -46 6147 -32
rect 6179 -46 6439 -32
rect -541 -90 -233 -76
rect -201 -90 347 -76
rect 379 -90 927 -76
rect 959 -90 1507 -76
rect 1539 -90 2087 -76
rect 2119 -90 2667 -76
rect 2699 -90 3247 -76
rect 3279 -90 3827 -76
rect 3859 -90 4407 -76
rect 4439 -90 4987 -76
rect 5019 -90 5567 -76
rect 5599 -90 6147 -76
rect 6179 -90 6439 -76
tri -58 -154 -24 -120 se
rect -24 -154 26 -120
tri 26 -154 60 -120 sw
tri 522 -154 556 -120 se
rect 556 -154 606 -120
tri 606 -154 640 -120 sw
tri 1102 -154 1136 -120 se
rect 1136 -154 1186 -120
tri 1186 -154 1220 -120 sw
tri 1682 -154 1716 -120 se
rect 1716 -154 1766 -120
tri 1766 -154 1800 -120 sw
tri 2262 -154 2296 -120 se
rect 2296 -154 2346 -120
tri 2346 -154 2380 -120 sw
tri 2842 -154 2876 -120 se
rect 2876 -154 2926 -120
tri 2926 -154 2960 -120 sw
tri 3422 -154 3456 -120 se
rect 3456 -154 3506 -120
tri 3506 -154 3540 -120 sw
tri 4002 -154 4036 -120 se
rect 4036 -154 4086 -120
tri 4086 -154 4120 -120 sw
tri 4582 -154 4616 -120 se
rect 4616 -154 4666 -120
tri 4666 -154 4700 -120 sw
tri 5162 -154 5196 -120 se
rect 5196 -154 5246 -120
tri 5246 -154 5280 -120 sw
tri 5742 -154 5776 -120 se
rect 5776 -154 5826 -120
tri 5826 -154 5860 -120 sw
tri 6322 -154 6356 -120 se
rect 6356 -154 6406 -120
tri 6406 -154 6440 -120 sw
tri -84 -180 -58 -154 se
rect -58 -180 -40 -154
tri -40 -180 -14 -154 nw
tri 16 -180 42 -154 ne
rect 42 -180 60 -154
tri 60 -180 86 -154 sw
tri 496 -180 522 -154 se
rect 522 -180 540 -154
tri 540 -180 566 -154 nw
tri 596 -180 622 -154 ne
rect 622 -180 640 -154
tri 640 -180 666 -154 sw
tri 1076 -180 1102 -154 se
rect 1102 -180 1120 -154
tri 1120 -180 1146 -154 nw
tri 1176 -180 1202 -154 ne
rect 1202 -180 1220 -154
tri 1220 -180 1246 -154 sw
tri 1656 -180 1682 -154 se
rect 1682 -180 1700 -154
tri 1700 -180 1726 -154 nw
tri 1756 -180 1782 -154 ne
rect 1782 -180 1800 -154
tri 1800 -180 1826 -154 sw
tri 2236 -180 2262 -154 se
rect 2262 -180 2280 -154
tri 2280 -180 2306 -154 nw
tri 2336 -180 2362 -154 ne
rect 2362 -180 2380 -154
tri 2380 -180 2406 -154 sw
tri 2816 -180 2842 -154 se
rect 2842 -180 2860 -154
tri 2860 -180 2886 -154 nw
tri 2916 -180 2942 -154 ne
rect 2942 -180 2960 -154
tri 2960 -180 2986 -154 sw
tri 3396 -180 3422 -154 se
rect 3422 -180 3440 -154
tri 3440 -180 3466 -154 nw
tri 3496 -180 3522 -154 ne
rect 3522 -180 3540 -154
tri 3540 -180 3566 -154 sw
tri 3976 -180 4002 -154 se
rect 4002 -180 4020 -154
tri 4020 -180 4046 -154 nw
tri 4076 -180 4102 -154 ne
rect 4102 -180 4120 -154
tri 4120 -180 4146 -154 sw
tri 4556 -180 4582 -154 se
rect 4582 -180 4600 -154
tri 4600 -180 4626 -154 nw
tri 4656 -180 4682 -154 ne
rect 4682 -180 4700 -154
tri 4700 -180 4726 -154 sw
tri 5136 -180 5162 -154 se
rect 5162 -180 5180 -154
tri 5180 -180 5206 -154 nw
tri 5236 -180 5262 -154 ne
rect 5262 -180 5280 -154
tri 5280 -180 5306 -154 sw
tri 5716 -180 5742 -154 se
rect 5742 -180 5760 -154
tri 5760 -180 5786 -154 nw
tri 5816 -180 5842 -154 ne
rect 5842 -180 5860 -154
tri 5860 -180 5886 -154 sw
tri 6296 -180 6322 -154 se
rect 6322 -180 6340 -154
tri 6340 -180 6366 -154 nw
tri 6396 -180 6422 -154 ne
rect 6422 -180 6440 -154
tri 6440 -180 6466 -154 sw
rect -541 -214 -450 -180
rect -420 -214 -74 -180
tri -74 -214 -40 -180 nw
tri 42 -214 76 -180 ne
rect 76 -214 130 -180
rect 160 -214 506 -180
tri 506 -214 540 -180 nw
rect 619 -214 710 -180
rect 740 -214 1086 -180
tri 1086 -214 1120 -180 nw
tri 1202 -214 1236 -180 ne
rect 1236 -214 1290 -180
rect 1320 -214 1666 -180
tri 1666 -214 1700 -180 nw
rect 1779 -214 1870 -180
rect 1900 -214 2246 -180
tri 2246 -214 2280 -180 nw
tri 2362 -214 2396 -180 ne
rect 2396 -214 2450 -180
rect 2480 -214 2826 -180
tri 2826 -214 2860 -180 nw
rect 2939 -214 3030 -180
rect 3060 -214 3406 -180
tri 3406 -214 3440 -180 nw
tri 3522 -214 3556 -180 ne
rect 3556 -214 3610 -180
rect 3640 -214 3986 -180
tri 3986 -214 4020 -180 nw
rect 4099 -214 4190 -180
rect 4220 -214 4566 -180
tri 4566 -214 4600 -180 nw
tri 4682 -214 4716 -180 ne
rect 4716 -214 4770 -180
rect 4800 -214 5146 -180
tri 5146 -214 5180 -180 nw
rect 5259 -214 5350 -180
rect 5380 -214 5726 -180
tri 5726 -214 5760 -180 nw
tri 5842 -214 5876 -180 ne
rect 5876 -214 5930 -180
rect 5960 -214 6306 -180
tri 6306 -214 6340 -180 nw
tri 6422 -214 6456 -180 ne
rect 6456 -214 6466 -180
rect -541 -316 -233 -302
rect -201 -316 347 -302
rect 379 -316 927 -302
rect 959 -316 1507 -302
rect 1539 -316 2087 -302
rect 2119 -316 2667 -302
rect 2699 -316 3247 -302
rect 3279 -316 3827 -302
rect 3859 -316 4407 -302
rect 4439 -316 4987 -302
rect 5019 -316 5567 -302
rect 5599 -316 6147 -302
rect 6179 -316 6439 -302
rect -541 -360 -233 -346
rect -201 -360 347 -346
rect 379 -360 927 -346
rect 959 -360 1507 -346
rect 1539 -360 2087 -346
rect 2119 -360 2667 -346
rect 2699 -360 3247 -346
rect 3279 -360 3827 -346
rect 3859 -360 4407 -346
rect 4439 -360 4987 -346
rect 5019 -360 5567 -346
rect 5599 -360 6147 -346
rect 6179 -360 6439 -346
tri -58 -424 -24 -390 se
rect -24 -424 26 -390
tri 26 -424 60 -390 sw
tri 522 -424 556 -390 se
rect 556 -424 606 -390
tri 606 -424 640 -390 sw
tri 1102 -424 1136 -390 se
rect 1136 -424 1186 -390
tri 1186 -424 1220 -390 sw
tri 1682 -424 1716 -390 se
rect 1716 -424 1766 -390
tri 1766 -424 1800 -390 sw
tri 2262 -424 2296 -390 se
rect 2296 -424 2346 -390
tri 2346 -424 2380 -390 sw
tri 2842 -424 2876 -390 se
rect 2876 -424 2926 -390
tri 2926 -424 2960 -390 sw
tri 3422 -424 3456 -390 se
rect 3456 -424 3506 -390
tri 3506 -424 3540 -390 sw
tri 4002 -424 4036 -390 se
rect 4036 -424 4086 -390
tri 4086 -424 4120 -390 sw
tri 4582 -424 4616 -390 se
rect 4616 -424 4666 -390
tri 4666 -424 4700 -390 sw
tri 5162 -424 5196 -390 se
rect 5196 -424 5246 -390
tri 5246 -424 5280 -390 sw
tri 5742 -424 5776 -390 se
rect 5776 -424 5826 -390
tri 5826 -424 5860 -390 sw
tri 6322 -424 6356 -390 se
rect 6356 -424 6406 -390
tri 6406 -424 6440 -390 sw
tri -84 -450 -58 -424 se
rect -58 -450 -40 -424
tri -40 -450 -14 -424 nw
tri 16 -450 42 -424 ne
rect 42 -450 60 -424
tri 60 -450 86 -424 sw
tri 496 -450 522 -424 se
rect 522 -450 540 -424
tri 540 -450 566 -424 nw
tri 596 -450 622 -424 ne
rect 622 -450 640 -424
tri 640 -450 666 -424 sw
tri 1076 -450 1102 -424 se
rect 1102 -450 1120 -424
tri 1120 -450 1146 -424 nw
tri 1176 -450 1202 -424 ne
rect 1202 -450 1220 -424
tri 1220 -450 1246 -424 sw
tri 1656 -450 1682 -424 se
rect 1682 -450 1700 -424
tri 1700 -450 1726 -424 nw
tri 1756 -450 1782 -424 ne
rect 1782 -450 1800 -424
tri 1800 -450 1826 -424 sw
tri 2236 -450 2262 -424 se
rect 2262 -450 2280 -424
tri 2280 -450 2306 -424 nw
tri 2336 -450 2362 -424 ne
rect 2362 -450 2380 -424
tri 2380 -450 2406 -424 sw
tri 2816 -450 2842 -424 se
rect 2842 -450 2860 -424
tri 2860 -450 2886 -424 nw
tri 2916 -450 2942 -424 ne
rect 2942 -450 2960 -424
tri 2960 -450 2986 -424 sw
tri 3396 -450 3422 -424 se
rect 3422 -450 3440 -424
tri 3440 -450 3466 -424 nw
tri 3496 -450 3522 -424 ne
rect 3522 -450 3540 -424
tri 3540 -450 3566 -424 sw
tri 3976 -450 4002 -424 se
rect 4002 -450 4020 -424
tri 4020 -450 4046 -424 nw
tri 4076 -450 4102 -424 ne
rect 4102 -450 4120 -424
tri 4120 -450 4146 -424 sw
tri 4556 -450 4582 -424 se
rect 4582 -450 4600 -424
tri 4600 -450 4626 -424 nw
tri 4656 -450 4682 -424 ne
rect 4682 -450 4700 -424
tri 4700 -450 4726 -424 sw
tri 5136 -450 5162 -424 se
rect 5162 -450 5180 -424
tri 5180 -450 5206 -424 nw
tri 5236 -450 5262 -424 ne
rect 5262 -450 5280 -424
tri 5280 -450 5306 -424 sw
tri 5716 -450 5742 -424 se
rect 5742 -450 5760 -424
tri 5760 -450 5786 -424 nw
tri 5816 -450 5842 -424 ne
rect 5842 -450 5860 -424
tri 5860 -450 5886 -424 sw
tri 6296 -450 6322 -424 se
rect 6322 -450 6340 -424
tri 6340 -450 6366 -424 nw
tri 6396 -450 6422 -424 ne
rect 6422 -450 6440 -424
tri 6440 -450 6466 -424 sw
rect -541 -484 -450 -450
rect -420 -484 -74 -450
tri -74 -484 -40 -450 nw
tri 42 -484 76 -450 ne
rect 76 -484 130 -450
rect 160 -484 506 -450
tri 506 -484 540 -450 nw
rect 619 -484 710 -450
rect 740 -484 1086 -450
tri 1086 -484 1120 -450 nw
tri 1202 -484 1236 -450 ne
rect 1236 -484 1290 -450
rect 1320 -484 1666 -450
tri 1666 -484 1700 -450 nw
rect 1779 -484 1870 -450
rect 1900 -484 2246 -450
tri 2246 -484 2280 -450 nw
tri 2362 -484 2396 -450 ne
rect 2396 -484 2450 -450
rect 2480 -484 2826 -450
tri 2826 -484 2860 -450 nw
rect 2939 -484 3030 -450
rect 3060 -484 3406 -450
tri 3406 -484 3440 -450 nw
tri 3522 -484 3556 -450 ne
rect 3556 -484 3610 -450
rect 3640 -484 3986 -450
tri 3986 -484 4020 -450 nw
rect 4099 -484 4190 -450
rect 4220 -484 4566 -450
tri 4566 -484 4600 -450 nw
tri 4682 -484 4716 -450 ne
rect 4716 -484 4770 -450
rect 4800 -484 5146 -450
tri 5146 -484 5180 -450 nw
rect 5259 -484 5350 -450
rect 5380 -484 5726 -450
tri 5726 -484 5760 -450 nw
tri 5842 -484 5876 -450 ne
rect 5876 -484 5930 -450
rect 5960 -484 6306 -450
tri 6306 -484 6340 -450 nw
tri 6422 -484 6456 -450 ne
rect 6456 -484 6466 -450
rect -541 -586 -233 -572
rect -201 -586 347 -572
rect 379 -586 927 -572
rect 959 -586 1507 -572
rect 1539 -586 2087 -572
rect 2119 -586 2667 -572
rect 2699 -586 3247 -572
rect 3279 -586 3827 -572
rect 3859 -586 4407 -572
rect 4439 -586 4987 -572
rect 5019 -586 5567 -572
rect 5599 -586 6147 -572
rect 6179 -586 6439 -572
rect -541 -630 -233 -616
rect -201 -630 347 -616
rect 379 -630 927 -616
rect 959 -630 1507 -616
rect 1539 -630 2087 -616
rect 2119 -630 2667 -616
rect 2699 -630 3247 -616
rect 3279 -630 3827 -616
rect 3859 -630 4407 -616
rect 4439 -630 4987 -616
rect 5019 -630 5567 -616
rect 5599 -630 6147 -616
rect 6179 -630 6439 -616
tri -58 -694 -24 -660 se
rect -24 -694 26 -660
tri 26 -694 60 -660 sw
tri 522 -694 556 -660 se
rect 556 -694 606 -660
tri 606 -694 640 -660 sw
tri 1102 -694 1136 -660 se
rect 1136 -694 1186 -660
tri 1186 -694 1220 -660 sw
tri 1682 -694 1716 -660 se
rect 1716 -694 1766 -660
tri 1766 -694 1800 -660 sw
tri 2262 -694 2296 -660 se
rect 2296 -694 2346 -660
tri 2346 -694 2380 -660 sw
tri 2842 -694 2876 -660 se
rect 2876 -694 2926 -660
tri 2926 -694 2960 -660 sw
tri 3422 -694 3456 -660 se
rect 3456 -694 3506 -660
tri 3506 -694 3540 -660 sw
tri 4002 -694 4036 -660 se
rect 4036 -694 4086 -660
tri 4086 -694 4120 -660 sw
tri 4582 -694 4616 -660 se
rect 4616 -694 4666 -660
tri 4666 -694 4700 -660 sw
tri 5162 -694 5196 -660 se
rect 5196 -694 5246 -660
tri 5246 -694 5280 -660 sw
tri 5742 -694 5776 -660 se
rect 5776 -694 5826 -660
tri 5826 -694 5860 -660 sw
tri 6322 -694 6356 -660 se
rect 6356 -694 6406 -660
tri 6406 -694 6440 -660 sw
tri -84 -720 -58 -694 se
rect -58 -720 -40 -694
tri -40 -720 -14 -694 nw
tri 16 -720 42 -694 ne
rect 42 -720 60 -694
tri 60 -720 86 -694 sw
tri 496 -720 522 -694 se
rect 522 -720 540 -694
tri 540 -720 566 -694 nw
tri 596 -720 622 -694 ne
rect 622 -720 640 -694
tri 640 -720 666 -694 sw
tri 1076 -720 1102 -694 se
rect 1102 -720 1120 -694
tri 1120 -720 1146 -694 nw
tri 1176 -720 1202 -694 ne
rect 1202 -720 1220 -694
tri 1220 -720 1246 -694 sw
tri 1656 -720 1682 -694 se
rect 1682 -720 1700 -694
tri 1700 -720 1726 -694 nw
tri 1756 -720 1782 -694 ne
rect 1782 -720 1800 -694
tri 1800 -720 1826 -694 sw
tri 2236 -720 2262 -694 se
rect 2262 -720 2280 -694
tri 2280 -720 2306 -694 nw
tri 2336 -720 2362 -694 ne
rect 2362 -720 2380 -694
tri 2380 -720 2406 -694 sw
tri 2816 -720 2842 -694 se
rect 2842 -720 2860 -694
tri 2860 -720 2886 -694 nw
tri 2916 -720 2942 -694 ne
rect 2942 -720 2960 -694
tri 2960 -720 2986 -694 sw
tri 3396 -720 3422 -694 se
rect 3422 -720 3440 -694
tri 3440 -720 3466 -694 nw
tri 3496 -720 3522 -694 ne
rect 3522 -720 3540 -694
tri 3540 -720 3566 -694 sw
tri 3976 -720 4002 -694 se
rect 4002 -720 4020 -694
tri 4020 -720 4046 -694 nw
tri 4076 -720 4102 -694 ne
rect 4102 -720 4120 -694
tri 4120 -720 4146 -694 sw
tri 4556 -720 4582 -694 se
rect 4582 -720 4600 -694
tri 4600 -720 4626 -694 nw
tri 4656 -720 4682 -694 ne
rect 4682 -720 4700 -694
tri 4700 -720 4726 -694 sw
tri 5136 -720 5162 -694 se
rect 5162 -720 5180 -694
tri 5180 -720 5206 -694 nw
tri 5236 -720 5262 -694 ne
rect 5262 -720 5280 -694
tri 5280 -720 5306 -694 sw
tri 5716 -720 5742 -694 se
rect 5742 -720 5760 -694
tri 5760 -720 5786 -694 nw
tri 5816 -720 5842 -694 ne
rect 5842 -720 5860 -694
tri 5860 -720 5886 -694 sw
tri 6296 -720 6322 -694 se
rect 6322 -720 6340 -694
tri 6340 -720 6366 -694 nw
tri 6396 -720 6422 -694 ne
rect 6422 -720 6440 -694
tri 6440 -720 6466 -694 sw
rect -541 -754 -450 -720
rect -420 -754 -74 -720
tri -74 -754 -40 -720 nw
tri 42 -754 76 -720 ne
rect 76 -754 130 -720
rect 160 -754 506 -720
tri 506 -754 540 -720 nw
rect 619 -754 710 -720
rect 740 -754 1086 -720
tri 1086 -754 1120 -720 nw
tri 1202 -754 1236 -720 ne
rect 1236 -754 1290 -720
rect 1320 -754 1666 -720
tri 1666 -754 1700 -720 nw
rect 1779 -754 1870 -720
rect 1900 -754 2246 -720
tri 2246 -754 2280 -720 nw
tri 2362 -754 2396 -720 ne
rect 2396 -754 2450 -720
rect 2480 -754 2826 -720
tri 2826 -754 2860 -720 nw
rect 2939 -754 3030 -720
rect 3060 -754 3406 -720
tri 3406 -754 3440 -720 nw
tri 3522 -754 3556 -720 ne
rect 3556 -754 3610 -720
rect 3640 -754 3986 -720
tri 3986 -754 4020 -720 nw
rect 4099 -754 4190 -720
rect 4220 -754 4566 -720
tri 4566 -754 4600 -720 nw
tri 4682 -754 4716 -720 ne
rect 4716 -754 4770 -720
rect 4800 -754 5146 -720
tri 5146 -754 5180 -720 nw
rect 5259 -754 5350 -720
rect 5380 -754 5726 -720
tri 5726 -754 5760 -720 nw
tri 5842 -754 5876 -720 ne
rect 5876 -754 5930 -720
rect 5960 -754 6306 -720
tri 6306 -754 6340 -720 nw
tri 6422 -754 6456 -720 ne
rect 6456 -754 6466 -720
rect -541 -856 -233 -842
rect -201 -856 347 -842
rect 379 -856 927 -842
rect 959 -856 1507 -842
rect 1539 -856 2087 -842
rect 2119 -856 2667 -842
rect 2699 -856 3247 -842
rect 3279 -856 3827 -842
rect 3859 -856 4407 -842
rect 4439 -856 4987 -842
rect 5019 -856 5567 -842
rect 5599 -856 6147 -842
rect 6179 -856 6439 -842
rect -541 -900 -233 -886
rect -201 -900 347 -886
rect 379 -900 927 -886
rect 959 -900 1507 -886
rect 1539 -900 2087 -886
rect 2119 -900 2667 -886
rect 2699 -900 3247 -886
rect 3279 -900 3827 -886
rect 3859 -900 4407 -886
rect 4439 -900 4987 -886
rect 5019 -900 5567 -886
rect 5599 -900 6147 -886
rect 6179 -900 6439 -886
tri -58 -964 -24 -930 se
rect -24 -964 26 -930
tri 26 -964 60 -930 sw
tri 522 -964 556 -930 se
rect 556 -964 606 -930
tri 606 -964 640 -930 sw
tri 1102 -964 1136 -930 se
rect 1136 -964 1186 -930
tri 1186 -964 1220 -930 sw
tri 1682 -964 1716 -930 se
rect 1716 -964 1766 -930
tri 1766 -964 1800 -930 sw
tri 2262 -964 2296 -930 se
rect 2296 -964 2346 -930
tri 2346 -964 2380 -930 sw
tri 2842 -964 2876 -930 se
rect 2876 -964 2926 -930
tri 2926 -964 2960 -930 sw
tri 3422 -964 3456 -930 se
rect 3456 -964 3506 -930
tri 3506 -964 3540 -930 sw
tri 4002 -964 4036 -930 se
rect 4036 -964 4086 -930
tri 4086 -964 4120 -930 sw
tri 4582 -964 4616 -930 se
rect 4616 -964 4666 -930
tri 4666 -964 4700 -930 sw
tri 5162 -964 5196 -930 se
rect 5196 -964 5246 -930
tri 5246 -964 5280 -930 sw
tri 5742 -964 5776 -930 se
rect 5776 -964 5826 -930
tri 5826 -964 5860 -930 sw
tri 6322 -964 6356 -930 se
rect 6356 -964 6406 -930
tri 6406 -964 6440 -930 sw
tri -84 -990 -58 -964 se
rect -58 -990 -40 -964
tri -40 -990 -14 -964 nw
tri 16 -990 42 -964 ne
rect 42 -990 60 -964
tri 60 -990 86 -964 sw
tri 496 -990 522 -964 se
rect 522 -990 540 -964
tri 540 -990 566 -964 nw
tri 596 -990 622 -964 ne
rect 622 -990 640 -964
tri 640 -990 666 -964 sw
tri 1076 -990 1102 -964 se
rect 1102 -990 1120 -964
tri 1120 -990 1146 -964 nw
tri 1176 -990 1202 -964 ne
rect 1202 -990 1220 -964
tri 1220 -990 1246 -964 sw
tri 1656 -990 1682 -964 se
rect 1682 -990 1700 -964
tri 1700 -990 1726 -964 nw
tri 1756 -990 1782 -964 ne
rect 1782 -990 1800 -964
tri 1800 -990 1826 -964 sw
tri 2236 -990 2262 -964 se
rect 2262 -990 2280 -964
tri 2280 -990 2306 -964 nw
tri 2336 -990 2362 -964 ne
rect 2362 -990 2380 -964
tri 2380 -990 2406 -964 sw
tri 2816 -990 2842 -964 se
rect 2842 -990 2860 -964
tri 2860 -990 2886 -964 nw
tri 2916 -990 2942 -964 ne
rect 2942 -990 2960 -964
tri 2960 -990 2986 -964 sw
tri 3396 -990 3422 -964 se
rect 3422 -990 3440 -964
tri 3440 -990 3466 -964 nw
tri 3496 -990 3522 -964 ne
rect 3522 -990 3540 -964
tri 3540 -990 3566 -964 sw
tri 3976 -990 4002 -964 se
rect 4002 -990 4020 -964
tri 4020 -990 4046 -964 nw
tri 4076 -990 4102 -964 ne
rect 4102 -990 4120 -964
tri 4120 -990 4146 -964 sw
tri 4556 -990 4582 -964 se
rect 4582 -990 4600 -964
tri 4600 -990 4626 -964 nw
tri 4656 -990 4682 -964 ne
rect 4682 -990 4700 -964
tri 4700 -990 4726 -964 sw
tri 5136 -990 5162 -964 se
rect 5162 -990 5180 -964
tri 5180 -990 5206 -964 nw
tri 5236 -990 5262 -964 ne
rect 5262 -990 5280 -964
tri 5280 -990 5306 -964 sw
tri 5716 -990 5742 -964 se
rect 5742 -990 5760 -964
tri 5760 -990 5786 -964 nw
tri 5816 -990 5842 -964 ne
rect 5842 -990 5860 -964
tri 5860 -990 5886 -964 sw
tri 6296 -990 6322 -964 se
rect 6322 -990 6340 -964
tri 6340 -990 6366 -964 nw
tri 6396 -990 6422 -964 ne
rect 6422 -990 6440 -964
tri 6440 -990 6466 -964 sw
rect -541 -1024 -450 -990
rect -420 -1024 -74 -990
tri -74 -1024 -40 -990 nw
tri 42 -1024 76 -990 ne
rect 76 -1024 130 -990
rect 160 -1024 506 -990
tri 506 -1024 540 -990 nw
rect 619 -1024 710 -990
rect 740 -1024 1086 -990
tri 1086 -1024 1120 -990 nw
tri 1202 -1024 1236 -990 ne
rect 1236 -1024 1290 -990
rect 1320 -1024 1666 -990
tri 1666 -1024 1700 -990 nw
rect 1779 -1024 1870 -990
rect 1900 -1024 2246 -990
tri 2246 -1024 2280 -990 nw
tri 2362 -1024 2396 -990 ne
rect 2396 -1024 2450 -990
rect 2480 -1024 2826 -990
tri 2826 -1024 2860 -990 nw
rect 2939 -1024 3030 -990
rect 3060 -1024 3406 -990
tri 3406 -1024 3440 -990 nw
tri 3522 -1024 3556 -990 ne
rect 3556 -1024 3610 -990
rect 3640 -1024 3986 -990
tri 3986 -1024 4020 -990 nw
rect 4099 -1024 4190 -990
rect 4220 -1024 4566 -990
tri 4566 -1024 4600 -990 nw
tri 4682 -1024 4716 -990 ne
rect 4716 -1024 4770 -990
rect 4800 -1024 5146 -990
tri 5146 -1024 5180 -990 nw
rect 5259 -1024 5350 -990
rect 5380 -1024 5726 -990
tri 5726 -1024 5760 -990 nw
tri 5842 -1024 5876 -990 ne
rect 5876 -1024 5930 -990
rect 5960 -1024 6306 -990
tri 6306 -1024 6340 -990 nw
tri 6422 -1024 6456 -990 ne
rect 6456 -1024 6466 -990
rect -541 -1126 -233 -1112
rect -201 -1126 347 -1112
rect 379 -1126 927 -1112
rect 959 -1126 1507 -1112
rect 1539 -1126 2087 -1112
rect 2119 -1126 2667 -1112
rect 2699 -1126 3247 -1112
rect 3279 -1126 3827 -1112
rect 3859 -1126 4407 -1112
rect 4439 -1126 4987 -1112
rect 5019 -1126 5567 -1112
rect 5599 -1126 6147 -1112
rect 6179 -1126 6439 -1112
rect -541 -1170 -233 -1156
rect -201 -1170 347 -1156
rect 379 -1170 927 -1156
rect 959 -1170 1507 -1156
rect 1539 -1170 2087 -1156
rect 2119 -1170 2667 -1156
rect 2699 -1170 3247 -1156
rect 3279 -1170 3827 -1156
rect 3859 -1170 4407 -1156
rect 4439 -1170 4987 -1156
rect 5019 -1170 5567 -1156
rect 5599 -1170 6147 -1156
rect 6179 -1170 6439 -1156
tri -58 -1234 -24 -1200 se
rect -24 -1234 26 -1200
tri 26 -1234 60 -1200 sw
tri 522 -1234 556 -1200 se
rect 556 -1234 606 -1200
tri 606 -1234 640 -1200 sw
tri 1102 -1234 1136 -1200 se
rect 1136 -1234 1186 -1200
tri 1186 -1234 1220 -1200 sw
tri 1682 -1234 1716 -1200 se
rect 1716 -1234 1766 -1200
tri 1766 -1234 1800 -1200 sw
tri 2262 -1234 2296 -1200 se
rect 2296 -1234 2346 -1200
tri 2346 -1234 2380 -1200 sw
tri 2842 -1234 2876 -1200 se
rect 2876 -1234 2926 -1200
tri 2926 -1234 2960 -1200 sw
tri 3422 -1234 3456 -1200 se
rect 3456 -1234 3506 -1200
tri 3506 -1234 3540 -1200 sw
tri 4002 -1234 4036 -1200 se
rect 4036 -1234 4086 -1200
tri 4086 -1234 4120 -1200 sw
tri 4582 -1234 4616 -1200 se
rect 4616 -1234 4666 -1200
tri 4666 -1234 4700 -1200 sw
tri 5162 -1234 5196 -1200 se
rect 5196 -1234 5246 -1200
tri 5246 -1234 5280 -1200 sw
tri 5742 -1234 5776 -1200 se
rect 5776 -1234 5826 -1200
tri 5826 -1234 5860 -1200 sw
tri 6322 -1234 6356 -1200 se
rect 6356 -1234 6406 -1200
tri 6406 -1234 6440 -1200 sw
tri -84 -1260 -58 -1234 se
rect -58 -1260 -40 -1234
tri -40 -1260 -14 -1234 nw
tri 16 -1260 42 -1234 ne
rect 42 -1260 60 -1234
tri 60 -1260 86 -1234 sw
tri 496 -1260 522 -1234 se
rect 522 -1260 540 -1234
tri 540 -1260 566 -1234 nw
tri 596 -1260 622 -1234 ne
rect 622 -1260 640 -1234
tri 640 -1260 666 -1234 sw
tri 1076 -1260 1102 -1234 se
rect 1102 -1260 1120 -1234
tri 1120 -1260 1146 -1234 nw
tri 1176 -1260 1202 -1234 ne
rect 1202 -1260 1220 -1234
tri 1220 -1260 1246 -1234 sw
tri 1656 -1260 1682 -1234 se
rect 1682 -1260 1700 -1234
tri 1700 -1260 1726 -1234 nw
tri 1756 -1260 1782 -1234 ne
rect 1782 -1260 1800 -1234
tri 1800 -1260 1826 -1234 sw
tri 2236 -1260 2262 -1234 se
rect 2262 -1260 2280 -1234
tri 2280 -1260 2306 -1234 nw
tri 2336 -1260 2362 -1234 ne
rect 2362 -1260 2380 -1234
tri 2380 -1260 2406 -1234 sw
tri 2816 -1260 2842 -1234 se
rect 2842 -1260 2860 -1234
tri 2860 -1260 2886 -1234 nw
tri 2916 -1260 2942 -1234 ne
rect 2942 -1260 2960 -1234
tri 2960 -1260 2986 -1234 sw
tri 3396 -1260 3422 -1234 se
rect 3422 -1260 3440 -1234
tri 3440 -1260 3466 -1234 nw
tri 3496 -1260 3522 -1234 ne
rect 3522 -1260 3540 -1234
tri 3540 -1260 3566 -1234 sw
tri 3976 -1260 4002 -1234 se
rect 4002 -1260 4020 -1234
tri 4020 -1260 4046 -1234 nw
tri 4076 -1260 4102 -1234 ne
rect 4102 -1260 4120 -1234
tri 4120 -1260 4146 -1234 sw
tri 4556 -1260 4582 -1234 se
rect 4582 -1260 4600 -1234
tri 4600 -1260 4626 -1234 nw
tri 4656 -1260 4682 -1234 ne
rect 4682 -1260 4700 -1234
tri 4700 -1260 4726 -1234 sw
tri 5136 -1260 5162 -1234 se
rect 5162 -1260 5180 -1234
tri 5180 -1260 5206 -1234 nw
tri 5236 -1260 5262 -1234 ne
rect 5262 -1260 5280 -1234
tri 5280 -1260 5306 -1234 sw
tri 5716 -1260 5742 -1234 se
rect 5742 -1260 5760 -1234
tri 5760 -1260 5786 -1234 nw
tri 5816 -1260 5842 -1234 ne
rect 5842 -1260 5860 -1234
tri 5860 -1260 5886 -1234 sw
tri 6296 -1260 6322 -1234 se
rect 6322 -1260 6340 -1234
tri 6340 -1260 6366 -1234 nw
tri 6396 -1260 6422 -1234 ne
rect 6422 -1260 6440 -1234
tri 6440 -1260 6466 -1234 sw
rect -541 -1294 -450 -1260
rect -420 -1294 -74 -1260
tri -74 -1294 -40 -1260 nw
tri 42 -1294 76 -1260 ne
rect 76 -1294 130 -1260
rect 160 -1294 506 -1260
tri 506 -1294 540 -1260 nw
rect 619 -1294 710 -1260
rect 740 -1294 1086 -1260
tri 1086 -1294 1120 -1260 nw
tri 1202 -1294 1236 -1260 ne
rect 1236 -1294 1290 -1260
rect 1320 -1294 1666 -1260
tri 1666 -1294 1700 -1260 nw
rect 1779 -1294 1870 -1260
rect 1900 -1294 2246 -1260
tri 2246 -1294 2280 -1260 nw
tri 2362 -1294 2396 -1260 ne
rect 2396 -1294 2450 -1260
rect 2480 -1294 2826 -1260
tri 2826 -1294 2860 -1260 nw
rect 2939 -1294 3030 -1260
rect 3060 -1294 3406 -1260
tri 3406 -1294 3440 -1260 nw
tri 3522 -1294 3556 -1260 ne
rect 3556 -1294 3610 -1260
rect 3640 -1294 3986 -1260
tri 3986 -1294 4020 -1260 nw
rect 4099 -1294 4190 -1260
rect 4220 -1294 4566 -1260
tri 4566 -1294 4600 -1260 nw
tri 4682 -1294 4716 -1260 ne
rect 4716 -1294 4770 -1260
rect 4800 -1294 5146 -1260
tri 5146 -1294 5180 -1260 nw
rect 5259 -1294 5350 -1260
rect 5380 -1294 5726 -1260
tri 5726 -1294 5760 -1260 nw
tri 5842 -1294 5876 -1260 ne
rect 5876 -1294 5930 -1260
rect 5960 -1294 6306 -1260
tri 6306 -1294 6340 -1260 nw
tri 6422 -1294 6456 -1260 ne
rect 6456 -1294 6466 -1260
rect -541 -1396 -233 -1382
rect -201 -1396 347 -1382
rect 379 -1396 927 -1382
rect 959 -1396 1507 -1382
rect 1539 -1396 2087 -1382
rect 2119 -1396 2667 -1382
rect 2699 -1396 3247 -1382
rect 3279 -1396 3827 -1382
rect 3859 -1396 4407 -1382
rect 4439 -1396 4987 -1382
rect 5019 -1396 5567 -1382
rect 5599 -1396 6147 -1382
rect 6179 -1396 6439 -1382
rect -541 -1440 -233 -1426
rect -201 -1440 347 -1426
rect 379 -1440 927 -1426
rect 959 -1440 1507 -1426
rect 1539 -1440 2087 -1426
rect 2119 -1440 2667 -1426
rect 2699 -1440 3247 -1426
rect 3279 -1440 3827 -1426
rect 3859 -1440 4407 -1426
rect 4439 -1440 4987 -1426
rect 5019 -1440 5567 -1426
rect 5599 -1440 6147 -1426
rect 6179 -1440 6439 -1426
tri -58 -1504 -24 -1470 se
rect -24 -1504 26 -1470
tri 26 -1504 60 -1470 sw
tri 522 -1504 556 -1470 se
rect 556 -1504 606 -1470
tri 606 -1504 640 -1470 sw
tri 1102 -1504 1136 -1470 se
rect 1136 -1504 1186 -1470
tri 1186 -1504 1220 -1470 sw
tri 1682 -1504 1716 -1470 se
rect 1716 -1504 1766 -1470
tri 1766 -1504 1800 -1470 sw
tri 2262 -1504 2296 -1470 se
rect 2296 -1504 2346 -1470
tri 2346 -1504 2380 -1470 sw
tri 2842 -1504 2876 -1470 se
rect 2876 -1504 2926 -1470
tri 2926 -1504 2960 -1470 sw
tri 3422 -1504 3456 -1470 se
rect 3456 -1504 3506 -1470
tri 3506 -1504 3540 -1470 sw
tri 4002 -1504 4036 -1470 se
rect 4036 -1504 4086 -1470
tri 4086 -1504 4120 -1470 sw
tri 4582 -1504 4616 -1470 se
rect 4616 -1504 4666 -1470
tri 4666 -1504 4700 -1470 sw
tri 5162 -1504 5196 -1470 se
rect 5196 -1504 5246 -1470
tri 5246 -1504 5280 -1470 sw
tri 5742 -1504 5776 -1470 se
rect 5776 -1504 5826 -1470
tri 5826 -1504 5860 -1470 sw
tri 6322 -1504 6356 -1470 se
rect 6356 -1504 6406 -1470
tri 6406 -1504 6440 -1470 sw
tri -84 -1530 -58 -1504 se
rect -58 -1530 -40 -1504
tri -40 -1530 -14 -1504 nw
tri 16 -1530 42 -1504 ne
rect 42 -1530 60 -1504
tri 60 -1530 86 -1504 sw
tri 496 -1530 522 -1504 se
rect 522 -1530 540 -1504
tri 540 -1530 566 -1504 nw
tri 596 -1530 622 -1504 ne
rect 622 -1530 640 -1504
tri 640 -1530 666 -1504 sw
tri 1076 -1530 1102 -1504 se
rect 1102 -1530 1120 -1504
tri 1120 -1530 1146 -1504 nw
tri 1176 -1530 1202 -1504 ne
rect 1202 -1530 1220 -1504
tri 1220 -1530 1246 -1504 sw
tri 1656 -1530 1682 -1504 se
rect 1682 -1530 1700 -1504
tri 1700 -1530 1726 -1504 nw
tri 1756 -1530 1782 -1504 ne
rect 1782 -1530 1800 -1504
tri 1800 -1530 1826 -1504 sw
tri 2236 -1530 2262 -1504 se
rect 2262 -1530 2280 -1504
tri 2280 -1530 2306 -1504 nw
tri 2336 -1530 2362 -1504 ne
rect 2362 -1530 2380 -1504
tri 2380 -1530 2406 -1504 sw
tri 2816 -1530 2842 -1504 se
rect 2842 -1530 2860 -1504
tri 2860 -1530 2886 -1504 nw
tri 2916 -1530 2942 -1504 ne
rect 2942 -1530 2960 -1504
tri 2960 -1530 2986 -1504 sw
tri 3396 -1530 3422 -1504 se
rect 3422 -1530 3440 -1504
tri 3440 -1530 3466 -1504 nw
tri 3496 -1530 3522 -1504 ne
rect 3522 -1530 3540 -1504
tri 3540 -1530 3566 -1504 sw
tri 3976 -1530 4002 -1504 se
rect 4002 -1530 4020 -1504
tri 4020 -1530 4046 -1504 nw
tri 4076 -1530 4102 -1504 ne
rect 4102 -1530 4120 -1504
tri 4120 -1530 4146 -1504 sw
tri 4556 -1530 4582 -1504 se
rect 4582 -1530 4600 -1504
tri 4600 -1530 4626 -1504 nw
tri 4656 -1530 4682 -1504 ne
rect 4682 -1530 4700 -1504
tri 4700 -1530 4726 -1504 sw
tri 5136 -1530 5162 -1504 se
rect 5162 -1530 5180 -1504
tri 5180 -1530 5206 -1504 nw
tri 5236 -1530 5262 -1504 ne
rect 5262 -1530 5280 -1504
tri 5280 -1530 5306 -1504 sw
tri 5716 -1530 5742 -1504 se
rect 5742 -1530 5760 -1504
tri 5760 -1530 5786 -1504 nw
tri 5816 -1530 5842 -1504 ne
rect 5842 -1530 5860 -1504
tri 5860 -1530 5886 -1504 sw
tri 6296 -1530 6322 -1504 se
rect 6322 -1530 6340 -1504
tri 6340 -1530 6366 -1504 nw
tri 6396 -1530 6422 -1504 ne
rect 6422 -1530 6440 -1504
tri 6440 -1530 6466 -1504 sw
rect -541 -1564 -450 -1530
rect -420 -1564 -74 -1530
tri -74 -1564 -40 -1530 nw
tri 42 -1564 76 -1530 ne
rect 76 -1564 130 -1530
rect 160 -1564 506 -1530
tri 506 -1564 540 -1530 nw
rect 619 -1564 710 -1530
rect 740 -1564 1086 -1530
tri 1086 -1564 1120 -1530 nw
tri 1202 -1564 1236 -1530 ne
rect 1236 -1564 1290 -1530
rect 1320 -1564 1666 -1530
tri 1666 -1564 1700 -1530 nw
rect 1779 -1564 1870 -1530
rect 1900 -1564 2246 -1530
tri 2246 -1564 2280 -1530 nw
tri 2362 -1564 2396 -1530 ne
rect 2396 -1564 2450 -1530
rect 2480 -1564 2826 -1530
tri 2826 -1564 2860 -1530 nw
rect 2939 -1564 3030 -1530
rect 3060 -1564 3406 -1530
tri 3406 -1564 3440 -1530 nw
tri 3522 -1564 3556 -1530 ne
rect 3556 -1564 3610 -1530
rect 3640 -1564 3986 -1530
tri 3986 -1564 4020 -1530 nw
rect 4099 -1564 4190 -1530
rect 4220 -1564 4566 -1530
tri 4566 -1564 4600 -1530 nw
tri 4682 -1564 4716 -1530 ne
rect 4716 -1564 4770 -1530
rect 4800 -1564 5146 -1530
tri 5146 -1564 5180 -1530 nw
rect 5259 -1564 5350 -1530
rect 5380 -1564 5726 -1530
tri 5726 -1564 5760 -1530 nw
tri 5842 -1564 5876 -1530 ne
rect 5876 -1564 5930 -1530
rect 5960 -1564 6306 -1530
tri 6306 -1564 6340 -1530 nw
tri 6422 -1564 6456 -1530 ne
rect 6456 -1564 6466 -1530
rect -541 -1666 -233 -1652
rect -201 -1666 347 -1652
rect 379 -1666 927 -1652
rect 959 -1666 1507 -1652
rect 1539 -1666 2087 -1652
rect 2119 -1666 2667 -1652
rect 2699 -1666 3247 -1652
rect 3279 -1666 3827 -1652
rect 3859 -1666 4407 -1652
rect 4439 -1666 4987 -1652
rect 5019 -1666 5567 -1652
rect 5599 -1666 6147 -1652
rect 6179 -1666 6439 -1652
rect -541 -1710 -233 -1696
rect -201 -1710 347 -1696
rect 379 -1710 927 -1696
rect 959 -1710 1507 -1696
rect 1539 -1710 2087 -1696
rect 2119 -1710 2667 -1696
rect 2699 -1710 3247 -1696
rect 3279 -1710 3827 -1696
rect 3859 -1710 4407 -1696
rect 4439 -1710 4987 -1696
rect 5019 -1710 5567 -1696
rect 5599 -1710 6147 -1696
rect 6179 -1710 6439 -1696
tri -58 -1774 -24 -1740 se
rect -24 -1774 26 -1740
tri 26 -1774 60 -1740 sw
tri 522 -1774 556 -1740 se
rect 556 -1774 606 -1740
tri 606 -1774 640 -1740 sw
tri 1102 -1774 1136 -1740 se
rect 1136 -1774 1186 -1740
tri 1186 -1774 1220 -1740 sw
tri 1682 -1774 1716 -1740 se
rect 1716 -1774 1766 -1740
tri 1766 -1774 1800 -1740 sw
tri 2262 -1774 2296 -1740 se
rect 2296 -1774 2346 -1740
tri 2346 -1774 2380 -1740 sw
tri 2842 -1774 2876 -1740 se
rect 2876 -1774 2926 -1740
tri 2926 -1774 2960 -1740 sw
tri 3422 -1774 3456 -1740 se
rect 3456 -1774 3506 -1740
tri 3506 -1774 3540 -1740 sw
tri 4002 -1774 4036 -1740 se
rect 4036 -1774 4086 -1740
tri 4086 -1774 4120 -1740 sw
tri 4582 -1774 4616 -1740 se
rect 4616 -1774 4666 -1740
tri 4666 -1774 4700 -1740 sw
tri 5162 -1774 5196 -1740 se
rect 5196 -1774 5246 -1740
tri 5246 -1774 5280 -1740 sw
tri 5742 -1774 5776 -1740 se
rect 5776 -1774 5826 -1740
tri 5826 -1774 5860 -1740 sw
tri 6322 -1774 6356 -1740 se
rect 6356 -1774 6406 -1740
tri 6406 -1774 6440 -1740 sw
tri -84 -1800 -58 -1774 se
rect -58 -1800 -40 -1774
tri -40 -1800 -14 -1774 nw
tri 16 -1800 42 -1774 ne
rect 42 -1800 60 -1774
tri 60 -1800 86 -1774 sw
tri 496 -1800 522 -1774 se
rect 522 -1800 540 -1774
tri 540 -1800 566 -1774 nw
tri 596 -1800 622 -1774 ne
rect 622 -1800 640 -1774
tri 640 -1800 666 -1774 sw
tri 1076 -1800 1102 -1774 se
rect 1102 -1800 1120 -1774
tri 1120 -1800 1146 -1774 nw
tri 1176 -1800 1202 -1774 ne
rect 1202 -1800 1220 -1774
tri 1220 -1800 1246 -1774 sw
tri 1656 -1800 1682 -1774 se
rect 1682 -1800 1700 -1774
tri 1700 -1800 1726 -1774 nw
tri 1756 -1800 1782 -1774 ne
rect 1782 -1800 1800 -1774
tri 1800 -1800 1826 -1774 sw
tri 2236 -1800 2262 -1774 se
rect 2262 -1800 2280 -1774
tri 2280 -1800 2306 -1774 nw
tri 2336 -1800 2362 -1774 ne
rect 2362 -1800 2380 -1774
tri 2380 -1800 2406 -1774 sw
tri 2816 -1800 2842 -1774 se
rect 2842 -1800 2860 -1774
tri 2860 -1800 2886 -1774 nw
tri 2916 -1800 2942 -1774 ne
rect 2942 -1800 2960 -1774
tri 2960 -1800 2986 -1774 sw
tri 3396 -1800 3422 -1774 se
rect 3422 -1800 3440 -1774
tri 3440 -1800 3466 -1774 nw
tri 3496 -1800 3522 -1774 ne
rect 3522 -1800 3540 -1774
tri 3540 -1800 3566 -1774 sw
tri 3976 -1800 4002 -1774 se
rect 4002 -1800 4020 -1774
tri 4020 -1800 4046 -1774 nw
tri 4076 -1800 4102 -1774 ne
rect 4102 -1800 4120 -1774
tri 4120 -1800 4146 -1774 sw
tri 4556 -1800 4582 -1774 se
rect 4582 -1800 4600 -1774
tri 4600 -1800 4626 -1774 nw
tri 4656 -1800 4682 -1774 ne
rect 4682 -1800 4700 -1774
tri 4700 -1800 4726 -1774 sw
tri 5136 -1800 5162 -1774 se
rect 5162 -1800 5180 -1774
tri 5180 -1800 5206 -1774 nw
tri 5236 -1800 5262 -1774 ne
rect 5262 -1800 5280 -1774
tri 5280 -1800 5306 -1774 sw
tri 5716 -1800 5742 -1774 se
rect 5742 -1800 5760 -1774
tri 5760 -1800 5786 -1774 nw
tri 5816 -1800 5842 -1774 ne
rect 5842 -1800 5860 -1774
tri 5860 -1800 5886 -1774 sw
tri 6296 -1800 6322 -1774 se
rect 6322 -1800 6340 -1774
tri 6340 -1800 6366 -1774 nw
tri 6396 -1800 6422 -1774 ne
rect 6422 -1800 6440 -1774
tri 6440 -1800 6466 -1774 sw
rect -541 -1834 -450 -1800
rect -420 -1834 -74 -1800
tri -74 -1834 -40 -1800 nw
tri 42 -1834 76 -1800 ne
rect 76 -1834 130 -1800
rect 160 -1834 506 -1800
tri 506 -1834 540 -1800 nw
rect 619 -1834 710 -1800
rect 740 -1834 1086 -1800
tri 1086 -1834 1120 -1800 nw
tri 1202 -1834 1236 -1800 ne
rect 1236 -1834 1290 -1800
rect 1320 -1834 1666 -1800
tri 1666 -1834 1700 -1800 nw
rect 1779 -1834 1870 -1800
rect 1900 -1834 2246 -1800
tri 2246 -1834 2280 -1800 nw
tri 2362 -1834 2396 -1800 ne
rect 2396 -1834 2450 -1800
rect 2480 -1834 2826 -1800
tri 2826 -1834 2860 -1800 nw
rect 2939 -1834 3030 -1800
rect 3060 -1834 3406 -1800
tri 3406 -1834 3440 -1800 nw
tri 3522 -1834 3556 -1800 ne
rect 3556 -1834 3610 -1800
rect 3640 -1834 3986 -1800
tri 3986 -1834 4020 -1800 nw
rect 4099 -1834 4190 -1800
rect 4220 -1834 4566 -1800
tri 4566 -1834 4600 -1800 nw
tri 4682 -1834 4716 -1800 ne
rect 4716 -1834 4770 -1800
rect 4800 -1834 5146 -1800
tri 5146 -1834 5180 -1800 nw
rect 5259 -1834 5350 -1800
rect 5380 -1834 5726 -1800
tri 5726 -1834 5760 -1800 nw
tri 5842 -1834 5876 -1800 ne
rect 5876 -1834 5930 -1800
rect 5960 -1834 6306 -1800
tri 6306 -1834 6340 -1800 nw
tri 6422 -1834 6456 -1800 ne
rect 6456 -1834 6466 -1800
rect -541 -1936 -233 -1922
rect -201 -1936 347 -1922
rect 379 -1936 927 -1922
rect 959 -1936 1507 -1922
rect 1539 -1936 2087 -1922
rect 2119 -1936 2667 -1922
rect 2699 -1936 3247 -1922
rect 3279 -1936 3827 -1922
rect 3859 -1936 4407 -1922
rect 4439 -1936 4987 -1922
rect 5019 -1936 5567 -1922
rect 5599 -1936 6147 -1922
rect 6179 -1936 6439 -1922
rect -541 -1980 -233 -1966
rect -201 -1980 347 -1966
rect 379 -1980 927 -1966
rect 959 -1980 1507 -1966
rect 1539 -1980 2087 -1966
rect 2119 -1980 2667 -1966
rect 2699 -1980 3247 -1966
rect 3279 -1980 3827 -1966
rect 3859 -1980 4407 -1966
rect 4439 -1980 4987 -1966
rect 5019 -1980 5567 -1966
rect 5599 -1980 6147 -1966
rect 6179 -1980 6439 -1966
tri -58 -2044 -24 -2010 se
rect -24 -2044 26 -2010
tri 26 -2044 60 -2010 sw
tri 522 -2044 556 -2010 se
rect 556 -2044 606 -2010
tri 606 -2044 640 -2010 sw
tri 1102 -2044 1136 -2010 se
rect 1136 -2044 1186 -2010
tri 1186 -2044 1220 -2010 sw
tri 1682 -2044 1716 -2010 se
rect 1716 -2044 1766 -2010
tri 1766 -2044 1800 -2010 sw
tri 2262 -2044 2296 -2010 se
rect 2296 -2044 2346 -2010
tri 2346 -2044 2380 -2010 sw
tri 2842 -2044 2876 -2010 se
rect 2876 -2044 2926 -2010
tri 2926 -2044 2960 -2010 sw
tri 3422 -2044 3456 -2010 se
rect 3456 -2044 3506 -2010
tri 3506 -2044 3540 -2010 sw
tri 4002 -2044 4036 -2010 se
rect 4036 -2044 4086 -2010
tri 4086 -2044 4120 -2010 sw
tri 4582 -2044 4616 -2010 se
rect 4616 -2044 4666 -2010
tri 4666 -2044 4700 -2010 sw
tri 5162 -2044 5196 -2010 se
rect 5196 -2044 5246 -2010
tri 5246 -2044 5280 -2010 sw
tri 5742 -2044 5776 -2010 se
rect 5776 -2044 5826 -2010
tri 5826 -2044 5860 -2010 sw
tri 6322 -2044 6356 -2010 se
rect 6356 -2044 6406 -2010
tri 6406 -2044 6440 -2010 sw
tri -84 -2070 -58 -2044 se
rect -58 -2070 -40 -2044
tri -40 -2070 -14 -2044 nw
tri 16 -2070 42 -2044 ne
rect 42 -2070 60 -2044
tri 60 -2070 86 -2044 sw
tri 496 -2070 522 -2044 se
rect 522 -2070 540 -2044
tri 540 -2070 566 -2044 nw
tri 596 -2070 622 -2044 ne
rect 622 -2070 640 -2044
tri 640 -2070 666 -2044 sw
tri 1076 -2070 1102 -2044 se
rect 1102 -2070 1120 -2044
tri 1120 -2070 1146 -2044 nw
tri 1176 -2070 1202 -2044 ne
rect 1202 -2070 1220 -2044
tri 1220 -2070 1246 -2044 sw
tri 1656 -2070 1682 -2044 se
rect 1682 -2070 1700 -2044
tri 1700 -2070 1726 -2044 nw
tri 1756 -2070 1782 -2044 ne
rect 1782 -2070 1800 -2044
tri 1800 -2070 1826 -2044 sw
tri 2236 -2070 2262 -2044 se
rect 2262 -2070 2280 -2044
tri 2280 -2070 2306 -2044 nw
tri 2336 -2070 2362 -2044 ne
rect 2362 -2070 2380 -2044
tri 2380 -2070 2406 -2044 sw
tri 2816 -2070 2842 -2044 se
rect 2842 -2070 2860 -2044
tri 2860 -2070 2886 -2044 nw
tri 2916 -2070 2942 -2044 ne
rect 2942 -2070 2960 -2044
tri 2960 -2070 2986 -2044 sw
tri 3396 -2070 3422 -2044 se
rect 3422 -2070 3440 -2044
tri 3440 -2070 3466 -2044 nw
tri 3496 -2070 3522 -2044 ne
rect 3522 -2070 3540 -2044
tri 3540 -2070 3566 -2044 sw
tri 3976 -2070 4002 -2044 se
rect 4002 -2070 4020 -2044
tri 4020 -2070 4046 -2044 nw
tri 4076 -2070 4102 -2044 ne
rect 4102 -2070 4120 -2044
tri 4120 -2070 4146 -2044 sw
tri 4556 -2070 4582 -2044 se
rect 4582 -2070 4600 -2044
tri 4600 -2070 4626 -2044 nw
tri 4656 -2070 4682 -2044 ne
rect 4682 -2070 4700 -2044
tri 4700 -2070 4726 -2044 sw
tri 5136 -2070 5162 -2044 se
rect 5162 -2070 5180 -2044
tri 5180 -2070 5206 -2044 nw
tri 5236 -2070 5262 -2044 ne
rect 5262 -2070 5280 -2044
tri 5280 -2070 5306 -2044 sw
tri 5716 -2070 5742 -2044 se
rect 5742 -2070 5760 -2044
tri 5760 -2070 5786 -2044 nw
tri 5816 -2070 5842 -2044 ne
rect 5842 -2070 5860 -2044
tri 5860 -2070 5886 -2044 sw
tri 6296 -2070 6322 -2044 se
rect 6322 -2070 6340 -2044
tri 6340 -2070 6366 -2044 nw
tri 6396 -2070 6422 -2044 ne
rect 6422 -2070 6440 -2044
tri 6440 -2070 6466 -2044 sw
rect -541 -2104 -450 -2070
rect -420 -2104 -74 -2070
tri -74 -2104 -40 -2070 nw
tri 42 -2104 76 -2070 ne
rect 76 -2104 130 -2070
rect 160 -2104 506 -2070
tri 506 -2104 540 -2070 nw
rect 619 -2104 710 -2070
rect 740 -2104 1086 -2070
tri 1086 -2104 1120 -2070 nw
tri 1202 -2104 1236 -2070 ne
rect 1236 -2104 1290 -2070
rect 1320 -2104 1666 -2070
tri 1666 -2104 1700 -2070 nw
rect 1779 -2104 1870 -2070
rect 1900 -2104 2246 -2070
tri 2246 -2104 2280 -2070 nw
tri 2362 -2104 2396 -2070 ne
rect 2396 -2104 2450 -2070
rect 2480 -2104 2826 -2070
tri 2826 -2104 2860 -2070 nw
rect 2939 -2104 3030 -2070
rect 3060 -2104 3406 -2070
tri 3406 -2104 3440 -2070 nw
tri 3522 -2104 3556 -2070 ne
rect 3556 -2104 3610 -2070
rect 3640 -2104 3986 -2070
tri 3986 -2104 4020 -2070 nw
rect 4099 -2104 4190 -2070
rect 4220 -2104 4566 -2070
tri 4566 -2104 4600 -2070 nw
tri 4682 -2104 4716 -2070 ne
rect 4716 -2104 4770 -2070
rect 4800 -2104 5146 -2070
tri 5146 -2104 5180 -2070 nw
rect 5259 -2104 5350 -2070
rect 5380 -2104 5726 -2070
tri 5726 -2104 5760 -2070 nw
tri 5842 -2104 5876 -2070 ne
rect 5876 -2104 5930 -2070
rect 5960 -2104 6306 -2070
tri 6306 -2104 6340 -2070 nw
tri 6422 -2104 6456 -2070 ne
rect 6456 -2104 6466 -2070
rect -541 -2206 -233 -2192
rect -201 -2206 347 -2192
rect 379 -2206 927 -2192
rect 959 -2206 1507 -2192
rect 1539 -2206 2087 -2192
rect 2119 -2206 2667 -2192
rect 2699 -2206 3247 -2192
rect 3279 -2206 3827 -2192
rect 3859 -2206 4407 -2192
rect 4439 -2206 4987 -2192
rect 5019 -2206 5567 -2192
rect 5599 -2206 6147 -2192
rect 6179 -2206 6439 -2192
rect -541 -2250 -233 -2236
rect -201 -2250 347 -2236
rect 379 -2250 927 -2236
rect 959 -2250 1507 -2236
rect 1539 -2250 2087 -2236
rect 2119 -2250 2667 -2236
rect 2699 -2250 3247 -2236
rect 3279 -2250 3827 -2236
rect 3859 -2250 4407 -2236
rect 4439 -2250 4987 -2236
rect 5019 -2250 5567 -2236
rect 5599 -2250 6147 -2236
rect 6179 -2250 6439 -2236
tri -58 -2314 -24 -2280 se
rect -24 -2314 26 -2280
tri 26 -2314 60 -2280 sw
tri 522 -2314 556 -2280 se
rect 556 -2314 606 -2280
tri 606 -2314 640 -2280 sw
tri 1102 -2314 1136 -2280 se
rect 1136 -2314 1186 -2280
tri 1186 -2314 1220 -2280 sw
tri 1682 -2314 1716 -2280 se
rect 1716 -2314 1766 -2280
tri 1766 -2314 1800 -2280 sw
tri 2262 -2314 2296 -2280 se
rect 2296 -2314 2346 -2280
tri 2346 -2314 2380 -2280 sw
tri 2842 -2314 2876 -2280 se
rect 2876 -2314 2926 -2280
tri 2926 -2314 2960 -2280 sw
tri 3422 -2314 3456 -2280 se
rect 3456 -2314 3506 -2280
tri 3506 -2314 3540 -2280 sw
tri 4002 -2314 4036 -2280 se
rect 4036 -2314 4086 -2280
tri 4086 -2314 4120 -2280 sw
tri 4582 -2314 4616 -2280 se
rect 4616 -2314 4666 -2280
tri 4666 -2314 4700 -2280 sw
tri 5162 -2314 5196 -2280 se
rect 5196 -2314 5246 -2280
tri 5246 -2314 5280 -2280 sw
tri 5742 -2314 5776 -2280 se
rect 5776 -2314 5826 -2280
tri 5826 -2314 5860 -2280 sw
tri 6322 -2314 6356 -2280 se
rect 6356 -2314 6406 -2280
tri 6406 -2314 6440 -2280 sw
tri -84 -2340 -58 -2314 se
rect -58 -2340 -40 -2314
tri -40 -2340 -14 -2314 nw
tri 16 -2340 42 -2314 ne
rect 42 -2340 60 -2314
tri 60 -2340 86 -2314 sw
tri 496 -2340 522 -2314 se
rect 522 -2340 540 -2314
tri 540 -2340 566 -2314 nw
tri 596 -2340 622 -2314 ne
rect 622 -2340 640 -2314
tri 640 -2340 666 -2314 sw
tri 1076 -2340 1102 -2314 se
rect 1102 -2340 1120 -2314
tri 1120 -2340 1146 -2314 nw
tri 1176 -2340 1202 -2314 ne
rect 1202 -2340 1220 -2314
tri 1220 -2340 1246 -2314 sw
tri 1656 -2340 1682 -2314 se
rect 1682 -2340 1700 -2314
tri 1700 -2340 1726 -2314 nw
tri 1756 -2340 1782 -2314 ne
rect 1782 -2340 1800 -2314
tri 1800 -2340 1826 -2314 sw
tri 2236 -2340 2262 -2314 se
rect 2262 -2340 2280 -2314
tri 2280 -2340 2306 -2314 nw
tri 2336 -2340 2362 -2314 ne
rect 2362 -2340 2380 -2314
tri 2380 -2340 2406 -2314 sw
tri 2816 -2340 2842 -2314 se
rect 2842 -2340 2860 -2314
tri 2860 -2340 2886 -2314 nw
tri 2916 -2340 2942 -2314 ne
rect 2942 -2340 2960 -2314
tri 2960 -2340 2986 -2314 sw
tri 3396 -2340 3422 -2314 se
rect 3422 -2340 3440 -2314
tri 3440 -2340 3466 -2314 nw
tri 3496 -2340 3522 -2314 ne
rect 3522 -2340 3540 -2314
tri 3540 -2340 3566 -2314 sw
tri 3976 -2340 4002 -2314 se
rect 4002 -2340 4020 -2314
tri 4020 -2340 4046 -2314 nw
tri 4076 -2340 4102 -2314 ne
rect 4102 -2340 4120 -2314
tri 4120 -2340 4146 -2314 sw
tri 4556 -2340 4582 -2314 se
rect 4582 -2340 4600 -2314
tri 4600 -2340 4626 -2314 nw
tri 4656 -2340 4682 -2314 ne
rect 4682 -2340 4700 -2314
tri 4700 -2340 4726 -2314 sw
tri 5136 -2340 5162 -2314 se
rect 5162 -2340 5180 -2314
tri 5180 -2340 5206 -2314 nw
tri 5236 -2340 5262 -2314 ne
rect 5262 -2340 5280 -2314
tri 5280 -2340 5306 -2314 sw
tri 5716 -2340 5742 -2314 se
rect 5742 -2340 5760 -2314
tri 5760 -2340 5786 -2314 nw
tri 5816 -2340 5842 -2314 ne
rect 5842 -2340 5860 -2314
tri 5860 -2340 5886 -2314 sw
tri 6296 -2340 6322 -2314 se
rect 6322 -2340 6340 -2314
tri 6340 -2340 6366 -2314 nw
tri 6396 -2340 6422 -2314 ne
rect 6422 -2340 6440 -2314
tri 6440 -2340 6466 -2314 sw
rect -541 -2374 -450 -2340
rect -420 -2374 -74 -2340
tri -74 -2374 -40 -2340 nw
tri 42 -2374 76 -2340 ne
rect 76 -2374 130 -2340
rect 160 -2374 506 -2340
tri 506 -2374 540 -2340 nw
rect 619 -2374 710 -2340
rect 740 -2374 1086 -2340
tri 1086 -2374 1120 -2340 nw
tri 1202 -2374 1236 -2340 ne
rect 1236 -2374 1290 -2340
rect 1320 -2374 1666 -2340
tri 1666 -2374 1700 -2340 nw
rect 1779 -2374 1870 -2340
rect 1900 -2374 2246 -2340
tri 2246 -2374 2280 -2340 nw
tri 2362 -2374 2396 -2340 ne
rect 2396 -2374 2450 -2340
rect 2480 -2374 2826 -2340
tri 2826 -2374 2860 -2340 nw
rect 2939 -2374 3030 -2340
rect 3060 -2374 3406 -2340
tri 3406 -2374 3440 -2340 nw
tri 3522 -2374 3556 -2340 ne
rect 3556 -2374 3610 -2340
rect 3640 -2374 3986 -2340
tri 3986 -2374 4020 -2340 nw
rect 4099 -2374 4190 -2340
rect 4220 -2374 4566 -2340
tri 4566 -2374 4600 -2340 nw
tri 4682 -2374 4716 -2340 ne
rect 4716 -2374 4770 -2340
rect 4800 -2374 5146 -2340
tri 5146 -2374 5180 -2340 nw
rect 5259 -2374 5350 -2340
rect 5380 -2374 5726 -2340
tri 5726 -2374 5760 -2340 nw
tri 5842 -2374 5876 -2340 ne
rect 5876 -2374 5930 -2340
rect 5960 -2374 6306 -2340
tri 6306 -2374 6340 -2340 nw
tri 6422 -2374 6456 -2340 ne
rect 6456 -2374 6466 -2340
rect -541 -2476 -233 -2462
rect -201 -2476 347 -2462
rect 379 -2476 927 -2462
rect 959 -2476 1507 -2462
rect 1539 -2476 2087 -2462
rect 2119 -2476 2667 -2462
rect 2699 -2476 3247 -2462
rect 3279 -2476 3827 -2462
rect 3859 -2476 4407 -2462
rect 4439 -2476 4987 -2462
rect 5019 -2476 5567 -2462
rect 5599 -2476 6147 -2462
rect 6179 -2476 6439 -2462
<< via1 >>
rect -14 1676 16 1710
rect 566 1676 596 1710
rect 1146 1677 1176 1710
rect 1146 1676 1176 1677
rect 1726 1676 1756 1710
rect 2306 1677 2336 1710
rect 2306 1676 2336 1677
rect 2886 1676 2916 1710
rect 3466 1677 3496 1710
rect 3466 1676 3496 1677
rect 4046 1676 4076 1710
rect 4626 1677 4656 1710
rect 4626 1676 4656 1677
rect 5206 1676 5236 1710
rect 5786 1677 5816 1710
rect 5786 1676 5816 1677
rect 6366 1676 6396 1710
rect -14 1407 16 1440
rect -14 1406 16 1407
rect 566 1406 596 1440
rect 1146 1407 1176 1440
rect 1146 1406 1176 1407
rect 1726 1406 1756 1440
rect 2306 1407 2336 1440
rect 2306 1406 2336 1407
rect 2886 1406 2916 1440
rect 3466 1407 3496 1440
rect 3466 1406 3496 1407
rect 4046 1406 4076 1440
rect 4626 1407 4656 1440
rect 4626 1406 4656 1407
rect 5206 1406 5236 1440
rect 5786 1407 5816 1440
rect 5786 1406 5816 1407
rect 6366 1406 6396 1440
rect -14 1137 16 1170
rect -14 1136 16 1137
rect 566 1136 596 1170
rect 1146 1137 1176 1170
rect 1146 1136 1176 1137
rect 1726 1136 1756 1170
rect 2306 1137 2336 1170
rect 2306 1136 2336 1137
rect 2886 1136 2916 1170
rect 3466 1137 3496 1170
rect 3466 1136 3496 1137
rect 4046 1136 4076 1170
rect 4626 1137 4656 1170
rect 4626 1136 4656 1137
rect 5206 1136 5236 1170
rect 5786 1137 5816 1170
rect 5786 1136 5816 1137
rect 6366 1136 6396 1170
rect -14 867 16 900
rect -14 866 16 867
rect 566 866 596 900
rect 1146 867 1176 900
rect 1146 866 1176 867
rect 1726 866 1756 900
rect 2306 867 2336 900
rect 2306 866 2336 867
rect 2886 866 2916 900
rect 3466 867 3496 900
rect 3466 866 3496 867
rect 4046 866 4076 900
rect 4626 867 4656 900
rect 4626 866 4656 867
rect 5206 866 5236 900
rect 5786 867 5816 900
rect 5786 866 5816 867
rect 6366 866 6396 900
rect -14 597 16 630
rect -14 596 16 597
rect 566 596 596 630
rect 1146 597 1176 630
rect 1146 596 1176 597
rect 1726 596 1756 630
rect 2306 597 2336 630
rect 2306 596 2336 597
rect 2886 596 2916 630
rect 3466 597 3496 630
rect 3466 596 3496 597
rect 4046 596 4076 630
rect 4626 597 4656 630
rect 4626 596 4656 597
rect 5206 596 5236 630
rect 5786 597 5816 630
rect 5786 596 5816 597
rect 6366 596 6396 630
rect -14 327 16 360
rect -14 326 16 327
rect 566 326 596 360
rect 1146 327 1176 360
rect 1146 326 1176 327
rect 1726 326 1756 360
rect 2306 327 2336 360
rect 2306 326 2336 327
rect 2886 326 2916 360
rect 3466 327 3496 360
rect 3466 326 3496 327
rect 4046 326 4076 360
rect 4626 327 4656 360
rect 4626 326 4656 327
rect 5206 326 5236 360
rect 5786 327 5816 360
rect 5786 326 5816 327
rect 6366 326 6396 360
rect -14 57 16 90
rect -14 56 16 57
rect 566 56 596 90
rect 1146 57 1176 90
rect 1146 56 1176 57
rect 1726 56 1756 90
rect 2306 57 2336 90
rect 2306 56 2336 57
rect 2886 56 2916 90
rect 3466 57 3496 90
rect 3466 56 3496 57
rect 4046 56 4076 90
rect 4626 57 4656 90
rect 4626 56 4656 57
rect 5206 56 5236 90
rect 5786 57 5816 90
rect 5786 56 5816 57
rect 6366 56 6396 90
rect -14 -213 16 -180
rect -14 -214 16 -213
rect 566 -214 596 -180
rect 1146 -213 1176 -180
rect 1146 -214 1176 -213
rect 1726 -214 1756 -180
rect 2306 -213 2336 -180
rect 2306 -214 2336 -213
rect 2886 -214 2916 -180
rect 3466 -213 3496 -180
rect 3466 -214 3496 -213
rect 4046 -214 4076 -180
rect 4626 -213 4656 -180
rect 4626 -214 4656 -213
rect 5206 -214 5236 -180
rect 5786 -213 5816 -180
rect 5786 -214 5816 -213
rect 6366 -214 6396 -180
rect -14 -483 16 -450
rect -14 -484 16 -483
rect 566 -484 596 -450
rect 1146 -483 1176 -450
rect 1146 -484 1176 -483
rect 1726 -484 1756 -450
rect 2306 -483 2336 -450
rect 2306 -484 2336 -483
rect 2886 -484 2916 -450
rect 3466 -483 3496 -450
rect 3466 -484 3496 -483
rect 4046 -484 4076 -450
rect 4626 -483 4656 -450
rect 4626 -484 4656 -483
rect 5206 -484 5236 -450
rect 5786 -483 5816 -450
rect 5786 -484 5816 -483
rect 6366 -484 6396 -450
rect -14 -753 16 -720
rect -14 -754 16 -753
rect 566 -754 596 -720
rect 1146 -753 1176 -720
rect 1146 -754 1176 -753
rect 1726 -754 1756 -720
rect 2306 -753 2336 -720
rect 2306 -754 2336 -753
rect 2886 -754 2916 -720
rect 3466 -753 3496 -720
rect 3466 -754 3496 -753
rect 4046 -754 4076 -720
rect 4626 -753 4656 -720
rect 4626 -754 4656 -753
rect 5206 -754 5236 -720
rect 5786 -753 5816 -720
rect 5786 -754 5816 -753
rect 6366 -754 6396 -720
rect -14 -1023 16 -990
rect -14 -1024 16 -1023
rect 566 -1024 596 -990
rect 1146 -1023 1176 -990
rect 1146 -1024 1176 -1023
rect 1726 -1024 1756 -990
rect 2306 -1023 2336 -990
rect 2306 -1024 2336 -1023
rect 2886 -1024 2916 -990
rect 3466 -1023 3496 -990
rect 3466 -1024 3496 -1023
rect 4046 -1024 4076 -990
rect 4626 -1023 4656 -990
rect 4626 -1024 4656 -1023
rect 5206 -1024 5236 -990
rect 5786 -1023 5816 -990
rect 5786 -1024 5816 -1023
rect 6366 -1024 6396 -990
rect -14 -1293 16 -1260
rect -14 -1294 16 -1293
rect 566 -1294 596 -1260
rect 1146 -1293 1176 -1260
rect 1146 -1294 1176 -1293
rect 1726 -1294 1756 -1260
rect 2306 -1293 2336 -1260
rect 2306 -1294 2336 -1293
rect 2886 -1294 2916 -1260
rect 3466 -1293 3496 -1260
rect 3466 -1294 3496 -1293
rect 4046 -1294 4076 -1260
rect 4626 -1293 4656 -1260
rect 4626 -1294 4656 -1293
rect 5206 -1294 5236 -1260
rect 5786 -1293 5816 -1260
rect 5786 -1294 5816 -1293
rect 6366 -1294 6396 -1260
rect -14 -1563 16 -1530
rect -14 -1564 16 -1563
rect 566 -1564 596 -1530
rect 1146 -1563 1176 -1530
rect 1146 -1564 1176 -1563
rect 1726 -1564 1756 -1530
rect 2306 -1563 2336 -1530
rect 2306 -1564 2336 -1563
rect 2886 -1564 2916 -1530
rect 3466 -1563 3496 -1530
rect 3466 -1564 3496 -1563
rect 4046 -1564 4076 -1530
rect 4626 -1563 4656 -1530
rect 4626 -1564 4656 -1563
rect 5206 -1564 5236 -1530
rect 5786 -1563 5816 -1530
rect 5786 -1564 5816 -1563
rect 6366 -1564 6396 -1530
rect -14 -1833 16 -1800
rect -14 -1834 16 -1833
rect 566 -1834 596 -1800
rect 1146 -1833 1176 -1800
rect 1146 -1834 1176 -1833
rect 1726 -1834 1756 -1800
rect 2306 -1833 2336 -1800
rect 2306 -1834 2336 -1833
rect 2886 -1834 2916 -1800
rect 3466 -1833 3496 -1800
rect 3466 -1834 3496 -1833
rect 4046 -1834 4076 -1800
rect 4626 -1833 4656 -1800
rect 4626 -1834 4656 -1833
rect 5206 -1834 5236 -1800
rect 5786 -1833 5816 -1800
rect 5786 -1834 5816 -1833
rect 6366 -1834 6396 -1800
rect -14 -2103 16 -2070
rect -14 -2104 16 -2103
rect 566 -2104 596 -2070
rect 1146 -2103 1176 -2070
rect 1146 -2104 1176 -2103
rect 1726 -2104 1756 -2070
rect 2306 -2103 2336 -2070
rect 2306 -2104 2336 -2103
rect 2886 -2104 2916 -2070
rect 3466 -2103 3496 -2070
rect 3466 -2104 3496 -2103
rect 4046 -2104 4076 -2070
rect 4626 -2103 4656 -2070
rect 4626 -2104 4656 -2103
rect 5206 -2104 5236 -2070
rect 5786 -2103 5816 -2070
rect 5786 -2104 5816 -2103
rect 6366 -2104 6396 -2070
rect -14 -2373 16 -2340
rect -14 -2374 16 -2373
rect 566 -2374 596 -2340
rect 1146 -2373 1176 -2340
rect 1146 -2374 1176 -2373
rect 1726 -2374 1756 -2340
rect 2306 -2373 2336 -2340
rect 2306 -2374 2336 -2373
rect 2886 -2374 2916 -2340
rect 3466 -2373 3496 -2340
rect 3466 -2374 3496 -2373
rect 4046 -2374 4076 -2340
rect 4626 -2373 4656 -2340
rect 4626 -2374 4656 -2373
rect 5206 -2374 5236 -2340
rect 5786 -2373 5816 -2340
rect 5786 -2374 5816 -2373
rect 6366 -2374 6396 -2340
<< metal2 >>
rect -541 1676 -14 1710
rect 16 1676 566 1710
rect 596 1676 1146 1710
rect 1176 1676 1726 1710
rect 1756 1676 2306 1710
rect 2336 1676 2886 1710
rect 2916 1676 3466 1710
rect 3496 1676 4046 1710
rect 4076 1676 4626 1710
rect 4656 1676 5206 1710
rect 5236 1676 5786 1710
rect 5816 1676 6366 1710
rect 6396 1676 6466 1710
rect -541 1406 -14 1440
rect 16 1406 566 1440
rect 596 1406 1146 1440
rect 1176 1406 1726 1440
rect 1756 1406 2306 1440
rect 2336 1406 2886 1440
rect 2916 1406 3466 1440
rect 3496 1406 4046 1440
rect 4076 1406 4626 1440
rect 4656 1406 5206 1440
rect 5236 1406 5786 1440
rect 5816 1406 6366 1440
rect 6396 1406 6466 1440
rect -541 1136 -14 1170
rect 16 1136 566 1170
rect 596 1136 1146 1170
rect 1176 1136 1726 1170
rect 1756 1136 2306 1170
rect 2336 1136 2886 1170
rect 2916 1136 3466 1170
rect 3496 1136 4046 1170
rect 4076 1136 4626 1170
rect 4656 1136 5206 1170
rect 5236 1136 5786 1170
rect 5816 1136 6366 1170
rect 6396 1136 6466 1170
rect -541 866 -14 900
rect 16 866 566 900
rect 596 866 1146 900
rect 1176 866 1726 900
rect 1756 866 2306 900
rect 2336 866 2886 900
rect 2916 866 3466 900
rect 3496 866 4046 900
rect 4076 866 4626 900
rect 4656 866 5206 900
rect 5236 866 5786 900
rect 5816 866 6366 900
rect 6396 866 6466 900
rect -541 596 -14 630
rect 16 596 566 630
rect 596 596 1146 630
rect 1176 596 1726 630
rect 1756 596 2306 630
rect 2336 596 2886 630
rect 2916 596 3466 630
rect 3496 596 4046 630
rect 4076 596 4626 630
rect 4656 596 5206 630
rect 5236 596 5786 630
rect 5816 596 6366 630
rect 6396 596 6466 630
rect -541 326 -14 360
rect 16 326 566 360
rect 596 326 1146 360
rect 1176 326 1726 360
rect 1756 326 2306 360
rect 2336 326 2886 360
rect 2916 326 3466 360
rect 3496 326 4046 360
rect 4076 326 4626 360
rect 4656 326 5206 360
rect 5236 326 5786 360
rect 5816 326 6366 360
rect 6396 326 6466 360
rect -541 56 -14 90
rect 16 56 566 90
rect 596 56 1146 90
rect 1176 56 1726 90
rect 1756 56 2306 90
rect 2336 56 2886 90
rect 2916 56 3466 90
rect 3496 56 4046 90
rect 4076 56 4626 90
rect 4656 56 5206 90
rect 5236 56 5786 90
rect 5816 56 6366 90
rect 6396 56 6466 90
rect -541 -214 -14 -180
rect 16 -214 566 -180
rect 596 -214 1146 -180
rect 1176 -214 1726 -180
rect 1756 -214 2306 -180
rect 2336 -214 2886 -180
rect 2916 -214 3466 -180
rect 3496 -214 4046 -180
rect 4076 -214 4626 -180
rect 4656 -214 5206 -180
rect 5236 -214 5786 -180
rect 5816 -214 6366 -180
rect 6396 -214 6466 -180
rect -541 -484 -14 -450
rect 16 -484 566 -450
rect 596 -484 1146 -450
rect 1176 -484 1726 -450
rect 1756 -484 2306 -450
rect 2336 -484 2886 -450
rect 2916 -484 3466 -450
rect 3496 -484 4046 -450
rect 4076 -484 4626 -450
rect 4656 -484 5206 -450
rect 5236 -484 5786 -450
rect 5816 -484 6366 -450
rect 6396 -484 6466 -450
rect -541 -754 -14 -720
rect 16 -754 566 -720
rect 596 -754 1146 -720
rect 1176 -754 1726 -720
rect 1756 -754 2306 -720
rect 2336 -754 2886 -720
rect 2916 -754 3466 -720
rect 3496 -754 4046 -720
rect 4076 -754 4626 -720
rect 4656 -754 5206 -720
rect 5236 -754 5786 -720
rect 5816 -754 6366 -720
rect 6396 -754 6466 -720
rect -541 -1024 -14 -990
rect 16 -1024 566 -990
rect 596 -1024 1146 -990
rect 1176 -1024 1726 -990
rect 1756 -1024 2306 -990
rect 2336 -1024 2886 -990
rect 2916 -1024 3466 -990
rect 3496 -1024 4046 -990
rect 4076 -1024 4626 -990
rect 4656 -1024 5206 -990
rect 5236 -1024 5786 -990
rect 5816 -1024 6366 -990
rect 6396 -1024 6466 -990
rect -541 -1294 -14 -1260
rect 16 -1294 566 -1260
rect 596 -1294 1146 -1260
rect 1176 -1294 1726 -1260
rect 1756 -1294 2306 -1260
rect 2336 -1294 2886 -1260
rect 2916 -1294 3466 -1260
rect 3496 -1294 4046 -1260
rect 4076 -1294 4626 -1260
rect 4656 -1294 5206 -1260
rect 5236 -1294 5786 -1260
rect 5816 -1294 6366 -1260
rect 6396 -1294 6466 -1260
rect -541 -1564 -14 -1530
rect 16 -1564 566 -1530
rect 596 -1564 1146 -1530
rect 1176 -1564 1726 -1530
rect 1756 -1564 2306 -1530
rect 2336 -1564 2886 -1530
rect 2916 -1564 3466 -1530
rect 3496 -1564 4046 -1530
rect 4076 -1564 4626 -1530
rect 4656 -1564 5206 -1530
rect 5236 -1564 5786 -1530
rect 5816 -1564 6366 -1530
rect 6396 -1564 6466 -1530
rect -541 -1834 -14 -1800
rect 16 -1834 566 -1800
rect 596 -1834 1146 -1800
rect 1176 -1834 1726 -1800
rect 1756 -1834 2306 -1800
rect 2336 -1834 2886 -1800
rect 2916 -1834 3466 -1800
rect 3496 -1834 4046 -1800
rect 4076 -1834 4626 -1800
rect 4656 -1834 5206 -1800
rect 5236 -1834 5786 -1800
rect 5816 -1834 6366 -1800
rect 6396 -1834 6466 -1800
rect -541 -2104 -14 -2070
rect 16 -2104 566 -2070
rect 596 -2104 1146 -2070
rect 1176 -2104 1726 -2070
rect 1756 -2104 2306 -2070
rect 2336 -2104 2886 -2070
rect 2916 -2104 3466 -2070
rect 3496 -2104 4046 -2070
rect 4076 -2104 4626 -2070
rect 4656 -2104 5206 -2070
rect 5236 -2104 5786 -2070
rect 5816 -2104 6366 -2070
rect 6396 -2104 6466 -2070
rect -541 -2374 -14 -2340
rect 16 -2374 566 -2340
rect 596 -2374 1146 -2340
rect 1176 -2374 1726 -2340
rect 1756 -2374 2306 -2340
rect 2336 -2374 2886 -2340
rect 2916 -2374 3466 -2340
rect 3496 -2374 4046 -2340
rect 4076 -2374 4626 -2340
rect 4656 -2374 5206 -2340
rect 5236 -2374 5786 -2340
rect 5816 -2374 6366 -2340
rect 6396 -2374 6466 -2340
<< labels >>
rlabel poly -541 1814 6439 1844 1 WWL_0
port 1 n
rlabel metal1 -233 1800 -201 1814 1 VDD
port 3 n
rlabel metal1 -233 1574 -201 1588 1 GND
port 9 n
rlabel metal1 -541 1676 -532 1710 3 RWL1_0
port 22 e
rlabel metal2 -529 1676 -520 1710 1 RWL0_0
port 23 n
rlabel metal1 -493 1881 -478 1892 1 RBL1_0
port 24 n
rlabel metal1 -391 1886 -376 1892 1 WBLb_0
port 25 n
rlabel metal1 -57 1887 -42 1893 1 WBL_0
port 26 n
rlabel metal1 44 1882 59 1892 1 RBL0_0
port 27 n
<< end >>
