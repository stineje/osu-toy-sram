VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 10T_toy_magic
  CLASS BLOCK ;
  FOREIGN 10T_toy_magic ;
  ORIGIN 0.500 0.095 ;
  SIZE 2.760 BY 1.350 ;
  PIN WBL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.024175 ;
    PORT
      LAYER li1 ;
        RECT 1.820 0.825 1.895 0.970 ;
    END
  END WBL
  PIN WBLb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.023100 ;
    PORT
      LAYER li1 ;
        RECT -0.130 0.825 -0.055 0.965 ;
    END
  END WBLb
  PIN RBL0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.045150 ;
    PORT
      LAYER li1 ;
        RECT 2.185 0.095 2.260 0.305 ;
    END
  END RBL0
  PIN RBL1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.045150 ;
    PORT
      LAYER li1 ;
        RECT -0.500 0.095 -0.425 0.305 ;
    END
  END RBL1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.490 0.625 1.255 1.105 ;
      LAYER li1 ;
        RECT 0.800 1.035 0.960 1.105 ;
        RECT 0.810 1.025 0.950 1.035 ;
      LAYER met1 ;
        RECT -0.500 1.035 2.260 1.105 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.500 0.395 0.350 1.255 ;
        RECT 1.410 0.395 2.260 1.255 ;
        RECT -0.500 -0.095 2.260 0.395 ;
      LAYER li1 ;
        RECT 0.810 -0.025 0.950 -0.015 ;
        RECT 0.800 -0.095 0.960 -0.025 ;
      LAYER met1 ;
        RECT -0.500 -0.095 2.260 -0.025 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 0.275 0.825 0.350 0.965 ;
        RECT 0.490 0.775 0.565 0.915 ;
        RECT 1.195 0.835 1.255 0.915 ;
        POLYGON 1.195 0.835 1.255 0.835 1.255 0.775 ;
        RECT 1.410 0.825 1.485 0.965 ;
        RECT -0.285 0.415 -0.135 0.585 ;
        RECT 0.220 0.305 0.370 0.475 ;
        RECT 0.610 0.440 0.760 0.610 ;
        RECT 1.000 0.440 1.150 0.610 ;
        RECT 1.390 0.305 1.540 0.475 ;
        RECT 1.895 0.415 2.045 0.585 ;
        RECT 0.485 0.220 0.535 0.255 ;
        POLYGON 0.535 0.255 0.570 0.220 0.535 0.220 ;
        RECT 0.485 0.095 0.570 0.220 ;
        RECT 1.190 0.095 1.275 0.255 ;
  END
END 10T_toy_magic
MACRO 10T_4x4_magic
  CLASS BLOCK ;
  FOREIGN 10T_4x4_magic ;
  ORIGIN 0.440 1.570 ;
  SIZE 6.205 BY 2.940 ;
  PIN RWL1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 0.185 -0.820 0.335 -0.650 ;
        RECT 3.085 -0.820 3.235 -0.650 ;
      LAYER met1 ;
        POLYGON 2.315 -0.350 2.315 -0.520 2.145 -0.520 ;
        RECT 2.315 -0.520 2.565 -0.350 ;
        POLYGON 2.565 -0.350 2.735 -0.520 2.565 -0.520 ;
        POLYGON 5.215 -0.350 5.215 -0.520 5.045 -0.520 ;
        RECT 5.215 -0.520 5.465 -0.350 ;
        POLYGON 5.465 -0.350 5.635 -0.520 5.465 -0.520 ;
        POLYGON 2.145 -0.520 2.145 -0.650 2.015 -0.650 ;
        RECT 2.145 -0.650 2.235 -0.520 ;
        POLYGON 2.235 -0.520 2.365 -0.520 2.235 -0.650 ;
        POLYGON 2.515 -0.520 2.645 -0.520 2.645 -0.650 ;
        RECT 2.645 -0.650 2.735 -0.520 ;
        POLYGON 2.735 -0.520 2.865 -0.650 2.735 -0.650 ;
        POLYGON 5.045 -0.520 5.045 -0.650 4.915 -0.650 ;
        RECT 5.045 -0.650 5.135 -0.520 ;
        POLYGON 5.135 -0.520 5.265 -0.520 5.135 -0.650 ;
        POLYGON 5.415 -0.520 5.545 -0.520 5.545 -0.650 ;
        RECT 5.545 -0.650 5.635 -0.520 ;
        POLYGON 5.635 -0.520 5.765 -0.650 5.635 -0.650 ;
        RECT -0.420 -0.820 2.065 -0.650 ;
        POLYGON 2.065 -0.650 2.235 -0.650 2.065 -0.820 ;
        POLYGON 2.645 -0.650 2.815 -0.650 2.815 -0.820 ;
        RECT 2.815 -0.820 4.965 -0.650 ;
        POLYGON 4.965 -0.650 5.135 -0.650 4.965 -0.820 ;
        POLYGON 5.545 -0.650 5.715 -0.650 5.715 -0.820 ;
        RECT 5.715 -0.820 5.765 -0.650 ;
    END
  END RWL1_0
  PIN RWL0_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 2.365 -0.820 2.515 -0.650 ;
        RECT 5.265 -0.820 5.415 -0.650 ;
      LAYER mcon ;
        RECT 2.365 -0.815 2.515 -0.650 ;
      LAYER met1 ;
        RECT 2.365 -0.820 2.515 -0.650 ;
        RECT 5.265 -0.820 5.415 -0.650 ;
      LAYER met2 ;
        RECT -0.420 -0.820 5.765 -0.650 ;
    END
  END RWL0_0
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.030 0.510 0.820 1.370 ;
        RECT 1.880 0.510 3.720 1.370 ;
        RECT 4.780 0.510 5.630 1.370 ;
        RECT -0.030 0.020 5.630 0.510 ;
        RECT -0.030 -0.840 0.820 0.020 ;
        RECT 1.880 -0.840 3.720 0.020 ;
        RECT 4.780 -0.840 5.630 0.020 ;
        RECT -0.030 -1.330 5.630 -0.840 ;
      LAYER li1 ;
        RECT 1.270 0.020 1.430 0.100 ;
        RECT 4.170 0.020 4.330 0.100 ;
        RECT 1.270 -1.330 1.430 -1.250 ;
        RECT 4.170 -1.330 4.330 -1.250 ;
      LAYER met1 ;
        RECT -0.270 0.020 5.630 0.090 ;
        RECT -0.270 -1.330 5.630 -1.260 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.960 0.740 1.725 1.220 ;
        RECT 3.860 0.740 4.625 1.220 ;
      LAYER li1 ;
        RECT 1.270 1.140 1.430 1.220 ;
        RECT 4.170 1.140 4.330 1.220 ;
      LAYER mcon ;
        RECT 1.270 1.150 1.430 1.220 ;
        RECT 4.170 1.150 4.330 1.220 ;
      LAYER met1 ;
        RECT -0.270 1.150 5.630 1.220 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.960 -0.610 1.725 -0.130 ;
        RECT 3.860 -0.610 4.625 -0.130 ;
      LAYER li1 ;
        RECT 1.270 -0.210 1.430 -0.130 ;
        RECT 4.170 -0.210 4.330 -0.130 ;
      LAYER mcon ;
        RECT 1.270 -0.200 1.430 -0.130 ;
        RECT 4.170 -0.200 4.330 -0.130 ;
      LAYER met1 ;
        RECT -0.270 -0.200 5.630 -0.130 ;
    END
  END VDD
  PIN WWL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.084000 ;
    PORT
      LAYER li1 ;
        RECT -0.420 -0.130 -0.270 0.020 ;
    END
  END WWL_0
  PIN RWL0_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 2.365 0.530 2.515 0.700 ;
        RECT 5.265 0.530 5.415 0.700 ;
      LAYER mcon ;
        RECT 2.365 0.535 2.515 0.700 ;
      LAYER met1 ;
        RECT 2.365 0.530 2.515 0.700 ;
        RECT 5.265 0.530 5.415 0.700 ;
      LAYER met2 ;
        RECT -0.440 0.530 5.765 0.700 ;
    END
  END RWL0_1
  PIN RWL1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 0.185 0.530 0.335 0.700 ;
        RECT 3.085 0.530 3.235 0.700 ;
      LAYER met1 ;
        POLYGON 2.315 1.000 2.315 0.830 2.145 0.830 ;
        RECT 2.315 0.830 2.565 1.000 ;
        POLYGON 2.565 1.000 2.735 0.830 2.565 0.830 ;
        POLYGON 5.215 1.000 5.215 0.830 5.045 0.830 ;
        RECT 5.215 0.830 5.465 1.000 ;
        POLYGON 5.465 1.000 5.635 0.830 5.465 0.830 ;
        POLYGON 2.145 0.830 2.145 0.700 2.015 0.700 ;
        RECT 2.145 0.700 2.235 0.830 ;
        POLYGON 2.235 0.830 2.365 0.830 2.235 0.700 ;
        POLYGON 2.515 0.830 2.645 0.830 2.645 0.700 ;
        RECT 2.645 0.700 2.735 0.830 ;
        POLYGON 2.735 0.830 2.865 0.700 2.735 0.700 ;
        POLYGON 5.045 0.830 5.045 0.700 4.915 0.700 ;
        RECT 5.045 0.700 5.135 0.830 ;
        POLYGON 5.135 0.830 5.265 0.830 5.135 0.700 ;
        POLYGON 5.415 0.830 5.545 0.830 5.545 0.700 ;
        RECT 5.545 0.700 5.635 0.830 ;
        POLYGON 5.635 0.830 5.765 0.700 5.635 0.700 ;
        RECT -0.440 0.530 2.065 0.700 ;
        POLYGON 2.065 0.700 2.235 0.700 2.065 0.530 ;
        POLYGON 2.645 0.700 2.815 0.700 2.815 0.530 ;
        RECT 2.815 0.530 4.965 0.700 ;
        POLYGON 4.965 0.700 5.135 0.700 4.965 0.530 ;
        POLYGON 5.545 0.700 5.715 0.700 5.715 0.530 ;
        RECT 5.715 0.530 5.765 0.700 ;
    END
  END RWL1_1
  PIN WWL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.084000 ;
    PORT
      LAYER li1 ;
        RECT -0.420 1.220 -0.270 1.370 ;
    END
  END WWL_1
  PIN RBL1_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.090300 ;
    PORT
      LAYER li1 ;
        RECT -0.030 0.210 0.045 0.420 ;
        RECT -0.030 -1.140 0.045 -0.930 ;
    END
  END RBL1_0
  PIN WBLb_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.046200 ;
    PORT
      LAYER li1 ;
        RECT 0.340 0.940 0.415 1.080 ;
        RECT 0.340 -0.410 0.415 -0.270 ;
    END
  END WBLb_0
  PIN WBL_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048350 ;
    PORT
      LAYER li1 ;
        RECT 2.290 0.940 2.365 1.085 ;
        RECT 2.290 -0.410 2.365 -0.265 ;
    END
  END WBL_0
  PIN RBL0_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.090300 ;
    PORT
      LAYER li1 ;
        RECT 2.655 0.210 2.730 0.420 ;
        RECT 2.655 -1.140 2.730 -0.930 ;
    END
  END RBL0_0
  PIN RBL1_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.090300 ;
    PORT
      LAYER li1 ;
        RECT 2.870 0.210 2.945 0.420 ;
        RECT 2.870 -1.140 2.945 -0.930 ;
    END
  END RBL1_1
  PIN WBLb_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.046200 ;
    PORT
      LAYER li1 ;
        RECT 3.240 0.940 3.315 1.080 ;
        RECT 3.240 -0.410 3.315 -0.270 ;
    END
  END WBLb_1
  PIN WBL_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048350 ;
    PORT
      LAYER li1 ;
        RECT 5.190 0.940 5.265 1.085 ;
        RECT 5.190 -0.410 5.265 -0.265 ;
    END
  END WBL_1
  PIN RBL0_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.090300 ;
    PORT
      LAYER li1 ;
        RECT 5.555 0.210 5.630 0.420 ;
        RECT 5.555 -1.140 5.630 -0.930 ;
    END
  END RBL0_1
  OBS
      LAYER li1 ;
        RECT 0.745 0.940 0.820 1.080 ;
        RECT 0.960 0.890 1.035 1.030 ;
        RECT 1.665 0.950 1.725 1.030 ;
        POLYGON 1.665 0.950 1.725 0.950 1.725 0.890 ;
        RECT 1.880 0.940 1.955 1.080 ;
        RECT 3.645 0.940 3.720 1.080 ;
        RECT 3.860 0.890 3.935 1.030 ;
        RECT 4.565 0.950 4.625 1.030 ;
        POLYGON 4.565 0.950 4.625 0.950 4.625 0.890 ;
        RECT 4.780 0.940 4.855 1.080 ;
        RECT 0.690 0.420 0.840 0.590 ;
        RECT 1.080 0.555 1.230 0.725 ;
        RECT 1.470 0.555 1.620 0.725 ;
        RECT 1.860 0.420 2.010 0.590 ;
        RECT 3.590 0.420 3.740 0.590 ;
        RECT 3.980 0.555 4.130 0.725 ;
        RECT 4.370 0.555 4.520 0.725 ;
        RECT 4.760 0.420 4.910 0.590 ;
        RECT 0.955 0.335 1.005 0.370 ;
        POLYGON 1.005 0.370 1.040 0.335 1.005 0.335 ;
        RECT 0.955 0.210 1.040 0.335 ;
        RECT 1.660 0.210 1.745 0.370 ;
        RECT 3.855 0.335 3.905 0.370 ;
        POLYGON 3.905 0.370 3.940 0.335 3.905 0.335 ;
        RECT 3.855 0.210 3.940 0.335 ;
        RECT 4.560 0.210 4.645 0.370 ;
        RECT 0.745 -0.410 0.820 -0.270 ;
        RECT 0.960 -0.460 1.035 -0.320 ;
        RECT 1.665 -0.400 1.725 -0.320 ;
        POLYGON 1.665 -0.400 1.725 -0.400 1.725 -0.460 ;
        RECT 1.880 -0.410 1.955 -0.270 ;
        RECT 3.645 -0.410 3.720 -0.270 ;
        RECT 3.860 -0.460 3.935 -0.320 ;
        RECT 4.565 -0.400 4.625 -0.320 ;
        POLYGON 4.565 -0.400 4.625 -0.400 4.625 -0.460 ;
        RECT 4.780 -0.410 4.855 -0.270 ;
        RECT 0.690 -0.930 0.840 -0.760 ;
        RECT 1.080 -0.795 1.230 -0.625 ;
        RECT 1.470 -0.795 1.620 -0.625 ;
        RECT 1.860 -0.930 2.010 -0.760 ;
        RECT 3.590 -0.930 3.740 -0.760 ;
        RECT 3.980 -0.795 4.130 -0.625 ;
        RECT 4.370 -0.795 4.520 -0.625 ;
        RECT 4.760 -0.930 4.910 -0.760 ;
        RECT 0.955 -1.015 1.005 -0.980 ;
        POLYGON 1.005 -0.980 1.040 -1.015 1.005 -1.015 ;
        RECT 0.955 -1.140 1.040 -1.015 ;
        RECT 1.660 -1.140 1.745 -0.980 ;
        RECT 3.855 -1.015 3.905 -0.980 ;
        POLYGON 3.905 -0.980 3.940 -1.015 3.905 -1.015 ;
        RECT 3.855 -1.140 3.940 -1.015 ;
        RECT 4.560 -1.140 4.645 -0.980 ;
  END
END 10T_4x4_magic
END LIBRARY

