** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_4x4.sch
**.subckt 10T_4x4
x1 WWL_0 WBL_0 RBL0_0 RBL1_0 WBLb_0 RWL_0 RWL_0 VDD GND 10T_toy_xschem
x2 WWL_1 WBL_0 RBL0_0 RBL1_0 WBLb_0 RWL_1 RWL_1 VDD GND 10T_toy_xschem
x3 WWL_1 WBL_1 RBL0_1 RBL1_1 WBLb_1 RWL_1 RWL_1 VDD GND 10T_toy_xschem
x4 WWL_0 WBL_1 RBL0_1 RBL1_1 WBLb_1 RWL_0 RWL_0 VDD GND 10T_toy_xschem
V1 VDD GND 3
VWWL WBL_1 GND pwl 0ns 0V 5n 0.0v 5.1n 1.8v 10n 1.8v 10.1n 0v
VWBL WBLb_1 GND pwl 0ns 0V
VWBLb WWL_1 GND pwl 0ns 0V
VRWL0 RWL_1 GND pwl 0ns 0v
VWWL1 WBL_0 GND pwl 0ns 0V 5n 0.0v 5.1n 1.8v 10n 1.8v 10.1n 0v
VWBL1 WBLb_0 GND pwl 0ns 0V
VWBLb1 WWL_0 GND pwl 0ns 0V 4.9n 0.0v 5n 1.8v 9.9n 1.8v 10n 0v
VRWL2 RWL_0 GND pwl 0ns 0V 10.5n 0v 10.6n 1.8v
**** begin user architecture code

.lib /import/angmar1/repos/openpdk/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  10T_toy_xschem.sym # of pins=7
** sym_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_toy_xschem.sym
** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_toy_xschem.sch
.subckt 10T_toy_xschem  WWL WBL RBL0 RBL1 WBLb RWL0 RWL1  VDD  GND
*.ipin WWL
*.ipin RWL0
*.ipin RWL1
*.ipin WBL
*.ipin WBLb
*.opin RBL0
*.opin RBL1
x1 net1 net2 VDD GND INVX1
x2 net2 net1 VDD GND INVX1
XM1 net2 WWL WBL GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 WBLb WWL net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 RBL0 RWL0 net3 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.21 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 RBL1 RWL1 net4 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.21 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  INVX1.sym # of pins=2
** sym_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/INVX1.sym
** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/INVX1.sch
.subckt INVX1  Y A  VDD  GND
*.ipin A
*.opin Y
XM1 Y A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.21 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

**** begin user architecture code


.tran 1ps 30ns
.save all



**** end user architecture code
.end
