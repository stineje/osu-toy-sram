magic
tech sky130A
magscale 1 2
timestamp 1679443242
<< nwell >>
rect 834 228 866 230
rect 834 -42 866 -40
<< pwell >>
rect 254 18 286 20
rect -6 4 164 18
rect 237 -266 303 -252
rect 546 -266 574 274
rect 834 18 866 20
rect 834 -252 866 -250
<< psubdiffcont >>
rect 254 18 286 20
rect 834 18 866 20
rect 254 -252 286 -250
rect 834 -252 866 -250
<< nsubdiffcont >>
rect 254 228 286 230
rect 834 228 866 230
rect 254 -42 286 -40
rect 834 -42 866 -40
<< poly >>
rect -54 244 -6 274
rect 546 244 574 274
rect -54 -26 -6 4
rect 546 -26 574 4
<< polycont >>
rect -84 244 -54 274
rect -84 -26 -54 4
<< locali >>
rect 473 106 503 107
rect 473 -164 503 -163
<< corelocali >>
rect -6 -314 9 -266
rect 95 -314 110 -266
rect 430 -314 445 -266
rect 531 -314 546 -266
rect 574 -314 589 -266
rect 675 -314 690 -266
rect 1010 -314 1025 -266
rect 1111 -314 1126 -266
<< viali >>
rect 37 106 67 140
rect 473 107 503 140
rect 617 106 647 140
rect 1053 106 1083 140
rect 37 -164 67 -130
rect 473 -163 503 -130
rect 617 -164 647 -130
rect 1053 -164 1083 -130
<< metal1 >>
rect -54 230 -6 244
rect 546 230 574 244
tri 429 166 463 200 se
rect 463 166 513 200
tri 513 166 547 200 sw
tri 1009 166 1043 200 se
rect 1043 166 1093 200
tri 1093 166 1127 200 sw
tri 403 140 429 166 se
rect 429 140 447 166
tri 447 140 473 166 nw
tri 503 140 529 166 ne
rect 529 140 547 166
tri 547 140 573 166 sw
tri 983 140 1009 166 se
rect 1009 140 1027 166
tri 1027 140 1053 166 nw
tri 1083 140 1109 166 ne
rect 1109 140 1127 166
tri 1127 140 1153 166 sw
rect -88 106 37 140
rect 67 106 413 140
tri 413 106 447 140 nw
tri 529 106 563 140 ne
rect 563 106 617 140
rect 647 106 993 140
tri 993 106 1027 140 nw
tri 1109 106 1143 140 ne
rect 1143 106 1153 140
rect -54 4 -6 18
rect 546 4 574 18
rect -54 -40 -6 -26
rect 546 -40 574 -26
tri 429 -104 463 -70 se
rect 463 -104 513 -70
tri 513 -104 547 -70 sw
tri 1009 -104 1043 -70 se
rect 1043 -104 1093 -70
tri 1093 -104 1127 -70 sw
tri 403 -130 429 -104 se
rect 429 -130 447 -104
tri 447 -130 473 -104 nw
tri 503 -130 529 -104 ne
rect 529 -130 547 -104
tri 547 -130 573 -104 sw
tri 983 -130 1009 -104 se
rect 1009 -130 1027 -104
tri 1027 -130 1053 -104 nw
tri 1083 -130 1109 -104 ne
rect 1109 -130 1127 -104
tri 1127 -130 1153 -104 sw
rect -84 -164 37 -130
rect 67 -164 413 -130
tri 413 -164 447 -130 nw
tri 529 -164 563 -130 ne
rect 563 -164 617 -130
rect 647 -164 993 -130
tri 993 -164 1027 -130 nw
tri 1109 -164 1143 -130 ne
rect 1143 -164 1153 -130
rect -54 -266 -6 -252
rect 546 -266 574 -252
<< via1 >>
rect 473 107 503 140
rect 473 106 503 107
rect 1053 106 1083 140
rect 473 -163 503 -130
rect 473 -164 503 -163
rect 1053 -164 1083 -130
<< metal2 >>
rect -88 106 473 140
rect 503 106 1053 140
rect 1083 106 1153 140
rect -84 -164 473 -130
rect 503 -164 1053 -130
rect 1083 -164 1153 -130
use 10T_toy_magic  10T_toy_magic_0
timestamp 1679443213
transform 1 0 94 0 1 23
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_1
timestamp 1679443213
transform 1 0 674 0 1 23
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_2
timestamp 1679443213
transform 1 0 94 0 1 -247
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_3
timestamp 1679443213
transform 1 0 674 0 1 -247
box -100 -19 452 251
<< labels >>
rlabel metal1 -54 230 -24 244 1 VDD
port 4 ew power bidirectional abutment
rlabel metal1 -54 -40 -24 -26 1 VDD
port 4 ew power bidirectional abutment
rlabel metal1 -54 4 -24 18 1 GND
port 3 ew ground bidirectional abutment
rlabel metal1 -54 -266 -24 -252 1 GND
port 3 ew ground bidirectional abutment
rlabel corelocali -6 -314 9 -284 1 RBL1_0
port 9 ns signal output
rlabel corelocali 531 -314 546 -284 1 RBL0_0
port 12 ns signal output
rlabel corelocali 574 -314 589 -284 1 RBL1_1
port 13 ns signal output
rlabel corelocali 1111 -314 1126 -284 1 RBL0_1
port 16 ns signal output
rlabel locali -84 -26 -54 4 1 WWL_0
port 5 ew signal input
rlabel metal2 -54 -164 -24 -130 1 RWL0_0
port 2 ew signal input
rlabel metal1 -84 -164 -54 -130 1 RWL1_0
port 1 ew signal input
rlabel metal1 -88 106 -54 140 1 RWL1_1
port 7 ew signal input
rlabel metal2 -54 106 -20 140 1 RWL0_1
port 6 ew signal input
rlabel locali -84 244 -54 274 1 WWL_1
port 8 ew signal input
rlabel corelocali 95 -314 110 -284 1 WBLb_0
port 10 ns signal output
rlabel corelocali 430 -314 445 -284 1 WBL_0
port 11 ns signal output
rlabel corelocali 675 -314 690 -284 1 WBLb_1
port 14 ns signal output
rlabel corelocali 1010 -314 1025 -284 1 WBL_1
port 15 ns signal output
<< end >>
