*
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/models.all"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/tt_discrete.cor"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/ttcell.cor"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/npd.pm3"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/npass.pm3"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/ppu.pm3"


*** Define power and ground
vvdd vdd 0 DC 1.8V
vgnd gnd 0 DC 0V

VWWL wwl 0 pwl (0 0 5n 0.0 5.5n 1.8 10n 1.8 10.5n 0 15n 0.0 15.5n 1.8 20n 1.8 20.5n 0)
VWBL wbl 0 pwl (0 0 5n 0.0 5.5n 1.8 10n 1.8 10.5n 0 20.5n 0)
VWBLB wblb 0 pwl (0 1.8 5n 1.8 5.5n 0.0 10n 0.0 10.5n 1.8 20.5n 1.8)

VRWL0 rwl0 0 pwl (0 0 5n 0.0 5.5n 0.0 10n 0.0 10.5n 0 15n 0.0 15.5n 1.8 20n 1.8 20.5n 0)
VRWL1 rwl1 0 pwl (0 0 5n 0.0 5.5n 0.0 10n 0.0 10.5n 0 20.5n 0.0)

* Test pulse
VWWL42 a 0 pwl (0 0 5n 0.0 5.5n 1.8 10n 1.8 10.5n 0 15n 0.0 15.5n 1.8 20n 1.8 20.5n 0)

M1000 out1 a vdd vdd pshort w=1.26 l=0.15
M1001 out1 a gnd gnd nshort w=0.52 l=0.15


.tran 1ns 45ns

.print tran V(vwl,0)  V(wwl,0)  V(rwl0,0) V(rwl1,0) V(rbl0,0) V(rbl1,0)
.probe V(wwl,0) V(wbl,0) V(wblb,0) V(rwl0,0) V(rwl1,0) V(rbl0,0) V(rbl1,0) V(out1, 0) V(a, 0)
.op
.options probe post measout captab
.end

