magic
tech sky130A
magscale 1 2
timestamp 1656019537
<< error_s >>
rect 15 254 28 270
rect 117 268 130 270
rect 83 254 98 268
rect 107 254 137 268
rect 198 266 351 312
rect 180 254 372 266
rect 415 254 445 268
rect 451 254 464 270
rect 552 254 565 270
rect 595 254 608 270
rect 697 268 710 270
rect 663 254 678 268
rect 687 254 717 268
rect 778 266 931 312
rect 760 254 952 266
rect 995 254 1025 268
rect 1031 254 1044 270
rect 1132 254 1145 270
rect 1175 254 1188 270
rect 1277 268 1290 270
rect 1243 254 1258 268
rect 1267 254 1297 268
rect 1358 266 1511 312
rect 1340 254 1532 266
rect 1575 254 1605 268
rect 1611 254 1624 270
rect 1712 254 1725 270
rect 1755 254 1768 270
rect 1857 268 1870 270
rect 1823 254 1838 268
rect 1847 254 1877 268
rect 1938 266 2091 312
rect 1920 254 2112 266
rect 2155 254 2185 268
rect 2191 254 2204 270
rect 2292 254 2305 270
rect 2335 254 2348 270
rect 2437 268 2450 270
rect 2403 254 2418 268
rect 2427 254 2457 268
rect 2518 266 2671 312
rect 2500 254 2692 266
rect 2735 254 2765 268
rect 2771 254 2784 270
rect 2872 254 2885 270
rect 2915 254 2928 270
rect 3017 268 3030 270
rect 2983 254 2998 268
rect 3007 254 3037 268
rect 3098 266 3251 312
rect 3080 254 3272 266
rect 3315 254 3345 268
rect 3351 254 3364 270
rect 3452 254 3465 270
rect 3495 254 3508 270
rect 3597 268 3610 270
rect 3563 254 3578 268
rect 3587 254 3617 268
rect 3678 266 3831 312
rect 3660 254 3852 266
rect 3895 254 3925 268
rect 3931 254 3944 270
rect 4032 254 4045 270
rect 4075 254 4088 270
rect 4177 268 4190 270
rect 4143 254 4158 268
rect 4167 254 4197 268
rect 4258 266 4411 312
rect 4240 254 4432 266
rect 4475 254 4505 268
rect 4511 254 4524 270
rect 4612 254 4625 270
rect 0 240 4625 254
rect 15 136 28 240
rect 73 218 74 228
rect 89 218 102 228
rect 73 214 102 218
rect 107 214 137 240
rect 155 226 171 228
rect 243 226 296 240
rect 244 224 308 226
rect 155 214 170 218
rect 73 212 170 214
rect 57 204 108 212
rect 57 192 82 204
rect 89 192 108 204
rect 139 204 189 212
rect 139 196 155 204
rect 162 202 189 204
rect 198 204 213 208
rect 260 204 292 224
rect 351 212 366 240
rect 415 237 445 240
rect 415 234 451 237
rect 381 226 397 228
rect 382 214 397 218
rect 415 215 454 234
rect 473 228 480 229
rect 479 221 480 228
rect 463 218 464 221
rect 479 218 492 221
rect 415 214 445 215
rect 454 214 460 215
rect 463 214 492 218
rect 382 213 492 214
rect 382 212 498 213
rect 351 204 419 212
rect 198 202 267 204
rect 285 202 419 204
rect 162 198 234 202
rect 162 196 287 198
rect 162 192 234 196
rect 57 184 108 192
rect 155 188 234 192
rect 315 188 419 202
rect 448 204 498 212
rect 448 195 464 204
rect 155 184 419 188
rect 445 192 464 195
rect 471 192 498 204
rect 445 184 498 192
rect 73 176 74 184
rect 89 176 102 184
rect 73 168 89 176
rect 70 161 89 164
rect 70 152 92 161
rect 43 142 92 152
rect 43 136 73 142
rect 92 137 97 142
rect 15 120 89 136
rect 107 128 137 184
rect 172 174 380 184
rect 415 180 460 184
rect 463 183 464 184
rect 479 183 492 184
rect 339 170 387 174
rect 222 148 252 157
rect 315 150 330 157
rect 351 148 387 170
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 15 118 28 120
rect 43 118 77 120
rect 15 102 89 118
rect 116 114 129 128
rect 144 114 160 130
rect 206 125 217 138
rect -1 80 0 96
rect 15 80 28 102
rect 43 80 73 102
rect 116 98 178 114
rect 206 107 217 123
rect 222 118 232 138
rect 242 118 256 138
rect 259 125 268 138
rect 284 125 293 138
rect 222 107 256 118
rect 259 107 268 123
rect 284 107 293 123
rect 300 118 310 138
rect 320 118 334 138
rect 335 125 346 138
rect 300 107 334 118
rect 335 107 346 123
rect 392 114 408 130
rect 415 128 445 180
rect 479 176 480 183
rect 464 168 480 176
rect 451 136 464 155
rect 479 136 509 152
rect 451 120 525 136
rect 451 118 464 120
rect 479 118 513 120
rect 116 96 129 98
rect 144 96 178 98
rect 116 80 178 96
rect 222 91 238 94
rect 300 91 330 102
rect 378 98 424 114
rect 451 102 525 118
rect 378 96 412 98
rect 377 80 424 96
rect 451 80 464 102
rect 479 80 509 102
rect 536 80 537 96
rect 552 80 565 240
rect 595 136 608 240
rect 653 218 654 228
rect 669 218 682 228
rect 653 214 682 218
rect 687 214 717 240
rect 735 226 751 228
rect 823 226 876 240
rect 824 224 888 226
rect 735 214 750 218
rect 653 212 750 214
rect 637 204 688 212
rect 637 192 662 204
rect 669 192 688 204
rect 719 204 769 212
rect 719 196 735 204
rect 742 202 769 204
rect 778 204 793 208
rect 840 204 872 224
rect 931 212 946 240
rect 995 237 1025 240
rect 995 234 1031 237
rect 961 226 977 228
rect 962 214 977 218
rect 995 215 1034 234
rect 1053 228 1060 229
rect 1059 221 1060 228
rect 1043 218 1044 221
rect 1059 218 1072 221
rect 995 214 1025 215
rect 1034 214 1040 215
rect 1043 214 1072 218
rect 962 213 1072 214
rect 962 212 1078 213
rect 931 204 999 212
rect 778 202 847 204
rect 865 202 999 204
rect 742 198 814 202
rect 742 196 867 198
rect 742 192 814 196
rect 637 184 688 192
rect 735 188 814 192
rect 895 188 999 202
rect 1028 204 1078 212
rect 1028 195 1044 204
rect 735 184 999 188
rect 1025 192 1044 195
rect 1051 192 1078 204
rect 1025 184 1078 192
rect 653 176 654 184
rect 669 176 682 184
rect 653 168 669 176
rect 650 161 669 164
rect 650 152 672 161
rect 623 142 672 152
rect 623 136 653 142
rect 672 137 677 142
rect 595 120 669 136
rect 687 128 717 184
rect 752 174 960 184
rect 995 180 1040 184
rect 1043 183 1044 184
rect 1059 183 1072 184
rect 919 170 967 174
rect 802 148 832 157
rect 895 150 910 157
rect 931 148 967 170
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 595 118 608 120
rect 623 118 657 120
rect 595 102 669 118
rect 696 114 709 128
rect 724 114 740 130
rect 786 125 797 138
rect 579 80 580 96
rect 595 80 608 102
rect 623 80 653 102
rect 696 98 758 114
rect 786 107 797 123
rect 802 118 812 138
rect 822 118 836 138
rect 839 125 848 138
rect 864 125 873 138
rect 802 107 836 118
rect 839 107 848 123
rect 864 107 873 123
rect 880 118 890 138
rect 900 118 914 138
rect 915 125 926 138
rect 880 107 914 118
rect 915 107 926 123
rect 972 114 988 130
rect 995 128 1025 180
rect 1059 176 1060 183
rect 1044 168 1060 176
rect 1031 136 1044 155
rect 1059 136 1089 152
rect 1031 120 1105 136
rect 1031 118 1044 120
rect 1059 118 1093 120
rect 696 96 709 98
rect 724 96 758 98
rect 696 80 758 96
rect 802 91 818 94
rect 880 91 910 102
rect 958 98 1004 114
rect 1031 102 1105 118
rect 958 96 992 98
rect 957 80 1004 96
rect 1031 80 1044 102
rect 1059 80 1089 102
rect 1116 80 1117 96
rect 1132 80 1145 240
rect 1175 136 1188 240
rect 1233 218 1234 228
rect 1249 218 1262 228
rect 1233 214 1262 218
rect 1267 214 1297 240
rect 1315 226 1331 228
rect 1403 226 1456 240
rect 1404 224 1468 226
rect 1315 214 1330 218
rect 1233 212 1330 214
rect 1217 204 1268 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1299 204 1349 212
rect 1299 196 1315 204
rect 1322 202 1349 204
rect 1358 204 1373 208
rect 1420 204 1452 224
rect 1511 212 1526 240
rect 1575 237 1605 240
rect 1575 234 1611 237
rect 1541 226 1557 228
rect 1542 214 1557 218
rect 1575 215 1614 234
rect 1633 228 1640 229
rect 1639 221 1640 228
rect 1623 218 1624 221
rect 1639 218 1652 221
rect 1575 214 1605 215
rect 1614 214 1620 215
rect 1623 214 1652 218
rect 1542 213 1652 214
rect 1542 212 1658 213
rect 1511 204 1579 212
rect 1358 202 1427 204
rect 1445 202 1579 204
rect 1322 198 1394 202
rect 1322 196 1447 198
rect 1322 192 1394 196
rect 1217 184 1268 192
rect 1315 188 1394 192
rect 1475 188 1579 202
rect 1608 204 1658 212
rect 1608 195 1624 204
rect 1315 184 1579 188
rect 1605 192 1624 195
rect 1631 192 1658 204
rect 1605 184 1658 192
rect 1233 176 1234 184
rect 1249 176 1262 184
rect 1233 168 1249 176
rect 1230 161 1249 164
rect 1230 152 1252 161
rect 1203 142 1252 152
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1175 120 1249 136
rect 1267 128 1297 184
rect 1332 174 1540 184
rect 1575 180 1620 184
rect 1623 183 1624 184
rect 1639 183 1652 184
rect 1499 170 1547 174
rect 1382 148 1412 157
rect 1475 150 1490 157
rect 1511 148 1547 170
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1175 118 1188 120
rect 1203 118 1237 120
rect 1175 102 1249 118
rect 1276 114 1289 128
rect 1304 114 1320 130
rect 1366 125 1377 138
rect 1159 80 1160 96
rect 1175 80 1188 102
rect 1203 80 1233 102
rect 1276 98 1338 114
rect 1366 107 1377 123
rect 1382 118 1392 138
rect 1402 118 1416 138
rect 1419 125 1428 138
rect 1444 125 1453 138
rect 1382 107 1416 118
rect 1419 107 1428 123
rect 1444 107 1453 123
rect 1460 118 1470 138
rect 1480 118 1494 138
rect 1495 125 1506 138
rect 1460 107 1494 118
rect 1495 107 1506 123
rect 1552 114 1568 130
rect 1575 128 1605 180
rect 1639 176 1640 183
rect 1624 168 1640 176
rect 1611 136 1624 155
rect 1639 136 1669 152
rect 1611 120 1685 136
rect 1611 118 1624 120
rect 1639 118 1673 120
rect 1276 96 1289 98
rect 1304 96 1338 98
rect 1276 80 1338 96
rect 1382 91 1398 94
rect 1460 91 1490 102
rect 1538 98 1584 114
rect 1611 102 1685 118
rect 1538 96 1572 98
rect 1537 80 1584 96
rect 1611 80 1624 102
rect 1639 80 1669 102
rect 1696 80 1697 96
rect 1712 80 1725 240
rect 1755 136 1768 240
rect 1813 218 1814 228
rect 1829 218 1842 228
rect 1813 214 1842 218
rect 1847 214 1877 240
rect 1895 226 1911 228
rect 1983 226 2036 240
rect 1984 224 2048 226
rect 1895 214 1910 218
rect 1813 212 1910 214
rect 1797 204 1848 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1879 204 1929 212
rect 1879 196 1895 204
rect 1902 202 1929 204
rect 1938 204 1953 208
rect 2000 204 2032 224
rect 2091 212 2106 240
rect 2155 237 2185 240
rect 2155 234 2191 237
rect 2121 226 2137 228
rect 2122 214 2137 218
rect 2155 215 2194 234
rect 2213 228 2220 229
rect 2219 221 2220 228
rect 2203 218 2204 221
rect 2219 218 2232 221
rect 2155 214 2185 215
rect 2194 214 2200 215
rect 2203 214 2232 218
rect 2122 213 2232 214
rect 2122 212 2238 213
rect 2091 204 2159 212
rect 1938 202 2007 204
rect 2025 202 2159 204
rect 1902 198 1974 202
rect 1902 196 2027 198
rect 1902 192 1974 196
rect 1797 184 1848 192
rect 1895 188 1974 192
rect 2055 188 2159 202
rect 2188 204 2238 212
rect 2188 195 2204 204
rect 1895 184 2159 188
rect 2185 192 2204 195
rect 2211 192 2238 204
rect 2185 184 2238 192
rect 1813 176 1814 184
rect 1829 176 1842 184
rect 1813 168 1829 176
rect 1810 161 1829 164
rect 1810 152 1832 161
rect 1783 142 1832 152
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1755 120 1829 136
rect 1847 128 1877 184
rect 1912 174 2120 184
rect 2155 180 2200 184
rect 2203 183 2204 184
rect 2219 183 2232 184
rect 2079 170 2127 174
rect 1962 148 1992 157
rect 2055 150 2070 157
rect 2091 148 2127 170
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 1755 118 1768 120
rect 1783 118 1817 120
rect 1755 102 1829 118
rect 1856 114 1869 128
rect 1884 114 1900 130
rect 1946 125 1957 138
rect 1739 80 1740 96
rect 1755 80 1768 102
rect 1783 80 1813 102
rect 1856 98 1918 114
rect 1946 107 1957 123
rect 1962 118 1972 138
rect 1982 118 1996 138
rect 1999 125 2008 138
rect 2024 125 2033 138
rect 1962 107 1996 118
rect 1999 107 2008 123
rect 2024 107 2033 123
rect 2040 118 2050 138
rect 2060 118 2074 138
rect 2075 125 2086 138
rect 2040 107 2074 118
rect 2075 107 2086 123
rect 2132 114 2148 130
rect 2155 128 2185 180
rect 2219 176 2220 183
rect 2204 168 2220 176
rect 2191 136 2204 155
rect 2219 136 2249 152
rect 2191 120 2265 136
rect 2191 118 2204 120
rect 2219 118 2253 120
rect 1856 96 1869 98
rect 1884 96 1918 98
rect 1856 80 1918 96
rect 1962 91 1978 94
rect 2040 91 2070 102
rect 2118 98 2164 114
rect 2191 102 2265 118
rect 2118 96 2152 98
rect 2117 80 2164 96
rect 2191 80 2204 102
rect 2219 80 2249 102
rect 2276 80 2277 96
rect 2292 80 2305 240
rect 2335 136 2348 240
rect 2393 218 2394 228
rect 2409 218 2422 228
rect 2393 214 2422 218
rect 2427 214 2457 240
rect 2475 226 2491 228
rect 2563 226 2616 240
rect 2564 224 2628 226
rect 2475 214 2490 218
rect 2393 212 2490 214
rect 2377 204 2428 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2459 204 2509 212
rect 2459 196 2475 204
rect 2482 202 2509 204
rect 2518 204 2533 208
rect 2580 204 2612 224
rect 2671 212 2686 240
rect 2735 237 2765 240
rect 2735 234 2771 237
rect 2701 226 2717 228
rect 2702 214 2717 218
rect 2735 215 2774 234
rect 2793 228 2800 229
rect 2799 221 2800 228
rect 2783 218 2784 221
rect 2799 218 2812 221
rect 2735 214 2765 215
rect 2774 214 2780 215
rect 2783 214 2812 218
rect 2702 213 2812 214
rect 2702 212 2818 213
rect 2671 204 2739 212
rect 2518 202 2587 204
rect 2605 202 2739 204
rect 2482 198 2554 202
rect 2482 196 2607 198
rect 2482 192 2554 196
rect 2377 184 2428 192
rect 2475 188 2554 192
rect 2635 188 2739 202
rect 2768 204 2818 212
rect 2768 195 2784 204
rect 2475 184 2739 188
rect 2765 192 2784 195
rect 2791 192 2818 204
rect 2765 184 2818 192
rect 2393 176 2394 184
rect 2409 176 2422 184
rect 2393 168 2409 176
rect 2390 161 2409 164
rect 2390 152 2412 161
rect 2363 142 2412 152
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2335 120 2409 136
rect 2427 128 2457 184
rect 2492 174 2700 184
rect 2735 180 2780 184
rect 2783 183 2784 184
rect 2799 183 2812 184
rect 2659 170 2707 174
rect 2542 148 2572 157
rect 2635 150 2650 157
rect 2671 148 2707 170
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2335 118 2348 120
rect 2363 118 2397 120
rect 2335 102 2409 118
rect 2436 114 2449 128
rect 2464 114 2480 130
rect 2526 125 2537 138
rect 2319 80 2320 96
rect 2335 80 2348 102
rect 2363 80 2393 102
rect 2436 98 2498 114
rect 2526 107 2537 123
rect 2542 118 2552 138
rect 2562 118 2576 138
rect 2579 125 2588 138
rect 2604 125 2613 138
rect 2542 107 2576 118
rect 2579 107 2588 123
rect 2604 107 2613 123
rect 2620 118 2630 138
rect 2640 118 2654 138
rect 2655 125 2666 138
rect 2620 107 2654 118
rect 2655 107 2666 123
rect 2712 114 2728 130
rect 2735 128 2765 180
rect 2799 176 2800 183
rect 2784 168 2800 176
rect 2771 136 2784 155
rect 2799 136 2829 152
rect 2771 120 2845 136
rect 2771 118 2784 120
rect 2799 118 2833 120
rect 2436 96 2449 98
rect 2464 96 2498 98
rect 2436 80 2498 96
rect 2542 91 2558 94
rect 2620 91 2650 102
rect 2698 98 2744 114
rect 2771 102 2845 118
rect 2698 96 2732 98
rect 2697 80 2744 96
rect 2771 80 2784 102
rect 2799 80 2829 102
rect 2856 80 2857 96
rect 2872 80 2885 240
rect 2915 136 2928 240
rect 2973 218 2974 228
rect 2989 218 3002 228
rect 2973 214 3002 218
rect 3007 214 3037 240
rect 3055 226 3071 228
rect 3143 226 3196 240
rect 3144 224 3208 226
rect 3055 214 3070 218
rect 2973 212 3070 214
rect 2957 204 3008 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3039 204 3089 212
rect 3039 196 3055 204
rect 3062 202 3089 204
rect 3098 204 3113 208
rect 3160 204 3192 224
rect 3251 212 3266 240
rect 3315 237 3345 240
rect 3315 234 3351 237
rect 3281 226 3297 228
rect 3282 214 3297 218
rect 3315 215 3354 234
rect 3373 228 3380 229
rect 3379 221 3380 228
rect 3363 218 3364 221
rect 3379 218 3392 221
rect 3315 214 3345 215
rect 3354 214 3360 215
rect 3363 214 3392 218
rect 3282 213 3392 214
rect 3282 212 3398 213
rect 3251 204 3319 212
rect 3098 202 3167 204
rect 3185 202 3319 204
rect 3062 198 3134 202
rect 3062 196 3187 198
rect 3062 192 3134 196
rect 2957 184 3008 192
rect 3055 188 3134 192
rect 3215 188 3319 202
rect 3348 204 3398 212
rect 3348 195 3364 204
rect 3055 184 3319 188
rect 3345 192 3364 195
rect 3371 192 3398 204
rect 3345 184 3398 192
rect 2973 176 2974 184
rect 2989 176 3002 184
rect 2973 168 2989 176
rect 2970 161 2989 164
rect 2970 152 2992 161
rect 2943 142 2992 152
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2915 120 2989 136
rect 3007 128 3037 184
rect 3072 174 3280 184
rect 3315 180 3360 184
rect 3363 183 3364 184
rect 3379 183 3392 184
rect 3239 170 3287 174
rect 3122 148 3152 157
rect 3215 150 3230 157
rect 3251 148 3287 170
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 2915 118 2928 120
rect 2943 118 2977 120
rect 2915 102 2989 118
rect 3016 114 3029 128
rect 3044 114 3060 130
rect 3106 125 3117 138
rect 2899 80 2900 96
rect 2915 80 2928 102
rect 2943 80 2973 102
rect 3016 98 3078 114
rect 3106 107 3117 123
rect 3122 118 3132 138
rect 3142 118 3156 138
rect 3159 125 3168 138
rect 3184 125 3193 138
rect 3122 107 3156 118
rect 3159 107 3168 123
rect 3184 107 3193 123
rect 3200 118 3210 138
rect 3220 118 3234 138
rect 3235 125 3246 138
rect 3200 107 3234 118
rect 3235 107 3246 123
rect 3292 114 3308 130
rect 3315 128 3345 180
rect 3379 176 3380 183
rect 3364 168 3380 176
rect 3351 136 3364 155
rect 3379 136 3409 152
rect 3351 120 3425 136
rect 3351 118 3364 120
rect 3379 118 3413 120
rect 3016 96 3029 98
rect 3044 96 3078 98
rect 3016 80 3078 96
rect 3122 91 3138 94
rect 3200 91 3230 102
rect 3278 98 3324 114
rect 3351 102 3425 118
rect 3278 96 3312 98
rect 3277 80 3324 96
rect 3351 80 3364 102
rect 3379 80 3409 102
rect 3436 80 3437 96
rect 3452 80 3465 240
rect 3495 136 3508 240
rect 3553 218 3554 228
rect 3569 218 3582 228
rect 3553 214 3582 218
rect 3587 214 3617 240
rect 3635 226 3651 228
rect 3723 226 3776 240
rect 3724 224 3788 226
rect 3635 214 3650 218
rect 3553 212 3650 214
rect 3537 204 3588 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3619 204 3669 212
rect 3619 196 3635 204
rect 3642 202 3669 204
rect 3678 204 3693 208
rect 3740 204 3772 224
rect 3831 212 3846 240
rect 3895 237 3925 240
rect 3895 234 3931 237
rect 3861 226 3877 228
rect 3862 214 3877 218
rect 3895 215 3934 234
rect 3953 228 3960 229
rect 3959 221 3960 228
rect 3943 218 3944 221
rect 3959 218 3972 221
rect 3895 214 3925 215
rect 3934 214 3940 215
rect 3943 214 3972 218
rect 3862 213 3972 214
rect 3862 212 3978 213
rect 3831 204 3899 212
rect 3678 202 3747 204
rect 3765 202 3899 204
rect 3642 198 3714 202
rect 3642 196 3767 198
rect 3642 192 3714 196
rect 3537 184 3588 192
rect 3635 188 3714 192
rect 3795 188 3899 202
rect 3928 204 3978 212
rect 3928 195 3944 204
rect 3635 184 3899 188
rect 3925 192 3944 195
rect 3951 192 3978 204
rect 3925 184 3978 192
rect 3553 176 3554 184
rect 3569 176 3582 184
rect 3553 168 3569 176
rect 3550 161 3569 164
rect 3550 152 3572 161
rect 3523 142 3572 152
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3495 120 3569 136
rect 3587 128 3617 184
rect 3652 174 3860 184
rect 3895 180 3940 184
rect 3943 183 3944 184
rect 3959 183 3972 184
rect 3819 170 3867 174
rect 3702 148 3732 157
rect 3795 150 3810 157
rect 3831 148 3867 170
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3495 118 3508 120
rect 3523 118 3557 120
rect 3495 102 3569 118
rect 3596 114 3609 128
rect 3624 114 3640 130
rect 3686 125 3697 138
rect 3479 80 3480 96
rect 3495 80 3508 102
rect 3523 80 3553 102
rect 3596 98 3658 114
rect 3686 107 3697 123
rect 3702 118 3712 138
rect 3722 118 3736 138
rect 3739 125 3748 138
rect 3764 125 3773 138
rect 3702 107 3736 118
rect 3739 107 3748 123
rect 3764 107 3773 123
rect 3780 118 3790 138
rect 3800 118 3814 138
rect 3815 125 3826 138
rect 3780 107 3814 118
rect 3815 107 3826 123
rect 3872 114 3888 130
rect 3895 128 3925 180
rect 3959 176 3960 183
rect 3944 168 3960 176
rect 3931 136 3944 155
rect 3959 136 3989 152
rect 3931 120 4005 136
rect 3931 118 3944 120
rect 3959 118 3993 120
rect 3596 96 3609 98
rect 3624 96 3658 98
rect 3596 80 3658 96
rect 3702 91 3718 94
rect 3780 91 3810 102
rect 3858 98 3904 114
rect 3931 102 4005 118
rect 3858 96 3892 98
rect 3857 80 3904 96
rect 3931 80 3944 102
rect 3959 80 3989 102
rect 4016 80 4017 96
rect 4032 80 4045 240
rect 4075 136 4088 240
rect 4133 218 4134 228
rect 4149 218 4162 228
rect 4133 214 4162 218
rect 4167 214 4197 240
rect 4215 226 4231 228
rect 4303 226 4356 240
rect 4304 224 4368 226
rect 4215 214 4230 218
rect 4133 212 4230 214
rect 4117 204 4168 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4199 204 4249 212
rect 4199 196 4215 204
rect 4222 202 4249 204
rect 4258 204 4273 208
rect 4320 204 4352 224
rect 4411 212 4426 240
rect 4475 237 4505 240
rect 4475 234 4511 237
rect 4441 226 4457 228
rect 4442 214 4457 218
rect 4475 215 4514 234
rect 4533 228 4540 229
rect 4539 221 4540 228
rect 4523 218 4524 221
rect 4539 218 4552 221
rect 4475 214 4505 215
rect 4514 214 4520 215
rect 4523 214 4552 218
rect 4442 213 4552 214
rect 4442 212 4558 213
rect 4411 204 4479 212
rect 4258 202 4327 204
rect 4345 202 4479 204
rect 4222 198 4294 202
rect 4222 196 4347 198
rect 4222 192 4294 196
rect 4117 184 4168 192
rect 4215 188 4294 192
rect 4375 188 4479 202
rect 4508 204 4558 212
rect 4508 195 4524 204
rect 4215 184 4479 188
rect 4505 192 4524 195
rect 4531 192 4558 204
rect 4505 184 4558 192
rect 4133 176 4134 184
rect 4149 176 4162 184
rect 4133 168 4149 176
rect 4130 161 4149 164
rect 4130 152 4152 161
rect 4103 142 4152 152
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4075 120 4149 136
rect 4167 128 4197 184
rect 4232 174 4440 184
rect 4475 180 4520 184
rect 4523 183 4524 184
rect 4539 183 4552 184
rect 4399 170 4447 174
rect 4282 148 4312 157
rect 4375 150 4390 157
rect 4411 148 4447 170
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4075 118 4088 120
rect 4103 118 4137 120
rect 4075 102 4149 118
rect 4176 114 4189 128
rect 4204 114 4220 130
rect 4266 125 4277 138
rect 4059 80 4060 96
rect 4075 80 4088 102
rect 4103 80 4133 102
rect 4176 98 4238 114
rect 4266 107 4277 123
rect 4282 118 4292 138
rect 4302 118 4316 138
rect 4319 125 4328 138
rect 4344 125 4353 138
rect 4282 107 4316 118
rect 4319 107 4328 123
rect 4344 107 4353 123
rect 4360 118 4370 138
rect 4380 118 4394 138
rect 4395 125 4406 138
rect 4360 107 4394 118
rect 4395 107 4406 123
rect 4452 114 4468 130
rect 4475 128 4505 180
rect 4539 176 4540 183
rect 4524 168 4540 176
rect 4511 136 4524 155
rect 4539 136 4569 152
rect 4511 120 4585 136
rect 4511 118 4524 120
rect 4539 118 4573 120
rect 4176 96 4189 98
rect 4204 96 4238 98
rect 4176 80 4238 96
rect 4282 91 4298 94
rect 4360 91 4390 102
rect 4438 98 4484 114
rect 4511 102 4585 118
rect 4438 96 4472 98
rect 4437 80 4484 96
rect 4511 80 4524 102
rect 4539 80 4569 102
rect 4596 80 4597 96
rect 4612 80 4625 240
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 160 80
rect 172 68 247 80
rect 305 68 380 80
rect 392 68 423 80
rect 429 68 464 80
rect 98 66 260 68
rect -7 38 34 46
rect 116 38 129 66
rect 144 64 159 66
rect 183 39 190 46
rect 193 38 260 66
rect 292 66 464 68
rect 262 44 290 48
rect 292 44 372 66
rect 393 64 408 66
rect 262 42 372 44
rect 262 38 290 42
rect 292 38 372 42
rect -1 28 0 38
rect 15 28 28 38
rect 43 28 73 38
rect 116 28 159 38
rect 166 28 174 38
rect 193 30 196 38
rect 260 30 292 38
rect 193 28 359 30
rect 378 28 389 38
rect 393 28 423 38
rect 451 28 464 66
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 740 80
rect 752 68 827 80
rect 885 68 960 80
rect 972 68 1003 80
rect 1009 68 1044 80
rect 678 66 840 68
rect 573 38 614 46
rect 696 38 709 66
rect 724 64 739 66
rect 763 39 770 46
rect 773 38 840 66
rect 872 66 1044 68
rect 842 44 870 48
rect 872 44 952 66
rect 973 64 988 66
rect 842 42 952 44
rect 842 38 870 42
rect 872 38 952 42
rect 479 28 509 38
rect 536 28 537 38
rect 552 28 565 38
rect 579 28 580 38
rect 595 28 608 38
rect 623 28 653 38
rect 696 28 739 38
rect 746 28 754 38
rect 773 30 776 38
rect 840 30 872 38
rect 773 28 939 30
rect 958 28 969 38
rect 973 28 1003 38
rect 1031 28 1044 66
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1320 80
rect 1332 68 1407 80
rect 1465 68 1540 80
rect 1552 68 1583 80
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1153 38 1194 46
rect 1276 38 1289 66
rect 1304 64 1319 66
rect 1343 39 1350 46
rect 1353 38 1420 66
rect 1452 66 1624 68
rect 1422 44 1450 48
rect 1452 44 1532 66
rect 1553 64 1568 66
rect 1422 42 1532 44
rect 1422 38 1450 42
rect 1452 38 1532 42
rect 1059 28 1089 38
rect 1116 28 1117 38
rect 1132 28 1145 38
rect 1159 28 1160 38
rect 1175 28 1188 38
rect 1203 28 1233 38
rect 1276 28 1319 38
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1420 30 1452 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1553 28 1583 38
rect 1611 28 1624 66
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1900 80
rect 1912 68 1987 80
rect 2045 68 2120 80
rect 2132 68 2163 80
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1733 38 1774 46
rect 1856 38 1869 66
rect 1884 64 1899 66
rect 1923 39 1930 46
rect 1933 38 2000 66
rect 2032 66 2204 68
rect 2002 44 2030 48
rect 2032 44 2112 66
rect 2133 64 2148 66
rect 2002 42 2112 44
rect 2002 38 2030 42
rect 2032 38 2112 42
rect 1639 28 1669 38
rect 1696 28 1697 38
rect 1712 28 1725 38
rect 1739 28 1740 38
rect 1755 28 1768 38
rect 1783 28 1813 38
rect 1856 28 1899 38
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 2000 30 2032 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2133 28 2163 38
rect 2191 28 2204 66
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2480 80
rect 2492 68 2567 80
rect 2625 68 2700 80
rect 2712 68 2743 80
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2313 38 2354 46
rect 2436 38 2449 66
rect 2464 64 2479 66
rect 2503 39 2510 46
rect 2513 38 2580 66
rect 2612 66 2784 68
rect 2582 44 2610 48
rect 2612 44 2692 66
rect 2713 64 2728 66
rect 2582 42 2692 44
rect 2582 38 2610 42
rect 2612 38 2692 42
rect 2219 28 2249 38
rect 2276 28 2277 38
rect 2292 28 2305 38
rect 2319 28 2320 38
rect 2335 28 2348 38
rect 2363 28 2393 38
rect 2436 28 2479 38
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2580 30 2612 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2713 28 2743 38
rect 2771 28 2784 66
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3060 80
rect 3072 68 3147 80
rect 3205 68 3280 80
rect 3292 68 3323 80
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 2893 38 2934 46
rect 3016 38 3029 66
rect 3044 64 3059 66
rect 3083 39 3090 46
rect 3093 38 3160 66
rect 3192 66 3364 68
rect 3162 44 3190 48
rect 3192 44 3272 66
rect 3293 64 3308 66
rect 3162 42 3272 44
rect 3162 38 3190 42
rect 3192 38 3272 42
rect 2799 28 2829 38
rect 2856 28 2857 38
rect 2872 28 2885 38
rect 2899 28 2900 38
rect 2915 28 2928 38
rect 2943 28 2973 38
rect 3016 28 3059 38
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3160 30 3192 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3293 28 3323 38
rect 3351 28 3364 66
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3640 80
rect 3652 68 3727 80
rect 3785 68 3860 80
rect 3872 68 3903 80
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3473 38 3514 46
rect 3596 38 3609 66
rect 3624 64 3639 66
rect 3663 39 3670 46
rect 3673 38 3740 66
rect 3772 66 3944 68
rect 3742 44 3770 48
rect 3772 44 3852 66
rect 3873 64 3888 66
rect 3742 42 3852 44
rect 3742 38 3770 42
rect 3772 38 3852 42
rect 3379 28 3409 38
rect 3436 28 3437 38
rect 3452 28 3465 38
rect 3479 28 3480 38
rect 3495 28 3508 38
rect 3523 28 3553 38
rect 3596 28 3639 38
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3740 30 3772 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3873 28 3903 38
rect 3931 28 3944 66
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4220 80
rect 4232 68 4307 80
rect 4365 68 4440 80
rect 4452 68 4483 80
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4053 38 4094 46
rect 4176 38 4189 66
rect 4204 64 4219 66
rect 4243 39 4250 46
rect 4253 38 4320 66
rect 4352 66 4524 68
rect 4322 44 4350 48
rect 4352 44 4432 66
rect 4453 64 4468 66
rect 4322 42 4432 44
rect 4322 38 4350 42
rect 4352 38 4432 42
rect 3959 28 3989 38
rect 4016 28 4017 38
rect 4032 28 4045 38
rect 4059 28 4060 38
rect 4075 28 4088 38
rect 4103 28 4133 38
rect 4176 28 4219 38
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4320 30 4352 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4453 28 4483 38
rect 4511 28 4524 66
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4539 28 4569 38
rect 4596 28 4597 38
rect 4612 28 4625 38
rect -1 22 4625 28
rect 0 14 4625 22
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 129 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 243 0 294 1
rect 451 0 464 14
rect 244 -2 308 0
rect 479 -4 509 14
rect 552 0 565 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 709 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 823 0 874 1
rect 1031 0 1044 14
rect 824 -2 888 0
rect 1059 -4 1089 14
rect 1132 0 1145 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1289 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1403 0 1454 1
rect 1611 0 1624 14
rect 1404 -2 1468 0
rect 1639 -4 1669 14
rect 1712 0 1725 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1869 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1983 0 2034 1
rect 2191 0 2204 14
rect 1984 -2 2048 0
rect 2219 -4 2249 14
rect 2292 0 2305 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2449 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2563 0 2614 1
rect 2771 0 2784 14
rect 2564 -2 2628 0
rect 2799 -4 2829 14
rect 2872 0 2885 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3029 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3143 0 3194 1
rect 3351 0 3364 14
rect 3144 -2 3208 0
rect 3379 -4 3409 14
rect 3452 0 3465 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3609 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3723 0 3774 1
rect 3931 0 3944 14
rect 3724 -2 3788 0
rect 3959 -4 3989 14
rect 4032 0 4045 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4189 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4303 0 4354 1
rect 4511 0 4524 14
rect 4304 -2 4368 0
rect 4539 -4 4569 14
rect 4612 0 4625 14
<< pwell >>
rect 552 0 580 270
rect 1132 0 1160 270
rect 1712 0 1740 270
rect 2292 0 2320 270
rect 2872 0 2900 270
rect 3452 0 3480 270
rect 4032 0 4060 270
<< poly >>
rect 552 240 580 270
rect 1132 240 1160 270
rect 1712 240 1740 270
rect 2292 240 2320 270
rect 2872 240 2900 270
rect 3452 240 3480 270
rect 4032 240 4060 270
<< polycont >>
rect 623 102 653 136
rect 1059 102 1089 136
rect 1203 102 1233 136
rect 1639 102 1669 136
rect 1783 102 1813 136
rect 2219 102 2249 136
rect 2363 102 2393 136
rect 2799 102 2829 136
rect 2943 102 2973 136
rect 3379 102 3409 136
rect 3523 102 3553 136
rect 3959 102 3989 136
rect 4103 102 4133 136
rect 4539 102 4569 136
<< viali >>
rect 43 102 73 136
rect 479 102 509 136
rect 623 102 653 136
rect 1059 102 1089 136
rect 1203 102 1233 136
rect 1639 102 1669 136
rect 1783 102 1813 136
rect 2219 102 2249 136
rect 2363 102 2393 136
rect 2799 102 2829 136
rect 2943 102 2973 136
rect 3379 102 3409 136
rect 3523 102 3553 136
rect 3959 102 3989 136
rect 4103 102 4133 136
rect 4539 102 4569 136
<< metal1 >>
rect 552 226 580 240
rect 1132 226 1160 240
rect 1712 226 1740 240
rect 2292 226 2320 240
rect 2872 226 2900 240
rect 3452 226 3480 240
rect 4032 226 4060 240
rect 0 102 43 136
rect 73 102 479 136
rect 509 102 623 136
rect 653 102 1059 136
rect 1089 102 1203 136
rect 1233 102 1639 136
rect 1669 102 1783 136
rect 1813 102 2219 136
rect 2249 102 2363 136
rect 2393 102 2799 136
rect 2829 102 2943 136
rect 2973 102 3379 136
rect 3409 102 3523 136
rect 3553 102 3959 136
rect 3989 102 4103 136
rect 4133 102 4539 136
rect 552 0 580 14
rect 1132 0 1160 14
rect 1712 0 1740 14
rect 2292 0 2320 14
rect 2872 0 2900 14
rect 3452 0 3480 14
rect 4032 0 4060 14
use 10T_toy_magic  10T_toy_magic_7
timestamp 1655238822
transform 1 0 100 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_6
timestamp 1655238822
transform 1 0 680 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_5
timestamp 1655238822
transform 1 0 1260 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_4
timestamp 1655238822
transform 1 0 1840 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_3
timestamp 1655238822
transform 1 0 2420 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_2
timestamp 1655238822
transform 1 0 3000 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_1
timestamp 1655238822
transform 1 0 4160 0 1 19
box -107 -23 471 293
use 10T_toy_magic  10T_toy_magic_0
timestamp 1655238822
transform 1 0 3580 0 1 19
box -107 -23 471 293
<< labels >>
rlabel poly 0 240 30 270 1 WWL
port 17 ew signal input
rlabel metal1 0 102 15 136 1 RWL
port 18 ew signal input
rlabel corelocali 74 184 89 212 1 WBLb_0
port 19 ns signal input
rlabel corelocali 464 184 479 213 1 WBL_0
port 20 ns signal input
rlabel corelocali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel corelocali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel corelocali 654 184 669 212 1 WBLb_1
port 21 ns signal input
rlabel corelocali 1044 184 1059 213 1 WBL_1
port 22 ns signal input
rlabel corelocali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel corelocali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel corelocali 1234 184 1249 212 1 WBLb_2
port 23 ns signal input
rlabel corelocali 1624 184 1639 213 1 WBL_2
port 24 ns signal input
rlabel corelocali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel corelocali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel corelocali 1814 184 1829 212 1 WBLb_3
port 25 ns signal input
rlabel corelocali 2204 184 2219 213 1 WBL_3
port 26 ns signal input
rlabel corelocali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel corelocali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel corelocali 2394 184 2409 212 1 WBLb_4
port 27 ns signal input
rlabel corelocali 2784 184 2799 213 1 WBL_4
port 28 ns signal input
rlabel corelocali 2320 38 2335 80 1 RBL1_4
port 8 ns signal output
rlabel corelocali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel corelocali 2974 184 2989 212 1 WBLb_5
port 29 ns signal input
rlabel corelocali 3364 184 3379 213 1 WBL_5
port 30 ns signal input
rlabel corelocali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel corelocali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel corelocali 3554 184 3569 212 1 WBLb_6
port 31 ns signal input
rlabel corelocali 3944 184 3959 213 1 WBL_6
port 32 ns signal input
rlabel corelocali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel corelocali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel corelocali 4134 184 4149 212 1 WBLb_7
port 33 ns signal input
rlabel corelocali 4524 184 4539 213 1 WBL_7
port 34 ns signal input
rlabel corelocali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel corelocali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel metal1 0 226 15 240 1 VDD
port 35 ns power bidirectional abutment
rlabel metal1 0 0 15 14 1 GND
port 36 ns ground bidirectional abutment
<< end >>
