magic
tech sky130A
magscale 1 2
timestamp 1668471109
<< error_s >>
rect 9 258 22 274
rect 77 258 92 272
rect 111 260 124 322
rect 192 270 345 316
rect 174 258 366 270
rect 445 258 458 322
rect 540 258 559 274
rect 574 258 580 274
rect 589 258 602 274
rect 657 258 672 272
rect 691 260 704 322
rect 772 270 925 316
rect 754 258 946 270
rect 1025 258 1038 322
rect 1126 258 1139 274
rect -54 244 1139 258
rect 9 174 22 244
rect 67 228 84 232
rect 88 230 96 232
rect 86 228 96 230
rect 67 218 96 228
rect 149 218 165 232
rect 203 228 209 230
rect 216 228 324 244
rect 331 228 337 230
rect 345 228 360 244
rect 426 238 445 241
rect 67 216 165 218
rect 192 216 360 228
rect 375 218 391 232
rect 426 219 448 238
rect 458 232 474 233
rect 457 230 474 232
rect 458 225 474 230
rect 448 218 454 219
rect 457 218 486 225
rect 375 217 486 218
rect 375 216 492 217
rect 51 208 102 216
rect 149 208 183 216
rect 51 196 76 208
rect 83 196 102 208
rect 156 206 183 208
rect 192 206 413 216
rect 448 213 454 216
rect 156 202 413 206
rect 51 188 102 196
rect 149 188 413 202
rect 457 208 492 216
rect 3 140 22 174
rect 67 180 96 188
rect 67 174 84 180
rect 67 172 101 174
rect 149 172 165 188
rect 166 178 374 188
rect 375 178 391 188
rect 439 184 454 199
rect 457 196 458 208
rect 465 196 492 208
rect 457 188 492 196
rect 457 187 486 188
rect 177 174 391 178
rect 192 172 391 174
rect 426 174 439 184
rect 457 174 474 187
rect 426 172 474 174
rect 68 168 101 172
rect 64 166 101 168
rect 64 165 131 166
rect 64 160 95 165
rect 101 160 131 165
rect 64 156 131 160
rect 37 153 131 156
rect 37 146 86 153
rect 37 140 67 146
rect 86 141 91 146
rect 3 124 83 140
rect 95 132 131 153
rect 192 148 381 172
rect 426 171 473 172
rect 439 166 473 171
rect 207 145 381 148
rect 200 142 381 145
rect 409 165 473 166
rect 3 122 22 124
rect 37 122 71 124
rect 3 106 83 122
rect 3 100 22 106
rect -7 84 22 100
rect 37 90 67 106
rect 95 84 101 132
rect 104 126 123 132
rect 138 126 168 134
rect 104 118 168 126
rect 104 102 184 118
rect 200 111 262 142
rect 278 111 340 142
rect 409 140 458 165
rect 473 140 503 158
rect 372 126 402 134
rect 409 132 519 140
rect 372 118 417 126
rect 104 100 123 102
rect 138 100 184 102
rect 104 84 184 100
rect 211 98 246 111
rect 287 108 324 111
rect 287 106 329 108
rect 216 95 246 98
rect 225 91 232 95
rect 232 90 233 91
rect 191 84 201 90
rect -13 76 28 84
rect -13 50 2 76
rect 9 50 28 76
rect 92 72 123 84
rect 138 72 241 84
rect 253 74 279 100
rect 294 95 324 106
rect 356 102 418 118
rect 356 100 402 102
rect 356 84 418 100
rect 430 84 436 132
rect 439 124 519 132
rect 439 122 458 124
rect 473 122 507 124
rect 439 107 519 122
rect 439 106 525 107
rect 439 84 458 106
rect 473 90 503 106
rect 531 100 537 174
rect 540 100 559 244
rect 574 100 580 244
rect 589 174 602 244
rect 647 228 664 232
rect 668 230 676 232
rect 666 228 676 230
rect 647 218 676 228
rect 729 218 745 232
rect 783 228 789 230
rect 796 228 904 244
rect 911 228 917 230
rect 925 228 940 244
rect 1006 238 1025 241
rect 647 216 745 218
rect 772 216 940 228
rect 955 218 971 232
rect 1006 219 1028 238
rect 1038 232 1054 233
rect 1037 230 1054 232
rect 1038 225 1054 230
rect 1028 218 1034 219
rect 1037 218 1066 225
rect 955 217 1066 218
rect 955 216 1072 217
rect 631 208 682 216
rect 729 208 763 216
rect 631 196 656 208
rect 663 196 682 208
rect 736 206 763 208
rect 772 206 993 216
rect 1028 213 1034 216
rect 736 202 993 206
rect 631 188 682 196
rect 729 188 993 202
rect 1037 208 1072 216
rect 583 140 602 174
rect 647 180 676 188
rect 647 174 664 180
rect 647 172 681 174
rect 729 172 745 188
rect 746 178 954 188
rect 955 178 971 188
rect 1019 184 1034 199
rect 1037 196 1038 208
rect 1045 196 1072 208
rect 1037 188 1072 196
rect 1037 187 1066 188
rect 757 174 971 178
rect 772 172 971 174
rect 1006 174 1019 184
rect 1037 174 1054 187
rect 1006 172 1054 174
rect 648 168 681 172
rect 644 166 681 168
rect 644 165 711 166
rect 644 160 675 165
rect 681 160 711 165
rect 644 156 711 160
rect 617 153 711 156
rect 617 146 666 153
rect 617 140 647 146
rect 666 141 671 146
rect 583 124 663 140
rect 675 132 711 153
rect 772 148 961 172
rect 1006 171 1053 172
rect 1019 166 1053 171
rect 787 145 961 148
rect 780 142 961 145
rect 989 165 1053 166
rect 583 122 602 124
rect 617 122 651 124
rect 583 106 663 122
rect 583 100 602 106
rect 299 74 402 84
rect 253 72 402 74
rect 423 72 458 84
rect 92 70 254 72
rect 104 50 123 70
rect 138 68 168 70
rect -13 42 28 50
rect 110 46 123 50
rect 175 54 254 70
rect 286 70 458 72
rect 286 54 365 70
rect 372 68 402 70
rect -7 32 22 42
rect 37 32 67 46
rect 110 32 153 46
rect 175 42 365 54
rect 430 50 436 70
rect 160 32 190 42
rect 191 32 349 42
rect 353 32 383 42
rect 387 32 417 46
rect 445 32 458 70
rect 530 84 559 100
rect 573 84 602 100
rect 617 90 647 106
rect 675 84 681 132
rect 684 126 703 132
rect 718 126 748 134
rect 684 118 748 126
rect 684 102 764 118
rect 780 111 842 142
rect 858 111 920 142
rect 989 140 1038 165
rect 1053 140 1083 156
rect 952 126 982 134
rect 989 132 1099 140
rect 952 118 997 126
rect 684 100 703 102
rect 718 100 764 102
rect 684 84 764 100
rect 791 98 826 111
rect 867 108 904 111
rect 867 106 909 108
rect 796 95 826 98
rect 805 91 812 95
rect 812 90 813 91
rect 771 84 781 90
rect 530 76 565 84
rect 530 50 531 76
rect 538 50 565 76
rect 473 32 503 46
rect 530 42 565 50
rect 567 76 608 84
rect 567 50 582 76
rect 589 50 608 76
rect 672 72 703 84
rect 718 72 821 84
rect 833 74 859 100
rect 874 95 904 106
rect 936 102 998 118
rect 936 100 982 102
rect 936 84 998 100
rect 1010 84 1016 132
rect 1019 124 1099 132
rect 1019 122 1038 124
rect 1053 122 1087 124
rect 1019 106 1099 122
rect 1019 84 1038 106
rect 1053 90 1083 106
rect 1111 100 1117 174
rect 1126 100 1139 244
rect 879 74 982 84
rect 833 72 982 74
rect 1003 72 1038 84
rect 672 70 834 72
rect 684 50 703 70
rect 718 68 748 70
rect 567 42 608 50
rect 690 46 703 50
rect 755 54 834 70
rect 866 70 1038 72
rect 866 54 945 70
rect 952 68 982 70
rect 530 32 559 42
rect 573 32 602 42
rect 617 32 647 46
rect 690 32 733 46
rect 755 42 945 54
rect 1010 50 1016 70
rect 740 32 770 42
rect 771 32 929 42
rect 933 32 963 42
rect 967 32 997 46
rect 1025 32 1038 70
rect 1110 84 1139 100
rect 1110 76 1145 84
rect 1110 50 1111 76
rect 1118 50 1145 76
rect 1053 32 1083 46
rect 1110 42 1145 50
rect 1110 32 1139 42
rect -54 18 1139 32
rect 9 -12 22 18
rect 37 4 67 18
rect 110 4 153 18
rect 160 4 380 18
rect 387 4 417 18
rect 77 -10 92 2
rect 111 -10 124 4
rect 192 0 345 4
rect 74 -12 96 -10
rect 174 -12 366 0
rect 445 -12 458 18
rect 473 4 503 18
rect 540 -12 559 18
rect 574 -12 580 18
rect 589 -12 602 18
rect 617 4 647 18
rect 690 4 733 18
rect 740 4 960 18
rect 967 4 997 18
rect 657 -10 672 2
rect 691 -10 704 4
rect 772 0 925 4
rect 654 -12 676 -10
rect 754 -12 946 0
rect 1025 -12 1038 18
rect 1053 4 1083 18
rect 1126 -12 1139 18
rect -54 -26 1139 -12
rect 9 -96 22 -26
rect 74 -30 96 -26
rect 67 -42 84 -38
rect 88 -40 96 -38
rect 86 -42 96 -40
rect 67 -52 96 -42
rect 149 -52 165 -38
rect 203 -48 209 -40
rect 216 -42 324 -26
rect 67 -54 165 -52
rect 51 -62 102 -54
rect 149 -62 183 -54
rect 51 -74 76 -62
rect 83 -74 102 -62
rect 156 -64 183 -62
rect 192 -62 209 -48
rect 254 -62 286 -42
rect 331 -48 337 -40
rect 345 -48 360 -26
rect 426 -32 445 -29
rect 331 -54 360 -48
rect 375 -52 391 -38
rect 426 -51 448 -32
rect 458 -38 474 -37
rect 457 -40 474 -38
rect 458 -45 474 -40
rect 448 -52 454 -51
rect 457 -52 486 -45
rect 375 -53 486 -52
rect 375 -54 492 -53
rect 331 -62 413 -54
rect 448 -57 454 -54
rect 192 -64 413 -62
rect 156 -68 228 -64
rect 256 -66 284 -64
rect 309 -68 413 -64
rect 51 -82 102 -74
rect 149 -76 281 -68
rect 286 -76 413 -68
rect 457 -62 492 -54
rect 149 -78 228 -76
rect 309 -78 413 -76
rect 149 -82 246 -78
rect 3 -130 22 -96
rect 67 -90 96 -82
rect 67 -96 84 -90
rect 67 -98 101 -96
rect 149 -98 165 -82
rect 166 -86 246 -82
rect 294 -82 413 -78
rect 294 -86 374 -82
rect 166 -92 374 -86
rect 375 -92 391 -82
rect 439 -86 454 -71
rect 457 -74 458 -62
rect 465 -74 492 -62
rect 457 -82 492 -74
rect 457 -83 486 -82
rect 177 -96 281 -92
rect 68 -102 101 -98
rect 64 -104 101 -102
rect 64 -105 131 -104
rect 64 -110 95 -105
rect 101 -110 131 -105
rect 192 -108 207 -96
rect 64 -114 131 -110
rect 37 -117 131 -114
rect 37 -124 86 -117
rect 37 -130 67 -124
rect 86 -129 91 -124
rect 3 -146 83 -130
rect 95 -138 131 -117
rect 216 -118 246 -109
rect 269 -114 287 -96
rect 345 -98 391 -92
rect 426 -96 439 -86
rect 457 -96 474 -83
rect 426 -98 474 -96
rect 307 -104 309 -102
rect 309 -109 321 -104
rect 294 -116 324 -109
rect 294 -118 325 -116
rect 345 -118 381 -98
rect 426 -99 473 -98
rect 439 -104 473 -99
rect 192 -122 381 -118
rect 207 -125 381 -122
rect 200 -128 381 -125
rect 409 -105 473 -104
rect 3 -148 22 -146
rect 37 -148 71 -146
rect 3 -164 83 -148
rect 3 -170 22 -164
rect -7 -186 22 -170
rect 37 -180 67 -164
rect 95 -186 101 -138
rect 104 -144 123 -138
rect 138 -144 168 -136
rect 104 -152 168 -144
rect 104 -168 184 -152
rect 200 -159 262 -128
rect 278 -159 340 -128
rect 409 -130 458 -105
rect 473 -130 503 -112
rect 372 -144 402 -136
rect 409 -138 519 -130
rect 372 -152 417 -144
rect 104 -170 123 -168
rect 138 -170 184 -168
rect 104 -186 184 -170
rect 211 -172 246 -159
rect 287 -162 324 -159
rect 287 -164 329 -162
rect 216 -175 246 -172
rect 225 -179 232 -175
rect 232 -180 233 -179
rect 191 -186 201 -180
rect -13 -194 28 -186
rect -13 -220 2 -194
rect 9 -220 28 -194
rect 92 -198 123 -186
rect 138 -198 241 -186
rect 253 -196 279 -170
rect 294 -175 324 -164
rect 356 -168 418 -152
rect 356 -170 402 -168
rect 356 -186 418 -170
rect 430 -186 436 -138
rect 439 -146 519 -138
rect 439 -148 458 -146
rect 473 -148 507 -146
rect 439 -163 519 -148
rect 439 -164 525 -163
rect 439 -186 458 -164
rect 473 -180 503 -164
rect 531 -170 537 -96
rect 540 -170 559 -26
rect 574 -170 580 -26
rect 589 -96 602 -26
rect 654 -30 676 -26
rect 647 -42 664 -38
rect 668 -40 676 -38
rect 666 -42 676 -40
rect 647 -52 676 -42
rect 729 -52 745 -38
rect 783 -48 789 -40
rect 796 -42 904 -26
rect 647 -54 745 -52
rect 631 -62 682 -54
rect 729 -62 763 -54
rect 631 -74 656 -62
rect 663 -74 682 -62
rect 736 -64 763 -62
rect 772 -62 789 -48
rect 834 -62 866 -42
rect 911 -48 917 -40
rect 925 -48 940 -26
rect 1006 -32 1025 -29
rect 911 -54 940 -48
rect 955 -52 971 -38
rect 1006 -51 1028 -32
rect 1038 -38 1054 -37
rect 1037 -40 1054 -38
rect 1038 -45 1054 -40
rect 1028 -52 1034 -51
rect 1037 -52 1066 -45
rect 955 -53 1066 -52
rect 955 -54 1072 -53
rect 911 -62 993 -54
rect 1028 -57 1034 -54
rect 772 -64 993 -62
rect 736 -68 808 -64
rect 836 -66 864 -64
rect 889 -68 993 -64
rect 631 -82 682 -74
rect 729 -76 861 -68
rect 866 -76 993 -68
rect 1037 -62 1072 -54
rect 729 -78 808 -76
rect 889 -78 993 -76
rect 729 -82 826 -78
rect 583 -130 602 -96
rect 647 -90 676 -82
rect 647 -96 664 -90
rect 647 -98 681 -96
rect 729 -98 745 -82
rect 746 -86 826 -82
rect 874 -82 993 -78
rect 874 -86 954 -82
rect 746 -92 954 -86
rect 955 -92 971 -82
rect 1019 -86 1034 -71
rect 1037 -74 1038 -62
rect 1045 -74 1072 -62
rect 1037 -82 1072 -74
rect 1037 -83 1066 -82
rect 757 -96 861 -92
rect 648 -102 681 -98
rect 644 -104 681 -102
rect 644 -105 711 -104
rect 644 -110 675 -105
rect 681 -110 711 -105
rect 772 -108 787 -96
rect 644 -114 711 -110
rect 617 -117 711 -114
rect 617 -124 666 -117
rect 617 -130 647 -124
rect 666 -129 671 -124
rect 583 -146 663 -130
rect 675 -138 711 -117
rect 796 -118 826 -109
rect 849 -114 867 -96
rect 925 -98 971 -92
rect 1006 -96 1019 -86
rect 1037 -96 1054 -83
rect 1006 -98 1054 -96
rect 887 -104 889 -102
rect 889 -109 901 -104
rect 874 -116 904 -109
rect 874 -118 905 -116
rect 925 -118 961 -98
rect 1006 -99 1053 -98
rect 1019 -104 1053 -99
rect 772 -122 961 -118
rect 787 -125 961 -122
rect 780 -128 961 -125
rect 989 -105 1053 -104
rect 583 -148 602 -146
rect 617 -148 651 -146
rect 583 -164 663 -148
rect 583 -170 602 -164
rect 299 -196 402 -186
rect 253 -198 402 -196
rect 423 -198 458 -186
rect 92 -200 254 -198
rect 104 -220 123 -200
rect 138 -202 168 -200
rect -13 -228 28 -220
rect -7 -238 22 -228
rect 110 -238 123 -220
rect 175 -216 254 -200
rect 286 -200 458 -198
rect 286 -216 365 -200
rect 372 -202 402 -200
rect 175 -228 365 -216
rect 430 -220 436 -200
rect 160 -238 168 -228
rect 187 -236 190 -228
rect 191 -236 209 -228
rect 254 -236 286 -228
rect 331 -236 349 -228
rect 187 -238 353 -236
rect 372 -238 383 -228
rect 445 -238 458 -200
rect 530 -186 559 -170
rect 573 -186 602 -170
rect 617 -180 647 -164
rect 675 -186 681 -138
rect 684 -144 703 -138
rect 718 -144 748 -136
rect 684 -152 748 -144
rect 684 -168 764 -152
rect 780 -159 842 -128
rect 858 -159 920 -128
rect 989 -130 1038 -105
rect 1053 -130 1083 -114
rect 952 -144 982 -136
rect 989 -138 1099 -130
rect 952 -152 997 -144
rect 684 -170 703 -168
rect 718 -170 764 -168
rect 684 -186 764 -170
rect 791 -172 826 -159
rect 867 -162 904 -159
rect 867 -164 909 -162
rect 796 -175 826 -172
rect 805 -179 812 -175
rect 812 -180 813 -179
rect 771 -186 781 -180
rect 530 -194 565 -186
rect 530 -220 531 -194
rect 538 -220 565 -194
rect 530 -228 565 -220
rect 567 -194 608 -186
rect 567 -220 582 -194
rect 589 -220 608 -194
rect 672 -198 703 -186
rect 718 -198 821 -186
rect 833 -196 859 -170
rect 874 -175 904 -164
rect 936 -168 998 -152
rect 936 -170 982 -168
rect 936 -186 998 -170
rect 1010 -186 1016 -138
rect 1019 -146 1099 -138
rect 1019 -148 1038 -146
rect 1053 -148 1087 -146
rect 1019 -164 1099 -148
rect 1019 -186 1038 -164
rect 1053 -180 1083 -164
rect 1111 -170 1117 -96
rect 1126 -170 1139 -26
rect 879 -196 982 -186
rect 833 -198 982 -196
rect 1003 -198 1038 -186
rect 672 -200 834 -198
rect 684 -220 703 -200
rect 718 -202 748 -200
rect 567 -228 608 -220
rect 530 -238 559 -228
rect 573 -238 602 -228
rect 690 -238 703 -220
rect 755 -216 834 -200
rect 866 -200 1038 -198
rect 866 -216 945 -200
rect 952 -202 982 -200
rect 755 -228 945 -216
rect 1010 -220 1016 -200
rect 740 -238 748 -228
rect 767 -236 770 -228
rect 771 -236 789 -228
rect 834 -236 866 -228
rect 911 -236 929 -228
rect 767 -238 933 -236
rect 952 -238 963 -228
rect 1025 -238 1038 -200
rect 1110 -186 1139 -170
rect 1110 -194 1145 -186
rect 1110 -220 1111 -194
rect 1118 -220 1145 -194
rect 1110 -228 1145 -220
rect 1110 -238 1139 -228
rect -54 -252 1139 -238
rect 9 -314 22 -252
rect 37 -270 67 -252
rect 110 -266 153 -252
rect 160 -265 168 -252
rect 201 -265 339 -252
rect 372 -265 380 -252
rect 123 -284 153 -266
rect 216 -266 324 -265
rect 216 -270 246 -266
rect 254 -268 286 -266
rect 294 -270 324 -266
rect 387 -284 417 -252
rect 445 -266 458 -252
rect 473 -270 503 -252
rect 540 -314 559 -252
rect 574 -314 580 -252
rect 589 -314 602 -252
rect 617 -270 647 -252
rect 690 -266 733 -252
rect 740 -265 748 -252
rect 781 -265 919 -252
rect 952 -265 960 -252
rect 703 -284 733 -266
rect 796 -266 904 -265
rect 796 -270 826 -266
rect 834 -268 866 -266
rect 874 -270 904 -266
rect 967 -284 997 -252
rect 1025 -266 1038 -252
rect 1053 -270 1083 -252
rect 1126 -314 1139 -252
<< nwell >>
rect 834 228 866 230
rect 834 -42 866 -40
<< pwell >>
rect 254 18 286 20
rect -6 4 164 18
rect 237 -266 303 -252
rect 546 -266 574 274
rect 834 18 866 20
rect 834 -252 866 -250
<< psubdiffcont >>
rect 254 18 286 20
rect 834 18 866 20
rect 254 -252 286 -250
rect 834 -252 866 -250
<< nsubdiffcont >>
rect 254 228 286 230
rect 834 228 866 230
rect 254 -42 286 -40
rect 834 -42 866 -40
<< poly >>
rect -54 244 -6 274
rect 546 244 574 274
rect -54 -26 -6 4
rect 546 -26 574 4
<< locali >>
rect 473 106 503 107
rect 473 -164 503 -163
<< corelocali >>
rect 96 274 111 322
rect 430 274 445 322
rect 676 274 691 322
rect 1010 274 1025 322
rect -6 -314 9 -266
rect 531 -314 546 -266
rect 574 -314 589 -266
rect 1111 -314 1126 -266
<< viali >>
rect 37 106 67 140
rect 473 107 503 140
rect 617 106 647 140
rect 1053 106 1083 140
rect 37 -164 67 -130
rect 473 -163 503 -130
rect 617 -164 647 -130
rect 1053 -164 1083 -130
<< metal1 >>
rect -54 230 -6 244
rect 546 230 574 244
tri 429 166 463 200 se
rect 463 166 513 200
tri 513 166 547 200 sw
tri 1009 166 1043 200 se
rect 1043 166 1093 200
tri 1093 166 1127 200 sw
tri 403 140 429 166 se
rect 429 140 447 166
tri 447 140 473 166 nw
tri 503 140 529 166 ne
rect 529 140 547 166
tri 547 140 573 166 sw
tri 983 140 1009 166 se
rect 1009 140 1027 166
tri 1027 140 1053 166 nw
tri 1083 140 1109 166 ne
rect 1109 140 1127 166
tri 1127 140 1153 166 sw
rect -54 106 37 140
rect 67 106 413 140
tri 413 106 447 140 nw
tri 529 106 563 140 ne
rect 563 106 617 140
rect 647 106 993 140
tri 993 106 1027 140 nw
tri 1109 106 1143 140 ne
rect 1143 106 1153 140
rect -54 4 -6 18
rect 546 4 574 18
rect -54 -40 -6 -26
rect 546 -40 574 -26
tri 429 -104 463 -70 se
rect 463 -104 513 -70
tri 513 -104 547 -70 sw
tri 1009 -104 1043 -70 se
rect 1043 -104 1093 -70
tri 1093 -104 1127 -70 sw
tri 403 -130 429 -104 se
rect 429 -130 447 -104
tri 447 -130 473 -104 nw
tri 503 -130 529 -104 ne
rect 529 -130 547 -104
tri 547 -130 573 -104 sw
tri 983 -130 1009 -104 se
rect 1009 -130 1027 -104
tri 1027 -130 1053 -104 nw
tri 1083 -130 1109 -104 ne
rect 1109 -130 1127 -104
tri 1127 -130 1153 -104 sw
rect -54 -164 37 -130
rect 67 -164 413 -130
tri 413 -164 447 -130 nw
tri 529 -164 563 -130 ne
rect 563 -164 617 -130
rect 647 -164 993 -130
tri 993 -164 1027 -130 nw
tri 1109 -164 1143 -130 ne
rect 1143 -164 1153 -130
rect -54 -266 -6 -252
rect 546 -266 574 -252
<< via1 >>
rect 473 107 503 140
rect 473 106 503 107
rect 1053 106 1083 140
rect 473 -163 503 -130
rect 473 -164 503 -163
rect 1053 -164 1083 -130
<< metal2 >>
rect -54 106 473 140
rect 503 106 1053 140
rect 1083 106 1153 140
rect -54 -164 473 -130
rect 503 -164 1053 -130
rect 1083 -164 1153 -130
use 10T_toy_magic  10T_toy_magic_0
timestamp 1658880696
transform 1 0 94 0 1 23
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_1
timestamp 1658880696
transform 1 0 674 0 1 23
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_2
timestamp 1658880696
transform 1 0 94 0 1 -247
box -100 -19 452 251
use 10T_toy_magic  10T_toy_magic_3
timestamp 1658880696
transform 1 0 674 0 1 -247
box -100 -19 452 251
<< labels >>
rlabel poly -54 244 -24 274 1 WWL_0
rlabel poly -54 -26 -24 4 1 WWL_1
rlabel metal1 -54 230 -24 244 1 VDD
rlabel metal1 -54 -40 -24 -26 1 VDD
rlabel metal1 -54 4 -24 18 1 GND
rlabel metal1 -54 -266 -24 -252 1 GND
rlabel corelocali -6 -314 9 -284 1 RBL1_0
rlabel corelocali 531 -314 546 -284 1 RBL0_0
rlabel corelocali 574 -314 589 -284 1 RBL1_1
rlabel corelocali 1111 -314 1126 -284 1 RBL0_1
rlabel metal1 -54 -164 -24 -130 1 RWL_1
rlabel metal1 -54 106 -20 140 1 RWL1_0
rlabel metal2 -54 106 -20 140 1 RWL0_0
<< end >>
