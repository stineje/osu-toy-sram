* HSPICE file created from 10T_toy_magic.ext - technology: sky130

.option scale=5000u

.subckt x10T_toy_magic WWL RWL0 RWL1 WBL WBLb RBL0 RBL1 VDD GND
X0 junc0 junc1 VDD VDD sky130_fd_pr__special_pfet_pass ad=0 pd=0 as=2504 ps=288 w=28 l=30
X1 GND junc0 junc1 GND sky130_fd_pr__special_nfet_latch ad=0 pd=0 as=0 ps=0 w=42 l=30
X2 RWL0_junc junc0 GND GND sky130_fd_pr__special_nfet_pass ad=0 pd=0 as=9008 ps=928 w=28 l=30
X3 VDD junc0 junc1 VDD sky130_fd_pr__special_pfet_pass ad=0 pd=0 as=0 ps=0 w=28 l=30
X4 WBL WWL junc0 GND sky130_fd_pr__nfet_01v8 ad=967 pd=126 as=0 ps=0 w=28 l=30
X5 junc1 WWL WBLb GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=924 ps=122 w=28 l=30
X6 GND junc1 RWL1_junc GND sky130_fd_pr__special_nfet_pass ad=0 pd=0 as=0 ps=0 w=28 l=30
X7 RBL0 RWL0 RWL0_junc GND sky130_fd_pr__nfet_01v8 ad=1806 pd=170 as=0 ps=0 w=42 l=30
X8 junc0 junc1 GND GND sky130_fd_pr__special_nfet_latch ad=0 pd=0 as=0 ps=0 w=42 l=30
X9 RWL1_junc RWL1 RBL1 GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1806 ps=170 w=42 l=30
.ends

** hspice subcircuit dictionary
