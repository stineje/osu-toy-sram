magic
tech sky130A
magscale 1 2
timestamp 1653598015
<< error_p >>
rect 38 373 80 388
rect 16 361 90 373
rect 16 360 96 361
rect 16 352 80 360
rect 16 349 46 352
rect 72 349 80 352
rect 16 345 80 349
rect 90 345 96 360
rect 22 344 96 345
rect 64 338 80 344
rect -4 334 38 338
rect 64 334 122 338
rect -4 329 122 334
rect 183 329 211 342
rect -4 308 73 329
rect 80 308 122 329
rect 152 317 226 329
rect 152 316 227 317
rect 152 308 217 316
rect 36 303 38 308
rect 73 307 89 308
rect 66 296 89 307
rect 91 296 107 308
rect 152 304 191 308
rect 203 304 217 308
rect 152 301 217 304
rect 226 301 227 316
rect 167 300 227 301
rect 66 292 107 296
rect 183 292 213 300
rect 24 271 38 292
rect 57 276 123 292
rect -16 255 38 271
rect -16 241 0 255
rect 1 254 38 255
rect 66 262 107 276
rect 127 262 267 292
rect 1 247 61 254
rect 37 244 61 247
rect 38 241 61 244
rect 66 246 89 262
rect 174 258 213 262
rect 174 251 217 258
rect 226 251 227 258
rect 240 251 266 254
rect 66 241 80 246
rect 14 227 30 241
rect 1 191 30 227
rect 0 190 30 191
rect -2 174 30 190
rect 38 217 80 241
rect 144 236 266 251
rect 107 217 123 228
rect 125 221 141 228
rect 144 221 148 236
rect 166 221 170 236
rect 125 217 148 221
rect 38 174 68 217
rect 69 212 80 217
rect 138 216 148 217
rect 107 212 148 216
rect 174 212 211 236
rect 91 196 98 212
rect 107 202 157 212
rect 107 192 118 202
rect 138 192 157 202
rect 107 182 157 192
rect 174 200 204 212
rect 174 182 188 200
rect 138 175 148 182
rect -2 172 38 174
rect -16 167 38 172
rect -16 149 34 167
rect -16 142 38 149
rect -2 126 30 142
rect 0 125 30 126
rect 1 91 30 125
rect 38 129 68 142
rect 69 134 80 172
rect 107 166 123 175
rect 125 166 148 175
rect 174 174 180 182
rect 174 172 188 174
rect 107 141 123 150
rect 138 138 148 166
rect 172 142 188 172
rect 195 142 198 200
rect 202 174 204 200
rect 240 191 312 236
rect 226 190 312 191
rect 224 175 312 190
rect 223 174 312 175
rect 202 167 312 174
rect 204 149 312 167
rect 202 142 312 149
rect 38 91 80 129
rect 91 104 102 134
rect 107 124 148 138
rect 107 114 118 124
rect 138 114 148 124
rect 174 119 188 142
rect 202 119 204 142
rect 223 141 312 142
rect 224 126 312 141
rect 226 125 312 126
rect 107 104 148 114
rect 150 104 157 119
rect 174 104 204 119
rect 138 99 148 104
rect 1 89 80 91
rect 14 75 80 89
rect 107 88 123 99
rect 125 88 148 99
rect 174 95 207 104
rect 35 70 80 75
rect 138 83 148 88
rect 170 83 207 95
rect 240 83 312 125
rect 138 77 207 83
rect 35 69 89 70
rect 1 61 89 69
rect 38 58 89 61
rect 138 62 213 77
rect 38 54 107 58
rect 138 54 202 62
rect 207 54 209 62
rect 24 51 38 54
rect 66 51 107 54
rect 16 40 107 51
rect 123 40 179 54
rect 16 34 179 40
rect 207 34 263 54
rect 16 24 263 34
rect 66 9 89 24
rect 91 9 107 24
rect 146 15 226 24
rect -4 -11 38 9
rect 73 8 122 9
rect 80 -11 122 8
rect 146 8 187 15
rect 199 8 213 15
rect 146 0 213 8
rect 163 -1 223 0
rect -4 -21 122 -11
rect 12 -29 90 -21
rect 179 -26 207 -1
rect 12 -30 96 -29
rect 12 -37 46 -30
rect 72 -37 80 -30
rect 12 -45 80 -37
rect 90 -45 96 -30
rect 22 -46 96 -45
rect 38 -71 80 -46
<< nwell >>
rect 144 83 240 236
<< pwell >>
rect 12 304 106 357
rect 12 263 92 304
rect 182 301 211 316
rect 12 257 106 263
rect 0 200 106 257
rect 183 258 207 260
rect 183 243 211 258
rect -26 116 106 200
rect 0 61 106 116
rect 12 53 106 61
rect 179 60 207 70
rect 12 14 92 53
rect 12 -45 106 14
rect 179 0 207 15
<< nmos >>
rect 38 308 80 338
rect 183 262 211 292
rect 179 24 207 54
rect 38 -21 80 9
<< npd >>
rect 38 182 80 212
rect 38 104 80 134
<< npass >>
rect 38 262 66 292
rect 38 24 66 54
<< ppu >>
rect 174 182 202 212
rect 174 104 202 134
<< ndiff >>
rect 38 338 80 345
rect 38 303 80 308
rect 38 292 66 303
rect 183 292 211 301
rect 38 255 66 262
rect 0 241 66 255
rect 183 258 211 262
rect 0 174 14 241
tri 61 220 71 230 se
rect 71 220 80 237
rect 38 212 80 220
rect 38 174 80 182
rect 14 142 80 174
rect 0 75 14 142
rect 38 134 80 142
rect 38 96 80 104
rect 70 79 80 96
rect 0 61 66 75
rect 38 54 66 61
rect 179 54 207 62
rect 38 14 66 24
rect 179 15 207 24
rect 38 9 80 14
rect 38 -30 80 -21
<< pdiff >>
rect 174 212 202 221
rect 174 174 202 182
rect 174 142 226 174
rect 174 134 202 142
rect 174 95 202 104
tri 174 83 186 95 nw
<< ndiffc >>
rect 38 345 80 360
rect 183 301 211 316
rect 183 243 211 258
rect 38 230 71 237
rect 38 220 61 230
tri 61 220 71 230 nw
rect 0 142 14 174
rect 38 79 70 96
rect 179 62 207 77
rect 179 0 207 15
rect 38 -45 80 -30
<< pdiffc >>
rect 174 221 202 236
rect 226 142 240 174
tri 174 83 186 95 se
rect 186 83 202 95
<< poly >>
rect 16 308 38 338
rect 80 308 98 338
rect 16 262 38 292
rect 66 262 73 292
rect 152 262 183 292
rect 211 262 270 292
rect 16 182 38 212
rect 80 182 107 212
rect 141 182 174 212
rect 202 182 224 212
rect 16 104 38 134
rect 80 104 107 134
rect 141 104 174 134
rect 202 104 224 134
rect 240 54 270 262
rect 16 24 38 54
rect 66 24 73 54
rect 146 24 179 54
rect 207 24 270 54
rect 16 -21 38 9
rect 80 -21 96 9
<< polycont >>
rect 73 262 107 292
rect 107 182 141 212
rect 107 104 141 134
rect 73 24 107 54
<< corelocali >>
rect 16 345 38 360
rect 80 345 90 360
rect 152 301 183 316
rect 211 301 226 316
rect 14 262 73 273
rect 107 262 226 273
rect 14 258 226 262
rect 14 245 183 258
rect 14 237 71 245
rect 14 220 38 237
tri 71 230 86 245 nw
rect 170 243 183 245
rect 211 243 226 258
rect 170 236 226 243
rect 170 221 174 236
rect 202 221 226 236
rect 14 219 60 220
tri 60 219 61 220 nw
rect 170 219 226 221
rect 0 174 14 191
tri 63 182 98 217 se
rect 98 212 142 217
rect 98 182 107 212
rect 141 182 142 212
rect 0 125 14 142
tri 42 161 63 182 se
rect 63 175 142 182
rect 63 161 70 175
rect 42 97 70 161
tri 70 149 96 175 nw
tri 152 141 170 159 se
rect 170 147 198 219
rect 226 175 240 191
rect 102 134 170 141
rect 102 104 107 134
rect 141 119 170 134
tri 170 119 198 147 nw
rect 226 125 240 141
rect 141 104 150 119
rect 102 99 150 104
tri 150 99 170 119 nw
rect 16 96 70 97
rect 16 79 38 96
tri 186 95 188 97 se
rect 188 95 226 97
rect 202 83 226 95
rect 16 71 70 79
tri 162 71 174 83 se
rect 174 77 226 83
rect 174 71 179 77
rect 16 62 179 71
rect 207 62 226 77
rect 16 54 226 62
rect 16 43 73 54
rect 107 43 226 54
rect 146 0 179 15
rect 207 0 226 15
rect 12 -45 38 -30
rect 80 -45 90 -30
<< viali >>
rect 223 174 240 175
rect 223 142 226 174
rect 226 142 240 174
rect 223 141 240 142
<< labels >>
rlabel poly 240 24 270 292 1 WWl
port 1 nsew signal input
rlabel poly 38 -21 80 9 1 RWL0
port 2 nsew signal input
rlabel poly 38 308 80 338 1 RWL1
port 3 nsew signal input
rlabel corelocali 146 0 179 15 1 WBL
port 4 nsew signal input
rlabel corelocali 152 301 183 316 1 WBLb
port 5 nsew signal input
rlabel corelocali 12 -45 38 -30 1 RBL0
port 6 nsew signal output
rlabel corelocali 16 345 38 360 1 RBL1
port 7 nsew signal output
rlabel locali 223 141 240 175 1 VDD
port 8 nsew power bidirectional
rlabel locali 0 142 14 174 1 GND
port 9 nsew ground bidirectional
<< end >>
