** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_32x32_xschem.sch
**.subckt 10T_32x32_xschem
x1 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_2 RWL_2 VDD GND 10T_1x32_xschem
x2 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_3 RWL_3 VDD GND 10T_1x32_xschem
x3 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_4 RWL_4 VDD GND 10T_1x32_xschem
x4 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_5 RWL_5 VDD GND 10T_1x32_xschem
x5 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_6 RWL_6 VDD GND 10T_1x32_xschem
x6 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 __UNCONNECTED_PIN__0 RWL_7 VDD GND 10T_1x32_xschem
x7 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_1 RWL_1 VDD GND 10T_1x32_xschem
x8 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_0 RWL_0 VDD GND 10T_1x32_xschem
x9 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_8 RWL_8 VDD GND 10T_1x32_xschem
x10 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_9 RWL_9 VDD GND 10T_1x32_xschem
x11 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_12 RWL_12 VDD GND 10T_1x32_xschem
x12 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_13 RWL_13 VDD GND 10T_1x32_xschem
x13 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_14 RWL_14 VDD GND 10T_1x32_xschem
x14 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_15 RWL_15 VDD GND 10T_1x32_xschem
x15 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_16 RWL_16 VDD GND 10T_1x32_xschem
x16 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_17 RWL_17 VDD GND 10T_1x32_xschem
x17 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_11 RWL_11 VDD GND 10T_1x32_xschem
x18 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_10 RWL_10 VDD GND 10T_1x32_xschem
x19 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_18 RWL_18 VDD GND 10T_1x32_xschem
x20 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_19 RWL_19 VDD GND 10T_1x32_xschem
x21 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_22 RWL_22 VDD GND 10T_1x32_xschem
x22 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_23 RWL_23 VDD GND 10T_1x32_xschem
x23 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_24 RWL_24 VDD GND 10T_1x32_xschem
x24 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_25 RWL_25 VDD GND 10T_1x32_xschem
x25 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_26 RWL_26 VDD GND 10T_1x32_xschem
x26 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_27 RWL_27 VDD GND 10T_1x32_xschem
x27 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_21 RWL_21 VDD GND 10T_1x32_xschem
x28 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_20 RWL_20 VDD GND 10T_1x32_xschem
x29 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_28 RWL_28 VDD GND 10T_1x32_xschem
x30 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_29 RWL_29 VDD GND 10T_1x32_xschem
x31 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_30 RWL_30 VDD GND 10T_1x32_xschem
x32 RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18 RBL0_26 WBL_26 WBL_2
+ RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11 WBLb_30 WBLb_22 RBL0_31
+ RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13 RBL1_5 WBL_4 RBL1_20
+ WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27 RBL1_3 WBLb_5 WBLb_13
+ RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29 WBLb_18 RBL0_21 WBLb_10
+ RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9 WBLb_24 WBLb_16 RBL1_23
+ RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1 WBL_13 RBL0_9 RBL0_28
+ WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19 WBL_14 RBL0_11 WBL_6
+ RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31 WBLb_23 RBL0_16 RBL0_8
+ WBLb_15 RBL0_0 WBLb_7 WWL_31 RWL_31 VDD GND 10T_1x32_xschem
**.ends

* expanding   symbol:  10T_1x32_xschem.sym # of pins=130
** sym_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_1x32_xschem.sym
** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_1x32_xschem.sch
.subckt 10T_1x32_xschem  RBL0_22 WBL_25 RBL0_30 WBL_17 WBL_9 WBL_1 RBL0_14 RBL0_6 WBL_18 RBL0_18
+ RBL0_26 WBL_26 WBL_2 RBL0_2 RBL0_10 WBL_10 WBL_19 WBL_27 RBL1_30 RBL1_22 RBL1_14 WBL_3 RBL1_6 WBL_11
+ WBLb_30 WBLb_22 RBL0_31 RBL0_23 RBL0_7 RBL0_15 WBLb_6 WBLb_14 RBL1_21 WBL_20 RBL1_29 WBL_28 WBL_12 RBL1_13
+ RBL1_5 WBL_4 RBL1_20 WBL_23 WBL_31 RBL1_28 WBL_15 RBL1_4 RBL1_12 WBL_7 WBLb_29 WBLb_21 RBL1_19 RBL1_27
+ RBL1_3 WBLb_5 WBLb_13 RBL1_11 WBL_24 WBL_16 RBL1_18 RBL1_26 WBL_8 RBL1_2 RBL1_10 WBL_0 WBLb_26 RBL0_29
+ WBLb_18 RBL0_21 WBLb_10 RBL0_5 RBL0_13 WBLb_2 RBL1_25 WBLb_25 WBLb_17 RBL1_17 WBLb_9 RBL1_1 WBLb_1 RBL1_9
+ WBLb_24 WBLb_16 RBL1_23 RBL1_31 WBLb_0 WBLb_8 RBL1_7 RBL1_15 WBL_29 WBL_21 RBL0_17 RBL0_25 WBL_5 RBL0_1
+ WBL_13 RBL0_9 RBL0_28 WBLb_28 WBLb_20 RBL0_20 WBLb_12 WBLb_4 RBL0_4 RBL0_12 RBL0_27 WBL_30 WBL_22 RBL0_19
+ WBL_14 RBL0_11 WBL_6 RBL0_3 RBL1_24 WBLb_27 WBLb_19 RBL1_16 WBLb_11 RBL1_8 WBLb_3 RBL1_0 RBL0_24 WBLb_31
+ WBLb_23 RBL0_16 RBL0_8 WBLb_15 RBL0_0 WBLb_7 WWL RWL  VDD  GND
*.ipin WBL_1
*.opin RBL0_6
*.ipin WBL_2
*.ipin WBL_3
*.ipin WBLb_6
*.ipin WBL_4
*.ipin WBL_7
*.ipin WBLb_5
*.ipin WBL_0
*.ipin WBLb_2
*.ipin WBLb_1
*.ipin WBLb_0
*.ipin WBL_5
*.ipin WBLb_4
*.ipin WBL_6
*.ipin WBLb_3
*.ipin WBLb_7
*.ipin WWL
*.ipin RWL
*.opin RBL0_2
*.opin RBL1_6
*.opin RBL0_7
*.opin RBL1_5
*.opin RBL1_4
*.opin RBL1_3
*.opin RBL1_2
*.opin RBL0_5
*.opin RBL1_1
*.opin RBL1_7
*.opin RBL0_1
*.opin RBL0_4
*.opin RBL0_3
*.opin RBL1_0
*.opin RBL0_0
*.opin RBL0_8
*.opin RBL0_9
*.opin RBL0_10
*.opin RBL0_11
*.opin RBL0_12
*.opin RBL0_13
*.opin RBL0_14
*.opin RBL0_15
*.opin RBL1_8
*.opin RBL1_9
*.opin RBL1_10
*.opin RBL1_11
*.opin RBL1_12
*.opin RBL1_13
*.opin RBL1_14
*.opin RBL1_15
*.ipin WBL_8
*.ipin WBL_9
*.ipin WBL_10
*.ipin WBL_11
*.ipin WBL_12
*.ipin WBL_13
*.ipin WBL_14
*.ipin WBL_15
*.ipin WBLb_8
*.ipin WBLb_9
*.ipin WBLb_10
*.ipin WBLb_11
*.ipin WBLb_12
*.ipin WBLb_13
*.ipin WBLb_14
*.ipin WBLb_15
*.opin RBL0_16
*.opin RBL0_18
*.opin RBL0_19
*.opin RBL0_20
*.opin RBL0_21
*.opin RBL0_22
*.opin RBL0_17
*.opin RBL0_23
*.opin RBL1_16
*.opin RBL1_17
*.opin RBL1_18
*.opin RBL1_19
*.opin RBL1_20
*.opin RBL1_21
*.opin RBL1_22
*.opin RBL1_23
*.ipin WBL_16
*.ipin WBL_17
*.ipin WBL_18
*.ipin WBL_19
*.ipin WBL_20
*.ipin WBL_21
*.ipin WBL_22
*.ipin WBL_23
*.ipin WBLb_16
*.ipin WBLb_17
*.ipin WBLb_18
*.ipin WBLb_19
*.ipin WBLb_20
*.ipin WBLb_21
*.ipin WBLb_22
*.ipin WBLb_23
*.ipin WBL_24
*.ipin WBL_25
*.ipin WBL_26
*.ipin WBL_27
*.ipin WBL_28
*.ipin WBL_29
*.ipin WBL_30
*.ipin WBL_31
*.ipin WBLb_24
*.ipin WBLb_25
*.ipin WBLb_26
*.ipin WBLb_27
*.ipin WBLb_28
*.ipin WBLb_29
*.ipin WBLb_30
*.ipin WBLb_31
*.opin RBL0_24
*.opin RBL0_26
*.opin RBL0_25
*.opin RBL0_27
*.opin RBL0_28
*.opin RBL0_29
*.opin RBL0_30
*.opin RBL0_31
*.opin RBL1_24
*.opin RBL1_25
*.opin RBL1_26
*.opin RBL1_27
*.opin RBL1_28
*.opin RBL1_29
*.opin RBL1_30
*.opin RBL1_31
x1 WBL_1 WBL_2 WBL_3 WBLb_6 WBL_4 WBL_7 WBLb_5 WBL_0 WBLb_2 WBLb_1 WBLb_0 WBL_5 WBLb_4 WBL_6 WBLb_3
+ WBLb_7 WWL RWL RBL0_6 RBL0_2 RBL1_6 RBL0_7 RBL1_5 RBL1_4 RBL1_3 RBL1_2 RBL0_5 RBL1_1 RBL1_7 RBL0_1 RBL0_4
+ RBL0_3 RBL1_0 RBL0_0 VDD GND 10T_1x8_xschem
x2 WBL_9 WBL_10 WBL_11 WBLb_14 WBL_12 WBL_15 WBLb_13 WBL_8 WBLb_10 WBLb_9 WBLb_8 WBL_13 WBLb_12
+ WBL_14 WBLb_11 WBLb_15 WWL RWL RBL0_14 RBL0_10 RBL1_14 RBL0_15 RBL1_13 RBL1_12 RBL1_11 RBL1_10 RBL0_13
+ RBL1_9 RBL1_15 RBL0_9 RBL0_12 RBL0_11 RBL1_8 RBL0_8 VDD GND 10T_1x8_xschem
x3 WBL_17 WBL_18 WBL_19 WBLb_22 WBL_20 WBL_23 WBLb_21 WBL_16 WBLb_18 WBLb_17 WBLb_16 WBL_21 WBLb_20
+ WBL_22 WBLb_19 WBLb_23 WWL RWL RBL0_22 RBL0_18 RBL1_22 RBL0_23 RBL1_21 RBL1_20 RBL1_19 RBL1_18 RBL0_21
+ RBL1_17 RBL1_23 RBL0_17 RBL0_20 RBL0_19 RBL1_16 RBL0_16 VDD GND 10T_1x8_xschem
x4 WBL_25 WBL_26 WBL_27 WBLb_30 WBL_28 WBL_31 WBLb_29 WBL_24 WBLb_26 WBLb_25 WBLb_24 WBL_29 WBLb_28
+ WBL_30 WBLb_27 WBLb_31 WWL RWL RBL0_30 RBL0_26 RBL1_30 RBL0_31 RBL1_29 RBL1_28 RBL1_27 RBL1_26 RBL0_29
+ RBL1_25 RBL1_31 RBL0_25 RBL0_28 RBL0_27 RBL1_24 RBL0_24 VDD GND 10T_1x8_xschem
.ends


* expanding   symbol:  10T_1x8_xschem.sym # of pins=34
** sym_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_1x8_xschem.sym
** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_1x8_xschem.sch
.subckt 10T_1x8_xschem  WBL_1 WBL_2 WBL_3 WBLb_6 WBL_4 WBL_7 WBLb_5 WBL_0 WBLb_2 WBLb_1 WBLb_0 WBL_5
+ WBLb_4 WBL_6 WBLb_3 WBLb_7 WWL RWL RBL0_6 RBL0_2 RBL1_6 RBL0_7 RBL1_5 RBL1_4 RBL1_3 RBL1_2 RBL0_5 RBL1_1
+ RBL1_7 RBL0_1 RBL0_4 RBL0_3 RBL1_0 RBL0_0  VDD  GND
*.ipin WBLb_0
*.opin RBL0_0
*.ipin WBL_0
*.ipin WBLb_1
*.ipin WBL_1
*.ipin WBLb_2
*.ipin WBL_2
*.ipin WBLb_3
*.ipin WBL_3
*.ipin WBLb_4
*.ipin WBL_4
*.ipin WBL_5
*.ipin WBLb_5
*.ipin WBL_6
*.ipin WBLb_6
*.ipin WBLb_7
*.ipin WBL_7
*.opin RBL1_0
*.opin RBL0_1
*.opin RBL1_1
*.opin RBL0_2
*.opin RBL1_2
*.opin RBL0_3
*.opin RBL1_3
*.opin RBL0_4
*.opin RBL1_4
*.opin RBL0_5
*.opin RBL1_5
*.opin RBL0_6
*.opin RBL1_6
*.opin RBL0_7
*.opin RBL1_7
*.ipin WWL
*.ipin RWL
*  x1 -  10T-toy  IS MISSING !!!!
x1 WWL WBL_0 RBL0_0 RBL1_0 WBLb_0 RWL RWL VDD GND 10T_toy_xschem
x2 WWL WBL_1 RBL0_1 RBL1_1 WBLb_1 RWL RWL VDD GND 10T_toy_xschem
x3 WWL WBL_2 RBL0_2 RBL1_2 WBLb_2 RWL RWL VDD GND 10T_toy_xschem
x4 WWL WBL_3 RBL0_3 RBL1_3 WBLb_3 RWL RWL VDD GND 10T_toy_xschem
x5 WWL WBL_4 RBL0_4 RBL1_4 WBLb_4 RWL RWL VDD GND 10T_toy_xschem
x6 WWL WBL_5 RBL0_5 RBL1_5 WBLb_5 RWL RWL VDD GND 10T_toy_xschem
x7 WWL WBL_6 RBL0_6 RBL1_6 WBLb_6 RWL RWL VDD GND 10T_toy_xschem
x8 WWL WBL_7 RBL0_7 RBL1_7 WBLb_7 RWL RWL VDD GND 10T_toy_xschem
.ends


* expanding   symbol:  10T_toy_xschem.sym # of pins=7
** sym_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_toy_xschem.sym
** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/10T_toy_xschem.sch
.subckt 10T_toy_xschem  WWL WBL RBL0 RBL1 WBLb RWL0 RWL1  VDD  GND
*.ipin WWL
*.ipin RWL0
*.ipin RWL1
*.ipin WBL
*.ipin WBLb
*.opin RBL0
*.opin RBL1
x1 net1 net2 VDD GND INVX1
x2 net2 net1 VDD GND INVX1
XM1 net2 WWL WBL GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 WBLb WWL net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 RBL0 RWL0 net3 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.21 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 RBL1 RWL1 net4 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.21 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  INVX1.sym # of pins=2
** sym_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/INVX1.sym
** sch_path: /home/abishek/SRAM_WORK/osu-toy-sram/custom_layout/INVX1.sch
.subckt INVX1  Y A  VDD  GND
*.ipin A
*.opin Y
XM1 Y A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.21 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.14 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
