magic
tech sky130A
magscale 1 2
timestamp 1654632733
<< error_s >>
rect 29 164 56 274
rect 28 152 56 164
rect 57 215 85 274
rect 94 231 100 274
rect 93 221 100 231
rect 109 271 122 274
rect 109 221 148 271
rect 174 270 327 316
rect 156 244 348 270
rect 152 230 168 231
rect 219 230 270 244
rect 220 228 284 230
rect 327 228 342 244
rect 93 217 148 221
rect 152 217 167 221
rect 93 215 167 217
rect 174 217 342 228
rect 174 215 348 217
rect 57 207 128 215
rect 57 195 102 207
rect 109 195 128 207
rect 57 187 128 195
rect 136 187 137 215
rect 148 213 348 215
rect 356 213 386 267
rect 394 217 395 227
rect 410 217 423 274
rect 394 213 423 217
rect 148 211 423 213
rect 148 203 436 211
rect 148 191 397 203
rect 402 191 436 203
rect 148 187 436 191
rect 57 152 85 187
rect 93 171 100 187
rect 28 136 85 152
rect 94 164 100 171
rect 109 183 436 187
rect 109 178 386 183
rect 94 139 108 164
rect 109 139 148 178
rect 174 148 386 178
rect 394 167 395 183
rect 410 162 423 183
rect 189 145 386 148
rect 94 136 148 139
rect 28 131 148 136
rect 182 142 386 145
rect 28 127 122 131
rect 182 129 193 142
rect 28 120 134 127
rect 28 118 85 120
rect 94 118 134 120
rect 28 111 134 118
rect 182 111 193 127
rect 198 122 208 142
rect 218 122 232 142
rect 235 129 244 142
rect 260 129 269 142
rect 198 111 232 122
rect 235 111 237 127
rect 260 111 269 127
rect 276 122 286 142
rect 296 122 310 142
rect 311 129 322 142
rect 356 127 386 142
rect 401 139 423 162
rect 276 111 310 122
rect 311 111 322 127
rect 370 111 386 127
rect 395 134 423 139
rect 429 134 439 150
rect 440 134 467 274
rect 468 134 496 274
rect 395 118 496 134
rect 395 116 423 118
rect 426 116 467 118
rect 468 116 496 118
rect 395 111 496 116
rect 28 102 152 111
rect 28 100 85 102
rect 27 84 85 100
rect 94 93 152 102
rect 198 95 205 102
rect 276 95 306 106
rect 356 100 496 111
rect 497 152 525 274
rect 526 215 554 274
rect 563 231 569 274
rect 562 221 569 231
rect 578 271 591 274
rect 578 221 617 271
rect 643 270 796 316
rect 625 244 817 270
rect 621 230 637 231
rect 688 230 739 244
rect 689 228 753 230
rect 796 228 811 244
rect 562 217 617 221
rect 621 217 636 221
rect 562 215 636 217
rect 643 217 811 228
rect 643 215 817 217
rect 526 207 597 215
rect 526 195 571 207
rect 578 195 597 207
rect 526 187 597 195
rect 605 187 606 215
rect 617 213 817 215
rect 825 213 855 267
rect 863 217 864 227
rect 879 217 892 274
rect 863 213 892 217
rect 617 211 892 213
rect 617 203 905 211
rect 617 191 866 203
rect 871 191 905 203
rect 617 187 905 191
rect 526 152 554 187
rect 562 171 569 187
rect 497 136 554 152
rect 563 164 569 171
rect 578 183 905 187
rect 578 178 855 183
rect 563 139 577 164
rect 578 139 617 178
rect 643 148 855 178
rect 863 167 864 183
rect 879 162 892 183
rect 658 145 855 148
rect 563 136 617 139
rect 497 131 617 136
rect 651 142 855 145
rect 497 127 591 131
rect 651 129 662 142
rect 497 120 603 127
rect 497 118 554 120
rect 563 118 603 120
rect 497 111 603 118
rect 651 111 662 127
rect 667 122 677 142
rect 687 122 701 142
rect 704 129 713 142
rect 729 129 738 142
rect 667 111 701 122
rect 704 111 706 127
rect 729 111 738 127
rect 745 122 755 142
rect 765 122 779 142
rect 780 129 791 142
rect 825 127 855 142
rect 870 139 892 162
rect 745 111 779 122
rect 780 111 791 127
rect 839 111 855 127
rect 864 134 892 139
rect 898 134 908 150
rect 909 134 936 274
rect 937 162 951 274
rect 952 162 965 274
rect 937 134 965 162
rect 864 118 965 134
rect 864 116 892 118
rect 895 116 936 118
rect 937 116 965 118
rect 864 111 965 116
rect 497 102 621 111
rect 497 100 554 102
rect 356 95 423 100
rect 356 93 390 95
rect 395 93 423 95
rect 94 84 164 93
rect 340 84 423 93
rect 429 84 554 100
rect 563 93 621 102
rect 667 95 674 102
rect 745 95 775 106
rect 825 100 965 111
rect 825 95 892 100
rect 825 93 859 95
rect 864 93 892 95
rect 563 84 633 93
rect 809 84 892 93
rect 898 84 965 100
rect 0 42 85 84
rect 89 72 223 84
rect 281 72 423 84
rect 89 70 236 72
rect 27 26 28 42
rect 29 0 85 42
rect 29 -106 56 0
rect 28 -118 56 -106
rect 57 -55 85 0
rect 94 61 134 70
rect 94 49 122 61
rect 94 -39 100 49
rect 93 -49 100 -39
rect 109 46 122 49
rect 109 20 148 46
rect 156 42 166 51
rect 169 46 236 70
rect 268 70 423 72
rect 268 46 348 70
rect 370 61 386 70
rect 395 49 423 70
rect 169 42 348 46
rect 356 42 386 46
rect 109 1 122 20
rect 155 18 327 42
rect 335 20 386 42
rect 335 18 365 20
rect 155 4 349 18
rect 109 -49 148 1
rect 174 0 327 4
rect 156 -26 348 0
rect 152 -40 168 -39
rect 219 -40 270 -26
rect 220 -42 284 -40
rect 235 -43 269 -42
rect 93 -53 148 -49
rect 152 -53 167 -49
rect 93 -55 167 -53
rect 57 -63 128 -55
rect 57 -75 102 -63
rect 109 -75 128 -63
rect 57 -83 128 -75
rect 136 -83 137 -55
rect 148 -62 198 -55
rect 236 -62 268 -43
rect 327 -53 342 -26
rect 327 -57 348 -53
rect 356 -57 386 -3
rect 394 -53 395 -43
rect 410 -53 423 49
rect 440 46 554 84
rect 558 72 692 84
rect 750 72 892 84
rect 558 70 705 72
rect 429 26 554 46
rect 429 0 467 26
rect 394 -57 423 -53
rect 327 -59 423 -57
rect 306 -62 436 -59
rect 148 -64 243 -62
rect 261 -64 436 -62
rect 148 -68 210 -64
rect 291 -67 436 -64
rect 148 -71 263 -68
rect 148 -78 210 -71
rect 291 -78 397 -67
rect 148 -79 397 -78
rect 402 -79 436 -67
rect 148 -83 436 -79
rect 57 -118 85 -83
rect 93 -99 100 -83
rect 28 -134 85 -118
rect 94 -106 100 -99
rect 109 -87 436 -83
rect 109 -92 386 -87
rect 94 -131 108 -106
rect 109 -131 148 -92
rect 315 -96 386 -92
rect 198 -118 228 -109
rect 291 -116 306 -109
rect 327 -118 386 -96
rect 394 -103 395 -87
rect 410 -108 423 -87
rect 174 -122 386 -118
rect 189 -125 386 -122
rect 94 -134 148 -131
rect 28 -139 148 -134
rect 182 -128 386 -125
rect 28 -143 122 -139
rect 182 -141 193 -128
rect 28 -150 134 -143
rect 28 -152 85 -150
rect 94 -152 134 -150
rect 28 -159 134 -152
rect 182 -159 193 -143
rect 198 -148 208 -128
rect 218 -148 232 -128
rect 235 -141 244 -128
rect 260 -141 269 -128
rect 198 -159 232 -148
rect 235 -159 237 -143
rect 260 -159 269 -143
rect 276 -148 286 -128
rect 296 -148 310 -128
rect 311 -141 322 -128
rect 356 -143 386 -128
rect 401 -131 423 -108
rect 276 -159 310 -148
rect 311 -159 322 -143
rect 370 -159 386 -143
rect 395 -136 423 -131
rect 429 -136 439 -120
rect 440 -136 467 0
rect 468 -136 496 26
rect 395 -152 496 -136
rect 395 -154 423 -152
rect 429 -154 463 -152
rect 468 -154 496 -152
rect 395 -159 496 -154
rect 28 -168 152 -159
rect 28 -170 85 -168
rect 27 -186 85 -170
rect 94 -177 152 -168
rect 198 -175 205 -168
rect 276 -175 306 -164
rect 356 -170 496 -159
rect 497 0 554 26
rect 497 -118 525 0
rect 526 -55 554 0
rect 563 61 603 70
rect 563 49 591 61
rect 563 -39 569 49
rect 562 -49 569 -39
rect 578 46 591 49
rect 578 20 617 46
rect 625 42 635 51
rect 638 46 705 70
rect 737 70 892 72
rect 737 46 817 70
rect 839 61 855 70
rect 864 49 892 70
rect 638 42 817 46
rect 825 42 855 46
rect 578 1 591 20
rect 624 18 796 42
rect 804 20 855 42
rect 804 18 834 20
rect 624 4 818 18
rect 578 -49 617 1
rect 643 0 796 4
rect 625 -26 817 0
rect 621 -40 637 -39
rect 688 -40 739 -26
rect 689 -42 753 -40
rect 704 -43 738 -42
rect 562 -53 617 -49
rect 621 -53 636 -49
rect 562 -55 636 -53
rect 526 -63 597 -55
rect 526 -75 571 -63
rect 578 -75 597 -63
rect 526 -83 597 -75
rect 605 -83 606 -55
rect 617 -62 667 -55
rect 705 -62 737 -43
rect 796 -53 811 -26
rect 796 -57 817 -53
rect 825 -57 855 -3
rect 863 -53 864 -43
rect 879 -53 892 49
rect 909 46 978 84
rect 898 42 978 46
rect 898 26 951 42
rect 898 0 936 26
rect 863 -57 892 -53
rect 796 -59 892 -57
rect 775 -62 905 -59
rect 617 -64 712 -62
rect 730 -64 905 -62
rect 617 -68 679 -64
rect 760 -67 905 -64
rect 617 -71 732 -68
rect 617 -78 679 -71
rect 760 -78 866 -67
rect 617 -79 866 -78
rect 871 -79 905 -67
rect 617 -83 905 -79
rect 526 -118 554 -83
rect 562 -99 569 -83
rect 497 -134 554 -118
rect 563 -106 569 -99
rect 578 -87 905 -83
rect 578 -92 855 -87
rect 563 -131 577 -106
rect 578 -131 617 -92
rect 784 -96 855 -92
rect 667 -118 697 -109
rect 760 -116 775 -109
rect 796 -118 855 -96
rect 863 -103 864 -87
rect 879 -108 892 -87
rect 643 -122 855 -118
rect 658 -125 855 -122
rect 563 -134 617 -131
rect 497 -139 617 -134
rect 651 -128 855 -125
rect 497 -143 591 -139
rect 651 -141 662 -128
rect 497 -150 603 -143
rect 497 -152 554 -150
rect 563 -152 603 -150
rect 497 -159 603 -152
rect 651 -159 662 -143
rect 667 -148 677 -128
rect 687 -148 701 -128
rect 704 -141 713 -128
rect 729 -141 738 -128
rect 667 -159 701 -148
rect 704 -159 706 -143
rect 729 -159 738 -143
rect 745 -148 755 -128
rect 765 -148 779 -128
rect 780 -141 791 -128
rect 825 -143 855 -128
rect 870 -131 892 -108
rect 745 -159 779 -148
rect 780 -159 791 -143
rect 839 -159 855 -143
rect 864 -136 892 -131
rect 898 -136 908 -120
rect 909 -136 936 0
rect 937 -108 951 26
rect 952 -108 965 42
rect 937 -136 965 -108
rect 864 -152 965 -136
rect 864 -154 892 -152
rect 898 -154 932 -152
rect 937 -154 965 -152
rect 864 -159 965 -154
rect 497 -168 621 -159
rect 497 -170 554 -168
rect 356 -175 423 -170
rect 356 -177 390 -175
rect 395 -177 423 -175
rect 94 -186 164 -177
rect 340 -186 423 -177
rect 429 -186 459 -170
rect 0 -228 85 -186
rect 89 -198 223 -186
rect 281 -198 423 -186
rect 89 -200 236 -198
rect 27 -244 28 -228
rect 29 -266 85 -228
rect 94 -209 134 -200
rect 94 -221 122 -209
rect 94 -266 100 -221
rect 109 -228 122 -221
rect 156 -228 166 -219
rect 109 -242 148 -228
rect 155 -229 166 -228
rect 169 -228 236 -200
rect 268 -200 423 -198
rect 268 -228 348 -200
rect 370 -209 386 -200
rect 395 -221 423 -200
rect 109 -266 122 -242
rect 155 -265 163 -229
rect 169 -236 185 -228
rect 236 -232 243 -228
rect 261 -232 268 -228
rect 236 -236 268 -232
rect 169 -252 335 -236
rect 341 -242 386 -228
rect 341 -252 365 -242
rect 183 -265 321 -252
rect 341 -265 349 -252
rect 219 -266 285 -265
rect 410 -266 423 -221
rect 467 -228 554 -170
rect 563 -177 621 -168
rect 667 -175 674 -168
rect 745 -175 775 -164
rect 825 -170 965 -159
rect 825 -175 892 -170
rect 825 -177 859 -175
rect 864 -177 892 -175
rect 563 -186 633 -177
rect 809 -186 892 -177
rect 898 -186 928 -170
rect 936 -186 965 -170
rect 558 -198 692 -186
rect 750 -198 892 -186
rect 558 -200 705 -198
rect 50 -270 80 -266
rect 220 -268 284 -266
rect 429 -270 459 -228
rect 467 -244 468 -228
rect 469 -244 554 -228
rect 469 -266 496 -244
rect 497 -266 554 -244
rect 563 -209 603 -200
rect 563 -221 591 -209
rect 563 -266 569 -221
rect 578 -228 591 -221
rect 625 -228 635 -219
rect 578 -242 617 -228
rect 624 -229 635 -228
rect 638 -228 705 -200
rect 737 -200 892 -198
rect 737 -228 817 -200
rect 839 -209 855 -200
rect 864 -221 892 -200
rect 578 -266 591 -242
rect 624 -265 632 -229
rect 638 -236 654 -228
rect 705 -232 712 -228
rect 730 -232 737 -228
rect 705 -236 737 -232
rect 638 -252 804 -236
rect 810 -242 855 -228
rect 810 -252 834 -242
rect 652 -265 790 -252
rect 810 -265 818 -252
rect 688 -266 754 -265
rect 879 -266 892 -221
rect 936 -204 978 -186
rect 936 -220 939 -204
rect 944 -220 978 -204
rect 936 -228 978 -220
rect 519 -270 549 -266
rect 689 -268 753 -266
rect 898 -270 928 -228
rect 936 -244 937 -228
rect 952 -266 965 -228
<< poly >>
rect 483 244 497 274
rect 483 -26 497 4
<< corelocali >>
rect 439 -59 454 135
rect 908 -62 923 135
use 10T_toy_magic  10T_toy_magic_3
timestamp 1654632086
transform 1 0 545 0 1 -247
box -76 -23 433 293
use 10T_toy_magic  10T_toy_magic_2
timestamp 1654632086
transform 1 0 76 0 1 -247
box -76 -23 433 293
use 10T_toy_magic  10T_toy_magic_1
timestamp 1654632086
transform 1 0 545 0 1 23
box -76 -23 433 293
use 10T_toy_magic  10T_toy_magic_0
timestamp 1654632086
transform 1 0 76 0 1 23
box -76 -23 433 293
<< end >>
