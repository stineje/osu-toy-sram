magic
tech sky130A
magscale 1 2
timestamp 1656028469
<< error_s >>
rect 15 4304 28 4320
rect 117 4318 130 4320
rect 83 4304 98 4318
rect 107 4304 137 4318
rect 198 4316 351 4362
rect 180 4304 372 4316
rect 415 4304 445 4318
rect 451 4304 464 4320
rect 552 4304 565 4320
rect 595 4304 608 4320
rect 697 4318 710 4320
rect 663 4304 678 4318
rect 687 4304 717 4318
rect 778 4316 931 4362
rect 760 4304 952 4316
rect 995 4304 1025 4318
rect 1031 4304 1044 4320
rect 1132 4304 1145 4320
rect 1175 4304 1188 4320
rect 1277 4318 1290 4320
rect 1243 4304 1258 4318
rect 1267 4304 1297 4318
rect 1358 4316 1511 4362
rect 1340 4304 1532 4316
rect 1575 4304 1605 4318
rect 1611 4304 1624 4320
rect 1712 4304 1725 4320
rect 1755 4304 1768 4320
rect 1857 4318 1870 4320
rect 1823 4304 1838 4318
rect 1847 4304 1877 4318
rect 1938 4316 2091 4362
rect 1920 4304 2112 4316
rect 2155 4304 2185 4318
rect 2191 4304 2204 4320
rect 2292 4304 2305 4320
rect 2335 4304 2348 4320
rect 2437 4318 2450 4320
rect 2403 4304 2418 4318
rect 2427 4304 2457 4318
rect 2518 4316 2671 4362
rect 2500 4304 2692 4316
rect 2735 4304 2765 4318
rect 2771 4304 2784 4320
rect 2872 4304 2885 4320
rect 2915 4304 2928 4320
rect 3017 4318 3030 4320
rect 2983 4304 2998 4318
rect 3007 4304 3037 4318
rect 3098 4316 3251 4362
rect 3080 4304 3272 4316
rect 3315 4304 3345 4318
rect 3351 4304 3364 4320
rect 3452 4304 3465 4320
rect 3495 4304 3508 4320
rect 3597 4318 3610 4320
rect 3563 4304 3578 4318
rect 3587 4304 3617 4318
rect 3678 4316 3831 4362
rect 3660 4304 3852 4316
rect 3895 4304 3925 4318
rect 3931 4304 3944 4320
rect 4032 4304 4045 4320
rect 4075 4304 4088 4320
rect 4177 4318 4190 4320
rect 4143 4304 4158 4318
rect 4167 4304 4197 4318
rect 4258 4316 4411 4362
rect 4240 4304 4432 4316
rect 4475 4304 4505 4318
rect 4511 4304 4524 4320
rect 4612 4304 4625 4320
rect 0 4290 4625 4304
rect 15 4186 28 4290
rect 73 4268 74 4278
rect 89 4268 102 4278
rect 73 4264 102 4268
rect 107 4264 137 4290
rect 155 4276 171 4278
rect 243 4276 296 4290
rect 244 4274 308 4276
rect 351 4274 366 4290
rect 415 4287 445 4290
rect 415 4284 451 4287
rect 381 4276 397 4278
rect 155 4264 170 4268
rect 73 4262 170 4264
rect 198 4262 366 4274
rect 382 4264 397 4268
rect 415 4265 454 4284
rect 473 4278 480 4279
rect 479 4271 480 4278
rect 463 4268 464 4271
rect 479 4268 492 4271
rect 415 4264 445 4265
rect 454 4264 460 4265
rect 463 4264 492 4268
rect 382 4263 492 4264
rect 382 4262 498 4263
rect 57 4254 108 4262
rect 57 4242 82 4254
rect 89 4242 108 4254
rect 139 4254 189 4262
rect 139 4246 155 4254
rect 162 4252 189 4254
rect 198 4252 419 4262
rect 162 4242 419 4252
rect 448 4254 498 4262
rect 448 4245 464 4254
rect 57 4234 108 4242
rect 155 4234 419 4242
rect 445 4242 464 4245
rect 471 4242 498 4254
rect 445 4234 498 4242
rect 73 4226 74 4234
rect 89 4226 102 4234
rect 73 4218 89 4226
rect 70 4211 89 4214
rect 70 4202 92 4211
rect 43 4192 92 4202
rect 43 4186 73 4192
rect 92 4187 97 4192
rect 15 4170 89 4186
rect 107 4178 137 4234
rect 172 4224 380 4234
rect 415 4230 460 4234
rect 463 4233 464 4234
rect 479 4233 492 4234
rect 198 4194 387 4224
rect 213 4191 387 4194
rect 206 4188 387 4191
rect 15 4168 28 4170
rect 43 4168 77 4170
rect 15 4152 89 4168
rect 116 4164 129 4178
rect 144 4164 160 4180
rect 206 4175 217 4188
rect -1 4130 0 4146
rect 15 4130 28 4152
rect 43 4130 73 4152
rect 116 4148 178 4164
rect 206 4157 217 4173
rect 222 4168 232 4188
rect 242 4168 256 4188
rect 259 4175 268 4188
rect 284 4175 293 4188
rect 222 4157 256 4168
rect 259 4157 268 4173
rect 284 4157 293 4173
rect 300 4168 310 4188
rect 320 4168 334 4188
rect 335 4175 346 4188
rect 300 4157 334 4168
rect 335 4157 346 4173
rect 392 4164 408 4180
rect 415 4178 445 4230
rect 479 4226 480 4233
rect 464 4218 480 4226
rect 451 4186 464 4205
rect 479 4186 509 4202
rect 451 4170 525 4186
rect 451 4168 464 4170
rect 479 4168 513 4170
rect 116 4146 129 4148
rect 144 4146 178 4148
rect 116 4130 178 4146
rect 222 4141 238 4144
rect 300 4141 330 4152
rect 378 4148 424 4164
rect 451 4152 525 4168
rect 378 4146 412 4148
rect 377 4130 424 4146
rect 451 4130 464 4152
rect 479 4130 509 4152
rect 536 4130 537 4146
rect 552 4130 565 4290
rect 595 4186 608 4290
rect 653 4268 654 4278
rect 669 4268 682 4278
rect 653 4264 682 4268
rect 687 4264 717 4290
rect 735 4276 751 4278
rect 823 4276 876 4290
rect 824 4274 888 4276
rect 931 4274 946 4290
rect 995 4287 1025 4290
rect 995 4284 1031 4287
rect 961 4276 977 4278
rect 735 4264 750 4268
rect 653 4262 750 4264
rect 778 4262 946 4274
rect 962 4264 977 4268
rect 995 4265 1034 4284
rect 1053 4278 1060 4279
rect 1059 4271 1060 4278
rect 1043 4268 1044 4271
rect 1059 4268 1072 4271
rect 995 4264 1025 4265
rect 1034 4264 1040 4265
rect 1043 4264 1072 4268
rect 962 4263 1072 4264
rect 962 4262 1078 4263
rect 637 4254 688 4262
rect 637 4242 662 4254
rect 669 4242 688 4254
rect 719 4254 769 4262
rect 719 4246 735 4254
rect 742 4252 769 4254
rect 778 4252 999 4262
rect 742 4242 999 4252
rect 1028 4254 1078 4262
rect 1028 4245 1044 4254
rect 637 4234 688 4242
rect 735 4234 999 4242
rect 1025 4242 1044 4245
rect 1051 4242 1078 4254
rect 1025 4234 1078 4242
rect 653 4226 654 4234
rect 669 4226 682 4234
rect 653 4218 669 4226
rect 650 4211 669 4214
rect 650 4202 672 4211
rect 623 4192 672 4202
rect 623 4186 653 4192
rect 672 4187 677 4192
rect 595 4170 669 4186
rect 687 4178 717 4234
rect 752 4224 960 4234
rect 995 4230 1040 4234
rect 1043 4233 1044 4234
rect 1059 4233 1072 4234
rect 778 4194 967 4224
rect 793 4191 967 4194
rect 786 4188 967 4191
rect 595 4168 608 4170
rect 623 4168 657 4170
rect 595 4152 669 4168
rect 696 4164 709 4178
rect 724 4164 740 4180
rect 786 4175 797 4188
rect 579 4130 580 4146
rect 595 4130 608 4152
rect 623 4130 653 4152
rect 696 4148 758 4164
rect 786 4157 797 4173
rect 802 4168 812 4188
rect 822 4168 836 4188
rect 839 4175 848 4188
rect 864 4175 873 4188
rect 802 4157 836 4168
rect 839 4157 848 4173
rect 864 4157 873 4173
rect 880 4168 890 4188
rect 900 4168 914 4188
rect 915 4175 926 4188
rect 880 4157 914 4168
rect 915 4157 926 4173
rect 972 4164 988 4180
rect 995 4178 1025 4230
rect 1059 4226 1060 4233
rect 1044 4218 1060 4226
rect 1031 4186 1044 4205
rect 1059 4186 1089 4202
rect 1031 4170 1105 4186
rect 1031 4168 1044 4170
rect 1059 4168 1093 4170
rect 696 4146 709 4148
rect 724 4146 758 4148
rect 696 4130 758 4146
rect 802 4141 818 4144
rect 880 4141 910 4152
rect 958 4148 1004 4164
rect 1031 4152 1105 4168
rect 958 4146 992 4148
rect 957 4130 1004 4146
rect 1031 4130 1044 4152
rect 1059 4130 1089 4152
rect 1116 4130 1117 4146
rect 1132 4130 1145 4290
rect 1175 4186 1188 4290
rect 1233 4268 1234 4278
rect 1249 4268 1262 4278
rect 1233 4264 1262 4268
rect 1267 4264 1297 4290
rect 1315 4276 1331 4278
rect 1403 4276 1456 4290
rect 1404 4274 1468 4276
rect 1511 4274 1526 4290
rect 1575 4287 1605 4290
rect 1575 4284 1611 4287
rect 1541 4276 1557 4278
rect 1315 4264 1330 4268
rect 1233 4262 1330 4264
rect 1358 4262 1526 4274
rect 1542 4264 1557 4268
rect 1575 4265 1614 4284
rect 1633 4278 1640 4279
rect 1639 4271 1640 4278
rect 1623 4268 1624 4271
rect 1639 4268 1652 4271
rect 1575 4264 1605 4265
rect 1614 4264 1620 4265
rect 1623 4264 1652 4268
rect 1542 4263 1652 4264
rect 1542 4262 1658 4263
rect 1217 4254 1268 4262
rect 1217 4242 1242 4254
rect 1249 4242 1268 4254
rect 1299 4254 1349 4262
rect 1299 4246 1315 4254
rect 1322 4252 1349 4254
rect 1358 4252 1579 4262
rect 1322 4242 1579 4252
rect 1608 4254 1658 4262
rect 1608 4245 1624 4254
rect 1217 4234 1268 4242
rect 1315 4234 1579 4242
rect 1605 4242 1624 4245
rect 1631 4242 1658 4254
rect 1605 4234 1658 4242
rect 1233 4226 1234 4234
rect 1249 4226 1262 4234
rect 1233 4218 1249 4226
rect 1230 4211 1249 4214
rect 1230 4202 1252 4211
rect 1203 4192 1252 4202
rect 1203 4186 1233 4192
rect 1252 4187 1257 4192
rect 1175 4170 1249 4186
rect 1267 4178 1297 4234
rect 1332 4224 1540 4234
rect 1575 4230 1620 4234
rect 1623 4233 1624 4234
rect 1639 4233 1652 4234
rect 1358 4194 1547 4224
rect 1373 4191 1547 4194
rect 1366 4188 1547 4191
rect 1175 4168 1188 4170
rect 1203 4168 1237 4170
rect 1175 4152 1249 4168
rect 1276 4164 1289 4178
rect 1304 4164 1320 4180
rect 1366 4175 1377 4188
rect 1159 4130 1160 4146
rect 1175 4130 1188 4152
rect 1203 4130 1233 4152
rect 1276 4148 1338 4164
rect 1366 4157 1377 4173
rect 1382 4168 1392 4188
rect 1402 4168 1416 4188
rect 1419 4175 1428 4188
rect 1444 4175 1453 4188
rect 1382 4157 1416 4168
rect 1419 4157 1428 4173
rect 1444 4157 1453 4173
rect 1460 4168 1470 4188
rect 1480 4168 1494 4188
rect 1495 4175 1506 4188
rect 1460 4157 1494 4168
rect 1495 4157 1506 4173
rect 1552 4164 1568 4180
rect 1575 4178 1605 4230
rect 1639 4226 1640 4233
rect 1624 4218 1640 4226
rect 1611 4186 1624 4205
rect 1639 4186 1669 4202
rect 1611 4170 1685 4186
rect 1611 4168 1624 4170
rect 1639 4168 1673 4170
rect 1276 4146 1289 4148
rect 1304 4146 1338 4148
rect 1276 4130 1338 4146
rect 1382 4141 1398 4144
rect 1460 4141 1490 4152
rect 1538 4148 1584 4164
rect 1611 4152 1685 4168
rect 1538 4146 1572 4148
rect 1537 4130 1584 4146
rect 1611 4130 1624 4152
rect 1639 4130 1669 4152
rect 1696 4130 1697 4146
rect 1712 4130 1725 4290
rect 1755 4186 1768 4290
rect 1813 4268 1814 4278
rect 1829 4268 1842 4278
rect 1813 4264 1842 4268
rect 1847 4264 1877 4290
rect 1895 4276 1911 4278
rect 1983 4276 2036 4290
rect 1984 4274 2048 4276
rect 2091 4274 2106 4290
rect 2155 4287 2185 4290
rect 2155 4284 2191 4287
rect 2121 4276 2137 4278
rect 1895 4264 1910 4268
rect 1813 4262 1910 4264
rect 1938 4262 2106 4274
rect 2122 4264 2137 4268
rect 2155 4265 2194 4284
rect 2213 4278 2220 4279
rect 2219 4271 2220 4278
rect 2203 4268 2204 4271
rect 2219 4268 2232 4271
rect 2155 4264 2185 4265
rect 2194 4264 2200 4265
rect 2203 4264 2232 4268
rect 2122 4263 2232 4264
rect 2122 4262 2238 4263
rect 1797 4254 1848 4262
rect 1797 4242 1822 4254
rect 1829 4242 1848 4254
rect 1879 4254 1929 4262
rect 1879 4246 1895 4254
rect 1902 4252 1929 4254
rect 1938 4252 2159 4262
rect 1902 4242 2159 4252
rect 2188 4254 2238 4262
rect 2188 4245 2204 4254
rect 1797 4234 1848 4242
rect 1895 4234 2159 4242
rect 2185 4242 2204 4245
rect 2211 4242 2238 4254
rect 2185 4234 2238 4242
rect 1813 4226 1814 4234
rect 1829 4226 1842 4234
rect 1813 4218 1829 4226
rect 1810 4211 1829 4214
rect 1810 4202 1832 4211
rect 1783 4192 1832 4202
rect 1783 4186 1813 4192
rect 1832 4187 1837 4192
rect 1755 4170 1829 4186
rect 1847 4178 1877 4234
rect 1912 4224 2120 4234
rect 2155 4230 2200 4234
rect 2203 4233 2204 4234
rect 2219 4233 2232 4234
rect 1938 4194 2127 4224
rect 1953 4191 2127 4194
rect 1946 4188 2127 4191
rect 1755 4168 1768 4170
rect 1783 4168 1817 4170
rect 1755 4152 1829 4168
rect 1856 4164 1869 4178
rect 1884 4164 1900 4180
rect 1946 4175 1957 4188
rect 1739 4130 1740 4146
rect 1755 4130 1768 4152
rect 1783 4130 1813 4152
rect 1856 4148 1918 4164
rect 1946 4157 1957 4173
rect 1962 4168 1972 4188
rect 1982 4168 1996 4188
rect 1999 4175 2008 4188
rect 2024 4175 2033 4188
rect 1962 4157 1996 4168
rect 1999 4157 2008 4173
rect 2024 4157 2033 4173
rect 2040 4168 2050 4188
rect 2060 4168 2074 4188
rect 2075 4175 2086 4188
rect 2040 4157 2074 4168
rect 2075 4157 2086 4173
rect 2132 4164 2148 4180
rect 2155 4178 2185 4230
rect 2219 4226 2220 4233
rect 2204 4218 2220 4226
rect 2191 4186 2204 4205
rect 2219 4186 2249 4202
rect 2191 4170 2265 4186
rect 2191 4168 2204 4170
rect 2219 4168 2253 4170
rect 1856 4146 1869 4148
rect 1884 4146 1918 4148
rect 1856 4130 1918 4146
rect 1962 4141 1978 4144
rect 2040 4141 2070 4152
rect 2118 4148 2164 4164
rect 2191 4152 2265 4168
rect 2118 4146 2152 4148
rect 2117 4130 2164 4146
rect 2191 4130 2204 4152
rect 2219 4130 2249 4152
rect 2276 4130 2277 4146
rect 2292 4130 2305 4290
rect 2335 4186 2348 4290
rect 2393 4268 2394 4278
rect 2409 4268 2422 4278
rect 2393 4264 2422 4268
rect 2427 4264 2457 4290
rect 2475 4276 2491 4278
rect 2563 4276 2616 4290
rect 2564 4274 2628 4276
rect 2671 4274 2686 4290
rect 2735 4287 2765 4290
rect 2735 4284 2771 4287
rect 2701 4276 2717 4278
rect 2475 4264 2490 4268
rect 2393 4262 2490 4264
rect 2518 4262 2686 4274
rect 2702 4264 2717 4268
rect 2735 4265 2774 4284
rect 2793 4278 2800 4279
rect 2799 4271 2800 4278
rect 2783 4268 2784 4271
rect 2799 4268 2812 4271
rect 2735 4264 2765 4265
rect 2774 4264 2780 4265
rect 2783 4264 2812 4268
rect 2702 4263 2812 4264
rect 2702 4262 2818 4263
rect 2377 4254 2428 4262
rect 2377 4242 2402 4254
rect 2409 4242 2428 4254
rect 2459 4254 2509 4262
rect 2459 4246 2475 4254
rect 2482 4252 2509 4254
rect 2518 4252 2739 4262
rect 2482 4242 2739 4252
rect 2768 4254 2818 4262
rect 2768 4245 2784 4254
rect 2377 4234 2428 4242
rect 2475 4234 2739 4242
rect 2765 4242 2784 4245
rect 2791 4242 2818 4254
rect 2765 4234 2818 4242
rect 2393 4226 2394 4234
rect 2409 4226 2422 4234
rect 2393 4218 2409 4226
rect 2390 4211 2409 4214
rect 2390 4202 2412 4211
rect 2363 4192 2412 4202
rect 2363 4186 2393 4192
rect 2412 4187 2417 4192
rect 2335 4170 2409 4186
rect 2427 4178 2457 4234
rect 2492 4224 2700 4234
rect 2735 4230 2780 4234
rect 2783 4233 2784 4234
rect 2799 4233 2812 4234
rect 2518 4194 2707 4224
rect 2533 4191 2707 4194
rect 2526 4188 2707 4191
rect 2335 4168 2348 4170
rect 2363 4168 2397 4170
rect 2335 4152 2409 4168
rect 2436 4164 2449 4178
rect 2464 4164 2480 4180
rect 2526 4175 2537 4188
rect 2319 4130 2320 4146
rect 2335 4130 2348 4152
rect 2363 4130 2393 4152
rect 2436 4148 2498 4164
rect 2526 4157 2537 4173
rect 2542 4168 2552 4188
rect 2562 4168 2576 4188
rect 2579 4175 2588 4188
rect 2604 4175 2613 4188
rect 2542 4157 2576 4168
rect 2579 4157 2588 4173
rect 2604 4157 2613 4173
rect 2620 4168 2630 4188
rect 2640 4168 2654 4188
rect 2655 4175 2666 4188
rect 2620 4157 2654 4168
rect 2655 4157 2666 4173
rect 2712 4164 2728 4180
rect 2735 4178 2765 4230
rect 2799 4226 2800 4233
rect 2784 4218 2800 4226
rect 2771 4186 2784 4205
rect 2799 4186 2829 4202
rect 2771 4170 2845 4186
rect 2771 4168 2784 4170
rect 2799 4168 2833 4170
rect 2436 4146 2449 4148
rect 2464 4146 2498 4148
rect 2436 4130 2498 4146
rect 2542 4141 2558 4144
rect 2620 4141 2650 4152
rect 2698 4148 2744 4164
rect 2771 4152 2845 4168
rect 2698 4146 2732 4148
rect 2697 4130 2744 4146
rect 2771 4130 2784 4152
rect 2799 4130 2829 4152
rect 2856 4130 2857 4146
rect 2872 4130 2885 4290
rect 2915 4186 2928 4290
rect 2973 4268 2974 4278
rect 2989 4268 3002 4278
rect 2973 4264 3002 4268
rect 3007 4264 3037 4290
rect 3055 4276 3071 4278
rect 3143 4276 3196 4290
rect 3144 4274 3208 4276
rect 3251 4274 3266 4290
rect 3315 4287 3345 4290
rect 3315 4284 3351 4287
rect 3281 4276 3297 4278
rect 3055 4264 3070 4268
rect 2973 4262 3070 4264
rect 3098 4262 3266 4274
rect 3282 4264 3297 4268
rect 3315 4265 3354 4284
rect 3373 4278 3380 4279
rect 3379 4271 3380 4278
rect 3363 4268 3364 4271
rect 3379 4268 3392 4271
rect 3315 4264 3345 4265
rect 3354 4264 3360 4265
rect 3363 4264 3392 4268
rect 3282 4263 3392 4264
rect 3282 4262 3398 4263
rect 2957 4254 3008 4262
rect 2957 4242 2982 4254
rect 2989 4242 3008 4254
rect 3039 4254 3089 4262
rect 3039 4246 3055 4254
rect 3062 4252 3089 4254
rect 3098 4252 3319 4262
rect 3062 4242 3319 4252
rect 3348 4254 3398 4262
rect 3348 4245 3364 4254
rect 2957 4234 3008 4242
rect 3055 4234 3319 4242
rect 3345 4242 3364 4245
rect 3371 4242 3398 4254
rect 3345 4234 3398 4242
rect 2973 4226 2974 4234
rect 2989 4226 3002 4234
rect 2973 4218 2989 4226
rect 2970 4211 2989 4214
rect 2970 4202 2992 4211
rect 2943 4192 2992 4202
rect 2943 4186 2973 4192
rect 2992 4187 2997 4192
rect 2915 4170 2989 4186
rect 3007 4178 3037 4234
rect 3072 4224 3280 4234
rect 3315 4230 3360 4234
rect 3363 4233 3364 4234
rect 3379 4233 3392 4234
rect 3098 4194 3287 4224
rect 3113 4191 3287 4194
rect 3106 4188 3287 4191
rect 2915 4168 2928 4170
rect 2943 4168 2977 4170
rect 2915 4152 2989 4168
rect 3016 4164 3029 4178
rect 3044 4164 3060 4180
rect 3106 4175 3117 4188
rect 2899 4130 2900 4146
rect 2915 4130 2928 4152
rect 2943 4130 2973 4152
rect 3016 4148 3078 4164
rect 3106 4157 3117 4173
rect 3122 4168 3132 4188
rect 3142 4168 3156 4188
rect 3159 4175 3168 4188
rect 3184 4175 3193 4188
rect 3122 4157 3156 4168
rect 3159 4157 3168 4173
rect 3184 4157 3193 4173
rect 3200 4168 3210 4188
rect 3220 4168 3234 4188
rect 3235 4175 3246 4188
rect 3200 4157 3234 4168
rect 3235 4157 3246 4173
rect 3292 4164 3308 4180
rect 3315 4178 3345 4230
rect 3379 4226 3380 4233
rect 3364 4218 3380 4226
rect 3351 4186 3364 4205
rect 3379 4186 3409 4202
rect 3351 4170 3425 4186
rect 3351 4168 3364 4170
rect 3379 4168 3413 4170
rect 3016 4146 3029 4148
rect 3044 4146 3078 4148
rect 3016 4130 3078 4146
rect 3122 4141 3138 4144
rect 3200 4141 3230 4152
rect 3278 4148 3324 4164
rect 3351 4152 3425 4168
rect 3278 4146 3312 4148
rect 3277 4130 3324 4146
rect 3351 4130 3364 4152
rect 3379 4130 3409 4152
rect 3436 4130 3437 4146
rect 3452 4130 3465 4290
rect 3495 4186 3508 4290
rect 3553 4268 3554 4278
rect 3569 4268 3582 4278
rect 3553 4264 3582 4268
rect 3587 4264 3617 4290
rect 3635 4276 3651 4278
rect 3723 4276 3776 4290
rect 3724 4274 3788 4276
rect 3831 4274 3846 4290
rect 3895 4287 3925 4290
rect 3895 4284 3931 4287
rect 3861 4276 3877 4278
rect 3635 4264 3650 4268
rect 3553 4262 3650 4264
rect 3678 4262 3846 4274
rect 3862 4264 3877 4268
rect 3895 4265 3934 4284
rect 3953 4278 3960 4279
rect 3959 4271 3960 4278
rect 3943 4268 3944 4271
rect 3959 4268 3972 4271
rect 3895 4264 3925 4265
rect 3934 4264 3940 4265
rect 3943 4264 3972 4268
rect 3862 4263 3972 4264
rect 3862 4262 3978 4263
rect 3537 4254 3588 4262
rect 3537 4242 3562 4254
rect 3569 4242 3588 4254
rect 3619 4254 3669 4262
rect 3619 4246 3635 4254
rect 3642 4252 3669 4254
rect 3678 4252 3899 4262
rect 3642 4242 3899 4252
rect 3928 4254 3978 4262
rect 3928 4245 3944 4254
rect 3537 4234 3588 4242
rect 3635 4234 3899 4242
rect 3925 4242 3944 4245
rect 3951 4242 3978 4254
rect 3925 4234 3978 4242
rect 3553 4226 3554 4234
rect 3569 4226 3582 4234
rect 3553 4218 3569 4226
rect 3550 4211 3569 4214
rect 3550 4202 3572 4211
rect 3523 4192 3572 4202
rect 3523 4186 3553 4192
rect 3572 4187 3577 4192
rect 3495 4170 3569 4186
rect 3587 4178 3617 4234
rect 3652 4224 3860 4234
rect 3895 4230 3940 4234
rect 3943 4233 3944 4234
rect 3959 4233 3972 4234
rect 3678 4194 3867 4224
rect 3693 4191 3867 4194
rect 3686 4188 3867 4191
rect 3495 4168 3508 4170
rect 3523 4168 3557 4170
rect 3495 4152 3569 4168
rect 3596 4164 3609 4178
rect 3624 4164 3640 4180
rect 3686 4175 3697 4188
rect 3479 4130 3480 4146
rect 3495 4130 3508 4152
rect 3523 4130 3553 4152
rect 3596 4148 3658 4164
rect 3686 4157 3697 4173
rect 3702 4168 3712 4188
rect 3722 4168 3736 4188
rect 3739 4175 3748 4188
rect 3764 4175 3773 4188
rect 3702 4157 3736 4168
rect 3739 4157 3748 4173
rect 3764 4157 3773 4173
rect 3780 4168 3790 4188
rect 3800 4168 3814 4188
rect 3815 4175 3826 4188
rect 3780 4157 3814 4168
rect 3815 4157 3826 4173
rect 3872 4164 3888 4180
rect 3895 4178 3925 4230
rect 3959 4226 3960 4233
rect 3944 4218 3960 4226
rect 3931 4186 3944 4205
rect 3959 4186 3989 4202
rect 3931 4170 4005 4186
rect 3931 4168 3944 4170
rect 3959 4168 3993 4170
rect 3596 4146 3609 4148
rect 3624 4146 3658 4148
rect 3596 4130 3658 4146
rect 3702 4141 3718 4144
rect 3780 4141 3810 4152
rect 3858 4148 3904 4164
rect 3931 4152 4005 4168
rect 3858 4146 3892 4148
rect 3857 4130 3904 4146
rect 3931 4130 3944 4152
rect 3959 4130 3989 4152
rect 4016 4130 4017 4146
rect 4032 4130 4045 4290
rect 4075 4186 4088 4290
rect 4133 4268 4134 4278
rect 4149 4268 4162 4278
rect 4133 4264 4162 4268
rect 4167 4264 4197 4290
rect 4215 4276 4231 4278
rect 4303 4276 4356 4290
rect 4304 4274 4368 4276
rect 4411 4274 4426 4290
rect 4475 4287 4505 4290
rect 4475 4284 4511 4287
rect 4441 4276 4457 4278
rect 4215 4264 4230 4268
rect 4133 4262 4230 4264
rect 4258 4262 4426 4274
rect 4442 4264 4457 4268
rect 4475 4265 4514 4284
rect 4533 4278 4540 4279
rect 4539 4271 4540 4278
rect 4523 4268 4524 4271
rect 4539 4268 4552 4271
rect 4475 4264 4505 4265
rect 4514 4264 4520 4265
rect 4523 4264 4552 4268
rect 4442 4263 4552 4264
rect 4442 4262 4558 4263
rect 4117 4254 4168 4262
rect 4117 4242 4142 4254
rect 4149 4242 4168 4254
rect 4199 4254 4249 4262
rect 4199 4246 4215 4254
rect 4222 4252 4249 4254
rect 4258 4252 4479 4262
rect 4222 4242 4479 4252
rect 4508 4254 4558 4262
rect 4508 4245 4524 4254
rect 4117 4234 4168 4242
rect 4215 4234 4479 4242
rect 4505 4242 4524 4245
rect 4531 4242 4558 4254
rect 4505 4234 4558 4242
rect 4133 4226 4134 4234
rect 4149 4226 4162 4234
rect 4133 4218 4149 4226
rect 4130 4211 4149 4214
rect 4130 4202 4152 4211
rect 4103 4192 4152 4202
rect 4103 4186 4133 4192
rect 4152 4187 4157 4192
rect 4075 4170 4149 4186
rect 4167 4178 4197 4234
rect 4232 4224 4440 4234
rect 4475 4230 4520 4234
rect 4523 4233 4524 4234
rect 4539 4233 4552 4234
rect 4258 4194 4447 4224
rect 4273 4191 4447 4194
rect 4266 4188 4447 4191
rect 4075 4168 4088 4170
rect 4103 4168 4137 4170
rect 4075 4152 4149 4168
rect 4176 4164 4189 4178
rect 4204 4164 4220 4180
rect 4266 4175 4277 4188
rect 4059 4130 4060 4146
rect 4075 4130 4088 4152
rect 4103 4130 4133 4152
rect 4176 4148 4238 4164
rect 4266 4157 4277 4173
rect 4282 4168 4292 4188
rect 4302 4168 4316 4188
rect 4319 4175 4328 4188
rect 4344 4175 4353 4188
rect 4282 4157 4316 4168
rect 4319 4157 4328 4173
rect 4344 4157 4353 4173
rect 4360 4168 4370 4188
rect 4380 4168 4394 4188
rect 4395 4175 4406 4188
rect 4360 4157 4394 4168
rect 4395 4157 4406 4173
rect 4452 4164 4468 4180
rect 4475 4178 4505 4230
rect 4539 4226 4540 4233
rect 4524 4218 4540 4226
rect 4511 4186 4524 4205
rect 4539 4186 4569 4202
rect 4511 4170 4585 4186
rect 4511 4168 4524 4170
rect 4539 4168 4573 4170
rect 4176 4146 4189 4148
rect 4204 4146 4238 4148
rect 4176 4130 4238 4146
rect 4282 4141 4298 4144
rect 4360 4141 4390 4152
rect 4438 4148 4484 4164
rect 4511 4152 4585 4168
rect 4438 4146 4472 4148
rect 4437 4130 4484 4146
rect 4511 4130 4524 4152
rect 4539 4130 4569 4152
rect 4596 4130 4597 4146
rect 4612 4130 4625 4290
rect -7 4122 34 4130
rect -7 4096 8 4122
rect 15 4096 34 4122
rect 98 4118 160 4130
rect 172 4118 247 4130
rect 305 4118 380 4130
rect 392 4118 423 4130
rect 429 4118 464 4130
rect 98 4116 260 4118
rect -7 4088 34 4096
rect 116 4092 129 4116
rect 144 4114 159 4116
rect -1 4078 0 4088
rect 15 4078 28 4088
rect 43 4078 73 4092
rect 116 4078 159 4092
rect 183 4089 190 4096
rect 193 4092 260 4116
rect 292 4116 464 4118
rect 262 4094 290 4098
rect 292 4094 372 4116
rect 393 4114 408 4116
rect 262 4092 372 4094
rect 193 4088 372 4092
rect 166 4078 196 4088
rect 198 4078 351 4088
rect 359 4078 389 4088
rect 393 4078 423 4092
rect 451 4078 464 4116
rect 536 4122 571 4130
rect 536 4096 537 4122
rect 544 4096 571 4122
rect 479 4078 509 4092
rect 536 4088 571 4096
rect 573 4122 614 4130
rect 573 4096 588 4122
rect 595 4096 614 4122
rect 678 4118 740 4130
rect 752 4118 827 4130
rect 885 4118 960 4130
rect 972 4118 1003 4130
rect 1009 4118 1044 4130
rect 678 4116 840 4118
rect 573 4088 614 4096
rect 696 4092 709 4116
rect 724 4114 739 4116
rect 536 4078 537 4088
rect 552 4078 565 4088
rect 579 4078 580 4088
rect 595 4078 608 4088
rect 623 4078 653 4092
rect 696 4078 739 4092
rect 763 4089 770 4096
rect 773 4092 840 4116
rect 872 4116 1044 4118
rect 842 4094 870 4098
rect 872 4094 952 4116
rect 973 4114 988 4116
rect 842 4092 952 4094
rect 773 4088 952 4092
rect 746 4078 776 4088
rect 778 4078 931 4088
rect 939 4078 969 4088
rect 973 4078 1003 4092
rect 1031 4078 1044 4116
rect 1116 4122 1151 4130
rect 1116 4096 1117 4122
rect 1124 4096 1151 4122
rect 1059 4078 1089 4092
rect 1116 4088 1151 4096
rect 1153 4122 1194 4130
rect 1153 4096 1168 4122
rect 1175 4096 1194 4122
rect 1258 4118 1320 4130
rect 1332 4118 1407 4130
rect 1465 4118 1540 4130
rect 1552 4118 1583 4130
rect 1589 4118 1624 4130
rect 1258 4116 1420 4118
rect 1153 4088 1194 4096
rect 1276 4092 1289 4116
rect 1304 4114 1319 4116
rect 1116 4078 1117 4088
rect 1132 4078 1145 4088
rect 1159 4078 1160 4088
rect 1175 4078 1188 4088
rect 1203 4078 1233 4092
rect 1276 4078 1319 4092
rect 1343 4089 1350 4096
rect 1353 4092 1420 4116
rect 1452 4116 1624 4118
rect 1422 4094 1450 4098
rect 1452 4094 1532 4116
rect 1553 4114 1568 4116
rect 1422 4092 1532 4094
rect 1353 4088 1532 4092
rect 1326 4078 1356 4088
rect 1358 4078 1511 4088
rect 1519 4078 1549 4088
rect 1553 4078 1583 4092
rect 1611 4078 1624 4116
rect 1696 4122 1731 4130
rect 1696 4096 1697 4122
rect 1704 4096 1731 4122
rect 1639 4078 1669 4092
rect 1696 4088 1731 4096
rect 1733 4122 1774 4130
rect 1733 4096 1748 4122
rect 1755 4096 1774 4122
rect 1838 4118 1900 4130
rect 1912 4118 1987 4130
rect 2045 4118 2120 4130
rect 2132 4118 2163 4130
rect 2169 4118 2204 4130
rect 1838 4116 2000 4118
rect 1733 4088 1774 4096
rect 1856 4092 1869 4116
rect 1884 4114 1899 4116
rect 1696 4078 1697 4088
rect 1712 4078 1725 4088
rect 1739 4078 1740 4088
rect 1755 4078 1768 4088
rect 1783 4078 1813 4092
rect 1856 4078 1899 4092
rect 1923 4089 1930 4096
rect 1933 4092 2000 4116
rect 2032 4116 2204 4118
rect 2002 4094 2030 4098
rect 2032 4094 2112 4116
rect 2133 4114 2148 4116
rect 2002 4092 2112 4094
rect 1933 4088 2112 4092
rect 1906 4078 1936 4088
rect 1938 4078 2091 4088
rect 2099 4078 2129 4088
rect 2133 4078 2163 4092
rect 2191 4078 2204 4116
rect 2276 4122 2311 4130
rect 2276 4096 2277 4122
rect 2284 4096 2311 4122
rect 2219 4078 2249 4092
rect 2276 4088 2311 4096
rect 2313 4122 2354 4130
rect 2313 4096 2328 4122
rect 2335 4096 2354 4122
rect 2418 4118 2480 4130
rect 2492 4118 2567 4130
rect 2625 4118 2700 4130
rect 2712 4118 2743 4130
rect 2749 4118 2784 4130
rect 2418 4116 2580 4118
rect 2313 4088 2354 4096
rect 2436 4092 2449 4116
rect 2464 4114 2479 4116
rect 2276 4078 2277 4088
rect 2292 4078 2305 4088
rect 2319 4078 2320 4088
rect 2335 4078 2348 4088
rect 2363 4078 2393 4092
rect 2436 4078 2479 4092
rect 2503 4089 2510 4096
rect 2513 4092 2580 4116
rect 2612 4116 2784 4118
rect 2582 4094 2610 4098
rect 2612 4094 2692 4116
rect 2713 4114 2728 4116
rect 2582 4092 2692 4094
rect 2513 4088 2692 4092
rect 2486 4078 2516 4088
rect 2518 4078 2671 4088
rect 2679 4078 2709 4088
rect 2713 4078 2743 4092
rect 2771 4078 2784 4116
rect 2856 4122 2891 4130
rect 2856 4096 2857 4122
rect 2864 4096 2891 4122
rect 2799 4078 2829 4092
rect 2856 4088 2891 4096
rect 2893 4122 2934 4130
rect 2893 4096 2908 4122
rect 2915 4096 2934 4122
rect 2998 4118 3060 4130
rect 3072 4118 3147 4130
rect 3205 4118 3280 4130
rect 3292 4118 3323 4130
rect 3329 4118 3364 4130
rect 2998 4116 3160 4118
rect 2893 4088 2934 4096
rect 3016 4092 3029 4116
rect 3044 4114 3059 4116
rect 2856 4078 2857 4088
rect 2872 4078 2885 4088
rect 2899 4078 2900 4088
rect 2915 4078 2928 4088
rect 2943 4078 2973 4092
rect 3016 4078 3059 4092
rect 3083 4089 3090 4096
rect 3093 4092 3160 4116
rect 3192 4116 3364 4118
rect 3162 4094 3190 4098
rect 3192 4094 3272 4116
rect 3293 4114 3308 4116
rect 3162 4092 3272 4094
rect 3093 4088 3272 4092
rect 3066 4078 3096 4088
rect 3098 4078 3251 4088
rect 3259 4078 3289 4088
rect 3293 4078 3323 4092
rect 3351 4078 3364 4116
rect 3436 4122 3471 4130
rect 3436 4096 3437 4122
rect 3444 4096 3471 4122
rect 3379 4078 3409 4092
rect 3436 4088 3471 4096
rect 3473 4122 3514 4130
rect 3473 4096 3488 4122
rect 3495 4096 3514 4122
rect 3578 4118 3640 4130
rect 3652 4118 3727 4130
rect 3785 4118 3860 4130
rect 3872 4118 3903 4130
rect 3909 4118 3944 4130
rect 3578 4116 3740 4118
rect 3473 4088 3514 4096
rect 3596 4092 3609 4116
rect 3624 4114 3639 4116
rect 3436 4078 3437 4088
rect 3452 4078 3465 4088
rect 3479 4078 3480 4088
rect 3495 4078 3508 4088
rect 3523 4078 3553 4092
rect 3596 4078 3639 4092
rect 3663 4089 3670 4096
rect 3673 4092 3740 4116
rect 3772 4116 3944 4118
rect 3742 4094 3770 4098
rect 3772 4094 3852 4116
rect 3873 4114 3888 4116
rect 3742 4092 3852 4094
rect 3673 4088 3852 4092
rect 3646 4078 3676 4088
rect 3678 4078 3831 4088
rect 3839 4078 3869 4088
rect 3873 4078 3903 4092
rect 3931 4078 3944 4116
rect 4016 4122 4051 4130
rect 4016 4096 4017 4122
rect 4024 4096 4051 4122
rect 3959 4078 3989 4092
rect 4016 4088 4051 4096
rect 4053 4122 4094 4130
rect 4053 4096 4068 4122
rect 4075 4096 4094 4122
rect 4158 4118 4220 4130
rect 4232 4118 4307 4130
rect 4365 4118 4440 4130
rect 4452 4118 4483 4130
rect 4489 4118 4524 4130
rect 4158 4116 4320 4118
rect 4053 4088 4094 4096
rect 4176 4092 4189 4116
rect 4204 4114 4219 4116
rect 4016 4078 4017 4088
rect 4032 4078 4045 4088
rect 4059 4078 4060 4088
rect 4075 4078 4088 4088
rect 4103 4078 4133 4092
rect 4176 4078 4219 4092
rect 4243 4089 4250 4096
rect 4253 4092 4320 4116
rect 4352 4116 4524 4118
rect 4322 4094 4350 4098
rect 4352 4094 4432 4116
rect 4453 4114 4468 4116
rect 4322 4092 4432 4094
rect 4253 4088 4432 4092
rect 4226 4078 4256 4088
rect 4258 4078 4411 4088
rect 4419 4078 4449 4088
rect 4453 4078 4483 4092
rect 4511 4078 4524 4116
rect 4596 4122 4631 4130
rect 4596 4096 4597 4122
rect 4604 4096 4631 4122
rect 4539 4078 4569 4092
rect 4596 4088 4631 4096
rect 4596 4078 4597 4088
rect 4612 4078 4625 4088
rect -1 4072 4625 4078
rect 0 4064 4625 4072
rect 15 4034 28 4064
rect 43 4046 73 4064
rect 116 4050 130 4064
rect 166 4050 386 4064
rect 117 4048 130 4050
rect 83 4036 98 4048
rect 80 4034 102 4036
rect 107 4034 137 4048
rect 198 4046 351 4050
rect 180 4034 372 4046
rect 415 4034 445 4048
rect 451 4034 464 4064
rect 479 4046 509 4064
rect 552 4034 565 4064
rect 595 4034 608 4064
rect 623 4046 653 4064
rect 696 4050 710 4064
rect 746 4050 966 4064
rect 697 4048 710 4050
rect 663 4036 678 4048
rect 660 4034 682 4036
rect 687 4034 717 4048
rect 778 4046 931 4050
rect 760 4034 952 4046
rect 995 4034 1025 4048
rect 1031 4034 1044 4064
rect 1059 4046 1089 4064
rect 1132 4034 1145 4064
rect 1175 4034 1188 4064
rect 1203 4046 1233 4064
rect 1276 4050 1290 4064
rect 1326 4050 1546 4064
rect 1277 4048 1290 4050
rect 1243 4036 1258 4048
rect 1240 4034 1262 4036
rect 1267 4034 1297 4048
rect 1358 4046 1511 4050
rect 1340 4034 1532 4046
rect 1575 4034 1605 4048
rect 1611 4034 1624 4064
rect 1639 4046 1669 4064
rect 1712 4034 1725 4064
rect 1755 4034 1768 4064
rect 1783 4046 1813 4064
rect 1856 4050 1870 4064
rect 1906 4050 2126 4064
rect 1857 4048 1870 4050
rect 1823 4036 1838 4048
rect 1820 4034 1842 4036
rect 1847 4034 1877 4048
rect 1938 4046 2091 4050
rect 1920 4034 2112 4046
rect 2155 4034 2185 4048
rect 2191 4034 2204 4064
rect 2219 4046 2249 4064
rect 2292 4034 2305 4064
rect 2335 4034 2348 4064
rect 2363 4046 2393 4064
rect 2436 4050 2450 4064
rect 2486 4050 2706 4064
rect 2437 4048 2450 4050
rect 2403 4036 2418 4048
rect 2400 4034 2422 4036
rect 2427 4034 2457 4048
rect 2518 4046 2671 4050
rect 2500 4034 2692 4046
rect 2735 4034 2765 4048
rect 2771 4034 2784 4064
rect 2799 4046 2829 4064
rect 2872 4034 2885 4064
rect 2915 4034 2928 4064
rect 2943 4046 2973 4064
rect 3016 4050 3030 4064
rect 3066 4050 3286 4064
rect 3017 4048 3030 4050
rect 2983 4036 2998 4048
rect 2980 4034 3002 4036
rect 3007 4034 3037 4048
rect 3098 4046 3251 4050
rect 3080 4034 3272 4046
rect 3315 4034 3345 4048
rect 3351 4034 3364 4064
rect 3379 4046 3409 4064
rect 3452 4034 3465 4064
rect 3495 4034 3508 4064
rect 3523 4046 3553 4064
rect 3596 4050 3610 4064
rect 3646 4050 3866 4064
rect 3597 4048 3610 4050
rect 3563 4036 3578 4048
rect 3560 4034 3582 4036
rect 3587 4034 3617 4048
rect 3678 4046 3831 4050
rect 3660 4034 3852 4046
rect 3895 4034 3925 4048
rect 3931 4034 3944 4064
rect 3959 4046 3989 4064
rect 4032 4034 4045 4064
rect 4075 4034 4088 4064
rect 4103 4046 4133 4064
rect 4176 4050 4190 4064
rect 4226 4050 4446 4064
rect 4177 4048 4190 4050
rect 4143 4036 4158 4048
rect 4140 4034 4162 4036
rect 4167 4034 4197 4048
rect 4258 4046 4411 4050
rect 4240 4034 4432 4046
rect 4475 4034 4505 4048
rect 4511 4034 4524 4064
rect 4539 4046 4569 4064
rect 4612 4034 4625 4064
rect 0 4020 4625 4034
rect 15 3916 28 4020
rect 73 3998 74 4008
rect 89 3998 102 4008
rect 73 3994 102 3998
rect 107 3994 137 4020
rect 155 4006 171 4008
rect 243 4006 296 4020
rect 244 4004 308 4006
rect 351 4004 366 4020
rect 415 4017 445 4020
rect 415 4014 451 4017
rect 381 4006 397 4008
rect 155 3994 170 3998
rect 73 3992 170 3994
rect 198 3992 366 4004
rect 382 3994 397 3998
rect 415 3995 454 4014
rect 473 4008 480 4009
rect 479 4001 480 4008
rect 463 3998 464 4001
rect 479 3998 492 4001
rect 415 3994 445 3995
rect 454 3994 460 3995
rect 463 3994 492 3998
rect 382 3993 492 3994
rect 382 3992 498 3993
rect 57 3984 108 3992
rect 57 3972 82 3984
rect 89 3972 108 3984
rect 139 3984 189 3992
rect 139 3976 155 3984
rect 162 3982 189 3984
rect 198 3982 419 3992
rect 162 3972 419 3982
rect 448 3984 498 3992
rect 448 3975 464 3984
rect 57 3964 108 3972
rect 155 3964 419 3972
rect 445 3972 464 3975
rect 471 3972 498 3984
rect 445 3964 498 3972
rect 73 3956 74 3964
rect 89 3956 102 3964
rect 73 3948 89 3956
rect 70 3941 89 3944
rect 70 3932 92 3941
rect 43 3922 92 3932
rect 43 3916 73 3922
rect 92 3917 97 3922
rect 15 3900 89 3916
rect 107 3908 137 3964
rect 172 3954 380 3964
rect 415 3960 460 3964
rect 463 3963 464 3964
rect 479 3963 492 3964
rect 198 3924 387 3954
rect 213 3921 387 3924
rect 206 3918 387 3921
rect 15 3898 28 3900
rect 43 3898 77 3900
rect 15 3882 89 3898
rect 116 3894 129 3908
rect 144 3894 160 3910
rect 206 3905 217 3918
rect -1 3860 0 3876
rect 15 3860 28 3882
rect 43 3860 73 3882
rect 116 3878 178 3894
rect 206 3887 217 3903
rect 222 3898 232 3918
rect 242 3898 256 3918
rect 259 3905 268 3918
rect 284 3905 293 3918
rect 222 3887 256 3898
rect 259 3887 268 3903
rect 284 3887 293 3903
rect 300 3898 310 3918
rect 320 3898 334 3918
rect 335 3905 346 3918
rect 300 3887 334 3898
rect 335 3887 346 3903
rect 392 3894 408 3910
rect 415 3908 445 3960
rect 479 3956 480 3963
rect 464 3948 480 3956
rect 451 3916 464 3935
rect 479 3916 509 3932
rect 451 3900 525 3916
rect 451 3898 464 3900
rect 479 3898 513 3900
rect 116 3876 129 3878
rect 144 3876 178 3878
rect 116 3860 178 3876
rect 222 3871 238 3874
rect 300 3871 330 3882
rect 378 3878 424 3894
rect 451 3882 525 3898
rect 378 3876 412 3878
rect 377 3860 424 3876
rect 451 3860 464 3882
rect 479 3860 509 3882
rect 536 3860 537 3876
rect 552 3860 565 4020
rect 595 3916 608 4020
rect 653 3998 654 4008
rect 669 3998 682 4008
rect 653 3994 682 3998
rect 687 3994 717 4020
rect 735 4006 751 4008
rect 823 4006 876 4020
rect 824 4004 888 4006
rect 931 4004 946 4020
rect 995 4017 1025 4020
rect 995 4014 1031 4017
rect 961 4006 977 4008
rect 735 3994 750 3998
rect 653 3992 750 3994
rect 778 3992 946 4004
rect 962 3994 977 3998
rect 995 3995 1034 4014
rect 1053 4008 1060 4009
rect 1059 4001 1060 4008
rect 1043 3998 1044 4001
rect 1059 3998 1072 4001
rect 995 3994 1025 3995
rect 1034 3994 1040 3995
rect 1043 3994 1072 3998
rect 962 3993 1072 3994
rect 962 3992 1078 3993
rect 637 3984 688 3992
rect 637 3972 662 3984
rect 669 3972 688 3984
rect 719 3984 769 3992
rect 719 3976 735 3984
rect 742 3982 769 3984
rect 778 3982 999 3992
rect 742 3972 999 3982
rect 1028 3984 1078 3992
rect 1028 3975 1044 3984
rect 637 3964 688 3972
rect 735 3964 999 3972
rect 1025 3972 1044 3975
rect 1051 3972 1078 3984
rect 1025 3964 1078 3972
rect 653 3956 654 3964
rect 669 3956 682 3964
rect 653 3948 669 3956
rect 650 3941 669 3944
rect 650 3932 672 3941
rect 623 3922 672 3932
rect 623 3916 653 3922
rect 672 3917 677 3922
rect 595 3900 669 3916
rect 687 3908 717 3964
rect 752 3954 960 3964
rect 995 3960 1040 3964
rect 1043 3963 1044 3964
rect 1059 3963 1072 3964
rect 778 3924 967 3954
rect 793 3921 967 3924
rect 786 3918 967 3921
rect 595 3898 608 3900
rect 623 3898 657 3900
rect 595 3882 669 3898
rect 696 3894 709 3908
rect 724 3894 740 3910
rect 786 3905 797 3918
rect 579 3860 580 3876
rect 595 3860 608 3882
rect 623 3860 653 3882
rect 696 3878 758 3894
rect 786 3887 797 3903
rect 802 3898 812 3918
rect 822 3898 836 3918
rect 839 3905 848 3918
rect 864 3905 873 3918
rect 802 3887 836 3898
rect 839 3887 848 3903
rect 864 3887 873 3903
rect 880 3898 890 3918
rect 900 3898 914 3918
rect 915 3905 926 3918
rect 880 3887 914 3898
rect 915 3887 926 3903
rect 972 3894 988 3910
rect 995 3908 1025 3960
rect 1059 3956 1060 3963
rect 1044 3948 1060 3956
rect 1031 3916 1044 3935
rect 1059 3916 1089 3932
rect 1031 3900 1105 3916
rect 1031 3898 1044 3900
rect 1059 3898 1093 3900
rect 696 3876 709 3878
rect 724 3876 758 3878
rect 696 3860 758 3876
rect 802 3871 818 3874
rect 880 3871 910 3882
rect 958 3878 1004 3894
rect 1031 3882 1105 3898
rect 958 3876 992 3878
rect 957 3860 1004 3876
rect 1031 3860 1044 3882
rect 1059 3860 1089 3882
rect 1116 3860 1117 3876
rect 1132 3860 1145 4020
rect 1175 3916 1188 4020
rect 1233 3998 1234 4008
rect 1249 3998 1262 4008
rect 1233 3994 1262 3998
rect 1267 3994 1297 4020
rect 1315 4006 1331 4008
rect 1403 4006 1456 4020
rect 1404 4004 1468 4006
rect 1511 4004 1526 4020
rect 1575 4017 1605 4020
rect 1575 4014 1611 4017
rect 1541 4006 1557 4008
rect 1315 3994 1330 3998
rect 1233 3992 1330 3994
rect 1358 3992 1526 4004
rect 1542 3994 1557 3998
rect 1575 3995 1614 4014
rect 1633 4008 1640 4009
rect 1639 4001 1640 4008
rect 1623 3998 1624 4001
rect 1639 3998 1652 4001
rect 1575 3994 1605 3995
rect 1614 3994 1620 3995
rect 1623 3994 1652 3998
rect 1542 3993 1652 3994
rect 1542 3992 1658 3993
rect 1217 3984 1268 3992
rect 1217 3972 1242 3984
rect 1249 3972 1268 3984
rect 1299 3984 1349 3992
rect 1299 3976 1315 3984
rect 1322 3982 1349 3984
rect 1358 3982 1579 3992
rect 1322 3972 1579 3982
rect 1608 3984 1658 3992
rect 1608 3975 1624 3984
rect 1217 3964 1268 3972
rect 1315 3964 1579 3972
rect 1605 3972 1624 3975
rect 1631 3972 1658 3984
rect 1605 3964 1658 3972
rect 1233 3956 1234 3964
rect 1249 3956 1262 3964
rect 1233 3948 1249 3956
rect 1230 3941 1249 3944
rect 1230 3932 1252 3941
rect 1203 3922 1252 3932
rect 1203 3916 1233 3922
rect 1252 3917 1257 3922
rect 1175 3900 1249 3916
rect 1267 3908 1297 3964
rect 1332 3954 1540 3964
rect 1575 3960 1620 3964
rect 1623 3963 1624 3964
rect 1639 3963 1652 3964
rect 1358 3924 1547 3954
rect 1373 3921 1547 3924
rect 1366 3918 1547 3921
rect 1175 3898 1188 3900
rect 1203 3898 1237 3900
rect 1175 3882 1249 3898
rect 1276 3894 1289 3908
rect 1304 3894 1320 3910
rect 1366 3905 1377 3918
rect 1159 3860 1160 3876
rect 1175 3860 1188 3882
rect 1203 3860 1233 3882
rect 1276 3878 1338 3894
rect 1366 3887 1377 3903
rect 1382 3898 1392 3918
rect 1402 3898 1416 3918
rect 1419 3905 1428 3918
rect 1444 3905 1453 3918
rect 1382 3887 1416 3898
rect 1419 3887 1428 3903
rect 1444 3887 1453 3903
rect 1460 3898 1470 3918
rect 1480 3898 1494 3918
rect 1495 3905 1506 3918
rect 1460 3887 1494 3898
rect 1495 3887 1506 3903
rect 1552 3894 1568 3910
rect 1575 3908 1605 3960
rect 1639 3956 1640 3963
rect 1624 3948 1640 3956
rect 1611 3916 1624 3935
rect 1639 3916 1669 3932
rect 1611 3900 1685 3916
rect 1611 3898 1624 3900
rect 1639 3898 1673 3900
rect 1276 3876 1289 3878
rect 1304 3876 1338 3878
rect 1276 3860 1338 3876
rect 1382 3871 1398 3874
rect 1460 3871 1490 3882
rect 1538 3878 1584 3894
rect 1611 3882 1685 3898
rect 1538 3876 1572 3878
rect 1537 3860 1584 3876
rect 1611 3860 1624 3882
rect 1639 3860 1669 3882
rect 1696 3860 1697 3876
rect 1712 3860 1725 4020
rect 1755 3916 1768 4020
rect 1813 3998 1814 4008
rect 1829 3998 1842 4008
rect 1813 3994 1842 3998
rect 1847 3994 1877 4020
rect 1895 4006 1911 4008
rect 1983 4006 2036 4020
rect 1984 4004 2048 4006
rect 2091 4004 2106 4020
rect 2155 4017 2185 4020
rect 2155 4014 2191 4017
rect 2121 4006 2137 4008
rect 1895 3994 1910 3998
rect 1813 3992 1910 3994
rect 1938 3992 2106 4004
rect 2122 3994 2137 3998
rect 2155 3995 2194 4014
rect 2213 4008 2220 4009
rect 2219 4001 2220 4008
rect 2203 3998 2204 4001
rect 2219 3998 2232 4001
rect 2155 3994 2185 3995
rect 2194 3994 2200 3995
rect 2203 3994 2232 3998
rect 2122 3993 2232 3994
rect 2122 3992 2238 3993
rect 1797 3984 1848 3992
rect 1797 3972 1822 3984
rect 1829 3972 1848 3984
rect 1879 3984 1929 3992
rect 1879 3976 1895 3984
rect 1902 3982 1929 3984
rect 1938 3982 2159 3992
rect 1902 3972 2159 3982
rect 2188 3984 2238 3992
rect 2188 3975 2204 3984
rect 1797 3964 1848 3972
rect 1895 3964 2159 3972
rect 2185 3972 2204 3975
rect 2211 3972 2238 3984
rect 2185 3964 2238 3972
rect 1813 3956 1814 3964
rect 1829 3956 1842 3964
rect 1813 3948 1829 3956
rect 1810 3941 1829 3944
rect 1810 3932 1832 3941
rect 1783 3922 1832 3932
rect 1783 3916 1813 3922
rect 1832 3917 1837 3922
rect 1755 3900 1829 3916
rect 1847 3908 1877 3964
rect 1912 3954 2120 3964
rect 2155 3960 2200 3964
rect 2203 3963 2204 3964
rect 2219 3963 2232 3964
rect 1938 3924 2127 3954
rect 1953 3921 2127 3924
rect 1946 3918 2127 3921
rect 1755 3898 1768 3900
rect 1783 3898 1817 3900
rect 1755 3882 1829 3898
rect 1856 3894 1869 3908
rect 1884 3894 1900 3910
rect 1946 3905 1957 3918
rect 1739 3860 1740 3876
rect 1755 3860 1768 3882
rect 1783 3860 1813 3882
rect 1856 3878 1918 3894
rect 1946 3887 1957 3903
rect 1962 3898 1972 3918
rect 1982 3898 1996 3918
rect 1999 3905 2008 3918
rect 2024 3905 2033 3918
rect 1962 3887 1996 3898
rect 1999 3887 2008 3903
rect 2024 3887 2033 3903
rect 2040 3898 2050 3918
rect 2060 3898 2074 3918
rect 2075 3905 2086 3918
rect 2040 3887 2074 3898
rect 2075 3887 2086 3903
rect 2132 3894 2148 3910
rect 2155 3908 2185 3960
rect 2219 3956 2220 3963
rect 2204 3948 2220 3956
rect 2191 3916 2204 3935
rect 2219 3916 2249 3932
rect 2191 3900 2265 3916
rect 2191 3898 2204 3900
rect 2219 3898 2253 3900
rect 1856 3876 1869 3878
rect 1884 3876 1918 3878
rect 1856 3860 1918 3876
rect 1962 3871 1978 3874
rect 2040 3871 2070 3882
rect 2118 3878 2164 3894
rect 2191 3882 2265 3898
rect 2118 3876 2152 3878
rect 2117 3860 2164 3876
rect 2191 3860 2204 3882
rect 2219 3860 2249 3882
rect 2276 3860 2277 3876
rect 2292 3860 2305 4020
rect 2335 3916 2348 4020
rect 2393 3998 2394 4008
rect 2409 3998 2422 4008
rect 2393 3994 2422 3998
rect 2427 3994 2457 4020
rect 2475 4006 2491 4008
rect 2563 4006 2616 4020
rect 2564 4004 2628 4006
rect 2671 4004 2686 4020
rect 2735 4017 2765 4020
rect 2735 4014 2771 4017
rect 2701 4006 2717 4008
rect 2475 3994 2490 3998
rect 2393 3992 2490 3994
rect 2518 3992 2686 4004
rect 2702 3994 2717 3998
rect 2735 3995 2774 4014
rect 2793 4008 2800 4009
rect 2799 4001 2800 4008
rect 2783 3998 2784 4001
rect 2799 3998 2812 4001
rect 2735 3994 2765 3995
rect 2774 3994 2780 3995
rect 2783 3994 2812 3998
rect 2702 3993 2812 3994
rect 2702 3992 2818 3993
rect 2377 3984 2428 3992
rect 2377 3972 2402 3984
rect 2409 3972 2428 3984
rect 2459 3984 2509 3992
rect 2459 3976 2475 3984
rect 2482 3982 2509 3984
rect 2518 3982 2739 3992
rect 2482 3972 2739 3982
rect 2768 3984 2818 3992
rect 2768 3975 2784 3984
rect 2377 3964 2428 3972
rect 2475 3964 2739 3972
rect 2765 3972 2784 3975
rect 2791 3972 2818 3984
rect 2765 3964 2818 3972
rect 2393 3956 2394 3964
rect 2409 3956 2422 3964
rect 2393 3948 2409 3956
rect 2390 3941 2409 3944
rect 2390 3932 2412 3941
rect 2363 3922 2412 3932
rect 2363 3916 2393 3922
rect 2412 3917 2417 3922
rect 2335 3900 2409 3916
rect 2427 3908 2457 3964
rect 2492 3954 2700 3964
rect 2735 3960 2780 3964
rect 2783 3963 2784 3964
rect 2799 3963 2812 3964
rect 2518 3924 2707 3954
rect 2533 3921 2707 3924
rect 2526 3918 2707 3921
rect 2335 3898 2348 3900
rect 2363 3898 2397 3900
rect 2335 3882 2409 3898
rect 2436 3894 2449 3908
rect 2464 3894 2480 3910
rect 2526 3905 2537 3918
rect 2319 3860 2320 3876
rect 2335 3860 2348 3882
rect 2363 3860 2393 3882
rect 2436 3878 2498 3894
rect 2526 3887 2537 3903
rect 2542 3898 2552 3918
rect 2562 3898 2576 3918
rect 2579 3905 2588 3918
rect 2604 3905 2613 3918
rect 2542 3887 2576 3898
rect 2579 3887 2588 3903
rect 2604 3887 2613 3903
rect 2620 3898 2630 3918
rect 2640 3898 2654 3918
rect 2655 3905 2666 3918
rect 2620 3887 2654 3898
rect 2655 3887 2666 3903
rect 2712 3894 2728 3910
rect 2735 3908 2765 3960
rect 2799 3956 2800 3963
rect 2784 3948 2800 3956
rect 2771 3916 2784 3935
rect 2799 3916 2829 3932
rect 2771 3900 2845 3916
rect 2771 3898 2784 3900
rect 2799 3898 2833 3900
rect 2436 3876 2449 3878
rect 2464 3876 2498 3878
rect 2436 3860 2498 3876
rect 2542 3871 2558 3874
rect 2620 3871 2650 3882
rect 2698 3878 2744 3894
rect 2771 3882 2845 3898
rect 2698 3876 2732 3878
rect 2697 3860 2744 3876
rect 2771 3860 2784 3882
rect 2799 3860 2829 3882
rect 2856 3860 2857 3876
rect 2872 3860 2885 4020
rect 2915 3916 2928 4020
rect 2973 3998 2974 4008
rect 2989 3998 3002 4008
rect 2973 3994 3002 3998
rect 3007 3994 3037 4020
rect 3055 4006 3071 4008
rect 3143 4006 3196 4020
rect 3144 4004 3208 4006
rect 3251 4004 3266 4020
rect 3315 4017 3345 4020
rect 3315 4014 3351 4017
rect 3281 4006 3297 4008
rect 3055 3994 3070 3998
rect 2973 3992 3070 3994
rect 3098 3992 3266 4004
rect 3282 3994 3297 3998
rect 3315 3995 3354 4014
rect 3373 4008 3380 4009
rect 3379 4001 3380 4008
rect 3363 3998 3364 4001
rect 3379 3998 3392 4001
rect 3315 3994 3345 3995
rect 3354 3994 3360 3995
rect 3363 3994 3392 3998
rect 3282 3993 3392 3994
rect 3282 3992 3398 3993
rect 2957 3984 3008 3992
rect 2957 3972 2982 3984
rect 2989 3972 3008 3984
rect 3039 3984 3089 3992
rect 3039 3976 3055 3984
rect 3062 3982 3089 3984
rect 3098 3982 3319 3992
rect 3062 3972 3319 3982
rect 3348 3984 3398 3992
rect 3348 3975 3364 3984
rect 2957 3964 3008 3972
rect 3055 3964 3319 3972
rect 3345 3972 3364 3975
rect 3371 3972 3398 3984
rect 3345 3964 3398 3972
rect 2973 3956 2974 3964
rect 2989 3956 3002 3964
rect 2973 3948 2989 3956
rect 2970 3941 2989 3944
rect 2970 3932 2992 3941
rect 2943 3922 2992 3932
rect 2943 3916 2973 3922
rect 2992 3917 2997 3922
rect 2915 3900 2989 3916
rect 3007 3908 3037 3964
rect 3072 3954 3280 3964
rect 3315 3960 3360 3964
rect 3363 3963 3364 3964
rect 3379 3963 3392 3964
rect 3098 3924 3287 3954
rect 3113 3921 3287 3924
rect 3106 3918 3287 3921
rect 2915 3898 2928 3900
rect 2943 3898 2977 3900
rect 2915 3882 2989 3898
rect 3016 3894 3029 3908
rect 3044 3894 3060 3910
rect 3106 3905 3117 3918
rect 2899 3860 2900 3876
rect 2915 3860 2928 3882
rect 2943 3860 2973 3882
rect 3016 3878 3078 3894
rect 3106 3887 3117 3903
rect 3122 3898 3132 3918
rect 3142 3898 3156 3918
rect 3159 3905 3168 3918
rect 3184 3905 3193 3918
rect 3122 3887 3156 3898
rect 3159 3887 3168 3903
rect 3184 3887 3193 3903
rect 3200 3898 3210 3918
rect 3220 3898 3234 3918
rect 3235 3905 3246 3918
rect 3200 3887 3234 3898
rect 3235 3887 3246 3903
rect 3292 3894 3308 3910
rect 3315 3908 3345 3960
rect 3379 3956 3380 3963
rect 3364 3948 3380 3956
rect 3351 3916 3364 3935
rect 3379 3916 3409 3932
rect 3351 3900 3425 3916
rect 3351 3898 3364 3900
rect 3379 3898 3413 3900
rect 3016 3876 3029 3878
rect 3044 3876 3078 3878
rect 3016 3860 3078 3876
rect 3122 3871 3138 3874
rect 3200 3871 3230 3882
rect 3278 3878 3324 3894
rect 3351 3882 3425 3898
rect 3278 3876 3312 3878
rect 3277 3860 3324 3876
rect 3351 3860 3364 3882
rect 3379 3860 3409 3882
rect 3436 3860 3437 3876
rect 3452 3860 3465 4020
rect 3495 3916 3508 4020
rect 3553 3998 3554 4008
rect 3569 3998 3582 4008
rect 3553 3994 3582 3998
rect 3587 3994 3617 4020
rect 3635 4006 3651 4008
rect 3723 4006 3776 4020
rect 3724 4004 3788 4006
rect 3831 4004 3846 4020
rect 3895 4017 3925 4020
rect 3895 4014 3931 4017
rect 3861 4006 3877 4008
rect 3635 3994 3650 3998
rect 3553 3992 3650 3994
rect 3678 3992 3846 4004
rect 3862 3994 3877 3998
rect 3895 3995 3934 4014
rect 3953 4008 3960 4009
rect 3959 4001 3960 4008
rect 3943 3998 3944 4001
rect 3959 3998 3972 4001
rect 3895 3994 3925 3995
rect 3934 3994 3940 3995
rect 3943 3994 3972 3998
rect 3862 3993 3972 3994
rect 3862 3992 3978 3993
rect 3537 3984 3588 3992
rect 3537 3972 3562 3984
rect 3569 3972 3588 3984
rect 3619 3984 3669 3992
rect 3619 3976 3635 3984
rect 3642 3982 3669 3984
rect 3678 3982 3899 3992
rect 3642 3972 3899 3982
rect 3928 3984 3978 3992
rect 3928 3975 3944 3984
rect 3537 3964 3588 3972
rect 3635 3964 3899 3972
rect 3925 3972 3944 3975
rect 3951 3972 3978 3984
rect 3925 3964 3978 3972
rect 3553 3956 3554 3964
rect 3569 3956 3582 3964
rect 3553 3948 3569 3956
rect 3550 3941 3569 3944
rect 3550 3932 3572 3941
rect 3523 3922 3572 3932
rect 3523 3916 3553 3922
rect 3572 3917 3577 3922
rect 3495 3900 3569 3916
rect 3587 3908 3617 3964
rect 3652 3954 3860 3964
rect 3895 3960 3940 3964
rect 3943 3963 3944 3964
rect 3959 3963 3972 3964
rect 3678 3924 3867 3954
rect 3693 3921 3867 3924
rect 3686 3918 3867 3921
rect 3495 3898 3508 3900
rect 3523 3898 3557 3900
rect 3495 3882 3569 3898
rect 3596 3894 3609 3908
rect 3624 3894 3640 3910
rect 3686 3905 3697 3918
rect 3479 3860 3480 3876
rect 3495 3860 3508 3882
rect 3523 3860 3553 3882
rect 3596 3878 3658 3894
rect 3686 3887 3697 3903
rect 3702 3898 3712 3918
rect 3722 3898 3736 3918
rect 3739 3905 3748 3918
rect 3764 3905 3773 3918
rect 3702 3887 3736 3898
rect 3739 3887 3748 3903
rect 3764 3887 3773 3903
rect 3780 3898 3790 3918
rect 3800 3898 3814 3918
rect 3815 3905 3826 3918
rect 3780 3887 3814 3898
rect 3815 3887 3826 3903
rect 3872 3894 3888 3910
rect 3895 3908 3925 3960
rect 3959 3956 3960 3963
rect 3944 3948 3960 3956
rect 3931 3916 3944 3935
rect 3959 3916 3989 3932
rect 3931 3900 4005 3916
rect 3931 3898 3944 3900
rect 3959 3898 3993 3900
rect 3596 3876 3609 3878
rect 3624 3876 3658 3878
rect 3596 3860 3658 3876
rect 3702 3871 3718 3874
rect 3780 3871 3810 3882
rect 3858 3878 3904 3894
rect 3931 3882 4005 3898
rect 3858 3876 3892 3878
rect 3857 3860 3904 3876
rect 3931 3860 3944 3882
rect 3959 3860 3989 3882
rect 4016 3860 4017 3876
rect 4032 3860 4045 4020
rect 4075 3916 4088 4020
rect 4133 3998 4134 4008
rect 4149 3998 4162 4008
rect 4133 3994 4162 3998
rect 4167 3994 4197 4020
rect 4215 4006 4231 4008
rect 4303 4006 4356 4020
rect 4304 4004 4368 4006
rect 4411 4004 4426 4020
rect 4475 4017 4505 4020
rect 4475 4014 4511 4017
rect 4441 4006 4457 4008
rect 4215 3994 4230 3998
rect 4133 3992 4230 3994
rect 4258 3992 4426 4004
rect 4442 3994 4457 3998
rect 4475 3995 4514 4014
rect 4533 4008 4540 4009
rect 4539 4001 4540 4008
rect 4523 3998 4524 4001
rect 4539 3998 4552 4001
rect 4475 3994 4505 3995
rect 4514 3994 4520 3995
rect 4523 3994 4552 3998
rect 4442 3993 4552 3994
rect 4442 3992 4558 3993
rect 4117 3984 4168 3992
rect 4117 3972 4142 3984
rect 4149 3972 4168 3984
rect 4199 3984 4249 3992
rect 4199 3976 4215 3984
rect 4222 3982 4249 3984
rect 4258 3982 4479 3992
rect 4222 3972 4479 3982
rect 4508 3984 4558 3992
rect 4508 3975 4524 3984
rect 4117 3964 4168 3972
rect 4215 3964 4479 3972
rect 4505 3972 4524 3975
rect 4531 3972 4558 3984
rect 4505 3964 4558 3972
rect 4133 3956 4134 3964
rect 4149 3956 4162 3964
rect 4133 3948 4149 3956
rect 4130 3941 4149 3944
rect 4130 3932 4152 3941
rect 4103 3922 4152 3932
rect 4103 3916 4133 3922
rect 4152 3917 4157 3922
rect 4075 3900 4149 3916
rect 4167 3908 4197 3964
rect 4232 3954 4440 3964
rect 4475 3960 4520 3964
rect 4523 3963 4524 3964
rect 4539 3963 4552 3964
rect 4258 3924 4447 3954
rect 4273 3921 4447 3924
rect 4266 3918 4447 3921
rect 4075 3898 4088 3900
rect 4103 3898 4137 3900
rect 4075 3882 4149 3898
rect 4176 3894 4189 3908
rect 4204 3894 4220 3910
rect 4266 3905 4277 3918
rect 4059 3860 4060 3876
rect 4075 3860 4088 3882
rect 4103 3860 4133 3882
rect 4176 3878 4238 3894
rect 4266 3887 4277 3903
rect 4282 3898 4292 3918
rect 4302 3898 4316 3918
rect 4319 3905 4328 3918
rect 4344 3905 4353 3918
rect 4282 3887 4316 3898
rect 4319 3887 4328 3903
rect 4344 3887 4353 3903
rect 4360 3898 4370 3918
rect 4380 3898 4394 3918
rect 4395 3905 4406 3918
rect 4360 3887 4394 3898
rect 4395 3887 4406 3903
rect 4452 3894 4468 3910
rect 4475 3908 4505 3960
rect 4539 3956 4540 3963
rect 4524 3948 4540 3956
rect 4511 3916 4524 3935
rect 4539 3916 4569 3932
rect 4511 3900 4585 3916
rect 4511 3898 4524 3900
rect 4539 3898 4573 3900
rect 4176 3876 4189 3878
rect 4204 3876 4238 3878
rect 4176 3860 4238 3876
rect 4282 3871 4298 3874
rect 4360 3871 4390 3882
rect 4438 3878 4484 3894
rect 4511 3882 4585 3898
rect 4438 3876 4472 3878
rect 4437 3860 4484 3876
rect 4511 3860 4524 3882
rect 4539 3860 4569 3882
rect 4596 3860 4597 3876
rect 4612 3860 4625 4020
rect -7 3852 34 3860
rect -7 3826 8 3852
rect 15 3826 34 3852
rect 98 3848 160 3860
rect 172 3848 247 3860
rect 305 3848 380 3860
rect 392 3848 423 3860
rect 429 3848 464 3860
rect 98 3846 260 3848
rect -7 3818 34 3826
rect 116 3822 129 3846
rect 144 3844 159 3846
rect -1 3808 0 3818
rect 15 3808 28 3818
rect 43 3808 73 3822
rect 116 3808 159 3822
rect 183 3819 190 3826
rect 193 3822 260 3846
rect 292 3846 464 3848
rect 262 3824 290 3828
rect 292 3824 372 3846
rect 393 3844 408 3846
rect 262 3822 372 3824
rect 193 3818 372 3822
rect 166 3808 196 3818
rect 198 3808 351 3818
rect 359 3808 389 3818
rect 393 3808 423 3822
rect 451 3808 464 3846
rect 536 3852 571 3860
rect 536 3826 537 3852
rect 544 3826 571 3852
rect 479 3808 509 3822
rect 536 3818 571 3826
rect 573 3852 614 3860
rect 573 3826 588 3852
rect 595 3826 614 3852
rect 678 3848 740 3860
rect 752 3848 827 3860
rect 885 3848 960 3860
rect 972 3848 1003 3860
rect 1009 3848 1044 3860
rect 678 3846 840 3848
rect 573 3818 614 3826
rect 696 3822 709 3846
rect 724 3844 739 3846
rect 536 3808 537 3818
rect 552 3808 565 3818
rect 579 3808 580 3818
rect 595 3808 608 3818
rect 623 3808 653 3822
rect 696 3808 739 3822
rect 763 3819 770 3826
rect 773 3822 840 3846
rect 872 3846 1044 3848
rect 842 3824 870 3828
rect 872 3824 952 3846
rect 973 3844 988 3846
rect 842 3822 952 3824
rect 773 3818 952 3822
rect 746 3808 776 3818
rect 778 3808 931 3818
rect 939 3808 969 3818
rect 973 3808 1003 3822
rect 1031 3808 1044 3846
rect 1116 3852 1151 3860
rect 1116 3826 1117 3852
rect 1124 3826 1151 3852
rect 1059 3808 1089 3822
rect 1116 3818 1151 3826
rect 1153 3852 1194 3860
rect 1153 3826 1168 3852
rect 1175 3826 1194 3852
rect 1258 3848 1320 3860
rect 1332 3848 1407 3860
rect 1465 3848 1540 3860
rect 1552 3848 1583 3860
rect 1589 3848 1624 3860
rect 1258 3846 1420 3848
rect 1153 3818 1194 3826
rect 1276 3822 1289 3846
rect 1304 3844 1319 3846
rect 1116 3808 1117 3818
rect 1132 3808 1145 3818
rect 1159 3808 1160 3818
rect 1175 3808 1188 3818
rect 1203 3808 1233 3822
rect 1276 3808 1319 3822
rect 1343 3819 1350 3826
rect 1353 3822 1420 3846
rect 1452 3846 1624 3848
rect 1422 3824 1450 3828
rect 1452 3824 1532 3846
rect 1553 3844 1568 3846
rect 1422 3822 1532 3824
rect 1353 3818 1532 3822
rect 1326 3808 1356 3818
rect 1358 3808 1511 3818
rect 1519 3808 1549 3818
rect 1553 3808 1583 3822
rect 1611 3808 1624 3846
rect 1696 3852 1731 3860
rect 1696 3826 1697 3852
rect 1704 3826 1731 3852
rect 1639 3808 1669 3822
rect 1696 3818 1731 3826
rect 1733 3852 1774 3860
rect 1733 3826 1748 3852
rect 1755 3826 1774 3852
rect 1838 3848 1900 3860
rect 1912 3848 1987 3860
rect 2045 3848 2120 3860
rect 2132 3848 2163 3860
rect 2169 3848 2204 3860
rect 1838 3846 2000 3848
rect 1733 3818 1774 3826
rect 1856 3822 1869 3846
rect 1884 3844 1899 3846
rect 1696 3808 1697 3818
rect 1712 3808 1725 3818
rect 1739 3808 1740 3818
rect 1755 3808 1768 3818
rect 1783 3808 1813 3822
rect 1856 3808 1899 3822
rect 1923 3819 1930 3826
rect 1933 3822 2000 3846
rect 2032 3846 2204 3848
rect 2002 3824 2030 3828
rect 2032 3824 2112 3846
rect 2133 3844 2148 3846
rect 2002 3822 2112 3824
rect 1933 3818 2112 3822
rect 1906 3808 1936 3818
rect 1938 3808 2091 3818
rect 2099 3808 2129 3818
rect 2133 3808 2163 3822
rect 2191 3808 2204 3846
rect 2276 3852 2311 3860
rect 2276 3826 2277 3852
rect 2284 3826 2311 3852
rect 2219 3808 2249 3822
rect 2276 3818 2311 3826
rect 2313 3852 2354 3860
rect 2313 3826 2328 3852
rect 2335 3826 2354 3852
rect 2418 3848 2480 3860
rect 2492 3848 2567 3860
rect 2625 3848 2700 3860
rect 2712 3848 2743 3860
rect 2749 3848 2784 3860
rect 2418 3846 2580 3848
rect 2313 3818 2354 3826
rect 2436 3822 2449 3846
rect 2464 3844 2479 3846
rect 2276 3808 2277 3818
rect 2292 3808 2305 3818
rect 2319 3808 2320 3818
rect 2335 3808 2348 3818
rect 2363 3808 2393 3822
rect 2436 3808 2479 3822
rect 2503 3819 2510 3826
rect 2513 3822 2580 3846
rect 2612 3846 2784 3848
rect 2582 3824 2610 3828
rect 2612 3824 2692 3846
rect 2713 3844 2728 3846
rect 2582 3822 2692 3824
rect 2513 3818 2692 3822
rect 2486 3808 2516 3818
rect 2518 3808 2671 3818
rect 2679 3808 2709 3818
rect 2713 3808 2743 3822
rect 2771 3808 2784 3846
rect 2856 3852 2891 3860
rect 2856 3826 2857 3852
rect 2864 3826 2891 3852
rect 2799 3808 2829 3822
rect 2856 3818 2891 3826
rect 2893 3852 2934 3860
rect 2893 3826 2908 3852
rect 2915 3826 2934 3852
rect 2998 3848 3060 3860
rect 3072 3848 3147 3860
rect 3205 3848 3280 3860
rect 3292 3848 3323 3860
rect 3329 3848 3364 3860
rect 2998 3846 3160 3848
rect 2893 3818 2934 3826
rect 3016 3822 3029 3846
rect 3044 3844 3059 3846
rect 2856 3808 2857 3818
rect 2872 3808 2885 3818
rect 2899 3808 2900 3818
rect 2915 3808 2928 3818
rect 2943 3808 2973 3822
rect 3016 3808 3059 3822
rect 3083 3819 3090 3826
rect 3093 3822 3160 3846
rect 3192 3846 3364 3848
rect 3162 3824 3190 3828
rect 3192 3824 3272 3846
rect 3293 3844 3308 3846
rect 3162 3822 3272 3824
rect 3093 3818 3272 3822
rect 3066 3808 3096 3818
rect 3098 3808 3251 3818
rect 3259 3808 3289 3818
rect 3293 3808 3323 3822
rect 3351 3808 3364 3846
rect 3436 3852 3471 3860
rect 3436 3826 3437 3852
rect 3444 3826 3471 3852
rect 3379 3808 3409 3822
rect 3436 3818 3471 3826
rect 3473 3852 3514 3860
rect 3473 3826 3488 3852
rect 3495 3826 3514 3852
rect 3578 3848 3640 3860
rect 3652 3848 3727 3860
rect 3785 3848 3860 3860
rect 3872 3848 3903 3860
rect 3909 3848 3944 3860
rect 3578 3846 3740 3848
rect 3473 3818 3514 3826
rect 3596 3822 3609 3846
rect 3624 3844 3639 3846
rect 3436 3808 3437 3818
rect 3452 3808 3465 3818
rect 3479 3808 3480 3818
rect 3495 3808 3508 3818
rect 3523 3808 3553 3822
rect 3596 3808 3639 3822
rect 3663 3819 3670 3826
rect 3673 3822 3740 3846
rect 3772 3846 3944 3848
rect 3742 3824 3770 3828
rect 3772 3824 3852 3846
rect 3873 3844 3888 3846
rect 3742 3822 3852 3824
rect 3673 3818 3852 3822
rect 3646 3808 3676 3818
rect 3678 3808 3831 3818
rect 3839 3808 3869 3818
rect 3873 3808 3903 3822
rect 3931 3808 3944 3846
rect 4016 3852 4051 3860
rect 4016 3826 4017 3852
rect 4024 3826 4051 3852
rect 3959 3808 3989 3822
rect 4016 3818 4051 3826
rect 4053 3852 4094 3860
rect 4053 3826 4068 3852
rect 4075 3826 4094 3852
rect 4158 3848 4220 3860
rect 4232 3848 4307 3860
rect 4365 3848 4440 3860
rect 4452 3848 4483 3860
rect 4489 3848 4524 3860
rect 4158 3846 4320 3848
rect 4053 3818 4094 3826
rect 4176 3822 4189 3846
rect 4204 3844 4219 3846
rect 4016 3808 4017 3818
rect 4032 3808 4045 3818
rect 4059 3808 4060 3818
rect 4075 3808 4088 3818
rect 4103 3808 4133 3822
rect 4176 3808 4219 3822
rect 4243 3819 4250 3826
rect 4253 3822 4320 3846
rect 4352 3846 4524 3848
rect 4322 3824 4350 3828
rect 4352 3824 4432 3846
rect 4453 3844 4468 3846
rect 4322 3822 4432 3824
rect 4253 3818 4432 3822
rect 4226 3808 4256 3818
rect 4258 3808 4411 3818
rect 4419 3808 4449 3818
rect 4453 3808 4483 3822
rect 4511 3808 4524 3846
rect 4596 3852 4631 3860
rect 4596 3826 4597 3852
rect 4604 3826 4631 3852
rect 4539 3808 4569 3822
rect 4596 3818 4631 3826
rect 4596 3808 4597 3818
rect 4612 3808 4625 3818
rect -1 3802 4625 3808
rect 0 3794 4625 3802
rect 15 3764 28 3794
rect 43 3776 73 3794
rect 116 3780 130 3794
rect 166 3780 386 3794
rect 117 3778 130 3780
rect 83 3766 98 3778
rect 80 3764 102 3766
rect 107 3764 137 3778
rect 198 3776 351 3780
rect 180 3764 372 3776
rect 415 3764 445 3778
rect 451 3764 464 3794
rect 479 3776 509 3794
rect 552 3764 565 3794
rect 595 3764 608 3794
rect 623 3776 653 3794
rect 696 3780 710 3794
rect 746 3780 966 3794
rect 697 3778 710 3780
rect 663 3766 678 3778
rect 660 3764 682 3766
rect 687 3764 717 3778
rect 778 3776 931 3780
rect 760 3764 952 3776
rect 995 3764 1025 3778
rect 1031 3764 1044 3794
rect 1059 3776 1089 3794
rect 1132 3764 1145 3794
rect 1175 3764 1188 3794
rect 1203 3776 1233 3794
rect 1276 3780 1290 3794
rect 1326 3780 1546 3794
rect 1277 3778 1290 3780
rect 1243 3766 1258 3778
rect 1240 3764 1262 3766
rect 1267 3764 1297 3778
rect 1358 3776 1511 3780
rect 1340 3764 1532 3776
rect 1575 3764 1605 3778
rect 1611 3764 1624 3794
rect 1639 3776 1669 3794
rect 1712 3764 1725 3794
rect 1755 3764 1768 3794
rect 1783 3776 1813 3794
rect 1856 3780 1870 3794
rect 1906 3780 2126 3794
rect 1857 3778 1870 3780
rect 1823 3766 1838 3778
rect 1820 3764 1842 3766
rect 1847 3764 1877 3778
rect 1938 3776 2091 3780
rect 1920 3764 2112 3776
rect 2155 3764 2185 3778
rect 2191 3764 2204 3794
rect 2219 3776 2249 3794
rect 2292 3764 2305 3794
rect 2335 3764 2348 3794
rect 2363 3776 2393 3794
rect 2436 3780 2450 3794
rect 2486 3780 2706 3794
rect 2437 3778 2450 3780
rect 2403 3766 2418 3778
rect 2400 3764 2422 3766
rect 2427 3764 2457 3778
rect 2518 3776 2671 3780
rect 2500 3764 2692 3776
rect 2735 3764 2765 3778
rect 2771 3764 2784 3794
rect 2799 3776 2829 3794
rect 2872 3764 2885 3794
rect 2915 3764 2928 3794
rect 2943 3776 2973 3794
rect 3016 3780 3030 3794
rect 3066 3780 3286 3794
rect 3017 3778 3030 3780
rect 2983 3766 2998 3778
rect 2980 3764 3002 3766
rect 3007 3764 3037 3778
rect 3098 3776 3251 3780
rect 3080 3764 3272 3776
rect 3315 3764 3345 3778
rect 3351 3764 3364 3794
rect 3379 3776 3409 3794
rect 3452 3764 3465 3794
rect 3495 3764 3508 3794
rect 3523 3776 3553 3794
rect 3596 3780 3610 3794
rect 3646 3780 3866 3794
rect 3597 3778 3610 3780
rect 3563 3766 3578 3778
rect 3560 3764 3582 3766
rect 3587 3764 3617 3778
rect 3678 3776 3831 3780
rect 3660 3764 3852 3776
rect 3895 3764 3925 3778
rect 3931 3764 3944 3794
rect 3959 3776 3989 3794
rect 4032 3764 4045 3794
rect 4075 3764 4088 3794
rect 4103 3776 4133 3794
rect 4176 3780 4190 3794
rect 4226 3780 4446 3794
rect 4177 3778 4190 3780
rect 4143 3766 4158 3778
rect 4140 3764 4162 3766
rect 4167 3764 4197 3778
rect 4258 3776 4411 3780
rect 4240 3764 4432 3776
rect 4475 3764 4505 3778
rect 4511 3764 4524 3794
rect 4539 3776 4569 3794
rect 4612 3764 4625 3794
rect 0 3750 4625 3764
rect 15 3646 28 3750
rect 73 3728 74 3738
rect 89 3728 102 3738
rect 73 3724 102 3728
rect 107 3724 137 3750
rect 155 3736 171 3738
rect 243 3736 296 3750
rect 244 3734 308 3736
rect 351 3734 366 3750
rect 415 3747 445 3750
rect 415 3744 451 3747
rect 381 3736 397 3738
rect 155 3724 170 3728
rect 73 3722 170 3724
rect 198 3722 366 3734
rect 382 3724 397 3728
rect 415 3725 454 3744
rect 473 3738 480 3739
rect 479 3731 480 3738
rect 463 3728 464 3731
rect 479 3728 492 3731
rect 415 3724 445 3725
rect 454 3724 460 3725
rect 463 3724 492 3728
rect 382 3723 492 3724
rect 382 3722 498 3723
rect 57 3714 108 3722
rect 57 3702 82 3714
rect 89 3702 108 3714
rect 139 3714 189 3722
rect 139 3706 155 3714
rect 162 3712 189 3714
rect 198 3712 419 3722
rect 162 3702 419 3712
rect 448 3714 498 3722
rect 448 3705 464 3714
rect 57 3694 108 3702
rect 155 3694 419 3702
rect 445 3702 464 3705
rect 471 3702 498 3714
rect 445 3694 498 3702
rect 73 3686 74 3694
rect 89 3686 102 3694
rect 73 3678 89 3686
rect 70 3671 89 3674
rect 70 3662 92 3671
rect 43 3652 92 3662
rect 43 3646 73 3652
rect 92 3647 97 3652
rect 15 3630 89 3646
rect 107 3638 137 3694
rect 172 3684 380 3694
rect 415 3690 460 3694
rect 463 3693 464 3694
rect 479 3693 492 3694
rect 198 3654 387 3684
rect 213 3651 387 3654
rect 206 3648 387 3651
rect 15 3628 28 3630
rect 43 3628 77 3630
rect 15 3612 89 3628
rect 116 3624 129 3638
rect 144 3624 160 3640
rect 206 3635 217 3648
rect -1 3590 0 3606
rect 15 3590 28 3612
rect 43 3590 73 3612
rect 116 3608 178 3624
rect 206 3617 217 3633
rect 222 3628 232 3648
rect 242 3628 256 3648
rect 259 3635 268 3648
rect 284 3635 293 3648
rect 222 3617 256 3628
rect 259 3617 268 3633
rect 284 3617 293 3633
rect 300 3628 310 3648
rect 320 3628 334 3648
rect 335 3635 346 3648
rect 300 3617 334 3628
rect 335 3617 346 3633
rect 392 3624 408 3640
rect 415 3638 445 3690
rect 479 3686 480 3693
rect 464 3678 480 3686
rect 451 3646 464 3665
rect 479 3646 509 3662
rect 451 3630 525 3646
rect 451 3628 464 3630
rect 479 3628 513 3630
rect 116 3606 129 3608
rect 144 3606 178 3608
rect 116 3590 178 3606
rect 222 3601 238 3604
rect 300 3601 330 3612
rect 378 3608 424 3624
rect 451 3612 525 3628
rect 378 3606 412 3608
rect 377 3590 424 3606
rect 451 3590 464 3612
rect 479 3590 509 3612
rect 536 3590 537 3606
rect 552 3590 565 3750
rect 595 3646 608 3750
rect 653 3728 654 3738
rect 669 3728 682 3738
rect 653 3724 682 3728
rect 687 3724 717 3750
rect 735 3736 751 3738
rect 823 3736 876 3750
rect 824 3734 888 3736
rect 931 3734 946 3750
rect 995 3747 1025 3750
rect 995 3744 1031 3747
rect 961 3736 977 3738
rect 735 3724 750 3728
rect 653 3722 750 3724
rect 778 3722 946 3734
rect 962 3724 977 3728
rect 995 3725 1034 3744
rect 1053 3738 1060 3739
rect 1059 3731 1060 3738
rect 1043 3728 1044 3731
rect 1059 3728 1072 3731
rect 995 3724 1025 3725
rect 1034 3724 1040 3725
rect 1043 3724 1072 3728
rect 962 3723 1072 3724
rect 962 3722 1078 3723
rect 637 3714 688 3722
rect 637 3702 662 3714
rect 669 3702 688 3714
rect 719 3714 769 3722
rect 719 3706 735 3714
rect 742 3712 769 3714
rect 778 3712 999 3722
rect 742 3702 999 3712
rect 1028 3714 1078 3722
rect 1028 3705 1044 3714
rect 637 3694 688 3702
rect 735 3694 999 3702
rect 1025 3702 1044 3705
rect 1051 3702 1078 3714
rect 1025 3694 1078 3702
rect 653 3686 654 3694
rect 669 3686 682 3694
rect 653 3678 669 3686
rect 650 3671 669 3674
rect 650 3662 672 3671
rect 623 3652 672 3662
rect 623 3646 653 3652
rect 672 3647 677 3652
rect 595 3630 669 3646
rect 687 3638 717 3694
rect 752 3684 960 3694
rect 995 3690 1040 3694
rect 1043 3693 1044 3694
rect 1059 3693 1072 3694
rect 778 3654 967 3684
rect 793 3651 967 3654
rect 786 3648 967 3651
rect 595 3628 608 3630
rect 623 3628 657 3630
rect 595 3612 669 3628
rect 696 3624 709 3638
rect 724 3624 740 3640
rect 786 3635 797 3648
rect 579 3590 580 3606
rect 595 3590 608 3612
rect 623 3590 653 3612
rect 696 3608 758 3624
rect 786 3617 797 3633
rect 802 3628 812 3648
rect 822 3628 836 3648
rect 839 3635 848 3648
rect 864 3635 873 3648
rect 802 3617 836 3628
rect 839 3617 848 3633
rect 864 3617 873 3633
rect 880 3628 890 3648
rect 900 3628 914 3648
rect 915 3635 926 3648
rect 880 3617 914 3628
rect 915 3617 926 3633
rect 972 3624 988 3640
rect 995 3638 1025 3690
rect 1059 3686 1060 3693
rect 1044 3678 1060 3686
rect 1031 3646 1044 3665
rect 1059 3646 1089 3662
rect 1031 3630 1105 3646
rect 1031 3628 1044 3630
rect 1059 3628 1093 3630
rect 696 3606 709 3608
rect 724 3606 758 3608
rect 696 3590 758 3606
rect 802 3601 818 3604
rect 880 3601 910 3612
rect 958 3608 1004 3624
rect 1031 3612 1105 3628
rect 958 3606 992 3608
rect 957 3590 1004 3606
rect 1031 3590 1044 3612
rect 1059 3590 1089 3612
rect 1116 3590 1117 3606
rect 1132 3590 1145 3750
rect 1175 3646 1188 3750
rect 1233 3728 1234 3738
rect 1249 3728 1262 3738
rect 1233 3724 1262 3728
rect 1267 3724 1297 3750
rect 1315 3736 1331 3738
rect 1403 3736 1456 3750
rect 1404 3734 1468 3736
rect 1511 3734 1526 3750
rect 1575 3747 1605 3750
rect 1575 3744 1611 3747
rect 1541 3736 1557 3738
rect 1315 3724 1330 3728
rect 1233 3722 1330 3724
rect 1358 3722 1526 3734
rect 1542 3724 1557 3728
rect 1575 3725 1614 3744
rect 1633 3738 1640 3739
rect 1639 3731 1640 3738
rect 1623 3728 1624 3731
rect 1639 3728 1652 3731
rect 1575 3724 1605 3725
rect 1614 3724 1620 3725
rect 1623 3724 1652 3728
rect 1542 3723 1652 3724
rect 1542 3722 1658 3723
rect 1217 3714 1268 3722
rect 1217 3702 1242 3714
rect 1249 3702 1268 3714
rect 1299 3714 1349 3722
rect 1299 3706 1315 3714
rect 1322 3712 1349 3714
rect 1358 3712 1579 3722
rect 1322 3702 1579 3712
rect 1608 3714 1658 3722
rect 1608 3705 1624 3714
rect 1217 3694 1268 3702
rect 1315 3694 1579 3702
rect 1605 3702 1624 3705
rect 1631 3702 1658 3714
rect 1605 3694 1658 3702
rect 1233 3686 1234 3694
rect 1249 3686 1262 3694
rect 1233 3678 1249 3686
rect 1230 3671 1249 3674
rect 1230 3662 1252 3671
rect 1203 3652 1252 3662
rect 1203 3646 1233 3652
rect 1252 3647 1257 3652
rect 1175 3630 1249 3646
rect 1267 3638 1297 3694
rect 1332 3684 1540 3694
rect 1575 3690 1620 3694
rect 1623 3693 1624 3694
rect 1639 3693 1652 3694
rect 1358 3654 1547 3684
rect 1373 3651 1547 3654
rect 1366 3648 1547 3651
rect 1175 3628 1188 3630
rect 1203 3628 1237 3630
rect 1175 3612 1249 3628
rect 1276 3624 1289 3638
rect 1304 3624 1320 3640
rect 1366 3635 1377 3648
rect 1159 3590 1160 3606
rect 1175 3590 1188 3612
rect 1203 3590 1233 3612
rect 1276 3608 1338 3624
rect 1366 3617 1377 3633
rect 1382 3628 1392 3648
rect 1402 3628 1416 3648
rect 1419 3635 1428 3648
rect 1444 3635 1453 3648
rect 1382 3617 1416 3628
rect 1419 3617 1428 3633
rect 1444 3617 1453 3633
rect 1460 3628 1470 3648
rect 1480 3628 1494 3648
rect 1495 3635 1506 3648
rect 1460 3617 1494 3628
rect 1495 3617 1506 3633
rect 1552 3624 1568 3640
rect 1575 3638 1605 3690
rect 1639 3686 1640 3693
rect 1624 3678 1640 3686
rect 1611 3646 1624 3665
rect 1639 3646 1669 3662
rect 1611 3630 1685 3646
rect 1611 3628 1624 3630
rect 1639 3628 1673 3630
rect 1276 3606 1289 3608
rect 1304 3606 1338 3608
rect 1276 3590 1338 3606
rect 1382 3601 1398 3604
rect 1460 3601 1490 3612
rect 1538 3608 1584 3624
rect 1611 3612 1685 3628
rect 1538 3606 1572 3608
rect 1537 3590 1584 3606
rect 1611 3590 1624 3612
rect 1639 3590 1669 3612
rect 1696 3590 1697 3606
rect 1712 3590 1725 3750
rect 1755 3646 1768 3750
rect 1813 3728 1814 3738
rect 1829 3728 1842 3738
rect 1813 3724 1842 3728
rect 1847 3724 1877 3750
rect 1895 3736 1911 3738
rect 1983 3736 2036 3750
rect 1984 3734 2048 3736
rect 2091 3734 2106 3750
rect 2155 3747 2185 3750
rect 2155 3744 2191 3747
rect 2121 3736 2137 3738
rect 1895 3724 1910 3728
rect 1813 3722 1910 3724
rect 1938 3722 2106 3734
rect 2122 3724 2137 3728
rect 2155 3725 2194 3744
rect 2213 3738 2220 3739
rect 2219 3731 2220 3738
rect 2203 3728 2204 3731
rect 2219 3728 2232 3731
rect 2155 3724 2185 3725
rect 2194 3724 2200 3725
rect 2203 3724 2232 3728
rect 2122 3723 2232 3724
rect 2122 3722 2238 3723
rect 1797 3714 1848 3722
rect 1797 3702 1822 3714
rect 1829 3702 1848 3714
rect 1879 3714 1929 3722
rect 1879 3706 1895 3714
rect 1902 3712 1929 3714
rect 1938 3712 2159 3722
rect 1902 3702 2159 3712
rect 2188 3714 2238 3722
rect 2188 3705 2204 3714
rect 1797 3694 1848 3702
rect 1895 3694 2159 3702
rect 2185 3702 2204 3705
rect 2211 3702 2238 3714
rect 2185 3694 2238 3702
rect 1813 3686 1814 3694
rect 1829 3686 1842 3694
rect 1813 3678 1829 3686
rect 1810 3671 1829 3674
rect 1810 3662 1832 3671
rect 1783 3652 1832 3662
rect 1783 3646 1813 3652
rect 1832 3647 1837 3652
rect 1755 3630 1829 3646
rect 1847 3638 1877 3694
rect 1912 3684 2120 3694
rect 2155 3690 2200 3694
rect 2203 3693 2204 3694
rect 2219 3693 2232 3694
rect 1938 3654 2127 3684
rect 1953 3651 2127 3654
rect 1946 3648 2127 3651
rect 1755 3628 1768 3630
rect 1783 3628 1817 3630
rect 1755 3612 1829 3628
rect 1856 3624 1869 3638
rect 1884 3624 1900 3640
rect 1946 3635 1957 3648
rect 1739 3590 1740 3606
rect 1755 3590 1768 3612
rect 1783 3590 1813 3612
rect 1856 3608 1918 3624
rect 1946 3617 1957 3633
rect 1962 3628 1972 3648
rect 1982 3628 1996 3648
rect 1999 3635 2008 3648
rect 2024 3635 2033 3648
rect 1962 3617 1996 3628
rect 1999 3617 2008 3633
rect 2024 3617 2033 3633
rect 2040 3628 2050 3648
rect 2060 3628 2074 3648
rect 2075 3635 2086 3648
rect 2040 3617 2074 3628
rect 2075 3617 2086 3633
rect 2132 3624 2148 3640
rect 2155 3638 2185 3690
rect 2219 3686 2220 3693
rect 2204 3678 2220 3686
rect 2191 3646 2204 3665
rect 2219 3646 2249 3662
rect 2191 3630 2265 3646
rect 2191 3628 2204 3630
rect 2219 3628 2253 3630
rect 1856 3606 1869 3608
rect 1884 3606 1918 3608
rect 1856 3590 1918 3606
rect 1962 3601 1978 3604
rect 2040 3601 2070 3612
rect 2118 3608 2164 3624
rect 2191 3612 2265 3628
rect 2118 3606 2152 3608
rect 2117 3590 2164 3606
rect 2191 3590 2204 3612
rect 2219 3590 2249 3612
rect 2276 3590 2277 3606
rect 2292 3590 2305 3750
rect 2335 3646 2348 3750
rect 2393 3728 2394 3738
rect 2409 3728 2422 3738
rect 2393 3724 2422 3728
rect 2427 3724 2457 3750
rect 2475 3736 2491 3738
rect 2563 3736 2616 3750
rect 2564 3734 2628 3736
rect 2671 3734 2686 3750
rect 2735 3747 2765 3750
rect 2735 3744 2771 3747
rect 2701 3736 2717 3738
rect 2475 3724 2490 3728
rect 2393 3722 2490 3724
rect 2518 3722 2686 3734
rect 2702 3724 2717 3728
rect 2735 3725 2774 3744
rect 2793 3738 2800 3739
rect 2799 3731 2800 3738
rect 2783 3728 2784 3731
rect 2799 3728 2812 3731
rect 2735 3724 2765 3725
rect 2774 3724 2780 3725
rect 2783 3724 2812 3728
rect 2702 3723 2812 3724
rect 2702 3722 2818 3723
rect 2377 3714 2428 3722
rect 2377 3702 2402 3714
rect 2409 3702 2428 3714
rect 2459 3714 2509 3722
rect 2459 3706 2475 3714
rect 2482 3712 2509 3714
rect 2518 3712 2739 3722
rect 2482 3702 2739 3712
rect 2768 3714 2818 3722
rect 2768 3705 2784 3714
rect 2377 3694 2428 3702
rect 2475 3694 2739 3702
rect 2765 3702 2784 3705
rect 2791 3702 2818 3714
rect 2765 3694 2818 3702
rect 2393 3686 2394 3694
rect 2409 3686 2422 3694
rect 2393 3678 2409 3686
rect 2390 3671 2409 3674
rect 2390 3662 2412 3671
rect 2363 3652 2412 3662
rect 2363 3646 2393 3652
rect 2412 3647 2417 3652
rect 2335 3630 2409 3646
rect 2427 3638 2457 3694
rect 2492 3684 2700 3694
rect 2735 3690 2780 3694
rect 2783 3693 2784 3694
rect 2799 3693 2812 3694
rect 2518 3654 2707 3684
rect 2533 3651 2707 3654
rect 2526 3648 2707 3651
rect 2335 3628 2348 3630
rect 2363 3628 2397 3630
rect 2335 3612 2409 3628
rect 2436 3624 2449 3638
rect 2464 3624 2480 3640
rect 2526 3635 2537 3648
rect 2319 3590 2320 3606
rect 2335 3590 2348 3612
rect 2363 3590 2393 3612
rect 2436 3608 2498 3624
rect 2526 3617 2537 3633
rect 2542 3628 2552 3648
rect 2562 3628 2576 3648
rect 2579 3635 2588 3648
rect 2604 3635 2613 3648
rect 2542 3617 2576 3628
rect 2579 3617 2588 3633
rect 2604 3617 2613 3633
rect 2620 3628 2630 3648
rect 2640 3628 2654 3648
rect 2655 3635 2666 3648
rect 2620 3617 2654 3628
rect 2655 3617 2666 3633
rect 2712 3624 2728 3640
rect 2735 3638 2765 3690
rect 2799 3686 2800 3693
rect 2784 3678 2800 3686
rect 2771 3646 2784 3665
rect 2799 3646 2829 3662
rect 2771 3630 2845 3646
rect 2771 3628 2784 3630
rect 2799 3628 2833 3630
rect 2436 3606 2449 3608
rect 2464 3606 2498 3608
rect 2436 3590 2498 3606
rect 2542 3601 2558 3604
rect 2620 3601 2650 3612
rect 2698 3608 2744 3624
rect 2771 3612 2845 3628
rect 2698 3606 2732 3608
rect 2697 3590 2744 3606
rect 2771 3590 2784 3612
rect 2799 3590 2829 3612
rect 2856 3590 2857 3606
rect 2872 3590 2885 3750
rect 2915 3646 2928 3750
rect 2973 3728 2974 3738
rect 2989 3728 3002 3738
rect 2973 3724 3002 3728
rect 3007 3724 3037 3750
rect 3055 3736 3071 3738
rect 3143 3736 3196 3750
rect 3144 3734 3208 3736
rect 3251 3734 3266 3750
rect 3315 3747 3345 3750
rect 3315 3744 3351 3747
rect 3281 3736 3297 3738
rect 3055 3724 3070 3728
rect 2973 3722 3070 3724
rect 3098 3722 3266 3734
rect 3282 3724 3297 3728
rect 3315 3725 3354 3744
rect 3373 3738 3380 3739
rect 3379 3731 3380 3738
rect 3363 3728 3364 3731
rect 3379 3728 3392 3731
rect 3315 3724 3345 3725
rect 3354 3724 3360 3725
rect 3363 3724 3392 3728
rect 3282 3723 3392 3724
rect 3282 3722 3398 3723
rect 2957 3714 3008 3722
rect 2957 3702 2982 3714
rect 2989 3702 3008 3714
rect 3039 3714 3089 3722
rect 3039 3706 3055 3714
rect 3062 3712 3089 3714
rect 3098 3712 3319 3722
rect 3062 3702 3319 3712
rect 3348 3714 3398 3722
rect 3348 3705 3364 3714
rect 2957 3694 3008 3702
rect 3055 3694 3319 3702
rect 3345 3702 3364 3705
rect 3371 3702 3398 3714
rect 3345 3694 3398 3702
rect 2973 3686 2974 3694
rect 2989 3686 3002 3694
rect 2973 3678 2989 3686
rect 2970 3671 2989 3674
rect 2970 3662 2992 3671
rect 2943 3652 2992 3662
rect 2943 3646 2973 3652
rect 2992 3647 2997 3652
rect 2915 3630 2989 3646
rect 3007 3638 3037 3694
rect 3072 3684 3280 3694
rect 3315 3690 3360 3694
rect 3363 3693 3364 3694
rect 3379 3693 3392 3694
rect 3098 3654 3287 3684
rect 3113 3651 3287 3654
rect 3106 3648 3287 3651
rect 2915 3628 2928 3630
rect 2943 3628 2977 3630
rect 2915 3612 2989 3628
rect 3016 3624 3029 3638
rect 3044 3624 3060 3640
rect 3106 3635 3117 3648
rect 2899 3590 2900 3606
rect 2915 3590 2928 3612
rect 2943 3590 2973 3612
rect 3016 3608 3078 3624
rect 3106 3617 3117 3633
rect 3122 3628 3132 3648
rect 3142 3628 3156 3648
rect 3159 3635 3168 3648
rect 3184 3635 3193 3648
rect 3122 3617 3156 3628
rect 3159 3617 3168 3633
rect 3184 3617 3193 3633
rect 3200 3628 3210 3648
rect 3220 3628 3234 3648
rect 3235 3635 3246 3648
rect 3200 3617 3234 3628
rect 3235 3617 3246 3633
rect 3292 3624 3308 3640
rect 3315 3638 3345 3690
rect 3379 3686 3380 3693
rect 3364 3678 3380 3686
rect 3351 3646 3364 3665
rect 3379 3646 3409 3662
rect 3351 3630 3425 3646
rect 3351 3628 3364 3630
rect 3379 3628 3413 3630
rect 3016 3606 3029 3608
rect 3044 3606 3078 3608
rect 3016 3590 3078 3606
rect 3122 3601 3138 3604
rect 3200 3601 3230 3612
rect 3278 3608 3324 3624
rect 3351 3612 3425 3628
rect 3278 3606 3312 3608
rect 3277 3590 3324 3606
rect 3351 3590 3364 3612
rect 3379 3590 3409 3612
rect 3436 3590 3437 3606
rect 3452 3590 3465 3750
rect 3495 3646 3508 3750
rect 3553 3728 3554 3738
rect 3569 3728 3582 3738
rect 3553 3724 3582 3728
rect 3587 3724 3617 3750
rect 3635 3736 3651 3738
rect 3723 3736 3776 3750
rect 3724 3734 3788 3736
rect 3831 3734 3846 3750
rect 3895 3747 3925 3750
rect 3895 3744 3931 3747
rect 3861 3736 3877 3738
rect 3635 3724 3650 3728
rect 3553 3722 3650 3724
rect 3678 3722 3846 3734
rect 3862 3724 3877 3728
rect 3895 3725 3934 3744
rect 3953 3738 3960 3739
rect 3959 3731 3960 3738
rect 3943 3728 3944 3731
rect 3959 3728 3972 3731
rect 3895 3724 3925 3725
rect 3934 3724 3940 3725
rect 3943 3724 3972 3728
rect 3862 3723 3972 3724
rect 3862 3722 3978 3723
rect 3537 3714 3588 3722
rect 3537 3702 3562 3714
rect 3569 3702 3588 3714
rect 3619 3714 3669 3722
rect 3619 3706 3635 3714
rect 3642 3712 3669 3714
rect 3678 3712 3899 3722
rect 3642 3702 3899 3712
rect 3928 3714 3978 3722
rect 3928 3705 3944 3714
rect 3537 3694 3588 3702
rect 3635 3694 3899 3702
rect 3925 3702 3944 3705
rect 3951 3702 3978 3714
rect 3925 3694 3978 3702
rect 3553 3686 3554 3694
rect 3569 3686 3582 3694
rect 3553 3678 3569 3686
rect 3550 3671 3569 3674
rect 3550 3662 3572 3671
rect 3523 3652 3572 3662
rect 3523 3646 3553 3652
rect 3572 3647 3577 3652
rect 3495 3630 3569 3646
rect 3587 3638 3617 3694
rect 3652 3684 3860 3694
rect 3895 3690 3940 3694
rect 3943 3693 3944 3694
rect 3959 3693 3972 3694
rect 3678 3654 3867 3684
rect 3693 3651 3867 3654
rect 3686 3648 3867 3651
rect 3495 3628 3508 3630
rect 3523 3628 3557 3630
rect 3495 3612 3569 3628
rect 3596 3624 3609 3638
rect 3624 3624 3640 3640
rect 3686 3635 3697 3648
rect 3479 3590 3480 3606
rect 3495 3590 3508 3612
rect 3523 3590 3553 3612
rect 3596 3608 3658 3624
rect 3686 3617 3697 3633
rect 3702 3628 3712 3648
rect 3722 3628 3736 3648
rect 3739 3635 3748 3648
rect 3764 3635 3773 3648
rect 3702 3617 3736 3628
rect 3739 3617 3748 3633
rect 3764 3617 3773 3633
rect 3780 3628 3790 3648
rect 3800 3628 3814 3648
rect 3815 3635 3826 3648
rect 3780 3617 3814 3628
rect 3815 3617 3826 3633
rect 3872 3624 3888 3640
rect 3895 3638 3925 3690
rect 3959 3686 3960 3693
rect 3944 3678 3960 3686
rect 3931 3646 3944 3665
rect 3959 3646 3989 3662
rect 3931 3630 4005 3646
rect 3931 3628 3944 3630
rect 3959 3628 3993 3630
rect 3596 3606 3609 3608
rect 3624 3606 3658 3608
rect 3596 3590 3658 3606
rect 3702 3601 3718 3604
rect 3780 3601 3810 3612
rect 3858 3608 3904 3624
rect 3931 3612 4005 3628
rect 3858 3606 3892 3608
rect 3857 3590 3904 3606
rect 3931 3590 3944 3612
rect 3959 3590 3989 3612
rect 4016 3590 4017 3606
rect 4032 3590 4045 3750
rect 4075 3646 4088 3750
rect 4133 3728 4134 3738
rect 4149 3728 4162 3738
rect 4133 3724 4162 3728
rect 4167 3724 4197 3750
rect 4215 3736 4231 3738
rect 4303 3736 4356 3750
rect 4304 3734 4368 3736
rect 4411 3734 4426 3750
rect 4475 3747 4505 3750
rect 4475 3744 4511 3747
rect 4441 3736 4457 3738
rect 4215 3724 4230 3728
rect 4133 3722 4230 3724
rect 4258 3722 4426 3734
rect 4442 3724 4457 3728
rect 4475 3725 4514 3744
rect 4533 3738 4540 3739
rect 4539 3731 4540 3738
rect 4523 3728 4524 3731
rect 4539 3728 4552 3731
rect 4475 3724 4505 3725
rect 4514 3724 4520 3725
rect 4523 3724 4552 3728
rect 4442 3723 4552 3724
rect 4442 3722 4558 3723
rect 4117 3714 4168 3722
rect 4117 3702 4142 3714
rect 4149 3702 4168 3714
rect 4199 3714 4249 3722
rect 4199 3706 4215 3714
rect 4222 3712 4249 3714
rect 4258 3712 4479 3722
rect 4222 3702 4479 3712
rect 4508 3714 4558 3722
rect 4508 3705 4524 3714
rect 4117 3694 4168 3702
rect 4215 3694 4479 3702
rect 4505 3702 4524 3705
rect 4531 3702 4558 3714
rect 4505 3694 4558 3702
rect 4133 3686 4134 3694
rect 4149 3686 4162 3694
rect 4133 3678 4149 3686
rect 4130 3671 4149 3674
rect 4130 3662 4152 3671
rect 4103 3652 4152 3662
rect 4103 3646 4133 3652
rect 4152 3647 4157 3652
rect 4075 3630 4149 3646
rect 4167 3638 4197 3694
rect 4232 3684 4440 3694
rect 4475 3690 4520 3694
rect 4523 3693 4524 3694
rect 4539 3693 4552 3694
rect 4258 3654 4447 3684
rect 4273 3651 4447 3654
rect 4266 3648 4447 3651
rect 4075 3628 4088 3630
rect 4103 3628 4137 3630
rect 4075 3612 4149 3628
rect 4176 3624 4189 3638
rect 4204 3624 4220 3640
rect 4266 3635 4277 3648
rect 4059 3590 4060 3606
rect 4075 3590 4088 3612
rect 4103 3590 4133 3612
rect 4176 3608 4238 3624
rect 4266 3617 4277 3633
rect 4282 3628 4292 3648
rect 4302 3628 4316 3648
rect 4319 3635 4328 3648
rect 4344 3635 4353 3648
rect 4282 3617 4316 3628
rect 4319 3617 4328 3633
rect 4344 3617 4353 3633
rect 4360 3628 4370 3648
rect 4380 3628 4394 3648
rect 4395 3635 4406 3648
rect 4360 3617 4394 3628
rect 4395 3617 4406 3633
rect 4452 3624 4468 3640
rect 4475 3638 4505 3690
rect 4539 3686 4540 3693
rect 4524 3678 4540 3686
rect 4511 3646 4524 3665
rect 4539 3646 4569 3662
rect 4511 3630 4585 3646
rect 4511 3628 4524 3630
rect 4539 3628 4573 3630
rect 4176 3606 4189 3608
rect 4204 3606 4238 3608
rect 4176 3590 4238 3606
rect 4282 3601 4298 3604
rect 4360 3601 4390 3612
rect 4438 3608 4484 3624
rect 4511 3612 4585 3628
rect 4438 3606 4472 3608
rect 4437 3590 4484 3606
rect 4511 3590 4524 3612
rect 4539 3590 4569 3612
rect 4596 3590 4597 3606
rect 4612 3590 4625 3750
rect -7 3582 34 3590
rect -7 3556 8 3582
rect 15 3556 34 3582
rect 98 3578 160 3590
rect 172 3578 247 3590
rect 305 3578 380 3590
rect 392 3578 423 3590
rect 429 3578 464 3590
rect 98 3576 260 3578
rect -7 3548 34 3556
rect 116 3552 129 3576
rect 144 3574 159 3576
rect -1 3538 0 3548
rect 15 3538 28 3548
rect 43 3538 73 3552
rect 116 3538 159 3552
rect 183 3549 190 3556
rect 193 3552 260 3576
rect 292 3576 464 3578
rect 262 3554 290 3558
rect 292 3554 372 3576
rect 393 3574 408 3576
rect 262 3552 372 3554
rect 193 3548 372 3552
rect 166 3538 196 3548
rect 198 3538 351 3548
rect 359 3538 389 3548
rect 393 3538 423 3552
rect 451 3538 464 3576
rect 536 3582 571 3590
rect 536 3556 537 3582
rect 544 3556 571 3582
rect 479 3538 509 3552
rect 536 3548 571 3556
rect 573 3582 614 3590
rect 573 3556 588 3582
rect 595 3556 614 3582
rect 678 3578 740 3590
rect 752 3578 827 3590
rect 885 3578 960 3590
rect 972 3578 1003 3590
rect 1009 3578 1044 3590
rect 678 3576 840 3578
rect 573 3548 614 3556
rect 696 3552 709 3576
rect 724 3574 739 3576
rect 536 3538 537 3548
rect 552 3538 565 3548
rect 579 3538 580 3548
rect 595 3538 608 3548
rect 623 3538 653 3552
rect 696 3538 739 3552
rect 763 3549 770 3556
rect 773 3552 840 3576
rect 872 3576 1044 3578
rect 842 3554 870 3558
rect 872 3554 952 3576
rect 973 3574 988 3576
rect 842 3552 952 3554
rect 773 3548 952 3552
rect 746 3538 776 3548
rect 778 3538 931 3548
rect 939 3538 969 3548
rect 973 3538 1003 3552
rect 1031 3538 1044 3576
rect 1116 3582 1151 3590
rect 1116 3556 1117 3582
rect 1124 3556 1151 3582
rect 1059 3538 1089 3552
rect 1116 3548 1151 3556
rect 1153 3582 1194 3590
rect 1153 3556 1168 3582
rect 1175 3556 1194 3582
rect 1258 3578 1320 3590
rect 1332 3578 1407 3590
rect 1465 3578 1540 3590
rect 1552 3578 1583 3590
rect 1589 3578 1624 3590
rect 1258 3576 1420 3578
rect 1153 3548 1194 3556
rect 1276 3552 1289 3576
rect 1304 3574 1319 3576
rect 1116 3538 1117 3548
rect 1132 3538 1145 3548
rect 1159 3538 1160 3548
rect 1175 3538 1188 3548
rect 1203 3538 1233 3552
rect 1276 3538 1319 3552
rect 1343 3549 1350 3556
rect 1353 3552 1420 3576
rect 1452 3576 1624 3578
rect 1422 3554 1450 3558
rect 1452 3554 1532 3576
rect 1553 3574 1568 3576
rect 1422 3552 1532 3554
rect 1353 3548 1532 3552
rect 1326 3538 1356 3548
rect 1358 3538 1511 3548
rect 1519 3538 1549 3548
rect 1553 3538 1583 3552
rect 1611 3538 1624 3576
rect 1696 3582 1731 3590
rect 1696 3556 1697 3582
rect 1704 3556 1731 3582
rect 1639 3538 1669 3552
rect 1696 3548 1731 3556
rect 1733 3582 1774 3590
rect 1733 3556 1748 3582
rect 1755 3556 1774 3582
rect 1838 3578 1900 3590
rect 1912 3578 1987 3590
rect 2045 3578 2120 3590
rect 2132 3578 2163 3590
rect 2169 3578 2204 3590
rect 1838 3576 2000 3578
rect 1733 3548 1774 3556
rect 1856 3552 1869 3576
rect 1884 3574 1899 3576
rect 1696 3538 1697 3548
rect 1712 3538 1725 3548
rect 1739 3538 1740 3548
rect 1755 3538 1768 3548
rect 1783 3538 1813 3552
rect 1856 3538 1899 3552
rect 1923 3549 1930 3556
rect 1933 3552 2000 3576
rect 2032 3576 2204 3578
rect 2002 3554 2030 3558
rect 2032 3554 2112 3576
rect 2133 3574 2148 3576
rect 2002 3552 2112 3554
rect 1933 3548 2112 3552
rect 1906 3538 1936 3548
rect 1938 3538 2091 3548
rect 2099 3538 2129 3548
rect 2133 3538 2163 3552
rect 2191 3538 2204 3576
rect 2276 3582 2311 3590
rect 2276 3556 2277 3582
rect 2284 3556 2311 3582
rect 2219 3538 2249 3552
rect 2276 3548 2311 3556
rect 2313 3582 2354 3590
rect 2313 3556 2328 3582
rect 2335 3556 2354 3582
rect 2418 3578 2480 3590
rect 2492 3578 2567 3590
rect 2625 3578 2700 3590
rect 2712 3578 2743 3590
rect 2749 3578 2784 3590
rect 2418 3576 2580 3578
rect 2313 3548 2354 3556
rect 2436 3552 2449 3576
rect 2464 3574 2479 3576
rect 2276 3538 2277 3548
rect 2292 3538 2305 3548
rect 2319 3538 2320 3548
rect 2335 3538 2348 3548
rect 2363 3538 2393 3552
rect 2436 3538 2479 3552
rect 2503 3549 2510 3556
rect 2513 3552 2580 3576
rect 2612 3576 2784 3578
rect 2582 3554 2610 3558
rect 2612 3554 2692 3576
rect 2713 3574 2728 3576
rect 2582 3552 2692 3554
rect 2513 3548 2692 3552
rect 2486 3538 2516 3548
rect 2518 3538 2671 3548
rect 2679 3538 2709 3548
rect 2713 3538 2743 3552
rect 2771 3538 2784 3576
rect 2856 3582 2891 3590
rect 2856 3556 2857 3582
rect 2864 3556 2891 3582
rect 2799 3538 2829 3552
rect 2856 3548 2891 3556
rect 2893 3582 2934 3590
rect 2893 3556 2908 3582
rect 2915 3556 2934 3582
rect 2998 3578 3060 3590
rect 3072 3578 3147 3590
rect 3205 3578 3280 3590
rect 3292 3578 3323 3590
rect 3329 3578 3364 3590
rect 2998 3576 3160 3578
rect 2893 3548 2934 3556
rect 3016 3552 3029 3576
rect 3044 3574 3059 3576
rect 2856 3538 2857 3548
rect 2872 3538 2885 3548
rect 2899 3538 2900 3548
rect 2915 3538 2928 3548
rect 2943 3538 2973 3552
rect 3016 3538 3059 3552
rect 3083 3549 3090 3556
rect 3093 3552 3160 3576
rect 3192 3576 3364 3578
rect 3162 3554 3190 3558
rect 3192 3554 3272 3576
rect 3293 3574 3308 3576
rect 3162 3552 3272 3554
rect 3093 3548 3272 3552
rect 3066 3538 3096 3548
rect 3098 3538 3251 3548
rect 3259 3538 3289 3548
rect 3293 3538 3323 3552
rect 3351 3538 3364 3576
rect 3436 3582 3471 3590
rect 3436 3556 3437 3582
rect 3444 3556 3471 3582
rect 3379 3538 3409 3552
rect 3436 3548 3471 3556
rect 3473 3582 3514 3590
rect 3473 3556 3488 3582
rect 3495 3556 3514 3582
rect 3578 3578 3640 3590
rect 3652 3578 3727 3590
rect 3785 3578 3860 3590
rect 3872 3578 3903 3590
rect 3909 3578 3944 3590
rect 3578 3576 3740 3578
rect 3473 3548 3514 3556
rect 3596 3552 3609 3576
rect 3624 3574 3639 3576
rect 3436 3538 3437 3548
rect 3452 3538 3465 3548
rect 3479 3538 3480 3548
rect 3495 3538 3508 3548
rect 3523 3538 3553 3552
rect 3596 3538 3639 3552
rect 3663 3549 3670 3556
rect 3673 3552 3740 3576
rect 3772 3576 3944 3578
rect 3742 3554 3770 3558
rect 3772 3554 3852 3576
rect 3873 3574 3888 3576
rect 3742 3552 3852 3554
rect 3673 3548 3852 3552
rect 3646 3538 3676 3548
rect 3678 3538 3831 3548
rect 3839 3538 3869 3548
rect 3873 3538 3903 3552
rect 3931 3538 3944 3576
rect 4016 3582 4051 3590
rect 4016 3556 4017 3582
rect 4024 3556 4051 3582
rect 3959 3538 3989 3552
rect 4016 3548 4051 3556
rect 4053 3582 4094 3590
rect 4053 3556 4068 3582
rect 4075 3556 4094 3582
rect 4158 3578 4220 3590
rect 4232 3578 4307 3590
rect 4365 3578 4440 3590
rect 4452 3578 4483 3590
rect 4489 3578 4524 3590
rect 4158 3576 4320 3578
rect 4053 3548 4094 3556
rect 4176 3552 4189 3576
rect 4204 3574 4219 3576
rect 4016 3538 4017 3548
rect 4032 3538 4045 3548
rect 4059 3538 4060 3548
rect 4075 3538 4088 3548
rect 4103 3538 4133 3552
rect 4176 3538 4219 3552
rect 4243 3549 4250 3556
rect 4253 3552 4320 3576
rect 4352 3576 4524 3578
rect 4322 3554 4350 3558
rect 4352 3554 4432 3576
rect 4453 3574 4468 3576
rect 4322 3552 4432 3554
rect 4253 3548 4432 3552
rect 4226 3538 4256 3548
rect 4258 3538 4411 3548
rect 4419 3538 4449 3548
rect 4453 3538 4483 3552
rect 4511 3538 4524 3576
rect 4596 3582 4631 3590
rect 4596 3556 4597 3582
rect 4604 3556 4631 3582
rect 4539 3538 4569 3552
rect 4596 3548 4631 3556
rect 4596 3538 4597 3548
rect 4612 3538 4625 3548
rect -1 3532 4625 3538
rect 0 3524 4625 3532
rect 15 3494 28 3524
rect 43 3506 73 3524
rect 116 3510 130 3524
rect 166 3510 386 3524
rect 117 3508 130 3510
rect 83 3496 98 3508
rect 80 3494 102 3496
rect 107 3494 137 3508
rect 198 3506 351 3510
rect 180 3494 372 3506
rect 415 3494 445 3508
rect 451 3494 464 3524
rect 479 3506 509 3524
rect 552 3494 565 3524
rect 595 3494 608 3524
rect 623 3506 653 3524
rect 696 3510 710 3524
rect 746 3510 966 3524
rect 697 3508 710 3510
rect 663 3496 678 3508
rect 660 3494 682 3496
rect 687 3494 717 3508
rect 778 3506 931 3510
rect 760 3494 952 3506
rect 995 3494 1025 3508
rect 1031 3494 1044 3524
rect 1059 3506 1089 3524
rect 1132 3494 1145 3524
rect 1175 3494 1188 3524
rect 1203 3506 1233 3524
rect 1276 3510 1290 3524
rect 1326 3510 1546 3524
rect 1277 3508 1290 3510
rect 1243 3496 1258 3508
rect 1240 3494 1262 3496
rect 1267 3494 1297 3508
rect 1358 3506 1511 3510
rect 1340 3494 1532 3506
rect 1575 3494 1605 3508
rect 1611 3494 1624 3524
rect 1639 3506 1669 3524
rect 1712 3494 1725 3524
rect 1755 3494 1768 3524
rect 1783 3506 1813 3524
rect 1856 3510 1870 3524
rect 1906 3510 2126 3524
rect 1857 3508 1870 3510
rect 1823 3496 1838 3508
rect 1820 3494 1842 3496
rect 1847 3494 1877 3508
rect 1938 3506 2091 3510
rect 1920 3494 2112 3506
rect 2155 3494 2185 3508
rect 2191 3494 2204 3524
rect 2219 3506 2249 3524
rect 2292 3494 2305 3524
rect 2335 3494 2348 3524
rect 2363 3506 2393 3524
rect 2436 3510 2450 3524
rect 2486 3510 2706 3524
rect 2437 3508 2450 3510
rect 2403 3496 2418 3508
rect 2400 3494 2422 3496
rect 2427 3494 2457 3508
rect 2518 3506 2671 3510
rect 2500 3494 2692 3506
rect 2735 3494 2765 3508
rect 2771 3494 2784 3524
rect 2799 3506 2829 3524
rect 2872 3494 2885 3524
rect 2915 3494 2928 3524
rect 2943 3506 2973 3524
rect 3016 3510 3030 3524
rect 3066 3510 3286 3524
rect 3017 3508 3030 3510
rect 2983 3496 2998 3508
rect 2980 3494 3002 3496
rect 3007 3494 3037 3508
rect 3098 3506 3251 3510
rect 3080 3494 3272 3506
rect 3315 3494 3345 3508
rect 3351 3494 3364 3524
rect 3379 3506 3409 3524
rect 3452 3494 3465 3524
rect 3495 3494 3508 3524
rect 3523 3506 3553 3524
rect 3596 3510 3610 3524
rect 3646 3510 3866 3524
rect 3597 3508 3610 3510
rect 3563 3496 3578 3508
rect 3560 3494 3582 3496
rect 3587 3494 3617 3508
rect 3678 3506 3831 3510
rect 3660 3494 3852 3506
rect 3895 3494 3925 3508
rect 3931 3494 3944 3524
rect 3959 3506 3989 3524
rect 4032 3494 4045 3524
rect 4075 3494 4088 3524
rect 4103 3506 4133 3524
rect 4176 3510 4190 3524
rect 4226 3510 4446 3524
rect 4177 3508 4190 3510
rect 4143 3496 4158 3508
rect 4140 3494 4162 3496
rect 4167 3494 4197 3508
rect 4258 3506 4411 3510
rect 4240 3494 4432 3506
rect 4475 3494 4505 3508
rect 4511 3494 4524 3524
rect 4539 3506 4569 3524
rect 4612 3494 4625 3524
rect 0 3480 4625 3494
rect 15 3376 28 3480
rect 73 3458 74 3468
rect 89 3458 102 3468
rect 73 3454 102 3458
rect 107 3454 137 3480
rect 155 3466 171 3468
rect 243 3466 296 3480
rect 244 3464 308 3466
rect 351 3464 366 3480
rect 415 3477 445 3480
rect 415 3474 451 3477
rect 381 3466 397 3468
rect 155 3454 170 3458
rect 73 3452 170 3454
rect 198 3452 366 3464
rect 382 3454 397 3458
rect 415 3455 454 3474
rect 473 3468 480 3469
rect 479 3461 480 3468
rect 463 3458 464 3461
rect 479 3458 492 3461
rect 415 3454 445 3455
rect 454 3454 460 3455
rect 463 3454 492 3458
rect 382 3453 492 3454
rect 382 3452 498 3453
rect 57 3444 108 3452
rect 57 3432 82 3444
rect 89 3432 108 3444
rect 139 3444 189 3452
rect 139 3436 155 3444
rect 162 3442 189 3444
rect 198 3442 419 3452
rect 162 3432 419 3442
rect 448 3444 498 3452
rect 448 3435 464 3444
rect 57 3424 108 3432
rect 155 3424 419 3432
rect 445 3432 464 3435
rect 471 3432 498 3444
rect 445 3424 498 3432
rect 73 3416 74 3424
rect 89 3416 102 3424
rect 73 3408 89 3416
rect 70 3401 89 3404
rect 70 3392 92 3401
rect 43 3382 92 3392
rect 43 3376 73 3382
rect 92 3377 97 3382
rect 15 3360 89 3376
rect 107 3368 137 3424
rect 172 3414 380 3424
rect 415 3420 460 3424
rect 463 3423 464 3424
rect 479 3423 492 3424
rect 198 3384 387 3414
rect 213 3381 387 3384
rect 206 3378 387 3381
rect 15 3358 28 3360
rect 43 3358 77 3360
rect 15 3342 89 3358
rect 116 3354 129 3368
rect 144 3354 160 3370
rect 206 3365 217 3378
rect -1 3320 0 3336
rect 15 3320 28 3342
rect 43 3320 73 3342
rect 116 3338 178 3354
rect 206 3347 217 3363
rect 222 3358 232 3378
rect 242 3358 256 3378
rect 259 3365 268 3378
rect 284 3365 293 3378
rect 222 3347 256 3358
rect 259 3347 268 3363
rect 284 3347 293 3363
rect 300 3358 310 3378
rect 320 3358 334 3378
rect 335 3365 346 3378
rect 300 3347 334 3358
rect 335 3347 346 3363
rect 392 3354 408 3370
rect 415 3368 445 3420
rect 479 3416 480 3423
rect 464 3408 480 3416
rect 451 3376 464 3395
rect 479 3376 509 3392
rect 451 3360 525 3376
rect 451 3358 464 3360
rect 479 3358 513 3360
rect 116 3336 129 3338
rect 144 3336 178 3338
rect 116 3320 178 3336
rect 222 3331 238 3334
rect 300 3331 330 3342
rect 378 3338 424 3354
rect 451 3342 525 3358
rect 378 3336 412 3338
rect 377 3320 424 3336
rect 451 3320 464 3342
rect 479 3320 509 3342
rect 536 3320 537 3336
rect 552 3320 565 3480
rect 595 3376 608 3480
rect 653 3458 654 3468
rect 669 3458 682 3468
rect 653 3454 682 3458
rect 687 3454 717 3480
rect 735 3466 751 3468
rect 823 3466 876 3480
rect 824 3464 888 3466
rect 931 3464 946 3480
rect 995 3477 1025 3480
rect 995 3474 1031 3477
rect 961 3466 977 3468
rect 735 3454 750 3458
rect 653 3452 750 3454
rect 778 3452 946 3464
rect 962 3454 977 3458
rect 995 3455 1034 3474
rect 1053 3468 1060 3469
rect 1059 3461 1060 3468
rect 1043 3458 1044 3461
rect 1059 3458 1072 3461
rect 995 3454 1025 3455
rect 1034 3454 1040 3455
rect 1043 3454 1072 3458
rect 962 3453 1072 3454
rect 962 3452 1078 3453
rect 637 3444 688 3452
rect 637 3432 662 3444
rect 669 3432 688 3444
rect 719 3444 769 3452
rect 719 3436 735 3444
rect 742 3442 769 3444
rect 778 3442 999 3452
rect 742 3432 999 3442
rect 1028 3444 1078 3452
rect 1028 3435 1044 3444
rect 637 3424 688 3432
rect 735 3424 999 3432
rect 1025 3432 1044 3435
rect 1051 3432 1078 3444
rect 1025 3424 1078 3432
rect 653 3416 654 3424
rect 669 3416 682 3424
rect 653 3408 669 3416
rect 650 3401 669 3404
rect 650 3392 672 3401
rect 623 3382 672 3392
rect 623 3376 653 3382
rect 672 3377 677 3382
rect 595 3360 669 3376
rect 687 3368 717 3424
rect 752 3414 960 3424
rect 995 3420 1040 3424
rect 1043 3423 1044 3424
rect 1059 3423 1072 3424
rect 778 3384 967 3414
rect 793 3381 967 3384
rect 786 3378 967 3381
rect 595 3358 608 3360
rect 623 3358 657 3360
rect 595 3342 669 3358
rect 696 3354 709 3368
rect 724 3354 740 3370
rect 786 3365 797 3378
rect 579 3320 580 3336
rect 595 3320 608 3342
rect 623 3320 653 3342
rect 696 3338 758 3354
rect 786 3347 797 3363
rect 802 3358 812 3378
rect 822 3358 836 3378
rect 839 3365 848 3378
rect 864 3365 873 3378
rect 802 3347 836 3358
rect 839 3347 848 3363
rect 864 3347 873 3363
rect 880 3358 890 3378
rect 900 3358 914 3378
rect 915 3365 926 3378
rect 880 3347 914 3358
rect 915 3347 926 3363
rect 972 3354 988 3370
rect 995 3368 1025 3420
rect 1059 3416 1060 3423
rect 1044 3408 1060 3416
rect 1031 3376 1044 3395
rect 1059 3376 1089 3392
rect 1031 3360 1105 3376
rect 1031 3358 1044 3360
rect 1059 3358 1093 3360
rect 696 3336 709 3338
rect 724 3336 758 3338
rect 696 3320 758 3336
rect 802 3331 818 3334
rect 880 3331 910 3342
rect 958 3338 1004 3354
rect 1031 3342 1105 3358
rect 958 3336 992 3338
rect 957 3320 1004 3336
rect 1031 3320 1044 3342
rect 1059 3320 1089 3342
rect 1116 3320 1117 3336
rect 1132 3320 1145 3480
rect 1175 3376 1188 3480
rect 1233 3458 1234 3468
rect 1249 3458 1262 3468
rect 1233 3454 1262 3458
rect 1267 3454 1297 3480
rect 1315 3466 1331 3468
rect 1403 3466 1456 3480
rect 1404 3464 1468 3466
rect 1511 3464 1526 3480
rect 1575 3477 1605 3480
rect 1575 3474 1611 3477
rect 1541 3466 1557 3468
rect 1315 3454 1330 3458
rect 1233 3452 1330 3454
rect 1358 3452 1526 3464
rect 1542 3454 1557 3458
rect 1575 3455 1614 3474
rect 1633 3468 1640 3469
rect 1639 3461 1640 3468
rect 1623 3458 1624 3461
rect 1639 3458 1652 3461
rect 1575 3454 1605 3455
rect 1614 3454 1620 3455
rect 1623 3454 1652 3458
rect 1542 3453 1652 3454
rect 1542 3452 1658 3453
rect 1217 3444 1268 3452
rect 1217 3432 1242 3444
rect 1249 3432 1268 3444
rect 1299 3444 1349 3452
rect 1299 3436 1315 3444
rect 1322 3442 1349 3444
rect 1358 3442 1579 3452
rect 1322 3432 1579 3442
rect 1608 3444 1658 3452
rect 1608 3435 1624 3444
rect 1217 3424 1268 3432
rect 1315 3424 1579 3432
rect 1605 3432 1624 3435
rect 1631 3432 1658 3444
rect 1605 3424 1658 3432
rect 1233 3416 1234 3424
rect 1249 3416 1262 3424
rect 1233 3408 1249 3416
rect 1230 3401 1249 3404
rect 1230 3392 1252 3401
rect 1203 3382 1252 3392
rect 1203 3376 1233 3382
rect 1252 3377 1257 3382
rect 1175 3360 1249 3376
rect 1267 3368 1297 3424
rect 1332 3414 1540 3424
rect 1575 3420 1620 3424
rect 1623 3423 1624 3424
rect 1639 3423 1652 3424
rect 1358 3384 1547 3414
rect 1373 3381 1547 3384
rect 1366 3378 1547 3381
rect 1175 3358 1188 3360
rect 1203 3358 1237 3360
rect 1175 3342 1249 3358
rect 1276 3354 1289 3368
rect 1304 3354 1320 3370
rect 1366 3365 1377 3378
rect 1159 3320 1160 3336
rect 1175 3320 1188 3342
rect 1203 3320 1233 3342
rect 1276 3338 1338 3354
rect 1366 3347 1377 3363
rect 1382 3358 1392 3378
rect 1402 3358 1416 3378
rect 1419 3365 1428 3378
rect 1444 3365 1453 3378
rect 1382 3347 1416 3358
rect 1419 3347 1428 3363
rect 1444 3347 1453 3363
rect 1460 3358 1470 3378
rect 1480 3358 1494 3378
rect 1495 3365 1506 3378
rect 1460 3347 1494 3358
rect 1495 3347 1506 3363
rect 1552 3354 1568 3370
rect 1575 3368 1605 3420
rect 1639 3416 1640 3423
rect 1624 3408 1640 3416
rect 1611 3376 1624 3395
rect 1639 3376 1669 3392
rect 1611 3360 1685 3376
rect 1611 3358 1624 3360
rect 1639 3358 1673 3360
rect 1276 3336 1289 3338
rect 1304 3336 1338 3338
rect 1276 3320 1338 3336
rect 1382 3331 1398 3334
rect 1460 3331 1490 3342
rect 1538 3338 1584 3354
rect 1611 3342 1685 3358
rect 1538 3336 1572 3338
rect 1537 3320 1584 3336
rect 1611 3320 1624 3342
rect 1639 3320 1669 3342
rect 1696 3320 1697 3336
rect 1712 3320 1725 3480
rect 1755 3376 1768 3480
rect 1813 3458 1814 3468
rect 1829 3458 1842 3468
rect 1813 3454 1842 3458
rect 1847 3454 1877 3480
rect 1895 3466 1911 3468
rect 1983 3466 2036 3480
rect 1984 3464 2048 3466
rect 2091 3464 2106 3480
rect 2155 3477 2185 3480
rect 2155 3474 2191 3477
rect 2121 3466 2137 3468
rect 1895 3454 1910 3458
rect 1813 3452 1910 3454
rect 1938 3452 2106 3464
rect 2122 3454 2137 3458
rect 2155 3455 2194 3474
rect 2213 3468 2220 3469
rect 2219 3461 2220 3468
rect 2203 3458 2204 3461
rect 2219 3458 2232 3461
rect 2155 3454 2185 3455
rect 2194 3454 2200 3455
rect 2203 3454 2232 3458
rect 2122 3453 2232 3454
rect 2122 3452 2238 3453
rect 1797 3444 1848 3452
rect 1797 3432 1822 3444
rect 1829 3432 1848 3444
rect 1879 3444 1929 3452
rect 1879 3436 1895 3444
rect 1902 3442 1929 3444
rect 1938 3442 2159 3452
rect 1902 3432 2159 3442
rect 2188 3444 2238 3452
rect 2188 3435 2204 3444
rect 1797 3424 1848 3432
rect 1895 3424 2159 3432
rect 2185 3432 2204 3435
rect 2211 3432 2238 3444
rect 2185 3424 2238 3432
rect 1813 3416 1814 3424
rect 1829 3416 1842 3424
rect 1813 3408 1829 3416
rect 1810 3401 1829 3404
rect 1810 3392 1832 3401
rect 1783 3382 1832 3392
rect 1783 3376 1813 3382
rect 1832 3377 1837 3382
rect 1755 3360 1829 3376
rect 1847 3368 1877 3424
rect 1912 3414 2120 3424
rect 2155 3420 2200 3424
rect 2203 3423 2204 3424
rect 2219 3423 2232 3424
rect 1938 3384 2127 3414
rect 1953 3381 2127 3384
rect 1946 3378 2127 3381
rect 1755 3358 1768 3360
rect 1783 3358 1817 3360
rect 1755 3342 1829 3358
rect 1856 3354 1869 3368
rect 1884 3354 1900 3370
rect 1946 3365 1957 3378
rect 1739 3320 1740 3336
rect 1755 3320 1768 3342
rect 1783 3320 1813 3342
rect 1856 3338 1918 3354
rect 1946 3347 1957 3363
rect 1962 3358 1972 3378
rect 1982 3358 1996 3378
rect 1999 3365 2008 3378
rect 2024 3365 2033 3378
rect 1962 3347 1996 3358
rect 1999 3347 2008 3363
rect 2024 3347 2033 3363
rect 2040 3358 2050 3378
rect 2060 3358 2074 3378
rect 2075 3365 2086 3378
rect 2040 3347 2074 3358
rect 2075 3347 2086 3363
rect 2132 3354 2148 3370
rect 2155 3368 2185 3420
rect 2219 3416 2220 3423
rect 2204 3408 2220 3416
rect 2191 3376 2204 3395
rect 2219 3376 2249 3392
rect 2191 3360 2265 3376
rect 2191 3358 2204 3360
rect 2219 3358 2253 3360
rect 1856 3336 1869 3338
rect 1884 3336 1918 3338
rect 1856 3320 1918 3336
rect 1962 3331 1978 3334
rect 2040 3331 2070 3342
rect 2118 3338 2164 3354
rect 2191 3342 2265 3358
rect 2118 3336 2152 3338
rect 2117 3320 2164 3336
rect 2191 3320 2204 3342
rect 2219 3320 2249 3342
rect 2276 3320 2277 3336
rect 2292 3320 2305 3480
rect 2335 3376 2348 3480
rect 2393 3458 2394 3468
rect 2409 3458 2422 3468
rect 2393 3454 2422 3458
rect 2427 3454 2457 3480
rect 2475 3466 2491 3468
rect 2563 3466 2616 3480
rect 2564 3464 2628 3466
rect 2671 3464 2686 3480
rect 2735 3477 2765 3480
rect 2735 3474 2771 3477
rect 2701 3466 2717 3468
rect 2475 3454 2490 3458
rect 2393 3452 2490 3454
rect 2518 3452 2686 3464
rect 2702 3454 2717 3458
rect 2735 3455 2774 3474
rect 2793 3468 2800 3469
rect 2799 3461 2800 3468
rect 2783 3458 2784 3461
rect 2799 3458 2812 3461
rect 2735 3454 2765 3455
rect 2774 3454 2780 3455
rect 2783 3454 2812 3458
rect 2702 3453 2812 3454
rect 2702 3452 2818 3453
rect 2377 3444 2428 3452
rect 2377 3432 2402 3444
rect 2409 3432 2428 3444
rect 2459 3444 2509 3452
rect 2459 3436 2475 3444
rect 2482 3442 2509 3444
rect 2518 3442 2739 3452
rect 2482 3432 2739 3442
rect 2768 3444 2818 3452
rect 2768 3435 2784 3444
rect 2377 3424 2428 3432
rect 2475 3424 2739 3432
rect 2765 3432 2784 3435
rect 2791 3432 2818 3444
rect 2765 3424 2818 3432
rect 2393 3416 2394 3424
rect 2409 3416 2422 3424
rect 2393 3408 2409 3416
rect 2390 3401 2409 3404
rect 2390 3392 2412 3401
rect 2363 3382 2412 3392
rect 2363 3376 2393 3382
rect 2412 3377 2417 3382
rect 2335 3360 2409 3376
rect 2427 3368 2457 3424
rect 2492 3414 2700 3424
rect 2735 3420 2780 3424
rect 2783 3423 2784 3424
rect 2799 3423 2812 3424
rect 2518 3384 2707 3414
rect 2533 3381 2707 3384
rect 2526 3378 2707 3381
rect 2335 3358 2348 3360
rect 2363 3358 2397 3360
rect 2335 3342 2409 3358
rect 2436 3354 2449 3368
rect 2464 3354 2480 3370
rect 2526 3365 2537 3378
rect 2319 3320 2320 3336
rect 2335 3320 2348 3342
rect 2363 3320 2393 3342
rect 2436 3338 2498 3354
rect 2526 3347 2537 3363
rect 2542 3358 2552 3378
rect 2562 3358 2576 3378
rect 2579 3365 2588 3378
rect 2604 3365 2613 3378
rect 2542 3347 2576 3358
rect 2579 3347 2588 3363
rect 2604 3347 2613 3363
rect 2620 3358 2630 3378
rect 2640 3358 2654 3378
rect 2655 3365 2666 3378
rect 2620 3347 2654 3358
rect 2655 3347 2666 3363
rect 2712 3354 2728 3370
rect 2735 3368 2765 3420
rect 2799 3416 2800 3423
rect 2784 3408 2800 3416
rect 2771 3376 2784 3395
rect 2799 3376 2829 3392
rect 2771 3360 2845 3376
rect 2771 3358 2784 3360
rect 2799 3358 2833 3360
rect 2436 3336 2449 3338
rect 2464 3336 2498 3338
rect 2436 3320 2498 3336
rect 2542 3331 2558 3334
rect 2620 3331 2650 3342
rect 2698 3338 2744 3354
rect 2771 3342 2845 3358
rect 2698 3336 2732 3338
rect 2697 3320 2744 3336
rect 2771 3320 2784 3342
rect 2799 3320 2829 3342
rect 2856 3320 2857 3336
rect 2872 3320 2885 3480
rect 2915 3376 2928 3480
rect 2973 3458 2974 3468
rect 2989 3458 3002 3468
rect 2973 3454 3002 3458
rect 3007 3454 3037 3480
rect 3055 3466 3071 3468
rect 3143 3466 3196 3480
rect 3144 3464 3208 3466
rect 3251 3464 3266 3480
rect 3315 3477 3345 3480
rect 3315 3474 3351 3477
rect 3281 3466 3297 3468
rect 3055 3454 3070 3458
rect 2973 3452 3070 3454
rect 3098 3452 3266 3464
rect 3282 3454 3297 3458
rect 3315 3455 3354 3474
rect 3373 3468 3380 3469
rect 3379 3461 3380 3468
rect 3363 3458 3364 3461
rect 3379 3458 3392 3461
rect 3315 3454 3345 3455
rect 3354 3454 3360 3455
rect 3363 3454 3392 3458
rect 3282 3453 3392 3454
rect 3282 3452 3398 3453
rect 2957 3444 3008 3452
rect 2957 3432 2982 3444
rect 2989 3432 3008 3444
rect 3039 3444 3089 3452
rect 3039 3436 3055 3444
rect 3062 3442 3089 3444
rect 3098 3442 3319 3452
rect 3062 3432 3319 3442
rect 3348 3444 3398 3452
rect 3348 3435 3364 3444
rect 2957 3424 3008 3432
rect 3055 3424 3319 3432
rect 3345 3432 3364 3435
rect 3371 3432 3398 3444
rect 3345 3424 3398 3432
rect 2973 3416 2974 3424
rect 2989 3416 3002 3424
rect 2973 3408 2989 3416
rect 2970 3401 2989 3404
rect 2970 3392 2992 3401
rect 2943 3382 2992 3392
rect 2943 3376 2973 3382
rect 2992 3377 2997 3382
rect 2915 3360 2989 3376
rect 3007 3368 3037 3424
rect 3072 3414 3280 3424
rect 3315 3420 3360 3424
rect 3363 3423 3364 3424
rect 3379 3423 3392 3424
rect 3098 3384 3287 3414
rect 3113 3381 3287 3384
rect 3106 3378 3287 3381
rect 2915 3358 2928 3360
rect 2943 3358 2977 3360
rect 2915 3342 2989 3358
rect 3016 3354 3029 3368
rect 3044 3354 3060 3370
rect 3106 3365 3117 3378
rect 2899 3320 2900 3336
rect 2915 3320 2928 3342
rect 2943 3320 2973 3342
rect 3016 3338 3078 3354
rect 3106 3347 3117 3363
rect 3122 3358 3132 3378
rect 3142 3358 3156 3378
rect 3159 3365 3168 3378
rect 3184 3365 3193 3378
rect 3122 3347 3156 3358
rect 3159 3347 3168 3363
rect 3184 3347 3193 3363
rect 3200 3358 3210 3378
rect 3220 3358 3234 3378
rect 3235 3365 3246 3378
rect 3200 3347 3234 3358
rect 3235 3347 3246 3363
rect 3292 3354 3308 3370
rect 3315 3368 3345 3420
rect 3379 3416 3380 3423
rect 3364 3408 3380 3416
rect 3351 3376 3364 3395
rect 3379 3376 3409 3392
rect 3351 3360 3425 3376
rect 3351 3358 3364 3360
rect 3379 3358 3413 3360
rect 3016 3336 3029 3338
rect 3044 3336 3078 3338
rect 3016 3320 3078 3336
rect 3122 3331 3138 3334
rect 3200 3331 3230 3342
rect 3278 3338 3324 3354
rect 3351 3342 3425 3358
rect 3278 3336 3312 3338
rect 3277 3320 3324 3336
rect 3351 3320 3364 3342
rect 3379 3320 3409 3342
rect 3436 3320 3437 3336
rect 3452 3320 3465 3480
rect 3495 3376 3508 3480
rect 3553 3458 3554 3468
rect 3569 3458 3582 3468
rect 3553 3454 3582 3458
rect 3587 3454 3617 3480
rect 3635 3466 3651 3468
rect 3723 3466 3776 3480
rect 3724 3464 3788 3466
rect 3831 3464 3846 3480
rect 3895 3477 3925 3480
rect 3895 3474 3931 3477
rect 3861 3466 3877 3468
rect 3635 3454 3650 3458
rect 3553 3452 3650 3454
rect 3678 3452 3846 3464
rect 3862 3454 3877 3458
rect 3895 3455 3934 3474
rect 3953 3468 3960 3469
rect 3959 3461 3960 3468
rect 3943 3458 3944 3461
rect 3959 3458 3972 3461
rect 3895 3454 3925 3455
rect 3934 3454 3940 3455
rect 3943 3454 3972 3458
rect 3862 3453 3972 3454
rect 3862 3452 3978 3453
rect 3537 3444 3588 3452
rect 3537 3432 3562 3444
rect 3569 3432 3588 3444
rect 3619 3444 3669 3452
rect 3619 3436 3635 3444
rect 3642 3442 3669 3444
rect 3678 3442 3899 3452
rect 3642 3432 3899 3442
rect 3928 3444 3978 3452
rect 3928 3435 3944 3444
rect 3537 3424 3588 3432
rect 3635 3424 3899 3432
rect 3925 3432 3944 3435
rect 3951 3432 3978 3444
rect 3925 3424 3978 3432
rect 3553 3416 3554 3424
rect 3569 3416 3582 3424
rect 3553 3408 3569 3416
rect 3550 3401 3569 3404
rect 3550 3392 3572 3401
rect 3523 3382 3572 3392
rect 3523 3376 3553 3382
rect 3572 3377 3577 3382
rect 3495 3360 3569 3376
rect 3587 3368 3617 3424
rect 3652 3414 3860 3424
rect 3895 3420 3940 3424
rect 3943 3423 3944 3424
rect 3959 3423 3972 3424
rect 3678 3384 3867 3414
rect 3693 3381 3867 3384
rect 3686 3378 3867 3381
rect 3495 3358 3508 3360
rect 3523 3358 3557 3360
rect 3495 3342 3569 3358
rect 3596 3354 3609 3368
rect 3624 3354 3640 3370
rect 3686 3365 3697 3378
rect 3479 3320 3480 3336
rect 3495 3320 3508 3342
rect 3523 3320 3553 3342
rect 3596 3338 3658 3354
rect 3686 3347 3697 3363
rect 3702 3358 3712 3378
rect 3722 3358 3736 3378
rect 3739 3365 3748 3378
rect 3764 3365 3773 3378
rect 3702 3347 3736 3358
rect 3739 3347 3748 3363
rect 3764 3347 3773 3363
rect 3780 3358 3790 3378
rect 3800 3358 3814 3378
rect 3815 3365 3826 3378
rect 3780 3347 3814 3358
rect 3815 3347 3826 3363
rect 3872 3354 3888 3370
rect 3895 3368 3925 3420
rect 3959 3416 3960 3423
rect 3944 3408 3960 3416
rect 3931 3376 3944 3395
rect 3959 3376 3989 3392
rect 3931 3360 4005 3376
rect 3931 3358 3944 3360
rect 3959 3358 3993 3360
rect 3596 3336 3609 3338
rect 3624 3336 3658 3338
rect 3596 3320 3658 3336
rect 3702 3331 3718 3334
rect 3780 3331 3810 3342
rect 3858 3338 3904 3354
rect 3931 3342 4005 3358
rect 3858 3336 3892 3338
rect 3857 3320 3904 3336
rect 3931 3320 3944 3342
rect 3959 3320 3989 3342
rect 4016 3320 4017 3336
rect 4032 3320 4045 3480
rect 4075 3376 4088 3480
rect 4133 3458 4134 3468
rect 4149 3458 4162 3468
rect 4133 3454 4162 3458
rect 4167 3454 4197 3480
rect 4215 3466 4231 3468
rect 4303 3466 4356 3480
rect 4304 3464 4368 3466
rect 4411 3464 4426 3480
rect 4475 3477 4505 3480
rect 4475 3474 4511 3477
rect 4441 3466 4457 3468
rect 4215 3454 4230 3458
rect 4133 3452 4230 3454
rect 4258 3452 4426 3464
rect 4442 3454 4457 3458
rect 4475 3455 4514 3474
rect 4533 3468 4540 3469
rect 4539 3461 4540 3468
rect 4523 3458 4524 3461
rect 4539 3458 4552 3461
rect 4475 3454 4505 3455
rect 4514 3454 4520 3455
rect 4523 3454 4552 3458
rect 4442 3453 4552 3454
rect 4442 3452 4558 3453
rect 4117 3444 4168 3452
rect 4117 3432 4142 3444
rect 4149 3432 4168 3444
rect 4199 3444 4249 3452
rect 4199 3436 4215 3444
rect 4222 3442 4249 3444
rect 4258 3442 4479 3452
rect 4222 3432 4479 3442
rect 4508 3444 4558 3452
rect 4508 3435 4524 3444
rect 4117 3424 4168 3432
rect 4215 3424 4479 3432
rect 4505 3432 4524 3435
rect 4531 3432 4558 3444
rect 4505 3424 4558 3432
rect 4133 3416 4134 3424
rect 4149 3416 4162 3424
rect 4133 3408 4149 3416
rect 4130 3401 4149 3404
rect 4130 3392 4152 3401
rect 4103 3382 4152 3392
rect 4103 3376 4133 3382
rect 4152 3377 4157 3382
rect 4075 3360 4149 3376
rect 4167 3368 4197 3424
rect 4232 3414 4440 3424
rect 4475 3420 4520 3424
rect 4523 3423 4524 3424
rect 4539 3423 4552 3424
rect 4258 3384 4447 3414
rect 4273 3381 4447 3384
rect 4266 3378 4447 3381
rect 4075 3358 4088 3360
rect 4103 3358 4137 3360
rect 4075 3342 4149 3358
rect 4176 3354 4189 3368
rect 4204 3354 4220 3370
rect 4266 3365 4277 3378
rect 4059 3320 4060 3336
rect 4075 3320 4088 3342
rect 4103 3320 4133 3342
rect 4176 3338 4238 3354
rect 4266 3347 4277 3363
rect 4282 3358 4292 3378
rect 4302 3358 4316 3378
rect 4319 3365 4328 3378
rect 4344 3365 4353 3378
rect 4282 3347 4316 3358
rect 4319 3347 4328 3363
rect 4344 3347 4353 3363
rect 4360 3358 4370 3378
rect 4380 3358 4394 3378
rect 4395 3365 4406 3378
rect 4360 3347 4394 3358
rect 4395 3347 4406 3363
rect 4452 3354 4468 3370
rect 4475 3368 4505 3420
rect 4539 3416 4540 3423
rect 4524 3408 4540 3416
rect 4511 3376 4524 3395
rect 4539 3376 4569 3392
rect 4511 3360 4585 3376
rect 4511 3358 4524 3360
rect 4539 3358 4573 3360
rect 4176 3336 4189 3338
rect 4204 3336 4238 3338
rect 4176 3320 4238 3336
rect 4282 3331 4298 3334
rect 4360 3331 4390 3342
rect 4438 3338 4484 3354
rect 4511 3342 4585 3358
rect 4438 3336 4472 3338
rect 4437 3320 4484 3336
rect 4511 3320 4524 3342
rect 4539 3320 4569 3342
rect 4596 3320 4597 3336
rect 4612 3320 4625 3480
rect -7 3312 34 3320
rect -7 3286 8 3312
rect 15 3286 34 3312
rect 98 3308 160 3320
rect 172 3308 247 3320
rect 305 3308 380 3320
rect 392 3308 423 3320
rect 429 3308 464 3320
rect 98 3306 260 3308
rect -7 3278 34 3286
rect 116 3282 129 3306
rect 144 3304 159 3306
rect -1 3268 0 3278
rect 15 3268 28 3278
rect 43 3268 73 3282
rect 116 3268 159 3282
rect 183 3279 190 3286
rect 193 3282 260 3306
rect 292 3306 464 3308
rect 262 3284 290 3288
rect 292 3284 372 3306
rect 393 3304 408 3306
rect 262 3282 372 3284
rect 193 3278 372 3282
rect 166 3268 196 3278
rect 198 3268 351 3278
rect 359 3268 389 3278
rect 393 3268 423 3282
rect 451 3268 464 3306
rect 536 3312 571 3320
rect 536 3286 537 3312
rect 544 3286 571 3312
rect 479 3268 509 3282
rect 536 3278 571 3286
rect 573 3312 614 3320
rect 573 3286 588 3312
rect 595 3286 614 3312
rect 678 3308 740 3320
rect 752 3308 827 3320
rect 885 3308 960 3320
rect 972 3308 1003 3320
rect 1009 3308 1044 3320
rect 678 3306 840 3308
rect 573 3278 614 3286
rect 696 3282 709 3306
rect 724 3304 739 3306
rect 536 3268 537 3278
rect 552 3268 565 3278
rect 579 3268 580 3278
rect 595 3268 608 3278
rect 623 3268 653 3282
rect 696 3268 739 3282
rect 763 3279 770 3286
rect 773 3282 840 3306
rect 872 3306 1044 3308
rect 842 3284 870 3288
rect 872 3284 952 3306
rect 973 3304 988 3306
rect 842 3282 952 3284
rect 773 3278 952 3282
rect 746 3268 776 3278
rect 778 3268 931 3278
rect 939 3268 969 3278
rect 973 3268 1003 3282
rect 1031 3268 1044 3306
rect 1116 3312 1151 3320
rect 1116 3286 1117 3312
rect 1124 3286 1151 3312
rect 1059 3268 1089 3282
rect 1116 3278 1151 3286
rect 1153 3312 1194 3320
rect 1153 3286 1168 3312
rect 1175 3286 1194 3312
rect 1258 3308 1320 3320
rect 1332 3308 1407 3320
rect 1465 3308 1540 3320
rect 1552 3308 1583 3320
rect 1589 3308 1624 3320
rect 1258 3306 1420 3308
rect 1153 3278 1194 3286
rect 1276 3282 1289 3306
rect 1304 3304 1319 3306
rect 1116 3268 1117 3278
rect 1132 3268 1145 3278
rect 1159 3268 1160 3278
rect 1175 3268 1188 3278
rect 1203 3268 1233 3282
rect 1276 3268 1319 3282
rect 1343 3279 1350 3286
rect 1353 3282 1420 3306
rect 1452 3306 1624 3308
rect 1422 3284 1450 3288
rect 1452 3284 1532 3306
rect 1553 3304 1568 3306
rect 1422 3282 1532 3284
rect 1353 3278 1532 3282
rect 1326 3268 1356 3278
rect 1358 3268 1511 3278
rect 1519 3268 1549 3278
rect 1553 3268 1583 3282
rect 1611 3268 1624 3306
rect 1696 3312 1731 3320
rect 1696 3286 1697 3312
rect 1704 3286 1731 3312
rect 1639 3268 1669 3282
rect 1696 3278 1731 3286
rect 1733 3312 1774 3320
rect 1733 3286 1748 3312
rect 1755 3286 1774 3312
rect 1838 3308 1900 3320
rect 1912 3308 1987 3320
rect 2045 3308 2120 3320
rect 2132 3308 2163 3320
rect 2169 3308 2204 3320
rect 1838 3306 2000 3308
rect 1733 3278 1774 3286
rect 1856 3282 1869 3306
rect 1884 3304 1899 3306
rect 1696 3268 1697 3278
rect 1712 3268 1725 3278
rect 1739 3268 1740 3278
rect 1755 3268 1768 3278
rect 1783 3268 1813 3282
rect 1856 3268 1899 3282
rect 1923 3279 1930 3286
rect 1933 3282 2000 3306
rect 2032 3306 2204 3308
rect 2002 3284 2030 3288
rect 2032 3284 2112 3306
rect 2133 3304 2148 3306
rect 2002 3282 2112 3284
rect 1933 3278 2112 3282
rect 1906 3268 1936 3278
rect 1938 3268 2091 3278
rect 2099 3268 2129 3278
rect 2133 3268 2163 3282
rect 2191 3268 2204 3306
rect 2276 3312 2311 3320
rect 2276 3286 2277 3312
rect 2284 3286 2311 3312
rect 2219 3268 2249 3282
rect 2276 3278 2311 3286
rect 2313 3312 2354 3320
rect 2313 3286 2328 3312
rect 2335 3286 2354 3312
rect 2418 3308 2480 3320
rect 2492 3308 2567 3320
rect 2625 3308 2700 3320
rect 2712 3308 2743 3320
rect 2749 3308 2784 3320
rect 2418 3306 2580 3308
rect 2313 3278 2354 3286
rect 2436 3282 2449 3306
rect 2464 3304 2479 3306
rect 2276 3268 2277 3278
rect 2292 3268 2305 3278
rect 2319 3268 2320 3278
rect 2335 3268 2348 3278
rect 2363 3268 2393 3282
rect 2436 3268 2479 3282
rect 2503 3279 2510 3286
rect 2513 3282 2580 3306
rect 2612 3306 2784 3308
rect 2582 3284 2610 3288
rect 2612 3284 2692 3306
rect 2713 3304 2728 3306
rect 2582 3282 2692 3284
rect 2513 3278 2692 3282
rect 2486 3268 2516 3278
rect 2518 3268 2671 3278
rect 2679 3268 2709 3278
rect 2713 3268 2743 3282
rect 2771 3268 2784 3306
rect 2856 3312 2891 3320
rect 2856 3286 2857 3312
rect 2864 3286 2891 3312
rect 2799 3268 2829 3282
rect 2856 3278 2891 3286
rect 2893 3312 2934 3320
rect 2893 3286 2908 3312
rect 2915 3286 2934 3312
rect 2998 3308 3060 3320
rect 3072 3308 3147 3320
rect 3205 3308 3280 3320
rect 3292 3308 3323 3320
rect 3329 3308 3364 3320
rect 2998 3306 3160 3308
rect 2893 3278 2934 3286
rect 3016 3282 3029 3306
rect 3044 3304 3059 3306
rect 2856 3268 2857 3278
rect 2872 3268 2885 3278
rect 2899 3268 2900 3278
rect 2915 3268 2928 3278
rect 2943 3268 2973 3282
rect 3016 3268 3059 3282
rect 3083 3279 3090 3286
rect 3093 3282 3160 3306
rect 3192 3306 3364 3308
rect 3162 3284 3190 3288
rect 3192 3284 3272 3306
rect 3293 3304 3308 3306
rect 3162 3282 3272 3284
rect 3093 3278 3272 3282
rect 3066 3268 3096 3278
rect 3098 3268 3251 3278
rect 3259 3268 3289 3278
rect 3293 3268 3323 3282
rect 3351 3268 3364 3306
rect 3436 3312 3471 3320
rect 3436 3286 3437 3312
rect 3444 3286 3471 3312
rect 3379 3268 3409 3282
rect 3436 3278 3471 3286
rect 3473 3312 3514 3320
rect 3473 3286 3488 3312
rect 3495 3286 3514 3312
rect 3578 3308 3640 3320
rect 3652 3308 3727 3320
rect 3785 3308 3860 3320
rect 3872 3308 3903 3320
rect 3909 3308 3944 3320
rect 3578 3306 3740 3308
rect 3473 3278 3514 3286
rect 3596 3282 3609 3306
rect 3624 3304 3639 3306
rect 3436 3268 3437 3278
rect 3452 3268 3465 3278
rect 3479 3268 3480 3278
rect 3495 3268 3508 3278
rect 3523 3268 3553 3282
rect 3596 3268 3639 3282
rect 3663 3279 3670 3286
rect 3673 3282 3740 3306
rect 3772 3306 3944 3308
rect 3742 3284 3770 3288
rect 3772 3284 3852 3306
rect 3873 3304 3888 3306
rect 3742 3282 3852 3284
rect 3673 3278 3852 3282
rect 3646 3268 3676 3278
rect 3678 3268 3831 3278
rect 3839 3268 3869 3278
rect 3873 3268 3903 3282
rect 3931 3268 3944 3306
rect 4016 3312 4051 3320
rect 4016 3286 4017 3312
rect 4024 3286 4051 3312
rect 3959 3268 3989 3282
rect 4016 3278 4051 3286
rect 4053 3312 4094 3320
rect 4053 3286 4068 3312
rect 4075 3286 4094 3312
rect 4158 3308 4220 3320
rect 4232 3308 4307 3320
rect 4365 3308 4440 3320
rect 4452 3308 4483 3320
rect 4489 3308 4524 3320
rect 4158 3306 4320 3308
rect 4053 3278 4094 3286
rect 4176 3282 4189 3306
rect 4204 3304 4219 3306
rect 4016 3268 4017 3278
rect 4032 3268 4045 3278
rect 4059 3268 4060 3278
rect 4075 3268 4088 3278
rect 4103 3268 4133 3282
rect 4176 3268 4219 3282
rect 4243 3279 4250 3286
rect 4253 3282 4320 3306
rect 4352 3306 4524 3308
rect 4322 3284 4350 3288
rect 4352 3284 4432 3306
rect 4453 3304 4468 3306
rect 4322 3282 4432 3284
rect 4253 3278 4432 3282
rect 4226 3268 4256 3278
rect 4258 3268 4411 3278
rect 4419 3268 4449 3278
rect 4453 3268 4483 3282
rect 4511 3268 4524 3306
rect 4596 3312 4631 3320
rect 4596 3286 4597 3312
rect 4604 3286 4631 3312
rect 4539 3268 4569 3282
rect 4596 3278 4631 3286
rect 4596 3268 4597 3278
rect 4612 3268 4625 3278
rect -1 3262 4625 3268
rect 0 3254 4625 3262
rect 15 3224 28 3254
rect 43 3236 73 3254
rect 116 3240 130 3254
rect 166 3240 386 3254
rect 117 3238 130 3240
rect 83 3226 98 3238
rect 80 3224 102 3226
rect 107 3224 137 3238
rect 198 3236 351 3240
rect 180 3224 372 3236
rect 415 3224 445 3238
rect 451 3224 464 3254
rect 479 3236 509 3254
rect 552 3224 565 3254
rect 595 3224 608 3254
rect 623 3236 653 3254
rect 696 3240 710 3254
rect 746 3240 966 3254
rect 697 3238 710 3240
rect 663 3226 678 3238
rect 660 3224 682 3226
rect 687 3224 717 3238
rect 778 3236 931 3240
rect 760 3224 952 3236
rect 995 3224 1025 3238
rect 1031 3224 1044 3254
rect 1059 3236 1089 3254
rect 1132 3224 1145 3254
rect 1175 3224 1188 3254
rect 1203 3236 1233 3254
rect 1276 3240 1290 3254
rect 1326 3240 1546 3254
rect 1277 3238 1290 3240
rect 1243 3226 1258 3238
rect 1240 3224 1262 3226
rect 1267 3224 1297 3238
rect 1358 3236 1511 3240
rect 1340 3224 1532 3236
rect 1575 3224 1605 3238
rect 1611 3224 1624 3254
rect 1639 3236 1669 3254
rect 1712 3224 1725 3254
rect 1755 3224 1768 3254
rect 1783 3236 1813 3254
rect 1856 3240 1870 3254
rect 1906 3240 2126 3254
rect 1857 3238 1870 3240
rect 1823 3226 1838 3238
rect 1820 3224 1842 3226
rect 1847 3224 1877 3238
rect 1938 3236 2091 3240
rect 1920 3224 2112 3236
rect 2155 3224 2185 3238
rect 2191 3224 2204 3254
rect 2219 3236 2249 3254
rect 2292 3224 2305 3254
rect 2335 3224 2348 3254
rect 2363 3236 2393 3254
rect 2436 3240 2450 3254
rect 2486 3240 2706 3254
rect 2437 3238 2450 3240
rect 2403 3226 2418 3238
rect 2400 3224 2422 3226
rect 2427 3224 2457 3238
rect 2518 3236 2671 3240
rect 2500 3224 2692 3236
rect 2735 3224 2765 3238
rect 2771 3224 2784 3254
rect 2799 3236 2829 3254
rect 2872 3224 2885 3254
rect 2915 3224 2928 3254
rect 2943 3236 2973 3254
rect 3016 3240 3030 3254
rect 3066 3240 3286 3254
rect 3017 3238 3030 3240
rect 2983 3226 2998 3238
rect 2980 3224 3002 3226
rect 3007 3224 3037 3238
rect 3098 3236 3251 3240
rect 3080 3224 3272 3236
rect 3315 3224 3345 3238
rect 3351 3224 3364 3254
rect 3379 3236 3409 3254
rect 3452 3224 3465 3254
rect 3495 3224 3508 3254
rect 3523 3236 3553 3254
rect 3596 3240 3610 3254
rect 3646 3240 3866 3254
rect 3597 3238 3610 3240
rect 3563 3226 3578 3238
rect 3560 3224 3582 3226
rect 3587 3224 3617 3238
rect 3678 3236 3831 3240
rect 3660 3224 3852 3236
rect 3895 3224 3925 3238
rect 3931 3224 3944 3254
rect 3959 3236 3989 3254
rect 4032 3224 4045 3254
rect 4075 3224 4088 3254
rect 4103 3236 4133 3254
rect 4176 3240 4190 3254
rect 4226 3240 4446 3254
rect 4177 3238 4190 3240
rect 4143 3226 4158 3238
rect 4140 3224 4162 3226
rect 4167 3224 4197 3238
rect 4258 3236 4411 3240
rect 4240 3224 4432 3236
rect 4475 3224 4505 3238
rect 4511 3224 4524 3254
rect 4539 3236 4569 3254
rect 4612 3224 4625 3254
rect 0 3210 4625 3224
rect 15 3106 28 3210
rect 73 3188 74 3198
rect 89 3188 102 3198
rect 73 3184 102 3188
rect 107 3184 137 3210
rect 155 3196 171 3198
rect 243 3196 296 3210
rect 244 3194 308 3196
rect 351 3194 366 3210
rect 415 3207 445 3210
rect 415 3204 451 3207
rect 381 3196 397 3198
rect 155 3184 170 3188
rect 73 3182 170 3184
rect 198 3182 366 3194
rect 382 3184 397 3188
rect 415 3185 454 3204
rect 473 3198 480 3199
rect 479 3191 480 3198
rect 463 3188 464 3191
rect 479 3188 492 3191
rect 415 3184 445 3185
rect 454 3184 460 3185
rect 463 3184 492 3188
rect 382 3183 492 3184
rect 382 3182 498 3183
rect 57 3174 108 3182
rect 57 3162 82 3174
rect 89 3162 108 3174
rect 139 3174 189 3182
rect 139 3166 155 3174
rect 162 3172 189 3174
rect 198 3172 419 3182
rect 162 3162 419 3172
rect 448 3174 498 3182
rect 448 3165 464 3174
rect 57 3154 108 3162
rect 155 3154 419 3162
rect 445 3162 464 3165
rect 471 3162 498 3174
rect 445 3154 498 3162
rect 73 3146 74 3154
rect 89 3146 102 3154
rect 73 3138 89 3146
rect 70 3131 89 3134
rect 70 3122 92 3131
rect 43 3112 92 3122
rect 43 3106 73 3112
rect 92 3107 97 3112
rect 15 3090 89 3106
rect 107 3098 137 3154
rect 172 3144 380 3154
rect 415 3150 460 3154
rect 463 3153 464 3154
rect 479 3153 492 3154
rect 198 3114 387 3144
rect 213 3111 387 3114
rect 206 3108 387 3111
rect 15 3088 28 3090
rect 43 3088 77 3090
rect 15 3072 89 3088
rect 116 3084 129 3098
rect 144 3084 160 3100
rect 206 3095 217 3108
rect -1 3050 0 3066
rect 15 3050 28 3072
rect 43 3050 73 3072
rect 116 3068 178 3084
rect 206 3077 217 3093
rect 222 3088 232 3108
rect 242 3088 256 3108
rect 259 3095 268 3108
rect 284 3095 293 3108
rect 222 3077 256 3088
rect 259 3077 268 3093
rect 284 3077 293 3093
rect 300 3088 310 3108
rect 320 3088 334 3108
rect 335 3095 346 3108
rect 300 3077 334 3088
rect 335 3077 346 3093
rect 392 3084 408 3100
rect 415 3098 445 3150
rect 479 3146 480 3153
rect 464 3138 480 3146
rect 451 3106 464 3125
rect 479 3106 509 3122
rect 451 3090 525 3106
rect 451 3088 464 3090
rect 479 3088 513 3090
rect 116 3066 129 3068
rect 144 3066 178 3068
rect 116 3050 178 3066
rect 222 3061 238 3064
rect 300 3061 330 3072
rect 378 3068 424 3084
rect 451 3072 525 3088
rect 378 3066 412 3068
rect 377 3050 424 3066
rect 451 3050 464 3072
rect 479 3050 509 3072
rect 536 3050 537 3066
rect 552 3050 565 3210
rect 595 3106 608 3210
rect 653 3188 654 3198
rect 669 3188 682 3198
rect 653 3184 682 3188
rect 687 3184 717 3210
rect 735 3196 751 3198
rect 823 3196 876 3210
rect 824 3194 888 3196
rect 931 3194 946 3210
rect 995 3207 1025 3210
rect 995 3204 1031 3207
rect 961 3196 977 3198
rect 735 3184 750 3188
rect 653 3182 750 3184
rect 778 3182 946 3194
rect 962 3184 977 3188
rect 995 3185 1034 3204
rect 1053 3198 1060 3199
rect 1059 3191 1060 3198
rect 1043 3188 1044 3191
rect 1059 3188 1072 3191
rect 995 3184 1025 3185
rect 1034 3184 1040 3185
rect 1043 3184 1072 3188
rect 962 3183 1072 3184
rect 962 3182 1078 3183
rect 637 3174 688 3182
rect 637 3162 662 3174
rect 669 3162 688 3174
rect 719 3174 769 3182
rect 719 3166 735 3174
rect 742 3172 769 3174
rect 778 3172 999 3182
rect 742 3162 999 3172
rect 1028 3174 1078 3182
rect 1028 3165 1044 3174
rect 637 3154 688 3162
rect 735 3154 999 3162
rect 1025 3162 1044 3165
rect 1051 3162 1078 3174
rect 1025 3154 1078 3162
rect 653 3146 654 3154
rect 669 3146 682 3154
rect 653 3138 669 3146
rect 650 3131 669 3134
rect 650 3122 672 3131
rect 623 3112 672 3122
rect 623 3106 653 3112
rect 672 3107 677 3112
rect 595 3090 669 3106
rect 687 3098 717 3154
rect 752 3144 960 3154
rect 995 3150 1040 3154
rect 1043 3153 1044 3154
rect 1059 3153 1072 3154
rect 778 3114 967 3144
rect 793 3111 967 3114
rect 786 3108 967 3111
rect 595 3088 608 3090
rect 623 3088 657 3090
rect 595 3072 669 3088
rect 696 3084 709 3098
rect 724 3084 740 3100
rect 786 3095 797 3108
rect 579 3050 580 3066
rect 595 3050 608 3072
rect 623 3050 653 3072
rect 696 3068 758 3084
rect 786 3077 797 3093
rect 802 3088 812 3108
rect 822 3088 836 3108
rect 839 3095 848 3108
rect 864 3095 873 3108
rect 802 3077 836 3088
rect 839 3077 848 3093
rect 864 3077 873 3093
rect 880 3088 890 3108
rect 900 3088 914 3108
rect 915 3095 926 3108
rect 880 3077 914 3088
rect 915 3077 926 3093
rect 972 3084 988 3100
rect 995 3098 1025 3150
rect 1059 3146 1060 3153
rect 1044 3138 1060 3146
rect 1031 3106 1044 3125
rect 1059 3106 1089 3122
rect 1031 3090 1105 3106
rect 1031 3088 1044 3090
rect 1059 3088 1093 3090
rect 696 3066 709 3068
rect 724 3066 758 3068
rect 696 3050 758 3066
rect 802 3061 818 3064
rect 880 3061 910 3072
rect 958 3068 1004 3084
rect 1031 3072 1105 3088
rect 958 3066 992 3068
rect 957 3050 1004 3066
rect 1031 3050 1044 3072
rect 1059 3050 1089 3072
rect 1116 3050 1117 3066
rect 1132 3050 1145 3210
rect 1175 3106 1188 3210
rect 1233 3188 1234 3198
rect 1249 3188 1262 3198
rect 1233 3184 1262 3188
rect 1267 3184 1297 3210
rect 1315 3196 1331 3198
rect 1403 3196 1456 3210
rect 1404 3194 1468 3196
rect 1511 3194 1526 3210
rect 1575 3207 1605 3210
rect 1575 3204 1611 3207
rect 1541 3196 1557 3198
rect 1315 3184 1330 3188
rect 1233 3182 1330 3184
rect 1358 3182 1526 3194
rect 1542 3184 1557 3188
rect 1575 3185 1614 3204
rect 1633 3198 1640 3199
rect 1639 3191 1640 3198
rect 1623 3188 1624 3191
rect 1639 3188 1652 3191
rect 1575 3184 1605 3185
rect 1614 3184 1620 3185
rect 1623 3184 1652 3188
rect 1542 3183 1652 3184
rect 1542 3182 1658 3183
rect 1217 3174 1268 3182
rect 1217 3162 1242 3174
rect 1249 3162 1268 3174
rect 1299 3174 1349 3182
rect 1299 3166 1315 3174
rect 1322 3172 1349 3174
rect 1358 3172 1579 3182
rect 1322 3162 1579 3172
rect 1608 3174 1658 3182
rect 1608 3165 1624 3174
rect 1217 3154 1268 3162
rect 1315 3154 1579 3162
rect 1605 3162 1624 3165
rect 1631 3162 1658 3174
rect 1605 3154 1658 3162
rect 1233 3146 1234 3154
rect 1249 3146 1262 3154
rect 1233 3138 1249 3146
rect 1230 3131 1249 3134
rect 1230 3122 1252 3131
rect 1203 3112 1252 3122
rect 1203 3106 1233 3112
rect 1252 3107 1257 3112
rect 1175 3090 1249 3106
rect 1267 3098 1297 3154
rect 1332 3144 1540 3154
rect 1575 3150 1620 3154
rect 1623 3153 1624 3154
rect 1639 3153 1652 3154
rect 1358 3114 1547 3144
rect 1373 3111 1547 3114
rect 1366 3108 1547 3111
rect 1175 3088 1188 3090
rect 1203 3088 1237 3090
rect 1175 3072 1249 3088
rect 1276 3084 1289 3098
rect 1304 3084 1320 3100
rect 1366 3095 1377 3108
rect 1159 3050 1160 3066
rect 1175 3050 1188 3072
rect 1203 3050 1233 3072
rect 1276 3068 1338 3084
rect 1366 3077 1377 3093
rect 1382 3088 1392 3108
rect 1402 3088 1416 3108
rect 1419 3095 1428 3108
rect 1444 3095 1453 3108
rect 1382 3077 1416 3088
rect 1419 3077 1428 3093
rect 1444 3077 1453 3093
rect 1460 3088 1470 3108
rect 1480 3088 1494 3108
rect 1495 3095 1506 3108
rect 1460 3077 1494 3088
rect 1495 3077 1506 3093
rect 1552 3084 1568 3100
rect 1575 3098 1605 3150
rect 1639 3146 1640 3153
rect 1624 3138 1640 3146
rect 1611 3106 1624 3125
rect 1639 3106 1669 3122
rect 1611 3090 1685 3106
rect 1611 3088 1624 3090
rect 1639 3088 1673 3090
rect 1276 3066 1289 3068
rect 1304 3066 1338 3068
rect 1276 3050 1338 3066
rect 1382 3061 1398 3064
rect 1460 3061 1490 3072
rect 1538 3068 1584 3084
rect 1611 3072 1685 3088
rect 1538 3066 1572 3068
rect 1537 3050 1584 3066
rect 1611 3050 1624 3072
rect 1639 3050 1669 3072
rect 1696 3050 1697 3066
rect 1712 3050 1725 3210
rect 1755 3106 1768 3210
rect 1813 3188 1814 3198
rect 1829 3188 1842 3198
rect 1813 3184 1842 3188
rect 1847 3184 1877 3210
rect 1895 3196 1911 3198
rect 1983 3196 2036 3210
rect 1984 3194 2048 3196
rect 2091 3194 2106 3210
rect 2155 3207 2185 3210
rect 2155 3204 2191 3207
rect 2121 3196 2137 3198
rect 1895 3184 1910 3188
rect 1813 3182 1910 3184
rect 1938 3182 2106 3194
rect 2122 3184 2137 3188
rect 2155 3185 2194 3204
rect 2213 3198 2220 3199
rect 2219 3191 2220 3198
rect 2203 3188 2204 3191
rect 2219 3188 2232 3191
rect 2155 3184 2185 3185
rect 2194 3184 2200 3185
rect 2203 3184 2232 3188
rect 2122 3183 2232 3184
rect 2122 3182 2238 3183
rect 1797 3174 1848 3182
rect 1797 3162 1822 3174
rect 1829 3162 1848 3174
rect 1879 3174 1929 3182
rect 1879 3166 1895 3174
rect 1902 3172 1929 3174
rect 1938 3172 2159 3182
rect 1902 3162 2159 3172
rect 2188 3174 2238 3182
rect 2188 3165 2204 3174
rect 1797 3154 1848 3162
rect 1895 3154 2159 3162
rect 2185 3162 2204 3165
rect 2211 3162 2238 3174
rect 2185 3154 2238 3162
rect 1813 3146 1814 3154
rect 1829 3146 1842 3154
rect 1813 3138 1829 3146
rect 1810 3131 1829 3134
rect 1810 3122 1832 3131
rect 1783 3112 1832 3122
rect 1783 3106 1813 3112
rect 1832 3107 1837 3112
rect 1755 3090 1829 3106
rect 1847 3098 1877 3154
rect 1912 3144 2120 3154
rect 2155 3150 2200 3154
rect 2203 3153 2204 3154
rect 2219 3153 2232 3154
rect 1938 3114 2127 3144
rect 1953 3111 2127 3114
rect 1946 3108 2127 3111
rect 1755 3088 1768 3090
rect 1783 3088 1817 3090
rect 1755 3072 1829 3088
rect 1856 3084 1869 3098
rect 1884 3084 1900 3100
rect 1946 3095 1957 3108
rect 1739 3050 1740 3066
rect 1755 3050 1768 3072
rect 1783 3050 1813 3072
rect 1856 3068 1918 3084
rect 1946 3077 1957 3093
rect 1962 3088 1972 3108
rect 1982 3088 1996 3108
rect 1999 3095 2008 3108
rect 2024 3095 2033 3108
rect 1962 3077 1996 3088
rect 1999 3077 2008 3093
rect 2024 3077 2033 3093
rect 2040 3088 2050 3108
rect 2060 3088 2074 3108
rect 2075 3095 2086 3108
rect 2040 3077 2074 3088
rect 2075 3077 2086 3093
rect 2132 3084 2148 3100
rect 2155 3098 2185 3150
rect 2219 3146 2220 3153
rect 2204 3138 2220 3146
rect 2191 3106 2204 3125
rect 2219 3106 2249 3122
rect 2191 3090 2265 3106
rect 2191 3088 2204 3090
rect 2219 3088 2253 3090
rect 1856 3066 1869 3068
rect 1884 3066 1918 3068
rect 1856 3050 1918 3066
rect 1962 3061 1978 3064
rect 2040 3061 2070 3072
rect 2118 3068 2164 3084
rect 2191 3072 2265 3088
rect 2118 3066 2152 3068
rect 2117 3050 2164 3066
rect 2191 3050 2204 3072
rect 2219 3050 2249 3072
rect 2276 3050 2277 3066
rect 2292 3050 2305 3210
rect 2335 3106 2348 3210
rect 2393 3188 2394 3198
rect 2409 3188 2422 3198
rect 2393 3184 2422 3188
rect 2427 3184 2457 3210
rect 2475 3196 2491 3198
rect 2563 3196 2616 3210
rect 2564 3194 2628 3196
rect 2671 3194 2686 3210
rect 2735 3207 2765 3210
rect 2735 3204 2771 3207
rect 2701 3196 2717 3198
rect 2475 3184 2490 3188
rect 2393 3182 2490 3184
rect 2518 3182 2686 3194
rect 2702 3184 2717 3188
rect 2735 3185 2774 3204
rect 2793 3198 2800 3199
rect 2799 3191 2800 3198
rect 2783 3188 2784 3191
rect 2799 3188 2812 3191
rect 2735 3184 2765 3185
rect 2774 3184 2780 3185
rect 2783 3184 2812 3188
rect 2702 3183 2812 3184
rect 2702 3182 2818 3183
rect 2377 3174 2428 3182
rect 2377 3162 2402 3174
rect 2409 3162 2428 3174
rect 2459 3174 2509 3182
rect 2459 3166 2475 3174
rect 2482 3172 2509 3174
rect 2518 3172 2739 3182
rect 2482 3162 2739 3172
rect 2768 3174 2818 3182
rect 2768 3165 2784 3174
rect 2377 3154 2428 3162
rect 2475 3154 2739 3162
rect 2765 3162 2784 3165
rect 2791 3162 2818 3174
rect 2765 3154 2818 3162
rect 2393 3146 2394 3154
rect 2409 3146 2422 3154
rect 2393 3138 2409 3146
rect 2390 3131 2409 3134
rect 2390 3122 2412 3131
rect 2363 3112 2412 3122
rect 2363 3106 2393 3112
rect 2412 3107 2417 3112
rect 2335 3090 2409 3106
rect 2427 3098 2457 3154
rect 2492 3144 2700 3154
rect 2735 3150 2780 3154
rect 2783 3153 2784 3154
rect 2799 3153 2812 3154
rect 2518 3114 2707 3144
rect 2533 3111 2707 3114
rect 2526 3108 2707 3111
rect 2335 3088 2348 3090
rect 2363 3088 2397 3090
rect 2335 3072 2409 3088
rect 2436 3084 2449 3098
rect 2464 3084 2480 3100
rect 2526 3095 2537 3108
rect 2319 3050 2320 3066
rect 2335 3050 2348 3072
rect 2363 3050 2393 3072
rect 2436 3068 2498 3084
rect 2526 3077 2537 3093
rect 2542 3088 2552 3108
rect 2562 3088 2576 3108
rect 2579 3095 2588 3108
rect 2604 3095 2613 3108
rect 2542 3077 2576 3088
rect 2579 3077 2588 3093
rect 2604 3077 2613 3093
rect 2620 3088 2630 3108
rect 2640 3088 2654 3108
rect 2655 3095 2666 3108
rect 2620 3077 2654 3088
rect 2655 3077 2666 3093
rect 2712 3084 2728 3100
rect 2735 3098 2765 3150
rect 2799 3146 2800 3153
rect 2784 3138 2800 3146
rect 2771 3106 2784 3125
rect 2799 3106 2829 3122
rect 2771 3090 2845 3106
rect 2771 3088 2784 3090
rect 2799 3088 2833 3090
rect 2436 3066 2449 3068
rect 2464 3066 2498 3068
rect 2436 3050 2498 3066
rect 2542 3061 2558 3064
rect 2620 3061 2650 3072
rect 2698 3068 2744 3084
rect 2771 3072 2845 3088
rect 2698 3066 2732 3068
rect 2697 3050 2744 3066
rect 2771 3050 2784 3072
rect 2799 3050 2829 3072
rect 2856 3050 2857 3066
rect 2872 3050 2885 3210
rect 2915 3106 2928 3210
rect 2973 3188 2974 3198
rect 2989 3188 3002 3198
rect 2973 3184 3002 3188
rect 3007 3184 3037 3210
rect 3055 3196 3071 3198
rect 3143 3196 3196 3210
rect 3144 3194 3208 3196
rect 3251 3194 3266 3210
rect 3315 3207 3345 3210
rect 3315 3204 3351 3207
rect 3281 3196 3297 3198
rect 3055 3184 3070 3188
rect 2973 3182 3070 3184
rect 3098 3182 3266 3194
rect 3282 3184 3297 3188
rect 3315 3185 3354 3204
rect 3373 3198 3380 3199
rect 3379 3191 3380 3198
rect 3363 3188 3364 3191
rect 3379 3188 3392 3191
rect 3315 3184 3345 3185
rect 3354 3184 3360 3185
rect 3363 3184 3392 3188
rect 3282 3183 3392 3184
rect 3282 3182 3398 3183
rect 2957 3174 3008 3182
rect 2957 3162 2982 3174
rect 2989 3162 3008 3174
rect 3039 3174 3089 3182
rect 3039 3166 3055 3174
rect 3062 3172 3089 3174
rect 3098 3172 3319 3182
rect 3062 3162 3319 3172
rect 3348 3174 3398 3182
rect 3348 3165 3364 3174
rect 2957 3154 3008 3162
rect 3055 3154 3319 3162
rect 3345 3162 3364 3165
rect 3371 3162 3398 3174
rect 3345 3154 3398 3162
rect 2973 3146 2974 3154
rect 2989 3146 3002 3154
rect 2973 3138 2989 3146
rect 2970 3131 2989 3134
rect 2970 3122 2992 3131
rect 2943 3112 2992 3122
rect 2943 3106 2973 3112
rect 2992 3107 2997 3112
rect 2915 3090 2989 3106
rect 3007 3098 3037 3154
rect 3072 3144 3280 3154
rect 3315 3150 3360 3154
rect 3363 3153 3364 3154
rect 3379 3153 3392 3154
rect 3098 3114 3287 3144
rect 3113 3111 3287 3114
rect 3106 3108 3287 3111
rect 2915 3088 2928 3090
rect 2943 3088 2977 3090
rect 2915 3072 2989 3088
rect 3016 3084 3029 3098
rect 3044 3084 3060 3100
rect 3106 3095 3117 3108
rect 2899 3050 2900 3066
rect 2915 3050 2928 3072
rect 2943 3050 2973 3072
rect 3016 3068 3078 3084
rect 3106 3077 3117 3093
rect 3122 3088 3132 3108
rect 3142 3088 3156 3108
rect 3159 3095 3168 3108
rect 3184 3095 3193 3108
rect 3122 3077 3156 3088
rect 3159 3077 3168 3093
rect 3184 3077 3193 3093
rect 3200 3088 3210 3108
rect 3220 3088 3234 3108
rect 3235 3095 3246 3108
rect 3200 3077 3234 3088
rect 3235 3077 3246 3093
rect 3292 3084 3308 3100
rect 3315 3098 3345 3150
rect 3379 3146 3380 3153
rect 3364 3138 3380 3146
rect 3351 3106 3364 3125
rect 3379 3106 3409 3122
rect 3351 3090 3425 3106
rect 3351 3088 3364 3090
rect 3379 3088 3413 3090
rect 3016 3066 3029 3068
rect 3044 3066 3078 3068
rect 3016 3050 3078 3066
rect 3122 3061 3138 3064
rect 3200 3061 3230 3072
rect 3278 3068 3324 3084
rect 3351 3072 3425 3088
rect 3278 3066 3312 3068
rect 3277 3050 3324 3066
rect 3351 3050 3364 3072
rect 3379 3050 3409 3072
rect 3436 3050 3437 3066
rect 3452 3050 3465 3210
rect 3495 3106 3508 3210
rect 3553 3188 3554 3198
rect 3569 3188 3582 3198
rect 3553 3184 3582 3188
rect 3587 3184 3617 3210
rect 3635 3196 3651 3198
rect 3723 3196 3776 3210
rect 3724 3194 3788 3196
rect 3831 3194 3846 3210
rect 3895 3207 3925 3210
rect 3895 3204 3931 3207
rect 3861 3196 3877 3198
rect 3635 3184 3650 3188
rect 3553 3182 3650 3184
rect 3678 3182 3846 3194
rect 3862 3184 3877 3188
rect 3895 3185 3934 3204
rect 3953 3198 3960 3199
rect 3959 3191 3960 3198
rect 3943 3188 3944 3191
rect 3959 3188 3972 3191
rect 3895 3184 3925 3185
rect 3934 3184 3940 3185
rect 3943 3184 3972 3188
rect 3862 3183 3972 3184
rect 3862 3182 3978 3183
rect 3537 3174 3588 3182
rect 3537 3162 3562 3174
rect 3569 3162 3588 3174
rect 3619 3174 3669 3182
rect 3619 3166 3635 3174
rect 3642 3172 3669 3174
rect 3678 3172 3899 3182
rect 3642 3162 3899 3172
rect 3928 3174 3978 3182
rect 3928 3165 3944 3174
rect 3537 3154 3588 3162
rect 3635 3154 3899 3162
rect 3925 3162 3944 3165
rect 3951 3162 3978 3174
rect 3925 3154 3978 3162
rect 3553 3146 3554 3154
rect 3569 3146 3582 3154
rect 3553 3138 3569 3146
rect 3550 3131 3569 3134
rect 3550 3122 3572 3131
rect 3523 3112 3572 3122
rect 3523 3106 3553 3112
rect 3572 3107 3577 3112
rect 3495 3090 3569 3106
rect 3587 3098 3617 3154
rect 3652 3144 3860 3154
rect 3895 3150 3940 3154
rect 3943 3153 3944 3154
rect 3959 3153 3972 3154
rect 3678 3114 3867 3144
rect 3693 3111 3867 3114
rect 3686 3108 3867 3111
rect 3495 3088 3508 3090
rect 3523 3088 3557 3090
rect 3495 3072 3569 3088
rect 3596 3084 3609 3098
rect 3624 3084 3640 3100
rect 3686 3095 3697 3108
rect 3479 3050 3480 3066
rect 3495 3050 3508 3072
rect 3523 3050 3553 3072
rect 3596 3068 3658 3084
rect 3686 3077 3697 3093
rect 3702 3088 3712 3108
rect 3722 3088 3736 3108
rect 3739 3095 3748 3108
rect 3764 3095 3773 3108
rect 3702 3077 3736 3088
rect 3739 3077 3748 3093
rect 3764 3077 3773 3093
rect 3780 3088 3790 3108
rect 3800 3088 3814 3108
rect 3815 3095 3826 3108
rect 3780 3077 3814 3088
rect 3815 3077 3826 3093
rect 3872 3084 3888 3100
rect 3895 3098 3925 3150
rect 3959 3146 3960 3153
rect 3944 3138 3960 3146
rect 3931 3106 3944 3125
rect 3959 3106 3989 3122
rect 3931 3090 4005 3106
rect 3931 3088 3944 3090
rect 3959 3088 3993 3090
rect 3596 3066 3609 3068
rect 3624 3066 3658 3068
rect 3596 3050 3658 3066
rect 3702 3061 3718 3064
rect 3780 3061 3810 3072
rect 3858 3068 3904 3084
rect 3931 3072 4005 3088
rect 3858 3066 3892 3068
rect 3857 3050 3904 3066
rect 3931 3050 3944 3072
rect 3959 3050 3989 3072
rect 4016 3050 4017 3066
rect 4032 3050 4045 3210
rect 4075 3106 4088 3210
rect 4133 3188 4134 3198
rect 4149 3188 4162 3198
rect 4133 3184 4162 3188
rect 4167 3184 4197 3210
rect 4215 3196 4231 3198
rect 4303 3196 4356 3210
rect 4304 3194 4368 3196
rect 4411 3194 4426 3210
rect 4475 3207 4505 3210
rect 4475 3204 4511 3207
rect 4441 3196 4457 3198
rect 4215 3184 4230 3188
rect 4133 3182 4230 3184
rect 4258 3182 4426 3194
rect 4442 3184 4457 3188
rect 4475 3185 4514 3204
rect 4533 3198 4540 3199
rect 4539 3191 4540 3198
rect 4523 3188 4524 3191
rect 4539 3188 4552 3191
rect 4475 3184 4505 3185
rect 4514 3184 4520 3185
rect 4523 3184 4552 3188
rect 4442 3183 4552 3184
rect 4442 3182 4558 3183
rect 4117 3174 4168 3182
rect 4117 3162 4142 3174
rect 4149 3162 4168 3174
rect 4199 3174 4249 3182
rect 4199 3166 4215 3174
rect 4222 3172 4249 3174
rect 4258 3172 4479 3182
rect 4222 3162 4479 3172
rect 4508 3174 4558 3182
rect 4508 3165 4524 3174
rect 4117 3154 4168 3162
rect 4215 3154 4479 3162
rect 4505 3162 4524 3165
rect 4531 3162 4558 3174
rect 4505 3154 4558 3162
rect 4133 3146 4134 3154
rect 4149 3146 4162 3154
rect 4133 3138 4149 3146
rect 4130 3131 4149 3134
rect 4130 3122 4152 3131
rect 4103 3112 4152 3122
rect 4103 3106 4133 3112
rect 4152 3107 4157 3112
rect 4075 3090 4149 3106
rect 4167 3098 4197 3154
rect 4232 3144 4440 3154
rect 4475 3150 4520 3154
rect 4523 3153 4524 3154
rect 4539 3153 4552 3154
rect 4258 3114 4447 3144
rect 4273 3111 4447 3114
rect 4266 3108 4447 3111
rect 4075 3088 4088 3090
rect 4103 3088 4137 3090
rect 4075 3072 4149 3088
rect 4176 3084 4189 3098
rect 4204 3084 4220 3100
rect 4266 3095 4277 3108
rect 4059 3050 4060 3066
rect 4075 3050 4088 3072
rect 4103 3050 4133 3072
rect 4176 3068 4238 3084
rect 4266 3077 4277 3093
rect 4282 3088 4292 3108
rect 4302 3088 4316 3108
rect 4319 3095 4328 3108
rect 4344 3095 4353 3108
rect 4282 3077 4316 3088
rect 4319 3077 4328 3093
rect 4344 3077 4353 3093
rect 4360 3088 4370 3108
rect 4380 3088 4394 3108
rect 4395 3095 4406 3108
rect 4360 3077 4394 3088
rect 4395 3077 4406 3093
rect 4452 3084 4468 3100
rect 4475 3098 4505 3150
rect 4539 3146 4540 3153
rect 4524 3138 4540 3146
rect 4511 3106 4524 3125
rect 4539 3106 4569 3122
rect 4511 3090 4585 3106
rect 4511 3088 4524 3090
rect 4539 3088 4573 3090
rect 4176 3066 4189 3068
rect 4204 3066 4238 3068
rect 4176 3050 4238 3066
rect 4282 3061 4298 3064
rect 4360 3061 4390 3072
rect 4438 3068 4484 3084
rect 4511 3072 4585 3088
rect 4438 3066 4472 3068
rect 4437 3050 4484 3066
rect 4511 3050 4524 3072
rect 4539 3050 4569 3072
rect 4596 3050 4597 3066
rect 4612 3050 4625 3210
rect -7 3042 34 3050
rect -7 3016 8 3042
rect 15 3016 34 3042
rect 98 3038 160 3050
rect 172 3038 247 3050
rect 305 3038 380 3050
rect 392 3038 423 3050
rect 429 3038 464 3050
rect 98 3036 260 3038
rect -7 3008 34 3016
rect 116 3012 129 3036
rect 144 3034 159 3036
rect -1 2998 0 3008
rect 15 2998 28 3008
rect 43 2998 73 3012
rect 116 2998 159 3012
rect 183 3009 190 3016
rect 193 3012 260 3036
rect 292 3036 464 3038
rect 262 3014 290 3018
rect 292 3014 372 3036
rect 393 3034 408 3036
rect 262 3012 372 3014
rect 193 3008 372 3012
rect 166 2998 196 3008
rect 198 2998 351 3008
rect 359 2998 389 3008
rect 393 2998 423 3012
rect 451 2998 464 3036
rect 536 3042 571 3050
rect 536 3016 537 3042
rect 544 3016 571 3042
rect 479 2998 509 3012
rect 536 3008 571 3016
rect 573 3042 614 3050
rect 573 3016 588 3042
rect 595 3016 614 3042
rect 678 3038 740 3050
rect 752 3038 827 3050
rect 885 3038 960 3050
rect 972 3038 1003 3050
rect 1009 3038 1044 3050
rect 678 3036 840 3038
rect 573 3008 614 3016
rect 696 3012 709 3036
rect 724 3034 739 3036
rect 536 2998 537 3008
rect 552 2998 565 3008
rect 579 2998 580 3008
rect 595 2998 608 3008
rect 623 2998 653 3012
rect 696 2998 739 3012
rect 763 3009 770 3016
rect 773 3012 840 3036
rect 872 3036 1044 3038
rect 842 3014 870 3018
rect 872 3014 952 3036
rect 973 3034 988 3036
rect 842 3012 952 3014
rect 773 3008 952 3012
rect 746 2998 776 3008
rect 778 2998 931 3008
rect 939 2998 969 3008
rect 973 2998 1003 3012
rect 1031 2998 1044 3036
rect 1116 3042 1151 3050
rect 1116 3016 1117 3042
rect 1124 3016 1151 3042
rect 1059 2998 1089 3012
rect 1116 3008 1151 3016
rect 1153 3042 1194 3050
rect 1153 3016 1168 3042
rect 1175 3016 1194 3042
rect 1258 3038 1320 3050
rect 1332 3038 1407 3050
rect 1465 3038 1540 3050
rect 1552 3038 1583 3050
rect 1589 3038 1624 3050
rect 1258 3036 1420 3038
rect 1153 3008 1194 3016
rect 1276 3012 1289 3036
rect 1304 3034 1319 3036
rect 1116 2998 1117 3008
rect 1132 2998 1145 3008
rect 1159 2998 1160 3008
rect 1175 2998 1188 3008
rect 1203 2998 1233 3012
rect 1276 2998 1319 3012
rect 1343 3009 1350 3016
rect 1353 3012 1420 3036
rect 1452 3036 1624 3038
rect 1422 3014 1450 3018
rect 1452 3014 1532 3036
rect 1553 3034 1568 3036
rect 1422 3012 1532 3014
rect 1353 3008 1532 3012
rect 1326 2998 1356 3008
rect 1358 2998 1511 3008
rect 1519 2998 1549 3008
rect 1553 2998 1583 3012
rect 1611 2998 1624 3036
rect 1696 3042 1731 3050
rect 1696 3016 1697 3042
rect 1704 3016 1731 3042
rect 1639 2998 1669 3012
rect 1696 3008 1731 3016
rect 1733 3042 1774 3050
rect 1733 3016 1748 3042
rect 1755 3016 1774 3042
rect 1838 3038 1900 3050
rect 1912 3038 1987 3050
rect 2045 3038 2120 3050
rect 2132 3038 2163 3050
rect 2169 3038 2204 3050
rect 1838 3036 2000 3038
rect 1733 3008 1774 3016
rect 1856 3012 1869 3036
rect 1884 3034 1899 3036
rect 1696 2998 1697 3008
rect 1712 2998 1725 3008
rect 1739 2998 1740 3008
rect 1755 2998 1768 3008
rect 1783 2998 1813 3012
rect 1856 2998 1899 3012
rect 1923 3009 1930 3016
rect 1933 3012 2000 3036
rect 2032 3036 2204 3038
rect 2002 3014 2030 3018
rect 2032 3014 2112 3036
rect 2133 3034 2148 3036
rect 2002 3012 2112 3014
rect 1933 3008 2112 3012
rect 1906 2998 1936 3008
rect 1938 2998 2091 3008
rect 2099 2998 2129 3008
rect 2133 2998 2163 3012
rect 2191 2998 2204 3036
rect 2276 3042 2311 3050
rect 2276 3016 2277 3042
rect 2284 3016 2311 3042
rect 2219 2998 2249 3012
rect 2276 3008 2311 3016
rect 2313 3042 2354 3050
rect 2313 3016 2328 3042
rect 2335 3016 2354 3042
rect 2418 3038 2480 3050
rect 2492 3038 2567 3050
rect 2625 3038 2700 3050
rect 2712 3038 2743 3050
rect 2749 3038 2784 3050
rect 2418 3036 2580 3038
rect 2313 3008 2354 3016
rect 2436 3012 2449 3036
rect 2464 3034 2479 3036
rect 2276 2998 2277 3008
rect 2292 2998 2305 3008
rect 2319 2998 2320 3008
rect 2335 2998 2348 3008
rect 2363 2998 2393 3012
rect 2436 2998 2479 3012
rect 2503 3009 2510 3016
rect 2513 3012 2580 3036
rect 2612 3036 2784 3038
rect 2582 3014 2610 3018
rect 2612 3014 2692 3036
rect 2713 3034 2728 3036
rect 2582 3012 2692 3014
rect 2513 3008 2692 3012
rect 2486 2998 2516 3008
rect 2518 2998 2671 3008
rect 2679 2998 2709 3008
rect 2713 2998 2743 3012
rect 2771 2998 2784 3036
rect 2856 3042 2891 3050
rect 2856 3016 2857 3042
rect 2864 3016 2891 3042
rect 2799 2998 2829 3012
rect 2856 3008 2891 3016
rect 2893 3042 2934 3050
rect 2893 3016 2908 3042
rect 2915 3016 2934 3042
rect 2998 3038 3060 3050
rect 3072 3038 3147 3050
rect 3205 3038 3280 3050
rect 3292 3038 3323 3050
rect 3329 3038 3364 3050
rect 2998 3036 3160 3038
rect 2893 3008 2934 3016
rect 3016 3012 3029 3036
rect 3044 3034 3059 3036
rect 2856 2998 2857 3008
rect 2872 2998 2885 3008
rect 2899 2998 2900 3008
rect 2915 2998 2928 3008
rect 2943 2998 2973 3012
rect 3016 2998 3059 3012
rect 3083 3009 3090 3016
rect 3093 3012 3160 3036
rect 3192 3036 3364 3038
rect 3162 3014 3190 3018
rect 3192 3014 3272 3036
rect 3293 3034 3308 3036
rect 3162 3012 3272 3014
rect 3093 3008 3272 3012
rect 3066 2998 3096 3008
rect 3098 2998 3251 3008
rect 3259 2998 3289 3008
rect 3293 2998 3323 3012
rect 3351 2998 3364 3036
rect 3436 3042 3471 3050
rect 3436 3016 3437 3042
rect 3444 3016 3471 3042
rect 3379 2998 3409 3012
rect 3436 3008 3471 3016
rect 3473 3042 3514 3050
rect 3473 3016 3488 3042
rect 3495 3016 3514 3042
rect 3578 3038 3640 3050
rect 3652 3038 3727 3050
rect 3785 3038 3860 3050
rect 3872 3038 3903 3050
rect 3909 3038 3944 3050
rect 3578 3036 3740 3038
rect 3473 3008 3514 3016
rect 3596 3012 3609 3036
rect 3624 3034 3639 3036
rect 3436 2998 3437 3008
rect 3452 2998 3465 3008
rect 3479 2998 3480 3008
rect 3495 2998 3508 3008
rect 3523 2998 3553 3012
rect 3596 2998 3639 3012
rect 3663 3009 3670 3016
rect 3673 3012 3740 3036
rect 3772 3036 3944 3038
rect 3742 3014 3770 3018
rect 3772 3014 3852 3036
rect 3873 3034 3888 3036
rect 3742 3012 3852 3014
rect 3673 3008 3852 3012
rect 3646 2998 3676 3008
rect 3678 2998 3831 3008
rect 3839 2998 3869 3008
rect 3873 2998 3903 3012
rect 3931 2998 3944 3036
rect 4016 3042 4051 3050
rect 4016 3016 4017 3042
rect 4024 3016 4051 3042
rect 3959 2998 3989 3012
rect 4016 3008 4051 3016
rect 4053 3042 4094 3050
rect 4053 3016 4068 3042
rect 4075 3016 4094 3042
rect 4158 3038 4220 3050
rect 4232 3038 4307 3050
rect 4365 3038 4440 3050
rect 4452 3038 4483 3050
rect 4489 3038 4524 3050
rect 4158 3036 4320 3038
rect 4053 3008 4094 3016
rect 4176 3012 4189 3036
rect 4204 3034 4219 3036
rect 4016 2998 4017 3008
rect 4032 2998 4045 3008
rect 4059 2998 4060 3008
rect 4075 2998 4088 3008
rect 4103 2998 4133 3012
rect 4176 2998 4219 3012
rect 4243 3009 4250 3016
rect 4253 3012 4320 3036
rect 4352 3036 4524 3038
rect 4322 3014 4350 3018
rect 4352 3014 4432 3036
rect 4453 3034 4468 3036
rect 4322 3012 4432 3014
rect 4253 3008 4432 3012
rect 4226 2998 4256 3008
rect 4258 2998 4411 3008
rect 4419 2998 4449 3008
rect 4453 2998 4483 3012
rect 4511 2998 4524 3036
rect 4596 3042 4631 3050
rect 4596 3016 4597 3042
rect 4604 3016 4631 3042
rect 4539 2998 4569 3012
rect 4596 3008 4631 3016
rect 4596 2998 4597 3008
rect 4612 2998 4625 3008
rect -1 2992 4625 2998
rect 0 2984 4625 2992
rect 15 2954 28 2984
rect 43 2966 73 2984
rect 116 2970 130 2984
rect 166 2970 386 2984
rect 117 2968 130 2970
rect 83 2956 98 2968
rect 80 2954 102 2956
rect 107 2954 137 2968
rect 198 2966 351 2970
rect 180 2954 372 2966
rect 415 2954 445 2968
rect 451 2954 464 2984
rect 479 2966 509 2984
rect 552 2954 565 2984
rect 595 2954 608 2984
rect 623 2966 653 2984
rect 696 2970 710 2984
rect 746 2970 966 2984
rect 697 2968 710 2970
rect 663 2956 678 2968
rect 660 2954 682 2956
rect 687 2954 717 2968
rect 778 2966 931 2970
rect 760 2954 952 2966
rect 995 2954 1025 2968
rect 1031 2954 1044 2984
rect 1059 2966 1089 2984
rect 1132 2954 1145 2984
rect 1175 2954 1188 2984
rect 1203 2966 1233 2984
rect 1276 2970 1290 2984
rect 1326 2970 1546 2984
rect 1277 2968 1290 2970
rect 1243 2956 1258 2968
rect 1240 2954 1262 2956
rect 1267 2954 1297 2968
rect 1358 2966 1511 2970
rect 1340 2954 1532 2966
rect 1575 2954 1605 2968
rect 1611 2954 1624 2984
rect 1639 2966 1669 2984
rect 1712 2954 1725 2984
rect 1755 2954 1768 2984
rect 1783 2966 1813 2984
rect 1856 2970 1870 2984
rect 1906 2970 2126 2984
rect 1857 2968 1870 2970
rect 1823 2956 1838 2968
rect 1820 2954 1842 2956
rect 1847 2954 1877 2968
rect 1938 2966 2091 2970
rect 1920 2954 2112 2966
rect 2155 2954 2185 2968
rect 2191 2954 2204 2984
rect 2219 2966 2249 2984
rect 2292 2954 2305 2984
rect 2335 2954 2348 2984
rect 2363 2966 2393 2984
rect 2436 2970 2450 2984
rect 2486 2970 2706 2984
rect 2437 2968 2450 2970
rect 2403 2956 2418 2968
rect 2400 2954 2422 2956
rect 2427 2954 2457 2968
rect 2518 2966 2671 2970
rect 2500 2954 2692 2966
rect 2735 2954 2765 2968
rect 2771 2954 2784 2984
rect 2799 2966 2829 2984
rect 2872 2954 2885 2984
rect 2915 2954 2928 2984
rect 2943 2966 2973 2984
rect 3016 2970 3030 2984
rect 3066 2970 3286 2984
rect 3017 2968 3030 2970
rect 2983 2956 2998 2968
rect 2980 2954 3002 2956
rect 3007 2954 3037 2968
rect 3098 2966 3251 2970
rect 3080 2954 3272 2966
rect 3315 2954 3345 2968
rect 3351 2954 3364 2984
rect 3379 2966 3409 2984
rect 3452 2954 3465 2984
rect 3495 2954 3508 2984
rect 3523 2966 3553 2984
rect 3596 2970 3610 2984
rect 3646 2970 3866 2984
rect 3597 2968 3610 2970
rect 3563 2956 3578 2968
rect 3560 2954 3582 2956
rect 3587 2954 3617 2968
rect 3678 2966 3831 2970
rect 3660 2954 3852 2966
rect 3895 2954 3925 2968
rect 3931 2954 3944 2984
rect 3959 2966 3989 2984
rect 4032 2954 4045 2984
rect 4075 2954 4088 2984
rect 4103 2966 4133 2984
rect 4176 2970 4190 2984
rect 4226 2970 4446 2984
rect 4177 2968 4190 2970
rect 4143 2956 4158 2968
rect 4140 2954 4162 2956
rect 4167 2954 4197 2968
rect 4258 2966 4411 2970
rect 4240 2954 4432 2966
rect 4475 2954 4505 2968
rect 4511 2954 4524 2984
rect 4539 2966 4569 2984
rect 4612 2954 4625 2984
rect 0 2940 4625 2954
rect 15 2836 28 2940
rect 73 2918 74 2928
rect 89 2918 102 2928
rect 73 2914 102 2918
rect 107 2914 137 2940
rect 155 2926 171 2928
rect 243 2926 296 2940
rect 244 2924 308 2926
rect 351 2924 366 2940
rect 415 2937 445 2940
rect 415 2934 451 2937
rect 381 2926 397 2928
rect 155 2914 170 2918
rect 73 2912 170 2914
rect 198 2912 366 2924
rect 382 2914 397 2918
rect 415 2915 454 2934
rect 473 2928 480 2929
rect 479 2921 480 2928
rect 463 2918 464 2921
rect 479 2918 492 2921
rect 415 2914 445 2915
rect 454 2914 460 2915
rect 463 2914 492 2918
rect 382 2913 492 2914
rect 382 2912 498 2913
rect 57 2904 108 2912
rect 57 2892 82 2904
rect 89 2892 108 2904
rect 139 2904 189 2912
rect 139 2896 155 2904
rect 162 2902 189 2904
rect 198 2902 419 2912
rect 162 2892 419 2902
rect 448 2904 498 2912
rect 448 2895 464 2904
rect 57 2884 108 2892
rect 155 2884 419 2892
rect 445 2892 464 2895
rect 471 2892 498 2904
rect 445 2884 498 2892
rect 73 2876 74 2884
rect 89 2876 102 2884
rect 73 2868 89 2876
rect 70 2861 89 2864
rect 70 2852 92 2861
rect 43 2842 92 2852
rect 43 2836 73 2842
rect 92 2837 97 2842
rect 15 2820 89 2836
rect 107 2828 137 2884
rect 172 2874 380 2884
rect 415 2880 460 2884
rect 463 2883 464 2884
rect 479 2883 492 2884
rect 198 2844 387 2874
rect 213 2841 387 2844
rect 206 2838 387 2841
rect 15 2818 28 2820
rect 43 2818 77 2820
rect 15 2802 89 2818
rect 116 2814 129 2828
rect 144 2814 160 2830
rect 206 2825 217 2838
rect -1 2780 0 2796
rect 15 2780 28 2802
rect 43 2780 73 2802
rect 116 2798 178 2814
rect 206 2807 217 2823
rect 222 2818 232 2838
rect 242 2818 256 2838
rect 259 2825 268 2838
rect 284 2825 293 2838
rect 222 2807 256 2818
rect 259 2807 268 2823
rect 284 2807 293 2823
rect 300 2818 310 2838
rect 320 2818 334 2838
rect 335 2825 346 2838
rect 300 2807 334 2818
rect 335 2807 346 2823
rect 392 2814 408 2830
rect 415 2828 445 2880
rect 479 2876 480 2883
rect 464 2868 480 2876
rect 451 2836 464 2855
rect 479 2836 509 2852
rect 451 2820 525 2836
rect 451 2818 464 2820
rect 479 2818 513 2820
rect 116 2796 129 2798
rect 144 2796 178 2798
rect 116 2780 178 2796
rect 222 2791 238 2794
rect 300 2791 330 2802
rect 378 2798 424 2814
rect 451 2802 525 2818
rect 378 2796 412 2798
rect 377 2780 424 2796
rect 451 2780 464 2802
rect 479 2780 509 2802
rect 536 2780 537 2796
rect 552 2780 565 2940
rect 595 2836 608 2940
rect 653 2918 654 2928
rect 669 2918 682 2928
rect 653 2914 682 2918
rect 687 2914 717 2940
rect 735 2926 751 2928
rect 823 2926 876 2940
rect 824 2924 888 2926
rect 931 2924 946 2940
rect 995 2937 1025 2940
rect 995 2934 1031 2937
rect 961 2926 977 2928
rect 735 2914 750 2918
rect 653 2912 750 2914
rect 778 2912 946 2924
rect 962 2914 977 2918
rect 995 2915 1034 2934
rect 1053 2928 1060 2929
rect 1059 2921 1060 2928
rect 1043 2918 1044 2921
rect 1059 2918 1072 2921
rect 995 2914 1025 2915
rect 1034 2914 1040 2915
rect 1043 2914 1072 2918
rect 962 2913 1072 2914
rect 962 2912 1078 2913
rect 637 2904 688 2912
rect 637 2892 662 2904
rect 669 2892 688 2904
rect 719 2904 769 2912
rect 719 2896 735 2904
rect 742 2902 769 2904
rect 778 2902 999 2912
rect 742 2892 999 2902
rect 1028 2904 1078 2912
rect 1028 2895 1044 2904
rect 637 2884 688 2892
rect 735 2884 999 2892
rect 1025 2892 1044 2895
rect 1051 2892 1078 2904
rect 1025 2884 1078 2892
rect 653 2876 654 2884
rect 669 2876 682 2884
rect 653 2868 669 2876
rect 650 2861 669 2864
rect 650 2852 672 2861
rect 623 2842 672 2852
rect 623 2836 653 2842
rect 672 2837 677 2842
rect 595 2820 669 2836
rect 687 2828 717 2884
rect 752 2874 960 2884
rect 995 2880 1040 2884
rect 1043 2883 1044 2884
rect 1059 2883 1072 2884
rect 778 2844 967 2874
rect 793 2841 967 2844
rect 786 2838 967 2841
rect 595 2818 608 2820
rect 623 2818 657 2820
rect 595 2802 669 2818
rect 696 2814 709 2828
rect 724 2814 740 2830
rect 786 2825 797 2838
rect 579 2780 580 2796
rect 595 2780 608 2802
rect 623 2780 653 2802
rect 696 2798 758 2814
rect 786 2807 797 2823
rect 802 2818 812 2838
rect 822 2818 836 2838
rect 839 2825 848 2838
rect 864 2825 873 2838
rect 802 2807 836 2818
rect 839 2807 848 2823
rect 864 2807 873 2823
rect 880 2818 890 2838
rect 900 2818 914 2838
rect 915 2825 926 2838
rect 880 2807 914 2818
rect 915 2807 926 2823
rect 972 2814 988 2830
rect 995 2828 1025 2880
rect 1059 2876 1060 2883
rect 1044 2868 1060 2876
rect 1031 2836 1044 2855
rect 1059 2836 1089 2852
rect 1031 2820 1105 2836
rect 1031 2818 1044 2820
rect 1059 2818 1093 2820
rect 696 2796 709 2798
rect 724 2796 758 2798
rect 696 2780 758 2796
rect 802 2791 818 2794
rect 880 2791 910 2802
rect 958 2798 1004 2814
rect 1031 2802 1105 2818
rect 958 2796 992 2798
rect 957 2780 1004 2796
rect 1031 2780 1044 2802
rect 1059 2780 1089 2802
rect 1116 2780 1117 2796
rect 1132 2780 1145 2940
rect 1175 2836 1188 2940
rect 1233 2918 1234 2928
rect 1249 2918 1262 2928
rect 1233 2914 1262 2918
rect 1267 2914 1297 2940
rect 1315 2926 1331 2928
rect 1403 2926 1456 2940
rect 1404 2924 1468 2926
rect 1511 2924 1526 2940
rect 1575 2937 1605 2940
rect 1575 2934 1611 2937
rect 1541 2926 1557 2928
rect 1315 2914 1330 2918
rect 1233 2912 1330 2914
rect 1358 2912 1526 2924
rect 1542 2914 1557 2918
rect 1575 2915 1614 2934
rect 1633 2928 1640 2929
rect 1639 2921 1640 2928
rect 1623 2918 1624 2921
rect 1639 2918 1652 2921
rect 1575 2914 1605 2915
rect 1614 2914 1620 2915
rect 1623 2914 1652 2918
rect 1542 2913 1652 2914
rect 1542 2912 1658 2913
rect 1217 2904 1268 2912
rect 1217 2892 1242 2904
rect 1249 2892 1268 2904
rect 1299 2904 1349 2912
rect 1299 2896 1315 2904
rect 1322 2902 1349 2904
rect 1358 2902 1579 2912
rect 1322 2892 1579 2902
rect 1608 2904 1658 2912
rect 1608 2895 1624 2904
rect 1217 2884 1268 2892
rect 1315 2884 1579 2892
rect 1605 2892 1624 2895
rect 1631 2892 1658 2904
rect 1605 2884 1658 2892
rect 1233 2876 1234 2884
rect 1249 2876 1262 2884
rect 1233 2868 1249 2876
rect 1230 2861 1249 2864
rect 1230 2852 1252 2861
rect 1203 2842 1252 2852
rect 1203 2836 1233 2842
rect 1252 2837 1257 2842
rect 1175 2820 1249 2836
rect 1267 2828 1297 2884
rect 1332 2874 1540 2884
rect 1575 2880 1620 2884
rect 1623 2883 1624 2884
rect 1639 2883 1652 2884
rect 1358 2844 1547 2874
rect 1373 2841 1547 2844
rect 1366 2838 1547 2841
rect 1175 2818 1188 2820
rect 1203 2818 1237 2820
rect 1175 2802 1249 2818
rect 1276 2814 1289 2828
rect 1304 2814 1320 2830
rect 1366 2825 1377 2838
rect 1159 2780 1160 2796
rect 1175 2780 1188 2802
rect 1203 2780 1233 2802
rect 1276 2798 1338 2814
rect 1366 2807 1377 2823
rect 1382 2818 1392 2838
rect 1402 2818 1416 2838
rect 1419 2825 1428 2838
rect 1444 2825 1453 2838
rect 1382 2807 1416 2818
rect 1419 2807 1428 2823
rect 1444 2807 1453 2823
rect 1460 2818 1470 2838
rect 1480 2818 1494 2838
rect 1495 2825 1506 2838
rect 1460 2807 1494 2818
rect 1495 2807 1506 2823
rect 1552 2814 1568 2830
rect 1575 2828 1605 2880
rect 1639 2876 1640 2883
rect 1624 2868 1640 2876
rect 1611 2836 1624 2855
rect 1639 2836 1669 2852
rect 1611 2820 1685 2836
rect 1611 2818 1624 2820
rect 1639 2818 1673 2820
rect 1276 2796 1289 2798
rect 1304 2796 1338 2798
rect 1276 2780 1338 2796
rect 1382 2791 1398 2794
rect 1460 2791 1490 2802
rect 1538 2798 1584 2814
rect 1611 2802 1685 2818
rect 1538 2796 1572 2798
rect 1537 2780 1584 2796
rect 1611 2780 1624 2802
rect 1639 2780 1669 2802
rect 1696 2780 1697 2796
rect 1712 2780 1725 2940
rect 1755 2836 1768 2940
rect 1813 2918 1814 2928
rect 1829 2918 1842 2928
rect 1813 2914 1842 2918
rect 1847 2914 1877 2940
rect 1895 2926 1911 2928
rect 1983 2926 2036 2940
rect 1984 2924 2048 2926
rect 2091 2924 2106 2940
rect 2155 2937 2185 2940
rect 2155 2934 2191 2937
rect 2121 2926 2137 2928
rect 1895 2914 1910 2918
rect 1813 2912 1910 2914
rect 1938 2912 2106 2924
rect 2122 2914 2137 2918
rect 2155 2915 2194 2934
rect 2213 2928 2220 2929
rect 2219 2921 2220 2928
rect 2203 2918 2204 2921
rect 2219 2918 2232 2921
rect 2155 2914 2185 2915
rect 2194 2914 2200 2915
rect 2203 2914 2232 2918
rect 2122 2913 2232 2914
rect 2122 2912 2238 2913
rect 1797 2904 1848 2912
rect 1797 2892 1822 2904
rect 1829 2892 1848 2904
rect 1879 2904 1929 2912
rect 1879 2896 1895 2904
rect 1902 2902 1929 2904
rect 1938 2902 2159 2912
rect 1902 2892 2159 2902
rect 2188 2904 2238 2912
rect 2188 2895 2204 2904
rect 1797 2884 1848 2892
rect 1895 2884 2159 2892
rect 2185 2892 2204 2895
rect 2211 2892 2238 2904
rect 2185 2884 2238 2892
rect 1813 2876 1814 2884
rect 1829 2876 1842 2884
rect 1813 2868 1829 2876
rect 1810 2861 1829 2864
rect 1810 2852 1832 2861
rect 1783 2842 1832 2852
rect 1783 2836 1813 2842
rect 1832 2837 1837 2842
rect 1755 2820 1829 2836
rect 1847 2828 1877 2884
rect 1912 2874 2120 2884
rect 2155 2880 2200 2884
rect 2203 2883 2204 2884
rect 2219 2883 2232 2884
rect 1938 2844 2127 2874
rect 1953 2841 2127 2844
rect 1946 2838 2127 2841
rect 1755 2818 1768 2820
rect 1783 2818 1817 2820
rect 1755 2802 1829 2818
rect 1856 2814 1869 2828
rect 1884 2814 1900 2830
rect 1946 2825 1957 2838
rect 1739 2780 1740 2796
rect 1755 2780 1768 2802
rect 1783 2780 1813 2802
rect 1856 2798 1918 2814
rect 1946 2807 1957 2823
rect 1962 2818 1972 2838
rect 1982 2818 1996 2838
rect 1999 2825 2008 2838
rect 2024 2825 2033 2838
rect 1962 2807 1996 2818
rect 1999 2807 2008 2823
rect 2024 2807 2033 2823
rect 2040 2818 2050 2838
rect 2060 2818 2074 2838
rect 2075 2825 2086 2838
rect 2040 2807 2074 2818
rect 2075 2807 2086 2823
rect 2132 2814 2148 2830
rect 2155 2828 2185 2880
rect 2219 2876 2220 2883
rect 2204 2868 2220 2876
rect 2191 2836 2204 2855
rect 2219 2836 2249 2852
rect 2191 2820 2265 2836
rect 2191 2818 2204 2820
rect 2219 2818 2253 2820
rect 1856 2796 1869 2798
rect 1884 2796 1918 2798
rect 1856 2780 1918 2796
rect 1962 2791 1978 2794
rect 2040 2791 2070 2802
rect 2118 2798 2164 2814
rect 2191 2802 2265 2818
rect 2118 2796 2152 2798
rect 2117 2780 2164 2796
rect 2191 2780 2204 2802
rect 2219 2780 2249 2802
rect 2276 2780 2277 2796
rect 2292 2780 2305 2940
rect 2335 2836 2348 2940
rect 2393 2918 2394 2928
rect 2409 2918 2422 2928
rect 2393 2914 2422 2918
rect 2427 2914 2457 2940
rect 2475 2926 2491 2928
rect 2563 2926 2616 2940
rect 2564 2924 2628 2926
rect 2671 2924 2686 2940
rect 2735 2937 2765 2940
rect 2735 2934 2771 2937
rect 2701 2926 2717 2928
rect 2475 2914 2490 2918
rect 2393 2912 2490 2914
rect 2518 2912 2686 2924
rect 2702 2914 2717 2918
rect 2735 2915 2774 2934
rect 2793 2928 2800 2929
rect 2799 2921 2800 2928
rect 2783 2918 2784 2921
rect 2799 2918 2812 2921
rect 2735 2914 2765 2915
rect 2774 2914 2780 2915
rect 2783 2914 2812 2918
rect 2702 2913 2812 2914
rect 2702 2912 2818 2913
rect 2377 2904 2428 2912
rect 2377 2892 2402 2904
rect 2409 2892 2428 2904
rect 2459 2904 2509 2912
rect 2459 2896 2475 2904
rect 2482 2902 2509 2904
rect 2518 2902 2739 2912
rect 2482 2892 2739 2902
rect 2768 2904 2818 2912
rect 2768 2895 2784 2904
rect 2377 2884 2428 2892
rect 2475 2884 2739 2892
rect 2765 2892 2784 2895
rect 2791 2892 2818 2904
rect 2765 2884 2818 2892
rect 2393 2876 2394 2884
rect 2409 2876 2422 2884
rect 2393 2868 2409 2876
rect 2390 2861 2409 2864
rect 2390 2852 2412 2861
rect 2363 2842 2412 2852
rect 2363 2836 2393 2842
rect 2412 2837 2417 2842
rect 2335 2820 2409 2836
rect 2427 2828 2457 2884
rect 2492 2874 2700 2884
rect 2735 2880 2780 2884
rect 2783 2883 2784 2884
rect 2799 2883 2812 2884
rect 2518 2844 2707 2874
rect 2533 2841 2707 2844
rect 2526 2838 2707 2841
rect 2335 2818 2348 2820
rect 2363 2818 2397 2820
rect 2335 2802 2409 2818
rect 2436 2814 2449 2828
rect 2464 2814 2480 2830
rect 2526 2825 2537 2838
rect 2319 2780 2320 2796
rect 2335 2780 2348 2802
rect 2363 2780 2393 2802
rect 2436 2798 2498 2814
rect 2526 2807 2537 2823
rect 2542 2818 2552 2838
rect 2562 2818 2576 2838
rect 2579 2825 2588 2838
rect 2604 2825 2613 2838
rect 2542 2807 2576 2818
rect 2579 2807 2588 2823
rect 2604 2807 2613 2823
rect 2620 2818 2630 2838
rect 2640 2818 2654 2838
rect 2655 2825 2666 2838
rect 2620 2807 2654 2818
rect 2655 2807 2666 2823
rect 2712 2814 2728 2830
rect 2735 2828 2765 2880
rect 2799 2876 2800 2883
rect 2784 2868 2800 2876
rect 2771 2836 2784 2855
rect 2799 2836 2829 2852
rect 2771 2820 2845 2836
rect 2771 2818 2784 2820
rect 2799 2818 2833 2820
rect 2436 2796 2449 2798
rect 2464 2796 2498 2798
rect 2436 2780 2498 2796
rect 2542 2791 2558 2794
rect 2620 2791 2650 2802
rect 2698 2798 2744 2814
rect 2771 2802 2845 2818
rect 2698 2796 2732 2798
rect 2697 2780 2744 2796
rect 2771 2780 2784 2802
rect 2799 2780 2829 2802
rect 2856 2780 2857 2796
rect 2872 2780 2885 2940
rect 2915 2836 2928 2940
rect 2973 2918 2974 2928
rect 2989 2918 3002 2928
rect 2973 2914 3002 2918
rect 3007 2914 3037 2940
rect 3055 2926 3071 2928
rect 3143 2926 3196 2940
rect 3144 2924 3208 2926
rect 3251 2924 3266 2940
rect 3315 2937 3345 2940
rect 3315 2934 3351 2937
rect 3281 2926 3297 2928
rect 3055 2914 3070 2918
rect 2973 2912 3070 2914
rect 3098 2912 3266 2924
rect 3282 2914 3297 2918
rect 3315 2915 3354 2934
rect 3373 2928 3380 2929
rect 3379 2921 3380 2928
rect 3363 2918 3364 2921
rect 3379 2918 3392 2921
rect 3315 2914 3345 2915
rect 3354 2914 3360 2915
rect 3363 2914 3392 2918
rect 3282 2913 3392 2914
rect 3282 2912 3398 2913
rect 2957 2904 3008 2912
rect 2957 2892 2982 2904
rect 2989 2892 3008 2904
rect 3039 2904 3089 2912
rect 3039 2896 3055 2904
rect 3062 2902 3089 2904
rect 3098 2902 3319 2912
rect 3062 2892 3319 2902
rect 3348 2904 3398 2912
rect 3348 2895 3364 2904
rect 2957 2884 3008 2892
rect 3055 2884 3319 2892
rect 3345 2892 3364 2895
rect 3371 2892 3398 2904
rect 3345 2884 3398 2892
rect 2973 2876 2974 2884
rect 2989 2876 3002 2884
rect 2973 2868 2989 2876
rect 2970 2861 2989 2864
rect 2970 2852 2992 2861
rect 2943 2842 2992 2852
rect 2943 2836 2973 2842
rect 2992 2837 2997 2842
rect 2915 2820 2989 2836
rect 3007 2828 3037 2884
rect 3072 2874 3280 2884
rect 3315 2880 3360 2884
rect 3363 2883 3364 2884
rect 3379 2883 3392 2884
rect 3098 2844 3287 2874
rect 3113 2841 3287 2844
rect 3106 2838 3287 2841
rect 2915 2818 2928 2820
rect 2943 2818 2977 2820
rect 2915 2802 2989 2818
rect 3016 2814 3029 2828
rect 3044 2814 3060 2830
rect 3106 2825 3117 2838
rect 2899 2780 2900 2796
rect 2915 2780 2928 2802
rect 2943 2780 2973 2802
rect 3016 2798 3078 2814
rect 3106 2807 3117 2823
rect 3122 2818 3132 2838
rect 3142 2818 3156 2838
rect 3159 2825 3168 2838
rect 3184 2825 3193 2838
rect 3122 2807 3156 2818
rect 3159 2807 3168 2823
rect 3184 2807 3193 2823
rect 3200 2818 3210 2838
rect 3220 2818 3234 2838
rect 3235 2825 3246 2838
rect 3200 2807 3234 2818
rect 3235 2807 3246 2823
rect 3292 2814 3308 2830
rect 3315 2828 3345 2880
rect 3379 2876 3380 2883
rect 3364 2868 3380 2876
rect 3351 2836 3364 2855
rect 3379 2836 3409 2852
rect 3351 2820 3425 2836
rect 3351 2818 3364 2820
rect 3379 2818 3413 2820
rect 3016 2796 3029 2798
rect 3044 2796 3078 2798
rect 3016 2780 3078 2796
rect 3122 2791 3138 2794
rect 3200 2791 3230 2802
rect 3278 2798 3324 2814
rect 3351 2802 3425 2818
rect 3278 2796 3312 2798
rect 3277 2780 3324 2796
rect 3351 2780 3364 2802
rect 3379 2780 3409 2802
rect 3436 2780 3437 2796
rect 3452 2780 3465 2940
rect 3495 2836 3508 2940
rect 3553 2918 3554 2928
rect 3569 2918 3582 2928
rect 3553 2914 3582 2918
rect 3587 2914 3617 2940
rect 3635 2926 3651 2928
rect 3723 2926 3776 2940
rect 3724 2924 3788 2926
rect 3831 2924 3846 2940
rect 3895 2937 3925 2940
rect 3895 2934 3931 2937
rect 3861 2926 3877 2928
rect 3635 2914 3650 2918
rect 3553 2912 3650 2914
rect 3678 2912 3846 2924
rect 3862 2914 3877 2918
rect 3895 2915 3934 2934
rect 3953 2928 3960 2929
rect 3959 2921 3960 2928
rect 3943 2918 3944 2921
rect 3959 2918 3972 2921
rect 3895 2914 3925 2915
rect 3934 2914 3940 2915
rect 3943 2914 3972 2918
rect 3862 2913 3972 2914
rect 3862 2912 3978 2913
rect 3537 2904 3588 2912
rect 3537 2892 3562 2904
rect 3569 2892 3588 2904
rect 3619 2904 3669 2912
rect 3619 2896 3635 2904
rect 3642 2902 3669 2904
rect 3678 2902 3899 2912
rect 3642 2892 3899 2902
rect 3928 2904 3978 2912
rect 3928 2895 3944 2904
rect 3537 2884 3588 2892
rect 3635 2884 3899 2892
rect 3925 2892 3944 2895
rect 3951 2892 3978 2904
rect 3925 2884 3978 2892
rect 3553 2876 3554 2884
rect 3569 2876 3582 2884
rect 3553 2868 3569 2876
rect 3550 2861 3569 2864
rect 3550 2852 3572 2861
rect 3523 2842 3572 2852
rect 3523 2836 3553 2842
rect 3572 2837 3577 2842
rect 3495 2820 3569 2836
rect 3587 2828 3617 2884
rect 3652 2874 3860 2884
rect 3895 2880 3940 2884
rect 3943 2883 3944 2884
rect 3959 2883 3972 2884
rect 3678 2844 3867 2874
rect 3693 2841 3867 2844
rect 3686 2838 3867 2841
rect 3495 2818 3508 2820
rect 3523 2818 3557 2820
rect 3495 2802 3569 2818
rect 3596 2814 3609 2828
rect 3624 2814 3640 2830
rect 3686 2825 3697 2838
rect 3479 2780 3480 2796
rect 3495 2780 3508 2802
rect 3523 2780 3553 2802
rect 3596 2798 3658 2814
rect 3686 2807 3697 2823
rect 3702 2818 3712 2838
rect 3722 2818 3736 2838
rect 3739 2825 3748 2838
rect 3764 2825 3773 2838
rect 3702 2807 3736 2818
rect 3739 2807 3748 2823
rect 3764 2807 3773 2823
rect 3780 2818 3790 2838
rect 3800 2818 3814 2838
rect 3815 2825 3826 2838
rect 3780 2807 3814 2818
rect 3815 2807 3826 2823
rect 3872 2814 3888 2830
rect 3895 2828 3925 2880
rect 3959 2876 3960 2883
rect 3944 2868 3960 2876
rect 3931 2836 3944 2855
rect 3959 2836 3989 2852
rect 3931 2820 4005 2836
rect 3931 2818 3944 2820
rect 3959 2818 3993 2820
rect 3596 2796 3609 2798
rect 3624 2796 3658 2798
rect 3596 2780 3658 2796
rect 3702 2791 3718 2794
rect 3780 2791 3810 2802
rect 3858 2798 3904 2814
rect 3931 2802 4005 2818
rect 3858 2796 3892 2798
rect 3857 2780 3904 2796
rect 3931 2780 3944 2802
rect 3959 2780 3989 2802
rect 4016 2780 4017 2796
rect 4032 2780 4045 2940
rect 4075 2836 4088 2940
rect 4133 2918 4134 2928
rect 4149 2918 4162 2928
rect 4133 2914 4162 2918
rect 4167 2914 4197 2940
rect 4215 2926 4231 2928
rect 4303 2926 4356 2940
rect 4304 2924 4368 2926
rect 4411 2924 4426 2940
rect 4475 2937 4505 2940
rect 4475 2934 4511 2937
rect 4441 2926 4457 2928
rect 4215 2914 4230 2918
rect 4133 2912 4230 2914
rect 4258 2912 4426 2924
rect 4442 2914 4457 2918
rect 4475 2915 4514 2934
rect 4533 2928 4540 2929
rect 4539 2921 4540 2928
rect 4523 2918 4524 2921
rect 4539 2918 4552 2921
rect 4475 2914 4505 2915
rect 4514 2914 4520 2915
rect 4523 2914 4552 2918
rect 4442 2913 4552 2914
rect 4442 2912 4558 2913
rect 4117 2904 4168 2912
rect 4117 2892 4142 2904
rect 4149 2892 4168 2904
rect 4199 2904 4249 2912
rect 4199 2896 4215 2904
rect 4222 2902 4249 2904
rect 4258 2902 4479 2912
rect 4222 2892 4479 2902
rect 4508 2904 4558 2912
rect 4508 2895 4524 2904
rect 4117 2884 4168 2892
rect 4215 2884 4479 2892
rect 4505 2892 4524 2895
rect 4531 2892 4558 2904
rect 4505 2884 4558 2892
rect 4133 2876 4134 2884
rect 4149 2876 4162 2884
rect 4133 2868 4149 2876
rect 4130 2861 4149 2864
rect 4130 2852 4152 2861
rect 4103 2842 4152 2852
rect 4103 2836 4133 2842
rect 4152 2837 4157 2842
rect 4075 2820 4149 2836
rect 4167 2828 4197 2884
rect 4232 2874 4440 2884
rect 4475 2880 4520 2884
rect 4523 2883 4524 2884
rect 4539 2883 4552 2884
rect 4258 2844 4447 2874
rect 4273 2841 4447 2844
rect 4266 2838 4447 2841
rect 4075 2818 4088 2820
rect 4103 2818 4137 2820
rect 4075 2802 4149 2818
rect 4176 2814 4189 2828
rect 4204 2814 4220 2830
rect 4266 2825 4277 2838
rect 4059 2780 4060 2796
rect 4075 2780 4088 2802
rect 4103 2780 4133 2802
rect 4176 2798 4238 2814
rect 4266 2807 4277 2823
rect 4282 2818 4292 2838
rect 4302 2818 4316 2838
rect 4319 2825 4328 2838
rect 4344 2825 4353 2838
rect 4282 2807 4316 2818
rect 4319 2807 4328 2823
rect 4344 2807 4353 2823
rect 4360 2818 4370 2838
rect 4380 2818 4394 2838
rect 4395 2825 4406 2838
rect 4360 2807 4394 2818
rect 4395 2807 4406 2823
rect 4452 2814 4468 2830
rect 4475 2828 4505 2880
rect 4539 2876 4540 2883
rect 4524 2868 4540 2876
rect 4511 2836 4524 2855
rect 4539 2836 4569 2852
rect 4511 2820 4585 2836
rect 4511 2818 4524 2820
rect 4539 2818 4573 2820
rect 4176 2796 4189 2798
rect 4204 2796 4238 2798
rect 4176 2780 4238 2796
rect 4282 2791 4298 2794
rect 4360 2791 4390 2802
rect 4438 2798 4484 2814
rect 4511 2802 4585 2818
rect 4438 2796 4472 2798
rect 4437 2780 4484 2796
rect 4511 2780 4524 2802
rect 4539 2780 4569 2802
rect 4596 2780 4597 2796
rect 4612 2780 4625 2940
rect -7 2772 34 2780
rect -7 2746 8 2772
rect 15 2746 34 2772
rect 98 2768 160 2780
rect 172 2768 247 2780
rect 305 2768 380 2780
rect 392 2768 423 2780
rect 429 2768 464 2780
rect 98 2766 260 2768
rect -7 2738 34 2746
rect 116 2742 129 2766
rect 144 2764 159 2766
rect -1 2728 0 2738
rect 15 2728 28 2738
rect 43 2728 73 2742
rect 116 2728 159 2742
rect 183 2739 190 2746
rect 193 2742 260 2766
rect 292 2766 464 2768
rect 262 2744 290 2748
rect 292 2744 372 2766
rect 393 2764 408 2766
rect 262 2742 372 2744
rect 193 2738 372 2742
rect 166 2728 196 2738
rect 198 2728 351 2738
rect 359 2728 389 2738
rect 393 2728 423 2742
rect 451 2728 464 2766
rect 536 2772 571 2780
rect 536 2746 537 2772
rect 544 2746 571 2772
rect 479 2728 509 2742
rect 536 2738 571 2746
rect 573 2772 614 2780
rect 573 2746 588 2772
rect 595 2746 614 2772
rect 678 2768 740 2780
rect 752 2768 827 2780
rect 885 2768 960 2780
rect 972 2768 1003 2780
rect 1009 2768 1044 2780
rect 678 2766 840 2768
rect 573 2738 614 2746
rect 696 2742 709 2766
rect 724 2764 739 2766
rect 536 2728 537 2738
rect 552 2728 565 2738
rect 579 2728 580 2738
rect 595 2728 608 2738
rect 623 2728 653 2742
rect 696 2728 739 2742
rect 763 2739 770 2746
rect 773 2742 840 2766
rect 872 2766 1044 2768
rect 842 2744 870 2748
rect 872 2744 952 2766
rect 973 2764 988 2766
rect 842 2742 952 2744
rect 773 2738 952 2742
rect 746 2728 776 2738
rect 778 2728 931 2738
rect 939 2728 969 2738
rect 973 2728 1003 2742
rect 1031 2728 1044 2766
rect 1116 2772 1151 2780
rect 1116 2746 1117 2772
rect 1124 2746 1151 2772
rect 1059 2728 1089 2742
rect 1116 2738 1151 2746
rect 1153 2772 1194 2780
rect 1153 2746 1168 2772
rect 1175 2746 1194 2772
rect 1258 2768 1320 2780
rect 1332 2768 1407 2780
rect 1465 2768 1540 2780
rect 1552 2768 1583 2780
rect 1589 2768 1624 2780
rect 1258 2766 1420 2768
rect 1153 2738 1194 2746
rect 1276 2742 1289 2766
rect 1304 2764 1319 2766
rect 1116 2728 1117 2738
rect 1132 2728 1145 2738
rect 1159 2728 1160 2738
rect 1175 2728 1188 2738
rect 1203 2728 1233 2742
rect 1276 2728 1319 2742
rect 1343 2739 1350 2746
rect 1353 2742 1420 2766
rect 1452 2766 1624 2768
rect 1422 2744 1450 2748
rect 1452 2744 1532 2766
rect 1553 2764 1568 2766
rect 1422 2742 1532 2744
rect 1353 2738 1532 2742
rect 1326 2728 1356 2738
rect 1358 2728 1511 2738
rect 1519 2728 1549 2738
rect 1553 2728 1583 2742
rect 1611 2728 1624 2766
rect 1696 2772 1731 2780
rect 1696 2746 1697 2772
rect 1704 2746 1731 2772
rect 1639 2728 1669 2742
rect 1696 2738 1731 2746
rect 1733 2772 1774 2780
rect 1733 2746 1748 2772
rect 1755 2746 1774 2772
rect 1838 2768 1900 2780
rect 1912 2768 1987 2780
rect 2045 2768 2120 2780
rect 2132 2768 2163 2780
rect 2169 2768 2204 2780
rect 1838 2766 2000 2768
rect 1733 2738 1774 2746
rect 1856 2742 1869 2766
rect 1884 2764 1899 2766
rect 1696 2728 1697 2738
rect 1712 2728 1725 2738
rect 1739 2728 1740 2738
rect 1755 2728 1768 2738
rect 1783 2728 1813 2742
rect 1856 2728 1899 2742
rect 1923 2739 1930 2746
rect 1933 2742 2000 2766
rect 2032 2766 2204 2768
rect 2002 2744 2030 2748
rect 2032 2744 2112 2766
rect 2133 2764 2148 2766
rect 2002 2742 2112 2744
rect 1933 2738 2112 2742
rect 1906 2728 1936 2738
rect 1938 2728 2091 2738
rect 2099 2728 2129 2738
rect 2133 2728 2163 2742
rect 2191 2728 2204 2766
rect 2276 2772 2311 2780
rect 2276 2746 2277 2772
rect 2284 2746 2311 2772
rect 2219 2728 2249 2742
rect 2276 2738 2311 2746
rect 2313 2772 2354 2780
rect 2313 2746 2328 2772
rect 2335 2746 2354 2772
rect 2418 2768 2480 2780
rect 2492 2768 2567 2780
rect 2625 2768 2700 2780
rect 2712 2768 2743 2780
rect 2749 2768 2784 2780
rect 2418 2766 2580 2768
rect 2313 2738 2354 2746
rect 2436 2742 2449 2766
rect 2464 2764 2479 2766
rect 2276 2728 2277 2738
rect 2292 2728 2305 2738
rect 2319 2728 2320 2738
rect 2335 2728 2348 2738
rect 2363 2728 2393 2742
rect 2436 2728 2479 2742
rect 2503 2739 2510 2746
rect 2513 2742 2580 2766
rect 2612 2766 2784 2768
rect 2582 2744 2610 2748
rect 2612 2744 2692 2766
rect 2713 2764 2728 2766
rect 2582 2742 2692 2744
rect 2513 2738 2692 2742
rect 2486 2728 2516 2738
rect 2518 2728 2671 2738
rect 2679 2728 2709 2738
rect 2713 2728 2743 2742
rect 2771 2728 2784 2766
rect 2856 2772 2891 2780
rect 2856 2746 2857 2772
rect 2864 2746 2891 2772
rect 2799 2728 2829 2742
rect 2856 2738 2891 2746
rect 2893 2772 2934 2780
rect 2893 2746 2908 2772
rect 2915 2746 2934 2772
rect 2998 2768 3060 2780
rect 3072 2768 3147 2780
rect 3205 2768 3280 2780
rect 3292 2768 3323 2780
rect 3329 2768 3364 2780
rect 2998 2766 3160 2768
rect 2893 2738 2934 2746
rect 3016 2742 3029 2766
rect 3044 2764 3059 2766
rect 2856 2728 2857 2738
rect 2872 2728 2885 2738
rect 2899 2728 2900 2738
rect 2915 2728 2928 2738
rect 2943 2728 2973 2742
rect 3016 2728 3059 2742
rect 3083 2739 3090 2746
rect 3093 2742 3160 2766
rect 3192 2766 3364 2768
rect 3162 2744 3190 2748
rect 3192 2744 3272 2766
rect 3293 2764 3308 2766
rect 3162 2742 3272 2744
rect 3093 2738 3272 2742
rect 3066 2728 3096 2738
rect 3098 2728 3251 2738
rect 3259 2728 3289 2738
rect 3293 2728 3323 2742
rect 3351 2728 3364 2766
rect 3436 2772 3471 2780
rect 3436 2746 3437 2772
rect 3444 2746 3471 2772
rect 3379 2728 3409 2742
rect 3436 2738 3471 2746
rect 3473 2772 3514 2780
rect 3473 2746 3488 2772
rect 3495 2746 3514 2772
rect 3578 2768 3640 2780
rect 3652 2768 3727 2780
rect 3785 2768 3860 2780
rect 3872 2768 3903 2780
rect 3909 2768 3944 2780
rect 3578 2766 3740 2768
rect 3473 2738 3514 2746
rect 3596 2742 3609 2766
rect 3624 2764 3639 2766
rect 3436 2728 3437 2738
rect 3452 2728 3465 2738
rect 3479 2728 3480 2738
rect 3495 2728 3508 2738
rect 3523 2728 3553 2742
rect 3596 2728 3639 2742
rect 3663 2739 3670 2746
rect 3673 2742 3740 2766
rect 3772 2766 3944 2768
rect 3742 2744 3770 2748
rect 3772 2744 3852 2766
rect 3873 2764 3888 2766
rect 3742 2742 3852 2744
rect 3673 2738 3852 2742
rect 3646 2728 3676 2738
rect 3678 2728 3831 2738
rect 3839 2728 3869 2738
rect 3873 2728 3903 2742
rect 3931 2728 3944 2766
rect 4016 2772 4051 2780
rect 4016 2746 4017 2772
rect 4024 2746 4051 2772
rect 3959 2728 3989 2742
rect 4016 2738 4051 2746
rect 4053 2772 4094 2780
rect 4053 2746 4068 2772
rect 4075 2746 4094 2772
rect 4158 2768 4220 2780
rect 4232 2768 4307 2780
rect 4365 2768 4440 2780
rect 4452 2768 4483 2780
rect 4489 2768 4524 2780
rect 4158 2766 4320 2768
rect 4053 2738 4094 2746
rect 4176 2742 4189 2766
rect 4204 2764 4219 2766
rect 4016 2728 4017 2738
rect 4032 2728 4045 2738
rect 4059 2728 4060 2738
rect 4075 2728 4088 2738
rect 4103 2728 4133 2742
rect 4176 2728 4219 2742
rect 4243 2739 4250 2746
rect 4253 2742 4320 2766
rect 4352 2766 4524 2768
rect 4322 2744 4350 2748
rect 4352 2744 4432 2766
rect 4453 2764 4468 2766
rect 4322 2742 4432 2744
rect 4253 2738 4432 2742
rect 4226 2728 4256 2738
rect 4258 2728 4411 2738
rect 4419 2728 4449 2738
rect 4453 2728 4483 2742
rect 4511 2728 4524 2766
rect 4596 2772 4631 2780
rect 4596 2746 4597 2772
rect 4604 2746 4631 2772
rect 4539 2728 4569 2742
rect 4596 2738 4631 2746
rect 4596 2728 4597 2738
rect 4612 2728 4625 2738
rect -1 2722 4625 2728
rect 0 2714 4625 2722
rect 15 2684 28 2714
rect 43 2696 73 2714
rect 116 2700 130 2714
rect 166 2700 386 2714
rect 117 2698 130 2700
rect 83 2686 98 2698
rect 80 2684 102 2686
rect 107 2684 137 2698
rect 198 2696 351 2700
rect 180 2684 372 2696
rect 415 2684 445 2698
rect 451 2684 464 2714
rect 479 2696 509 2714
rect 552 2684 565 2714
rect 595 2684 608 2714
rect 623 2696 653 2714
rect 696 2700 710 2714
rect 746 2700 966 2714
rect 697 2698 710 2700
rect 663 2686 678 2698
rect 660 2684 682 2686
rect 687 2684 717 2698
rect 778 2696 931 2700
rect 760 2684 952 2696
rect 995 2684 1025 2698
rect 1031 2684 1044 2714
rect 1059 2696 1089 2714
rect 1132 2684 1145 2714
rect 1175 2684 1188 2714
rect 1203 2696 1233 2714
rect 1276 2700 1290 2714
rect 1326 2700 1546 2714
rect 1277 2698 1290 2700
rect 1243 2686 1258 2698
rect 1240 2684 1262 2686
rect 1267 2684 1297 2698
rect 1358 2696 1511 2700
rect 1340 2684 1532 2696
rect 1575 2684 1605 2698
rect 1611 2684 1624 2714
rect 1639 2696 1669 2714
rect 1712 2684 1725 2714
rect 1755 2684 1768 2714
rect 1783 2696 1813 2714
rect 1856 2700 1870 2714
rect 1906 2700 2126 2714
rect 1857 2698 1870 2700
rect 1823 2686 1838 2698
rect 1820 2684 1842 2686
rect 1847 2684 1877 2698
rect 1938 2696 2091 2700
rect 1920 2684 2112 2696
rect 2155 2684 2185 2698
rect 2191 2684 2204 2714
rect 2219 2696 2249 2714
rect 2292 2684 2305 2714
rect 2335 2684 2348 2714
rect 2363 2696 2393 2714
rect 2436 2700 2450 2714
rect 2486 2700 2706 2714
rect 2437 2698 2450 2700
rect 2403 2686 2418 2698
rect 2400 2684 2422 2686
rect 2427 2684 2457 2698
rect 2518 2696 2671 2700
rect 2500 2684 2692 2696
rect 2735 2684 2765 2698
rect 2771 2684 2784 2714
rect 2799 2696 2829 2714
rect 2872 2684 2885 2714
rect 2915 2684 2928 2714
rect 2943 2696 2973 2714
rect 3016 2700 3030 2714
rect 3066 2700 3286 2714
rect 3017 2698 3030 2700
rect 2983 2686 2998 2698
rect 2980 2684 3002 2686
rect 3007 2684 3037 2698
rect 3098 2696 3251 2700
rect 3080 2684 3272 2696
rect 3315 2684 3345 2698
rect 3351 2684 3364 2714
rect 3379 2696 3409 2714
rect 3452 2684 3465 2714
rect 3495 2684 3508 2714
rect 3523 2696 3553 2714
rect 3596 2700 3610 2714
rect 3646 2700 3866 2714
rect 3597 2698 3610 2700
rect 3563 2686 3578 2698
rect 3560 2684 3582 2686
rect 3587 2684 3617 2698
rect 3678 2696 3831 2700
rect 3660 2684 3852 2696
rect 3895 2684 3925 2698
rect 3931 2684 3944 2714
rect 3959 2696 3989 2714
rect 4032 2684 4045 2714
rect 4075 2684 4088 2714
rect 4103 2696 4133 2714
rect 4176 2700 4190 2714
rect 4226 2700 4446 2714
rect 4177 2698 4190 2700
rect 4143 2686 4158 2698
rect 4140 2684 4162 2686
rect 4167 2684 4197 2698
rect 4258 2696 4411 2700
rect 4240 2684 4432 2696
rect 4475 2684 4505 2698
rect 4511 2684 4524 2714
rect 4539 2696 4569 2714
rect 4612 2684 4625 2714
rect 0 2670 4625 2684
rect 15 2566 28 2670
rect 73 2648 74 2658
rect 89 2648 102 2658
rect 73 2644 102 2648
rect 107 2644 137 2670
rect 155 2656 171 2658
rect 243 2656 296 2670
rect 244 2654 308 2656
rect 351 2654 366 2670
rect 415 2667 445 2670
rect 415 2664 451 2667
rect 381 2656 397 2658
rect 155 2644 170 2648
rect 73 2642 170 2644
rect 198 2642 366 2654
rect 382 2644 397 2648
rect 415 2645 454 2664
rect 473 2658 480 2659
rect 479 2651 480 2658
rect 463 2648 464 2651
rect 479 2648 492 2651
rect 415 2644 445 2645
rect 454 2644 460 2645
rect 463 2644 492 2648
rect 382 2643 492 2644
rect 382 2642 498 2643
rect 57 2634 108 2642
rect 57 2622 82 2634
rect 89 2622 108 2634
rect 139 2634 189 2642
rect 139 2626 155 2634
rect 162 2632 189 2634
rect 198 2632 419 2642
rect 162 2622 419 2632
rect 448 2634 498 2642
rect 448 2625 464 2634
rect 57 2614 108 2622
rect 155 2614 419 2622
rect 445 2622 464 2625
rect 471 2622 498 2634
rect 445 2614 498 2622
rect 73 2606 74 2614
rect 89 2606 102 2614
rect 73 2598 89 2606
rect 70 2591 89 2594
rect 70 2582 92 2591
rect 43 2572 92 2582
rect 43 2566 73 2572
rect 92 2567 97 2572
rect 15 2550 89 2566
rect 107 2558 137 2614
rect 172 2604 380 2614
rect 415 2610 460 2614
rect 463 2613 464 2614
rect 479 2613 492 2614
rect 198 2574 387 2604
rect 213 2571 387 2574
rect 206 2568 387 2571
rect 15 2548 28 2550
rect 43 2548 77 2550
rect 15 2532 89 2548
rect 116 2544 129 2558
rect 144 2544 160 2560
rect 206 2555 217 2568
rect -1 2510 0 2526
rect 15 2510 28 2532
rect 43 2510 73 2532
rect 116 2528 178 2544
rect 206 2537 217 2553
rect 222 2548 232 2568
rect 242 2548 256 2568
rect 259 2555 268 2568
rect 284 2555 293 2568
rect 222 2537 256 2548
rect 259 2537 268 2553
rect 284 2537 293 2553
rect 300 2548 310 2568
rect 320 2548 334 2568
rect 335 2555 346 2568
rect 300 2537 334 2548
rect 335 2537 346 2553
rect 392 2544 408 2560
rect 415 2558 445 2610
rect 479 2606 480 2613
rect 464 2598 480 2606
rect 451 2566 464 2585
rect 479 2566 509 2582
rect 451 2550 525 2566
rect 451 2548 464 2550
rect 479 2548 513 2550
rect 116 2526 129 2528
rect 144 2526 178 2528
rect 116 2510 178 2526
rect 222 2521 238 2524
rect 300 2521 330 2532
rect 378 2528 424 2544
rect 451 2532 525 2548
rect 378 2526 412 2528
rect 377 2510 424 2526
rect 451 2510 464 2532
rect 479 2510 509 2532
rect 536 2510 537 2526
rect 552 2510 565 2670
rect 595 2566 608 2670
rect 653 2648 654 2658
rect 669 2648 682 2658
rect 653 2644 682 2648
rect 687 2644 717 2670
rect 735 2656 751 2658
rect 823 2656 876 2670
rect 824 2654 888 2656
rect 931 2654 946 2670
rect 995 2667 1025 2670
rect 995 2664 1031 2667
rect 961 2656 977 2658
rect 735 2644 750 2648
rect 653 2642 750 2644
rect 778 2642 946 2654
rect 962 2644 977 2648
rect 995 2645 1034 2664
rect 1053 2658 1060 2659
rect 1059 2651 1060 2658
rect 1043 2648 1044 2651
rect 1059 2648 1072 2651
rect 995 2644 1025 2645
rect 1034 2644 1040 2645
rect 1043 2644 1072 2648
rect 962 2643 1072 2644
rect 962 2642 1078 2643
rect 637 2634 688 2642
rect 637 2622 662 2634
rect 669 2622 688 2634
rect 719 2634 769 2642
rect 719 2626 735 2634
rect 742 2632 769 2634
rect 778 2632 999 2642
rect 742 2622 999 2632
rect 1028 2634 1078 2642
rect 1028 2625 1044 2634
rect 637 2614 688 2622
rect 735 2614 999 2622
rect 1025 2622 1044 2625
rect 1051 2622 1078 2634
rect 1025 2614 1078 2622
rect 653 2606 654 2614
rect 669 2606 682 2614
rect 653 2598 669 2606
rect 650 2591 669 2594
rect 650 2582 672 2591
rect 623 2572 672 2582
rect 623 2566 653 2572
rect 672 2567 677 2572
rect 595 2550 669 2566
rect 687 2558 717 2614
rect 752 2604 960 2614
rect 995 2610 1040 2614
rect 1043 2613 1044 2614
rect 1059 2613 1072 2614
rect 778 2574 967 2604
rect 793 2571 967 2574
rect 786 2568 967 2571
rect 595 2548 608 2550
rect 623 2548 657 2550
rect 595 2532 669 2548
rect 696 2544 709 2558
rect 724 2544 740 2560
rect 786 2555 797 2568
rect 579 2510 580 2526
rect 595 2510 608 2532
rect 623 2510 653 2532
rect 696 2528 758 2544
rect 786 2537 797 2553
rect 802 2548 812 2568
rect 822 2548 836 2568
rect 839 2555 848 2568
rect 864 2555 873 2568
rect 802 2537 836 2548
rect 839 2537 848 2553
rect 864 2537 873 2553
rect 880 2548 890 2568
rect 900 2548 914 2568
rect 915 2555 926 2568
rect 880 2537 914 2548
rect 915 2537 926 2553
rect 972 2544 988 2560
rect 995 2558 1025 2610
rect 1059 2606 1060 2613
rect 1044 2598 1060 2606
rect 1031 2566 1044 2585
rect 1059 2566 1089 2582
rect 1031 2550 1105 2566
rect 1031 2548 1044 2550
rect 1059 2548 1093 2550
rect 696 2526 709 2528
rect 724 2526 758 2528
rect 696 2510 758 2526
rect 802 2521 818 2524
rect 880 2521 910 2532
rect 958 2528 1004 2544
rect 1031 2532 1105 2548
rect 958 2526 992 2528
rect 957 2510 1004 2526
rect 1031 2510 1044 2532
rect 1059 2510 1089 2532
rect 1116 2510 1117 2526
rect 1132 2510 1145 2670
rect 1175 2566 1188 2670
rect 1233 2648 1234 2658
rect 1249 2648 1262 2658
rect 1233 2644 1262 2648
rect 1267 2644 1297 2670
rect 1315 2656 1331 2658
rect 1403 2656 1456 2670
rect 1404 2654 1468 2656
rect 1511 2654 1526 2670
rect 1575 2667 1605 2670
rect 1575 2664 1611 2667
rect 1541 2656 1557 2658
rect 1315 2644 1330 2648
rect 1233 2642 1330 2644
rect 1358 2642 1526 2654
rect 1542 2644 1557 2648
rect 1575 2645 1614 2664
rect 1633 2658 1640 2659
rect 1639 2651 1640 2658
rect 1623 2648 1624 2651
rect 1639 2648 1652 2651
rect 1575 2644 1605 2645
rect 1614 2644 1620 2645
rect 1623 2644 1652 2648
rect 1542 2643 1652 2644
rect 1542 2642 1658 2643
rect 1217 2634 1268 2642
rect 1217 2622 1242 2634
rect 1249 2622 1268 2634
rect 1299 2634 1349 2642
rect 1299 2626 1315 2634
rect 1322 2632 1349 2634
rect 1358 2632 1579 2642
rect 1322 2622 1579 2632
rect 1608 2634 1658 2642
rect 1608 2625 1624 2634
rect 1217 2614 1268 2622
rect 1315 2614 1579 2622
rect 1605 2622 1624 2625
rect 1631 2622 1658 2634
rect 1605 2614 1658 2622
rect 1233 2606 1234 2614
rect 1249 2606 1262 2614
rect 1233 2598 1249 2606
rect 1230 2591 1249 2594
rect 1230 2582 1252 2591
rect 1203 2572 1252 2582
rect 1203 2566 1233 2572
rect 1252 2567 1257 2572
rect 1175 2550 1249 2566
rect 1267 2558 1297 2614
rect 1332 2604 1540 2614
rect 1575 2610 1620 2614
rect 1623 2613 1624 2614
rect 1639 2613 1652 2614
rect 1358 2574 1547 2604
rect 1373 2571 1547 2574
rect 1366 2568 1547 2571
rect 1175 2548 1188 2550
rect 1203 2548 1237 2550
rect 1175 2532 1249 2548
rect 1276 2544 1289 2558
rect 1304 2544 1320 2560
rect 1366 2555 1377 2568
rect 1159 2510 1160 2526
rect 1175 2510 1188 2532
rect 1203 2510 1233 2532
rect 1276 2528 1338 2544
rect 1366 2537 1377 2553
rect 1382 2548 1392 2568
rect 1402 2548 1416 2568
rect 1419 2555 1428 2568
rect 1444 2555 1453 2568
rect 1382 2537 1416 2548
rect 1419 2537 1428 2553
rect 1444 2537 1453 2553
rect 1460 2548 1470 2568
rect 1480 2548 1494 2568
rect 1495 2555 1506 2568
rect 1460 2537 1494 2548
rect 1495 2537 1506 2553
rect 1552 2544 1568 2560
rect 1575 2558 1605 2610
rect 1639 2606 1640 2613
rect 1624 2598 1640 2606
rect 1611 2566 1624 2585
rect 1639 2566 1669 2582
rect 1611 2550 1685 2566
rect 1611 2548 1624 2550
rect 1639 2548 1673 2550
rect 1276 2526 1289 2528
rect 1304 2526 1338 2528
rect 1276 2510 1338 2526
rect 1382 2521 1398 2524
rect 1460 2521 1490 2532
rect 1538 2528 1584 2544
rect 1611 2532 1685 2548
rect 1538 2526 1572 2528
rect 1537 2510 1584 2526
rect 1611 2510 1624 2532
rect 1639 2510 1669 2532
rect 1696 2510 1697 2526
rect 1712 2510 1725 2670
rect 1755 2566 1768 2670
rect 1813 2648 1814 2658
rect 1829 2648 1842 2658
rect 1813 2644 1842 2648
rect 1847 2644 1877 2670
rect 1895 2656 1911 2658
rect 1983 2656 2036 2670
rect 1984 2654 2048 2656
rect 2091 2654 2106 2670
rect 2155 2667 2185 2670
rect 2155 2664 2191 2667
rect 2121 2656 2137 2658
rect 1895 2644 1910 2648
rect 1813 2642 1910 2644
rect 1938 2642 2106 2654
rect 2122 2644 2137 2648
rect 2155 2645 2194 2664
rect 2213 2658 2220 2659
rect 2219 2651 2220 2658
rect 2203 2648 2204 2651
rect 2219 2648 2232 2651
rect 2155 2644 2185 2645
rect 2194 2644 2200 2645
rect 2203 2644 2232 2648
rect 2122 2643 2232 2644
rect 2122 2642 2238 2643
rect 1797 2634 1848 2642
rect 1797 2622 1822 2634
rect 1829 2622 1848 2634
rect 1879 2634 1929 2642
rect 1879 2626 1895 2634
rect 1902 2632 1929 2634
rect 1938 2632 2159 2642
rect 1902 2622 2159 2632
rect 2188 2634 2238 2642
rect 2188 2625 2204 2634
rect 1797 2614 1848 2622
rect 1895 2614 2159 2622
rect 2185 2622 2204 2625
rect 2211 2622 2238 2634
rect 2185 2614 2238 2622
rect 1813 2606 1814 2614
rect 1829 2606 1842 2614
rect 1813 2598 1829 2606
rect 1810 2591 1829 2594
rect 1810 2582 1832 2591
rect 1783 2572 1832 2582
rect 1783 2566 1813 2572
rect 1832 2567 1837 2572
rect 1755 2550 1829 2566
rect 1847 2558 1877 2614
rect 1912 2604 2120 2614
rect 2155 2610 2200 2614
rect 2203 2613 2204 2614
rect 2219 2613 2232 2614
rect 1938 2574 2127 2604
rect 1953 2571 2127 2574
rect 1946 2568 2127 2571
rect 1755 2548 1768 2550
rect 1783 2548 1817 2550
rect 1755 2532 1829 2548
rect 1856 2544 1869 2558
rect 1884 2544 1900 2560
rect 1946 2555 1957 2568
rect 1739 2510 1740 2526
rect 1755 2510 1768 2532
rect 1783 2510 1813 2532
rect 1856 2528 1918 2544
rect 1946 2537 1957 2553
rect 1962 2548 1972 2568
rect 1982 2548 1996 2568
rect 1999 2555 2008 2568
rect 2024 2555 2033 2568
rect 1962 2537 1996 2548
rect 1999 2537 2008 2553
rect 2024 2537 2033 2553
rect 2040 2548 2050 2568
rect 2060 2548 2074 2568
rect 2075 2555 2086 2568
rect 2040 2537 2074 2548
rect 2075 2537 2086 2553
rect 2132 2544 2148 2560
rect 2155 2558 2185 2610
rect 2219 2606 2220 2613
rect 2204 2598 2220 2606
rect 2191 2566 2204 2585
rect 2219 2566 2249 2582
rect 2191 2550 2265 2566
rect 2191 2548 2204 2550
rect 2219 2548 2253 2550
rect 1856 2526 1869 2528
rect 1884 2526 1918 2528
rect 1856 2510 1918 2526
rect 1962 2521 1978 2524
rect 2040 2521 2070 2532
rect 2118 2528 2164 2544
rect 2191 2532 2265 2548
rect 2118 2526 2152 2528
rect 2117 2510 2164 2526
rect 2191 2510 2204 2532
rect 2219 2510 2249 2532
rect 2276 2510 2277 2526
rect 2292 2510 2305 2670
rect 2335 2566 2348 2670
rect 2393 2648 2394 2658
rect 2409 2648 2422 2658
rect 2393 2644 2422 2648
rect 2427 2644 2457 2670
rect 2475 2656 2491 2658
rect 2563 2656 2616 2670
rect 2564 2654 2628 2656
rect 2671 2654 2686 2670
rect 2735 2667 2765 2670
rect 2735 2664 2771 2667
rect 2701 2656 2717 2658
rect 2475 2644 2490 2648
rect 2393 2642 2490 2644
rect 2518 2642 2686 2654
rect 2702 2644 2717 2648
rect 2735 2645 2774 2664
rect 2793 2658 2800 2659
rect 2799 2651 2800 2658
rect 2783 2648 2784 2651
rect 2799 2648 2812 2651
rect 2735 2644 2765 2645
rect 2774 2644 2780 2645
rect 2783 2644 2812 2648
rect 2702 2643 2812 2644
rect 2702 2642 2818 2643
rect 2377 2634 2428 2642
rect 2377 2622 2402 2634
rect 2409 2622 2428 2634
rect 2459 2634 2509 2642
rect 2459 2626 2475 2634
rect 2482 2632 2509 2634
rect 2518 2632 2739 2642
rect 2482 2622 2739 2632
rect 2768 2634 2818 2642
rect 2768 2625 2784 2634
rect 2377 2614 2428 2622
rect 2475 2614 2739 2622
rect 2765 2622 2784 2625
rect 2791 2622 2818 2634
rect 2765 2614 2818 2622
rect 2393 2606 2394 2614
rect 2409 2606 2422 2614
rect 2393 2598 2409 2606
rect 2390 2591 2409 2594
rect 2390 2582 2412 2591
rect 2363 2572 2412 2582
rect 2363 2566 2393 2572
rect 2412 2567 2417 2572
rect 2335 2550 2409 2566
rect 2427 2558 2457 2614
rect 2492 2604 2700 2614
rect 2735 2610 2780 2614
rect 2783 2613 2784 2614
rect 2799 2613 2812 2614
rect 2518 2574 2707 2604
rect 2533 2571 2707 2574
rect 2526 2568 2707 2571
rect 2335 2548 2348 2550
rect 2363 2548 2397 2550
rect 2335 2532 2409 2548
rect 2436 2544 2449 2558
rect 2464 2544 2480 2560
rect 2526 2555 2537 2568
rect 2319 2510 2320 2526
rect 2335 2510 2348 2532
rect 2363 2510 2393 2532
rect 2436 2528 2498 2544
rect 2526 2537 2537 2553
rect 2542 2548 2552 2568
rect 2562 2548 2576 2568
rect 2579 2555 2588 2568
rect 2604 2555 2613 2568
rect 2542 2537 2576 2548
rect 2579 2537 2588 2553
rect 2604 2537 2613 2553
rect 2620 2548 2630 2568
rect 2640 2548 2654 2568
rect 2655 2555 2666 2568
rect 2620 2537 2654 2548
rect 2655 2537 2666 2553
rect 2712 2544 2728 2560
rect 2735 2558 2765 2610
rect 2799 2606 2800 2613
rect 2784 2598 2800 2606
rect 2771 2566 2784 2585
rect 2799 2566 2829 2582
rect 2771 2550 2845 2566
rect 2771 2548 2784 2550
rect 2799 2548 2833 2550
rect 2436 2526 2449 2528
rect 2464 2526 2498 2528
rect 2436 2510 2498 2526
rect 2542 2521 2558 2524
rect 2620 2521 2650 2532
rect 2698 2528 2744 2544
rect 2771 2532 2845 2548
rect 2698 2526 2732 2528
rect 2697 2510 2744 2526
rect 2771 2510 2784 2532
rect 2799 2510 2829 2532
rect 2856 2510 2857 2526
rect 2872 2510 2885 2670
rect 2915 2566 2928 2670
rect 2973 2648 2974 2658
rect 2989 2648 3002 2658
rect 2973 2644 3002 2648
rect 3007 2644 3037 2670
rect 3055 2656 3071 2658
rect 3143 2656 3196 2670
rect 3144 2654 3208 2656
rect 3251 2654 3266 2670
rect 3315 2667 3345 2670
rect 3315 2664 3351 2667
rect 3281 2656 3297 2658
rect 3055 2644 3070 2648
rect 2973 2642 3070 2644
rect 3098 2642 3266 2654
rect 3282 2644 3297 2648
rect 3315 2645 3354 2664
rect 3373 2658 3380 2659
rect 3379 2651 3380 2658
rect 3363 2648 3364 2651
rect 3379 2648 3392 2651
rect 3315 2644 3345 2645
rect 3354 2644 3360 2645
rect 3363 2644 3392 2648
rect 3282 2643 3392 2644
rect 3282 2642 3398 2643
rect 2957 2634 3008 2642
rect 2957 2622 2982 2634
rect 2989 2622 3008 2634
rect 3039 2634 3089 2642
rect 3039 2626 3055 2634
rect 3062 2632 3089 2634
rect 3098 2632 3319 2642
rect 3062 2622 3319 2632
rect 3348 2634 3398 2642
rect 3348 2625 3364 2634
rect 2957 2614 3008 2622
rect 3055 2614 3319 2622
rect 3345 2622 3364 2625
rect 3371 2622 3398 2634
rect 3345 2614 3398 2622
rect 2973 2606 2974 2614
rect 2989 2606 3002 2614
rect 2973 2598 2989 2606
rect 2970 2591 2989 2594
rect 2970 2582 2992 2591
rect 2943 2572 2992 2582
rect 2943 2566 2973 2572
rect 2992 2567 2997 2572
rect 2915 2550 2989 2566
rect 3007 2558 3037 2614
rect 3072 2604 3280 2614
rect 3315 2610 3360 2614
rect 3363 2613 3364 2614
rect 3379 2613 3392 2614
rect 3098 2574 3287 2604
rect 3113 2571 3287 2574
rect 3106 2568 3287 2571
rect 2915 2548 2928 2550
rect 2943 2548 2977 2550
rect 2915 2532 2989 2548
rect 3016 2544 3029 2558
rect 3044 2544 3060 2560
rect 3106 2555 3117 2568
rect 2899 2510 2900 2526
rect 2915 2510 2928 2532
rect 2943 2510 2973 2532
rect 3016 2528 3078 2544
rect 3106 2537 3117 2553
rect 3122 2548 3132 2568
rect 3142 2548 3156 2568
rect 3159 2555 3168 2568
rect 3184 2555 3193 2568
rect 3122 2537 3156 2548
rect 3159 2537 3168 2553
rect 3184 2537 3193 2553
rect 3200 2548 3210 2568
rect 3220 2548 3234 2568
rect 3235 2555 3246 2568
rect 3200 2537 3234 2548
rect 3235 2537 3246 2553
rect 3292 2544 3308 2560
rect 3315 2558 3345 2610
rect 3379 2606 3380 2613
rect 3364 2598 3380 2606
rect 3351 2566 3364 2585
rect 3379 2566 3409 2582
rect 3351 2550 3425 2566
rect 3351 2548 3364 2550
rect 3379 2548 3413 2550
rect 3016 2526 3029 2528
rect 3044 2526 3078 2528
rect 3016 2510 3078 2526
rect 3122 2521 3138 2524
rect 3200 2521 3230 2532
rect 3278 2528 3324 2544
rect 3351 2532 3425 2548
rect 3278 2526 3312 2528
rect 3277 2510 3324 2526
rect 3351 2510 3364 2532
rect 3379 2510 3409 2532
rect 3436 2510 3437 2526
rect 3452 2510 3465 2670
rect 3495 2566 3508 2670
rect 3553 2648 3554 2658
rect 3569 2648 3582 2658
rect 3553 2644 3582 2648
rect 3587 2644 3617 2670
rect 3635 2656 3651 2658
rect 3723 2656 3776 2670
rect 3724 2654 3788 2656
rect 3831 2654 3846 2670
rect 3895 2667 3925 2670
rect 3895 2664 3931 2667
rect 3861 2656 3877 2658
rect 3635 2644 3650 2648
rect 3553 2642 3650 2644
rect 3678 2642 3846 2654
rect 3862 2644 3877 2648
rect 3895 2645 3934 2664
rect 3953 2658 3960 2659
rect 3959 2651 3960 2658
rect 3943 2648 3944 2651
rect 3959 2648 3972 2651
rect 3895 2644 3925 2645
rect 3934 2644 3940 2645
rect 3943 2644 3972 2648
rect 3862 2643 3972 2644
rect 3862 2642 3978 2643
rect 3537 2634 3588 2642
rect 3537 2622 3562 2634
rect 3569 2622 3588 2634
rect 3619 2634 3669 2642
rect 3619 2626 3635 2634
rect 3642 2632 3669 2634
rect 3678 2632 3899 2642
rect 3642 2622 3899 2632
rect 3928 2634 3978 2642
rect 3928 2625 3944 2634
rect 3537 2614 3588 2622
rect 3635 2614 3899 2622
rect 3925 2622 3944 2625
rect 3951 2622 3978 2634
rect 3925 2614 3978 2622
rect 3553 2606 3554 2614
rect 3569 2606 3582 2614
rect 3553 2598 3569 2606
rect 3550 2591 3569 2594
rect 3550 2582 3572 2591
rect 3523 2572 3572 2582
rect 3523 2566 3553 2572
rect 3572 2567 3577 2572
rect 3495 2550 3569 2566
rect 3587 2558 3617 2614
rect 3652 2604 3860 2614
rect 3895 2610 3940 2614
rect 3943 2613 3944 2614
rect 3959 2613 3972 2614
rect 3678 2574 3867 2604
rect 3693 2571 3867 2574
rect 3686 2568 3867 2571
rect 3495 2548 3508 2550
rect 3523 2548 3557 2550
rect 3495 2532 3569 2548
rect 3596 2544 3609 2558
rect 3624 2544 3640 2560
rect 3686 2555 3697 2568
rect 3479 2510 3480 2526
rect 3495 2510 3508 2532
rect 3523 2510 3553 2532
rect 3596 2528 3658 2544
rect 3686 2537 3697 2553
rect 3702 2548 3712 2568
rect 3722 2548 3736 2568
rect 3739 2555 3748 2568
rect 3764 2555 3773 2568
rect 3702 2537 3736 2548
rect 3739 2537 3748 2553
rect 3764 2537 3773 2553
rect 3780 2548 3790 2568
rect 3800 2548 3814 2568
rect 3815 2555 3826 2568
rect 3780 2537 3814 2548
rect 3815 2537 3826 2553
rect 3872 2544 3888 2560
rect 3895 2558 3925 2610
rect 3959 2606 3960 2613
rect 3944 2598 3960 2606
rect 3931 2566 3944 2585
rect 3959 2566 3989 2582
rect 3931 2550 4005 2566
rect 3931 2548 3944 2550
rect 3959 2548 3993 2550
rect 3596 2526 3609 2528
rect 3624 2526 3658 2528
rect 3596 2510 3658 2526
rect 3702 2521 3718 2524
rect 3780 2521 3810 2532
rect 3858 2528 3904 2544
rect 3931 2532 4005 2548
rect 3858 2526 3892 2528
rect 3857 2510 3904 2526
rect 3931 2510 3944 2532
rect 3959 2510 3989 2532
rect 4016 2510 4017 2526
rect 4032 2510 4045 2670
rect 4075 2566 4088 2670
rect 4133 2648 4134 2658
rect 4149 2648 4162 2658
rect 4133 2644 4162 2648
rect 4167 2644 4197 2670
rect 4215 2656 4231 2658
rect 4303 2656 4356 2670
rect 4304 2654 4368 2656
rect 4411 2654 4426 2670
rect 4475 2667 4505 2670
rect 4475 2664 4511 2667
rect 4441 2656 4457 2658
rect 4215 2644 4230 2648
rect 4133 2642 4230 2644
rect 4258 2642 4426 2654
rect 4442 2644 4457 2648
rect 4475 2645 4514 2664
rect 4533 2658 4540 2659
rect 4539 2651 4540 2658
rect 4523 2648 4524 2651
rect 4539 2648 4552 2651
rect 4475 2644 4505 2645
rect 4514 2644 4520 2645
rect 4523 2644 4552 2648
rect 4442 2643 4552 2644
rect 4442 2642 4558 2643
rect 4117 2634 4168 2642
rect 4117 2622 4142 2634
rect 4149 2622 4168 2634
rect 4199 2634 4249 2642
rect 4199 2626 4215 2634
rect 4222 2632 4249 2634
rect 4258 2632 4479 2642
rect 4222 2622 4479 2632
rect 4508 2634 4558 2642
rect 4508 2625 4524 2634
rect 4117 2614 4168 2622
rect 4215 2614 4479 2622
rect 4505 2622 4524 2625
rect 4531 2622 4558 2634
rect 4505 2614 4558 2622
rect 4133 2606 4134 2614
rect 4149 2606 4162 2614
rect 4133 2598 4149 2606
rect 4130 2591 4149 2594
rect 4130 2582 4152 2591
rect 4103 2572 4152 2582
rect 4103 2566 4133 2572
rect 4152 2567 4157 2572
rect 4075 2550 4149 2566
rect 4167 2558 4197 2614
rect 4232 2604 4440 2614
rect 4475 2610 4520 2614
rect 4523 2613 4524 2614
rect 4539 2613 4552 2614
rect 4258 2574 4447 2604
rect 4273 2571 4447 2574
rect 4266 2568 4447 2571
rect 4075 2548 4088 2550
rect 4103 2548 4137 2550
rect 4075 2532 4149 2548
rect 4176 2544 4189 2558
rect 4204 2544 4220 2560
rect 4266 2555 4277 2568
rect 4059 2510 4060 2526
rect 4075 2510 4088 2532
rect 4103 2510 4133 2532
rect 4176 2528 4238 2544
rect 4266 2537 4277 2553
rect 4282 2548 4292 2568
rect 4302 2548 4316 2568
rect 4319 2555 4328 2568
rect 4344 2555 4353 2568
rect 4282 2537 4316 2548
rect 4319 2537 4328 2553
rect 4344 2537 4353 2553
rect 4360 2548 4370 2568
rect 4380 2548 4394 2568
rect 4395 2555 4406 2568
rect 4360 2537 4394 2548
rect 4395 2537 4406 2553
rect 4452 2544 4468 2560
rect 4475 2558 4505 2610
rect 4539 2606 4540 2613
rect 4524 2598 4540 2606
rect 4511 2566 4524 2585
rect 4539 2566 4569 2582
rect 4511 2550 4585 2566
rect 4511 2548 4524 2550
rect 4539 2548 4573 2550
rect 4176 2526 4189 2528
rect 4204 2526 4238 2528
rect 4176 2510 4238 2526
rect 4282 2521 4298 2524
rect 4360 2521 4390 2532
rect 4438 2528 4484 2544
rect 4511 2532 4585 2548
rect 4438 2526 4472 2528
rect 4437 2510 4484 2526
rect 4511 2510 4524 2532
rect 4539 2510 4569 2532
rect 4596 2510 4597 2526
rect 4612 2510 4625 2670
rect -7 2502 34 2510
rect -7 2476 8 2502
rect 15 2476 34 2502
rect 98 2498 160 2510
rect 172 2498 247 2510
rect 305 2498 380 2510
rect 392 2498 423 2510
rect 429 2498 464 2510
rect 98 2496 260 2498
rect -7 2468 34 2476
rect 116 2472 129 2496
rect 144 2494 159 2496
rect -1 2458 0 2468
rect 15 2458 28 2468
rect 43 2458 73 2472
rect 116 2458 159 2472
rect 183 2469 190 2476
rect 193 2472 260 2496
rect 292 2496 464 2498
rect 262 2474 290 2478
rect 292 2474 372 2496
rect 393 2494 408 2496
rect 262 2472 372 2474
rect 193 2468 372 2472
rect 166 2458 196 2468
rect 198 2458 351 2468
rect 359 2458 389 2468
rect 393 2458 423 2472
rect 451 2458 464 2496
rect 536 2502 571 2510
rect 536 2476 537 2502
rect 544 2476 571 2502
rect 479 2458 509 2472
rect 536 2468 571 2476
rect 573 2502 614 2510
rect 573 2476 588 2502
rect 595 2476 614 2502
rect 678 2498 740 2510
rect 752 2498 827 2510
rect 885 2498 960 2510
rect 972 2498 1003 2510
rect 1009 2498 1044 2510
rect 678 2496 840 2498
rect 573 2468 614 2476
rect 696 2472 709 2496
rect 724 2494 739 2496
rect 536 2458 537 2468
rect 552 2458 565 2468
rect 579 2458 580 2468
rect 595 2458 608 2468
rect 623 2458 653 2472
rect 696 2458 739 2472
rect 763 2469 770 2476
rect 773 2472 840 2496
rect 872 2496 1044 2498
rect 842 2474 870 2478
rect 872 2474 952 2496
rect 973 2494 988 2496
rect 842 2472 952 2474
rect 773 2468 952 2472
rect 746 2458 776 2468
rect 778 2458 931 2468
rect 939 2458 969 2468
rect 973 2458 1003 2472
rect 1031 2458 1044 2496
rect 1116 2502 1151 2510
rect 1116 2476 1117 2502
rect 1124 2476 1151 2502
rect 1059 2458 1089 2472
rect 1116 2468 1151 2476
rect 1153 2502 1194 2510
rect 1153 2476 1168 2502
rect 1175 2476 1194 2502
rect 1258 2498 1320 2510
rect 1332 2498 1407 2510
rect 1465 2498 1540 2510
rect 1552 2498 1583 2510
rect 1589 2498 1624 2510
rect 1258 2496 1420 2498
rect 1153 2468 1194 2476
rect 1276 2472 1289 2496
rect 1304 2494 1319 2496
rect 1116 2458 1117 2468
rect 1132 2458 1145 2468
rect 1159 2458 1160 2468
rect 1175 2458 1188 2468
rect 1203 2458 1233 2472
rect 1276 2458 1319 2472
rect 1343 2469 1350 2476
rect 1353 2472 1420 2496
rect 1452 2496 1624 2498
rect 1422 2474 1450 2478
rect 1452 2474 1532 2496
rect 1553 2494 1568 2496
rect 1422 2472 1532 2474
rect 1353 2468 1532 2472
rect 1326 2458 1356 2468
rect 1358 2458 1511 2468
rect 1519 2458 1549 2468
rect 1553 2458 1583 2472
rect 1611 2458 1624 2496
rect 1696 2502 1731 2510
rect 1696 2476 1697 2502
rect 1704 2476 1731 2502
rect 1639 2458 1669 2472
rect 1696 2468 1731 2476
rect 1733 2502 1774 2510
rect 1733 2476 1748 2502
rect 1755 2476 1774 2502
rect 1838 2498 1900 2510
rect 1912 2498 1987 2510
rect 2045 2498 2120 2510
rect 2132 2498 2163 2510
rect 2169 2498 2204 2510
rect 1838 2496 2000 2498
rect 1733 2468 1774 2476
rect 1856 2472 1869 2496
rect 1884 2494 1899 2496
rect 1696 2458 1697 2468
rect 1712 2458 1725 2468
rect 1739 2458 1740 2468
rect 1755 2458 1768 2468
rect 1783 2458 1813 2472
rect 1856 2458 1899 2472
rect 1923 2469 1930 2476
rect 1933 2472 2000 2496
rect 2032 2496 2204 2498
rect 2002 2474 2030 2478
rect 2032 2474 2112 2496
rect 2133 2494 2148 2496
rect 2002 2472 2112 2474
rect 1933 2468 2112 2472
rect 1906 2458 1936 2468
rect 1938 2458 2091 2468
rect 2099 2458 2129 2468
rect 2133 2458 2163 2472
rect 2191 2458 2204 2496
rect 2276 2502 2311 2510
rect 2276 2476 2277 2502
rect 2284 2476 2311 2502
rect 2219 2458 2249 2472
rect 2276 2468 2311 2476
rect 2313 2502 2354 2510
rect 2313 2476 2328 2502
rect 2335 2476 2354 2502
rect 2418 2498 2480 2510
rect 2492 2498 2567 2510
rect 2625 2498 2700 2510
rect 2712 2498 2743 2510
rect 2749 2498 2784 2510
rect 2418 2496 2580 2498
rect 2313 2468 2354 2476
rect 2436 2472 2449 2496
rect 2464 2494 2479 2496
rect 2276 2458 2277 2468
rect 2292 2458 2305 2468
rect 2319 2458 2320 2468
rect 2335 2458 2348 2468
rect 2363 2458 2393 2472
rect 2436 2458 2479 2472
rect 2503 2469 2510 2476
rect 2513 2472 2580 2496
rect 2612 2496 2784 2498
rect 2582 2474 2610 2478
rect 2612 2474 2692 2496
rect 2713 2494 2728 2496
rect 2582 2472 2692 2474
rect 2513 2468 2692 2472
rect 2486 2458 2516 2468
rect 2518 2458 2671 2468
rect 2679 2458 2709 2468
rect 2713 2458 2743 2472
rect 2771 2458 2784 2496
rect 2856 2502 2891 2510
rect 2856 2476 2857 2502
rect 2864 2476 2891 2502
rect 2799 2458 2829 2472
rect 2856 2468 2891 2476
rect 2893 2502 2934 2510
rect 2893 2476 2908 2502
rect 2915 2476 2934 2502
rect 2998 2498 3060 2510
rect 3072 2498 3147 2510
rect 3205 2498 3280 2510
rect 3292 2498 3323 2510
rect 3329 2498 3364 2510
rect 2998 2496 3160 2498
rect 2893 2468 2934 2476
rect 3016 2472 3029 2496
rect 3044 2494 3059 2496
rect 2856 2458 2857 2468
rect 2872 2458 2885 2468
rect 2899 2458 2900 2468
rect 2915 2458 2928 2468
rect 2943 2458 2973 2472
rect 3016 2458 3059 2472
rect 3083 2469 3090 2476
rect 3093 2472 3160 2496
rect 3192 2496 3364 2498
rect 3162 2474 3190 2478
rect 3192 2474 3272 2496
rect 3293 2494 3308 2496
rect 3162 2472 3272 2474
rect 3093 2468 3272 2472
rect 3066 2458 3096 2468
rect 3098 2458 3251 2468
rect 3259 2458 3289 2468
rect 3293 2458 3323 2472
rect 3351 2458 3364 2496
rect 3436 2502 3471 2510
rect 3436 2476 3437 2502
rect 3444 2476 3471 2502
rect 3379 2458 3409 2472
rect 3436 2468 3471 2476
rect 3473 2502 3514 2510
rect 3473 2476 3488 2502
rect 3495 2476 3514 2502
rect 3578 2498 3640 2510
rect 3652 2498 3727 2510
rect 3785 2498 3860 2510
rect 3872 2498 3903 2510
rect 3909 2498 3944 2510
rect 3578 2496 3740 2498
rect 3473 2468 3514 2476
rect 3596 2472 3609 2496
rect 3624 2494 3639 2496
rect 3436 2458 3437 2468
rect 3452 2458 3465 2468
rect 3479 2458 3480 2468
rect 3495 2458 3508 2468
rect 3523 2458 3553 2472
rect 3596 2458 3639 2472
rect 3663 2469 3670 2476
rect 3673 2472 3740 2496
rect 3772 2496 3944 2498
rect 3742 2474 3770 2478
rect 3772 2474 3852 2496
rect 3873 2494 3888 2496
rect 3742 2472 3852 2474
rect 3673 2468 3852 2472
rect 3646 2458 3676 2468
rect 3678 2458 3831 2468
rect 3839 2458 3869 2468
rect 3873 2458 3903 2472
rect 3931 2458 3944 2496
rect 4016 2502 4051 2510
rect 4016 2476 4017 2502
rect 4024 2476 4051 2502
rect 3959 2458 3989 2472
rect 4016 2468 4051 2476
rect 4053 2502 4094 2510
rect 4053 2476 4068 2502
rect 4075 2476 4094 2502
rect 4158 2498 4220 2510
rect 4232 2498 4307 2510
rect 4365 2498 4440 2510
rect 4452 2498 4483 2510
rect 4489 2498 4524 2510
rect 4158 2496 4320 2498
rect 4053 2468 4094 2476
rect 4176 2472 4189 2496
rect 4204 2494 4219 2496
rect 4016 2458 4017 2468
rect 4032 2458 4045 2468
rect 4059 2458 4060 2468
rect 4075 2458 4088 2468
rect 4103 2458 4133 2472
rect 4176 2458 4219 2472
rect 4243 2469 4250 2476
rect 4253 2472 4320 2496
rect 4352 2496 4524 2498
rect 4322 2474 4350 2478
rect 4352 2474 4432 2496
rect 4453 2494 4468 2496
rect 4322 2472 4432 2474
rect 4253 2468 4432 2472
rect 4226 2458 4256 2468
rect 4258 2458 4411 2468
rect 4419 2458 4449 2468
rect 4453 2458 4483 2472
rect 4511 2458 4524 2496
rect 4596 2502 4631 2510
rect 4596 2476 4597 2502
rect 4604 2476 4631 2502
rect 4539 2458 4569 2472
rect 4596 2468 4631 2476
rect 4596 2458 4597 2468
rect 4612 2458 4625 2468
rect -1 2452 4625 2458
rect 0 2444 4625 2452
rect 15 2414 28 2444
rect 43 2426 73 2444
rect 116 2430 130 2444
rect 166 2430 386 2444
rect 117 2428 130 2430
rect 83 2416 98 2428
rect 80 2414 102 2416
rect 107 2414 137 2428
rect 198 2426 351 2430
rect 180 2414 372 2426
rect 415 2414 445 2428
rect 451 2414 464 2444
rect 479 2426 509 2444
rect 552 2414 565 2444
rect 595 2414 608 2444
rect 623 2426 653 2444
rect 696 2430 710 2444
rect 746 2430 966 2444
rect 697 2428 710 2430
rect 663 2416 678 2428
rect 660 2414 682 2416
rect 687 2414 717 2428
rect 778 2426 931 2430
rect 760 2414 952 2426
rect 995 2414 1025 2428
rect 1031 2414 1044 2444
rect 1059 2426 1089 2444
rect 1132 2414 1145 2444
rect 1175 2414 1188 2444
rect 1203 2426 1233 2444
rect 1276 2430 1290 2444
rect 1326 2430 1546 2444
rect 1277 2428 1290 2430
rect 1243 2416 1258 2428
rect 1240 2414 1262 2416
rect 1267 2414 1297 2428
rect 1358 2426 1511 2430
rect 1340 2414 1532 2426
rect 1575 2414 1605 2428
rect 1611 2414 1624 2444
rect 1639 2426 1669 2444
rect 1712 2414 1725 2444
rect 1755 2414 1768 2444
rect 1783 2426 1813 2444
rect 1856 2430 1870 2444
rect 1906 2430 2126 2444
rect 1857 2428 1870 2430
rect 1823 2416 1838 2428
rect 1820 2414 1842 2416
rect 1847 2414 1877 2428
rect 1938 2426 2091 2430
rect 1920 2414 2112 2426
rect 2155 2414 2185 2428
rect 2191 2414 2204 2444
rect 2219 2426 2249 2444
rect 2292 2414 2305 2444
rect 2335 2414 2348 2444
rect 2363 2426 2393 2444
rect 2436 2430 2450 2444
rect 2486 2430 2706 2444
rect 2437 2428 2450 2430
rect 2403 2416 2418 2428
rect 2400 2414 2422 2416
rect 2427 2414 2457 2428
rect 2518 2426 2671 2430
rect 2500 2414 2692 2426
rect 2735 2414 2765 2428
rect 2771 2414 2784 2444
rect 2799 2426 2829 2444
rect 2872 2414 2885 2444
rect 2915 2414 2928 2444
rect 2943 2426 2973 2444
rect 3016 2430 3030 2444
rect 3066 2430 3286 2444
rect 3017 2428 3030 2430
rect 2983 2416 2998 2428
rect 2980 2414 3002 2416
rect 3007 2414 3037 2428
rect 3098 2426 3251 2430
rect 3080 2414 3272 2426
rect 3315 2414 3345 2428
rect 3351 2414 3364 2444
rect 3379 2426 3409 2444
rect 3452 2414 3465 2444
rect 3495 2414 3508 2444
rect 3523 2426 3553 2444
rect 3596 2430 3610 2444
rect 3646 2430 3866 2444
rect 3597 2428 3610 2430
rect 3563 2416 3578 2428
rect 3560 2414 3582 2416
rect 3587 2414 3617 2428
rect 3678 2426 3831 2430
rect 3660 2414 3852 2426
rect 3895 2414 3925 2428
rect 3931 2414 3944 2444
rect 3959 2426 3989 2444
rect 4032 2414 4045 2444
rect 4075 2414 4088 2444
rect 4103 2426 4133 2444
rect 4176 2430 4190 2444
rect 4226 2430 4446 2444
rect 4177 2428 4190 2430
rect 4143 2416 4158 2428
rect 4140 2414 4162 2416
rect 4167 2414 4197 2428
rect 4258 2426 4411 2430
rect 4240 2414 4432 2426
rect 4475 2414 4505 2428
rect 4511 2414 4524 2444
rect 4539 2426 4569 2444
rect 4612 2414 4625 2444
rect 0 2400 4625 2414
rect 15 2296 28 2400
rect 73 2378 74 2388
rect 89 2378 102 2388
rect 73 2374 102 2378
rect 107 2374 137 2400
rect 155 2386 171 2388
rect 243 2386 296 2400
rect 244 2384 308 2386
rect 351 2384 366 2400
rect 415 2397 445 2400
rect 415 2394 451 2397
rect 381 2386 397 2388
rect 155 2374 170 2378
rect 73 2372 170 2374
rect 198 2372 366 2384
rect 382 2374 397 2378
rect 415 2375 454 2394
rect 473 2388 480 2389
rect 479 2381 480 2388
rect 463 2378 464 2381
rect 479 2378 492 2381
rect 415 2374 445 2375
rect 454 2374 460 2375
rect 463 2374 492 2378
rect 382 2373 492 2374
rect 382 2372 498 2373
rect 57 2364 108 2372
rect 57 2352 82 2364
rect 89 2352 108 2364
rect 139 2364 189 2372
rect 139 2356 155 2364
rect 162 2362 189 2364
rect 198 2362 419 2372
rect 162 2352 419 2362
rect 448 2364 498 2372
rect 448 2355 464 2364
rect 57 2344 108 2352
rect 155 2344 419 2352
rect 445 2352 464 2355
rect 471 2352 498 2364
rect 445 2344 498 2352
rect 73 2336 74 2344
rect 89 2336 102 2344
rect 73 2328 89 2336
rect 70 2321 89 2324
rect 70 2312 92 2321
rect 43 2302 92 2312
rect 43 2296 73 2302
rect 92 2297 97 2302
rect 15 2280 89 2296
rect 107 2288 137 2344
rect 172 2334 380 2344
rect 415 2340 460 2344
rect 463 2343 464 2344
rect 479 2343 492 2344
rect 198 2304 387 2334
rect 213 2301 387 2304
rect 206 2298 387 2301
rect 15 2278 28 2280
rect 43 2278 77 2280
rect 15 2262 89 2278
rect 116 2274 129 2288
rect 144 2274 160 2290
rect 206 2285 217 2298
rect -1 2240 0 2256
rect 15 2240 28 2262
rect 43 2240 73 2262
rect 116 2258 178 2274
rect 206 2267 217 2283
rect 222 2278 232 2298
rect 242 2278 256 2298
rect 259 2285 268 2298
rect 284 2285 293 2298
rect 222 2267 256 2278
rect 259 2267 268 2283
rect 284 2267 293 2283
rect 300 2278 310 2298
rect 320 2278 334 2298
rect 335 2285 346 2298
rect 300 2267 334 2278
rect 335 2267 346 2283
rect 392 2274 408 2290
rect 415 2288 445 2340
rect 479 2336 480 2343
rect 464 2328 480 2336
rect 451 2296 464 2315
rect 479 2296 509 2312
rect 451 2280 525 2296
rect 451 2278 464 2280
rect 479 2278 513 2280
rect 116 2256 129 2258
rect 144 2256 178 2258
rect 116 2240 178 2256
rect 222 2251 238 2254
rect 300 2251 330 2262
rect 378 2258 424 2274
rect 451 2262 525 2278
rect 378 2256 412 2258
rect 377 2240 424 2256
rect 451 2240 464 2262
rect 479 2240 509 2262
rect 536 2240 537 2256
rect 552 2240 565 2400
rect 595 2296 608 2400
rect 653 2378 654 2388
rect 669 2378 682 2388
rect 653 2374 682 2378
rect 687 2374 717 2400
rect 735 2386 751 2388
rect 823 2386 876 2400
rect 824 2384 888 2386
rect 931 2384 946 2400
rect 995 2397 1025 2400
rect 995 2394 1031 2397
rect 961 2386 977 2388
rect 735 2374 750 2378
rect 653 2372 750 2374
rect 778 2372 946 2384
rect 962 2374 977 2378
rect 995 2375 1034 2394
rect 1053 2388 1060 2389
rect 1059 2381 1060 2388
rect 1043 2378 1044 2381
rect 1059 2378 1072 2381
rect 995 2374 1025 2375
rect 1034 2374 1040 2375
rect 1043 2374 1072 2378
rect 962 2373 1072 2374
rect 962 2372 1078 2373
rect 637 2364 688 2372
rect 637 2352 662 2364
rect 669 2352 688 2364
rect 719 2364 769 2372
rect 719 2356 735 2364
rect 742 2362 769 2364
rect 778 2362 999 2372
rect 742 2352 999 2362
rect 1028 2364 1078 2372
rect 1028 2355 1044 2364
rect 637 2344 688 2352
rect 735 2344 999 2352
rect 1025 2352 1044 2355
rect 1051 2352 1078 2364
rect 1025 2344 1078 2352
rect 653 2336 654 2344
rect 669 2336 682 2344
rect 653 2328 669 2336
rect 650 2321 669 2324
rect 650 2312 672 2321
rect 623 2302 672 2312
rect 623 2296 653 2302
rect 672 2297 677 2302
rect 595 2280 669 2296
rect 687 2288 717 2344
rect 752 2334 960 2344
rect 995 2340 1040 2344
rect 1043 2343 1044 2344
rect 1059 2343 1072 2344
rect 778 2304 967 2334
rect 793 2301 967 2304
rect 786 2298 967 2301
rect 595 2278 608 2280
rect 623 2278 657 2280
rect 595 2262 669 2278
rect 696 2274 709 2288
rect 724 2274 740 2290
rect 786 2285 797 2298
rect 579 2240 580 2256
rect 595 2240 608 2262
rect 623 2240 653 2262
rect 696 2258 758 2274
rect 786 2267 797 2283
rect 802 2278 812 2298
rect 822 2278 836 2298
rect 839 2285 848 2298
rect 864 2285 873 2298
rect 802 2267 836 2278
rect 839 2267 848 2283
rect 864 2267 873 2283
rect 880 2278 890 2298
rect 900 2278 914 2298
rect 915 2285 926 2298
rect 880 2267 914 2278
rect 915 2267 926 2283
rect 972 2274 988 2290
rect 995 2288 1025 2340
rect 1059 2336 1060 2343
rect 1044 2328 1060 2336
rect 1031 2296 1044 2315
rect 1059 2296 1089 2312
rect 1031 2280 1105 2296
rect 1031 2278 1044 2280
rect 1059 2278 1093 2280
rect 696 2256 709 2258
rect 724 2256 758 2258
rect 696 2240 758 2256
rect 802 2251 818 2254
rect 880 2251 910 2262
rect 958 2258 1004 2274
rect 1031 2262 1105 2278
rect 958 2256 992 2258
rect 957 2240 1004 2256
rect 1031 2240 1044 2262
rect 1059 2240 1089 2262
rect 1116 2240 1117 2256
rect 1132 2240 1145 2400
rect 1175 2296 1188 2400
rect 1233 2378 1234 2388
rect 1249 2378 1262 2388
rect 1233 2374 1262 2378
rect 1267 2374 1297 2400
rect 1315 2386 1331 2388
rect 1403 2386 1456 2400
rect 1404 2384 1468 2386
rect 1511 2384 1526 2400
rect 1575 2397 1605 2400
rect 1575 2394 1611 2397
rect 1541 2386 1557 2388
rect 1315 2374 1330 2378
rect 1233 2372 1330 2374
rect 1358 2372 1526 2384
rect 1542 2374 1557 2378
rect 1575 2375 1614 2394
rect 1633 2388 1640 2389
rect 1639 2381 1640 2388
rect 1623 2378 1624 2381
rect 1639 2378 1652 2381
rect 1575 2374 1605 2375
rect 1614 2374 1620 2375
rect 1623 2374 1652 2378
rect 1542 2373 1652 2374
rect 1542 2372 1658 2373
rect 1217 2364 1268 2372
rect 1217 2352 1242 2364
rect 1249 2352 1268 2364
rect 1299 2364 1349 2372
rect 1299 2356 1315 2364
rect 1322 2362 1349 2364
rect 1358 2362 1579 2372
rect 1322 2352 1579 2362
rect 1608 2364 1658 2372
rect 1608 2355 1624 2364
rect 1217 2344 1268 2352
rect 1315 2344 1579 2352
rect 1605 2352 1624 2355
rect 1631 2352 1658 2364
rect 1605 2344 1658 2352
rect 1233 2336 1234 2344
rect 1249 2336 1262 2344
rect 1233 2328 1249 2336
rect 1230 2321 1249 2324
rect 1230 2312 1252 2321
rect 1203 2302 1252 2312
rect 1203 2296 1233 2302
rect 1252 2297 1257 2302
rect 1175 2280 1249 2296
rect 1267 2288 1297 2344
rect 1332 2334 1540 2344
rect 1575 2340 1620 2344
rect 1623 2343 1624 2344
rect 1639 2343 1652 2344
rect 1358 2304 1547 2334
rect 1373 2301 1547 2304
rect 1366 2298 1547 2301
rect 1175 2278 1188 2280
rect 1203 2278 1237 2280
rect 1175 2262 1249 2278
rect 1276 2274 1289 2288
rect 1304 2274 1320 2290
rect 1366 2285 1377 2298
rect 1159 2240 1160 2256
rect 1175 2240 1188 2262
rect 1203 2240 1233 2262
rect 1276 2258 1338 2274
rect 1366 2267 1377 2283
rect 1382 2278 1392 2298
rect 1402 2278 1416 2298
rect 1419 2285 1428 2298
rect 1444 2285 1453 2298
rect 1382 2267 1416 2278
rect 1419 2267 1428 2283
rect 1444 2267 1453 2283
rect 1460 2278 1470 2298
rect 1480 2278 1494 2298
rect 1495 2285 1506 2298
rect 1460 2267 1494 2278
rect 1495 2267 1506 2283
rect 1552 2274 1568 2290
rect 1575 2288 1605 2340
rect 1639 2336 1640 2343
rect 1624 2328 1640 2336
rect 1611 2296 1624 2315
rect 1639 2296 1669 2312
rect 1611 2280 1685 2296
rect 1611 2278 1624 2280
rect 1639 2278 1673 2280
rect 1276 2256 1289 2258
rect 1304 2256 1338 2258
rect 1276 2240 1338 2256
rect 1382 2251 1398 2254
rect 1460 2251 1490 2262
rect 1538 2258 1584 2274
rect 1611 2262 1685 2278
rect 1538 2256 1572 2258
rect 1537 2240 1584 2256
rect 1611 2240 1624 2262
rect 1639 2240 1669 2262
rect 1696 2240 1697 2256
rect 1712 2240 1725 2400
rect 1755 2296 1768 2400
rect 1813 2378 1814 2388
rect 1829 2378 1842 2388
rect 1813 2374 1842 2378
rect 1847 2374 1877 2400
rect 1895 2386 1911 2388
rect 1983 2386 2036 2400
rect 1984 2384 2048 2386
rect 2091 2384 2106 2400
rect 2155 2397 2185 2400
rect 2155 2394 2191 2397
rect 2121 2386 2137 2388
rect 1895 2374 1910 2378
rect 1813 2372 1910 2374
rect 1938 2372 2106 2384
rect 2122 2374 2137 2378
rect 2155 2375 2194 2394
rect 2213 2388 2220 2389
rect 2219 2381 2220 2388
rect 2203 2378 2204 2381
rect 2219 2378 2232 2381
rect 2155 2374 2185 2375
rect 2194 2374 2200 2375
rect 2203 2374 2232 2378
rect 2122 2373 2232 2374
rect 2122 2372 2238 2373
rect 1797 2364 1848 2372
rect 1797 2352 1822 2364
rect 1829 2352 1848 2364
rect 1879 2364 1929 2372
rect 1879 2356 1895 2364
rect 1902 2362 1929 2364
rect 1938 2362 2159 2372
rect 1902 2352 2159 2362
rect 2188 2364 2238 2372
rect 2188 2355 2204 2364
rect 1797 2344 1848 2352
rect 1895 2344 2159 2352
rect 2185 2352 2204 2355
rect 2211 2352 2238 2364
rect 2185 2344 2238 2352
rect 1813 2336 1814 2344
rect 1829 2336 1842 2344
rect 1813 2328 1829 2336
rect 1810 2321 1829 2324
rect 1810 2312 1832 2321
rect 1783 2302 1832 2312
rect 1783 2296 1813 2302
rect 1832 2297 1837 2302
rect 1755 2280 1829 2296
rect 1847 2288 1877 2344
rect 1912 2334 2120 2344
rect 2155 2340 2200 2344
rect 2203 2343 2204 2344
rect 2219 2343 2232 2344
rect 1938 2304 2127 2334
rect 1953 2301 2127 2304
rect 1946 2298 2127 2301
rect 1755 2278 1768 2280
rect 1783 2278 1817 2280
rect 1755 2262 1829 2278
rect 1856 2274 1869 2288
rect 1884 2274 1900 2290
rect 1946 2285 1957 2298
rect 1739 2240 1740 2256
rect 1755 2240 1768 2262
rect 1783 2240 1813 2262
rect 1856 2258 1918 2274
rect 1946 2267 1957 2283
rect 1962 2278 1972 2298
rect 1982 2278 1996 2298
rect 1999 2285 2008 2298
rect 2024 2285 2033 2298
rect 1962 2267 1996 2278
rect 1999 2267 2008 2283
rect 2024 2267 2033 2283
rect 2040 2278 2050 2298
rect 2060 2278 2074 2298
rect 2075 2285 2086 2298
rect 2040 2267 2074 2278
rect 2075 2267 2086 2283
rect 2132 2274 2148 2290
rect 2155 2288 2185 2340
rect 2219 2336 2220 2343
rect 2204 2328 2220 2336
rect 2191 2296 2204 2315
rect 2219 2296 2249 2312
rect 2191 2280 2265 2296
rect 2191 2278 2204 2280
rect 2219 2278 2253 2280
rect 1856 2256 1869 2258
rect 1884 2256 1918 2258
rect 1856 2240 1918 2256
rect 1962 2251 1978 2254
rect 2040 2251 2070 2262
rect 2118 2258 2164 2274
rect 2191 2262 2265 2278
rect 2118 2256 2152 2258
rect 2117 2240 2164 2256
rect 2191 2240 2204 2262
rect 2219 2240 2249 2262
rect 2276 2240 2277 2256
rect 2292 2240 2305 2400
rect 2335 2296 2348 2400
rect 2393 2378 2394 2388
rect 2409 2378 2422 2388
rect 2393 2374 2422 2378
rect 2427 2374 2457 2400
rect 2475 2386 2491 2388
rect 2563 2386 2616 2400
rect 2564 2384 2628 2386
rect 2671 2384 2686 2400
rect 2735 2397 2765 2400
rect 2735 2394 2771 2397
rect 2701 2386 2717 2388
rect 2475 2374 2490 2378
rect 2393 2372 2490 2374
rect 2518 2372 2686 2384
rect 2702 2374 2717 2378
rect 2735 2375 2774 2394
rect 2793 2388 2800 2389
rect 2799 2381 2800 2388
rect 2783 2378 2784 2381
rect 2799 2378 2812 2381
rect 2735 2374 2765 2375
rect 2774 2374 2780 2375
rect 2783 2374 2812 2378
rect 2702 2373 2812 2374
rect 2702 2372 2818 2373
rect 2377 2364 2428 2372
rect 2377 2352 2402 2364
rect 2409 2352 2428 2364
rect 2459 2364 2509 2372
rect 2459 2356 2475 2364
rect 2482 2362 2509 2364
rect 2518 2362 2739 2372
rect 2482 2352 2739 2362
rect 2768 2364 2818 2372
rect 2768 2355 2784 2364
rect 2377 2344 2428 2352
rect 2475 2344 2739 2352
rect 2765 2352 2784 2355
rect 2791 2352 2818 2364
rect 2765 2344 2818 2352
rect 2393 2336 2394 2344
rect 2409 2336 2422 2344
rect 2393 2328 2409 2336
rect 2390 2321 2409 2324
rect 2390 2312 2412 2321
rect 2363 2302 2412 2312
rect 2363 2296 2393 2302
rect 2412 2297 2417 2302
rect 2335 2280 2409 2296
rect 2427 2288 2457 2344
rect 2492 2334 2700 2344
rect 2735 2340 2780 2344
rect 2783 2343 2784 2344
rect 2799 2343 2812 2344
rect 2518 2304 2707 2334
rect 2533 2301 2707 2304
rect 2526 2298 2707 2301
rect 2335 2278 2348 2280
rect 2363 2278 2397 2280
rect 2335 2262 2409 2278
rect 2436 2274 2449 2288
rect 2464 2274 2480 2290
rect 2526 2285 2537 2298
rect 2319 2240 2320 2256
rect 2335 2240 2348 2262
rect 2363 2240 2393 2262
rect 2436 2258 2498 2274
rect 2526 2267 2537 2283
rect 2542 2278 2552 2298
rect 2562 2278 2576 2298
rect 2579 2285 2588 2298
rect 2604 2285 2613 2298
rect 2542 2267 2576 2278
rect 2579 2267 2588 2283
rect 2604 2267 2613 2283
rect 2620 2278 2630 2298
rect 2640 2278 2654 2298
rect 2655 2285 2666 2298
rect 2620 2267 2654 2278
rect 2655 2267 2666 2283
rect 2712 2274 2728 2290
rect 2735 2288 2765 2340
rect 2799 2336 2800 2343
rect 2784 2328 2800 2336
rect 2771 2296 2784 2315
rect 2799 2296 2829 2312
rect 2771 2280 2845 2296
rect 2771 2278 2784 2280
rect 2799 2278 2833 2280
rect 2436 2256 2449 2258
rect 2464 2256 2498 2258
rect 2436 2240 2498 2256
rect 2542 2251 2558 2254
rect 2620 2251 2650 2262
rect 2698 2258 2744 2274
rect 2771 2262 2845 2278
rect 2698 2256 2732 2258
rect 2697 2240 2744 2256
rect 2771 2240 2784 2262
rect 2799 2240 2829 2262
rect 2856 2240 2857 2256
rect 2872 2240 2885 2400
rect 2915 2296 2928 2400
rect 2973 2378 2974 2388
rect 2989 2378 3002 2388
rect 2973 2374 3002 2378
rect 3007 2374 3037 2400
rect 3055 2386 3071 2388
rect 3143 2386 3196 2400
rect 3144 2384 3208 2386
rect 3251 2384 3266 2400
rect 3315 2397 3345 2400
rect 3315 2394 3351 2397
rect 3281 2386 3297 2388
rect 3055 2374 3070 2378
rect 2973 2372 3070 2374
rect 3098 2372 3266 2384
rect 3282 2374 3297 2378
rect 3315 2375 3354 2394
rect 3373 2388 3380 2389
rect 3379 2381 3380 2388
rect 3363 2378 3364 2381
rect 3379 2378 3392 2381
rect 3315 2374 3345 2375
rect 3354 2374 3360 2375
rect 3363 2374 3392 2378
rect 3282 2373 3392 2374
rect 3282 2372 3398 2373
rect 2957 2364 3008 2372
rect 2957 2352 2982 2364
rect 2989 2352 3008 2364
rect 3039 2364 3089 2372
rect 3039 2356 3055 2364
rect 3062 2362 3089 2364
rect 3098 2362 3319 2372
rect 3062 2352 3319 2362
rect 3348 2364 3398 2372
rect 3348 2355 3364 2364
rect 2957 2344 3008 2352
rect 3055 2344 3319 2352
rect 3345 2352 3364 2355
rect 3371 2352 3398 2364
rect 3345 2344 3398 2352
rect 2973 2336 2974 2344
rect 2989 2336 3002 2344
rect 2973 2328 2989 2336
rect 2970 2321 2989 2324
rect 2970 2312 2992 2321
rect 2943 2302 2992 2312
rect 2943 2296 2973 2302
rect 2992 2297 2997 2302
rect 2915 2280 2989 2296
rect 3007 2288 3037 2344
rect 3072 2334 3280 2344
rect 3315 2340 3360 2344
rect 3363 2343 3364 2344
rect 3379 2343 3392 2344
rect 3098 2304 3287 2334
rect 3113 2301 3287 2304
rect 3106 2298 3287 2301
rect 2915 2278 2928 2280
rect 2943 2278 2977 2280
rect 2915 2262 2989 2278
rect 3016 2274 3029 2288
rect 3044 2274 3060 2290
rect 3106 2285 3117 2298
rect 2899 2240 2900 2256
rect 2915 2240 2928 2262
rect 2943 2240 2973 2262
rect 3016 2258 3078 2274
rect 3106 2267 3117 2283
rect 3122 2278 3132 2298
rect 3142 2278 3156 2298
rect 3159 2285 3168 2298
rect 3184 2285 3193 2298
rect 3122 2267 3156 2278
rect 3159 2267 3168 2283
rect 3184 2267 3193 2283
rect 3200 2278 3210 2298
rect 3220 2278 3234 2298
rect 3235 2285 3246 2298
rect 3200 2267 3234 2278
rect 3235 2267 3246 2283
rect 3292 2274 3308 2290
rect 3315 2288 3345 2340
rect 3379 2336 3380 2343
rect 3364 2328 3380 2336
rect 3351 2296 3364 2315
rect 3379 2296 3409 2312
rect 3351 2280 3425 2296
rect 3351 2278 3364 2280
rect 3379 2278 3413 2280
rect 3016 2256 3029 2258
rect 3044 2256 3078 2258
rect 3016 2240 3078 2256
rect 3122 2251 3138 2254
rect 3200 2251 3230 2262
rect 3278 2258 3324 2274
rect 3351 2262 3425 2278
rect 3278 2256 3312 2258
rect 3277 2240 3324 2256
rect 3351 2240 3364 2262
rect 3379 2240 3409 2262
rect 3436 2240 3437 2256
rect 3452 2240 3465 2400
rect 3495 2296 3508 2400
rect 3553 2378 3554 2388
rect 3569 2378 3582 2388
rect 3553 2374 3582 2378
rect 3587 2374 3617 2400
rect 3635 2386 3651 2388
rect 3723 2386 3776 2400
rect 3724 2384 3788 2386
rect 3831 2384 3846 2400
rect 3895 2397 3925 2400
rect 3895 2394 3931 2397
rect 3861 2386 3877 2388
rect 3635 2374 3650 2378
rect 3553 2372 3650 2374
rect 3678 2372 3846 2384
rect 3862 2374 3877 2378
rect 3895 2375 3934 2394
rect 3953 2388 3960 2389
rect 3959 2381 3960 2388
rect 3943 2378 3944 2381
rect 3959 2378 3972 2381
rect 3895 2374 3925 2375
rect 3934 2374 3940 2375
rect 3943 2374 3972 2378
rect 3862 2373 3972 2374
rect 3862 2372 3978 2373
rect 3537 2364 3588 2372
rect 3537 2352 3562 2364
rect 3569 2352 3588 2364
rect 3619 2364 3669 2372
rect 3619 2356 3635 2364
rect 3642 2362 3669 2364
rect 3678 2362 3899 2372
rect 3642 2352 3899 2362
rect 3928 2364 3978 2372
rect 3928 2355 3944 2364
rect 3537 2344 3588 2352
rect 3635 2344 3899 2352
rect 3925 2352 3944 2355
rect 3951 2352 3978 2364
rect 3925 2344 3978 2352
rect 3553 2336 3554 2344
rect 3569 2336 3582 2344
rect 3553 2328 3569 2336
rect 3550 2321 3569 2324
rect 3550 2312 3572 2321
rect 3523 2302 3572 2312
rect 3523 2296 3553 2302
rect 3572 2297 3577 2302
rect 3495 2280 3569 2296
rect 3587 2288 3617 2344
rect 3652 2334 3860 2344
rect 3895 2340 3940 2344
rect 3943 2343 3944 2344
rect 3959 2343 3972 2344
rect 3678 2304 3867 2334
rect 3693 2301 3867 2304
rect 3686 2298 3867 2301
rect 3495 2278 3508 2280
rect 3523 2278 3557 2280
rect 3495 2262 3569 2278
rect 3596 2274 3609 2288
rect 3624 2274 3640 2290
rect 3686 2285 3697 2298
rect 3479 2240 3480 2256
rect 3495 2240 3508 2262
rect 3523 2240 3553 2262
rect 3596 2258 3658 2274
rect 3686 2267 3697 2283
rect 3702 2278 3712 2298
rect 3722 2278 3736 2298
rect 3739 2285 3748 2298
rect 3764 2285 3773 2298
rect 3702 2267 3736 2278
rect 3739 2267 3748 2283
rect 3764 2267 3773 2283
rect 3780 2278 3790 2298
rect 3800 2278 3814 2298
rect 3815 2285 3826 2298
rect 3780 2267 3814 2278
rect 3815 2267 3826 2283
rect 3872 2274 3888 2290
rect 3895 2288 3925 2340
rect 3959 2336 3960 2343
rect 3944 2328 3960 2336
rect 3931 2296 3944 2315
rect 3959 2296 3989 2312
rect 3931 2280 4005 2296
rect 3931 2278 3944 2280
rect 3959 2278 3993 2280
rect 3596 2256 3609 2258
rect 3624 2256 3658 2258
rect 3596 2240 3658 2256
rect 3702 2251 3718 2254
rect 3780 2251 3810 2262
rect 3858 2258 3904 2274
rect 3931 2262 4005 2278
rect 3858 2256 3892 2258
rect 3857 2240 3904 2256
rect 3931 2240 3944 2262
rect 3959 2240 3989 2262
rect 4016 2240 4017 2256
rect 4032 2240 4045 2400
rect 4075 2296 4088 2400
rect 4133 2378 4134 2388
rect 4149 2378 4162 2388
rect 4133 2374 4162 2378
rect 4167 2374 4197 2400
rect 4215 2386 4231 2388
rect 4303 2386 4356 2400
rect 4304 2384 4368 2386
rect 4411 2384 4426 2400
rect 4475 2397 4505 2400
rect 4475 2394 4511 2397
rect 4441 2386 4457 2388
rect 4215 2374 4230 2378
rect 4133 2372 4230 2374
rect 4258 2372 4426 2384
rect 4442 2374 4457 2378
rect 4475 2375 4514 2394
rect 4533 2388 4540 2389
rect 4539 2381 4540 2388
rect 4523 2378 4524 2381
rect 4539 2378 4552 2381
rect 4475 2374 4505 2375
rect 4514 2374 4520 2375
rect 4523 2374 4552 2378
rect 4442 2373 4552 2374
rect 4442 2372 4558 2373
rect 4117 2364 4168 2372
rect 4117 2352 4142 2364
rect 4149 2352 4168 2364
rect 4199 2364 4249 2372
rect 4199 2356 4215 2364
rect 4222 2362 4249 2364
rect 4258 2362 4479 2372
rect 4222 2352 4479 2362
rect 4508 2364 4558 2372
rect 4508 2355 4524 2364
rect 4117 2344 4168 2352
rect 4215 2344 4479 2352
rect 4505 2352 4524 2355
rect 4531 2352 4558 2364
rect 4505 2344 4558 2352
rect 4133 2336 4134 2344
rect 4149 2336 4162 2344
rect 4133 2328 4149 2336
rect 4130 2321 4149 2324
rect 4130 2312 4152 2321
rect 4103 2302 4152 2312
rect 4103 2296 4133 2302
rect 4152 2297 4157 2302
rect 4075 2280 4149 2296
rect 4167 2288 4197 2344
rect 4232 2334 4440 2344
rect 4475 2340 4520 2344
rect 4523 2343 4524 2344
rect 4539 2343 4552 2344
rect 4258 2304 4447 2334
rect 4273 2301 4447 2304
rect 4266 2298 4447 2301
rect 4075 2278 4088 2280
rect 4103 2278 4137 2280
rect 4075 2262 4149 2278
rect 4176 2274 4189 2288
rect 4204 2274 4220 2290
rect 4266 2285 4277 2298
rect 4059 2240 4060 2256
rect 4075 2240 4088 2262
rect 4103 2240 4133 2262
rect 4176 2258 4238 2274
rect 4266 2267 4277 2283
rect 4282 2278 4292 2298
rect 4302 2278 4316 2298
rect 4319 2285 4328 2298
rect 4344 2285 4353 2298
rect 4282 2267 4316 2278
rect 4319 2267 4328 2283
rect 4344 2267 4353 2283
rect 4360 2278 4370 2298
rect 4380 2278 4394 2298
rect 4395 2285 4406 2298
rect 4360 2267 4394 2278
rect 4395 2267 4406 2283
rect 4452 2274 4468 2290
rect 4475 2288 4505 2340
rect 4539 2336 4540 2343
rect 4524 2328 4540 2336
rect 4511 2296 4524 2315
rect 4539 2296 4569 2312
rect 4511 2280 4585 2296
rect 4511 2278 4524 2280
rect 4539 2278 4573 2280
rect 4176 2256 4189 2258
rect 4204 2256 4238 2258
rect 4176 2240 4238 2256
rect 4282 2251 4298 2254
rect 4360 2251 4390 2262
rect 4438 2258 4484 2274
rect 4511 2262 4585 2278
rect 4438 2256 4472 2258
rect 4437 2240 4484 2256
rect 4511 2240 4524 2262
rect 4539 2240 4569 2262
rect 4596 2240 4597 2256
rect 4612 2240 4625 2400
rect -7 2232 34 2240
rect -7 2206 8 2232
rect 15 2206 34 2232
rect 98 2228 160 2240
rect 172 2228 247 2240
rect 305 2228 380 2240
rect 392 2228 423 2240
rect 429 2228 464 2240
rect 98 2226 260 2228
rect -7 2198 34 2206
rect 116 2202 129 2226
rect 144 2224 159 2226
rect -1 2188 0 2198
rect 15 2188 28 2198
rect 43 2188 73 2202
rect 116 2188 159 2202
rect 183 2199 190 2206
rect 193 2202 260 2226
rect 292 2226 464 2228
rect 262 2204 290 2208
rect 292 2204 372 2226
rect 393 2224 408 2226
rect 262 2202 372 2204
rect 193 2198 372 2202
rect 166 2188 196 2198
rect 198 2188 351 2198
rect 359 2188 389 2198
rect 393 2188 423 2202
rect 451 2188 464 2226
rect 536 2232 571 2240
rect 536 2206 537 2232
rect 544 2206 571 2232
rect 479 2188 509 2202
rect 536 2198 571 2206
rect 573 2232 614 2240
rect 573 2206 588 2232
rect 595 2206 614 2232
rect 678 2228 740 2240
rect 752 2228 827 2240
rect 885 2228 960 2240
rect 972 2228 1003 2240
rect 1009 2228 1044 2240
rect 678 2226 840 2228
rect 573 2198 614 2206
rect 696 2202 709 2226
rect 724 2224 739 2226
rect 536 2188 537 2198
rect 552 2188 565 2198
rect 579 2188 580 2198
rect 595 2188 608 2198
rect 623 2188 653 2202
rect 696 2188 739 2202
rect 763 2199 770 2206
rect 773 2202 840 2226
rect 872 2226 1044 2228
rect 842 2204 870 2208
rect 872 2204 952 2226
rect 973 2224 988 2226
rect 842 2202 952 2204
rect 773 2198 952 2202
rect 746 2188 776 2198
rect 778 2188 931 2198
rect 939 2188 969 2198
rect 973 2188 1003 2202
rect 1031 2188 1044 2226
rect 1116 2232 1151 2240
rect 1116 2206 1117 2232
rect 1124 2206 1151 2232
rect 1059 2188 1089 2202
rect 1116 2198 1151 2206
rect 1153 2232 1194 2240
rect 1153 2206 1168 2232
rect 1175 2206 1194 2232
rect 1258 2228 1320 2240
rect 1332 2228 1407 2240
rect 1465 2228 1540 2240
rect 1552 2228 1583 2240
rect 1589 2228 1624 2240
rect 1258 2226 1420 2228
rect 1153 2198 1194 2206
rect 1276 2202 1289 2226
rect 1304 2224 1319 2226
rect 1116 2188 1117 2198
rect 1132 2188 1145 2198
rect 1159 2188 1160 2198
rect 1175 2188 1188 2198
rect 1203 2188 1233 2202
rect 1276 2188 1319 2202
rect 1343 2199 1350 2206
rect 1353 2202 1420 2226
rect 1452 2226 1624 2228
rect 1422 2204 1450 2208
rect 1452 2204 1532 2226
rect 1553 2224 1568 2226
rect 1422 2202 1532 2204
rect 1353 2198 1532 2202
rect 1326 2188 1356 2198
rect 1358 2188 1511 2198
rect 1519 2188 1549 2198
rect 1553 2188 1583 2202
rect 1611 2188 1624 2226
rect 1696 2232 1731 2240
rect 1696 2206 1697 2232
rect 1704 2206 1731 2232
rect 1639 2188 1669 2202
rect 1696 2198 1731 2206
rect 1733 2232 1774 2240
rect 1733 2206 1748 2232
rect 1755 2206 1774 2232
rect 1838 2228 1900 2240
rect 1912 2228 1987 2240
rect 2045 2228 2120 2240
rect 2132 2228 2163 2240
rect 2169 2228 2204 2240
rect 1838 2226 2000 2228
rect 1733 2198 1774 2206
rect 1856 2202 1869 2226
rect 1884 2224 1899 2226
rect 1696 2188 1697 2198
rect 1712 2188 1725 2198
rect 1739 2188 1740 2198
rect 1755 2188 1768 2198
rect 1783 2188 1813 2202
rect 1856 2188 1899 2202
rect 1923 2199 1930 2206
rect 1933 2202 2000 2226
rect 2032 2226 2204 2228
rect 2002 2204 2030 2208
rect 2032 2204 2112 2226
rect 2133 2224 2148 2226
rect 2002 2202 2112 2204
rect 1933 2198 2112 2202
rect 1906 2188 1936 2198
rect 1938 2188 2091 2198
rect 2099 2188 2129 2198
rect 2133 2188 2163 2202
rect 2191 2188 2204 2226
rect 2276 2232 2311 2240
rect 2276 2206 2277 2232
rect 2284 2206 2311 2232
rect 2219 2188 2249 2202
rect 2276 2198 2311 2206
rect 2313 2232 2354 2240
rect 2313 2206 2328 2232
rect 2335 2206 2354 2232
rect 2418 2228 2480 2240
rect 2492 2228 2567 2240
rect 2625 2228 2700 2240
rect 2712 2228 2743 2240
rect 2749 2228 2784 2240
rect 2418 2226 2580 2228
rect 2313 2198 2354 2206
rect 2436 2202 2449 2226
rect 2464 2224 2479 2226
rect 2276 2188 2277 2198
rect 2292 2188 2305 2198
rect 2319 2188 2320 2198
rect 2335 2188 2348 2198
rect 2363 2188 2393 2202
rect 2436 2188 2479 2202
rect 2503 2199 2510 2206
rect 2513 2202 2580 2226
rect 2612 2226 2784 2228
rect 2582 2204 2610 2208
rect 2612 2204 2692 2226
rect 2713 2224 2728 2226
rect 2582 2202 2692 2204
rect 2513 2198 2692 2202
rect 2486 2188 2516 2198
rect 2518 2188 2671 2198
rect 2679 2188 2709 2198
rect 2713 2188 2743 2202
rect 2771 2188 2784 2226
rect 2856 2232 2891 2240
rect 2856 2206 2857 2232
rect 2864 2206 2891 2232
rect 2799 2188 2829 2202
rect 2856 2198 2891 2206
rect 2893 2232 2934 2240
rect 2893 2206 2908 2232
rect 2915 2206 2934 2232
rect 2998 2228 3060 2240
rect 3072 2228 3147 2240
rect 3205 2228 3280 2240
rect 3292 2228 3323 2240
rect 3329 2228 3364 2240
rect 2998 2226 3160 2228
rect 2893 2198 2934 2206
rect 3016 2202 3029 2226
rect 3044 2224 3059 2226
rect 2856 2188 2857 2198
rect 2872 2188 2885 2198
rect 2899 2188 2900 2198
rect 2915 2188 2928 2198
rect 2943 2188 2973 2202
rect 3016 2188 3059 2202
rect 3083 2199 3090 2206
rect 3093 2202 3160 2226
rect 3192 2226 3364 2228
rect 3162 2204 3190 2208
rect 3192 2204 3272 2226
rect 3293 2224 3308 2226
rect 3162 2202 3272 2204
rect 3093 2198 3272 2202
rect 3066 2188 3096 2198
rect 3098 2188 3251 2198
rect 3259 2188 3289 2198
rect 3293 2188 3323 2202
rect 3351 2188 3364 2226
rect 3436 2232 3471 2240
rect 3436 2206 3437 2232
rect 3444 2206 3471 2232
rect 3379 2188 3409 2202
rect 3436 2198 3471 2206
rect 3473 2232 3514 2240
rect 3473 2206 3488 2232
rect 3495 2206 3514 2232
rect 3578 2228 3640 2240
rect 3652 2228 3727 2240
rect 3785 2228 3860 2240
rect 3872 2228 3903 2240
rect 3909 2228 3944 2240
rect 3578 2226 3740 2228
rect 3473 2198 3514 2206
rect 3596 2202 3609 2226
rect 3624 2224 3639 2226
rect 3436 2188 3437 2198
rect 3452 2188 3465 2198
rect 3479 2188 3480 2198
rect 3495 2188 3508 2198
rect 3523 2188 3553 2202
rect 3596 2188 3639 2202
rect 3663 2199 3670 2206
rect 3673 2202 3740 2226
rect 3772 2226 3944 2228
rect 3742 2204 3770 2208
rect 3772 2204 3852 2226
rect 3873 2224 3888 2226
rect 3742 2202 3852 2204
rect 3673 2198 3852 2202
rect 3646 2188 3676 2198
rect 3678 2188 3831 2198
rect 3839 2188 3869 2198
rect 3873 2188 3903 2202
rect 3931 2188 3944 2226
rect 4016 2232 4051 2240
rect 4016 2206 4017 2232
rect 4024 2206 4051 2232
rect 3959 2188 3989 2202
rect 4016 2198 4051 2206
rect 4053 2232 4094 2240
rect 4053 2206 4068 2232
rect 4075 2206 4094 2232
rect 4158 2228 4220 2240
rect 4232 2228 4307 2240
rect 4365 2228 4440 2240
rect 4452 2228 4483 2240
rect 4489 2228 4524 2240
rect 4158 2226 4320 2228
rect 4053 2198 4094 2206
rect 4176 2202 4189 2226
rect 4204 2224 4219 2226
rect 4016 2188 4017 2198
rect 4032 2188 4045 2198
rect 4059 2188 4060 2198
rect 4075 2188 4088 2198
rect 4103 2188 4133 2202
rect 4176 2188 4219 2202
rect 4243 2199 4250 2206
rect 4253 2202 4320 2226
rect 4352 2226 4524 2228
rect 4322 2204 4350 2208
rect 4352 2204 4432 2226
rect 4453 2224 4468 2226
rect 4322 2202 4432 2204
rect 4253 2198 4432 2202
rect 4226 2188 4256 2198
rect 4258 2188 4411 2198
rect 4419 2188 4449 2198
rect 4453 2188 4483 2202
rect 4511 2188 4524 2226
rect 4596 2232 4631 2240
rect 4596 2206 4597 2232
rect 4604 2206 4631 2232
rect 4539 2188 4569 2202
rect 4596 2198 4631 2206
rect 4596 2188 4597 2198
rect 4612 2188 4625 2198
rect -1 2182 4625 2188
rect 0 2174 4625 2182
rect 15 2144 28 2174
rect 43 2156 73 2174
rect 116 2160 130 2174
rect 166 2160 386 2174
rect 117 2158 130 2160
rect 83 2146 98 2158
rect 80 2144 102 2146
rect 107 2144 137 2158
rect 198 2156 351 2160
rect 180 2144 372 2156
rect 415 2144 445 2158
rect 451 2144 464 2174
rect 479 2156 509 2174
rect 552 2144 565 2174
rect 595 2144 608 2174
rect 623 2156 653 2174
rect 696 2160 710 2174
rect 746 2160 966 2174
rect 697 2158 710 2160
rect 663 2146 678 2158
rect 660 2144 682 2146
rect 687 2144 717 2158
rect 778 2156 931 2160
rect 760 2144 952 2156
rect 995 2144 1025 2158
rect 1031 2144 1044 2174
rect 1059 2156 1089 2174
rect 1132 2144 1145 2174
rect 1175 2144 1188 2174
rect 1203 2156 1233 2174
rect 1276 2160 1290 2174
rect 1326 2160 1546 2174
rect 1277 2158 1290 2160
rect 1243 2146 1258 2158
rect 1240 2144 1262 2146
rect 1267 2144 1297 2158
rect 1358 2156 1511 2160
rect 1340 2144 1532 2156
rect 1575 2144 1605 2158
rect 1611 2144 1624 2174
rect 1639 2156 1669 2174
rect 1712 2144 1725 2174
rect 1755 2144 1768 2174
rect 1783 2156 1813 2174
rect 1856 2160 1870 2174
rect 1906 2160 2126 2174
rect 1857 2158 1870 2160
rect 1823 2146 1838 2158
rect 1820 2144 1842 2146
rect 1847 2144 1877 2158
rect 1938 2156 2091 2160
rect 1920 2144 2112 2156
rect 2155 2144 2185 2158
rect 2191 2144 2204 2174
rect 2219 2156 2249 2174
rect 2292 2144 2305 2174
rect 2335 2144 2348 2174
rect 2363 2156 2393 2174
rect 2436 2160 2450 2174
rect 2486 2160 2706 2174
rect 2437 2158 2450 2160
rect 2403 2146 2418 2158
rect 2400 2144 2422 2146
rect 2427 2144 2457 2158
rect 2518 2156 2671 2160
rect 2500 2144 2692 2156
rect 2735 2144 2765 2158
rect 2771 2144 2784 2174
rect 2799 2156 2829 2174
rect 2872 2144 2885 2174
rect 2915 2144 2928 2174
rect 2943 2156 2973 2174
rect 3016 2160 3030 2174
rect 3066 2160 3286 2174
rect 3017 2158 3030 2160
rect 2983 2146 2998 2158
rect 2980 2144 3002 2146
rect 3007 2144 3037 2158
rect 3098 2156 3251 2160
rect 3080 2144 3272 2156
rect 3315 2144 3345 2158
rect 3351 2144 3364 2174
rect 3379 2156 3409 2174
rect 3452 2144 3465 2174
rect 3495 2144 3508 2174
rect 3523 2156 3553 2174
rect 3596 2160 3610 2174
rect 3646 2160 3866 2174
rect 3597 2158 3610 2160
rect 3563 2146 3578 2158
rect 3560 2144 3582 2146
rect 3587 2144 3617 2158
rect 3678 2156 3831 2160
rect 3660 2144 3852 2156
rect 3895 2144 3925 2158
rect 3931 2144 3944 2174
rect 3959 2156 3989 2174
rect 4032 2144 4045 2174
rect 4075 2144 4088 2174
rect 4103 2156 4133 2174
rect 4176 2160 4190 2174
rect 4226 2160 4446 2174
rect 4177 2158 4190 2160
rect 4143 2146 4158 2158
rect 4140 2144 4162 2146
rect 4167 2144 4197 2158
rect 4258 2156 4411 2160
rect 4240 2144 4432 2156
rect 4475 2144 4505 2158
rect 4511 2144 4524 2174
rect 4539 2156 4569 2174
rect 4612 2144 4625 2174
rect 0 2130 4625 2144
rect 15 2026 28 2130
rect 73 2108 74 2118
rect 89 2108 102 2118
rect 73 2104 102 2108
rect 107 2104 137 2130
rect 155 2116 171 2118
rect 243 2116 296 2130
rect 244 2114 308 2116
rect 351 2114 366 2130
rect 415 2127 445 2130
rect 415 2124 451 2127
rect 381 2116 397 2118
rect 155 2104 170 2108
rect 73 2102 170 2104
rect 198 2102 366 2114
rect 382 2104 397 2108
rect 415 2105 454 2124
rect 473 2118 480 2119
rect 479 2111 480 2118
rect 463 2108 464 2111
rect 479 2108 492 2111
rect 415 2104 445 2105
rect 454 2104 460 2105
rect 463 2104 492 2108
rect 382 2103 492 2104
rect 382 2102 498 2103
rect 57 2094 108 2102
rect 57 2082 82 2094
rect 89 2082 108 2094
rect 139 2094 189 2102
rect 139 2086 155 2094
rect 162 2092 189 2094
rect 198 2092 419 2102
rect 162 2082 419 2092
rect 448 2094 498 2102
rect 448 2085 464 2094
rect 57 2074 108 2082
rect 155 2074 419 2082
rect 445 2082 464 2085
rect 471 2082 498 2094
rect 445 2074 498 2082
rect 73 2066 74 2074
rect 89 2066 102 2074
rect 73 2058 89 2066
rect 70 2051 89 2054
rect 70 2042 92 2051
rect 43 2032 92 2042
rect 43 2026 73 2032
rect 92 2027 97 2032
rect 15 2010 89 2026
rect 107 2018 137 2074
rect 172 2064 380 2074
rect 415 2070 460 2074
rect 463 2073 464 2074
rect 479 2073 492 2074
rect 198 2034 387 2064
rect 213 2031 387 2034
rect 206 2028 387 2031
rect 15 2008 28 2010
rect 43 2008 77 2010
rect 15 1992 89 2008
rect 116 2004 129 2018
rect 144 2004 160 2020
rect 206 2015 217 2028
rect -1 1970 0 1986
rect 15 1970 28 1992
rect 43 1970 73 1992
rect 116 1988 178 2004
rect 206 1997 217 2013
rect 222 2008 232 2028
rect 242 2008 256 2028
rect 259 2015 268 2028
rect 284 2015 293 2028
rect 222 1997 256 2008
rect 259 1997 268 2013
rect 284 1997 293 2013
rect 300 2008 310 2028
rect 320 2008 334 2028
rect 335 2015 346 2028
rect 300 1997 334 2008
rect 335 1997 346 2013
rect 392 2004 408 2020
rect 415 2018 445 2070
rect 479 2066 480 2073
rect 464 2058 480 2066
rect 451 2026 464 2045
rect 479 2026 509 2042
rect 451 2010 525 2026
rect 451 2008 464 2010
rect 479 2008 513 2010
rect 116 1986 129 1988
rect 144 1986 178 1988
rect 116 1970 178 1986
rect 222 1981 238 1984
rect 300 1981 330 1992
rect 378 1988 424 2004
rect 451 1992 525 2008
rect 378 1986 412 1988
rect 377 1970 424 1986
rect 451 1970 464 1992
rect 479 1970 509 1992
rect 536 1970 537 1986
rect 552 1970 565 2130
rect 595 2026 608 2130
rect 653 2108 654 2118
rect 669 2108 682 2118
rect 653 2104 682 2108
rect 687 2104 717 2130
rect 735 2116 751 2118
rect 823 2116 876 2130
rect 824 2114 888 2116
rect 931 2114 946 2130
rect 995 2127 1025 2130
rect 995 2124 1031 2127
rect 961 2116 977 2118
rect 735 2104 750 2108
rect 653 2102 750 2104
rect 778 2102 946 2114
rect 962 2104 977 2108
rect 995 2105 1034 2124
rect 1053 2118 1060 2119
rect 1059 2111 1060 2118
rect 1043 2108 1044 2111
rect 1059 2108 1072 2111
rect 995 2104 1025 2105
rect 1034 2104 1040 2105
rect 1043 2104 1072 2108
rect 962 2103 1072 2104
rect 962 2102 1078 2103
rect 637 2094 688 2102
rect 637 2082 662 2094
rect 669 2082 688 2094
rect 719 2094 769 2102
rect 719 2086 735 2094
rect 742 2092 769 2094
rect 778 2092 999 2102
rect 742 2082 999 2092
rect 1028 2094 1078 2102
rect 1028 2085 1044 2094
rect 637 2074 688 2082
rect 735 2074 999 2082
rect 1025 2082 1044 2085
rect 1051 2082 1078 2094
rect 1025 2074 1078 2082
rect 653 2066 654 2074
rect 669 2066 682 2074
rect 653 2058 669 2066
rect 650 2051 669 2054
rect 650 2042 672 2051
rect 623 2032 672 2042
rect 623 2026 653 2032
rect 672 2027 677 2032
rect 595 2010 669 2026
rect 687 2018 717 2074
rect 752 2064 960 2074
rect 995 2070 1040 2074
rect 1043 2073 1044 2074
rect 1059 2073 1072 2074
rect 778 2034 967 2064
rect 793 2031 967 2034
rect 786 2028 967 2031
rect 595 2008 608 2010
rect 623 2008 657 2010
rect 595 1992 669 2008
rect 696 2004 709 2018
rect 724 2004 740 2020
rect 786 2015 797 2028
rect 579 1970 580 1986
rect 595 1970 608 1992
rect 623 1970 653 1992
rect 696 1988 758 2004
rect 786 1997 797 2013
rect 802 2008 812 2028
rect 822 2008 836 2028
rect 839 2015 848 2028
rect 864 2015 873 2028
rect 802 1997 836 2008
rect 839 1997 848 2013
rect 864 1997 873 2013
rect 880 2008 890 2028
rect 900 2008 914 2028
rect 915 2015 926 2028
rect 880 1997 914 2008
rect 915 1997 926 2013
rect 972 2004 988 2020
rect 995 2018 1025 2070
rect 1059 2066 1060 2073
rect 1044 2058 1060 2066
rect 1031 2026 1044 2045
rect 1059 2026 1089 2042
rect 1031 2010 1105 2026
rect 1031 2008 1044 2010
rect 1059 2008 1093 2010
rect 696 1986 709 1988
rect 724 1986 758 1988
rect 696 1970 758 1986
rect 802 1981 818 1984
rect 880 1981 910 1992
rect 958 1988 1004 2004
rect 1031 1992 1105 2008
rect 958 1986 992 1988
rect 957 1970 1004 1986
rect 1031 1970 1044 1992
rect 1059 1970 1089 1992
rect 1116 1970 1117 1986
rect 1132 1970 1145 2130
rect 1175 2026 1188 2130
rect 1233 2108 1234 2118
rect 1249 2108 1262 2118
rect 1233 2104 1262 2108
rect 1267 2104 1297 2130
rect 1315 2116 1331 2118
rect 1403 2116 1456 2130
rect 1404 2114 1468 2116
rect 1511 2114 1526 2130
rect 1575 2127 1605 2130
rect 1575 2124 1611 2127
rect 1541 2116 1557 2118
rect 1315 2104 1330 2108
rect 1233 2102 1330 2104
rect 1358 2102 1526 2114
rect 1542 2104 1557 2108
rect 1575 2105 1614 2124
rect 1633 2118 1640 2119
rect 1639 2111 1640 2118
rect 1623 2108 1624 2111
rect 1639 2108 1652 2111
rect 1575 2104 1605 2105
rect 1614 2104 1620 2105
rect 1623 2104 1652 2108
rect 1542 2103 1652 2104
rect 1542 2102 1658 2103
rect 1217 2094 1268 2102
rect 1217 2082 1242 2094
rect 1249 2082 1268 2094
rect 1299 2094 1349 2102
rect 1299 2086 1315 2094
rect 1322 2092 1349 2094
rect 1358 2092 1579 2102
rect 1322 2082 1579 2092
rect 1608 2094 1658 2102
rect 1608 2085 1624 2094
rect 1217 2074 1268 2082
rect 1315 2074 1579 2082
rect 1605 2082 1624 2085
rect 1631 2082 1658 2094
rect 1605 2074 1658 2082
rect 1233 2066 1234 2074
rect 1249 2066 1262 2074
rect 1233 2058 1249 2066
rect 1230 2051 1249 2054
rect 1230 2042 1252 2051
rect 1203 2032 1252 2042
rect 1203 2026 1233 2032
rect 1252 2027 1257 2032
rect 1175 2010 1249 2026
rect 1267 2018 1297 2074
rect 1332 2064 1540 2074
rect 1575 2070 1620 2074
rect 1623 2073 1624 2074
rect 1639 2073 1652 2074
rect 1358 2034 1547 2064
rect 1373 2031 1547 2034
rect 1366 2028 1547 2031
rect 1175 2008 1188 2010
rect 1203 2008 1237 2010
rect 1175 1992 1249 2008
rect 1276 2004 1289 2018
rect 1304 2004 1320 2020
rect 1366 2015 1377 2028
rect 1159 1970 1160 1986
rect 1175 1970 1188 1992
rect 1203 1970 1233 1992
rect 1276 1988 1338 2004
rect 1366 1997 1377 2013
rect 1382 2008 1392 2028
rect 1402 2008 1416 2028
rect 1419 2015 1428 2028
rect 1444 2015 1453 2028
rect 1382 1997 1416 2008
rect 1419 1997 1428 2013
rect 1444 1997 1453 2013
rect 1460 2008 1470 2028
rect 1480 2008 1494 2028
rect 1495 2015 1506 2028
rect 1460 1997 1494 2008
rect 1495 1997 1506 2013
rect 1552 2004 1568 2020
rect 1575 2018 1605 2070
rect 1639 2066 1640 2073
rect 1624 2058 1640 2066
rect 1611 2026 1624 2045
rect 1639 2026 1669 2042
rect 1611 2010 1685 2026
rect 1611 2008 1624 2010
rect 1639 2008 1673 2010
rect 1276 1986 1289 1988
rect 1304 1986 1338 1988
rect 1276 1970 1338 1986
rect 1382 1981 1398 1984
rect 1460 1981 1490 1992
rect 1538 1988 1584 2004
rect 1611 1992 1685 2008
rect 1538 1986 1572 1988
rect 1537 1970 1584 1986
rect 1611 1970 1624 1992
rect 1639 1970 1669 1992
rect 1696 1970 1697 1986
rect 1712 1970 1725 2130
rect 1755 2026 1768 2130
rect 1813 2108 1814 2118
rect 1829 2108 1842 2118
rect 1813 2104 1842 2108
rect 1847 2104 1877 2130
rect 1895 2116 1911 2118
rect 1983 2116 2036 2130
rect 1984 2114 2048 2116
rect 2091 2114 2106 2130
rect 2155 2127 2185 2130
rect 2155 2124 2191 2127
rect 2121 2116 2137 2118
rect 1895 2104 1910 2108
rect 1813 2102 1910 2104
rect 1938 2102 2106 2114
rect 2122 2104 2137 2108
rect 2155 2105 2194 2124
rect 2213 2118 2220 2119
rect 2219 2111 2220 2118
rect 2203 2108 2204 2111
rect 2219 2108 2232 2111
rect 2155 2104 2185 2105
rect 2194 2104 2200 2105
rect 2203 2104 2232 2108
rect 2122 2103 2232 2104
rect 2122 2102 2238 2103
rect 1797 2094 1848 2102
rect 1797 2082 1822 2094
rect 1829 2082 1848 2094
rect 1879 2094 1929 2102
rect 1879 2086 1895 2094
rect 1902 2092 1929 2094
rect 1938 2092 2159 2102
rect 1902 2082 2159 2092
rect 2188 2094 2238 2102
rect 2188 2085 2204 2094
rect 1797 2074 1848 2082
rect 1895 2074 2159 2082
rect 2185 2082 2204 2085
rect 2211 2082 2238 2094
rect 2185 2074 2238 2082
rect 1813 2066 1814 2074
rect 1829 2066 1842 2074
rect 1813 2058 1829 2066
rect 1810 2051 1829 2054
rect 1810 2042 1832 2051
rect 1783 2032 1832 2042
rect 1783 2026 1813 2032
rect 1832 2027 1837 2032
rect 1755 2010 1829 2026
rect 1847 2018 1877 2074
rect 1912 2064 2120 2074
rect 2155 2070 2200 2074
rect 2203 2073 2204 2074
rect 2219 2073 2232 2074
rect 1938 2034 2127 2064
rect 1953 2031 2127 2034
rect 1946 2028 2127 2031
rect 1755 2008 1768 2010
rect 1783 2008 1817 2010
rect 1755 1992 1829 2008
rect 1856 2004 1869 2018
rect 1884 2004 1900 2020
rect 1946 2015 1957 2028
rect 1739 1970 1740 1986
rect 1755 1970 1768 1992
rect 1783 1970 1813 1992
rect 1856 1988 1918 2004
rect 1946 1997 1957 2013
rect 1962 2008 1972 2028
rect 1982 2008 1996 2028
rect 1999 2015 2008 2028
rect 2024 2015 2033 2028
rect 1962 1997 1996 2008
rect 1999 1997 2008 2013
rect 2024 1997 2033 2013
rect 2040 2008 2050 2028
rect 2060 2008 2074 2028
rect 2075 2015 2086 2028
rect 2040 1997 2074 2008
rect 2075 1997 2086 2013
rect 2132 2004 2148 2020
rect 2155 2018 2185 2070
rect 2219 2066 2220 2073
rect 2204 2058 2220 2066
rect 2191 2026 2204 2045
rect 2219 2026 2249 2042
rect 2191 2010 2265 2026
rect 2191 2008 2204 2010
rect 2219 2008 2253 2010
rect 1856 1986 1869 1988
rect 1884 1986 1918 1988
rect 1856 1970 1918 1986
rect 1962 1981 1978 1984
rect 2040 1981 2070 1992
rect 2118 1988 2164 2004
rect 2191 1992 2265 2008
rect 2118 1986 2152 1988
rect 2117 1970 2164 1986
rect 2191 1970 2204 1992
rect 2219 1970 2249 1992
rect 2276 1970 2277 1986
rect 2292 1970 2305 2130
rect 2335 2026 2348 2130
rect 2393 2108 2394 2118
rect 2409 2108 2422 2118
rect 2393 2104 2422 2108
rect 2427 2104 2457 2130
rect 2475 2116 2491 2118
rect 2563 2116 2616 2130
rect 2564 2114 2628 2116
rect 2671 2114 2686 2130
rect 2735 2127 2765 2130
rect 2735 2124 2771 2127
rect 2701 2116 2717 2118
rect 2475 2104 2490 2108
rect 2393 2102 2490 2104
rect 2518 2102 2686 2114
rect 2702 2104 2717 2108
rect 2735 2105 2774 2124
rect 2793 2118 2800 2119
rect 2799 2111 2800 2118
rect 2783 2108 2784 2111
rect 2799 2108 2812 2111
rect 2735 2104 2765 2105
rect 2774 2104 2780 2105
rect 2783 2104 2812 2108
rect 2702 2103 2812 2104
rect 2702 2102 2818 2103
rect 2377 2094 2428 2102
rect 2377 2082 2402 2094
rect 2409 2082 2428 2094
rect 2459 2094 2509 2102
rect 2459 2086 2475 2094
rect 2482 2092 2509 2094
rect 2518 2092 2739 2102
rect 2482 2082 2739 2092
rect 2768 2094 2818 2102
rect 2768 2085 2784 2094
rect 2377 2074 2428 2082
rect 2475 2074 2739 2082
rect 2765 2082 2784 2085
rect 2791 2082 2818 2094
rect 2765 2074 2818 2082
rect 2393 2066 2394 2074
rect 2409 2066 2422 2074
rect 2393 2058 2409 2066
rect 2390 2051 2409 2054
rect 2390 2042 2412 2051
rect 2363 2032 2412 2042
rect 2363 2026 2393 2032
rect 2412 2027 2417 2032
rect 2335 2010 2409 2026
rect 2427 2018 2457 2074
rect 2492 2064 2700 2074
rect 2735 2070 2780 2074
rect 2783 2073 2784 2074
rect 2799 2073 2812 2074
rect 2518 2034 2707 2064
rect 2533 2031 2707 2034
rect 2526 2028 2707 2031
rect 2335 2008 2348 2010
rect 2363 2008 2397 2010
rect 2335 1992 2409 2008
rect 2436 2004 2449 2018
rect 2464 2004 2480 2020
rect 2526 2015 2537 2028
rect 2319 1970 2320 1986
rect 2335 1970 2348 1992
rect 2363 1970 2393 1992
rect 2436 1988 2498 2004
rect 2526 1997 2537 2013
rect 2542 2008 2552 2028
rect 2562 2008 2576 2028
rect 2579 2015 2588 2028
rect 2604 2015 2613 2028
rect 2542 1997 2576 2008
rect 2579 1997 2588 2013
rect 2604 1997 2613 2013
rect 2620 2008 2630 2028
rect 2640 2008 2654 2028
rect 2655 2015 2666 2028
rect 2620 1997 2654 2008
rect 2655 1997 2666 2013
rect 2712 2004 2728 2020
rect 2735 2018 2765 2070
rect 2799 2066 2800 2073
rect 2784 2058 2800 2066
rect 2771 2026 2784 2045
rect 2799 2026 2829 2042
rect 2771 2010 2845 2026
rect 2771 2008 2784 2010
rect 2799 2008 2833 2010
rect 2436 1986 2449 1988
rect 2464 1986 2498 1988
rect 2436 1970 2498 1986
rect 2542 1981 2558 1984
rect 2620 1981 2650 1992
rect 2698 1988 2744 2004
rect 2771 1992 2845 2008
rect 2698 1986 2732 1988
rect 2697 1970 2744 1986
rect 2771 1970 2784 1992
rect 2799 1970 2829 1992
rect 2856 1970 2857 1986
rect 2872 1970 2885 2130
rect 2915 2026 2928 2130
rect 2973 2108 2974 2118
rect 2989 2108 3002 2118
rect 2973 2104 3002 2108
rect 3007 2104 3037 2130
rect 3055 2116 3071 2118
rect 3143 2116 3196 2130
rect 3144 2114 3208 2116
rect 3251 2114 3266 2130
rect 3315 2127 3345 2130
rect 3315 2124 3351 2127
rect 3281 2116 3297 2118
rect 3055 2104 3070 2108
rect 2973 2102 3070 2104
rect 3098 2102 3266 2114
rect 3282 2104 3297 2108
rect 3315 2105 3354 2124
rect 3373 2118 3380 2119
rect 3379 2111 3380 2118
rect 3363 2108 3364 2111
rect 3379 2108 3392 2111
rect 3315 2104 3345 2105
rect 3354 2104 3360 2105
rect 3363 2104 3392 2108
rect 3282 2103 3392 2104
rect 3282 2102 3398 2103
rect 2957 2094 3008 2102
rect 2957 2082 2982 2094
rect 2989 2082 3008 2094
rect 3039 2094 3089 2102
rect 3039 2086 3055 2094
rect 3062 2092 3089 2094
rect 3098 2092 3319 2102
rect 3062 2082 3319 2092
rect 3348 2094 3398 2102
rect 3348 2085 3364 2094
rect 2957 2074 3008 2082
rect 3055 2074 3319 2082
rect 3345 2082 3364 2085
rect 3371 2082 3398 2094
rect 3345 2074 3398 2082
rect 2973 2066 2974 2074
rect 2989 2066 3002 2074
rect 2973 2058 2989 2066
rect 2970 2051 2989 2054
rect 2970 2042 2992 2051
rect 2943 2032 2992 2042
rect 2943 2026 2973 2032
rect 2992 2027 2997 2032
rect 2915 2010 2989 2026
rect 3007 2018 3037 2074
rect 3072 2064 3280 2074
rect 3315 2070 3360 2074
rect 3363 2073 3364 2074
rect 3379 2073 3392 2074
rect 3098 2034 3287 2064
rect 3113 2031 3287 2034
rect 3106 2028 3287 2031
rect 2915 2008 2928 2010
rect 2943 2008 2977 2010
rect 2915 1992 2989 2008
rect 3016 2004 3029 2018
rect 3044 2004 3060 2020
rect 3106 2015 3117 2028
rect 2899 1970 2900 1986
rect 2915 1970 2928 1992
rect 2943 1970 2973 1992
rect 3016 1988 3078 2004
rect 3106 1997 3117 2013
rect 3122 2008 3132 2028
rect 3142 2008 3156 2028
rect 3159 2015 3168 2028
rect 3184 2015 3193 2028
rect 3122 1997 3156 2008
rect 3159 1997 3168 2013
rect 3184 1997 3193 2013
rect 3200 2008 3210 2028
rect 3220 2008 3234 2028
rect 3235 2015 3246 2028
rect 3200 1997 3234 2008
rect 3235 1997 3246 2013
rect 3292 2004 3308 2020
rect 3315 2018 3345 2070
rect 3379 2066 3380 2073
rect 3364 2058 3380 2066
rect 3351 2026 3364 2045
rect 3379 2026 3409 2042
rect 3351 2010 3425 2026
rect 3351 2008 3364 2010
rect 3379 2008 3413 2010
rect 3016 1986 3029 1988
rect 3044 1986 3078 1988
rect 3016 1970 3078 1986
rect 3122 1981 3138 1984
rect 3200 1981 3230 1992
rect 3278 1988 3324 2004
rect 3351 1992 3425 2008
rect 3278 1986 3312 1988
rect 3277 1970 3324 1986
rect 3351 1970 3364 1992
rect 3379 1970 3409 1992
rect 3436 1970 3437 1986
rect 3452 1970 3465 2130
rect 3495 2026 3508 2130
rect 3553 2108 3554 2118
rect 3569 2108 3582 2118
rect 3553 2104 3582 2108
rect 3587 2104 3617 2130
rect 3635 2116 3651 2118
rect 3723 2116 3776 2130
rect 3724 2114 3788 2116
rect 3831 2114 3846 2130
rect 3895 2127 3925 2130
rect 3895 2124 3931 2127
rect 3861 2116 3877 2118
rect 3635 2104 3650 2108
rect 3553 2102 3650 2104
rect 3678 2102 3846 2114
rect 3862 2104 3877 2108
rect 3895 2105 3934 2124
rect 3953 2118 3960 2119
rect 3959 2111 3960 2118
rect 3943 2108 3944 2111
rect 3959 2108 3972 2111
rect 3895 2104 3925 2105
rect 3934 2104 3940 2105
rect 3943 2104 3972 2108
rect 3862 2103 3972 2104
rect 3862 2102 3978 2103
rect 3537 2094 3588 2102
rect 3537 2082 3562 2094
rect 3569 2082 3588 2094
rect 3619 2094 3669 2102
rect 3619 2086 3635 2094
rect 3642 2092 3669 2094
rect 3678 2092 3899 2102
rect 3642 2082 3899 2092
rect 3928 2094 3978 2102
rect 3928 2085 3944 2094
rect 3537 2074 3588 2082
rect 3635 2074 3899 2082
rect 3925 2082 3944 2085
rect 3951 2082 3978 2094
rect 3925 2074 3978 2082
rect 3553 2066 3554 2074
rect 3569 2066 3582 2074
rect 3553 2058 3569 2066
rect 3550 2051 3569 2054
rect 3550 2042 3572 2051
rect 3523 2032 3572 2042
rect 3523 2026 3553 2032
rect 3572 2027 3577 2032
rect 3495 2010 3569 2026
rect 3587 2018 3617 2074
rect 3652 2064 3860 2074
rect 3895 2070 3940 2074
rect 3943 2073 3944 2074
rect 3959 2073 3972 2074
rect 3678 2034 3867 2064
rect 3693 2031 3867 2034
rect 3686 2028 3867 2031
rect 3495 2008 3508 2010
rect 3523 2008 3557 2010
rect 3495 1992 3569 2008
rect 3596 2004 3609 2018
rect 3624 2004 3640 2020
rect 3686 2015 3697 2028
rect 3479 1970 3480 1986
rect 3495 1970 3508 1992
rect 3523 1970 3553 1992
rect 3596 1988 3658 2004
rect 3686 1997 3697 2013
rect 3702 2008 3712 2028
rect 3722 2008 3736 2028
rect 3739 2015 3748 2028
rect 3764 2015 3773 2028
rect 3702 1997 3736 2008
rect 3739 1997 3748 2013
rect 3764 1997 3773 2013
rect 3780 2008 3790 2028
rect 3800 2008 3814 2028
rect 3815 2015 3826 2028
rect 3780 1997 3814 2008
rect 3815 1997 3826 2013
rect 3872 2004 3888 2020
rect 3895 2018 3925 2070
rect 3959 2066 3960 2073
rect 3944 2058 3960 2066
rect 3931 2026 3944 2045
rect 3959 2026 3989 2042
rect 3931 2010 4005 2026
rect 3931 2008 3944 2010
rect 3959 2008 3993 2010
rect 3596 1986 3609 1988
rect 3624 1986 3658 1988
rect 3596 1970 3658 1986
rect 3702 1981 3718 1984
rect 3780 1981 3810 1992
rect 3858 1988 3904 2004
rect 3931 1992 4005 2008
rect 3858 1986 3892 1988
rect 3857 1970 3904 1986
rect 3931 1970 3944 1992
rect 3959 1970 3989 1992
rect 4016 1970 4017 1986
rect 4032 1970 4045 2130
rect 4075 2026 4088 2130
rect 4133 2108 4134 2118
rect 4149 2108 4162 2118
rect 4133 2104 4162 2108
rect 4167 2104 4197 2130
rect 4215 2116 4231 2118
rect 4303 2116 4356 2130
rect 4304 2114 4368 2116
rect 4411 2114 4426 2130
rect 4475 2127 4505 2130
rect 4475 2124 4511 2127
rect 4441 2116 4457 2118
rect 4215 2104 4230 2108
rect 4133 2102 4230 2104
rect 4258 2102 4426 2114
rect 4442 2104 4457 2108
rect 4475 2105 4514 2124
rect 4533 2118 4540 2119
rect 4539 2111 4540 2118
rect 4523 2108 4524 2111
rect 4539 2108 4552 2111
rect 4475 2104 4505 2105
rect 4514 2104 4520 2105
rect 4523 2104 4552 2108
rect 4442 2103 4552 2104
rect 4442 2102 4558 2103
rect 4117 2094 4168 2102
rect 4117 2082 4142 2094
rect 4149 2082 4168 2094
rect 4199 2094 4249 2102
rect 4199 2086 4215 2094
rect 4222 2092 4249 2094
rect 4258 2092 4479 2102
rect 4222 2082 4479 2092
rect 4508 2094 4558 2102
rect 4508 2085 4524 2094
rect 4117 2074 4168 2082
rect 4215 2074 4479 2082
rect 4505 2082 4524 2085
rect 4531 2082 4558 2094
rect 4505 2074 4558 2082
rect 4133 2066 4134 2074
rect 4149 2066 4162 2074
rect 4133 2058 4149 2066
rect 4130 2051 4149 2054
rect 4130 2042 4152 2051
rect 4103 2032 4152 2042
rect 4103 2026 4133 2032
rect 4152 2027 4157 2032
rect 4075 2010 4149 2026
rect 4167 2018 4197 2074
rect 4232 2064 4440 2074
rect 4475 2070 4520 2074
rect 4523 2073 4524 2074
rect 4539 2073 4552 2074
rect 4258 2034 4447 2064
rect 4273 2031 4447 2034
rect 4266 2028 4447 2031
rect 4075 2008 4088 2010
rect 4103 2008 4137 2010
rect 4075 1992 4149 2008
rect 4176 2004 4189 2018
rect 4204 2004 4220 2020
rect 4266 2015 4277 2028
rect 4059 1970 4060 1986
rect 4075 1970 4088 1992
rect 4103 1970 4133 1992
rect 4176 1988 4238 2004
rect 4266 1997 4277 2013
rect 4282 2008 4292 2028
rect 4302 2008 4316 2028
rect 4319 2015 4328 2028
rect 4344 2015 4353 2028
rect 4282 1997 4316 2008
rect 4319 1997 4328 2013
rect 4344 1997 4353 2013
rect 4360 2008 4370 2028
rect 4380 2008 4394 2028
rect 4395 2015 4406 2028
rect 4360 1997 4394 2008
rect 4395 1997 4406 2013
rect 4452 2004 4468 2020
rect 4475 2018 4505 2070
rect 4539 2066 4540 2073
rect 4524 2058 4540 2066
rect 4511 2026 4524 2045
rect 4539 2026 4569 2042
rect 4511 2010 4585 2026
rect 4511 2008 4524 2010
rect 4539 2008 4573 2010
rect 4176 1986 4189 1988
rect 4204 1986 4238 1988
rect 4176 1970 4238 1986
rect 4282 1981 4298 1984
rect 4360 1981 4390 1992
rect 4438 1988 4484 2004
rect 4511 1992 4585 2008
rect 4438 1986 4472 1988
rect 4437 1970 4484 1986
rect 4511 1970 4524 1992
rect 4539 1970 4569 1992
rect 4596 1970 4597 1986
rect 4612 1970 4625 2130
rect -7 1962 34 1970
rect -7 1936 8 1962
rect 15 1936 34 1962
rect 98 1958 160 1970
rect 172 1958 247 1970
rect 305 1958 380 1970
rect 392 1958 423 1970
rect 429 1958 464 1970
rect 98 1956 260 1958
rect -7 1928 34 1936
rect 116 1932 129 1956
rect 144 1954 159 1956
rect -1 1918 0 1928
rect 15 1918 28 1928
rect 43 1918 73 1932
rect 116 1918 159 1932
rect 183 1929 190 1936
rect 193 1932 260 1956
rect 292 1956 464 1958
rect 262 1934 290 1938
rect 292 1934 372 1956
rect 393 1954 408 1956
rect 262 1932 372 1934
rect 193 1928 372 1932
rect 166 1918 196 1928
rect 198 1918 351 1928
rect 359 1918 389 1928
rect 393 1918 423 1932
rect 451 1918 464 1956
rect 536 1962 571 1970
rect 536 1936 537 1962
rect 544 1936 571 1962
rect 479 1918 509 1932
rect 536 1928 571 1936
rect 573 1962 614 1970
rect 573 1936 588 1962
rect 595 1936 614 1962
rect 678 1958 740 1970
rect 752 1958 827 1970
rect 885 1958 960 1970
rect 972 1958 1003 1970
rect 1009 1958 1044 1970
rect 678 1956 840 1958
rect 573 1928 614 1936
rect 696 1932 709 1956
rect 724 1954 739 1956
rect 536 1918 537 1928
rect 552 1918 565 1928
rect 579 1918 580 1928
rect 595 1918 608 1928
rect 623 1918 653 1932
rect 696 1918 739 1932
rect 763 1929 770 1936
rect 773 1932 840 1956
rect 872 1956 1044 1958
rect 842 1934 870 1938
rect 872 1934 952 1956
rect 973 1954 988 1956
rect 842 1932 952 1934
rect 773 1928 952 1932
rect 746 1918 776 1928
rect 778 1918 931 1928
rect 939 1918 969 1928
rect 973 1918 1003 1932
rect 1031 1918 1044 1956
rect 1116 1962 1151 1970
rect 1116 1936 1117 1962
rect 1124 1936 1151 1962
rect 1059 1918 1089 1932
rect 1116 1928 1151 1936
rect 1153 1962 1194 1970
rect 1153 1936 1168 1962
rect 1175 1936 1194 1962
rect 1258 1958 1320 1970
rect 1332 1958 1407 1970
rect 1465 1958 1540 1970
rect 1552 1958 1583 1970
rect 1589 1958 1624 1970
rect 1258 1956 1420 1958
rect 1153 1928 1194 1936
rect 1276 1932 1289 1956
rect 1304 1954 1319 1956
rect 1116 1918 1117 1928
rect 1132 1918 1145 1928
rect 1159 1918 1160 1928
rect 1175 1918 1188 1928
rect 1203 1918 1233 1932
rect 1276 1918 1319 1932
rect 1343 1929 1350 1936
rect 1353 1932 1420 1956
rect 1452 1956 1624 1958
rect 1422 1934 1450 1938
rect 1452 1934 1532 1956
rect 1553 1954 1568 1956
rect 1422 1932 1532 1934
rect 1353 1928 1532 1932
rect 1326 1918 1356 1928
rect 1358 1918 1511 1928
rect 1519 1918 1549 1928
rect 1553 1918 1583 1932
rect 1611 1918 1624 1956
rect 1696 1962 1731 1970
rect 1696 1936 1697 1962
rect 1704 1936 1731 1962
rect 1639 1918 1669 1932
rect 1696 1928 1731 1936
rect 1733 1962 1774 1970
rect 1733 1936 1748 1962
rect 1755 1936 1774 1962
rect 1838 1958 1900 1970
rect 1912 1958 1987 1970
rect 2045 1958 2120 1970
rect 2132 1958 2163 1970
rect 2169 1958 2204 1970
rect 1838 1956 2000 1958
rect 1733 1928 1774 1936
rect 1856 1932 1869 1956
rect 1884 1954 1899 1956
rect 1696 1918 1697 1928
rect 1712 1918 1725 1928
rect 1739 1918 1740 1928
rect 1755 1918 1768 1928
rect 1783 1918 1813 1932
rect 1856 1918 1899 1932
rect 1923 1929 1930 1936
rect 1933 1932 2000 1956
rect 2032 1956 2204 1958
rect 2002 1934 2030 1938
rect 2032 1934 2112 1956
rect 2133 1954 2148 1956
rect 2002 1932 2112 1934
rect 1933 1928 2112 1932
rect 1906 1918 1936 1928
rect 1938 1918 2091 1928
rect 2099 1918 2129 1928
rect 2133 1918 2163 1932
rect 2191 1918 2204 1956
rect 2276 1962 2311 1970
rect 2276 1936 2277 1962
rect 2284 1936 2311 1962
rect 2219 1918 2249 1932
rect 2276 1928 2311 1936
rect 2313 1962 2354 1970
rect 2313 1936 2328 1962
rect 2335 1936 2354 1962
rect 2418 1958 2480 1970
rect 2492 1958 2567 1970
rect 2625 1958 2700 1970
rect 2712 1958 2743 1970
rect 2749 1958 2784 1970
rect 2418 1956 2580 1958
rect 2313 1928 2354 1936
rect 2436 1932 2449 1956
rect 2464 1954 2479 1956
rect 2276 1918 2277 1928
rect 2292 1918 2305 1928
rect 2319 1918 2320 1928
rect 2335 1918 2348 1928
rect 2363 1918 2393 1932
rect 2436 1918 2479 1932
rect 2503 1929 2510 1936
rect 2513 1932 2580 1956
rect 2612 1956 2784 1958
rect 2582 1934 2610 1938
rect 2612 1934 2692 1956
rect 2713 1954 2728 1956
rect 2582 1932 2692 1934
rect 2513 1928 2692 1932
rect 2486 1918 2516 1928
rect 2518 1918 2671 1928
rect 2679 1918 2709 1928
rect 2713 1918 2743 1932
rect 2771 1918 2784 1956
rect 2856 1962 2891 1970
rect 2856 1936 2857 1962
rect 2864 1936 2891 1962
rect 2799 1918 2829 1932
rect 2856 1928 2891 1936
rect 2893 1962 2934 1970
rect 2893 1936 2908 1962
rect 2915 1936 2934 1962
rect 2998 1958 3060 1970
rect 3072 1958 3147 1970
rect 3205 1958 3280 1970
rect 3292 1958 3323 1970
rect 3329 1958 3364 1970
rect 2998 1956 3160 1958
rect 2893 1928 2934 1936
rect 3016 1932 3029 1956
rect 3044 1954 3059 1956
rect 2856 1918 2857 1928
rect 2872 1918 2885 1928
rect 2899 1918 2900 1928
rect 2915 1918 2928 1928
rect 2943 1918 2973 1932
rect 3016 1918 3059 1932
rect 3083 1929 3090 1936
rect 3093 1932 3160 1956
rect 3192 1956 3364 1958
rect 3162 1934 3190 1938
rect 3192 1934 3272 1956
rect 3293 1954 3308 1956
rect 3162 1932 3272 1934
rect 3093 1928 3272 1932
rect 3066 1918 3096 1928
rect 3098 1918 3251 1928
rect 3259 1918 3289 1928
rect 3293 1918 3323 1932
rect 3351 1918 3364 1956
rect 3436 1962 3471 1970
rect 3436 1936 3437 1962
rect 3444 1936 3471 1962
rect 3379 1918 3409 1932
rect 3436 1928 3471 1936
rect 3473 1962 3514 1970
rect 3473 1936 3488 1962
rect 3495 1936 3514 1962
rect 3578 1958 3640 1970
rect 3652 1958 3727 1970
rect 3785 1958 3860 1970
rect 3872 1958 3903 1970
rect 3909 1958 3944 1970
rect 3578 1956 3740 1958
rect 3473 1928 3514 1936
rect 3596 1932 3609 1956
rect 3624 1954 3639 1956
rect 3436 1918 3437 1928
rect 3452 1918 3465 1928
rect 3479 1918 3480 1928
rect 3495 1918 3508 1928
rect 3523 1918 3553 1932
rect 3596 1918 3639 1932
rect 3663 1929 3670 1936
rect 3673 1932 3740 1956
rect 3772 1956 3944 1958
rect 3742 1934 3770 1938
rect 3772 1934 3852 1956
rect 3873 1954 3888 1956
rect 3742 1932 3852 1934
rect 3673 1928 3852 1932
rect 3646 1918 3676 1928
rect 3678 1918 3831 1928
rect 3839 1918 3869 1928
rect 3873 1918 3903 1932
rect 3931 1918 3944 1956
rect 4016 1962 4051 1970
rect 4016 1936 4017 1962
rect 4024 1936 4051 1962
rect 3959 1918 3989 1932
rect 4016 1928 4051 1936
rect 4053 1962 4094 1970
rect 4053 1936 4068 1962
rect 4075 1936 4094 1962
rect 4158 1958 4220 1970
rect 4232 1958 4307 1970
rect 4365 1958 4440 1970
rect 4452 1958 4483 1970
rect 4489 1958 4524 1970
rect 4158 1956 4320 1958
rect 4053 1928 4094 1936
rect 4176 1932 4189 1956
rect 4204 1954 4219 1956
rect 4016 1918 4017 1928
rect 4032 1918 4045 1928
rect 4059 1918 4060 1928
rect 4075 1918 4088 1928
rect 4103 1918 4133 1932
rect 4176 1918 4219 1932
rect 4243 1929 4250 1936
rect 4253 1932 4320 1956
rect 4352 1956 4524 1958
rect 4322 1934 4350 1938
rect 4352 1934 4432 1956
rect 4453 1954 4468 1956
rect 4322 1932 4432 1934
rect 4253 1928 4432 1932
rect 4226 1918 4256 1928
rect 4258 1918 4411 1928
rect 4419 1918 4449 1928
rect 4453 1918 4483 1932
rect 4511 1918 4524 1956
rect 4596 1962 4631 1970
rect 4596 1936 4597 1962
rect 4604 1936 4631 1962
rect 4539 1918 4569 1932
rect 4596 1928 4631 1936
rect 4596 1918 4597 1928
rect 4612 1918 4625 1928
rect -1 1912 4625 1918
rect 0 1904 4625 1912
rect 15 1874 28 1904
rect 43 1886 73 1904
rect 116 1890 130 1904
rect 166 1890 386 1904
rect 117 1888 130 1890
rect 83 1876 98 1888
rect 80 1874 102 1876
rect 107 1874 137 1888
rect 198 1886 351 1890
rect 180 1874 372 1886
rect 415 1874 445 1888
rect 451 1874 464 1904
rect 479 1886 509 1904
rect 552 1874 565 1904
rect 595 1874 608 1904
rect 623 1886 653 1904
rect 696 1890 710 1904
rect 746 1890 966 1904
rect 697 1888 710 1890
rect 663 1876 678 1888
rect 660 1874 682 1876
rect 687 1874 717 1888
rect 778 1886 931 1890
rect 760 1874 952 1886
rect 995 1874 1025 1888
rect 1031 1874 1044 1904
rect 1059 1886 1089 1904
rect 1132 1874 1145 1904
rect 1175 1874 1188 1904
rect 1203 1886 1233 1904
rect 1276 1890 1290 1904
rect 1326 1890 1546 1904
rect 1277 1888 1290 1890
rect 1243 1876 1258 1888
rect 1240 1874 1262 1876
rect 1267 1874 1297 1888
rect 1358 1886 1511 1890
rect 1340 1874 1532 1886
rect 1575 1874 1605 1888
rect 1611 1874 1624 1904
rect 1639 1886 1669 1904
rect 1712 1874 1725 1904
rect 1755 1874 1768 1904
rect 1783 1886 1813 1904
rect 1856 1890 1870 1904
rect 1906 1890 2126 1904
rect 1857 1888 1870 1890
rect 1823 1876 1838 1888
rect 1820 1874 1842 1876
rect 1847 1874 1877 1888
rect 1938 1886 2091 1890
rect 1920 1874 2112 1886
rect 2155 1874 2185 1888
rect 2191 1874 2204 1904
rect 2219 1886 2249 1904
rect 2292 1874 2305 1904
rect 2335 1874 2348 1904
rect 2363 1886 2393 1904
rect 2436 1890 2450 1904
rect 2486 1890 2706 1904
rect 2437 1888 2450 1890
rect 2403 1876 2418 1888
rect 2400 1874 2422 1876
rect 2427 1874 2457 1888
rect 2518 1886 2671 1890
rect 2500 1874 2692 1886
rect 2735 1874 2765 1888
rect 2771 1874 2784 1904
rect 2799 1886 2829 1904
rect 2872 1874 2885 1904
rect 2915 1874 2928 1904
rect 2943 1886 2973 1904
rect 3016 1890 3030 1904
rect 3066 1890 3286 1904
rect 3017 1888 3030 1890
rect 2983 1876 2998 1888
rect 2980 1874 3002 1876
rect 3007 1874 3037 1888
rect 3098 1886 3251 1890
rect 3080 1874 3272 1886
rect 3315 1874 3345 1888
rect 3351 1874 3364 1904
rect 3379 1886 3409 1904
rect 3452 1874 3465 1904
rect 3495 1874 3508 1904
rect 3523 1886 3553 1904
rect 3596 1890 3610 1904
rect 3646 1890 3866 1904
rect 3597 1888 3610 1890
rect 3563 1876 3578 1888
rect 3560 1874 3582 1876
rect 3587 1874 3617 1888
rect 3678 1886 3831 1890
rect 3660 1874 3852 1886
rect 3895 1874 3925 1888
rect 3931 1874 3944 1904
rect 3959 1886 3989 1904
rect 4032 1874 4045 1904
rect 4075 1874 4088 1904
rect 4103 1886 4133 1904
rect 4176 1890 4190 1904
rect 4226 1890 4446 1904
rect 4177 1888 4190 1890
rect 4143 1876 4158 1888
rect 4140 1874 4162 1876
rect 4167 1874 4197 1888
rect 4258 1886 4411 1890
rect 4240 1874 4432 1886
rect 4475 1874 4505 1888
rect 4511 1874 4524 1904
rect 4539 1886 4569 1904
rect 4612 1874 4625 1904
rect 0 1860 4625 1874
rect 15 1756 28 1860
rect 73 1838 74 1848
rect 89 1838 102 1848
rect 73 1834 102 1838
rect 107 1834 137 1860
rect 155 1846 171 1848
rect 243 1846 296 1860
rect 244 1844 308 1846
rect 351 1844 366 1860
rect 415 1857 445 1860
rect 415 1854 451 1857
rect 381 1846 397 1848
rect 155 1834 170 1838
rect 73 1832 170 1834
rect 198 1832 366 1844
rect 382 1834 397 1838
rect 415 1835 454 1854
rect 473 1848 480 1849
rect 479 1841 480 1848
rect 463 1838 464 1841
rect 479 1838 492 1841
rect 415 1834 445 1835
rect 454 1834 460 1835
rect 463 1834 492 1838
rect 382 1833 492 1834
rect 382 1832 498 1833
rect 57 1824 108 1832
rect 57 1812 82 1824
rect 89 1812 108 1824
rect 139 1824 189 1832
rect 139 1816 155 1824
rect 162 1822 189 1824
rect 198 1822 419 1832
rect 162 1812 419 1822
rect 448 1824 498 1832
rect 448 1815 464 1824
rect 57 1804 108 1812
rect 155 1804 419 1812
rect 445 1812 464 1815
rect 471 1812 498 1824
rect 445 1804 498 1812
rect 73 1796 74 1804
rect 89 1796 102 1804
rect 73 1788 89 1796
rect 70 1781 89 1784
rect 70 1772 92 1781
rect 43 1762 92 1772
rect 43 1756 73 1762
rect 92 1757 97 1762
rect 15 1740 89 1756
rect 107 1748 137 1804
rect 172 1794 380 1804
rect 415 1800 460 1804
rect 463 1803 464 1804
rect 479 1803 492 1804
rect 198 1764 387 1794
rect 213 1761 387 1764
rect 206 1758 387 1761
rect 15 1738 28 1740
rect 43 1738 77 1740
rect 15 1722 89 1738
rect 116 1734 129 1748
rect 144 1734 160 1750
rect 206 1745 217 1758
rect -1 1700 0 1716
rect 15 1700 28 1722
rect 43 1700 73 1722
rect 116 1718 178 1734
rect 206 1727 217 1743
rect 222 1738 232 1758
rect 242 1738 256 1758
rect 259 1745 268 1758
rect 284 1745 293 1758
rect 222 1727 256 1738
rect 259 1727 268 1743
rect 284 1727 293 1743
rect 300 1738 310 1758
rect 320 1738 334 1758
rect 335 1745 346 1758
rect 300 1727 334 1738
rect 335 1727 346 1743
rect 392 1734 408 1750
rect 415 1748 445 1800
rect 479 1796 480 1803
rect 464 1788 480 1796
rect 451 1756 464 1775
rect 479 1756 509 1772
rect 451 1740 525 1756
rect 451 1738 464 1740
rect 479 1738 513 1740
rect 116 1716 129 1718
rect 144 1716 178 1718
rect 116 1700 178 1716
rect 222 1711 238 1714
rect 300 1711 330 1722
rect 378 1718 424 1734
rect 451 1722 525 1738
rect 378 1716 412 1718
rect 377 1700 424 1716
rect 451 1700 464 1722
rect 479 1700 509 1722
rect 536 1700 537 1716
rect 552 1700 565 1860
rect 595 1756 608 1860
rect 653 1838 654 1848
rect 669 1838 682 1848
rect 653 1834 682 1838
rect 687 1834 717 1860
rect 735 1846 751 1848
rect 823 1846 876 1860
rect 824 1844 888 1846
rect 931 1844 946 1860
rect 995 1857 1025 1860
rect 995 1854 1031 1857
rect 961 1846 977 1848
rect 735 1834 750 1838
rect 653 1832 750 1834
rect 778 1832 946 1844
rect 962 1834 977 1838
rect 995 1835 1034 1854
rect 1053 1848 1060 1849
rect 1059 1841 1060 1848
rect 1043 1838 1044 1841
rect 1059 1838 1072 1841
rect 995 1834 1025 1835
rect 1034 1834 1040 1835
rect 1043 1834 1072 1838
rect 962 1833 1072 1834
rect 962 1832 1078 1833
rect 637 1824 688 1832
rect 637 1812 662 1824
rect 669 1812 688 1824
rect 719 1824 769 1832
rect 719 1816 735 1824
rect 742 1822 769 1824
rect 778 1822 999 1832
rect 742 1812 999 1822
rect 1028 1824 1078 1832
rect 1028 1815 1044 1824
rect 637 1804 688 1812
rect 735 1804 999 1812
rect 1025 1812 1044 1815
rect 1051 1812 1078 1824
rect 1025 1804 1078 1812
rect 653 1796 654 1804
rect 669 1796 682 1804
rect 653 1788 669 1796
rect 650 1781 669 1784
rect 650 1772 672 1781
rect 623 1762 672 1772
rect 623 1756 653 1762
rect 672 1757 677 1762
rect 595 1740 669 1756
rect 687 1748 717 1804
rect 752 1794 960 1804
rect 995 1800 1040 1804
rect 1043 1803 1044 1804
rect 1059 1803 1072 1804
rect 778 1764 967 1794
rect 793 1761 967 1764
rect 786 1758 967 1761
rect 595 1738 608 1740
rect 623 1738 657 1740
rect 595 1722 669 1738
rect 696 1734 709 1748
rect 724 1734 740 1750
rect 786 1745 797 1758
rect 579 1700 580 1716
rect 595 1700 608 1722
rect 623 1700 653 1722
rect 696 1718 758 1734
rect 786 1727 797 1743
rect 802 1738 812 1758
rect 822 1738 836 1758
rect 839 1745 848 1758
rect 864 1745 873 1758
rect 802 1727 836 1738
rect 839 1727 848 1743
rect 864 1727 873 1743
rect 880 1738 890 1758
rect 900 1738 914 1758
rect 915 1745 926 1758
rect 880 1727 914 1738
rect 915 1727 926 1743
rect 972 1734 988 1750
rect 995 1748 1025 1800
rect 1059 1796 1060 1803
rect 1044 1788 1060 1796
rect 1031 1756 1044 1775
rect 1059 1756 1089 1772
rect 1031 1740 1105 1756
rect 1031 1738 1044 1740
rect 1059 1738 1093 1740
rect 696 1716 709 1718
rect 724 1716 758 1718
rect 696 1700 758 1716
rect 802 1711 818 1714
rect 880 1711 910 1722
rect 958 1718 1004 1734
rect 1031 1722 1105 1738
rect 958 1716 992 1718
rect 957 1700 1004 1716
rect 1031 1700 1044 1722
rect 1059 1700 1089 1722
rect 1116 1700 1117 1716
rect 1132 1700 1145 1860
rect 1175 1756 1188 1860
rect 1233 1838 1234 1848
rect 1249 1838 1262 1848
rect 1233 1834 1262 1838
rect 1267 1834 1297 1860
rect 1315 1846 1331 1848
rect 1403 1846 1456 1860
rect 1404 1844 1468 1846
rect 1511 1844 1526 1860
rect 1575 1857 1605 1860
rect 1575 1854 1611 1857
rect 1541 1846 1557 1848
rect 1315 1834 1330 1838
rect 1233 1832 1330 1834
rect 1358 1832 1526 1844
rect 1542 1834 1557 1838
rect 1575 1835 1614 1854
rect 1633 1848 1640 1849
rect 1639 1841 1640 1848
rect 1623 1838 1624 1841
rect 1639 1838 1652 1841
rect 1575 1834 1605 1835
rect 1614 1834 1620 1835
rect 1623 1834 1652 1838
rect 1542 1833 1652 1834
rect 1542 1832 1658 1833
rect 1217 1824 1268 1832
rect 1217 1812 1242 1824
rect 1249 1812 1268 1824
rect 1299 1824 1349 1832
rect 1299 1816 1315 1824
rect 1322 1822 1349 1824
rect 1358 1822 1579 1832
rect 1322 1812 1579 1822
rect 1608 1824 1658 1832
rect 1608 1815 1624 1824
rect 1217 1804 1268 1812
rect 1315 1804 1579 1812
rect 1605 1812 1624 1815
rect 1631 1812 1658 1824
rect 1605 1804 1658 1812
rect 1233 1796 1234 1804
rect 1249 1796 1262 1804
rect 1233 1788 1249 1796
rect 1230 1781 1249 1784
rect 1230 1772 1252 1781
rect 1203 1762 1252 1772
rect 1203 1756 1233 1762
rect 1252 1757 1257 1762
rect 1175 1740 1249 1756
rect 1267 1748 1297 1804
rect 1332 1794 1540 1804
rect 1575 1800 1620 1804
rect 1623 1803 1624 1804
rect 1639 1803 1652 1804
rect 1358 1764 1547 1794
rect 1373 1761 1547 1764
rect 1366 1758 1547 1761
rect 1175 1738 1188 1740
rect 1203 1738 1237 1740
rect 1175 1722 1249 1738
rect 1276 1734 1289 1748
rect 1304 1734 1320 1750
rect 1366 1745 1377 1758
rect 1159 1700 1160 1716
rect 1175 1700 1188 1722
rect 1203 1700 1233 1722
rect 1276 1718 1338 1734
rect 1366 1727 1377 1743
rect 1382 1738 1392 1758
rect 1402 1738 1416 1758
rect 1419 1745 1428 1758
rect 1444 1745 1453 1758
rect 1382 1727 1416 1738
rect 1419 1727 1428 1743
rect 1444 1727 1453 1743
rect 1460 1738 1470 1758
rect 1480 1738 1494 1758
rect 1495 1745 1506 1758
rect 1460 1727 1494 1738
rect 1495 1727 1506 1743
rect 1552 1734 1568 1750
rect 1575 1748 1605 1800
rect 1639 1796 1640 1803
rect 1624 1788 1640 1796
rect 1611 1756 1624 1775
rect 1639 1756 1669 1772
rect 1611 1740 1685 1756
rect 1611 1738 1624 1740
rect 1639 1738 1673 1740
rect 1276 1716 1289 1718
rect 1304 1716 1338 1718
rect 1276 1700 1338 1716
rect 1382 1711 1398 1714
rect 1460 1711 1490 1722
rect 1538 1718 1584 1734
rect 1611 1722 1685 1738
rect 1538 1716 1572 1718
rect 1537 1700 1584 1716
rect 1611 1700 1624 1722
rect 1639 1700 1669 1722
rect 1696 1700 1697 1716
rect 1712 1700 1725 1860
rect 1755 1756 1768 1860
rect 1813 1838 1814 1848
rect 1829 1838 1842 1848
rect 1813 1834 1842 1838
rect 1847 1834 1877 1860
rect 1895 1846 1911 1848
rect 1983 1846 2036 1860
rect 1984 1844 2048 1846
rect 2091 1844 2106 1860
rect 2155 1857 2185 1860
rect 2155 1854 2191 1857
rect 2121 1846 2137 1848
rect 1895 1834 1910 1838
rect 1813 1832 1910 1834
rect 1938 1832 2106 1844
rect 2122 1834 2137 1838
rect 2155 1835 2194 1854
rect 2213 1848 2220 1849
rect 2219 1841 2220 1848
rect 2203 1838 2204 1841
rect 2219 1838 2232 1841
rect 2155 1834 2185 1835
rect 2194 1834 2200 1835
rect 2203 1834 2232 1838
rect 2122 1833 2232 1834
rect 2122 1832 2238 1833
rect 1797 1824 1848 1832
rect 1797 1812 1822 1824
rect 1829 1812 1848 1824
rect 1879 1824 1929 1832
rect 1879 1816 1895 1824
rect 1902 1822 1929 1824
rect 1938 1822 2159 1832
rect 1902 1812 2159 1822
rect 2188 1824 2238 1832
rect 2188 1815 2204 1824
rect 1797 1804 1848 1812
rect 1895 1804 2159 1812
rect 2185 1812 2204 1815
rect 2211 1812 2238 1824
rect 2185 1804 2238 1812
rect 1813 1796 1814 1804
rect 1829 1796 1842 1804
rect 1813 1788 1829 1796
rect 1810 1781 1829 1784
rect 1810 1772 1832 1781
rect 1783 1762 1832 1772
rect 1783 1756 1813 1762
rect 1832 1757 1837 1762
rect 1755 1740 1829 1756
rect 1847 1748 1877 1804
rect 1912 1794 2120 1804
rect 2155 1800 2200 1804
rect 2203 1803 2204 1804
rect 2219 1803 2232 1804
rect 1938 1764 2127 1794
rect 1953 1761 2127 1764
rect 1946 1758 2127 1761
rect 1755 1738 1768 1740
rect 1783 1738 1817 1740
rect 1755 1722 1829 1738
rect 1856 1734 1869 1748
rect 1884 1734 1900 1750
rect 1946 1745 1957 1758
rect 1739 1700 1740 1716
rect 1755 1700 1768 1722
rect 1783 1700 1813 1722
rect 1856 1718 1918 1734
rect 1946 1727 1957 1743
rect 1962 1738 1972 1758
rect 1982 1738 1996 1758
rect 1999 1745 2008 1758
rect 2024 1745 2033 1758
rect 1962 1727 1996 1738
rect 1999 1727 2008 1743
rect 2024 1727 2033 1743
rect 2040 1738 2050 1758
rect 2060 1738 2074 1758
rect 2075 1745 2086 1758
rect 2040 1727 2074 1738
rect 2075 1727 2086 1743
rect 2132 1734 2148 1750
rect 2155 1748 2185 1800
rect 2219 1796 2220 1803
rect 2204 1788 2220 1796
rect 2191 1756 2204 1775
rect 2219 1756 2249 1772
rect 2191 1740 2265 1756
rect 2191 1738 2204 1740
rect 2219 1738 2253 1740
rect 1856 1716 1869 1718
rect 1884 1716 1918 1718
rect 1856 1700 1918 1716
rect 1962 1711 1978 1714
rect 2040 1711 2070 1722
rect 2118 1718 2164 1734
rect 2191 1722 2265 1738
rect 2118 1716 2152 1718
rect 2117 1700 2164 1716
rect 2191 1700 2204 1722
rect 2219 1700 2249 1722
rect 2276 1700 2277 1716
rect 2292 1700 2305 1860
rect 2335 1756 2348 1860
rect 2393 1838 2394 1848
rect 2409 1838 2422 1848
rect 2393 1834 2422 1838
rect 2427 1834 2457 1860
rect 2475 1846 2491 1848
rect 2563 1846 2616 1860
rect 2564 1844 2628 1846
rect 2671 1844 2686 1860
rect 2735 1857 2765 1860
rect 2735 1854 2771 1857
rect 2701 1846 2717 1848
rect 2475 1834 2490 1838
rect 2393 1832 2490 1834
rect 2518 1832 2686 1844
rect 2702 1834 2717 1838
rect 2735 1835 2774 1854
rect 2793 1848 2800 1849
rect 2799 1841 2800 1848
rect 2783 1838 2784 1841
rect 2799 1838 2812 1841
rect 2735 1834 2765 1835
rect 2774 1834 2780 1835
rect 2783 1834 2812 1838
rect 2702 1833 2812 1834
rect 2702 1832 2818 1833
rect 2377 1824 2428 1832
rect 2377 1812 2402 1824
rect 2409 1812 2428 1824
rect 2459 1824 2509 1832
rect 2459 1816 2475 1824
rect 2482 1822 2509 1824
rect 2518 1822 2739 1832
rect 2482 1812 2739 1822
rect 2768 1824 2818 1832
rect 2768 1815 2784 1824
rect 2377 1804 2428 1812
rect 2475 1804 2739 1812
rect 2765 1812 2784 1815
rect 2791 1812 2818 1824
rect 2765 1804 2818 1812
rect 2393 1796 2394 1804
rect 2409 1796 2422 1804
rect 2393 1788 2409 1796
rect 2390 1781 2409 1784
rect 2390 1772 2412 1781
rect 2363 1762 2412 1772
rect 2363 1756 2393 1762
rect 2412 1757 2417 1762
rect 2335 1740 2409 1756
rect 2427 1748 2457 1804
rect 2492 1794 2700 1804
rect 2735 1800 2780 1804
rect 2783 1803 2784 1804
rect 2799 1803 2812 1804
rect 2518 1764 2707 1794
rect 2533 1761 2707 1764
rect 2526 1758 2707 1761
rect 2335 1738 2348 1740
rect 2363 1738 2397 1740
rect 2335 1722 2409 1738
rect 2436 1734 2449 1748
rect 2464 1734 2480 1750
rect 2526 1745 2537 1758
rect 2319 1700 2320 1716
rect 2335 1700 2348 1722
rect 2363 1700 2393 1722
rect 2436 1718 2498 1734
rect 2526 1727 2537 1743
rect 2542 1738 2552 1758
rect 2562 1738 2576 1758
rect 2579 1745 2588 1758
rect 2604 1745 2613 1758
rect 2542 1727 2576 1738
rect 2579 1727 2588 1743
rect 2604 1727 2613 1743
rect 2620 1738 2630 1758
rect 2640 1738 2654 1758
rect 2655 1745 2666 1758
rect 2620 1727 2654 1738
rect 2655 1727 2666 1743
rect 2712 1734 2728 1750
rect 2735 1748 2765 1800
rect 2799 1796 2800 1803
rect 2784 1788 2800 1796
rect 2771 1756 2784 1775
rect 2799 1756 2829 1772
rect 2771 1740 2845 1756
rect 2771 1738 2784 1740
rect 2799 1738 2833 1740
rect 2436 1716 2449 1718
rect 2464 1716 2498 1718
rect 2436 1700 2498 1716
rect 2542 1711 2558 1714
rect 2620 1711 2650 1722
rect 2698 1718 2744 1734
rect 2771 1722 2845 1738
rect 2698 1716 2732 1718
rect 2697 1700 2744 1716
rect 2771 1700 2784 1722
rect 2799 1700 2829 1722
rect 2856 1700 2857 1716
rect 2872 1700 2885 1860
rect 2915 1756 2928 1860
rect 2973 1838 2974 1848
rect 2989 1838 3002 1848
rect 2973 1834 3002 1838
rect 3007 1834 3037 1860
rect 3055 1846 3071 1848
rect 3143 1846 3196 1860
rect 3144 1844 3208 1846
rect 3251 1844 3266 1860
rect 3315 1857 3345 1860
rect 3315 1854 3351 1857
rect 3281 1846 3297 1848
rect 3055 1834 3070 1838
rect 2973 1832 3070 1834
rect 3098 1832 3266 1844
rect 3282 1834 3297 1838
rect 3315 1835 3354 1854
rect 3373 1848 3380 1849
rect 3379 1841 3380 1848
rect 3363 1838 3364 1841
rect 3379 1838 3392 1841
rect 3315 1834 3345 1835
rect 3354 1834 3360 1835
rect 3363 1834 3392 1838
rect 3282 1833 3392 1834
rect 3282 1832 3398 1833
rect 2957 1824 3008 1832
rect 2957 1812 2982 1824
rect 2989 1812 3008 1824
rect 3039 1824 3089 1832
rect 3039 1816 3055 1824
rect 3062 1822 3089 1824
rect 3098 1822 3319 1832
rect 3062 1812 3319 1822
rect 3348 1824 3398 1832
rect 3348 1815 3364 1824
rect 2957 1804 3008 1812
rect 3055 1804 3319 1812
rect 3345 1812 3364 1815
rect 3371 1812 3398 1824
rect 3345 1804 3398 1812
rect 2973 1796 2974 1804
rect 2989 1796 3002 1804
rect 2973 1788 2989 1796
rect 2970 1781 2989 1784
rect 2970 1772 2992 1781
rect 2943 1762 2992 1772
rect 2943 1756 2973 1762
rect 2992 1757 2997 1762
rect 2915 1740 2989 1756
rect 3007 1748 3037 1804
rect 3072 1794 3280 1804
rect 3315 1800 3360 1804
rect 3363 1803 3364 1804
rect 3379 1803 3392 1804
rect 3098 1764 3287 1794
rect 3113 1761 3287 1764
rect 3106 1758 3287 1761
rect 2915 1738 2928 1740
rect 2943 1738 2977 1740
rect 2915 1722 2989 1738
rect 3016 1734 3029 1748
rect 3044 1734 3060 1750
rect 3106 1745 3117 1758
rect 2899 1700 2900 1716
rect 2915 1700 2928 1722
rect 2943 1700 2973 1722
rect 3016 1718 3078 1734
rect 3106 1727 3117 1743
rect 3122 1738 3132 1758
rect 3142 1738 3156 1758
rect 3159 1745 3168 1758
rect 3184 1745 3193 1758
rect 3122 1727 3156 1738
rect 3159 1727 3168 1743
rect 3184 1727 3193 1743
rect 3200 1738 3210 1758
rect 3220 1738 3234 1758
rect 3235 1745 3246 1758
rect 3200 1727 3234 1738
rect 3235 1727 3246 1743
rect 3292 1734 3308 1750
rect 3315 1748 3345 1800
rect 3379 1796 3380 1803
rect 3364 1788 3380 1796
rect 3351 1756 3364 1775
rect 3379 1756 3409 1772
rect 3351 1740 3425 1756
rect 3351 1738 3364 1740
rect 3379 1738 3413 1740
rect 3016 1716 3029 1718
rect 3044 1716 3078 1718
rect 3016 1700 3078 1716
rect 3122 1711 3138 1714
rect 3200 1711 3230 1722
rect 3278 1718 3324 1734
rect 3351 1722 3425 1738
rect 3278 1716 3312 1718
rect 3277 1700 3324 1716
rect 3351 1700 3364 1722
rect 3379 1700 3409 1722
rect 3436 1700 3437 1716
rect 3452 1700 3465 1860
rect 3495 1756 3508 1860
rect 3553 1838 3554 1848
rect 3569 1838 3582 1848
rect 3553 1834 3582 1838
rect 3587 1834 3617 1860
rect 3635 1846 3651 1848
rect 3723 1846 3776 1860
rect 3724 1844 3788 1846
rect 3831 1844 3846 1860
rect 3895 1857 3925 1860
rect 3895 1854 3931 1857
rect 3861 1846 3877 1848
rect 3635 1834 3650 1838
rect 3553 1832 3650 1834
rect 3678 1832 3846 1844
rect 3862 1834 3877 1838
rect 3895 1835 3934 1854
rect 3953 1848 3960 1849
rect 3959 1841 3960 1848
rect 3943 1838 3944 1841
rect 3959 1838 3972 1841
rect 3895 1834 3925 1835
rect 3934 1834 3940 1835
rect 3943 1834 3972 1838
rect 3862 1833 3972 1834
rect 3862 1832 3978 1833
rect 3537 1824 3588 1832
rect 3537 1812 3562 1824
rect 3569 1812 3588 1824
rect 3619 1824 3669 1832
rect 3619 1816 3635 1824
rect 3642 1822 3669 1824
rect 3678 1822 3899 1832
rect 3642 1812 3899 1822
rect 3928 1824 3978 1832
rect 3928 1815 3944 1824
rect 3537 1804 3588 1812
rect 3635 1804 3899 1812
rect 3925 1812 3944 1815
rect 3951 1812 3978 1824
rect 3925 1804 3978 1812
rect 3553 1796 3554 1804
rect 3569 1796 3582 1804
rect 3553 1788 3569 1796
rect 3550 1781 3569 1784
rect 3550 1772 3572 1781
rect 3523 1762 3572 1772
rect 3523 1756 3553 1762
rect 3572 1757 3577 1762
rect 3495 1740 3569 1756
rect 3587 1748 3617 1804
rect 3652 1794 3860 1804
rect 3895 1800 3940 1804
rect 3943 1803 3944 1804
rect 3959 1803 3972 1804
rect 3678 1764 3867 1794
rect 3693 1761 3867 1764
rect 3686 1758 3867 1761
rect 3495 1738 3508 1740
rect 3523 1738 3557 1740
rect 3495 1722 3569 1738
rect 3596 1734 3609 1748
rect 3624 1734 3640 1750
rect 3686 1745 3697 1758
rect 3479 1700 3480 1716
rect 3495 1700 3508 1722
rect 3523 1700 3553 1722
rect 3596 1718 3658 1734
rect 3686 1727 3697 1743
rect 3702 1738 3712 1758
rect 3722 1738 3736 1758
rect 3739 1745 3748 1758
rect 3764 1745 3773 1758
rect 3702 1727 3736 1738
rect 3739 1727 3748 1743
rect 3764 1727 3773 1743
rect 3780 1738 3790 1758
rect 3800 1738 3814 1758
rect 3815 1745 3826 1758
rect 3780 1727 3814 1738
rect 3815 1727 3826 1743
rect 3872 1734 3888 1750
rect 3895 1748 3925 1800
rect 3959 1796 3960 1803
rect 3944 1788 3960 1796
rect 3931 1756 3944 1775
rect 3959 1756 3989 1772
rect 3931 1740 4005 1756
rect 3931 1738 3944 1740
rect 3959 1738 3993 1740
rect 3596 1716 3609 1718
rect 3624 1716 3658 1718
rect 3596 1700 3658 1716
rect 3702 1711 3718 1714
rect 3780 1711 3810 1722
rect 3858 1718 3904 1734
rect 3931 1722 4005 1738
rect 3858 1716 3892 1718
rect 3857 1700 3904 1716
rect 3931 1700 3944 1722
rect 3959 1700 3989 1722
rect 4016 1700 4017 1716
rect 4032 1700 4045 1860
rect 4075 1756 4088 1860
rect 4133 1838 4134 1848
rect 4149 1838 4162 1848
rect 4133 1834 4162 1838
rect 4167 1834 4197 1860
rect 4215 1846 4231 1848
rect 4303 1846 4356 1860
rect 4304 1844 4368 1846
rect 4411 1844 4426 1860
rect 4475 1857 4505 1860
rect 4475 1854 4511 1857
rect 4441 1846 4457 1848
rect 4215 1834 4230 1838
rect 4133 1832 4230 1834
rect 4258 1832 4426 1844
rect 4442 1834 4457 1838
rect 4475 1835 4514 1854
rect 4533 1848 4540 1849
rect 4539 1841 4540 1848
rect 4523 1838 4524 1841
rect 4539 1838 4552 1841
rect 4475 1834 4505 1835
rect 4514 1834 4520 1835
rect 4523 1834 4552 1838
rect 4442 1833 4552 1834
rect 4442 1832 4558 1833
rect 4117 1824 4168 1832
rect 4117 1812 4142 1824
rect 4149 1812 4168 1824
rect 4199 1824 4249 1832
rect 4199 1816 4215 1824
rect 4222 1822 4249 1824
rect 4258 1822 4479 1832
rect 4222 1812 4479 1822
rect 4508 1824 4558 1832
rect 4508 1815 4524 1824
rect 4117 1804 4168 1812
rect 4215 1804 4479 1812
rect 4505 1812 4524 1815
rect 4531 1812 4558 1824
rect 4505 1804 4558 1812
rect 4133 1796 4134 1804
rect 4149 1796 4162 1804
rect 4133 1788 4149 1796
rect 4130 1781 4149 1784
rect 4130 1772 4152 1781
rect 4103 1762 4152 1772
rect 4103 1756 4133 1762
rect 4152 1757 4157 1762
rect 4075 1740 4149 1756
rect 4167 1748 4197 1804
rect 4232 1794 4440 1804
rect 4475 1800 4520 1804
rect 4523 1803 4524 1804
rect 4539 1803 4552 1804
rect 4258 1764 4447 1794
rect 4273 1761 4447 1764
rect 4266 1758 4447 1761
rect 4075 1738 4088 1740
rect 4103 1738 4137 1740
rect 4075 1722 4149 1738
rect 4176 1734 4189 1748
rect 4204 1734 4220 1750
rect 4266 1745 4277 1758
rect 4059 1700 4060 1716
rect 4075 1700 4088 1722
rect 4103 1700 4133 1722
rect 4176 1718 4238 1734
rect 4266 1727 4277 1743
rect 4282 1738 4292 1758
rect 4302 1738 4316 1758
rect 4319 1745 4328 1758
rect 4344 1745 4353 1758
rect 4282 1727 4316 1738
rect 4319 1727 4328 1743
rect 4344 1727 4353 1743
rect 4360 1738 4370 1758
rect 4380 1738 4394 1758
rect 4395 1745 4406 1758
rect 4360 1727 4394 1738
rect 4395 1727 4406 1743
rect 4452 1734 4468 1750
rect 4475 1748 4505 1800
rect 4539 1796 4540 1803
rect 4524 1788 4540 1796
rect 4511 1756 4524 1775
rect 4539 1756 4569 1772
rect 4511 1740 4585 1756
rect 4511 1738 4524 1740
rect 4539 1738 4573 1740
rect 4176 1716 4189 1718
rect 4204 1716 4238 1718
rect 4176 1700 4238 1716
rect 4282 1711 4298 1714
rect 4360 1711 4390 1722
rect 4438 1718 4484 1734
rect 4511 1722 4585 1738
rect 4438 1716 4472 1718
rect 4437 1700 4484 1716
rect 4511 1700 4524 1722
rect 4539 1700 4569 1722
rect 4596 1700 4597 1716
rect 4612 1700 4625 1860
rect -7 1692 34 1700
rect -7 1666 8 1692
rect 15 1666 34 1692
rect 98 1688 160 1700
rect 172 1688 247 1700
rect 305 1688 380 1700
rect 392 1688 423 1700
rect 429 1688 464 1700
rect 98 1686 260 1688
rect -7 1658 34 1666
rect 116 1662 129 1686
rect 144 1684 159 1686
rect -1 1648 0 1658
rect 15 1648 28 1658
rect 43 1648 73 1662
rect 116 1648 159 1662
rect 183 1659 190 1666
rect 193 1662 260 1686
rect 292 1686 464 1688
rect 262 1664 290 1668
rect 292 1664 372 1686
rect 393 1684 408 1686
rect 262 1662 372 1664
rect 193 1658 372 1662
rect 166 1648 196 1658
rect 198 1648 351 1658
rect 359 1648 389 1658
rect 393 1648 423 1662
rect 451 1648 464 1686
rect 536 1692 571 1700
rect 536 1666 537 1692
rect 544 1666 571 1692
rect 479 1648 509 1662
rect 536 1658 571 1666
rect 573 1692 614 1700
rect 573 1666 588 1692
rect 595 1666 614 1692
rect 678 1688 740 1700
rect 752 1688 827 1700
rect 885 1688 960 1700
rect 972 1688 1003 1700
rect 1009 1688 1044 1700
rect 678 1686 840 1688
rect 573 1658 614 1666
rect 696 1662 709 1686
rect 724 1684 739 1686
rect 536 1648 537 1658
rect 552 1648 565 1658
rect 579 1648 580 1658
rect 595 1648 608 1658
rect 623 1648 653 1662
rect 696 1648 739 1662
rect 763 1659 770 1666
rect 773 1662 840 1686
rect 872 1686 1044 1688
rect 842 1664 870 1668
rect 872 1664 952 1686
rect 973 1684 988 1686
rect 842 1662 952 1664
rect 773 1658 952 1662
rect 746 1648 776 1658
rect 778 1648 931 1658
rect 939 1648 969 1658
rect 973 1648 1003 1662
rect 1031 1648 1044 1686
rect 1116 1692 1151 1700
rect 1116 1666 1117 1692
rect 1124 1666 1151 1692
rect 1059 1648 1089 1662
rect 1116 1658 1151 1666
rect 1153 1692 1194 1700
rect 1153 1666 1168 1692
rect 1175 1666 1194 1692
rect 1258 1688 1320 1700
rect 1332 1688 1407 1700
rect 1465 1688 1540 1700
rect 1552 1688 1583 1700
rect 1589 1688 1624 1700
rect 1258 1686 1420 1688
rect 1153 1658 1194 1666
rect 1276 1662 1289 1686
rect 1304 1684 1319 1686
rect 1116 1648 1117 1658
rect 1132 1648 1145 1658
rect 1159 1648 1160 1658
rect 1175 1648 1188 1658
rect 1203 1648 1233 1662
rect 1276 1648 1319 1662
rect 1343 1659 1350 1666
rect 1353 1662 1420 1686
rect 1452 1686 1624 1688
rect 1422 1664 1450 1668
rect 1452 1664 1532 1686
rect 1553 1684 1568 1686
rect 1422 1662 1532 1664
rect 1353 1658 1532 1662
rect 1326 1648 1356 1658
rect 1358 1648 1511 1658
rect 1519 1648 1549 1658
rect 1553 1648 1583 1662
rect 1611 1648 1624 1686
rect 1696 1692 1731 1700
rect 1696 1666 1697 1692
rect 1704 1666 1731 1692
rect 1639 1648 1669 1662
rect 1696 1658 1731 1666
rect 1733 1692 1774 1700
rect 1733 1666 1748 1692
rect 1755 1666 1774 1692
rect 1838 1688 1900 1700
rect 1912 1688 1987 1700
rect 2045 1688 2120 1700
rect 2132 1688 2163 1700
rect 2169 1688 2204 1700
rect 1838 1686 2000 1688
rect 1733 1658 1774 1666
rect 1856 1662 1869 1686
rect 1884 1684 1899 1686
rect 1696 1648 1697 1658
rect 1712 1648 1725 1658
rect 1739 1648 1740 1658
rect 1755 1648 1768 1658
rect 1783 1648 1813 1662
rect 1856 1648 1899 1662
rect 1923 1659 1930 1666
rect 1933 1662 2000 1686
rect 2032 1686 2204 1688
rect 2002 1664 2030 1668
rect 2032 1664 2112 1686
rect 2133 1684 2148 1686
rect 2002 1662 2112 1664
rect 1933 1658 2112 1662
rect 1906 1648 1936 1658
rect 1938 1648 2091 1658
rect 2099 1648 2129 1658
rect 2133 1648 2163 1662
rect 2191 1648 2204 1686
rect 2276 1692 2311 1700
rect 2276 1666 2277 1692
rect 2284 1666 2311 1692
rect 2219 1648 2249 1662
rect 2276 1658 2311 1666
rect 2313 1692 2354 1700
rect 2313 1666 2328 1692
rect 2335 1666 2354 1692
rect 2418 1688 2480 1700
rect 2492 1688 2567 1700
rect 2625 1688 2700 1700
rect 2712 1688 2743 1700
rect 2749 1688 2784 1700
rect 2418 1686 2580 1688
rect 2313 1658 2354 1666
rect 2436 1662 2449 1686
rect 2464 1684 2479 1686
rect 2276 1648 2277 1658
rect 2292 1648 2305 1658
rect 2319 1648 2320 1658
rect 2335 1648 2348 1658
rect 2363 1648 2393 1662
rect 2436 1648 2479 1662
rect 2503 1659 2510 1666
rect 2513 1662 2580 1686
rect 2612 1686 2784 1688
rect 2582 1664 2610 1668
rect 2612 1664 2692 1686
rect 2713 1684 2728 1686
rect 2582 1662 2692 1664
rect 2513 1658 2692 1662
rect 2486 1648 2516 1658
rect 2518 1648 2671 1658
rect 2679 1648 2709 1658
rect 2713 1648 2743 1662
rect 2771 1648 2784 1686
rect 2856 1692 2891 1700
rect 2856 1666 2857 1692
rect 2864 1666 2891 1692
rect 2799 1648 2829 1662
rect 2856 1658 2891 1666
rect 2893 1692 2934 1700
rect 2893 1666 2908 1692
rect 2915 1666 2934 1692
rect 2998 1688 3060 1700
rect 3072 1688 3147 1700
rect 3205 1688 3280 1700
rect 3292 1688 3323 1700
rect 3329 1688 3364 1700
rect 2998 1686 3160 1688
rect 2893 1658 2934 1666
rect 3016 1662 3029 1686
rect 3044 1684 3059 1686
rect 2856 1648 2857 1658
rect 2872 1648 2885 1658
rect 2899 1648 2900 1658
rect 2915 1648 2928 1658
rect 2943 1648 2973 1662
rect 3016 1648 3059 1662
rect 3083 1659 3090 1666
rect 3093 1662 3160 1686
rect 3192 1686 3364 1688
rect 3162 1664 3190 1668
rect 3192 1664 3272 1686
rect 3293 1684 3308 1686
rect 3162 1662 3272 1664
rect 3093 1658 3272 1662
rect 3066 1648 3096 1658
rect 3098 1648 3251 1658
rect 3259 1648 3289 1658
rect 3293 1648 3323 1662
rect 3351 1648 3364 1686
rect 3436 1692 3471 1700
rect 3436 1666 3437 1692
rect 3444 1666 3471 1692
rect 3379 1648 3409 1662
rect 3436 1658 3471 1666
rect 3473 1692 3514 1700
rect 3473 1666 3488 1692
rect 3495 1666 3514 1692
rect 3578 1688 3640 1700
rect 3652 1688 3727 1700
rect 3785 1688 3860 1700
rect 3872 1688 3903 1700
rect 3909 1688 3944 1700
rect 3578 1686 3740 1688
rect 3473 1658 3514 1666
rect 3596 1662 3609 1686
rect 3624 1684 3639 1686
rect 3436 1648 3437 1658
rect 3452 1648 3465 1658
rect 3479 1648 3480 1658
rect 3495 1648 3508 1658
rect 3523 1648 3553 1662
rect 3596 1648 3639 1662
rect 3663 1659 3670 1666
rect 3673 1662 3740 1686
rect 3772 1686 3944 1688
rect 3742 1664 3770 1668
rect 3772 1664 3852 1686
rect 3873 1684 3888 1686
rect 3742 1662 3852 1664
rect 3673 1658 3852 1662
rect 3646 1648 3676 1658
rect 3678 1648 3831 1658
rect 3839 1648 3869 1658
rect 3873 1648 3903 1662
rect 3931 1648 3944 1686
rect 4016 1692 4051 1700
rect 4016 1666 4017 1692
rect 4024 1666 4051 1692
rect 3959 1648 3989 1662
rect 4016 1658 4051 1666
rect 4053 1692 4094 1700
rect 4053 1666 4068 1692
rect 4075 1666 4094 1692
rect 4158 1688 4220 1700
rect 4232 1688 4307 1700
rect 4365 1688 4440 1700
rect 4452 1688 4483 1700
rect 4489 1688 4524 1700
rect 4158 1686 4320 1688
rect 4053 1658 4094 1666
rect 4176 1662 4189 1686
rect 4204 1684 4219 1686
rect 4016 1648 4017 1658
rect 4032 1648 4045 1658
rect 4059 1648 4060 1658
rect 4075 1648 4088 1658
rect 4103 1648 4133 1662
rect 4176 1648 4219 1662
rect 4243 1659 4250 1666
rect 4253 1662 4320 1686
rect 4352 1686 4524 1688
rect 4322 1664 4350 1668
rect 4352 1664 4432 1686
rect 4453 1684 4468 1686
rect 4322 1662 4432 1664
rect 4253 1658 4432 1662
rect 4226 1648 4256 1658
rect 4258 1648 4411 1658
rect 4419 1648 4449 1658
rect 4453 1648 4483 1662
rect 4511 1648 4524 1686
rect 4596 1692 4631 1700
rect 4596 1666 4597 1692
rect 4604 1666 4631 1692
rect 4539 1648 4569 1662
rect 4596 1658 4631 1666
rect 4596 1648 4597 1658
rect 4612 1648 4625 1658
rect -1 1642 4625 1648
rect 0 1634 4625 1642
rect 15 1604 28 1634
rect 43 1616 73 1634
rect 116 1620 130 1634
rect 166 1620 386 1634
rect 117 1618 130 1620
rect 83 1606 98 1618
rect 80 1604 102 1606
rect 107 1604 137 1618
rect 198 1616 351 1620
rect 180 1604 372 1616
rect 415 1604 445 1618
rect 451 1604 464 1634
rect 479 1616 509 1634
rect 552 1604 565 1634
rect 595 1604 608 1634
rect 623 1616 653 1634
rect 696 1620 710 1634
rect 746 1620 966 1634
rect 697 1618 710 1620
rect 663 1606 678 1618
rect 660 1604 682 1606
rect 687 1604 717 1618
rect 778 1616 931 1620
rect 760 1604 952 1616
rect 995 1604 1025 1618
rect 1031 1604 1044 1634
rect 1059 1616 1089 1634
rect 1132 1604 1145 1634
rect 1175 1604 1188 1634
rect 1203 1616 1233 1634
rect 1276 1620 1290 1634
rect 1326 1620 1546 1634
rect 1277 1618 1290 1620
rect 1243 1606 1258 1618
rect 1240 1604 1262 1606
rect 1267 1604 1297 1618
rect 1358 1616 1511 1620
rect 1340 1604 1532 1616
rect 1575 1604 1605 1618
rect 1611 1604 1624 1634
rect 1639 1616 1669 1634
rect 1712 1604 1725 1634
rect 1755 1604 1768 1634
rect 1783 1616 1813 1634
rect 1856 1620 1870 1634
rect 1906 1620 2126 1634
rect 1857 1618 1870 1620
rect 1823 1606 1838 1618
rect 1820 1604 1842 1606
rect 1847 1604 1877 1618
rect 1938 1616 2091 1620
rect 1920 1604 2112 1616
rect 2155 1604 2185 1618
rect 2191 1604 2204 1634
rect 2219 1616 2249 1634
rect 2292 1604 2305 1634
rect 2335 1604 2348 1634
rect 2363 1616 2393 1634
rect 2436 1620 2450 1634
rect 2486 1620 2706 1634
rect 2437 1618 2450 1620
rect 2403 1606 2418 1618
rect 2400 1604 2422 1606
rect 2427 1604 2457 1618
rect 2518 1616 2671 1620
rect 2500 1604 2692 1616
rect 2735 1604 2765 1618
rect 2771 1604 2784 1634
rect 2799 1616 2829 1634
rect 2872 1604 2885 1634
rect 2915 1604 2928 1634
rect 2943 1616 2973 1634
rect 3016 1620 3030 1634
rect 3066 1620 3286 1634
rect 3017 1618 3030 1620
rect 2983 1606 2998 1618
rect 2980 1604 3002 1606
rect 3007 1604 3037 1618
rect 3098 1616 3251 1620
rect 3080 1604 3272 1616
rect 3315 1604 3345 1618
rect 3351 1604 3364 1634
rect 3379 1616 3409 1634
rect 3452 1604 3465 1634
rect 3495 1604 3508 1634
rect 3523 1616 3553 1634
rect 3596 1620 3610 1634
rect 3646 1620 3866 1634
rect 3597 1618 3610 1620
rect 3563 1606 3578 1618
rect 3560 1604 3582 1606
rect 3587 1604 3617 1618
rect 3678 1616 3831 1620
rect 3660 1604 3852 1616
rect 3895 1604 3925 1618
rect 3931 1604 3944 1634
rect 3959 1616 3989 1634
rect 4032 1604 4045 1634
rect 4075 1604 4088 1634
rect 4103 1616 4133 1634
rect 4176 1620 4190 1634
rect 4226 1620 4446 1634
rect 4177 1618 4190 1620
rect 4143 1606 4158 1618
rect 4140 1604 4162 1606
rect 4167 1604 4197 1618
rect 4258 1616 4411 1620
rect 4240 1604 4432 1616
rect 4475 1604 4505 1618
rect 4511 1604 4524 1634
rect 4539 1616 4569 1634
rect 4612 1604 4625 1634
rect 0 1590 4625 1604
rect 15 1486 28 1590
rect 73 1568 74 1578
rect 89 1568 102 1578
rect 73 1564 102 1568
rect 107 1564 137 1590
rect 155 1576 171 1578
rect 243 1576 296 1590
rect 244 1574 308 1576
rect 351 1574 366 1590
rect 415 1587 445 1590
rect 415 1584 451 1587
rect 381 1576 397 1578
rect 155 1564 170 1568
rect 73 1562 170 1564
rect 198 1562 366 1574
rect 382 1564 397 1568
rect 415 1565 454 1584
rect 473 1578 480 1579
rect 479 1571 480 1578
rect 463 1568 464 1571
rect 479 1568 492 1571
rect 415 1564 445 1565
rect 454 1564 460 1565
rect 463 1564 492 1568
rect 382 1563 492 1564
rect 382 1562 498 1563
rect 57 1554 108 1562
rect 57 1542 82 1554
rect 89 1542 108 1554
rect 139 1554 189 1562
rect 139 1546 155 1554
rect 162 1552 189 1554
rect 198 1552 419 1562
rect 162 1542 419 1552
rect 448 1554 498 1562
rect 448 1545 464 1554
rect 57 1534 108 1542
rect 155 1534 419 1542
rect 445 1542 464 1545
rect 471 1542 498 1554
rect 445 1534 498 1542
rect 73 1526 74 1534
rect 89 1526 102 1534
rect 73 1518 89 1526
rect 70 1511 89 1514
rect 70 1502 92 1511
rect 43 1492 92 1502
rect 43 1486 73 1492
rect 92 1487 97 1492
rect 15 1470 89 1486
rect 107 1478 137 1534
rect 172 1524 380 1534
rect 415 1530 460 1534
rect 463 1533 464 1534
rect 479 1533 492 1534
rect 198 1494 387 1524
rect 213 1491 387 1494
rect 206 1488 387 1491
rect 15 1468 28 1470
rect 43 1468 77 1470
rect 15 1452 89 1468
rect 116 1464 129 1478
rect 144 1464 160 1480
rect 206 1475 217 1488
rect -1 1430 0 1446
rect 15 1430 28 1452
rect 43 1430 73 1452
rect 116 1448 178 1464
rect 206 1457 217 1473
rect 222 1468 232 1488
rect 242 1468 256 1488
rect 259 1475 268 1488
rect 284 1475 293 1488
rect 222 1457 256 1468
rect 259 1457 268 1473
rect 284 1457 293 1473
rect 300 1468 310 1488
rect 320 1468 334 1488
rect 335 1475 346 1488
rect 300 1457 334 1468
rect 335 1457 346 1473
rect 392 1464 408 1480
rect 415 1478 445 1530
rect 479 1526 480 1533
rect 464 1518 480 1526
rect 451 1486 464 1505
rect 479 1486 509 1502
rect 451 1470 525 1486
rect 451 1468 464 1470
rect 479 1468 513 1470
rect 116 1446 129 1448
rect 144 1446 178 1448
rect 116 1430 178 1446
rect 222 1441 238 1444
rect 300 1441 330 1452
rect 378 1448 424 1464
rect 451 1452 525 1468
rect 378 1446 412 1448
rect 377 1430 424 1446
rect 451 1430 464 1452
rect 479 1430 509 1452
rect 536 1430 537 1446
rect 552 1430 565 1590
rect 595 1486 608 1590
rect 653 1568 654 1578
rect 669 1568 682 1578
rect 653 1564 682 1568
rect 687 1564 717 1590
rect 735 1576 751 1578
rect 823 1576 876 1590
rect 824 1574 888 1576
rect 931 1574 946 1590
rect 995 1587 1025 1590
rect 995 1584 1031 1587
rect 961 1576 977 1578
rect 735 1564 750 1568
rect 653 1562 750 1564
rect 778 1562 946 1574
rect 962 1564 977 1568
rect 995 1565 1034 1584
rect 1053 1578 1060 1579
rect 1059 1571 1060 1578
rect 1043 1568 1044 1571
rect 1059 1568 1072 1571
rect 995 1564 1025 1565
rect 1034 1564 1040 1565
rect 1043 1564 1072 1568
rect 962 1563 1072 1564
rect 962 1562 1078 1563
rect 637 1554 688 1562
rect 637 1542 662 1554
rect 669 1542 688 1554
rect 719 1554 769 1562
rect 719 1546 735 1554
rect 742 1552 769 1554
rect 778 1552 999 1562
rect 742 1542 999 1552
rect 1028 1554 1078 1562
rect 1028 1545 1044 1554
rect 637 1534 688 1542
rect 735 1534 999 1542
rect 1025 1542 1044 1545
rect 1051 1542 1078 1554
rect 1025 1534 1078 1542
rect 653 1526 654 1534
rect 669 1526 682 1534
rect 653 1518 669 1526
rect 650 1511 669 1514
rect 650 1502 672 1511
rect 623 1492 672 1502
rect 623 1486 653 1492
rect 672 1487 677 1492
rect 595 1470 669 1486
rect 687 1478 717 1534
rect 752 1524 960 1534
rect 995 1530 1040 1534
rect 1043 1533 1044 1534
rect 1059 1533 1072 1534
rect 778 1494 967 1524
rect 793 1491 967 1494
rect 786 1488 967 1491
rect 595 1468 608 1470
rect 623 1468 657 1470
rect 595 1452 669 1468
rect 696 1464 709 1478
rect 724 1464 740 1480
rect 786 1475 797 1488
rect 579 1430 580 1446
rect 595 1430 608 1452
rect 623 1430 653 1452
rect 696 1448 758 1464
rect 786 1457 797 1473
rect 802 1468 812 1488
rect 822 1468 836 1488
rect 839 1475 848 1488
rect 864 1475 873 1488
rect 802 1457 836 1468
rect 839 1457 848 1473
rect 864 1457 873 1473
rect 880 1468 890 1488
rect 900 1468 914 1488
rect 915 1475 926 1488
rect 880 1457 914 1468
rect 915 1457 926 1473
rect 972 1464 988 1480
rect 995 1478 1025 1530
rect 1059 1526 1060 1533
rect 1044 1518 1060 1526
rect 1031 1486 1044 1505
rect 1059 1486 1089 1502
rect 1031 1470 1105 1486
rect 1031 1468 1044 1470
rect 1059 1468 1093 1470
rect 696 1446 709 1448
rect 724 1446 758 1448
rect 696 1430 758 1446
rect 802 1441 818 1444
rect 880 1441 910 1452
rect 958 1448 1004 1464
rect 1031 1452 1105 1468
rect 958 1446 992 1448
rect 957 1430 1004 1446
rect 1031 1430 1044 1452
rect 1059 1430 1089 1452
rect 1116 1430 1117 1446
rect 1132 1430 1145 1590
rect 1175 1486 1188 1590
rect 1233 1568 1234 1578
rect 1249 1568 1262 1578
rect 1233 1564 1262 1568
rect 1267 1564 1297 1590
rect 1315 1576 1331 1578
rect 1403 1576 1456 1590
rect 1404 1574 1468 1576
rect 1511 1574 1526 1590
rect 1575 1587 1605 1590
rect 1575 1584 1611 1587
rect 1541 1576 1557 1578
rect 1315 1564 1330 1568
rect 1233 1562 1330 1564
rect 1358 1562 1526 1574
rect 1542 1564 1557 1568
rect 1575 1565 1614 1584
rect 1633 1578 1640 1579
rect 1639 1571 1640 1578
rect 1623 1568 1624 1571
rect 1639 1568 1652 1571
rect 1575 1564 1605 1565
rect 1614 1564 1620 1565
rect 1623 1564 1652 1568
rect 1542 1563 1652 1564
rect 1542 1562 1658 1563
rect 1217 1554 1268 1562
rect 1217 1542 1242 1554
rect 1249 1542 1268 1554
rect 1299 1554 1349 1562
rect 1299 1546 1315 1554
rect 1322 1552 1349 1554
rect 1358 1552 1579 1562
rect 1322 1542 1579 1552
rect 1608 1554 1658 1562
rect 1608 1545 1624 1554
rect 1217 1534 1268 1542
rect 1315 1534 1579 1542
rect 1605 1542 1624 1545
rect 1631 1542 1658 1554
rect 1605 1534 1658 1542
rect 1233 1526 1234 1534
rect 1249 1526 1262 1534
rect 1233 1518 1249 1526
rect 1230 1511 1249 1514
rect 1230 1502 1252 1511
rect 1203 1492 1252 1502
rect 1203 1486 1233 1492
rect 1252 1487 1257 1492
rect 1175 1470 1249 1486
rect 1267 1478 1297 1534
rect 1332 1524 1540 1534
rect 1575 1530 1620 1534
rect 1623 1533 1624 1534
rect 1639 1533 1652 1534
rect 1358 1494 1547 1524
rect 1373 1491 1547 1494
rect 1366 1488 1547 1491
rect 1175 1468 1188 1470
rect 1203 1468 1237 1470
rect 1175 1452 1249 1468
rect 1276 1464 1289 1478
rect 1304 1464 1320 1480
rect 1366 1475 1377 1488
rect 1159 1430 1160 1446
rect 1175 1430 1188 1452
rect 1203 1430 1233 1452
rect 1276 1448 1338 1464
rect 1366 1457 1377 1473
rect 1382 1468 1392 1488
rect 1402 1468 1416 1488
rect 1419 1475 1428 1488
rect 1444 1475 1453 1488
rect 1382 1457 1416 1468
rect 1419 1457 1428 1473
rect 1444 1457 1453 1473
rect 1460 1468 1470 1488
rect 1480 1468 1494 1488
rect 1495 1475 1506 1488
rect 1460 1457 1494 1468
rect 1495 1457 1506 1473
rect 1552 1464 1568 1480
rect 1575 1478 1605 1530
rect 1639 1526 1640 1533
rect 1624 1518 1640 1526
rect 1611 1486 1624 1505
rect 1639 1486 1669 1502
rect 1611 1470 1685 1486
rect 1611 1468 1624 1470
rect 1639 1468 1673 1470
rect 1276 1446 1289 1448
rect 1304 1446 1338 1448
rect 1276 1430 1338 1446
rect 1382 1441 1398 1444
rect 1460 1441 1490 1452
rect 1538 1448 1584 1464
rect 1611 1452 1685 1468
rect 1538 1446 1572 1448
rect 1537 1430 1584 1446
rect 1611 1430 1624 1452
rect 1639 1430 1669 1452
rect 1696 1430 1697 1446
rect 1712 1430 1725 1590
rect 1755 1486 1768 1590
rect 1813 1568 1814 1578
rect 1829 1568 1842 1578
rect 1813 1564 1842 1568
rect 1847 1564 1877 1590
rect 1895 1576 1911 1578
rect 1983 1576 2036 1590
rect 1984 1574 2048 1576
rect 2091 1574 2106 1590
rect 2155 1587 2185 1590
rect 2155 1584 2191 1587
rect 2121 1576 2137 1578
rect 1895 1564 1910 1568
rect 1813 1562 1910 1564
rect 1938 1562 2106 1574
rect 2122 1564 2137 1568
rect 2155 1565 2194 1584
rect 2213 1578 2220 1579
rect 2219 1571 2220 1578
rect 2203 1568 2204 1571
rect 2219 1568 2232 1571
rect 2155 1564 2185 1565
rect 2194 1564 2200 1565
rect 2203 1564 2232 1568
rect 2122 1563 2232 1564
rect 2122 1562 2238 1563
rect 1797 1554 1848 1562
rect 1797 1542 1822 1554
rect 1829 1542 1848 1554
rect 1879 1554 1929 1562
rect 1879 1546 1895 1554
rect 1902 1552 1929 1554
rect 1938 1552 2159 1562
rect 1902 1542 2159 1552
rect 2188 1554 2238 1562
rect 2188 1545 2204 1554
rect 1797 1534 1848 1542
rect 1895 1534 2159 1542
rect 2185 1542 2204 1545
rect 2211 1542 2238 1554
rect 2185 1534 2238 1542
rect 1813 1526 1814 1534
rect 1829 1526 1842 1534
rect 1813 1518 1829 1526
rect 1810 1511 1829 1514
rect 1810 1502 1832 1511
rect 1783 1492 1832 1502
rect 1783 1486 1813 1492
rect 1832 1487 1837 1492
rect 1755 1470 1829 1486
rect 1847 1478 1877 1534
rect 1912 1524 2120 1534
rect 2155 1530 2200 1534
rect 2203 1533 2204 1534
rect 2219 1533 2232 1534
rect 1938 1494 2127 1524
rect 1953 1491 2127 1494
rect 1946 1488 2127 1491
rect 1755 1468 1768 1470
rect 1783 1468 1817 1470
rect 1755 1452 1829 1468
rect 1856 1464 1869 1478
rect 1884 1464 1900 1480
rect 1946 1475 1957 1488
rect 1739 1430 1740 1446
rect 1755 1430 1768 1452
rect 1783 1430 1813 1452
rect 1856 1448 1918 1464
rect 1946 1457 1957 1473
rect 1962 1468 1972 1488
rect 1982 1468 1996 1488
rect 1999 1475 2008 1488
rect 2024 1475 2033 1488
rect 1962 1457 1996 1468
rect 1999 1457 2008 1473
rect 2024 1457 2033 1473
rect 2040 1468 2050 1488
rect 2060 1468 2074 1488
rect 2075 1475 2086 1488
rect 2040 1457 2074 1468
rect 2075 1457 2086 1473
rect 2132 1464 2148 1480
rect 2155 1478 2185 1530
rect 2219 1526 2220 1533
rect 2204 1518 2220 1526
rect 2191 1486 2204 1505
rect 2219 1486 2249 1502
rect 2191 1470 2265 1486
rect 2191 1468 2204 1470
rect 2219 1468 2253 1470
rect 1856 1446 1869 1448
rect 1884 1446 1918 1448
rect 1856 1430 1918 1446
rect 1962 1441 1978 1444
rect 2040 1441 2070 1452
rect 2118 1448 2164 1464
rect 2191 1452 2265 1468
rect 2118 1446 2152 1448
rect 2117 1430 2164 1446
rect 2191 1430 2204 1452
rect 2219 1430 2249 1452
rect 2276 1430 2277 1446
rect 2292 1430 2305 1590
rect 2335 1486 2348 1590
rect 2393 1568 2394 1578
rect 2409 1568 2422 1578
rect 2393 1564 2422 1568
rect 2427 1564 2457 1590
rect 2475 1576 2491 1578
rect 2563 1576 2616 1590
rect 2564 1574 2628 1576
rect 2671 1574 2686 1590
rect 2735 1587 2765 1590
rect 2735 1584 2771 1587
rect 2701 1576 2717 1578
rect 2475 1564 2490 1568
rect 2393 1562 2490 1564
rect 2518 1562 2686 1574
rect 2702 1564 2717 1568
rect 2735 1565 2774 1584
rect 2793 1578 2800 1579
rect 2799 1571 2800 1578
rect 2783 1568 2784 1571
rect 2799 1568 2812 1571
rect 2735 1564 2765 1565
rect 2774 1564 2780 1565
rect 2783 1564 2812 1568
rect 2702 1563 2812 1564
rect 2702 1562 2818 1563
rect 2377 1554 2428 1562
rect 2377 1542 2402 1554
rect 2409 1542 2428 1554
rect 2459 1554 2509 1562
rect 2459 1546 2475 1554
rect 2482 1552 2509 1554
rect 2518 1552 2739 1562
rect 2482 1542 2739 1552
rect 2768 1554 2818 1562
rect 2768 1545 2784 1554
rect 2377 1534 2428 1542
rect 2475 1534 2739 1542
rect 2765 1542 2784 1545
rect 2791 1542 2818 1554
rect 2765 1534 2818 1542
rect 2393 1526 2394 1534
rect 2409 1526 2422 1534
rect 2393 1518 2409 1526
rect 2390 1511 2409 1514
rect 2390 1502 2412 1511
rect 2363 1492 2412 1502
rect 2363 1486 2393 1492
rect 2412 1487 2417 1492
rect 2335 1470 2409 1486
rect 2427 1478 2457 1534
rect 2492 1524 2700 1534
rect 2735 1530 2780 1534
rect 2783 1533 2784 1534
rect 2799 1533 2812 1534
rect 2518 1494 2707 1524
rect 2533 1491 2707 1494
rect 2526 1488 2707 1491
rect 2335 1468 2348 1470
rect 2363 1468 2397 1470
rect 2335 1452 2409 1468
rect 2436 1464 2449 1478
rect 2464 1464 2480 1480
rect 2526 1475 2537 1488
rect 2319 1430 2320 1446
rect 2335 1430 2348 1452
rect 2363 1430 2393 1452
rect 2436 1448 2498 1464
rect 2526 1457 2537 1473
rect 2542 1468 2552 1488
rect 2562 1468 2576 1488
rect 2579 1475 2588 1488
rect 2604 1475 2613 1488
rect 2542 1457 2576 1468
rect 2579 1457 2588 1473
rect 2604 1457 2613 1473
rect 2620 1468 2630 1488
rect 2640 1468 2654 1488
rect 2655 1475 2666 1488
rect 2620 1457 2654 1468
rect 2655 1457 2666 1473
rect 2712 1464 2728 1480
rect 2735 1478 2765 1530
rect 2799 1526 2800 1533
rect 2784 1518 2800 1526
rect 2771 1486 2784 1505
rect 2799 1486 2829 1502
rect 2771 1470 2845 1486
rect 2771 1468 2784 1470
rect 2799 1468 2833 1470
rect 2436 1446 2449 1448
rect 2464 1446 2498 1448
rect 2436 1430 2498 1446
rect 2542 1441 2558 1444
rect 2620 1441 2650 1452
rect 2698 1448 2744 1464
rect 2771 1452 2845 1468
rect 2698 1446 2732 1448
rect 2697 1430 2744 1446
rect 2771 1430 2784 1452
rect 2799 1430 2829 1452
rect 2856 1430 2857 1446
rect 2872 1430 2885 1590
rect 2915 1486 2928 1590
rect 2973 1568 2974 1578
rect 2989 1568 3002 1578
rect 2973 1564 3002 1568
rect 3007 1564 3037 1590
rect 3055 1576 3071 1578
rect 3143 1576 3196 1590
rect 3144 1574 3208 1576
rect 3251 1574 3266 1590
rect 3315 1587 3345 1590
rect 3315 1584 3351 1587
rect 3281 1576 3297 1578
rect 3055 1564 3070 1568
rect 2973 1562 3070 1564
rect 3098 1562 3266 1574
rect 3282 1564 3297 1568
rect 3315 1565 3354 1584
rect 3373 1578 3380 1579
rect 3379 1571 3380 1578
rect 3363 1568 3364 1571
rect 3379 1568 3392 1571
rect 3315 1564 3345 1565
rect 3354 1564 3360 1565
rect 3363 1564 3392 1568
rect 3282 1563 3392 1564
rect 3282 1562 3398 1563
rect 2957 1554 3008 1562
rect 2957 1542 2982 1554
rect 2989 1542 3008 1554
rect 3039 1554 3089 1562
rect 3039 1546 3055 1554
rect 3062 1552 3089 1554
rect 3098 1552 3319 1562
rect 3062 1542 3319 1552
rect 3348 1554 3398 1562
rect 3348 1545 3364 1554
rect 2957 1534 3008 1542
rect 3055 1534 3319 1542
rect 3345 1542 3364 1545
rect 3371 1542 3398 1554
rect 3345 1534 3398 1542
rect 2973 1526 2974 1534
rect 2989 1526 3002 1534
rect 2973 1518 2989 1526
rect 2970 1511 2989 1514
rect 2970 1502 2992 1511
rect 2943 1492 2992 1502
rect 2943 1486 2973 1492
rect 2992 1487 2997 1492
rect 2915 1470 2989 1486
rect 3007 1478 3037 1534
rect 3072 1524 3280 1534
rect 3315 1530 3360 1534
rect 3363 1533 3364 1534
rect 3379 1533 3392 1534
rect 3098 1494 3287 1524
rect 3113 1491 3287 1494
rect 3106 1488 3287 1491
rect 2915 1468 2928 1470
rect 2943 1468 2977 1470
rect 2915 1452 2989 1468
rect 3016 1464 3029 1478
rect 3044 1464 3060 1480
rect 3106 1475 3117 1488
rect 2899 1430 2900 1446
rect 2915 1430 2928 1452
rect 2943 1430 2973 1452
rect 3016 1448 3078 1464
rect 3106 1457 3117 1473
rect 3122 1468 3132 1488
rect 3142 1468 3156 1488
rect 3159 1475 3168 1488
rect 3184 1475 3193 1488
rect 3122 1457 3156 1468
rect 3159 1457 3168 1473
rect 3184 1457 3193 1473
rect 3200 1468 3210 1488
rect 3220 1468 3234 1488
rect 3235 1475 3246 1488
rect 3200 1457 3234 1468
rect 3235 1457 3246 1473
rect 3292 1464 3308 1480
rect 3315 1478 3345 1530
rect 3379 1526 3380 1533
rect 3364 1518 3380 1526
rect 3351 1486 3364 1505
rect 3379 1486 3409 1502
rect 3351 1470 3425 1486
rect 3351 1468 3364 1470
rect 3379 1468 3413 1470
rect 3016 1446 3029 1448
rect 3044 1446 3078 1448
rect 3016 1430 3078 1446
rect 3122 1441 3138 1444
rect 3200 1441 3230 1452
rect 3278 1448 3324 1464
rect 3351 1452 3425 1468
rect 3278 1446 3312 1448
rect 3277 1430 3324 1446
rect 3351 1430 3364 1452
rect 3379 1430 3409 1452
rect 3436 1430 3437 1446
rect 3452 1430 3465 1590
rect 3495 1486 3508 1590
rect 3553 1568 3554 1578
rect 3569 1568 3582 1578
rect 3553 1564 3582 1568
rect 3587 1564 3617 1590
rect 3635 1576 3651 1578
rect 3723 1576 3776 1590
rect 3724 1574 3788 1576
rect 3831 1574 3846 1590
rect 3895 1587 3925 1590
rect 3895 1584 3931 1587
rect 3861 1576 3877 1578
rect 3635 1564 3650 1568
rect 3553 1562 3650 1564
rect 3678 1562 3846 1574
rect 3862 1564 3877 1568
rect 3895 1565 3934 1584
rect 3953 1578 3960 1579
rect 3959 1571 3960 1578
rect 3943 1568 3944 1571
rect 3959 1568 3972 1571
rect 3895 1564 3925 1565
rect 3934 1564 3940 1565
rect 3943 1564 3972 1568
rect 3862 1563 3972 1564
rect 3862 1562 3978 1563
rect 3537 1554 3588 1562
rect 3537 1542 3562 1554
rect 3569 1542 3588 1554
rect 3619 1554 3669 1562
rect 3619 1546 3635 1554
rect 3642 1552 3669 1554
rect 3678 1552 3899 1562
rect 3642 1542 3899 1552
rect 3928 1554 3978 1562
rect 3928 1545 3944 1554
rect 3537 1534 3588 1542
rect 3635 1534 3899 1542
rect 3925 1542 3944 1545
rect 3951 1542 3978 1554
rect 3925 1534 3978 1542
rect 3553 1526 3554 1534
rect 3569 1526 3582 1534
rect 3553 1518 3569 1526
rect 3550 1511 3569 1514
rect 3550 1502 3572 1511
rect 3523 1492 3572 1502
rect 3523 1486 3553 1492
rect 3572 1487 3577 1492
rect 3495 1470 3569 1486
rect 3587 1478 3617 1534
rect 3652 1524 3860 1534
rect 3895 1530 3940 1534
rect 3943 1533 3944 1534
rect 3959 1533 3972 1534
rect 3678 1494 3867 1524
rect 3693 1491 3867 1494
rect 3686 1488 3867 1491
rect 3495 1468 3508 1470
rect 3523 1468 3557 1470
rect 3495 1452 3569 1468
rect 3596 1464 3609 1478
rect 3624 1464 3640 1480
rect 3686 1475 3697 1488
rect 3479 1430 3480 1446
rect 3495 1430 3508 1452
rect 3523 1430 3553 1452
rect 3596 1448 3658 1464
rect 3686 1457 3697 1473
rect 3702 1468 3712 1488
rect 3722 1468 3736 1488
rect 3739 1475 3748 1488
rect 3764 1475 3773 1488
rect 3702 1457 3736 1468
rect 3739 1457 3748 1473
rect 3764 1457 3773 1473
rect 3780 1468 3790 1488
rect 3800 1468 3814 1488
rect 3815 1475 3826 1488
rect 3780 1457 3814 1468
rect 3815 1457 3826 1473
rect 3872 1464 3888 1480
rect 3895 1478 3925 1530
rect 3959 1526 3960 1533
rect 3944 1518 3960 1526
rect 3931 1486 3944 1505
rect 3959 1486 3989 1502
rect 3931 1470 4005 1486
rect 3931 1468 3944 1470
rect 3959 1468 3993 1470
rect 3596 1446 3609 1448
rect 3624 1446 3658 1448
rect 3596 1430 3658 1446
rect 3702 1441 3718 1444
rect 3780 1441 3810 1452
rect 3858 1448 3904 1464
rect 3931 1452 4005 1468
rect 3858 1446 3892 1448
rect 3857 1430 3904 1446
rect 3931 1430 3944 1452
rect 3959 1430 3989 1452
rect 4016 1430 4017 1446
rect 4032 1430 4045 1590
rect 4075 1486 4088 1590
rect 4133 1568 4134 1578
rect 4149 1568 4162 1578
rect 4133 1564 4162 1568
rect 4167 1564 4197 1590
rect 4215 1576 4231 1578
rect 4303 1576 4356 1590
rect 4304 1574 4368 1576
rect 4411 1574 4426 1590
rect 4475 1587 4505 1590
rect 4475 1584 4511 1587
rect 4441 1576 4457 1578
rect 4215 1564 4230 1568
rect 4133 1562 4230 1564
rect 4258 1562 4426 1574
rect 4442 1564 4457 1568
rect 4475 1565 4514 1584
rect 4533 1578 4540 1579
rect 4539 1571 4540 1578
rect 4523 1568 4524 1571
rect 4539 1568 4552 1571
rect 4475 1564 4505 1565
rect 4514 1564 4520 1565
rect 4523 1564 4552 1568
rect 4442 1563 4552 1564
rect 4442 1562 4558 1563
rect 4117 1554 4168 1562
rect 4117 1542 4142 1554
rect 4149 1542 4168 1554
rect 4199 1554 4249 1562
rect 4199 1546 4215 1554
rect 4222 1552 4249 1554
rect 4258 1552 4479 1562
rect 4222 1542 4479 1552
rect 4508 1554 4558 1562
rect 4508 1545 4524 1554
rect 4117 1534 4168 1542
rect 4215 1534 4479 1542
rect 4505 1542 4524 1545
rect 4531 1542 4558 1554
rect 4505 1534 4558 1542
rect 4133 1526 4134 1534
rect 4149 1526 4162 1534
rect 4133 1518 4149 1526
rect 4130 1511 4149 1514
rect 4130 1502 4152 1511
rect 4103 1492 4152 1502
rect 4103 1486 4133 1492
rect 4152 1487 4157 1492
rect 4075 1470 4149 1486
rect 4167 1478 4197 1534
rect 4232 1524 4440 1534
rect 4475 1530 4520 1534
rect 4523 1533 4524 1534
rect 4539 1533 4552 1534
rect 4258 1494 4447 1524
rect 4273 1491 4447 1494
rect 4266 1488 4447 1491
rect 4075 1468 4088 1470
rect 4103 1468 4137 1470
rect 4075 1452 4149 1468
rect 4176 1464 4189 1478
rect 4204 1464 4220 1480
rect 4266 1475 4277 1488
rect 4059 1430 4060 1446
rect 4075 1430 4088 1452
rect 4103 1430 4133 1452
rect 4176 1448 4238 1464
rect 4266 1457 4277 1473
rect 4282 1468 4292 1488
rect 4302 1468 4316 1488
rect 4319 1475 4328 1488
rect 4344 1475 4353 1488
rect 4282 1457 4316 1468
rect 4319 1457 4328 1473
rect 4344 1457 4353 1473
rect 4360 1468 4370 1488
rect 4380 1468 4394 1488
rect 4395 1475 4406 1488
rect 4360 1457 4394 1468
rect 4395 1457 4406 1473
rect 4452 1464 4468 1480
rect 4475 1478 4505 1530
rect 4539 1526 4540 1533
rect 4524 1518 4540 1526
rect 4511 1486 4524 1505
rect 4539 1486 4569 1502
rect 4511 1470 4585 1486
rect 4511 1468 4524 1470
rect 4539 1468 4573 1470
rect 4176 1446 4189 1448
rect 4204 1446 4238 1448
rect 4176 1430 4238 1446
rect 4282 1441 4298 1444
rect 4360 1441 4390 1452
rect 4438 1448 4484 1464
rect 4511 1452 4585 1468
rect 4438 1446 4472 1448
rect 4437 1430 4484 1446
rect 4511 1430 4524 1452
rect 4539 1430 4569 1452
rect 4596 1430 4597 1446
rect 4612 1430 4625 1590
rect -7 1422 34 1430
rect -7 1396 8 1422
rect 15 1396 34 1422
rect 98 1418 160 1430
rect 172 1418 247 1430
rect 305 1418 380 1430
rect 392 1418 423 1430
rect 429 1418 464 1430
rect 98 1416 260 1418
rect -7 1388 34 1396
rect 116 1392 129 1416
rect 144 1414 159 1416
rect -1 1378 0 1388
rect 15 1378 28 1388
rect 43 1378 73 1392
rect 116 1378 159 1392
rect 183 1389 190 1396
rect 193 1392 260 1416
rect 292 1416 464 1418
rect 262 1394 290 1398
rect 292 1394 372 1416
rect 393 1414 408 1416
rect 262 1392 372 1394
rect 193 1388 372 1392
rect 166 1378 196 1388
rect 198 1378 351 1388
rect 359 1378 389 1388
rect 393 1378 423 1392
rect 451 1378 464 1416
rect 536 1422 571 1430
rect 536 1396 537 1422
rect 544 1396 571 1422
rect 479 1378 509 1392
rect 536 1388 571 1396
rect 573 1422 614 1430
rect 573 1396 588 1422
rect 595 1396 614 1422
rect 678 1418 740 1430
rect 752 1418 827 1430
rect 885 1418 960 1430
rect 972 1418 1003 1430
rect 1009 1418 1044 1430
rect 678 1416 840 1418
rect 573 1388 614 1396
rect 696 1392 709 1416
rect 724 1414 739 1416
rect 536 1378 537 1388
rect 552 1378 565 1388
rect 579 1378 580 1388
rect 595 1378 608 1388
rect 623 1378 653 1392
rect 696 1378 739 1392
rect 763 1389 770 1396
rect 773 1392 840 1416
rect 872 1416 1044 1418
rect 842 1394 870 1398
rect 872 1394 952 1416
rect 973 1414 988 1416
rect 842 1392 952 1394
rect 773 1388 952 1392
rect 746 1378 776 1388
rect 778 1378 931 1388
rect 939 1378 969 1388
rect 973 1378 1003 1392
rect 1031 1378 1044 1416
rect 1116 1422 1151 1430
rect 1116 1396 1117 1422
rect 1124 1396 1151 1422
rect 1059 1378 1089 1392
rect 1116 1388 1151 1396
rect 1153 1422 1194 1430
rect 1153 1396 1168 1422
rect 1175 1396 1194 1422
rect 1258 1418 1320 1430
rect 1332 1418 1407 1430
rect 1465 1418 1540 1430
rect 1552 1418 1583 1430
rect 1589 1418 1624 1430
rect 1258 1416 1420 1418
rect 1153 1388 1194 1396
rect 1276 1392 1289 1416
rect 1304 1414 1319 1416
rect 1116 1378 1117 1388
rect 1132 1378 1145 1388
rect 1159 1378 1160 1388
rect 1175 1378 1188 1388
rect 1203 1378 1233 1392
rect 1276 1378 1319 1392
rect 1343 1389 1350 1396
rect 1353 1392 1420 1416
rect 1452 1416 1624 1418
rect 1422 1394 1450 1398
rect 1452 1394 1532 1416
rect 1553 1414 1568 1416
rect 1422 1392 1532 1394
rect 1353 1388 1532 1392
rect 1326 1378 1356 1388
rect 1358 1378 1511 1388
rect 1519 1378 1549 1388
rect 1553 1378 1583 1392
rect 1611 1378 1624 1416
rect 1696 1422 1731 1430
rect 1696 1396 1697 1422
rect 1704 1396 1731 1422
rect 1639 1378 1669 1392
rect 1696 1388 1731 1396
rect 1733 1422 1774 1430
rect 1733 1396 1748 1422
rect 1755 1396 1774 1422
rect 1838 1418 1900 1430
rect 1912 1418 1987 1430
rect 2045 1418 2120 1430
rect 2132 1418 2163 1430
rect 2169 1418 2204 1430
rect 1838 1416 2000 1418
rect 1733 1388 1774 1396
rect 1856 1392 1869 1416
rect 1884 1414 1899 1416
rect 1696 1378 1697 1388
rect 1712 1378 1725 1388
rect 1739 1378 1740 1388
rect 1755 1378 1768 1388
rect 1783 1378 1813 1392
rect 1856 1378 1899 1392
rect 1923 1389 1930 1396
rect 1933 1392 2000 1416
rect 2032 1416 2204 1418
rect 2002 1394 2030 1398
rect 2032 1394 2112 1416
rect 2133 1414 2148 1416
rect 2002 1392 2112 1394
rect 1933 1388 2112 1392
rect 1906 1378 1936 1388
rect 1938 1378 2091 1388
rect 2099 1378 2129 1388
rect 2133 1378 2163 1392
rect 2191 1378 2204 1416
rect 2276 1422 2311 1430
rect 2276 1396 2277 1422
rect 2284 1396 2311 1422
rect 2219 1378 2249 1392
rect 2276 1388 2311 1396
rect 2313 1422 2354 1430
rect 2313 1396 2328 1422
rect 2335 1396 2354 1422
rect 2418 1418 2480 1430
rect 2492 1418 2567 1430
rect 2625 1418 2700 1430
rect 2712 1418 2743 1430
rect 2749 1418 2784 1430
rect 2418 1416 2580 1418
rect 2313 1388 2354 1396
rect 2436 1392 2449 1416
rect 2464 1414 2479 1416
rect 2276 1378 2277 1388
rect 2292 1378 2305 1388
rect 2319 1378 2320 1388
rect 2335 1378 2348 1388
rect 2363 1378 2393 1392
rect 2436 1378 2479 1392
rect 2503 1389 2510 1396
rect 2513 1392 2580 1416
rect 2612 1416 2784 1418
rect 2582 1394 2610 1398
rect 2612 1394 2692 1416
rect 2713 1414 2728 1416
rect 2582 1392 2692 1394
rect 2513 1388 2692 1392
rect 2486 1378 2516 1388
rect 2518 1378 2671 1388
rect 2679 1378 2709 1388
rect 2713 1378 2743 1392
rect 2771 1378 2784 1416
rect 2856 1422 2891 1430
rect 2856 1396 2857 1422
rect 2864 1396 2891 1422
rect 2799 1378 2829 1392
rect 2856 1388 2891 1396
rect 2893 1422 2934 1430
rect 2893 1396 2908 1422
rect 2915 1396 2934 1422
rect 2998 1418 3060 1430
rect 3072 1418 3147 1430
rect 3205 1418 3280 1430
rect 3292 1418 3323 1430
rect 3329 1418 3364 1430
rect 2998 1416 3160 1418
rect 2893 1388 2934 1396
rect 3016 1392 3029 1416
rect 3044 1414 3059 1416
rect 2856 1378 2857 1388
rect 2872 1378 2885 1388
rect 2899 1378 2900 1388
rect 2915 1378 2928 1388
rect 2943 1378 2973 1392
rect 3016 1378 3059 1392
rect 3083 1389 3090 1396
rect 3093 1392 3160 1416
rect 3192 1416 3364 1418
rect 3162 1394 3190 1398
rect 3192 1394 3272 1416
rect 3293 1414 3308 1416
rect 3162 1392 3272 1394
rect 3093 1388 3272 1392
rect 3066 1378 3096 1388
rect 3098 1378 3251 1388
rect 3259 1378 3289 1388
rect 3293 1378 3323 1392
rect 3351 1378 3364 1416
rect 3436 1422 3471 1430
rect 3436 1396 3437 1422
rect 3444 1396 3471 1422
rect 3379 1378 3409 1392
rect 3436 1388 3471 1396
rect 3473 1422 3514 1430
rect 3473 1396 3488 1422
rect 3495 1396 3514 1422
rect 3578 1418 3640 1430
rect 3652 1418 3727 1430
rect 3785 1418 3860 1430
rect 3872 1418 3903 1430
rect 3909 1418 3944 1430
rect 3578 1416 3740 1418
rect 3473 1388 3514 1396
rect 3596 1392 3609 1416
rect 3624 1414 3639 1416
rect 3436 1378 3437 1388
rect 3452 1378 3465 1388
rect 3479 1378 3480 1388
rect 3495 1378 3508 1388
rect 3523 1378 3553 1392
rect 3596 1378 3639 1392
rect 3663 1389 3670 1396
rect 3673 1392 3740 1416
rect 3772 1416 3944 1418
rect 3742 1394 3770 1398
rect 3772 1394 3852 1416
rect 3873 1414 3888 1416
rect 3742 1392 3852 1394
rect 3673 1388 3852 1392
rect 3646 1378 3676 1388
rect 3678 1378 3831 1388
rect 3839 1378 3869 1388
rect 3873 1378 3903 1392
rect 3931 1378 3944 1416
rect 4016 1422 4051 1430
rect 4016 1396 4017 1422
rect 4024 1396 4051 1422
rect 3959 1378 3989 1392
rect 4016 1388 4051 1396
rect 4053 1422 4094 1430
rect 4053 1396 4068 1422
rect 4075 1396 4094 1422
rect 4158 1418 4220 1430
rect 4232 1418 4307 1430
rect 4365 1418 4440 1430
rect 4452 1418 4483 1430
rect 4489 1418 4524 1430
rect 4158 1416 4320 1418
rect 4053 1388 4094 1396
rect 4176 1392 4189 1416
rect 4204 1414 4219 1416
rect 4016 1378 4017 1388
rect 4032 1378 4045 1388
rect 4059 1378 4060 1388
rect 4075 1378 4088 1388
rect 4103 1378 4133 1392
rect 4176 1378 4219 1392
rect 4243 1389 4250 1396
rect 4253 1392 4320 1416
rect 4352 1416 4524 1418
rect 4322 1394 4350 1398
rect 4352 1394 4432 1416
rect 4453 1414 4468 1416
rect 4322 1392 4432 1394
rect 4253 1388 4432 1392
rect 4226 1378 4256 1388
rect 4258 1378 4411 1388
rect 4419 1378 4449 1388
rect 4453 1378 4483 1392
rect 4511 1378 4524 1416
rect 4596 1422 4631 1430
rect 4596 1396 4597 1422
rect 4604 1396 4631 1422
rect 4539 1378 4569 1392
rect 4596 1388 4631 1396
rect 4596 1378 4597 1388
rect 4612 1378 4625 1388
rect -1 1372 4625 1378
rect 0 1364 4625 1372
rect 15 1334 28 1364
rect 43 1346 73 1364
rect 116 1350 130 1364
rect 166 1350 386 1364
rect 117 1348 130 1350
rect 83 1336 98 1348
rect 80 1334 102 1336
rect 107 1334 137 1348
rect 198 1346 351 1350
rect 180 1334 372 1346
rect 415 1334 445 1348
rect 451 1334 464 1364
rect 479 1346 509 1364
rect 552 1334 565 1364
rect 595 1334 608 1364
rect 623 1346 653 1364
rect 696 1350 710 1364
rect 746 1350 966 1364
rect 697 1348 710 1350
rect 663 1336 678 1348
rect 660 1334 682 1336
rect 687 1334 717 1348
rect 778 1346 931 1350
rect 760 1334 952 1346
rect 995 1334 1025 1348
rect 1031 1334 1044 1364
rect 1059 1346 1089 1364
rect 1132 1334 1145 1364
rect 1175 1334 1188 1364
rect 1203 1346 1233 1364
rect 1276 1350 1290 1364
rect 1326 1350 1546 1364
rect 1277 1348 1290 1350
rect 1243 1336 1258 1348
rect 1240 1334 1262 1336
rect 1267 1334 1297 1348
rect 1358 1346 1511 1350
rect 1340 1334 1532 1346
rect 1575 1334 1605 1348
rect 1611 1334 1624 1364
rect 1639 1346 1669 1364
rect 1712 1334 1725 1364
rect 1755 1334 1768 1364
rect 1783 1346 1813 1364
rect 1856 1350 1870 1364
rect 1906 1350 2126 1364
rect 1857 1348 1870 1350
rect 1823 1336 1838 1348
rect 1820 1334 1842 1336
rect 1847 1334 1877 1348
rect 1938 1346 2091 1350
rect 1920 1334 2112 1346
rect 2155 1334 2185 1348
rect 2191 1334 2204 1364
rect 2219 1346 2249 1364
rect 2292 1334 2305 1364
rect 2335 1334 2348 1364
rect 2363 1346 2393 1364
rect 2436 1350 2450 1364
rect 2486 1350 2706 1364
rect 2437 1348 2450 1350
rect 2403 1336 2418 1348
rect 2400 1334 2422 1336
rect 2427 1334 2457 1348
rect 2518 1346 2671 1350
rect 2500 1334 2692 1346
rect 2735 1334 2765 1348
rect 2771 1334 2784 1364
rect 2799 1346 2829 1364
rect 2872 1334 2885 1364
rect 2915 1334 2928 1364
rect 2943 1346 2973 1364
rect 3016 1350 3030 1364
rect 3066 1350 3286 1364
rect 3017 1348 3030 1350
rect 2983 1336 2998 1348
rect 2980 1334 3002 1336
rect 3007 1334 3037 1348
rect 3098 1346 3251 1350
rect 3080 1334 3272 1346
rect 3315 1334 3345 1348
rect 3351 1334 3364 1364
rect 3379 1346 3409 1364
rect 3452 1334 3465 1364
rect 3495 1334 3508 1364
rect 3523 1346 3553 1364
rect 3596 1350 3610 1364
rect 3646 1350 3866 1364
rect 3597 1348 3610 1350
rect 3563 1336 3578 1348
rect 3560 1334 3582 1336
rect 3587 1334 3617 1348
rect 3678 1346 3831 1350
rect 3660 1334 3852 1346
rect 3895 1334 3925 1348
rect 3931 1334 3944 1364
rect 3959 1346 3989 1364
rect 4032 1334 4045 1364
rect 4075 1334 4088 1364
rect 4103 1346 4133 1364
rect 4176 1350 4190 1364
rect 4226 1350 4446 1364
rect 4177 1348 4190 1350
rect 4143 1336 4158 1348
rect 4140 1334 4162 1336
rect 4167 1334 4197 1348
rect 4258 1346 4411 1350
rect 4240 1334 4432 1346
rect 4475 1334 4505 1348
rect 4511 1334 4524 1364
rect 4539 1346 4569 1364
rect 4612 1334 4625 1364
rect 0 1320 4625 1334
rect 15 1216 28 1320
rect 73 1298 74 1308
rect 89 1298 102 1308
rect 73 1294 102 1298
rect 107 1294 137 1320
rect 155 1306 171 1308
rect 243 1306 296 1320
rect 244 1304 308 1306
rect 351 1304 366 1320
rect 415 1317 445 1320
rect 415 1314 451 1317
rect 381 1306 397 1308
rect 155 1294 170 1298
rect 73 1292 170 1294
rect 198 1292 366 1304
rect 382 1294 397 1298
rect 415 1295 454 1314
rect 473 1308 480 1309
rect 479 1301 480 1308
rect 463 1298 464 1301
rect 479 1298 492 1301
rect 415 1294 445 1295
rect 454 1294 460 1295
rect 463 1294 492 1298
rect 382 1293 492 1294
rect 382 1292 498 1293
rect 57 1284 108 1292
rect 57 1272 82 1284
rect 89 1272 108 1284
rect 139 1284 189 1292
rect 139 1276 155 1284
rect 162 1282 189 1284
rect 198 1282 419 1292
rect 162 1272 419 1282
rect 448 1284 498 1292
rect 448 1275 464 1284
rect 57 1264 108 1272
rect 155 1264 419 1272
rect 445 1272 464 1275
rect 471 1272 498 1284
rect 445 1264 498 1272
rect 73 1256 74 1264
rect 89 1256 102 1264
rect 73 1248 89 1256
rect 70 1241 89 1244
rect 70 1232 92 1241
rect 43 1222 92 1232
rect 43 1216 73 1222
rect 92 1217 97 1222
rect 15 1200 89 1216
rect 107 1208 137 1264
rect 172 1254 380 1264
rect 415 1260 460 1264
rect 463 1263 464 1264
rect 479 1263 492 1264
rect 198 1224 387 1254
rect 213 1221 387 1224
rect 206 1218 387 1221
rect 15 1198 28 1200
rect 43 1198 77 1200
rect 15 1182 89 1198
rect 116 1194 129 1208
rect 144 1194 160 1210
rect 206 1205 217 1218
rect -1 1160 0 1176
rect 15 1160 28 1182
rect 43 1160 73 1182
rect 116 1178 178 1194
rect 206 1187 217 1203
rect 222 1198 232 1218
rect 242 1198 256 1218
rect 259 1205 268 1218
rect 284 1205 293 1218
rect 222 1187 256 1198
rect 259 1187 268 1203
rect 284 1187 293 1203
rect 300 1198 310 1218
rect 320 1198 334 1218
rect 335 1205 346 1218
rect 300 1187 334 1198
rect 335 1187 346 1203
rect 392 1194 408 1210
rect 415 1208 445 1260
rect 479 1256 480 1263
rect 464 1248 480 1256
rect 451 1216 464 1235
rect 479 1216 509 1232
rect 451 1200 525 1216
rect 451 1198 464 1200
rect 479 1198 513 1200
rect 116 1176 129 1178
rect 144 1176 178 1178
rect 116 1160 178 1176
rect 222 1171 238 1174
rect 300 1171 330 1182
rect 378 1178 424 1194
rect 451 1182 525 1198
rect 378 1176 412 1178
rect 377 1160 424 1176
rect 451 1160 464 1182
rect 479 1160 509 1182
rect 536 1160 537 1176
rect 552 1160 565 1320
rect 595 1216 608 1320
rect 653 1298 654 1308
rect 669 1298 682 1308
rect 653 1294 682 1298
rect 687 1294 717 1320
rect 735 1306 751 1308
rect 823 1306 876 1320
rect 824 1304 888 1306
rect 931 1304 946 1320
rect 995 1317 1025 1320
rect 995 1314 1031 1317
rect 961 1306 977 1308
rect 735 1294 750 1298
rect 653 1292 750 1294
rect 778 1292 946 1304
rect 962 1294 977 1298
rect 995 1295 1034 1314
rect 1053 1308 1060 1309
rect 1059 1301 1060 1308
rect 1043 1298 1044 1301
rect 1059 1298 1072 1301
rect 995 1294 1025 1295
rect 1034 1294 1040 1295
rect 1043 1294 1072 1298
rect 962 1293 1072 1294
rect 962 1292 1078 1293
rect 637 1284 688 1292
rect 637 1272 662 1284
rect 669 1272 688 1284
rect 719 1284 769 1292
rect 719 1276 735 1284
rect 742 1282 769 1284
rect 778 1282 999 1292
rect 742 1272 999 1282
rect 1028 1284 1078 1292
rect 1028 1275 1044 1284
rect 637 1264 688 1272
rect 735 1264 999 1272
rect 1025 1272 1044 1275
rect 1051 1272 1078 1284
rect 1025 1264 1078 1272
rect 653 1256 654 1264
rect 669 1256 682 1264
rect 653 1248 669 1256
rect 650 1241 669 1244
rect 650 1232 672 1241
rect 623 1222 672 1232
rect 623 1216 653 1222
rect 672 1217 677 1222
rect 595 1200 669 1216
rect 687 1208 717 1264
rect 752 1254 960 1264
rect 995 1260 1040 1264
rect 1043 1263 1044 1264
rect 1059 1263 1072 1264
rect 778 1224 967 1254
rect 793 1221 967 1224
rect 786 1218 967 1221
rect 595 1198 608 1200
rect 623 1198 657 1200
rect 595 1182 669 1198
rect 696 1194 709 1208
rect 724 1194 740 1210
rect 786 1205 797 1218
rect 579 1160 580 1176
rect 595 1160 608 1182
rect 623 1160 653 1182
rect 696 1178 758 1194
rect 786 1187 797 1203
rect 802 1198 812 1218
rect 822 1198 836 1218
rect 839 1205 848 1218
rect 864 1205 873 1218
rect 802 1187 836 1198
rect 839 1187 848 1203
rect 864 1187 873 1203
rect 880 1198 890 1218
rect 900 1198 914 1218
rect 915 1205 926 1218
rect 880 1187 914 1198
rect 915 1187 926 1203
rect 972 1194 988 1210
rect 995 1208 1025 1260
rect 1059 1256 1060 1263
rect 1044 1248 1060 1256
rect 1031 1216 1044 1235
rect 1059 1216 1089 1232
rect 1031 1200 1105 1216
rect 1031 1198 1044 1200
rect 1059 1198 1093 1200
rect 696 1176 709 1178
rect 724 1176 758 1178
rect 696 1160 758 1176
rect 802 1171 818 1174
rect 880 1171 910 1182
rect 958 1178 1004 1194
rect 1031 1182 1105 1198
rect 958 1176 992 1178
rect 957 1160 1004 1176
rect 1031 1160 1044 1182
rect 1059 1160 1089 1182
rect 1116 1160 1117 1176
rect 1132 1160 1145 1320
rect 1175 1216 1188 1320
rect 1233 1298 1234 1308
rect 1249 1298 1262 1308
rect 1233 1294 1262 1298
rect 1267 1294 1297 1320
rect 1315 1306 1331 1308
rect 1403 1306 1456 1320
rect 1404 1304 1468 1306
rect 1511 1304 1526 1320
rect 1575 1317 1605 1320
rect 1575 1314 1611 1317
rect 1541 1306 1557 1308
rect 1315 1294 1330 1298
rect 1233 1292 1330 1294
rect 1358 1292 1526 1304
rect 1542 1294 1557 1298
rect 1575 1295 1614 1314
rect 1633 1308 1640 1309
rect 1639 1301 1640 1308
rect 1623 1298 1624 1301
rect 1639 1298 1652 1301
rect 1575 1294 1605 1295
rect 1614 1294 1620 1295
rect 1623 1294 1652 1298
rect 1542 1293 1652 1294
rect 1542 1292 1658 1293
rect 1217 1284 1268 1292
rect 1217 1272 1242 1284
rect 1249 1272 1268 1284
rect 1299 1284 1349 1292
rect 1299 1276 1315 1284
rect 1322 1282 1349 1284
rect 1358 1282 1579 1292
rect 1322 1272 1579 1282
rect 1608 1284 1658 1292
rect 1608 1275 1624 1284
rect 1217 1264 1268 1272
rect 1315 1264 1579 1272
rect 1605 1272 1624 1275
rect 1631 1272 1658 1284
rect 1605 1264 1658 1272
rect 1233 1256 1234 1264
rect 1249 1256 1262 1264
rect 1233 1248 1249 1256
rect 1230 1241 1249 1244
rect 1230 1232 1252 1241
rect 1203 1222 1252 1232
rect 1203 1216 1233 1222
rect 1252 1217 1257 1222
rect 1175 1200 1249 1216
rect 1267 1208 1297 1264
rect 1332 1254 1540 1264
rect 1575 1260 1620 1264
rect 1623 1263 1624 1264
rect 1639 1263 1652 1264
rect 1358 1224 1547 1254
rect 1373 1221 1547 1224
rect 1366 1218 1547 1221
rect 1175 1198 1188 1200
rect 1203 1198 1237 1200
rect 1175 1182 1249 1198
rect 1276 1194 1289 1208
rect 1304 1194 1320 1210
rect 1366 1205 1377 1218
rect 1159 1160 1160 1176
rect 1175 1160 1188 1182
rect 1203 1160 1233 1182
rect 1276 1178 1338 1194
rect 1366 1187 1377 1203
rect 1382 1198 1392 1218
rect 1402 1198 1416 1218
rect 1419 1205 1428 1218
rect 1444 1205 1453 1218
rect 1382 1187 1416 1198
rect 1419 1187 1428 1203
rect 1444 1187 1453 1203
rect 1460 1198 1470 1218
rect 1480 1198 1494 1218
rect 1495 1205 1506 1218
rect 1460 1187 1494 1198
rect 1495 1187 1506 1203
rect 1552 1194 1568 1210
rect 1575 1208 1605 1260
rect 1639 1256 1640 1263
rect 1624 1248 1640 1256
rect 1611 1216 1624 1235
rect 1639 1216 1669 1232
rect 1611 1200 1685 1216
rect 1611 1198 1624 1200
rect 1639 1198 1673 1200
rect 1276 1176 1289 1178
rect 1304 1176 1338 1178
rect 1276 1160 1338 1176
rect 1382 1171 1398 1174
rect 1460 1171 1490 1182
rect 1538 1178 1584 1194
rect 1611 1182 1685 1198
rect 1538 1176 1572 1178
rect 1537 1160 1584 1176
rect 1611 1160 1624 1182
rect 1639 1160 1669 1182
rect 1696 1160 1697 1176
rect 1712 1160 1725 1320
rect 1755 1216 1768 1320
rect 1813 1298 1814 1308
rect 1829 1298 1842 1308
rect 1813 1294 1842 1298
rect 1847 1294 1877 1320
rect 1895 1306 1911 1308
rect 1983 1306 2036 1320
rect 1984 1304 2048 1306
rect 2091 1304 2106 1320
rect 2155 1317 2185 1320
rect 2155 1314 2191 1317
rect 2121 1306 2137 1308
rect 1895 1294 1910 1298
rect 1813 1292 1910 1294
rect 1938 1292 2106 1304
rect 2122 1294 2137 1298
rect 2155 1295 2194 1314
rect 2213 1308 2220 1309
rect 2219 1301 2220 1308
rect 2203 1298 2204 1301
rect 2219 1298 2232 1301
rect 2155 1294 2185 1295
rect 2194 1294 2200 1295
rect 2203 1294 2232 1298
rect 2122 1293 2232 1294
rect 2122 1292 2238 1293
rect 1797 1284 1848 1292
rect 1797 1272 1822 1284
rect 1829 1272 1848 1284
rect 1879 1284 1929 1292
rect 1879 1276 1895 1284
rect 1902 1282 1929 1284
rect 1938 1282 2159 1292
rect 1902 1272 2159 1282
rect 2188 1284 2238 1292
rect 2188 1275 2204 1284
rect 1797 1264 1848 1272
rect 1895 1264 2159 1272
rect 2185 1272 2204 1275
rect 2211 1272 2238 1284
rect 2185 1264 2238 1272
rect 1813 1256 1814 1264
rect 1829 1256 1842 1264
rect 1813 1248 1829 1256
rect 1810 1241 1829 1244
rect 1810 1232 1832 1241
rect 1783 1222 1832 1232
rect 1783 1216 1813 1222
rect 1832 1217 1837 1222
rect 1755 1200 1829 1216
rect 1847 1208 1877 1264
rect 1912 1254 2120 1264
rect 2155 1260 2200 1264
rect 2203 1263 2204 1264
rect 2219 1263 2232 1264
rect 1938 1224 2127 1254
rect 1953 1221 2127 1224
rect 1946 1218 2127 1221
rect 1755 1198 1768 1200
rect 1783 1198 1817 1200
rect 1755 1182 1829 1198
rect 1856 1194 1869 1208
rect 1884 1194 1900 1210
rect 1946 1205 1957 1218
rect 1739 1160 1740 1176
rect 1755 1160 1768 1182
rect 1783 1160 1813 1182
rect 1856 1178 1918 1194
rect 1946 1187 1957 1203
rect 1962 1198 1972 1218
rect 1982 1198 1996 1218
rect 1999 1205 2008 1218
rect 2024 1205 2033 1218
rect 1962 1187 1996 1198
rect 1999 1187 2008 1203
rect 2024 1187 2033 1203
rect 2040 1198 2050 1218
rect 2060 1198 2074 1218
rect 2075 1205 2086 1218
rect 2040 1187 2074 1198
rect 2075 1187 2086 1203
rect 2132 1194 2148 1210
rect 2155 1208 2185 1260
rect 2219 1256 2220 1263
rect 2204 1248 2220 1256
rect 2191 1216 2204 1235
rect 2219 1216 2249 1232
rect 2191 1200 2265 1216
rect 2191 1198 2204 1200
rect 2219 1198 2253 1200
rect 1856 1176 1869 1178
rect 1884 1176 1918 1178
rect 1856 1160 1918 1176
rect 1962 1171 1978 1174
rect 2040 1171 2070 1182
rect 2118 1178 2164 1194
rect 2191 1182 2265 1198
rect 2118 1176 2152 1178
rect 2117 1160 2164 1176
rect 2191 1160 2204 1182
rect 2219 1160 2249 1182
rect 2276 1160 2277 1176
rect 2292 1160 2305 1320
rect 2335 1216 2348 1320
rect 2393 1298 2394 1308
rect 2409 1298 2422 1308
rect 2393 1294 2422 1298
rect 2427 1294 2457 1320
rect 2475 1306 2491 1308
rect 2563 1306 2616 1320
rect 2564 1304 2628 1306
rect 2671 1304 2686 1320
rect 2735 1317 2765 1320
rect 2735 1314 2771 1317
rect 2701 1306 2717 1308
rect 2475 1294 2490 1298
rect 2393 1292 2490 1294
rect 2518 1292 2686 1304
rect 2702 1294 2717 1298
rect 2735 1295 2774 1314
rect 2793 1308 2800 1309
rect 2799 1301 2800 1308
rect 2783 1298 2784 1301
rect 2799 1298 2812 1301
rect 2735 1294 2765 1295
rect 2774 1294 2780 1295
rect 2783 1294 2812 1298
rect 2702 1293 2812 1294
rect 2702 1292 2818 1293
rect 2377 1284 2428 1292
rect 2377 1272 2402 1284
rect 2409 1272 2428 1284
rect 2459 1284 2509 1292
rect 2459 1276 2475 1284
rect 2482 1282 2509 1284
rect 2518 1282 2739 1292
rect 2482 1272 2739 1282
rect 2768 1284 2818 1292
rect 2768 1275 2784 1284
rect 2377 1264 2428 1272
rect 2475 1264 2739 1272
rect 2765 1272 2784 1275
rect 2791 1272 2818 1284
rect 2765 1264 2818 1272
rect 2393 1256 2394 1264
rect 2409 1256 2422 1264
rect 2393 1248 2409 1256
rect 2390 1241 2409 1244
rect 2390 1232 2412 1241
rect 2363 1222 2412 1232
rect 2363 1216 2393 1222
rect 2412 1217 2417 1222
rect 2335 1200 2409 1216
rect 2427 1208 2457 1264
rect 2492 1254 2700 1264
rect 2735 1260 2780 1264
rect 2783 1263 2784 1264
rect 2799 1263 2812 1264
rect 2518 1224 2707 1254
rect 2533 1221 2707 1224
rect 2526 1218 2707 1221
rect 2335 1198 2348 1200
rect 2363 1198 2397 1200
rect 2335 1182 2409 1198
rect 2436 1194 2449 1208
rect 2464 1194 2480 1210
rect 2526 1205 2537 1218
rect 2319 1160 2320 1176
rect 2335 1160 2348 1182
rect 2363 1160 2393 1182
rect 2436 1178 2498 1194
rect 2526 1187 2537 1203
rect 2542 1198 2552 1218
rect 2562 1198 2576 1218
rect 2579 1205 2588 1218
rect 2604 1205 2613 1218
rect 2542 1187 2576 1198
rect 2579 1187 2588 1203
rect 2604 1187 2613 1203
rect 2620 1198 2630 1218
rect 2640 1198 2654 1218
rect 2655 1205 2666 1218
rect 2620 1187 2654 1198
rect 2655 1187 2666 1203
rect 2712 1194 2728 1210
rect 2735 1208 2765 1260
rect 2799 1256 2800 1263
rect 2784 1248 2800 1256
rect 2771 1216 2784 1235
rect 2799 1216 2829 1232
rect 2771 1200 2845 1216
rect 2771 1198 2784 1200
rect 2799 1198 2833 1200
rect 2436 1176 2449 1178
rect 2464 1176 2498 1178
rect 2436 1160 2498 1176
rect 2542 1171 2558 1174
rect 2620 1171 2650 1182
rect 2698 1178 2744 1194
rect 2771 1182 2845 1198
rect 2698 1176 2732 1178
rect 2697 1160 2744 1176
rect 2771 1160 2784 1182
rect 2799 1160 2829 1182
rect 2856 1160 2857 1176
rect 2872 1160 2885 1320
rect 2915 1216 2928 1320
rect 2973 1298 2974 1308
rect 2989 1298 3002 1308
rect 2973 1294 3002 1298
rect 3007 1294 3037 1320
rect 3055 1306 3071 1308
rect 3143 1306 3196 1320
rect 3144 1304 3208 1306
rect 3251 1304 3266 1320
rect 3315 1317 3345 1320
rect 3315 1314 3351 1317
rect 3281 1306 3297 1308
rect 3055 1294 3070 1298
rect 2973 1292 3070 1294
rect 3098 1292 3266 1304
rect 3282 1294 3297 1298
rect 3315 1295 3354 1314
rect 3373 1308 3380 1309
rect 3379 1301 3380 1308
rect 3363 1298 3364 1301
rect 3379 1298 3392 1301
rect 3315 1294 3345 1295
rect 3354 1294 3360 1295
rect 3363 1294 3392 1298
rect 3282 1293 3392 1294
rect 3282 1292 3398 1293
rect 2957 1284 3008 1292
rect 2957 1272 2982 1284
rect 2989 1272 3008 1284
rect 3039 1284 3089 1292
rect 3039 1276 3055 1284
rect 3062 1282 3089 1284
rect 3098 1282 3319 1292
rect 3062 1272 3319 1282
rect 3348 1284 3398 1292
rect 3348 1275 3364 1284
rect 2957 1264 3008 1272
rect 3055 1264 3319 1272
rect 3345 1272 3364 1275
rect 3371 1272 3398 1284
rect 3345 1264 3398 1272
rect 2973 1256 2974 1264
rect 2989 1256 3002 1264
rect 2973 1248 2989 1256
rect 2970 1241 2989 1244
rect 2970 1232 2992 1241
rect 2943 1222 2992 1232
rect 2943 1216 2973 1222
rect 2992 1217 2997 1222
rect 2915 1200 2989 1216
rect 3007 1208 3037 1264
rect 3072 1254 3280 1264
rect 3315 1260 3360 1264
rect 3363 1263 3364 1264
rect 3379 1263 3392 1264
rect 3098 1224 3287 1254
rect 3113 1221 3287 1224
rect 3106 1218 3287 1221
rect 2915 1198 2928 1200
rect 2943 1198 2977 1200
rect 2915 1182 2989 1198
rect 3016 1194 3029 1208
rect 3044 1194 3060 1210
rect 3106 1205 3117 1218
rect 2899 1160 2900 1176
rect 2915 1160 2928 1182
rect 2943 1160 2973 1182
rect 3016 1178 3078 1194
rect 3106 1187 3117 1203
rect 3122 1198 3132 1218
rect 3142 1198 3156 1218
rect 3159 1205 3168 1218
rect 3184 1205 3193 1218
rect 3122 1187 3156 1198
rect 3159 1187 3168 1203
rect 3184 1187 3193 1203
rect 3200 1198 3210 1218
rect 3220 1198 3234 1218
rect 3235 1205 3246 1218
rect 3200 1187 3234 1198
rect 3235 1187 3246 1203
rect 3292 1194 3308 1210
rect 3315 1208 3345 1260
rect 3379 1256 3380 1263
rect 3364 1248 3380 1256
rect 3351 1216 3364 1235
rect 3379 1216 3409 1232
rect 3351 1200 3425 1216
rect 3351 1198 3364 1200
rect 3379 1198 3413 1200
rect 3016 1176 3029 1178
rect 3044 1176 3078 1178
rect 3016 1160 3078 1176
rect 3122 1171 3138 1174
rect 3200 1171 3230 1182
rect 3278 1178 3324 1194
rect 3351 1182 3425 1198
rect 3278 1176 3312 1178
rect 3277 1160 3324 1176
rect 3351 1160 3364 1182
rect 3379 1160 3409 1182
rect 3436 1160 3437 1176
rect 3452 1160 3465 1320
rect 3495 1216 3508 1320
rect 3553 1298 3554 1308
rect 3569 1298 3582 1308
rect 3553 1294 3582 1298
rect 3587 1294 3617 1320
rect 3635 1306 3651 1308
rect 3723 1306 3776 1320
rect 3724 1304 3788 1306
rect 3831 1304 3846 1320
rect 3895 1317 3925 1320
rect 3895 1314 3931 1317
rect 3861 1306 3877 1308
rect 3635 1294 3650 1298
rect 3553 1292 3650 1294
rect 3678 1292 3846 1304
rect 3862 1294 3877 1298
rect 3895 1295 3934 1314
rect 3953 1308 3960 1309
rect 3959 1301 3960 1308
rect 3943 1298 3944 1301
rect 3959 1298 3972 1301
rect 3895 1294 3925 1295
rect 3934 1294 3940 1295
rect 3943 1294 3972 1298
rect 3862 1293 3972 1294
rect 3862 1292 3978 1293
rect 3537 1284 3588 1292
rect 3537 1272 3562 1284
rect 3569 1272 3588 1284
rect 3619 1284 3669 1292
rect 3619 1276 3635 1284
rect 3642 1282 3669 1284
rect 3678 1282 3899 1292
rect 3642 1272 3899 1282
rect 3928 1284 3978 1292
rect 3928 1275 3944 1284
rect 3537 1264 3588 1272
rect 3635 1264 3899 1272
rect 3925 1272 3944 1275
rect 3951 1272 3978 1284
rect 3925 1264 3978 1272
rect 3553 1256 3554 1264
rect 3569 1256 3582 1264
rect 3553 1248 3569 1256
rect 3550 1241 3569 1244
rect 3550 1232 3572 1241
rect 3523 1222 3572 1232
rect 3523 1216 3553 1222
rect 3572 1217 3577 1222
rect 3495 1200 3569 1216
rect 3587 1208 3617 1264
rect 3652 1254 3860 1264
rect 3895 1260 3940 1264
rect 3943 1263 3944 1264
rect 3959 1263 3972 1264
rect 3678 1224 3867 1254
rect 3693 1221 3867 1224
rect 3686 1218 3867 1221
rect 3495 1198 3508 1200
rect 3523 1198 3557 1200
rect 3495 1182 3569 1198
rect 3596 1194 3609 1208
rect 3624 1194 3640 1210
rect 3686 1205 3697 1218
rect 3479 1160 3480 1176
rect 3495 1160 3508 1182
rect 3523 1160 3553 1182
rect 3596 1178 3658 1194
rect 3686 1187 3697 1203
rect 3702 1198 3712 1218
rect 3722 1198 3736 1218
rect 3739 1205 3748 1218
rect 3764 1205 3773 1218
rect 3702 1187 3736 1198
rect 3739 1187 3748 1203
rect 3764 1187 3773 1203
rect 3780 1198 3790 1218
rect 3800 1198 3814 1218
rect 3815 1205 3826 1218
rect 3780 1187 3814 1198
rect 3815 1187 3826 1203
rect 3872 1194 3888 1210
rect 3895 1208 3925 1260
rect 3959 1256 3960 1263
rect 3944 1248 3960 1256
rect 3931 1216 3944 1235
rect 3959 1216 3989 1232
rect 3931 1200 4005 1216
rect 3931 1198 3944 1200
rect 3959 1198 3993 1200
rect 3596 1176 3609 1178
rect 3624 1176 3658 1178
rect 3596 1160 3658 1176
rect 3702 1171 3718 1174
rect 3780 1171 3810 1182
rect 3858 1178 3904 1194
rect 3931 1182 4005 1198
rect 3858 1176 3892 1178
rect 3857 1160 3904 1176
rect 3931 1160 3944 1182
rect 3959 1160 3989 1182
rect 4016 1160 4017 1176
rect 4032 1160 4045 1320
rect 4075 1216 4088 1320
rect 4133 1298 4134 1308
rect 4149 1298 4162 1308
rect 4133 1294 4162 1298
rect 4167 1294 4197 1320
rect 4215 1306 4231 1308
rect 4303 1306 4356 1320
rect 4304 1304 4368 1306
rect 4411 1304 4426 1320
rect 4475 1317 4505 1320
rect 4475 1314 4511 1317
rect 4441 1306 4457 1308
rect 4215 1294 4230 1298
rect 4133 1292 4230 1294
rect 4258 1292 4426 1304
rect 4442 1294 4457 1298
rect 4475 1295 4514 1314
rect 4533 1308 4540 1309
rect 4539 1301 4540 1308
rect 4523 1298 4524 1301
rect 4539 1298 4552 1301
rect 4475 1294 4505 1295
rect 4514 1294 4520 1295
rect 4523 1294 4552 1298
rect 4442 1293 4552 1294
rect 4442 1292 4558 1293
rect 4117 1284 4168 1292
rect 4117 1272 4142 1284
rect 4149 1272 4168 1284
rect 4199 1284 4249 1292
rect 4199 1276 4215 1284
rect 4222 1282 4249 1284
rect 4258 1282 4479 1292
rect 4222 1272 4479 1282
rect 4508 1284 4558 1292
rect 4508 1275 4524 1284
rect 4117 1264 4168 1272
rect 4215 1264 4479 1272
rect 4505 1272 4524 1275
rect 4531 1272 4558 1284
rect 4505 1264 4558 1272
rect 4133 1256 4134 1264
rect 4149 1256 4162 1264
rect 4133 1248 4149 1256
rect 4130 1241 4149 1244
rect 4130 1232 4152 1241
rect 4103 1222 4152 1232
rect 4103 1216 4133 1222
rect 4152 1217 4157 1222
rect 4075 1200 4149 1216
rect 4167 1208 4197 1264
rect 4232 1254 4440 1264
rect 4475 1260 4520 1264
rect 4523 1263 4524 1264
rect 4539 1263 4552 1264
rect 4258 1224 4447 1254
rect 4273 1221 4447 1224
rect 4266 1218 4447 1221
rect 4075 1198 4088 1200
rect 4103 1198 4137 1200
rect 4075 1182 4149 1198
rect 4176 1194 4189 1208
rect 4204 1194 4220 1210
rect 4266 1205 4277 1218
rect 4059 1160 4060 1176
rect 4075 1160 4088 1182
rect 4103 1160 4133 1182
rect 4176 1178 4238 1194
rect 4266 1187 4277 1203
rect 4282 1198 4292 1218
rect 4302 1198 4316 1218
rect 4319 1205 4328 1218
rect 4344 1205 4353 1218
rect 4282 1187 4316 1198
rect 4319 1187 4328 1203
rect 4344 1187 4353 1203
rect 4360 1198 4370 1218
rect 4380 1198 4394 1218
rect 4395 1205 4406 1218
rect 4360 1187 4394 1198
rect 4395 1187 4406 1203
rect 4452 1194 4468 1210
rect 4475 1208 4505 1260
rect 4539 1256 4540 1263
rect 4524 1248 4540 1256
rect 4511 1216 4524 1235
rect 4539 1216 4569 1232
rect 4511 1200 4585 1216
rect 4511 1198 4524 1200
rect 4539 1198 4573 1200
rect 4176 1176 4189 1178
rect 4204 1176 4238 1178
rect 4176 1160 4238 1176
rect 4282 1171 4298 1174
rect 4360 1171 4390 1182
rect 4438 1178 4484 1194
rect 4511 1182 4585 1198
rect 4438 1176 4472 1178
rect 4437 1160 4484 1176
rect 4511 1160 4524 1182
rect 4539 1160 4569 1182
rect 4596 1160 4597 1176
rect 4612 1160 4625 1320
rect -7 1152 34 1160
rect -7 1126 8 1152
rect 15 1126 34 1152
rect 98 1148 160 1160
rect 172 1148 247 1160
rect 305 1148 380 1160
rect 392 1148 423 1160
rect 429 1148 464 1160
rect 98 1146 260 1148
rect -7 1118 34 1126
rect 116 1122 129 1146
rect 144 1144 159 1146
rect -1 1108 0 1118
rect 15 1108 28 1118
rect 43 1108 73 1122
rect 116 1108 159 1122
rect 183 1119 190 1126
rect 193 1122 260 1146
rect 292 1146 464 1148
rect 262 1124 290 1128
rect 292 1124 372 1146
rect 393 1144 408 1146
rect 262 1122 372 1124
rect 193 1118 372 1122
rect 166 1108 196 1118
rect 198 1108 351 1118
rect 359 1108 389 1118
rect 393 1108 423 1122
rect 451 1108 464 1146
rect 536 1152 571 1160
rect 536 1126 537 1152
rect 544 1126 571 1152
rect 479 1108 509 1122
rect 536 1118 571 1126
rect 573 1152 614 1160
rect 573 1126 588 1152
rect 595 1126 614 1152
rect 678 1148 740 1160
rect 752 1148 827 1160
rect 885 1148 960 1160
rect 972 1148 1003 1160
rect 1009 1148 1044 1160
rect 678 1146 840 1148
rect 573 1118 614 1126
rect 696 1122 709 1146
rect 724 1144 739 1146
rect 536 1108 537 1118
rect 552 1108 565 1118
rect 579 1108 580 1118
rect 595 1108 608 1118
rect 623 1108 653 1122
rect 696 1108 739 1122
rect 763 1119 770 1126
rect 773 1122 840 1146
rect 872 1146 1044 1148
rect 842 1124 870 1128
rect 872 1124 952 1146
rect 973 1144 988 1146
rect 842 1122 952 1124
rect 773 1118 952 1122
rect 746 1108 776 1118
rect 778 1108 931 1118
rect 939 1108 969 1118
rect 973 1108 1003 1122
rect 1031 1108 1044 1146
rect 1116 1152 1151 1160
rect 1116 1126 1117 1152
rect 1124 1126 1151 1152
rect 1059 1108 1089 1122
rect 1116 1118 1151 1126
rect 1153 1152 1194 1160
rect 1153 1126 1168 1152
rect 1175 1126 1194 1152
rect 1258 1148 1320 1160
rect 1332 1148 1407 1160
rect 1465 1148 1540 1160
rect 1552 1148 1583 1160
rect 1589 1148 1624 1160
rect 1258 1146 1420 1148
rect 1153 1118 1194 1126
rect 1276 1122 1289 1146
rect 1304 1144 1319 1146
rect 1116 1108 1117 1118
rect 1132 1108 1145 1118
rect 1159 1108 1160 1118
rect 1175 1108 1188 1118
rect 1203 1108 1233 1122
rect 1276 1108 1319 1122
rect 1343 1119 1350 1126
rect 1353 1122 1420 1146
rect 1452 1146 1624 1148
rect 1422 1124 1450 1128
rect 1452 1124 1532 1146
rect 1553 1144 1568 1146
rect 1422 1122 1532 1124
rect 1353 1118 1532 1122
rect 1326 1108 1356 1118
rect 1358 1108 1511 1118
rect 1519 1108 1549 1118
rect 1553 1108 1583 1122
rect 1611 1108 1624 1146
rect 1696 1152 1731 1160
rect 1696 1126 1697 1152
rect 1704 1126 1731 1152
rect 1639 1108 1669 1122
rect 1696 1118 1731 1126
rect 1733 1152 1774 1160
rect 1733 1126 1748 1152
rect 1755 1126 1774 1152
rect 1838 1148 1900 1160
rect 1912 1148 1987 1160
rect 2045 1148 2120 1160
rect 2132 1148 2163 1160
rect 2169 1148 2204 1160
rect 1838 1146 2000 1148
rect 1733 1118 1774 1126
rect 1856 1122 1869 1146
rect 1884 1144 1899 1146
rect 1696 1108 1697 1118
rect 1712 1108 1725 1118
rect 1739 1108 1740 1118
rect 1755 1108 1768 1118
rect 1783 1108 1813 1122
rect 1856 1108 1899 1122
rect 1923 1119 1930 1126
rect 1933 1122 2000 1146
rect 2032 1146 2204 1148
rect 2002 1124 2030 1128
rect 2032 1124 2112 1146
rect 2133 1144 2148 1146
rect 2002 1122 2112 1124
rect 1933 1118 2112 1122
rect 1906 1108 1936 1118
rect 1938 1108 2091 1118
rect 2099 1108 2129 1118
rect 2133 1108 2163 1122
rect 2191 1108 2204 1146
rect 2276 1152 2311 1160
rect 2276 1126 2277 1152
rect 2284 1126 2311 1152
rect 2219 1108 2249 1122
rect 2276 1118 2311 1126
rect 2313 1152 2354 1160
rect 2313 1126 2328 1152
rect 2335 1126 2354 1152
rect 2418 1148 2480 1160
rect 2492 1148 2567 1160
rect 2625 1148 2700 1160
rect 2712 1148 2743 1160
rect 2749 1148 2784 1160
rect 2418 1146 2580 1148
rect 2313 1118 2354 1126
rect 2436 1122 2449 1146
rect 2464 1144 2479 1146
rect 2276 1108 2277 1118
rect 2292 1108 2305 1118
rect 2319 1108 2320 1118
rect 2335 1108 2348 1118
rect 2363 1108 2393 1122
rect 2436 1108 2479 1122
rect 2503 1119 2510 1126
rect 2513 1122 2580 1146
rect 2612 1146 2784 1148
rect 2582 1124 2610 1128
rect 2612 1124 2692 1146
rect 2713 1144 2728 1146
rect 2582 1122 2692 1124
rect 2513 1118 2692 1122
rect 2486 1108 2516 1118
rect 2518 1108 2671 1118
rect 2679 1108 2709 1118
rect 2713 1108 2743 1122
rect 2771 1108 2784 1146
rect 2856 1152 2891 1160
rect 2856 1126 2857 1152
rect 2864 1126 2891 1152
rect 2799 1108 2829 1122
rect 2856 1118 2891 1126
rect 2893 1152 2934 1160
rect 2893 1126 2908 1152
rect 2915 1126 2934 1152
rect 2998 1148 3060 1160
rect 3072 1148 3147 1160
rect 3205 1148 3280 1160
rect 3292 1148 3323 1160
rect 3329 1148 3364 1160
rect 2998 1146 3160 1148
rect 2893 1118 2934 1126
rect 3016 1122 3029 1146
rect 3044 1144 3059 1146
rect 2856 1108 2857 1118
rect 2872 1108 2885 1118
rect 2899 1108 2900 1118
rect 2915 1108 2928 1118
rect 2943 1108 2973 1122
rect 3016 1108 3059 1122
rect 3083 1119 3090 1126
rect 3093 1122 3160 1146
rect 3192 1146 3364 1148
rect 3162 1124 3190 1128
rect 3192 1124 3272 1146
rect 3293 1144 3308 1146
rect 3162 1122 3272 1124
rect 3093 1118 3272 1122
rect 3066 1108 3096 1118
rect 3098 1108 3251 1118
rect 3259 1108 3289 1118
rect 3293 1108 3323 1122
rect 3351 1108 3364 1146
rect 3436 1152 3471 1160
rect 3436 1126 3437 1152
rect 3444 1126 3471 1152
rect 3379 1108 3409 1122
rect 3436 1118 3471 1126
rect 3473 1152 3514 1160
rect 3473 1126 3488 1152
rect 3495 1126 3514 1152
rect 3578 1148 3640 1160
rect 3652 1148 3727 1160
rect 3785 1148 3860 1160
rect 3872 1148 3903 1160
rect 3909 1148 3944 1160
rect 3578 1146 3740 1148
rect 3473 1118 3514 1126
rect 3596 1122 3609 1146
rect 3624 1144 3639 1146
rect 3436 1108 3437 1118
rect 3452 1108 3465 1118
rect 3479 1108 3480 1118
rect 3495 1108 3508 1118
rect 3523 1108 3553 1122
rect 3596 1108 3639 1122
rect 3663 1119 3670 1126
rect 3673 1122 3740 1146
rect 3772 1146 3944 1148
rect 3742 1124 3770 1128
rect 3772 1124 3852 1146
rect 3873 1144 3888 1146
rect 3742 1122 3852 1124
rect 3673 1118 3852 1122
rect 3646 1108 3676 1118
rect 3678 1108 3831 1118
rect 3839 1108 3869 1118
rect 3873 1108 3903 1122
rect 3931 1108 3944 1146
rect 4016 1152 4051 1160
rect 4016 1126 4017 1152
rect 4024 1126 4051 1152
rect 3959 1108 3989 1122
rect 4016 1118 4051 1126
rect 4053 1152 4094 1160
rect 4053 1126 4068 1152
rect 4075 1126 4094 1152
rect 4158 1148 4220 1160
rect 4232 1148 4307 1160
rect 4365 1148 4440 1160
rect 4452 1148 4483 1160
rect 4489 1148 4524 1160
rect 4158 1146 4320 1148
rect 4053 1118 4094 1126
rect 4176 1122 4189 1146
rect 4204 1144 4219 1146
rect 4016 1108 4017 1118
rect 4032 1108 4045 1118
rect 4059 1108 4060 1118
rect 4075 1108 4088 1118
rect 4103 1108 4133 1122
rect 4176 1108 4219 1122
rect 4243 1119 4250 1126
rect 4253 1122 4320 1146
rect 4352 1146 4524 1148
rect 4322 1124 4350 1128
rect 4352 1124 4432 1146
rect 4453 1144 4468 1146
rect 4322 1122 4432 1124
rect 4253 1118 4432 1122
rect 4226 1108 4256 1118
rect 4258 1108 4411 1118
rect 4419 1108 4449 1118
rect 4453 1108 4483 1122
rect 4511 1108 4524 1146
rect 4596 1152 4631 1160
rect 4596 1126 4597 1152
rect 4604 1126 4631 1152
rect 4539 1108 4569 1122
rect 4596 1118 4631 1126
rect 4596 1108 4597 1118
rect 4612 1108 4625 1118
rect -1 1102 4625 1108
rect 0 1094 4625 1102
rect 15 1064 28 1094
rect 43 1076 73 1094
rect 116 1080 130 1094
rect 166 1080 386 1094
rect 117 1078 130 1080
rect 83 1066 98 1078
rect 80 1064 102 1066
rect 107 1064 137 1078
rect 198 1076 351 1080
rect 180 1064 372 1076
rect 415 1064 445 1078
rect 451 1064 464 1094
rect 479 1076 509 1094
rect 552 1064 565 1094
rect 595 1064 608 1094
rect 623 1076 653 1094
rect 696 1080 710 1094
rect 746 1080 966 1094
rect 697 1078 710 1080
rect 663 1066 678 1078
rect 660 1064 682 1066
rect 687 1064 717 1078
rect 778 1076 931 1080
rect 760 1064 952 1076
rect 995 1064 1025 1078
rect 1031 1064 1044 1094
rect 1059 1076 1089 1094
rect 1132 1064 1145 1094
rect 1175 1064 1188 1094
rect 1203 1076 1233 1094
rect 1276 1080 1290 1094
rect 1326 1080 1546 1094
rect 1277 1078 1290 1080
rect 1243 1066 1258 1078
rect 1240 1064 1262 1066
rect 1267 1064 1297 1078
rect 1358 1076 1511 1080
rect 1340 1064 1532 1076
rect 1575 1064 1605 1078
rect 1611 1064 1624 1094
rect 1639 1076 1669 1094
rect 1712 1064 1725 1094
rect 1755 1064 1768 1094
rect 1783 1076 1813 1094
rect 1856 1080 1870 1094
rect 1906 1080 2126 1094
rect 1857 1078 1870 1080
rect 1823 1066 1838 1078
rect 1820 1064 1842 1066
rect 1847 1064 1877 1078
rect 1938 1076 2091 1080
rect 1920 1064 2112 1076
rect 2155 1064 2185 1078
rect 2191 1064 2204 1094
rect 2219 1076 2249 1094
rect 2292 1064 2305 1094
rect 2335 1064 2348 1094
rect 2363 1076 2393 1094
rect 2436 1080 2450 1094
rect 2486 1080 2706 1094
rect 2437 1078 2450 1080
rect 2403 1066 2418 1078
rect 2400 1064 2422 1066
rect 2427 1064 2457 1078
rect 2518 1076 2671 1080
rect 2500 1064 2692 1076
rect 2735 1064 2765 1078
rect 2771 1064 2784 1094
rect 2799 1076 2829 1094
rect 2872 1064 2885 1094
rect 2915 1064 2928 1094
rect 2943 1076 2973 1094
rect 3016 1080 3030 1094
rect 3066 1080 3286 1094
rect 3017 1078 3030 1080
rect 2983 1066 2998 1078
rect 2980 1064 3002 1066
rect 3007 1064 3037 1078
rect 3098 1076 3251 1080
rect 3080 1064 3272 1076
rect 3315 1064 3345 1078
rect 3351 1064 3364 1094
rect 3379 1076 3409 1094
rect 3452 1064 3465 1094
rect 3495 1064 3508 1094
rect 3523 1076 3553 1094
rect 3596 1080 3610 1094
rect 3646 1080 3866 1094
rect 3597 1078 3610 1080
rect 3563 1066 3578 1078
rect 3560 1064 3582 1066
rect 3587 1064 3617 1078
rect 3678 1076 3831 1080
rect 3660 1064 3852 1076
rect 3895 1064 3925 1078
rect 3931 1064 3944 1094
rect 3959 1076 3989 1094
rect 4032 1064 4045 1094
rect 4075 1064 4088 1094
rect 4103 1076 4133 1094
rect 4176 1080 4190 1094
rect 4226 1080 4446 1094
rect 4177 1078 4190 1080
rect 4143 1066 4158 1078
rect 4140 1064 4162 1066
rect 4167 1064 4197 1078
rect 4258 1076 4411 1080
rect 4240 1064 4432 1076
rect 4475 1064 4505 1078
rect 4511 1064 4524 1094
rect 4539 1076 4569 1094
rect 4612 1064 4625 1094
rect 0 1050 4625 1064
rect 15 946 28 1050
rect 73 1028 74 1038
rect 89 1028 102 1038
rect 73 1024 102 1028
rect 107 1024 137 1050
rect 155 1036 171 1038
rect 243 1036 296 1050
rect 244 1034 308 1036
rect 351 1034 366 1050
rect 415 1047 445 1050
rect 415 1044 451 1047
rect 381 1036 397 1038
rect 155 1024 170 1028
rect 73 1022 170 1024
rect 198 1022 366 1034
rect 382 1024 397 1028
rect 415 1025 454 1044
rect 473 1038 480 1039
rect 479 1031 480 1038
rect 463 1028 464 1031
rect 479 1028 492 1031
rect 415 1024 445 1025
rect 454 1024 460 1025
rect 463 1024 492 1028
rect 382 1023 492 1024
rect 382 1022 498 1023
rect 57 1014 108 1022
rect 57 1002 82 1014
rect 89 1002 108 1014
rect 139 1014 189 1022
rect 139 1006 155 1014
rect 162 1012 189 1014
rect 198 1012 419 1022
rect 162 1002 419 1012
rect 448 1014 498 1022
rect 448 1005 464 1014
rect 57 994 108 1002
rect 155 994 419 1002
rect 445 1002 464 1005
rect 471 1002 498 1014
rect 445 994 498 1002
rect 73 986 74 994
rect 89 986 102 994
rect 73 978 89 986
rect 70 971 89 974
rect 70 962 92 971
rect 43 952 92 962
rect 43 946 73 952
rect 92 947 97 952
rect 15 930 89 946
rect 107 938 137 994
rect 172 984 380 994
rect 415 990 460 994
rect 463 993 464 994
rect 479 993 492 994
rect 198 954 387 984
rect 213 951 387 954
rect 206 948 387 951
rect 15 928 28 930
rect 43 928 77 930
rect 15 912 89 928
rect 116 924 129 938
rect 144 924 160 940
rect 206 935 217 948
rect -1 890 0 906
rect 15 890 28 912
rect 43 890 73 912
rect 116 908 178 924
rect 206 917 217 933
rect 222 928 232 948
rect 242 928 256 948
rect 259 935 268 948
rect 284 935 293 948
rect 222 917 256 928
rect 259 917 268 933
rect 284 917 293 933
rect 300 928 310 948
rect 320 928 334 948
rect 335 935 346 948
rect 300 917 334 928
rect 335 917 346 933
rect 392 924 408 940
rect 415 938 445 990
rect 479 986 480 993
rect 464 978 480 986
rect 451 946 464 965
rect 479 946 509 962
rect 451 930 525 946
rect 451 928 464 930
rect 479 928 513 930
rect 116 906 129 908
rect 144 906 178 908
rect 116 890 178 906
rect 222 901 238 904
rect 300 901 330 912
rect 378 908 424 924
rect 451 912 525 928
rect 378 906 412 908
rect 377 890 424 906
rect 451 890 464 912
rect 479 890 509 912
rect 536 890 537 906
rect 552 890 565 1050
rect 595 946 608 1050
rect 653 1028 654 1038
rect 669 1028 682 1038
rect 653 1024 682 1028
rect 687 1024 717 1050
rect 735 1036 751 1038
rect 823 1036 876 1050
rect 824 1034 888 1036
rect 931 1034 946 1050
rect 995 1047 1025 1050
rect 995 1044 1031 1047
rect 961 1036 977 1038
rect 735 1024 750 1028
rect 653 1022 750 1024
rect 778 1022 946 1034
rect 962 1024 977 1028
rect 995 1025 1034 1044
rect 1053 1038 1060 1039
rect 1059 1031 1060 1038
rect 1043 1028 1044 1031
rect 1059 1028 1072 1031
rect 995 1024 1025 1025
rect 1034 1024 1040 1025
rect 1043 1024 1072 1028
rect 962 1023 1072 1024
rect 962 1022 1078 1023
rect 637 1014 688 1022
rect 637 1002 662 1014
rect 669 1002 688 1014
rect 719 1014 769 1022
rect 719 1006 735 1014
rect 742 1012 769 1014
rect 778 1012 999 1022
rect 742 1002 999 1012
rect 1028 1014 1078 1022
rect 1028 1005 1044 1014
rect 637 994 688 1002
rect 735 994 999 1002
rect 1025 1002 1044 1005
rect 1051 1002 1078 1014
rect 1025 994 1078 1002
rect 653 986 654 994
rect 669 986 682 994
rect 653 978 669 986
rect 650 971 669 974
rect 650 962 672 971
rect 623 952 672 962
rect 623 946 653 952
rect 672 947 677 952
rect 595 930 669 946
rect 687 938 717 994
rect 752 984 960 994
rect 995 990 1040 994
rect 1043 993 1044 994
rect 1059 993 1072 994
rect 778 954 967 984
rect 793 951 967 954
rect 786 948 967 951
rect 595 928 608 930
rect 623 928 657 930
rect 595 912 669 928
rect 696 924 709 938
rect 724 924 740 940
rect 786 935 797 948
rect 579 890 580 906
rect 595 890 608 912
rect 623 890 653 912
rect 696 908 758 924
rect 786 917 797 933
rect 802 928 812 948
rect 822 928 836 948
rect 839 935 848 948
rect 864 935 873 948
rect 802 917 836 928
rect 839 917 848 933
rect 864 917 873 933
rect 880 928 890 948
rect 900 928 914 948
rect 915 935 926 948
rect 880 917 914 928
rect 915 917 926 933
rect 972 924 988 940
rect 995 938 1025 990
rect 1059 986 1060 993
rect 1044 978 1060 986
rect 1031 946 1044 965
rect 1059 946 1089 962
rect 1031 930 1105 946
rect 1031 928 1044 930
rect 1059 928 1093 930
rect 696 906 709 908
rect 724 906 758 908
rect 696 890 758 906
rect 802 901 818 904
rect 880 901 910 912
rect 958 908 1004 924
rect 1031 912 1105 928
rect 958 906 992 908
rect 957 890 1004 906
rect 1031 890 1044 912
rect 1059 890 1089 912
rect 1116 890 1117 906
rect 1132 890 1145 1050
rect 1175 946 1188 1050
rect 1233 1028 1234 1038
rect 1249 1028 1262 1038
rect 1233 1024 1262 1028
rect 1267 1024 1297 1050
rect 1315 1036 1331 1038
rect 1403 1036 1456 1050
rect 1404 1034 1468 1036
rect 1511 1034 1526 1050
rect 1575 1047 1605 1050
rect 1575 1044 1611 1047
rect 1541 1036 1557 1038
rect 1315 1024 1330 1028
rect 1233 1022 1330 1024
rect 1358 1022 1526 1034
rect 1542 1024 1557 1028
rect 1575 1025 1614 1044
rect 1633 1038 1640 1039
rect 1639 1031 1640 1038
rect 1623 1028 1624 1031
rect 1639 1028 1652 1031
rect 1575 1024 1605 1025
rect 1614 1024 1620 1025
rect 1623 1024 1652 1028
rect 1542 1023 1652 1024
rect 1542 1022 1658 1023
rect 1217 1014 1268 1022
rect 1217 1002 1242 1014
rect 1249 1002 1268 1014
rect 1299 1014 1349 1022
rect 1299 1006 1315 1014
rect 1322 1012 1349 1014
rect 1358 1012 1579 1022
rect 1322 1002 1579 1012
rect 1608 1014 1658 1022
rect 1608 1005 1624 1014
rect 1217 994 1268 1002
rect 1315 994 1579 1002
rect 1605 1002 1624 1005
rect 1631 1002 1658 1014
rect 1605 994 1658 1002
rect 1233 986 1234 994
rect 1249 986 1262 994
rect 1233 978 1249 986
rect 1230 971 1249 974
rect 1230 962 1252 971
rect 1203 952 1252 962
rect 1203 946 1233 952
rect 1252 947 1257 952
rect 1175 930 1249 946
rect 1267 938 1297 994
rect 1332 984 1540 994
rect 1575 990 1620 994
rect 1623 993 1624 994
rect 1639 993 1652 994
rect 1358 954 1547 984
rect 1373 951 1547 954
rect 1366 948 1547 951
rect 1175 928 1188 930
rect 1203 928 1237 930
rect 1175 912 1249 928
rect 1276 924 1289 938
rect 1304 924 1320 940
rect 1366 935 1377 948
rect 1159 890 1160 906
rect 1175 890 1188 912
rect 1203 890 1233 912
rect 1276 908 1338 924
rect 1366 917 1377 933
rect 1382 928 1392 948
rect 1402 928 1416 948
rect 1419 935 1428 948
rect 1444 935 1453 948
rect 1382 917 1416 928
rect 1419 917 1428 933
rect 1444 917 1453 933
rect 1460 928 1470 948
rect 1480 928 1494 948
rect 1495 935 1506 948
rect 1460 917 1494 928
rect 1495 917 1506 933
rect 1552 924 1568 940
rect 1575 938 1605 990
rect 1639 986 1640 993
rect 1624 978 1640 986
rect 1611 946 1624 965
rect 1639 946 1669 962
rect 1611 930 1685 946
rect 1611 928 1624 930
rect 1639 928 1673 930
rect 1276 906 1289 908
rect 1304 906 1338 908
rect 1276 890 1338 906
rect 1382 901 1398 904
rect 1460 901 1490 912
rect 1538 908 1584 924
rect 1611 912 1685 928
rect 1538 906 1572 908
rect 1537 890 1584 906
rect 1611 890 1624 912
rect 1639 890 1669 912
rect 1696 890 1697 906
rect 1712 890 1725 1050
rect 1755 946 1768 1050
rect 1813 1028 1814 1038
rect 1829 1028 1842 1038
rect 1813 1024 1842 1028
rect 1847 1024 1877 1050
rect 1895 1036 1911 1038
rect 1983 1036 2036 1050
rect 1984 1034 2048 1036
rect 2091 1034 2106 1050
rect 2155 1047 2185 1050
rect 2155 1044 2191 1047
rect 2121 1036 2137 1038
rect 1895 1024 1910 1028
rect 1813 1022 1910 1024
rect 1938 1022 2106 1034
rect 2122 1024 2137 1028
rect 2155 1025 2194 1044
rect 2213 1038 2220 1039
rect 2219 1031 2220 1038
rect 2203 1028 2204 1031
rect 2219 1028 2232 1031
rect 2155 1024 2185 1025
rect 2194 1024 2200 1025
rect 2203 1024 2232 1028
rect 2122 1023 2232 1024
rect 2122 1022 2238 1023
rect 1797 1014 1848 1022
rect 1797 1002 1822 1014
rect 1829 1002 1848 1014
rect 1879 1014 1929 1022
rect 1879 1006 1895 1014
rect 1902 1012 1929 1014
rect 1938 1012 2159 1022
rect 1902 1002 2159 1012
rect 2188 1014 2238 1022
rect 2188 1005 2204 1014
rect 1797 994 1848 1002
rect 1895 994 2159 1002
rect 2185 1002 2204 1005
rect 2211 1002 2238 1014
rect 2185 994 2238 1002
rect 1813 986 1814 994
rect 1829 986 1842 994
rect 1813 978 1829 986
rect 1810 971 1829 974
rect 1810 962 1832 971
rect 1783 952 1832 962
rect 1783 946 1813 952
rect 1832 947 1837 952
rect 1755 930 1829 946
rect 1847 938 1877 994
rect 1912 984 2120 994
rect 2155 990 2200 994
rect 2203 993 2204 994
rect 2219 993 2232 994
rect 1938 954 2127 984
rect 1953 951 2127 954
rect 1946 948 2127 951
rect 1755 928 1768 930
rect 1783 928 1817 930
rect 1755 912 1829 928
rect 1856 924 1869 938
rect 1884 924 1900 940
rect 1946 935 1957 948
rect 1739 890 1740 906
rect 1755 890 1768 912
rect 1783 890 1813 912
rect 1856 908 1918 924
rect 1946 917 1957 933
rect 1962 928 1972 948
rect 1982 928 1996 948
rect 1999 935 2008 948
rect 2024 935 2033 948
rect 1962 917 1996 928
rect 1999 917 2008 933
rect 2024 917 2033 933
rect 2040 928 2050 948
rect 2060 928 2074 948
rect 2075 935 2086 948
rect 2040 917 2074 928
rect 2075 917 2086 933
rect 2132 924 2148 940
rect 2155 938 2185 990
rect 2219 986 2220 993
rect 2204 978 2220 986
rect 2191 946 2204 965
rect 2219 946 2249 962
rect 2191 930 2265 946
rect 2191 928 2204 930
rect 2219 928 2253 930
rect 1856 906 1869 908
rect 1884 906 1918 908
rect 1856 890 1918 906
rect 1962 901 1978 904
rect 2040 901 2070 912
rect 2118 908 2164 924
rect 2191 912 2265 928
rect 2118 906 2152 908
rect 2117 890 2164 906
rect 2191 890 2204 912
rect 2219 890 2249 912
rect 2276 890 2277 906
rect 2292 890 2305 1050
rect 2335 946 2348 1050
rect 2393 1028 2394 1038
rect 2409 1028 2422 1038
rect 2393 1024 2422 1028
rect 2427 1024 2457 1050
rect 2475 1036 2491 1038
rect 2563 1036 2616 1050
rect 2564 1034 2628 1036
rect 2671 1034 2686 1050
rect 2735 1047 2765 1050
rect 2735 1044 2771 1047
rect 2701 1036 2717 1038
rect 2475 1024 2490 1028
rect 2393 1022 2490 1024
rect 2518 1022 2686 1034
rect 2702 1024 2717 1028
rect 2735 1025 2774 1044
rect 2793 1038 2800 1039
rect 2799 1031 2800 1038
rect 2783 1028 2784 1031
rect 2799 1028 2812 1031
rect 2735 1024 2765 1025
rect 2774 1024 2780 1025
rect 2783 1024 2812 1028
rect 2702 1023 2812 1024
rect 2702 1022 2818 1023
rect 2377 1014 2428 1022
rect 2377 1002 2402 1014
rect 2409 1002 2428 1014
rect 2459 1014 2509 1022
rect 2459 1006 2475 1014
rect 2482 1012 2509 1014
rect 2518 1012 2739 1022
rect 2482 1002 2739 1012
rect 2768 1014 2818 1022
rect 2768 1005 2784 1014
rect 2377 994 2428 1002
rect 2475 994 2739 1002
rect 2765 1002 2784 1005
rect 2791 1002 2818 1014
rect 2765 994 2818 1002
rect 2393 986 2394 994
rect 2409 986 2422 994
rect 2393 978 2409 986
rect 2390 971 2409 974
rect 2390 962 2412 971
rect 2363 952 2412 962
rect 2363 946 2393 952
rect 2412 947 2417 952
rect 2335 930 2409 946
rect 2427 938 2457 994
rect 2492 984 2700 994
rect 2735 990 2780 994
rect 2783 993 2784 994
rect 2799 993 2812 994
rect 2518 954 2707 984
rect 2533 951 2707 954
rect 2526 948 2707 951
rect 2335 928 2348 930
rect 2363 928 2397 930
rect 2335 912 2409 928
rect 2436 924 2449 938
rect 2464 924 2480 940
rect 2526 935 2537 948
rect 2319 890 2320 906
rect 2335 890 2348 912
rect 2363 890 2393 912
rect 2436 908 2498 924
rect 2526 917 2537 933
rect 2542 928 2552 948
rect 2562 928 2576 948
rect 2579 935 2588 948
rect 2604 935 2613 948
rect 2542 917 2576 928
rect 2579 917 2588 933
rect 2604 917 2613 933
rect 2620 928 2630 948
rect 2640 928 2654 948
rect 2655 935 2666 948
rect 2620 917 2654 928
rect 2655 917 2666 933
rect 2712 924 2728 940
rect 2735 938 2765 990
rect 2799 986 2800 993
rect 2784 978 2800 986
rect 2771 946 2784 965
rect 2799 946 2829 962
rect 2771 930 2845 946
rect 2771 928 2784 930
rect 2799 928 2833 930
rect 2436 906 2449 908
rect 2464 906 2498 908
rect 2436 890 2498 906
rect 2542 901 2558 904
rect 2620 901 2650 912
rect 2698 908 2744 924
rect 2771 912 2845 928
rect 2698 906 2732 908
rect 2697 890 2744 906
rect 2771 890 2784 912
rect 2799 890 2829 912
rect 2856 890 2857 906
rect 2872 890 2885 1050
rect 2915 946 2928 1050
rect 2973 1028 2974 1038
rect 2989 1028 3002 1038
rect 2973 1024 3002 1028
rect 3007 1024 3037 1050
rect 3055 1036 3071 1038
rect 3143 1036 3196 1050
rect 3144 1034 3208 1036
rect 3251 1034 3266 1050
rect 3315 1047 3345 1050
rect 3315 1044 3351 1047
rect 3281 1036 3297 1038
rect 3055 1024 3070 1028
rect 2973 1022 3070 1024
rect 3098 1022 3266 1034
rect 3282 1024 3297 1028
rect 3315 1025 3354 1044
rect 3373 1038 3380 1039
rect 3379 1031 3380 1038
rect 3363 1028 3364 1031
rect 3379 1028 3392 1031
rect 3315 1024 3345 1025
rect 3354 1024 3360 1025
rect 3363 1024 3392 1028
rect 3282 1023 3392 1024
rect 3282 1022 3398 1023
rect 2957 1014 3008 1022
rect 2957 1002 2982 1014
rect 2989 1002 3008 1014
rect 3039 1014 3089 1022
rect 3039 1006 3055 1014
rect 3062 1012 3089 1014
rect 3098 1012 3319 1022
rect 3062 1002 3319 1012
rect 3348 1014 3398 1022
rect 3348 1005 3364 1014
rect 2957 994 3008 1002
rect 3055 994 3319 1002
rect 3345 1002 3364 1005
rect 3371 1002 3398 1014
rect 3345 994 3398 1002
rect 2973 986 2974 994
rect 2989 986 3002 994
rect 2973 978 2989 986
rect 2970 971 2989 974
rect 2970 962 2992 971
rect 2943 952 2992 962
rect 2943 946 2973 952
rect 2992 947 2997 952
rect 2915 930 2989 946
rect 3007 938 3037 994
rect 3072 984 3280 994
rect 3315 990 3360 994
rect 3363 993 3364 994
rect 3379 993 3392 994
rect 3098 954 3287 984
rect 3113 951 3287 954
rect 3106 948 3287 951
rect 2915 928 2928 930
rect 2943 928 2977 930
rect 2915 912 2989 928
rect 3016 924 3029 938
rect 3044 924 3060 940
rect 3106 935 3117 948
rect 2899 890 2900 906
rect 2915 890 2928 912
rect 2943 890 2973 912
rect 3016 908 3078 924
rect 3106 917 3117 933
rect 3122 928 3132 948
rect 3142 928 3156 948
rect 3159 935 3168 948
rect 3184 935 3193 948
rect 3122 917 3156 928
rect 3159 917 3168 933
rect 3184 917 3193 933
rect 3200 928 3210 948
rect 3220 928 3234 948
rect 3235 935 3246 948
rect 3200 917 3234 928
rect 3235 917 3246 933
rect 3292 924 3308 940
rect 3315 938 3345 990
rect 3379 986 3380 993
rect 3364 978 3380 986
rect 3351 946 3364 965
rect 3379 946 3409 962
rect 3351 930 3425 946
rect 3351 928 3364 930
rect 3379 928 3413 930
rect 3016 906 3029 908
rect 3044 906 3078 908
rect 3016 890 3078 906
rect 3122 901 3138 904
rect 3200 901 3230 912
rect 3278 908 3324 924
rect 3351 912 3425 928
rect 3278 906 3312 908
rect 3277 890 3324 906
rect 3351 890 3364 912
rect 3379 890 3409 912
rect 3436 890 3437 906
rect 3452 890 3465 1050
rect 3495 946 3508 1050
rect 3553 1028 3554 1038
rect 3569 1028 3582 1038
rect 3553 1024 3582 1028
rect 3587 1024 3617 1050
rect 3635 1036 3651 1038
rect 3723 1036 3776 1050
rect 3724 1034 3788 1036
rect 3831 1034 3846 1050
rect 3895 1047 3925 1050
rect 3895 1044 3931 1047
rect 3861 1036 3877 1038
rect 3635 1024 3650 1028
rect 3553 1022 3650 1024
rect 3678 1022 3846 1034
rect 3862 1024 3877 1028
rect 3895 1025 3934 1044
rect 3953 1038 3960 1039
rect 3959 1031 3960 1038
rect 3943 1028 3944 1031
rect 3959 1028 3972 1031
rect 3895 1024 3925 1025
rect 3934 1024 3940 1025
rect 3943 1024 3972 1028
rect 3862 1023 3972 1024
rect 3862 1022 3978 1023
rect 3537 1014 3588 1022
rect 3537 1002 3562 1014
rect 3569 1002 3588 1014
rect 3619 1014 3669 1022
rect 3619 1006 3635 1014
rect 3642 1012 3669 1014
rect 3678 1012 3899 1022
rect 3642 1002 3899 1012
rect 3928 1014 3978 1022
rect 3928 1005 3944 1014
rect 3537 994 3588 1002
rect 3635 994 3899 1002
rect 3925 1002 3944 1005
rect 3951 1002 3978 1014
rect 3925 994 3978 1002
rect 3553 986 3554 994
rect 3569 986 3582 994
rect 3553 978 3569 986
rect 3550 971 3569 974
rect 3550 962 3572 971
rect 3523 952 3572 962
rect 3523 946 3553 952
rect 3572 947 3577 952
rect 3495 930 3569 946
rect 3587 938 3617 994
rect 3652 984 3860 994
rect 3895 990 3940 994
rect 3943 993 3944 994
rect 3959 993 3972 994
rect 3678 954 3867 984
rect 3693 951 3867 954
rect 3686 948 3867 951
rect 3495 928 3508 930
rect 3523 928 3557 930
rect 3495 912 3569 928
rect 3596 924 3609 938
rect 3624 924 3640 940
rect 3686 935 3697 948
rect 3479 890 3480 906
rect 3495 890 3508 912
rect 3523 890 3553 912
rect 3596 908 3658 924
rect 3686 917 3697 933
rect 3702 928 3712 948
rect 3722 928 3736 948
rect 3739 935 3748 948
rect 3764 935 3773 948
rect 3702 917 3736 928
rect 3739 917 3748 933
rect 3764 917 3773 933
rect 3780 928 3790 948
rect 3800 928 3814 948
rect 3815 935 3826 948
rect 3780 917 3814 928
rect 3815 917 3826 933
rect 3872 924 3888 940
rect 3895 938 3925 990
rect 3959 986 3960 993
rect 3944 978 3960 986
rect 3931 946 3944 965
rect 3959 946 3989 962
rect 3931 930 4005 946
rect 3931 928 3944 930
rect 3959 928 3993 930
rect 3596 906 3609 908
rect 3624 906 3658 908
rect 3596 890 3658 906
rect 3702 901 3718 904
rect 3780 901 3810 912
rect 3858 908 3904 924
rect 3931 912 4005 928
rect 3858 906 3892 908
rect 3857 890 3904 906
rect 3931 890 3944 912
rect 3959 890 3989 912
rect 4016 890 4017 906
rect 4032 890 4045 1050
rect 4075 946 4088 1050
rect 4133 1028 4134 1038
rect 4149 1028 4162 1038
rect 4133 1024 4162 1028
rect 4167 1024 4197 1050
rect 4215 1036 4231 1038
rect 4303 1036 4356 1050
rect 4304 1034 4368 1036
rect 4411 1034 4426 1050
rect 4475 1047 4505 1050
rect 4475 1044 4511 1047
rect 4441 1036 4457 1038
rect 4215 1024 4230 1028
rect 4133 1022 4230 1024
rect 4258 1022 4426 1034
rect 4442 1024 4457 1028
rect 4475 1025 4514 1044
rect 4533 1038 4540 1039
rect 4539 1031 4540 1038
rect 4523 1028 4524 1031
rect 4539 1028 4552 1031
rect 4475 1024 4505 1025
rect 4514 1024 4520 1025
rect 4523 1024 4552 1028
rect 4442 1023 4552 1024
rect 4442 1022 4558 1023
rect 4117 1014 4168 1022
rect 4117 1002 4142 1014
rect 4149 1002 4168 1014
rect 4199 1014 4249 1022
rect 4199 1006 4215 1014
rect 4222 1012 4249 1014
rect 4258 1012 4479 1022
rect 4222 1002 4479 1012
rect 4508 1014 4558 1022
rect 4508 1005 4524 1014
rect 4117 994 4168 1002
rect 4215 994 4479 1002
rect 4505 1002 4524 1005
rect 4531 1002 4558 1014
rect 4505 994 4558 1002
rect 4133 986 4134 994
rect 4149 986 4162 994
rect 4133 978 4149 986
rect 4130 971 4149 974
rect 4130 962 4152 971
rect 4103 952 4152 962
rect 4103 946 4133 952
rect 4152 947 4157 952
rect 4075 930 4149 946
rect 4167 938 4197 994
rect 4232 984 4440 994
rect 4475 990 4520 994
rect 4523 993 4524 994
rect 4539 993 4552 994
rect 4258 954 4447 984
rect 4273 951 4447 954
rect 4266 948 4447 951
rect 4075 928 4088 930
rect 4103 928 4137 930
rect 4075 912 4149 928
rect 4176 924 4189 938
rect 4204 924 4220 940
rect 4266 935 4277 948
rect 4059 890 4060 906
rect 4075 890 4088 912
rect 4103 890 4133 912
rect 4176 908 4238 924
rect 4266 917 4277 933
rect 4282 928 4292 948
rect 4302 928 4316 948
rect 4319 935 4328 948
rect 4344 935 4353 948
rect 4282 917 4316 928
rect 4319 917 4328 933
rect 4344 917 4353 933
rect 4360 928 4370 948
rect 4380 928 4394 948
rect 4395 935 4406 948
rect 4360 917 4394 928
rect 4395 917 4406 933
rect 4452 924 4468 940
rect 4475 938 4505 990
rect 4539 986 4540 993
rect 4524 978 4540 986
rect 4511 946 4524 965
rect 4539 946 4569 962
rect 4511 930 4585 946
rect 4511 928 4524 930
rect 4539 928 4573 930
rect 4176 906 4189 908
rect 4204 906 4238 908
rect 4176 890 4238 906
rect 4282 901 4298 904
rect 4360 901 4390 912
rect 4438 908 4484 924
rect 4511 912 4585 928
rect 4438 906 4472 908
rect 4437 890 4484 906
rect 4511 890 4524 912
rect 4539 890 4569 912
rect 4596 890 4597 906
rect 4612 890 4625 1050
rect -7 882 34 890
rect -7 856 8 882
rect 15 856 34 882
rect 98 878 160 890
rect 172 878 247 890
rect 305 878 380 890
rect 392 878 423 890
rect 429 878 464 890
rect 98 876 260 878
rect -7 848 34 856
rect 116 852 129 876
rect 144 874 159 876
rect -1 838 0 848
rect 15 838 28 848
rect 43 838 73 852
rect 116 838 159 852
rect 183 849 190 856
rect 193 852 260 876
rect 292 876 464 878
rect 262 854 290 858
rect 292 854 372 876
rect 393 874 408 876
rect 262 852 372 854
rect 193 848 372 852
rect 166 838 196 848
rect 198 838 351 848
rect 359 838 389 848
rect 393 838 423 852
rect 451 838 464 876
rect 536 882 571 890
rect 536 856 537 882
rect 544 856 571 882
rect 479 838 509 852
rect 536 848 571 856
rect 573 882 614 890
rect 573 856 588 882
rect 595 856 614 882
rect 678 878 740 890
rect 752 878 827 890
rect 885 878 960 890
rect 972 878 1003 890
rect 1009 878 1044 890
rect 678 876 840 878
rect 573 848 614 856
rect 696 852 709 876
rect 724 874 739 876
rect 536 838 537 848
rect 552 838 565 848
rect 579 838 580 848
rect 595 838 608 848
rect 623 838 653 852
rect 696 838 739 852
rect 763 849 770 856
rect 773 852 840 876
rect 872 876 1044 878
rect 842 854 870 858
rect 872 854 952 876
rect 973 874 988 876
rect 842 852 952 854
rect 773 848 952 852
rect 746 838 776 848
rect 778 838 931 848
rect 939 838 969 848
rect 973 838 1003 852
rect 1031 838 1044 876
rect 1116 882 1151 890
rect 1116 856 1117 882
rect 1124 856 1151 882
rect 1059 838 1089 852
rect 1116 848 1151 856
rect 1153 882 1194 890
rect 1153 856 1168 882
rect 1175 856 1194 882
rect 1258 878 1320 890
rect 1332 878 1407 890
rect 1465 878 1540 890
rect 1552 878 1583 890
rect 1589 878 1624 890
rect 1258 876 1420 878
rect 1153 848 1194 856
rect 1276 852 1289 876
rect 1304 874 1319 876
rect 1116 838 1117 848
rect 1132 838 1145 848
rect 1159 838 1160 848
rect 1175 838 1188 848
rect 1203 838 1233 852
rect 1276 838 1319 852
rect 1343 849 1350 856
rect 1353 852 1420 876
rect 1452 876 1624 878
rect 1422 854 1450 858
rect 1452 854 1532 876
rect 1553 874 1568 876
rect 1422 852 1532 854
rect 1353 848 1532 852
rect 1326 838 1356 848
rect 1358 838 1511 848
rect 1519 838 1549 848
rect 1553 838 1583 852
rect 1611 838 1624 876
rect 1696 882 1731 890
rect 1696 856 1697 882
rect 1704 856 1731 882
rect 1639 838 1669 852
rect 1696 848 1731 856
rect 1733 882 1774 890
rect 1733 856 1748 882
rect 1755 856 1774 882
rect 1838 878 1900 890
rect 1912 878 1987 890
rect 2045 878 2120 890
rect 2132 878 2163 890
rect 2169 878 2204 890
rect 1838 876 2000 878
rect 1733 848 1774 856
rect 1856 852 1869 876
rect 1884 874 1899 876
rect 1696 838 1697 848
rect 1712 838 1725 848
rect 1739 838 1740 848
rect 1755 838 1768 848
rect 1783 838 1813 852
rect 1856 838 1899 852
rect 1923 849 1930 856
rect 1933 852 2000 876
rect 2032 876 2204 878
rect 2002 854 2030 858
rect 2032 854 2112 876
rect 2133 874 2148 876
rect 2002 852 2112 854
rect 1933 848 2112 852
rect 1906 838 1936 848
rect 1938 838 2091 848
rect 2099 838 2129 848
rect 2133 838 2163 852
rect 2191 838 2204 876
rect 2276 882 2311 890
rect 2276 856 2277 882
rect 2284 856 2311 882
rect 2219 838 2249 852
rect 2276 848 2311 856
rect 2313 882 2354 890
rect 2313 856 2328 882
rect 2335 856 2354 882
rect 2418 878 2480 890
rect 2492 878 2567 890
rect 2625 878 2700 890
rect 2712 878 2743 890
rect 2749 878 2784 890
rect 2418 876 2580 878
rect 2313 848 2354 856
rect 2436 852 2449 876
rect 2464 874 2479 876
rect 2276 838 2277 848
rect 2292 838 2305 848
rect 2319 838 2320 848
rect 2335 838 2348 848
rect 2363 838 2393 852
rect 2436 838 2479 852
rect 2503 849 2510 856
rect 2513 852 2580 876
rect 2612 876 2784 878
rect 2582 854 2610 858
rect 2612 854 2692 876
rect 2713 874 2728 876
rect 2582 852 2692 854
rect 2513 848 2692 852
rect 2486 838 2516 848
rect 2518 838 2671 848
rect 2679 838 2709 848
rect 2713 838 2743 852
rect 2771 838 2784 876
rect 2856 882 2891 890
rect 2856 856 2857 882
rect 2864 856 2891 882
rect 2799 838 2829 852
rect 2856 848 2891 856
rect 2893 882 2934 890
rect 2893 856 2908 882
rect 2915 856 2934 882
rect 2998 878 3060 890
rect 3072 878 3147 890
rect 3205 878 3280 890
rect 3292 878 3323 890
rect 3329 878 3364 890
rect 2998 876 3160 878
rect 2893 848 2934 856
rect 3016 852 3029 876
rect 3044 874 3059 876
rect 2856 838 2857 848
rect 2872 838 2885 848
rect 2899 838 2900 848
rect 2915 838 2928 848
rect 2943 838 2973 852
rect 3016 838 3059 852
rect 3083 849 3090 856
rect 3093 852 3160 876
rect 3192 876 3364 878
rect 3162 854 3190 858
rect 3192 854 3272 876
rect 3293 874 3308 876
rect 3162 852 3272 854
rect 3093 848 3272 852
rect 3066 838 3096 848
rect 3098 838 3251 848
rect 3259 838 3289 848
rect 3293 838 3323 852
rect 3351 838 3364 876
rect 3436 882 3471 890
rect 3436 856 3437 882
rect 3444 856 3471 882
rect 3379 838 3409 852
rect 3436 848 3471 856
rect 3473 882 3514 890
rect 3473 856 3488 882
rect 3495 856 3514 882
rect 3578 878 3640 890
rect 3652 878 3727 890
rect 3785 878 3860 890
rect 3872 878 3903 890
rect 3909 878 3944 890
rect 3578 876 3740 878
rect 3473 848 3514 856
rect 3596 852 3609 876
rect 3624 874 3639 876
rect 3436 838 3437 848
rect 3452 838 3465 848
rect 3479 838 3480 848
rect 3495 838 3508 848
rect 3523 838 3553 852
rect 3596 838 3639 852
rect 3663 849 3670 856
rect 3673 852 3740 876
rect 3772 876 3944 878
rect 3742 854 3770 858
rect 3772 854 3852 876
rect 3873 874 3888 876
rect 3742 852 3852 854
rect 3673 848 3852 852
rect 3646 838 3676 848
rect 3678 838 3831 848
rect 3839 838 3869 848
rect 3873 838 3903 852
rect 3931 838 3944 876
rect 4016 882 4051 890
rect 4016 856 4017 882
rect 4024 856 4051 882
rect 3959 838 3989 852
rect 4016 848 4051 856
rect 4053 882 4094 890
rect 4053 856 4068 882
rect 4075 856 4094 882
rect 4158 878 4220 890
rect 4232 878 4307 890
rect 4365 878 4440 890
rect 4452 878 4483 890
rect 4489 878 4524 890
rect 4158 876 4320 878
rect 4053 848 4094 856
rect 4176 852 4189 876
rect 4204 874 4219 876
rect 4016 838 4017 848
rect 4032 838 4045 848
rect 4059 838 4060 848
rect 4075 838 4088 848
rect 4103 838 4133 852
rect 4176 838 4219 852
rect 4243 849 4250 856
rect 4253 852 4320 876
rect 4352 876 4524 878
rect 4322 854 4350 858
rect 4352 854 4432 876
rect 4453 874 4468 876
rect 4322 852 4432 854
rect 4253 848 4432 852
rect 4226 838 4256 848
rect 4258 838 4411 848
rect 4419 838 4449 848
rect 4453 838 4483 852
rect 4511 838 4524 876
rect 4596 882 4631 890
rect 4596 856 4597 882
rect 4604 856 4631 882
rect 4539 838 4569 852
rect 4596 848 4631 856
rect 4596 838 4597 848
rect 4612 838 4625 848
rect -1 832 4625 838
rect 0 824 4625 832
rect 15 794 28 824
rect 43 806 73 824
rect 116 810 130 824
rect 166 810 386 824
rect 117 808 130 810
rect 83 796 98 808
rect 80 794 102 796
rect 107 794 137 808
rect 198 806 351 810
rect 180 794 372 806
rect 415 794 445 808
rect 451 794 464 824
rect 479 806 509 824
rect 552 794 565 824
rect 595 794 608 824
rect 623 806 653 824
rect 696 810 710 824
rect 746 810 966 824
rect 697 808 710 810
rect 663 796 678 808
rect 660 794 682 796
rect 687 794 717 808
rect 778 806 931 810
rect 760 794 952 806
rect 995 794 1025 808
rect 1031 794 1044 824
rect 1059 806 1089 824
rect 1132 794 1145 824
rect 1175 794 1188 824
rect 1203 806 1233 824
rect 1276 810 1290 824
rect 1326 810 1546 824
rect 1277 808 1290 810
rect 1243 796 1258 808
rect 1240 794 1262 796
rect 1267 794 1297 808
rect 1358 806 1511 810
rect 1340 794 1532 806
rect 1575 794 1605 808
rect 1611 794 1624 824
rect 1639 806 1669 824
rect 1712 794 1725 824
rect 1755 794 1768 824
rect 1783 806 1813 824
rect 1856 810 1870 824
rect 1906 810 2126 824
rect 1857 808 1870 810
rect 1823 796 1838 808
rect 1820 794 1842 796
rect 1847 794 1877 808
rect 1938 806 2091 810
rect 1920 794 2112 806
rect 2155 794 2185 808
rect 2191 794 2204 824
rect 2219 806 2249 824
rect 2292 794 2305 824
rect 2335 794 2348 824
rect 2363 806 2393 824
rect 2436 810 2450 824
rect 2486 810 2706 824
rect 2437 808 2450 810
rect 2403 796 2418 808
rect 2400 794 2422 796
rect 2427 794 2457 808
rect 2518 806 2671 810
rect 2500 794 2692 806
rect 2735 794 2765 808
rect 2771 794 2784 824
rect 2799 806 2829 824
rect 2872 794 2885 824
rect 2915 794 2928 824
rect 2943 806 2973 824
rect 3016 810 3030 824
rect 3066 810 3286 824
rect 3017 808 3030 810
rect 2983 796 2998 808
rect 2980 794 3002 796
rect 3007 794 3037 808
rect 3098 806 3251 810
rect 3080 794 3272 806
rect 3315 794 3345 808
rect 3351 794 3364 824
rect 3379 806 3409 824
rect 3452 794 3465 824
rect 3495 794 3508 824
rect 3523 806 3553 824
rect 3596 810 3610 824
rect 3646 810 3866 824
rect 3597 808 3610 810
rect 3563 796 3578 808
rect 3560 794 3582 796
rect 3587 794 3617 808
rect 3678 806 3831 810
rect 3660 794 3852 806
rect 3895 794 3925 808
rect 3931 794 3944 824
rect 3959 806 3989 824
rect 4032 794 4045 824
rect 4075 794 4088 824
rect 4103 806 4133 824
rect 4176 810 4190 824
rect 4226 810 4446 824
rect 4177 808 4190 810
rect 4143 796 4158 808
rect 4140 794 4162 796
rect 4167 794 4197 808
rect 4258 806 4411 810
rect 4240 794 4432 806
rect 4475 794 4505 808
rect 4511 794 4524 824
rect 4539 806 4569 824
rect 4612 794 4625 824
rect 0 780 4625 794
rect 15 676 28 780
rect 73 758 74 768
rect 89 758 102 768
rect 73 754 102 758
rect 107 754 137 780
rect 155 766 171 768
rect 243 766 296 780
rect 244 764 308 766
rect 351 764 366 780
rect 415 777 445 780
rect 415 774 451 777
rect 381 766 397 768
rect 155 754 170 758
rect 73 752 170 754
rect 198 752 366 764
rect 382 754 397 758
rect 415 755 454 774
rect 473 768 480 769
rect 479 761 480 768
rect 463 758 464 761
rect 479 758 492 761
rect 415 754 445 755
rect 454 754 460 755
rect 463 754 492 758
rect 382 753 492 754
rect 382 752 498 753
rect 57 744 108 752
rect 57 732 82 744
rect 89 732 108 744
rect 139 744 189 752
rect 139 736 155 744
rect 162 742 189 744
rect 198 742 419 752
rect 162 732 419 742
rect 448 744 498 752
rect 448 735 464 744
rect 57 724 108 732
rect 155 724 419 732
rect 445 732 464 735
rect 471 732 498 744
rect 445 724 498 732
rect 73 716 74 724
rect 89 716 102 724
rect 73 708 89 716
rect 70 701 89 704
rect 70 692 92 701
rect 43 682 92 692
rect 43 676 73 682
rect 92 677 97 682
rect 15 660 89 676
rect 107 668 137 724
rect 172 714 380 724
rect 415 720 460 724
rect 463 723 464 724
rect 479 723 492 724
rect 198 684 387 714
rect 213 681 387 684
rect 206 678 387 681
rect 15 658 28 660
rect 43 658 77 660
rect 15 642 89 658
rect 116 654 129 668
rect 144 654 160 670
rect 206 665 217 678
rect -1 620 0 636
rect 15 620 28 642
rect 43 620 73 642
rect 116 638 178 654
rect 206 647 217 663
rect 222 658 232 678
rect 242 658 256 678
rect 259 665 268 678
rect 284 665 293 678
rect 222 647 256 658
rect 259 647 268 663
rect 284 647 293 663
rect 300 658 310 678
rect 320 658 334 678
rect 335 665 346 678
rect 300 647 334 658
rect 335 647 346 663
rect 392 654 408 670
rect 415 668 445 720
rect 479 716 480 723
rect 464 708 480 716
rect 451 676 464 695
rect 479 676 509 692
rect 451 660 525 676
rect 451 658 464 660
rect 479 658 513 660
rect 116 636 129 638
rect 144 636 178 638
rect 116 620 178 636
rect 222 631 238 634
rect 300 631 330 642
rect 378 638 424 654
rect 451 642 525 658
rect 378 636 412 638
rect 377 620 424 636
rect 451 620 464 642
rect 479 620 509 642
rect 536 620 537 636
rect 552 620 565 780
rect 595 676 608 780
rect 653 758 654 768
rect 669 758 682 768
rect 653 754 682 758
rect 687 754 717 780
rect 735 766 751 768
rect 823 766 876 780
rect 824 764 888 766
rect 931 764 946 780
rect 995 777 1025 780
rect 995 774 1031 777
rect 961 766 977 768
rect 735 754 750 758
rect 653 752 750 754
rect 778 752 946 764
rect 962 754 977 758
rect 995 755 1034 774
rect 1053 768 1060 769
rect 1059 761 1060 768
rect 1043 758 1044 761
rect 1059 758 1072 761
rect 995 754 1025 755
rect 1034 754 1040 755
rect 1043 754 1072 758
rect 962 753 1072 754
rect 962 752 1078 753
rect 637 744 688 752
rect 637 732 662 744
rect 669 732 688 744
rect 719 744 769 752
rect 719 736 735 744
rect 742 742 769 744
rect 778 742 999 752
rect 742 732 999 742
rect 1028 744 1078 752
rect 1028 735 1044 744
rect 637 724 688 732
rect 735 724 999 732
rect 1025 732 1044 735
rect 1051 732 1078 744
rect 1025 724 1078 732
rect 653 716 654 724
rect 669 716 682 724
rect 653 708 669 716
rect 650 701 669 704
rect 650 692 672 701
rect 623 682 672 692
rect 623 676 653 682
rect 672 677 677 682
rect 595 660 669 676
rect 687 668 717 724
rect 752 714 960 724
rect 995 720 1040 724
rect 1043 723 1044 724
rect 1059 723 1072 724
rect 778 684 967 714
rect 793 681 967 684
rect 786 678 967 681
rect 595 658 608 660
rect 623 658 657 660
rect 595 642 669 658
rect 696 654 709 668
rect 724 654 740 670
rect 786 665 797 678
rect 579 620 580 636
rect 595 620 608 642
rect 623 620 653 642
rect 696 638 758 654
rect 786 647 797 663
rect 802 658 812 678
rect 822 658 836 678
rect 839 665 848 678
rect 864 665 873 678
rect 802 647 836 658
rect 839 647 848 663
rect 864 647 873 663
rect 880 658 890 678
rect 900 658 914 678
rect 915 665 926 678
rect 880 647 914 658
rect 915 647 926 663
rect 972 654 988 670
rect 995 668 1025 720
rect 1059 716 1060 723
rect 1044 708 1060 716
rect 1031 676 1044 695
rect 1059 676 1089 692
rect 1031 660 1105 676
rect 1031 658 1044 660
rect 1059 658 1093 660
rect 696 636 709 638
rect 724 636 758 638
rect 696 620 758 636
rect 802 631 818 634
rect 880 631 910 642
rect 958 638 1004 654
rect 1031 642 1105 658
rect 958 636 992 638
rect 957 620 1004 636
rect 1031 620 1044 642
rect 1059 620 1089 642
rect 1116 620 1117 636
rect 1132 620 1145 780
rect 1175 676 1188 780
rect 1233 758 1234 768
rect 1249 758 1262 768
rect 1233 754 1262 758
rect 1267 754 1297 780
rect 1315 766 1331 768
rect 1403 766 1456 780
rect 1404 764 1468 766
rect 1511 764 1526 780
rect 1575 777 1605 780
rect 1575 774 1611 777
rect 1541 766 1557 768
rect 1315 754 1330 758
rect 1233 752 1330 754
rect 1358 752 1526 764
rect 1542 754 1557 758
rect 1575 755 1614 774
rect 1633 768 1640 769
rect 1639 761 1640 768
rect 1623 758 1624 761
rect 1639 758 1652 761
rect 1575 754 1605 755
rect 1614 754 1620 755
rect 1623 754 1652 758
rect 1542 753 1652 754
rect 1542 752 1658 753
rect 1217 744 1268 752
rect 1217 732 1242 744
rect 1249 732 1268 744
rect 1299 744 1349 752
rect 1299 736 1315 744
rect 1322 742 1349 744
rect 1358 742 1579 752
rect 1322 732 1579 742
rect 1608 744 1658 752
rect 1608 735 1624 744
rect 1217 724 1268 732
rect 1315 724 1579 732
rect 1605 732 1624 735
rect 1631 732 1658 744
rect 1605 724 1658 732
rect 1233 716 1234 724
rect 1249 716 1262 724
rect 1233 708 1249 716
rect 1230 701 1249 704
rect 1230 692 1252 701
rect 1203 682 1252 692
rect 1203 676 1233 682
rect 1252 677 1257 682
rect 1175 660 1249 676
rect 1267 668 1297 724
rect 1332 714 1540 724
rect 1575 720 1620 724
rect 1623 723 1624 724
rect 1639 723 1652 724
rect 1358 684 1547 714
rect 1373 681 1547 684
rect 1366 678 1547 681
rect 1175 658 1188 660
rect 1203 658 1237 660
rect 1175 642 1249 658
rect 1276 654 1289 668
rect 1304 654 1320 670
rect 1366 665 1377 678
rect 1159 620 1160 636
rect 1175 620 1188 642
rect 1203 620 1233 642
rect 1276 638 1338 654
rect 1366 647 1377 663
rect 1382 658 1392 678
rect 1402 658 1416 678
rect 1419 665 1428 678
rect 1444 665 1453 678
rect 1382 647 1416 658
rect 1419 647 1428 663
rect 1444 647 1453 663
rect 1460 658 1470 678
rect 1480 658 1494 678
rect 1495 665 1506 678
rect 1460 647 1494 658
rect 1495 647 1506 663
rect 1552 654 1568 670
rect 1575 668 1605 720
rect 1639 716 1640 723
rect 1624 708 1640 716
rect 1611 676 1624 695
rect 1639 676 1669 692
rect 1611 660 1685 676
rect 1611 658 1624 660
rect 1639 658 1673 660
rect 1276 636 1289 638
rect 1304 636 1338 638
rect 1276 620 1338 636
rect 1382 631 1398 634
rect 1460 631 1490 642
rect 1538 638 1584 654
rect 1611 642 1685 658
rect 1538 636 1572 638
rect 1537 620 1584 636
rect 1611 620 1624 642
rect 1639 620 1669 642
rect 1696 620 1697 636
rect 1712 620 1725 780
rect 1755 676 1768 780
rect 1813 758 1814 768
rect 1829 758 1842 768
rect 1813 754 1842 758
rect 1847 754 1877 780
rect 1895 766 1911 768
rect 1983 766 2036 780
rect 1984 764 2048 766
rect 2091 764 2106 780
rect 2155 777 2185 780
rect 2155 774 2191 777
rect 2121 766 2137 768
rect 1895 754 1910 758
rect 1813 752 1910 754
rect 1938 752 2106 764
rect 2122 754 2137 758
rect 2155 755 2194 774
rect 2213 768 2220 769
rect 2219 761 2220 768
rect 2203 758 2204 761
rect 2219 758 2232 761
rect 2155 754 2185 755
rect 2194 754 2200 755
rect 2203 754 2232 758
rect 2122 753 2232 754
rect 2122 752 2238 753
rect 1797 744 1848 752
rect 1797 732 1822 744
rect 1829 732 1848 744
rect 1879 744 1929 752
rect 1879 736 1895 744
rect 1902 742 1929 744
rect 1938 742 2159 752
rect 1902 732 2159 742
rect 2188 744 2238 752
rect 2188 735 2204 744
rect 1797 724 1848 732
rect 1895 724 2159 732
rect 2185 732 2204 735
rect 2211 732 2238 744
rect 2185 724 2238 732
rect 1813 716 1814 724
rect 1829 716 1842 724
rect 1813 708 1829 716
rect 1810 701 1829 704
rect 1810 692 1832 701
rect 1783 682 1832 692
rect 1783 676 1813 682
rect 1832 677 1837 682
rect 1755 660 1829 676
rect 1847 668 1877 724
rect 1912 714 2120 724
rect 2155 720 2200 724
rect 2203 723 2204 724
rect 2219 723 2232 724
rect 1938 684 2127 714
rect 1953 681 2127 684
rect 1946 678 2127 681
rect 1755 658 1768 660
rect 1783 658 1817 660
rect 1755 642 1829 658
rect 1856 654 1869 668
rect 1884 654 1900 670
rect 1946 665 1957 678
rect 1739 620 1740 636
rect 1755 620 1768 642
rect 1783 620 1813 642
rect 1856 638 1918 654
rect 1946 647 1957 663
rect 1962 658 1972 678
rect 1982 658 1996 678
rect 1999 665 2008 678
rect 2024 665 2033 678
rect 1962 647 1996 658
rect 1999 647 2008 663
rect 2024 647 2033 663
rect 2040 658 2050 678
rect 2060 658 2074 678
rect 2075 665 2086 678
rect 2040 647 2074 658
rect 2075 647 2086 663
rect 2132 654 2148 670
rect 2155 668 2185 720
rect 2219 716 2220 723
rect 2204 708 2220 716
rect 2191 676 2204 695
rect 2219 676 2249 692
rect 2191 660 2265 676
rect 2191 658 2204 660
rect 2219 658 2253 660
rect 1856 636 1869 638
rect 1884 636 1918 638
rect 1856 620 1918 636
rect 1962 631 1978 634
rect 2040 631 2070 642
rect 2118 638 2164 654
rect 2191 642 2265 658
rect 2118 636 2152 638
rect 2117 620 2164 636
rect 2191 620 2204 642
rect 2219 620 2249 642
rect 2276 620 2277 636
rect 2292 620 2305 780
rect 2335 676 2348 780
rect 2393 758 2394 768
rect 2409 758 2422 768
rect 2393 754 2422 758
rect 2427 754 2457 780
rect 2475 766 2491 768
rect 2563 766 2616 780
rect 2564 764 2628 766
rect 2671 764 2686 780
rect 2735 777 2765 780
rect 2735 774 2771 777
rect 2701 766 2717 768
rect 2475 754 2490 758
rect 2393 752 2490 754
rect 2518 752 2686 764
rect 2702 754 2717 758
rect 2735 755 2774 774
rect 2793 768 2800 769
rect 2799 761 2800 768
rect 2783 758 2784 761
rect 2799 758 2812 761
rect 2735 754 2765 755
rect 2774 754 2780 755
rect 2783 754 2812 758
rect 2702 753 2812 754
rect 2702 752 2818 753
rect 2377 744 2428 752
rect 2377 732 2402 744
rect 2409 732 2428 744
rect 2459 744 2509 752
rect 2459 736 2475 744
rect 2482 742 2509 744
rect 2518 742 2739 752
rect 2482 732 2739 742
rect 2768 744 2818 752
rect 2768 735 2784 744
rect 2377 724 2428 732
rect 2475 724 2739 732
rect 2765 732 2784 735
rect 2791 732 2818 744
rect 2765 724 2818 732
rect 2393 716 2394 724
rect 2409 716 2422 724
rect 2393 708 2409 716
rect 2390 701 2409 704
rect 2390 692 2412 701
rect 2363 682 2412 692
rect 2363 676 2393 682
rect 2412 677 2417 682
rect 2335 660 2409 676
rect 2427 668 2457 724
rect 2492 714 2700 724
rect 2735 720 2780 724
rect 2783 723 2784 724
rect 2799 723 2812 724
rect 2518 684 2707 714
rect 2533 681 2707 684
rect 2526 678 2707 681
rect 2335 658 2348 660
rect 2363 658 2397 660
rect 2335 642 2409 658
rect 2436 654 2449 668
rect 2464 654 2480 670
rect 2526 665 2537 678
rect 2319 620 2320 636
rect 2335 620 2348 642
rect 2363 620 2393 642
rect 2436 638 2498 654
rect 2526 647 2537 663
rect 2542 658 2552 678
rect 2562 658 2576 678
rect 2579 665 2588 678
rect 2604 665 2613 678
rect 2542 647 2576 658
rect 2579 647 2588 663
rect 2604 647 2613 663
rect 2620 658 2630 678
rect 2640 658 2654 678
rect 2655 665 2666 678
rect 2620 647 2654 658
rect 2655 647 2666 663
rect 2712 654 2728 670
rect 2735 668 2765 720
rect 2799 716 2800 723
rect 2784 708 2800 716
rect 2771 676 2784 695
rect 2799 676 2829 692
rect 2771 660 2845 676
rect 2771 658 2784 660
rect 2799 658 2833 660
rect 2436 636 2449 638
rect 2464 636 2498 638
rect 2436 620 2498 636
rect 2542 631 2558 634
rect 2620 631 2650 642
rect 2698 638 2744 654
rect 2771 642 2845 658
rect 2698 636 2732 638
rect 2697 620 2744 636
rect 2771 620 2784 642
rect 2799 620 2829 642
rect 2856 620 2857 636
rect 2872 620 2885 780
rect 2915 676 2928 780
rect 2973 758 2974 768
rect 2989 758 3002 768
rect 2973 754 3002 758
rect 3007 754 3037 780
rect 3055 766 3071 768
rect 3143 766 3196 780
rect 3144 764 3208 766
rect 3251 764 3266 780
rect 3315 777 3345 780
rect 3315 774 3351 777
rect 3281 766 3297 768
rect 3055 754 3070 758
rect 2973 752 3070 754
rect 3098 752 3266 764
rect 3282 754 3297 758
rect 3315 755 3354 774
rect 3373 768 3380 769
rect 3379 761 3380 768
rect 3363 758 3364 761
rect 3379 758 3392 761
rect 3315 754 3345 755
rect 3354 754 3360 755
rect 3363 754 3392 758
rect 3282 753 3392 754
rect 3282 752 3398 753
rect 2957 744 3008 752
rect 2957 732 2982 744
rect 2989 732 3008 744
rect 3039 744 3089 752
rect 3039 736 3055 744
rect 3062 742 3089 744
rect 3098 742 3319 752
rect 3062 732 3319 742
rect 3348 744 3398 752
rect 3348 735 3364 744
rect 2957 724 3008 732
rect 3055 724 3319 732
rect 3345 732 3364 735
rect 3371 732 3398 744
rect 3345 724 3398 732
rect 2973 716 2974 724
rect 2989 716 3002 724
rect 2973 708 2989 716
rect 2970 701 2989 704
rect 2970 692 2992 701
rect 2943 682 2992 692
rect 2943 676 2973 682
rect 2992 677 2997 682
rect 2915 660 2989 676
rect 3007 668 3037 724
rect 3072 714 3280 724
rect 3315 720 3360 724
rect 3363 723 3364 724
rect 3379 723 3392 724
rect 3098 684 3287 714
rect 3113 681 3287 684
rect 3106 678 3287 681
rect 2915 658 2928 660
rect 2943 658 2977 660
rect 2915 642 2989 658
rect 3016 654 3029 668
rect 3044 654 3060 670
rect 3106 665 3117 678
rect 2899 620 2900 636
rect 2915 620 2928 642
rect 2943 620 2973 642
rect 3016 638 3078 654
rect 3106 647 3117 663
rect 3122 658 3132 678
rect 3142 658 3156 678
rect 3159 665 3168 678
rect 3184 665 3193 678
rect 3122 647 3156 658
rect 3159 647 3168 663
rect 3184 647 3193 663
rect 3200 658 3210 678
rect 3220 658 3234 678
rect 3235 665 3246 678
rect 3200 647 3234 658
rect 3235 647 3246 663
rect 3292 654 3308 670
rect 3315 668 3345 720
rect 3379 716 3380 723
rect 3364 708 3380 716
rect 3351 676 3364 695
rect 3379 676 3409 692
rect 3351 660 3425 676
rect 3351 658 3364 660
rect 3379 658 3413 660
rect 3016 636 3029 638
rect 3044 636 3078 638
rect 3016 620 3078 636
rect 3122 631 3138 634
rect 3200 631 3230 642
rect 3278 638 3324 654
rect 3351 642 3425 658
rect 3278 636 3312 638
rect 3277 620 3324 636
rect 3351 620 3364 642
rect 3379 620 3409 642
rect 3436 620 3437 636
rect 3452 620 3465 780
rect 3495 676 3508 780
rect 3553 758 3554 768
rect 3569 758 3582 768
rect 3553 754 3582 758
rect 3587 754 3617 780
rect 3635 766 3651 768
rect 3723 766 3776 780
rect 3724 764 3788 766
rect 3831 764 3846 780
rect 3895 777 3925 780
rect 3895 774 3931 777
rect 3861 766 3877 768
rect 3635 754 3650 758
rect 3553 752 3650 754
rect 3678 752 3846 764
rect 3862 754 3877 758
rect 3895 755 3934 774
rect 3953 768 3960 769
rect 3959 761 3960 768
rect 3943 758 3944 761
rect 3959 758 3972 761
rect 3895 754 3925 755
rect 3934 754 3940 755
rect 3943 754 3972 758
rect 3862 753 3972 754
rect 3862 752 3978 753
rect 3537 744 3588 752
rect 3537 732 3562 744
rect 3569 732 3588 744
rect 3619 744 3669 752
rect 3619 736 3635 744
rect 3642 742 3669 744
rect 3678 742 3899 752
rect 3642 732 3899 742
rect 3928 744 3978 752
rect 3928 735 3944 744
rect 3537 724 3588 732
rect 3635 724 3899 732
rect 3925 732 3944 735
rect 3951 732 3978 744
rect 3925 724 3978 732
rect 3553 716 3554 724
rect 3569 716 3582 724
rect 3553 708 3569 716
rect 3550 701 3569 704
rect 3550 692 3572 701
rect 3523 682 3572 692
rect 3523 676 3553 682
rect 3572 677 3577 682
rect 3495 660 3569 676
rect 3587 668 3617 724
rect 3652 714 3860 724
rect 3895 720 3940 724
rect 3943 723 3944 724
rect 3959 723 3972 724
rect 3678 684 3867 714
rect 3693 681 3867 684
rect 3686 678 3867 681
rect 3495 658 3508 660
rect 3523 658 3557 660
rect 3495 642 3569 658
rect 3596 654 3609 668
rect 3624 654 3640 670
rect 3686 665 3697 678
rect 3479 620 3480 636
rect 3495 620 3508 642
rect 3523 620 3553 642
rect 3596 638 3658 654
rect 3686 647 3697 663
rect 3702 658 3712 678
rect 3722 658 3736 678
rect 3739 665 3748 678
rect 3764 665 3773 678
rect 3702 647 3736 658
rect 3739 647 3748 663
rect 3764 647 3773 663
rect 3780 658 3790 678
rect 3800 658 3814 678
rect 3815 665 3826 678
rect 3780 647 3814 658
rect 3815 647 3826 663
rect 3872 654 3888 670
rect 3895 668 3925 720
rect 3959 716 3960 723
rect 3944 708 3960 716
rect 3931 676 3944 695
rect 3959 676 3989 692
rect 3931 660 4005 676
rect 3931 658 3944 660
rect 3959 658 3993 660
rect 3596 636 3609 638
rect 3624 636 3658 638
rect 3596 620 3658 636
rect 3702 631 3718 634
rect 3780 631 3810 642
rect 3858 638 3904 654
rect 3931 642 4005 658
rect 3858 636 3892 638
rect 3857 620 3904 636
rect 3931 620 3944 642
rect 3959 620 3989 642
rect 4016 620 4017 636
rect 4032 620 4045 780
rect 4075 676 4088 780
rect 4133 758 4134 768
rect 4149 758 4162 768
rect 4133 754 4162 758
rect 4167 754 4197 780
rect 4215 766 4231 768
rect 4303 766 4356 780
rect 4304 764 4368 766
rect 4411 764 4426 780
rect 4475 777 4505 780
rect 4475 774 4511 777
rect 4441 766 4457 768
rect 4215 754 4230 758
rect 4133 752 4230 754
rect 4258 752 4426 764
rect 4442 754 4457 758
rect 4475 755 4514 774
rect 4533 768 4540 769
rect 4539 761 4540 768
rect 4523 758 4524 761
rect 4539 758 4552 761
rect 4475 754 4505 755
rect 4514 754 4520 755
rect 4523 754 4552 758
rect 4442 753 4552 754
rect 4442 752 4558 753
rect 4117 744 4168 752
rect 4117 732 4142 744
rect 4149 732 4168 744
rect 4199 744 4249 752
rect 4199 736 4215 744
rect 4222 742 4249 744
rect 4258 742 4479 752
rect 4222 732 4479 742
rect 4508 744 4558 752
rect 4508 735 4524 744
rect 4117 724 4168 732
rect 4215 724 4479 732
rect 4505 732 4524 735
rect 4531 732 4558 744
rect 4505 724 4558 732
rect 4133 716 4134 724
rect 4149 716 4162 724
rect 4133 708 4149 716
rect 4130 701 4149 704
rect 4130 692 4152 701
rect 4103 682 4152 692
rect 4103 676 4133 682
rect 4152 677 4157 682
rect 4075 660 4149 676
rect 4167 668 4197 724
rect 4232 714 4440 724
rect 4475 720 4520 724
rect 4523 723 4524 724
rect 4539 723 4552 724
rect 4258 684 4447 714
rect 4273 681 4447 684
rect 4266 678 4447 681
rect 4075 658 4088 660
rect 4103 658 4137 660
rect 4075 642 4149 658
rect 4176 654 4189 668
rect 4204 654 4220 670
rect 4266 665 4277 678
rect 4059 620 4060 636
rect 4075 620 4088 642
rect 4103 620 4133 642
rect 4176 638 4238 654
rect 4266 647 4277 663
rect 4282 658 4292 678
rect 4302 658 4316 678
rect 4319 665 4328 678
rect 4344 665 4353 678
rect 4282 647 4316 658
rect 4319 647 4328 663
rect 4344 647 4353 663
rect 4360 658 4370 678
rect 4380 658 4394 678
rect 4395 665 4406 678
rect 4360 647 4394 658
rect 4395 647 4406 663
rect 4452 654 4468 670
rect 4475 668 4505 720
rect 4539 716 4540 723
rect 4524 708 4540 716
rect 4511 676 4524 695
rect 4539 676 4569 692
rect 4511 660 4585 676
rect 4511 658 4524 660
rect 4539 658 4573 660
rect 4176 636 4189 638
rect 4204 636 4238 638
rect 4176 620 4238 636
rect 4282 631 4298 634
rect 4360 631 4390 642
rect 4438 638 4484 654
rect 4511 642 4585 658
rect 4438 636 4472 638
rect 4437 620 4484 636
rect 4511 620 4524 642
rect 4539 620 4569 642
rect 4596 620 4597 636
rect 4612 620 4625 780
rect -7 612 34 620
rect -7 586 8 612
rect 15 586 34 612
rect 98 608 160 620
rect 172 608 247 620
rect 305 608 380 620
rect 392 608 423 620
rect 429 608 464 620
rect 98 606 260 608
rect -7 578 34 586
rect 116 582 129 606
rect 144 604 159 606
rect -1 568 0 578
rect 15 568 28 578
rect 43 568 73 582
rect 116 568 159 582
rect 183 579 190 586
rect 193 582 260 606
rect 292 606 464 608
rect 262 584 290 588
rect 292 584 372 606
rect 393 604 408 606
rect 262 582 372 584
rect 193 578 372 582
rect 166 568 196 578
rect 198 568 351 578
rect 359 568 389 578
rect 393 568 423 582
rect 451 568 464 606
rect 536 612 571 620
rect 536 586 537 612
rect 544 586 571 612
rect 479 568 509 582
rect 536 578 571 586
rect 573 612 614 620
rect 573 586 588 612
rect 595 586 614 612
rect 678 608 740 620
rect 752 608 827 620
rect 885 608 960 620
rect 972 608 1003 620
rect 1009 608 1044 620
rect 678 606 840 608
rect 573 578 614 586
rect 696 582 709 606
rect 724 604 739 606
rect 536 568 537 578
rect 552 568 565 578
rect 579 568 580 578
rect 595 568 608 578
rect 623 568 653 582
rect 696 568 739 582
rect 763 579 770 586
rect 773 582 840 606
rect 872 606 1044 608
rect 842 584 870 588
rect 872 584 952 606
rect 973 604 988 606
rect 842 582 952 584
rect 773 578 952 582
rect 746 568 776 578
rect 778 568 931 578
rect 939 568 969 578
rect 973 568 1003 582
rect 1031 568 1044 606
rect 1116 612 1151 620
rect 1116 586 1117 612
rect 1124 586 1151 612
rect 1059 568 1089 582
rect 1116 578 1151 586
rect 1153 612 1194 620
rect 1153 586 1168 612
rect 1175 586 1194 612
rect 1258 608 1320 620
rect 1332 608 1407 620
rect 1465 608 1540 620
rect 1552 608 1583 620
rect 1589 608 1624 620
rect 1258 606 1420 608
rect 1153 578 1194 586
rect 1276 582 1289 606
rect 1304 604 1319 606
rect 1116 568 1117 578
rect 1132 568 1145 578
rect 1159 568 1160 578
rect 1175 568 1188 578
rect 1203 568 1233 582
rect 1276 568 1319 582
rect 1343 579 1350 586
rect 1353 582 1420 606
rect 1452 606 1624 608
rect 1422 584 1450 588
rect 1452 584 1532 606
rect 1553 604 1568 606
rect 1422 582 1532 584
rect 1353 578 1532 582
rect 1326 568 1356 578
rect 1358 568 1511 578
rect 1519 568 1549 578
rect 1553 568 1583 582
rect 1611 568 1624 606
rect 1696 612 1731 620
rect 1696 586 1697 612
rect 1704 586 1731 612
rect 1639 568 1669 582
rect 1696 578 1731 586
rect 1733 612 1774 620
rect 1733 586 1748 612
rect 1755 586 1774 612
rect 1838 608 1900 620
rect 1912 608 1987 620
rect 2045 608 2120 620
rect 2132 608 2163 620
rect 2169 608 2204 620
rect 1838 606 2000 608
rect 1733 578 1774 586
rect 1856 582 1869 606
rect 1884 604 1899 606
rect 1696 568 1697 578
rect 1712 568 1725 578
rect 1739 568 1740 578
rect 1755 568 1768 578
rect 1783 568 1813 582
rect 1856 568 1899 582
rect 1923 579 1930 586
rect 1933 582 2000 606
rect 2032 606 2204 608
rect 2002 584 2030 588
rect 2032 584 2112 606
rect 2133 604 2148 606
rect 2002 582 2112 584
rect 1933 578 2112 582
rect 1906 568 1936 578
rect 1938 568 2091 578
rect 2099 568 2129 578
rect 2133 568 2163 582
rect 2191 568 2204 606
rect 2276 612 2311 620
rect 2276 586 2277 612
rect 2284 586 2311 612
rect 2219 568 2249 582
rect 2276 578 2311 586
rect 2313 612 2354 620
rect 2313 586 2328 612
rect 2335 586 2354 612
rect 2418 608 2480 620
rect 2492 608 2567 620
rect 2625 608 2700 620
rect 2712 608 2743 620
rect 2749 608 2784 620
rect 2418 606 2580 608
rect 2313 578 2354 586
rect 2436 582 2449 606
rect 2464 604 2479 606
rect 2276 568 2277 578
rect 2292 568 2305 578
rect 2319 568 2320 578
rect 2335 568 2348 578
rect 2363 568 2393 582
rect 2436 568 2479 582
rect 2503 579 2510 586
rect 2513 582 2580 606
rect 2612 606 2784 608
rect 2582 584 2610 588
rect 2612 584 2692 606
rect 2713 604 2728 606
rect 2582 582 2692 584
rect 2513 578 2692 582
rect 2486 568 2516 578
rect 2518 568 2671 578
rect 2679 568 2709 578
rect 2713 568 2743 582
rect 2771 568 2784 606
rect 2856 612 2891 620
rect 2856 586 2857 612
rect 2864 586 2891 612
rect 2799 568 2829 582
rect 2856 578 2891 586
rect 2893 612 2934 620
rect 2893 586 2908 612
rect 2915 586 2934 612
rect 2998 608 3060 620
rect 3072 608 3147 620
rect 3205 608 3280 620
rect 3292 608 3323 620
rect 3329 608 3364 620
rect 2998 606 3160 608
rect 2893 578 2934 586
rect 3016 582 3029 606
rect 3044 604 3059 606
rect 2856 568 2857 578
rect 2872 568 2885 578
rect 2899 568 2900 578
rect 2915 568 2928 578
rect 2943 568 2973 582
rect 3016 568 3059 582
rect 3083 579 3090 586
rect 3093 582 3160 606
rect 3192 606 3364 608
rect 3162 584 3190 588
rect 3192 584 3272 606
rect 3293 604 3308 606
rect 3162 582 3272 584
rect 3093 578 3272 582
rect 3066 568 3096 578
rect 3098 568 3251 578
rect 3259 568 3289 578
rect 3293 568 3323 582
rect 3351 568 3364 606
rect 3436 612 3471 620
rect 3436 586 3437 612
rect 3444 586 3471 612
rect 3379 568 3409 582
rect 3436 578 3471 586
rect 3473 612 3514 620
rect 3473 586 3488 612
rect 3495 586 3514 612
rect 3578 608 3640 620
rect 3652 608 3727 620
rect 3785 608 3860 620
rect 3872 608 3903 620
rect 3909 608 3944 620
rect 3578 606 3740 608
rect 3473 578 3514 586
rect 3596 582 3609 606
rect 3624 604 3639 606
rect 3436 568 3437 578
rect 3452 568 3465 578
rect 3479 568 3480 578
rect 3495 568 3508 578
rect 3523 568 3553 582
rect 3596 568 3639 582
rect 3663 579 3670 586
rect 3673 582 3740 606
rect 3772 606 3944 608
rect 3742 584 3770 588
rect 3772 584 3852 606
rect 3873 604 3888 606
rect 3742 582 3852 584
rect 3673 578 3852 582
rect 3646 568 3676 578
rect 3678 568 3831 578
rect 3839 568 3869 578
rect 3873 568 3903 582
rect 3931 568 3944 606
rect 4016 612 4051 620
rect 4016 586 4017 612
rect 4024 586 4051 612
rect 3959 568 3989 582
rect 4016 578 4051 586
rect 4053 612 4094 620
rect 4053 586 4068 612
rect 4075 586 4094 612
rect 4158 608 4220 620
rect 4232 608 4307 620
rect 4365 608 4440 620
rect 4452 608 4483 620
rect 4489 608 4524 620
rect 4158 606 4320 608
rect 4053 578 4094 586
rect 4176 582 4189 606
rect 4204 604 4219 606
rect 4016 568 4017 578
rect 4032 568 4045 578
rect 4059 568 4060 578
rect 4075 568 4088 578
rect 4103 568 4133 582
rect 4176 568 4219 582
rect 4243 579 4250 586
rect 4253 582 4320 606
rect 4352 606 4524 608
rect 4322 584 4350 588
rect 4352 584 4432 606
rect 4453 604 4468 606
rect 4322 582 4432 584
rect 4253 578 4432 582
rect 4226 568 4256 578
rect 4258 568 4411 578
rect 4419 568 4449 578
rect 4453 568 4483 582
rect 4511 568 4524 606
rect 4596 612 4631 620
rect 4596 586 4597 612
rect 4604 586 4631 612
rect 4539 568 4569 582
rect 4596 578 4631 586
rect 4596 568 4597 578
rect 4612 568 4625 578
rect -1 562 4625 568
rect 0 554 4625 562
rect 15 524 28 554
rect 43 536 73 554
rect 116 540 130 554
rect 166 540 386 554
rect 117 538 130 540
rect 83 526 98 538
rect 80 524 102 526
rect 107 524 137 538
rect 198 536 351 540
rect 180 524 372 536
rect 415 524 445 538
rect 451 524 464 554
rect 479 536 509 554
rect 552 524 565 554
rect 595 524 608 554
rect 623 536 653 554
rect 696 540 710 554
rect 746 540 966 554
rect 697 538 710 540
rect 663 526 678 538
rect 660 524 682 526
rect 687 524 717 538
rect 778 536 931 540
rect 760 524 952 536
rect 995 524 1025 538
rect 1031 524 1044 554
rect 1059 536 1089 554
rect 1132 524 1145 554
rect 1175 524 1188 554
rect 1203 536 1233 554
rect 1276 540 1290 554
rect 1326 540 1546 554
rect 1277 538 1290 540
rect 1243 526 1258 538
rect 1240 524 1262 526
rect 1267 524 1297 538
rect 1358 536 1511 540
rect 1340 524 1532 536
rect 1575 524 1605 538
rect 1611 524 1624 554
rect 1639 536 1669 554
rect 1712 524 1725 554
rect 1755 524 1768 554
rect 1783 536 1813 554
rect 1856 540 1870 554
rect 1906 540 2126 554
rect 1857 538 1870 540
rect 1823 526 1838 538
rect 1820 524 1842 526
rect 1847 524 1877 538
rect 1938 536 2091 540
rect 1920 524 2112 536
rect 2155 524 2185 538
rect 2191 524 2204 554
rect 2219 536 2249 554
rect 2292 524 2305 554
rect 2335 524 2348 554
rect 2363 536 2393 554
rect 2436 540 2450 554
rect 2486 540 2706 554
rect 2437 538 2450 540
rect 2403 526 2418 538
rect 2400 524 2422 526
rect 2427 524 2457 538
rect 2518 536 2671 540
rect 2500 524 2692 536
rect 2735 524 2765 538
rect 2771 524 2784 554
rect 2799 536 2829 554
rect 2872 524 2885 554
rect 2915 524 2928 554
rect 2943 536 2973 554
rect 3016 540 3030 554
rect 3066 540 3286 554
rect 3017 538 3030 540
rect 2983 526 2998 538
rect 2980 524 3002 526
rect 3007 524 3037 538
rect 3098 536 3251 540
rect 3080 524 3272 536
rect 3315 524 3345 538
rect 3351 524 3364 554
rect 3379 536 3409 554
rect 3452 524 3465 554
rect 3495 524 3508 554
rect 3523 536 3553 554
rect 3596 540 3610 554
rect 3646 540 3866 554
rect 3597 538 3610 540
rect 3563 526 3578 538
rect 3560 524 3582 526
rect 3587 524 3617 538
rect 3678 536 3831 540
rect 3660 524 3852 536
rect 3895 524 3925 538
rect 3931 524 3944 554
rect 3959 536 3989 554
rect 4032 524 4045 554
rect 4075 524 4088 554
rect 4103 536 4133 554
rect 4176 540 4190 554
rect 4226 540 4446 554
rect 4177 538 4190 540
rect 4143 526 4158 538
rect 4140 524 4162 526
rect 4167 524 4197 538
rect 4258 536 4411 540
rect 4240 524 4432 536
rect 4475 524 4505 538
rect 4511 524 4524 554
rect 4539 536 4569 554
rect 4612 524 4625 554
rect 0 510 4625 524
rect 15 406 28 510
rect 73 488 74 498
rect 89 488 102 498
rect 73 484 102 488
rect 107 484 137 510
rect 155 496 171 498
rect 243 496 296 510
rect 244 494 308 496
rect 351 494 366 510
rect 415 507 445 510
rect 415 504 451 507
rect 381 496 397 498
rect 155 484 170 488
rect 73 482 170 484
rect 198 482 366 494
rect 382 484 397 488
rect 415 485 454 504
rect 473 498 480 499
rect 479 491 480 498
rect 463 488 464 491
rect 479 488 492 491
rect 415 484 445 485
rect 454 484 460 485
rect 463 484 492 488
rect 382 483 492 484
rect 382 482 498 483
rect 57 474 108 482
rect 57 462 82 474
rect 89 462 108 474
rect 139 474 189 482
rect 139 466 155 474
rect 162 472 189 474
rect 198 472 419 482
rect 162 462 419 472
rect 448 474 498 482
rect 448 465 464 474
rect 57 454 108 462
rect 155 454 419 462
rect 445 462 464 465
rect 471 462 498 474
rect 445 454 498 462
rect 73 446 74 454
rect 89 446 102 454
rect 73 438 89 446
rect 70 431 89 434
rect 70 422 92 431
rect 43 412 92 422
rect 43 406 73 412
rect 92 407 97 412
rect 15 390 89 406
rect 107 398 137 454
rect 172 444 380 454
rect 415 450 460 454
rect 463 453 464 454
rect 479 453 492 454
rect 198 414 387 444
rect 213 411 387 414
rect 206 408 387 411
rect 15 388 28 390
rect 43 388 77 390
rect 15 372 89 388
rect 116 384 129 398
rect 144 384 160 400
rect 206 395 217 408
rect -1 350 0 366
rect 15 350 28 372
rect 43 350 73 372
rect 116 368 178 384
rect 206 377 217 393
rect 222 388 232 408
rect 242 388 256 408
rect 259 395 268 408
rect 284 395 293 408
rect 222 377 256 388
rect 259 377 268 393
rect 284 377 293 393
rect 300 388 310 408
rect 320 388 334 408
rect 335 395 346 408
rect 300 377 334 388
rect 335 377 346 393
rect 392 384 408 400
rect 415 398 445 450
rect 479 446 480 453
rect 464 438 480 446
rect 451 406 464 425
rect 479 406 509 422
rect 451 390 525 406
rect 451 388 464 390
rect 479 388 513 390
rect 116 366 129 368
rect 144 366 178 368
rect 116 350 178 366
rect 222 361 238 364
rect 300 361 330 372
rect 378 368 424 384
rect 451 372 525 388
rect 378 366 412 368
rect 377 350 424 366
rect 451 350 464 372
rect 479 350 509 372
rect 536 350 537 366
rect 552 350 565 510
rect 595 406 608 510
rect 653 488 654 498
rect 669 488 682 498
rect 653 484 682 488
rect 687 484 717 510
rect 735 496 751 498
rect 823 496 876 510
rect 824 494 888 496
rect 931 494 946 510
rect 995 507 1025 510
rect 995 504 1031 507
rect 961 496 977 498
rect 735 484 750 488
rect 653 482 750 484
rect 778 482 946 494
rect 962 484 977 488
rect 995 485 1034 504
rect 1053 498 1060 499
rect 1059 491 1060 498
rect 1043 488 1044 491
rect 1059 488 1072 491
rect 995 484 1025 485
rect 1034 484 1040 485
rect 1043 484 1072 488
rect 962 483 1072 484
rect 962 482 1078 483
rect 637 474 688 482
rect 637 462 662 474
rect 669 462 688 474
rect 719 474 769 482
rect 719 466 735 474
rect 742 472 769 474
rect 778 472 999 482
rect 742 462 999 472
rect 1028 474 1078 482
rect 1028 465 1044 474
rect 637 454 688 462
rect 735 454 999 462
rect 1025 462 1044 465
rect 1051 462 1078 474
rect 1025 454 1078 462
rect 653 446 654 454
rect 669 446 682 454
rect 653 438 669 446
rect 650 431 669 434
rect 650 422 672 431
rect 623 412 672 422
rect 623 406 653 412
rect 672 407 677 412
rect 595 390 669 406
rect 687 398 717 454
rect 752 444 960 454
rect 995 450 1040 454
rect 1043 453 1044 454
rect 1059 453 1072 454
rect 778 414 967 444
rect 793 411 967 414
rect 786 408 967 411
rect 595 388 608 390
rect 623 388 657 390
rect 595 372 669 388
rect 696 384 709 398
rect 724 384 740 400
rect 786 395 797 408
rect 579 350 580 366
rect 595 350 608 372
rect 623 350 653 372
rect 696 368 758 384
rect 786 377 797 393
rect 802 388 812 408
rect 822 388 836 408
rect 839 395 848 408
rect 864 395 873 408
rect 802 377 836 388
rect 839 377 848 393
rect 864 377 873 393
rect 880 388 890 408
rect 900 388 914 408
rect 915 395 926 408
rect 880 377 914 388
rect 915 377 926 393
rect 972 384 988 400
rect 995 398 1025 450
rect 1059 446 1060 453
rect 1044 438 1060 446
rect 1031 406 1044 425
rect 1059 406 1089 422
rect 1031 390 1105 406
rect 1031 388 1044 390
rect 1059 388 1093 390
rect 696 366 709 368
rect 724 366 758 368
rect 696 350 758 366
rect 802 361 818 364
rect 880 361 910 372
rect 958 368 1004 384
rect 1031 372 1105 388
rect 958 366 992 368
rect 957 350 1004 366
rect 1031 350 1044 372
rect 1059 350 1089 372
rect 1116 350 1117 366
rect 1132 350 1145 510
rect 1175 406 1188 510
rect 1233 488 1234 498
rect 1249 488 1262 498
rect 1233 484 1262 488
rect 1267 484 1297 510
rect 1315 496 1331 498
rect 1403 496 1456 510
rect 1404 494 1468 496
rect 1511 494 1526 510
rect 1575 507 1605 510
rect 1575 504 1611 507
rect 1541 496 1557 498
rect 1315 484 1330 488
rect 1233 482 1330 484
rect 1358 482 1526 494
rect 1542 484 1557 488
rect 1575 485 1614 504
rect 1633 498 1640 499
rect 1639 491 1640 498
rect 1623 488 1624 491
rect 1639 488 1652 491
rect 1575 484 1605 485
rect 1614 484 1620 485
rect 1623 484 1652 488
rect 1542 483 1652 484
rect 1542 482 1658 483
rect 1217 474 1268 482
rect 1217 462 1242 474
rect 1249 462 1268 474
rect 1299 474 1349 482
rect 1299 466 1315 474
rect 1322 472 1349 474
rect 1358 472 1579 482
rect 1322 462 1579 472
rect 1608 474 1658 482
rect 1608 465 1624 474
rect 1217 454 1268 462
rect 1315 454 1579 462
rect 1605 462 1624 465
rect 1631 462 1658 474
rect 1605 454 1658 462
rect 1233 446 1234 454
rect 1249 446 1262 454
rect 1233 438 1249 446
rect 1230 431 1249 434
rect 1230 422 1252 431
rect 1203 412 1252 422
rect 1203 406 1233 412
rect 1252 407 1257 412
rect 1175 390 1249 406
rect 1267 398 1297 454
rect 1332 444 1540 454
rect 1575 450 1620 454
rect 1623 453 1624 454
rect 1639 453 1652 454
rect 1358 414 1547 444
rect 1373 411 1547 414
rect 1366 408 1547 411
rect 1175 388 1188 390
rect 1203 388 1237 390
rect 1175 372 1249 388
rect 1276 384 1289 398
rect 1304 384 1320 400
rect 1366 395 1377 408
rect 1159 350 1160 366
rect 1175 350 1188 372
rect 1203 350 1233 372
rect 1276 368 1338 384
rect 1366 377 1377 393
rect 1382 388 1392 408
rect 1402 388 1416 408
rect 1419 395 1428 408
rect 1444 395 1453 408
rect 1382 377 1416 388
rect 1419 377 1428 393
rect 1444 377 1453 393
rect 1460 388 1470 408
rect 1480 388 1494 408
rect 1495 395 1506 408
rect 1460 377 1494 388
rect 1495 377 1506 393
rect 1552 384 1568 400
rect 1575 398 1605 450
rect 1639 446 1640 453
rect 1624 438 1640 446
rect 1611 406 1624 425
rect 1639 406 1669 422
rect 1611 390 1685 406
rect 1611 388 1624 390
rect 1639 388 1673 390
rect 1276 366 1289 368
rect 1304 366 1338 368
rect 1276 350 1338 366
rect 1382 361 1398 364
rect 1460 361 1490 372
rect 1538 368 1584 384
rect 1611 372 1685 388
rect 1538 366 1572 368
rect 1537 350 1584 366
rect 1611 350 1624 372
rect 1639 350 1669 372
rect 1696 350 1697 366
rect 1712 350 1725 510
rect 1755 406 1768 510
rect 1813 488 1814 498
rect 1829 488 1842 498
rect 1813 484 1842 488
rect 1847 484 1877 510
rect 1895 496 1911 498
rect 1983 496 2036 510
rect 1984 494 2048 496
rect 2091 494 2106 510
rect 2155 507 2185 510
rect 2155 504 2191 507
rect 2121 496 2137 498
rect 1895 484 1910 488
rect 1813 482 1910 484
rect 1938 482 2106 494
rect 2122 484 2137 488
rect 2155 485 2194 504
rect 2213 498 2220 499
rect 2219 491 2220 498
rect 2203 488 2204 491
rect 2219 488 2232 491
rect 2155 484 2185 485
rect 2194 484 2200 485
rect 2203 484 2232 488
rect 2122 483 2232 484
rect 2122 482 2238 483
rect 1797 474 1848 482
rect 1797 462 1822 474
rect 1829 462 1848 474
rect 1879 474 1929 482
rect 1879 466 1895 474
rect 1902 472 1929 474
rect 1938 472 2159 482
rect 1902 462 2159 472
rect 2188 474 2238 482
rect 2188 465 2204 474
rect 1797 454 1848 462
rect 1895 454 2159 462
rect 2185 462 2204 465
rect 2211 462 2238 474
rect 2185 454 2238 462
rect 1813 446 1814 454
rect 1829 446 1842 454
rect 1813 438 1829 446
rect 1810 431 1829 434
rect 1810 422 1832 431
rect 1783 412 1832 422
rect 1783 406 1813 412
rect 1832 407 1837 412
rect 1755 390 1829 406
rect 1847 398 1877 454
rect 1912 444 2120 454
rect 2155 450 2200 454
rect 2203 453 2204 454
rect 2219 453 2232 454
rect 1938 414 2127 444
rect 1953 411 2127 414
rect 1946 408 2127 411
rect 1755 388 1768 390
rect 1783 388 1817 390
rect 1755 372 1829 388
rect 1856 384 1869 398
rect 1884 384 1900 400
rect 1946 395 1957 408
rect 1739 350 1740 366
rect 1755 350 1768 372
rect 1783 350 1813 372
rect 1856 368 1918 384
rect 1946 377 1957 393
rect 1962 388 1972 408
rect 1982 388 1996 408
rect 1999 395 2008 408
rect 2024 395 2033 408
rect 1962 377 1996 388
rect 1999 377 2008 393
rect 2024 377 2033 393
rect 2040 388 2050 408
rect 2060 388 2074 408
rect 2075 395 2086 408
rect 2040 377 2074 388
rect 2075 377 2086 393
rect 2132 384 2148 400
rect 2155 398 2185 450
rect 2219 446 2220 453
rect 2204 438 2220 446
rect 2191 406 2204 425
rect 2219 406 2249 422
rect 2191 390 2265 406
rect 2191 388 2204 390
rect 2219 388 2253 390
rect 1856 366 1869 368
rect 1884 366 1918 368
rect 1856 350 1918 366
rect 1962 361 1978 364
rect 2040 361 2070 372
rect 2118 368 2164 384
rect 2191 372 2265 388
rect 2118 366 2152 368
rect 2117 350 2164 366
rect 2191 350 2204 372
rect 2219 350 2249 372
rect 2276 350 2277 366
rect 2292 350 2305 510
rect 2335 406 2348 510
rect 2393 488 2394 498
rect 2409 488 2422 498
rect 2393 484 2422 488
rect 2427 484 2457 510
rect 2475 496 2491 498
rect 2563 496 2616 510
rect 2564 494 2628 496
rect 2671 494 2686 510
rect 2735 507 2765 510
rect 2735 504 2771 507
rect 2701 496 2717 498
rect 2475 484 2490 488
rect 2393 482 2490 484
rect 2518 482 2686 494
rect 2702 484 2717 488
rect 2735 485 2774 504
rect 2793 498 2800 499
rect 2799 491 2800 498
rect 2783 488 2784 491
rect 2799 488 2812 491
rect 2735 484 2765 485
rect 2774 484 2780 485
rect 2783 484 2812 488
rect 2702 483 2812 484
rect 2702 482 2818 483
rect 2377 474 2428 482
rect 2377 462 2402 474
rect 2409 462 2428 474
rect 2459 474 2509 482
rect 2459 466 2475 474
rect 2482 472 2509 474
rect 2518 472 2739 482
rect 2482 462 2739 472
rect 2768 474 2818 482
rect 2768 465 2784 474
rect 2377 454 2428 462
rect 2475 454 2739 462
rect 2765 462 2784 465
rect 2791 462 2818 474
rect 2765 454 2818 462
rect 2393 446 2394 454
rect 2409 446 2422 454
rect 2393 438 2409 446
rect 2390 431 2409 434
rect 2390 422 2412 431
rect 2363 412 2412 422
rect 2363 406 2393 412
rect 2412 407 2417 412
rect 2335 390 2409 406
rect 2427 398 2457 454
rect 2492 444 2700 454
rect 2735 450 2780 454
rect 2783 453 2784 454
rect 2799 453 2812 454
rect 2518 414 2707 444
rect 2533 411 2707 414
rect 2526 408 2707 411
rect 2335 388 2348 390
rect 2363 388 2397 390
rect 2335 372 2409 388
rect 2436 384 2449 398
rect 2464 384 2480 400
rect 2526 395 2537 408
rect 2319 350 2320 366
rect 2335 350 2348 372
rect 2363 350 2393 372
rect 2436 368 2498 384
rect 2526 377 2537 393
rect 2542 388 2552 408
rect 2562 388 2576 408
rect 2579 395 2588 408
rect 2604 395 2613 408
rect 2542 377 2576 388
rect 2579 377 2588 393
rect 2604 377 2613 393
rect 2620 388 2630 408
rect 2640 388 2654 408
rect 2655 395 2666 408
rect 2620 377 2654 388
rect 2655 377 2666 393
rect 2712 384 2728 400
rect 2735 398 2765 450
rect 2799 446 2800 453
rect 2784 438 2800 446
rect 2771 406 2784 425
rect 2799 406 2829 422
rect 2771 390 2845 406
rect 2771 388 2784 390
rect 2799 388 2833 390
rect 2436 366 2449 368
rect 2464 366 2498 368
rect 2436 350 2498 366
rect 2542 361 2558 364
rect 2620 361 2650 372
rect 2698 368 2744 384
rect 2771 372 2845 388
rect 2698 366 2732 368
rect 2697 350 2744 366
rect 2771 350 2784 372
rect 2799 350 2829 372
rect 2856 350 2857 366
rect 2872 350 2885 510
rect 2915 406 2928 510
rect 2973 488 2974 498
rect 2989 488 3002 498
rect 2973 484 3002 488
rect 3007 484 3037 510
rect 3055 496 3071 498
rect 3143 496 3196 510
rect 3144 494 3208 496
rect 3251 494 3266 510
rect 3315 507 3345 510
rect 3315 504 3351 507
rect 3281 496 3297 498
rect 3055 484 3070 488
rect 2973 482 3070 484
rect 3098 482 3266 494
rect 3282 484 3297 488
rect 3315 485 3354 504
rect 3373 498 3380 499
rect 3379 491 3380 498
rect 3363 488 3364 491
rect 3379 488 3392 491
rect 3315 484 3345 485
rect 3354 484 3360 485
rect 3363 484 3392 488
rect 3282 483 3392 484
rect 3282 482 3398 483
rect 2957 474 3008 482
rect 2957 462 2982 474
rect 2989 462 3008 474
rect 3039 474 3089 482
rect 3039 466 3055 474
rect 3062 472 3089 474
rect 3098 472 3319 482
rect 3062 462 3319 472
rect 3348 474 3398 482
rect 3348 465 3364 474
rect 2957 454 3008 462
rect 3055 454 3319 462
rect 3345 462 3364 465
rect 3371 462 3398 474
rect 3345 454 3398 462
rect 2973 446 2974 454
rect 2989 446 3002 454
rect 2973 438 2989 446
rect 2970 431 2989 434
rect 2970 422 2992 431
rect 2943 412 2992 422
rect 2943 406 2973 412
rect 2992 407 2997 412
rect 2915 390 2989 406
rect 3007 398 3037 454
rect 3072 444 3280 454
rect 3315 450 3360 454
rect 3363 453 3364 454
rect 3379 453 3392 454
rect 3098 414 3287 444
rect 3113 411 3287 414
rect 3106 408 3287 411
rect 2915 388 2928 390
rect 2943 388 2977 390
rect 2915 372 2989 388
rect 3016 384 3029 398
rect 3044 384 3060 400
rect 3106 395 3117 408
rect 2899 350 2900 366
rect 2915 350 2928 372
rect 2943 350 2973 372
rect 3016 368 3078 384
rect 3106 377 3117 393
rect 3122 388 3132 408
rect 3142 388 3156 408
rect 3159 395 3168 408
rect 3184 395 3193 408
rect 3122 377 3156 388
rect 3159 377 3168 393
rect 3184 377 3193 393
rect 3200 388 3210 408
rect 3220 388 3234 408
rect 3235 395 3246 408
rect 3200 377 3234 388
rect 3235 377 3246 393
rect 3292 384 3308 400
rect 3315 398 3345 450
rect 3379 446 3380 453
rect 3364 438 3380 446
rect 3351 406 3364 425
rect 3379 406 3409 422
rect 3351 390 3425 406
rect 3351 388 3364 390
rect 3379 388 3413 390
rect 3016 366 3029 368
rect 3044 366 3078 368
rect 3016 350 3078 366
rect 3122 361 3138 364
rect 3200 361 3230 372
rect 3278 368 3324 384
rect 3351 372 3425 388
rect 3278 366 3312 368
rect 3277 350 3324 366
rect 3351 350 3364 372
rect 3379 350 3409 372
rect 3436 350 3437 366
rect 3452 350 3465 510
rect 3495 406 3508 510
rect 3553 488 3554 498
rect 3569 488 3582 498
rect 3553 484 3582 488
rect 3587 484 3617 510
rect 3635 496 3651 498
rect 3723 496 3776 510
rect 3724 494 3788 496
rect 3831 494 3846 510
rect 3895 507 3925 510
rect 3895 504 3931 507
rect 3861 496 3877 498
rect 3635 484 3650 488
rect 3553 482 3650 484
rect 3678 482 3846 494
rect 3862 484 3877 488
rect 3895 485 3934 504
rect 3953 498 3960 499
rect 3959 491 3960 498
rect 3943 488 3944 491
rect 3959 488 3972 491
rect 3895 484 3925 485
rect 3934 484 3940 485
rect 3943 484 3972 488
rect 3862 483 3972 484
rect 3862 482 3978 483
rect 3537 474 3588 482
rect 3537 462 3562 474
rect 3569 462 3588 474
rect 3619 474 3669 482
rect 3619 466 3635 474
rect 3642 472 3669 474
rect 3678 472 3899 482
rect 3642 462 3899 472
rect 3928 474 3978 482
rect 3928 465 3944 474
rect 3537 454 3588 462
rect 3635 454 3899 462
rect 3925 462 3944 465
rect 3951 462 3978 474
rect 3925 454 3978 462
rect 3553 446 3554 454
rect 3569 446 3582 454
rect 3553 438 3569 446
rect 3550 431 3569 434
rect 3550 422 3572 431
rect 3523 412 3572 422
rect 3523 406 3553 412
rect 3572 407 3577 412
rect 3495 390 3569 406
rect 3587 398 3617 454
rect 3652 444 3860 454
rect 3895 450 3940 454
rect 3943 453 3944 454
rect 3959 453 3972 454
rect 3678 414 3867 444
rect 3693 411 3867 414
rect 3686 408 3867 411
rect 3495 388 3508 390
rect 3523 388 3557 390
rect 3495 372 3569 388
rect 3596 384 3609 398
rect 3624 384 3640 400
rect 3686 395 3697 408
rect 3479 350 3480 366
rect 3495 350 3508 372
rect 3523 350 3553 372
rect 3596 368 3658 384
rect 3686 377 3697 393
rect 3702 388 3712 408
rect 3722 388 3736 408
rect 3739 395 3748 408
rect 3764 395 3773 408
rect 3702 377 3736 388
rect 3739 377 3748 393
rect 3764 377 3773 393
rect 3780 388 3790 408
rect 3800 388 3814 408
rect 3815 395 3826 408
rect 3780 377 3814 388
rect 3815 377 3826 393
rect 3872 384 3888 400
rect 3895 398 3925 450
rect 3959 446 3960 453
rect 3944 438 3960 446
rect 3931 406 3944 425
rect 3959 406 3989 422
rect 3931 390 4005 406
rect 3931 388 3944 390
rect 3959 388 3993 390
rect 3596 366 3609 368
rect 3624 366 3658 368
rect 3596 350 3658 366
rect 3702 361 3718 364
rect 3780 361 3810 372
rect 3858 368 3904 384
rect 3931 372 4005 388
rect 3858 366 3892 368
rect 3857 350 3904 366
rect 3931 350 3944 372
rect 3959 350 3989 372
rect 4016 350 4017 366
rect 4032 350 4045 510
rect 4075 406 4088 510
rect 4133 488 4134 498
rect 4149 488 4162 498
rect 4133 484 4162 488
rect 4167 484 4197 510
rect 4215 496 4231 498
rect 4303 496 4356 510
rect 4304 494 4368 496
rect 4411 494 4426 510
rect 4475 507 4505 510
rect 4475 504 4511 507
rect 4441 496 4457 498
rect 4215 484 4230 488
rect 4133 482 4230 484
rect 4258 482 4426 494
rect 4442 484 4457 488
rect 4475 485 4514 504
rect 4533 498 4540 499
rect 4539 491 4540 498
rect 4523 488 4524 491
rect 4539 488 4552 491
rect 4475 484 4505 485
rect 4514 484 4520 485
rect 4523 484 4552 488
rect 4442 483 4552 484
rect 4442 482 4558 483
rect 4117 474 4168 482
rect 4117 462 4142 474
rect 4149 462 4168 474
rect 4199 474 4249 482
rect 4199 466 4215 474
rect 4222 472 4249 474
rect 4258 472 4479 482
rect 4222 462 4479 472
rect 4508 474 4558 482
rect 4508 465 4524 474
rect 4117 454 4168 462
rect 4215 454 4479 462
rect 4505 462 4524 465
rect 4531 462 4558 474
rect 4505 454 4558 462
rect 4133 446 4134 454
rect 4149 446 4162 454
rect 4133 438 4149 446
rect 4130 431 4149 434
rect 4130 422 4152 431
rect 4103 412 4152 422
rect 4103 406 4133 412
rect 4152 407 4157 412
rect 4075 390 4149 406
rect 4167 398 4197 454
rect 4232 444 4440 454
rect 4475 450 4520 454
rect 4523 453 4524 454
rect 4539 453 4552 454
rect 4258 414 4447 444
rect 4273 411 4447 414
rect 4266 408 4447 411
rect 4075 388 4088 390
rect 4103 388 4137 390
rect 4075 372 4149 388
rect 4176 384 4189 398
rect 4204 384 4220 400
rect 4266 395 4277 408
rect 4059 350 4060 366
rect 4075 350 4088 372
rect 4103 350 4133 372
rect 4176 368 4238 384
rect 4266 377 4277 393
rect 4282 388 4292 408
rect 4302 388 4316 408
rect 4319 395 4328 408
rect 4344 395 4353 408
rect 4282 377 4316 388
rect 4319 377 4328 393
rect 4344 377 4353 393
rect 4360 388 4370 408
rect 4380 388 4394 408
rect 4395 395 4406 408
rect 4360 377 4394 388
rect 4395 377 4406 393
rect 4452 384 4468 400
rect 4475 398 4505 450
rect 4539 446 4540 453
rect 4524 438 4540 446
rect 4511 406 4524 425
rect 4539 406 4569 422
rect 4511 390 4585 406
rect 4511 388 4524 390
rect 4539 388 4573 390
rect 4176 366 4189 368
rect 4204 366 4238 368
rect 4176 350 4238 366
rect 4282 361 4298 364
rect 4360 361 4390 372
rect 4438 368 4484 384
rect 4511 372 4585 388
rect 4438 366 4472 368
rect 4437 350 4484 366
rect 4511 350 4524 372
rect 4539 350 4569 372
rect 4596 350 4597 366
rect 4612 350 4625 510
rect -7 342 34 350
rect -7 316 8 342
rect 15 316 34 342
rect 98 338 160 350
rect 172 338 247 350
rect 305 338 380 350
rect 392 338 423 350
rect 429 338 464 350
rect 98 336 260 338
rect -7 308 34 316
rect 116 312 129 336
rect 144 334 159 336
rect -1 298 0 308
rect 15 298 28 308
rect 43 298 73 312
rect 116 298 159 312
rect 183 309 190 316
rect 193 312 260 336
rect 292 336 464 338
rect 262 314 290 318
rect 292 314 372 336
rect 393 334 408 336
rect 262 312 372 314
rect 193 308 372 312
rect 166 298 196 308
rect 198 298 351 308
rect 359 298 389 308
rect 393 298 423 312
rect 451 298 464 336
rect 536 342 571 350
rect 536 316 537 342
rect 544 316 571 342
rect 479 298 509 312
rect 536 308 571 316
rect 573 342 614 350
rect 573 316 588 342
rect 595 316 614 342
rect 678 338 740 350
rect 752 338 827 350
rect 885 338 960 350
rect 972 338 1003 350
rect 1009 338 1044 350
rect 678 336 840 338
rect 573 308 614 316
rect 696 312 709 336
rect 724 334 739 336
rect 536 298 537 308
rect 552 298 565 308
rect 579 298 580 308
rect 595 298 608 308
rect 623 298 653 312
rect 696 298 739 312
rect 763 309 770 316
rect 773 312 840 336
rect 872 336 1044 338
rect 842 314 870 318
rect 872 314 952 336
rect 973 334 988 336
rect 842 312 952 314
rect 773 308 952 312
rect 746 298 776 308
rect 778 298 931 308
rect 939 298 969 308
rect 973 298 1003 312
rect 1031 298 1044 336
rect 1116 342 1151 350
rect 1116 316 1117 342
rect 1124 316 1151 342
rect 1059 298 1089 312
rect 1116 308 1151 316
rect 1153 342 1194 350
rect 1153 316 1168 342
rect 1175 316 1194 342
rect 1258 338 1320 350
rect 1332 338 1407 350
rect 1465 338 1540 350
rect 1552 338 1583 350
rect 1589 338 1624 350
rect 1258 336 1420 338
rect 1153 308 1194 316
rect 1276 312 1289 336
rect 1304 334 1319 336
rect 1116 298 1117 308
rect 1132 298 1145 308
rect 1159 298 1160 308
rect 1175 298 1188 308
rect 1203 298 1233 312
rect 1276 298 1319 312
rect 1343 309 1350 316
rect 1353 312 1420 336
rect 1452 336 1624 338
rect 1422 314 1450 318
rect 1452 314 1532 336
rect 1553 334 1568 336
rect 1422 312 1532 314
rect 1353 308 1532 312
rect 1326 298 1356 308
rect 1358 298 1511 308
rect 1519 298 1549 308
rect 1553 298 1583 312
rect 1611 298 1624 336
rect 1696 342 1731 350
rect 1696 316 1697 342
rect 1704 316 1731 342
rect 1639 298 1669 312
rect 1696 308 1731 316
rect 1733 342 1774 350
rect 1733 316 1748 342
rect 1755 316 1774 342
rect 1838 338 1900 350
rect 1912 338 1987 350
rect 2045 338 2120 350
rect 2132 338 2163 350
rect 2169 338 2204 350
rect 1838 336 2000 338
rect 1733 308 1774 316
rect 1856 312 1869 336
rect 1884 334 1899 336
rect 1696 298 1697 308
rect 1712 298 1725 308
rect 1739 298 1740 308
rect 1755 298 1768 308
rect 1783 298 1813 312
rect 1856 298 1899 312
rect 1923 309 1930 316
rect 1933 312 2000 336
rect 2032 336 2204 338
rect 2002 314 2030 318
rect 2032 314 2112 336
rect 2133 334 2148 336
rect 2002 312 2112 314
rect 1933 308 2112 312
rect 1906 298 1936 308
rect 1938 298 2091 308
rect 2099 298 2129 308
rect 2133 298 2163 312
rect 2191 298 2204 336
rect 2276 342 2311 350
rect 2276 316 2277 342
rect 2284 316 2311 342
rect 2219 298 2249 312
rect 2276 308 2311 316
rect 2313 342 2354 350
rect 2313 316 2328 342
rect 2335 316 2354 342
rect 2418 338 2480 350
rect 2492 338 2567 350
rect 2625 338 2700 350
rect 2712 338 2743 350
rect 2749 338 2784 350
rect 2418 336 2580 338
rect 2313 308 2354 316
rect 2436 312 2449 336
rect 2464 334 2479 336
rect 2276 298 2277 308
rect 2292 298 2305 308
rect 2319 298 2320 308
rect 2335 298 2348 308
rect 2363 298 2393 312
rect 2436 298 2479 312
rect 2503 309 2510 316
rect 2513 312 2580 336
rect 2612 336 2784 338
rect 2582 314 2610 318
rect 2612 314 2692 336
rect 2713 334 2728 336
rect 2582 312 2692 314
rect 2513 308 2692 312
rect 2486 298 2516 308
rect 2518 298 2671 308
rect 2679 298 2709 308
rect 2713 298 2743 312
rect 2771 298 2784 336
rect 2856 342 2891 350
rect 2856 316 2857 342
rect 2864 316 2891 342
rect 2799 298 2829 312
rect 2856 308 2891 316
rect 2893 342 2934 350
rect 2893 316 2908 342
rect 2915 316 2934 342
rect 2998 338 3060 350
rect 3072 338 3147 350
rect 3205 338 3280 350
rect 3292 338 3323 350
rect 3329 338 3364 350
rect 2998 336 3160 338
rect 2893 308 2934 316
rect 3016 312 3029 336
rect 3044 334 3059 336
rect 2856 298 2857 308
rect 2872 298 2885 308
rect 2899 298 2900 308
rect 2915 298 2928 308
rect 2943 298 2973 312
rect 3016 298 3059 312
rect 3083 309 3090 316
rect 3093 312 3160 336
rect 3192 336 3364 338
rect 3162 314 3190 318
rect 3192 314 3272 336
rect 3293 334 3308 336
rect 3162 312 3272 314
rect 3093 308 3272 312
rect 3066 298 3096 308
rect 3098 298 3251 308
rect 3259 298 3289 308
rect 3293 298 3323 312
rect 3351 298 3364 336
rect 3436 342 3471 350
rect 3436 316 3437 342
rect 3444 316 3471 342
rect 3379 298 3409 312
rect 3436 308 3471 316
rect 3473 342 3514 350
rect 3473 316 3488 342
rect 3495 316 3514 342
rect 3578 338 3640 350
rect 3652 338 3727 350
rect 3785 338 3860 350
rect 3872 338 3903 350
rect 3909 338 3944 350
rect 3578 336 3740 338
rect 3473 308 3514 316
rect 3596 312 3609 336
rect 3624 334 3639 336
rect 3436 298 3437 308
rect 3452 298 3465 308
rect 3479 298 3480 308
rect 3495 298 3508 308
rect 3523 298 3553 312
rect 3596 298 3639 312
rect 3663 309 3670 316
rect 3673 312 3740 336
rect 3772 336 3944 338
rect 3742 314 3770 318
rect 3772 314 3852 336
rect 3873 334 3888 336
rect 3742 312 3852 314
rect 3673 308 3852 312
rect 3646 298 3676 308
rect 3678 298 3831 308
rect 3839 298 3869 308
rect 3873 298 3903 312
rect 3931 298 3944 336
rect 4016 342 4051 350
rect 4016 316 4017 342
rect 4024 316 4051 342
rect 3959 298 3989 312
rect 4016 308 4051 316
rect 4053 342 4094 350
rect 4053 316 4068 342
rect 4075 316 4094 342
rect 4158 338 4220 350
rect 4232 338 4307 350
rect 4365 338 4440 350
rect 4452 338 4483 350
rect 4489 338 4524 350
rect 4158 336 4320 338
rect 4053 308 4094 316
rect 4176 312 4189 336
rect 4204 334 4219 336
rect 4016 298 4017 308
rect 4032 298 4045 308
rect 4059 298 4060 308
rect 4075 298 4088 308
rect 4103 298 4133 312
rect 4176 298 4219 312
rect 4243 309 4250 316
rect 4253 312 4320 336
rect 4352 336 4524 338
rect 4322 314 4350 318
rect 4352 314 4432 336
rect 4453 334 4468 336
rect 4322 312 4432 314
rect 4253 308 4432 312
rect 4226 298 4256 308
rect 4258 298 4411 308
rect 4419 298 4449 308
rect 4453 298 4483 312
rect 4511 298 4524 336
rect 4596 342 4631 350
rect 4596 316 4597 342
rect 4604 316 4631 342
rect 4539 298 4569 312
rect 4596 308 4631 316
rect 4596 298 4597 308
rect 4612 298 4625 308
rect -1 292 4625 298
rect 0 284 4625 292
rect 15 254 28 284
rect 43 266 73 284
rect 116 270 130 284
rect 166 270 386 284
rect 117 268 130 270
rect 83 256 98 268
rect 80 254 102 256
rect 107 254 137 268
rect 198 266 351 270
rect 180 254 372 266
rect 415 254 445 268
rect 451 254 464 284
rect 479 266 509 284
rect 552 254 565 284
rect 595 254 608 284
rect 623 266 653 284
rect 696 270 710 284
rect 746 270 966 284
rect 697 268 710 270
rect 663 256 678 268
rect 660 254 682 256
rect 687 254 717 268
rect 778 266 931 270
rect 760 254 952 266
rect 995 254 1025 268
rect 1031 254 1044 284
rect 1059 266 1089 284
rect 1132 254 1145 284
rect 1175 254 1188 284
rect 1203 266 1233 284
rect 1276 270 1290 284
rect 1326 270 1546 284
rect 1277 268 1290 270
rect 1243 256 1258 268
rect 1240 254 1262 256
rect 1267 254 1297 268
rect 1358 266 1511 270
rect 1340 254 1532 266
rect 1575 254 1605 268
rect 1611 254 1624 284
rect 1639 266 1669 284
rect 1712 254 1725 284
rect 1755 254 1768 284
rect 1783 266 1813 284
rect 1856 270 1870 284
rect 1906 270 2126 284
rect 1857 268 1870 270
rect 1823 256 1838 268
rect 1820 254 1842 256
rect 1847 254 1877 268
rect 1938 266 2091 270
rect 1920 254 2112 266
rect 2155 254 2185 268
rect 2191 254 2204 284
rect 2219 266 2249 284
rect 2292 254 2305 284
rect 2335 254 2348 284
rect 2363 266 2393 284
rect 2436 270 2450 284
rect 2486 270 2706 284
rect 2437 268 2450 270
rect 2403 256 2418 268
rect 2400 254 2422 256
rect 2427 254 2457 268
rect 2518 266 2671 270
rect 2500 254 2692 266
rect 2735 254 2765 268
rect 2771 254 2784 284
rect 2799 266 2829 284
rect 2872 254 2885 284
rect 2915 254 2928 284
rect 2943 266 2973 284
rect 3016 270 3030 284
rect 3066 270 3286 284
rect 3017 268 3030 270
rect 2983 256 2998 268
rect 2980 254 3002 256
rect 3007 254 3037 268
rect 3098 266 3251 270
rect 3080 254 3272 266
rect 3315 254 3345 268
rect 3351 254 3364 284
rect 3379 266 3409 284
rect 3452 254 3465 284
rect 3495 254 3508 284
rect 3523 266 3553 284
rect 3596 270 3610 284
rect 3646 270 3866 284
rect 3597 268 3610 270
rect 3563 256 3578 268
rect 3560 254 3582 256
rect 3587 254 3617 268
rect 3678 266 3831 270
rect 3660 254 3852 266
rect 3895 254 3925 268
rect 3931 254 3944 284
rect 3959 266 3989 284
rect 4032 254 4045 284
rect 4075 254 4088 284
rect 4103 266 4133 284
rect 4176 270 4190 284
rect 4226 270 4446 284
rect 4177 268 4190 270
rect 4143 256 4158 268
rect 4140 254 4162 256
rect 4167 254 4197 268
rect 4258 266 4411 270
rect 4240 254 4432 266
rect 4475 254 4505 268
rect 4511 254 4524 284
rect 4539 266 4569 284
rect 4612 254 4625 284
rect 0 240 4625 254
rect 15 136 28 240
rect 73 218 74 228
rect 89 218 102 228
rect 73 214 102 218
rect 107 214 137 240
rect 155 226 171 228
rect 243 226 296 240
rect 244 224 308 226
rect 155 214 170 218
rect 73 212 170 214
rect 57 204 108 212
rect 57 192 82 204
rect 89 192 108 204
rect 139 204 189 212
rect 139 196 155 204
rect 162 202 189 204
rect 198 204 213 208
rect 260 204 292 224
rect 351 212 366 240
rect 415 237 445 240
rect 415 234 451 237
rect 381 226 397 228
rect 382 214 397 218
rect 415 215 454 234
rect 473 228 480 229
rect 479 221 480 228
rect 463 218 464 221
rect 479 218 492 221
rect 415 214 445 215
rect 454 214 460 215
rect 463 214 492 218
rect 382 213 492 214
rect 382 212 498 213
rect 351 204 419 212
rect 198 202 267 204
rect 285 202 419 204
rect 162 198 234 202
rect 162 196 287 198
rect 162 192 234 196
rect 57 184 108 192
rect 155 188 234 192
rect 315 188 419 202
rect 448 204 498 212
rect 448 195 464 204
rect 155 184 419 188
rect 445 192 464 195
rect 471 192 498 204
rect 445 184 498 192
rect 73 176 74 184
rect 89 176 102 184
rect 73 168 89 176
rect 70 161 89 164
rect 70 152 92 161
rect 43 142 92 152
rect 43 136 73 142
rect 92 137 97 142
rect 15 120 89 136
rect 107 128 137 184
rect 172 174 380 184
rect 415 180 460 184
rect 463 183 464 184
rect 479 183 492 184
rect 339 170 387 174
rect 222 148 252 157
rect 315 150 330 157
rect 351 148 387 170
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 15 118 28 120
rect 43 118 77 120
rect 15 102 89 118
rect 116 114 129 128
rect 144 114 160 130
rect 206 125 217 138
rect -1 80 0 96
rect 15 80 28 102
rect 43 80 73 102
rect 116 98 178 114
rect 206 107 217 123
rect 222 118 232 138
rect 242 118 256 138
rect 259 125 268 138
rect 284 125 293 138
rect 222 107 256 118
rect 259 107 267 123
rect 284 107 293 123
rect 300 118 310 138
rect 320 118 334 138
rect 335 125 346 138
rect 300 107 334 118
rect 335 107 346 123
rect 392 114 408 130
rect 415 128 445 180
rect 479 176 480 183
rect 464 168 480 176
rect 451 136 464 155
rect 479 136 509 152
rect 451 120 525 136
rect 451 118 464 120
rect 479 118 513 120
rect 116 96 129 98
rect 144 96 178 98
rect 116 80 178 96
rect 222 91 235 94
rect 300 91 330 102
rect 378 98 424 114
rect 451 102 525 118
rect 378 96 412 98
rect 377 80 424 96
rect 451 80 464 102
rect 479 80 509 102
rect 536 80 537 96
rect 552 80 565 240
rect 595 136 608 240
rect 653 218 654 228
rect 669 218 682 228
rect 653 214 682 218
rect 687 214 717 240
rect 735 226 751 228
rect 823 226 876 240
rect 824 224 888 226
rect 735 214 750 218
rect 653 212 750 214
rect 637 204 688 212
rect 637 192 662 204
rect 669 192 688 204
rect 719 204 769 212
rect 719 196 735 204
rect 742 202 769 204
rect 778 204 793 208
rect 840 204 872 224
rect 931 212 946 240
rect 995 237 1025 240
rect 995 234 1031 237
rect 961 226 977 228
rect 962 214 977 218
rect 995 215 1034 234
rect 1053 228 1060 229
rect 1059 221 1060 228
rect 1043 218 1044 221
rect 1059 218 1072 221
rect 995 214 1025 215
rect 1034 214 1040 215
rect 1043 214 1072 218
rect 962 213 1072 214
rect 962 212 1078 213
rect 931 204 999 212
rect 778 202 847 204
rect 865 202 999 204
rect 742 198 814 202
rect 742 196 867 198
rect 742 192 814 196
rect 637 184 688 192
rect 735 188 814 192
rect 895 188 999 202
rect 1028 204 1078 212
rect 1028 195 1044 204
rect 735 184 999 188
rect 1025 192 1044 195
rect 1051 192 1078 204
rect 1025 184 1078 192
rect 653 176 654 184
rect 669 176 682 184
rect 653 168 669 176
rect 650 161 669 164
rect 650 152 672 161
rect 623 142 672 152
rect 623 136 653 142
rect 672 137 677 142
rect 595 120 669 136
rect 687 128 717 184
rect 752 174 960 184
rect 995 180 1040 184
rect 1043 183 1044 184
rect 1059 183 1072 184
rect 919 170 967 174
rect 802 148 832 157
rect 895 150 910 157
rect 931 148 967 170
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 595 118 608 120
rect 623 118 657 120
rect 595 102 669 118
rect 696 114 709 128
rect 724 114 740 130
rect 786 125 797 138
rect 579 80 580 96
rect 595 80 608 102
rect 623 80 653 102
rect 696 98 758 114
rect 786 107 797 123
rect 802 118 812 138
rect 822 118 836 138
rect 839 125 848 138
rect 864 125 873 138
rect 802 107 836 118
rect 839 107 847 123
rect 864 107 873 123
rect 880 118 890 138
rect 900 118 914 138
rect 915 125 926 138
rect 880 107 914 118
rect 915 107 926 123
rect 972 114 988 130
rect 995 128 1025 180
rect 1059 176 1060 183
rect 1044 168 1060 176
rect 1031 136 1044 155
rect 1059 136 1089 152
rect 1031 120 1105 136
rect 1031 118 1044 120
rect 1059 118 1093 120
rect 696 96 709 98
rect 724 96 758 98
rect 696 80 758 96
rect 802 91 815 94
rect 880 91 910 102
rect 958 98 1004 114
rect 1031 102 1105 118
rect 958 96 992 98
rect 957 80 1004 96
rect 1031 80 1044 102
rect 1059 80 1089 102
rect 1116 80 1117 96
rect 1132 80 1145 240
rect 1175 136 1188 240
rect 1233 218 1234 228
rect 1249 218 1262 228
rect 1233 214 1262 218
rect 1267 214 1297 240
rect 1315 226 1331 228
rect 1403 226 1456 240
rect 1404 224 1468 226
rect 1315 214 1330 218
rect 1233 212 1330 214
rect 1217 204 1268 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1299 204 1349 212
rect 1299 196 1315 204
rect 1322 202 1349 204
rect 1358 204 1373 208
rect 1420 204 1452 224
rect 1511 212 1526 240
rect 1575 237 1605 240
rect 1575 234 1611 237
rect 1541 226 1557 228
rect 1542 214 1557 218
rect 1575 215 1614 234
rect 1633 228 1640 229
rect 1639 221 1640 228
rect 1623 218 1624 221
rect 1639 218 1652 221
rect 1575 214 1605 215
rect 1614 214 1620 215
rect 1623 214 1652 218
rect 1542 213 1652 214
rect 1542 212 1658 213
rect 1511 204 1579 212
rect 1358 202 1427 204
rect 1445 202 1579 204
rect 1322 198 1394 202
rect 1322 196 1447 198
rect 1322 192 1394 196
rect 1217 184 1268 192
rect 1315 188 1394 192
rect 1475 188 1579 202
rect 1608 204 1658 212
rect 1608 195 1624 204
rect 1315 184 1579 188
rect 1605 192 1624 195
rect 1631 192 1658 204
rect 1605 184 1658 192
rect 1233 176 1234 184
rect 1249 176 1262 184
rect 1233 168 1249 176
rect 1230 161 1249 164
rect 1230 152 1252 161
rect 1203 142 1252 152
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1175 120 1249 136
rect 1267 128 1297 184
rect 1332 174 1540 184
rect 1575 180 1620 184
rect 1623 183 1624 184
rect 1639 183 1652 184
rect 1499 170 1547 174
rect 1382 148 1412 157
rect 1475 150 1490 157
rect 1511 148 1547 170
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1175 118 1188 120
rect 1203 118 1237 120
rect 1175 102 1249 118
rect 1276 114 1289 128
rect 1304 114 1320 130
rect 1366 125 1377 138
rect 1159 80 1160 96
rect 1175 80 1188 102
rect 1203 80 1233 102
rect 1276 98 1338 114
rect 1366 107 1377 123
rect 1382 118 1392 138
rect 1402 118 1416 138
rect 1419 125 1428 138
rect 1444 125 1453 138
rect 1382 107 1416 118
rect 1419 107 1427 123
rect 1444 107 1453 123
rect 1460 118 1470 138
rect 1480 118 1494 138
rect 1495 125 1506 138
rect 1460 107 1494 118
rect 1495 107 1506 123
rect 1552 114 1568 130
rect 1575 128 1605 180
rect 1639 176 1640 183
rect 1624 168 1640 176
rect 1611 136 1624 155
rect 1639 136 1669 152
rect 1611 120 1685 136
rect 1611 118 1624 120
rect 1639 118 1673 120
rect 1276 96 1289 98
rect 1304 96 1338 98
rect 1276 80 1338 96
rect 1382 91 1395 94
rect 1460 91 1490 102
rect 1538 98 1584 114
rect 1611 102 1685 118
rect 1538 96 1572 98
rect 1537 80 1584 96
rect 1611 80 1624 102
rect 1639 80 1669 102
rect 1696 80 1697 96
rect 1712 80 1725 240
rect 1755 136 1768 240
rect 1813 218 1814 228
rect 1829 218 1842 228
rect 1813 214 1842 218
rect 1847 214 1877 240
rect 1895 226 1911 228
rect 1983 226 2036 240
rect 1984 224 2048 226
rect 1895 214 1910 218
rect 1813 212 1910 214
rect 1797 204 1848 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1879 204 1929 212
rect 1879 196 1895 204
rect 1902 202 1929 204
rect 1938 204 1953 208
rect 2000 204 2032 224
rect 2091 212 2106 240
rect 2155 237 2185 240
rect 2155 234 2191 237
rect 2121 226 2137 228
rect 2122 214 2137 218
rect 2155 215 2194 234
rect 2213 228 2220 229
rect 2219 221 2220 228
rect 2203 218 2204 221
rect 2219 218 2232 221
rect 2155 214 2185 215
rect 2194 214 2200 215
rect 2203 214 2232 218
rect 2122 213 2232 214
rect 2122 212 2238 213
rect 2091 204 2159 212
rect 1938 202 2007 204
rect 2025 202 2159 204
rect 1902 198 1974 202
rect 1902 196 2027 198
rect 1902 192 1974 196
rect 1797 184 1848 192
rect 1895 188 1974 192
rect 2055 188 2159 202
rect 2188 204 2238 212
rect 2188 195 2204 204
rect 1895 184 2159 188
rect 2185 192 2204 195
rect 2211 192 2238 204
rect 2185 184 2238 192
rect 1813 176 1814 184
rect 1829 176 1842 184
rect 1813 168 1829 176
rect 1810 161 1829 164
rect 1810 152 1832 161
rect 1783 142 1832 152
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1755 120 1829 136
rect 1847 128 1877 184
rect 1912 174 2120 184
rect 2155 180 2200 184
rect 2203 183 2204 184
rect 2219 183 2232 184
rect 2079 170 2127 174
rect 1962 148 1992 157
rect 2055 150 2070 157
rect 2091 148 2127 170
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 1755 118 1768 120
rect 1783 118 1817 120
rect 1755 102 1829 118
rect 1856 114 1869 128
rect 1884 114 1900 130
rect 1946 125 1957 138
rect 1739 80 1740 96
rect 1755 80 1768 102
rect 1783 80 1813 102
rect 1856 98 1918 114
rect 1946 107 1957 123
rect 1962 118 1972 138
rect 1982 118 1996 138
rect 1999 125 2008 138
rect 2024 125 2033 138
rect 1962 107 1996 118
rect 1999 107 2007 123
rect 2024 107 2033 123
rect 2040 118 2050 138
rect 2060 118 2074 138
rect 2075 125 2086 138
rect 2040 107 2074 118
rect 2075 107 2086 123
rect 2132 114 2148 130
rect 2155 128 2185 180
rect 2219 176 2220 183
rect 2204 168 2220 176
rect 2191 136 2204 155
rect 2219 136 2249 152
rect 2191 120 2265 136
rect 2191 118 2204 120
rect 2219 118 2253 120
rect 1856 96 1869 98
rect 1884 96 1918 98
rect 1856 80 1918 96
rect 1962 91 1975 94
rect 2040 91 2070 102
rect 2118 98 2164 114
rect 2191 102 2265 118
rect 2118 96 2152 98
rect 2117 80 2164 96
rect 2191 80 2204 102
rect 2219 80 2249 102
rect 2276 80 2277 96
rect 2292 80 2305 240
rect 2335 136 2348 240
rect 2393 218 2394 228
rect 2409 218 2422 228
rect 2393 214 2422 218
rect 2427 214 2457 240
rect 2475 226 2491 228
rect 2563 226 2616 240
rect 2564 224 2628 226
rect 2475 214 2490 218
rect 2393 212 2490 214
rect 2377 204 2428 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2459 204 2509 212
rect 2459 196 2475 204
rect 2482 202 2509 204
rect 2518 204 2533 208
rect 2580 204 2612 224
rect 2671 212 2686 240
rect 2735 237 2765 240
rect 2735 234 2771 237
rect 2701 226 2717 228
rect 2702 214 2717 218
rect 2735 215 2774 234
rect 2793 228 2800 229
rect 2799 221 2800 228
rect 2783 218 2784 221
rect 2799 218 2812 221
rect 2735 214 2765 215
rect 2774 214 2780 215
rect 2783 214 2812 218
rect 2702 213 2812 214
rect 2702 212 2818 213
rect 2671 204 2739 212
rect 2518 202 2587 204
rect 2605 202 2739 204
rect 2482 198 2554 202
rect 2482 196 2607 198
rect 2482 192 2554 196
rect 2377 184 2428 192
rect 2475 188 2554 192
rect 2635 188 2739 202
rect 2768 204 2818 212
rect 2768 195 2784 204
rect 2475 184 2739 188
rect 2765 192 2784 195
rect 2791 192 2818 204
rect 2765 184 2818 192
rect 2393 176 2394 184
rect 2409 176 2422 184
rect 2393 168 2409 176
rect 2390 161 2409 164
rect 2390 152 2412 161
rect 2363 142 2412 152
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2335 120 2409 136
rect 2427 128 2457 184
rect 2492 174 2700 184
rect 2735 180 2780 184
rect 2783 183 2784 184
rect 2799 183 2812 184
rect 2659 170 2707 174
rect 2542 148 2572 157
rect 2635 150 2650 157
rect 2671 148 2707 170
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2335 118 2348 120
rect 2363 118 2397 120
rect 2335 102 2409 118
rect 2436 114 2449 128
rect 2464 114 2480 130
rect 2526 125 2537 138
rect 2319 80 2320 96
rect 2335 80 2348 102
rect 2363 80 2393 102
rect 2436 98 2498 114
rect 2526 107 2537 123
rect 2542 118 2552 138
rect 2562 118 2576 138
rect 2579 125 2588 138
rect 2604 125 2613 138
rect 2542 107 2576 118
rect 2579 107 2587 123
rect 2604 107 2613 123
rect 2620 118 2630 138
rect 2640 118 2654 138
rect 2655 125 2666 138
rect 2620 107 2654 118
rect 2655 107 2666 123
rect 2712 114 2728 130
rect 2735 128 2765 180
rect 2799 176 2800 183
rect 2784 168 2800 176
rect 2771 136 2784 155
rect 2799 136 2829 152
rect 2771 120 2845 136
rect 2771 118 2784 120
rect 2799 118 2833 120
rect 2436 96 2449 98
rect 2464 96 2498 98
rect 2436 80 2498 96
rect 2542 91 2555 94
rect 2620 91 2650 102
rect 2698 98 2744 114
rect 2771 102 2845 118
rect 2698 96 2732 98
rect 2697 80 2744 96
rect 2771 80 2784 102
rect 2799 80 2829 102
rect 2856 80 2857 96
rect 2872 80 2885 240
rect 2915 136 2928 240
rect 2973 218 2974 228
rect 2989 218 3002 228
rect 2973 214 3002 218
rect 3007 214 3037 240
rect 3055 226 3071 228
rect 3143 226 3196 240
rect 3144 224 3208 226
rect 3055 214 3070 218
rect 2973 212 3070 214
rect 2957 204 3008 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3039 204 3089 212
rect 3039 196 3055 204
rect 3062 202 3089 204
rect 3098 204 3113 208
rect 3160 204 3192 224
rect 3251 212 3266 240
rect 3315 237 3345 240
rect 3315 234 3351 237
rect 3281 226 3297 228
rect 3282 214 3297 218
rect 3315 215 3354 234
rect 3373 228 3380 229
rect 3379 221 3380 228
rect 3363 218 3364 221
rect 3379 218 3392 221
rect 3315 214 3345 215
rect 3354 214 3360 215
rect 3363 214 3392 218
rect 3282 213 3392 214
rect 3282 212 3398 213
rect 3251 204 3319 212
rect 3098 202 3167 204
rect 3185 202 3319 204
rect 3062 198 3134 202
rect 3062 196 3187 198
rect 3062 192 3134 196
rect 2957 184 3008 192
rect 3055 188 3134 192
rect 3215 188 3319 202
rect 3348 204 3398 212
rect 3348 195 3364 204
rect 3055 184 3319 188
rect 3345 192 3364 195
rect 3371 192 3398 204
rect 3345 184 3398 192
rect 2973 176 2974 184
rect 2989 176 3002 184
rect 2973 168 2989 176
rect 2970 161 2989 164
rect 2970 152 2992 161
rect 2943 142 2992 152
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2915 120 2989 136
rect 3007 128 3037 184
rect 3072 174 3280 184
rect 3315 180 3360 184
rect 3363 183 3364 184
rect 3379 183 3392 184
rect 3239 170 3287 174
rect 3122 148 3152 157
rect 3215 150 3230 157
rect 3251 148 3287 170
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 2915 118 2928 120
rect 2943 118 2977 120
rect 2915 102 2989 118
rect 3016 114 3029 128
rect 3044 114 3060 130
rect 3106 125 3117 138
rect 2899 80 2900 96
rect 2915 80 2928 102
rect 2943 80 2973 102
rect 3016 98 3078 114
rect 3106 107 3117 123
rect 3122 118 3132 138
rect 3142 118 3156 138
rect 3159 125 3168 138
rect 3184 125 3193 138
rect 3122 107 3156 118
rect 3159 107 3167 123
rect 3184 107 3193 123
rect 3200 118 3210 138
rect 3220 118 3234 138
rect 3235 125 3246 138
rect 3200 107 3234 118
rect 3235 107 3246 123
rect 3292 114 3308 130
rect 3315 128 3345 180
rect 3379 176 3380 183
rect 3364 168 3380 176
rect 3351 136 3364 155
rect 3379 136 3409 152
rect 3351 120 3425 136
rect 3351 118 3364 120
rect 3379 118 3413 120
rect 3016 96 3029 98
rect 3044 96 3078 98
rect 3016 80 3078 96
rect 3122 91 3135 94
rect 3200 91 3230 102
rect 3278 98 3324 114
rect 3351 102 3425 118
rect 3278 96 3312 98
rect 3277 80 3324 96
rect 3351 80 3364 102
rect 3379 80 3409 102
rect 3436 80 3437 96
rect 3452 80 3465 240
rect 3495 136 3508 240
rect 3553 218 3554 228
rect 3569 218 3582 228
rect 3553 214 3582 218
rect 3587 214 3617 240
rect 3635 226 3651 228
rect 3723 226 3776 240
rect 3724 224 3788 226
rect 3635 214 3650 218
rect 3553 212 3650 214
rect 3537 204 3588 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3619 204 3669 212
rect 3619 196 3635 204
rect 3642 202 3669 204
rect 3678 204 3693 208
rect 3740 204 3772 224
rect 3831 212 3846 240
rect 3895 237 3925 240
rect 3895 234 3931 237
rect 3861 226 3877 228
rect 3862 214 3877 218
rect 3895 215 3934 234
rect 3953 228 3960 229
rect 3959 221 3960 228
rect 3943 218 3944 221
rect 3959 218 3972 221
rect 3895 214 3925 215
rect 3934 214 3940 215
rect 3943 214 3972 218
rect 3862 213 3972 214
rect 3862 212 3978 213
rect 3831 204 3899 212
rect 3678 202 3747 204
rect 3765 202 3899 204
rect 3642 198 3714 202
rect 3642 196 3767 198
rect 3642 192 3714 196
rect 3537 184 3588 192
rect 3635 188 3714 192
rect 3795 188 3899 202
rect 3928 204 3978 212
rect 3928 195 3944 204
rect 3635 184 3899 188
rect 3925 192 3944 195
rect 3951 192 3978 204
rect 3925 184 3978 192
rect 3553 176 3554 184
rect 3569 176 3582 184
rect 3553 168 3569 176
rect 3550 161 3569 164
rect 3550 152 3572 161
rect 3523 142 3572 152
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3495 120 3569 136
rect 3587 128 3617 184
rect 3652 174 3860 184
rect 3895 180 3940 184
rect 3943 183 3944 184
rect 3959 183 3972 184
rect 3819 170 3867 174
rect 3702 148 3732 157
rect 3795 150 3810 157
rect 3831 148 3867 170
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3495 118 3508 120
rect 3523 118 3557 120
rect 3495 102 3569 118
rect 3596 114 3609 128
rect 3624 114 3640 130
rect 3686 125 3697 138
rect 3479 80 3480 96
rect 3495 80 3508 102
rect 3523 80 3553 102
rect 3596 98 3658 114
rect 3686 107 3697 123
rect 3702 118 3712 138
rect 3722 118 3736 138
rect 3739 125 3748 138
rect 3764 125 3773 138
rect 3702 107 3736 118
rect 3739 107 3747 123
rect 3764 107 3773 123
rect 3780 118 3790 138
rect 3800 118 3814 138
rect 3815 125 3826 138
rect 3780 107 3814 118
rect 3815 107 3826 123
rect 3872 114 3888 130
rect 3895 128 3925 180
rect 3959 176 3960 183
rect 3944 168 3960 176
rect 3931 136 3944 155
rect 3959 136 3989 152
rect 3931 120 4005 136
rect 3931 118 3944 120
rect 3959 118 3993 120
rect 3596 96 3609 98
rect 3624 96 3658 98
rect 3596 80 3658 96
rect 3702 91 3715 94
rect 3780 91 3810 102
rect 3858 98 3904 114
rect 3931 102 4005 118
rect 3858 96 3892 98
rect 3857 80 3904 96
rect 3931 80 3944 102
rect 3959 80 3989 102
rect 4016 80 4017 96
rect 4032 80 4045 240
rect 4075 136 4088 240
rect 4133 218 4134 228
rect 4149 218 4162 228
rect 4133 214 4162 218
rect 4167 214 4197 240
rect 4215 226 4231 228
rect 4303 226 4356 240
rect 4304 224 4368 226
rect 4215 214 4230 218
rect 4133 212 4230 214
rect 4117 204 4168 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4199 204 4249 212
rect 4199 196 4215 204
rect 4222 202 4249 204
rect 4258 204 4273 208
rect 4320 204 4352 224
rect 4411 212 4426 240
rect 4475 237 4505 240
rect 4475 234 4511 237
rect 4441 226 4457 228
rect 4442 214 4457 218
rect 4475 215 4514 234
rect 4533 228 4540 229
rect 4539 221 4540 228
rect 4523 218 4524 221
rect 4539 218 4552 221
rect 4475 214 4505 215
rect 4514 214 4520 215
rect 4523 214 4552 218
rect 4442 213 4552 214
rect 4442 212 4558 213
rect 4411 204 4479 212
rect 4258 202 4327 204
rect 4345 202 4479 204
rect 4222 198 4294 202
rect 4222 196 4347 198
rect 4222 192 4294 196
rect 4117 184 4168 192
rect 4215 188 4294 192
rect 4375 188 4479 202
rect 4508 204 4558 212
rect 4508 195 4524 204
rect 4215 184 4479 188
rect 4505 192 4524 195
rect 4531 192 4558 204
rect 4505 184 4558 192
rect 4133 176 4134 184
rect 4149 176 4162 184
rect 4133 168 4149 176
rect 4130 161 4149 164
rect 4130 152 4152 161
rect 4103 142 4152 152
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4075 120 4149 136
rect 4167 128 4197 184
rect 4232 174 4440 184
rect 4475 180 4520 184
rect 4523 183 4524 184
rect 4539 183 4552 184
rect 4399 170 4447 174
rect 4282 148 4312 157
rect 4375 150 4390 157
rect 4411 148 4447 170
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4075 118 4088 120
rect 4103 118 4137 120
rect 4075 102 4149 118
rect 4176 114 4189 128
rect 4204 114 4220 130
rect 4266 125 4277 138
rect 4059 80 4060 96
rect 4075 80 4088 102
rect 4103 80 4133 102
rect 4176 98 4238 114
rect 4266 107 4277 123
rect 4282 118 4292 138
rect 4302 118 4316 138
rect 4319 125 4328 138
rect 4344 125 4353 138
rect 4282 107 4316 118
rect 4319 107 4327 123
rect 4344 107 4353 123
rect 4360 118 4370 138
rect 4380 118 4394 138
rect 4395 125 4406 138
rect 4360 107 4394 118
rect 4395 107 4406 123
rect 4452 114 4468 130
rect 4475 128 4505 180
rect 4539 176 4540 183
rect 4524 168 4540 176
rect 4511 136 4524 155
rect 4539 136 4569 152
rect 4511 120 4585 136
rect 4511 118 4524 120
rect 4539 118 4573 120
rect 4176 96 4189 98
rect 4204 96 4238 98
rect 4176 80 4238 96
rect 4282 91 4295 94
rect 4360 91 4390 102
rect 4438 98 4484 114
rect 4511 102 4585 118
rect 4438 96 4472 98
rect 4437 80 4484 96
rect 4511 80 4524 102
rect 4539 80 4569 102
rect 4596 80 4597 96
rect 4612 80 4625 240
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 160 80
rect 172 68 247 80
rect 305 68 380 80
rect 392 68 423 80
rect 429 68 464 80
rect 98 66 260 68
rect -7 38 34 46
rect 116 38 129 66
rect 144 64 159 66
rect 183 39 190 46
rect 193 38 260 66
rect 292 66 464 68
rect 262 44 290 48
rect 292 44 372 66
rect 393 64 408 66
rect 262 42 372 44
rect 262 38 290 42
rect 292 38 372 42
rect -1 28 0 38
rect 15 28 28 38
rect 43 28 73 38
rect 116 28 159 38
rect 166 28 174 38
rect 193 30 196 38
rect 260 30 292 38
rect 193 28 359 30
rect 378 28 389 38
rect 393 28 423 38
rect 451 28 464 66
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 740 80
rect 752 68 827 80
rect 885 68 960 80
rect 972 68 1003 80
rect 1009 68 1044 80
rect 678 66 840 68
rect 573 38 614 46
rect 696 38 709 66
rect 724 64 739 66
rect 763 39 770 46
rect 773 38 840 66
rect 872 66 1044 68
rect 842 44 870 48
rect 872 44 952 66
rect 973 64 988 66
rect 842 42 952 44
rect 842 38 870 42
rect 872 38 952 42
rect 479 28 509 38
rect 536 28 537 38
rect 552 28 565 38
rect 579 28 580 38
rect 595 28 608 38
rect 623 28 653 38
rect 696 28 739 38
rect 746 28 754 38
rect 773 30 776 38
rect 840 30 872 38
rect 773 28 939 30
rect 958 28 969 38
rect 973 28 1003 38
rect 1031 28 1044 66
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1320 80
rect 1332 68 1407 80
rect 1465 68 1540 80
rect 1552 68 1583 80
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1153 38 1194 46
rect 1276 38 1289 66
rect 1304 64 1319 66
rect 1343 39 1350 46
rect 1353 38 1420 66
rect 1452 66 1624 68
rect 1422 44 1450 48
rect 1452 44 1532 66
rect 1553 64 1568 66
rect 1422 42 1532 44
rect 1422 38 1450 42
rect 1452 38 1532 42
rect 1059 28 1089 38
rect 1116 28 1117 38
rect 1132 28 1145 38
rect 1159 28 1160 38
rect 1175 28 1188 38
rect 1203 28 1233 38
rect 1276 28 1319 38
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1420 30 1452 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1553 28 1583 38
rect 1611 28 1624 66
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1900 80
rect 1912 68 1987 80
rect 2045 68 2120 80
rect 2132 68 2163 80
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1733 38 1774 46
rect 1856 38 1869 66
rect 1884 64 1899 66
rect 1923 39 1930 46
rect 1933 38 2000 66
rect 2032 66 2204 68
rect 2002 44 2030 48
rect 2032 44 2112 66
rect 2133 64 2148 66
rect 2002 42 2112 44
rect 2002 38 2030 42
rect 2032 38 2112 42
rect 1639 28 1669 38
rect 1696 28 1697 38
rect 1712 28 1725 38
rect 1739 28 1740 38
rect 1755 28 1768 38
rect 1783 28 1813 38
rect 1856 28 1899 38
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 2000 30 2032 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2133 28 2163 38
rect 2191 28 2204 66
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2480 80
rect 2492 68 2567 80
rect 2625 68 2700 80
rect 2712 68 2743 80
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2313 38 2354 46
rect 2436 38 2449 66
rect 2464 64 2479 66
rect 2503 39 2510 46
rect 2513 38 2580 66
rect 2612 66 2784 68
rect 2582 44 2610 48
rect 2612 44 2692 66
rect 2713 64 2728 66
rect 2582 42 2692 44
rect 2582 38 2610 42
rect 2612 38 2692 42
rect 2219 28 2249 38
rect 2276 28 2277 38
rect 2292 28 2305 38
rect 2319 28 2320 38
rect 2335 28 2348 38
rect 2363 28 2393 38
rect 2436 28 2479 38
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2580 30 2612 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2713 28 2743 38
rect 2771 28 2784 66
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3060 80
rect 3072 68 3147 80
rect 3205 68 3280 80
rect 3292 68 3323 80
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 2893 38 2934 46
rect 3016 38 3029 66
rect 3044 64 3059 66
rect 3083 39 3090 46
rect 3093 38 3160 66
rect 3192 66 3364 68
rect 3162 44 3190 48
rect 3192 44 3272 66
rect 3293 64 3308 66
rect 3162 42 3272 44
rect 3162 38 3190 42
rect 3192 38 3272 42
rect 2799 28 2829 38
rect 2856 28 2857 38
rect 2872 28 2885 38
rect 2899 28 2900 38
rect 2915 28 2928 38
rect 2943 28 2973 38
rect 3016 28 3059 38
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3160 30 3192 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3293 28 3323 38
rect 3351 28 3364 66
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3640 80
rect 3652 68 3727 80
rect 3785 68 3860 80
rect 3872 68 3903 80
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3473 38 3514 46
rect 3596 38 3609 66
rect 3624 64 3639 66
rect 3663 39 3670 46
rect 3673 38 3740 66
rect 3772 66 3944 68
rect 3742 44 3770 48
rect 3772 44 3852 66
rect 3873 64 3888 66
rect 3742 42 3852 44
rect 3742 38 3770 42
rect 3772 38 3852 42
rect 3379 28 3409 38
rect 3436 28 3437 38
rect 3452 28 3465 38
rect 3479 28 3480 38
rect 3495 28 3508 38
rect 3523 28 3553 38
rect 3596 28 3639 38
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3740 30 3772 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3873 28 3903 38
rect 3931 28 3944 66
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4220 80
rect 4232 68 4307 80
rect 4365 68 4440 80
rect 4452 68 4483 80
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4053 38 4094 46
rect 4176 38 4189 66
rect 4204 64 4219 66
rect 4243 39 4250 46
rect 4253 38 4320 66
rect 4352 66 4524 68
rect 4322 44 4350 48
rect 4352 44 4432 66
rect 4453 64 4468 66
rect 4322 42 4432 44
rect 4322 38 4350 42
rect 4352 38 4432 42
rect 3959 28 3989 38
rect 4016 28 4017 38
rect 4032 28 4045 38
rect 4059 28 4060 38
rect 4075 28 4088 38
rect 4103 28 4133 38
rect 4176 28 4219 38
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4320 30 4352 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4453 28 4483 38
rect 4511 28 4524 66
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4539 28 4569 38
rect 4596 28 4597 38
rect 4612 28 4625 38
rect -1 22 4625 28
rect 0 14 4625 22
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 129 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 243 0 294 1
rect 451 0 464 14
rect 244 -2 308 0
rect 479 -4 509 14
rect 552 0 565 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 709 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 823 0 874 1
rect 1031 0 1044 14
rect 824 -2 888 0
rect 1059 -4 1089 14
rect 1132 0 1145 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1289 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1403 0 1454 1
rect 1611 0 1624 14
rect 1404 -2 1468 0
rect 1639 -4 1669 14
rect 1712 0 1725 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1869 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1983 0 2034 1
rect 2191 0 2204 14
rect 1984 -2 2048 0
rect 2219 -4 2249 14
rect 2292 0 2305 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2449 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2563 0 2614 1
rect 2771 0 2784 14
rect 2564 -2 2628 0
rect 2799 -4 2829 14
rect 2872 0 2885 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3029 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3143 0 3194 1
rect 3351 0 3364 14
rect 3144 -2 3208 0
rect 3379 -4 3409 14
rect 3452 0 3465 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3609 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3723 0 3774 1
rect 3931 0 3944 14
rect 3724 -2 3788 0
rect 3959 -4 3989 14
rect 4032 0 4045 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4189 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4303 0 4354 1
rect 4511 0 4524 14
rect 4304 -2 4368 0
rect 4539 -4 4569 14
rect 4612 0 4625 14
<< pwell >>
rect 74 184 89 212
rect 464 184 479 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
<< ndiffc >>
rect 74 184 89 212
rect 464 184 479 213
rect 654 184 669 212
rect 1044 184 1059 213
rect 1234 184 1249 212
rect 1624 184 1639 213
rect 1814 184 1829 212
rect 2204 184 2219 213
rect 2394 184 2409 212
rect 2784 184 2799 213
rect 2974 184 2989 212
rect 3364 184 3379 213
rect 3554 184 3569 212
rect 3944 184 3959 213
rect 4134 184 4149 212
rect 4524 184 4539 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 1117 38 1132 80
rect 1160 38 1175 80
rect 1697 38 1712 80
rect 1740 38 1755 80
rect 2277 38 2292 80
rect 2320 38 2335 80
rect 2857 38 2872 80
rect 2900 38 2915 80
rect 3437 38 3452 80
rect 3480 38 3495 80
rect 4017 38 4032 80
rect 4060 38 4075 80
rect 4597 38 4612 80
<< poly >>
rect 0 4290 30 4320
rect 0 4020 30 4050
rect 0 3750 30 3780
rect 0 3480 30 3510
rect 0 3210 30 3240
rect 0 2940 30 2970
rect 0 2670 30 2700
rect 0 2400 30 2430
rect 0 2130 30 2160
rect 0 1860 30 1890
rect 0 1590 30 1620
rect 0 1320 30 1350
rect 0 1050 30 1080
rect 0 780 30 810
rect 0 510 30 540
rect 0 240 30 270
<< metal1 >>
rect 0 4276 15 4290
rect 0 4152 15 4186
rect 0 4050 15 4064
rect 0 4006 15 4020
rect 0 3882 15 3916
rect 0 3780 15 3794
rect 0 3736 15 3750
rect 0 3612 15 3646
rect 0 3510 15 3524
rect 0 3466 15 3480
rect 0 3342 15 3376
rect 0 3240 15 3254
rect 0 3196 15 3210
rect 0 3072 15 3106
rect 0 2970 15 2984
rect 0 2926 15 2940
rect 0 2802 15 2836
rect 0 2700 15 2714
rect 0 2656 15 2670
rect 0 2532 15 2566
rect 0 2430 15 2444
rect 0 2386 15 2400
rect 0 2262 15 2296
rect 0 2160 15 2174
rect 0 2116 15 2130
rect 0 1992 15 2026
rect 0 1890 15 1904
rect 0 1846 15 1860
rect 0 1722 15 1756
rect 0 1620 15 1634
rect 0 1576 15 1590
rect 0 1452 15 1486
rect 0 1350 15 1364
rect 0 1306 15 1320
rect 0 1182 15 1216
rect 0 1080 15 1094
rect 0 1036 15 1050
rect 0 912 15 946
rect 0 810 15 824
rect 0 766 15 780
rect 0 642 15 676
rect 0 540 15 554
rect 0 496 15 510
rect 0 372 15 406
rect 0 270 15 284
rect 0 226 15 240
rect 0 102 15 136
rect 0 0 15 14
use 10T_1x8_magic  10T_1x8_magic_8
timestamp 1656019537
transform 1 0 0 0 1 270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_9
timestamp 1656019537
transform 1 0 0 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_10
timestamp 1656019537
transform 1 0 0 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_11
timestamp 1656019537
transform 1 0 0 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_12
timestamp 1656019537
transform 1 0 0 0 1 1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_13
timestamp 1656019537
transform 1 0 0 0 1 1350
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_14
timestamp 1656019537
transform 1 0 0 0 1 1890
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_15
timestamp 1656019537
transform 1 0 0 0 1 1620
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1656019537
transform 1 0 0 0 1 2430
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1656019537
transform 1 0 0 0 1 2160
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1656019537
transform 1 0 0 0 1 2700
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1656019537
transform 1 0 0 0 1 2970
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1656019537
transform 1 0 0 0 1 3510
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1656019537
transform 1 0 0 0 1 3240
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1656019537
transform 1 0 0 0 1 4050
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1656019537
transform 1 0 0 0 1 3780
box -7 -4 4631 312
<< labels >>
rlabel metal1 0 4152 15 4186 1 RWL_0
port 34 ew signal input
rlabel poly 0 4020 30 4050 1 WWL_1
port 35 ew signal input
rlabel metal1 0 3882 15 3916 1 RWL_1
port 36 ew signal input
rlabel poly 0 3750 30 3780 1 WWL_2
port 37 ew signal input
rlabel metal1 0 3612 15 3646 1 RWL_2
port 38 ew signal input
rlabel poly 0 3480 30 3510 1 WWL_3
port 39 ew signal input
rlabel metal1 0 3342 15 3376 1 RWL_3
port 40 ew signal input
rlabel poly 0 3210 30 3240 1 WWL_4
port 41 ew signal input
rlabel metal1 0 3072 15 3106 1 RWL_4
port 42 ew signal input
rlabel poly 0 2940 30 2970 1 WWL_5
port 43 ew signal input
rlabel metal1 0 2802 15 2836 1 RWL_5
port 44 ew signal input
rlabel poly 0 2670 30 2700 1 WWL_6
port 45 ew signal input
rlabel metal1 0 2532 15 2566 1 RWL_6
port 46 ew signal input
rlabel poly 0 2400 30 2430 1 WWL_7
port 47 ew signal input
rlabel metal1 0 2262 15 2296 1 RWL_7
port 48 ew signal input
rlabel metal1 0 4276 15 4290 1 VDD
port 65 ew power bidirectional abutment
rlabel metal1 0 4050 15 4064 1 GND
port 66 ew ground bidirectional abutment
rlabel metal1 0 3736 15 3750 1 VDD
rlabel metal1 0 3466 15 3480 1 VDD
rlabel metal1 0 4006 15 4020 1 VDD
rlabel metal1 0 3196 15 3210 1 VDD
rlabel metal1 0 2656 15 2670 1 VDD
rlabel metal1 0 2386 15 2400 1 VDD
rlabel metal1 0 2926 15 2940 1 VDD
rlabel metal1 0 3240 15 3254 1 GND
rlabel metal1 0 3510 15 3524 1 GND
rlabel metal1 0 3780 15 3794 1 GND
rlabel metal1 0 2970 15 2984 1 GND
rlabel metal1 0 2160 15 2174 1 GND
rlabel metal1 0 2430 15 2444 1 GND
rlabel metal1 0 2700 15 2714 1 GND
rlabel poly 0 4290 30 4320 1 WWL_0
port 33 ew signal input
rlabel metal1 0 540 15 554 1 GND
rlabel metal1 0 270 15 284 1 GND
rlabel metal1 0 0 15 14 1 GND
rlabel metal1 0 810 15 824 1 GND
rlabel metal1 0 1620 15 1634 1 GND
rlabel metal1 0 1350 15 1364 1 GND
rlabel metal1 0 1080 15 1094 1 GND
rlabel metal1 0 766 15 780 1 VDD
rlabel metal1 0 226 15 240 1 VDD
rlabel metal1 0 496 15 510 1 VDD
rlabel metal1 0 1036 15 1050 1 VDD
rlabel metal1 0 1846 15 1860 1 VDD
rlabel metal1 0 1306 15 1320 1 VDD
rlabel metal1 0 1576 15 1590 1 VDD
rlabel metal1 0 1890 15 1904 1 GND
rlabel metal1 0 2116 15 2130 1 VDD
rlabel locali 4134 184 4149 212 1 WBLb_7
port 32 ns signal input
rlabel locali 4524 184 4539 213 1 WBL_7
port 31 ns signal input
rlabel locali 3554 184 3569 212 1 WBLb_6
port 30 ns signal input
rlabel locali 3944 184 3959 213 1 WBL_6
port 29 ns signal input
rlabel locali 2974 184 2989 212 1 WBLb_5
port 28 ns signal input
rlabel locali 3364 184 3379 213 1 WBL_5
port 27 ns signal input
rlabel locali 2394 184 2409 212 1 WBLb_4
port 26 ns signal input
rlabel locali 2784 184 2799 213 1 WBL_4
port 25 ns signal input
rlabel locali 1814 184 1829 212 1 WBLb_3
port 24 ns signal input
rlabel locali 2204 184 2219 213 1 WBL_3
port 23 ns signal input
rlabel locali 1234 184 1249 212 1 WBLb_2
port 22 ns signal input
rlabel locali 1624 184 1639 213 1 WBL_2
port 21 ns signal input
rlabel locali 654 184 669 212 1 WBLb_1
port 20 ns signal input
rlabel locali 1044 184 1059 213 1 WBL_1
port 19 ns signal input
rlabel locali 74 184 89 212 1 WBLb_0
port 18 ns signal input
rlabel locali 464 184 479 213 1 WBL_0
port 17 ns signal input
rlabel locali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel locali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel locali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel locali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel locali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel locali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel locali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel locali 2320 38 2335 80 1 RBL1_4
port 9 ns signal output
rlabel locali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel locali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel locali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel locali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel locali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel locali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel locali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel locali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel poly 0 2130 30 2160 1 WWL_8
port 49 ew signal input
rlabel metal1 0 1992 15 2026 1 RWL_8
port 50 ew signal input
rlabel poly 0 1860 30 1890 1 WWL_9
port 51 ew signal input
rlabel metal1 0 1722 15 1756 1 RWL_9
port 52 ew signal input
rlabel poly 0 1590 30 1620 1 WWL_10
port 53 ew signal input
rlabel metal1 0 1452 15 1486 1 RWL_10
port 54 ew signal input
rlabel poly 0 1320 30 1350 1 WWL_11
port 55 ew signal input
rlabel metal1 0 1182 15 1216 1 RWL_11
port 56 ew signal input
rlabel poly 0 1050 30 1080 1 WWL_12
port 57 ew signal input
rlabel metal1 0 912 15 946 1 RWL_12
port 58 ew signal input
rlabel poly 0 780 30 810 1 WWL_13
port 59 ew signal input
rlabel metal1 0 642 15 676 1 RWL_13
port 60 ew signal input
rlabel poly 0 510 30 540 1 WWL_14
port 61 ew signal input
rlabel metal1 0 372 15 406 1 RWL_14
port 62 ew signal input
rlabel poly 0 240 30 270 1 WWL_15
port 63 ew signal input
rlabel metal1 0 102 15 136 1 RWL_15
port 64 ew signal input
<< end >>
