* FILE: 10T-toy.sp

********************** begin header *****************************

* SPICE Header file for TSMC 3.3 0.35 process (scn4me_subm)

.OPTIONS post NOMOD probe measout captab 

**################################################
* Only Typical/Typical spice models included
.include '/programs/micromagic/mmi_local/ami05.mod'
**################################################

.param ln_min   =  0.4u
.param lp_min   =  0.4u

.PARAM vddp=3.30	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 25
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "10T-toy" generated by MMI_SUE5.6.37 on Sat Nov 13 
*+ 12:31:23 CST 2021.

.SUBCKT invM A1 O 
M_1 O A1 Vdd vdd p W='0.14*1u' L='0.15*1u' 
M_2 O A1 Gnd gnd n W='0.21*1u' L='0.15*1u' 
.ENDS	$ invM

* start main CELL 10T-toy
* .SUBCKT 10T-toy BL BLb WL1 WL2 
XinvM net_2 net_1 invM 
M_1 net_2 WL1 BL gnd n W='0.14*1u' L='0.15*1u' 
M_2 BLb WL2 net_1 gnd n W='0.14*1u' L='0.15*1u' 
M_3 net_3 uc_net_4 uc_net_7 gnd n W='0.14*1u' L='0.025*1u' 
M_4 gnd net_2 net_3 gnd n W='0.42*1u' L='0.15*1u' 
M_5 uc_net_5 uc_net_8 net_6 gnd n W='0.14*1u' L='0.025*1u' 
M_6 net_6 net_1 gnd gnd n W='0.42*1u' L='0.15*1u' 
XInv net_1 net_2 invM 
* .ENDS	$ 10T-toy

.GLOBAL gnd vdd

.END

