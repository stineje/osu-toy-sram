magic
tech sky130A
magscale 1 2
timestamp 1652384410
<< error_p >>
rect 38 329 66 342
rect 14 316 226 329
rect 22 308 82 316
rect 22 307 46 308
rect 58 307 82 308
rect 14 301 226 307
rect 22 300 82 301
rect -18 273 16 292
rect 66 273 68 300
rect 138 293 148 301
rect 138 292 228 293
rect 138 273 148 292
rect -18 267 226 273
rect -18 262 16 267
rect 38 262 68 267
rect 38 254 80 262
rect 138 255 148 267
rect 174 255 204 267
rect 22 247 46 254
rect 52 251 82 254
rect 144 251 148 255
rect 158 251 218 255
rect 52 249 218 251
rect 58 247 218 249
rect 22 245 218 247
rect 22 237 86 245
rect 22 230 87 237
rect 22 225 71 230
rect 14 220 71 225
rect 107 221 141 228
rect 144 221 148 245
rect 158 225 218 245
rect 158 221 226 225
rect 14 219 61 220
rect -4 191 16 212
rect 38 204 61 219
rect 107 217 148 221
rect 63 212 148 217
rect 170 219 226 221
rect -4 182 28 191
rect 63 185 157 212
rect 91 182 157 185
rect 170 205 204 219
rect 240 212 312 316
rect 170 182 188 205
rect -2 174 28 182
rect -2 167 38 174
rect -2 149 34 167
rect -2 142 38 149
rect -2 134 28 142
rect -4 125 28 134
rect -4 104 16 125
rect 42 112 48 174
rect 70 161 96 175
rect 107 166 148 182
rect 68 149 96 161
rect 138 150 148 166
rect 170 159 180 182
rect 68 112 70 149
rect 107 141 148 150
rect 160 149 180 159
rect 152 147 180 149
rect 152 141 170 147
rect 172 142 180 147
rect 102 134 148 141
rect 174 134 180 142
rect 38 106 70 112
rect 91 131 157 134
rect 174 131 188 134
rect 189 131 198 205
rect 202 174 204 205
rect 224 175 312 212
rect 223 174 312 175
rect 202 167 312 174
rect 204 149 312 167
rect 91 119 198 131
rect 202 142 312 149
rect 38 104 80 106
rect 91 104 170 119
rect 38 97 70 104
rect 102 99 170 104
rect 174 111 188 119
rect 202 111 204 142
rect 223 141 312 142
rect 14 96 70 97
rect 14 91 46 96
rect 22 71 46 91
rect 68 87 70 96
rect 107 88 148 99
rect 58 79 70 87
rect 138 83 148 88
rect 174 97 204 111
rect 224 104 312 141
rect 174 91 226 97
rect 174 83 218 91
rect 144 79 148 83
rect 58 71 82 79
rect 158 71 218 83
rect 22 65 218 71
rect 22 62 82 65
rect 38 54 80 62
rect 158 61 218 65
rect -18 49 16 54
rect 38 49 68 54
rect 138 49 144 61
rect 174 49 204 61
rect -18 43 226 49
rect -18 28 16 43
rect 66 34 68 43
rect 38 28 68 34
rect 138 28 144 43
rect -18 24 226 28
rect 14 23 228 24
rect 14 9 226 23
rect 22 8 46 9
rect 58 8 82 9
rect 22 -1 82 8
rect 240 0 312 104
rect 38 -26 66 -1
<< nwell >>
rect 144 0 240 316
<< pwell >>
rect 12 263 92 342
rect 12 200 106 263
rect -26 116 106 200
rect 12 53 106 116
rect 12 -26 92 53
<< npd >>
rect 38 182 80 212
rect 38 104 80 134
<< npass >>
rect 38 262 66 292
rect 38 24 66 54
<< ppu >>
rect 174 262 202 267
rect 174 182 202 212
rect 174 104 202 134
rect 174 49 202 54
<< ndiff >>
rect 38 292 66 301
rect 38 254 66 262
tri 61 220 71 230 se
rect 71 220 80 237
rect 38 212 80 220
rect 38 174 80 182
rect 14 142 80 174
rect 38 134 80 142
rect 38 96 80 104
rect 70 79 80 96
rect 38 54 66 62
rect 38 15 66 24
<< pdiff >>
rect 174 255 202 262
rect 174 212 202 221
rect 174 174 202 182
rect 174 142 226 174
rect 174 134 202 142
rect 174 95 202 104
tri 174 83 186 95 nw
rect 174 54 202 61
<< ndiffc >>
rect 38 301 66 316
rect 38 237 66 254
rect 38 230 71 237
rect 38 220 61 230
tri 61 220 71 230 nw
rect 0 142 14 174
rect 38 79 70 96
rect 38 62 66 79
rect 38 0 66 15
<< pdiffc >>
rect 174 221 202 255
rect 226 142 240 174
tri 174 83 186 95 se
rect 186 83 202 95
rect 174 61 202 83
<< poly >>
rect 16 262 38 292
rect 66 267 240 292
rect 66 262 174 267
rect 202 262 240 267
rect 16 182 38 212
rect 80 182 107 212
rect 141 182 174 212
rect 202 182 224 212
rect 16 104 38 134
rect 80 104 107 134
rect 141 104 174 134
rect 202 104 224 134
rect 16 24 38 54
rect 66 49 174 54
rect 202 49 240 54
rect 66 24 240 49
<< polycont >>
rect 107 182 141 212
rect 107 104 141 134
<< corelocali >>
rect 14 301 38 316
rect 66 301 226 316
rect 14 255 226 273
rect 14 254 174 255
rect 14 220 38 254
rect 66 245 174 254
rect 66 237 71 245
tri 71 230 86 245 nw
rect 170 221 174 245
rect 202 221 226 255
rect 14 219 60 220
tri 60 219 61 220 nw
rect 170 219 226 221
rect 0 174 14 191
tri 63 182 98 217 se
rect 98 212 142 217
rect 98 182 107 212
rect 141 182 142 212
rect 0 125 14 142
tri 42 161 63 182 se
rect 63 175 142 182
rect 63 161 70 175
rect 42 97 70 161
tri 70 149 96 175 nw
tri 160 149 170 159 se
rect 170 149 198 219
rect 226 175 240 191
tri 152 141 160 149 se
rect 160 147 198 149
rect 160 141 170 147
rect 102 134 170 141
rect 102 104 107 134
rect 141 119 170 134
tri 170 119 198 147 nw
rect 226 125 240 141
rect 141 104 150 119
rect 102 99 150 104
tri 150 99 170 119 nw
rect 14 96 70 97
rect 14 62 38 96
tri 186 95 188 97 se
rect 188 95 226 97
rect 66 71 70 79
tri 162 71 174 83 se
rect 66 62 174 71
rect 14 61 174 62
rect 202 61 226 95
rect 14 43 226 61
rect 14 0 38 15
rect 66 0 226 15
<< viali >>
rect 223 174 240 175
rect 223 142 226 174
rect 226 142 240 174
rect 223 141 240 142
<< labels >>
rlabel corelocali 107 182 141 212 1 left_net
rlabel corelocali 107 104 141 134 1 right_net

rlabel poly 16 262 240 292 1 WL2
port 1 nsew signal input
rlabel poly 16 24 240 54 1 WL1
port 2 nsew signal input
rlabel corelocali 14 0 226 15 1 bit_v
port 3 nsew signal bidirectional
rlabel corelocali 14 301 226 316 1 bit_b_v
port 4 nsew signal bidirectional
rlabel corelocali 226 125 240 191 1 VPWR
port 5 nsew power bidirectional
rlabel corelocali 0 125 14 191 1 VGND
port 5 nsew ground bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
