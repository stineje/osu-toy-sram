* FILE: 10tcell.sp

********************** begin header *****************************

* SPICE Header file for TSMC 3.3 0.35 process (scn4me_subm)

.OPTIONS post NOMOD probe measout captab 

**################################################
* Only Typical/Typical spice models included
.include '/programs/micromagic/mmi_local/ami05.mod'
**################################################

.param ln_min   =  0.4u
.param lp_min   =  0.4u

.PARAM vddp=3.30	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 25
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "10tcell" generated by MMI_SUE5.6.37 on Fri Nov 12 
*+ 13:58:31 CST 2021.

* start main CELL 10tcell
* .SUBCKT 10tcell  
M_1 net_3 net_7 uc_net_9 gnd n W='0.42*1u' L='0.15*1u' 
M_2 net_8 net_2 net_3 gnd n W='0.42*1u' L='0.15*1u' 
M_3 net_4 net_2 net_5 gnd n W='0.42*1u' L='0.15*1u' 
M_4 uc_net_6 net_7 net_4 gnd n W='0.42*1u' L='0.15*1u' 
M_5 net_10 net_8 net_3 gnd n W='0.42*1u' L='0.15*1u' 
M_6 net_4 net_5 net_10 gnd n W='0.42*1u' L='0.15*1u' 
M_7 net_5 net_8 gnd gnd n W='0.42*1u' L='0.15*1u' 
M_8 gnd net_5 net_8 gnd n W='0.42*1u' L='0.15*1u' 
M_9 uc_net_1 net_8 vdd vdd p W='0.42*1u' L='0.15*1u' 
M_10 vdd net_5 net_8 vdd p W='0.42*1u' L='0.15*1u' 
* .ENDS	$ 10tcell

.GLOBAL gnd vdd

.END

