VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO toysram_16x12
  CLASS BLOCK ;
  FOREIGN toysram_16x12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.000 BY 22.000 ;
  PIN RWL0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500 1.200 2.700 2.400 ;
    END
  END RWL0[0]
  PIN RWL0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000 1.200 4.200 2.400 ;
    END
  END RWL0[1]
  PIN RWL0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.500 1.200 5.700 2.400 ;
    END
  END RWL0[2]
  PIN RWL0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.000 1.200 7.200 2.400 ;
    END
  END RWL0[3]
  PIN RWL0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.500 1.200 8.700 2.400 ;
    END
  END RWL0[4]
  PIN RWL0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.000 1.200 10.200 2.400 ;
    END
  END RWL0[5]
  PIN RWL0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500 1.200 11.700 2.400 ;
    END
  END RWL0[6]
  PIN RWL0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.000 1.200 13.200 2.400 ;
    END
  END RWL0[7]
  PIN RWL0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.500 1.200 14.700 2.400 ;
    END
  END RWL0[8]
  PIN RWL0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.000 1.200 16.200 2.400 ;
    END
  END RWL0[9]
  PIN RWL0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.500 1.200 17.700 2.400 ;
    END
  END RWL0[10]
  PIN RWL0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.000 1.200 19.200 2.400 ;
    END
  END RWL0[11]
  PIN RWL0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.500 1.200 20.700 2.400 ;
    END
  END RWL0[12]
  PIN RWL0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.000 1.200 22.200 2.400 ;
    END
  END RWL0[13]
  PIN RWL0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.500 1.200 23.700 2.400 ;
    END
  END RWL0[14]
  PIN RWL0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.000 1.200 25.200 2.400 ;
    END
  END RWL0[15]
  PIN RWL1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500 3.200 2.700 4.400 ;
    END
  END RWL1[0]
  PIN RWL1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000 3.200 4.200 4.400 ;
    END
  END RWL1[1]
  PIN RWL1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.500 3.200 5.700 4.400 ;
    END
  END RWL1[2]
  PIN RWL1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.000 3.200 7.200 4.400 ;
    END
  END RWL1[3]
  PIN RWL1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.500 3.200 8.700 4.400 ;
    END
  END RWL1[4]
  PIN RWL1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.000 3.200 10.200 4.400 ;
    END
  END RWL1[5]
  PIN RWL1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500 3.200 11.700 4.400 ;
    END
  END RWL1[6]
  PIN RWL1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.000 3.200 13.200 4.400 ;
    END
  END RWL1[7]
  PIN RWL1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.500 3.200 14.700 4.400 ;
    END
  END RWL1[8]
  PIN RWL1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.000 3.200 16.200 4.400 ;
    END
  END RWL1[9]
  PIN RWL1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.500 3.200 17.700 4.400 ;
    END
  END RWL1[10]
  PIN RWL1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.000 3.200 19.200 4.400 ;
    END
  END RWL1[11]
  PIN RWL1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.500 3.200 20.700 4.400 ;
    END
  END RWL1[12]
  PIN RWL1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.000 3.200 22.200 4.400 ;
    END
  END RWL1[13]
  PIN RWL1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.500 3.200 23.700 4.400 ;
    END
  END RWL1[14]
  PIN RWL1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.000 3.200 25.200 4.400 ;
    END
  END RWL1[15]
  PIN WWL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500 5.200 2.700 6.400 ;
    END
  END WWL[0]
  PIN WWL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.000 5.200 4.200 6.400 ;
    END
  END WWL[1]
  PIN WWL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.500 5.200 5.700 6.400 ;
    END
  END WWL[2]
  PIN WWL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.000 5.200 7.200 6.400 ;
    END
  END WWL[3]
  PIN WWL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.500 5.200 8.700 6.400 ;
    END
  END WWL[4]
  PIN WWL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.000 5.200 10.200 6.400 ;
    END
  END WWL[5]
  PIN WWL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500 5.200 11.700 6.400 ;
    END
  END WWL[6]
  PIN WWL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.000 5.200 13.200 6.400 ;
    END
  END WWL[7]
  PIN WWL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.500 5.200 14.700 6.400 ;
    END
  END WWL[8]
  PIN WWL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.000 5.200 16.200 6.400 ;
    END
  END WWL[9]
  PIN WWL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.500 5.200 17.700 6.400 ;
    END
  END WWL[10]
  PIN WWL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.000 5.200 19.200 6.400 ;
    END
  END WWL[11]
  PIN WWL[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.500 5.200 20.700 6.400 ;
    END
  END WWL[12]
  PIN WWL[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.000 5.200 22.200 6.400 ;
    END
  END WWL[13]
  PIN WWL[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.500 5.200 23.700 6.400 ;
    END
  END WWL[14]
  PIN WWL[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.000 5.200 25.200 6.400 ;
    END
  END WWL[15]
  PIN RBL0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 1.400 33.000 2.600 ;
    END
  END RBL0[0]
  PIN RBL0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 2.800 33.000 4.000 ;
    END
  END RBL0[1]
  PIN RBL0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 4.200 33.000 5.400 ;
    END
  END RBL0[2]
  PIN RBL0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 5.600 33.000 6.800 ;
    END
  END RBL0[3]
  PIN RBL0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 7.000 33.000 8.200 ;
    END
  END RBL0[4]
  PIN RBL0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 8.400 33.000 9.600 ;
    END
  END RBL0[5]
  PIN RBL0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 9.800 33.000 11.000 ;
    END
  END RBL0[6]
  PIN RBL0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 11.200 33.000 12.400 ;
    END
  END RBL0[7]
  PIN RBL0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 12.600 33.000 13.800 ;
    END
  END RBL0[8]
  PIN RBL0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 14.000 33.000 15.200 ;
    END
  END RBL0[9]
  PIN RBL0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 15.400 33.000 16.600 ;
    END
  END RBL0[10]
  PIN RBL0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 31.800 16.800 33.000 18.000 ;
    END
  END RBL0[11]
  PIN RBL1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 1.400 31.000 2.600 ;
    END
  END RBL1[0]
  PIN RBL1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 2.800 31.000 4.000 ;
    END
  END RBL1[1]
  PIN RBL1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 4.200 31.000 5.400 ;
    END
  END RBL1[2]
  PIN RBL1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 5.600 31.000 6.800 ;
    END
  END RBL1[3]
  PIN RBL1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 7.000 31.000 8.200 ;
    END
  END RBL1[4]
  PIN RBL1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 8.400 31.000 9.600 ;
    END
  END RBL1[5]
  PIN RBL1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 9.800 31.000 11.000 ;
    END
  END RBL1[6]
  PIN RBL1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 11.200 31.000 12.400 ;
    END
  END RBL1[7]
  PIN RBL1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 12.600 31.000 13.800 ;
    END
  END RBL1[8]
  PIN RBL1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 14.000 31.000 15.200 ;
    END
  END RBL1[9]
  PIN RBL1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 15.400 31.000 16.600 ;
    END
  END RBL1[10]
  PIN RBL1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.800 16.800 31.000 18.000 ;
    END
  END RBL1[11]
  PIN WBL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 1.400 29.000 2.600 ;
    END
  END WBL[0]
  PIN WBL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 2.800 29.000 4.000 ;
    END
  END WBL[1]
  PIN WBL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 4.200 29.000 5.400 ;
    END
  END WBL[2]
  PIN WBL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 5.600 29.000 6.800 ;
    END
  END WBL[3]
  PIN WBL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 7.000 29.000 8.200 ;
    END
  END WBL[4]
  PIN WBL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 8.400 29.000 9.600 ;
    END
  END WBL[5]
  PIN WBL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 9.800 29.000 11.000 ;
    END
  END WBL[6]
  PIN WBL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 11.200 29.000 12.400 ;
    END
  END WBL[7]
  PIN WBL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 12.600 29.000 13.800 ;
    END
  END WBL[8]
  PIN WBL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 14.000 29.000 15.200 ;
    END
  END WBL[9]
  PIN WBL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 15.400 29.000 16.600 ;
    END
  END WBL[10]
  PIN WBL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 27.800 16.800 29.000 18.000 ;
    END
  END WBL[11]
  PIN WBLb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 1.400 27.000 2.600 ;
    END
  END WBLb[0]
  PIN WBLb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 2.800 27.000 4.000 ;
    END
  END WBLb[1]
  PIN WBLb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 4.200 27.000 5.400 ;
    END
  END WBLb[2]
  PIN WBLb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 5.600 27.000 6.800 ;
    END
  END WBLb[3]
  PIN WBLb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 7.000 27.000 8.200 ;
    END
  END WBLb[4]
  PIN WBLb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 8.400 27.000 9.600 ;
    END
  END WBLb[5]
  PIN WBLb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 9.800 27.000 11.000 ;
    END
  END WBLb[6]
  PIN WBLb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 11.200 27.000 12.400 ;
    END
  END WBLb[7]
  PIN WBLb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 12.600 27.000 13.800 ;
    END
  END WBLb[8]
  PIN WBLb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 14.000 27.000 15.200 ;
    END
  END WBLb[9]
  PIN WBLb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 15.400 27.000 16.600 ;
    END
  END WBLb[10]
  PIN WBLb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.800 16.800 27.000 18.000 ;
    END
  END WBLb[11]
END toysram_16x12
END LIBRARY

