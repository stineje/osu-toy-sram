VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 10T_16x12_2r1w_magic_flattened
  CLASS BLOCK ;
  FOREIGN 10T_16x12_2r1w_magic_flattened ;
  ORIGIN 0.275 0.275 ;
  SIZE 35.035 BY 22.085 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 0.955 0.685 1.720 1.165 ;
        RECT 3.855 0.685 4.620 1.165 ;
        RECT 6.755 0.685 7.520 1.165 ;
        RECT 9.655 0.685 10.420 1.165 ;
        RECT 12.555 0.685 13.320 1.165 ;
        RECT 15.455 0.685 16.220 1.165 ;
        RECT 18.355 0.685 19.120 1.165 ;
        RECT 21.255 0.685 22.020 1.165 ;
        RECT 24.155 0.685 24.920 1.165 ;
        RECT 27.055 0.685 27.820 1.165 ;
        RECT 29.955 0.685 30.720 1.165 ;
        RECT 32.855 0.685 33.620 1.165 ;
      LAYER li1 ;
        RECT 1.265 1.095 1.425 1.165 ;
        RECT 4.165 1.095 4.325 1.165 ;
        RECT 7.065 1.095 7.225 1.165 ;
        RECT 9.965 1.095 10.125 1.165 ;
        RECT 12.865 1.095 13.025 1.165 ;
        RECT 15.765 1.095 15.925 1.165 ;
        RECT 18.665 1.095 18.825 1.165 ;
        RECT 21.565 1.095 21.725 1.165 ;
        RECT 24.465 1.095 24.625 1.165 ;
        RECT 27.365 1.095 27.525 1.165 ;
        RECT 30.265 1.095 30.425 1.165 ;
        RECT 33.165 1.095 33.325 1.165 ;
        RECT 1.275 1.085 1.415 1.095 ;
        RECT 4.175 1.085 4.315 1.095 ;
        RECT 7.075 1.085 7.215 1.095 ;
        RECT 9.975 1.085 10.115 1.095 ;
        RECT 12.875 1.085 13.015 1.095 ;
        RECT 15.775 1.085 15.915 1.095 ;
        RECT 18.675 1.085 18.815 1.095 ;
        RECT 21.575 1.085 21.715 1.095 ;
        RECT 24.475 1.085 24.615 1.095 ;
        RECT 27.375 1.085 27.515 1.095 ;
        RECT 30.275 1.085 30.415 1.095 ;
        RECT 33.175 1.085 33.315 1.095 ;
      LAYER met1 ;
        RECT -0.275 1.095 34.625 1.165 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 2.035 1.720 2.515 ;
        RECT 3.855 2.035 4.620 2.515 ;
        RECT 6.755 2.035 7.520 2.515 ;
        RECT 9.655 2.035 10.420 2.515 ;
        RECT 12.555 2.035 13.320 2.515 ;
        RECT 15.455 2.035 16.220 2.515 ;
        RECT 18.355 2.035 19.120 2.515 ;
        RECT 21.255 2.035 22.020 2.515 ;
        RECT 24.155 2.035 24.920 2.515 ;
        RECT 27.055 2.035 27.820 2.515 ;
        RECT 29.955 2.035 30.720 2.515 ;
        RECT 32.855 2.035 33.620 2.515 ;
      LAYER li1 ;
        RECT 1.265 2.445 1.425 2.515 ;
        RECT 4.165 2.445 4.325 2.515 ;
        RECT 7.065 2.445 7.225 2.515 ;
        RECT 9.965 2.445 10.125 2.515 ;
        RECT 12.865 2.445 13.025 2.515 ;
        RECT 15.765 2.445 15.925 2.515 ;
        RECT 18.665 2.445 18.825 2.515 ;
        RECT 21.565 2.445 21.725 2.515 ;
        RECT 24.465 2.445 24.625 2.515 ;
        RECT 27.365 2.445 27.525 2.515 ;
        RECT 30.265 2.445 30.425 2.515 ;
        RECT 33.165 2.445 33.325 2.515 ;
        RECT 1.275 2.435 1.415 2.445 ;
        RECT 4.175 2.435 4.315 2.445 ;
        RECT 7.075 2.435 7.215 2.445 ;
        RECT 9.975 2.435 10.115 2.445 ;
        RECT 12.875 2.435 13.015 2.445 ;
        RECT 15.775 2.435 15.915 2.445 ;
        RECT 18.675 2.435 18.815 2.445 ;
        RECT 21.575 2.435 21.715 2.445 ;
        RECT 24.475 2.435 24.615 2.445 ;
        RECT 27.375 2.435 27.515 2.445 ;
        RECT 30.275 2.435 30.415 2.445 ;
        RECT 33.175 2.435 33.315 2.445 ;
      LAYER met1 ;
        RECT -0.275 2.445 34.625 2.515 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 3.385 1.720 3.865 ;
        RECT 3.855 3.385 4.620 3.865 ;
        RECT 6.755 3.385 7.520 3.865 ;
        RECT 9.655 3.385 10.420 3.865 ;
        RECT 12.555 3.385 13.320 3.865 ;
        RECT 15.455 3.385 16.220 3.865 ;
        RECT 18.355 3.385 19.120 3.865 ;
        RECT 21.255 3.385 22.020 3.865 ;
        RECT 24.155 3.385 24.920 3.865 ;
        RECT 27.055 3.385 27.820 3.865 ;
        RECT 29.955 3.385 30.720 3.865 ;
        RECT 32.855 3.385 33.620 3.865 ;
      LAYER li1 ;
        RECT 1.265 3.795 1.425 3.865 ;
        RECT 4.165 3.795 4.325 3.865 ;
        RECT 7.065 3.795 7.225 3.865 ;
        RECT 9.965 3.795 10.125 3.865 ;
        RECT 12.865 3.795 13.025 3.865 ;
        RECT 15.765 3.795 15.925 3.865 ;
        RECT 18.665 3.795 18.825 3.865 ;
        RECT 21.565 3.795 21.725 3.865 ;
        RECT 24.465 3.795 24.625 3.865 ;
        RECT 27.365 3.795 27.525 3.865 ;
        RECT 30.265 3.795 30.425 3.865 ;
        RECT 33.165 3.795 33.325 3.865 ;
        RECT 1.275 3.785 1.415 3.795 ;
        RECT 4.175 3.785 4.315 3.795 ;
        RECT 7.075 3.785 7.215 3.795 ;
        RECT 9.975 3.785 10.115 3.795 ;
        RECT 12.875 3.785 13.015 3.795 ;
        RECT 15.775 3.785 15.915 3.795 ;
        RECT 18.675 3.785 18.815 3.795 ;
        RECT 21.575 3.785 21.715 3.795 ;
        RECT 24.475 3.785 24.615 3.795 ;
        RECT 27.375 3.785 27.515 3.795 ;
        RECT 30.275 3.785 30.415 3.795 ;
        RECT 33.175 3.785 33.315 3.795 ;
      LAYER met1 ;
        RECT -0.275 3.795 34.625 3.865 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 4.735 1.720 5.215 ;
        RECT 3.855 4.735 4.620 5.215 ;
        RECT 6.755 4.735 7.520 5.215 ;
        RECT 9.655 4.735 10.420 5.215 ;
        RECT 12.555 4.735 13.320 5.215 ;
        RECT 15.455 4.735 16.220 5.215 ;
        RECT 18.355 4.735 19.120 5.215 ;
        RECT 21.255 4.735 22.020 5.215 ;
        RECT 24.155 4.735 24.920 5.215 ;
        RECT 27.055 4.735 27.820 5.215 ;
        RECT 29.955 4.735 30.720 5.215 ;
        RECT 32.855 4.735 33.620 5.215 ;
      LAYER li1 ;
        RECT 1.265 5.145 1.425 5.215 ;
        RECT 4.165 5.145 4.325 5.215 ;
        RECT 7.065 5.145 7.225 5.215 ;
        RECT 9.965 5.145 10.125 5.215 ;
        RECT 12.865 5.145 13.025 5.215 ;
        RECT 15.765 5.145 15.925 5.215 ;
        RECT 18.665 5.145 18.825 5.215 ;
        RECT 21.565 5.145 21.725 5.215 ;
        RECT 24.465 5.145 24.625 5.215 ;
        RECT 27.365 5.145 27.525 5.215 ;
        RECT 30.265 5.145 30.425 5.215 ;
        RECT 33.165 5.145 33.325 5.215 ;
        RECT 1.275 5.135 1.415 5.145 ;
        RECT 4.175 5.135 4.315 5.145 ;
        RECT 7.075 5.135 7.215 5.145 ;
        RECT 9.975 5.135 10.115 5.145 ;
        RECT 12.875 5.135 13.015 5.145 ;
        RECT 15.775 5.135 15.915 5.145 ;
        RECT 18.675 5.135 18.815 5.145 ;
        RECT 21.575 5.135 21.715 5.145 ;
        RECT 24.475 5.135 24.615 5.145 ;
        RECT 27.375 5.135 27.515 5.145 ;
        RECT 30.275 5.135 30.415 5.145 ;
        RECT 33.175 5.135 33.315 5.145 ;
      LAYER met1 ;
        RECT -0.275 5.145 34.625 5.215 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 6.085 1.720 6.565 ;
        RECT 3.855 6.085 4.620 6.565 ;
        RECT 6.755 6.085 7.520 6.565 ;
        RECT 9.655 6.085 10.420 6.565 ;
        RECT 12.555 6.085 13.320 6.565 ;
        RECT 15.455 6.085 16.220 6.565 ;
        RECT 18.355 6.085 19.120 6.565 ;
        RECT 21.255 6.085 22.020 6.565 ;
        RECT 24.155 6.085 24.920 6.565 ;
        RECT 27.055 6.085 27.820 6.565 ;
        RECT 29.955 6.085 30.720 6.565 ;
        RECT 32.855 6.085 33.620 6.565 ;
      LAYER li1 ;
        RECT 1.265 6.495 1.425 6.565 ;
        RECT 4.165 6.495 4.325 6.565 ;
        RECT 7.065 6.495 7.225 6.565 ;
        RECT 9.965 6.495 10.125 6.565 ;
        RECT 12.865 6.495 13.025 6.565 ;
        RECT 15.765 6.495 15.925 6.565 ;
        RECT 18.665 6.495 18.825 6.565 ;
        RECT 21.565 6.495 21.725 6.565 ;
        RECT 24.465 6.495 24.625 6.565 ;
        RECT 27.365 6.495 27.525 6.565 ;
        RECT 30.265 6.495 30.425 6.565 ;
        RECT 33.165 6.495 33.325 6.565 ;
        RECT 1.275 6.485 1.415 6.495 ;
        RECT 4.175 6.485 4.315 6.495 ;
        RECT 7.075 6.485 7.215 6.495 ;
        RECT 9.975 6.485 10.115 6.495 ;
        RECT 12.875 6.485 13.015 6.495 ;
        RECT 15.775 6.485 15.915 6.495 ;
        RECT 18.675 6.485 18.815 6.495 ;
        RECT 21.575 6.485 21.715 6.495 ;
        RECT 24.475 6.485 24.615 6.495 ;
        RECT 27.375 6.485 27.515 6.495 ;
        RECT 30.275 6.485 30.415 6.495 ;
        RECT 33.175 6.485 33.315 6.495 ;
      LAYER met1 ;
        RECT -0.275 6.495 34.625 6.565 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 7.435 1.720 7.915 ;
        RECT 3.855 7.435 4.620 7.915 ;
        RECT 6.755 7.435 7.520 7.915 ;
        RECT 9.655 7.435 10.420 7.915 ;
        RECT 12.555 7.435 13.320 7.915 ;
        RECT 15.455 7.435 16.220 7.915 ;
        RECT 18.355 7.435 19.120 7.915 ;
        RECT 21.255 7.435 22.020 7.915 ;
        RECT 24.155 7.435 24.920 7.915 ;
        RECT 27.055 7.435 27.820 7.915 ;
        RECT 29.955 7.435 30.720 7.915 ;
        RECT 32.855 7.435 33.620 7.915 ;
      LAYER li1 ;
        RECT 1.265 7.845 1.425 7.915 ;
        RECT 4.165 7.845 4.325 7.915 ;
        RECT 7.065 7.845 7.225 7.915 ;
        RECT 9.965 7.845 10.125 7.915 ;
        RECT 12.865 7.845 13.025 7.915 ;
        RECT 15.765 7.845 15.925 7.915 ;
        RECT 18.665 7.845 18.825 7.915 ;
        RECT 21.565 7.845 21.725 7.915 ;
        RECT 24.465 7.845 24.625 7.915 ;
        RECT 27.365 7.845 27.525 7.915 ;
        RECT 30.265 7.845 30.425 7.915 ;
        RECT 33.165 7.845 33.325 7.915 ;
        RECT 1.275 7.835 1.415 7.845 ;
        RECT 4.175 7.835 4.315 7.845 ;
        RECT 7.075 7.835 7.215 7.845 ;
        RECT 9.975 7.835 10.115 7.845 ;
        RECT 12.875 7.835 13.015 7.845 ;
        RECT 15.775 7.835 15.915 7.845 ;
        RECT 18.675 7.835 18.815 7.845 ;
        RECT 21.575 7.835 21.715 7.845 ;
        RECT 24.475 7.835 24.615 7.845 ;
        RECT 27.375 7.835 27.515 7.845 ;
        RECT 30.275 7.835 30.415 7.845 ;
        RECT 33.175 7.835 33.315 7.845 ;
      LAYER met1 ;
        RECT -0.275 7.845 34.625 7.915 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 8.785 1.720 9.265 ;
        RECT 3.855 8.785 4.620 9.265 ;
        RECT 6.755 8.785 7.520 9.265 ;
        RECT 9.655 8.785 10.420 9.265 ;
        RECT 12.555 8.785 13.320 9.265 ;
        RECT 15.455 8.785 16.220 9.265 ;
        RECT 18.355 8.785 19.120 9.265 ;
        RECT 21.255 8.785 22.020 9.265 ;
        RECT 24.155 8.785 24.920 9.265 ;
        RECT 27.055 8.785 27.820 9.265 ;
        RECT 29.955 8.785 30.720 9.265 ;
        RECT 32.855 8.785 33.620 9.265 ;
      LAYER li1 ;
        RECT 1.265 9.195 1.425 9.265 ;
        RECT 4.165 9.195 4.325 9.265 ;
        RECT 7.065 9.195 7.225 9.265 ;
        RECT 9.965 9.195 10.125 9.265 ;
        RECT 12.865 9.195 13.025 9.265 ;
        RECT 15.765 9.195 15.925 9.265 ;
        RECT 18.665 9.195 18.825 9.265 ;
        RECT 21.565 9.195 21.725 9.265 ;
        RECT 24.465 9.195 24.625 9.265 ;
        RECT 27.365 9.195 27.525 9.265 ;
        RECT 30.265 9.195 30.425 9.265 ;
        RECT 33.165 9.195 33.325 9.265 ;
        RECT 1.275 9.185 1.415 9.195 ;
        RECT 4.175 9.185 4.315 9.195 ;
        RECT 7.075 9.185 7.215 9.195 ;
        RECT 9.975 9.185 10.115 9.195 ;
        RECT 12.875 9.185 13.015 9.195 ;
        RECT 15.775 9.185 15.915 9.195 ;
        RECT 18.675 9.185 18.815 9.195 ;
        RECT 21.575 9.185 21.715 9.195 ;
        RECT 24.475 9.185 24.615 9.195 ;
        RECT 27.375 9.185 27.515 9.195 ;
        RECT 30.275 9.185 30.415 9.195 ;
        RECT 33.175 9.185 33.315 9.195 ;
      LAYER met1 ;
        RECT -0.275 9.195 34.625 9.265 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 10.135 1.720 10.615 ;
        RECT 3.855 10.135 4.620 10.615 ;
        RECT 6.755 10.135 7.520 10.615 ;
        RECT 9.655 10.135 10.420 10.615 ;
        RECT 12.555 10.135 13.320 10.615 ;
        RECT 15.455 10.135 16.220 10.615 ;
        RECT 18.355 10.135 19.120 10.615 ;
        RECT 21.255 10.135 22.020 10.615 ;
        RECT 24.155 10.135 24.920 10.615 ;
        RECT 27.055 10.135 27.820 10.615 ;
        RECT 29.955 10.135 30.720 10.615 ;
        RECT 32.855 10.135 33.620 10.615 ;
      LAYER li1 ;
        RECT 1.265 10.545 1.425 10.615 ;
        RECT 4.165 10.545 4.325 10.615 ;
        RECT 7.065 10.545 7.225 10.615 ;
        RECT 9.965 10.545 10.125 10.615 ;
        RECT 12.865 10.545 13.025 10.615 ;
        RECT 15.765 10.545 15.925 10.615 ;
        RECT 18.665 10.545 18.825 10.615 ;
        RECT 21.565 10.545 21.725 10.615 ;
        RECT 24.465 10.545 24.625 10.615 ;
        RECT 27.365 10.545 27.525 10.615 ;
        RECT 30.265 10.545 30.425 10.615 ;
        RECT 33.165 10.545 33.325 10.615 ;
        RECT 1.275 10.535 1.415 10.545 ;
        RECT 4.175 10.535 4.315 10.545 ;
        RECT 7.075 10.535 7.215 10.545 ;
        RECT 9.975 10.535 10.115 10.545 ;
        RECT 12.875 10.535 13.015 10.545 ;
        RECT 15.775 10.535 15.915 10.545 ;
        RECT 18.675 10.535 18.815 10.545 ;
        RECT 21.575 10.535 21.715 10.545 ;
        RECT 24.475 10.535 24.615 10.545 ;
        RECT 27.375 10.535 27.515 10.545 ;
        RECT 30.275 10.535 30.415 10.545 ;
        RECT 33.175 10.535 33.315 10.545 ;
      LAYER met1 ;
        RECT -0.275 10.545 34.625 10.615 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 11.485 1.720 11.965 ;
        RECT 3.855 11.485 4.620 11.965 ;
        RECT 6.755 11.485 7.520 11.965 ;
        RECT 9.655 11.485 10.420 11.965 ;
        RECT 12.555 11.485 13.320 11.965 ;
        RECT 15.455 11.485 16.220 11.965 ;
        RECT 18.355 11.485 19.120 11.965 ;
        RECT 21.255 11.485 22.020 11.965 ;
        RECT 24.155 11.485 24.920 11.965 ;
        RECT 27.055 11.485 27.820 11.965 ;
        RECT 29.955 11.485 30.720 11.965 ;
        RECT 32.855 11.485 33.620 11.965 ;
      LAYER li1 ;
        RECT 1.265 11.895 1.425 11.965 ;
        RECT 4.165 11.895 4.325 11.965 ;
        RECT 7.065 11.895 7.225 11.965 ;
        RECT 9.965 11.895 10.125 11.965 ;
        RECT 12.865 11.895 13.025 11.965 ;
        RECT 15.765 11.895 15.925 11.965 ;
        RECT 18.665 11.895 18.825 11.965 ;
        RECT 21.565 11.895 21.725 11.965 ;
        RECT 24.465 11.895 24.625 11.965 ;
        RECT 27.365 11.895 27.525 11.965 ;
        RECT 30.265 11.895 30.425 11.965 ;
        RECT 33.165 11.895 33.325 11.965 ;
        RECT 1.275 11.885 1.415 11.895 ;
        RECT 4.175 11.885 4.315 11.895 ;
        RECT 7.075 11.885 7.215 11.895 ;
        RECT 9.975 11.885 10.115 11.895 ;
        RECT 12.875 11.885 13.015 11.895 ;
        RECT 15.775 11.885 15.915 11.895 ;
        RECT 18.675 11.885 18.815 11.895 ;
        RECT 21.575 11.885 21.715 11.895 ;
        RECT 24.475 11.885 24.615 11.895 ;
        RECT 27.375 11.885 27.515 11.895 ;
        RECT 30.275 11.885 30.415 11.895 ;
        RECT 33.175 11.885 33.315 11.895 ;
      LAYER met1 ;
        RECT -0.275 11.895 34.625 11.965 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 12.835 1.720 13.315 ;
        RECT 3.855 12.835 4.620 13.315 ;
        RECT 6.755 12.835 7.520 13.315 ;
        RECT 9.655 12.835 10.420 13.315 ;
        RECT 12.555 12.835 13.320 13.315 ;
        RECT 15.455 12.835 16.220 13.315 ;
        RECT 18.355 12.835 19.120 13.315 ;
        RECT 21.255 12.835 22.020 13.315 ;
        RECT 24.155 12.835 24.920 13.315 ;
        RECT 27.055 12.835 27.820 13.315 ;
        RECT 29.955 12.835 30.720 13.315 ;
        RECT 32.855 12.835 33.620 13.315 ;
      LAYER li1 ;
        RECT 1.265 13.245 1.425 13.315 ;
        RECT 4.165 13.245 4.325 13.315 ;
        RECT 7.065 13.245 7.225 13.315 ;
        RECT 9.965 13.245 10.125 13.315 ;
        RECT 12.865 13.245 13.025 13.315 ;
        RECT 15.765 13.245 15.925 13.315 ;
        RECT 18.665 13.245 18.825 13.315 ;
        RECT 21.565 13.245 21.725 13.315 ;
        RECT 24.465 13.245 24.625 13.315 ;
        RECT 27.365 13.245 27.525 13.315 ;
        RECT 30.265 13.245 30.425 13.315 ;
        RECT 33.165 13.245 33.325 13.315 ;
        RECT 1.275 13.235 1.415 13.245 ;
        RECT 4.175 13.235 4.315 13.245 ;
        RECT 7.075 13.235 7.215 13.245 ;
        RECT 9.975 13.235 10.115 13.245 ;
        RECT 12.875 13.235 13.015 13.245 ;
        RECT 15.775 13.235 15.915 13.245 ;
        RECT 18.675 13.235 18.815 13.245 ;
        RECT 21.575 13.235 21.715 13.245 ;
        RECT 24.475 13.235 24.615 13.245 ;
        RECT 27.375 13.235 27.515 13.245 ;
        RECT 30.275 13.235 30.415 13.245 ;
        RECT 33.175 13.235 33.315 13.245 ;
      LAYER met1 ;
        RECT -0.275 13.245 34.625 13.315 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 14.185 1.720 14.665 ;
        RECT 3.855 14.185 4.620 14.665 ;
        RECT 6.755 14.185 7.520 14.665 ;
        RECT 9.655 14.185 10.420 14.665 ;
        RECT 12.555 14.185 13.320 14.665 ;
        RECT 15.455 14.185 16.220 14.665 ;
        RECT 18.355 14.185 19.120 14.665 ;
        RECT 21.255 14.185 22.020 14.665 ;
        RECT 24.155 14.185 24.920 14.665 ;
        RECT 27.055 14.185 27.820 14.665 ;
        RECT 29.955 14.185 30.720 14.665 ;
        RECT 32.855 14.185 33.620 14.665 ;
      LAYER li1 ;
        RECT 1.265 14.595 1.425 14.665 ;
        RECT 4.165 14.595 4.325 14.665 ;
        RECT 7.065 14.595 7.225 14.665 ;
        RECT 9.965 14.595 10.125 14.665 ;
        RECT 12.865 14.595 13.025 14.665 ;
        RECT 15.765 14.595 15.925 14.665 ;
        RECT 18.665 14.595 18.825 14.665 ;
        RECT 21.565 14.595 21.725 14.665 ;
        RECT 24.465 14.595 24.625 14.665 ;
        RECT 27.365 14.595 27.525 14.665 ;
        RECT 30.265 14.595 30.425 14.665 ;
        RECT 33.165 14.595 33.325 14.665 ;
        RECT 1.275 14.585 1.415 14.595 ;
        RECT 4.175 14.585 4.315 14.595 ;
        RECT 7.075 14.585 7.215 14.595 ;
        RECT 9.975 14.585 10.115 14.595 ;
        RECT 12.875 14.585 13.015 14.595 ;
        RECT 15.775 14.585 15.915 14.595 ;
        RECT 18.675 14.585 18.815 14.595 ;
        RECT 21.575 14.585 21.715 14.595 ;
        RECT 24.475 14.585 24.615 14.595 ;
        RECT 27.375 14.585 27.515 14.595 ;
        RECT 30.275 14.585 30.415 14.595 ;
        RECT 33.175 14.585 33.315 14.595 ;
      LAYER met1 ;
        RECT -0.275 14.595 34.625 14.665 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 15.535 1.720 16.015 ;
        RECT 3.855 15.535 4.620 16.015 ;
        RECT 6.755 15.535 7.520 16.015 ;
        RECT 9.655 15.535 10.420 16.015 ;
        RECT 12.555 15.535 13.320 16.015 ;
        RECT 15.455 15.535 16.220 16.015 ;
        RECT 18.355 15.535 19.120 16.015 ;
        RECT 21.255 15.535 22.020 16.015 ;
        RECT 24.155 15.535 24.920 16.015 ;
        RECT 27.055 15.535 27.820 16.015 ;
        RECT 29.955 15.535 30.720 16.015 ;
        RECT 32.855 15.535 33.620 16.015 ;
      LAYER li1 ;
        RECT 1.265 15.945 1.425 16.015 ;
        RECT 4.165 15.945 4.325 16.015 ;
        RECT 7.065 15.945 7.225 16.015 ;
        RECT 9.965 15.945 10.125 16.015 ;
        RECT 12.865 15.945 13.025 16.015 ;
        RECT 15.765 15.945 15.925 16.015 ;
        RECT 18.665 15.945 18.825 16.015 ;
        RECT 21.565 15.945 21.725 16.015 ;
        RECT 24.465 15.945 24.625 16.015 ;
        RECT 27.365 15.945 27.525 16.015 ;
        RECT 30.265 15.945 30.425 16.015 ;
        RECT 33.165 15.945 33.325 16.015 ;
        RECT 1.275 15.935 1.415 15.945 ;
        RECT 4.175 15.935 4.315 15.945 ;
        RECT 7.075 15.935 7.215 15.945 ;
        RECT 9.975 15.935 10.115 15.945 ;
        RECT 12.875 15.935 13.015 15.945 ;
        RECT 15.775 15.935 15.915 15.945 ;
        RECT 18.675 15.935 18.815 15.945 ;
        RECT 21.575 15.935 21.715 15.945 ;
        RECT 24.475 15.935 24.615 15.945 ;
        RECT 27.375 15.935 27.515 15.945 ;
        RECT 30.275 15.935 30.415 15.945 ;
        RECT 33.175 15.935 33.315 15.945 ;
      LAYER met1 ;
        RECT -0.275 15.945 34.625 16.015 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 16.885 1.720 17.365 ;
        RECT 3.855 16.885 4.620 17.365 ;
        RECT 6.755 16.885 7.520 17.365 ;
        RECT 9.655 16.885 10.420 17.365 ;
        RECT 12.555 16.885 13.320 17.365 ;
        RECT 15.455 16.885 16.220 17.365 ;
        RECT 18.355 16.885 19.120 17.365 ;
        RECT 21.255 16.885 22.020 17.365 ;
        RECT 24.155 16.885 24.920 17.365 ;
        RECT 27.055 16.885 27.820 17.365 ;
        RECT 29.955 16.885 30.720 17.365 ;
        RECT 32.855 16.885 33.620 17.365 ;
      LAYER li1 ;
        RECT 1.265 17.295 1.425 17.365 ;
        RECT 4.165 17.295 4.325 17.365 ;
        RECT 7.065 17.295 7.225 17.365 ;
        RECT 9.965 17.295 10.125 17.365 ;
        RECT 12.865 17.295 13.025 17.365 ;
        RECT 15.765 17.295 15.925 17.365 ;
        RECT 18.665 17.295 18.825 17.365 ;
        RECT 21.565 17.295 21.725 17.365 ;
        RECT 24.465 17.295 24.625 17.365 ;
        RECT 27.365 17.295 27.525 17.365 ;
        RECT 30.265 17.295 30.425 17.365 ;
        RECT 33.165 17.295 33.325 17.365 ;
        RECT 1.275 17.285 1.415 17.295 ;
        RECT 4.175 17.285 4.315 17.295 ;
        RECT 7.075 17.285 7.215 17.295 ;
        RECT 9.975 17.285 10.115 17.295 ;
        RECT 12.875 17.285 13.015 17.295 ;
        RECT 15.775 17.285 15.915 17.295 ;
        RECT 18.675 17.285 18.815 17.295 ;
        RECT 21.575 17.285 21.715 17.295 ;
        RECT 24.475 17.285 24.615 17.295 ;
        RECT 27.375 17.285 27.515 17.295 ;
        RECT 30.275 17.285 30.415 17.295 ;
        RECT 33.175 17.285 33.315 17.295 ;
      LAYER met1 ;
        RECT -0.275 17.295 34.625 17.365 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 18.235 1.720 18.715 ;
        RECT 3.855 18.235 4.620 18.715 ;
        RECT 6.755 18.235 7.520 18.715 ;
        RECT 9.655 18.235 10.420 18.715 ;
        RECT 12.555 18.235 13.320 18.715 ;
        RECT 15.455 18.235 16.220 18.715 ;
        RECT 18.355 18.235 19.120 18.715 ;
        RECT 21.255 18.235 22.020 18.715 ;
        RECT 24.155 18.235 24.920 18.715 ;
        RECT 27.055 18.235 27.820 18.715 ;
        RECT 29.955 18.235 30.720 18.715 ;
        RECT 32.855 18.235 33.620 18.715 ;
      LAYER li1 ;
        RECT 1.265 18.645 1.425 18.715 ;
        RECT 4.165 18.645 4.325 18.715 ;
        RECT 7.065 18.645 7.225 18.715 ;
        RECT 9.965 18.645 10.125 18.715 ;
        RECT 12.865 18.645 13.025 18.715 ;
        RECT 15.765 18.645 15.925 18.715 ;
        RECT 18.665 18.645 18.825 18.715 ;
        RECT 21.565 18.645 21.725 18.715 ;
        RECT 24.465 18.645 24.625 18.715 ;
        RECT 27.365 18.645 27.525 18.715 ;
        RECT 30.265 18.645 30.425 18.715 ;
        RECT 33.165 18.645 33.325 18.715 ;
        RECT 1.275 18.635 1.415 18.645 ;
        RECT 4.175 18.635 4.315 18.645 ;
        RECT 7.075 18.635 7.215 18.645 ;
        RECT 9.975 18.635 10.115 18.645 ;
        RECT 12.875 18.635 13.015 18.645 ;
        RECT 15.775 18.635 15.915 18.645 ;
        RECT 18.675 18.635 18.815 18.645 ;
        RECT 21.575 18.635 21.715 18.645 ;
        RECT 24.475 18.635 24.615 18.645 ;
        RECT 27.375 18.635 27.515 18.645 ;
        RECT 30.275 18.635 30.415 18.645 ;
        RECT 33.175 18.635 33.315 18.645 ;
      LAYER met1 ;
        RECT -0.275 18.645 34.625 18.715 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 19.585 1.720 20.065 ;
        RECT 3.855 19.585 4.620 20.065 ;
        RECT 6.755 19.585 7.520 20.065 ;
        RECT 9.655 19.585 10.420 20.065 ;
        RECT 12.555 19.585 13.320 20.065 ;
        RECT 15.455 19.585 16.220 20.065 ;
        RECT 18.355 19.585 19.120 20.065 ;
        RECT 21.255 19.585 22.020 20.065 ;
        RECT 24.155 19.585 24.920 20.065 ;
        RECT 27.055 19.585 27.820 20.065 ;
        RECT 29.955 19.585 30.720 20.065 ;
        RECT 32.855 19.585 33.620 20.065 ;
      LAYER li1 ;
        RECT 1.265 19.995 1.425 20.065 ;
        RECT 4.165 19.995 4.325 20.065 ;
        RECT 7.065 19.995 7.225 20.065 ;
        RECT 9.965 19.995 10.125 20.065 ;
        RECT 12.865 19.995 13.025 20.065 ;
        RECT 15.765 19.995 15.925 20.065 ;
        RECT 18.665 19.995 18.825 20.065 ;
        RECT 21.565 19.995 21.725 20.065 ;
        RECT 24.465 19.995 24.625 20.065 ;
        RECT 27.365 19.995 27.525 20.065 ;
        RECT 30.265 19.995 30.425 20.065 ;
        RECT 33.165 19.995 33.325 20.065 ;
        RECT 1.275 19.985 1.415 19.995 ;
        RECT 4.175 19.985 4.315 19.995 ;
        RECT 7.075 19.985 7.215 19.995 ;
        RECT 9.975 19.985 10.115 19.995 ;
        RECT 12.875 19.985 13.015 19.995 ;
        RECT 15.775 19.985 15.915 19.995 ;
        RECT 18.675 19.985 18.815 19.995 ;
        RECT 21.575 19.985 21.715 19.995 ;
        RECT 24.475 19.985 24.615 19.995 ;
        RECT 27.375 19.985 27.515 19.995 ;
        RECT 30.275 19.985 30.415 19.995 ;
        RECT 33.175 19.985 33.315 19.995 ;
      LAYER met1 ;
        RECT -0.275 19.995 34.625 20.065 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.955 20.935 1.720 21.415 ;
        RECT 3.855 20.935 4.620 21.415 ;
        RECT 6.755 20.935 7.520 21.415 ;
        RECT 9.655 20.935 10.420 21.415 ;
        RECT 12.555 20.935 13.320 21.415 ;
        RECT 15.455 20.935 16.220 21.415 ;
        RECT 18.355 20.935 19.120 21.415 ;
        RECT 21.255 20.935 22.020 21.415 ;
        RECT 24.155 20.935 24.920 21.415 ;
        RECT 27.055 20.935 27.820 21.415 ;
        RECT 29.955 20.935 30.720 21.415 ;
        RECT 32.855 20.935 33.620 21.415 ;
      LAYER li1 ;
        RECT 1.265 21.345 1.425 21.415 ;
        RECT 4.165 21.345 4.325 21.415 ;
        RECT 7.065 21.345 7.225 21.415 ;
        RECT 9.965 21.345 10.125 21.415 ;
        RECT 12.865 21.345 13.025 21.415 ;
        RECT 15.765 21.345 15.925 21.415 ;
        RECT 18.665 21.345 18.825 21.415 ;
        RECT 21.565 21.345 21.725 21.415 ;
        RECT 24.465 21.345 24.625 21.415 ;
        RECT 27.365 21.345 27.525 21.415 ;
        RECT 30.265 21.345 30.425 21.415 ;
        RECT 33.165 21.345 33.325 21.415 ;
        RECT 1.275 21.335 1.415 21.345 ;
        RECT 4.175 21.335 4.315 21.345 ;
        RECT 7.075 21.335 7.215 21.345 ;
        RECT 9.975 21.335 10.115 21.345 ;
        RECT 12.875 21.335 13.015 21.345 ;
        RECT 15.775 21.335 15.915 21.345 ;
        RECT 18.675 21.335 18.815 21.345 ;
        RECT 21.575 21.335 21.715 21.345 ;
        RECT 24.475 21.335 24.615 21.345 ;
        RECT 27.375 21.335 27.515 21.345 ;
        RECT 30.275 21.335 30.415 21.345 ;
        RECT 33.175 21.335 33.315 21.345 ;
      LAYER met1 ;
        RECT -0.275 21.345 34.625 21.415 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.035 20.705 0.815 21.565 ;
        RECT 1.875 20.705 3.715 21.565 ;
        RECT 4.775 20.705 5.625 21.565 ;
        RECT -0.035 20.215 5.625 20.705 ;
        RECT -0.035 19.355 0.815 20.215 ;
        RECT 1.875 19.355 3.715 20.215 ;
        RECT 4.775 19.355 5.625 20.215 ;
        RECT -0.035 18.865 5.625 19.355 ;
        RECT -0.035 18.005 0.815 18.865 ;
        RECT 1.875 18.005 3.715 18.865 ;
        RECT 4.775 18.005 5.625 18.865 ;
        RECT -0.035 17.515 5.625 18.005 ;
        RECT -0.035 16.655 0.815 17.515 ;
        RECT 1.875 16.655 3.715 17.515 ;
        RECT 4.775 16.655 5.625 17.515 ;
        RECT -0.035 16.165 5.625 16.655 ;
        RECT -0.035 15.305 0.815 16.165 ;
        RECT 1.875 15.305 3.715 16.165 ;
        RECT 4.775 15.305 5.625 16.165 ;
        RECT -0.035 14.815 5.625 15.305 ;
        RECT -0.035 13.955 0.815 14.815 ;
        RECT 1.875 13.955 3.715 14.815 ;
        RECT 4.775 13.955 5.625 14.815 ;
        RECT -0.035 13.465 5.625 13.955 ;
        RECT -0.035 12.605 0.815 13.465 ;
        RECT 1.875 12.605 3.715 13.465 ;
        RECT 4.775 12.605 5.625 13.465 ;
        RECT -0.035 12.115 5.625 12.605 ;
        RECT -0.035 11.255 0.815 12.115 ;
        RECT 1.875 11.255 3.715 12.115 ;
        RECT 4.775 11.255 5.625 12.115 ;
        RECT -0.035 10.765 5.625 11.255 ;
        RECT -0.035 9.905 0.815 10.765 ;
        RECT 1.875 9.905 3.715 10.765 ;
        RECT 4.775 9.905 5.625 10.765 ;
        RECT -0.035 9.415 5.625 9.905 ;
        RECT -0.035 8.555 0.815 9.415 ;
        RECT 1.875 8.555 3.715 9.415 ;
        RECT 4.775 8.555 5.625 9.415 ;
        RECT -0.035 8.065 5.625 8.555 ;
        RECT -0.035 7.205 0.815 8.065 ;
        RECT 1.875 7.205 3.715 8.065 ;
        RECT 4.775 7.205 5.625 8.065 ;
        RECT -0.035 6.715 5.625 7.205 ;
        RECT -0.035 5.855 0.815 6.715 ;
        RECT 1.875 5.855 3.715 6.715 ;
        RECT 4.775 5.855 5.625 6.715 ;
        RECT -0.035 5.365 5.625 5.855 ;
        RECT -0.035 4.505 0.815 5.365 ;
        RECT 1.875 4.505 3.715 5.365 ;
        RECT 4.775 4.505 5.625 5.365 ;
        RECT -0.035 4.015 5.625 4.505 ;
        RECT -0.035 3.155 0.815 4.015 ;
        RECT 1.875 3.155 3.715 4.015 ;
        RECT 4.775 3.155 5.625 4.015 ;
        RECT -0.035 2.665 5.625 3.155 ;
        RECT -0.035 1.805 0.815 2.665 ;
        RECT 1.875 1.805 3.715 2.665 ;
        RECT 4.775 1.805 5.625 2.665 ;
        RECT -0.035 1.315 5.625 1.805 ;
        RECT -0.035 0.455 0.815 1.315 ;
        RECT 1.875 0.455 3.715 1.315 ;
        RECT 4.775 0.455 5.625 1.315 ;
        RECT -0.035 -0.035 5.625 0.455 ;
        RECT 5.765 20.705 6.615 21.565 ;
        RECT 7.675 20.705 9.515 21.565 ;
        RECT 10.575 20.705 11.425 21.565 ;
        RECT 5.765 20.215 11.425 20.705 ;
        RECT 5.765 19.355 6.615 20.215 ;
        RECT 7.675 19.355 9.515 20.215 ;
        RECT 10.575 19.355 11.425 20.215 ;
        RECT 5.765 18.865 11.425 19.355 ;
        RECT 5.765 18.005 6.615 18.865 ;
        RECT 7.675 18.005 9.515 18.865 ;
        RECT 10.575 18.005 11.425 18.865 ;
        RECT 5.765 17.515 11.425 18.005 ;
        RECT 5.765 16.655 6.615 17.515 ;
        RECT 7.675 16.655 9.515 17.515 ;
        RECT 10.575 16.655 11.425 17.515 ;
        RECT 5.765 16.165 11.425 16.655 ;
        RECT 5.765 15.305 6.615 16.165 ;
        RECT 7.675 15.305 9.515 16.165 ;
        RECT 10.575 15.305 11.425 16.165 ;
        RECT 5.765 14.815 11.425 15.305 ;
        RECT 5.765 13.955 6.615 14.815 ;
        RECT 7.675 13.955 9.515 14.815 ;
        RECT 10.575 13.955 11.425 14.815 ;
        RECT 5.765 13.465 11.425 13.955 ;
        RECT 5.765 12.605 6.615 13.465 ;
        RECT 7.675 12.605 9.515 13.465 ;
        RECT 10.575 12.605 11.425 13.465 ;
        RECT 5.765 12.115 11.425 12.605 ;
        RECT 5.765 11.255 6.615 12.115 ;
        RECT 7.675 11.255 9.515 12.115 ;
        RECT 10.575 11.255 11.425 12.115 ;
        RECT 5.765 10.765 11.425 11.255 ;
        RECT 5.765 9.905 6.615 10.765 ;
        RECT 7.675 9.905 9.515 10.765 ;
        RECT 10.575 9.905 11.425 10.765 ;
        RECT 5.765 9.415 11.425 9.905 ;
        RECT 5.765 8.555 6.615 9.415 ;
        RECT 7.675 8.555 9.515 9.415 ;
        RECT 10.575 8.555 11.425 9.415 ;
        RECT 5.765 8.065 11.425 8.555 ;
        RECT 5.765 7.205 6.615 8.065 ;
        RECT 7.675 7.205 9.515 8.065 ;
        RECT 10.575 7.205 11.425 8.065 ;
        RECT 5.765 6.715 11.425 7.205 ;
        RECT 5.765 5.855 6.615 6.715 ;
        RECT 7.675 5.855 9.515 6.715 ;
        RECT 10.575 5.855 11.425 6.715 ;
        RECT 5.765 5.365 11.425 5.855 ;
        RECT 5.765 4.505 6.615 5.365 ;
        RECT 7.675 4.505 9.515 5.365 ;
        RECT 10.575 4.505 11.425 5.365 ;
        RECT 5.765 4.015 11.425 4.505 ;
        RECT 5.765 3.155 6.615 4.015 ;
        RECT 7.675 3.155 9.515 4.015 ;
        RECT 10.575 3.155 11.425 4.015 ;
        RECT 5.765 2.665 11.425 3.155 ;
        RECT 5.765 1.805 6.615 2.665 ;
        RECT 7.675 1.805 9.515 2.665 ;
        RECT 10.575 1.805 11.425 2.665 ;
        RECT 5.765 1.315 11.425 1.805 ;
        RECT 5.765 0.455 6.615 1.315 ;
        RECT 7.675 0.455 9.515 1.315 ;
        RECT 10.575 0.455 11.425 1.315 ;
        RECT 5.765 -0.035 11.425 0.455 ;
        RECT 11.565 20.705 12.415 21.565 ;
        RECT 13.475 20.705 15.315 21.565 ;
        RECT 16.375 20.705 17.225 21.565 ;
        RECT 11.565 20.215 17.225 20.705 ;
        RECT 11.565 19.355 12.415 20.215 ;
        RECT 13.475 19.355 15.315 20.215 ;
        RECT 16.375 19.355 17.225 20.215 ;
        RECT 11.565 18.865 17.225 19.355 ;
        RECT 11.565 18.005 12.415 18.865 ;
        RECT 13.475 18.005 15.315 18.865 ;
        RECT 16.375 18.005 17.225 18.865 ;
        RECT 11.565 17.515 17.225 18.005 ;
        RECT 11.565 16.655 12.415 17.515 ;
        RECT 13.475 16.655 15.315 17.515 ;
        RECT 16.375 16.655 17.225 17.515 ;
        RECT 11.565 16.165 17.225 16.655 ;
        RECT 11.565 15.305 12.415 16.165 ;
        RECT 13.475 15.305 15.315 16.165 ;
        RECT 16.375 15.305 17.225 16.165 ;
        RECT 11.565 14.815 17.225 15.305 ;
        RECT 11.565 13.955 12.415 14.815 ;
        RECT 13.475 13.955 15.315 14.815 ;
        RECT 16.375 13.955 17.225 14.815 ;
        RECT 11.565 13.465 17.225 13.955 ;
        RECT 11.565 12.605 12.415 13.465 ;
        RECT 13.475 12.605 15.315 13.465 ;
        RECT 16.375 12.605 17.225 13.465 ;
        RECT 11.565 12.115 17.225 12.605 ;
        RECT 11.565 11.255 12.415 12.115 ;
        RECT 13.475 11.255 15.315 12.115 ;
        RECT 16.375 11.255 17.225 12.115 ;
        RECT 11.565 10.765 17.225 11.255 ;
        RECT 11.565 9.905 12.415 10.765 ;
        RECT 13.475 9.905 15.315 10.765 ;
        RECT 16.375 9.905 17.225 10.765 ;
        RECT 11.565 9.415 17.225 9.905 ;
        RECT 11.565 8.555 12.415 9.415 ;
        RECT 13.475 8.555 15.315 9.415 ;
        RECT 16.375 8.555 17.225 9.415 ;
        RECT 11.565 8.065 17.225 8.555 ;
        RECT 11.565 7.205 12.415 8.065 ;
        RECT 13.475 7.205 15.315 8.065 ;
        RECT 16.375 7.205 17.225 8.065 ;
        RECT 11.565 6.715 17.225 7.205 ;
        RECT 11.565 5.855 12.415 6.715 ;
        RECT 13.475 5.855 15.315 6.715 ;
        RECT 16.375 5.855 17.225 6.715 ;
        RECT 11.565 5.365 17.225 5.855 ;
        RECT 11.565 4.505 12.415 5.365 ;
        RECT 13.475 4.505 15.315 5.365 ;
        RECT 16.375 4.505 17.225 5.365 ;
        RECT 11.565 4.015 17.225 4.505 ;
        RECT 11.565 3.155 12.415 4.015 ;
        RECT 13.475 3.155 15.315 4.015 ;
        RECT 16.375 3.155 17.225 4.015 ;
        RECT 11.565 2.665 17.225 3.155 ;
        RECT 11.565 1.805 12.415 2.665 ;
        RECT 13.475 1.805 15.315 2.665 ;
        RECT 16.375 1.805 17.225 2.665 ;
        RECT 11.565 1.315 17.225 1.805 ;
        RECT 11.565 0.455 12.415 1.315 ;
        RECT 13.475 0.455 15.315 1.315 ;
        RECT 16.375 0.455 17.225 1.315 ;
        RECT 11.565 -0.035 17.225 0.455 ;
        RECT 17.365 20.705 18.215 21.565 ;
        RECT 19.275 20.705 21.115 21.565 ;
        RECT 22.175 20.705 23.025 21.565 ;
        RECT 17.365 20.215 23.025 20.705 ;
        RECT 17.365 19.355 18.215 20.215 ;
        RECT 19.275 19.355 21.115 20.215 ;
        RECT 22.175 19.355 23.025 20.215 ;
        RECT 17.365 18.865 23.025 19.355 ;
        RECT 17.365 18.005 18.215 18.865 ;
        RECT 19.275 18.005 21.115 18.865 ;
        RECT 22.175 18.005 23.025 18.865 ;
        RECT 17.365 17.515 23.025 18.005 ;
        RECT 17.365 16.655 18.215 17.515 ;
        RECT 19.275 16.655 21.115 17.515 ;
        RECT 22.175 16.655 23.025 17.515 ;
        RECT 17.365 16.165 23.025 16.655 ;
        RECT 17.365 15.305 18.215 16.165 ;
        RECT 19.275 15.305 21.115 16.165 ;
        RECT 22.175 15.305 23.025 16.165 ;
        RECT 17.365 14.815 23.025 15.305 ;
        RECT 17.365 13.955 18.215 14.815 ;
        RECT 19.275 13.955 21.115 14.815 ;
        RECT 22.175 13.955 23.025 14.815 ;
        RECT 17.365 13.465 23.025 13.955 ;
        RECT 17.365 12.605 18.215 13.465 ;
        RECT 19.275 12.605 21.115 13.465 ;
        RECT 22.175 12.605 23.025 13.465 ;
        RECT 17.365 12.115 23.025 12.605 ;
        RECT 17.365 11.255 18.215 12.115 ;
        RECT 19.275 11.255 21.115 12.115 ;
        RECT 22.175 11.255 23.025 12.115 ;
        RECT 17.365 10.765 23.025 11.255 ;
        RECT 17.365 9.905 18.215 10.765 ;
        RECT 19.275 9.905 21.115 10.765 ;
        RECT 22.175 9.905 23.025 10.765 ;
        RECT 17.365 9.415 23.025 9.905 ;
        RECT 17.365 8.555 18.215 9.415 ;
        RECT 19.275 8.555 21.115 9.415 ;
        RECT 22.175 8.555 23.025 9.415 ;
        RECT 17.365 8.065 23.025 8.555 ;
        RECT 17.365 7.205 18.215 8.065 ;
        RECT 19.275 7.205 21.115 8.065 ;
        RECT 22.175 7.205 23.025 8.065 ;
        RECT 17.365 6.715 23.025 7.205 ;
        RECT 17.365 5.855 18.215 6.715 ;
        RECT 19.275 5.855 21.115 6.715 ;
        RECT 22.175 5.855 23.025 6.715 ;
        RECT 17.365 5.365 23.025 5.855 ;
        RECT 17.365 4.505 18.215 5.365 ;
        RECT 19.275 4.505 21.115 5.365 ;
        RECT 22.175 4.505 23.025 5.365 ;
        RECT 17.365 4.015 23.025 4.505 ;
        RECT 17.365 3.155 18.215 4.015 ;
        RECT 19.275 3.155 21.115 4.015 ;
        RECT 22.175 3.155 23.025 4.015 ;
        RECT 17.365 2.665 23.025 3.155 ;
        RECT 17.365 1.805 18.215 2.665 ;
        RECT 19.275 1.805 21.115 2.665 ;
        RECT 22.175 1.805 23.025 2.665 ;
        RECT 17.365 1.315 23.025 1.805 ;
        RECT 17.365 0.455 18.215 1.315 ;
        RECT 19.275 0.455 21.115 1.315 ;
        RECT 22.175 0.455 23.025 1.315 ;
        RECT 17.365 -0.035 23.025 0.455 ;
        RECT 23.165 20.705 24.015 21.565 ;
        RECT 25.075 20.705 26.915 21.565 ;
        RECT 27.975 20.705 28.825 21.565 ;
        RECT 23.165 20.215 28.825 20.705 ;
        RECT 23.165 19.355 24.015 20.215 ;
        RECT 25.075 19.355 26.915 20.215 ;
        RECT 27.975 19.355 28.825 20.215 ;
        RECT 23.165 18.865 28.825 19.355 ;
        RECT 23.165 18.005 24.015 18.865 ;
        RECT 25.075 18.005 26.915 18.865 ;
        RECT 27.975 18.005 28.825 18.865 ;
        RECT 23.165 17.515 28.825 18.005 ;
        RECT 23.165 16.655 24.015 17.515 ;
        RECT 25.075 16.655 26.915 17.515 ;
        RECT 27.975 16.655 28.825 17.515 ;
        RECT 23.165 16.165 28.825 16.655 ;
        RECT 23.165 15.305 24.015 16.165 ;
        RECT 25.075 15.305 26.915 16.165 ;
        RECT 27.975 15.305 28.825 16.165 ;
        RECT 23.165 14.815 28.825 15.305 ;
        RECT 23.165 13.955 24.015 14.815 ;
        RECT 25.075 13.955 26.915 14.815 ;
        RECT 27.975 13.955 28.825 14.815 ;
        RECT 23.165 13.465 28.825 13.955 ;
        RECT 23.165 12.605 24.015 13.465 ;
        RECT 25.075 12.605 26.915 13.465 ;
        RECT 27.975 12.605 28.825 13.465 ;
        RECT 23.165 12.115 28.825 12.605 ;
        RECT 23.165 11.255 24.015 12.115 ;
        RECT 25.075 11.255 26.915 12.115 ;
        RECT 27.975 11.255 28.825 12.115 ;
        RECT 23.165 10.765 28.825 11.255 ;
        RECT 23.165 9.905 24.015 10.765 ;
        RECT 25.075 9.905 26.915 10.765 ;
        RECT 27.975 9.905 28.825 10.765 ;
        RECT 23.165 9.415 28.825 9.905 ;
        RECT 23.165 8.555 24.015 9.415 ;
        RECT 25.075 8.555 26.915 9.415 ;
        RECT 27.975 8.555 28.825 9.415 ;
        RECT 23.165 8.065 28.825 8.555 ;
        RECT 23.165 7.205 24.015 8.065 ;
        RECT 25.075 7.205 26.915 8.065 ;
        RECT 27.975 7.205 28.825 8.065 ;
        RECT 23.165 6.715 28.825 7.205 ;
        RECT 23.165 5.855 24.015 6.715 ;
        RECT 25.075 5.855 26.915 6.715 ;
        RECT 27.975 5.855 28.825 6.715 ;
        RECT 23.165 5.365 28.825 5.855 ;
        RECT 23.165 4.505 24.015 5.365 ;
        RECT 25.075 4.505 26.915 5.365 ;
        RECT 27.975 4.505 28.825 5.365 ;
        RECT 23.165 4.015 28.825 4.505 ;
        RECT 23.165 3.155 24.015 4.015 ;
        RECT 25.075 3.155 26.915 4.015 ;
        RECT 27.975 3.155 28.825 4.015 ;
        RECT 23.165 2.665 28.825 3.155 ;
        RECT 23.165 1.805 24.015 2.665 ;
        RECT 25.075 1.805 26.915 2.665 ;
        RECT 27.975 1.805 28.825 2.665 ;
        RECT 23.165 1.315 28.825 1.805 ;
        RECT 23.165 0.455 24.015 1.315 ;
        RECT 25.075 0.455 26.915 1.315 ;
        RECT 27.975 0.455 28.825 1.315 ;
        RECT 23.165 -0.035 28.825 0.455 ;
        RECT 28.965 20.705 29.815 21.565 ;
        RECT 30.875 20.705 32.715 21.565 ;
        RECT 33.775 20.705 34.625 21.565 ;
        RECT 28.965 20.215 34.625 20.705 ;
        RECT 28.965 19.355 29.815 20.215 ;
        RECT 30.875 19.355 32.715 20.215 ;
        RECT 33.775 19.355 34.625 20.215 ;
        RECT 28.965 18.865 34.625 19.355 ;
        RECT 28.965 18.005 29.815 18.865 ;
        RECT 30.875 18.005 32.715 18.865 ;
        RECT 33.775 18.005 34.625 18.865 ;
        RECT 28.965 17.515 34.625 18.005 ;
        RECT 28.965 16.655 29.815 17.515 ;
        RECT 30.875 16.655 32.715 17.515 ;
        RECT 33.775 16.655 34.625 17.515 ;
        RECT 28.965 16.165 34.625 16.655 ;
        RECT 28.965 15.305 29.815 16.165 ;
        RECT 30.875 15.305 32.715 16.165 ;
        RECT 33.775 15.305 34.625 16.165 ;
        RECT 28.965 14.815 34.625 15.305 ;
        RECT 28.965 13.955 29.815 14.815 ;
        RECT 30.875 13.955 32.715 14.815 ;
        RECT 33.775 13.955 34.625 14.815 ;
        RECT 28.965 13.465 34.625 13.955 ;
        RECT 28.965 12.605 29.815 13.465 ;
        RECT 30.875 12.605 32.715 13.465 ;
        RECT 33.775 12.605 34.625 13.465 ;
        RECT 28.965 12.115 34.625 12.605 ;
        RECT 28.965 11.255 29.815 12.115 ;
        RECT 30.875 11.255 32.715 12.115 ;
        RECT 33.775 11.255 34.625 12.115 ;
        RECT 28.965 10.765 34.625 11.255 ;
        RECT 28.965 9.905 29.815 10.765 ;
        RECT 30.875 9.905 32.715 10.765 ;
        RECT 33.775 9.905 34.625 10.765 ;
        RECT 28.965 9.415 34.625 9.905 ;
        RECT 28.965 8.555 29.815 9.415 ;
        RECT 30.875 8.555 32.715 9.415 ;
        RECT 33.775 8.555 34.625 9.415 ;
        RECT 28.965 8.065 34.625 8.555 ;
        RECT 28.965 7.205 29.815 8.065 ;
        RECT 30.875 7.205 32.715 8.065 ;
        RECT 33.775 7.205 34.625 8.065 ;
        RECT 28.965 6.715 34.625 7.205 ;
        RECT 28.965 5.855 29.815 6.715 ;
        RECT 30.875 5.855 32.715 6.715 ;
        RECT 33.775 5.855 34.625 6.715 ;
        RECT 28.965 5.365 34.625 5.855 ;
        RECT 28.965 4.505 29.815 5.365 ;
        RECT 30.875 4.505 32.715 5.365 ;
        RECT 33.775 4.505 34.625 5.365 ;
        RECT 28.965 4.015 34.625 4.505 ;
        RECT 28.965 3.155 29.815 4.015 ;
        RECT 30.875 3.155 32.715 4.015 ;
        RECT 33.775 3.155 34.625 4.015 ;
        RECT 28.965 2.665 34.625 3.155 ;
        RECT 28.965 1.805 29.815 2.665 ;
        RECT 30.875 1.805 32.715 2.665 ;
        RECT 33.775 1.805 34.625 2.665 ;
        RECT 28.965 1.315 34.625 1.805 ;
        RECT 28.965 0.455 29.815 1.315 ;
        RECT 30.875 0.455 32.715 1.315 ;
        RECT 33.775 0.455 34.625 1.315 ;
        RECT 28.965 -0.035 34.625 0.455 ;
      LAYER li1 ;
        RECT 1.275 20.285 1.415 20.295 ;
        RECT 4.175 20.285 4.315 20.295 ;
        RECT 7.075 20.285 7.215 20.295 ;
        RECT 9.975 20.285 10.115 20.295 ;
        RECT 12.875 20.285 13.015 20.295 ;
        RECT 15.775 20.285 15.915 20.295 ;
        RECT 18.675 20.285 18.815 20.295 ;
        RECT 21.575 20.285 21.715 20.295 ;
        RECT 24.475 20.285 24.615 20.295 ;
        RECT 27.375 20.285 27.515 20.295 ;
        RECT 30.275 20.285 30.415 20.295 ;
        RECT 33.175 20.285 33.315 20.295 ;
        RECT 1.265 20.215 1.425 20.285 ;
        RECT 4.165 20.215 4.325 20.285 ;
        RECT 7.065 20.215 7.225 20.285 ;
        RECT 9.965 20.215 10.125 20.285 ;
        RECT 12.865 20.215 13.025 20.285 ;
        RECT 15.765 20.215 15.925 20.285 ;
        RECT 18.665 20.215 18.825 20.285 ;
        RECT 21.565 20.215 21.725 20.285 ;
        RECT 24.465 20.215 24.625 20.285 ;
        RECT 27.365 20.215 27.525 20.285 ;
        RECT 30.265 20.215 30.425 20.285 ;
        RECT 33.165 20.215 33.325 20.285 ;
        RECT 1.275 18.935 1.415 18.945 ;
        RECT 4.175 18.935 4.315 18.945 ;
        RECT 7.075 18.935 7.215 18.945 ;
        RECT 9.975 18.935 10.115 18.945 ;
        RECT 12.875 18.935 13.015 18.945 ;
        RECT 15.775 18.935 15.915 18.945 ;
        RECT 18.675 18.935 18.815 18.945 ;
        RECT 21.575 18.935 21.715 18.945 ;
        RECT 24.475 18.935 24.615 18.945 ;
        RECT 27.375 18.935 27.515 18.945 ;
        RECT 30.275 18.935 30.415 18.945 ;
        RECT 33.175 18.935 33.315 18.945 ;
        RECT 1.265 18.865 1.425 18.935 ;
        RECT 4.165 18.865 4.325 18.935 ;
        RECT 7.065 18.865 7.225 18.935 ;
        RECT 9.965 18.865 10.125 18.935 ;
        RECT 12.865 18.865 13.025 18.935 ;
        RECT 15.765 18.865 15.925 18.935 ;
        RECT 18.665 18.865 18.825 18.935 ;
        RECT 21.565 18.865 21.725 18.935 ;
        RECT 24.465 18.865 24.625 18.935 ;
        RECT 27.365 18.865 27.525 18.935 ;
        RECT 30.265 18.865 30.425 18.935 ;
        RECT 33.165 18.865 33.325 18.935 ;
        RECT 1.275 17.585 1.415 17.595 ;
        RECT 4.175 17.585 4.315 17.595 ;
        RECT 7.075 17.585 7.215 17.595 ;
        RECT 9.975 17.585 10.115 17.595 ;
        RECT 12.875 17.585 13.015 17.595 ;
        RECT 15.775 17.585 15.915 17.595 ;
        RECT 18.675 17.585 18.815 17.595 ;
        RECT 21.575 17.585 21.715 17.595 ;
        RECT 24.475 17.585 24.615 17.595 ;
        RECT 27.375 17.585 27.515 17.595 ;
        RECT 30.275 17.585 30.415 17.595 ;
        RECT 33.175 17.585 33.315 17.595 ;
        RECT 1.265 17.515 1.425 17.585 ;
        RECT 4.165 17.515 4.325 17.585 ;
        RECT 7.065 17.515 7.225 17.585 ;
        RECT 9.965 17.515 10.125 17.585 ;
        RECT 12.865 17.515 13.025 17.585 ;
        RECT 15.765 17.515 15.925 17.585 ;
        RECT 18.665 17.515 18.825 17.585 ;
        RECT 21.565 17.515 21.725 17.585 ;
        RECT 24.465 17.515 24.625 17.585 ;
        RECT 27.365 17.515 27.525 17.585 ;
        RECT 30.265 17.515 30.425 17.585 ;
        RECT 33.165 17.515 33.325 17.585 ;
        RECT 1.275 16.235 1.415 16.245 ;
        RECT 4.175 16.235 4.315 16.245 ;
        RECT 7.075 16.235 7.215 16.245 ;
        RECT 9.975 16.235 10.115 16.245 ;
        RECT 12.875 16.235 13.015 16.245 ;
        RECT 15.775 16.235 15.915 16.245 ;
        RECT 18.675 16.235 18.815 16.245 ;
        RECT 21.575 16.235 21.715 16.245 ;
        RECT 24.475 16.235 24.615 16.245 ;
        RECT 27.375 16.235 27.515 16.245 ;
        RECT 30.275 16.235 30.415 16.245 ;
        RECT 33.175 16.235 33.315 16.245 ;
        RECT 1.265 16.165 1.425 16.235 ;
        RECT 4.165 16.165 4.325 16.235 ;
        RECT 7.065 16.165 7.225 16.235 ;
        RECT 9.965 16.165 10.125 16.235 ;
        RECT 12.865 16.165 13.025 16.235 ;
        RECT 15.765 16.165 15.925 16.235 ;
        RECT 18.665 16.165 18.825 16.235 ;
        RECT 21.565 16.165 21.725 16.235 ;
        RECT 24.465 16.165 24.625 16.235 ;
        RECT 27.365 16.165 27.525 16.235 ;
        RECT 30.265 16.165 30.425 16.235 ;
        RECT 33.165 16.165 33.325 16.235 ;
        RECT 1.275 14.885 1.415 14.895 ;
        RECT 4.175 14.885 4.315 14.895 ;
        RECT 7.075 14.885 7.215 14.895 ;
        RECT 9.975 14.885 10.115 14.895 ;
        RECT 12.875 14.885 13.015 14.895 ;
        RECT 15.775 14.885 15.915 14.895 ;
        RECT 18.675 14.885 18.815 14.895 ;
        RECT 21.575 14.885 21.715 14.895 ;
        RECT 24.475 14.885 24.615 14.895 ;
        RECT 27.375 14.885 27.515 14.895 ;
        RECT 30.275 14.885 30.415 14.895 ;
        RECT 33.175 14.885 33.315 14.895 ;
        RECT 1.265 14.815 1.425 14.885 ;
        RECT 4.165 14.815 4.325 14.885 ;
        RECT 7.065 14.815 7.225 14.885 ;
        RECT 9.965 14.815 10.125 14.885 ;
        RECT 12.865 14.815 13.025 14.885 ;
        RECT 15.765 14.815 15.925 14.885 ;
        RECT 18.665 14.815 18.825 14.885 ;
        RECT 21.565 14.815 21.725 14.885 ;
        RECT 24.465 14.815 24.625 14.885 ;
        RECT 27.365 14.815 27.525 14.885 ;
        RECT 30.265 14.815 30.425 14.885 ;
        RECT 33.165 14.815 33.325 14.885 ;
        RECT 1.275 13.535 1.415 13.545 ;
        RECT 4.175 13.535 4.315 13.545 ;
        RECT 7.075 13.535 7.215 13.545 ;
        RECT 9.975 13.535 10.115 13.545 ;
        RECT 12.875 13.535 13.015 13.545 ;
        RECT 15.775 13.535 15.915 13.545 ;
        RECT 18.675 13.535 18.815 13.545 ;
        RECT 21.575 13.535 21.715 13.545 ;
        RECT 24.475 13.535 24.615 13.545 ;
        RECT 27.375 13.535 27.515 13.545 ;
        RECT 30.275 13.535 30.415 13.545 ;
        RECT 33.175 13.535 33.315 13.545 ;
        RECT 1.265 13.465 1.425 13.535 ;
        RECT 4.165 13.465 4.325 13.535 ;
        RECT 7.065 13.465 7.225 13.535 ;
        RECT 9.965 13.465 10.125 13.535 ;
        RECT 12.865 13.465 13.025 13.535 ;
        RECT 15.765 13.465 15.925 13.535 ;
        RECT 18.665 13.465 18.825 13.535 ;
        RECT 21.565 13.465 21.725 13.535 ;
        RECT 24.465 13.465 24.625 13.535 ;
        RECT 27.365 13.465 27.525 13.535 ;
        RECT 30.265 13.465 30.425 13.535 ;
        RECT 33.165 13.465 33.325 13.535 ;
        RECT 1.275 12.185 1.415 12.195 ;
        RECT 4.175 12.185 4.315 12.195 ;
        RECT 7.075 12.185 7.215 12.195 ;
        RECT 9.975 12.185 10.115 12.195 ;
        RECT 12.875 12.185 13.015 12.195 ;
        RECT 15.775 12.185 15.915 12.195 ;
        RECT 18.675 12.185 18.815 12.195 ;
        RECT 21.575 12.185 21.715 12.195 ;
        RECT 24.475 12.185 24.615 12.195 ;
        RECT 27.375 12.185 27.515 12.195 ;
        RECT 30.275 12.185 30.415 12.195 ;
        RECT 33.175 12.185 33.315 12.195 ;
        RECT 1.265 12.115 1.425 12.185 ;
        RECT 4.165 12.115 4.325 12.185 ;
        RECT 7.065 12.115 7.225 12.185 ;
        RECT 9.965 12.115 10.125 12.185 ;
        RECT 12.865 12.115 13.025 12.185 ;
        RECT 15.765 12.115 15.925 12.185 ;
        RECT 18.665 12.115 18.825 12.185 ;
        RECT 21.565 12.115 21.725 12.185 ;
        RECT 24.465 12.115 24.625 12.185 ;
        RECT 27.365 12.115 27.525 12.185 ;
        RECT 30.265 12.115 30.425 12.185 ;
        RECT 33.165 12.115 33.325 12.185 ;
        RECT 1.275 10.835 1.415 10.845 ;
        RECT 4.175 10.835 4.315 10.845 ;
        RECT 7.075 10.835 7.215 10.845 ;
        RECT 9.975 10.835 10.115 10.845 ;
        RECT 12.875 10.835 13.015 10.845 ;
        RECT 15.775 10.835 15.915 10.845 ;
        RECT 18.675 10.835 18.815 10.845 ;
        RECT 21.575 10.835 21.715 10.845 ;
        RECT 24.475 10.835 24.615 10.845 ;
        RECT 27.375 10.835 27.515 10.845 ;
        RECT 30.275 10.835 30.415 10.845 ;
        RECT 33.175 10.835 33.315 10.845 ;
        RECT 1.265 10.765 1.425 10.835 ;
        RECT 4.165 10.765 4.325 10.835 ;
        RECT 7.065 10.765 7.225 10.835 ;
        RECT 9.965 10.765 10.125 10.835 ;
        RECT 12.865 10.765 13.025 10.835 ;
        RECT 15.765 10.765 15.925 10.835 ;
        RECT 18.665 10.765 18.825 10.835 ;
        RECT 21.565 10.765 21.725 10.835 ;
        RECT 24.465 10.765 24.625 10.835 ;
        RECT 27.365 10.765 27.525 10.835 ;
        RECT 30.265 10.765 30.425 10.835 ;
        RECT 33.165 10.765 33.325 10.835 ;
        RECT 1.275 9.485 1.415 9.495 ;
        RECT 4.175 9.485 4.315 9.495 ;
        RECT 7.075 9.485 7.215 9.495 ;
        RECT 9.975 9.485 10.115 9.495 ;
        RECT 12.875 9.485 13.015 9.495 ;
        RECT 15.775 9.485 15.915 9.495 ;
        RECT 18.675 9.485 18.815 9.495 ;
        RECT 21.575 9.485 21.715 9.495 ;
        RECT 24.475 9.485 24.615 9.495 ;
        RECT 27.375 9.485 27.515 9.495 ;
        RECT 30.275 9.485 30.415 9.495 ;
        RECT 33.175 9.485 33.315 9.495 ;
        RECT 1.265 9.415 1.425 9.485 ;
        RECT 4.165 9.415 4.325 9.485 ;
        RECT 7.065 9.415 7.225 9.485 ;
        RECT 9.965 9.415 10.125 9.485 ;
        RECT 12.865 9.415 13.025 9.485 ;
        RECT 15.765 9.415 15.925 9.485 ;
        RECT 18.665 9.415 18.825 9.485 ;
        RECT 21.565 9.415 21.725 9.485 ;
        RECT 24.465 9.415 24.625 9.485 ;
        RECT 27.365 9.415 27.525 9.485 ;
        RECT 30.265 9.415 30.425 9.485 ;
        RECT 33.165 9.415 33.325 9.485 ;
        RECT 1.275 8.135 1.415 8.145 ;
        RECT 4.175 8.135 4.315 8.145 ;
        RECT 7.075 8.135 7.215 8.145 ;
        RECT 9.975 8.135 10.115 8.145 ;
        RECT 12.875 8.135 13.015 8.145 ;
        RECT 15.775 8.135 15.915 8.145 ;
        RECT 18.675 8.135 18.815 8.145 ;
        RECT 21.575 8.135 21.715 8.145 ;
        RECT 24.475 8.135 24.615 8.145 ;
        RECT 27.375 8.135 27.515 8.145 ;
        RECT 30.275 8.135 30.415 8.145 ;
        RECT 33.175 8.135 33.315 8.145 ;
        RECT 1.265 8.065 1.425 8.135 ;
        RECT 4.165 8.065 4.325 8.135 ;
        RECT 7.065 8.065 7.225 8.135 ;
        RECT 9.965 8.065 10.125 8.135 ;
        RECT 12.865 8.065 13.025 8.135 ;
        RECT 15.765 8.065 15.925 8.135 ;
        RECT 18.665 8.065 18.825 8.135 ;
        RECT 21.565 8.065 21.725 8.135 ;
        RECT 24.465 8.065 24.625 8.135 ;
        RECT 27.365 8.065 27.525 8.135 ;
        RECT 30.265 8.065 30.425 8.135 ;
        RECT 33.165 8.065 33.325 8.135 ;
        RECT 1.275 6.785 1.415 6.795 ;
        RECT 4.175 6.785 4.315 6.795 ;
        RECT 7.075 6.785 7.215 6.795 ;
        RECT 9.975 6.785 10.115 6.795 ;
        RECT 12.875 6.785 13.015 6.795 ;
        RECT 15.775 6.785 15.915 6.795 ;
        RECT 18.675 6.785 18.815 6.795 ;
        RECT 21.575 6.785 21.715 6.795 ;
        RECT 24.475 6.785 24.615 6.795 ;
        RECT 27.375 6.785 27.515 6.795 ;
        RECT 30.275 6.785 30.415 6.795 ;
        RECT 33.175 6.785 33.315 6.795 ;
        RECT 1.265 6.715 1.425 6.785 ;
        RECT 4.165 6.715 4.325 6.785 ;
        RECT 7.065 6.715 7.225 6.785 ;
        RECT 9.965 6.715 10.125 6.785 ;
        RECT 12.865 6.715 13.025 6.785 ;
        RECT 15.765 6.715 15.925 6.785 ;
        RECT 18.665 6.715 18.825 6.785 ;
        RECT 21.565 6.715 21.725 6.785 ;
        RECT 24.465 6.715 24.625 6.785 ;
        RECT 27.365 6.715 27.525 6.785 ;
        RECT 30.265 6.715 30.425 6.785 ;
        RECT 33.165 6.715 33.325 6.785 ;
        RECT 1.275 5.435 1.415 5.445 ;
        RECT 4.175 5.435 4.315 5.445 ;
        RECT 7.075 5.435 7.215 5.445 ;
        RECT 9.975 5.435 10.115 5.445 ;
        RECT 12.875 5.435 13.015 5.445 ;
        RECT 15.775 5.435 15.915 5.445 ;
        RECT 18.675 5.435 18.815 5.445 ;
        RECT 21.575 5.435 21.715 5.445 ;
        RECT 24.475 5.435 24.615 5.445 ;
        RECT 27.375 5.435 27.515 5.445 ;
        RECT 30.275 5.435 30.415 5.445 ;
        RECT 33.175 5.435 33.315 5.445 ;
        RECT 1.265 5.365 1.425 5.435 ;
        RECT 4.165 5.365 4.325 5.435 ;
        RECT 7.065 5.365 7.225 5.435 ;
        RECT 9.965 5.365 10.125 5.435 ;
        RECT 12.865 5.365 13.025 5.435 ;
        RECT 15.765 5.365 15.925 5.435 ;
        RECT 18.665 5.365 18.825 5.435 ;
        RECT 21.565 5.365 21.725 5.435 ;
        RECT 24.465 5.365 24.625 5.435 ;
        RECT 27.365 5.365 27.525 5.435 ;
        RECT 30.265 5.365 30.425 5.435 ;
        RECT 33.165 5.365 33.325 5.435 ;
        RECT 1.275 4.085 1.415 4.095 ;
        RECT 4.175 4.085 4.315 4.095 ;
        RECT 7.075 4.085 7.215 4.095 ;
        RECT 9.975 4.085 10.115 4.095 ;
        RECT 12.875 4.085 13.015 4.095 ;
        RECT 15.775 4.085 15.915 4.095 ;
        RECT 18.675 4.085 18.815 4.095 ;
        RECT 21.575 4.085 21.715 4.095 ;
        RECT 24.475 4.085 24.615 4.095 ;
        RECT 27.375 4.085 27.515 4.095 ;
        RECT 30.275 4.085 30.415 4.095 ;
        RECT 33.175 4.085 33.315 4.095 ;
        RECT 1.265 4.015 1.425 4.085 ;
        RECT 4.165 4.015 4.325 4.085 ;
        RECT 7.065 4.015 7.225 4.085 ;
        RECT 9.965 4.015 10.125 4.085 ;
        RECT 12.865 4.015 13.025 4.085 ;
        RECT 15.765 4.015 15.925 4.085 ;
        RECT 18.665 4.015 18.825 4.085 ;
        RECT 21.565 4.015 21.725 4.085 ;
        RECT 24.465 4.015 24.625 4.085 ;
        RECT 27.365 4.015 27.525 4.085 ;
        RECT 30.265 4.015 30.425 4.085 ;
        RECT 33.165 4.015 33.325 4.085 ;
        RECT 1.275 2.735 1.415 2.745 ;
        RECT 4.175 2.735 4.315 2.745 ;
        RECT 7.075 2.735 7.215 2.745 ;
        RECT 9.975 2.735 10.115 2.745 ;
        RECT 12.875 2.735 13.015 2.745 ;
        RECT 15.775 2.735 15.915 2.745 ;
        RECT 18.675 2.735 18.815 2.745 ;
        RECT 21.575 2.735 21.715 2.745 ;
        RECT 24.475 2.735 24.615 2.745 ;
        RECT 27.375 2.735 27.515 2.745 ;
        RECT 30.275 2.735 30.415 2.745 ;
        RECT 33.175 2.735 33.315 2.745 ;
        RECT 1.265 2.665 1.425 2.735 ;
        RECT 4.165 2.665 4.325 2.735 ;
        RECT 7.065 2.665 7.225 2.735 ;
        RECT 9.965 2.665 10.125 2.735 ;
        RECT 12.865 2.665 13.025 2.735 ;
        RECT 15.765 2.665 15.925 2.735 ;
        RECT 18.665 2.665 18.825 2.735 ;
        RECT 21.565 2.665 21.725 2.735 ;
        RECT 24.465 2.665 24.625 2.735 ;
        RECT 27.365 2.665 27.525 2.735 ;
        RECT 30.265 2.665 30.425 2.735 ;
        RECT 33.165 2.665 33.325 2.735 ;
        RECT 1.275 1.385 1.415 1.395 ;
        RECT 4.175 1.385 4.315 1.395 ;
        RECT 7.075 1.385 7.215 1.395 ;
        RECT 9.975 1.385 10.115 1.395 ;
        RECT 12.875 1.385 13.015 1.395 ;
        RECT 15.775 1.385 15.915 1.395 ;
        RECT 18.675 1.385 18.815 1.395 ;
        RECT 21.575 1.385 21.715 1.395 ;
        RECT 24.475 1.385 24.615 1.395 ;
        RECT 27.375 1.385 27.515 1.395 ;
        RECT 30.275 1.385 30.415 1.395 ;
        RECT 33.175 1.385 33.315 1.395 ;
        RECT 1.265 1.315 1.425 1.385 ;
        RECT 4.165 1.315 4.325 1.385 ;
        RECT 7.065 1.315 7.225 1.385 ;
        RECT 9.965 1.315 10.125 1.385 ;
        RECT 12.865 1.315 13.025 1.385 ;
        RECT 15.765 1.315 15.925 1.385 ;
        RECT 18.665 1.315 18.825 1.385 ;
        RECT 21.565 1.315 21.725 1.385 ;
        RECT 24.465 1.315 24.625 1.385 ;
        RECT 27.365 1.315 27.525 1.385 ;
        RECT 30.265 1.315 30.425 1.385 ;
        RECT 33.165 1.315 33.325 1.385 ;
        RECT 1.275 0.035 1.415 0.045 ;
        RECT 4.175 0.035 4.315 0.045 ;
        RECT 7.075 0.035 7.215 0.045 ;
        RECT 9.975 0.035 10.115 0.045 ;
        RECT 12.875 0.035 13.015 0.045 ;
        RECT 15.775 0.035 15.915 0.045 ;
        RECT 18.675 0.035 18.815 0.045 ;
        RECT 21.575 0.035 21.715 0.045 ;
        RECT 24.475 0.035 24.615 0.045 ;
        RECT 27.375 0.035 27.515 0.045 ;
        RECT 30.275 0.035 30.415 0.045 ;
        RECT 33.175 0.035 33.315 0.045 ;
        RECT 1.265 -0.035 1.425 0.035 ;
        RECT 4.165 -0.035 4.325 0.035 ;
        RECT 7.065 -0.035 7.225 0.035 ;
        RECT 9.965 -0.035 10.125 0.035 ;
        RECT 12.865 -0.035 13.025 0.035 ;
        RECT 15.765 -0.035 15.925 0.035 ;
        RECT 18.665 -0.035 18.825 0.035 ;
        RECT 21.565 -0.035 21.725 0.035 ;
        RECT 24.465 -0.035 24.625 0.035 ;
        RECT 27.365 -0.035 27.525 0.035 ;
        RECT 30.265 -0.035 30.425 0.035 ;
        RECT 33.165 -0.035 33.325 0.035 ;
      LAYER met1 ;
        RECT -0.275 20.215 34.625 20.285 ;
        RECT -0.275 18.865 34.625 18.935 ;
        RECT -0.275 17.515 34.625 17.585 ;
        RECT -0.275 16.165 34.625 16.235 ;
        RECT -0.275 14.815 34.625 14.885 ;
        RECT -0.275 13.465 34.625 13.535 ;
        RECT -0.275 12.115 34.625 12.185 ;
        RECT -0.275 10.765 34.625 10.835 ;
        RECT -0.275 9.415 34.625 9.485 ;
        RECT -0.275 8.065 34.625 8.135 ;
        RECT -0.275 6.715 34.625 6.785 ;
        RECT -0.275 5.365 34.625 5.435 ;
        RECT -0.275 4.015 34.625 4.085 ;
        RECT -0.275 2.665 34.625 2.735 ;
        RECT -0.275 1.315 34.625 1.385 ;
        RECT -0.275 -0.035 34.625 0.035 ;
    END
  END GND
  PIN RWL0_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 0.475 2.510 0.645 ;
        RECT 5.260 0.475 5.410 0.645 ;
        RECT 8.160 0.475 8.310 0.645 ;
        RECT 11.060 0.475 11.210 0.645 ;
        RECT 13.960 0.475 14.110 0.645 ;
        RECT 16.860 0.475 17.010 0.645 ;
        RECT 19.760 0.475 19.910 0.645 ;
        RECT 22.660 0.475 22.810 0.645 ;
        RECT 25.560 0.475 25.710 0.645 ;
        RECT 28.460 0.475 28.610 0.645 ;
        RECT 31.360 0.475 31.510 0.645 ;
        RECT 34.260 0.475 34.410 0.645 ;
      LAYER mcon ;
        RECT 2.360 0.480 2.510 0.645 ;
        RECT 8.160 0.480 8.310 0.645 ;
        RECT 13.960 0.480 14.110 0.645 ;
        RECT 19.760 0.480 19.910 0.645 ;
        RECT 25.560 0.480 25.710 0.645 ;
        RECT 31.360 0.480 31.510 0.645 ;
      LAYER met1 ;
        RECT 2.360 0.475 2.510 0.645 ;
        RECT 5.260 0.475 5.410 0.645 ;
        RECT 8.160 0.475 8.310 0.645 ;
        RECT 11.060 0.475 11.210 0.645 ;
        RECT 13.960 0.475 14.110 0.645 ;
        RECT 16.860 0.475 17.010 0.645 ;
        RECT 19.760 0.475 19.910 0.645 ;
        RECT 22.660 0.475 22.810 0.645 ;
        RECT 25.560 0.475 25.710 0.645 ;
        RECT 28.460 0.475 28.610 0.645 ;
        RECT 31.360 0.475 31.510 0.645 ;
        RECT 34.260 0.475 34.410 0.645 ;
      LAYER met2 ;
        RECT -0.275 0.475 34.760 0.645 ;
    END
  END RWL0_0
  PIN RWL1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 0.475 0.330 0.645 ;
        RECT 3.080 0.475 3.230 0.645 ;
        RECT 5.980 0.475 6.130 0.645 ;
        RECT 8.880 0.475 9.030 0.645 ;
        RECT 11.780 0.475 11.930 0.645 ;
        RECT 14.680 0.475 14.830 0.645 ;
        RECT 17.580 0.475 17.730 0.645 ;
        RECT 20.480 0.475 20.630 0.645 ;
        RECT 23.380 0.475 23.530 0.645 ;
        RECT 26.280 0.475 26.430 0.645 ;
        RECT 29.180 0.475 29.330 0.645 ;
        RECT 32.080 0.475 32.230 0.645 ;
      LAYER met1 ;
        POLYGON 2.310 0.945 2.310 0.775 2.140 0.775 ;
        RECT 2.310 0.775 2.560 0.945 ;
        POLYGON 2.560 0.945 2.730 0.775 2.560 0.775 ;
        POLYGON 5.210 0.945 5.210 0.775 5.040 0.775 ;
        RECT 5.210 0.775 5.460 0.945 ;
        POLYGON 5.460 0.945 5.630 0.775 5.460 0.775 ;
        POLYGON 8.110 0.945 8.110 0.775 7.940 0.775 ;
        RECT 8.110 0.775 8.360 0.945 ;
        POLYGON 8.360 0.945 8.530 0.775 8.360 0.775 ;
        POLYGON 11.010 0.945 11.010 0.775 10.840 0.775 ;
        RECT 11.010 0.775 11.260 0.945 ;
        POLYGON 11.260 0.945 11.430 0.775 11.260 0.775 ;
        POLYGON 13.910 0.945 13.910 0.775 13.740 0.775 ;
        RECT 13.910 0.775 14.160 0.945 ;
        POLYGON 14.160 0.945 14.330 0.775 14.160 0.775 ;
        POLYGON 16.810 0.945 16.810 0.775 16.640 0.775 ;
        RECT 16.810 0.775 17.060 0.945 ;
        POLYGON 17.060 0.945 17.230 0.775 17.060 0.775 ;
        POLYGON 19.710 0.945 19.710 0.775 19.540 0.775 ;
        RECT 19.710 0.775 19.960 0.945 ;
        POLYGON 19.960 0.945 20.130 0.775 19.960 0.775 ;
        POLYGON 22.610 0.945 22.610 0.775 22.440 0.775 ;
        RECT 22.610 0.775 22.860 0.945 ;
        POLYGON 22.860 0.945 23.030 0.775 22.860 0.775 ;
        POLYGON 25.510 0.945 25.510 0.775 25.340 0.775 ;
        RECT 25.510 0.775 25.760 0.945 ;
        POLYGON 25.760 0.945 25.930 0.775 25.760 0.775 ;
        POLYGON 28.410 0.945 28.410 0.775 28.240 0.775 ;
        RECT 28.410 0.775 28.660 0.945 ;
        POLYGON 28.660 0.945 28.830 0.775 28.660 0.775 ;
        POLYGON 31.310 0.945 31.310 0.775 31.140 0.775 ;
        RECT 31.310 0.775 31.560 0.945 ;
        POLYGON 31.560 0.945 31.730 0.775 31.560 0.775 ;
        POLYGON 34.210 0.945 34.210 0.775 34.040 0.775 ;
        RECT 34.210 0.775 34.460 0.945 ;
        POLYGON 34.460 0.945 34.630 0.775 34.460 0.775 ;
        POLYGON 2.140 0.775 2.140 0.645 2.010 0.645 ;
        RECT 2.140 0.645 2.230 0.775 ;
        POLYGON 2.230 0.775 2.360 0.775 2.230 0.645 ;
        POLYGON 2.510 0.775 2.640 0.775 2.640 0.645 ;
        RECT 2.640 0.645 2.730 0.775 ;
        POLYGON 2.730 0.775 2.860 0.645 2.730 0.645 ;
        POLYGON 5.040 0.775 5.040 0.645 4.910 0.645 ;
        RECT 5.040 0.645 5.130 0.775 ;
        POLYGON 5.130 0.775 5.260 0.775 5.130 0.645 ;
        POLYGON 5.410 0.775 5.540 0.775 5.540 0.645 ;
        RECT 5.540 0.645 5.630 0.775 ;
        POLYGON 5.630 0.775 5.760 0.645 5.630 0.645 ;
        POLYGON 7.940 0.775 7.940 0.645 7.810 0.645 ;
        RECT 7.940 0.645 8.030 0.775 ;
        POLYGON 8.030 0.775 8.160 0.775 8.030 0.645 ;
        POLYGON 8.310 0.775 8.440 0.775 8.440 0.645 ;
        RECT 8.440 0.645 8.530 0.775 ;
        POLYGON 8.530 0.775 8.660 0.645 8.530 0.645 ;
        POLYGON 10.840 0.775 10.840 0.645 10.710 0.645 ;
        RECT 10.840 0.645 10.930 0.775 ;
        POLYGON 10.930 0.775 11.060 0.775 10.930 0.645 ;
        POLYGON 11.210 0.775 11.340 0.775 11.340 0.645 ;
        RECT 11.340 0.645 11.430 0.775 ;
        POLYGON 11.430 0.775 11.560 0.645 11.430 0.645 ;
        POLYGON 13.740 0.775 13.740 0.645 13.610 0.645 ;
        RECT 13.740 0.645 13.830 0.775 ;
        POLYGON 13.830 0.775 13.960 0.775 13.830 0.645 ;
        POLYGON 14.110 0.775 14.240 0.775 14.240 0.645 ;
        RECT 14.240 0.645 14.330 0.775 ;
        POLYGON 14.330 0.775 14.460 0.645 14.330 0.645 ;
        POLYGON 16.640 0.775 16.640 0.645 16.510 0.645 ;
        RECT 16.640 0.645 16.730 0.775 ;
        POLYGON 16.730 0.775 16.860 0.775 16.730 0.645 ;
        POLYGON 17.010 0.775 17.140 0.775 17.140 0.645 ;
        RECT 17.140 0.645 17.230 0.775 ;
        POLYGON 17.230 0.775 17.360 0.645 17.230 0.645 ;
        POLYGON 19.540 0.775 19.540 0.645 19.410 0.645 ;
        RECT 19.540 0.645 19.630 0.775 ;
        POLYGON 19.630 0.775 19.760 0.775 19.630 0.645 ;
        POLYGON 19.910 0.775 20.040 0.775 20.040 0.645 ;
        RECT 20.040 0.645 20.130 0.775 ;
        POLYGON 20.130 0.775 20.260 0.645 20.130 0.645 ;
        POLYGON 22.440 0.775 22.440 0.645 22.310 0.645 ;
        RECT 22.440 0.645 22.530 0.775 ;
        POLYGON 22.530 0.775 22.660 0.775 22.530 0.645 ;
        POLYGON 22.810 0.775 22.940 0.775 22.940 0.645 ;
        RECT 22.940 0.645 23.030 0.775 ;
        POLYGON 23.030 0.775 23.160 0.645 23.030 0.645 ;
        POLYGON 25.340 0.775 25.340 0.645 25.210 0.645 ;
        RECT 25.340 0.645 25.430 0.775 ;
        POLYGON 25.430 0.775 25.560 0.775 25.430 0.645 ;
        POLYGON 25.710 0.775 25.840 0.775 25.840 0.645 ;
        RECT 25.840 0.645 25.930 0.775 ;
        POLYGON 25.930 0.775 26.060 0.645 25.930 0.645 ;
        POLYGON 28.240 0.775 28.240 0.645 28.110 0.645 ;
        RECT 28.240 0.645 28.330 0.775 ;
        POLYGON 28.330 0.775 28.460 0.775 28.330 0.645 ;
        POLYGON 28.610 0.775 28.740 0.775 28.740 0.645 ;
        RECT 28.740 0.645 28.830 0.775 ;
        POLYGON 28.830 0.775 28.960 0.645 28.830 0.645 ;
        POLYGON 31.140 0.775 31.140 0.645 31.010 0.645 ;
        RECT 31.140 0.645 31.230 0.775 ;
        POLYGON 31.230 0.775 31.360 0.775 31.230 0.645 ;
        POLYGON 31.510 0.775 31.640 0.775 31.640 0.645 ;
        RECT 31.640 0.645 31.730 0.775 ;
        POLYGON 31.730 0.775 31.860 0.645 31.730 0.645 ;
        POLYGON 34.040 0.775 34.040 0.645 33.910 0.645 ;
        RECT 34.040 0.645 34.130 0.775 ;
        POLYGON 34.130 0.775 34.260 0.775 34.130 0.645 ;
        POLYGON 34.410 0.775 34.540 0.775 34.540 0.645 ;
        RECT 34.540 0.645 34.630 0.775 ;
        POLYGON 34.630 0.775 34.760 0.645 34.630 0.645 ;
        RECT -0.275 0.475 2.060 0.645 ;
        POLYGON 2.060 0.645 2.230 0.645 2.060 0.475 ;
        POLYGON 2.640 0.645 2.810 0.645 2.810 0.475 ;
        RECT 2.810 0.475 4.960 0.645 ;
        POLYGON 4.960 0.645 5.130 0.645 4.960 0.475 ;
        RECT 5.525 0.475 7.860 0.645 ;
        POLYGON 7.860 0.645 8.030 0.645 7.860 0.475 ;
        POLYGON 8.440 0.645 8.610 0.645 8.610 0.475 ;
        RECT 8.610 0.475 10.760 0.645 ;
        POLYGON 10.760 0.645 10.930 0.645 10.760 0.475 ;
        RECT 11.325 0.475 13.660 0.645 ;
        POLYGON 13.660 0.645 13.830 0.645 13.660 0.475 ;
        POLYGON 14.240 0.645 14.410 0.645 14.410 0.475 ;
        RECT 14.410 0.475 16.560 0.645 ;
        POLYGON 16.560 0.645 16.730 0.645 16.560 0.475 ;
        RECT 17.125 0.475 19.460 0.645 ;
        POLYGON 19.460 0.645 19.630 0.645 19.460 0.475 ;
        POLYGON 20.040 0.645 20.210 0.645 20.210 0.475 ;
        RECT 20.210 0.475 22.360 0.645 ;
        POLYGON 22.360 0.645 22.530 0.645 22.360 0.475 ;
        RECT 22.925 0.475 25.260 0.645 ;
        POLYGON 25.260 0.645 25.430 0.645 25.260 0.475 ;
        POLYGON 25.840 0.645 26.010 0.645 26.010 0.475 ;
        RECT 26.010 0.475 28.160 0.645 ;
        POLYGON 28.160 0.645 28.330 0.645 28.160 0.475 ;
        RECT 28.725 0.475 31.060 0.645 ;
        POLYGON 31.060 0.645 31.230 0.645 31.060 0.475 ;
        POLYGON 31.640 0.645 31.810 0.645 31.810 0.475 ;
        RECT 31.810 0.475 33.960 0.645 ;
        POLYGON 33.960 0.645 34.130 0.645 33.960 0.475 ;
        POLYGON 34.540 0.645 34.710 0.645 34.710 0.475 ;
        RECT 34.710 0.475 34.760 0.645 ;
    END
  END RWL1_0
  PIN RBL0_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 2.650 20.405 2.725 20.615 ;
        RECT 2.650 19.055 2.725 19.265 ;
        RECT 2.650 17.705 2.725 17.915 ;
        RECT 2.650 16.355 2.725 16.565 ;
        RECT 2.650 15.005 2.725 15.215 ;
        RECT 2.650 13.655 2.725 13.865 ;
        RECT 2.650 12.305 2.725 12.515 ;
        RECT 2.650 10.955 2.725 11.165 ;
        RECT 2.650 9.605 2.725 9.815 ;
        RECT 2.650 8.255 2.725 8.465 ;
        RECT 2.650 6.905 2.725 7.115 ;
        RECT 2.650 5.555 2.725 5.765 ;
        RECT 2.650 4.205 2.725 4.415 ;
        RECT 2.650 2.855 2.725 3.065 ;
        RECT 2.650 1.505 2.725 1.715 ;
        RECT 2.650 0.155 2.725 0.365 ;
    END
  END RBL0_0
  PIN RBL1_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT -0.035 20.405 0.040 20.615 ;
        RECT -0.035 19.055 0.040 19.265 ;
        RECT -0.035 17.705 0.040 17.915 ;
        RECT -0.035 16.355 0.040 16.565 ;
        RECT -0.035 15.005 0.040 15.215 ;
        RECT -0.035 13.655 0.040 13.865 ;
        RECT -0.035 12.305 0.040 12.515 ;
        RECT -0.035 10.955 0.040 11.165 ;
        RECT -0.035 9.605 0.040 9.815 ;
        RECT -0.035 8.255 0.040 8.465 ;
        RECT -0.035 6.905 0.040 7.115 ;
        RECT -0.035 5.555 0.040 5.765 ;
        RECT -0.035 4.205 0.040 4.415 ;
        RECT -0.035 2.855 0.040 3.065 ;
        RECT -0.035 1.505 0.040 1.715 ;
        RECT -0.035 0.155 0.040 0.365 ;
    END
  END RBL1_0
  PIN WBL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 2.285 21.135 2.360 21.280 ;
        RECT 2.285 19.785 2.360 19.930 ;
        RECT 2.285 18.435 2.360 18.580 ;
        RECT 2.285 17.085 2.360 17.230 ;
        RECT 2.285 15.735 2.360 15.880 ;
        RECT 2.285 14.385 2.360 14.530 ;
        RECT 2.285 13.035 2.360 13.180 ;
        RECT 2.285 11.685 2.360 11.830 ;
        RECT 2.285 10.335 2.360 10.480 ;
        RECT 2.285 8.985 2.360 9.130 ;
        RECT 2.285 7.635 2.360 7.780 ;
        RECT 2.285 6.285 2.360 6.430 ;
        RECT 2.285 4.935 2.360 5.080 ;
        RECT 2.285 3.585 2.360 3.730 ;
        RECT 2.285 2.235 2.360 2.380 ;
        RECT 2.285 0.885 2.360 1.030 ;
    END
  END WBL_0
  PIN WBLb_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 0.335 21.135 0.410 21.275 ;
        RECT 0.335 19.785 0.410 19.925 ;
        RECT 0.335 18.435 0.410 18.575 ;
        RECT 0.335 17.085 0.410 17.225 ;
        RECT 0.335 15.735 0.410 15.875 ;
        RECT 0.335 14.385 0.410 14.525 ;
        RECT 0.335 13.035 0.410 13.175 ;
        RECT 0.335 11.685 0.410 11.825 ;
        RECT 0.335 10.335 0.410 10.475 ;
        RECT 0.335 8.985 0.410 9.125 ;
        RECT 0.335 7.635 0.410 7.775 ;
        RECT 0.335 6.285 0.410 6.425 ;
        RECT 0.335 4.935 0.410 5.075 ;
        RECT 0.335 3.585 0.410 3.725 ;
        RECT 0.335 2.235 0.410 2.375 ;
        RECT 0.335 0.885 0.410 1.025 ;
    END
  END WBLb_0
  PIN RWL0_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 1.825 2.510 1.995 ;
        RECT 5.260 1.825 5.410 1.995 ;
        RECT 8.160 1.825 8.310 1.995 ;
        RECT 11.060 1.825 11.210 1.995 ;
        RECT 13.960 1.825 14.110 1.995 ;
        RECT 16.860 1.825 17.010 1.995 ;
        RECT 19.760 1.825 19.910 1.995 ;
        RECT 22.660 1.825 22.810 1.995 ;
        RECT 25.560 1.825 25.710 1.995 ;
        RECT 28.460 1.825 28.610 1.995 ;
        RECT 31.360 1.825 31.510 1.995 ;
        RECT 34.260 1.825 34.410 1.995 ;
      LAYER mcon ;
        RECT 2.360 1.830 2.510 1.995 ;
        RECT 8.160 1.830 8.310 1.995 ;
        RECT 13.960 1.830 14.110 1.995 ;
        RECT 19.760 1.830 19.910 1.995 ;
        RECT 25.560 1.830 25.710 1.995 ;
        RECT 31.360 1.830 31.510 1.995 ;
      LAYER met1 ;
        RECT 2.360 1.825 2.510 1.995 ;
        RECT 5.260 1.825 5.410 1.995 ;
        RECT 8.160 1.825 8.310 1.995 ;
        RECT 11.060 1.825 11.210 1.995 ;
        RECT 13.960 1.825 14.110 1.995 ;
        RECT 16.860 1.825 17.010 1.995 ;
        RECT 19.760 1.825 19.910 1.995 ;
        RECT 22.660 1.825 22.810 1.995 ;
        RECT 25.560 1.825 25.710 1.995 ;
        RECT 28.460 1.825 28.610 1.995 ;
        RECT 31.360 1.825 31.510 1.995 ;
        RECT 34.260 1.825 34.410 1.995 ;
      LAYER met2 ;
        RECT -0.275 1.825 34.760 1.995 ;
    END
  END RWL0_1
  PIN RWL1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 1.825 0.330 1.995 ;
        RECT 3.080 1.825 3.230 1.995 ;
        RECT 5.980 1.825 6.130 1.995 ;
        RECT 8.880 1.825 9.030 1.995 ;
        RECT 11.780 1.825 11.930 1.995 ;
        RECT 14.680 1.825 14.830 1.995 ;
        RECT 17.580 1.825 17.730 1.995 ;
        RECT 20.480 1.825 20.630 1.995 ;
        RECT 23.380 1.825 23.530 1.995 ;
        RECT 26.280 1.825 26.430 1.995 ;
        RECT 29.180 1.825 29.330 1.995 ;
        RECT 32.080 1.825 32.230 1.995 ;
      LAYER met1 ;
        POLYGON 2.310 2.295 2.310 2.125 2.140 2.125 ;
        RECT 2.310 2.125 2.560 2.295 ;
        POLYGON 2.560 2.295 2.730 2.125 2.560 2.125 ;
        POLYGON 5.210 2.295 5.210 2.125 5.040 2.125 ;
        RECT 5.210 2.125 5.460 2.295 ;
        POLYGON 5.460 2.295 5.630 2.125 5.460 2.125 ;
        POLYGON 8.110 2.295 8.110 2.125 7.940 2.125 ;
        RECT 8.110 2.125 8.360 2.295 ;
        POLYGON 8.360 2.295 8.530 2.125 8.360 2.125 ;
        POLYGON 11.010 2.295 11.010 2.125 10.840 2.125 ;
        RECT 11.010 2.125 11.260 2.295 ;
        POLYGON 11.260 2.295 11.430 2.125 11.260 2.125 ;
        POLYGON 13.910 2.295 13.910 2.125 13.740 2.125 ;
        RECT 13.910 2.125 14.160 2.295 ;
        POLYGON 14.160 2.295 14.330 2.125 14.160 2.125 ;
        POLYGON 16.810 2.295 16.810 2.125 16.640 2.125 ;
        RECT 16.810 2.125 17.060 2.295 ;
        POLYGON 17.060 2.295 17.230 2.125 17.060 2.125 ;
        POLYGON 19.710 2.295 19.710 2.125 19.540 2.125 ;
        RECT 19.710 2.125 19.960 2.295 ;
        POLYGON 19.960 2.295 20.130 2.125 19.960 2.125 ;
        POLYGON 22.610 2.295 22.610 2.125 22.440 2.125 ;
        RECT 22.610 2.125 22.860 2.295 ;
        POLYGON 22.860 2.295 23.030 2.125 22.860 2.125 ;
        POLYGON 25.510 2.295 25.510 2.125 25.340 2.125 ;
        RECT 25.510 2.125 25.760 2.295 ;
        POLYGON 25.760 2.295 25.930 2.125 25.760 2.125 ;
        POLYGON 28.410 2.295 28.410 2.125 28.240 2.125 ;
        RECT 28.410 2.125 28.660 2.295 ;
        POLYGON 28.660 2.295 28.830 2.125 28.660 2.125 ;
        POLYGON 31.310 2.295 31.310 2.125 31.140 2.125 ;
        RECT 31.310 2.125 31.560 2.295 ;
        POLYGON 31.560 2.295 31.730 2.125 31.560 2.125 ;
        POLYGON 34.210 2.295 34.210 2.125 34.040 2.125 ;
        RECT 34.210 2.125 34.460 2.295 ;
        POLYGON 34.460 2.295 34.630 2.125 34.460 2.125 ;
        POLYGON 2.140 2.125 2.140 1.995 2.010 1.995 ;
        RECT 2.140 1.995 2.230 2.125 ;
        POLYGON 2.230 2.125 2.360 2.125 2.230 1.995 ;
        POLYGON 2.510 2.125 2.640 2.125 2.640 1.995 ;
        RECT 2.640 1.995 2.730 2.125 ;
        POLYGON 2.730 2.125 2.860 1.995 2.730 1.995 ;
        POLYGON 5.040 2.125 5.040 1.995 4.910 1.995 ;
        RECT 5.040 1.995 5.130 2.125 ;
        POLYGON 5.130 2.125 5.260 2.125 5.130 1.995 ;
        POLYGON 5.410 2.125 5.540 2.125 5.540 1.995 ;
        RECT 5.540 1.995 5.630 2.125 ;
        POLYGON 5.630 2.125 5.760 1.995 5.630 1.995 ;
        POLYGON 7.940 2.125 7.940 1.995 7.810 1.995 ;
        RECT 7.940 1.995 8.030 2.125 ;
        POLYGON 8.030 2.125 8.160 2.125 8.030 1.995 ;
        POLYGON 8.310 2.125 8.440 2.125 8.440 1.995 ;
        RECT 8.440 1.995 8.530 2.125 ;
        POLYGON 8.530 2.125 8.660 1.995 8.530 1.995 ;
        POLYGON 10.840 2.125 10.840 1.995 10.710 1.995 ;
        RECT 10.840 1.995 10.930 2.125 ;
        POLYGON 10.930 2.125 11.060 2.125 10.930 1.995 ;
        POLYGON 11.210 2.125 11.340 2.125 11.340 1.995 ;
        RECT 11.340 1.995 11.430 2.125 ;
        POLYGON 11.430 2.125 11.560 1.995 11.430 1.995 ;
        POLYGON 13.740 2.125 13.740 1.995 13.610 1.995 ;
        RECT 13.740 1.995 13.830 2.125 ;
        POLYGON 13.830 2.125 13.960 2.125 13.830 1.995 ;
        POLYGON 14.110 2.125 14.240 2.125 14.240 1.995 ;
        RECT 14.240 1.995 14.330 2.125 ;
        POLYGON 14.330 2.125 14.460 1.995 14.330 1.995 ;
        POLYGON 16.640 2.125 16.640 1.995 16.510 1.995 ;
        RECT 16.640 1.995 16.730 2.125 ;
        POLYGON 16.730 2.125 16.860 2.125 16.730 1.995 ;
        POLYGON 17.010 2.125 17.140 2.125 17.140 1.995 ;
        RECT 17.140 1.995 17.230 2.125 ;
        POLYGON 17.230 2.125 17.360 1.995 17.230 1.995 ;
        POLYGON 19.540 2.125 19.540 1.995 19.410 1.995 ;
        RECT 19.540 1.995 19.630 2.125 ;
        POLYGON 19.630 2.125 19.760 2.125 19.630 1.995 ;
        POLYGON 19.910 2.125 20.040 2.125 20.040 1.995 ;
        RECT 20.040 1.995 20.130 2.125 ;
        POLYGON 20.130 2.125 20.260 1.995 20.130 1.995 ;
        POLYGON 22.440 2.125 22.440 1.995 22.310 1.995 ;
        RECT 22.440 1.995 22.530 2.125 ;
        POLYGON 22.530 2.125 22.660 2.125 22.530 1.995 ;
        POLYGON 22.810 2.125 22.940 2.125 22.940 1.995 ;
        RECT 22.940 1.995 23.030 2.125 ;
        POLYGON 23.030 2.125 23.160 1.995 23.030 1.995 ;
        POLYGON 25.340 2.125 25.340 1.995 25.210 1.995 ;
        RECT 25.340 1.995 25.430 2.125 ;
        POLYGON 25.430 2.125 25.560 2.125 25.430 1.995 ;
        POLYGON 25.710 2.125 25.840 2.125 25.840 1.995 ;
        RECT 25.840 1.995 25.930 2.125 ;
        POLYGON 25.930 2.125 26.060 1.995 25.930 1.995 ;
        POLYGON 28.240 2.125 28.240 1.995 28.110 1.995 ;
        RECT 28.240 1.995 28.330 2.125 ;
        POLYGON 28.330 2.125 28.460 2.125 28.330 1.995 ;
        POLYGON 28.610 2.125 28.740 2.125 28.740 1.995 ;
        RECT 28.740 1.995 28.830 2.125 ;
        POLYGON 28.830 2.125 28.960 1.995 28.830 1.995 ;
        POLYGON 31.140 2.125 31.140 1.995 31.010 1.995 ;
        RECT 31.140 1.995 31.230 2.125 ;
        POLYGON 31.230 2.125 31.360 2.125 31.230 1.995 ;
        POLYGON 31.510 2.125 31.640 2.125 31.640 1.995 ;
        RECT 31.640 1.995 31.730 2.125 ;
        POLYGON 31.730 2.125 31.860 1.995 31.730 1.995 ;
        POLYGON 34.040 2.125 34.040 1.995 33.910 1.995 ;
        RECT 34.040 1.995 34.130 2.125 ;
        POLYGON 34.130 2.125 34.260 2.125 34.130 1.995 ;
        POLYGON 34.410 2.125 34.540 2.125 34.540 1.995 ;
        RECT 34.540 1.995 34.630 2.125 ;
        POLYGON 34.630 2.125 34.760 1.995 34.630 1.995 ;
        RECT -0.275 1.825 2.060 1.995 ;
        POLYGON 2.060 1.995 2.230 1.995 2.060 1.825 ;
        POLYGON 2.640 1.995 2.810 1.995 2.810 1.825 ;
        RECT 2.810 1.825 4.960 1.995 ;
        POLYGON 4.960 1.995 5.130 1.995 4.960 1.825 ;
        RECT 5.525 1.825 7.860 1.995 ;
        POLYGON 7.860 1.995 8.030 1.995 7.860 1.825 ;
        POLYGON 8.440 1.995 8.610 1.995 8.610 1.825 ;
        RECT 8.610 1.825 10.760 1.995 ;
        POLYGON 10.760 1.995 10.930 1.995 10.760 1.825 ;
        RECT 11.325 1.825 13.660 1.995 ;
        POLYGON 13.660 1.995 13.830 1.995 13.660 1.825 ;
        POLYGON 14.240 1.995 14.410 1.995 14.410 1.825 ;
        RECT 14.410 1.825 16.560 1.995 ;
        POLYGON 16.560 1.995 16.730 1.995 16.560 1.825 ;
        RECT 17.125 1.825 19.460 1.995 ;
        POLYGON 19.460 1.995 19.630 1.995 19.460 1.825 ;
        POLYGON 20.040 1.995 20.210 1.995 20.210 1.825 ;
        RECT 20.210 1.825 22.360 1.995 ;
        POLYGON 22.360 1.995 22.530 1.995 22.360 1.825 ;
        RECT 22.925 1.825 25.260 1.995 ;
        POLYGON 25.260 1.995 25.430 1.995 25.260 1.825 ;
        POLYGON 25.840 1.995 26.010 1.995 26.010 1.825 ;
        RECT 26.010 1.825 28.160 1.995 ;
        POLYGON 28.160 1.995 28.330 1.995 28.160 1.825 ;
        RECT 28.725 1.825 31.060 1.995 ;
        POLYGON 31.060 1.995 31.230 1.995 31.060 1.825 ;
        POLYGON 31.640 1.995 31.810 1.995 31.810 1.825 ;
        RECT 31.810 1.825 33.960 1.995 ;
        POLYGON 33.960 1.995 34.130 1.995 33.960 1.825 ;
        POLYGON 34.540 1.995 34.710 1.995 34.710 1.825 ;
        RECT 34.710 1.825 34.760 1.995 ;
    END
  END RWL1_1
  PIN RWL0_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 3.175 2.510 3.345 ;
        RECT 5.260 3.175 5.410 3.345 ;
        RECT 8.160 3.175 8.310 3.345 ;
        RECT 11.060 3.175 11.210 3.345 ;
        RECT 13.960 3.175 14.110 3.345 ;
        RECT 16.860 3.175 17.010 3.345 ;
        RECT 19.760 3.175 19.910 3.345 ;
        RECT 22.660 3.175 22.810 3.345 ;
        RECT 25.560 3.175 25.710 3.345 ;
        RECT 28.460 3.175 28.610 3.345 ;
        RECT 31.360 3.175 31.510 3.345 ;
        RECT 34.260 3.175 34.410 3.345 ;
      LAYER mcon ;
        RECT 2.360 3.180 2.510 3.345 ;
        RECT 8.160 3.180 8.310 3.345 ;
        RECT 13.960 3.180 14.110 3.345 ;
        RECT 19.760 3.180 19.910 3.345 ;
        RECT 25.560 3.180 25.710 3.345 ;
        RECT 31.360 3.180 31.510 3.345 ;
      LAYER met1 ;
        RECT 2.360 3.175 2.510 3.345 ;
        RECT 5.260 3.175 5.410 3.345 ;
        RECT 8.160 3.175 8.310 3.345 ;
        RECT 11.060 3.175 11.210 3.345 ;
        RECT 13.960 3.175 14.110 3.345 ;
        RECT 16.860 3.175 17.010 3.345 ;
        RECT 19.760 3.175 19.910 3.345 ;
        RECT 22.660 3.175 22.810 3.345 ;
        RECT 25.560 3.175 25.710 3.345 ;
        RECT 28.460 3.175 28.610 3.345 ;
        RECT 31.360 3.175 31.510 3.345 ;
        RECT 34.260 3.175 34.410 3.345 ;
      LAYER met2 ;
        RECT -0.275 3.175 34.760 3.345 ;
    END
  END RWL0_2
  PIN RWL1_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 3.175 0.330 3.345 ;
        RECT 3.080 3.175 3.230 3.345 ;
        RECT 5.980 3.175 6.130 3.345 ;
        RECT 8.880 3.175 9.030 3.345 ;
        RECT 11.780 3.175 11.930 3.345 ;
        RECT 14.680 3.175 14.830 3.345 ;
        RECT 17.580 3.175 17.730 3.345 ;
        RECT 20.480 3.175 20.630 3.345 ;
        RECT 23.380 3.175 23.530 3.345 ;
        RECT 26.280 3.175 26.430 3.345 ;
        RECT 29.180 3.175 29.330 3.345 ;
        RECT 32.080 3.175 32.230 3.345 ;
      LAYER met1 ;
        POLYGON 2.310 3.645 2.310 3.475 2.140 3.475 ;
        RECT 2.310 3.475 2.560 3.645 ;
        POLYGON 2.560 3.645 2.730 3.475 2.560 3.475 ;
        POLYGON 5.210 3.645 5.210 3.475 5.040 3.475 ;
        RECT 5.210 3.475 5.460 3.645 ;
        POLYGON 5.460 3.645 5.630 3.475 5.460 3.475 ;
        POLYGON 8.110 3.645 8.110 3.475 7.940 3.475 ;
        RECT 8.110 3.475 8.360 3.645 ;
        POLYGON 8.360 3.645 8.530 3.475 8.360 3.475 ;
        POLYGON 11.010 3.645 11.010 3.475 10.840 3.475 ;
        RECT 11.010 3.475 11.260 3.645 ;
        POLYGON 11.260 3.645 11.430 3.475 11.260 3.475 ;
        POLYGON 13.910 3.645 13.910 3.475 13.740 3.475 ;
        RECT 13.910 3.475 14.160 3.645 ;
        POLYGON 14.160 3.645 14.330 3.475 14.160 3.475 ;
        POLYGON 16.810 3.645 16.810 3.475 16.640 3.475 ;
        RECT 16.810 3.475 17.060 3.645 ;
        POLYGON 17.060 3.645 17.230 3.475 17.060 3.475 ;
        POLYGON 19.710 3.645 19.710 3.475 19.540 3.475 ;
        RECT 19.710 3.475 19.960 3.645 ;
        POLYGON 19.960 3.645 20.130 3.475 19.960 3.475 ;
        POLYGON 22.610 3.645 22.610 3.475 22.440 3.475 ;
        RECT 22.610 3.475 22.860 3.645 ;
        POLYGON 22.860 3.645 23.030 3.475 22.860 3.475 ;
        POLYGON 25.510 3.645 25.510 3.475 25.340 3.475 ;
        RECT 25.510 3.475 25.760 3.645 ;
        POLYGON 25.760 3.645 25.930 3.475 25.760 3.475 ;
        POLYGON 28.410 3.645 28.410 3.475 28.240 3.475 ;
        RECT 28.410 3.475 28.660 3.645 ;
        POLYGON 28.660 3.645 28.830 3.475 28.660 3.475 ;
        POLYGON 31.310 3.645 31.310 3.475 31.140 3.475 ;
        RECT 31.310 3.475 31.560 3.645 ;
        POLYGON 31.560 3.645 31.730 3.475 31.560 3.475 ;
        POLYGON 34.210 3.645 34.210 3.475 34.040 3.475 ;
        RECT 34.210 3.475 34.460 3.645 ;
        POLYGON 34.460 3.645 34.630 3.475 34.460 3.475 ;
        POLYGON 2.140 3.475 2.140 3.345 2.010 3.345 ;
        RECT 2.140 3.345 2.230 3.475 ;
        POLYGON 2.230 3.475 2.360 3.475 2.230 3.345 ;
        POLYGON 2.510 3.475 2.640 3.475 2.640 3.345 ;
        RECT 2.640 3.345 2.730 3.475 ;
        POLYGON 2.730 3.475 2.860 3.345 2.730 3.345 ;
        POLYGON 5.040 3.475 5.040 3.345 4.910 3.345 ;
        RECT 5.040 3.345 5.130 3.475 ;
        POLYGON 5.130 3.475 5.260 3.475 5.130 3.345 ;
        POLYGON 5.410 3.475 5.540 3.475 5.540 3.345 ;
        RECT 5.540 3.345 5.630 3.475 ;
        POLYGON 5.630 3.475 5.760 3.345 5.630 3.345 ;
        POLYGON 7.940 3.475 7.940 3.345 7.810 3.345 ;
        RECT 7.940 3.345 8.030 3.475 ;
        POLYGON 8.030 3.475 8.160 3.475 8.030 3.345 ;
        POLYGON 8.310 3.475 8.440 3.475 8.440 3.345 ;
        RECT 8.440 3.345 8.530 3.475 ;
        POLYGON 8.530 3.475 8.660 3.345 8.530 3.345 ;
        POLYGON 10.840 3.475 10.840 3.345 10.710 3.345 ;
        RECT 10.840 3.345 10.930 3.475 ;
        POLYGON 10.930 3.475 11.060 3.475 10.930 3.345 ;
        POLYGON 11.210 3.475 11.340 3.475 11.340 3.345 ;
        RECT 11.340 3.345 11.430 3.475 ;
        POLYGON 11.430 3.475 11.560 3.345 11.430 3.345 ;
        POLYGON 13.740 3.475 13.740 3.345 13.610 3.345 ;
        RECT 13.740 3.345 13.830 3.475 ;
        POLYGON 13.830 3.475 13.960 3.475 13.830 3.345 ;
        POLYGON 14.110 3.475 14.240 3.475 14.240 3.345 ;
        RECT 14.240 3.345 14.330 3.475 ;
        POLYGON 14.330 3.475 14.460 3.345 14.330 3.345 ;
        POLYGON 16.640 3.475 16.640 3.345 16.510 3.345 ;
        RECT 16.640 3.345 16.730 3.475 ;
        POLYGON 16.730 3.475 16.860 3.475 16.730 3.345 ;
        POLYGON 17.010 3.475 17.140 3.475 17.140 3.345 ;
        RECT 17.140 3.345 17.230 3.475 ;
        POLYGON 17.230 3.475 17.360 3.345 17.230 3.345 ;
        POLYGON 19.540 3.475 19.540 3.345 19.410 3.345 ;
        RECT 19.540 3.345 19.630 3.475 ;
        POLYGON 19.630 3.475 19.760 3.475 19.630 3.345 ;
        POLYGON 19.910 3.475 20.040 3.475 20.040 3.345 ;
        RECT 20.040 3.345 20.130 3.475 ;
        POLYGON 20.130 3.475 20.260 3.345 20.130 3.345 ;
        POLYGON 22.440 3.475 22.440 3.345 22.310 3.345 ;
        RECT 22.440 3.345 22.530 3.475 ;
        POLYGON 22.530 3.475 22.660 3.475 22.530 3.345 ;
        POLYGON 22.810 3.475 22.940 3.475 22.940 3.345 ;
        RECT 22.940 3.345 23.030 3.475 ;
        POLYGON 23.030 3.475 23.160 3.345 23.030 3.345 ;
        POLYGON 25.340 3.475 25.340 3.345 25.210 3.345 ;
        RECT 25.340 3.345 25.430 3.475 ;
        POLYGON 25.430 3.475 25.560 3.475 25.430 3.345 ;
        POLYGON 25.710 3.475 25.840 3.475 25.840 3.345 ;
        RECT 25.840 3.345 25.930 3.475 ;
        POLYGON 25.930 3.475 26.060 3.345 25.930 3.345 ;
        POLYGON 28.240 3.475 28.240 3.345 28.110 3.345 ;
        RECT 28.240 3.345 28.330 3.475 ;
        POLYGON 28.330 3.475 28.460 3.475 28.330 3.345 ;
        POLYGON 28.610 3.475 28.740 3.475 28.740 3.345 ;
        RECT 28.740 3.345 28.830 3.475 ;
        POLYGON 28.830 3.475 28.960 3.345 28.830 3.345 ;
        POLYGON 31.140 3.475 31.140 3.345 31.010 3.345 ;
        RECT 31.140 3.345 31.230 3.475 ;
        POLYGON 31.230 3.475 31.360 3.475 31.230 3.345 ;
        POLYGON 31.510 3.475 31.640 3.475 31.640 3.345 ;
        RECT 31.640 3.345 31.730 3.475 ;
        POLYGON 31.730 3.475 31.860 3.345 31.730 3.345 ;
        POLYGON 34.040 3.475 34.040 3.345 33.910 3.345 ;
        RECT 34.040 3.345 34.130 3.475 ;
        POLYGON 34.130 3.475 34.260 3.475 34.130 3.345 ;
        POLYGON 34.410 3.475 34.540 3.475 34.540 3.345 ;
        RECT 34.540 3.345 34.630 3.475 ;
        POLYGON 34.630 3.475 34.760 3.345 34.630 3.345 ;
        RECT -0.275 3.175 2.060 3.345 ;
        POLYGON 2.060 3.345 2.230 3.345 2.060 3.175 ;
        POLYGON 2.640 3.345 2.810 3.345 2.810 3.175 ;
        RECT 2.810 3.175 4.960 3.345 ;
        POLYGON 4.960 3.345 5.130 3.345 4.960 3.175 ;
        RECT 5.525 3.175 7.860 3.345 ;
        POLYGON 7.860 3.345 8.030 3.345 7.860 3.175 ;
        POLYGON 8.440 3.345 8.610 3.345 8.610 3.175 ;
        RECT 8.610 3.175 10.760 3.345 ;
        POLYGON 10.760 3.345 10.930 3.345 10.760 3.175 ;
        RECT 11.325 3.175 13.660 3.345 ;
        POLYGON 13.660 3.345 13.830 3.345 13.660 3.175 ;
        POLYGON 14.240 3.345 14.410 3.345 14.410 3.175 ;
        RECT 14.410 3.175 16.560 3.345 ;
        POLYGON 16.560 3.345 16.730 3.345 16.560 3.175 ;
        RECT 17.125 3.175 19.460 3.345 ;
        POLYGON 19.460 3.345 19.630 3.345 19.460 3.175 ;
        POLYGON 20.040 3.345 20.210 3.345 20.210 3.175 ;
        RECT 20.210 3.175 22.360 3.345 ;
        POLYGON 22.360 3.345 22.530 3.345 22.360 3.175 ;
        RECT 22.925 3.175 25.260 3.345 ;
        POLYGON 25.260 3.345 25.430 3.345 25.260 3.175 ;
        POLYGON 25.840 3.345 26.010 3.345 26.010 3.175 ;
        RECT 26.010 3.175 28.160 3.345 ;
        POLYGON 28.160 3.345 28.330 3.345 28.160 3.175 ;
        RECT 28.725 3.175 31.060 3.345 ;
        POLYGON 31.060 3.345 31.230 3.345 31.060 3.175 ;
        POLYGON 31.640 3.345 31.810 3.345 31.810 3.175 ;
        RECT 31.810 3.175 33.960 3.345 ;
        POLYGON 33.960 3.345 34.130 3.345 33.960 3.175 ;
        POLYGON 34.540 3.345 34.710 3.345 34.710 3.175 ;
        RECT 34.710 3.175 34.760 3.345 ;
    END
  END RWL1_2
  PIN RWL0_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 4.525 2.510 4.695 ;
        RECT 5.260 4.525 5.410 4.695 ;
        RECT 8.160 4.525 8.310 4.695 ;
        RECT 11.060 4.525 11.210 4.695 ;
        RECT 13.960 4.525 14.110 4.695 ;
        RECT 16.860 4.525 17.010 4.695 ;
        RECT 19.760 4.525 19.910 4.695 ;
        RECT 22.660 4.525 22.810 4.695 ;
        RECT 25.560 4.525 25.710 4.695 ;
        RECT 28.460 4.525 28.610 4.695 ;
        RECT 31.360 4.525 31.510 4.695 ;
        RECT 34.260 4.525 34.410 4.695 ;
      LAYER mcon ;
        RECT 2.360 4.530 2.510 4.695 ;
        RECT 8.160 4.530 8.310 4.695 ;
        RECT 13.960 4.530 14.110 4.695 ;
        RECT 19.760 4.530 19.910 4.695 ;
        RECT 25.560 4.530 25.710 4.695 ;
        RECT 31.360 4.530 31.510 4.695 ;
      LAYER met1 ;
        RECT 2.360 4.525 2.510 4.695 ;
        RECT 5.260 4.525 5.410 4.695 ;
        RECT 8.160 4.525 8.310 4.695 ;
        RECT 11.060 4.525 11.210 4.695 ;
        RECT 13.960 4.525 14.110 4.695 ;
        RECT 16.860 4.525 17.010 4.695 ;
        RECT 19.760 4.525 19.910 4.695 ;
        RECT 22.660 4.525 22.810 4.695 ;
        RECT 25.560 4.525 25.710 4.695 ;
        RECT 28.460 4.525 28.610 4.695 ;
        RECT 31.360 4.525 31.510 4.695 ;
        RECT 34.260 4.525 34.410 4.695 ;
      LAYER met2 ;
        RECT -0.275 4.525 34.760 4.695 ;
    END
  END RWL0_3
  PIN RWL1_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 4.525 0.330 4.695 ;
        RECT 3.080 4.525 3.230 4.695 ;
        RECT 5.980 4.525 6.130 4.695 ;
        RECT 8.880 4.525 9.030 4.695 ;
        RECT 11.780 4.525 11.930 4.695 ;
        RECT 14.680 4.525 14.830 4.695 ;
        RECT 17.580 4.525 17.730 4.695 ;
        RECT 20.480 4.525 20.630 4.695 ;
        RECT 23.380 4.525 23.530 4.695 ;
        RECT 26.280 4.525 26.430 4.695 ;
        RECT 29.180 4.525 29.330 4.695 ;
        RECT 32.080 4.525 32.230 4.695 ;
      LAYER met1 ;
        POLYGON 2.310 4.995 2.310 4.825 2.140 4.825 ;
        RECT 2.310 4.825 2.560 4.995 ;
        POLYGON 2.560 4.995 2.730 4.825 2.560 4.825 ;
        POLYGON 5.210 4.995 5.210 4.825 5.040 4.825 ;
        RECT 5.210 4.825 5.460 4.995 ;
        POLYGON 5.460 4.995 5.630 4.825 5.460 4.825 ;
        POLYGON 8.110 4.995 8.110 4.825 7.940 4.825 ;
        RECT 8.110 4.825 8.360 4.995 ;
        POLYGON 8.360 4.995 8.530 4.825 8.360 4.825 ;
        POLYGON 11.010 4.995 11.010 4.825 10.840 4.825 ;
        RECT 11.010 4.825 11.260 4.995 ;
        POLYGON 11.260 4.995 11.430 4.825 11.260 4.825 ;
        POLYGON 13.910 4.995 13.910 4.825 13.740 4.825 ;
        RECT 13.910 4.825 14.160 4.995 ;
        POLYGON 14.160 4.995 14.330 4.825 14.160 4.825 ;
        POLYGON 16.810 4.995 16.810 4.825 16.640 4.825 ;
        RECT 16.810 4.825 17.060 4.995 ;
        POLYGON 17.060 4.995 17.230 4.825 17.060 4.825 ;
        POLYGON 19.710 4.995 19.710 4.825 19.540 4.825 ;
        RECT 19.710 4.825 19.960 4.995 ;
        POLYGON 19.960 4.995 20.130 4.825 19.960 4.825 ;
        POLYGON 22.610 4.995 22.610 4.825 22.440 4.825 ;
        RECT 22.610 4.825 22.860 4.995 ;
        POLYGON 22.860 4.995 23.030 4.825 22.860 4.825 ;
        POLYGON 25.510 4.995 25.510 4.825 25.340 4.825 ;
        RECT 25.510 4.825 25.760 4.995 ;
        POLYGON 25.760 4.995 25.930 4.825 25.760 4.825 ;
        POLYGON 28.410 4.995 28.410 4.825 28.240 4.825 ;
        RECT 28.410 4.825 28.660 4.995 ;
        POLYGON 28.660 4.995 28.830 4.825 28.660 4.825 ;
        POLYGON 31.310 4.995 31.310 4.825 31.140 4.825 ;
        RECT 31.310 4.825 31.560 4.995 ;
        POLYGON 31.560 4.995 31.730 4.825 31.560 4.825 ;
        POLYGON 34.210 4.995 34.210 4.825 34.040 4.825 ;
        RECT 34.210 4.825 34.460 4.995 ;
        POLYGON 34.460 4.995 34.630 4.825 34.460 4.825 ;
        POLYGON 2.140 4.825 2.140 4.695 2.010 4.695 ;
        RECT 2.140 4.695 2.230 4.825 ;
        POLYGON 2.230 4.825 2.360 4.825 2.230 4.695 ;
        POLYGON 2.510 4.825 2.640 4.825 2.640 4.695 ;
        RECT 2.640 4.695 2.730 4.825 ;
        POLYGON 2.730 4.825 2.860 4.695 2.730 4.695 ;
        POLYGON 5.040 4.825 5.040 4.695 4.910 4.695 ;
        RECT 5.040 4.695 5.130 4.825 ;
        POLYGON 5.130 4.825 5.260 4.825 5.130 4.695 ;
        POLYGON 5.410 4.825 5.540 4.825 5.540 4.695 ;
        RECT 5.540 4.695 5.630 4.825 ;
        POLYGON 5.630 4.825 5.760 4.695 5.630 4.695 ;
        POLYGON 7.940 4.825 7.940 4.695 7.810 4.695 ;
        RECT 7.940 4.695 8.030 4.825 ;
        POLYGON 8.030 4.825 8.160 4.825 8.030 4.695 ;
        POLYGON 8.310 4.825 8.440 4.825 8.440 4.695 ;
        RECT 8.440 4.695 8.530 4.825 ;
        POLYGON 8.530 4.825 8.660 4.695 8.530 4.695 ;
        POLYGON 10.840 4.825 10.840 4.695 10.710 4.695 ;
        RECT 10.840 4.695 10.930 4.825 ;
        POLYGON 10.930 4.825 11.060 4.825 10.930 4.695 ;
        POLYGON 11.210 4.825 11.340 4.825 11.340 4.695 ;
        RECT 11.340 4.695 11.430 4.825 ;
        POLYGON 11.430 4.825 11.560 4.695 11.430 4.695 ;
        POLYGON 13.740 4.825 13.740 4.695 13.610 4.695 ;
        RECT 13.740 4.695 13.830 4.825 ;
        POLYGON 13.830 4.825 13.960 4.825 13.830 4.695 ;
        POLYGON 14.110 4.825 14.240 4.825 14.240 4.695 ;
        RECT 14.240 4.695 14.330 4.825 ;
        POLYGON 14.330 4.825 14.460 4.695 14.330 4.695 ;
        POLYGON 16.640 4.825 16.640 4.695 16.510 4.695 ;
        RECT 16.640 4.695 16.730 4.825 ;
        POLYGON 16.730 4.825 16.860 4.825 16.730 4.695 ;
        POLYGON 17.010 4.825 17.140 4.825 17.140 4.695 ;
        RECT 17.140 4.695 17.230 4.825 ;
        POLYGON 17.230 4.825 17.360 4.695 17.230 4.695 ;
        POLYGON 19.540 4.825 19.540 4.695 19.410 4.695 ;
        RECT 19.540 4.695 19.630 4.825 ;
        POLYGON 19.630 4.825 19.760 4.825 19.630 4.695 ;
        POLYGON 19.910 4.825 20.040 4.825 20.040 4.695 ;
        RECT 20.040 4.695 20.130 4.825 ;
        POLYGON 20.130 4.825 20.260 4.695 20.130 4.695 ;
        POLYGON 22.440 4.825 22.440 4.695 22.310 4.695 ;
        RECT 22.440 4.695 22.530 4.825 ;
        POLYGON 22.530 4.825 22.660 4.825 22.530 4.695 ;
        POLYGON 22.810 4.825 22.940 4.825 22.940 4.695 ;
        RECT 22.940 4.695 23.030 4.825 ;
        POLYGON 23.030 4.825 23.160 4.695 23.030 4.695 ;
        POLYGON 25.340 4.825 25.340 4.695 25.210 4.695 ;
        RECT 25.340 4.695 25.430 4.825 ;
        POLYGON 25.430 4.825 25.560 4.825 25.430 4.695 ;
        POLYGON 25.710 4.825 25.840 4.825 25.840 4.695 ;
        RECT 25.840 4.695 25.930 4.825 ;
        POLYGON 25.930 4.825 26.060 4.695 25.930 4.695 ;
        POLYGON 28.240 4.825 28.240 4.695 28.110 4.695 ;
        RECT 28.240 4.695 28.330 4.825 ;
        POLYGON 28.330 4.825 28.460 4.825 28.330 4.695 ;
        POLYGON 28.610 4.825 28.740 4.825 28.740 4.695 ;
        RECT 28.740 4.695 28.830 4.825 ;
        POLYGON 28.830 4.825 28.960 4.695 28.830 4.695 ;
        POLYGON 31.140 4.825 31.140 4.695 31.010 4.695 ;
        RECT 31.140 4.695 31.230 4.825 ;
        POLYGON 31.230 4.825 31.360 4.825 31.230 4.695 ;
        POLYGON 31.510 4.825 31.640 4.825 31.640 4.695 ;
        RECT 31.640 4.695 31.730 4.825 ;
        POLYGON 31.730 4.825 31.860 4.695 31.730 4.695 ;
        POLYGON 34.040 4.825 34.040 4.695 33.910 4.695 ;
        RECT 34.040 4.695 34.130 4.825 ;
        POLYGON 34.130 4.825 34.260 4.825 34.130 4.695 ;
        POLYGON 34.410 4.825 34.540 4.825 34.540 4.695 ;
        RECT 34.540 4.695 34.630 4.825 ;
        POLYGON 34.630 4.825 34.760 4.695 34.630 4.695 ;
        RECT -0.275 4.525 2.060 4.695 ;
        POLYGON 2.060 4.695 2.230 4.695 2.060 4.525 ;
        POLYGON 2.640 4.695 2.810 4.695 2.810 4.525 ;
        RECT 2.810 4.525 4.960 4.695 ;
        POLYGON 4.960 4.695 5.130 4.695 4.960 4.525 ;
        RECT 5.525 4.525 7.860 4.695 ;
        POLYGON 7.860 4.695 8.030 4.695 7.860 4.525 ;
        POLYGON 8.440 4.695 8.610 4.695 8.610 4.525 ;
        RECT 8.610 4.525 10.760 4.695 ;
        POLYGON 10.760 4.695 10.930 4.695 10.760 4.525 ;
        RECT 11.325 4.525 13.660 4.695 ;
        POLYGON 13.660 4.695 13.830 4.695 13.660 4.525 ;
        POLYGON 14.240 4.695 14.410 4.695 14.410 4.525 ;
        RECT 14.410 4.525 16.560 4.695 ;
        POLYGON 16.560 4.695 16.730 4.695 16.560 4.525 ;
        RECT 17.125 4.525 19.460 4.695 ;
        POLYGON 19.460 4.695 19.630 4.695 19.460 4.525 ;
        POLYGON 20.040 4.695 20.210 4.695 20.210 4.525 ;
        RECT 20.210 4.525 22.360 4.695 ;
        POLYGON 22.360 4.695 22.530 4.695 22.360 4.525 ;
        RECT 22.925 4.525 25.260 4.695 ;
        POLYGON 25.260 4.695 25.430 4.695 25.260 4.525 ;
        POLYGON 25.840 4.695 26.010 4.695 26.010 4.525 ;
        RECT 26.010 4.525 28.160 4.695 ;
        POLYGON 28.160 4.695 28.330 4.695 28.160 4.525 ;
        RECT 28.725 4.525 31.060 4.695 ;
        POLYGON 31.060 4.695 31.230 4.695 31.060 4.525 ;
        POLYGON 31.640 4.695 31.810 4.695 31.810 4.525 ;
        RECT 31.810 4.525 33.960 4.695 ;
        POLYGON 33.960 4.695 34.130 4.695 33.960 4.525 ;
        POLYGON 34.540 4.695 34.710 4.695 34.710 4.525 ;
        RECT 34.710 4.525 34.760 4.695 ;
    END
  END RWL1_3
  PIN RWL0_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 5.875 2.510 6.045 ;
        RECT 5.260 5.875 5.410 6.045 ;
        RECT 8.160 5.875 8.310 6.045 ;
        RECT 11.060 5.875 11.210 6.045 ;
        RECT 13.960 5.875 14.110 6.045 ;
        RECT 16.860 5.875 17.010 6.045 ;
        RECT 19.760 5.875 19.910 6.045 ;
        RECT 22.660 5.875 22.810 6.045 ;
        RECT 25.560 5.875 25.710 6.045 ;
        RECT 28.460 5.875 28.610 6.045 ;
        RECT 31.360 5.875 31.510 6.045 ;
        RECT 34.260 5.875 34.410 6.045 ;
      LAYER mcon ;
        RECT 2.360 5.880 2.510 6.045 ;
        RECT 8.160 5.880 8.310 6.045 ;
        RECT 13.960 5.880 14.110 6.045 ;
        RECT 19.760 5.880 19.910 6.045 ;
        RECT 25.560 5.880 25.710 6.045 ;
        RECT 31.360 5.880 31.510 6.045 ;
      LAYER met1 ;
        RECT 2.360 5.875 2.510 6.045 ;
        RECT 5.260 5.875 5.410 6.045 ;
        RECT 8.160 5.875 8.310 6.045 ;
        RECT 11.060 5.875 11.210 6.045 ;
        RECT 13.960 5.875 14.110 6.045 ;
        RECT 16.860 5.875 17.010 6.045 ;
        RECT 19.760 5.875 19.910 6.045 ;
        RECT 22.660 5.875 22.810 6.045 ;
        RECT 25.560 5.875 25.710 6.045 ;
        RECT 28.460 5.875 28.610 6.045 ;
        RECT 31.360 5.875 31.510 6.045 ;
        RECT 34.260 5.875 34.410 6.045 ;
      LAYER met2 ;
        RECT -0.275 5.875 34.760 6.045 ;
    END
  END RWL0_4
  PIN RWL1_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 5.875 0.330 6.045 ;
        RECT 3.080 5.875 3.230 6.045 ;
        RECT 5.980 5.875 6.130 6.045 ;
        RECT 8.880 5.875 9.030 6.045 ;
        RECT 11.780 5.875 11.930 6.045 ;
        RECT 14.680 5.875 14.830 6.045 ;
        RECT 17.580 5.875 17.730 6.045 ;
        RECT 20.480 5.875 20.630 6.045 ;
        RECT 23.380 5.875 23.530 6.045 ;
        RECT 26.280 5.875 26.430 6.045 ;
        RECT 29.180 5.875 29.330 6.045 ;
        RECT 32.080 5.875 32.230 6.045 ;
      LAYER met1 ;
        POLYGON 2.310 6.345 2.310 6.175 2.140 6.175 ;
        RECT 2.310 6.175 2.560 6.345 ;
        POLYGON 2.560 6.345 2.730 6.175 2.560 6.175 ;
        POLYGON 5.210 6.345 5.210 6.175 5.040 6.175 ;
        RECT 5.210 6.175 5.460 6.345 ;
        POLYGON 5.460 6.345 5.630 6.175 5.460 6.175 ;
        POLYGON 8.110 6.345 8.110 6.175 7.940 6.175 ;
        RECT 8.110 6.175 8.360 6.345 ;
        POLYGON 8.360 6.345 8.530 6.175 8.360 6.175 ;
        POLYGON 11.010 6.345 11.010 6.175 10.840 6.175 ;
        RECT 11.010 6.175 11.260 6.345 ;
        POLYGON 11.260 6.345 11.430 6.175 11.260 6.175 ;
        POLYGON 13.910 6.345 13.910 6.175 13.740 6.175 ;
        RECT 13.910 6.175 14.160 6.345 ;
        POLYGON 14.160 6.345 14.330 6.175 14.160 6.175 ;
        POLYGON 16.810 6.345 16.810 6.175 16.640 6.175 ;
        RECT 16.810 6.175 17.060 6.345 ;
        POLYGON 17.060 6.345 17.230 6.175 17.060 6.175 ;
        POLYGON 19.710 6.345 19.710 6.175 19.540 6.175 ;
        RECT 19.710 6.175 19.960 6.345 ;
        POLYGON 19.960 6.345 20.130 6.175 19.960 6.175 ;
        POLYGON 22.610 6.345 22.610 6.175 22.440 6.175 ;
        RECT 22.610 6.175 22.860 6.345 ;
        POLYGON 22.860 6.345 23.030 6.175 22.860 6.175 ;
        POLYGON 25.510 6.345 25.510 6.175 25.340 6.175 ;
        RECT 25.510 6.175 25.760 6.345 ;
        POLYGON 25.760 6.345 25.930 6.175 25.760 6.175 ;
        POLYGON 28.410 6.345 28.410 6.175 28.240 6.175 ;
        RECT 28.410 6.175 28.660 6.345 ;
        POLYGON 28.660 6.345 28.830 6.175 28.660 6.175 ;
        POLYGON 31.310 6.345 31.310 6.175 31.140 6.175 ;
        RECT 31.310 6.175 31.560 6.345 ;
        POLYGON 31.560 6.345 31.730 6.175 31.560 6.175 ;
        POLYGON 34.210 6.345 34.210 6.175 34.040 6.175 ;
        RECT 34.210 6.175 34.460 6.345 ;
        POLYGON 34.460 6.345 34.630 6.175 34.460 6.175 ;
        POLYGON 2.140 6.175 2.140 6.045 2.010 6.045 ;
        RECT 2.140 6.045 2.230 6.175 ;
        POLYGON 2.230 6.175 2.360 6.175 2.230 6.045 ;
        POLYGON 2.510 6.175 2.640 6.175 2.640 6.045 ;
        RECT 2.640 6.045 2.730 6.175 ;
        POLYGON 2.730 6.175 2.860 6.045 2.730 6.045 ;
        POLYGON 5.040 6.175 5.040 6.045 4.910 6.045 ;
        RECT 5.040 6.045 5.130 6.175 ;
        POLYGON 5.130 6.175 5.260 6.175 5.130 6.045 ;
        POLYGON 5.410 6.175 5.540 6.175 5.540 6.045 ;
        RECT 5.540 6.045 5.630 6.175 ;
        POLYGON 5.630 6.175 5.760 6.045 5.630 6.045 ;
        POLYGON 7.940 6.175 7.940 6.045 7.810 6.045 ;
        RECT 7.940 6.045 8.030 6.175 ;
        POLYGON 8.030 6.175 8.160 6.175 8.030 6.045 ;
        POLYGON 8.310 6.175 8.440 6.175 8.440 6.045 ;
        RECT 8.440 6.045 8.530 6.175 ;
        POLYGON 8.530 6.175 8.660 6.045 8.530 6.045 ;
        POLYGON 10.840 6.175 10.840 6.045 10.710 6.045 ;
        RECT 10.840 6.045 10.930 6.175 ;
        POLYGON 10.930 6.175 11.060 6.175 10.930 6.045 ;
        POLYGON 11.210 6.175 11.340 6.175 11.340 6.045 ;
        RECT 11.340 6.045 11.430 6.175 ;
        POLYGON 11.430 6.175 11.560 6.045 11.430 6.045 ;
        POLYGON 13.740 6.175 13.740 6.045 13.610 6.045 ;
        RECT 13.740 6.045 13.830 6.175 ;
        POLYGON 13.830 6.175 13.960 6.175 13.830 6.045 ;
        POLYGON 14.110 6.175 14.240 6.175 14.240 6.045 ;
        RECT 14.240 6.045 14.330 6.175 ;
        POLYGON 14.330 6.175 14.460 6.045 14.330 6.045 ;
        POLYGON 16.640 6.175 16.640 6.045 16.510 6.045 ;
        RECT 16.640 6.045 16.730 6.175 ;
        POLYGON 16.730 6.175 16.860 6.175 16.730 6.045 ;
        POLYGON 17.010 6.175 17.140 6.175 17.140 6.045 ;
        RECT 17.140 6.045 17.230 6.175 ;
        POLYGON 17.230 6.175 17.360 6.045 17.230 6.045 ;
        POLYGON 19.540 6.175 19.540 6.045 19.410 6.045 ;
        RECT 19.540 6.045 19.630 6.175 ;
        POLYGON 19.630 6.175 19.760 6.175 19.630 6.045 ;
        POLYGON 19.910 6.175 20.040 6.175 20.040 6.045 ;
        RECT 20.040 6.045 20.130 6.175 ;
        POLYGON 20.130 6.175 20.260 6.045 20.130 6.045 ;
        POLYGON 22.440 6.175 22.440 6.045 22.310 6.045 ;
        RECT 22.440 6.045 22.530 6.175 ;
        POLYGON 22.530 6.175 22.660 6.175 22.530 6.045 ;
        POLYGON 22.810 6.175 22.940 6.175 22.940 6.045 ;
        RECT 22.940 6.045 23.030 6.175 ;
        POLYGON 23.030 6.175 23.160 6.045 23.030 6.045 ;
        POLYGON 25.340 6.175 25.340 6.045 25.210 6.045 ;
        RECT 25.340 6.045 25.430 6.175 ;
        POLYGON 25.430 6.175 25.560 6.175 25.430 6.045 ;
        POLYGON 25.710 6.175 25.840 6.175 25.840 6.045 ;
        RECT 25.840 6.045 25.930 6.175 ;
        POLYGON 25.930 6.175 26.060 6.045 25.930 6.045 ;
        POLYGON 28.240 6.175 28.240 6.045 28.110 6.045 ;
        RECT 28.240 6.045 28.330 6.175 ;
        POLYGON 28.330 6.175 28.460 6.175 28.330 6.045 ;
        POLYGON 28.610 6.175 28.740 6.175 28.740 6.045 ;
        RECT 28.740 6.045 28.830 6.175 ;
        POLYGON 28.830 6.175 28.960 6.045 28.830 6.045 ;
        POLYGON 31.140 6.175 31.140 6.045 31.010 6.045 ;
        RECT 31.140 6.045 31.230 6.175 ;
        POLYGON 31.230 6.175 31.360 6.175 31.230 6.045 ;
        POLYGON 31.510 6.175 31.640 6.175 31.640 6.045 ;
        RECT 31.640 6.045 31.730 6.175 ;
        POLYGON 31.730 6.175 31.860 6.045 31.730 6.045 ;
        POLYGON 34.040 6.175 34.040 6.045 33.910 6.045 ;
        RECT 34.040 6.045 34.130 6.175 ;
        POLYGON 34.130 6.175 34.260 6.175 34.130 6.045 ;
        POLYGON 34.410 6.175 34.540 6.175 34.540 6.045 ;
        RECT 34.540 6.045 34.630 6.175 ;
        POLYGON 34.630 6.175 34.760 6.045 34.630 6.045 ;
        RECT -0.275 5.875 2.060 6.045 ;
        POLYGON 2.060 6.045 2.230 6.045 2.060 5.875 ;
        POLYGON 2.640 6.045 2.810 6.045 2.810 5.875 ;
        RECT 2.810 5.875 4.960 6.045 ;
        POLYGON 4.960 6.045 5.130 6.045 4.960 5.875 ;
        RECT 5.525 5.875 7.860 6.045 ;
        POLYGON 7.860 6.045 8.030 6.045 7.860 5.875 ;
        POLYGON 8.440 6.045 8.610 6.045 8.610 5.875 ;
        RECT 8.610 5.875 10.760 6.045 ;
        POLYGON 10.760 6.045 10.930 6.045 10.760 5.875 ;
        RECT 11.325 5.875 13.660 6.045 ;
        POLYGON 13.660 6.045 13.830 6.045 13.660 5.875 ;
        POLYGON 14.240 6.045 14.410 6.045 14.410 5.875 ;
        RECT 14.410 5.875 16.560 6.045 ;
        POLYGON 16.560 6.045 16.730 6.045 16.560 5.875 ;
        RECT 17.125 5.875 19.460 6.045 ;
        POLYGON 19.460 6.045 19.630 6.045 19.460 5.875 ;
        POLYGON 20.040 6.045 20.210 6.045 20.210 5.875 ;
        RECT 20.210 5.875 22.360 6.045 ;
        POLYGON 22.360 6.045 22.530 6.045 22.360 5.875 ;
        RECT 22.925 5.875 25.260 6.045 ;
        POLYGON 25.260 6.045 25.430 6.045 25.260 5.875 ;
        POLYGON 25.840 6.045 26.010 6.045 26.010 5.875 ;
        RECT 26.010 5.875 28.160 6.045 ;
        POLYGON 28.160 6.045 28.330 6.045 28.160 5.875 ;
        RECT 28.725 5.875 31.060 6.045 ;
        POLYGON 31.060 6.045 31.230 6.045 31.060 5.875 ;
        POLYGON 31.640 6.045 31.810 6.045 31.810 5.875 ;
        RECT 31.810 5.875 33.960 6.045 ;
        POLYGON 33.960 6.045 34.130 6.045 33.960 5.875 ;
        POLYGON 34.540 6.045 34.710 6.045 34.710 5.875 ;
        RECT 34.710 5.875 34.760 6.045 ;
    END
  END RWL1_4
  PIN RWL0_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 7.225 2.510 7.395 ;
        RECT 5.260 7.225 5.410 7.395 ;
        RECT 8.160 7.225 8.310 7.395 ;
        RECT 11.060 7.225 11.210 7.395 ;
        RECT 13.960 7.225 14.110 7.395 ;
        RECT 16.860 7.225 17.010 7.395 ;
        RECT 19.760 7.225 19.910 7.395 ;
        RECT 22.660 7.225 22.810 7.395 ;
        RECT 25.560 7.225 25.710 7.395 ;
        RECT 28.460 7.225 28.610 7.395 ;
        RECT 31.360 7.225 31.510 7.395 ;
        RECT 34.260 7.225 34.410 7.395 ;
      LAYER mcon ;
        RECT 2.360 7.230 2.510 7.395 ;
        RECT 8.160 7.230 8.310 7.395 ;
        RECT 13.960 7.230 14.110 7.395 ;
        RECT 19.760 7.230 19.910 7.395 ;
        RECT 25.560 7.230 25.710 7.395 ;
        RECT 31.360 7.230 31.510 7.395 ;
      LAYER met1 ;
        RECT 2.360 7.225 2.510 7.395 ;
        RECT 5.260 7.225 5.410 7.395 ;
        RECT 8.160 7.225 8.310 7.395 ;
        RECT 11.060 7.225 11.210 7.395 ;
        RECT 13.960 7.225 14.110 7.395 ;
        RECT 16.860 7.225 17.010 7.395 ;
        RECT 19.760 7.225 19.910 7.395 ;
        RECT 22.660 7.225 22.810 7.395 ;
        RECT 25.560 7.225 25.710 7.395 ;
        RECT 28.460 7.225 28.610 7.395 ;
        RECT 31.360 7.225 31.510 7.395 ;
        RECT 34.260 7.225 34.410 7.395 ;
      LAYER met2 ;
        RECT -0.275 7.225 34.760 7.395 ;
    END
  END RWL0_5
  PIN RWL1_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 7.225 0.330 7.395 ;
        RECT 3.080 7.225 3.230 7.395 ;
        RECT 5.980 7.225 6.130 7.395 ;
        RECT 8.880 7.225 9.030 7.395 ;
        RECT 11.780 7.225 11.930 7.395 ;
        RECT 14.680 7.225 14.830 7.395 ;
        RECT 17.580 7.225 17.730 7.395 ;
        RECT 20.480 7.225 20.630 7.395 ;
        RECT 23.380 7.225 23.530 7.395 ;
        RECT 26.280 7.225 26.430 7.395 ;
        RECT 29.180 7.225 29.330 7.395 ;
        RECT 32.080 7.225 32.230 7.395 ;
      LAYER met1 ;
        POLYGON 2.310 7.695 2.310 7.525 2.140 7.525 ;
        RECT 2.310 7.525 2.560 7.695 ;
        POLYGON 2.560 7.695 2.730 7.525 2.560 7.525 ;
        POLYGON 5.210 7.695 5.210 7.525 5.040 7.525 ;
        RECT 5.210 7.525 5.460 7.695 ;
        POLYGON 5.460 7.695 5.630 7.525 5.460 7.525 ;
        POLYGON 8.110 7.695 8.110 7.525 7.940 7.525 ;
        RECT 8.110 7.525 8.360 7.695 ;
        POLYGON 8.360 7.695 8.530 7.525 8.360 7.525 ;
        POLYGON 11.010 7.695 11.010 7.525 10.840 7.525 ;
        RECT 11.010 7.525 11.260 7.695 ;
        POLYGON 11.260 7.695 11.430 7.525 11.260 7.525 ;
        POLYGON 13.910 7.695 13.910 7.525 13.740 7.525 ;
        RECT 13.910 7.525 14.160 7.695 ;
        POLYGON 14.160 7.695 14.330 7.525 14.160 7.525 ;
        POLYGON 16.810 7.695 16.810 7.525 16.640 7.525 ;
        RECT 16.810 7.525 17.060 7.695 ;
        POLYGON 17.060 7.695 17.230 7.525 17.060 7.525 ;
        POLYGON 19.710 7.695 19.710 7.525 19.540 7.525 ;
        RECT 19.710 7.525 19.960 7.695 ;
        POLYGON 19.960 7.695 20.130 7.525 19.960 7.525 ;
        POLYGON 22.610 7.695 22.610 7.525 22.440 7.525 ;
        RECT 22.610 7.525 22.860 7.695 ;
        POLYGON 22.860 7.695 23.030 7.525 22.860 7.525 ;
        POLYGON 25.510 7.695 25.510 7.525 25.340 7.525 ;
        RECT 25.510 7.525 25.760 7.695 ;
        POLYGON 25.760 7.695 25.930 7.525 25.760 7.525 ;
        POLYGON 28.410 7.695 28.410 7.525 28.240 7.525 ;
        RECT 28.410 7.525 28.660 7.695 ;
        POLYGON 28.660 7.695 28.830 7.525 28.660 7.525 ;
        POLYGON 31.310 7.695 31.310 7.525 31.140 7.525 ;
        RECT 31.310 7.525 31.560 7.695 ;
        POLYGON 31.560 7.695 31.730 7.525 31.560 7.525 ;
        POLYGON 34.210 7.695 34.210 7.525 34.040 7.525 ;
        RECT 34.210 7.525 34.460 7.695 ;
        POLYGON 34.460 7.695 34.630 7.525 34.460 7.525 ;
        POLYGON 2.140 7.525 2.140 7.395 2.010 7.395 ;
        RECT 2.140 7.395 2.230 7.525 ;
        POLYGON 2.230 7.525 2.360 7.525 2.230 7.395 ;
        POLYGON 2.510 7.525 2.640 7.525 2.640 7.395 ;
        RECT 2.640 7.395 2.730 7.525 ;
        POLYGON 2.730 7.525 2.860 7.395 2.730 7.395 ;
        POLYGON 5.040 7.525 5.040 7.395 4.910 7.395 ;
        RECT 5.040 7.395 5.130 7.525 ;
        POLYGON 5.130 7.525 5.260 7.525 5.130 7.395 ;
        POLYGON 5.410 7.525 5.540 7.525 5.540 7.395 ;
        RECT 5.540 7.395 5.630 7.525 ;
        POLYGON 5.630 7.525 5.760 7.395 5.630 7.395 ;
        POLYGON 7.940 7.525 7.940 7.395 7.810 7.395 ;
        RECT 7.940 7.395 8.030 7.525 ;
        POLYGON 8.030 7.525 8.160 7.525 8.030 7.395 ;
        POLYGON 8.310 7.525 8.440 7.525 8.440 7.395 ;
        RECT 8.440 7.395 8.530 7.525 ;
        POLYGON 8.530 7.525 8.660 7.395 8.530 7.395 ;
        POLYGON 10.840 7.525 10.840 7.395 10.710 7.395 ;
        RECT 10.840 7.395 10.930 7.525 ;
        POLYGON 10.930 7.525 11.060 7.525 10.930 7.395 ;
        POLYGON 11.210 7.525 11.340 7.525 11.340 7.395 ;
        RECT 11.340 7.395 11.430 7.525 ;
        POLYGON 11.430 7.525 11.560 7.395 11.430 7.395 ;
        POLYGON 13.740 7.525 13.740 7.395 13.610 7.395 ;
        RECT 13.740 7.395 13.830 7.525 ;
        POLYGON 13.830 7.525 13.960 7.525 13.830 7.395 ;
        POLYGON 14.110 7.525 14.240 7.525 14.240 7.395 ;
        RECT 14.240 7.395 14.330 7.525 ;
        POLYGON 14.330 7.525 14.460 7.395 14.330 7.395 ;
        POLYGON 16.640 7.525 16.640 7.395 16.510 7.395 ;
        RECT 16.640 7.395 16.730 7.525 ;
        POLYGON 16.730 7.525 16.860 7.525 16.730 7.395 ;
        POLYGON 17.010 7.525 17.140 7.525 17.140 7.395 ;
        RECT 17.140 7.395 17.230 7.525 ;
        POLYGON 17.230 7.525 17.360 7.395 17.230 7.395 ;
        POLYGON 19.540 7.525 19.540 7.395 19.410 7.395 ;
        RECT 19.540 7.395 19.630 7.525 ;
        POLYGON 19.630 7.525 19.760 7.525 19.630 7.395 ;
        POLYGON 19.910 7.525 20.040 7.525 20.040 7.395 ;
        RECT 20.040 7.395 20.130 7.525 ;
        POLYGON 20.130 7.525 20.260 7.395 20.130 7.395 ;
        POLYGON 22.440 7.525 22.440 7.395 22.310 7.395 ;
        RECT 22.440 7.395 22.530 7.525 ;
        POLYGON 22.530 7.525 22.660 7.525 22.530 7.395 ;
        POLYGON 22.810 7.525 22.940 7.525 22.940 7.395 ;
        RECT 22.940 7.395 23.030 7.525 ;
        POLYGON 23.030 7.525 23.160 7.395 23.030 7.395 ;
        POLYGON 25.340 7.525 25.340 7.395 25.210 7.395 ;
        RECT 25.340 7.395 25.430 7.525 ;
        POLYGON 25.430 7.525 25.560 7.525 25.430 7.395 ;
        POLYGON 25.710 7.525 25.840 7.525 25.840 7.395 ;
        RECT 25.840 7.395 25.930 7.525 ;
        POLYGON 25.930 7.525 26.060 7.395 25.930 7.395 ;
        POLYGON 28.240 7.525 28.240 7.395 28.110 7.395 ;
        RECT 28.240 7.395 28.330 7.525 ;
        POLYGON 28.330 7.525 28.460 7.525 28.330 7.395 ;
        POLYGON 28.610 7.525 28.740 7.525 28.740 7.395 ;
        RECT 28.740 7.395 28.830 7.525 ;
        POLYGON 28.830 7.525 28.960 7.395 28.830 7.395 ;
        POLYGON 31.140 7.525 31.140 7.395 31.010 7.395 ;
        RECT 31.140 7.395 31.230 7.525 ;
        POLYGON 31.230 7.525 31.360 7.525 31.230 7.395 ;
        POLYGON 31.510 7.525 31.640 7.525 31.640 7.395 ;
        RECT 31.640 7.395 31.730 7.525 ;
        POLYGON 31.730 7.525 31.860 7.395 31.730 7.395 ;
        POLYGON 34.040 7.525 34.040 7.395 33.910 7.395 ;
        RECT 34.040 7.395 34.130 7.525 ;
        POLYGON 34.130 7.525 34.260 7.525 34.130 7.395 ;
        POLYGON 34.410 7.525 34.540 7.525 34.540 7.395 ;
        RECT 34.540 7.395 34.630 7.525 ;
        POLYGON 34.630 7.525 34.760 7.395 34.630 7.395 ;
        RECT -0.275 7.225 2.060 7.395 ;
        POLYGON 2.060 7.395 2.230 7.395 2.060 7.225 ;
        POLYGON 2.640 7.395 2.810 7.395 2.810 7.225 ;
        RECT 2.810 7.225 4.960 7.395 ;
        POLYGON 4.960 7.395 5.130 7.395 4.960 7.225 ;
        RECT 5.525 7.225 7.860 7.395 ;
        POLYGON 7.860 7.395 8.030 7.395 7.860 7.225 ;
        POLYGON 8.440 7.395 8.610 7.395 8.610 7.225 ;
        RECT 8.610 7.225 10.760 7.395 ;
        POLYGON 10.760 7.395 10.930 7.395 10.760 7.225 ;
        RECT 11.325 7.225 13.660 7.395 ;
        POLYGON 13.660 7.395 13.830 7.395 13.660 7.225 ;
        POLYGON 14.240 7.395 14.410 7.395 14.410 7.225 ;
        RECT 14.410 7.225 16.560 7.395 ;
        POLYGON 16.560 7.395 16.730 7.395 16.560 7.225 ;
        RECT 17.125 7.225 19.460 7.395 ;
        POLYGON 19.460 7.395 19.630 7.395 19.460 7.225 ;
        POLYGON 20.040 7.395 20.210 7.395 20.210 7.225 ;
        RECT 20.210 7.225 22.360 7.395 ;
        POLYGON 22.360 7.395 22.530 7.395 22.360 7.225 ;
        RECT 22.925 7.225 25.260 7.395 ;
        POLYGON 25.260 7.395 25.430 7.395 25.260 7.225 ;
        POLYGON 25.840 7.395 26.010 7.395 26.010 7.225 ;
        RECT 26.010 7.225 28.160 7.395 ;
        POLYGON 28.160 7.395 28.330 7.395 28.160 7.225 ;
        RECT 28.725 7.225 31.060 7.395 ;
        POLYGON 31.060 7.395 31.230 7.395 31.060 7.225 ;
        POLYGON 31.640 7.395 31.810 7.395 31.810 7.225 ;
        RECT 31.810 7.225 33.960 7.395 ;
        POLYGON 33.960 7.395 34.130 7.395 33.960 7.225 ;
        POLYGON 34.540 7.395 34.710 7.395 34.710 7.225 ;
        RECT 34.710 7.225 34.760 7.395 ;
    END
  END RWL1_5
  PIN RWL0_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 8.575 2.510 8.745 ;
        RECT 5.260 8.575 5.410 8.745 ;
        RECT 8.160 8.575 8.310 8.745 ;
        RECT 11.060 8.575 11.210 8.745 ;
        RECT 13.960 8.575 14.110 8.745 ;
        RECT 16.860 8.575 17.010 8.745 ;
        RECT 19.760 8.575 19.910 8.745 ;
        RECT 22.660 8.575 22.810 8.745 ;
        RECT 25.560 8.575 25.710 8.745 ;
        RECT 28.460 8.575 28.610 8.745 ;
        RECT 31.360 8.575 31.510 8.745 ;
        RECT 34.260 8.575 34.410 8.745 ;
      LAYER mcon ;
        RECT 2.360 8.580 2.510 8.745 ;
        RECT 8.160 8.580 8.310 8.745 ;
        RECT 13.960 8.580 14.110 8.745 ;
        RECT 19.760 8.580 19.910 8.745 ;
        RECT 25.560 8.580 25.710 8.745 ;
        RECT 31.360 8.580 31.510 8.745 ;
      LAYER met1 ;
        RECT 2.360 8.575 2.510 8.745 ;
        RECT 5.260 8.575 5.410 8.745 ;
        RECT 8.160 8.575 8.310 8.745 ;
        RECT 11.060 8.575 11.210 8.745 ;
        RECT 13.960 8.575 14.110 8.745 ;
        RECT 16.860 8.575 17.010 8.745 ;
        RECT 19.760 8.575 19.910 8.745 ;
        RECT 22.660 8.575 22.810 8.745 ;
        RECT 25.560 8.575 25.710 8.745 ;
        RECT 28.460 8.575 28.610 8.745 ;
        RECT 31.360 8.575 31.510 8.745 ;
        RECT 34.260 8.575 34.410 8.745 ;
      LAYER met2 ;
        RECT -0.275 8.575 34.760 8.745 ;
    END
  END RWL0_6
  PIN RWL1_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 8.575 0.330 8.745 ;
        RECT 3.080 8.575 3.230 8.745 ;
        RECT 5.980 8.575 6.130 8.745 ;
        RECT 8.880 8.575 9.030 8.745 ;
        RECT 11.780 8.575 11.930 8.745 ;
        RECT 14.680 8.575 14.830 8.745 ;
        RECT 17.580 8.575 17.730 8.745 ;
        RECT 20.480 8.575 20.630 8.745 ;
        RECT 23.380 8.575 23.530 8.745 ;
        RECT 26.280 8.575 26.430 8.745 ;
        RECT 29.180 8.575 29.330 8.745 ;
        RECT 32.080 8.575 32.230 8.745 ;
      LAYER met1 ;
        POLYGON 2.310 9.045 2.310 8.875 2.140 8.875 ;
        RECT 2.310 8.875 2.560 9.045 ;
        POLYGON 2.560 9.045 2.730 8.875 2.560 8.875 ;
        POLYGON 5.210 9.045 5.210 8.875 5.040 8.875 ;
        RECT 5.210 8.875 5.460 9.045 ;
        POLYGON 5.460 9.045 5.630 8.875 5.460 8.875 ;
        POLYGON 8.110 9.045 8.110 8.875 7.940 8.875 ;
        RECT 8.110 8.875 8.360 9.045 ;
        POLYGON 8.360 9.045 8.530 8.875 8.360 8.875 ;
        POLYGON 11.010 9.045 11.010 8.875 10.840 8.875 ;
        RECT 11.010 8.875 11.260 9.045 ;
        POLYGON 11.260 9.045 11.430 8.875 11.260 8.875 ;
        POLYGON 13.910 9.045 13.910 8.875 13.740 8.875 ;
        RECT 13.910 8.875 14.160 9.045 ;
        POLYGON 14.160 9.045 14.330 8.875 14.160 8.875 ;
        POLYGON 16.810 9.045 16.810 8.875 16.640 8.875 ;
        RECT 16.810 8.875 17.060 9.045 ;
        POLYGON 17.060 9.045 17.230 8.875 17.060 8.875 ;
        POLYGON 19.710 9.045 19.710 8.875 19.540 8.875 ;
        RECT 19.710 8.875 19.960 9.045 ;
        POLYGON 19.960 9.045 20.130 8.875 19.960 8.875 ;
        POLYGON 22.610 9.045 22.610 8.875 22.440 8.875 ;
        RECT 22.610 8.875 22.860 9.045 ;
        POLYGON 22.860 9.045 23.030 8.875 22.860 8.875 ;
        POLYGON 25.510 9.045 25.510 8.875 25.340 8.875 ;
        RECT 25.510 8.875 25.760 9.045 ;
        POLYGON 25.760 9.045 25.930 8.875 25.760 8.875 ;
        POLYGON 28.410 9.045 28.410 8.875 28.240 8.875 ;
        RECT 28.410 8.875 28.660 9.045 ;
        POLYGON 28.660 9.045 28.830 8.875 28.660 8.875 ;
        POLYGON 31.310 9.045 31.310 8.875 31.140 8.875 ;
        RECT 31.310 8.875 31.560 9.045 ;
        POLYGON 31.560 9.045 31.730 8.875 31.560 8.875 ;
        POLYGON 34.210 9.045 34.210 8.875 34.040 8.875 ;
        RECT 34.210 8.875 34.460 9.045 ;
        POLYGON 34.460 9.045 34.630 8.875 34.460 8.875 ;
        POLYGON 2.140 8.875 2.140 8.745 2.010 8.745 ;
        RECT 2.140 8.745 2.230 8.875 ;
        POLYGON 2.230 8.875 2.360 8.875 2.230 8.745 ;
        POLYGON 2.510 8.875 2.640 8.875 2.640 8.745 ;
        RECT 2.640 8.745 2.730 8.875 ;
        POLYGON 2.730 8.875 2.860 8.745 2.730 8.745 ;
        POLYGON 5.040 8.875 5.040 8.745 4.910 8.745 ;
        RECT 5.040 8.745 5.130 8.875 ;
        POLYGON 5.130 8.875 5.260 8.875 5.130 8.745 ;
        POLYGON 5.410 8.875 5.540 8.875 5.540 8.745 ;
        RECT 5.540 8.745 5.630 8.875 ;
        POLYGON 5.630 8.875 5.760 8.745 5.630 8.745 ;
        POLYGON 7.940 8.875 7.940 8.745 7.810 8.745 ;
        RECT 7.940 8.745 8.030 8.875 ;
        POLYGON 8.030 8.875 8.160 8.875 8.030 8.745 ;
        POLYGON 8.310 8.875 8.440 8.875 8.440 8.745 ;
        RECT 8.440 8.745 8.530 8.875 ;
        POLYGON 8.530 8.875 8.660 8.745 8.530 8.745 ;
        POLYGON 10.840 8.875 10.840 8.745 10.710 8.745 ;
        RECT 10.840 8.745 10.930 8.875 ;
        POLYGON 10.930 8.875 11.060 8.875 10.930 8.745 ;
        POLYGON 11.210 8.875 11.340 8.875 11.340 8.745 ;
        RECT 11.340 8.745 11.430 8.875 ;
        POLYGON 11.430 8.875 11.560 8.745 11.430 8.745 ;
        POLYGON 13.740 8.875 13.740 8.745 13.610 8.745 ;
        RECT 13.740 8.745 13.830 8.875 ;
        POLYGON 13.830 8.875 13.960 8.875 13.830 8.745 ;
        POLYGON 14.110 8.875 14.240 8.875 14.240 8.745 ;
        RECT 14.240 8.745 14.330 8.875 ;
        POLYGON 14.330 8.875 14.460 8.745 14.330 8.745 ;
        POLYGON 16.640 8.875 16.640 8.745 16.510 8.745 ;
        RECT 16.640 8.745 16.730 8.875 ;
        POLYGON 16.730 8.875 16.860 8.875 16.730 8.745 ;
        POLYGON 17.010 8.875 17.140 8.875 17.140 8.745 ;
        RECT 17.140 8.745 17.230 8.875 ;
        POLYGON 17.230 8.875 17.360 8.745 17.230 8.745 ;
        POLYGON 19.540 8.875 19.540 8.745 19.410 8.745 ;
        RECT 19.540 8.745 19.630 8.875 ;
        POLYGON 19.630 8.875 19.760 8.875 19.630 8.745 ;
        POLYGON 19.910 8.875 20.040 8.875 20.040 8.745 ;
        RECT 20.040 8.745 20.130 8.875 ;
        POLYGON 20.130 8.875 20.260 8.745 20.130 8.745 ;
        POLYGON 22.440 8.875 22.440 8.745 22.310 8.745 ;
        RECT 22.440 8.745 22.530 8.875 ;
        POLYGON 22.530 8.875 22.660 8.875 22.530 8.745 ;
        POLYGON 22.810 8.875 22.940 8.875 22.940 8.745 ;
        RECT 22.940 8.745 23.030 8.875 ;
        POLYGON 23.030 8.875 23.160 8.745 23.030 8.745 ;
        POLYGON 25.340 8.875 25.340 8.745 25.210 8.745 ;
        RECT 25.340 8.745 25.430 8.875 ;
        POLYGON 25.430 8.875 25.560 8.875 25.430 8.745 ;
        POLYGON 25.710 8.875 25.840 8.875 25.840 8.745 ;
        RECT 25.840 8.745 25.930 8.875 ;
        POLYGON 25.930 8.875 26.060 8.745 25.930 8.745 ;
        POLYGON 28.240 8.875 28.240 8.745 28.110 8.745 ;
        RECT 28.240 8.745 28.330 8.875 ;
        POLYGON 28.330 8.875 28.460 8.875 28.330 8.745 ;
        POLYGON 28.610 8.875 28.740 8.875 28.740 8.745 ;
        RECT 28.740 8.745 28.830 8.875 ;
        POLYGON 28.830 8.875 28.960 8.745 28.830 8.745 ;
        POLYGON 31.140 8.875 31.140 8.745 31.010 8.745 ;
        RECT 31.140 8.745 31.230 8.875 ;
        POLYGON 31.230 8.875 31.360 8.875 31.230 8.745 ;
        POLYGON 31.510 8.875 31.640 8.875 31.640 8.745 ;
        RECT 31.640 8.745 31.730 8.875 ;
        POLYGON 31.730 8.875 31.860 8.745 31.730 8.745 ;
        POLYGON 34.040 8.875 34.040 8.745 33.910 8.745 ;
        RECT 34.040 8.745 34.130 8.875 ;
        POLYGON 34.130 8.875 34.260 8.875 34.130 8.745 ;
        POLYGON 34.410 8.875 34.540 8.875 34.540 8.745 ;
        RECT 34.540 8.745 34.630 8.875 ;
        POLYGON 34.630 8.875 34.760 8.745 34.630 8.745 ;
        RECT -0.275 8.575 2.060 8.745 ;
        POLYGON 2.060 8.745 2.230 8.745 2.060 8.575 ;
        POLYGON 2.640 8.745 2.810 8.745 2.810 8.575 ;
        RECT 2.810 8.575 4.960 8.745 ;
        POLYGON 4.960 8.745 5.130 8.745 4.960 8.575 ;
        RECT 5.525 8.575 7.860 8.745 ;
        POLYGON 7.860 8.745 8.030 8.745 7.860 8.575 ;
        POLYGON 8.440 8.745 8.610 8.745 8.610 8.575 ;
        RECT 8.610 8.575 10.760 8.745 ;
        POLYGON 10.760 8.745 10.930 8.745 10.760 8.575 ;
        RECT 11.325 8.575 13.660 8.745 ;
        POLYGON 13.660 8.745 13.830 8.745 13.660 8.575 ;
        POLYGON 14.240 8.745 14.410 8.745 14.410 8.575 ;
        RECT 14.410 8.575 16.560 8.745 ;
        POLYGON 16.560 8.745 16.730 8.745 16.560 8.575 ;
        RECT 17.125 8.575 19.460 8.745 ;
        POLYGON 19.460 8.745 19.630 8.745 19.460 8.575 ;
        POLYGON 20.040 8.745 20.210 8.745 20.210 8.575 ;
        RECT 20.210 8.575 22.360 8.745 ;
        POLYGON 22.360 8.745 22.530 8.745 22.360 8.575 ;
        RECT 22.925 8.575 25.260 8.745 ;
        POLYGON 25.260 8.745 25.430 8.745 25.260 8.575 ;
        POLYGON 25.840 8.745 26.010 8.745 26.010 8.575 ;
        RECT 26.010 8.575 28.160 8.745 ;
        POLYGON 28.160 8.745 28.330 8.745 28.160 8.575 ;
        RECT 28.725 8.575 31.060 8.745 ;
        POLYGON 31.060 8.745 31.230 8.745 31.060 8.575 ;
        POLYGON 31.640 8.745 31.810 8.745 31.810 8.575 ;
        RECT 31.810 8.575 33.960 8.745 ;
        POLYGON 33.960 8.745 34.130 8.745 33.960 8.575 ;
        POLYGON 34.540 8.745 34.710 8.745 34.710 8.575 ;
        RECT 34.710 8.575 34.760 8.745 ;
    END
  END RWL1_6
  PIN RWL0_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 9.925 2.510 10.095 ;
        RECT 5.260 9.925 5.410 10.095 ;
        RECT 8.160 9.925 8.310 10.095 ;
        RECT 11.060 9.925 11.210 10.095 ;
        RECT 13.960 9.925 14.110 10.095 ;
        RECT 16.860 9.925 17.010 10.095 ;
        RECT 19.760 9.925 19.910 10.095 ;
        RECT 22.660 9.925 22.810 10.095 ;
        RECT 25.560 9.925 25.710 10.095 ;
        RECT 28.460 9.925 28.610 10.095 ;
        RECT 31.360 9.925 31.510 10.095 ;
        RECT 34.260 9.925 34.410 10.095 ;
      LAYER mcon ;
        RECT 2.360 9.930 2.510 10.095 ;
        RECT 8.160 9.930 8.310 10.095 ;
        RECT 13.960 9.930 14.110 10.095 ;
        RECT 19.760 9.930 19.910 10.095 ;
        RECT 25.560 9.930 25.710 10.095 ;
        RECT 31.360 9.930 31.510 10.095 ;
      LAYER met1 ;
        RECT 2.360 9.925 2.510 10.095 ;
        RECT 5.260 9.925 5.410 10.095 ;
        RECT 8.160 9.925 8.310 10.095 ;
        RECT 11.060 9.925 11.210 10.095 ;
        RECT 13.960 9.925 14.110 10.095 ;
        RECT 16.860 9.925 17.010 10.095 ;
        RECT 19.760 9.925 19.910 10.095 ;
        RECT 22.660 9.925 22.810 10.095 ;
        RECT 25.560 9.925 25.710 10.095 ;
        RECT 28.460 9.925 28.610 10.095 ;
        RECT 31.360 9.925 31.510 10.095 ;
        RECT 34.260 9.925 34.410 10.095 ;
      LAYER met2 ;
        RECT -0.275 9.925 34.760 10.095 ;
    END
  END RWL0_7
  PIN RWL1_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 9.925 0.330 10.095 ;
        RECT 3.080 9.925 3.230 10.095 ;
        RECT 5.980 9.925 6.130 10.095 ;
        RECT 8.880 9.925 9.030 10.095 ;
        RECT 11.780 9.925 11.930 10.095 ;
        RECT 14.680 9.925 14.830 10.095 ;
        RECT 17.580 9.925 17.730 10.095 ;
        RECT 20.480 9.925 20.630 10.095 ;
        RECT 23.380 9.925 23.530 10.095 ;
        RECT 26.280 9.925 26.430 10.095 ;
        RECT 29.180 9.925 29.330 10.095 ;
        RECT 32.080 9.925 32.230 10.095 ;
      LAYER met1 ;
        POLYGON 2.310 10.395 2.310 10.225 2.140 10.225 ;
        RECT 2.310 10.225 2.560 10.395 ;
        POLYGON 2.560 10.395 2.730 10.225 2.560 10.225 ;
        POLYGON 5.210 10.395 5.210 10.225 5.040 10.225 ;
        RECT 5.210 10.225 5.460 10.395 ;
        POLYGON 5.460 10.395 5.630 10.225 5.460 10.225 ;
        POLYGON 8.110 10.395 8.110 10.225 7.940 10.225 ;
        RECT 8.110 10.225 8.360 10.395 ;
        POLYGON 8.360 10.395 8.530 10.225 8.360 10.225 ;
        POLYGON 11.010 10.395 11.010 10.225 10.840 10.225 ;
        RECT 11.010 10.225 11.260 10.395 ;
        POLYGON 11.260 10.395 11.430 10.225 11.260 10.225 ;
        POLYGON 13.910 10.395 13.910 10.225 13.740 10.225 ;
        RECT 13.910 10.225 14.160 10.395 ;
        POLYGON 14.160 10.395 14.330 10.225 14.160 10.225 ;
        POLYGON 16.810 10.395 16.810 10.225 16.640 10.225 ;
        RECT 16.810 10.225 17.060 10.395 ;
        POLYGON 17.060 10.395 17.230 10.225 17.060 10.225 ;
        POLYGON 19.710 10.395 19.710 10.225 19.540 10.225 ;
        RECT 19.710 10.225 19.960 10.395 ;
        POLYGON 19.960 10.395 20.130 10.225 19.960 10.225 ;
        POLYGON 22.610 10.395 22.610 10.225 22.440 10.225 ;
        RECT 22.610 10.225 22.860 10.395 ;
        POLYGON 22.860 10.395 23.030 10.225 22.860 10.225 ;
        POLYGON 25.510 10.395 25.510 10.225 25.340 10.225 ;
        RECT 25.510 10.225 25.760 10.395 ;
        POLYGON 25.760 10.395 25.930 10.225 25.760 10.225 ;
        POLYGON 28.410 10.395 28.410 10.225 28.240 10.225 ;
        RECT 28.410 10.225 28.660 10.395 ;
        POLYGON 28.660 10.395 28.830 10.225 28.660 10.225 ;
        POLYGON 31.310 10.395 31.310 10.225 31.140 10.225 ;
        RECT 31.310 10.225 31.560 10.395 ;
        POLYGON 31.560 10.395 31.730 10.225 31.560 10.225 ;
        POLYGON 34.210 10.395 34.210 10.225 34.040 10.225 ;
        RECT 34.210 10.225 34.460 10.395 ;
        POLYGON 34.460 10.395 34.630 10.225 34.460 10.225 ;
        POLYGON 2.140 10.225 2.140 10.095 2.010 10.095 ;
        RECT 2.140 10.095 2.230 10.225 ;
        POLYGON 2.230 10.225 2.360 10.225 2.230 10.095 ;
        POLYGON 2.510 10.225 2.640 10.225 2.640 10.095 ;
        RECT 2.640 10.095 2.730 10.225 ;
        POLYGON 2.730 10.225 2.860 10.095 2.730 10.095 ;
        POLYGON 5.040 10.225 5.040 10.095 4.910 10.095 ;
        RECT 5.040 10.095 5.130 10.225 ;
        POLYGON 5.130 10.225 5.260 10.225 5.130 10.095 ;
        POLYGON 5.410 10.225 5.540 10.225 5.540 10.095 ;
        RECT 5.540 10.095 5.630 10.225 ;
        POLYGON 5.630 10.225 5.760 10.095 5.630 10.095 ;
        POLYGON 7.940 10.225 7.940 10.095 7.810 10.095 ;
        RECT 7.940 10.095 8.030 10.225 ;
        POLYGON 8.030 10.225 8.160 10.225 8.030 10.095 ;
        POLYGON 8.310 10.225 8.440 10.225 8.440 10.095 ;
        RECT 8.440 10.095 8.530 10.225 ;
        POLYGON 8.530 10.225 8.660 10.095 8.530 10.095 ;
        POLYGON 10.840 10.225 10.840 10.095 10.710 10.095 ;
        RECT 10.840 10.095 10.930 10.225 ;
        POLYGON 10.930 10.225 11.060 10.225 10.930 10.095 ;
        POLYGON 11.210 10.225 11.340 10.225 11.340 10.095 ;
        RECT 11.340 10.095 11.430 10.225 ;
        POLYGON 11.430 10.225 11.560 10.095 11.430 10.095 ;
        POLYGON 13.740 10.225 13.740 10.095 13.610 10.095 ;
        RECT 13.740 10.095 13.830 10.225 ;
        POLYGON 13.830 10.225 13.960 10.225 13.830 10.095 ;
        POLYGON 14.110 10.225 14.240 10.225 14.240 10.095 ;
        RECT 14.240 10.095 14.330 10.225 ;
        POLYGON 14.330 10.225 14.460 10.095 14.330 10.095 ;
        POLYGON 16.640 10.225 16.640 10.095 16.510 10.095 ;
        RECT 16.640 10.095 16.730 10.225 ;
        POLYGON 16.730 10.225 16.860 10.225 16.730 10.095 ;
        POLYGON 17.010 10.225 17.140 10.225 17.140 10.095 ;
        RECT 17.140 10.095 17.230 10.225 ;
        POLYGON 17.230 10.225 17.360 10.095 17.230 10.095 ;
        POLYGON 19.540 10.225 19.540 10.095 19.410 10.095 ;
        RECT 19.540 10.095 19.630 10.225 ;
        POLYGON 19.630 10.225 19.760 10.225 19.630 10.095 ;
        POLYGON 19.910 10.225 20.040 10.225 20.040 10.095 ;
        RECT 20.040 10.095 20.130 10.225 ;
        POLYGON 20.130 10.225 20.260 10.095 20.130 10.095 ;
        POLYGON 22.440 10.225 22.440 10.095 22.310 10.095 ;
        RECT 22.440 10.095 22.530 10.225 ;
        POLYGON 22.530 10.225 22.660 10.225 22.530 10.095 ;
        POLYGON 22.810 10.225 22.940 10.225 22.940 10.095 ;
        RECT 22.940 10.095 23.030 10.225 ;
        POLYGON 23.030 10.225 23.160 10.095 23.030 10.095 ;
        POLYGON 25.340 10.225 25.340 10.095 25.210 10.095 ;
        RECT 25.340 10.095 25.430 10.225 ;
        POLYGON 25.430 10.225 25.560 10.225 25.430 10.095 ;
        POLYGON 25.710 10.225 25.840 10.225 25.840 10.095 ;
        RECT 25.840 10.095 25.930 10.225 ;
        POLYGON 25.930 10.225 26.060 10.095 25.930 10.095 ;
        POLYGON 28.240 10.225 28.240 10.095 28.110 10.095 ;
        RECT 28.240 10.095 28.330 10.225 ;
        POLYGON 28.330 10.225 28.460 10.225 28.330 10.095 ;
        POLYGON 28.610 10.225 28.740 10.225 28.740 10.095 ;
        RECT 28.740 10.095 28.830 10.225 ;
        POLYGON 28.830 10.225 28.960 10.095 28.830 10.095 ;
        POLYGON 31.140 10.225 31.140 10.095 31.010 10.095 ;
        RECT 31.140 10.095 31.230 10.225 ;
        POLYGON 31.230 10.225 31.360 10.225 31.230 10.095 ;
        POLYGON 31.510 10.225 31.640 10.225 31.640 10.095 ;
        RECT 31.640 10.095 31.730 10.225 ;
        POLYGON 31.730 10.225 31.860 10.095 31.730 10.095 ;
        POLYGON 34.040 10.225 34.040 10.095 33.910 10.095 ;
        RECT 34.040 10.095 34.130 10.225 ;
        POLYGON 34.130 10.225 34.260 10.225 34.130 10.095 ;
        POLYGON 34.410 10.225 34.540 10.225 34.540 10.095 ;
        RECT 34.540 10.095 34.630 10.225 ;
        POLYGON 34.630 10.225 34.760 10.095 34.630 10.095 ;
        RECT -0.275 9.925 2.060 10.095 ;
        POLYGON 2.060 10.095 2.230 10.095 2.060 9.925 ;
        POLYGON 2.640 10.095 2.810 10.095 2.810 9.925 ;
        RECT 2.810 9.925 4.960 10.095 ;
        POLYGON 4.960 10.095 5.130 10.095 4.960 9.925 ;
        RECT 5.525 9.925 7.860 10.095 ;
        POLYGON 7.860 10.095 8.030 10.095 7.860 9.925 ;
        POLYGON 8.440 10.095 8.610 10.095 8.610 9.925 ;
        RECT 8.610 9.925 10.760 10.095 ;
        POLYGON 10.760 10.095 10.930 10.095 10.760 9.925 ;
        RECT 11.325 9.925 13.660 10.095 ;
        POLYGON 13.660 10.095 13.830 10.095 13.660 9.925 ;
        POLYGON 14.240 10.095 14.410 10.095 14.410 9.925 ;
        RECT 14.410 9.925 16.560 10.095 ;
        POLYGON 16.560 10.095 16.730 10.095 16.560 9.925 ;
        RECT 17.125 9.925 19.460 10.095 ;
        POLYGON 19.460 10.095 19.630 10.095 19.460 9.925 ;
        POLYGON 20.040 10.095 20.210 10.095 20.210 9.925 ;
        RECT 20.210 9.925 22.360 10.095 ;
        POLYGON 22.360 10.095 22.530 10.095 22.360 9.925 ;
        RECT 22.925 9.925 25.260 10.095 ;
        POLYGON 25.260 10.095 25.430 10.095 25.260 9.925 ;
        POLYGON 25.840 10.095 26.010 10.095 26.010 9.925 ;
        RECT 26.010 9.925 28.160 10.095 ;
        POLYGON 28.160 10.095 28.330 10.095 28.160 9.925 ;
        RECT 28.725 9.925 31.060 10.095 ;
        POLYGON 31.060 10.095 31.230 10.095 31.060 9.925 ;
        POLYGON 31.640 10.095 31.810 10.095 31.810 9.925 ;
        RECT 31.810 9.925 33.960 10.095 ;
        POLYGON 33.960 10.095 34.130 10.095 33.960 9.925 ;
        POLYGON 34.540 10.095 34.710 10.095 34.710 9.925 ;
        RECT 34.710 9.925 34.760 10.095 ;
    END
  END RWL1_7
  PIN RWL0_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 11.275 2.510 11.445 ;
        RECT 5.260 11.275 5.410 11.445 ;
        RECT 8.160 11.275 8.310 11.445 ;
        RECT 11.060 11.275 11.210 11.445 ;
        RECT 13.960 11.275 14.110 11.445 ;
        RECT 16.860 11.275 17.010 11.445 ;
        RECT 19.760 11.275 19.910 11.445 ;
        RECT 22.660 11.275 22.810 11.445 ;
        RECT 25.560 11.275 25.710 11.445 ;
        RECT 28.460 11.275 28.610 11.445 ;
        RECT 31.360 11.275 31.510 11.445 ;
        RECT 34.260 11.275 34.410 11.445 ;
      LAYER mcon ;
        RECT 2.360 11.280 2.510 11.445 ;
        RECT 8.160 11.280 8.310 11.445 ;
        RECT 13.960 11.280 14.110 11.445 ;
        RECT 19.760 11.280 19.910 11.445 ;
        RECT 25.560 11.280 25.710 11.445 ;
        RECT 31.360 11.280 31.510 11.445 ;
      LAYER met1 ;
        RECT 2.360 11.275 2.510 11.445 ;
        RECT 5.260 11.275 5.410 11.445 ;
        RECT 8.160 11.275 8.310 11.445 ;
        RECT 11.060 11.275 11.210 11.445 ;
        RECT 13.960 11.275 14.110 11.445 ;
        RECT 16.860 11.275 17.010 11.445 ;
        RECT 19.760 11.275 19.910 11.445 ;
        RECT 22.660 11.275 22.810 11.445 ;
        RECT 25.560 11.275 25.710 11.445 ;
        RECT 28.460 11.275 28.610 11.445 ;
        RECT 31.360 11.275 31.510 11.445 ;
        RECT 34.260 11.275 34.410 11.445 ;
      LAYER met2 ;
        RECT -0.275 11.275 34.760 11.445 ;
    END
  END RWL0_8
  PIN RWL1_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 11.275 0.330 11.445 ;
        RECT 3.080 11.275 3.230 11.445 ;
        RECT 5.980 11.275 6.130 11.445 ;
        RECT 8.880 11.275 9.030 11.445 ;
        RECT 11.780 11.275 11.930 11.445 ;
        RECT 14.680 11.275 14.830 11.445 ;
        RECT 17.580 11.275 17.730 11.445 ;
        RECT 20.480 11.275 20.630 11.445 ;
        RECT 23.380 11.275 23.530 11.445 ;
        RECT 26.280 11.275 26.430 11.445 ;
        RECT 29.180 11.275 29.330 11.445 ;
        RECT 32.080 11.275 32.230 11.445 ;
      LAYER met1 ;
        POLYGON 2.310 11.745 2.310 11.575 2.140 11.575 ;
        RECT 2.310 11.575 2.560 11.745 ;
        POLYGON 2.560 11.745 2.730 11.575 2.560 11.575 ;
        POLYGON 5.210 11.745 5.210 11.575 5.040 11.575 ;
        RECT 5.210 11.575 5.460 11.745 ;
        POLYGON 5.460 11.745 5.630 11.575 5.460 11.575 ;
        POLYGON 8.110 11.745 8.110 11.575 7.940 11.575 ;
        RECT 8.110 11.575 8.360 11.745 ;
        POLYGON 8.360 11.745 8.530 11.575 8.360 11.575 ;
        POLYGON 11.010 11.745 11.010 11.575 10.840 11.575 ;
        RECT 11.010 11.575 11.260 11.745 ;
        POLYGON 11.260 11.745 11.430 11.575 11.260 11.575 ;
        POLYGON 13.910 11.745 13.910 11.575 13.740 11.575 ;
        RECT 13.910 11.575 14.160 11.745 ;
        POLYGON 14.160 11.745 14.330 11.575 14.160 11.575 ;
        POLYGON 16.810 11.745 16.810 11.575 16.640 11.575 ;
        RECT 16.810 11.575 17.060 11.745 ;
        POLYGON 17.060 11.745 17.230 11.575 17.060 11.575 ;
        POLYGON 19.710 11.745 19.710 11.575 19.540 11.575 ;
        RECT 19.710 11.575 19.960 11.745 ;
        POLYGON 19.960 11.745 20.130 11.575 19.960 11.575 ;
        POLYGON 22.610 11.745 22.610 11.575 22.440 11.575 ;
        RECT 22.610 11.575 22.860 11.745 ;
        POLYGON 22.860 11.745 23.030 11.575 22.860 11.575 ;
        POLYGON 25.510 11.745 25.510 11.575 25.340 11.575 ;
        RECT 25.510 11.575 25.760 11.745 ;
        POLYGON 25.760 11.745 25.930 11.575 25.760 11.575 ;
        POLYGON 28.410 11.745 28.410 11.575 28.240 11.575 ;
        RECT 28.410 11.575 28.660 11.745 ;
        POLYGON 28.660 11.745 28.830 11.575 28.660 11.575 ;
        POLYGON 31.310 11.745 31.310 11.575 31.140 11.575 ;
        RECT 31.310 11.575 31.560 11.745 ;
        POLYGON 31.560 11.745 31.730 11.575 31.560 11.575 ;
        POLYGON 34.210 11.745 34.210 11.575 34.040 11.575 ;
        RECT 34.210 11.575 34.460 11.745 ;
        POLYGON 34.460 11.745 34.630 11.575 34.460 11.575 ;
        POLYGON 2.140 11.575 2.140 11.445 2.010 11.445 ;
        RECT 2.140 11.445 2.230 11.575 ;
        POLYGON 2.230 11.575 2.360 11.575 2.230 11.445 ;
        POLYGON 2.510 11.575 2.640 11.575 2.640 11.445 ;
        RECT 2.640 11.445 2.730 11.575 ;
        POLYGON 2.730 11.575 2.860 11.445 2.730 11.445 ;
        POLYGON 5.040 11.575 5.040 11.445 4.910 11.445 ;
        RECT 5.040 11.445 5.130 11.575 ;
        POLYGON 5.130 11.575 5.260 11.575 5.130 11.445 ;
        POLYGON 5.410 11.575 5.540 11.575 5.540 11.445 ;
        RECT 5.540 11.445 5.630 11.575 ;
        POLYGON 5.630 11.575 5.760 11.445 5.630 11.445 ;
        POLYGON 7.940 11.575 7.940 11.445 7.810 11.445 ;
        RECT 7.940 11.445 8.030 11.575 ;
        POLYGON 8.030 11.575 8.160 11.575 8.030 11.445 ;
        POLYGON 8.310 11.575 8.440 11.575 8.440 11.445 ;
        RECT 8.440 11.445 8.530 11.575 ;
        POLYGON 8.530 11.575 8.660 11.445 8.530 11.445 ;
        POLYGON 10.840 11.575 10.840 11.445 10.710 11.445 ;
        RECT 10.840 11.445 10.930 11.575 ;
        POLYGON 10.930 11.575 11.060 11.575 10.930 11.445 ;
        POLYGON 11.210 11.575 11.340 11.575 11.340 11.445 ;
        RECT 11.340 11.445 11.430 11.575 ;
        POLYGON 11.430 11.575 11.560 11.445 11.430 11.445 ;
        POLYGON 13.740 11.575 13.740 11.445 13.610 11.445 ;
        RECT 13.740 11.445 13.830 11.575 ;
        POLYGON 13.830 11.575 13.960 11.575 13.830 11.445 ;
        POLYGON 14.110 11.575 14.240 11.575 14.240 11.445 ;
        RECT 14.240 11.445 14.330 11.575 ;
        POLYGON 14.330 11.575 14.460 11.445 14.330 11.445 ;
        POLYGON 16.640 11.575 16.640 11.445 16.510 11.445 ;
        RECT 16.640 11.445 16.730 11.575 ;
        POLYGON 16.730 11.575 16.860 11.575 16.730 11.445 ;
        POLYGON 17.010 11.575 17.140 11.575 17.140 11.445 ;
        RECT 17.140 11.445 17.230 11.575 ;
        POLYGON 17.230 11.575 17.360 11.445 17.230 11.445 ;
        POLYGON 19.540 11.575 19.540 11.445 19.410 11.445 ;
        RECT 19.540 11.445 19.630 11.575 ;
        POLYGON 19.630 11.575 19.760 11.575 19.630 11.445 ;
        POLYGON 19.910 11.575 20.040 11.575 20.040 11.445 ;
        RECT 20.040 11.445 20.130 11.575 ;
        POLYGON 20.130 11.575 20.260 11.445 20.130 11.445 ;
        POLYGON 22.440 11.575 22.440 11.445 22.310 11.445 ;
        RECT 22.440 11.445 22.530 11.575 ;
        POLYGON 22.530 11.575 22.660 11.575 22.530 11.445 ;
        POLYGON 22.810 11.575 22.940 11.575 22.940 11.445 ;
        RECT 22.940 11.445 23.030 11.575 ;
        POLYGON 23.030 11.575 23.160 11.445 23.030 11.445 ;
        POLYGON 25.340 11.575 25.340 11.445 25.210 11.445 ;
        RECT 25.340 11.445 25.430 11.575 ;
        POLYGON 25.430 11.575 25.560 11.575 25.430 11.445 ;
        POLYGON 25.710 11.575 25.840 11.575 25.840 11.445 ;
        RECT 25.840 11.445 25.930 11.575 ;
        POLYGON 25.930 11.575 26.060 11.445 25.930 11.445 ;
        POLYGON 28.240 11.575 28.240 11.445 28.110 11.445 ;
        RECT 28.240 11.445 28.330 11.575 ;
        POLYGON 28.330 11.575 28.460 11.575 28.330 11.445 ;
        POLYGON 28.610 11.575 28.740 11.575 28.740 11.445 ;
        RECT 28.740 11.445 28.830 11.575 ;
        POLYGON 28.830 11.575 28.960 11.445 28.830 11.445 ;
        POLYGON 31.140 11.575 31.140 11.445 31.010 11.445 ;
        RECT 31.140 11.445 31.230 11.575 ;
        POLYGON 31.230 11.575 31.360 11.575 31.230 11.445 ;
        POLYGON 31.510 11.575 31.640 11.575 31.640 11.445 ;
        RECT 31.640 11.445 31.730 11.575 ;
        POLYGON 31.730 11.575 31.860 11.445 31.730 11.445 ;
        POLYGON 34.040 11.575 34.040 11.445 33.910 11.445 ;
        RECT 34.040 11.445 34.130 11.575 ;
        POLYGON 34.130 11.575 34.260 11.575 34.130 11.445 ;
        POLYGON 34.410 11.575 34.540 11.575 34.540 11.445 ;
        RECT 34.540 11.445 34.630 11.575 ;
        POLYGON 34.630 11.575 34.760 11.445 34.630 11.445 ;
        RECT -0.275 11.275 2.060 11.445 ;
        POLYGON 2.060 11.445 2.230 11.445 2.060 11.275 ;
        POLYGON 2.640 11.445 2.810 11.445 2.810 11.275 ;
        RECT 2.810 11.275 4.960 11.445 ;
        POLYGON 4.960 11.445 5.130 11.445 4.960 11.275 ;
        RECT 5.525 11.275 7.860 11.445 ;
        POLYGON 7.860 11.445 8.030 11.445 7.860 11.275 ;
        POLYGON 8.440 11.445 8.610 11.445 8.610 11.275 ;
        RECT 8.610 11.275 10.760 11.445 ;
        POLYGON 10.760 11.445 10.930 11.445 10.760 11.275 ;
        RECT 11.325 11.275 13.660 11.445 ;
        POLYGON 13.660 11.445 13.830 11.445 13.660 11.275 ;
        POLYGON 14.240 11.445 14.410 11.445 14.410 11.275 ;
        RECT 14.410 11.275 16.560 11.445 ;
        POLYGON 16.560 11.445 16.730 11.445 16.560 11.275 ;
        RECT 17.125 11.275 19.460 11.445 ;
        POLYGON 19.460 11.445 19.630 11.445 19.460 11.275 ;
        POLYGON 20.040 11.445 20.210 11.445 20.210 11.275 ;
        RECT 20.210 11.275 22.360 11.445 ;
        POLYGON 22.360 11.445 22.530 11.445 22.360 11.275 ;
        RECT 22.925 11.275 25.260 11.445 ;
        POLYGON 25.260 11.445 25.430 11.445 25.260 11.275 ;
        POLYGON 25.840 11.445 26.010 11.445 26.010 11.275 ;
        RECT 26.010 11.275 28.160 11.445 ;
        POLYGON 28.160 11.445 28.330 11.445 28.160 11.275 ;
        RECT 28.725 11.275 31.060 11.445 ;
        POLYGON 31.060 11.445 31.230 11.445 31.060 11.275 ;
        POLYGON 31.640 11.445 31.810 11.445 31.810 11.275 ;
        RECT 31.810 11.275 33.960 11.445 ;
        POLYGON 33.960 11.445 34.130 11.445 33.960 11.275 ;
        POLYGON 34.540 11.445 34.710 11.445 34.710 11.275 ;
        RECT 34.710 11.275 34.760 11.445 ;
    END
  END RWL1_8
  PIN RWL0_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 12.625 2.510 12.795 ;
        RECT 5.260 12.625 5.410 12.795 ;
        RECT 8.160 12.625 8.310 12.795 ;
        RECT 11.060 12.625 11.210 12.795 ;
        RECT 13.960 12.625 14.110 12.795 ;
        RECT 16.860 12.625 17.010 12.795 ;
        RECT 19.760 12.625 19.910 12.795 ;
        RECT 22.660 12.625 22.810 12.795 ;
        RECT 25.560 12.625 25.710 12.795 ;
        RECT 28.460 12.625 28.610 12.795 ;
        RECT 31.360 12.625 31.510 12.795 ;
        RECT 34.260 12.625 34.410 12.795 ;
      LAYER mcon ;
        RECT 2.360 12.630 2.510 12.795 ;
        RECT 8.160 12.630 8.310 12.795 ;
        RECT 13.960 12.630 14.110 12.795 ;
        RECT 19.760 12.630 19.910 12.795 ;
        RECT 25.560 12.630 25.710 12.795 ;
        RECT 31.360 12.630 31.510 12.795 ;
      LAYER met1 ;
        RECT 2.360 12.625 2.510 12.795 ;
        RECT 5.260 12.625 5.410 12.795 ;
        RECT 8.160 12.625 8.310 12.795 ;
        RECT 11.060 12.625 11.210 12.795 ;
        RECT 13.960 12.625 14.110 12.795 ;
        RECT 16.860 12.625 17.010 12.795 ;
        RECT 19.760 12.625 19.910 12.795 ;
        RECT 22.660 12.625 22.810 12.795 ;
        RECT 25.560 12.625 25.710 12.795 ;
        RECT 28.460 12.625 28.610 12.795 ;
        RECT 31.360 12.625 31.510 12.795 ;
        RECT 34.260 12.625 34.410 12.795 ;
      LAYER met2 ;
        RECT -0.275 12.625 34.760 12.795 ;
    END
  END RWL0_9
  PIN RWL1_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 12.625 0.330 12.795 ;
        RECT 3.080 12.625 3.230 12.795 ;
        RECT 5.980 12.625 6.130 12.795 ;
        RECT 8.880 12.625 9.030 12.795 ;
        RECT 11.780 12.625 11.930 12.795 ;
        RECT 14.680 12.625 14.830 12.795 ;
        RECT 17.580 12.625 17.730 12.795 ;
        RECT 20.480 12.625 20.630 12.795 ;
        RECT 23.380 12.625 23.530 12.795 ;
        RECT 26.280 12.625 26.430 12.795 ;
        RECT 29.180 12.625 29.330 12.795 ;
        RECT 32.080 12.625 32.230 12.795 ;
      LAYER met1 ;
        POLYGON 2.310 13.095 2.310 12.925 2.140 12.925 ;
        RECT 2.310 12.925 2.560 13.095 ;
        POLYGON 2.560 13.095 2.730 12.925 2.560 12.925 ;
        POLYGON 5.210 13.095 5.210 12.925 5.040 12.925 ;
        RECT 5.210 12.925 5.460 13.095 ;
        POLYGON 5.460 13.095 5.630 12.925 5.460 12.925 ;
        POLYGON 8.110 13.095 8.110 12.925 7.940 12.925 ;
        RECT 8.110 12.925 8.360 13.095 ;
        POLYGON 8.360 13.095 8.530 12.925 8.360 12.925 ;
        POLYGON 11.010 13.095 11.010 12.925 10.840 12.925 ;
        RECT 11.010 12.925 11.260 13.095 ;
        POLYGON 11.260 13.095 11.430 12.925 11.260 12.925 ;
        POLYGON 13.910 13.095 13.910 12.925 13.740 12.925 ;
        RECT 13.910 12.925 14.160 13.095 ;
        POLYGON 14.160 13.095 14.330 12.925 14.160 12.925 ;
        POLYGON 16.810 13.095 16.810 12.925 16.640 12.925 ;
        RECT 16.810 12.925 17.060 13.095 ;
        POLYGON 17.060 13.095 17.230 12.925 17.060 12.925 ;
        POLYGON 19.710 13.095 19.710 12.925 19.540 12.925 ;
        RECT 19.710 12.925 19.960 13.095 ;
        POLYGON 19.960 13.095 20.130 12.925 19.960 12.925 ;
        POLYGON 22.610 13.095 22.610 12.925 22.440 12.925 ;
        RECT 22.610 12.925 22.860 13.095 ;
        POLYGON 22.860 13.095 23.030 12.925 22.860 12.925 ;
        POLYGON 25.510 13.095 25.510 12.925 25.340 12.925 ;
        RECT 25.510 12.925 25.760 13.095 ;
        POLYGON 25.760 13.095 25.930 12.925 25.760 12.925 ;
        POLYGON 28.410 13.095 28.410 12.925 28.240 12.925 ;
        RECT 28.410 12.925 28.660 13.095 ;
        POLYGON 28.660 13.095 28.830 12.925 28.660 12.925 ;
        POLYGON 31.310 13.095 31.310 12.925 31.140 12.925 ;
        RECT 31.310 12.925 31.560 13.095 ;
        POLYGON 31.560 13.095 31.730 12.925 31.560 12.925 ;
        POLYGON 34.210 13.095 34.210 12.925 34.040 12.925 ;
        RECT 34.210 12.925 34.460 13.095 ;
        POLYGON 34.460 13.095 34.630 12.925 34.460 12.925 ;
        POLYGON 2.140 12.925 2.140 12.795 2.010 12.795 ;
        RECT 2.140 12.795 2.230 12.925 ;
        POLYGON 2.230 12.925 2.360 12.925 2.230 12.795 ;
        POLYGON 2.510 12.925 2.640 12.925 2.640 12.795 ;
        RECT 2.640 12.795 2.730 12.925 ;
        POLYGON 2.730 12.925 2.860 12.795 2.730 12.795 ;
        POLYGON 5.040 12.925 5.040 12.795 4.910 12.795 ;
        RECT 5.040 12.795 5.130 12.925 ;
        POLYGON 5.130 12.925 5.260 12.925 5.130 12.795 ;
        POLYGON 5.410 12.925 5.540 12.925 5.540 12.795 ;
        RECT 5.540 12.795 5.630 12.925 ;
        POLYGON 5.630 12.925 5.760 12.795 5.630 12.795 ;
        POLYGON 7.940 12.925 7.940 12.795 7.810 12.795 ;
        RECT 7.940 12.795 8.030 12.925 ;
        POLYGON 8.030 12.925 8.160 12.925 8.030 12.795 ;
        POLYGON 8.310 12.925 8.440 12.925 8.440 12.795 ;
        RECT 8.440 12.795 8.530 12.925 ;
        POLYGON 8.530 12.925 8.660 12.795 8.530 12.795 ;
        POLYGON 10.840 12.925 10.840 12.795 10.710 12.795 ;
        RECT 10.840 12.795 10.930 12.925 ;
        POLYGON 10.930 12.925 11.060 12.925 10.930 12.795 ;
        POLYGON 11.210 12.925 11.340 12.925 11.340 12.795 ;
        RECT 11.340 12.795 11.430 12.925 ;
        POLYGON 11.430 12.925 11.560 12.795 11.430 12.795 ;
        POLYGON 13.740 12.925 13.740 12.795 13.610 12.795 ;
        RECT 13.740 12.795 13.830 12.925 ;
        POLYGON 13.830 12.925 13.960 12.925 13.830 12.795 ;
        POLYGON 14.110 12.925 14.240 12.925 14.240 12.795 ;
        RECT 14.240 12.795 14.330 12.925 ;
        POLYGON 14.330 12.925 14.460 12.795 14.330 12.795 ;
        POLYGON 16.640 12.925 16.640 12.795 16.510 12.795 ;
        RECT 16.640 12.795 16.730 12.925 ;
        POLYGON 16.730 12.925 16.860 12.925 16.730 12.795 ;
        POLYGON 17.010 12.925 17.140 12.925 17.140 12.795 ;
        RECT 17.140 12.795 17.230 12.925 ;
        POLYGON 17.230 12.925 17.360 12.795 17.230 12.795 ;
        POLYGON 19.540 12.925 19.540 12.795 19.410 12.795 ;
        RECT 19.540 12.795 19.630 12.925 ;
        POLYGON 19.630 12.925 19.760 12.925 19.630 12.795 ;
        POLYGON 19.910 12.925 20.040 12.925 20.040 12.795 ;
        RECT 20.040 12.795 20.130 12.925 ;
        POLYGON 20.130 12.925 20.260 12.795 20.130 12.795 ;
        POLYGON 22.440 12.925 22.440 12.795 22.310 12.795 ;
        RECT 22.440 12.795 22.530 12.925 ;
        POLYGON 22.530 12.925 22.660 12.925 22.530 12.795 ;
        POLYGON 22.810 12.925 22.940 12.925 22.940 12.795 ;
        RECT 22.940 12.795 23.030 12.925 ;
        POLYGON 23.030 12.925 23.160 12.795 23.030 12.795 ;
        POLYGON 25.340 12.925 25.340 12.795 25.210 12.795 ;
        RECT 25.340 12.795 25.430 12.925 ;
        POLYGON 25.430 12.925 25.560 12.925 25.430 12.795 ;
        POLYGON 25.710 12.925 25.840 12.925 25.840 12.795 ;
        RECT 25.840 12.795 25.930 12.925 ;
        POLYGON 25.930 12.925 26.060 12.795 25.930 12.795 ;
        POLYGON 28.240 12.925 28.240 12.795 28.110 12.795 ;
        RECT 28.240 12.795 28.330 12.925 ;
        POLYGON 28.330 12.925 28.460 12.925 28.330 12.795 ;
        POLYGON 28.610 12.925 28.740 12.925 28.740 12.795 ;
        RECT 28.740 12.795 28.830 12.925 ;
        POLYGON 28.830 12.925 28.960 12.795 28.830 12.795 ;
        POLYGON 31.140 12.925 31.140 12.795 31.010 12.795 ;
        RECT 31.140 12.795 31.230 12.925 ;
        POLYGON 31.230 12.925 31.360 12.925 31.230 12.795 ;
        POLYGON 31.510 12.925 31.640 12.925 31.640 12.795 ;
        RECT 31.640 12.795 31.730 12.925 ;
        POLYGON 31.730 12.925 31.860 12.795 31.730 12.795 ;
        POLYGON 34.040 12.925 34.040 12.795 33.910 12.795 ;
        RECT 34.040 12.795 34.130 12.925 ;
        POLYGON 34.130 12.925 34.260 12.925 34.130 12.795 ;
        POLYGON 34.410 12.925 34.540 12.925 34.540 12.795 ;
        RECT 34.540 12.795 34.630 12.925 ;
        POLYGON 34.630 12.925 34.760 12.795 34.630 12.795 ;
        RECT -0.275 12.625 2.060 12.795 ;
        POLYGON 2.060 12.795 2.230 12.795 2.060 12.625 ;
        POLYGON 2.640 12.795 2.810 12.795 2.810 12.625 ;
        RECT 2.810 12.625 4.960 12.795 ;
        POLYGON 4.960 12.795 5.130 12.795 4.960 12.625 ;
        RECT 5.525 12.625 7.860 12.795 ;
        POLYGON 7.860 12.795 8.030 12.795 7.860 12.625 ;
        POLYGON 8.440 12.795 8.610 12.795 8.610 12.625 ;
        RECT 8.610 12.625 10.760 12.795 ;
        POLYGON 10.760 12.795 10.930 12.795 10.760 12.625 ;
        RECT 11.325 12.625 13.660 12.795 ;
        POLYGON 13.660 12.795 13.830 12.795 13.660 12.625 ;
        POLYGON 14.240 12.795 14.410 12.795 14.410 12.625 ;
        RECT 14.410 12.625 16.560 12.795 ;
        POLYGON 16.560 12.795 16.730 12.795 16.560 12.625 ;
        RECT 17.125 12.625 19.460 12.795 ;
        POLYGON 19.460 12.795 19.630 12.795 19.460 12.625 ;
        POLYGON 20.040 12.795 20.210 12.795 20.210 12.625 ;
        RECT 20.210 12.625 22.360 12.795 ;
        POLYGON 22.360 12.795 22.530 12.795 22.360 12.625 ;
        RECT 22.925 12.625 25.260 12.795 ;
        POLYGON 25.260 12.795 25.430 12.795 25.260 12.625 ;
        POLYGON 25.840 12.795 26.010 12.795 26.010 12.625 ;
        RECT 26.010 12.625 28.160 12.795 ;
        POLYGON 28.160 12.795 28.330 12.795 28.160 12.625 ;
        RECT 28.725 12.625 31.060 12.795 ;
        POLYGON 31.060 12.795 31.230 12.795 31.060 12.625 ;
        POLYGON 31.640 12.795 31.810 12.795 31.810 12.625 ;
        RECT 31.810 12.625 33.960 12.795 ;
        POLYGON 33.960 12.795 34.130 12.795 33.960 12.625 ;
        POLYGON 34.540 12.795 34.710 12.795 34.710 12.625 ;
        RECT 34.710 12.625 34.760 12.795 ;
    END
  END RWL1_9
  PIN RWL0_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 13.975 2.510 14.145 ;
        RECT 5.260 13.975 5.410 14.145 ;
        RECT 8.160 13.975 8.310 14.145 ;
        RECT 11.060 13.975 11.210 14.145 ;
        RECT 13.960 13.975 14.110 14.145 ;
        RECT 16.860 13.975 17.010 14.145 ;
        RECT 19.760 13.975 19.910 14.145 ;
        RECT 22.660 13.975 22.810 14.145 ;
        RECT 25.560 13.975 25.710 14.145 ;
        RECT 28.460 13.975 28.610 14.145 ;
        RECT 31.360 13.975 31.510 14.145 ;
        RECT 34.260 13.975 34.410 14.145 ;
      LAYER mcon ;
        RECT 2.360 13.980 2.510 14.145 ;
        RECT 8.160 13.980 8.310 14.145 ;
        RECT 13.960 13.980 14.110 14.145 ;
        RECT 19.760 13.980 19.910 14.145 ;
        RECT 25.560 13.980 25.710 14.145 ;
        RECT 31.360 13.980 31.510 14.145 ;
      LAYER met1 ;
        RECT 2.360 13.975 2.510 14.145 ;
        RECT 5.260 13.975 5.410 14.145 ;
        RECT 8.160 13.975 8.310 14.145 ;
        RECT 11.060 13.975 11.210 14.145 ;
        RECT 13.960 13.975 14.110 14.145 ;
        RECT 16.860 13.975 17.010 14.145 ;
        RECT 19.760 13.975 19.910 14.145 ;
        RECT 22.660 13.975 22.810 14.145 ;
        RECT 25.560 13.975 25.710 14.145 ;
        RECT 28.460 13.975 28.610 14.145 ;
        RECT 31.360 13.975 31.510 14.145 ;
        RECT 34.260 13.975 34.410 14.145 ;
      LAYER met2 ;
        RECT -0.275 13.975 34.760 14.145 ;
    END
  END RWL0_10
  PIN RWL1_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 13.975 0.330 14.145 ;
        RECT 3.080 13.975 3.230 14.145 ;
        RECT 5.980 13.975 6.130 14.145 ;
        RECT 8.880 13.975 9.030 14.145 ;
        RECT 11.780 13.975 11.930 14.145 ;
        RECT 14.680 13.975 14.830 14.145 ;
        RECT 17.580 13.975 17.730 14.145 ;
        RECT 20.480 13.975 20.630 14.145 ;
        RECT 23.380 13.975 23.530 14.145 ;
        RECT 26.280 13.975 26.430 14.145 ;
        RECT 29.180 13.975 29.330 14.145 ;
        RECT 32.080 13.975 32.230 14.145 ;
      LAYER met1 ;
        POLYGON 2.310 14.445 2.310 14.275 2.140 14.275 ;
        RECT 2.310 14.275 2.560 14.445 ;
        POLYGON 2.560 14.445 2.730 14.275 2.560 14.275 ;
        POLYGON 5.210 14.445 5.210 14.275 5.040 14.275 ;
        RECT 5.210 14.275 5.460 14.445 ;
        POLYGON 5.460 14.445 5.630 14.275 5.460 14.275 ;
        POLYGON 8.110 14.445 8.110 14.275 7.940 14.275 ;
        RECT 8.110 14.275 8.360 14.445 ;
        POLYGON 8.360 14.445 8.530 14.275 8.360 14.275 ;
        POLYGON 11.010 14.445 11.010 14.275 10.840 14.275 ;
        RECT 11.010 14.275 11.260 14.445 ;
        POLYGON 11.260 14.445 11.430 14.275 11.260 14.275 ;
        POLYGON 13.910 14.445 13.910 14.275 13.740 14.275 ;
        RECT 13.910 14.275 14.160 14.445 ;
        POLYGON 14.160 14.445 14.330 14.275 14.160 14.275 ;
        POLYGON 16.810 14.445 16.810 14.275 16.640 14.275 ;
        RECT 16.810 14.275 17.060 14.445 ;
        POLYGON 17.060 14.445 17.230 14.275 17.060 14.275 ;
        POLYGON 19.710 14.445 19.710 14.275 19.540 14.275 ;
        RECT 19.710 14.275 19.960 14.445 ;
        POLYGON 19.960 14.445 20.130 14.275 19.960 14.275 ;
        POLYGON 22.610 14.445 22.610 14.275 22.440 14.275 ;
        RECT 22.610 14.275 22.860 14.445 ;
        POLYGON 22.860 14.445 23.030 14.275 22.860 14.275 ;
        POLYGON 25.510 14.445 25.510 14.275 25.340 14.275 ;
        RECT 25.510 14.275 25.760 14.445 ;
        POLYGON 25.760 14.445 25.930 14.275 25.760 14.275 ;
        POLYGON 28.410 14.445 28.410 14.275 28.240 14.275 ;
        RECT 28.410 14.275 28.660 14.445 ;
        POLYGON 28.660 14.445 28.830 14.275 28.660 14.275 ;
        POLYGON 31.310 14.445 31.310 14.275 31.140 14.275 ;
        RECT 31.310 14.275 31.560 14.445 ;
        POLYGON 31.560 14.445 31.730 14.275 31.560 14.275 ;
        POLYGON 34.210 14.445 34.210 14.275 34.040 14.275 ;
        RECT 34.210 14.275 34.460 14.445 ;
        POLYGON 34.460 14.445 34.630 14.275 34.460 14.275 ;
        POLYGON 2.140 14.275 2.140 14.145 2.010 14.145 ;
        RECT 2.140 14.145 2.230 14.275 ;
        POLYGON 2.230 14.275 2.360 14.275 2.230 14.145 ;
        POLYGON 2.510 14.275 2.640 14.275 2.640 14.145 ;
        RECT 2.640 14.145 2.730 14.275 ;
        POLYGON 2.730 14.275 2.860 14.145 2.730 14.145 ;
        POLYGON 5.040 14.275 5.040 14.145 4.910 14.145 ;
        RECT 5.040 14.145 5.130 14.275 ;
        POLYGON 5.130 14.275 5.260 14.275 5.130 14.145 ;
        POLYGON 5.410 14.275 5.540 14.275 5.540 14.145 ;
        RECT 5.540 14.145 5.630 14.275 ;
        POLYGON 5.630 14.275 5.760 14.145 5.630 14.145 ;
        POLYGON 7.940 14.275 7.940 14.145 7.810 14.145 ;
        RECT 7.940 14.145 8.030 14.275 ;
        POLYGON 8.030 14.275 8.160 14.275 8.030 14.145 ;
        POLYGON 8.310 14.275 8.440 14.275 8.440 14.145 ;
        RECT 8.440 14.145 8.530 14.275 ;
        POLYGON 8.530 14.275 8.660 14.145 8.530 14.145 ;
        POLYGON 10.840 14.275 10.840 14.145 10.710 14.145 ;
        RECT 10.840 14.145 10.930 14.275 ;
        POLYGON 10.930 14.275 11.060 14.275 10.930 14.145 ;
        POLYGON 11.210 14.275 11.340 14.275 11.340 14.145 ;
        RECT 11.340 14.145 11.430 14.275 ;
        POLYGON 11.430 14.275 11.560 14.145 11.430 14.145 ;
        POLYGON 13.740 14.275 13.740 14.145 13.610 14.145 ;
        RECT 13.740 14.145 13.830 14.275 ;
        POLYGON 13.830 14.275 13.960 14.275 13.830 14.145 ;
        POLYGON 14.110 14.275 14.240 14.275 14.240 14.145 ;
        RECT 14.240 14.145 14.330 14.275 ;
        POLYGON 14.330 14.275 14.460 14.145 14.330 14.145 ;
        POLYGON 16.640 14.275 16.640 14.145 16.510 14.145 ;
        RECT 16.640 14.145 16.730 14.275 ;
        POLYGON 16.730 14.275 16.860 14.275 16.730 14.145 ;
        POLYGON 17.010 14.275 17.140 14.275 17.140 14.145 ;
        RECT 17.140 14.145 17.230 14.275 ;
        POLYGON 17.230 14.275 17.360 14.145 17.230 14.145 ;
        POLYGON 19.540 14.275 19.540 14.145 19.410 14.145 ;
        RECT 19.540 14.145 19.630 14.275 ;
        POLYGON 19.630 14.275 19.760 14.275 19.630 14.145 ;
        POLYGON 19.910 14.275 20.040 14.275 20.040 14.145 ;
        RECT 20.040 14.145 20.130 14.275 ;
        POLYGON 20.130 14.275 20.260 14.145 20.130 14.145 ;
        POLYGON 22.440 14.275 22.440 14.145 22.310 14.145 ;
        RECT 22.440 14.145 22.530 14.275 ;
        POLYGON 22.530 14.275 22.660 14.275 22.530 14.145 ;
        POLYGON 22.810 14.275 22.940 14.275 22.940 14.145 ;
        RECT 22.940 14.145 23.030 14.275 ;
        POLYGON 23.030 14.275 23.160 14.145 23.030 14.145 ;
        POLYGON 25.340 14.275 25.340 14.145 25.210 14.145 ;
        RECT 25.340 14.145 25.430 14.275 ;
        POLYGON 25.430 14.275 25.560 14.275 25.430 14.145 ;
        POLYGON 25.710 14.275 25.840 14.275 25.840 14.145 ;
        RECT 25.840 14.145 25.930 14.275 ;
        POLYGON 25.930 14.275 26.060 14.145 25.930 14.145 ;
        POLYGON 28.240 14.275 28.240 14.145 28.110 14.145 ;
        RECT 28.240 14.145 28.330 14.275 ;
        POLYGON 28.330 14.275 28.460 14.275 28.330 14.145 ;
        POLYGON 28.610 14.275 28.740 14.275 28.740 14.145 ;
        RECT 28.740 14.145 28.830 14.275 ;
        POLYGON 28.830 14.275 28.960 14.145 28.830 14.145 ;
        POLYGON 31.140 14.275 31.140 14.145 31.010 14.145 ;
        RECT 31.140 14.145 31.230 14.275 ;
        POLYGON 31.230 14.275 31.360 14.275 31.230 14.145 ;
        POLYGON 31.510 14.275 31.640 14.275 31.640 14.145 ;
        RECT 31.640 14.145 31.730 14.275 ;
        POLYGON 31.730 14.275 31.860 14.145 31.730 14.145 ;
        POLYGON 34.040 14.275 34.040 14.145 33.910 14.145 ;
        RECT 34.040 14.145 34.130 14.275 ;
        POLYGON 34.130 14.275 34.260 14.275 34.130 14.145 ;
        POLYGON 34.410 14.275 34.540 14.275 34.540 14.145 ;
        RECT 34.540 14.145 34.630 14.275 ;
        POLYGON 34.630 14.275 34.760 14.145 34.630 14.145 ;
        RECT -0.275 13.975 2.060 14.145 ;
        POLYGON 2.060 14.145 2.230 14.145 2.060 13.975 ;
        POLYGON 2.640 14.145 2.810 14.145 2.810 13.975 ;
        RECT 2.810 13.975 4.960 14.145 ;
        POLYGON 4.960 14.145 5.130 14.145 4.960 13.975 ;
        RECT 5.525 13.975 7.860 14.145 ;
        POLYGON 7.860 14.145 8.030 14.145 7.860 13.975 ;
        POLYGON 8.440 14.145 8.610 14.145 8.610 13.975 ;
        RECT 8.610 13.975 10.760 14.145 ;
        POLYGON 10.760 14.145 10.930 14.145 10.760 13.975 ;
        RECT 11.325 13.975 13.660 14.145 ;
        POLYGON 13.660 14.145 13.830 14.145 13.660 13.975 ;
        POLYGON 14.240 14.145 14.410 14.145 14.410 13.975 ;
        RECT 14.410 13.975 16.560 14.145 ;
        POLYGON 16.560 14.145 16.730 14.145 16.560 13.975 ;
        RECT 17.125 13.975 19.460 14.145 ;
        POLYGON 19.460 14.145 19.630 14.145 19.460 13.975 ;
        POLYGON 20.040 14.145 20.210 14.145 20.210 13.975 ;
        RECT 20.210 13.975 22.360 14.145 ;
        POLYGON 22.360 14.145 22.530 14.145 22.360 13.975 ;
        RECT 22.925 13.975 25.260 14.145 ;
        POLYGON 25.260 14.145 25.430 14.145 25.260 13.975 ;
        POLYGON 25.840 14.145 26.010 14.145 26.010 13.975 ;
        RECT 26.010 13.975 28.160 14.145 ;
        POLYGON 28.160 14.145 28.330 14.145 28.160 13.975 ;
        RECT 28.725 13.975 31.060 14.145 ;
        POLYGON 31.060 14.145 31.230 14.145 31.060 13.975 ;
        POLYGON 31.640 14.145 31.810 14.145 31.810 13.975 ;
        RECT 31.810 13.975 33.960 14.145 ;
        POLYGON 33.960 14.145 34.130 14.145 33.960 13.975 ;
        POLYGON 34.540 14.145 34.710 14.145 34.710 13.975 ;
        RECT 34.710 13.975 34.760 14.145 ;
    END
  END RWL1_10
  PIN RWL0_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 15.325 2.510 15.495 ;
        RECT 5.260 15.325 5.410 15.495 ;
        RECT 8.160 15.325 8.310 15.495 ;
        RECT 11.060 15.325 11.210 15.495 ;
        RECT 13.960 15.325 14.110 15.495 ;
        RECT 16.860 15.325 17.010 15.495 ;
        RECT 19.760 15.325 19.910 15.495 ;
        RECT 22.660 15.325 22.810 15.495 ;
        RECT 25.560 15.325 25.710 15.495 ;
        RECT 28.460 15.325 28.610 15.495 ;
        RECT 31.360 15.325 31.510 15.495 ;
        RECT 34.260 15.325 34.410 15.495 ;
      LAYER mcon ;
        RECT 2.360 15.330 2.510 15.495 ;
        RECT 8.160 15.330 8.310 15.495 ;
        RECT 13.960 15.330 14.110 15.495 ;
        RECT 19.760 15.330 19.910 15.495 ;
        RECT 25.560 15.330 25.710 15.495 ;
        RECT 31.360 15.330 31.510 15.495 ;
      LAYER met1 ;
        RECT 2.360 15.325 2.510 15.495 ;
        RECT 5.260 15.325 5.410 15.495 ;
        RECT 8.160 15.325 8.310 15.495 ;
        RECT 11.060 15.325 11.210 15.495 ;
        RECT 13.960 15.325 14.110 15.495 ;
        RECT 16.860 15.325 17.010 15.495 ;
        RECT 19.760 15.325 19.910 15.495 ;
        RECT 22.660 15.325 22.810 15.495 ;
        RECT 25.560 15.325 25.710 15.495 ;
        RECT 28.460 15.325 28.610 15.495 ;
        RECT 31.360 15.325 31.510 15.495 ;
        RECT 34.260 15.325 34.410 15.495 ;
      LAYER met2 ;
        RECT -0.275 15.325 34.760 15.495 ;
    END
  END RWL0_11
  PIN RWL1_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 15.325 0.330 15.495 ;
        RECT 3.080 15.325 3.230 15.495 ;
        RECT 5.980 15.325 6.130 15.495 ;
        RECT 8.880 15.325 9.030 15.495 ;
        RECT 11.780 15.325 11.930 15.495 ;
        RECT 14.680 15.325 14.830 15.495 ;
        RECT 17.580 15.325 17.730 15.495 ;
        RECT 20.480 15.325 20.630 15.495 ;
        RECT 23.380 15.325 23.530 15.495 ;
        RECT 26.280 15.325 26.430 15.495 ;
        RECT 29.180 15.325 29.330 15.495 ;
        RECT 32.080 15.325 32.230 15.495 ;
      LAYER met1 ;
        POLYGON 2.310 15.795 2.310 15.625 2.140 15.625 ;
        RECT 2.310 15.625 2.560 15.795 ;
        POLYGON 2.560 15.795 2.730 15.625 2.560 15.625 ;
        POLYGON 5.210 15.795 5.210 15.625 5.040 15.625 ;
        RECT 5.210 15.625 5.460 15.795 ;
        POLYGON 5.460 15.795 5.630 15.625 5.460 15.625 ;
        POLYGON 8.110 15.795 8.110 15.625 7.940 15.625 ;
        RECT 8.110 15.625 8.360 15.795 ;
        POLYGON 8.360 15.795 8.530 15.625 8.360 15.625 ;
        POLYGON 11.010 15.795 11.010 15.625 10.840 15.625 ;
        RECT 11.010 15.625 11.260 15.795 ;
        POLYGON 11.260 15.795 11.430 15.625 11.260 15.625 ;
        POLYGON 13.910 15.795 13.910 15.625 13.740 15.625 ;
        RECT 13.910 15.625 14.160 15.795 ;
        POLYGON 14.160 15.795 14.330 15.625 14.160 15.625 ;
        POLYGON 16.810 15.795 16.810 15.625 16.640 15.625 ;
        RECT 16.810 15.625 17.060 15.795 ;
        POLYGON 17.060 15.795 17.230 15.625 17.060 15.625 ;
        POLYGON 19.710 15.795 19.710 15.625 19.540 15.625 ;
        RECT 19.710 15.625 19.960 15.795 ;
        POLYGON 19.960 15.795 20.130 15.625 19.960 15.625 ;
        POLYGON 22.610 15.795 22.610 15.625 22.440 15.625 ;
        RECT 22.610 15.625 22.860 15.795 ;
        POLYGON 22.860 15.795 23.030 15.625 22.860 15.625 ;
        POLYGON 25.510 15.795 25.510 15.625 25.340 15.625 ;
        RECT 25.510 15.625 25.760 15.795 ;
        POLYGON 25.760 15.795 25.930 15.625 25.760 15.625 ;
        POLYGON 28.410 15.795 28.410 15.625 28.240 15.625 ;
        RECT 28.410 15.625 28.660 15.795 ;
        POLYGON 28.660 15.795 28.830 15.625 28.660 15.625 ;
        POLYGON 31.310 15.795 31.310 15.625 31.140 15.625 ;
        RECT 31.310 15.625 31.560 15.795 ;
        POLYGON 31.560 15.795 31.730 15.625 31.560 15.625 ;
        POLYGON 34.210 15.795 34.210 15.625 34.040 15.625 ;
        RECT 34.210 15.625 34.460 15.795 ;
        POLYGON 34.460 15.795 34.630 15.625 34.460 15.625 ;
        POLYGON 2.140 15.625 2.140 15.495 2.010 15.495 ;
        RECT 2.140 15.495 2.230 15.625 ;
        POLYGON 2.230 15.625 2.360 15.625 2.230 15.495 ;
        POLYGON 2.510 15.625 2.640 15.625 2.640 15.495 ;
        RECT 2.640 15.495 2.730 15.625 ;
        POLYGON 2.730 15.625 2.860 15.495 2.730 15.495 ;
        POLYGON 5.040 15.625 5.040 15.495 4.910 15.495 ;
        RECT 5.040 15.495 5.130 15.625 ;
        POLYGON 5.130 15.625 5.260 15.625 5.130 15.495 ;
        POLYGON 5.410 15.625 5.540 15.625 5.540 15.495 ;
        RECT 5.540 15.495 5.630 15.625 ;
        POLYGON 5.630 15.625 5.760 15.495 5.630 15.495 ;
        POLYGON 7.940 15.625 7.940 15.495 7.810 15.495 ;
        RECT 7.940 15.495 8.030 15.625 ;
        POLYGON 8.030 15.625 8.160 15.625 8.030 15.495 ;
        POLYGON 8.310 15.625 8.440 15.625 8.440 15.495 ;
        RECT 8.440 15.495 8.530 15.625 ;
        POLYGON 8.530 15.625 8.660 15.495 8.530 15.495 ;
        POLYGON 10.840 15.625 10.840 15.495 10.710 15.495 ;
        RECT 10.840 15.495 10.930 15.625 ;
        POLYGON 10.930 15.625 11.060 15.625 10.930 15.495 ;
        POLYGON 11.210 15.625 11.340 15.625 11.340 15.495 ;
        RECT 11.340 15.495 11.430 15.625 ;
        POLYGON 11.430 15.625 11.560 15.495 11.430 15.495 ;
        POLYGON 13.740 15.625 13.740 15.495 13.610 15.495 ;
        RECT 13.740 15.495 13.830 15.625 ;
        POLYGON 13.830 15.625 13.960 15.625 13.830 15.495 ;
        POLYGON 14.110 15.625 14.240 15.625 14.240 15.495 ;
        RECT 14.240 15.495 14.330 15.625 ;
        POLYGON 14.330 15.625 14.460 15.495 14.330 15.495 ;
        POLYGON 16.640 15.625 16.640 15.495 16.510 15.495 ;
        RECT 16.640 15.495 16.730 15.625 ;
        POLYGON 16.730 15.625 16.860 15.625 16.730 15.495 ;
        POLYGON 17.010 15.625 17.140 15.625 17.140 15.495 ;
        RECT 17.140 15.495 17.230 15.625 ;
        POLYGON 17.230 15.625 17.360 15.495 17.230 15.495 ;
        POLYGON 19.540 15.625 19.540 15.495 19.410 15.495 ;
        RECT 19.540 15.495 19.630 15.625 ;
        POLYGON 19.630 15.625 19.760 15.625 19.630 15.495 ;
        POLYGON 19.910 15.625 20.040 15.625 20.040 15.495 ;
        RECT 20.040 15.495 20.130 15.625 ;
        POLYGON 20.130 15.625 20.260 15.495 20.130 15.495 ;
        POLYGON 22.440 15.625 22.440 15.495 22.310 15.495 ;
        RECT 22.440 15.495 22.530 15.625 ;
        POLYGON 22.530 15.625 22.660 15.625 22.530 15.495 ;
        POLYGON 22.810 15.625 22.940 15.625 22.940 15.495 ;
        RECT 22.940 15.495 23.030 15.625 ;
        POLYGON 23.030 15.625 23.160 15.495 23.030 15.495 ;
        POLYGON 25.340 15.625 25.340 15.495 25.210 15.495 ;
        RECT 25.340 15.495 25.430 15.625 ;
        POLYGON 25.430 15.625 25.560 15.625 25.430 15.495 ;
        POLYGON 25.710 15.625 25.840 15.625 25.840 15.495 ;
        RECT 25.840 15.495 25.930 15.625 ;
        POLYGON 25.930 15.625 26.060 15.495 25.930 15.495 ;
        POLYGON 28.240 15.625 28.240 15.495 28.110 15.495 ;
        RECT 28.240 15.495 28.330 15.625 ;
        POLYGON 28.330 15.625 28.460 15.625 28.330 15.495 ;
        POLYGON 28.610 15.625 28.740 15.625 28.740 15.495 ;
        RECT 28.740 15.495 28.830 15.625 ;
        POLYGON 28.830 15.625 28.960 15.495 28.830 15.495 ;
        POLYGON 31.140 15.625 31.140 15.495 31.010 15.495 ;
        RECT 31.140 15.495 31.230 15.625 ;
        POLYGON 31.230 15.625 31.360 15.625 31.230 15.495 ;
        POLYGON 31.510 15.625 31.640 15.625 31.640 15.495 ;
        RECT 31.640 15.495 31.730 15.625 ;
        POLYGON 31.730 15.625 31.860 15.495 31.730 15.495 ;
        POLYGON 34.040 15.625 34.040 15.495 33.910 15.495 ;
        RECT 34.040 15.495 34.130 15.625 ;
        POLYGON 34.130 15.625 34.260 15.625 34.130 15.495 ;
        POLYGON 34.410 15.625 34.540 15.625 34.540 15.495 ;
        RECT 34.540 15.495 34.630 15.625 ;
        POLYGON 34.630 15.625 34.760 15.495 34.630 15.495 ;
        RECT -0.275 15.325 2.060 15.495 ;
        POLYGON 2.060 15.495 2.230 15.495 2.060 15.325 ;
        POLYGON 2.640 15.495 2.810 15.495 2.810 15.325 ;
        RECT 2.810 15.325 4.960 15.495 ;
        POLYGON 4.960 15.495 5.130 15.495 4.960 15.325 ;
        RECT 5.525 15.325 7.860 15.495 ;
        POLYGON 7.860 15.495 8.030 15.495 7.860 15.325 ;
        POLYGON 8.440 15.495 8.610 15.495 8.610 15.325 ;
        RECT 8.610 15.325 10.760 15.495 ;
        POLYGON 10.760 15.495 10.930 15.495 10.760 15.325 ;
        RECT 11.325 15.325 13.660 15.495 ;
        POLYGON 13.660 15.495 13.830 15.495 13.660 15.325 ;
        POLYGON 14.240 15.495 14.410 15.495 14.410 15.325 ;
        RECT 14.410 15.325 16.560 15.495 ;
        POLYGON 16.560 15.495 16.730 15.495 16.560 15.325 ;
        RECT 17.125 15.325 19.460 15.495 ;
        POLYGON 19.460 15.495 19.630 15.495 19.460 15.325 ;
        POLYGON 20.040 15.495 20.210 15.495 20.210 15.325 ;
        RECT 20.210 15.325 22.360 15.495 ;
        POLYGON 22.360 15.495 22.530 15.495 22.360 15.325 ;
        RECT 22.925 15.325 25.260 15.495 ;
        POLYGON 25.260 15.495 25.430 15.495 25.260 15.325 ;
        POLYGON 25.840 15.495 26.010 15.495 26.010 15.325 ;
        RECT 26.010 15.325 28.160 15.495 ;
        POLYGON 28.160 15.495 28.330 15.495 28.160 15.325 ;
        RECT 28.725 15.325 31.060 15.495 ;
        POLYGON 31.060 15.495 31.230 15.495 31.060 15.325 ;
        POLYGON 31.640 15.495 31.810 15.495 31.810 15.325 ;
        RECT 31.810 15.325 33.960 15.495 ;
        POLYGON 33.960 15.495 34.130 15.495 33.960 15.325 ;
        POLYGON 34.540 15.495 34.710 15.495 34.710 15.325 ;
        RECT 34.710 15.325 34.760 15.495 ;
    END
  END RWL1_11
  PIN RWL0_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 16.675 2.510 16.845 ;
        RECT 5.260 16.675 5.410 16.845 ;
        RECT 8.160 16.675 8.310 16.845 ;
        RECT 11.060 16.675 11.210 16.845 ;
        RECT 13.960 16.675 14.110 16.845 ;
        RECT 16.860 16.675 17.010 16.845 ;
        RECT 19.760 16.675 19.910 16.845 ;
        RECT 22.660 16.675 22.810 16.845 ;
        RECT 25.560 16.675 25.710 16.845 ;
        RECT 28.460 16.675 28.610 16.845 ;
        RECT 31.360 16.675 31.510 16.845 ;
        RECT 34.260 16.675 34.410 16.845 ;
      LAYER mcon ;
        RECT 2.360 16.680 2.510 16.845 ;
        RECT 8.160 16.680 8.310 16.845 ;
        RECT 13.960 16.680 14.110 16.845 ;
        RECT 19.760 16.680 19.910 16.845 ;
        RECT 25.560 16.680 25.710 16.845 ;
        RECT 31.360 16.680 31.510 16.845 ;
      LAYER met1 ;
        RECT 2.360 16.675 2.510 16.845 ;
        RECT 5.260 16.675 5.410 16.845 ;
        RECT 8.160 16.675 8.310 16.845 ;
        RECT 11.060 16.675 11.210 16.845 ;
        RECT 13.960 16.675 14.110 16.845 ;
        RECT 16.860 16.675 17.010 16.845 ;
        RECT 19.760 16.675 19.910 16.845 ;
        RECT 22.660 16.675 22.810 16.845 ;
        RECT 25.560 16.675 25.710 16.845 ;
        RECT 28.460 16.675 28.610 16.845 ;
        RECT 31.360 16.675 31.510 16.845 ;
        RECT 34.260 16.675 34.410 16.845 ;
      LAYER met2 ;
        RECT -0.275 16.675 34.760 16.845 ;
    END
  END RWL0_12
  PIN RWL1_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 16.675 0.330 16.845 ;
        RECT 3.080 16.675 3.230 16.845 ;
        RECT 5.980 16.675 6.130 16.845 ;
        RECT 8.880 16.675 9.030 16.845 ;
        RECT 11.780 16.675 11.930 16.845 ;
        RECT 14.680 16.675 14.830 16.845 ;
        RECT 17.580 16.675 17.730 16.845 ;
        RECT 20.480 16.675 20.630 16.845 ;
        RECT 23.380 16.675 23.530 16.845 ;
        RECT 26.280 16.675 26.430 16.845 ;
        RECT 29.180 16.675 29.330 16.845 ;
        RECT 32.080 16.675 32.230 16.845 ;
      LAYER met1 ;
        POLYGON 2.310 17.145 2.310 16.975 2.140 16.975 ;
        RECT 2.310 16.975 2.560 17.145 ;
        POLYGON 2.560 17.145 2.730 16.975 2.560 16.975 ;
        POLYGON 5.210 17.145 5.210 16.975 5.040 16.975 ;
        RECT 5.210 16.975 5.460 17.145 ;
        POLYGON 5.460 17.145 5.630 16.975 5.460 16.975 ;
        POLYGON 8.110 17.145 8.110 16.975 7.940 16.975 ;
        RECT 8.110 16.975 8.360 17.145 ;
        POLYGON 8.360 17.145 8.530 16.975 8.360 16.975 ;
        POLYGON 11.010 17.145 11.010 16.975 10.840 16.975 ;
        RECT 11.010 16.975 11.260 17.145 ;
        POLYGON 11.260 17.145 11.430 16.975 11.260 16.975 ;
        POLYGON 13.910 17.145 13.910 16.975 13.740 16.975 ;
        RECT 13.910 16.975 14.160 17.145 ;
        POLYGON 14.160 17.145 14.330 16.975 14.160 16.975 ;
        POLYGON 16.810 17.145 16.810 16.975 16.640 16.975 ;
        RECT 16.810 16.975 17.060 17.145 ;
        POLYGON 17.060 17.145 17.230 16.975 17.060 16.975 ;
        POLYGON 19.710 17.145 19.710 16.975 19.540 16.975 ;
        RECT 19.710 16.975 19.960 17.145 ;
        POLYGON 19.960 17.145 20.130 16.975 19.960 16.975 ;
        POLYGON 22.610 17.145 22.610 16.975 22.440 16.975 ;
        RECT 22.610 16.975 22.860 17.145 ;
        POLYGON 22.860 17.145 23.030 16.975 22.860 16.975 ;
        POLYGON 25.510 17.145 25.510 16.975 25.340 16.975 ;
        RECT 25.510 16.975 25.760 17.145 ;
        POLYGON 25.760 17.145 25.930 16.975 25.760 16.975 ;
        POLYGON 28.410 17.145 28.410 16.975 28.240 16.975 ;
        RECT 28.410 16.975 28.660 17.145 ;
        POLYGON 28.660 17.145 28.830 16.975 28.660 16.975 ;
        POLYGON 31.310 17.145 31.310 16.975 31.140 16.975 ;
        RECT 31.310 16.975 31.560 17.145 ;
        POLYGON 31.560 17.145 31.730 16.975 31.560 16.975 ;
        POLYGON 34.210 17.145 34.210 16.975 34.040 16.975 ;
        RECT 34.210 16.975 34.460 17.145 ;
        POLYGON 34.460 17.145 34.630 16.975 34.460 16.975 ;
        POLYGON 2.140 16.975 2.140 16.845 2.010 16.845 ;
        RECT 2.140 16.845 2.230 16.975 ;
        POLYGON 2.230 16.975 2.360 16.975 2.230 16.845 ;
        POLYGON 2.510 16.975 2.640 16.975 2.640 16.845 ;
        RECT 2.640 16.845 2.730 16.975 ;
        POLYGON 2.730 16.975 2.860 16.845 2.730 16.845 ;
        POLYGON 5.040 16.975 5.040 16.845 4.910 16.845 ;
        RECT 5.040 16.845 5.130 16.975 ;
        POLYGON 5.130 16.975 5.260 16.975 5.130 16.845 ;
        POLYGON 5.410 16.975 5.540 16.975 5.540 16.845 ;
        RECT 5.540 16.845 5.630 16.975 ;
        POLYGON 5.630 16.975 5.760 16.845 5.630 16.845 ;
        POLYGON 7.940 16.975 7.940 16.845 7.810 16.845 ;
        RECT 7.940 16.845 8.030 16.975 ;
        POLYGON 8.030 16.975 8.160 16.975 8.030 16.845 ;
        POLYGON 8.310 16.975 8.440 16.975 8.440 16.845 ;
        RECT 8.440 16.845 8.530 16.975 ;
        POLYGON 8.530 16.975 8.660 16.845 8.530 16.845 ;
        POLYGON 10.840 16.975 10.840 16.845 10.710 16.845 ;
        RECT 10.840 16.845 10.930 16.975 ;
        POLYGON 10.930 16.975 11.060 16.975 10.930 16.845 ;
        POLYGON 11.210 16.975 11.340 16.975 11.340 16.845 ;
        RECT 11.340 16.845 11.430 16.975 ;
        POLYGON 11.430 16.975 11.560 16.845 11.430 16.845 ;
        POLYGON 13.740 16.975 13.740 16.845 13.610 16.845 ;
        RECT 13.740 16.845 13.830 16.975 ;
        POLYGON 13.830 16.975 13.960 16.975 13.830 16.845 ;
        POLYGON 14.110 16.975 14.240 16.975 14.240 16.845 ;
        RECT 14.240 16.845 14.330 16.975 ;
        POLYGON 14.330 16.975 14.460 16.845 14.330 16.845 ;
        POLYGON 16.640 16.975 16.640 16.845 16.510 16.845 ;
        RECT 16.640 16.845 16.730 16.975 ;
        POLYGON 16.730 16.975 16.860 16.975 16.730 16.845 ;
        POLYGON 17.010 16.975 17.140 16.975 17.140 16.845 ;
        RECT 17.140 16.845 17.230 16.975 ;
        POLYGON 17.230 16.975 17.360 16.845 17.230 16.845 ;
        POLYGON 19.540 16.975 19.540 16.845 19.410 16.845 ;
        RECT 19.540 16.845 19.630 16.975 ;
        POLYGON 19.630 16.975 19.760 16.975 19.630 16.845 ;
        POLYGON 19.910 16.975 20.040 16.975 20.040 16.845 ;
        RECT 20.040 16.845 20.130 16.975 ;
        POLYGON 20.130 16.975 20.260 16.845 20.130 16.845 ;
        POLYGON 22.440 16.975 22.440 16.845 22.310 16.845 ;
        RECT 22.440 16.845 22.530 16.975 ;
        POLYGON 22.530 16.975 22.660 16.975 22.530 16.845 ;
        POLYGON 22.810 16.975 22.940 16.975 22.940 16.845 ;
        RECT 22.940 16.845 23.030 16.975 ;
        POLYGON 23.030 16.975 23.160 16.845 23.030 16.845 ;
        POLYGON 25.340 16.975 25.340 16.845 25.210 16.845 ;
        RECT 25.340 16.845 25.430 16.975 ;
        POLYGON 25.430 16.975 25.560 16.975 25.430 16.845 ;
        POLYGON 25.710 16.975 25.840 16.975 25.840 16.845 ;
        RECT 25.840 16.845 25.930 16.975 ;
        POLYGON 25.930 16.975 26.060 16.845 25.930 16.845 ;
        POLYGON 28.240 16.975 28.240 16.845 28.110 16.845 ;
        RECT 28.240 16.845 28.330 16.975 ;
        POLYGON 28.330 16.975 28.460 16.975 28.330 16.845 ;
        POLYGON 28.610 16.975 28.740 16.975 28.740 16.845 ;
        RECT 28.740 16.845 28.830 16.975 ;
        POLYGON 28.830 16.975 28.960 16.845 28.830 16.845 ;
        POLYGON 31.140 16.975 31.140 16.845 31.010 16.845 ;
        RECT 31.140 16.845 31.230 16.975 ;
        POLYGON 31.230 16.975 31.360 16.975 31.230 16.845 ;
        POLYGON 31.510 16.975 31.640 16.975 31.640 16.845 ;
        RECT 31.640 16.845 31.730 16.975 ;
        POLYGON 31.730 16.975 31.860 16.845 31.730 16.845 ;
        POLYGON 34.040 16.975 34.040 16.845 33.910 16.845 ;
        RECT 34.040 16.845 34.130 16.975 ;
        POLYGON 34.130 16.975 34.260 16.975 34.130 16.845 ;
        POLYGON 34.410 16.975 34.540 16.975 34.540 16.845 ;
        RECT 34.540 16.845 34.630 16.975 ;
        POLYGON 34.630 16.975 34.760 16.845 34.630 16.845 ;
        RECT -0.275 16.675 2.060 16.845 ;
        POLYGON 2.060 16.845 2.230 16.845 2.060 16.675 ;
        POLYGON 2.640 16.845 2.810 16.845 2.810 16.675 ;
        RECT 2.810 16.675 4.960 16.845 ;
        POLYGON 4.960 16.845 5.130 16.845 4.960 16.675 ;
        RECT 5.525 16.675 7.860 16.845 ;
        POLYGON 7.860 16.845 8.030 16.845 7.860 16.675 ;
        POLYGON 8.440 16.845 8.610 16.845 8.610 16.675 ;
        RECT 8.610 16.675 10.760 16.845 ;
        POLYGON 10.760 16.845 10.930 16.845 10.760 16.675 ;
        RECT 11.325 16.675 13.660 16.845 ;
        POLYGON 13.660 16.845 13.830 16.845 13.660 16.675 ;
        POLYGON 14.240 16.845 14.410 16.845 14.410 16.675 ;
        RECT 14.410 16.675 16.560 16.845 ;
        POLYGON 16.560 16.845 16.730 16.845 16.560 16.675 ;
        RECT 17.125 16.675 19.460 16.845 ;
        POLYGON 19.460 16.845 19.630 16.845 19.460 16.675 ;
        POLYGON 20.040 16.845 20.210 16.845 20.210 16.675 ;
        RECT 20.210 16.675 22.360 16.845 ;
        POLYGON 22.360 16.845 22.530 16.845 22.360 16.675 ;
        RECT 22.925 16.675 25.260 16.845 ;
        POLYGON 25.260 16.845 25.430 16.845 25.260 16.675 ;
        POLYGON 25.840 16.845 26.010 16.845 26.010 16.675 ;
        RECT 26.010 16.675 28.160 16.845 ;
        POLYGON 28.160 16.845 28.330 16.845 28.160 16.675 ;
        RECT 28.725 16.675 31.060 16.845 ;
        POLYGON 31.060 16.845 31.230 16.845 31.060 16.675 ;
        POLYGON 31.640 16.845 31.810 16.845 31.810 16.675 ;
        RECT 31.810 16.675 33.960 16.845 ;
        POLYGON 33.960 16.845 34.130 16.845 33.960 16.675 ;
        POLYGON 34.540 16.845 34.710 16.845 34.710 16.675 ;
        RECT 34.710 16.675 34.760 16.845 ;
    END
  END RWL1_12
  PIN RWL0_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 18.025 2.510 18.195 ;
        RECT 5.260 18.025 5.410 18.195 ;
        RECT 8.160 18.025 8.310 18.195 ;
        RECT 11.060 18.025 11.210 18.195 ;
        RECT 13.960 18.025 14.110 18.195 ;
        RECT 16.860 18.025 17.010 18.195 ;
        RECT 19.760 18.025 19.910 18.195 ;
        RECT 22.660 18.025 22.810 18.195 ;
        RECT 25.560 18.025 25.710 18.195 ;
        RECT 28.460 18.025 28.610 18.195 ;
        RECT 31.360 18.025 31.510 18.195 ;
        RECT 34.260 18.025 34.410 18.195 ;
      LAYER mcon ;
        RECT 2.360 18.030 2.510 18.195 ;
        RECT 8.160 18.030 8.310 18.195 ;
        RECT 13.960 18.030 14.110 18.195 ;
        RECT 19.760 18.030 19.910 18.195 ;
        RECT 25.560 18.030 25.710 18.195 ;
        RECT 31.360 18.030 31.510 18.195 ;
      LAYER met1 ;
        RECT 2.360 18.025 2.510 18.195 ;
        RECT 5.260 18.025 5.410 18.195 ;
        RECT 8.160 18.025 8.310 18.195 ;
        RECT 11.060 18.025 11.210 18.195 ;
        RECT 13.960 18.025 14.110 18.195 ;
        RECT 16.860 18.025 17.010 18.195 ;
        RECT 19.760 18.025 19.910 18.195 ;
        RECT 22.660 18.025 22.810 18.195 ;
        RECT 25.560 18.025 25.710 18.195 ;
        RECT 28.460 18.025 28.610 18.195 ;
        RECT 31.360 18.025 31.510 18.195 ;
        RECT 34.260 18.025 34.410 18.195 ;
      LAYER met2 ;
        RECT -0.275 18.025 34.760 18.195 ;
    END
  END RWL0_13
  PIN RWL1_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 18.025 0.330 18.195 ;
        RECT 3.080 18.025 3.230 18.195 ;
        RECT 5.980 18.025 6.130 18.195 ;
        RECT 8.880 18.025 9.030 18.195 ;
        RECT 11.780 18.025 11.930 18.195 ;
        RECT 14.680 18.025 14.830 18.195 ;
        RECT 17.580 18.025 17.730 18.195 ;
        RECT 20.480 18.025 20.630 18.195 ;
        RECT 23.380 18.025 23.530 18.195 ;
        RECT 26.280 18.025 26.430 18.195 ;
        RECT 29.180 18.025 29.330 18.195 ;
        RECT 32.080 18.025 32.230 18.195 ;
      LAYER met1 ;
        POLYGON 2.310 18.495 2.310 18.325 2.140 18.325 ;
        RECT 2.310 18.325 2.560 18.495 ;
        POLYGON 2.560 18.495 2.730 18.325 2.560 18.325 ;
        POLYGON 5.210 18.495 5.210 18.325 5.040 18.325 ;
        RECT 5.210 18.325 5.460 18.495 ;
        POLYGON 5.460 18.495 5.630 18.325 5.460 18.325 ;
        POLYGON 8.110 18.495 8.110 18.325 7.940 18.325 ;
        RECT 8.110 18.325 8.360 18.495 ;
        POLYGON 8.360 18.495 8.530 18.325 8.360 18.325 ;
        POLYGON 11.010 18.495 11.010 18.325 10.840 18.325 ;
        RECT 11.010 18.325 11.260 18.495 ;
        POLYGON 11.260 18.495 11.430 18.325 11.260 18.325 ;
        POLYGON 13.910 18.495 13.910 18.325 13.740 18.325 ;
        RECT 13.910 18.325 14.160 18.495 ;
        POLYGON 14.160 18.495 14.330 18.325 14.160 18.325 ;
        POLYGON 16.810 18.495 16.810 18.325 16.640 18.325 ;
        RECT 16.810 18.325 17.060 18.495 ;
        POLYGON 17.060 18.495 17.230 18.325 17.060 18.325 ;
        POLYGON 19.710 18.495 19.710 18.325 19.540 18.325 ;
        RECT 19.710 18.325 19.960 18.495 ;
        POLYGON 19.960 18.495 20.130 18.325 19.960 18.325 ;
        POLYGON 22.610 18.495 22.610 18.325 22.440 18.325 ;
        RECT 22.610 18.325 22.860 18.495 ;
        POLYGON 22.860 18.495 23.030 18.325 22.860 18.325 ;
        POLYGON 25.510 18.495 25.510 18.325 25.340 18.325 ;
        RECT 25.510 18.325 25.760 18.495 ;
        POLYGON 25.760 18.495 25.930 18.325 25.760 18.325 ;
        POLYGON 28.410 18.495 28.410 18.325 28.240 18.325 ;
        RECT 28.410 18.325 28.660 18.495 ;
        POLYGON 28.660 18.495 28.830 18.325 28.660 18.325 ;
        POLYGON 31.310 18.495 31.310 18.325 31.140 18.325 ;
        RECT 31.310 18.325 31.560 18.495 ;
        POLYGON 31.560 18.495 31.730 18.325 31.560 18.325 ;
        POLYGON 34.210 18.495 34.210 18.325 34.040 18.325 ;
        RECT 34.210 18.325 34.460 18.495 ;
        POLYGON 34.460 18.495 34.630 18.325 34.460 18.325 ;
        POLYGON 2.140 18.325 2.140 18.195 2.010 18.195 ;
        RECT 2.140 18.195 2.230 18.325 ;
        POLYGON 2.230 18.325 2.360 18.325 2.230 18.195 ;
        POLYGON 2.510 18.325 2.640 18.325 2.640 18.195 ;
        RECT 2.640 18.195 2.730 18.325 ;
        POLYGON 2.730 18.325 2.860 18.195 2.730 18.195 ;
        POLYGON 5.040 18.325 5.040 18.195 4.910 18.195 ;
        RECT 5.040 18.195 5.130 18.325 ;
        POLYGON 5.130 18.325 5.260 18.325 5.130 18.195 ;
        POLYGON 5.410 18.325 5.540 18.325 5.540 18.195 ;
        RECT 5.540 18.195 5.630 18.325 ;
        POLYGON 5.630 18.325 5.760 18.195 5.630 18.195 ;
        POLYGON 7.940 18.325 7.940 18.195 7.810 18.195 ;
        RECT 7.940 18.195 8.030 18.325 ;
        POLYGON 8.030 18.325 8.160 18.325 8.030 18.195 ;
        POLYGON 8.310 18.325 8.440 18.325 8.440 18.195 ;
        RECT 8.440 18.195 8.530 18.325 ;
        POLYGON 8.530 18.325 8.660 18.195 8.530 18.195 ;
        POLYGON 10.840 18.325 10.840 18.195 10.710 18.195 ;
        RECT 10.840 18.195 10.930 18.325 ;
        POLYGON 10.930 18.325 11.060 18.325 10.930 18.195 ;
        POLYGON 11.210 18.325 11.340 18.325 11.340 18.195 ;
        RECT 11.340 18.195 11.430 18.325 ;
        POLYGON 11.430 18.325 11.560 18.195 11.430 18.195 ;
        POLYGON 13.740 18.325 13.740 18.195 13.610 18.195 ;
        RECT 13.740 18.195 13.830 18.325 ;
        POLYGON 13.830 18.325 13.960 18.325 13.830 18.195 ;
        POLYGON 14.110 18.325 14.240 18.325 14.240 18.195 ;
        RECT 14.240 18.195 14.330 18.325 ;
        POLYGON 14.330 18.325 14.460 18.195 14.330 18.195 ;
        POLYGON 16.640 18.325 16.640 18.195 16.510 18.195 ;
        RECT 16.640 18.195 16.730 18.325 ;
        POLYGON 16.730 18.325 16.860 18.325 16.730 18.195 ;
        POLYGON 17.010 18.325 17.140 18.325 17.140 18.195 ;
        RECT 17.140 18.195 17.230 18.325 ;
        POLYGON 17.230 18.325 17.360 18.195 17.230 18.195 ;
        POLYGON 19.540 18.325 19.540 18.195 19.410 18.195 ;
        RECT 19.540 18.195 19.630 18.325 ;
        POLYGON 19.630 18.325 19.760 18.325 19.630 18.195 ;
        POLYGON 19.910 18.325 20.040 18.325 20.040 18.195 ;
        RECT 20.040 18.195 20.130 18.325 ;
        POLYGON 20.130 18.325 20.260 18.195 20.130 18.195 ;
        POLYGON 22.440 18.325 22.440 18.195 22.310 18.195 ;
        RECT 22.440 18.195 22.530 18.325 ;
        POLYGON 22.530 18.325 22.660 18.325 22.530 18.195 ;
        POLYGON 22.810 18.325 22.940 18.325 22.940 18.195 ;
        RECT 22.940 18.195 23.030 18.325 ;
        POLYGON 23.030 18.325 23.160 18.195 23.030 18.195 ;
        POLYGON 25.340 18.325 25.340 18.195 25.210 18.195 ;
        RECT 25.340 18.195 25.430 18.325 ;
        POLYGON 25.430 18.325 25.560 18.325 25.430 18.195 ;
        POLYGON 25.710 18.325 25.840 18.325 25.840 18.195 ;
        RECT 25.840 18.195 25.930 18.325 ;
        POLYGON 25.930 18.325 26.060 18.195 25.930 18.195 ;
        POLYGON 28.240 18.325 28.240 18.195 28.110 18.195 ;
        RECT 28.240 18.195 28.330 18.325 ;
        POLYGON 28.330 18.325 28.460 18.325 28.330 18.195 ;
        POLYGON 28.610 18.325 28.740 18.325 28.740 18.195 ;
        RECT 28.740 18.195 28.830 18.325 ;
        POLYGON 28.830 18.325 28.960 18.195 28.830 18.195 ;
        POLYGON 31.140 18.325 31.140 18.195 31.010 18.195 ;
        RECT 31.140 18.195 31.230 18.325 ;
        POLYGON 31.230 18.325 31.360 18.325 31.230 18.195 ;
        POLYGON 31.510 18.325 31.640 18.325 31.640 18.195 ;
        RECT 31.640 18.195 31.730 18.325 ;
        POLYGON 31.730 18.325 31.860 18.195 31.730 18.195 ;
        POLYGON 34.040 18.325 34.040 18.195 33.910 18.195 ;
        RECT 34.040 18.195 34.130 18.325 ;
        POLYGON 34.130 18.325 34.260 18.325 34.130 18.195 ;
        POLYGON 34.410 18.325 34.540 18.325 34.540 18.195 ;
        RECT 34.540 18.195 34.630 18.325 ;
        POLYGON 34.630 18.325 34.760 18.195 34.630 18.195 ;
        RECT -0.275 18.025 2.060 18.195 ;
        POLYGON 2.060 18.195 2.230 18.195 2.060 18.025 ;
        POLYGON 2.640 18.195 2.810 18.195 2.810 18.025 ;
        RECT 2.810 18.025 4.960 18.195 ;
        POLYGON 4.960 18.195 5.130 18.195 4.960 18.025 ;
        RECT 5.525 18.025 7.860 18.195 ;
        POLYGON 7.860 18.195 8.030 18.195 7.860 18.025 ;
        POLYGON 8.440 18.195 8.610 18.195 8.610 18.025 ;
        RECT 8.610 18.025 10.760 18.195 ;
        POLYGON 10.760 18.195 10.930 18.195 10.760 18.025 ;
        RECT 11.325 18.025 13.660 18.195 ;
        POLYGON 13.660 18.195 13.830 18.195 13.660 18.025 ;
        POLYGON 14.240 18.195 14.410 18.195 14.410 18.025 ;
        RECT 14.410 18.025 16.560 18.195 ;
        POLYGON 16.560 18.195 16.730 18.195 16.560 18.025 ;
        RECT 17.125 18.025 19.460 18.195 ;
        POLYGON 19.460 18.195 19.630 18.195 19.460 18.025 ;
        POLYGON 20.040 18.195 20.210 18.195 20.210 18.025 ;
        RECT 20.210 18.025 22.360 18.195 ;
        POLYGON 22.360 18.195 22.530 18.195 22.360 18.025 ;
        RECT 22.925 18.025 25.260 18.195 ;
        POLYGON 25.260 18.195 25.430 18.195 25.260 18.025 ;
        POLYGON 25.840 18.195 26.010 18.195 26.010 18.025 ;
        RECT 26.010 18.025 28.160 18.195 ;
        POLYGON 28.160 18.195 28.330 18.195 28.160 18.025 ;
        RECT 28.725 18.025 31.060 18.195 ;
        POLYGON 31.060 18.195 31.230 18.195 31.060 18.025 ;
        POLYGON 31.640 18.195 31.810 18.195 31.810 18.025 ;
        RECT 31.810 18.025 33.960 18.195 ;
        POLYGON 33.960 18.195 34.130 18.195 33.960 18.025 ;
        POLYGON 34.540 18.195 34.710 18.195 34.710 18.025 ;
        RECT 34.710 18.025 34.760 18.195 ;
    END
  END RWL1_13
  PIN RWL0_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 19.375 2.510 19.545 ;
        RECT 5.260 19.375 5.410 19.545 ;
        RECT 8.160 19.375 8.310 19.545 ;
        RECT 11.060 19.375 11.210 19.545 ;
        RECT 13.960 19.375 14.110 19.545 ;
        RECT 16.860 19.375 17.010 19.545 ;
        RECT 19.760 19.375 19.910 19.545 ;
        RECT 22.660 19.375 22.810 19.545 ;
        RECT 25.560 19.375 25.710 19.545 ;
        RECT 28.460 19.375 28.610 19.545 ;
        RECT 31.360 19.375 31.510 19.545 ;
        RECT 34.260 19.375 34.410 19.545 ;
      LAYER mcon ;
        RECT 2.360 19.380 2.510 19.545 ;
        RECT 8.160 19.380 8.310 19.545 ;
        RECT 13.960 19.380 14.110 19.545 ;
        RECT 19.760 19.380 19.910 19.545 ;
        RECT 25.560 19.380 25.710 19.545 ;
        RECT 31.360 19.380 31.510 19.545 ;
      LAYER met1 ;
        RECT 2.360 19.375 2.510 19.545 ;
        RECT 5.260 19.375 5.410 19.545 ;
        RECT 8.160 19.375 8.310 19.545 ;
        RECT 11.060 19.375 11.210 19.545 ;
        RECT 13.960 19.375 14.110 19.545 ;
        RECT 16.860 19.375 17.010 19.545 ;
        RECT 19.760 19.375 19.910 19.545 ;
        RECT 22.660 19.375 22.810 19.545 ;
        RECT 25.560 19.375 25.710 19.545 ;
        RECT 28.460 19.375 28.610 19.545 ;
        RECT 31.360 19.375 31.510 19.545 ;
        RECT 34.260 19.375 34.410 19.545 ;
      LAYER met2 ;
        RECT -0.275 19.375 34.760 19.545 ;
    END
  END RWL0_14
  PIN RWL1_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 19.375 0.330 19.545 ;
        RECT 3.080 19.375 3.230 19.545 ;
        RECT 5.980 19.375 6.130 19.545 ;
        RECT 8.880 19.375 9.030 19.545 ;
        RECT 11.780 19.375 11.930 19.545 ;
        RECT 14.680 19.375 14.830 19.545 ;
        RECT 17.580 19.375 17.730 19.545 ;
        RECT 20.480 19.375 20.630 19.545 ;
        RECT 23.380 19.375 23.530 19.545 ;
        RECT 26.280 19.375 26.430 19.545 ;
        RECT 29.180 19.375 29.330 19.545 ;
        RECT 32.080 19.375 32.230 19.545 ;
      LAYER met1 ;
        POLYGON 2.310 19.845 2.310 19.675 2.140 19.675 ;
        RECT 2.310 19.675 2.560 19.845 ;
        POLYGON 2.560 19.845 2.730 19.675 2.560 19.675 ;
        POLYGON 5.210 19.845 5.210 19.675 5.040 19.675 ;
        RECT 5.210 19.675 5.460 19.845 ;
        POLYGON 5.460 19.845 5.630 19.675 5.460 19.675 ;
        POLYGON 8.110 19.845 8.110 19.675 7.940 19.675 ;
        RECT 8.110 19.675 8.360 19.845 ;
        POLYGON 8.360 19.845 8.530 19.675 8.360 19.675 ;
        POLYGON 11.010 19.845 11.010 19.675 10.840 19.675 ;
        RECT 11.010 19.675 11.260 19.845 ;
        POLYGON 11.260 19.845 11.430 19.675 11.260 19.675 ;
        POLYGON 13.910 19.845 13.910 19.675 13.740 19.675 ;
        RECT 13.910 19.675 14.160 19.845 ;
        POLYGON 14.160 19.845 14.330 19.675 14.160 19.675 ;
        POLYGON 16.810 19.845 16.810 19.675 16.640 19.675 ;
        RECT 16.810 19.675 17.060 19.845 ;
        POLYGON 17.060 19.845 17.230 19.675 17.060 19.675 ;
        POLYGON 19.710 19.845 19.710 19.675 19.540 19.675 ;
        RECT 19.710 19.675 19.960 19.845 ;
        POLYGON 19.960 19.845 20.130 19.675 19.960 19.675 ;
        POLYGON 22.610 19.845 22.610 19.675 22.440 19.675 ;
        RECT 22.610 19.675 22.860 19.845 ;
        POLYGON 22.860 19.845 23.030 19.675 22.860 19.675 ;
        POLYGON 25.510 19.845 25.510 19.675 25.340 19.675 ;
        RECT 25.510 19.675 25.760 19.845 ;
        POLYGON 25.760 19.845 25.930 19.675 25.760 19.675 ;
        POLYGON 28.410 19.845 28.410 19.675 28.240 19.675 ;
        RECT 28.410 19.675 28.660 19.845 ;
        POLYGON 28.660 19.845 28.830 19.675 28.660 19.675 ;
        POLYGON 31.310 19.845 31.310 19.675 31.140 19.675 ;
        RECT 31.310 19.675 31.560 19.845 ;
        POLYGON 31.560 19.845 31.730 19.675 31.560 19.675 ;
        POLYGON 34.210 19.845 34.210 19.675 34.040 19.675 ;
        RECT 34.210 19.675 34.460 19.845 ;
        POLYGON 34.460 19.845 34.630 19.675 34.460 19.675 ;
        POLYGON 2.140 19.675 2.140 19.545 2.010 19.545 ;
        RECT 2.140 19.545 2.230 19.675 ;
        POLYGON 2.230 19.675 2.360 19.675 2.230 19.545 ;
        POLYGON 2.510 19.675 2.640 19.675 2.640 19.545 ;
        RECT 2.640 19.545 2.730 19.675 ;
        POLYGON 2.730 19.675 2.860 19.545 2.730 19.545 ;
        POLYGON 5.040 19.675 5.040 19.545 4.910 19.545 ;
        RECT 5.040 19.545 5.130 19.675 ;
        POLYGON 5.130 19.675 5.260 19.675 5.130 19.545 ;
        POLYGON 5.410 19.675 5.540 19.675 5.540 19.545 ;
        RECT 5.540 19.545 5.630 19.675 ;
        POLYGON 5.630 19.675 5.760 19.545 5.630 19.545 ;
        POLYGON 7.940 19.675 7.940 19.545 7.810 19.545 ;
        RECT 7.940 19.545 8.030 19.675 ;
        POLYGON 8.030 19.675 8.160 19.675 8.030 19.545 ;
        POLYGON 8.310 19.675 8.440 19.675 8.440 19.545 ;
        RECT 8.440 19.545 8.530 19.675 ;
        POLYGON 8.530 19.675 8.660 19.545 8.530 19.545 ;
        POLYGON 10.840 19.675 10.840 19.545 10.710 19.545 ;
        RECT 10.840 19.545 10.930 19.675 ;
        POLYGON 10.930 19.675 11.060 19.675 10.930 19.545 ;
        POLYGON 11.210 19.675 11.340 19.675 11.340 19.545 ;
        RECT 11.340 19.545 11.430 19.675 ;
        POLYGON 11.430 19.675 11.560 19.545 11.430 19.545 ;
        POLYGON 13.740 19.675 13.740 19.545 13.610 19.545 ;
        RECT 13.740 19.545 13.830 19.675 ;
        POLYGON 13.830 19.675 13.960 19.675 13.830 19.545 ;
        POLYGON 14.110 19.675 14.240 19.675 14.240 19.545 ;
        RECT 14.240 19.545 14.330 19.675 ;
        POLYGON 14.330 19.675 14.460 19.545 14.330 19.545 ;
        POLYGON 16.640 19.675 16.640 19.545 16.510 19.545 ;
        RECT 16.640 19.545 16.730 19.675 ;
        POLYGON 16.730 19.675 16.860 19.675 16.730 19.545 ;
        POLYGON 17.010 19.675 17.140 19.675 17.140 19.545 ;
        RECT 17.140 19.545 17.230 19.675 ;
        POLYGON 17.230 19.675 17.360 19.545 17.230 19.545 ;
        POLYGON 19.540 19.675 19.540 19.545 19.410 19.545 ;
        RECT 19.540 19.545 19.630 19.675 ;
        POLYGON 19.630 19.675 19.760 19.675 19.630 19.545 ;
        POLYGON 19.910 19.675 20.040 19.675 20.040 19.545 ;
        RECT 20.040 19.545 20.130 19.675 ;
        POLYGON 20.130 19.675 20.260 19.545 20.130 19.545 ;
        POLYGON 22.440 19.675 22.440 19.545 22.310 19.545 ;
        RECT 22.440 19.545 22.530 19.675 ;
        POLYGON 22.530 19.675 22.660 19.675 22.530 19.545 ;
        POLYGON 22.810 19.675 22.940 19.675 22.940 19.545 ;
        RECT 22.940 19.545 23.030 19.675 ;
        POLYGON 23.030 19.675 23.160 19.545 23.030 19.545 ;
        POLYGON 25.340 19.675 25.340 19.545 25.210 19.545 ;
        RECT 25.340 19.545 25.430 19.675 ;
        POLYGON 25.430 19.675 25.560 19.675 25.430 19.545 ;
        POLYGON 25.710 19.675 25.840 19.675 25.840 19.545 ;
        RECT 25.840 19.545 25.930 19.675 ;
        POLYGON 25.930 19.675 26.060 19.545 25.930 19.545 ;
        POLYGON 28.240 19.675 28.240 19.545 28.110 19.545 ;
        RECT 28.240 19.545 28.330 19.675 ;
        POLYGON 28.330 19.675 28.460 19.675 28.330 19.545 ;
        POLYGON 28.610 19.675 28.740 19.675 28.740 19.545 ;
        RECT 28.740 19.545 28.830 19.675 ;
        POLYGON 28.830 19.675 28.960 19.545 28.830 19.545 ;
        POLYGON 31.140 19.675 31.140 19.545 31.010 19.545 ;
        RECT 31.140 19.545 31.230 19.675 ;
        POLYGON 31.230 19.675 31.360 19.675 31.230 19.545 ;
        POLYGON 31.510 19.675 31.640 19.675 31.640 19.545 ;
        RECT 31.640 19.545 31.730 19.675 ;
        POLYGON 31.730 19.675 31.860 19.545 31.730 19.545 ;
        POLYGON 34.040 19.675 34.040 19.545 33.910 19.545 ;
        RECT 34.040 19.545 34.130 19.675 ;
        POLYGON 34.130 19.675 34.260 19.675 34.130 19.545 ;
        POLYGON 34.410 19.675 34.540 19.675 34.540 19.545 ;
        RECT 34.540 19.545 34.630 19.675 ;
        POLYGON 34.630 19.675 34.760 19.545 34.630 19.545 ;
        RECT -0.275 19.375 2.060 19.545 ;
        POLYGON 2.060 19.545 2.230 19.545 2.060 19.375 ;
        POLYGON 2.640 19.545 2.810 19.545 2.810 19.375 ;
        RECT 2.810 19.375 4.960 19.545 ;
        POLYGON 4.960 19.545 5.130 19.545 4.960 19.375 ;
        RECT 5.525 19.375 7.860 19.545 ;
        POLYGON 7.860 19.545 8.030 19.545 7.860 19.375 ;
        POLYGON 8.440 19.545 8.610 19.545 8.610 19.375 ;
        RECT 8.610 19.375 10.760 19.545 ;
        POLYGON 10.760 19.545 10.930 19.545 10.760 19.375 ;
        RECT 11.325 19.375 13.660 19.545 ;
        POLYGON 13.660 19.545 13.830 19.545 13.660 19.375 ;
        POLYGON 14.240 19.545 14.410 19.545 14.410 19.375 ;
        RECT 14.410 19.375 16.560 19.545 ;
        POLYGON 16.560 19.545 16.730 19.545 16.560 19.375 ;
        RECT 17.125 19.375 19.460 19.545 ;
        POLYGON 19.460 19.545 19.630 19.545 19.460 19.375 ;
        POLYGON 20.040 19.545 20.210 19.545 20.210 19.375 ;
        RECT 20.210 19.375 22.360 19.545 ;
        POLYGON 22.360 19.545 22.530 19.545 22.360 19.375 ;
        RECT 22.925 19.375 25.260 19.545 ;
        POLYGON 25.260 19.545 25.430 19.545 25.260 19.375 ;
        POLYGON 25.840 19.545 26.010 19.545 26.010 19.375 ;
        RECT 26.010 19.375 28.160 19.545 ;
        POLYGON 28.160 19.545 28.330 19.545 28.160 19.375 ;
        RECT 28.725 19.375 31.060 19.545 ;
        POLYGON 31.060 19.545 31.230 19.545 31.060 19.375 ;
        POLYGON 31.640 19.545 31.810 19.545 31.810 19.375 ;
        RECT 31.810 19.375 33.960 19.545 ;
        POLYGON 33.960 19.545 34.130 19.545 33.960 19.375 ;
        POLYGON 34.540 19.545 34.710 19.545 34.710 19.375 ;
        RECT 34.710 19.375 34.760 19.545 ;
    END
  END RWL1_14
  PIN RWL0_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 2.360 20.725 2.510 20.895 ;
        RECT 5.260 20.725 5.410 20.895 ;
        RECT 8.160 20.725 8.310 20.895 ;
        RECT 11.060 20.725 11.210 20.895 ;
        RECT 13.960 20.725 14.110 20.895 ;
        RECT 16.860 20.725 17.010 20.895 ;
        RECT 19.760 20.725 19.910 20.895 ;
        RECT 22.660 20.725 22.810 20.895 ;
        RECT 25.560 20.725 25.710 20.895 ;
        RECT 28.460 20.725 28.610 20.895 ;
        RECT 31.360 20.725 31.510 20.895 ;
        RECT 34.260 20.725 34.410 20.895 ;
      LAYER mcon ;
        RECT 8.160 20.730 8.310 20.895 ;
        RECT 13.960 20.730 14.110 20.895 ;
        RECT 19.760 20.730 19.910 20.895 ;
        RECT 25.560 20.730 25.710 20.895 ;
        RECT 31.360 20.730 31.510 20.895 ;
      LAYER met1 ;
        RECT 2.360 20.725 2.510 20.895 ;
        RECT 5.260 20.725 5.410 20.895 ;
        RECT 8.160 20.725 8.310 20.895 ;
        RECT 11.060 20.725 11.210 20.895 ;
        RECT 13.960 20.725 14.110 20.895 ;
        RECT 16.860 20.725 17.010 20.895 ;
        RECT 19.760 20.725 19.910 20.895 ;
        RECT 22.660 20.725 22.810 20.895 ;
        RECT 25.560 20.725 25.710 20.895 ;
        RECT 28.460 20.725 28.610 20.895 ;
        RECT 31.360 20.725 31.510 20.895 ;
        RECT 34.260 20.725 34.410 20.895 ;
      LAYER met2 ;
        RECT -0.275 20.725 34.760 20.895 ;
    END
  END RWL0_15
  PIN RWL1_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 20.725 0.330 20.895 ;
        RECT 3.080 20.725 3.230 20.895 ;
        RECT 5.980 20.725 6.130 20.895 ;
        RECT 8.880 20.725 9.030 20.895 ;
        RECT 11.780 20.725 11.930 20.895 ;
        RECT 14.680 20.725 14.830 20.895 ;
        RECT 17.580 20.725 17.730 20.895 ;
        RECT 20.480 20.725 20.630 20.895 ;
        RECT 23.380 20.725 23.530 20.895 ;
        RECT 26.280 20.725 26.430 20.895 ;
        RECT 29.180 20.725 29.330 20.895 ;
        RECT 32.080 20.725 32.230 20.895 ;
      LAYER met1 ;
        POLYGON 2.310 21.195 2.310 21.025 2.140 21.025 ;
        RECT 2.310 21.025 2.560 21.195 ;
        POLYGON 2.560 21.195 2.730 21.025 2.560 21.025 ;
        POLYGON 5.210 21.195 5.210 21.025 5.040 21.025 ;
        RECT 5.210 21.025 5.460 21.195 ;
        POLYGON 5.460 21.195 5.630 21.025 5.460 21.025 ;
        POLYGON 8.110 21.195 8.110 21.025 7.940 21.025 ;
        RECT 8.110 21.025 8.360 21.195 ;
        POLYGON 8.360 21.195 8.530 21.025 8.360 21.025 ;
        POLYGON 11.010 21.195 11.010 21.025 10.840 21.025 ;
        RECT 11.010 21.025 11.260 21.195 ;
        POLYGON 11.260 21.195 11.430 21.025 11.260 21.025 ;
        POLYGON 13.910 21.195 13.910 21.025 13.740 21.025 ;
        RECT 13.910 21.025 14.160 21.195 ;
        POLYGON 14.160 21.195 14.330 21.025 14.160 21.025 ;
        POLYGON 16.810 21.195 16.810 21.025 16.640 21.025 ;
        RECT 16.810 21.025 17.060 21.195 ;
        POLYGON 17.060 21.195 17.230 21.025 17.060 21.025 ;
        POLYGON 19.710 21.195 19.710 21.025 19.540 21.025 ;
        RECT 19.710 21.025 19.960 21.195 ;
        POLYGON 19.960 21.195 20.130 21.025 19.960 21.025 ;
        POLYGON 22.610 21.195 22.610 21.025 22.440 21.025 ;
        RECT 22.610 21.025 22.860 21.195 ;
        POLYGON 22.860 21.195 23.030 21.025 22.860 21.025 ;
        POLYGON 25.510 21.195 25.510 21.025 25.340 21.025 ;
        RECT 25.510 21.025 25.760 21.195 ;
        POLYGON 25.760 21.195 25.930 21.025 25.760 21.025 ;
        POLYGON 28.410 21.195 28.410 21.025 28.240 21.025 ;
        RECT 28.410 21.025 28.660 21.195 ;
        POLYGON 28.660 21.195 28.830 21.025 28.660 21.025 ;
        POLYGON 31.310 21.195 31.310 21.025 31.140 21.025 ;
        RECT 31.310 21.025 31.560 21.195 ;
        POLYGON 31.560 21.195 31.730 21.025 31.560 21.025 ;
        POLYGON 34.210 21.195 34.210 21.025 34.040 21.025 ;
        RECT 34.210 21.025 34.460 21.195 ;
        POLYGON 34.460 21.195 34.630 21.025 34.460 21.025 ;
        POLYGON 2.140 21.025 2.140 20.895 2.010 20.895 ;
        RECT 2.140 20.895 2.230 21.025 ;
        POLYGON 2.230 21.025 2.360 21.025 2.230 20.895 ;
        POLYGON 2.510 21.025 2.640 21.025 2.640 20.895 ;
        RECT 2.640 20.895 2.730 21.025 ;
        POLYGON 2.730 21.025 2.860 20.895 2.730 20.895 ;
        POLYGON 5.040 21.025 5.040 20.895 4.910 20.895 ;
        RECT 5.040 20.895 5.130 21.025 ;
        POLYGON 5.130 21.025 5.260 21.025 5.130 20.895 ;
        POLYGON 5.410 21.025 5.540 21.025 5.540 20.895 ;
        RECT 5.540 20.895 5.630 21.025 ;
        POLYGON 5.630 21.025 5.760 20.895 5.630 20.895 ;
        POLYGON 7.940 21.025 7.940 20.895 7.810 20.895 ;
        RECT 7.940 20.895 8.030 21.025 ;
        POLYGON 8.030 21.025 8.160 21.025 8.030 20.895 ;
        POLYGON 8.310 21.025 8.440 21.025 8.440 20.895 ;
        RECT 8.440 20.895 8.530 21.025 ;
        POLYGON 8.530 21.025 8.660 20.895 8.530 20.895 ;
        POLYGON 10.840 21.025 10.840 20.895 10.710 20.895 ;
        RECT 10.840 20.895 10.930 21.025 ;
        POLYGON 10.930 21.025 11.060 21.025 10.930 20.895 ;
        POLYGON 11.210 21.025 11.340 21.025 11.340 20.895 ;
        RECT 11.340 20.895 11.430 21.025 ;
        POLYGON 11.430 21.025 11.560 20.895 11.430 20.895 ;
        POLYGON 13.740 21.025 13.740 20.895 13.610 20.895 ;
        RECT 13.740 20.895 13.830 21.025 ;
        POLYGON 13.830 21.025 13.960 21.025 13.830 20.895 ;
        POLYGON 14.110 21.025 14.240 21.025 14.240 20.895 ;
        RECT 14.240 20.895 14.330 21.025 ;
        POLYGON 14.330 21.025 14.460 20.895 14.330 20.895 ;
        POLYGON 16.640 21.025 16.640 20.895 16.510 20.895 ;
        RECT 16.640 20.895 16.730 21.025 ;
        POLYGON 16.730 21.025 16.860 21.025 16.730 20.895 ;
        POLYGON 17.010 21.025 17.140 21.025 17.140 20.895 ;
        RECT 17.140 20.895 17.230 21.025 ;
        POLYGON 17.230 21.025 17.360 20.895 17.230 20.895 ;
        POLYGON 19.540 21.025 19.540 20.895 19.410 20.895 ;
        RECT 19.540 20.895 19.630 21.025 ;
        POLYGON 19.630 21.025 19.760 21.025 19.630 20.895 ;
        POLYGON 19.910 21.025 20.040 21.025 20.040 20.895 ;
        RECT 20.040 20.895 20.130 21.025 ;
        POLYGON 20.130 21.025 20.260 20.895 20.130 20.895 ;
        POLYGON 22.440 21.025 22.440 20.895 22.310 20.895 ;
        RECT 22.440 20.895 22.530 21.025 ;
        POLYGON 22.530 21.025 22.660 21.025 22.530 20.895 ;
        POLYGON 22.810 21.025 22.940 21.025 22.940 20.895 ;
        RECT 22.940 20.895 23.030 21.025 ;
        POLYGON 23.030 21.025 23.160 20.895 23.030 20.895 ;
        POLYGON 25.340 21.025 25.340 20.895 25.210 20.895 ;
        RECT 25.340 20.895 25.430 21.025 ;
        POLYGON 25.430 21.025 25.560 21.025 25.430 20.895 ;
        POLYGON 25.710 21.025 25.840 21.025 25.840 20.895 ;
        RECT 25.840 20.895 25.930 21.025 ;
        POLYGON 25.930 21.025 26.060 20.895 25.930 20.895 ;
        POLYGON 28.240 21.025 28.240 20.895 28.110 20.895 ;
        RECT 28.240 20.895 28.330 21.025 ;
        POLYGON 28.330 21.025 28.460 21.025 28.330 20.895 ;
        POLYGON 28.610 21.025 28.740 21.025 28.740 20.895 ;
        RECT 28.740 20.895 28.830 21.025 ;
        POLYGON 28.830 21.025 28.960 20.895 28.830 20.895 ;
        POLYGON 31.140 21.025 31.140 20.895 31.010 20.895 ;
        RECT 31.140 20.895 31.230 21.025 ;
        POLYGON 31.230 21.025 31.360 21.025 31.230 20.895 ;
        POLYGON 31.510 21.025 31.640 21.025 31.640 20.895 ;
        RECT 31.640 20.895 31.730 21.025 ;
        POLYGON 31.730 21.025 31.860 20.895 31.730 20.895 ;
        POLYGON 34.040 21.025 34.040 20.895 33.910 20.895 ;
        RECT 34.040 20.895 34.130 21.025 ;
        POLYGON 34.130 21.025 34.260 21.025 34.130 20.895 ;
        POLYGON 34.410 21.025 34.540 21.025 34.540 20.895 ;
        RECT 34.540 20.895 34.630 21.025 ;
        POLYGON 34.630 21.025 34.760 20.895 34.630 20.895 ;
        RECT -0.275 20.725 2.060 20.895 ;
        POLYGON 2.060 20.895 2.230 20.895 2.060 20.725 ;
        POLYGON 2.640 20.895 2.810 20.895 2.810 20.725 ;
        RECT 2.810 20.725 4.960 20.895 ;
        POLYGON 4.960 20.895 5.130 20.895 4.960 20.725 ;
        RECT 5.525 20.725 7.860 20.895 ;
        POLYGON 7.860 20.895 8.030 20.895 7.860 20.725 ;
        POLYGON 8.440 20.895 8.610 20.895 8.610 20.725 ;
        RECT 8.610 20.725 10.760 20.895 ;
        POLYGON 10.760 20.895 10.930 20.895 10.760 20.725 ;
        RECT 11.325 20.725 13.660 20.895 ;
        POLYGON 13.660 20.895 13.830 20.895 13.660 20.725 ;
        POLYGON 14.240 20.895 14.410 20.895 14.410 20.725 ;
        RECT 14.410 20.725 16.560 20.895 ;
        POLYGON 16.560 20.895 16.730 20.895 16.560 20.725 ;
        RECT 17.125 20.725 19.460 20.895 ;
        POLYGON 19.460 20.895 19.630 20.895 19.460 20.725 ;
        POLYGON 20.040 20.895 20.210 20.895 20.210 20.725 ;
        RECT 20.210 20.725 22.360 20.895 ;
        POLYGON 22.360 20.895 22.530 20.895 22.360 20.725 ;
        RECT 22.925 20.725 25.260 20.895 ;
        POLYGON 25.260 20.895 25.430 20.895 25.260 20.725 ;
        POLYGON 25.840 20.895 26.010 20.895 26.010 20.725 ;
        RECT 26.010 20.725 28.160 20.895 ;
        POLYGON 28.160 20.895 28.330 20.895 28.160 20.725 ;
        RECT 28.725 20.725 31.060 20.895 ;
        POLYGON 31.060 20.895 31.230 20.895 31.060 20.725 ;
        POLYGON 31.640 20.895 31.810 20.895 31.810 20.725 ;
        RECT 31.810 20.725 33.960 20.895 ;
        POLYGON 33.960 20.895 34.130 20.895 33.960 20.725 ;
        POLYGON 34.540 20.895 34.710 20.895 34.710 20.725 ;
        RECT 34.710 20.725 34.760 20.895 ;
    END
  END RWL1_15
  PIN RBL0_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 5.550 20.405 5.625 20.615 ;
        RECT 5.550 19.055 5.625 19.265 ;
        RECT 5.550 17.705 5.625 17.915 ;
        RECT 5.550 16.355 5.625 16.565 ;
        RECT 5.550 15.005 5.625 15.215 ;
        RECT 5.550 13.655 5.625 13.865 ;
        RECT 5.550 12.305 5.625 12.515 ;
        RECT 5.550 10.955 5.625 11.165 ;
        RECT 5.550 9.605 5.625 9.815 ;
        RECT 5.550 8.255 5.625 8.465 ;
        RECT 5.550 6.905 5.625 7.115 ;
        RECT 5.550 5.555 5.625 5.765 ;
        RECT 5.550 4.205 5.625 4.415 ;
        RECT 5.550 2.855 5.625 3.065 ;
        RECT 5.550 1.505 5.625 1.715 ;
        RECT 5.550 0.155 5.625 0.365 ;
    END
  END RBL0_1
  PIN RBL1_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 2.865 20.405 2.940 20.615 ;
        RECT 2.865 19.055 2.940 19.265 ;
        RECT 2.865 17.705 2.940 17.915 ;
        RECT 2.865 16.355 2.940 16.565 ;
        RECT 2.865 15.005 2.940 15.215 ;
        RECT 2.865 13.655 2.940 13.865 ;
        RECT 2.865 12.305 2.940 12.515 ;
        RECT 2.865 10.955 2.940 11.165 ;
        RECT 2.865 9.605 2.940 9.815 ;
        RECT 2.865 8.255 2.940 8.465 ;
        RECT 2.865 6.905 2.940 7.115 ;
        RECT 2.865 5.555 2.940 5.765 ;
        RECT 2.865 4.205 2.940 4.415 ;
        RECT 2.865 2.855 2.940 3.065 ;
        RECT 2.865 1.505 2.940 1.715 ;
        RECT 2.865 0.155 2.940 0.365 ;
    END
  END RBL1_1
  PIN WBL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 5.185 21.135 5.260 21.280 ;
        RECT 5.185 19.785 5.260 19.930 ;
        RECT 5.185 18.435 5.260 18.580 ;
        RECT 5.185 17.085 5.260 17.230 ;
        RECT 5.185 15.735 5.260 15.880 ;
        RECT 5.185 14.385 5.260 14.530 ;
        RECT 5.185 13.035 5.260 13.180 ;
        RECT 5.185 11.685 5.260 11.830 ;
        RECT 5.185 10.335 5.260 10.480 ;
        RECT 5.185 8.985 5.260 9.130 ;
        RECT 5.185 7.635 5.260 7.780 ;
        RECT 5.185 6.285 5.260 6.430 ;
        RECT 5.185 4.935 5.260 5.080 ;
        RECT 5.185 3.585 5.260 3.730 ;
        RECT 5.185 2.235 5.260 2.380 ;
        RECT 5.185 0.885 5.260 1.030 ;
    END
  END WBL_1
  PIN WBLb_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 3.235 21.135 3.310 21.275 ;
        RECT 3.235 19.785 3.310 19.925 ;
        RECT 3.235 18.435 3.310 18.575 ;
        RECT 3.235 17.085 3.310 17.225 ;
        RECT 3.235 15.735 3.310 15.875 ;
        RECT 3.235 14.385 3.310 14.525 ;
        RECT 3.235 13.035 3.310 13.175 ;
        RECT 3.235 11.685 3.310 11.825 ;
        RECT 3.235 10.335 3.310 10.475 ;
        RECT 3.235 8.985 3.310 9.125 ;
        RECT 3.235 7.635 3.310 7.775 ;
        RECT 3.235 6.285 3.310 6.425 ;
        RECT 3.235 4.935 3.310 5.075 ;
        RECT 3.235 3.585 3.310 3.725 ;
        RECT 3.235 2.235 3.310 2.375 ;
        RECT 3.235 0.885 3.310 1.025 ;
    END
  END WBLb_1
  PIN RBL0_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 8.450 20.405 8.525 20.615 ;
        RECT 8.450 19.055 8.525 19.265 ;
        RECT 8.450 17.705 8.525 17.915 ;
        RECT 8.450 16.355 8.525 16.565 ;
        RECT 8.450 15.005 8.525 15.215 ;
        RECT 8.450 13.655 8.525 13.865 ;
        RECT 8.450 12.305 8.525 12.515 ;
        RECT 8.450 10.955 8.525 11.165 ;
        RECT 8.450 9.605 8.525 9.815 ;
        RECT 8.450 8.255 8.525 8.465 ;
        RECT 8.450 6.905 8.525 7.115 ;
        RECT 8.450 5.555 8.525 5.765 ;
        RECT 8.450 4.205 8.525 4.415 ;
        RECT 8.450 2.855 8.525 3.065 ;
        RECT 8.450 1.505 8.525 1.715 ;
        RECT 8.450 0.155 8.525 0.365 ;
    END
  END RBL0_2
  PIN RBL1_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 5.765 20.405 5.840 20.615 ;
        RECT 5.765 19.055 5.840 19.265 ;
        RECT 5.765 17.705 5.840 17.915 ;
        RECT 5.765 16.355 5.840 16.565 ;
        RECT 5.765 15.005 5.840 15.215 ;
        RECT 5.765 13.655 5.840 13.865 ;
        RECT 5.765 12.305 5.840 12.515 ;
        RECT 5.765 10.955 5.840 11.165 ;
        RECT 5.765 9.605 5.840 9.815 ;
        RECT 5.765 8.255 5.840 8.465 ;
        RECT 5.765 6.905 5.840 7.115 ;
        RECT 5.765 5.555 5.840 5.765 ;
        RECT 5.765 4.205 5.840 4.415 ;
        RECT 5.765 2.855 5.840 3.065 ;
        RECT 5.765 1.505 5.840 1.715 ;
        RECT 5.765 0.155 5.840 0.365 ;
    END
  END RBL1_2
  PIN WBL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 8.085 21.135 8.160 21.280 ;
        RECT 8.085 19.785 8.160 19.930 ;
        RECT 8.085 18.435 8.160 18.580 ;
        RECT 8.085 17.085 8.160 17.230 ;
        RECT 8.085 15.735 8.160 15.880 ;
        RECT 8.085 14.385 8.160 14.530 ;
        RECT 8.085 13.035 8.160 13.180 ;
        RECT 8.085 11.685 8.160 11.830 ;
        RECT 8.085 10.335 8.160 10.480 ;
        RECT 8.085 8.985 8.160 9.130 ;
        RECT 8.085 7.635 8.160 7.780 ;
        RECT 8.085 6.285 8.160 6.430 ;
        RECT 8.085 4.935 8.160 5.080 ;
        RECT 8.085 3.585 8.160 3.730 ;
        RECT 8.085 2.235 8.160 2.380 ;
        RECT 8.085 0.885 8.160 1.030 ;
    END
  END WBL_2
  PIN WBLb_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 6.135 21.135 6.210 21.275 ;
        RECT 6.135 19.785 6.210 19.925 ;
        RECT 6.135 18.435 6.210 18.575 ;
        RECT 6.135 17.085 6.210 17.225 ;
        RECT 6.135 15.735 6.210 15.875 ;
        RECT 6.135 14.385 6.210 14.525 ;
        RECT 6.135 13.035 6.210 13.175 ;
        RECT 6.135 11.685 6.210 11.825 ;
        RECT 6.135 10.335 6.210 10.475 ;
        RECT 6.135 8.985 6.210 9.125 ;
        RECT 6.135 7.635 6.210 7.775 ;
        RECT 6.135 6.285 6.210 6.425 ;
        RECT 6.135 4.935 6.210 5.075 ;
        RECT 6.135 3.585 6.210 3.725 ;
        RECT 6.135 2.235 6.210 2.375 ;
        RECT 6.135 0.885 6.210 1.025 ;
    END
  END WBLb_2
  PIN RBL0_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 11.350 20.405 11.425 20.615 ;
        RECT 11.350 19.055 11.425 19.265 ;
        RECT 11.350 17.705 11.425 17.915 ;
        RECT 11.350 16.355 11.425 16.565 ;
        RECT 11.350 15.005 11.425 15.215 ;
        RECT 11.350 13.655 11.425 13.865 ;
        RECT 11.350 12.305 11.425 12.515 ;
        RECT 11.350 10.955 11.425 11.165 ;
        RECT 11.350 9.605 11.425 9.815 ;
        RECT 11.350 8.255 11.425 8.465 ;
        RECT 11.350 6.905 11.425 7.115 ;
        RECT 11.350 5.555 11.425 5.765 ;
        RECT 11.350 4.205 11.425 4.415 ;
        RECT 11.350 2.855 11.425 3.065 ;
        RECT 11.350 1.505 11.425 1.715 ;
        RECT 11.350 0.155 11.425 0.365 ;
    END
  END RBL0_3
  PIN RBL1_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 8.665 20.405 8.740 20.615 ;
        RECT 8.665 19.055 8.740 19.265 ;
        RECT 8.665 17.705 8.740 17.915 ;
        RECT 8.665 16.355 8.740 16.565 ;
        RECT 8.665 15.005 8.740 15.215 ;
        RECT 8.665 13.655 8.740 13.865 ;
        RECT 8.665 12.305 8.740 12.515 ;
        RECT 8.665 10.955 8.740 11.165 ;
        RECT 8.665 9.605 8.740 9.815 ;
        RECT 8.665 8.255 8.740 8.465 ;
        RECT 8.665 6.905 8.740 7.115 ;
        RECT 8.665 5.555 8.740 5.765 ;
        RECT 8.665 4.205 8.740 4.415 ;
        RECT 8.665 2.855 8.740 3.065 ;
        RECT 8.665 1.505 8.740 1.715 ;
        RECT 8.665 0.155 8.740 0.365 ;
    END
  END RBL1_3
  PIN WBL_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 10.985 21.135 11.060 21.280 ;
        RECT 10.985 19.785 11.060 19.930 ;
        RECT 10.985 18.435 11.060 18.580 ;
        RECT 10.985 17.085 11.060 17.230 ;
        RECT 10.985 15.735 11.060 15.880 ;
        RECT 10.985 14.385 11.060 14.530 ;
        RECT 10.985 13.035 11.060 13.180 ;
        RECT 10.985 11.685 11.060 11.830 ;
        RECT 10.985 10.335 11.060 10.480 ;
        RECT 10.985 8.985 11.060 9.130 ;
        RECT 10.985 7.635 11.060 7.780 ;
        RECT 10.985 6.285 11.060 6.430 ;
        RECT 10.985 4.935 11.060 5.080 ;
        RECT 10.985 3.585 11.060 3.730 ;
        RECT 10.985 2.235 11.060 2.380 ;
        RECT 10.985 0.885 11.060 1.030 ;
    END
  END WBL_3
  PIN WBLb_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 9.035 21.135 9.110 21.275 ;
        RECT 9.035 19.785 9.110 19.925 ;
        RECT 9.035 18.435 9.110 18.575 ;
        RECT 9.035 17.085 9.110 17.225 ;
        RECT 9.035 15.735 9.110 15.875 ;
        RECT 9.035 14.385 9.110 14.525 ;
        RECT 9.035 13.035 9.110 13.175 ;
        RECT 9.035 11.685 9.110 11.825 ;
        RECT 9.035 10.335 9.110 10.475 ;
        RECT 9.035 8.985 9.110 9.125 ;
        RECT 9.035 7.635 9.110 7.775 ;
        RECT 9.035 6.285 9.110 6.425 ;
        RECT 9.035 4.935 9.110 5.075 ;
        RECT 9.035 3.585 9.110 3.725 ;
        RECT 9.035 2.235 9.110 2.375 ;
        RECT 9.035 0.885 9.110 1.025 ;
    END
  END WBLb_3
  PIN RBL0_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 14.250 20.405 14.325 20.615 ;
        RECT 14.250 19.055 14.325 19.265 ;
        RECT 14.250 17.705 14.325 17.915 ;
        RECT 14.250 16.355 14.325 16.565 ;
        RECT 14.250 15.005 14.325 15.215 ;
        RECT 14.250 13.655 14.325 13.865 ;
        RECT 14.250 12.305 14.325 12.515 ;
        RECT 14.250 10.955 14.325 11.165 ;
        RECT 14.250 9.605 14.325 9.815 ;
        RECT 14.250 8.255 14.325 8.465 ;
        RECT 14.250 6.905 14.325 7.115 ;
        RECT 14.250 5.555 14.325 5.765 ;
        RECT 14.250 4.205 14.325 4.415 ;
        RECT 14.250 2.855 14.325 3.065 ;
        RECT 14.250 1.505 14.325 1.715 ;
        RECT 14.250 0.155 14.325 0.365 ;
    END
  END RBL0_4
  PIN RBL1_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 11.565 20.405 11.640 20.615 ;
        RECT 11.565 19.055 11.640 19.265 ;
        RECT 11.565 17.705 11.640 17.915 ;
        RECT 11.565 16.355 11.640 16.565 ;
        RECT 11.565 15.005 11.640 15.215 ;
        RECT 11.565 13.655 11.640 13.865 ;
        RECT 11.565 12.305 11.640 12.515 ;
        RECT 11.565 10.955 11.640 11.165 ;
        RECT 11.565 9.605 11.640 9.815 ;
        RECT 11.565 8.255 11.640 8.465 ;
        RECT 11.565 6.905 11.640 7.115 ;
        RECT 11.565 5.555 11.640 5.765 ;
        RECT 11.565 4.205 11.640 4.415 ;
        RECT 11.565 2.855 11.640 3.065 ;
        RECT 11.565 1.505 11.640 1.715 ;
        RECT 11.565 0.155 11.640 0.365 ;
    END
  END RBL1_4
  PIN WBL_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 13.885 21.135 13.960 21.280 ;
        RECT 13.885 19.785 13.960 19.930 ;
        RECT 13.885 18.435 13.960 18.580 ;
        RECT 13.885 17.085 13.960 17.230 ;
        RECT 13.885 15.735 13.960 15.880 ;
        RECT 13.885 14.385 13.960 14.530 ;
        RECT 13.885 13.035 13.960 13.180 ;
        RECT 13.885 11.685 13.960 11.830 ;
        RECT 13.885 10.335 13.960 10.480 ;
        RECT 13.885 8.985 13.960 9.130 ;
        RECT 13.885 7.635 13.960 7.780 ;
        RECT 13.885 6.285 13.960 6.430 ;
        RECT 13.885 4.935 13.960 5.080 ;
        RECT 13.885 3.585 13.960 3.730 ;
        RECT 13.885 2.235 13.960 2.380 ;
        RECT 13.885 0.885 13.960 1.030 ;
    END
  END WBL_4
  PIN WBLb_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 11.935 21.135 12.010 21.275 ;
        RECT 11.935 19.785 12.010 19.925 ;
        RECT 11.935 18.435 12.010 18.575 ;
        RECT 11.935 17.085 12.010 17.225 ;
        RECT 11.935 15.735 12.010 15.875 ;
        RECT 11.935 14.385 12.010 14.525 ;
        RECT 11.935 13.035 12.010 13.175 ;
        RECT 11.935 11.685 12.010 11.825 ;
        RECT 11.935 10.335 12.010 10.475 ;
        RECT 11.935 8.985 12.010 9.125 ;
        RECT 11.935 7.635 12.010 7.775 ;
        RECT 11.935 6.285 12.010 6.425 ;
        RECT 11.935 4.935 12.010 5.075 ;
        RECT 11.935 3.585 12.010 3.725 ;
        RECT 11.935 2.235 12.010 2.375 ;
        RECT 11.935 0.885 12.010 1.025 ;
    END
  END WBLb_4
  PIN RBL0_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 17.150 20.405 17.225 20.615 ;
        RECT 17.150 19.055 17.225 19.265 ;
        RECT 17.150 17.705 17.225 17.915 ;
        RECT 17.150 16.355 17.225 16.565 ;
        RECT 17.150 15.005 17.225 15.215 ;
        RECT 17.150 13.655 17.225 13.865 ;
        RECT 17.150 12.305 17.225 12.515 ;
        RECT 17.150 10.955 17.225 11.165 ;
        RECT 17.150 9.605 17.225 9.815 ;
        RECT 17.150 8.255 17.225 8.465 ;
        RECT 17.150 6.905 17.225 7.115 ;
        RECT 17.150 5.555 17.225 5.765 ;
        RECT 17.150 4.205 17.225 4.415 ;
        RECT 17.150 2.855 17.225 3.065 ;
        RECT 17.150 1.505 17.225 1.715 ;
        RECT 17.150 0.155 17.225 0.365 ;
    END
  END RBL0_5
  PIN RBL1_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 14.465 20.405 14.540 20.615 ;
        RECT 14.465 19.055 14.540 19.265 ;
        RECT 14.465 17.705 14.540 17.915 ;
        RECT 14.465 16.355 14.540 16.565 ;
        RECT 14.465 15.005 14.540 15.215 ;
        RECT 14.465 13.655 14.540 13.865 ;
        RECT 14.465 12.305 14.540 12.515 ;
        RECT 14.465 10.955 14.540 11.165 ;
        RECT 14.465 9.605 14.540 9.815 ;
        RECT 14.465 8.255 14.540 8.465 ;
        RECT 14.465 6.905 14.540 7.115 ;
        RECT 14.465 5.555 14.540 5.765 ;
        RECT 14.465 4.205 14.540 4.415 ;
        RECT 14.465 2.855 14.540 3.065 ;
        RECT 14.465 1.505 14.540 1.715 ;
        RECT 14.465 0.155 14.540 0.365 ;
    END
  END RBL1_5
  PIN WBL_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 16.785 21.135 16.860 21.280 ;
        RECT 16.785 19.785 16.860 19.930 ;
        RECT 16.785 18.435 16.860 18.580 ;
        RECT 16.785 17.085 16.860 17.230 ;
        RECT 16.785 15.735 16.860 15.880 ;
        RECT 16.785 14.385 16.860 14.530 ;
        RECT 16.785 13.035 16.860 13.180 ;
        RECT 16.785 11.685 16.860 11.830 ;
        RECT 16.785 10.335 16.860 10.480 ;
        RECT 16.785 8.985 16.860 9.130 ;
        RECT 16.785 7.635 16.860 7.780 ;
        RECT 16.785 6.285 16.860 6.430 ;
        RECT 16.785 4.935 16.860 5.080 ;
        RECT 16.785 3.585 16.860 3.730 ;
        RECT 16.785 2.235 16.860 2.380 ;
        RECT 16.785 0.885 16.860 1.030 ;
    END
  END WBL_5
  PIN WBLb_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 14.835 21.135 14.910 21.275 ;
        RECT 14.835 19.785 14.910 19.925 ;
        RECT 14.835 18.435 14.910 18.575 ;
        RECT 14.835 17.085 14.910 17.225 ;
        RECT 14.835 15.735 14.910 15.875 ;
        RECT 14.835 14.385 14.910 14.525 ;
        RECT 14.835 13.035 14.910 13.175 ;
        RECT 14.835 11.685 14.910 11.825 ;
        RECT 14.835 10.335 14.910 10.475 ;
        RECT 14.835 8.985 14.910 9.125 ;
        RECT 14.835 7.635 14.910 7.775 ;
        RECT 14.835 6.285 14.910 6.425 ;
        RECT 14.835 4.935 14.910 5.075 ;
        RECT 14.835 3.585 14.910 3.725 ;
        RECT 14.835 2.235 14.910 2.375 ;
        RECT 14.835 0.885 14.910 1.025 ;
    END
  END WBLb_5
  PIN RBL0_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 20.050 20.405 20.125 20.615 ;
        RECT 20.050 19.055 20.125 19.265 ;
        RECT 20.050 17.705 20.125 17.915 ;
        RECT 20.050 16.355 20.125 16.565 ;
        RECT 20.050 15.005 20.125 15.215 ;
        RECT 20.050 13.655 20.125 13.865 ;
        RECT 20.050 12.305 20.125 12.515 ;
        RECT 20.050 10.955 20.125 11.165 ;
        RECT 20.050 9.605 20.125 9.815 ;
        RECT 20.050 8.255 20.125 8.465 ;
        RECT 20.050 6.905 20.125 7.115 ;
        RECT 20.050 5.555 20.125 5.765 ;
        RECT 20.050 4.205 20.125 4.415 ;
        RECT 20.050 2.855 20.125 3.065 ;
        RECT 20.050 1.505 20.125 1.715 ;
        RECT 20.050 0.155 20.125 0.365 ;
    END
  END RBL0_6
  PIN RBL1_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 17.365 20.405 17.440 20.615 ;
        RECT 17.365 19.055 17.440 19.265 ;
        RECT 17.365 17.705 17.440 17.915 ;
        RECT 17.365 16.355 17.440 16.565 ;
        RECT 17.365 15.005 17.440 15.215 ;
        RECT 17.365 13.655 17.440 13.865 ;
        RECT 17.365 12.305 17.440 12.515 ;
        RECT 17.365 10.955 17.440 11.165 ;
        RECT 17.365 9.605 17.440 9.815 ;
        RECT 17.365 8.255 17.440 8.465 ;
        RECT 17.365 6.905 17.440 7.115 ;
        RECT 17.365 5.555 17.440 5.765 ;
        RECT 17.365 4.205 17.440 4.415 ;
        RECT 17.365 2.855 17.440 3.065 ;
        RECT 17.365 1.505 17.440 1.715 ;
        RECT 17.365 0.155 17.440 0.365 ;
    END
  END RBL1_6
  PIN WBL_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 19.685 21.135 19.760 21.280 ;
        RECT 19.685 19.785 19.760 19.930 ;
        RECT 19.685 18.435 19.760 18.580 ;
        RECT 19.685 17.085 19.760 17.230 ;
        RECT 19.685 15.735 19.760 15.880 ;
        RECT 19.685 14.385 19.760 14.530 ;
        RECT 19.685 13.035 19.760 13.180 ;
        RECT 19.685 11.685 19.760 11.830 ;
        RECT 19.685 10.335 19.760 10.480 ;
        RECT 19.685 8.985 19.760 9.130 ;
        RECT 19.685 7.635 19.760 7.780 ;
        RECT 19.685 6.285 19.760 6.430 ;
        RECT 19.685 4.935 19.760 5.080 ;
        RECT 19.685 3.585 19.760 3.730 ;
        RECT 19.685 2.235 19.760 2.380 ;
        RECT 19.685 0.885 19.760 1.030 ;
    END
  END WBL_6
  PIN WBLb_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 17.735 21.135 17.810 21.275 ;
        RECT 17.735 19.785 17.810 19.925 ;
        RECT 17.735 18.435 17.810 18.575 ;
        RECT 17.735 17.085 17.810 17.225 ;
        RECT 17.735 15.735 17.810 15.875 ;
        RECT 17.735 14.385 17.810 14.525 ;
        RECT 17.735 13.035 17.810 13.175 ;
        RECT 17.735 11.685 17.810 11.825 ;
        RECT 17.735 10.335 17.810 10.475 ;
        RECT 17.735 8.985 17.810 9.125 ;
        RECT 17.735 7.635 17.810 7.775 ;
        RECT 17.735 6.285 17.810 6.425 ;
        RECT 17.735 4.935 17.810 5.075 ;
        RECT 17.735 3.585 17.810 3.725 ;
        RECT 17.735 2.235 17.810 2.375 ;
        RECT 17.735 0.885 17.810 1.025 ;
    END
  END WBLb_6
  PIN RBL0_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 22.950 20.405 23.025 20.615 ;
        RECT 22.950 19.055 23.025 19.265 ;
        RECT 22.950 17.705 23.025 17.915 ;
        RECT 22.950 16.355 23.025 16.565 ;
        RECT 22.950 15.005 23.025 15.215 ;
        RECT 22.950 13.655 23.025 13.865 ;
        RECT 22.950 12.305 23.025 12.515 ;
        RECT 22.950 10.955 23.025 11.165 ;
        RECT 22.950 9.605 23.025 9.815 ;
        RECT 22.950 8.255 23.025 8.465 ;
        RECT 22.950 6.905 23.025 7.115 ;
        RECT 22.950 5.555 23.025 5.765 ;
        RECT 22.950 4.205 23.025 4.415 ;
        RECT 22.950 2.855 23.025 3.065 ;
        RECT 22.950 1.505 23.025 1.715 ;
        RECT 22.950 0.155 23.025 0.365 ;
    END
  END RBL0_7
  PIN RBL1_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 20.265 20.405 20.340 20.615 ;
        RECT 20.265 19.055 20.340 19.265 ;
        RECT 20.265 17.705 20.340 17.915 ;
        RECT 20.265 16.355 20.340 16.565 ;
        RECT 20.265 15.005 20.340 15.215 ;
        RECT 20.265 13.655 20.340 13.865 ;
        RECT 20.265 12.305 20.340 12.515 ;
        RECT 20.265 10.955 20.340 11.165 ;
        RECT 20.265 9.605 20.340 9.815 ;
        RECT 20.265 8.255 20.340 8.465 ;
        RECT 20.265 6.905 20.340 7.115 ;
        RECT 20.265 5.555 20.340 5.765 ;
        RECT 20.265 4.205 20.340 4.415 ;
        RECT 20.265 2.855 20.340 3.065 ;
        RECT 20.265 1.505 20.340 1.715 ;
        RECT 20.265 0.155 20.340 0.365 ;
    END
  END RBL1_7
  PIN WBL_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 22.585 21.135 22.660 21.280 ;
        RECT 22.585 19.785 22.660 19.930 ;
        RECT 22.585 18.435 22.660 18.580 ;
        RECT 22.585 17.085 22.660 17.230 ;
        RECT 22.585 15.735 22.660 15.880 ;
        RECT 22.585 14.385 22.660 14.530 ;
        RECT 22.585 13.035 22.660 13.180 ;
        RECT 22.585 11.685 22.660 11.830 ;
        RECT 22.585 10.335 22.660 10.480 ;
        RECT 22.585 8.985 22.660 9.130 ;
        RECT 22.585 7.635 22.660 7.780 ;
        RECT 22.585 6.285 22.660 6.430 ;
        RECT 22.585 4.935 22.660 5.080 ;
        RECT 22.585 3.585 22.660 3.730 ;
        RECT 22.585 2.235 22.660 2.380 ;
        RECT 22.585 0.885 22.660 1.030 ;
    END
  END WBL_7
  PIN WBLb_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 20.635 21.135 20.710 21.275 ;
        RECT 20.635 19.785 20.710 19.925 ;
        RECT 20.635 18.435 20.710 18.575 ;
        RECT 20.635 17.085 20.710 17.225 ;
        RECT 20.635 15.735 20.710 15.875 ;
        RECT 20.635 14.385 20.710 14.525 ;
        RECT 20.635 13.035 20.710 13.175 ;
        RECT 20.635 11.685 20.710 11.825 ;
        RECT 20.635 10.335 20.710 10.475 ;
        RECT 20.635 8.985 20.710 9.125 ;
        RECT 20.635 7.635 20.710 7.775 ;
        RECT 20.635 6.285 20.710 6.425 ;
        RECT 20.635 4.935 20.710 5.075 ;
        RECT 20.635 3.585 20.710 3.725 ;
        RECT 20.635 2.235 20.710 2.375 ;
        RECT 20.635 0.885 20.710 1.025 ;
    END
  END WBLb_7
  PIN RBL0_8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 25.850 20.405 25.925 20.615 ;
        RECT 25.850 19.055 25.925 19.265 ;
        RECT 25.850 17.705 25.925 17.915 ;
        RECT 25.850 16.355 25.925 16.565 ;
        RECT 25.850 15.005 25.925 15.215 ;
        RECT 25.850 13.655 25.925 13.865 ;
        RECT 25.850 12.305 25.925 12.515 ;
        RECT 25.850 10.955 25.925 11.165 ;
        RECT 25.850 9.605 25.925 9.815 ;
        RECT 25.850 8.255 25.925 8.465 ;
        RECT 25.850 6.905 25.925 7.115 ;
        RECT 25.850 5.555 25.925 5.765 ;
        RECT 25.850 4.205 25.925 4.415 ;
        RECT 25.850 2.855 25.925 3.065 ;
        RECT 25.850 1.505 25.925 1.715 ;
        RECT 25.850 0.155 25.925 0.365 ;
    END
  END RBL0_8
  PIN RBL1_8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 23.165 20.405 23.240 20.615 ;
        RECT 23.165 19.055 23.240 19.265 ;
        RECT 23.165 17.705 23.240 17.915 ;
        RECT 23.165 16.355 23.240 16.565 ;
        RECT 23.165 15.005 23.240 15.215 ;
        RECT 23.165 13.655 23.240 13.865 ;
        RECT 23.165 12.305 23.240 12.515 ;
        RECT 23.165 10.955 23.240 11.165 ;
        RECT 23.165 9.605 23.240 9.815 ;
        RECT 23.165 8.255 23.240 8.465 ;
        RECT 23.165 6.905 23.240 7.115 ;
        RECT 23.165 5.555 23.240 5.765 ;
        RECT 23.165 4.205 23.240 4.415 ;
        RECT 23.165 2.855 23.240 3.065 ;
        RECT 23.165 1.505 23.240 1.715 ;
        RECT 23.165 0.155 23.240 0.365 ;
    END
  END RBL1_8
  PIN WBL_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 25.485 21.135 25.560 21.280 ;
        RECT 25.485 19.785 25.560 19.930 ;
        RECT 25.485 18.435 25.560 18.580 ;
        RECT 25.485 17.085 25.560 17.230 ;
        RECT 25.485 15.735 25.560 15.880 ;
        RECT 25.485 14.385 25.560 14.530 ;
        RECT 25.485 13.035 25.560 13.180 ;
        RECT 25.485 11.685 25.560 11.830 ;
        RECT 25.485 10.335 25.560 10.480 ;
        RECT 25.485 8.985 25.560 9.130 ;
        RECT 25.485 7.635 25.560 7.780 ;
        RECT 25.485 6.285 25.560 6.430 ;
        RECT 25.485 4.935 25.560 5.080 ;
        RECT 25.485 3.585 25.560 3.730 ;
        RECT 25.485 2.235 25.560 2.380 ;
        RECT 25.485 0.885 25.560 1.030 ;
    END
  END WBL_8
  PIN WBLb_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 23.535 21.135 23.610 21.275 ;
        RECT 23.535 19.785 23.610 19.925 ;
        RECT 23.535 18.435 23.610 18.575 ;
        RECT 23.535 17.085 23.610 17.225 ;
        RECT 23.535 15.735 23.610 15.875 ;
        RECT 23.535 14.385 23.610 14.525 ;
        RECT 23.535 13.035 23.610 13.175 ;
        RECT 23.535 11.685 23.610 11.825 ;
        RECT 23.535 10.335 23.610 10.475 ;
        RECT 23.535 8.985 23.610 9.125 ;
        RECT 23.535 7.635 23.610 7.775 ;
        RECT 23.535 6.285 23.610 6.425 ;
        RECT 23.535 4.935 23.610 5.075 ;
        RECT 23.535 3.585 23.610 3.725 ;
        RECT 23.535 2.235 23.610 2.375 ;
        RECT 23.535 0.885 23.610 1.025 ;
    END
  END WBLb_8
  PIN RBL0_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 28.750 20.405 28.825 20.615 ;
        RECT 28.750 19.055 28.825 19.265 ;
        RECT 28.750 17.705 28.825 17.915 ;
        RECT 28.750 16.355 28.825 16.565 ;
        RECT 28.750 15.005 28.825 15.215 ;
        RECT 28.750 13.655 28.825 13.865 ;
        RECT 28.750 12.305 28.825 12.515 ;
        RECT 28.750 10.955 28.825 11.165 ;
        RECT 28.750 9.605 28.825 9.815 ;
        RECT 28.750 8.255 28.825 8.465 ;
        RECT 28.750 6.905 28.825 7.115 ;
        RECT 28.750 5.555 28.825 5.765 ;
        RECT 28.750 4.205 28.825 4.415 ;
        RECT 28.750 2.855 28.825 3.065 ;
        RECT 28.750 1.505 28.825 1.715 ;
        RECT 28.750 0.155 28.825 0.365 ;
    END
  END RBL0_9
  PIN RBL1_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 26.065 20.405 26.140 20.615 ;
        RECT 26.065 19.055 26.140 19.265 ;
        RECT 26.065 17.705 26.140 17.915 ;
        RECT 26.065 16.355 26.140 16.565 ;
        RECT 26.065 15.005 26.140 15.215 ;
        RECT 26.065 13.655 26.140 13.865 ;
        RECT 26.065 12.305 26.140 12.515 ;
        RECT 26.065 10.955 26.140 11.165 ;
        RECT 26.065 9.605 26.140 9.815 ;
        RECT 26.065 8.255 26.140 8.465 ;
        RECT 26.065 6.905 26.140 7.115 ;
        RECT 26.065 5.555 26.140 5.765 ;
        RECT 26.065 4.205 26.140 4.415 ;
        RECT 26.065 2.855 26.140 3.065 ;
        RECT 26.065 1.505 26.140 1.715 ;
        RECT 26.065 0.155 26.140 0.365 ;
    END
  END RBL1_9
  PIN WBL_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 28.385 21.135 28.460 21.280 ;
        RECT 28.385 19.785 28.460 19.930 ;
        RECT 28.385 18.435 28.460 18.580 ;
        RECT 28.385 17.085 28.460 17.230 ;
        RECT 28.385 15.735 28.460 15.880 ;
        RECT 28.385 14.385 28.460 14.530 ;
        RECT 28.385 13.035 28.460 13.180 ;
        RECT 28.385 11.685 28.460 11.830 ;
        RECT 28.385 10.335 28.460 10.480 ;
        RECT 28.385 8.985 28.460 9.130 ;
        RECT 28.385 7.635 28.460 7.780 ;
        RECT 28.385 6.285 28.460 6.430 ;
        RECT 28.385 4.935 28.460 5.080 ;
        RECT 28.385 3.585 28.460 3.730 ;
        RECT 28.385 2.235 28.460 2.380 ;
        RECT 28.385 0.885 28.460 1.030 ;
    END
  END WBL_9
  PIN WBLb_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 26.435 21.135 26.510 21.275 ;
        RECT 26.435 19.785 26.510 19.925 ;
        RECT 26.435 18.435 26.510 18.575 ;
        RECT 26.435 17.085 26.510 17.225 ;
        RECT 26.435 15.735 26.510 15.875 ;
        RECT 26.435 14.385 26.510 14.525 ;
        RECT 26.435 13.035 26.510 13.175 ;
        RECT 26.435 11.685 26.510 11.825 ;
        RECT 26.435 10.335 26.510 10.475 ;
        RECT 26.435 8.985 26.510 9.125 ;
        RECT 26.435 7.635 26.510 7.775 ;
        RECT 26.435 6.285 26.510 6.425 ;
        RECT 26.435 4.935 26.510 5.075 ;
        RECT 26.435 3.585 26.510 3.725 ;
        RECT 26.435 2.235 26.510 2.375 ;
        RECT 26.435 0.885 26.510 1.025 ;
    END
  END WBLb_9
  PIN RBL0_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 31.650 20.405 31.725 20.615 ;
        RECT 31.650 19.055 31.725 19.265 ;
        RECT 31.650 17.705 31.725 17.915 ;
        RECT 31.650 16.355 31.725 16.565 ;
        RECT 31.650 15.005 31.725 15.215 ;
        RECT 31.650 13.655 31.725 13.865 ;
        RECT 31.650 12.305 31.725 12.515 ;
        RECT 31.650 10.955 31.725 11.165 ;
        RECT 31.650 9.605 31.725 9.815 ;
        RECT 31.650 8.255 31.725 8.465 ;
        RECT 31.650 6.905 31.725 7.115 ;
        RECT 31.650 5.555 31.725 5.765 ;
        RECT 31.650 4.205 31.725 4.415 ;
        RECT 31.650 2.855 31.725 3.065 ;
        RECT 31.650 1.505 31.725 1.715 ;
        RECT 31.650 0.155 31.725 0.365 ;
    END
  END RBL0_10
  PIN RBL1_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 28.965 20.405 29.040 20.615 ;
        RECT 28.965 19.055 29.040 19.265 ;
        RECT 28.965 17.705 29.040 17.915 ;
        RECT 28.965 16.355 29.040 16.565 ;
        RECT 28.965 15.005 29.040 15.215 ;
        RECT 28.965 13.655 29.040 13.865 ;
        RECT 28.965 12.305 29.040 12.515 ;
        RECT 28.965 10.955 29.040 11.165 ;
        RECT 28.965 9.605 29.040 9.815 ;
        RECT 28.965 8.255 29.040 8.465 ;
        RECT 28.965 6.905 29.040 7.115 ;
        RECT 28.965 5.555 29.040 5.765 ;
        RECT 28.965 4.205 29.040 4.415 ;
        RECT 28.965 2.855 29.040 3.065 ;
        RECT 28.965 1.505 29.040 1.715 ;
        RECT 28.965 0.155 29.040 0.365 ;
    END
  END RBL1_10
  PIN WBL_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 31.285 21.135 31.360 21.280 ;
        RECT 31.285 19.785 31.360 19.930 ;
        RECT 31.285 18.435 31.360 18.580 ;
        RECT 31.285 17.085 31.360 17.230 ;
        RECT 31.285 15.735 31.360 15.880 ;
        RECT 31.285 14.385 31.360 14.530 ;
        RECT 31.285 13.035 31.360 13.180 ;
        RECT 31.285 11.685 31.360 11.830 ;
        RECT 31.285 10.335 31.360 10.480 ;
        RECT 31.285 8.985 31.360 9.130 ;
        RECT 31.285 7.635 31.360 7.780 ;
        RECT 31.285 6.285 31.360 6.430 ;
        RECT 31.285 4.935 31.360 5.080 ;
        RECT 31.285 3.585 31.360 3.730 ;
        RECT 31.285 2.235 31.360 2.380 ;
        RECT 31.285 0.885 31.360 1.030 ;
    END
  END WBL_10
  PIN WBLb_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 29.335 21.135 29.410 21.275 ;
        RECT 29.335 19.785 29.410 19.925 ;
        RECT 29.335 18.435 29.410 18.575 ;
        RECT 29.335 17.085 29.410 17.225 ;
        RECT 29.335 15.735 29.410 15.875 ;
        RECT 29.335 14.385 29.410 14.525 ;
        RECT 29.335 13.035 29.410 13.175 ;
        RECT 29.335 11.685 29.410 11.825 ;
        RECT 29.335 10.335 29.410 10.475 ;
        RECT 29.335 8.985 29.410 9.125 ;
        RECT 29.335 7.635 29.410 7.775 ;
        RECT 29.335 6.285 29.410 6.425 ;
        RECT 29.335 4.935 29.410 5.075 ;
        RECT 29.335 3.585 29.410 3.725 ;
        RECT 29.335 2.235 29.410 2.375 ;
        RECT 29.335 0.885 29.410 1.025 ;
    END
  END WBLb_10
  PIN RBL0_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 34.550 20.405 34.625 20.615 ;
        RECT 34.550 19.055 34.625 19.265 ;
        RECT 34.550 17.705 34.625 17.915 ;
        RECT 34.550 16.355 34.625 16.565 ;
        RECT 34.550 15.005 34.625 15.215 ;
        RECT 34.550 13.655 34.625 13.865 ;
        RECT 34.550 12.305 34.625 12.515 ;
        RECT 34.550 10.955 34.625 11.165 ;
        RECT 34.550 9.605 34.625 9.815 ;
        RECT 34.550 8.255 34.625 8.465 ;
        RECT 34.550 6.905 34.625 7.115 ;
        RECT 34.550 5.555 34.625 5.765 ;
        RECT 34.550 4.205 34.625 4.415 ;
        RECT 34.550 2.855 34.625 3.065 ;
        RECT 34.550 1.505 34.625 1.715 ;
        RECT 34.550 0.155 34.625 0.365 ;
    END
  END RBL0_11
  PIN RBL1_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.722400 ;
    PORT
      LAYER li1 ;
        RECT 31.865 20.405 31.940 20.615 ;
        RECT 31.865 19.055 31.940 19.265 ;
        RECT 31.865 17.705 31.940 17.915 ;
        RECT 31.865 16.355 31.940 16.565 ;
        RECT 31.865 15.005 31.940 15.215 ;
        RECT 31.865 13.655 31.940 13.865 ;
        RECT 31.865 12.305 31.940 12.515 ;
        RECT 31.865 10.955 31.940 11.165 ;
        RECT 31.865 9.605 31.940 9.815 ;
        RECT 31.865 8.255 31.940 8.465 ;
        RECT 31.865 6.905 31.940 7.115 ;
        RECT 31.865 5.555 31.940 5.765 ;
        RECT 31.865 4.205 31.940 4.415 ;
        RECT 31.865 2.855 31.940 3.065 ;
        RECT 31.865 1.505 31.940 1.715 ;
        RECT 31.865 0.155 31.940 0.365 ;
    END
  END RBL1_11
  PIN WBL_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.386800 ;
    PORT
      LAYER li1 ;
        RECT 34.185 21.135 34.260 21.280 ;
        RECT 34.185 19.785 34.260 19.930 ;
        RECT 34.185 18.435 34.260 18.580 ;
        RECT 34.185 17.085 34.260 17.230 ;
        RECT 34.185 15.735 34.260 15.880 ;
        RECT 34.185 14.385 34.260 14.530 ;
        RECT 34.185 13.035 34.260 13.180 ;
        RECT 34.185 11.685 34.260 11.830 ;
        RECT 34.185 10.335 34.260 10.480 ;
        RECT 34.185 8.985 34.260 9.130 ;
        RECT 34.185 7.635 34.260 7.780 ;
        RECT 34.185 6.285 34.260 6.430 ;
        RECT 34.185 4.935 34.260 5.080 ;
        RECT 34.185 3.585 34.260 3.730 ;
        RECT 34.185 2.235 34.260 2.380 ;
        RECT 34.185 0.885 34.260 1.030 ;
    END
  END WBL_11
  PIN WBLb_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.369600 ;
    PORT
      LAYER li1 ;
        RECT 32.235 21.135 32.310 21.275 ;
        RECT 32.235 19.785 32.310 19.925 ;
        RECT 32.235 18.435 32.310 18.575 ;
        RECT 32.235 17.085 32.310 17.225 ;
        RECT 32.235 15.735 32.310 15.875 ;
        RECT 32.235 14.385 32.310 14.525 ;
        RECT 32.235 13.035 32.310 13.175 ;
        RECT 32.235 11.685 32.310 11.825 ;
        RECT 32.235 10.335 32.310 10.475 ;
        RECT 32.235 8.985 32.310 9.125 ;
        RECT 32.235 7.635 32.310 7.775 ;
        RECT 32.235 6.285 32.310 6.425 ;
        RECT 32.235 4.935 32.310 5.075 ;
        RECT 32.235 3.585 32.310 3.725 ;
        RECT 32.235 2.235 32.310 2.375 ;
        RECT 32.235 0.885 32.310 1.025 ;
    END
  END WBLb_11
  OBS
      LAYER li1 ;
        RECT 0.740 21.135 0.815 21.275 ;
        RECT 0.955 21.085 1.030 21.225 ;
        RECT 1.660 21.145 1.720 21.225 ;
        POLYGON 1.660 21.145 1.720 21.145 1.720 21.085 ;
        RECT 1.875 21.135 1.950 21.275 ;
        RECT 3.640 21.135 3.715 21.275 ;
        RECT 3.855 21.085 3.930 21.225 ;
        RECT 4.560 21.145 4.620 21.225 ;
        POLYGON 4.560 21.145 4.620 21.145 4.620 21.085 ;
        RECT 4.775 21.135 4.850 21.275 ;
        RECT 6.540 21.135 6.615 21.275 ;
        RECT 6.755 21.085 6.830 21.225 ;
        RECT 7.460 21.145 7.520 21.225 ;
        POLYGON 7.460 21.145 7.520 21.145 7.520 21.085 ;
        RECT 7.675 21.135 7.750 21.275 ;
        RECT 9.440 21.135 9.515 21.275 ;
        RECT 9.655 21.085 9.730 21.225 ;
        RECT 10.360 21.145 10.420 21.225 ;
        POLYGON 10.360 21.145 10.420 21.145 10.420 21.085 ;
        RECT 10.575 21.135 10.650 21.275 ;
        RECT 12.340 21.135 12.415 21.275 ;
        RECT 12.555 21.085 12.630 21.225 ;
        RECT 13.260 21.145 13.320 21.225 ;
        POLYGON 13.260 21.145 13.320 21.145 13.320 21.085 ;
        RECT 13.475 21.135 13.550 21.275 ;
        RECT 15.240 21.135 15.315 21.275 ;
        RECT 15.455 21.085 15.530 21.225 ;
        RECT 16.160 21.145 16.220 21.225 ;
        POLYGON 16.160 21.145 16.220 21.145 16.220 21.085 ;
        RECT 16.375 21.135 16.450 21.275 ;
        RECT 18.140 21.135 18.215 21.275 ;
        RECT 18.355 21.085 18.430 21.225 ;
        RECT 19.060 21.145 19.120 21.225 ;
        POLYGON 19.060 21.145 19.120 21.145 19.120 21.085 ;
        RECT 19.275 21.135 19.350 21.275 ;
        RECT 21.040 21.135 21.115 21.275 ;
        RECT 21.255 21.085 21.330 21.225 ;
        RECT 21.960 21.145 22.020 21.225 ;
        POLYGON 21.960 21.145 22.020 21.145 22.020 21.085 ;
        RECT 22.175 21.135 22.250 21.275 ;
        RECT 23.940 21.135 24.015 21.275 ;
        RECT 24.155 21.085 24.230 21.225 ;
        RECT 24.860 21.145 24.920 21.225 ;
        POLYGON 24.860 21.145 24.920 21.145 24.920 21.085 ;
        RECT 25.075 21.135 25.150 21.275 ;
        RECT 26.840 21.135 26.915 21.275 ;
        RECT 27.055 21.085 27.130 21.225 ;
        RECT 27.760 21.145 27.820 21.225 ;
        POLYGON 27.760 21.145 27.820 21.145 27.820 21.085 ;
        RECT 27.975 21.135 28.050 21.275 ;
        RECT 29.740 21.135 29.815 21.275 ;
        RECT 29.955 21.085 30.030 21.225 ;
        RECT 30.660 21.145 30.720 21.225 ;
        POLYGON 30.660 21.145 30.720 21.145 30.720 21.085 ;
        RECT 30.875 21.135 30.950 21.275 ;
        RECT 32.640 21.135 32.715 21.275 ;
        RECT 32.855 21.085 32.930 21.225 ;
        RECT 33.560 21.145 33.620 21.225 ;
        POLYGON 33.560 21.145 33.620 21.145 33.620 21.085 ;
        RECT 33.775 21.135 33.850 21.275 ;
        RECT 0.685 20.615 0.835 20.785 ;
        RECT 1.075 20.750 1.225 20.920 ;
        RECT 1.465 20.750 1.615 20.920 ;
        RECT 1.855 20.615 2.005 20.785 ;
        RECT 3.585 20.615 3.735 20.785 ;
        RECT 3.975 20.750 4.125 20.920 ;
        RECT 4.365 20.750 4.515 20.920 ;
        RECT 4.755 20.615 4.905 20.785 ;
        RECT 6.485 20.615 6.635 20.785 ;
        RECT 6.875 20.750 7.025 20.920 ;
        RECT 7.265 20.750 7.415 20.920 ;
        RECT 7.655 20.615 7.805 20.785 ;
        RECT 9.385 20.615 9.535 20.785 ;
        RECT 9.775 20.750 9.925 20.920 ;
        RECT 10.165 20.750 10.315 20.920 ;
        RECT 10.555 20.615 10.705 20.785 ;
        RECT 12.285 20.615 12.435 20.785 ;
        RECT 12.675 20.750 12.825 20.920 ;
        RECT 13.065 20.750 13.215 20.920 ;
        RECT 13.455 20.615 13.605 20.785 ;
        RECT 15.185 20.615 15.335 20.785 ;
        RECT 15.575 20.750 15.725 20.920 ;
        RECT 15.965 20.750 16.115 20.920 ;
        RECT 16.355 20.615 16.505 20.785 ;
        RECT 18.085 20.615 18.235 20.785 ;
        RECT 18.475 20.750 18.625 20.920 ;
        RECT 18.865 20.750 19.015 20.920 ;
        RECT 19.255 20.615 19.405 20.785 ;
        RECT 20.985 20.615 21.135 20.785 ;
        RECT 21.375 20.750 21.525 20.920 ;
        RECT 21.765 20.750 21.915 20.920 ;
        RECT 22.155 20.615 22.305 20.785 ;
        RECT 23.885 20.615 24.035 20.785 ;
        RECT 24.275 20.750 24.425 20.920 ;
        RECT 24.665 20.750 24.815 20.920 ;
        RECT 25.055 20.615 25.205 20.785 ;
        RECT 26.785 20.615 26.935 20.785 ;
        RECT 27.175 20.750 27.325 20.920 ;
        RECT 27.565 20.750 27.715 20.920 ;
        RECT 27.955 20.615 28.105 20.785 ;
        RECT 29.685 20.615 29.835 20.785 ;
        RECT 30.075 20.750 30.225 20.920 ;
        RECT 30.465 20.750 30.615 20.920 ;
        RECT 30.855 20.615 31.005 20.785 ;
        RECT 32.585 20.615 32.735 20.785 ;
        RECT 32.975 20.750 33.125 20.920 ;
        RECT 33.365 20.750 33.515 20.920 ;
        RECT 33.755 20.615 33.905 20.785 ;
        RECT 0.950 20.530 1.000 20.565 ;
        POLYGON 1.000 20.565 1.035 20.530 1.000 20.530 ;
        RECT 0.950 20.405 1.035 20.530 ;
        RECT 1.655 20.405 1.740 20.565 ;
        RECT 3.850 20.530 3.900 20.565 ;
        POLYGON 3.900 20.565 3.935 20.530 3.900 20.530 ;
        RECT 3.850 20.405 3.935 20.530 ;
        RECT 4.555 20.405 4.640 20.565 ;
        RECT 6.750 20.530 6.800 20.565 ;
        POLYGON 6.800 20.565 6.835 20.530 6.800 20.530 ;
        RECT 6.750 20.405 6.835 20.530 ;
        RECT 7.455 20.405 7.540 20.565 ;
        RECT 9.650 20.530 9.700 20.565 ;
        POLYGON 9.700 20.565 9.735 20.530 9.700 20.530 ;
        RECT 9.650 20.405 9.735 20.530 ;
        RECT 10.355 20.405 10.440 20.565 ;
        RECT 12.550 20.530 12.600 20.565 ;
        POLYGON 12.600 20.565 12.635 20.530 12.600 20.530 ;
        RECT 12.550 20.405 12.635 20.530 ;
        RECT 13.255 20.405 13.340 20.565 ;
        RECT 15.450 20.530 15.500 20.565 ;
        POLYGON 15.500 20.565 15.535 20.530 15.500 20.530 ;
        RECT 15.450 20.405 15.535 20.530 ;
        RECT 16.155 20.405 16.240 20.565 ;
        RECT 18.350 20.530 18.400 20.565 ;
        POLYGON 18.400 20.565 18.435 20.530 18.400 20.530 ;
        RECT 18.350 20.405 18.435 20.530 ;
        RECT 19.055 20.405 19.140 20.565 ;
        RECT 21.250 20.530 21.300 20.565 ;
        POLYGON 21.300 20.565 21.335 20.530 21.300 20.530 ;
        RECT 21.250 20.405 21.335 20.530 ;
        RECT 21.955 20.405 22.040 20.565 ;
        RECT 24.150 20.530 24.200 20.565 ;
        POLYGON 24.200 20.565 24.235 20.530 24.200 20.530 ;
        RECT 24.150 20.405 24.235 20.530 ;
        RECT 24.855 20.405 24.940 20.565 ;
        RECT 27.050 20.530 27.100 20.565 ;
        POLYGON 27.100 20.565 27.135 20.530 27.100 20.530 ;
        RECT 27.050 20.405 27.135 20.530 ;
        RECT 27.755 20.405 27.840 20.565 ;
        RECT 29.950 20.530 30.000 20.565 ;
        POLYGON 30.000 20.565 30.035 20.530 30.000 20.530 ;
        RECT 29.950 20.405 30.035 20.530 ;
        RECT 30.655 20.405 30.740 20.565 ;
        RECT 32.850 20.530 32.900 20.565 ;
        POLYGON 32.900 20.565 32.935 20.530 32.900 20.530 ;
        RECT 32.850 20.405 32.935 20.530 ;
        RECT 33.555 20.405 33.640 20.565 ;
        RECT 0.740 19.785 0.815 19.925 ;
        RECT 0.955 19.735 1.030 19.875 ;
        RECT 1.660 19.795 1.720 19.875 ;
        POLYGON 1.660 19.795 1.720 19.795 1.720 19.735 ;
        RECT 1.875 19.785 1.950 19.925 ;
        RECT 3.640 19.785 3.715 19.925 ;
        RECT 3.855 19.735 3.930 19.875 ;
        RECT 4.560 19.795 4.620 19.875 ;
        POLYGON 4.560 19.795 4.620 19.795 4.620 19.735 ;
        RECT 4.775 19.785 4.850 19.925 ;
        RECT 6.540 19.785 6.615 19.925 ;
        RECT 6.755 19.735 6.830 19.875 ;
        RECT 7.460 19.795 7.520 19.875 ;
        POLYGON 7.460 19.795 7.520 19.795 7.520 19.735 ;
        RECT 7.675 19.785 7.750 19.925 ;
        RECT 9.440 19.785 9.515 19.925 ;
        RECT 9.655 19.735 9.730 19.875 ;
        RECT 10.360 19.795 10.420 19.875 ;
        POLYGON 10.360 19.795 10.420 19.795 10.420 19.735 ;
        RECT 10.575 19.785 10.650 19.925 ;
        RECT 12.340 19.785 12.415 19.925 ;
        RECT 12.555 19.735 12.630 19.875 ;
        RECT 13.260 19.795 13.320 19.875 ;
        POLYGON 13.260 19.795 13.320 19.795 13.320 19.735 ;
        RECT 13.475 19.785 13.550 19.925 ;
        RECT 15.240 19.785 15.315 19.925 ;
        RECT 15.455 19.735 15.530 19.875 ;
        RECT 16.160 19.795 16.220 19.875 ;
        POLYGON 16.160 19.795 16.220 19.795 16.220 19.735 ;
        RECT 16.375 19.785 16.450 19.925 ;
        RECT 18.140 19.785 18.215 19.925 ;
        RECT 18.355 19.735 18.430 19.875 ;
        RECT 19.060 19.795 19.120 19.875 ;
        POLYGON 19.060 19.795 19.120 19.795 19.120 19.735 ;
        RECT 19.275 19.785 19.350 19.925 ;
        RECT 21.040 19.785 21.115 19.925 ;
        RECT 21.255 19.735 21.330 19.875 ;
        RECT 21.960 19.795 22.020 19.875 ;
        POLYGON 21.960 19.795 22.020 19.795 22.020 19.735 ;
        RECT 22.175 19.785 22.250 19.925 ;
        RECT 23.940 19.785 24.015 19.925 ;
        RECT 24.155 19.735 24.230 19.875 ;
        RECT 24.860 19.795 24.920 19.875 ;
        POLYGON 24.860 19.795 24.920 19.795 24.920 19.735 ;
        RECT 25.075 19.785 25.150 19.925 ;
        RECT 26.840 19.785 26.915 19.925 ;
        RECT 27.055 19.735 27.130 19.875 ;
        RECT 27.760 19.795 27.820 19.875 ;
        POLYGON 27.760 19.795 27.820 19.795 27.820 19.735 ;
        RECT 27.975 19.785 28.050 19.925 ;
        RECT 29.740 19.785 29.815 19.925 ;
        RECT 29.955 19.735 30.030 19.875 ;
        RECT 30.660 19.795 30.720 19.875 ;
        POLYGON 30.660 19.795 30.720 19.795 30.720 19.735 ;
        RECT 30.875 19.785 30.950 19.925 ;
        RECT 32.640 19.785 32.715 19.925 ;
        RECT 32.855 19.735 32.930 19.875 ;
        RECT 33.560 19.795 33.620 19.875 ;
        POLYGON 33.560 19.795 33.620 19.795 33.620 19.735 ;
        RECT 33.775 19.785 33.850 19.925 ;
        RECT 0.685 19.265 0.835 19.435 ;
        RECT 1.075 19.400 1.225 19.570 ;
        RECT 1.465 19.400 1.615 19.570 ;
        RECT 1.855 19.265 2.005 19.435 ;
        RECT 3.585 19.265 3.735 19.435 ;
        RECT 3.975 19.400 4.125 19.570 ;
        RECT 4.365 19.400 4.515 19.570 ;
        RECT 4.755 19.265 4.905 19.435 ;
        RECT 6.485 19.265 6.635 19.435 ;
        RECT 6.875 19.400 7.025 19.570 ;
        RECT 7.265 19.400 7.415 19.570 ;
        RECT 7.655 19.265 7.805 19.435 ;
        RECT 9.385 19.265 9.535 19.435 ;
        RECT 9.775 19.400 9.925 19.570 ;
        RECT 10.165 19.400 10.315 19.570 ;
        RECT 10.555 19.265 10.705 19.435 ;
        RECT 12.285 19.265 12.435 19.435 ;
        RECT 12.675 19.400 12.825 19.570 ;
        RECT 13.065 19.400 13.215 19.570 ;
        RECT 13.455 19.265 13.605 19.435 ;
        RECT 15.185 19.265 15.335 19.435 ;
        RECT 15.575 19.400 15.725 19.570 ;
        RECT 15.965 19.400 16.115 19.570 ;
        RECT 16.355 19.265 16.505 19.435 ;
        RECT 18.085 19.265 18.235 19.435 ;
        RECT 18.475 19.400 18.625 19.570 ;
        RECT 18.865 19.400 19.015 19.570 ;
        RECT 19.255 19.265 19.405 19.435 ;
        RECT 20.985 19.265 21.135 19.435 ;
        RECT 21.375 19.400 21.525 19.570 ;
        RECT 21.765 19.400 21.915 19.570 ;
        RECT 22.155 19.265 22.305 19.435 ;
        RECT 23.885 19.265 24.035 19.435 ;
        RECT 24.275 19.400 24.425 19.570 ;
        RECT 24.665 19.400 24.815 19.570 ;
        RECT 25.055 19.265 25.205 19.435 ;
        RECT 26.785 19.265 26.935 19.435 ;
        RECT 27.175 19.400 27.325 19.570 ;
        RECT 27.565 19.400 27.715 19.570 ;
        RECT 27.955 19.265 28.105 19.435 ;
        RECT 29.685 19.265 29.835 19.435 ;
        RECT 30.075 19.400 30.225 19.570 ;
        RECT 30.465 19.400 30.615 19.570 ;
        RECT 30.855 19.265 31.005 19.435 ;
        RECT 32.585 19.265 32.735 19.435 ;
        RECT 32.975 19.400 33.125 19.570 ;
        RECT 33.365 19.400 33.515 19.570 ;
        RECT 33.755 19.265 33.905 19.435 ;
        RECT 0.950 19.180 1.000 19.215 ;
        POLYGON 1.000 19.215 1.035 19.180 1.000 19.180 ;
        RECT 0.950 19.055 1.035 19.180 ;
        RECT 1.655 19.055 1.740 19.215 ;
        RECT 3.850 19.180 3.900 19.215 ;
        POLYGON 3.900 19.215 3.935 19.180 3.900 19.180 ;
        RECT 3.850 19.055 3.935 19.180 ;
        RECT 4.555 19.055 4.640 19.215 ;
        RECT 6.750 19.180 6.800 19.215 ;
        POLYGON 6.800 19.215 6.835 19.180 6.800 19.180 ;
        RECT 6.750 19.055 6.835 19.180 ;
        RECT 7.455 19.055 7.540 19.215 ;
        RECT 9.650 19.180 9.700 19.215 ;
        POLYGON 9.700 19.215 9.735 19.180 9.700 19.180 ;
        RECT 9.650 19.055 9.735 19.180 ;
        RECT 10.355 19.055 10.440 19.215 ;
        RECT 12.550 19.180 12.600 19.215 ;
        POLYGON 12.600 19.215 12.635 19.180 12.600 19.180 ;
        RECT 12.550 19.055 12.635 19.180 ;
        RECT 13.255 19.055 13.340 19.215 ;
        RECT 15.450 19.180 15.500 19.215 ;
        POLYGON 15.500 19.215 15.535 19.180 15.500 19.180 ;
        RECT 15.450 19.055 15.535 19.180 ;
        RECT 16.155 19.055 16.240 19.215 ;
        RECT 18.350 19.180 18.400 19.215 ;
        POLYGON 18.400 19.215 18.435 19.180 18.400 19.180 ;
        RECT 18.350 19.055 18.435 19.180 ;
        RECT 19.055 19.055 19.140 19.215 ;
        RECT 21.250 19.180 21.300 19.215 ;
        POLYGON 21.300 19.215 21.335 19.180 21.300 19.180 ;
        RECT 21.250 19.055 21.335 19.180 ;
        RECT 21.955 19.055 22.040 19.215 ;
        RECT 24.150 19.180 24.200 19.215 ;
        POLYGON 24.200 19.215 24.235 19.180 24.200 19.180 ;
        RECT 24.150 19.055 24.235 19.180 ;
        RECT 24.855 19.055 24.940 19.215 ;
        RECT 27.050 19.180 27.100 19.215 ;
        POLYGON 27.100 19.215 27.135 19.180 27.100 19.180 ;
        RECT 27.050 19.055 27.135 19.180 ;
        RECT 27.755 19.055 27.840 19.215 ;
        RECT 29.950 19.180 30.000 19.215 ;
        POLYGON 30.000 19.215 30.035 19.180 30.000 19.180 ;
        RECT 29.950 19.055 30.035 19.180 ;
        RECT 30.655 19.055 30.740 19.215 ;
        RECT 32.850 19.180 32.900 19.215 ;
        POLYGON 32.900 19.215 32.935 19.180 32.900 19.180 ;
        RECT 32.850 19.055 32.935 19.180 ;
        RECT 33.555 19.055 33.640 19.215 ;
        RECT 0.740 18.435 0.815 18.575 ;
        RECT 0.955 18.385 1.030 18.525 ;
        RECT 1.660 18.445 1.720 18.525 ;
        POLYGON 1.660 18.445 1.720 18.445 1.720 18.385 ;
        RECT 1.875 18.435 1.950 18.575 ;
        RECT 3.640 18.435 3.715 18.575 ;
        RECT 3.855 18.385 3.930 18.525 ;
        RECT 4.560 18.445 4.620 18.525 ;
        POLYGON 4.560 18.445 4.620 18.445 4.620 18.385 ;
        RECT 4.775 18.435 4.850 18.575 ;
        RECT 6.540 18.435 6.615 18.575 ;
        RECT 6.755 18.385 6.830 18.525 ;
        RECT 7.460 18.445 7.520 18.525 ;
        POLYGON 7.460 18.445 7.520 18.445 7.520 18.385 ;
        RECT 7.675 18.435 7.750 18.575 ;
        RECT 9.440 18.435 9.515 18.575 ;
        RECT 9.655 18.385 9.730 18.525 ;
        RECT 10.360 18.445 10.420 18.525 ;
        POLYGON 10.360 18.445 10.420 18.445 10.420 18.385 ;
        RECT 10.575 18.435 10.650 18.575 ;
        RECT 12.340 18.435 12.415 18.575 ;
        RECT 12.555 18.385 12.630 18.525 ;
        RECT 13.260 18.445 13.320 18.525 ;
        POLYGON 13.260 18.445 13.320 18.445 13.320 18.385 ;
        RECT 13.475 18.435 13.550 18.575 ;
        RECT 15.240 18.435 15.315 18.575 ;
        RECT 15.455 18.385 15.530 18.525 ;
        RECT 16.160 18.445 16.220 18.525 ;
        POLYGON 16.160 18.445 16.220 18.445 16.220 18.385 ;
        RECT 16.375 18.435 16.450 18.575 ;
        RECT 18.140 18.435 18.215 18.575 ;
        RECT 18.355 18.385 18.430 18.525 ;
        RECT 19.060 18.445 19.120 18.525 ;
        POLYGON 19.060 18.445 19.120 18.445 19.120 18.385 ;
        RECT 19.275 18.435 19.350 18.575 ;
        RECT 21.040 18.435 21.115 18.575 ;
        RECT 21.255 18.385 21.330 18.525 ;
        RECT 21.960 18.445 22.020 18.525 ;
        POLYGON 21.960 18.445 22.020 18.445 22.020 18.385 ;
        RECT 22.175 18.435 22.250 18.575 ;
        RECT 23.940 18.435 24.015 18.575 ;
        RECT 24.155 18.385 24.230 18.525 ;
        RECT 24.860 18.445 24.920 18.525 ;
        POLYGON 24.860 18.445 24.920 18.445 24.920 18.385 ;
        RECT 25.075 18.435 25.150 18.575 ;
        RECT 26.840 18.435 26.915 18.575 ;
        RECT 27.055 18.385 27.130 18.525 ;
        RECT 27.760 18.445 27.820 18.525 ;
        POLYGON 27.760 18.445 27.820 18.445 27.820 18.385 ;
        RECT 27.975 18.435 28.050 18.575 ;
        RECT 29.740 18.435 29.815 18.575 ;
        RECT 29.955 18.385 30.030 18.525 ;
        RECT 30.660 18.445 30.720 18.525 ;
        POLYGON 30.660 18.445 30.720 18.445 30.720 18.385 ;
        RECT 30.875 18.435 30.950 18.575 ;
        RECT 32.640 18.435 32.715 18.575 ;
        RECT 32.855 18.385 32.930 18.525 ;
        RECT 33.560 18.445 33.620 18.525 ;
        POLYGON 33.560 18.445 33.620 18.445 33.620 18.385 ;
        RECT 33.775 18.435 33.850 18.575 ;
        RECT 0.685 17.915 0.835 18.085 ;
        RECT 1.075 18.050 1.225 18.220 ;
        RECT 1.465 18.050 1.615 18.220 ;
        RECT 1.855 17.915 2.005 18.085 ;
        RECT 3.585 17.915 3.735 18.085 ;
        RECT 3.975 18.050 4.125 18.220 ;
        RECT 4.365 18.050 4.515 18.220 ;
        RECT 4.755 17.915 4.905 18.085 ;
        RECT 6.485 17.915 6.635 18.085 ;
        RECT 6.875 18.050 7.025 18.220 ;
        RECT 7.265 18.050 7.415 18.220 ;
        RECT 7.655 17.915 7.805 18.085 ;
        RECT 9.385 17.915 9.535 18.085 ;
        RECT 9.775 18.050 9.925 18.220 ;
        RECT 10.165 18.050 10.315 18.220 ;
        RECT 10.555 17.915 10.705 18.085 ;
        RECT 12.285 17.915 12.435 18.085 ;
        RECT 12.675 18.050 12.825 18.220 ;
        RECT 13.065 18.050 13.215 18.220 ;
        RECT 13.455 17.915 13.605 18.085 ;
        RECT 15.185 17.915 15.335 18.085 ;
        RECT 15.575 18.050 15.725 18.220 ;
        RECT 15.965 18.050 16.115 18.220 ;
        RECT 16.355 17.915 16.505 18.085 ;
        RECT 18.085 17.915 18.235 18.085 ;
        RECT 18.475 18.050 18.625 18.220 ;
        RECT 18.865 18.050 19.015 18.220 ;
        RECT 19.255 17.915 19.405 18.085 ;
        RECT 20.985 17.915 21.135 18.085 ;
        RECT 21.375 18.050 21.525 18.220 ;
        RECT 21.765 18.050 21.915 18.220 ;
        RECT 22.155 17.915 22.305 18.085 ;
        RECT 23.885 17.915 24.035 18.085 ;
        RECT 24.275 18.050 24.425 18.220 ;
        RECT 24.665 18.050 24.815 18.220 ;
        RECT 25.055 17.915 25.205 18.085 ;
        RECT 26.785 17.915 26.935 18.085 ;
        RECT 27.175 18.050 27.325 18.220 ;
        RECT 27.565 18.050 27.715 18.220 ;
        RECT 27.955 17.915 28.105 18.085 ;
        RECT 29.685 17.915 29.835 18.085 ;
        RECT 30.075 18.050 30.225 18.220 ;
        RECT 30.465 18.050 30.615 18.220 ;
        RECT 30.855 17.915 31.005 18.085 ;
        RECT 32.585 17.915 32.735 18.085 ;
        RECT 32.975 18.050 33.125 18.220 ;
        RECT 33.365 18.050 33.515 18.220 ;
        RECT 33.755 17.915 33.905 18.085 ;
        RECT 0.950 17.830 1.000 17.865 ;
        POLYGON 1.000 17.865 1.035 17.830 1.000 17.830 ;
        RECT 0.950 17.705 1.035 17.830 ;
        RECT 1.655 17.705 1.740 17.865 ;
        RECT 3.850 17.830 3.900 17.865 ;
        POLYGON 3.900 17.865 3.935 17.830 3.900 17.830 ;
        RECT 3.850 17.705 3.935 17.830 ;
        RECT 4.555 17.705 4.640 17.865 ;
        RECT 6.750 17.830 6.800 17.865 ;
        POLYGON 6.800 17.865 6.835 17.830 6.800 17.830 ;
        RECT 6.750 17.705 6.835 17.830 ;
        RECT 7.455 17.705 7.540 17.865 ;
        RECT 9.650 17.830 9.700 17.865 ;
        POLYGON 9.700 17.865 9.735 17.830 9.700 17.830 ;
        RECT 9.650 17.705 9.735 17.830 ;
        RECT 10.355 17.705 10.440 17.865 ;
        RECT 12.550 17.830 12.600 17.865 ;
        POLYGON 12.600 17.865 12.635 17.830 12.600 17.830 ;
        RECT 12.550 17.705 12.635 17.830 ;
        RECT 13.255 17.705 13.340 17.865 ;
        RECT 15.450 17.830 15.500 17.865 ;
        POLYGON 15.500 17.865 15.535 17.830 15.500 17.830 ;
        RECT 15.450 17.705 15.535 17.830 ;
        RECT 16.155 17.705 16.240 17.865 ;
        RECT 18.350 17.830 18.400 17.865 ;
        POLYGON 18.400 17.865 18.435 17.830 18.400 17.830 ;
        RECT 18.350 17.705 18.435 17.830 ;
        RECT 19.055 17.705 19.140 17.865 ;
        RECT 21.250 17.830 21.300 17.865 ;
        POLYGON 21.300 17.865 21.335 17.830 21.300 17.830 ;
        RECT 21.250 17.705 21.335 17.830 ;
        RECT 21.955 17.705 22.040 17.865 ;
        RECT 24.150 17.830 24.200 17.865 ;
        POLYGON 24.200 17.865 24.235 17.830 24.200 17.830 ;
        RECT 24.150 17.705 24.235 17.830 ;
        RECT 24.855 17.705 24.940 17.865 ;
        RECT 27.050 17.830 27.100 17.865 ;
        POLYGON 27.100 17.865 27.135 17.830 27.100 17.830 ;
        RECT 27.050 17.705 27.135 17.830 ;
        RECT 27.755 17.705 27.840 17.865 ;
        RECT 29.950 17.830 30.000 17.865 ;
        POLYGON 30.000 17.865 30.035 17.830 30.000 17.830 ;
        RECT 29.950 17.705 30.035 17.830 ;
        RECT 30.655 17.705 30.740 17.865 ;
        RECT 32.850 17.830 32.900 17.865 ;
        POLYGON 32.900 17.865 32.935 17.830 32.900 17.830 ;
        RECT 32.850 17.705 32.935 17.830 ;
        RECT 33.555 17.705 33.640 17.865 ;
        RECT 0.740 17.085 0.815 17.225 ;
        RECT 0.955 17.035 1.030 17.175 ;
        RECT 1.660 17.095 1.720 17.175 ;
        POLYGON 1.660 17.095 1.720 17.095 1.720 17.035 ;
        RECT 1.875 17.085 1.950 17.225 ;
        RECT 3.640 17.085 3.715 17.225 ;
        RECT 3.855 17.035 3.930 17.175 ;
        RECT 4.560 17.095 4.620 17.175 ;
        POLYGON 4.560 17.095 4.620 17.095 4.620 17.035 ;
        RECT 4.775 17.085 4.850 17.225 ;
        RECT 6.540 17.085 6.615 17.225 ;
        RECT 6.755 17.035 6.830 17.175 ;
        RECT 7.460 17.095 7.520 17.175 ;
        POLYGON 7.460 17.095 7.520 17.095 7.520 17.035 ;
        RECT 7.675 17.085 7.750 17.225 ;
        RECT 9.440 17.085 9.515 17.225 ;
        RECT 9.655 17.035 9.730 17.175 ;
        RECT 10.360 17.095 10.420 17.175 ;
        POLYGON 10.360 17.095 10.420 17.095 10.420 17.035 ;
        RECT 10.575 17.085 10.650 17.225 ;
        RECT 12.340 17.085 12.415 17.225 ;
        RECT 12.555 17.035 12.630 17.175 ;
        RECT 13.260 17.095 13.320 17.175 ;
        POLYGON 13.260 17.095 13.320 17.095 13.320 17.035 ;
        RECT 13.475 17.085 13.550 17.225 ;
        RECT 15.240 17.085 15.315 17.225 ;
        RECT 15.455 17.035 15.530 17.175 ;
        RECT 16.160 17.095 16.220 17.175 ;
        POLYGON 16.160 17.095 16.220 17.095 16.220 17.035 ;
        RECT 16.375 17.085 16.450 17.225 ;
        RECT 18.140 17.085 18.215 17.225 ;
        RECT 18.355 17.035 18.430 17.175 ;
        RECT 19.060 17.095 19.120 17.175 ;
        POLYGON 19.060 17.095 19.120 17.095 19.120 17.035 ;
        RECT 19.275 17.085 19.350 17.225 ;
        RECT 21.040 17.085 21.115 17.225 ;
        RECT 21.255 17.035 21.330 17.175 ;
        RECT 21.960 17.095 22.020 17.175 ;
        POLYGON 21.960 17.095 22.020 17.095 22.020 17.035 ;
        RECT 22.175 17.085 22.250 17.225 ;
        RECT 23.940 17.085 24.015 17.225 ;
        RECT 24.155 17.035 24.230 17.175 ;
        RECT 24.860 17.095 24.920 17.175 ;
        POLYGON 24.860 17.095 24.920 17.095 24.920 17.035 ;
        RECT 25.075 17.085 25.150 17.225 ;
        RECT 26.840 17.085 26.915 17.225 ;
        RECT 27.055 17.035 27.130 17.175 ;
        RECT 27.760 17.095 27.820 17.175 ;
        POLYGON 27.760 17.095 27.820 17.095 27.820 17.035 ;
        RECT 27.975 17.085 28.050 17.225 ;
        RECT 29.740 17.085 29.815 17.225 ;
        RECT 29.955 17.035 30.030 17.175 ;
        RECT 30.660 17.095 30.720 17.175 ;
        POLYGON 30.660 17.095 30.720 17.095 30.720 17.035 ;
        RECT 30.875 17.085 30.950 17.225 ;
        RECT 32.640 17.085 32.715 17.225 ;
        RECT 32.855 17.035 32.930 17.175 ;
        RECT 33.560 17.095 33.620 17.175 ;
        POLYGON 33.560 17.095 33.620 17.095 33.620 17.035 ;
        RECT 33.775 17.085 33.850 17.225 ;
        RECT 0.685 16.565 0.835 16.735 ;
        RECT 1.075 16.700 1.225 16.870 ;
        RECT 1.465 16.700 1.615 16.870 ;
        RECT 1.855 16.565 2.005 16.735 ;
        RECT 3.585 16.565 3.735 16.735 ;
        RECT 3.975 16.700 4.125 16.870 ;
        RECT 4.365 16.700 4.515 16.870 ;
        RECT 4.755 16.565 4.905 16.735 ;
        RECT 6.485 16.565 6.635 16.735 ;
        RECT 6.875 16.700 7.025 16.870 ;
        RECT 7.265 16.700 7.415 16.870 ;
        RECT 7.655 16.565 7.805 16.735 ;
        RECT 9.385 16.565 9.535 16.735 ;
        RECT 9.775 16.700 9.925 16.870 ;
        RECT 10.165 16.700 10.315 16.870 ;
        RECT 10.555 16.565 10.705 16.735 ;
        RECT 12.285 16.565 12.435 16.735 ;
        RECT 12.675 16.700 12.825 16.870 ;
        RECT 13.065 16.700 13.215 16.870 ;
        RECT 13.455 16.565 13.605 16.735 ;
        RECT 15.185 16.565 15.335 16.735 ;
        RECT 15.575 16.700 15.725 16.870 ;
        RECT 15.965 16.700 16.115 16.870 ;
        RECT 16.355 16.565 16.505 16.735 ;
        RECT 18.085 16.565 18.235 16.735 ;
        RECT 18.475 16.700 18.625 16.870 ;
        RECT 18.865 16.700 19.015 16.870 ;
        RECT 19.255 16.565 19.405 16.735 ;
        RECT 20.985 16.565 21.135 16.735 ;
        RECT 21.375 16.700 21.525 16.870 ;
        RECT 21.765 16.700 21.915 16.870 ;
        RECT 22.155 16.565 22.305 16.735 ;
        RECT 23.885 16.565 24.035 16.735 ;
        RECT 24.275 16.700 24.425 16.870 ;
        RECT 24.665 16.700 24.815 16.870 ;
        RECT 25.055 16.565 25.205 16.735 ;
        RECT 26.785 16.565 26.935 16.735 ;
        RECT 27.175 16.700 27.325 16.870 ;
        RECT 27.565 16.700 27.715 16.870 ;
        RECT 27.955 16.565 28.105 16.735 ;
        RECT 29.685 16.565 29.835 16.735 ;
        RECT 30.075 16.700 30.225 16.870 ;
        RECT 30.465 16.700 30.615 16.870 ;
        RECT 30.855 16.565 31.005 16.735 ;
        RECT 32.585 16.565 32.735 16.735 ;
        RECT 32.975 16.700 33.125 16.870 ;
        RECT 33.365 16.700 33.515 16.870 ;
        RECT 33.755 16.565 33.905 16.735 ;
        RECT 0.950 16.480 1.000 16.515 ;
        POLYGON 1.000 16.515 1.035 16.480 1.000 16.480 ;
        RECT 0.950 16.355 1.035 16.480 ;
        RECT 1.655 16.355 1.740 16.515 ;
        RECT 3.850 16.480 3.900 16.515 ;
        POLYGON 3.900 16.515 3.935 16.480 3.900 16.480 ;
        RECT 3.850 16.355 3.935 16.480 ;
        RECT 4.555 16.355 4.640 16.515 ;
        RECT 6.750 16.480 6.800 16.515 ;
        POLYGON 6.800 16.515 6.835 16.480 6.800 16.480 ;
        RECT 6.750 16.355 6.835 16.480 ;
        RECT 7.455 16.355 7.540 16.515 ;
        RECT 9.650 16.480 9.700 16.515 ;
        POLYGON 9.700 16.515 9.735 16.480 9.700 16.480 ;
        RECT 9.650 16.355 9.735 16.480 ;
        RECT 10.355 16.355 10.440 16.515 ;
        RECT 12.550 16.480 12.600 16.515 ;
        POLYGON 12.600 16.515 12.635 16.480 12.600 16.480 ;
        RECT 12.550 16.355 12.635 16.480 ;
        RECT 13.255 16.355 13.340 16.515 ;
        RECT 15.450 16.480 15.500 16.515 ;
        POLYGON 15.500 16.515 15.535 16.480 15.500 16.480 ;
        RECT 15.450 16.355 15.535 16.480 ;
        RECT 16.155 16.355 16.240 16.515 ;
        RECT 18.350 16.480 18.400 16.515 ;
        POLYGON 18.400 16.515 18.435 16.480 18.400 16.480 ;
        RECT 18.350 16.355 18.435 16.480 ;
        RECT 19.055 16.355 19.140 16.515 ;
        RECT 21.250 16.480 21.300 16.515 ;
        POLYGON 21.300 16.515 21.335 16.480 21.300 16.480 ;
        RECT 21.250 16.355 21.335 16.480 ;
        RECT 21.955 16.355 22.040 16.515 ;
        RECT 24.150 16.480 24.200 16.515 ;
        POLYGON 24.200 16.515 24.235 16.480 24.200 16.480 ;
        RECT 24.150 16.355 24.235 16.480 ;
        RECT 24.855 16.355 24.940 16.515 ;
        RECT 27.050 16.480 27.100 16.515 ;
        POLYGON 27.100 16.515 27.135 16.480 27.100 16.480 ;
        RECT 27.050 16.355 27.135 16.480 ;
        RECT 27.755 16.355 27.840 16.515 ;
        RECT 29.950 16.480 30.000 16.515 ;
        POLYGON 30.000 16.515 30.035 16.480 30.000 16.480 ;
        RECT 29.950 16.355 30.035 16.480 ;
        RECT 30.655 16.355 30.740 16.515 ;
        RECT 32.850 16.480 32.900 16.515 ;
        POLYGON 32.900 16.515 32.935 16.480 32.900 16.480 ;
        RECT 32.850 16.355 32.935 16.480 ;
        RECT 33.555 16.355 33.640 16.515 ;
        RECT 0.740 15.735 0.815 15.875 ;
        RECT 0.955 15.685 1.030 15.825 ;
        RECT 1.660 15.745 1.720 15.825 ;
        POLYGON 1.660 15.745 1.720 15.745 1.720 15.685 ;
        RECT 1.875 15.735 1.950 15.875 ;
        RECT 3.640 15.735 3.715 15.875 ;
        RECT 3.855 15.685 3.930 15.825 ;
        RECT 4.560 15.745 4.620 15.825 ;
        POLYGON 4.560 15.745 4.620 15.745 4.620 15.685 ;
        RECT 4.775 15.735 4.850 15.875 ;
        RECT 6.540 15.735 6.615 15.875 ;
        RECT 6.755 15.685 6.830 15.825 ;
        RECT 7.460 15.745 7.520 15.825 ;
        POLYGON 7.460 15.745 7.520 15.745 7.520 15.685 ;
        RECT 7.675 15.735 7.750 15.875 ;
        RECT 9.440 15.735 9.515 15.875 ;
        RECT 9.655 15.685 9.730 15.825 ;
        RECT 10.360 15.745 10.420 15.825 ;
        POLYGON 10.360 15.745 10.420 15.745 10.420 15.685 ;
        RECT 10.575 15.735 10.650 15.875 ;
        RECT 12.340 15.735 12.415 15.875 ;
        RECT 12.555 15.685 12.630 15.825 ;
        RECT 13.260 15.745 13.320 15.825 ;
        POLYGON 13.260 15.745 13.320 15.745 13.320 15.685 ;
        RECT 13.475 15.735 13.550 15.875 ;
        RECT 15.240 15.735 15.315 15.875 ;
        RECT 15.455 15.685 15.530 15.825 ;
        RECT 16.160 15.745 16.220 15.825 ;
        POLYGON 16.160 15.745 16.220 15.745 16.220 15.685 ;
        RECT 16.375 15.735 16.450 15.875 ;
        RECT 18.140 15.735 18.215 15.875 ;
        RECT 18.355 15.685 18.430 15.825 ;
        RECT 19.060 15.745 19.120 15.825 ;
        POLYGON 19.060 15.745 19.120 15.745 19.120 15.685 ;
        RECT 19.275 15.735 19.350 15.875 ;
        RECT 21.040 15.735 21.115 15.875 ;
        RECT 21.255 15.685 21.330 15.825 ;
        RECT 21.960 15.745 22.020 15.825 ;
        POLYGON 21.960 15.745 22.020 15.745 22.020 15.685 ;
        RECT 22.175 15.735 22.250 15.875 ;
        RECT 23.940 15.735 24.015 15.875 ;
        RECT 24.155 15.685 24.230 15.825 ;
        RECT 24.860 15.745 24.920 15.825 ;
        POLYGON 24.860 15.745 24.920 15.745 24.920 15.685 ;
        RECT 25.075 15.735 25.150 15.875 ;
        RECT 26.840 15.735 26.915 15.875 ;
        RECT 27.055 15.685 27.130 15.825 ;
        RECT 27.760 15.745 27.820 15.825 ;
        POLYGON 27.760 15.745 27.820 15.745 27.820 15.685 ;
        RECT 27.975 15.735 28.050 15.875 ;
        RECT 29.740 15.735 29.815 15.875 ;
        RECT 29.955 15.685 30.030 15.825 ;
        RECT 30.660 15.745 30.720 15.825 ;
        POLYGON 30.660 15.745 30.720 15.745 30.720 15.685 ;
        RECT 30.875 15.735 30.950 15.875 ;
        RECT 32.640 15.735 32.715 15.875 ;
        RECT 32.855 15.685 32.930 15.825 ;
        RECT 33.560 15.745 33.620 15.825 ;
        POLYGON 33.560 15.745 33.620 15.745 33.620 15.685 ;
        RECT 33.775 15.735 33.850 15.875 ;
        RECT 0.685 15.215 0.835 15.385 ;
        RECT 1.075 15.350 1.225 15.520 ;
        RECT 1.465 15.350 1.615 15.520 ;
        RECT 1.855 15.215 2.005 15.385 ;
        RECT 3.585 15.215 3.735 15.385 ;
        RECT 3.975 15.350 4.125 15.520 ;
        RECT 4.365 15.350 4.515 15.520 ;
        RECT 4.755 15.215 4.905 15.385 ;
        RECT 6.485 15.215 6.635 15.385 ;
        RECT 6.875 15.350 7.025 15.520 ;
        RECT 7.265 15.350 7.415 15.520 ;
        RECT 7.655 15.215 7.805 15.385 ;
        RECT 9.385 15.215 9.535 15.385 ;
        RECT 9.775 15.350 9.925 15.520 ;
        RECT 10.165 15.350 10.315 15.520 ;
        RECT 10.555 15.215 10.705 15.385 ;
        RECT 12.285 15.215 12.435 15.385 ;
        RECT 12.675 15.350 12.825 15.520 ;
        RECT 13.065 15.350 13.215 15.520 ;
        RECT 13.455 15.215 13.605 15.385 ;
        RECT 15.185 15.215 15.335 15.385 ;
        RECT 15.575 15.350 15.725 15.520 ;
        RECT 15.965 15.350 16.115 15.520 ;
        RECT 16.355 15.215 16.505 15.385 ;
        RECT 18.085 15.215 18.235 15.385 ;
        RECT 18.475 15.350 18.625 15.520 ;
        RECT 18.865 15.350 19.015 15.520 ;
        RECT 19.255 15.215 19.405 15.385 ;
        RECT 20.985 15.215 21.135 15.385 ;
        RECT 21.375 15.350 21.525 15.520 ;
        RECT 21.765 15.350 21.915 15.520 ;
        RECT 22.155 15.215 22.305 15.385 ;
        RECT 23.885 15.215 24.035 15.385 ;
        RECT 24.275 15.350 24.425 15.520 ;
        RECT 24.665 15.350 24.815 15.520 ;
        RECT 25.055 15.215 25.205 15.385 ;
        RECT 26.785 15.215 26.935 15.385 ;
        RECT 27.175 15.350 27.325 15.520 ;
        RECT 27.565 15.350 27.715 15.520 ;
        RECT 27.955 15.215 28.105 15.385 ;
        RECT 29.685 15.215 29.835 15.385 ;
        RECT 30.075 15.350 30.225 15.520 ;
        RECT 30.465 15.350 30.615 15.520 ;
        RECT 30.855 15.215 31.005 15.385 ;
        RECT 32.585 15.215 32.735 15.385 ;
        RECT 32.975 15.350 33.125 15.520 ;
        RECT 33.365 15.350 33.515 15.520 ;
        RECT 33.755 15.215 33.905 15.385 ;
        RECT 0.950 15.130 1.000 15.165 ;
        POLYGON 1.000 15.165 1.035 15.130 1.000 15.130 ;
        RECT 0.950 15.005 1.035 15.130 ;
        RECT 1.655 15.005 1.740 15.165 ;
        RECT 3.850 15.130 3.900 15.165 ;
        POLYGON 3.900 15.165 3.935 15.130 3.900 15.130 ;
        RECT 3.850 15.005 3.935 15.130 ;
        RECT 4.555 15.005 4.640 15.165 ;
        RECT 6.750 15.130 6.800 15.165 ;
        POLYGON 6.800 15.165 6.835 15.130 6.800 15.130 ;
        RECT 6.750 15.005 6.835 15.130 ;
        RECT 7.455 15.005 7.540 15.165 ;
        RECT 9.650 15.130 9.700 15.165 ;
        POLYGON 9.700 15.165 9.735 15.130 9.700 15.130 ;
        RECT 9.650 15.005 9.735 15.130 ;
        RECT 10.355 15.005 10.440 15.165 ;
        RECT 12.550 15.130 12.600 15.165 ;
        POLYGON 12.600 15.165 12.635 15.130 12.600 15.130 ;
        RECT 12.550 15.005 12.635 15.130 ;
        RECT 13.255 15.005 13.340 15.165 ;
        RECT 15.450 15.130 15.500 15.165 ;
        POLYGON 15.500 15.165 15.535 15.130 15.500 15.130 ;
        RECT 15.450 15.005 15.535 15.130 ;
        RECT 16.155 15.005 16.240 15.165 ;
        RECT 18.350 15.130 18.400 15.165 ;
        POLYGON 18.400 15.165 18.435 15.130 18.400 15.130 ;
        RECT 18.350 15.005 18.435 15.130 ;
        RECT 19.055 15.005 19.140 15.165 ;
        RECT 21.250 15.130 21.300 15.165 ;
        POLYGON 21.300 15.165 21.335 15.130 21.300 15.130 ;
        RECT 21.250 15.005 21.335 15.130 ;
        RECT 21.955 15.005 22.040 15.165 ;
        RECT 24.150 15.130 24.200 15.165 ;
        POLYGON 24.200 15.165 24.235 15.130 24.200 15.130 ;
        RECT 24.150 15.005 24.235 15.130 ;
        RECT 24.855 15.005 24.940 15.165 ;
        RECT 27.050 15.130 27.100 15.165 ;
        POLYGON 27.100 15.165 27.135 15.130 27.100 15.130 ;
        RECT 27.050 15.005 27.135 15.130 ;
        RECT 27.755 15.005 27.840 15.165 ;
        RECT 29.950 15.130 30.000 15.165 ;
        POLYGON 30.000 15.165 30.035 15.130 30.000 15.130 ;
        RECT 29.950 15.005 30.035 15.130 ;
        RECT 30.655 15.005 30.740 15.165 ;
        RECT 32.850 15.130 32.900 15.165 ;
        POLYGON 32.900 15.165 32.935 15.130 32.900 15.130 ;
        RECT 32.850 15.005 32.935 15.130 ;
        RECT 33.555 15.005 33.640 15.165 ;
        RECT 0.740 14.385 0.815 14.525 ;
        RECT 0.955 14.335 1.030 14.475 ;
        RECT 1.660 14.395 1.720 14.475 ;
        POLYGON 1.660 14.395 1.720 14.395 1.720 14.335 ;
        RECT 1.875 14.385 1.950 14.525 ;
        RECT 3.640 14.385 3.715 14.525 ;
        RECT 3.855 14.335 3.930 14.475 ;
        RECT 4.560 14.395 4.620 14.475 ;
        POLYGON 4.560 14.395 4.620 14.395 4.620 14.335 ;
        RECT 4.775 14.385 4.850 14.525 ;
        RECT 6.540 14.385 6.615 14.525 ;
        RECT 6.755 14.335 6.830 14.475 ;
        RECT 7.460 14.395 7.520 14.475 ;
        POLYGON 7.460 14.395 7.520 14.395 7.520 14.335 ;
        RECT 7.675 14.385 7.750 14.525 ;
        RECT 9.440 14.385 9.515 14.525 ;
        RECT 9.655 14.335 9.730 14.475 ;
        RECT 10.360 14.395 10.420 14.475 ;
        POLYGON 10.360 14.395 10.420 14.395 10.420 14.335 ;
        RECT 10.575 14.385 10.650 14.525 ;
        RECT 12.340 14.385 12.415 14.525 ;
        RECT 12.555 14.335 12.630 14.475 ;
        RECT 13.260 14.395 13.320 14.475 ;
        POLYGON 13.260 14.395 13.320 14.395 13.320 14.335 ;
        RECT 13.475 14.385 13.550 14.525 ;
        RECT 15.240 14.385 15.315 14.525 ;
        RECT 15.455 14.335 15.530 14.475 ;
        RECT 16.160 14.395 16.220 14.475 ;
        POLYGON 16.160 14.395 16.220 14.395 16.220 14.335 ;
        RECT 16.375 14.385 16.450 14.525 ;
        RECT 18.140 14.385 18.215 14.525 ;
        RECT 18.355 14.335 18.430 14.475 ;
        RECT 19.060 14.395 19.120 14.475 ;
        POLYGON 19.060 14.395 19.120 14.395 19.120 14.335 ;
        RECT 19.275 14.385 19.350 14.525 ;
        RECT 21.040 14.385 21.115 14.525 ;
        RECT 21.255 14.335 21.330 14.475 ;
        RECT 21.960 14.395 22.020 14.475 ;
        POLYGON 21.960 14.395 22.020 14.395 22.020 14.335 ;
        RECT 22.175 14.385 22.250 14.525 ;
        RECT 23.940 14.385 24.015 14.525 ;
        RECT 24.155 14.335 24.230 14.475 ;
        RECT 24.860 14.395 24.920 14.475 ;
        POLYGON 24.860 14.395 24.920 14.395 24.920 14.335 ;
        RECT 25.075 14.385 25.150 14.525 ;
        RECT 26.840 14.385 26.915 14.525 ;
        RECT 27.055 14.335 27.130 14.475 ;
        RECT 27.760 14.395 27.820 14.475 ;
        POLYGON 27.760 14.395 27.820 14.395 27.820 14.335 ;
        RECT 27.975 14.385 28.050 14.525 ;
        RECT 29.740 14.385 29.815 14.525 ;
        RECT 29.955 14.335 30.030 14.475 ;
        RECT 30.660 14.395 30.720 14.475 ;
        POLYGON 30.660 14.395 30.720 14.395 30.720 14.335 ;
        RECT 30.875 14.385 30.950 14.525 ;
        RECT 32.640 14.385 32.715 14.525 ;
        RECT 32.855 14.335 32.930 14.475 ;
        RECT 33.560 14.395 33.620 14.475 ;
        POLYGON 33.560 14.395 33.620 14.395 33.620 14.335 ;
        RECT 33.775 14.385 33.850 14.525 ;
        RECT 0.685 13.865 0.835 14.035 ;
        RECT 1.075 14.000 1.225 14.170 ;
        RECT 1.465 14.000 1.615 14.170 ;
        RECT 1.855 13.865 2.005 14.035 ;
        RECT 3.585 13.865 3.735 14.035 ;
        RECT 3.975 14.000 4.125 14.170 ;
        RECT 4.365 14.000 4.515 14.170 ;
        RECT 4.755 13.865 4.905 14.035 ;
        RECT 6.485 13.865 6.635 14.035 ;
        RECT 6.875 14.000 7.025 14.170 ;
        RECT 7.265 14.000 7.415 14.170 ;
        RECT 7.655 13.865 7.805 14.035 ;
        RECT 9.385 13.865 9.535 14.035 ;
        RECT 9.775 14.000 9.925 14.170 ;
        RECT 10.165 14.000 10.315 14.170 ;
        RECT 10.555 13.865 10.705 14.035 ;
        RECT 12.285 13.865 12.435 14.035 ;
        RECT 12.675 14.000 12.825 14.170 ;
        RECT 13.065 14.000 13.215 14.170 ;
        RECT 13.455 13.865 13.605 14.035 ;
        RECT 15.185 13.865 15.335 14.035 ;
        RECT 15.575 14.000 15.725 14.170 ;
        RECT 15.965 14.000 16.115 14.170 ;
        RECT 16.355 13.865 16.505 14.035 ;
        RECT 18.085 13.865 18.235 14.035 ;
        RECT 18.475 14.000 18.625 14.170 ;
        RECT 18.865 14.000 19.015 14.170 ;
        RECT 19.255 13.865 19.405 14.035 ;
        RECT 20.985 13.865 21.135 14.035 ;
        RECT 21.375 14.000 21.525 14.170 ;
        RECT 21.765 14.000 21.915 14.170 ;
        RECT 22.155 13.865 22.305 14.035 ;
        RECT 23.885 13.865 24.035 14.035 ;
        RECT 24.275 14.000 24.425 14.170 ;
        RECT 24.665 14.000 24.815 14.170 ;
        RECT 25.055 13.865 25.205 14.035 ;
        RECT 26.785 13.865 26.935 14.035 ;
        RECT 27.175 14.000 27.325 14.170 ;
        RECT 27.565 14.000 27.715 14.170 ;
        RECT 27.955 13.865 28.105 14.035 ;
        RECT 29.685 13.865 29.835 14.035 ;
        RECT 30.075 14.000 30.225 14.170 ;
        RECT 30.465 14.000 30.615 14.170 ;
        RECT 30.855 13.865 31.005 14.035 ;
        RECT 32.585 13.865 32.735 14.035 ;
        RECT 32.975 14.000 33.125 14.170 ;
        RECT 33.365 14.000 33.515 14.170 ;
        RECT 33.755 13.865 33.905 14.035 ;
        RECT 0.950 13.780 1.000 13.815 ;
        POLYGON 1.000 13.815 1.035 13.780 1.000 13.780 ;
        RECT 0.950 13.655 1.035 13.780 ;
        RECT 1.655 13.655 1.740 13.815 ;
        RECT 3.850 13.780 3.900 13.815 ;
        POLYGON 3.900 13.815 3.935 13.780 3.900 13.780 ;
        RECT 3.850 13.655 3.935 13.780 ;
        RECT 4.555 13.655 4.640 13.815 ;
        RECT 6.750 13.780 6.800 13.815 ;
        POLYGON 6.800 13.815 6.835 13.780 6.800 13.780 ;
        RECT 6.750 13.655 6.835 13.780 ;
        RECT 7.455 13.655 7.540 13.815 ;
        RECT 9.650 13.780 9.700 13.815 ;
        POLYGON 9.700 13.815 9.735 13.780 9.700 13.780 ;
        RECT 9.650 13.655 9.735 13.780 ;
        RECT 10.355 13.655 10.440 13.815 ;
        RECT 12.550 13.780 12.600 13.815 ;
        POLYGON 12.600 13.815 12.635 13.780 12.600 13.780 ;
        RECT 12.550 13.655 12.635 13.780 ;
        RECT 13.255 13.655 13.340 13.815 ;
        RECT 15.450 13.780 15.500 13.815 ;
        POLYGON 15.500 13.815 15.535 13.780 15.500 13.780 ;
        RECT 15.450 13.655 15.535 13.780 ;
        RECT 16.155 13.655 16.240 13.815 ;
        RECT 18.350 13.780 18.400 13.815 ;
        POLYGON 18.400 13.815 18.435 13.780 18.400 13.780 ;
        RECT 18.350 13.655 18.435 13.780 ;
        RECT 19.055 13.655 19.140 13.815 ;
        RECT 21.250 13.780 21.300 13.815 ;
        POLYGON 21.300 13.815 21.335 13.780 21.300 13.780 ;
        RECT 21.250 13.655 21.335 13.780 ;
        RECT 21.955 13.655 22.040 13.815 ;
        RECT 24.150 13.780 24.200 13.815 ;
        POLYGON 24.200 13.815 24.235 13.780 24.200 13.780 ;
        RECT 24.150 13.655 24.235 13.780 ;
        RECT 24.855 13.655 24.940 13.815 ;
        RECT 27.050 13.780 27.100 13.815 ;
        POLYGON 27.100 13.815 27.135 13.780 27.100 13.780 ;
        RECT 27.050 13.655 27.135 13.780 ;
        RECT 27.755 13.655 27.840 13.815 ;
        RECT 29.950 13.780 30.000 13.815 ;
        POLYGON 30.000 13.815 30.035 13.780 30.000 13.780 ;
        RECT 29.950 13.655 30.035 13.780 ;
        RECT 30.655 13.655 30.740 13.815 ;
        RECT 32.850 13.780 32.900 13.815 ;
        POLYGON 32.900 13.815 32.935 13.780 32.900 13.780 ;
        RECT 32.850 13.655 32.935 13.780 ;
        RECT 33.555 13.655 33.640 13.815 ;
        RECT 0.740 13.035 0.815 13.175 ;
        RECT 0.955 12.985 1.030 13.125 ;
        RECT 1.660 13.045 1.720 13.125 ;
        POLYGON 1.660 13.045 1.720 13.045 1.720 12.985 ;
        RECT 1.875 13.035 1.950 13.175 ;
        RECT 3.640 13.035 3.715 13.175 ;
        RECT 3.855 12.985 3.930 13.125 ;
        RECT 4.560 13.045 4.620 13.125 ;
        POLYGON 4.560 13.045 4.620 13.045 4.620 12.985 ;
        RECT 4.775 13.035 4.850 13.175 ;
        RECT 6.540 13.035 6.615 13.175 ;
        RECT 6.755 12.985 6.830 13.125 ;
        RECT 7.460 13.045 7.520 13.125 ;
        POLYGON 7.460 13.045 7.520 13.045 7.520 12.985 ;
        RECT 7.675 13.035 7.750 13.175 ;
        RECT 9.440 13.035 9.515 13.175 ;
        RECT 9.655 12.985 9.730 13.125 ;
        RECT 10.360 13.045 10.420 13.125 ;
        POLYGON 10.360 13.045 10.420 13.045 10.420 12.985 ;
        RECT 10.575 13.035 10.650 13.175 ;
        RECT 12.340 13.035 12.415 13.175 ;
        RECT 12.555 12.985 12.630 13.125 ;
        RECT 13.260 13.045 13.320 13.125 ;
        POLYGON 13.260 13.045 13.320 13.045 13.320 12.985 ;
        RECT 13.475 13.035 13.550 13.175 ;
        RECT 15.240 13.035 15.315 13.175 ;
        RECT 15.455 12.985 15.530 13.125 ;
        RECT 16.160 13.045 16.220 13.125 ;
        POLYGON 16.160 13.045 16.220 13.045 16.220 12.985 ;
        RECT 16.375 13.035 16.450 13.175 ;
        RECT 18.140 13.035 18.215 13.175 ;
        RECT 18.355 12.985 18.430 13.125 ;
        RECT 19.060 13.045 19.120 13.125 ;
        POLYGON 19.060 13.045 19.120 13.045 19.120 12.985 ;
        RECT 19.275 13.035 19.350 13.175 ;
        RECT 21.040 13.035 21.115 13.175 ;
        RECT 21.255 12.985 21.330 13.125 ;
        RECT 21.960 13.045 22.020 13.125 ;
        POLYGON 21.960 13.045 22.020 13.045 22.020 12.985 ;
        RECT 22.175 13.035 22.250 13.175 ;
        RECT 23.940 13.035 24.015 13.175 ;
        RECT 24.155 12.985 24.230 13.125 ;
        RECT 24.860 13.045 24.920 13.125 ;
        POLYGON 24.860 13.045 24.920 13.045 24.920 12.985 ;
        RECT 25.075 13.035 25.150 13.175 ;
        RECT 26.840 13.035 26.915 13.175 ;
        RECT 27.055 12.985 27.130 13.125 ;
        RECT 27.760 13.045 27.820 13.125 ;
        POLYGON 27.760 13.045 27.820 13.045 27.820 12.985 ;
        RECT 27.975 13.035 28.050 13.175 ;
        RECT 29.740 13.035 29.815 13.175 ;
        RECT 29.955 12.985 30.030 13.125 ;
        RECT 30.660 13.045 30.720 13.125 ;
        POLYGON 30.660 13.045 30.720 13.045 30.720 12.985 ;
        RECT 30.875 13.035 30.950 13.175 ;
        RECT 32.640 13.035 32.715 13.175 ;
        RECT 32.855 12.985 32.930 13.125 ;
        RECT 33.560 13.045 33.620 13.125 ;
        POLYGON 33.560 13.045 33.620 13.045 33.620 12.985 ;
        RECT 33.775 13.035 33.850 13.175 ;
        RECT 0.685 12.515 0.835 12.685 ;
        RECT 1.075 12.650 1.225 12.820 ;
        RECT 1.465 12.650 1.615 12.820 ;
        RECT 1.855 12.515 2.005 12.685 ;
        RECT 3.585 12.515 3.735 12.685 ;
        RECT 3.975 12.650 4.125 12.820 ;
        RECT 4.365 12.650 4.515 12.820 ;
        RECT 4.755 12.515 4.905 12.685 ;
        RECT 6.485 12.515 6.635 12.685 ;
        RECT 6.875 12.650 7.025 12.820 ;
        RECT 7.265 12.650 7.415 12.820 ;
        RECT 7.655 12.515 7.805 12.685 ;
        RECT 9.385 12.515 9.535 12.685 ;
        RECT 9.775 12.650 9.925 12.820 ;
        RECT 10.165 12.650 10.315 12.820 ;
        RECT 10.555 12.515 10.705 12.685 ;
        RECT 12.285 12.515 12.435 12.685 ;
        RECT 12.675 12.650 12.825 12.820 ;
        RECT 13.065 12.650 13.215 12.820 ;
        RECT 13.455 12.515 13.605 12.685 ;
        RECT 15.185 12.515 15.335 12.685 ;
        RECT 15.575 12.650 15.725 12.820 ;
        RECT 15.965 12.650 16.115 12.820 ;
        RECT 16.355 12.515 16.505 12.685 ;
        RECT 18.085 12.515 18.235 12.685 ;
        RECT 18.475 12.650 18.625 12.820 ;
        RECT 18.865 12.650 19.015 12.820 ;
        RECT 19.255 12.515 19.405 12.685 ;
        RECT 20.985 12.515 21.135 12.685 ;
        RECT 21.375 12.650 21.525 12.820 ;
        RECT 21.765 12.650 21.915 12.820 ;
        RECT 22.155 12.515 22.305 12.685 ;
        RECT 23.885 12.515 24.035 12.685 ;
        RECT 24.275 12.650 24.425 12.820 ;
        RECT 24.665 12.650 24.815 12.820 ;
        RECT 25.055 12.515 25.205 12.685 ;
        RECT 26.785 12.515 26.935 12.685 ;
        RECT 27.175 12.650 27.325 12.820 ;
        RECT 27.565 12.650 27.715 12.820 ;
        RECT 27.955 12.515 28.105 12.685 ;
        RECT 29.685 12.515 29.835 12.685 ;
        RECT 30.075 12.650 30.225 12.820 ;
        RECT 30.465 12.650 30.615 12.820 ;
        RECT 30.855 12.515 31.005 12.685 ;
        RECT 32.585 12.515 32.735 12.685 ;
        RECT 32.975 12.650 33.125 12.820 ;
        RECT 33.365 12.650 33.515 12.820 ;
        RECT 33.755 12.515 33.905 12.685 ;
        RECT 0.950 12.430 1.000 12.465 ;
        POLYGON 1.000 12.465 1.035 12.430 1.000 12.430 ;
        RECT 0.950 12.305 1.035 12.430 ;
        RECT 1.655 12.305 1.740 12.465 ;
        RECT 3.850 12.430 3.900 12.465 ;
        POLYGON 3.900 12.465 3.935 12.430 3.900 12.430 ;
        RECT 3.850 12.305 3.935 12.430 ;
        RECT 4.555 12.305 4.640 12.465 ;
        RECT 6.750 12.430 6.800 12.465 ;
        POLYGON 6.800 12.465 6.835 12.430 6.800 12.430 ;
        RECT 6.750 12.305 6.835 12.430 ;
        RECT 7.455 12.305 7.540 12.465 ;
        RECT 9.650 12.430 9.700 12.465 ;
        POLYGON 9.700 12.465 9.735 12.430 9.700 12.430 ;
        RECT 9.650 12.305 9.735 12.430 ;
        RECT 10.355 12.305 10.440 12.465 ;
        RECT 12.550 12.430 12.600 12.465 ;
        POLYGON 12.600 12.465 12.635 12.430 12.600 12.430 ;
        RECT 12.550 12.305 12.635 12.430 ;
        RECT 13.255 12.305 13.340 12.465 ;
        RECT 15.450 12.430 15.500 12.465 ;
        POLYGON 15.500 12.465 15.535 12.430 15.500 12.430 ;
        RECT 15.450 12.305 15.535 12.430 ;
        RECT 16.155 12.305 16.240 12.465 ;
        RECT 18.350 12.430 18.400 12.465 ;
        POLYGON 18.400 12.465 18.435 12.430 18.400 12.430 ;
        RECT 18.350 12.305 18.435 12.430 ;
        RECT 19.055 12.305 19.140 12.465 ;
        RECT 21.250 12.430 21.300 12.465 ;
        POLYGON 21.300 12.465 21.335 12.430 21.300 12.430 ;
        RECT 21.250 12.305 21.335 12.430 ;
        RECT 21.955 12.305 22.040 12.465 ;
        RECT 24.150 12.430 24.200 12.465 ;
        POLYGON 24.200 12.465 24.235 12.430 24.200 12.430 ;
        RECT 24.150 12.305 24.235 12.430 ;
        RECT 24.855 12.305 24.940 12.465 ;
        RECT 27.050 12.430 27.100 12.465 ;
        POLYGON 27.100 12.465 27.135 12.430 27.100 12.430 ;
        RECT 27.050 12.305 27.135 12.430 ;
        RECT 27.755 12.305 27.840 12.465 ;
        RECT 29.950 12.430 30.000 12.465 ;
        POLYGON 30.000 12.465 30.035 12.430 30.000 12.430 ;
        RECT 29.950 12.305 30.035 12.430 ;
        RECT 30.655 12.305 30.740 12.465 ;
        RECT 32.850 12.430 32.900 12.465 ;
        POLYGON 32.900 12.465 32.935 12.430 32.900 12.430 ;
        RECT 32.850 12.305 32.935 12.430 ;
        RECT 33.555 12.305 33.640 12.465 ;
        RECT 0.740 11.685 0.815 11.825 ;
        RECT 0.955 11.635 1.030 11.775 ;
        RECT 1.660 11.695 1.720 11.775 ;
        POLYGON 1.660 11.695 1.720 11.695 1.720 11.635 ;
        RECT 1.875 11.685 1.950 11.825 ;
        RECT 3.640 11.685 3.715 11.825 ;
        RECT 3.855 11.635 3.930 11.775 ;
        RECT 4.560 11.695 4.620 11.775 ;
        POLYGON 4.560 11.695 4.620 11.695 4.620 11.635 ;
        RECT 4.775 11.685 4.850 11.825 ;
        RECT 6.540 11.685 6.615 11.825 ;
        RECT 6.755 11.635 6.830 11.775 ;
        RECT 7.460 11.695 7.520 11.775 ;
        POLYGON 7.460 11.695 7.520 11.695 7.520 11.635 ;
        RECT 7.675 11.685 7.750 11.825 ;
        RECT 9.440 11.685 9.515 11.825 ;
        RECT 9.655 11.635 9.730 11.775 ;
        RECT 10.360 11.695 10.420 11.775 ;
        POLYGON 10.360 11.695 10.420 11.695 10.420 11.635 ;
        RECT 10.575 11.685 10.650 11.825 ;
        RECT 12.340 11.685 12.415 11.825 ;
        RECT 12.555 11.635 12.630 11.775 ;
        RECT 13.260 11.695 13.320 11.775 ;
        POLYGON 13.260 11.695 13.320 11.695 13.320 11.635 ;
        RECT 13.475 11.685 13.550 11.825 ;
        RECT 15.240 11.685 15.315 11.825 ;
        RECT 15.455 11.635 15.530 11.775 ;
        RECT 16.160 11.695 16.220 11.775 ;
        POLYGON 16.160 11.695 16.220 11.695 16.220 11.635 ;
        RECT 16.375 11.685 16.450 11.825 ;
        RECT 18.140 11.685 18.215 11.825 ;
        RECT 18.355 11.635 18.430 11.775 ;
        RECT 19.060 11.695 19.120 11.775 ;
        POLYGON 19.060 11.695 19.120 11.695 19.120 11.635 ;
        RECT 19.275 11.685 19.350 11.825 ;
        RECT 21.040 11.685 21.115 11.825 ;
        RECT 21.255 11.635 21.330 11.775 ;
        RECT 21.960 11.695 22.020 11.775 ;
        POLYGON 21.960 11.695 22.020 11.695 22.020 11.635 ;
        RECT 22.175 11.685 22.250 11.825 ;
        RECT 23.940 11.685 24.015 11.825 ;
        RECT 24.155 11.635 24.230 11.775 ;
        RECT 24.860 11.695 24.920 11.775 ;
        POLYGON 24.860 11.695 24.920 11.695 24.920 11.635 ;
        RECT 25.075 11.685 25.150 11.825 ;
        RECT 26.840 11.685 26.915 11.825 ;
        RECT 27.055 11.635 27.130 11.775 ;
        RECT 27.760 11.695 27.820 11.775 ;
        POLYGON 27.760 11.695 27.820 11.695 27.820 11.635 ;
        RECT 27.975 11.685 28.050 11.825 ;
        RECT 29.740 11.685 29.815 11.825 ;
        RECT 29.955 11.635 30.030 11.775 ;
        RECT 30.660 11.695 30.720 11.775 ;
        POLYGON 30.660 11.695 30.720 11.695 30.720 11.635 ;
        RECT 30.875 11.685 30.950 11.825 ;
        RECT 32.640 11.685 32.715 11.825 ;
        RECT 32.855 11.635 32.930 11.775 ;
        RECT 33.560 11.695 33.620 11.775 ;
        POLYGON 33.560 11.695 33.620 11.695 33.620 11.635 ;
        RECT 33.775 11.685 33.850 11.825 ;
        RECT 0.685 11.165 0.835 11.335 ;
        RECT 1.075 11.300 1.225 11.470 ;
        RECT 1.465 11.300 1.615 11.470 ;
        RECT 1.855 11.165 2.005 11.335 ;
        RECT 3.585 11.165 3.735 11.335 ;
        RECT 3.975 11.300 4.125 11.470 ;
        RECT 4.365 11.300 4.515 11.470 ;
        RECT 4.755 11.165 4.905 11.335 ;
        RECT 6.485 11.165 6.635 11.335 ;
        RECT 6.875 11.300 7.025 11.470 ;
        RECT 7.265 11.300 7.415 11.470 ;
        RECT 7.655 11.165 7.805 11.335 ;
        RECT 9.385 11.165 9.535 11.335 ;
        RECT 9.775 11.300 9.925 11.470 ;
        RECT 10.165 11.300 10.315 11.470 ;
        RECT 10.555 11.165 10.705 11.335 ;
        RECT 12.285 11.165 12.435 11.335 ;
        RECT 12.675 11.300 12.825 11.470 ;
        RECT 13.065 11.300 13.215 11.470 ;
        RECT 13.455 11.165 13.605 11.335 ;
        RECT 15.185 11.165 15.335 11.335 ;
        RECT 15.575 11.300 15.725 11.470 ;
        RECT 15.965 11.300 16.115 11.470 ;
        RECT 16.355 11.165 16.505 11.335 ;
        RECT 18.085 11.165 18.235 11.335 ;
        RECT 18.475 11.300 18.625 11.470 ;
        RECT 18.865 11.300 19.015 11.470 ;
        RECT 19.255 11.165 19.405 11.335 ;
        RECT 20.985 11.165 21.135 11.335 ;
        RECT 21.375 11.300 21.525 11.470 ;
        RECT 21.765 11.300 21.915 11.470 ;
        RECT 22.155 11.165 22.305 11.335 ;
        RECT 23.885 11.165 24.035 11.335 ;
        RECT 24.275 11.300 24.425 11.470 ;
        RECT 24.665 11.300 24.815 11.470 ;
        RECT 25.055 11.165 25.205 11.335 ;
        RECT 26.785 11.165 26.935 11.335 ;
        RECT 27.175 11.300 27.325 11.470 ;
        RECT 27.565 11.300 27.715 11.470 ;
        RECT 27.955 11.165 28.105 11.335 ;
        RECT 29.685 11.165 29.835 11.335 ;
        RECT 30.075 11.300 30.225 11.470 ;
        RECT 30.465 11.300 30.615 11.470 ;
        RECT 30.855 11.165 31.005 11.335 ;
        RECT 32.585 11.165 32.735 11.335 ;
        RECT 32.975 11.300 33.125 11.470 ;
        RECT 33.365 11.300 33.515 11.470 ;
        RECT 33.755 11.165 33.905 11.335 ;
        RECT 0.950 11.080 1.000 11.115 ;
        POLYGON 1.000 11.115 1.035 11.080 1.000 11.080 ;
        RECT 0.950 10.955 1.035 11.080 ;
        RECT 1.655 10.955 1.740 11.115 ;
        RECT 3.850 11.080 3.900 11.115 ;
        POLYGON 3.900 11.115 3.935 11.080 3.900 11.080 ;
        RECT 3.850 10.955 3.935 11.080 ;
        RECT 4.555 10.955 4.640 11.115 ;
        RECT 6.750 11.080 6.800 11.115 ;
        POLYGON 6.800 11.115 6.835 11.080 6.800 11.080 ;
        RECT 6.750 10.955 6.835 11.080 ;
        RECT 7.455 10.955 7.540 11.115 ;
        RECT 9.650 11.080 9.700 11.115 ;
        POLYGON 9.700 11.115 9.735 11.080 9.700 11.080 ;
        RECT 9.650 10.955 9.735 11.080 ;
        RECT 10.355 10.955 10.440 11.115 ;
        RECT 12.550 11.080 12.600 11.115 ;
        POLYGON 12.600 11.115 12.635 11.080 12.600 11.080 ;
        RECT 12.550 10.955 12.635 11.080 ;
        RECT 13.255 10.955 13.340 11.115 ;
        RECT 15.450 11.080 15.500 11.115 ;
        POLYGON 15.500 11.115 15.535 11.080 15.500 11.080 ;
        RECT 15.450 10.955 15.535 11.080 ;
        RECT 16.155 10.955 16.240 11.115 ;
        RECT 18.350 11.080 18.400 11.115 ;
        POLYGON 18.400 11.115 18.435 11.080 18.400 11.080 ;
        RECT 18.350 10.955 18.435 11.080 ;
        RECT 19.055 10.955 19.140 11.115 ;
        RECT 21.250 11.080 21.300 11.115 ;
        POLYGON 21.300 11.115 21.335 11.080 21.300 11.080 ;
        RECT 21.250 10.955 21.335 11.080 ;
        RECT 21.955 10.955 22.040 11.115 ;
        RECT 24.150 11.080 24.200 11.115 ;
        POLYGON 24.200 11.115 24.235 11.080 24.200 11.080 ;
        RECT 24.150 10.955 24.235 11.080 ;
        RECT 24.855 10.955 24.940 11.115 ;
        RECT 27.050 11.080 27.100 11.115 ;
        POLYGON 27.100 11.115 27.135 11.080 27.100 11.080 ;
        RECT 27.050 10.955 27.135 11.080 ;
        RECT 27.755 10.955 27.840 11.115 ;
        RECT 29.950 11.080 30.000 11.115 ;
        POLYGON 30.000 11.115 30.035 11.080 30.000 11.080 ;
        RECT 29.950 10.955 30.035 11.080 ;
        RECT 30.655 10.955 30.740 11.115 ;
        RECT 32.850 11.080 32.900 11.115 ;
        POLYGON 32.900 11.115 32.935 11.080 32.900 11.080 ;
        RECT 32.850 10.955 32.935 11.080 ;
        RECT 33.555 10.955 33.640 11.115 ;
        RECT 0.740 10.335 0.815 10.475 ;
        RECT 0.955 10.285 1.030 10.425 ;
        RECT 1.660 10.345 1.720 10.425 ;
        POLYGON 1.660 10.345 1.720 10.345 1.720 10.285 ;
        RECT 1.875 10.335 1.950 10.475 ;
        RECT 3.640 10.335 3.715 10.475 ;
        RECT 3.855 10.285 3.930 10.425 ;
        RECT 4.560 10.345 4.620 10.425 ;
        POLYGON 4.560 10.345 4.620 10.345 4.620 10.285 ;
        RECT 4.775 10.335 4.850 10.475 ;
        RECT 6.540 10.335 6.615 10.475 ;
        RECT 6.755 10.285 6.830 10.425 ;
        RECT 7.460 10.345 7.520 10.425 ;
        POLYGON 7.460 10.345 7.520 10.345 7.520 10.285 ;
        RECT 7.675 10.335 7.750 10.475 ;
        RECT 9.440 10.335 9.515 10.475 ;
        RECT 9.655 10.285 9.730 10.425 ;
        RECT 10.360 10.345 10.420 10.425 ;
        POLYGON 10.360 10.345 10.420 10.345 10.420 10.285 ;
        RECT 10.575 10.335 10.650 10.475 ;
        RECT 12.340 10.335 12.415 10.475 ;
        RECT 12.555 10.285 12.630 10.425 ;
        RECT 13.260 10.345 13.320 10.425 ;
        POLYGON 13.260 10.345 13.320 10.345 13.320 10.285 ;
        RECT 13.475 10.335 13.550 10.475 ;
        RECT 15.240 10.335 15.315 10.475 ;
        RECT 15.455 10.285 15.530 10.425 ;
        RECT 16.160 10.345 16.220 10.425 ;
        POLYGON 16.160 10.345 16.220 10.345 16.220 10.285 ;
        RECT 16.375 10.335 16.450 10.475 ;
        RECT 18.140 10.335 18.215 10.475 ;
        RECT 18.355 10.285 18.430 10.425 ;
        RECT 19.060 10.345 19.120 10.425 ;
        POLYGON 19.060 10.345 19.120 10.345 19.120 10.285 ;
        RECT 19.275 10.335 19.350 10.475 ;
        RECT 21.040 10.335 21.115 10.475 ;
        RECT 21.255 10.285 21.330 10.425 ;
        RECT 21.960 10.345 22.020 10.425 ;
        POLYGON 21.960 10.345 22.020 10.345 22.020 10.285 ;
        RECT 22.175 10.335 22.250 10.475 ;
        RECT 23.940 10.335 24.015 10.475 ;
        RECT 24.155 10.285 24.230 10.425 ;
        RECT 24.860 10.345 24.920 10.425 ;
        POLYGON 24.860 10.345 24.920 10.345 24.920 10.285 ;
        RECT 25.075 10.335 25.150 10.475 ;
        RECT 26.840 10.335 26.915 10.475 ;
        RECT 27.055 10.285 27.130 10.425 ;
        RECT 27.760 10.345 27.820 10.425 ;
        POLYGON 27.760 10.345 27.820 10.345 27.820 10.285 ;
        RECT 27.975 10.335 28.050 10.475 ;
        RECT 29.740 10.335 29.815 10.475 ;
        RECT 29.955 10.285 30.030 10.425 ;
        RECT 30.660 10.345 30.720 10.425 ;
        POLYGON 30.660 10.345 30.720 10.345 30.720 10.285 ;
        RECT 30.875 10.335 30.950 10.475 ;
        RECT 32.640 10.335 32.715 10.475 ;
        RECT 32.855 10.285 32.930 10.425 ;
        RECT 33.560 10.345 33.620 10.425 ;
        POLYGON 33.560 10.345 33.620 10.345 33.620 10.285 ;
        RECT 33.775 10.335 33.850 10.475 ;
        RECT 0.685 9.815 0.835 9.985 ;
        RECT 1.075 9.950 1.225 10.120 ;
        RECT 1.465 9.950 1.615 10.120 ;
        RECT 1.855 9.815 2.005 9.985 ;
        RECT 3.585 9.815 3.735 9.985 ;
        RECT 3.975 9.950 4.125 10.120 ;
        RECT 4.365 9.950 4.515 10.120 ;
        RECT 4.755 9.815 4.905 9.985 ;
        RECT 6.485 9.815 6.635 9.985 ;
        RECT 6.875 9.950 7.025 10.120 ;
        RECT 7.265 9.950 7.415 10.120 ;
        RECT 7.655 9.815 7.805 9.985 ;
        RECT 9.385 9.815 9.535 9.985 ;
        RECT 9.775 9.950 9.925 10.120 ;
        RECT 10.165 9.950 10.315 10.120 ;
        RECT 10.555 9.815 10.705 9.985 ;
        RECT 12.285 9.815 12.435 9.985 ;
        RECT 12.675 9.950 12.825 10.120 ;
        RECT 13.065 9.950 13.215 10.120 ;
        RECT 13.455 9.815 13.605 9.985 ;
        RECT 15.185 9.815 15.335 9.985 ;
        RECT 15.575 9.950 15.725 10.120 ;
        RECT 15.965 9.950 16.115 10.120 ;
        RECT 16.355 9.815 16.505 9.985 ;
        RECT 18.085 9.815 18.235 9.985 ;
        RECT 18.475 9.950 18.625 10.120 ;
        RECT 18.865 9.950 19.015 10.120 ;
        RECT 19.255 9.815 19.405 9.985 ;
        RECT 20.985 9.815 21.135 9.985 ;
        RECT 21.375 9.950 21.525 10.120 ;
        RECT 21.765 9.950 21.915 10.120 ;
        RECT 22.155 9.815 22.305 9.985 ;
        RECT 23.885 9.815 24.035 9.985 ;
        RECT 24.275 9.950 24.425 10.120 ;
        RECT 24.665 9.950 24.815 10.120 ;
        RECT 25.055 9.815 25.205 9.985 ;
        RECT 26.785 9.815 26.935 9.985 ;
        RECT 27.175 9.950 27.325 10.120 ;
        RECT 27.565 9.950 27.715 10.120 ;
        RECT 27.955 9.815 28.105 9.985 ;
        RECT 29.685 9.815 29.835 9.985 ;
        RECT 30.075 9.950 30.225 10.120 ;
        RECT 30.465 9.950 30.615 10.120 ;
        RECT 30.855 9.815 31.005 9.985 ;
        RECT 32.585 9.815 32.735 9.985 ;
        RECT 32.975 9.950 33.125 10.120 ;
        RECT 33.365 9.950 33.515 10.120 ;
        RECT 33.755 9.815 33.905 9.985 ;
        RECT 0.950 9.730 1.000 9.765 ;
        POLYGON 1.000 9.765 1.035 9.730 1.000 9.730 ;
        RECT 0.950 9.605 1.035 9.730 ;
        RECT 1.655 9.605 1.740 9.765 ;
        RECT 3.850 9.730 3.900 9.765 ;
        POLYGON 3.900 9.765 3.935 9.730 3.900 9.730 ;
        RECT 3.850 9.605 3.935 9.730 ;
        RECT 4.555 9.605 4.640 9.765 ;
        RECT 6.750 9.730 6.800 9.765 ;
        POLYGON 6.800 9.765 6.835 9.730 6.800 9.730 ;
        RECT 6.750 9.605 6.835 9.730 ;
        RECT 7.455 9.605 7.540 9.765 ;
        RECT 9.650 9.730 9.700 9.765 ;
        POLYGON 9.700 9.765 9.735 9.730 9.700 9.730 ;
        RECT 9.650 9.605 9.735 9.730 ;
        RECT 10.355 9.605 10.440 9.765 ;
        RECT 12.550 9.730 12.600 9.765 ;
        POLYGON 12.600 9.765 12.635 9.730 12.600 9.730 ;
        RECT 12.550 9.605 12.635 9.730 ;
        RECT 13.255 9.605 13.340 9.765 ;
        RECT 15.450 9.730 15.500 9.765 ;
        POLYGON 15.500 9.765 15.535 9.730 15.500 9.730 ;
        RECT 15.450 9.605 15.535 9.730 ;
        RECT 16.155 9.605 16.240 9.765 ;
        RECT 18.350 9.730 18.400 9.765 ;
        POLYGON 18.400 9.765 18.435 9.730 18.400 9.730 ;
        RECT 18.350 9.605 18.435 9.730 ;
        RECT 19.055 9.605 19.140 9.765 ;
        RECT 21.250 9.730 21.300 9.765 ;
        POLYGON 21.300 9.765 21.335 9.730 21.300 9.730 ;
        RECT 21.250 9.605 21.335 9.730 ;
        RECT 21.955 9.605 22.040 9.765 ;
        RECT 24.150 9.730 24.200 9.765 ;
        POLYGON 24.200 9.765 24.235 9.730 24.200 9.730 ;
        RECT 24.150 9.605 24.235 9.730 ;
        RECT 24.855 9.605 24.940 9.765 ;
        RECT 27.050 9.730 27.100 9.765 ;
        POLYGON 27.100 9.765 27.135 9.730 27.100 9.730 ;
        RECT 27.050 9.605 27.135 9.730 ;
        RECT 27.755 9.605 27.840 9.765 ;
        RECT 29.950 9.730 30.000 9.765 ;
        POLYGON 30.000 9.765 30.035 9.730 30.000 9.730 ;
        RECT 29.950 9.605 30.035 9.730 ;
        RECT 30.655 9.605 30.740 9.765 ;
        RECT 32.850 9.730 32.900 9.765 ;
        POLYGON 32.900 9.765 32.935 9.730 32.900 9.730 ;
        RECT 32.850 9.605 32.935 9.730 ;
        RECT 33.555 9.605 33.640 9.765 ;
        RECT 0.740 8.985 0.815 9.125 ;
        RECT 0.955 8.935 1.030 9.075 ;
        RECT 1.660 8.995 1.720 9.075 ;
        POLYGON 1.660 8.995 1.720 8.995 1.720 8.935 ;
        RECT 1.875 8.985 1.950 9.125 ;
        RECT 3.640 8.985 3.715 9.125 ;
        RECT 3.855 8.935 3.930 9.075 ;
        RECT 4.560 8.995 4.620 9.075 ;
        POLYGON 4.560 8.995 4.620 8.995 4.620 8.935 ;
        RECT 4.775 8.985 4.850 9.125 ;
        RECT 6.540 8.985 6.615 9.125 ;
        RECT 6.755 8.935 6.830 9.075 ;
        RECT 7.460 8.995 7.520 9.075 ;
        POLYGON 7.460 8.995 7.520 8.995 7.520 8.935 ;
        RECT 7.675 8.985 7.750 9.125 ;
        RECT 9.440 8.985 9.515 9.125 ;
        RECT 9.655 8.935 9.730 9.075 ;
        RECT 10.360 8.995 10.420 9.075 ;
        POLYGON 10.360 8.995 10.420 8.995 10.420 8.935 ;
        RECT 10.575 8.985 10.650 9.125 ;
        RECT 12.340 8.985 12.415 9.125 ;
        RECT 12.555 8.935 12.630 9.075 ;
        RECT 13.260 8.995 13.320 9.075 ;
        POLYGON 13.260 8.995 13.320 8.995 13.320 8.935 ;
        RECT 13.475 8.985 13.550 9.125 ;
        RECT 15.240 8.985 15.315 9.125 ;
        RECT 15.455 8.935 15.530 9.075 ;
        RECT 16.160 8.995 16.220 9.075 ;
        POLYGON 16.160 8.995 16.220 8.995 16.220 8.935 ;
        RECT 16.375 8.985 16.450 9.125 ;
        RECT 18.140 8.985 18.215 9.125 ;
        RECT 18.355 8.935 18.430 9.075 ;
        RECT 19.060 8.995 19.120 9.075 ;
        POLYGON 19.060 8.995 19.120 8.995 19.120 8.935 ;
        RECT 19.275 8.985 19.350 9.125 ;
        RECT 21.040 8.985 21.115 9.125 ;
        RECT 21.255 8.935 21.330 9.075 ;
        RECT 21.960 8.995 22.020 9.075 ;
        POLYGON 21.960 8.995 22.020 8.995 22.020 8.935 ;
        RECT 22.175 8.985 22.250 9.125 ;
        RECT 23.940 8.985 24.015 9.125 ;
        RECT 24.155 8.935 24.230 9.075 ;
        RECT 24.860 8.995 24.920 9.075 ;
        POLYGON 24.860 8.995 24.920 8.995 24.920 8.935 ;
        RECT 25.075 8.985 25.150 9.125 ;
        RECT 26.840 8.985 26.915 9.125 ;
        RECT 27.055 8.935 27.130 9.075 ;
        RECT 27.760 8.995 27.820 9.075 ;
        POLYGON 27.760 8.995 27.820 8.995 27.820 8.935 ;
        RECT 27.975 8.985 28.050 9.125 ;
        RECT 29.740 8.985 29.815 9.125 ;
        RECT 29.955 8.935 30.030 9.075 ;
        RECT 30.660 8.995 30.720 9.075 ;
        POLYGON 30.660 8.995 30.720 8.995 30.720 8.935 ;
        RECT 30.875 8.985 30.950 9.125 ;
        RECT 32.640 8.985 32.715 9.125 ;
        RECT 32.855 8.935 32.930 9.075 ;
        RECT 33.560 8.995 33.620 9.075 ;
        POLYGON 33.560 8.995 33.620 8.995 33.620 8.935 ;
        RECT 33.775 8.985 33.850 9.125 ;
        RECT 0.685 8.465 0.835 8.635 ;
        RECT 1.075 8.600 1.225 8.770 ;
        RECT 1.465 8.600 1.615 8.770 ;
        RECT 1.855 8.465 2.005 8.635 ;
        RECT 3.585 8.465 3.735 8.635 ;
        RECT 3.975 8.600 4.125 8.770 ;
        RECT 4.365 8.600 4.515 8.770 ;
        RECT 4.755 8.465 4.905 8.635 ;
        RECT 6.485 8.465 6.635 8.635 ;
        RECT 6.875 8.600 7.025 8.770 ;
        RECT 7.265 8.600 7.415 8.770 ;
        RECT 7.655 8.465 7.805 8.635 ;
        RECT 9.385 8.465 9.535 8.635 ;
        RECT 9.775 8.600 9.925 8.770 ;
        RECT 10.165 8.600 10.315 8.770 ;
        RECT 10.555 8.465 10.705 8.635 ;
        RECT 12.285 8.465 12.435 8.635 ;
        RECT 12.675 8.600 12.825 8.770 ;
        RECT 13.065 8.600 13.215 8.770 ;
        RECT 13.455 8.465 13.605 8.635 ;
        RECT 15.185 8.465 15.335 8.635 ;
        RECT 15.575 8.600 15.725 8.770 ;
        RECT 15.965 8.600 16.115 8.770 ;
        RECT 16.355 8.465 16.505 8.635 ;
        RECT 18.085 8.465 18.235 8.635 ;
        RECT 18.475 8.600 18.625 8.770 ;
        RECT 18.865 8.600 19.015 8.770 ;
        RECT 19.255 8.465 19.405 8.635 ;
        RECT 20.985 8.465 21.135 8.635 ;
        RECT 21.375 8.600 21.525 8.770 ;
        RECT 21.765 8.600 21.915 8.770 ;
        RECT 22.155 8.465 22.305 8.635 ;
        RECT 23.885 8.465 24.035 8.635 ;
        RECT 24.275 8.600 24.425 8.770 ;
        RECT 24.665 8.600 24.815 8.770 ;
        RECT 25.055 8.465 25.205 8.635 ;
        RECT 26.785 8.465 26.935 8.635 ;
        RECT 27.175 8.600 27.325 8.770 ;
        RECT 27.565 8.600 27.715 8.770 ;
        RECT 27.955 8.465 28.105 8.635 ;
        RECT 29.685 8.465 29.835 8.635 ;
        RECT 30.075 8.600 30.225 8.770 ;
        RECT 30.465 8.600 30.615 8.770 ;
        RECT 30.855 8.465 31.005 8.635 ;
        RECT 32.585 8.465 32.735 8.635 ;
        RECT 32.975 8.600 33.125 8.770 ;
        RECT 33.365 8.600 33.515 8.770 ;
        RECT 33.755 8.465 33.905 8.635 ;
        RECT 0.950 8.380 1.000 8.415 ;
        POLYGON 1.000 8.415 1.035 8.380 1.000 8.380 ;
        RECT 0.950 8.255 1.035 8.380 ;
        RECT 1.655 8.255 1.740 8.415 ;
        RECT 3.850 8.380 3.900 8.415 ;
        POLYGON 3.900 8.415 3.935 8.380 3.900 8.380 ;
        RECT 3.850 8.255 3.935 8.380 ;
        RECT 4.555 8.255 4.640 8.415 ;
        RECT 6.750 8.380 6.800 8.415 ;
        POLYGON 6.800 8.415 6.835 8.380 6.800 8.380 ;
        RECT 6.750 8.255 6.835 8.380 ;
        RECT 7.455 8.255 7.540 8.415 ;
        RECT 9.650 8.380 9.700 8.415 ;
        POLYGON 9.700 8.415 9.735 8.380 9.700 8.380 ;
        RECT 9.650 8.255 9.735 8.380 ;
        RECT 10.355 8.255 10.440 8.415 ;
        RECT 12.550 8.380 12.600 8.415 ;
        POLYGON 12.600 8.415 12.635 8.380 12.600 8.380 ;
        RECT 12.550 8.255 12.635 8.380 ;
        RECT 13.255 8.255 13.340 8.415 ;
        RECT 15.450 8.380 15.500 8.415 ;
        POLYGON 15.500 8.415 15.535 8.380 15.500 8.380 ;
        RECT 15.450 8.255 15.535 8.380 ;
        RECT 16.155 8.255 16.240 8.415 ;
        RECT 18.350 8.380 18.400 8.415 ;
        POLYGON 18.400 8.415 18.435 8.380 18.400 8.380 ;
        RECT 18.350 8.255 18.435 8.380 ;
        RECT 19.055 8.255 19.140 8.415 ;
        RECT 21.250 8.380 21.300 8.415 ;
        POLYGON 21.300 8.415 21.335 8.380 21.300 8.380 ;
        RECT 21.250 8.255 21.335 8.380 ;
        RECT 21.955 8.255 22.040 8.415 ;
        RECT 24.150 8.380 24.200 8.415 ;
        POLYGON 24.200 8.415 24.235 8.380 24.200 8.380 ;
        RECT 24.150 8.255 24.235 8.380 ;
        RECT 24.855 8.255 24.940 8.415 ;
        RECT 27.050 8.380 27.100 8.415 ;
        POLYGON 27.100 8.415 27.135 8.380 27.100 8.380 ;
        RECT 27.050 8.255 27.135 8.380 ;
        RECT 27.755 8.255 27.840 8.415 ;
        RECT 29.950 8.380 30.000 8.415 ;
        POLYGON 30.000 8.415 30.035 8.380 30.000 8.380 ;
        RECT 29.950 8.255 30.035 8.380 ;
        RECT 30.655 8.255 30.740 8.415 ;
        RECT 32.850 8.380 32.900 8.415 ;
        POLYGON 32.900 8.415 32.935 8.380 32.900 8.380 ;
        RECT 32.850 8.255 32.935 8.380 ;
        RECT 33.555 8.255 33.640 8.415 ;
        RECT 0.740 7.635 0.815 7.775 ;
        RECT 0.955 7.585 1.030 7.725 ;
        RECT 1.660 7.645 1.720 7.725 ;
        POLYGON 1.660 7.645 1.720 7.645 1.720 7.585 ;
        RECT 1.875 7.635 1.950 7.775 ;
        RECT 3.640 7.635 3.715 7.775 ;
        RECT 3.855 7.585 3.930 7.725 ;
        RECT 4.560 7.645 4.620 7.725 ;
        POLYGON 4.560 7.645 4.620 7.645 4.620 7.585 ;
        RECT 4.775 7.635 4.850 7.775 ;
        RECT 6.540 7.635 6.615 7.775 ;
        RECT 6.755 7.585 6.830 7.725 ;
        RECT 7.460 7.645 7.520 7.725 ;
        POLYGON 7.460 7.645 7.520 7.645 7.520 7.585 ;
        RECT 7.675 7.635 7.750 7.775 ;
        RECT 9.440 7.635 9.515 7.775 ;
        RECT 9.655 7.585 9.730 7.725 ;
        RECT 10.360 7.645 10.420 7.725 ;
        POLYGON 10.360 7.645 10.420 7.645 10.420 7.585 ;
        RECT 10.575 7.635 10.650 7.775 ;
        RECT 12.340 7.635 12.415 7.775 ;
        RECT 12.555 7.585 12.630 7.725 ;
        RECT 13.260 7.645 13.320 7.725 ;
        POLYGON 13.260 7.645 13.320 7.645 13.320 7.585 ;
        RECT 13.475 7.635 13.550 7.775 ;
        RECT 15.240 7.635 15.315 7.775 ;
        RECT 15.455 7.585 15.530 7.725 ;
        RECT 16.160 7.645 16.220 7.725 ;
        POLYGON 16.160 7.645 16.220 7.645 16.220 7.585 ;
        RECT 16.375 7.635 16.450 7.775 ;
        RECT 18.140 7.635 18.215 7.775 ;
        RECT 18.355 7.585 18.430 7.725 ;
        RECT 19.060 7.645 19.120 7.725 ;
        POLYGON 19.060 7.645 19.120 7.645 19.120 7.585 ;
        RECT 19.275 7.635 19.350 7.775 ;
        RECT 21.040 7.635 21.115 7.775 ;
        RECT 21.255 7.585 21.330 7.725 ;
        RECT 21.960 7.645 22.020 7.725 ;
        POLYGON 21.960 7.645 22.020 7.645 22.020 7.585 ;
        RECT 22.175 7.635 22.250 7.775 ;
        RECT 23.940 7.635 24.015 7.775 ;
        RECT 24.155 7.585 24.230 7.725 ;
        RECT 24.860 7.645 24.920 7.725 ;
        POLYGON 24.860 7.645 24.920 7.645 24.920 7.585 ;
        RECT 25.075 7.635 25.150 7.775 ;
        RECT 26.840 7.635 26.915 7.775 ;
        RECT 27.055 7.585 27.130 7.725 ;
        RECT 27.760 7.645 27.820 7.725 ;
        POLYGON 27.760 7.645 27.820 7.645 27.820 7.585 ;
        RECT 27.975 7.635 28.050 7.775 ;
        RECT 29.740 7.635 29.815 7.775 ;
        RECT 29.955 7.585 30.030 7.725 ;
        RECT 30.660 7.645 30.720 7.725 ;
        POLYGON 30.660 7.645 30.720 7.645 30.720 7.585 ;
        RECT 30.875 7.635 30.950 7.775 ;
        RECT 32.640 7.635 32.715 7.775 ;
        RECT 32.855 7.585 32.930 7.725 ;
        RECT 33.560 7.645 33.620 7.725 ;
        POLYGON 33.560 7.645 33.620 7.645 33.620 7.585 ;
        RECT 33.775 7.635 33.850 7.775 ;
        RECT 0.685 7.115 0.835 7.285 ;
        RECT 1.075 7.250 1.225 7.420 ;
        RECT 1.465 7.250 1.615 7.420 ;
        RECT 1.855 7.115 2.005 7.285 ;
        RECT 3.585 7.115 3.735 7.285 ;
        RECT 3.975 7.250 4.125 7.420 ;
        RECT 4.365 7.250 4.515 7.420 ;
        RECT 4.755 7.115 4.905 7.285 ;
        RECT 6.485 7.115 6.635 7.285 ;
        RECT 6.875 7.250 7.025 7.420 ;
        RECT 7.265 7.250 7.415 7.420 ;
        RECT 7.655 7.115 7.805 7.285 ;
        RECT 9.385 7.115 9.535 7.285 ;
        RECT 9.775 7.250 9.925 7.420 ;
        RECT 10.165 7.250 10.315 7.420 ;
        RECT 10.555 7.115 10.705 7.285 ;
        RECT 12.285 7.115 12.435 7.285 ;
        RECT 12.675 7.250 12.825 7.420 ;
        RECT 13.065 7.250 13.215 7.420 ;
        RECT 13.455 7.115 13.605 7.285 ;
        RECT 15.185 7.115 15.335 7.285 ;
        RECT 15.575 7.250 15.725 7.420 ;
        RECT 15.965 7.250 16.115 7.420 ;
        RECT 16.355 7.115 16.505 7.285 ;
        RECT 18.085 7.115 18.235 7.285 ;
        RECT 18.475 7.250 18.625 7.420 ;
        RECT 18.865 7.250 19.015 7.420 ;
        RECT 19.255 7.115 19.405 7.285 ;
        RECT 20.985 7.115 21.135 7.285 ;
        RECT 21.375 7.250 21.525 7.420 ;
        RECT 21.765 7.250 21.915 7.420 ;
        RECT 22.155 7.115 22.305 7.285 ;
        RECT 23.885 7.115 24.035 7.285 ;
        RECT 24.275 7.250 24.425 7.420 ;
        RECT 24.665 7.250 24.815 7.420 ;
        RECT 25.055 7.115 25.205 7.285 ;
        RECT 26.785 7.115 26.935 7.285 ;
        RECT 27.175 7.250 27.325 7.420 ;
        RECT 27.565 7.250 27.715 7.420 ;
        RECT 27.955 7.115 28.105 7.285 ;
        RECT 29.685 7.115 29.835 7.285 ;
        RECT 30.075 7.250 30.225 7.420 ;
        RECT 30.465 7.250 30.615 7.420 ;
        RECT 30.855 7.115 31.005 7.285 ;
        RECT 32.585 7.115 32.735 7.285 ;
        RECT 32.975 7.250 33.125 7.420 ;
        RECT 33.365 7.250 33.515 7.420 ;
        RECT 33.755 7.115 33.905 7.285 ;
        RECT 0.950 7.030 1.000 7.065 ;
        POLYGON 1.000 7.065 1.035 7.030 1.000 7.030 ;
        RECT 0.950 6.905 1.035 7.030 ;
        RECT 1.655 6.905 1.740 7.065 ;
        RECT 3.850 7.030 3.900 7.065 ;
        POLYGON 3.900 7.065 3.935 7.030 3.900 7.030 ;
        RECT 3.850 6.905 3.935 7.030 ;
        RECT 4.555 6.905 4.640 7.065 ;
        RECT 6.750 7.030 6.800 7.065 ;
        POLYGON 6.800 7.065 6.835 7.030 6.800 7.030 ;
        RECT 6.750 6.905 6.835 7.030 ;
        RECT 7.455 6.905 7.540 7.065 ;
        RECT 9.650 7.030 9.700 7.065 ;
        POLYGON 9.700 7.065 9.735 7.030 9.700 7.030 ;
        RECT 9.650 6.905 9.735 7.030 ;
        RECT 10.355 6.905 10.440 7.065 ;
        RECT 12.550 7.030 12.600 7.065 ;
        POLYGON 12.600 7.065 12.635 7.030 12.600 7.030 ;
        RECT 12.550 6.905 12.635 7.030 ;
        RECT 13.255 6.905 13.340 7.065 ;
        RECT 15.450 7.030 15.500 7.065 ;
        POLYGON 15.500 7.065 15.535 7.030 15.500 7.030 ;
        RECT 15.450 6.905 15.535 7.030 ;
        RECT 16.155 6.905 16.240 7.065 ;
        RECT 18.350 7.030 18.400 7.065 ;
        POLYGON 18.400 7.065 18.435 7.030 18.400 7.030 ;
        RECT 18.350 6.905 18.435 7.030 ;
        RECT 19.055 6.905 19.140 7.065 ;
        RECT 21.250 7.030 21.300 7.065 ;
        POLYGON 21.300 7.065 21.335 7.030 21.300 7.030 ;
        RECT 21.250 6.905 21.335 7.030 ;
        RECT 21.955 6.905 22.040 7.065 ;
        RECT 24.150 7.030 24.200 7.065 ;
        POLYGON 24.200 7.065 24.235 7.030 24.200 7.030 ;
        RECT 24.150 6.905 24.235 7.030 ;
        RECT 24.855 6.905 24.940 7.065 ;
        RECT 27.050 7.030 27.100 7.065 ;
        POLYGON 27.100 7.065 27.135 7.030 27.100 7.030 ;
        RECT 27.050 6.905 27.135 7.030 ;
        RECT 27.755 6.905 27.840 7.065 ;
        RECT 29.950 7.030 30.000 7.065 ;
        POLYGON 30.000 7.065 30.035 7.030 30.000 7.030 ;
        RECT 29.950 6.905 30.035 7.030 ;
        RECT 30.655 6.905 30.740 7.065 ;
        RECT 32.850 7.030 32.900 7.065 ;
        POLYGON 32.900 7.065 32.935 7.030 32.900 7.030 ;
        RECT 32.850 6.905 32.935 7.030 ;
        RECT 33.555 6.905 33.640 7.065 ;
        RECT 0.740 6.285 0.815 6.425 ;
        RECT 0.955 6.235 1.030 6.375 ;
        RECT 1.660 6.295 1.720 6.375 ;
        POLYGON 1.660 6.295 1.720 6.295 1.720 6.235 ;
        RECT 1.875 6.285 1.950 6.425 ;
        RECT 3.640 6.285 3.715 6.425 ;
        RECT 3.855 6.235 3.930 6.375 ;
        RECT 4.560 6.295 4.620 6.375 ;
        POLYGON 4.560 6.295 4.620 6.295 4.620 6.235 ;
        RECT 4.775 6.285 4.850 6.425 ;
        RECT 6.540 6.285 6.615 6.425 ;
        RECT 6.755 6.235 6.830 6.375 ;
        RECT 7.460 6.295 7.520 6.375 ;
        POLYGON 7.460 6.295 7.520 6.295 7.520 6.235 ;
        RECT 7.675 6.285 7.750 6.425 ;
        RECT 9.440 6.285 9.515 6.425 ;
        RECT 9.655 6.235 9.730 6.375 ;
        RECT 10.360 6.295 10.420 6.375 ;
        POLYGON 10.360 6.295 10.420 6.295 10.420 6.235 ;
        RECT 10.575 6.285 10.650 6.425 ;
        RECT 12.340 6.285 12.415 6.425 ;
        RECT 12.555 6.235 12.630 6.375 ;
        RECT 13.260 6.295 13.320 6.375 ;
        POLYGON 13.260 6.295 13.320 6.295 13.320 6.235 ;
        RECT 13.475 6.285 13.550 6.425 ;
        RECT 15.240 6.285 15.315 6.425 ;
        RECT 15.455 6.235 15.530 6.375 ;
        RECT 16.160 6.295 16.220 6.375 ;
        POLYGON 16.160 6.295 16.220 6.295 16.220 6.235 ;
        RECT 16.375 6.285 16.450 6.425 ;
        RECT 18.140 6.285 18.215 6.425 ;
        RECT 18.355 6.235 18.430 6.375 ;
        RECT 19.060 6.295 19.120 6.375 ;
        POLYGON 19.060 6.295 19.120 6.295 19.120 6.235 ;
        RECT 19.275 6.285 19.350 6.425 ;
        RECT 21.040 6.285 21.115 6.425 ;
        RECT 21.255 6.235 21.330 6.375 ;
        RECT 21.960 6.295 22.020 6.375 ;
        POLYGON 21.960 6.295 22.020 6.295 22.020 6.235 ;
        RECT 22.175 6.285 22.250 6.425 ;
        RECT 23.940 6.285 24.015 6.425 ;
        RECT 24.155 6.235 24.230 6.375 ;
        RECT 24.860 6.295 24.920 6.375 ;
        POLYGON 24.860 6.295 24.920 6.295 24.920 6.235 ;
        RECT 25.075 6.285 25.150 6.425 ;
        RECT 26.840 6.285 26.915 6.425 ;
        RECT 27.055 6.235 27.130 6.375 ;
        RECT 27.760 6.295 27.820 6.375 ;
        POLYGON 27.760 6.295 27.820 6.295 27.820 6.235 ;
        RECT 27.975 6.285 28.050 6.425 ;
        RECT 29.740 6.285 29.815 6.425 ;
        RECT 29.955 6.235 30.030 6.375 ;
        RECT 30.660 6.295 30.720 6.375 ;
        POLYGON 30.660 6.295 30.720 6.295 30.720 6.235 ;
        RECT 30.875 6.285 30.950 6.425 ;
        RECT 32.640 6.285 32.715 6.425 ;
        RECT 32.855 6.235 32.930 6.375 ;
        RECT 33.560 6.295 33.620 6.375 ;
        POLYGON 33.560 6.295 33.620 6.295 33.620 6.235 ;
        RECT 33.775 6.285 33.850 6.425 ;
        RECT 0.685 5.765 0.835 5.935 ;
        RECT 1.075 5.900 1.225 6.070 ;
        RECT 1.465 5.900 1.615 6.070 ;
        RECT 1.855 5.765 2.005 5.935 ;
        RECT 3.585 5.765 3.735 5.935 ;
        RECT 3.975 5.900 4.125 6.070 ;
        RECT 4.365 5.900 4.515 6.070 ;
        RECT 4.755 5.765 4.905 5.935 ;
        RECT 6.485 5.765 6.635 5.935 ;
        RECT 6.875 5.900 7.025 6.070 ;
        RECT 7.265 5.900 7.415 6.070 ;
        RECT 7.655 5.765 7.805 5.935 ;
        RECT 9.385 5.765 9.535 5.935 ;
        RECT 9.775 5.900 9.925 6.070 ;
        RECT 10.165 5.900 10.315 6.070 ;
        RECT 10.555 5.765 10.705 5.935 ;
        RECT 12.285 5.765 12.435 5.935 ;
        RECT 12.675 5.900 12.825 6.070 ;
        RECT 13.065 5.900 13.215 6.070 ;
        RECT 13.455 5.765 13.605 5.935 ;
        RECT 15.185 5.765 15.335 5.935 ;
        RECT 15.575 5.900 15.725 6.070 ;
        RECT 15.965 5.900 16.115 6.070 ;
        RECT 16.355 5.765 16.505 5.935 ;
        RECT 18.085 5.765 18.235 5.935 ;
        RECT 18.475 5.900 18.625 6.070 ;
        RECT 18.865 5.900 19.015 6.070 ;
        RECT 19.255 5.765 19.405 5.935 ;
        RECT 20.985 5.765 21.135 5.935 ;
        RECT 21.375 5.900 21.525 6.070 ;
        RECT 21.765 5.900 21.915 6.070 ;
        RECT 22.155 5.765 22.305 5.935 ;
        RECT 23.885 5.765 24.035 5.935 ;
        RECT 24.275 5.900 24.425 6.070 ;
        RECT 24.665 5.900 24.815 6.070 ;
        RECT 25.055 5.765 25.205 5.935 ;
        RECT 26.785 5.765 26.935 5.935 ;
        RECT 27.175 5.900 27.325 6.070 ;
        RECT 27.565 5.900 27.715 6.070 ;
        RECT 27.955 5.765 28.105 5.935 ;
        RECT 29.685 5.765 29.835 5.935 ;
        RECT 30.075 5.900 30.225 6.070 ;
        RECT 30.465 5.900 30.615 6.070 ;
        RECT 30.855 5.765 31.005 5.935 ;
        RECT 32.585 5.765 32.735 5.935 ;
        RECT 32.975 5.900 33.125 6.070 ;
        RECT 33.365 5.900 33.515 6.070 ;
        RECT 33.755 5.765 33.905 5.935 ;
        RECT 0.950 5.680 1.000 5.715 ;
        POLYGON 1.000 5.715 1.035 5.680 1.000 5.680 ;
        RECT 0.950 5.555 1.035 5.680 ;
        RECT 1.655 5.555 1.740 5.715 ;
        RECT 3.850 5.680 3.900 5.715 ;
        POLYGON 3.900 5.715 3.935 5.680 3.900 5.680 ;
        RECT 3.850 5.555 3.935 5.680 ;
        RECT 4.555 5.555 4.640 5.715 ;
        RECT 6.750 5.680 6.800 5.715 ;
        POLYGON 6.800 5.715 6.835 5.680 6.800 5.680 ;
        RECT 6.750 5.555 6.835 5.680 ;
        RECT 7.455 5.555 7.540 5.715 ;
        RECT 9.650 5.680 9.700 5.715 ;
        POLYGON 9.700 5.715 9.735 5.680 9.700 5.680 ;
        RECT 9.650 5.555 9.735 5.680 ;
        RECT 10.355 5.555 10.440 5.715 ;
        RECT 12.550 5.680 12.600 5.715 ;
        POLYGON 12.600 5.715 12.635 5.680 12.600 5.680 ;
        RECT 12.550 5.555 12.635 5.680 ;
        RECT 13.255 5.555 13.340 5.715 ;
        RECT 15.450 5.680 15.500 5.715 ;
        POLYGON 15.500 5.715 15.535 5.680 15.500 5.680 ;
        RECT 15.450 5.555 15.535 5.680 ;
        RECT 16.155 5.555 16.240 5.715 ;
        RECT 18.350 5.680 18.400 5.715 ;
        POLYGON 18.400 5.715 18.435 5.680 18.400 5.680 ;
        RECT 18.350 5.555 18.435 5.680 ;
        RECT 19.055 5.555 19.140 5.715 ;
        RECT 21.250 5.680 21.300 5.715 ;
        POLYGON 21.300 5.715 21.335 5.680 21.300 5.680 ;
        RECT 21.250 5.555 21.335 5.680 ;
        RECT 21.955 5.555 22.040 5.715 ;
        RECT 24.150 5.680 24.200 5.715 ;
        POLYGON 24.200 5.715 24.235 5.680 24.200 5.680 ;
        RECT 24.150 5.555 24.235 5.680 ;
        RECT 24.855 5.555 24.940 5.715 ;
        RECT 27.050 5.680 27.100 5.715 ;
        POLYGON 27.100 5.715 27.135 5.680 27.100 5.680 ;
        RECT 27.050 5.555 27.135 5.680 ;
        RECT 27.755 5.555 27.840 5.715 ;
        RECT 29.950 5.680 30.000 5.715 ;
        POLYGON 30.000 5.715 30.035 5.680 30.000 5.680 ;
        RECT 29.950 5.555 30.035 5.680 ;
        RECT 30.655 5.555 30.740 5.715 ;
        RECT 32.850 5.680 32.900 5.715 ;
        POLYGON 32.900 5.715 32.935 5.680 32.900 5.680 ;
        RECT 32.850 5.555 32.935 5.680 ;
        RECT 33.555 5.555 33.640 5.715 ;
        RECT 0.740 4.935 0.815 5.075 ;
        RECT 0.955 4.885 1.030 5.025 ;
        RECT 1.660 4.945 1.720 5.025 ;
        POLYGON 1.660 4.945 1.720 4.945 1.720 4.885 ;
        RECT 1.875 4.935 1.950 5.075 ;
        RECT 3.640 4.935 3.715 5.075 ;
        RECT 3.855 4.885 3.930 5.025 ;
        RECT 4.560 4.945 4.620 5.025 ;
        POLYGON 4.560 4.945 4.620 4.945 4.620 4.885 ;
        RECT 4.775 4.935 4.850 5.075 ;
        RECT 6.540 4.935 6.615 5.075 ;
        RECT 6.755 4.885 6.830 5.025 ;
        RECT 7.460 4.945 7.520 5.025 ;
        POLYGON 7.460 4.945 7.520 4.945 7.520 4.885 ;
        RECT 7.675 4.935 7.750 5.075 ;
        RECT 9.440 4.935 9.515 5.075 ;
        RECT 9.655 4.885 9.730 5.025 ;
        RECT 10.360 4.945 10.420 5.025 ;
        POLYGON 10.360 4.945 10.420 4.945 10.420 4.885 ;
        RECT 10.575 4.935 10.650 5.075 ;
        RECT 12.340 4.935 12.415 5.075 ;
        RECT 12.555 4.885 12.630 5.025 ;
        RECT 13.260 4.945 13.320 5.025 ;
        POLYGON 13.260 4.945 13.320 4.945 13.320 4.885 ;
        RECT 13.475 4.935 13.550 5.075 ;
        RECT 15.240 4.935 15.315 5.075 ;
        RECT 15.455 4.885 15.530 5.025 ;
        RECT 16.160 4.945 16.220 5.025 ;
        POLYGON 16.160 4.945 16.220 4.945 16.220 4.885 ;
        RECT 16.375 4.935 16.450 5.075 ;
        RECT 18.140 4.935 18.215 5.075 ;
        RECT 18.355 4.885 18.430 5.025 ;
        RECT 19.060 4.945 19.120 5.025 ;
        POLYGON 19.060 4.945 19.120 4.945 19.120 4.885 ;
        RECT 19.275 4.935 19.350 5.075 ;
        RECT 21.040 4.935 21.115 5.075 ;
        RECT 21.255 4.885 21.330 5.025 ;
        RECT 21.960 4.945 22.020 5.025 ;
        POLYGON 21.960 4.945 22.020 4.945 22.020 4.885 ;
        RECT 22.175 4.935 22.250 5.075 ;
        RECT 23.940 4.935 24.015 5.075 ;
        RECT 24.155 4.885 24.230 5.025 ;
        RECT 24.860 4.945 24.920 5.025 ;
        POLYGON 24.860 4.945 24.920 4.945 24.920 4.885 ;
        RECT 25.075 4.935 25.150 5.075 ;
        RECT 26.840 4.935 26.915 5.075 ;
        RECT 27.055 4.885 27.130 5.025 ;
        RECT 27.760 4.945 27.820 5.025 ;
        POLYGON 27.760 4.945 27.820 4.945 27.820 4.885 ;
        RECT 27.975 4.935 28.050 5.075 ;
        RECT 29.740 4.935 29.815 5.075 ;
        RECT 29.955 4.885 30.030 5.025 ;
        RECT 30.660 4.945 30.720 5.025 ;
        POLYGON 30.660 4.945 30.720 4.945 30.720 4.885 ;
        RECT 30.875 4.935 30.950 5.075 ;
        RECT 32.640 4.935 32.715 5.075 ;
        RECT 32.855 4.885 32.930 5.025 ;
        RECT 33.560 4.945 33.620 5.025 ;
        POLYGON 33.560 4.945 33.620 4.945 33.620 4.885 ;
        RECT 33.775 4.935 33.850 5.075 ;
        RECT 0.685 4.415 0.835 4.585 ;
        RECT 1.075 4.550 1.225 4.720 ;
        RECT 1.465 4.550 1.615 4.720 ;
        RECT 1.855 4.415 2.005 4.585 ;
        RECT 3.585 4.415 3.735 4.585 ;
        RECT 3.975 4.550 4.125 4.720 ;
        RECT 4.365 4.550 4.515 4.720 ;
        RECT 4.755 4.415 4.905 4.585 ;
        RECT 6.485 4.415 6.635 4.585 ;
        RECT 6.875 4.550 7.025 4.720 ;
        RECT 7.265 4.550 7.415 4.720 ;
        RECT 7.655 4.415 7.805 4.585 ;
        RECT 9.385 4.415 9.535 4.585 ;
        RECT 9.775 4.550 9.925 4.720 ;
        RECT 10.165 4.550 10.315 4.720 ;
        RECT 10.555 4.415 10.705 4.585 ;
        RECT 12.285 4.415 12.435 4.585 ;
        RECT 12.675 4.550 12.825 4.720 ;
        RECT 13.065 4.550 13.215 4.720 ;
        RECT 13.455 4.415 13.605 4.585 ;
        RECT 15.185 4.415 15.335 4.585 ;
        RECT 15.575 4.550 15.725 4.720 ;
        RECT 15.965 4.550 16.115 4.720 ;
        RECT 16.355 4.415 16.505 4.585 ;
        RECT 18.085 4.415 18.235 4.585 ;
        RECT 18.475 4.550 18.625 4.720 ;
        RECT 18.865 4.550 19.015 4.720 ;
        RECT 19.255 4.415 19.405 4.585 ;
        RECT 20.985 4.415 21.135 4.585 ;
        RECT 21.375 4.550 21.525 4.720 ;
        RECT 21.765 4.550 21.915 4.720 ;
        RECT 22.155 4.415 22.305 4.585 ;
        RECT 23.885 4.415 24.035 4.585 ;
        RECT 24.275 4.550 24.425 4.720 ;
        RECT 24.665 4.550 24.815 4.720 ;
        RECT 25.055 4.415 25.205 4.585 ;
        RECT 26.785 4.415 26.935 4.585 ;
        RECT 27.175 4.550 27.325 4.720 ;
        RECT 27.565 4.550 27.715 4.720 ;
        RECT 27.955 4.415 28.105 4.585 ;
        RECT 29.685 4.415 29.835 4.585 ;
        RECT 30.075 4.550 30.225 4.720 ;
        RECT 30.465 4.550 30.615 4.720 ;
        RECT 30.855 4.415 31.005 4.585 ;
        RECT 32.585 4.415 32.735 4.585 ;
        RECT 32.975 4.550 33.125 4.720 ;
        RECT 33.365 4.550 33.515 4.720 ;
        RECT 33.755 4.415 33.905 4.585 ;
        RECT 0.950 4.330 1.000 4.365 ;
        POLYGON 1.000 4.365 1.035 4.330 1.000 4.330 ;
        RECT 0.950 4.205 1.035 4.330 ;
        RECT 1.655 4.205 1.740 4.365 ;
        RECT 3.850 4.330 3.900 4.365 ;
        POLYGON 3.900 4.365 3.935 4.330 3.900 4.330 ;
        RECT 3.850 4.205 3.935 4.330 ;
        RECT 4.555 4.205 4.640 4.365 ;
        RECT 6.750 4.330 6.800 4.365 ;
        POLYGON 6.800 4.365 6.835 4.330 6.800 4.330 ;
        RECT 6.750 4.205 6.835 4.330 ;
        RECT 7.455 4.205 7.540 4.365 ;
        RECT 9.650 4.330 9.700 4.365 ;
        POLYGON 9.700 4.365 9.735 4.330 9.700 4.330 ;
        RECT 9.650 4.205 9.735 4.330 ;
        RECT 10.355 4.205 10.440 4.365 ;
        RECT 12.550 4.330 12.600 4.365 ;
        POLYGON 12.600 4.365 12.635 4.330 12.600 4.330 ;
        RECT 12.550 4.205 12.635 4.330 ;
        RECT 13.255 4.205 13.340 4.365 ;
        RECT 15.450 4.330 15.500 4.365 ;
        POLYGON 15.500 4.365 15.535 4.330 15.500 4.330 ;
        RECT 15.450 4.205 15.535 4.330 ;
        RECT 16.155 4.205 16.240 4.365 ;
        RECT 18.350 4.330 18.400 4.365 ;
        POLYGON 18.400 4.365 18.435 4.330 18.400 4.330 ;
        RECT 18.350 4.205 18.435 4.330 ;
        RECT 19.055 4.205 19.140 4.365 ;
        RECT 21.250 4.330 21.300 4.365 ;
        POLYGON 21.300 4.365 21.335 4.330 21.300 4.330 ;
        RECT 21.250 4.205 21.335 4.330 ;
        RECT 21.955 4.205 22.040 4.365 ;
        RECT 24.150 4.330 24.200 4.365 ;
        POLYGON 24.200 4.365 24.235 4.330 24.200 4.330 ;
        RECT 24.150 4.205 24.235 4.330 ;
        RECT 24.855 4.205 24.940 4.365 ;
        RECT 27.050 4.330 27.100 4.365 ;
        POLYGON 27.100 4.365 27.135 4.330 27.100 4.330 ;
        RECT 27.050 4.205 27.135 4.330 ;
        RECT 27.755 4.205 27.840 4.365 ;
        RECT 29.950 4.330 30.000 4.365 ;
        POLYGON 30.000 4.365 30.035 4.330 30.000 4.330 ;
        RECT 29.950 4.205 30.035 4.330 ;
        RECT 30.655 4.205 30.740 4.365 ;
        RECT 32.850 4.330 32.900 4.365 ;
        POLYGON 32.900 4.365 32.935 4.330 32.900 4.330 ;
        RECT 32.850 4.205 32.935 4.330 ;
        RECT 33.555 4.205 33.640 4.365 ;
        RECT 0.740 3.585 0.815 3.725 ;
        RECT 0.955 3.535 1.030 3.675 ;
        RECT 1.660 3.595 1.720 3.675 ;
        POLYGON 1.660 3.595 1.720 3.595 1.720 3.535 ;
        RECT 1.875 3.585 1.950 3.725 ;
        RECT 3.640 3.585 3.715 3.725 ;
        RECT 3.855 3.535 3.930 3.675 ;
        RECT 4.560 3.595 4.620 3.675 ;
        POLYGON 4.560 3.595 4.620 3.595 4.620 3.535 ;
        RECT 4.775 3.585 4.850 3.725 ;
        RECT 6.540 3.585 6.615 3.725 ;
        RECT 6.755 3.535 6.830 3.675 ;
        RECT 7.460 3.595 7.520 3.675 ;
        POLYGON 7.460 3.595 7.520 3.595 7.520 3.535 ;
        RECT 7.675 3.585 7.750 3.725 ;
        RECT 9.440 3.585 9.515 3.725 ;
        RECT 9.655 3.535 9.730 3.675 ;
        RECT 10.360 3.595 10.420 3.675 ;
        POLYGON 10.360 3.595 10.420 3.595 10.420 3.535 ;
        RECT 10.575 3.585 10.650 3.725 ;
        RECT 12.340 3.585 12.415 3.725 ;
        RECT 12.555 3.535 12.630 3.675 ;
        RECT 13.260 3.595 13.320 3.675 ;
        POLYGON 13.260 3.595 13.320 3.595 13.320 3.535 ;
        RECT 13.475 3.585 13.550 3.725 ;
        RECT 15.240 3.585 15.315 3.725 ;
        RECT 15.455 3.535 15.530 3.675 ;
        RECT 16.160 3.595 16.220 3.675 ;
        POLYGON 16.160 3.595 16.220 3.595 16.220 3.535 ;
        RECT 16.375 3.585 16.450 3.725 ;
        RECT 18.140 3.585 18.215 3.725 ;
        RECT 18.355 3.535 18.430 3.675 ;
        RECT 19.060 3.595 19.120 3.675 ;
        POLYGON 19.060 3.595 19.120 3.595 19.120 3.535 ;
        RECT 19.275 3.585 19.350 3.725 ;
        RECT 21.040 3.585 21.115 3.725 ;
        RECT 21.255 3.535 21.330 3.675 ;
        RECT 21.960 3.595 22.020 3.675 ;
        POLYGON 21.960 3.595 22.020 3.595 22.020 3.535 ;
        RECT 22.175 3.585 22.250 3.725 ;
        RECT 23.940 3.585 24.015 3.725 ;
        RECT 24.155 3.535 24.230 3.675 ;
        RECT 24.860 3.595 24.920 3.675 ;
        POLYGON 24.860 3.595 24.920 3.595 24.920 3.535 ;
        RECT 25.075 3.585 25.150 3.725 ;
        RECT 26.840 3.585 26.915 3.725 ;
        RECT 27.055 3.535 27.130 3.675 ;
        RECT 27.760 3.595 27.820 3.675 ;
        POLYGON 27.760 3.595 27.820 3.595 27.820 3.535 ;
        RECT 27.975 3.585 28.050 3.725 ;
        RECT 29.740 3.585 29.815 3.725 ;
        RECT 29.955 3.535 30.030 3.675 ;
        RECT 30.660 3.595 30.720 3.675 ;
        POLYGON 30.660 3.595 30.720 3.595 30.720 3.535 ;
        RECT 30.875 3.585 30.950 3.725 ;
        RECT 32.640 3.585 32.715 3.725 ;
        RECT 32.855 3.535 32.930 3.675 ;
        RECT 33.560 3.595 33.620 3.675 ;
        POLYGON 33.560 3.595 33.620 3.595 33.620 3.535 ;
        RECT 33.775 3.585 33.850 3.725 ;
        RECT 0.685 3.065 0.835 3.235 ;
        RECT 1.075 3.200 1.225 3.370 ;
        RECT 1.465 3.200 1.615 3.370 ;
        RECT 1.855 3.065 2.005 3.235 ;
        RECT 3.585 3.065 3.735 3.235 ;
        RECT 3.975 3.200 4.125 3.370 ;
        RECT 4.365 3.200 4.515 3.370 ;
        RECT 4.755 3.065 4.905 3.235 ;
        RECT 6.485 3.065 6.635 3.235 ;
        RECT 6.875 3.200 7.025 3.370 ;
        RECT 7.265 3.200 7.415 3.370 ;
        RECT 7.655 3.065 7.805 3.235 ;
        RECT 9.385 3.065 9.535 3.235 ;
        RECT 9.775 3.200 9.925 3.370 ;
        RECT 10.165 3.200 10.315 3.370 ;
        RECT 10.555 3.065 10.705 3.235 ;
        RECT 12.285 3.065 12.435 3.235 ;
        RECT 12.675 3.200 12.825 3.370 ;
        RECT 13.065 3.200 13.215 3.370 ;
        RECT 13.455 3.065 13.605 3.235 ;
        RECT 15.185 3.065 15.335 3.235 ;
        RECT 15.575 3.200 15.725 3.370 ;
        RECT 15.965 3.200 16.115 3.370 ;
        RECT 16.355 3.065 16.505 3.235 ;
        RECT 18.085 3.065 18.235 3.235 ;
        RECT 18.475 3.200 18.625 3.370 ;
        RECT 18.865 3.200 19.015 3.370 ;
        RECT 19.255 3.065 19.405 3.235 ;
        RECT 20.985 3.065 21.135 3.235 ;
        RECT 21.375 3.200 21.525 3.370 ;
        RECT 21.765 3.200 21.915 3.370 ;
        RECT 22.155 3.065 22.305 3.235 ;
        RECT 23.885 3.065 24.035 3.235 ;
        RECT 24.275 3.200 24.425 3.370 ;
        RECT 24.665 3.200 24.815 3.370 ;
        RECT 25.055 3.065 25.205 3.235 ;
        RECT 26.785 3.065 26.935 3.235 ;
        RECT 27.175 3.200 27.325 3.370 ;
        RECT 27.565 3.200 27.715 3.370 ;
        RECT 27.955 3.065 28.105 3.235 ;
        RECT 29.685 3.065 29.835 3.235 ;
        RECT 30.075 3.200 30.225 3.370 ;
        RECT 30.465 3.200 30.615 3.370 ;
        RECT 30.855 3.065 31.005 3.235 ;
        RECT 32.585 3.065 32.735 3.235 ;
        RECT 32.975 3.200 33.125 3.370 ;
        RECT 33.365 3.200 33.515 3.370 ;
        RECT 33.755 3.065 33.905 3.235 ;
        RECT 0.950 2.980 1.000 3.015 ;
        POLYGON 1.000 3.015 1.035 2.980 1.000 2.980 ;
        RECT 0.950 2.855 1.035 2.980 ;
        RECT 1.655 2.855 1.740 3.015 ;
        RECT 3.850 2.980 3.900 3.015 ;
        POLYGON 3.900 3.015 3.935 2.980 3.900 2.980 ;
        RECT 3.850 2.855 3.935 2.980 ;
        RECT 4.555 2.855 4.640 3.015 ;
        RECT 6.750 2.980 6.800 3.015 ;
        POLYGON 6.800 3.015 6.835 2.980 6.800 2.980 ;
        RECT 6.750 2.855 6.835 2.980 ;
        RECT 7.455 2.855 7.540 3.015 ;
        RECT 9.650 2.980 9.700 3.015 ;
        POLYGON 9.700 3.015 9.735 2.980 9.700 2.980 ;
        RECT 9.650 2.855 9.735 2.980 ;
        RECT 10.355 2.855 10.440 3.015 ;
        RECT 12.550 2.980 12.600 3.015 ;
        POLYGON 12.600 3.015 12.635 2.980 12.600 2.980 ;
        RECT 12.550 2.855 12.635 2.980 ;
        RECT 13.255 2.855 13.340 3.015 ;
        RECT 15.450 2.980 15.500 3.015 ;
        POLYGON 15.500 3.015 15.535 2.980 15.500 2.980 ;
        RECT 15.450 2.855 15.535 2.980 ;
        RECT 16.155 2.855 16.240 3.015 ;
        RECT 18.350 2.980 18.400 3.015 ;
        POLYGON 18.400 3.015 18.435 2.980 18.400 2.980 ;
        RECT 18.350 2.855 18.435 2.980 ;
        RECT 19.055 2.855 19.140 3.015 ;
        RECT 21.250 2.980 21.300 3.015 ;
        POLYGON 21.300 3.015 21.335 2.980 21.300 2.980 ;
        RECT 21.250 2.855 21.335 2.980 ;
        RECT 21.955 2.855 22.040 3.015 ;
        RECT 24.150 2.980 24.200 3.015 ;
        POLYGON 24.200 3.015 24.235 2.980 24.200 2.980 ;
        RECT 24.150 2.855 24.235 2.980 ;
        RECT 24.855 2.855 24.940 3.015 ;
        RECT 27.050 2.980 27.100 3.015 ;
        POLYGON 27.100 3.015 27.135 2.980 27.100 2.980 ;
        RECT 27.050 2.855 27.135 2.980 ;
        RECT 27.755 2.855 27.840 3.015 ;
        RECT 29.950 2.980 30.000 3.015 ;
        POLYGON 30.000 3.015 30.035 2.980 30.000 2.980 ;
        RECT 29.950 2.855 30.035 2.980 ;
        RECT 30.655 2.855 30.740 3.015 ;
        RECT 32.850 2.980 32.900 3.015 ;
        POLYGON 32.900 3.015 32.935 2.980 32.900 2.980 ;
        RECT 32.850 2.855 32.935 2.980 ;
        RECT 33.555 2.855 33.640 3.015 ;
        RECT 0.740 2.235 0.815 2.375 ;
        RECT 0.955 2.185 1.030 2.325 ;
        RECT 1.660 2.245 1.720 2.325 ;
        POLYGON 1.660 2.245 1.720 2.245 1.720 2.185 ;
        RECT 1.875 2.235 1.950 2.375 ;
        RECT 3.640 2.235 3.715 2.375 ;
        RECT 3.855 2.185 3.930 2.325 ;
        RECT 4.560 2.245 4.620 2.325 ;
        POLYGON 4.560 2.245 4.620 2.245 4.620 2.185 ;
        RECT 4.775 2.235 4.850 2.375 ;
        RECT 6.540 2.235 6.615 2.375 ;
        RECT 6.755 2.185 6.830 2.325 ;
        RECT 7.460 2.245 7.520 2.325 ;
        POLYGON 7.460 2.245 7.520 2.245 7.520 2.185 ;
        RECT 7.675 2.235 7.750 2.375 ;
        RECT 9.440 2.235 9.515 2.375 ;
        RECT 9.655 2.185 9.730 2.325 ;
        RECT 10.360 2.245 10.420 2.325 ;
        POLYGON 10.360 2.245 10.420 2.245 10.420 2.185 ;
        RECT 10.575 2.235 10.650 2.375 ;
        RECT 12.340 2.235 12.415 2.375 ;
        RECT 12.555 2.185 12.630 2.325 ;
        RECT 13.260 2.245 13.320 2.325 ;
        POLYGON 13.260 2.245 13.320 2.245 13.320 2.185 ;
        RECT 13.475 2.235 13.550 2.375 ;
        RECT 15.240 2.235 15.315 2.375 ;
        RECT 15.455 2.185 15.530 2.325 ;
        RECT 16.160 2.245 16.220 2.325 ;
        POLYGON 16.160 2.245 16.220 2.245 16.220 2.185 ;
        RECT 16.375 2.235 16.450 2.375 ;
        RECT 18.140 2.235 18.215 2.375 ;
        RECT 18.355 2.185 18.430 2.325 ;
        RECT 19.060 2.245 19.120 2.325 ;
        POLYGON 19.060 2.245 19.120 2.245 19.120 2.185 ;
        RECT 19.275 2.235 19.350 2.375 ;
        RECT 21.040 2.235 21.115 2.375 ;
        RECT 21.255 2.185 21.330 2.325 ;
        RECT 21.960 2.245 22.020 2.325 ;
        POLYGON 21.960 2.245 22.020 2.245 22.020 2.185 ;
        RECT 22.175 2.235 22.250 2.375 ;
        RECT 23.940 2.235 24.015 2.375 ;
        RECT 24.155 2.185 24.230 2.325 ;
        RECT 24.860 2.245 24.920 2.325 ;
        POLYGON 24.860 2.245 24.920 2.245 24.920 2.185 ;
        RECT 25.075 2.235 25.150 2.375 ;
        RECT 26.840 2.235 26.915 2.375 ;
        RECT 27.055 2.185 27.130 2.325 ;
        RECT 27.760 2.245 27.820 2.325 ;
        POLYGON 27.760 2.245 27.820 2.245 27.820 2.185 ;
        RECT 27.975 2.235 28.050 2.375 ;
        RECT 29.740 2.235 29.815 2.375 ;
        RECT 29.955 2.185 30.030 2.325 ;
        RECT 30.660 2.245 30.720 2.325 ;
        POLYGON 30.660 2.245 30.720 2.245 30.720 2.185 ;
        RECT 30.875 2.235 30.950 2.375 ;
        RECT 32.640 2.235 32.715 2.375 ;
        RECT 32.855 2.185 32.930 2.325 ;
        RECT 33.560 2.245 33.620 2.325 ;
        POLYGON 33.560 2.245 33.620 2.245 33.620 2.185 ;
        RECT 33.775 2.235 33.850 2.375 ;
        RECT 0.685 1.715 0.835 1.885 ;
        RECT 1.075 1.850 1.225 2.020 ;
        RECT 1.465 1.850 1.615 2.020 ;
        RECT 1.855 1.715 2.005 1.885 ;
        RECT 3.585 1.715 3.735 1.885 ;
        RECT 3.975 1.850 4.125 2.020 ;
        RECT 4.365 1.850 4.515 2.020 ;
        RECT 4.755 1.715 4.905 1.885 ;
        RECT 6.485 1.715 6.635 1.885 ;
        RECT 6.875 1.850 7.025 2.020 ;
        RECT 7.265 1.850 7.415 2.020 ;
        RECT 7.655 1.715 7.805 1.885 ;
        RECT 9.385 1.715 9.535 1.885 ;
        RECT 9.775 1.850 9.925 2.020 ;
        RECT 10.165 1.850 10.315 2.020 ;
        RECT 10.555 1.715 10.705 1.885 ;
        RECT 12.285 1.715 12.435 1.885 ;
        RECT 12.675 1.850 12.825 2.020 ;
        RECT 13.065 1.850 13.215 2.020 ;
        RECT 13.455 1.715 13.605 1.885 ;
        RECT 15.185 1.715 15.335 1.885 ;
        RECT 15.575 1.850 15.725 2.020 ;
        RECT 15.965 1.850 16.115 2.020 ;
        RECT 16.355 1.715 16.505 1.885 ;
        RECT 18.085 1.715 18.235 1.885 ;
        RECT 18.475 1.850 18.625 2.020 ;
        RECT 18.865 1.850 19.015 2.020 ;
        RECT 19.255 1.715 19.405 1.885 ;
        RECT 20.985 1.715 21.135 1.885 ;
        RECT 21.375 1.850 21.525 2.020 ;
        RECT 21.765 1.850 21.915 2.020 ;
        RECT 22.155 1.715 22.305 1.885 ;
        RECT 23.885 1.715 24.035 1.885 ;
        RECT 24.275 1.850 24.425 2.020 ;
        RECT 24.665 1.850 24.815 2.020 ;
        RECT 25.055 1.715 25.205 1.885 ;
        RECT 26.785 1.715 26.935 1.885 ;
        RECT 27.175 1.850 27.325 2.020 ;
        RECT 27.565 1.850 27.715 2.020 ;
        RECT 27.955 1.715 28.105 1.885 ;
        RECT 29.685 1.715 29.835 1.885 ;
        RECT 30.075 1.850 30.225 2.020 ;
        RECT 30.465 1.850 30.615 2.020 ;
        RECT 30.855 1.715 31.005 1.885 ;
        RECT 32.585 1.715 32.735 1.885 ;
        RECT 32.975 1.850 33.125 2.020 ;
        RECT 33.365 1.850 33.515 2.020 ;
        RECT 33.755 1.715 33.905 1.885 ;
        RECT 0.950 1.630 1.000 1.665 ;
        POLYGON 1.000 1.665 1.035 1.630 1.000 1.630 ;
        RECT 0.950 1.505 1.035 1.630 ;
        RECT 1.655 1.505 1.740 1.665 ;
        RECT 3.850 1.630 3.900 1.665 ;
        POLYGON 3.900 1.665 3.935 1.630 3.900 1.630 ;
        RECT 3.850 1.505 3.935 1.630 ;
        RECT 4.555 1.505 4.640 1.665 ;
        RECT 6.750 1.630 6.800 1.665 ;
        POLYGON 6.800 1.665 6.835 1.630 6.800 1.630 ;
        RECT 6.750 1.505 6.835 1.630 ;
        RECT 7.455 1.505 7.540 1.665 ;
        RECT 9.650 1.630 9.700 1.665 ;
        POLYGON 9.700 1.665 9.735 1.630 9.700 1.630 ;
        RECT 9.650 1.505 9.735 1.630 ;
        RECT 10.355 1.505 10.440 1.665 ;
        RECT 12.550 1.630 12.600 1.665 ;
        POLYGON 12.600 1.665 12.635 1.630 12.600 1.630 ;
        RECT 12.550 1.505 12.635 1.630 ;
        RECT 13.255 1.505 13.340 1.665 ;
        RECT 15.450 1.630 15.500 1.665 ;
        POLYGON 15.500 1.665 15.535 1.630 15.500 1.630 ;
        RECT 15.450 1.505 15.535 1.630 ;
        RECT 16.155 1.505 16.240 1.665 ;
        RECT 18.350 1.630 18.400 1.665 ;
        POLYGON 18.400 1.665 18.435 1.630 18.400 1.630 ;
        RECT 18.350 1.505 18.435 1.630 ;
        RECT 19.055 1.505 19.140 1.665 ;
        RECT 21.250 1.630 21.300 1.665 ;
        POLYGON 21.300 1.665 21.335 1.630 21.300 1.630 ;
        RECT 21.250 1.505 21.335 1.630 ;
        RECT 21.955 1.505 22.040 1.665 ;
        RECT 24.150 1.630 24.200 1.665 ;
        POLYGON 24.200 1.665 24.235 1.630 24.200 1.630 ;
        RECT 24.150 1.505 24.235 1.630 ;
        RECT 24.855 1.505 24.940 1.665 ;
        RECT 27.050 1.630 27.100 1.665 ;
        POLYGON 27.100 1.665 27.135 1.630 27.100 1.630 ;
        RECT 27.050 1.505 27.135 1.630 ;
        RECT 27.755 1.505 27.840 1.665 ;
        RECT 29.950 1.630 30.000 1.665 ;
        POLYGON 30.000 1.665 30.035 1.630 30.000 1.630 ;
        RECT 29.950 1.505 30.035 1.630 ;
        RECT 30.655 1.505 30.740 1.665 ;
        RECT 32.850 1.630 32.900 1.665 ;
        POLYGON 32.900 1.665 32.935 1.630 32.900 1.630 ;
        RECT 32.850 1.505 32.935 1.630 ;
        RECT 33.555 1.505 33.640 1.665 ;
        RECT 0.740 0.885 0.815 1.025 ;
        RECT 0.955 0.835 1.030 0.975 ;
        RECT 1.660 0.895 1.720 0.975 ;
        POLYGON 1.660 0.895 1.720 0.895 1.720 0.835 ;
        RECT 1.875 0.885 1.950 1.025 ;
        RECT 3.640 0.885 3.715 1.025 ;
        RECT 3.855 0.835 3.930 0.975 ;
        RECT 4.560 0.895 4.620 0.975 ;
        POLYGON 4.560 0.895 4.620 0.895 4.620 0.835 ;
        RECT 4.775 0.885 4.850 1.025 ;
        RECT 6.540 0.885 6.615 1.025 ;
        RECT 6.755 0.835 6.830 0.975 ;
        RECT 7.460 0.895 7.520 0.975 ;
        POLYGON 7.460 0.895 7.520 0.895 7.520 0.835 ;
        RECT 7.675 0.885 7.750 1.025 ;
        RECT 9.440 0.885 9.515 1.025 ;
        RECT 9.655 0.835 9.730 0.975 ;
        RECT 10.360 0.895 10.420 0.975 ;
        POLYGON 10.360 0.895 10.420 0.895 10.420 0.835 ;
        RECT 10.575 0.885 10.650 1.025 ;
        RECT 12.340 0.885 12.415 1.025 ;
        RECT 12.555 0.835 12.630 0.975 ;
        RECT 13.260 0.895 13.320 0.975 ;
        POLYGON 13.260 0.895 13.320 0.895 13.320 0.835 ;
        RECT 13.475 0.885 13.550 1.025 ;
        RECT 15.240 0.885 15.315 1.025 ;
        RECT 15.455 0.835 15.530 0.975 ;
        RECT 16.160 0.895 16.220 0.975 ;
        POLYGON 16.160 0.895 16.220 0.895 16.220 0.835 ;
        RECT 16.375 0.885 16.450 1.025 ;
        RECT 18.140 0.885 18.215 1.025 ;
        RECT 18.355 0.835 18.430 0.975 ;
        RECT 19.060 0.895 19.120 0.975 ;
        POLYGON 19.060 0.895 19.120 0.895 19.120 0.835 ;
        RECT 19.275 0.885 19.350 1.025 ;
        RECT 21.040 0.885 21.115 1.025 ;
        RECT 21.255 0.835 21.330 0.975 ;
        RECT 21.960 0.895 22.020 0.975 ;
        POLYGON 21.960 0.895 22.020 0.895 22.020 0.835 ;
        RECT 22.175 0.885 22.250 1.025 ;
        RECT 23.940 0.885 24.015 1.025 ;
        RECT 24.155 0.835 24.230 0.975 ;
        RECT 24.860 0.895 24.920 0.975 ;
        POLYGON 24.860 0.895 24.920 0.895 24.920 0.835 ;
        RECT 25.075 0.885 25.150 1.025 ;
        RECT 26.840 0.885 26.915 1.025 ;
        RECT 27.055 0.835 27.130 0.975 ;
        RECT 27.760 0.895 27.820 0.975 ;
        POLYGON 27.760 0.895 27.820 0.895 27.820 0.835 ;
        RECT 27.975 0.885 28.050 1.025 ;
        RECT 29.740 0.885 29.815 1.025 ;
        RECT 29.955 0.835 30.030 0.975 ;
        RECT 30.660 0.895 30.720 0.975 ;
        POLYGON 30.660 0.895 30.720 0.895 30.720 0.835 ;
        RECT 30.875 0.885 30.950 1.025 ;
        RECT 32.640 0.885 32.715 1.025 ;
        RECT 32.855 0.835 32.930 0.975 ;
        RECT 33.560 0.895 33.620 0.975 ;
        POLYGON 33.560 0.895 33.620 0.895 33.620 0.835 ;
        RECT 33.775 0.885 33.850 1.025 ;
        RECT 0.685 0.365 0.835 0.535 ;
        RECT 1.075 0.500 1.225 0.670 ;
        RECT 1.465 0.500 1.615 0.670 ;
        RECT 1.855 0.365 2.005 0.535 ;
        RECT 3.585 0.365 3.735 0.535 ;
        RECT 3.975 0.500 4.125 0.670 ;
        RECT 4.365 0.500 4.515 0.670 ;
        RECT 4.755 0.365 4.905 0.535 ;
        RECT 6.485 0.365 6.635 0.535 ;
        RECT 6.875 0.500 7.025 0.670 ;
        RECT 7.265 0.500 7.415 0.670 ;
        RECT 7.655 0.365 7.805 0.535 ;
        RECT 9.385 0.365 9.535 0.535 ;
        RECT 9.775 0.500 9.925 0.670 ;
        RECT 10.165 0.500 10.315 0.670 ;
        RECT 10.555 0.365 10.705 0.535 ;
        RECT 12.285 0.365 12.435 0.535 ;
        RECT 12.675 0.500 12.825 0.670 ;
        RECT 13.065 0.500 13.215 0.670 ;
        RECT 13.455 0.365 13.605 0.535 ;
        RECT 15.185 0.365 15.335 0.535 ;
        RECT 15.575 0.500 15.725 0.670 ;
        RECT 15.965 0.500 16.115 0.670 ;
        RECT 16.355 0.365 16.505 0.535 ;
        RECT 18.085 0.365 18.235 0.535 ;
        RECT 18.475 0.500 18.625 0.670 ;
        RECT 18.865 0.500 19.015 0.670 ;
        RECT 19.255 0.365 19.405 0.535 ;
        RECT 20.985 0.365 21.135 0.535 ;
        RECT 21.375 0.500 21.525 0.670 ;
        RECT 21.765 0.500 21.915 0.670 ;
        RECT 22.155 0.365 22.305 0.535 ;
        RECT 23.885 0.365 24.035 0.535 ;
        RECT 24.275 0.500 24.425 0.670 ;
        RECT 24.665 0.500 24.815 0.670 ;
        RECT 25.055 0.365 25.205 0.535 ;
        RECT 26.785 0.365 26.935 0.535 ;
        RECT 27.175 0.500 27.325 0.670 ;
        RECT 27.565 0.500 27.715 0.670 ;
        RECT 27.955 0.365 28.105 0.535 ;
        RECT 29.685 0.365 29.835 0.535 ;
        RECT 30.075 0.500 30.225 0.670 ;
        RECT 30.465 0.500 30.615 0.670 ;
        RECT 30.855 0.365 31.005 0.535 ;
        RECT 32.585 0.365 32.735 0.535 ;
        RECT 32.975 0.500 33.125 0.670 ;
        RECT 33.365 0.500 33.515 0.670 ;
        RECT 33.755 0.365 33.905 0.535 ;
        RECT 0.950 0.280 1.000 0.315 ;
        POLYGON 1.000 0.315 1.035 0.280 1.000 0.280 ;
        RECT 0.950 0.155 1.035 0.280 ;
        RECT 1.655 0.155 1.740 0.315 ;
        RECT 3.850 0.280 3.900 0.315 ;
        POLYGON 3.900 0.315 3.935 0.280 3.900 0.280 ;
        RECT 3.850 0.155 3.935 0.280 ;
        RECT 4.555 0.155 4.640 0.315 ;
        RECT 6.750 0.280 6.800 0.315 ;
        POLYGON 6.800 0.315 6.835 0.280 6.800 0.280 ;
        RECT 6.750 0.155 6.835 0.280 ;
        RECT 7.455 0.155 7.540 0.315 ;
        RECT 9.650 0.280 9.700 0.315 ;
        POLYGON 9.700 0.315 9.735 0.280 9.700 0.280 ;
        RECT 9.650 0.155 9.735 0.280 ;
        RECT 10.355 0.155 10.440 0.315 ;
        RECT 12.550 0.280 12.600 0.315 ;
        POLYGON 12.600 0.315 12.635 0.280 12.600 0.280 ;
        RECT 12.550 0.155 12.635 0.280 ;
        RECT 13.255 0.155 13.340 0.315 ;
        RECT 15.450 0.280 15.500 0.315 ;
        POLYGON 15.500 0.315 15.535 0.280 15.500 0.280 ;
        RECT 15.450 0.155 15.535 0.280 ;
        RECT 16.155 0.155 16.240 0.315 ;
        RECT 18.350 0.280 18.400 0.315 ;
        POLYGON 18.400 0.315 18.435 0.280 18.400 0.280 ;
        RECT 18.350 0.155 18.435 0.280 ;
        RECT 19.055 0.155 19.140 0.315 ;
        RECT 21.250 0.280 21.300 0.315 ;
        POLYGON 21.300 0.315 21.335 0.280 21.300 0.280 ;
        RECT 21.250 0.155 21.335 0.280 ;
        RECT 21.955 0.155 22.040 0.315 ;
        RECT 24.150 0.280 24.200 0.315 ;
        POLYGON 24.200 0.315 24.235 0.280 24.200 0.280 ;
        RECT 24.150 0.155 24.235 0.280 ;
        RECT 24.855 0.155 24.940 0.315 ;
        RECT 27.050 0.280 27.100 0.315 ;
        POLYGON 27.100 0.315 27.135 0.280 27.100 0.280 ;
        RECT 27.050 0.155 27.135 0.280 ;
        RECT 27.755 0.155 27.840 0.315 ;
        RECT 29.950 0.280 30.000 0.315 ;
        POLYGON 30.000 0.315 30.035 0.280 30.000 0.280 ;
        RECT 29.950 0.155 30.035 0.280 ;
        RECT 30.655 0.155 30.740 0.315 ;
        RECT 32.850 0.280 32.900 0.315 ;
        POLYGON 32.900 0.315 32.935 0.280 32.900 0.280 ;
        RECT 32.850 0.155 32.935 0.280 ;
        RECT 33.555 0.155 33.640 0.315 ;
  END
END 10T_16x12_2r1w_magic_flattened
END LIBRARY

