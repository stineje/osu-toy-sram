magic
tech sky130A
magscale 1 2
timestamp 1658445342
<< error_s >>
rect 15 8624 28 8640
rect 117 8638 130 8640
rect 83 8624 98 8638
rect 107 8624 137 8638
rect 198 8636 351 8682
rect 180 8624 372 8636
rect 415 8624 445 8638
rect 451 8624 464 8640
rect 552 8624 565 8640
rect 595 8624 608 8640
rect 697 8638 710 8640
rect 663 8624 678 8638
rect 687 8624 717 8638
rect 778 8636 931 8682
rect 760 8624 952 8636
rect 995 8624 1025 8638
rect 1031 8624 1044 8640
rect 1132 8624 1145 8640
rect 1175 8624 1188 8640
rect 1277 8638 1290 8640
rect 1243 8624 1258 8638
rect 1267 8624 1297 8638
rect 1358 8636 1511 8682
rect 1340 8624 1532 8636
rect 1575 8624 1605 8638
rect 1611 8624 1624 8640
rect 1712 8624 1725 8640
rect 1755 8624 1768 8640
rect 1857 8638 1870 8640
rect 1823 8624 1838 8638
rect 1847 8624 1877 8638
rect 1938 8636 2091 8682
rect 1920 8624 2112 8636
rect 2155 8624 2185 8638
rect 2191 8624 2204 8640
rect 2292 8624 2305 8640
rect 2335 8624 2348 8640
rect 2437 8638 2450 8640
rect 2403 8624 2418 8638
rect 2427 8624 2457 8638
rect 2518 8636 2671 8682
rect 2500 8624 2692 8636
rect 2735 8624 2765 8638
rect 2771 8624 2784 8640
rect 2872 8624 2885 8640
rect 2915 8624 2928 8640
rect 3017 8638 3030 8640
rect 2983 8624 2998 8638
rect 3007 8624 3037 8638
rect 3098 8636 3251 8682
rect 3080 8624 3272 8636
rect 3315 8624 3345 8638
rect 3351 8624 3364 8640
rect 3452 8624 3465 8640
rect 3495 8624 3508 8640
rect 3597 8638 3610 8640
rect 3563 8624 3578 8638
rect 3587 8624 3617 8638
rect 3678 8636 3831 8682
rect 3660 8624 3852 8636
rect 3895 8624 3925 8638
rect 3931 8624 3944 8640
rect 4032 8624 4045 8640
rect 4075 8624 4088 8640
rect 4177 8638 4190 8640
rect 4143 8624 4158 8638
rect 4167 8624 4197 8638
rect 4258 8636 4411 8682
rect 4240 8624 4432 8636
rect 4475 8624 4505 8638
rect 4511 8624 4524 8640
rect 4612 8624 4625 8640
rect 4655 8624 4668 8640
rect 4757 8638 4770 8640
rect 4723 8624 4738 8638
rect 4747 8624 4777 8638
rect 4838 8636 4991 8682
rect 4820 8624 5012 8636
rect 5055 8624 5085 8638
rect 5091 8624 5104 8640
rect 5192 8624 5205 8640
rect 5235 8624 5248 8640
rect 5337 8638 5350 8640
rect 5303 8624 5318 8638
rect 5327 8624 5357 8638
rect 5418 8636 5571 8682
rect 5400 8624 5592 8636
rect 5635 8624 5665 8638
rect 5671 8624 5684 8640
rect 5772 8624 5785 8640
rect 5815 8624 5828 8640
rect 5917 8638 5930 8640
rect 5883 8624 5898 8638
rect 5907 8624 5937 8638
rect 5998 8636 6151 8682
rect 5980 8624 6172 8636
rect 6215 8624 6245 8638
rect 6251 8624 6264 8640
rect 6352 8624 6365 8640
rect 6395 8624 6408 8640
rect 6497 8638 6510 8640
rect 6463 8624 6478 8638
rect 6487 8624 6517 8638
rect 6578 8636 6731 8682
rect 6560 8624 6752 8636
rect 6795 8624 6825 8638
rect 6831 8624 6844 8640
rect 6932 8624 6945 8640
rect 6975 8624 6988 8640
rect 7077 8638 7090 8640
rect 7043 8624 7058 8638
rect 7067 8624 7097 8638
rect 7158 8636 7311 8682
rect 7140 8624 7332 8636
rect 7375 8624 7405 8638
rect 7411 8624 7424 8640
rect 7512 8624 7525 8640
rect 7555 8624 7568 8640
rect 7657 8638 7670 8640
rect 7623 8624 7638 8638
rect 7647 8624 7677 8638
rect 7738 8636 7891 8682
rect 7720 8624 7912 8636
rect 7955 8624 7985 8638
rect 7991 8624 8004 8640
rect 8092 8624 8105 8640
rect 8135 8624 8148 8640
rect 8237 8638 8250 8640
rect 8203 8624 8218 8638
rect 8227 8624 8257 8638
rect 8318 8636 8471 8682
rect 8300 8624 8492 8636
rect 8535 8624 8565 8638
rect 8571 8624 8584 8640
rect 8672 8624 8685 8640
rect 8715 8624 8728 8640
rect 8817 8638 8830 8640
rect 8783 8624 8798 8638
rect 8807 8624 8837 8638
rect 8898 8636 9051 8682
rect 8880 8624 9072 8636
rect 9115 8624 9145 8638
rect 9151 8624 9164 8640
rect 9252 8624 9265 8640
rect 0 8610 9265 8624
rect 15 8506 28 8610
rect 73 8588 74 8598
rect 89 8588 102 8598
rect 73 8584 102 8588
rect 107 8584 137 8610
rect 155 8596 171 8598
rect 243 8596 296 8610
rect 244 8594 308 8596
rect 351 8594 366 8610
rect 415 8607 445 8610
rect 415 8604 451 8607
rect 381 8596 397 8598
rect 155 8584 170 8588
rect 73 8582 170 8584
rect 198 8582 366 8594
rect 382 8584 397 8588
rect 415 8585 454 8604
rect 473 8598 480 8599
rect 479 8591 480 8598
rect 463 8588 464 8591
rect 479 8588 492 8591
rect 415 8584 445 8585
rect 454 8584 460 8585
rect 463 8584 492 8588
rect 382 8583 492 8584
rect 382 8582 498 8583
rect 57 8574 108 8582
rect 57 8562 82 8574
rect 89 8562 108 8574
rect 139 8574 189 8582
rect 139 8566 155 8574
rect 162 8572 189 8574
rect 198 8572 419 8582
rect 162 8562 419 8572
rect 448 8574 498 8582
rect 448 8565 464 8574
rect 57 8554 108 8562
rect 155 8554 419 8562
rect 445 8562 464 8565
rect 471 8562 498 8574
rect 445 8554 498 8562
rect 73 8546 74 8554
rect 89 8546 102 8554
rect 73 8538 89 8546
rect 70 8531 89 8534
rect 70 8522 92 8531
rect 43 8512 92 8522
rect 43 8506 73 8512
rect 92 8507 97 8512
rect 15 8490 89 8506
rect 107 8498 137 8554
rect 172 8544 380 8554
rect 415 8550 460 8554
rect 463 8553 464 8554
rect 479 8553 492 8554
rect 198 8514 387 8544
rect 213 8511 387 8514
rect 206 8508 387 8511
rect 15 8488 28 8490
rect 43 8488 77 8490
rect 15 8472 89 8488
rect 116 8484 129 8498
rect 144 8484 160 8500
rect 206 8495 217 8508
rect -1 8450 0 8466
rect 15 8450 28 8472
rect 43 8450 73 8472
rect 116 8468 178 8484
rect 206 8477 217 8493
rect 222 8488 232 8508
rect 242 8488 256 8508
rect 259 8495 268 8508
rect 284 8495 293 8508
rect 222 8477 256 8488
rect 259 8477 268 8493
rect 284 8477 293 8493
rect 300 8488 310 8508
rect 320 8488 334 8508
rect 335 8495 346 8508
rect 300 8477 334 8488
rect 335 8477 346 8493
rect 392 8484 408 8500
rect 415 8498 445 8550
rect 479 8546 480 8553
rect 464 8538 480 8546
rect 451 8506 464 8525
rect 479 8506 509 8522
rect 451 8490 525 8506
rect 451 8488 464 8490
rect 479 8488 513 8490
rect 116 8466 129 8468
rect 144 8466 178 8468
rect 116 8450 178 8466
rect 222 8461 238 8464
rect 300 8461 330 8472
rect 378 8468 424 8484
rect 451 8472 525 8488
rect 378 8466 412 8468
rect 377 8450 424 8466
rect 451 8450 464 8472
rect 479 8450 509 8472
rect 536 8450 537 8466
rect 552 8450 565 8610
rect 595 8506 608 8610
rect 653 8588 654 8598
rect 669 8588 682 8598
rect 653 8584 682 8588
rect 687 8584 717 8610
rect 735 8596 751 8598
rect 823 8596 876 8610
rect 824 8594 888 8596
rect 931 8594 946 8610
rect 995 8607 1025 8610
rect 995 8604 1031 8607
rect 961 8596 977 8598
rect 735 8584 750 8588
rect 653 8582 750 8584
rect 778 8582 946 8594
rect 962 8584 977 8588
rect 995 8585 1034 8604
rect 1053 8598 1060 8599
rect 1059 8591 1060 8598
rect 1043 8588 1044 8591
rect 1059 8588 1072 8591
rect 995 8584 1025 8585
rect 1034 8584 1040 8585
rect 1043 8584 1072 8588
rect 962 8583 1072 8584
rect 962 8582 1078 8583
rect 637 8574 688 8582
rect 637 8562 662 8574
rect 669 8562 688 8574
rect 719 8574 769 8582
rect 719 8566 735 8574
rect 742 8572 769 8574
rect 778 8572 999 8582
rect 742 8562 999 8572
rect 1028 8574 1078 8582
rect 1028 8565 1044 8574
rect 637 8554 688 8562
rect 735 8554 999 8562
rect 1025 8562 1044 8565
rect 1051 8562 1078 8574
rect 1025 8554 1078 8562
rect 653 8546 654 8554
rect 669 8546 682 8554
rect 653 8538 669 8546
rect 650 8531 669 8534
rect 650 8522 672 8531
rect 623 8512 672 8522
rect 623 8506 653 8512
rect 672 8507 677 8512
rect 595 8490 669 8506
rect 687 8498 717 8554
rect 752 8544 960 8554
rect 995 8550 1040 8554
rect 1043 8553 1044 8554
rect 1059 8553 1072 8554
rect 778 8514 967 8544
rect 793 8511 967 8514
rect 786 8508 967 8511
rect 595 8488 608 8490
rect 623 8488 657 8490
rect 595 8472 669 8488
rect 696 8484 709 8498
rect 724 8484 740 8500
rect 786 8495 797 8508
rect 579 8450 580 8466
rect 595 8450 608 8472
rect 623 8450 653 8472
rect 696 8468 758 8484
rect 786 8477 797 8493
rect 802 8488 812 8508
rect 822 8488 836 8508
rect 839 8495 848 8508
rect 864 8495 873 8508
rect 802 8477 836 8488
rect 839 8477 848 8493
rect 864 8477 873 8493
rect 880 8488 890 8508
rect 900 8488 914 8508
rect 915 8495 926 8508
rect 880 8477 914 8488
rect 915 8477 926 8493
rect 972 8484 988 8500
rect 995 8498 1025 8550
rect 1059 8546 1060 8553
rect 1044 8538 1060 8546
rect 1031 8506 1044 8525
rect 1059 8506 1089 8522
rect 1031 8490 1105 8506
rect 1031 8488 1044 8490
rect 1059 8488 1093 8490
rect 696 8466 709 8468
rect 724 8466 758 8468
rect 696 8450 758 8466
rect 802 8461 818 8464
rect 880 8461 910 8472
rect 958 8468 1004 8484
rect 1031 8472 1105 8488
rect 958 8466 992 8468
rect 957 8450 1004 8466
rect 1031 8450 1044 8472
rect 1059 8450 1089 8472
rect 1116 8450 1117 8466
rect 1132 8450 1145 8610
rect 1175 8506 1188 8610
rect 1233 8588 1234 8598
rect 1249 8588 1262 8598
rect 1233 8584 1262 8588
rect 1267 8584 1297 8610
rect 1315 8596 1331 8598
rect 1403 8596 1456 8610
rect 1404 8594 1468 8596
rect 1511 8594 1526 8610
rect 1575 8607 1605 8610
rect 1575 8604 1611 8607
rect 1541 8596 1557 8598
rect 1315 8584 1330 8588
rect 1233 8582 1330 8584
rect 1358 8582 1526 8594
rect 1542 8584 1557 8588
rect 1575 8585 1614 8604
rect 1633 8598 1640 8599
rect 1639 8591 1640 8598
rect 1623 8588 1624 8591
rect 1639 8588 1652 8591
rect 1575 8584 1605 8585
rect 1614 8584 1620 8585
rect 1623 8584 1652 8588
rect 1542 8583 1652 8584
rect 1542 8582 1658 8583
rect 1217 8574 1268 8582
rect 1217 8562 1242 8574
rect 1249 8562 1268 8574
rect 1299 8574 1349 8582
rect 1299 8566 1315 8574
rect 1322 8572 1349 8574
rect 1358 8572 1579 8582
rect 1322 8562 1579 8572
rect 1608 8574 1658 8582
rect 1608 8565 1624 8574
rect 1217 8554 1268 8562
rect 1315 8554 1579 8562
rect 1605 8562 1624 8565
rect 1631 8562 1658 8574
rect 1605 8554 1658 8562
rect 1233 8546 1234 8554
rect 1249 8546 1262 8554
rect 1233 8538 1249 8546
rect 1230 8531 1249 8534
rect 1230 8522 1252 8531
rect 1203 8512 1252 8522
rect 1203 8506 1233 8512
rect 1252 8507 1257 8512
rect 1175 8490 1249 8506
rect 1267 8498 1297 8554
rect 1332 8544 1540 8554
rect 1575 8550 1620 8554
rect 1623 8553 1624 8554
rect 1639 8553 1652 8554
rect 1358 8514 1547 8544
rect 1373 8511 1547 8514
rect 1366 8508 1547 8511
rect 1175 8488 1188 8490
rect 1203 8488 1237 8490
rect 1175 8472 1249 8488
rect 1276 8484 1289 8498
rect 1304 8484 1320 8500
rect 1366 8495 1377 8508
rect 1159 8450 1160 8466
rect 1175 8450 1188 8472
rect 1203 8450 1233 8472
rect 1276 8468 1338 8484
rect 1366 8477 1377 8493
rect 1382 8488 1392 8508
rect 1402 8488 1416 8508
rect 1419 8495 1428 8508
rect 1444 8495 1453 8508
rect 1382 8477 1416 8488
rect 1419 8477 1428 8493
rect 1444 8477 1453 8493
rect 1460 8488 1470 8508
rect 1480 8488 1494 8508
rect 1495 8495 1506 8508
rect 1460 8477 1494 8488
rect 1495 8477 1506 8493
rect 1552 8484 1568 8500
rect 1575 8498 1605 8550
rect 1639 8546 1640 8553
rect 1624 8538 1640 8546
rect 1611 8506 1624 8525
rect 1639 8506 1669 8522
rect 1611 8490 1685 8506
rect 1611 8488 1624 8490
rect 1639 8488 1673 8490
rect 1276 8466 1289 8468
rect 1304 8466 1338 8468
rect 1276 8450 1338 8466
rect 1382 8461 1398 8464
rect 1460 8461 1490 8472
rect 1538 8468 1584 8484
rect 1611 8472 1685 8488
rect 1538 8466 1572 8468
rect 1537 8450 1584 8466
rect 1611 8450 1624 8472
rect 1639 8450 1669 8472
rect 1696 8450 1697 8466
rect 1712 8450 1725 8610
rect 1755 8506 1768 8610
rect 1813 8588 1814 8598
rect 1829 8588 1842 8598
rect 1813 8584 1842 8588
rect 1847 8584 1877 8610
rect 1895 8596 1911 8598
rect 1983 8596 2036 8610
rect 1984 8594 2048 8596
rect 2091 8594 2106 8610
rect 2155 8607 2185 8610
rect 2155 8604 2191 8607
rect 2121 8596 2137 8598
rect 1895 8584 1910 8588
rect 1813 8582 1910 8584
rect 1938 8582 2106 8594
rect 2122 8584 2137 8588
rect 2155 8585 2194 8604
rect 2213 8598 2220 8599
rect 2219 8591 2220 8598
rect 2203 8588 2204 8591
rect 2219 8588 2232 8591
rect 2155 8584 2185 8585
rect 2194 8584 2200 8585
rect 2203 8584 2232 8588
rect 2122 8583 2232 8584
rect 2122 8582 2238 8583
rect 1797 8574 1848 8582
rect 1797 8562 1822 8574
rect 1829 8562 1848 8574
rect 1879 8574 1929 8582
rect 1879 8566 1895 8574
rect 1902 8572 1929 8574
rect 1938 8572 2159 8582
rect 1902 8562 2159 8572
rect 2188 8574 2238 8582
rect 2188 8565 2204 8574
rect 1797 8554 1848 8562
rect 1895 8554 2159 8562
rect 2185 8562 2204 8565
rect 2211 8562 2238 8574
rect 2185 8554 2238 8562
rect 1813 8546 1814 8554
rect 1829 8546 1842 8554
rect 1813 8538 1829 8546
rect 1810 8531 1829 8534
rect 1810 8522 1832 8531
rect 1783 8512 1832 8522
rect 1783 8506 1813 8512
rect 1832 8507 1837 8512
rect 1755 8490 1829 8506
rect 1847 8498 1877 8554
rect 1912 8544 2120 8554
rect 2155 8550 2200 8554
rect 2203 8553 2204 8554
rect 2219 8553 2232 8554
rect 1938 8514 2127 8544
rect 1953 8511 2127 8514
rect 1946 8508 2127 8511
rect 1755 8488 1768 8490
rect 1783 8488 1817 8490
rect 1755 8472 1829 8488
rect 1856 8484 1869 8498
rect 1884 8484 1900 8500
rect 1946 8495 1957 8508
rect 1739 8450 1740 8466
rect 1755 8450 1768 8472
rect 1783 8451 1813 8472
rect 1856 8468 1918 8484
rect 1946 8477 1957 8493
rect 1962 8488 1972 8508
rect 1982 8488 1996 8508
rect 1999 8495 2008 8508
rect 2024 8495 2033 8508
rect 1962 8477 1996 8488
rect 1999 8477 2008 8493
rect 2024 8477 2033 8493
rect 2040 8488 2050 8508
rect 2060 8488 2074 8508
rect 2075 8495 2086 8508
rect 2040 8477 2074 8488
rect 2075 8477 2086 8493
rect 2132 8484 2148 8500
rect 2155 8498 2185 8550
rect 2219 8546 2220 8553
rect 2204 8538 2220 8546
rect 2191 8506 2204 8525
rect 2219 8506 2249 8522
rect 2191 8490 2265 8506
rect 2191 8488 2204 8490
rect 2219 8488 2253 8490
rect 1856 8466 1869 8468
rect 1884 8466 1918 8468
rect 1856 8451 1918 8466
rect 1962 8461 1976 8464
rect 2040 8461 2070 8472
rect 2118 8468 2164 8484
rect 2191 8472 2265 8488
rect 2118 8466 2152 8468
rect 2117 8451 2164 8466
rect 1850 8450 1930 8451
rect 1937 8450 1947 8451
rect -7 8442 34 8450
rect -7 8416 8 8442
rect 15 8416 34 8442
rect 98 8438 160 8450
rect 172 8438 247 8450
rect 305 8438 380 8450
rect 392 8438 423 8450
rect 429 8438 464 8450
rect 98 8436 260 8438
rect -7 8408 34 8416
rect 116 8412 129 8436
rect 144 8434 159 8436
rect -1 8398 0 8408
rect 15 8398 28 8408
rect 43 8398 73 8412
rect 116 8398 159 8412
rect 183 8409 190 8416
rect 193 8412 260 8436
rect 292 8436 464 8438
rect 262 8414 290 8418
rect 292 8414 372 8436
rect 393 8434 408 8436
rect 262 8412 372 8414
rect 193 8408 372 8412
rect 166 8398 196 8408
rect 198 8398 351 8408
rect 359 8398 389 8408
rect 393 8398 423 8412
rect 451 8398 464 8436
rect 536 8442 571 8450
rect 536 8416 537 8442
rect 544 8416 571 8442
rect 479 8398 509 8412
rect 536 8408 571 8416
rect 573 8442 614 8450
rect 573 8416 588 8442
rect 595 8416 614 8442
rect 678 8438 740 8450
rect 752 8438 827 8450
rect 885 8438 960 8450
rect 972 8438 1003 8450
rect 1009 8438 1044 8450
rect 678 8436 840 8438
rect 573 8408 614 8416
rect 696 8412 709 8436
rect 724 8434 739 8436
rect 536 8398 537 8408
rect 552 8398 565 8408
rect 579 8398 580 8408
rect 595 8398 608 8408
rect 623 8398 653 8412
rect 696 8398 739 8412
rect 763 8409 770 8416
rect 773 8412 840 8436
rect 872 8436 1044 8438
rect 842 8414 870 8418
rect 872 8414 952 8436
rect 973 8434 988 8436
rect 842 8412 952 8414
rect 773 8408 952 8412
rect 746 8398 776 8408
rect 778 8398 931 8408
rect 939 8398 969 8408
rect 973 8398 1003 8412
rect 1031 8398 1044 8436
rect 1116 8442 1151 8450
rect 1116 8416 1117 8442
rect 1124 8416 1151 8442
rect 1059 8398 1089 8412
rect 1116 8408 1151 8416
rect 1153 8442 1194 8450
rect 1153 8416 1168 8442
rect 1175 8416 1194 8442
rect 1258 8438 1320 8450
rect 1332 8438 1407 8450
rect 1465 8438 1540 8450
rect 1552 8438 1583 8450
rect 1589 8438 1624 8450
rect 1258 8436 1420 8438
rect 1153 8408 1194 8416
rect 1276 8412 1289 8436
rect 1304 8434 1319 8436
rect 1116 8398 1117 8408
rect 1132 8398 1145 8408
rect 1159 8398 1160 8408
rect 1175 8398 1188 8408
rect 1203 8398 1233 8412
rect 1276 8398 1319 8412
rect 1343 8409 1350 8416
rect 1353 8412 1420 8436
rect 1452 8436 1624 8438
rect 1422 8414 1450 8418
rect 1452 8414 1532 8436
rect 1553 8434 1568 8436
rect 1422 8412 1532 8414
rect 1353 8408 1532 8412
rect 1326 8398 1356 8408
rect 1358 8398 1511 8408
rect 1519 8398 1549 8408
rect 1553 8398 1583 8412
rect 1611 8398 1624 8436
rect 1696 8442 1731 8450
rect 1696 8416 1697 8442
rect 1704 8416 1731 8442
rect 1639 8398 1669 8412
rect 1696 8408 1731 8416
rect 1733 8442 1774 8450
rect 1733 8416 1748 8442
rect 1755 8416 1774 8442
rect 1838 8438 1869 8450
rect 1884 8438 1987 8450
rect 1999 8440 2025 8451
rect 2102 8450 2164 8451
rect 2176 8450 2182 8451
rect 2191 8450 2204 8472
rect 2219 8451 2249 8472
rect 2276 8451 2277 8466
rect 2292 8451 2305 8610
rect 2335 8506 2348 8610
rect 2393 8588 2394 8598
rect 2409 8588 2422 8598
rect 2393 8584 2422 8588
rect 2427 8584 2457 8610
rect 2475 8596 2491 8598
rect 2563 8596 2616 8610
rect 2564 8594 2628 8596
rect 2671 8594 2686 8610
rect 2735 8607 2765 8610
rect 2735 8604 2771 8607
rect 2701 8596 2717 8598
rect 2475 8584 2490 8588
rect 2393 8582 2490 8584
rect 2518 8582 2686 8594
rect 2702 8584 2717 8588
rect 2735 8585 2774 8604
rect 2793 8598 2800 8599
rect 2799 8591 2800 8598
rect 2783 8588 2784 8591
rect 2799 8588 2812 8591
rect 2735 8584 2765 8585
rect 2774 8584 2780 8585
rect 2783 8584 2812 8588
rect 2702 8583 2812 8584
rect 2702 8582 2818 8583
rect 2377 8574 2428 8582
rect 2377 8562 2402 8574
rect 2409 8562 2428 8574
rect 2459 8574 2509 8582
rect 2459 8566 2475 8574
rect 2482 8572 2509 8574
rect 2518 8572 2739 8582
rect 2482 8562 2739 8572
rect 2768 8574 2818 8582
rect 2768 8565 2784 8574
rect 2377 8554 2428 8562
rect 2475 8554 2739 8562
rect 2765 8562 2784 8565
rect 2791 8562 2818 8574
rect 2765 8554 2818 8562
rect 2393 8546 2394 8554
rect 2409 8546 2422 8554
rect 2393 8538 2409 8546
rect 2390 8531 2409 8534
rect 2390 8522 2412 8531
rect 2363 8512 2412 8522
rect 2363 8506 2393 8512
rect 2412 8507 2417 8512
rect 2335 8490 2409 8506
rect 2427 8498 2457 8554
rect 2492 8544 2700 8554
rect 2735 8550 2780 8554
rect 2783 8553 2784 8554
rect 2799 8553 2812 8554
rect 2518 8514 2707 8544
rect 2533 8511 2707 8514
rect 2526 8508 2707 8511
rect 2335 8488 2348 8490
rect 2363 8488 2397 8490
rect 2335 8472 2409 8488
rect 2436 8484 2449 8498
rect 2464 8484 2480 8500
rect 2526 8495 2537 8508
rect 2045 8440 2148 8450
rect 1999 8438 2148 8440
rect 2169 8438 2204 8450
rect 1838 8436 2000 8438
rect 1850 8416 1869 8436
rect 1884 8434 1914 8436
rect 1733 8408 1774 8416
rect 1856 8412 1869 8416
rect 1921 8420 2000 8436
rect 2032 8436 2204 8438
rect 2032 8420 2111 8436
rect 2118 8434 2148 8436
rect 1696 8398 1697 8408
rect 1712 8398 1725 8408
rect 1739 8398 1740 8408
rect 1755 8398 1768 8408
rect 1783 8398 1813 8412
rect 1856 8398 1899 8412
rect 1921 8408 2111 8420
rect 2176 8416 2182 8436
rect 1906 8398 1936 8408
rect 1937 8398 2095 8408
rect 2099 8398 2129 8408
rect 2133 8398 2163 8412
rect 2191 8398 2204 8436
rect 2276 8450 2305 8451
rect 2319 8451 2320 8466
rect 2335 8451 2348 8472
rect 2363 8451 2393 8472
rect 2436 8468 2498 8484
rect 2526 8477 2537 8493
rect 2542 8488 2552 8508
rect 2562 8488 2576 8508
rect 2579 8495 2588 8508
rect 2604 8495 2613 8508
rect 2542 8477 2576 8488
rect 2579 8477 2588 8493
rect 2604 8477 2613 8493
rect 2620 8488 2630 8508
rect 2640 8488 2654 8508
rect 2655 8495 2666 8508
rect 2620 8477 2654 8488
rect 2655 8477 2666 8493
rect 2712 8484 2728 8500
rect 2735 8498 2765 8550
rect 2799 8546 2800 8553
rect 2784 8538 2800 8546
rect 2771 8506 2784 8525
rect 2799 8506 2829 8522
rect 2771 8490 2845 8506
rect 2771 8488 2784 8490
rect 2799 8488 2833 8490
rect 2436 8466 2449 8468
rect 2464 8466 2498 8468
rect 2436 8451 2498 8466
rect 2542 8461 2558 8464
rect 2620 8461 2650 8472
rect 2698 8468 2744 8484
rect 2771 8472 2845 8488
rect 2698 8466 2732 8468
rect 2697 8451 2744 8466
rect 2319 8450 2348 8451
rect 2430 8450 2510 8451
rect 2517 8450 2527 8451
rect 2276 8442 2311 8450
rect 2276 8416 2277 8442
rect 2284 8416 2311 8442
rect 2219 8398 2249 8412
rect 2276 8408 2311 8416
rect 2313 8442 2354 8450
rect 2313 8416 2328 8442
rect 2335 8416 2354 8442
rect 2418 8438 2449 8450
rect 2464 8438 2567 8450
rect 2579 8440 2605 8451
rect 2682 8450 2744 8451
rect 2756 8450 2762 8451
rect 2771 8450 2784 8472
rect 2799 8451 2829 8472
rect 2856 8451 2857 8466
rect 2872 8451 2885 8610
rect 2915 8506 2928 8610
rect 2973 8588 2974 8598
rect 2989 8588 3002 8598
rect 2973 8584 3002 8588
rect 3007 8584 3037 8610
rect 3055 8596 3071 8598
rect 3143 8596 3196 8610
rect 3144 8594 3208 8596
rect 3251 8594 3266 8610
rect 3315 8607 3345 8610
rect 3315 8604 3351 8607
rect 3281 8596 3297 8598
rect 3055 8584 3070 8588
rect 2973 8582 3070 8584
rect 3098 8582 3266 8594
rect 3282 8584 3297 8588
rect 3315 8585 3354 8604
rect 3373 8598 3380 8599
rect 3379 8591 3380 8598
rect 3363 8588 3364 8591
rect 3379 8588 3392 8591
rect 3315 8584 3345 8585
rect 3354 8584 3360 8585
rect 3363 8584 3392 8588
rect 3282 8583 3392 8584
rect 3282 8582 3398 8583
rect 2957 8574 3008 8582
rect 2957 8562 2982 8574
rect 2989 8562 3008 8574
rect 3039 8574 3089 8582
rect 3039 8566 3055 8574
rect 3062 8572 3089 8574
rect 3098 8572 3319 8582
rect 3062 8562 3319 8572
rect 3348 8574 3398 8582
rect 3348 8565 3364 8574
rect 2957 8554 3008 8562
rect 3055 8554 3319 8562
rect 3345 8562 3364 8565
rect 3371 8562 3398 8574
rect 3345 8554 3398 8562
rect 2973 8546 2974 8554
rect 2989 8546 3002 8554
rect 2973 8538 2989 8546
rect 2970 8531 2989 8534
rect 2970 8522 2992 8531
rect 2943 8512 2992 8522
rect 2943 8506 2973 8512
rect 2992 8507 2997 8512
rect 2915 8490 2989 8506
rect 3007 8498 3037 8554
rect 3072 8544 3280 8554
rect 3315 8550 3360 8554
rect 3363 8553 3364 8554
rect 3379 8553 3392 8554
rect 3098 8514 3287 8544
rect 3113 8511 3287 8514
rect 3106 8508 3287 8511
rect 2915 8488 2928 8490
rect 2943 8488 2977 8490
rect 2915 8472 2989 8488
rect 3016 8484 3029 8498
rect 3044 8484 3060 8500
rect 3106 8495 3117 8508
rect 2625 8440 2728 8450
rect 2579 8438 2728 8440
rect 2749 8438 2784 8450
rect 2418 8436 2580 8438
rect 2430 8416 2449 8436
rect 2464 8434 2494 8436
rect 2313 8408 2354 8416
rect 2436 8412 2449 8416
rect 2501 8420 2580 8436
rect 2612 8436 2784 8438
rect 2612 8420 2691 8436
rect 2698 8434 2728 8436
rect 2276 8398 2305 8408
rect 2319 8398 2348 8408
rect 2363 8398 2393 8412
rect 2436 8398 2479 8412
rect 2501 8408 2691 8420
rect 2756 8416 2762 8436
rect 2486 8398 2516 8408
rect 2517 8398 2675 8408
rect 2679 8398 2709 8408
rect 2713 8398 2743 8412
rect 2771 8398 2784 8436
rect 2856 8450 2885 8451
rect 2899 8451 2900 8466
rect 2915 8451 2928 8472
rect 2943 8451 2973 8472
rect 3016 8468 3078 8484
rect 3106 8477 3117 8493
rect 3122 8488 3132 8508
rect 3142 8488 3156 8508
rect 3159 8495 3168 8508
rect 3184 8495 3193 8508
rect 3122 8477 3156 8488
rect 3159 8477 3168 8493
rect 3184 8477 3193 8493
rect 3200 8488 3210 8508
rect 3220 8488 3234 8508
rect 3235 8495 3246 8508
rect 3200 8477 3234 8488
rect 3235 8477 3246 8493
rect 3292 8484 3308 8500
rect 3315 8498 3345 8550
rect 3379 8546 3380 8553
rect 3364 8538 3380 8546
rect 3351 8506 3364 8525
rect 3379 8506 3409 8522
rect 3351 8490 3425 8506
rect 3351 8488 3364 8490
rect 3379 8488 3413 8490
rect 3016 8466 3029 8468
rect 3044 8466 3078 8468
rect 3016 8451 3078 8466
rect 3122 8461 3138 8464
rect 3200 8461 3230 8472
rect 3278 8468 3324 8484
rect 3351 8472 3425 8488
rect 3278 8466 3312 8468
rect 3277 8451 3324 8466
rect 2899 8450 2928 8451
rect 3010 8450 3090 8451
rect 3097 8450 3107 8451
rect 2856 8442 2891 8450
rect 2856 8416 2857 8442
rect 2864 8416 2891 8442
rect 2799 8398 2829 8412
rect 2856 8408 2891 8416
rect 2893 8442 2934 8450
rect 2893 8416 2908 8442
rect 2915 8416 2934 8442
rect 2998 8438 3029 8450
rect 3044 8438 3147 8450
rect 3159 8440 3185 8451
rect 3262 8450 3324 8451
rect 3336 8450 3342 8451
rect 3351 8450 3364 8472
rect 3379 8451 3409 8472
rect 3436 8451 3437 8466
rect 3452 8451 3465 8610
rect 3495 8506 3508 8610
rect 3553 8588 3554 8598
rect 3569 8588 3582 8598
rect 3553 8584 3582 8588
rect 3587 8584 3617 8610
rect 3635 8596 3651 8598
rect 3723 8596 3776 8610
rect 3724 8594 3788 8596
rect 3831 8594 3846 8610
rect 3895 8607 3925 8610
rect 3895 8604 3931 8607
rect 3861 8596 3877 8598
rect 3635 8584 3650 8588
rect 3553 8582 3650 8584
rect 3678 8582 3846 8594
rect 3862 8584 3877 8588
rect 3895 8585 3934 8604
rect 3953 8598 3960 8599
rect 3959 8591 3960 8598
rect 3943 8588 3944 8591
rect 3959 8588 3972 8591
rect 3895 8584 3925 8585
rect 3934 8584 3940 8585
rect 3943 8584 3972 8588
rect 3862 8583 3972 8584
rect 3862 8582 3978 8583
rect 3537 8574 3588 8582
rect 3537 8562 3562 8574
rect 3569 8562 3588 8574
rect 3619 8574 3669 8582
rect 3619 8566 3635 8574
rect 3642 8572 3669 8574
rect 3678 8572 3899 8582
rect 3642 8562 3899 8572
rect 3928 8574 3978 8582
rect 3928 8565 3944 8574
rect 3537 8554 3588 8562
rect 3635 8554 3899 8562
rect 3925 8562 3944 8565
rect 3951 8562 3978 8574
rect 3925 8554 3978 8562
rect 3553 8546 3554 8554
rect 3569 8546 3582 8554
rect 3553 8538 3569 8546
rect 3550 8531 3569 8534
rect 3550 8522 3572 8531
rect 3523 8512 3572 8522
rect 3523 8506 3553 8512
rect 3572 8507 3577 8512
rect 3495 8490 3569 8506
rect 3587 8498 3617 8554
rect 3652 8544 3860 8554
rect 3895 8550 3940 8554
rect 3943 8553 3944 8554
rect 3959 8553 3972 8554
rect 3678 8514 3867 8544
rect 3693 8511 3867 8514
rect 3686 8508 3867 8511
rect 3495 8488 3508 8490
rect 3523 8488 3557 8490
rect 3495 8472 3569 8488
rect 3596 8484 3609 8498
rect 3624 8484 3640 8500
rect 3686 8495 3697 8508
rect 3205 8440 3308 8450
rect 3159 8438 3308 8440
rect 3329 8438 3364 8450
rect 2998 8436 3160 8438
rect 3010 8416 3029 8436
rect 3044 8434 3074 8436
rect 2893 8408 2934 8416
rect 3016 8412 3029 8416
rect 3081 8420 3160 8436
rect 3192 8436 3364 8438
rect 3192 8420 3271 8436
rect 3278 8434 3308 8436
rect 2856 8398 2885 8408
rect 2899 8398 2928 8408
rect 2943 8398 2973 8412
rect 3016 8398 3059 8412
rect 3081 8408 3271 8420
rect 3336 8416 3342 8436
rect 3066 8398 3096 8408
rect 3097 8398 3255 8408
rect 3259 8398 3289 8408
rect 3293 8398 3323 8412
rect 3351 8398 3364 8436
rect 3436 8450 3465 8451
rect 3479 8451 3480 8466
rect 3495 8451 3508 8472
rect 3523 8451 3553 8472
rect 3596 8468 3658 8484
rect 3686 8477 3697 8493
rect 3702 8488 3712 8508
rect 3722 8488 3736 8508
rect 3739 8495 3748 8508
rect 3764 8495 3773 8508
rect 3702 8477 3736 8488
rect 3739 8477 3748 8493
rect 3764 8477 3773 8493
rect 3780 8488 3790 8508
rect 3800 8488 3814 8508
rect 3815 8495 3826 8508
rect 3780 8477 3814 8488
rect 3815 8477 3826 8493
rect 3872 8484 3888 8500
rect 3895 8498 3925 8550
rect 3959 8546 3960 8553
rect 3944 8538 3960 8546
rect 3931 8506 3944 8525
rect 3959 8506 3989 8522
rect 3931 8490 4005 8506
rect 3931 8488 3944 8490
rect 3959 8488 3993 8490
rect 3596 8466 3609 8468
rect 3624 8466 3658 8468
rect 3596 8451 3658 8466
rect 3702 8461 3718 8464
rect 3780 8461 3810 8472
rect 3858 8468 3904 8484
rect 3931 8472 4005 8488
rect 3858 8466 3892 8468
rect 3857 8451 3904 8466
rect 3479 8450 3508 8451
rect 3590 8450 3670 8451
rect 3677 8450 3687 8451
rect 3436 8442 3471 8450
rect 3436 8416 3437 8442
rect 3444 8416 3471 8442
rect 3379 8398 3409 8412
rect 3436 8408 3471 8416
rect 3473 8442 3514 8450
rect 3473 8416 3488 8442
rect 3495 8416 3514 8442
rect 3578 8438 3609 8450
rect 3624 8438 3727 8450
rect 3739 8440 3765 8451
rect 3842 8450 3904 8451
rect 3916 8450 3922 8451
rect 3931 8450 3944 8472
rect 3959 8451 3989 8472
rect 4016 8451 4017 8466
rect 4032 8451 4045 8610
rect 4075 8506 4088 8610
rect 4133 8588 4134 8598
rect 4149 8588 4162 8598
rect 4133 8584 4162 8588
rect 4167 8584 4197 8610
rect 4215 8596 4231 8598
rect 4303 8596 4356 8610
rect 4304 8594 4368 8596
rect 4411 8594 4426 8610
rect 4475 8607 4505 8610
rect 4475 8604 4511 8607
rect 4441 8596 4457 8598
rect 4215 8584 4230 8588
rect 4133 8582 4230 8584
rect 4258 8582 4426 8594
rect 4442 8584 4457 8588
rect 4475 8585 4514 8604
rect 4533 8598 4540 8599
rect 4539 8591 4540 8598
rect 4523 8588 4524 8591
rect 4539 8588 4552 8591
rect 4475 8584 4505 8585
rect 4514 8584 4520 8585
rect 4523 8584 4552 8588
rect 4442 8583 4552 8584
rect 4442 8582 4558 8583
rect 4117 8574 4168 8582
rect 4117 8562 4142 8574
rect 4149 8562 4168 8574
rect 4199 8574 4249 8582
rect 4199 8566 4215 8574
rect 4222 8572 4249 8574
rect 4258 8572 4479 8582
rect 4222 8562 4479 8572
rect 4508 8574 4558 8582
rect 4508 8565 4524 8574
rect 4117 8554 4168 8562
rect 4215 8554 4479 8562
rect 4505 8562 4524 8565
rect 4531 8562 4558 8574
rect 4505 8554 4558 8562
rect 4133 8546 4134 8554
rect 4149 8546 4162 8554
rect 4133 8538 4149 8546
rect 4130 8531 4149 8534
rect 4130 8522 4152 8531
rect 4103 8512 4152 8522
rect 4103 8506 4133 8512
rect 4152 8507 4157 8512
rect 4075 8490 4149 8506
rect 4167 8498 4197 8554
rect 4232 8544 4440 8554
rect 4475 8550 4520 8554
rect 4523 8553 4524 8554
rect 4539 8553 4552 8554
rect 4258 8514 4447 8544
rect 4273 8511 4447 8514
rect 4266 8508 4447 8511
rect 4075 8488 4088 8490
rect 4103 8488 4137 8490
rect 4075 8472 4149 8488
rect 4176 8484 4189 8498
rect 4204 8484 4220 8500
rect 4266 8495 4277 8508
rect 3785 8440 3888 8450
rect 3739 8438 3888 8440
rect 3909 8438 3944 8450
rect 3578 8436 3740 8438
rect 3590 8416 3609 8436
rect 3624 8434 3654 8436
rect 3473 8408 3514 8416
rect 3596 8412 3609 8416
rect 3661 8420 3740 8436
rect 3772 8436 3944 8438
rect 3772 8420 3851 8436
rect 3858 8434 3888 8436
rect 3436 8398 3465 8408
rect 3479 8398 3508 8408
rect 3523 8398 3553 8412
rect 3596 8398 3639 8412
rect 3661 8408 3851 8420
rect 3916 8416 3922 8436
rect 3646 8398 3676 8408
rect 3677 8398 3835 8408
rect 3839 8398 3869 8408
rect 3873 8398 3903 8412
rect 3931 8398 3944 8436
rect 4016 8450 4045 8451
rect 4059 8451 4060 8466
rect 4075 8451 4088 8472
rect 4103 8451 4133 8472
rect 4176 8468 4238 8484
rect 4266 8477 4277 8493
rect 4282 8488 4292 8508
rect 4302 8488 4316 8508
rect 4319 8495 4328 8508
rect 4344 8495 4353 8508
rect 4282 8477 4316 8488
rect 4319 8477 4328 8493
rect 4344 8477 4353 8493
rect 4360 8488 4370 8508
rect 4380 8488 4394 8508
rect 4395 8495 4406 8508
rect 4360 8477 4394 8488
rect 4395 8477 4406 8493
rect 4452 8484 4468 8500
rect 4475 8498 4505 8550
rect 4539 8546 4540 8553
rect 4524 8538 4540 8546
rect 4511 8506 4524 8525
rect 4539 8506 4569 8522
rect 4511 8490 4585 8506
rect 4511 8488 4524 8490
rect 4539 8488 4573 8490
rect 4176 8466 4189 8468
rect 4204 8466 4238 8468
rect 4176 8451 4238 8466
rect 4282 8461 4298 8464
rect 4360 8461 4390 8472
rect 4438 8468 4484 8484
rect 4511 8472 4585 8488
rect 4438 8466 4472 8468
rect 4437 8451 4484 8466
rect 4059 8450 4088 8451
rect 4170 8450 4250 8451
rect 4257 8450 4267 8451
rect 4016 8442 4051 8450
rect 4016 8416 4017 8442
rect 4024 8416 4051 8442
rect 3959 8398 3989 8412
rect 4016 8408 4051 8416
rect 4053 8442 4094 8450
rect 4053 8416 4068 8442
rect 4075 8416 4094 8442
rect 4158 8438 4189 8450
rect 4204 8438 4307 8450
rect 4319 8440 4345 8451
rect 4422 8450 4484 8451
rect 4496 8450 4502 8451
rect 4511 8450 4524 8472
rect 4539 8451 4569 8472
rect 4596 8451 4597 8466
rect 4612 8451 4625 8610
rect 4655 8506 4668 8610
rect 4713 8588 4714 8598
rect 4729 8588 4742 8598
rect 4713 8584 4742 8588
rect 4747 8584 4777 8610
rect 4795 8596 4811 8598
rect 4883 8596 4936 8610
rect 4884 8594 4948 8596
rect 4991 8594 5006 8610
rect 5055 8607 5085 8610
rect 5055 8604 5091 8607
rect 5021 8596 5037 8598
rect 4795 8584 4810 8588
rect 4713 8582 4810 8584
rect 4838 8582 5006 8594
rect 5022 8584 5037 8588
rect 5055 8585 5094 8604
rect 5113 8598 5120 8599
rect 5119 8591 5120 8598
rect 5103 8588 5104 8591
rect 5119 8588 5132 8591
rect 5055 8584 5085 8585
rect 5094 8584 5100 8585
rect 5103 8584 5132 8588
rect 5022 8583 5132 8584
rect 5022 8582 5138 8583
rect 4697 8574 4748 8582
rect 4697 8562 4722 8574
rect 4729 8562 4748 8574
rect 4779 8574 4829 8582
rect 4779 8566 4795 8574
rect 4802 8572 4829 8574
rect 4838 8572 5059 8582
rect 4802 8562 5059 8572
rect 5088 8574 5138 8582
rect 5088 8565 5104 8574
rect 4697 8554 4748 8562
rect 4795 8554 5059 8562
rect 5085 8562 5104 8565
rect 5111 8562 5138 8574
rect 5085 8554 5138 8562
rect 4713 8546 4714 8554
rect 4729 8546 4742 8554
rect 4713 8538 4729 8546
rect 4710 8531 4729 8534
rect 4710 8522 4732 8531
rect 4683 8512 4732 8522
rect 4683 8506 4713 8512
rect 4732 8507 4737 8512
rect 4655 8490 4729 8506
rect 4747 8498 4777 8554
rect 4812 8544 5020 8554
rect 5055 8550 5100 8554
rect 5103 8553 5104 8554
rect 5119 8553 5132 8554
rect 4838 8514 5027 8544
rect 4853 8511 5027 8514
rect 4846 8508 5027 8511
rect 4655 8488 4668 8490
rect 4683 8488 4717 8490
rect 4655 8472 4729 8488
rect 4756 8484 4769 8498
rect 4784 8484 4800 8500
rect 4846 8495 4857 8508
rect 4365 8440 4468 8450
rect 4319 8438 4468 8440
rect 4489 8438 4524 8450
rect 4158 8436 4320 8438
rect 4170 8416 4189 8436
rect 4204 8434 4234 8436
rect 4053 8408 4094 8416
rect 4176 8412 4189 8416
rect 4241 8420 4320 8436
rect 4352 8436 4524 8438
rect 4352 8420 4431 8436
rect 4438 8434 4468 8436
rect 4016 8398 4045 8408
rect 4059 8398 4088 8408
rect 4103 8398 4133 8412
rect 4176 8398 4219 8412
rect 4241 8408 4431 8420
rect 4496 8416 4502 8436
rect 4226 8398 4256 8408
rect 4257 8398 4415 8408
rect 4419 8398 4449 8408
rect 4453 8398 4483 8412
rect 4511 8398 4524 8436
rect 4596 8450 4625 8451
rect 4639 8451 4640 8466
rect 4655 8451 4668 8472
rect 4683 8451 4713 8472
rect 4756 8468 4818 8484
rect 4846 8477 4857 8493
rect 4862 8488 4872 8508
rect 4882 8488 4896 8508
rect 4899 8495 4908 8508
rect 4924 8495 4933 8508
rect 4862 8477 4896 8488
rect 4899 8477 4908 8493
rect 4924 8477 4933 8493
rect 4940 8488 4950 8508
rect 4960 8488 4974 8508
rect 4975 8495 4986 8508
rect 4940 8477 4974 8488
rect 4975 8477 4986 8493
rect 5032 8484 5048 8500
rect 5055 8498 5085 8550
rect 5119 8546 5120 8553
rect 5104 8538 5120 8546
rect 5091 8506 5104 8525
rect 5119 8506 5149 8522
rect 5091 8490 5165 8506
rect 5091 8488 5104 8490
rect 5119 8488 5153 8490
rect 4756 8466 4769 8468
rect 4784 8466 4818 8468
rect 4756 8451 4818 8466
rect 4862 8461 4878 8464
rect 4940 8461 4970 8472
rect 5018 8468 5064 8484
rect 5091 8472 5165 8488
rect 5018 8466 5052 8468
rect 5017 8451 5064 8466
rect 4639 8450 4668 8451
rect 4750 8450 4830 8451
rect 4837 8450 4847 8451
rect 4596 8442 4631 8450
rect 4596 8416 4597 8442
rect 4604 8416 4631 8442
rect 4539 8398 4569 8412
rect 4596 8408 4631 8416
rect 4633 8442 4674 8450
rect 4633 8416 4648 8442
rect 4655 8416 4674 8442
rect 4738 8438 4769 8450
rect 4784 8438 4887 8450
rect 4899 8440 4925 8451
rect 5002 8450 5064 8451
rect 5076 8450 5082 8451
rect 5091 8450 5104 8472
rect 5119 8451 5149 8472
rect 5176 8451 5177 8466
rect 5192 8451 5205 8610
rect 5235 8506 5248 8610
rect 5293 8588 5294 8598
rect 5309 8588 5322 8598
rect 5293 8584 5322 8588
rect 5327 8584 5357 8610
rect 5375 8596 5391 8598
rect 5463 8596 5516 8610
rect 5464 8594 5528 8596
rect 5571 8594 5586 8610
rect 5635 8607 5665 8610
rect 5635 8604 5671 8607
rect 5601 8596 5617 8598
rect 5375 8584 5390 8588
rect 5293 8582 5390 8584
rect 5418 8582 5586 8594
rect 5602 8584 5617 8588
rect 5635 8585 5674 8604
rect 5693 8598 5700 8599
rect 5699 8591 5700 8598
rect 5683 8588 5684 8591
rect 5699 8588 5712 8591
rect 5635 8584 5665 8585
rect 5674 8584 5680 8585
rect 5683 8584 5712 8588
rect 5602 8583 5712 8584
rect 5602 8582 5718 8583
rect 5277 8574 5328 8582
rect 5277 8562 5302 8574
rect 5309 8562 5328 8574
rect 5359 8574 5409 8582
rect 5359 8566 5375 8574
rect 5382 8572 5409 8574
rect 5418 8572 5639 8582
rect 5382 8562 5639 8572
rect 5668 8574 5718 8582
rect 5668 8565 5684 8574
rect 5277 8554 5328 8562
rect 5375 8554 5639 8562
rect 5665 8562 5684 8565
rect 5691 8562 5718 8574
rect 5665 8554 5718 8562
rect 5293 8546 5294 8554
rect 5309 8546 5322 8554
rect 5293 8538 5309 8546
rect 5290 8531 5309 8534
rect 5290 8522 5312 8531
rect 5263 8512 5312 8522
rect 5263 8506 5293 8512
rect 5312 8507 5317 8512
rect 5235 8490 5309 8506
rect 5327 8498 5357 8554
rect 5392 8544 5600 8554
rect 5635 8550 5680 8554
rect 5683 8553 5684 8554
rect 5699 8553 5712 8554
rect 5418 8514 5607 8544
rect 5433 8511 5607 8514
rect 5426 8508 5607 8511
rect 5235 8488 5248 8490
rect 5263 8488 5297 8490
rect 5235 8472 5309 8488
rect 5336 8484 5349 8498
rect 5364 8484 5380 8500
rect 5426 8495 5437 8508
rect 4945 8440 5048 8450
rect 4899 8438 5048 8440
rect 5069 8438 5104 8450
rect 4738 8436 4900 8438
rect 4750 8416 4769 8436
rect 4784 8434 4814 8436
rect 4633 8408 4674 8416
rect 4756 8412 4769 8416
rect 4821 8420 4900 8436
rect 4932 8436 5104 8438
rect 4932 8420 5011 8436
rect 5018 8434 5048 8436
rect 4596 8398 4625 8408
rect 4639 8398 4668 8408
rect 4683 8398 4713 8412
rect 4756 8398 4799 8412
rect 4821 8408 5011 8420
rect 5076 8416 5082 8436
rect 4806 8398 4836 8408
rect 4837 8398 4995 8408
rect 4999 8398 5029 8408
rect 5033 8398 5063 8412
rect 5091 8398 5104 8436
rect 5176 8450 5205 8451
rect 5219 8451 5220 8466
rect 5235 8451 5248 8472
rect 5263 8451 5293 8472
rect 5336 8468 5398 8484
rect 5426 8477 5437 8493
rect 5442 8488 5452 8508
rect 5462 8488 5476 8508
rect 5479 8495 5488 8508
rect 5504 8495 5513 8508
rect 5442 8477 5476 8488
rect 5479 8477 5488 8493
rect 5504 8477 5513 8493
rect 5520 8488 5530 8508
rect 5540 8488 5554 8508
rect 5555 8495 5566 8508
rect 5520 8477 5554 8488
rect 5555 8477 5566 8493
rect 5612 8484 5628 8500
rect 5635 8498 5665 8550
rect 5699 8546 5700 8553
rect 5684 8538 5700 8546
rect 5671 8506 5684 8525
rect 5699 8506 5729 8522
rect 5671 8490 5745 8506
rect 5671 8488 5684 8490
rect 5699 8488 5733 8490
rect 5336 8466 5349 8468
rect 5364 8466 5398 8468
rect 5336 8451 5398 8466
rect 5442 8461 5458 8464
rect 5520 8461 5550 8472
rect 5598 8468 5644 8484
rect 5671 8472 5745 8488
rect 5598 8466 5632 8468
rect 5597 8451 5644 8466
rect 5219 8450 5248 8451
rect 5330 8450 5410 8451
rect 5417 8450 5427 8451
rect 5176 8442 5211 8450
rect 5176 8416 5177 8442
rect 5184 8416 5211 8442
rect 5119 8398 5149 8412
rect 5176 8408 5211 8416
rect 5213 8442 5254 8450
rect 5213 8416 5228 8442
rect 5235 8416 5254 8442
rect 5318 8438 5349 8450
rect 5364 8438 5467 8450
rect 5479 8440 5505 8451
rect 5582 8450 5644 8451
rect 5656 8450 5662 8451
rect 5671 8450 5684 8472
rect 5699 8451 5729 8472
rect 5756 8451 5757 8466
rect 5772 8451 5785 8610
rect 5815 8506 5828 8610
rect 5873 8588 5874 8598
rect 5889 8588 5902 8598
rect 5873 8584 5902 8588
rect 5907 8584 5937 8610
rect 5955 8596 5971 8598
rect 6043 8596 6096 8610
rect 6044 8594 6108 8596
rect 6151 8594 6166 8610
rect 6215 8607 6245 8610
rect 6215 8604 6251 8607
rect 6181 8596 6197 8598
rect 5955 8584 5970 8588
rect 5873 8582 5970 8584
rect 5998 8582 6166 8594
rect 6182 8584 6197 8588
rect 6215 8585 6254 8604
rect 6273 8598 6280 8599
rect 6279 8591 6280 8598
rect 6263 8588 6264 8591
rect 6279 8588 6292 8591
rect 6215 8584 6245 8585
rect 6254 8584 6260 8585
rect 6263 8584 6292 8588
rect 6182 8583 6292 8584
rect 6182 8582 6298 8583
rect 5857 8574 5908 8582
rect 5857 8562 5882 8574
rect 5889 8562 5908 8574
rect 5939 8574 5989 8582
rect 5939 8566 5955 8574
rect 5962 8572 5989 8574
rect 5998 8572 6219 8582
rect 5962 8562 6219 8572
rect 6248 8574 6298 8582
rect 6248 8565 6264 8574
rect 5857 8554 5908 8562
rect 5955 8554 6219 8562
rect 6245 8562 6264 8565
rect 6271 8562 6298 8574
rect 6245 8554 6298 8562
rect 5873 8546 5874 8554
rect 5889 8546 5902 8554
rect 5873 8538 5889 8546
rect 5870 8531 5889 8534
rect 5870 8522 5892 8531
rect 5843 8512 5892 8522
rect 5843 8506 5873 8512
rect 5892 8507 5897 8512
rect 5815 8490 5889 8506
rect 5907 8498 5937 8554
rect 5972 8544 6180 8554
rect 6215 8550 6260 8554
rect 6263 8553 6264 8554
rect 6279 8553 6292 8554
rect 5998 8514 6187 8544
rect 6013 8511 6187 8514
rect 6006 8508 6187 8511
rect 5815 8488 5828 8490
rect 5843 8488 5877 8490
rect 5815 8472 5889 8488
rect 5916 8484 5929 8498
rect 5944 8484 5960 8500
rect 6006 8495 6017 8508
rect 5525 8440 5628 8450
rect 5479 8438 5628 8440
rect 5649 8438 5684 8450
rect 5318 8436 5480 8438
rect 5330 8416 5349 8436
rect 5364 8434 5394 8436
rect 5213 8408 5254 8416
rect 5336 8412 5349 8416
rect 5401 8420 5480 8436
rect 5512 8436 5684 8438
rect 5512 8420 5591 8436
rect 5598 8434 5628 8436
rect 5176 8398 5205 8408
rect 5219 8398 5248 8408
rect 5263 8398 5293 8412
rect 5336 8398 5379 8412
rect 5401 8408 5591 8420
rect 5656 8416 5662 8436
rect 5386 8398 5416 8408
rect 5417 8398 5575 8408
rect 5579 8398 5609 8408
rect 5613 8398 5643 8412
rect 5671 8398 5684 8436
rect 5756 8450 5785 8451
rect 5799 8451 5800 8466
rect 5815 8451 5828 8472
rect 5843 8451 5873 8472
rect 5916 8468 5978 8484
rect 6006 8477 6017 8493
rect 6022 8488 6032 8508
rect 6042 8488 6056 8508
rect 6059 8495 6068 8508
rect 6084 8495 6093 8508
rect 6022 8477 6056 8488
rect 6059 8477 6068 8493
rect 6084 8477 6093 8493
rect 6100 8488 6110 8508
rect 6120 8488 6134 8508
rect 6135 8495 6146 8508
rect 6100 8477 6134 8488
rect 6135 8477 6146 8493
rect 6192 8484 6208 8500
rect 6215 8498 6245 8550
rect 6279 8546 6280 8553
rect 6264 8538 6280 8546
rect 6251 8506 6264 8525
rect 6279 8506 6309 8522
rect 6251 8490 6325 8506
rect 6251 8488 6264 8490
rect 6279 8488 6313 8490
rect 5916 8466 5929 8468
rect 5944 8466 5978 8468
rect 5916 8451 5978 8466
rect 6022 8461 6038 8464
rect 6100 8461 6130 8472
rect 6178 8468 6224 8484
rect 6251 8472 6325 8488
rect 6178 8466 6212 8468
rect 6177 8451 6224 8466
rect 5799 8450 5828 8451
rect 5910 8450 5990 8451
rect 5997 8450 6007 8451
rect 5756 8442 5791 8450
rect 5756 8416 5757 8442
rect 5764 8416 5791 8442
rect 5699 8398 5729 8412
rect 5756 8408 5791 8416
rect 5793 8442 5834 8450
rect 5793 8416 5808 8442
rect 5815 8416 5834 8442
rect 5898 8438 5929 8450
rect 5944 8438 6047 8450
rect 6059 8440 6085 8451
rect 6162 8450 6224 8451
rect 6236 8450 6242 8451
rect 6251 8450 6264 8472
rect 6279 8451 6309 8472
rect 6336 8451 6337 8466
rect 6352 8451 6365 8610
rect 6395 8506 6408 8610
rect 6453 8588 6454 8598
rect 6469 8588 6482 8598
rect 6453 8584 6482 8588
rect 6487 8584 6517 8610
rect 6535 8596 6551 8598
rect 6623 8596 6676 8610
rect 6624 8594 6688 8596
rect 6731 8594 6746 8610
rect 6795 8607 6825 8610
rect 6795 8604 6831 8607
rect 6761 8596 6777 8598
rect 6535 8584 6550 8588
rect 6453 8582 6550 8584
rect 6578 8582 6746 8594
rect 6762 8584 6777 8588
rect 6795 8585 6834 8604
rect 6853 8598 6860 8599
rect 6859 8591 6860 8598
rect 6843 8588 6844 8591
rect 6859 8588 6872 8591
rect 6795 8584 6825 8585
rect 6834 8584 6840 8585
rect 6843 8584 6872 8588
rect 6762 8583 6872 8584
rect 6762 8582 6878 8583
rect 6437 8574 6488 8582
rect 6437 8562 6462 8574
rect 6469 8562 6488 8574
rect 6519 8574 6569 8582
rect 6519 8566 6535 8574
rect 6542 8572 6569 8574
rect 6578 8572 6799 8582
rect 6542 8562 6799 8572
rect 6828 8574 6878 8582
rect 6828 8565 6844 8574
rect 6437 8554 6488 8562
rect 6535 8554 6799 8562
rect 6825 8562 6844 8565
rect 6851 8562 6878 8574
rect 6825 8554 6878 8562
rect 6453 8546 6454 8554
rect 6469 8546 6482 8554
rect 6453 8538 6469 8546
rect 6450 8531 6469 8534
rect 6450 8522 6472 8531
rect 6423 8512 6472 8522
rect 6423 8506 6453 8512
rect 6472 8507 6477 8512
rect 6395 8490 6469 8506
rect 6487 8498 6517 8554
rect 6552 8544 6760 8554
rect 6795 8550 6840 8554
rect 6843 8553 6844 8554
rect 6859 8553 6872 8554
rect 6578 8514 6767 8544
rect 6593 8511 6767 8514
rect 6586 8508 6767 8511
rect 6395 8488 6408 8490
rect 6423 8488 6457 8490
rect 6395 8472 6469 8488
rect 6496 8484 6509 8498
rect 6524 8484 6540 8500
rect 6586 8495 6597 8508
rect 6105 8440 6208 8450
rect 6059 8438 6208 8440
rect 6229 8438 6264 8450
rect 5898 8436 6060 8438
rect 5910 8416 5929 8436
rect 5944 8434 5974 8436
rect 5793 8408 5834 8416
rect 5916 8412 5929 8416
rect 5981 8420 6060 8436
rect 6092 8436 6264 8438
rect 6092 8420 6171 8436
rect 6178 8434 6208 8436
rect 5756 8398 5785 8408
rect 5799 8398 5828 8408
rect 5843 8398 5873 8412
rect 5916 8398 5959 8412
rect 5981 8408 6171 8420
rect 6236 8416 6242 8436
rect 5966 8398 5996 8408
rect 5997 8398 6155 8408
rect 6159 8398 6189 8408
rect 6193 8398 6223 8412
rect 6251 8398 6264 8436
rect 6336 8450 6365 8451
rect 6379 8451 6380 8466
rect 6395 8451 6408 8472
rect 6423 8451 6453 8472
rect 6496 8468 6558 8484
rect 6586 8477 6597 8493
rect 6602 8488 6612 8508
rect 6622 8488 6636 8508
rect 6639 8495 6648 8508
rect 6664 8495 6673 8508
rect 6602 8477 6636 8488
rect 6639 8477 6648 8493
rect 6664 8477 6673 8493
rect 6680 8488 6690 8508
rect 6700 8488 6714 8508
rect 6715 8495 6726 8508
rect 6680 8477 6714 8488
rect 6715 8477 6726 8493
rect 6772 8484 6788 8500
rect 6795 8498 6825 8550
rect 6859 8546 6860 8553
rect 6844 8538 6860 8546
rect 6831 8506 6844 8525
rect 6859 8506 6889 8522
rect 6831 8490 6905 8506
rect 6831 8488 6844 8490
rect 6859 8488 6893 8490
rect 6496 8466 6509 8468
rect 6524 8466 6558 8468
rect 6496 8451 6558 8466
rect 6602 8461 6618 8464
rect 6680 8461 6710 8472
rect 6758 8468 6804 8484
rect 6831 8472 6905 8488
rect 6758 8466 6792 8468
rect 6757 8451 6804 8466
rect 6379 8450 6408 8451
rect 6490 8450 6570 8451
rect 6577 8450 6587 8451
rect 6336 8442 6371 8450
rect 6336 8416 6337 8442
rect 6344 8416 6371 8442
rect 6279 8398 6309 8412
rect 6336 8408 6371 8416
rect 6373 8442 6414 8450
rect 6373 8416 6388 8442
rect 6395 8416 6414 8442
rect 6478 8438 6509 8450
rect 6524 8438 6627 8450
rect 6639 8440 6665 8451
rect 6742 8450 6804 8451
rect 6816 8450 6822 8451
rect 6831 8450 6844 8472
rect 6859 8451 6889 8472
rect 6916 8451 6917 8466
rect 6932 8451 6945 8610
rect 6975 8506 6988 8610
rect 7033 8588 7034 8598
rect 7049 8588 7062 8598
rect 7033 8584 7062 8588
rect 7067 8584 7097 8610
rect 7115 8596 7131 8598
rect 7203 8596 7256 8610
rect 7204 8594 7268 8596
rect 7311 8594 7326 8610
rect 7375 8607 7405 8610
rect 7375 8604 7411 8607
rect 7341 8596 7357 8598
rect 7115 8584 7130 8588
rect 7033 8582 7130 8584
rect 7158 8582 7326 8594
rect 7342 8584 7357 8588
rect 7375 8585 7414 8604
rect 7433 8598 7440 8599
rect 7439 8591 7440 8598
rect 7423 8588 7424 8591
rect 7439 8588 7452 8591
rect 7375 8584 7405 8585
rect 7414 8584 7420 8585
rect 7423 8584 7452 8588
rect 7342 8583 7452 8584
rect 7342 8582 7458 8583
rect 7017 8574 7068 8582
rect 7017 8562 7042 8574
rect 7049 8562 7068 8574
rect 7099 8574 7149 8582
rect 7099 8566 7115 8574
rect 7122 8572 7149 8574
rect 7158 8572 7379 8582
rect 7122 8562 7379 8572
rect 7408 8574 7458 8582
rect 7408 8565 7424 8574
rect 7017 8554 7068 8562
rect 7115 8554 7379 8562
rect 7405 8562 7424 8565
rect 7431 8562 7458 8574
rect 7405 8554 7458 8562
rect 7033 8546 7034 8554
rect 7049 8546 7062 8554
rect 7033 8538 7049 8546
rect 7030 8531 7049 8534
rect 7030 8522 7052 8531
rect 7003 8512 7052 8522
rect 7003 8506 7033 8512
rect 7052 8507 7057 8512
rect 6975 8490 7049 8506
rect 7067 8498 7097 8554
rect 7132 8544 7340 8554
rect 7375 8550 7420 8554
rect 7423 8553 7424 8554
rect 7439 8553 7452 8554
rect 7158 8514 7347 8544
rect 7173 8511 7347 8514
rect 7166 8508 7347 8511
rect 6975 8488 6988 8490
rect 7003 8488 7037 8490
rect 6975 8472 7049 8488
rect 7076 8484 7089 8498
rect 7104 8484 7120 8500
rect 7166 8495 7177 8508
rect 6685 8440 6788 8450
rect 6639 8438 6788 8440
rect 6809 8438 6844 8450
rect 6478 8436 6640 8438
rect 6490 8416 6509 8436
rect 6524 8434 6554 8436
rect 6373 8408 6414 8416
rect 6496 8412 6509 8416
rect 6561 8420 6640 8436
rect 6672 8436 6844 8438
rect 6672 8420 6751 8436
rect 6758 8434 6788 8436
rect 6336 8398 6365 8408
rect 6379 8398 6408 8408
rect 6423 8398 6453 8412
rect 6496 8398 6539 8412
rect 6561 8408 6751 8420
rect 6816 8416 6822 8436
rect 6546 8398 6576 8408
rect 6577 8398 6735 8408
rect 6739 8398 6769 8408
rect 6773 8398 6803 8412
rect 6831 8398 6844 8436
rect 6916 8450 6945 8451
rect 6959 8451 6960 8466
rect 6975 8451 6988 8472
rect 7003 8451 7033 8472
rect 7076 8468 7138 8484
rect 7166 8477 7177 8493
rect 7182 8488 7192 8508
rect 7202 8488 7216 8508
rect 7219 8495 7228 8508
rect 7244 8495 7253 8508
rect 7182 8477 7216 8488
rect 7219 8477 7228 8493
rect 7244 8477 7253 8493
rect 7260 8488 7270 8508
rect 7280 8488 7294 8508
rect 7295 8495 7306 8508
rect 7260 8477 7294 8488
rect 7295 8477 7306 8493
rect 7352 8484 7368 8500
rect 7375 8498 7405 8550
rect 7439 8546 7440 8553
rect 7424 8538 7440 8546
rect 7411 8506 7424 8525
rect 7439 8506 7469 8522
rect 7411 8490 7485 8506
rect 7411 8488 7424 8490
rect 7439 8488 7473 8490
rect 7076 8466 7089 8468
rect 7104 8466 7138 8468
rect 7076 8451 7138 8466
rect 7182 8461 7198 8464
rect 7260 8461 7290 8472
rect 7338 8468 7384 8484
rect 7411 8472 7485 8488
rect 7338 8466 7372 8468
rect 7337 8451 7384 8466
rect 6959 8450 6988 8451
rect 7070 8450 7150 8451
rect 7157 8450 7167 8451
rect 6916 8442 6951 8450
rect 6916 8416 6917 8442
rect 6924 8416 6951 8442
rect 6859 8398 6889 8412
rect 6916 8408 6951 8416
rect 6953 8442 6994 8450
rect 6953 8416 6968 8442
rect 6975 8416 6994 8442
rect 7058 8438 7089 8450
rect 7104 8438 7207 8450
rect 7219 8440 7245 8451
rect 7322 8450 7384 8451
rect 7396 8450 7402 8451
rect 7411 8450 7424 8472
rect 7439 8451 7469 8472
rect 7496 8451 7497 8466
rect 7512 8451 7525 8610
rect 7555 8506 7568 8610
rect 7613 8588 7614 8598
rect 7629 8588 7642 8598
rect 7613 8584 7642 8588
rect 7647 8584 7677 8610
rect 7695 8596 7711 8598
rect 7783 8596 7836 8610
rect 7784 8594 7848 8596
rect 7891 8594 7906 8610
rect 7955 8607 7985 8610
rect 7955 8604 7991 8607
rect 7921 8596 7937 8598
rect 7695 8584 7710 8588
rect 7613 8582 7710 8584
rect 7738 8582 7906 8594
rect 7922 8584 7937 8588
rect 7955 8585 7994 8604
rect 8013 8598 8020 8599
rect 8019 8591 8020 8598
rect 8003 8588 8004 8591
rect 8019 8588 8032 8591
rect 7955 8584 7985 8585
rect 7994 8584 8000 8585
rect 8003 8584 8032 8588
rect 7922 8583 8032 8584
rect 7922 8582 8038 8583
rect 7597 8574 7648 8582
rect 7597 8562 7622 8574
rect 7629 8562 7648 8574
rect 7679 8574 7729 8582
rect 7679 8566 7695 8574
rect 7702 8572 7729 8574
rect 7738 8572 7959 8582
rect 7702 8562 7959 8572
rect 7988 8574 8038 8582
rect 7988 8565 8004 8574
rect 7597 8554 7648 8562
rect 7695 8554 7959 8562
rect 7985 8562 8004 8565
rect 8011 8562 8038 8574
rect 7985 8554 8038 8562
rect 7613 8546 7614 8554
rect 7629 8546 7642 8554
rect 7613 8538 7629 8546
rect 7610 8531 7629 8534
rect 7610 8522 7632 8531
rect 7583 8512 7632 8522
rect 7583 8506 7613 8512
rect 7632 8507 7637 8512
rect 7555 8490 7629 8506
rect 7647 8498 7677 8554
rect 7712 8544 7920 8554
rect 7955 8550 8000 8554
rect 8003 8553 8004 8554
rect 8019 8553 8032 8554
rect 7738 8514 7927 8544
rect 7753 8511 7927 8514
rect 7746 8508 7927 8511
rect 7555 8488 7568 8490
rect 7583 8488 7617 8490
rect 7555 8472 7629 8488
rect 7656 8484 7669 8498
rect 7684 8484 7700 8500
rect 7746 8495 7757 8508
rect 7265 8440 7368 8450
rect 7219 8438 7368 8440
rect 7389 8438 7424 8450
rect 7058 8436 7220 8438
rect 7070 8416 7089 8436
rect 7104 8434 7134 8436
rect 6953 8408 6994 8416
rect 7076 8412 7089 8416
rect 7141 8420 7220 8436
rect 7252 8436 7424 8438
rect 7252 8420 7331 8436
rect 7338 8434 7368 8436
rect 6916 8398 6945 8408
rect 6959 8398 6988 8408
rect 7003 8398 7033 8412
rect 7076 8398 7119 8412
rect 7141 8408 7331 8420
rect 7396 8416 7402 8436
rect 7126 8398 7156 8408
rect 7157 8398 7315 8408
rect 7319 8398 7349 8408
rect 7353 8398 7383 8412
rect 7411 8398 7424 8436
rect 7496 8450 7525 8451
rect 7539 8451 7540 8466
rect 7555 8451 7568 8472
rect 7539 8450 7568 8451
rect 7583 8450 7613 8472
rect 7656 8468 7718 8484
rect 7746 8477 7757 8493
rect 7762 8488 7772 8508
rect 7782 8488 7796 8508
rect 7799 8495 7808 8508
rect 7824 8495 7833 8508
rect 7762 8477 7796 8488
rect 7799 8477 7808 8493
rect 7824 8477 7833 8493
rect 7840 8488 7850 8508
rect 7860 8488 7874 8508
rect 7875 8495 7886 8508
rect 7840 8477 7874 8488
rect 7875 8477 7886 8493
rect 7932 8484 7948 8500
rect 7955 8498 7985 8550
rect 8019 8546 8020 8553
rect 8004 8538 8020 8546
rect 7991 8506 8004 8525
rect 8019 8506 8049 8522
rect 7991 8490 8065 8506
rect 7991 8488 8004 8490
rect 8019 8488 8053 8490
rect 7656 8466 7669 8468
rect 7684 8466 7718 8468
rect 7656 8450 7718 8466
rect 7762 8461 7778 8464
rect 7840 8461 7870 8472
rect 7918 8468 7964 8484
rect 7991 8472 8065 8488
rect 7918 8466 7952 8468
rect 7917 8450 7964 8466
rect 7991 8450 8004 8472
rect 8019 8450 8049 8472
rect 8076 8450 8077 8466
rect 8092 8450 8105 8610
rect 8135 8506 8148 8610
rect 8193 8588 8194 8598
rect 8209 8588 8222 8598
rect 8193 8584 8222 8588
rect 8227 8584 8257 8610
rect 8275 8596 8291 8598
rect 8363 8596 8416 8610
rect 8364 8594 8428 8596
rect 8471 8594 8486 8610
rect 8535 8607 8565 8610
rect 8535 8604 8571 8607
rect 8501 8596 8517 8598
rect 8275 8584 8290 8588
rect 8193 8582 8290 8584
rect 8318 8582 8486 8594
rect 8502 8584 8517 8588
rect 8535 8585 8574 8604
rect 8593 8598 8600 8599
rect 8599 8591 8600 8598
rect 8583 8588 8584 8591
rect 8599 8588 8612 8591
rect 8535 8584 8565 8585
rect 8574 8584 8580 8585
rect 8583 8584 8612 8588
rect 8502 8583 8612 8584
rect 8502 8582 8618 8583
rect 8177 8574 8228 8582
rect 8177 8562 8202 8574
rect 8209 8562 8228 8574
rect 8259 8574 8309 8582
rect 8259 8566 8275 8574
rect 8282 8572 8309 8574
rect 8318 8572 8539 8582
rect 8282 8562 8539 8572
rect 8568 8574 8618 8582
rect 8568 8565 8584 8574
rect 8177 8554 8228 8562
rect 8275 8554 8539 8562
rect 8565 8562 8584 8565
rect 8591 8562 8618 8574
rect 8565 8554 8618 8562
rect 8193 8546 8194 8554
rect 8209 8546 8222 8554
rect 8193 8538 8209 8546
rect 8190 8531 8209 8534
rect 8190 8522 8212 8531
rect 8163 8512 8212 8522
rect 8163 8506 8193 8512
rect 8212 8507 8217 8512
rect 8135 8490 8209 8506
rect 8227 8498 8257 8554
rect 8292 8544 8500 8554
rect 8535 8550 8580 8554
rect 8583 8553 8584 8554
rect 8599 8553 8612 8554
rect 8318 8514 8507 8544
rect 8333 8511 8507 8514
rect 8326 8508 8507 8511
rect 8135 8488 8148 8490
rect 8163 8488 8197 8490
rect 8135 8472 8209 8488
rect 8236 8484 8249 8498
rect 8264 8484 8280 8500
rect 8326 8495 8337 8508
rect 8119 8450 8120 8466
rect 8135 8450 8148 8472
rect 8163 8450 8193 8472
rect 8236 8468 8298 8484
rect 8326 8477 8337 8493
rect 8342 8488 8352 8508
rect 8362 8488 8376 8508
rect 8379 8495 8388 8508
rect 8404 8495 8413 8508
rect 8342 8477 8376 8488
rect 8379 8477 8388 8493
rect 8404 8477 8413 8493
rect 8420 8488 8430 8508
rect 8440 8488 8454 8508
rect 8455 8495 8466 8508
rect 8420 8477 8454 8488
rect 8455 8477 8466 8493
rect 8512 8484 8528 8500
rect 8535 8498 8565 8550
rect 8599 8546 8600 8553
rect 8584 8538 8600 8546
rect 8571 8506 8584 8525
rect 8599 8506 8629 8522
rect 8571 8490 8645 8506
rect 8571 8488 8584 8490
rect 8599 8488 8633 8490
rect 8236 8466 8249 8468
rect 8264 8466 8298 8468
rect 8236 8450 8298 8466
rect 8342 8461 8358 8464
rect 8420 8461 8450 8472
rect 8498 8468 8544 8484
rect 8571 8472 8645 8488
rect 8498 8466 8532 8468
rect 8497 8450 8544 8466
rect 8571 8450 8584 8472
rect 8599 8450 8629 8472
rect 8656 8450 8657 8466
rect 8672 8450 8685 8610
rect 8715 8506 8728 8610
rect 8773 8588 8774 8598
rect 8789 8588 8802 8598
rect 8773 8584 8802 8588
rect 8807 8584 8837 8610
rect 8855 8596 8871 8598
rect 8943 8596 8996 8610
rect 8944 8594 9008 8596
rect 9051 8594 9066 8610
rect 9115 8607 9145 8610
rect 9115 8604 9151 8607
rect 9081 8596 9097 8598
rect 8855 8584 8870 8588
rect 8773 8582 8870 8584
rect 8898 8582 9066 8594
rect 9082 8584 9097 8588
rect 9115 8585 9154 8604
rect 9173 8598 9180 8599
rect 9179 8591 9180 8598
rect 9163 8588 9164 8591
rect 9179 8588 9192 8591
rect 9115 8584 9145 8585
rect 9154 8584 9160 8585
rect 9163 8584 9192 8588
rect 9082 8583 9192 8584
rect 9082 8582 9198 8583
rect 8757 8574 8808 8582
rect 8757 8562 8782 8574
rect 8789 8562 8808 8574
rect 8839 8574 8889 8582
rect 8839 8566 8855 8574
rect 8862 8572 8889 8574
rect 8898 8572 9119 8582
rect 8862 8562 9119 8572
rect 9148 8574 9198 8582
rect 9148 8565 9164 8574
rect 8757 8554 8808 8562
rect 8855 8554 9119 8562
rect 9145 8562 9164 8565
rect 9171 8562 9198 8574
rect 9145 8554 9198 8562
rect 8773 8546 8774 8554
rect 8789 8546 8802 8554
rect 8773 8538 8789 8546
rect 8770 8531 8789 8534
rect 8770 8522 8792 8531
rect 8743 8512 8792 8522
rect 8743 8506 8773 8512
rect 8792 8507 8797 8512
rect 8715 8490 8789 8506
rect 8807 8498 8837 8554
rect 8872 8544 9080 8554
rect 9115 8550 9160 8554
rect 9163 8553 9164 8554
rect 9179 8553 9192 8554
rect 8898 8514 9087 8544
rect 8913 8511 9087 8514
rect 8906 8508 9087 8511
rect 8715 8488 8728 8490
rect 8743 8488 8777 8490
rect 8715 8472 8789 8488
rect 8816 8484 8829 8498
rect 8844 8484 8860 8500
rect 8906 8495 8917 8508
rect 8699 8450 8700 8466
rect 8715 8450 8728 8472
rect 8743 8450 8773 8472
rect 8816 8468 8878 8484
rect 8906 8477 8917 8493
rect 8922 8488 8932 8508
rect 8942 8488 8956 8508
rect 8959 8495 8968 8508
rect 8984 8495 8993 8508
rect 8922 8477 8956 8488
rect 8959 8477 8968 8493
rect 8984 8477 8993 8493
rect 9000 8488 9010 8508
rect 9020 8488 9034 8508
rect 9035 8495 9046 8508
rect 9000 8477 9034 8488
rect 9035 8477 9046 8493
rect 9092 8484 9108 8500
rect 9115 8498 9145 8550
rect 9179 8546 9180 8553
rect 9164 8538 9180 8546
rect 9151 8506 9164 8525
rect 9179 8506 9209 8522
rect 9151 8490 9225 8506
rect 9151 8488 9164 8490
rect 9179 8488 9213 8490
rect 8816 8466 8829 8468
rect 8844 8466 8878 8468
rect 8816 8450 8878 8466
rect 8922 8461 8938 8464
rect 9000 8461 9030 8472
rect 9078 8468 9124 8484
rect 9151 8472 9225 8488
rect 9078 8466 9112 8468
rect 9077 8450 9124 8466
rect 9151 8450 9164 8472
rect 9179 8450 9209 8472
rect 9236 8450 9237 8466
rect 9252 8450 9265 8610
rect 7496 8442 7531 8450
rect 7496 8416 7497 8442
rect 7504 8416 7531 8442
rect 7439 8398 7469 8412
rect 7496 8408 7531 8416
rect 7533 8442 7574 8450
rect 7533 8416 7548 8442
rect 7555 8416 7574 8442
rect 7638 8438 7700 8450
rect 7712 8438 7787 8450
rect 7845 8438 7920 8450
rect 7932 8438 7963 8450
rect 7969 8438 8004 8450
rect 7638 8436 7800 8438
rect 7533 8408 7574 8416
rect 7656 8412 7669 8436
rect 7684 8434 7699 8436
rect 7496 8398 7525 8408
rect 7539 8398 7568 8408
rect 7583 8398 7613 8412
rect 7656 8398 7699 8412
rect 7723 8409 7730 8416
rect 7733 8412 7800 8436
rect 7832 8436 8004 8438
rect 7802 8414 7830 8418
rect 7832 8414 7912 8436
rect 7933 8434 7948 8436
rect 7802 8412 7912 8414
rect 7733 8408 7912 8412
rect 7706 8398 7736 8408
rect 7738 8398 7891 8408
rect 7899 8398 7929 8408
rect 7933 8398 7963 8412
rect 7991 8398 8004 8436
rect 8076 8442 8111 8450
rect 8076 8416 8077 8442
rect 8084 8416 8111 8442
rect 8019 8398 8049 8412
rect 8076 8408 8111 8416
rect 8113 8442 8154 8450
rect 8113 8416 8128 8442
rect 8135 8416 8154 8442
rect 8218 8438 8280 8450
rect 8292 8438 8367 8450
rect 8425 8438 8500 8450
rect 8512 8438 8543 8450
rect 8549 8438 8584 8450
rect 8218 8436 8380 8438
rect 8113 8408 8154 8416
rect 8236 8412 8249 8436
rect 8264 8434 8279 8436
rect 8076 8398 8077 8408
rect 8092 8398 8105 8408
rect 8119 8398 8120 8408
rect 8135 8398 8148 8408
rect 8163 8398 8193 8412
rect 8236 8398 8279 8412
rect 8303 8409 8310 8416
rect 8313 8412 8380 8436
rect 8412 8436 8584 8438
rect 8382 8414 8410 8418
rect 8412 8414 8492 8436
rect 8513 8434 8528 8436
rect 8382 8412 8492 8414
rect 8313 8408 8492 8412
rect 8286 8398 8316 8408
rect 8318 8398 8471 8408
rect 8479 8398 8509 8408
rect 8513 8398 8543 8412
rect 8571 8398 8584 8436
rect 8656 8442 8691 8450
rect 8656 8416 8657 8442
rect 8664 8416 8691 8442
rect 8599 8398 8629 8412
rect 8656 8408 8691 8416
rect 8693 8442 8734 8450
rect 8693 8416 8708 8442
rect 8715 8416 8734 8442
rect 8798 8438 8860 8450
rect 8872 8438 8947 8450
rect 9005 8438 9080 8450
rect 9092 8438 9123 8450
rect 9129 8438 9164 8450
rect 8798 8436 8960 8438
rect 8693 8408 8734 8416
rect 8816 8412 8829 8436
rect 8844 8434 8859 8436
rect 8656 8398 8657 8408
rect 8672 8398 8685 8408
rect 8699 8398 8700 8408
rect 8715 8398 8728 8408
rect 8743 8398 8773 8412
rect 8816 8398 8859 8412
rect 8883 8409 8890 8416
rect 8893 8412 8960 8436
rect 8992 8436 9164 8438
rect 8962 8414 8990 8418
rect 8992 8414 9072 8436
rect 9093 8434 9108 8436
rect 8962 8412 9072 8414
rect 8893 8408 9072 8412
rect 8866 8398 8896 8408
rect 8898 8398 9051 8408
rect 9059 8398 9089 8408
rect 9093 8398 9123 8412
rect 9151 8398 9164 8436
rect 9236 8442 9271 8450
rect 9236 8416 9237 8442
rect 9244 8416 9271 8442
rect 9179 8398 9209 8412
rect 9236 8408 9271 8416
rect 9236 8398 9237 8408
rect 9252 8398 9265 8408
rect -1 8392 9265 8398
rect 0 8384 9265 8392
rect 15 8354 28 8384
rect 43 8366 73 8384
rect 116 8370 130 8384
rect 166 8370 386 8384
rect 117 8368 130 8370
rect 83 8356 98 8368
rect 80 8354 102 8356
rect 107 8354 137 8368
rect 198 8366 351 8370
rect 180 8354 372 8366
rect 415 8354 445 8368
rect 451 8354 464 8384
rect 479 8366 509 8384
rect 552 8354 565 8384
rect 595 8354 608 8384
rect 623 8366 653 8384
rect 696 8370 710 8384
rect 746 8370 966 8384
rect 697 8368 710 8370
rect 663 8356 678 8368
rect 660 8354 682 8356
rect 687 8354 717 8368
rect 778 8366 931 8370
rect 760 8354 952 8366
rect 995 8354 1025 8368
rect 1031 8354 1044 8384
rect 1059 8366 1089 8384
rect 1132 8354 1145 8384
rect 1175 8354 1188 8384
rect 1203 8366 1233 8384
rect 1276 8370 1290 8384
rect 1326 8370 1546 8384
rect 1277 8368 1290 8370
rect 1243 8356 1258 8368
rect 1240 8354 1262 8356
rect 1267 8354 1297 8368
rect 1358 8366 1511 8370
rect 1340 8354 1532 8366
rect 1575 8354 1605 8368
rect 1611 8354 1624 8384
rect 1639 8366 1669 8384
rect 1712 8354 1725 8384
rect 1755 8354 1768 8384
rect 1783 8370 1813 8384
rect 1856 8370 1899 8384
rect 1906 8370 2126 8384
rect 2133 8370 2163 8384
rect 1823 8356 1838 8368
rect 1857 8356 1870 8370
rect 1938 8366 2091 8370
rect 1820 8354 1842 8356
rect 1920 8354 2112 8366
rect 2191 8354 2204 8384
rect 2219 8370 2249 8384
rect 2286 8354 2305 8384
rect 2320 8354 2326 8384
rect 2335 8354 2348 8384
rect 2363 8370 2393 8384
rect 2436 8370 2479 8384
rect 2486 8370 2706 8384
rect 2713 8370 2743 8384
rect 2403 8356 2418 8368
rect 2437 8356 2450 8370
rect 2518 8366 2671 8370
rect 2400 8354 2422 8356
rect 2500 8354 2692 8366
rect 2771 8354 2784 8384
rect 2799 8370 2829 8384
rect 2866 8354 2885 8384
rect 2900 8354 2906 8384
rect 2915 8354 2928 8384
rect 2943 8370 2973 8384
rect 3016 8370 3059 8384
rect 3066 8370 3286 8384
rect 3293 8370 3323 8384
rect 2983 8356 2998 8368
rect 3017 8356 3030 8370
rect 3098 8366 3251 8370
rect 2980 8354 3002 8356
rect 3080 8354 3272 8366
rect 3351 8354 3364 8384
rect 3379 8370 3409 8384
rect 3446 8354 3465 8384
rect 3480 8354 3486 8384
rect 3495 8354 3508 8384
rect 3523 8370 3553 8384
rect 3596 8370 3639 8384
rect 3646 8370 3866 8384
rect 3873 8370 3903 8384
rect 3563 8356 3578 8368
rect 3597 8356 3610 8370
rect 3678 8366 3831 8370
rect 3560 8354 3582 8356
rect 3660 8354 3852 8366
rect 3931 8354 3944 8384
rect 3959 8370 3989 8384
rect 4026 8354 4045 8384
rect 4060 8354 4066 8384
rect 4075 8354 4088 8384
rect 4103 8370 4133 8384
rect 4176 8370 4219 8384
rect 4226 8370 4446 8384
rect 4453 8370 4483 8384
rect 4143 8356 4158 8368
rect 4177 8356 4190 8370
rect 4258 8366 4411 8370
rect 4140 8354 4162 8356
rect 4240 8354 4432 8366
rect 4511 8354 4524 8384
rect 4539 8370 4569 8384
rect 4606 8354 4625 8384
rect 4640 8354 4646 8384
rect 4655 8354 4668 8384
rect 4683 8370 4713 8384
rect 4756 8370 4799 8384
rect 4806 8370 5026 8384
rect 5033 8370 5063 8384
rect 4723 8356 4738 8368
rect 4757 8356 4770 8370
rect 4838 8366 4991 8370
rect 4720 8354 4742 8356
rect 4820 8354 5012 8366
rect 5091 8354 5104 8384
rect 5119 8370 5149 8384
rect 5186 8354 5205 8384
rect 5220 8354 5226 8384
rect 5235 8354 5248 8384
rect 5263 8370 5293 8384
rect 5336 8370 5379 8384
rect 5386 8370 5606 8384
rect 5613 8370 5643 8384
rect 5303 8356 5318 8368
rect 5337 8356 5350 8370
rect 5418 8366 5571 8370
rect 5300 8354 5322 8356
rect 5400 8354 5592 8366
rect 5671 8354 5684 8384
rect 5699 8370 5729 8384
rect 5766 8354 5785 8384
rect 5800 8354 5806 8384
rect 5815 8354 5828 8384
rect 5843 8370 5873 8384
rect 5916 8370 5959 8384
rect 5966 8370 6186 8384
rect 6193 8370 6223 8384
rect 5883 8356 5898 8368
rect 5917 8356 5930 8370
rect 5998 8366 6151 8370
rect 5880 8354 5902 8356
rect 5980 8354 6172 8366
rect 6251 8354 6264 8384
rect 6279 8370 6309 8384
rect 6346 8354 6365 8384
rect 6380 8354 6386 8384
rect 6395 8354 6408 8384
rect 6423 8370 6453 8384
rect 6496 8370 6539 8384
rect 6546 8370 6766 8384
rect 6773 8370 6803 8384
rect 6463 8356 6478 8368
rect 6497 8356 6510 8370
rect 6578 8366 6731 8370
rect 6460 8354 6482 8356
rect 6560 8354 6752 8366
rect 6831 8354 6844 8384
rect 6859 8370 6889 8384
rect 6926 8354 6945 8384
rect 6960 8354 6966 8384
rect 6975 8354 6988 8384
rect 7003 8370 7033 8384
rect 7076 8370 7119 8384
rect 7126 8370 7346 8384
rect 7353 8370 7383 8384
rect 7043 8356 7058 8368
rect 7077 8356 7090 8370
rect 7158 8366 7311 8370
rect 7040 8354 7062 8356
rect 7140 8354 7332 8366
rect 7411 8354 7424 8384
rect 7439 8370 7469 8384
rect 7506 8354 7525 8384
rect 7540 8354 7546 8384
rect 7555 8354 7568 8384
rect 7583 8366 7613 8384
rect 7656 8370 7670 8384
rect 7706 8370 7926 8384
rect 7657 8368 7670 8370
rect 7623 8356 7638 8368
rect 7620 8354 7642 8356
rect 7647 8354 7677 8368
rect 7738 8366 7891 8370
rect 7720 8354 7912 8366
rect 7955 8354 7985 8368
rect 7991 8354 8004 8384
rect 8019 8366 8049 8384
rect 8092 8354 8105 8384
rect 8135 8354 8148 8384
rect 8163 8366 8193 8384
rect 8236 8370 8250 8384
rect 8286 8370 8506 8384
rect 8237 8368 8250 8370
rect 8203 8356 8218 8368
rect 8200 8354 8222 8356
rect 8227 8354 8257 8368
rect 8318 8366 8471 8370
rect 8300 8354 8492 8366
rect 8535 8354 8565 8368
rect 8571 8354 8584 8384
rect 8599 8366 8629 8384
rect 8672 8354 8685 8384
rect 8715 8354 8728 8384
rect 8743 8366 8773 8384
rect 8816 8370 8830 8384
rect 8866 8370 9086 8384
rect 8817 8368 8830 8370
rect 8783 8356 8798 8368
rect 8780 8354 8802 8356
rect 8807 8354 8837 8368
rect 8898 8366 9051 8370
rect 8880 8354 9072 8366
rect 9115 8354 9145 8368
rect 9151 8354 9164 8384
rect 9179 8366 9209 8384
rect 9252 8354 9265 8384
rect 0 8340 9265 8354
rect 15 8236 28 8340
rect 73 8318 74 8328
rect 89 8318 102 8328
rect 73 8314 102 8318
rect 107 8314 137 8340
rect 155 8326 171 8328
rect 243 8326 296 8340
rect 244 8324 308 8326
rect 351 8324 366 8340
rect 415 8337 445 8340
rect 415 8334 451 8337
rect 381 8326 397 8328
rect 155 8314 170 8318
rect 73 8312 170 8314
rect 198 8312 366 8324
rect 382 8314 397 8318
rect 415 8315 454 8334
rect 473 8328 480 8329
rect 479 8321 480 8328
rect 463 8318 464 8321
rect 479 8318 492 8321
rect 415 8314 445 8315
rect 454 8314 460 8315
rect 463 8314 492 8318
rect 382 8313 492 8314
rect 382 8312 498 8313
rect 57 8304 108 8312
rect 57 8292 82 8304
rect 89 8292 108 8304
rect 139 8304 189 8312
rect 139 8296 155 8304
rect 162 8302 189 8304
rect 198 8302 419 8312
rect 162 8292 419 8302
rect 448 8304 498 8312
rect 448 8295 464 8304
rect 57 8284 108 8292
rect 155 8284 419 8292
rect 445 8292 464 8295
rect 471 8292 498 8304
rect 445 8284 498 8292
rect 73 8276 74 8284
rect 89 8276 102 8284
rect 73 8268 89 8276
rect 70 8261 89 8264
rect 70 8252 92 8261
rect 43 8242 92 8252
rect 43 8236 73 8242
rect 92 8237 97 8242
rect 15 8220 89 8236
rect 107 8228 137 8284
rect 172 8274 380 8284
rect 415 8280 460 8284
rect 463 8283 464 8284
rect 479 8283 492 8284
rect 198 8244 387 8274
rect 213 8241 387 8244
rect 206 8238 387 8241
rect 15 8218 28 8220
rect 43 8218 77 8220
rect 15 8202 89 8218
rect 116 8214 129 8228
rect 144 8214 160 8230
rect 206 8225 217 8238
rect -1 8180 0 8196
rect 15 8180 28 8202
rect 43 8180 73 8202
rect 116 8198 178 8214
rect 206 8207 217 8223
rect 222 8218 232 8238
rect 242 8218 256 8238
rect 259 8225 268 8238
rect 284 8225 293 8238
rect 222 8207 256 8218
rect 259 8207 268 8223
rect 284 8207 293 8223
rect 300 8218 310 8238
rect 320 8218 334 8238
rect 335 8225 346 8238
rect 300 8207 334 8218
rect 335 8207 346 8223
rect 392 8214 408 8230
rect 415 8228 445 8280
rect 479 8276 480 8283
rect 464 8268 480 8276
rect 451 8236 464 8255
rect 479 8236 509 8252
rect 451 8220 525 8236
rect 451 8218 464 8220
rect 479 8218 513 8220
rect 116 8196 129 8198
rect 144 8196 178 8198
rect 116 8180 178 8196
rect 222 8191 238 8194
rect 300 8191 330 8202
rect 378 8198 424 8214
rect 451 8202 525 8218
rect 378 8196 412 8198
rect 377 8180 424 8196
rect 451 8180 464 8202
rect 479 8180 509 8202
rect 536 8180 537 8196
rect 552 8180 565 8340
rect 595 8236 608 8340
rect 653 8318 654 8328
rect 669 8318 682 8328
rect 653 8314 682 8318
rect 687 8314 717 8340
rect 735 8326 751 8328
rect 823 8326 876 8340
rect 824 8324 888 8326
rect 931 8324 946 8340
rect 995 8337 1025 8340
rect 995 8334 1031 8337
rect 961 8326 977 8328
rect 735 8314 750 8318
rect 653 8312 750 8314
rect 778 8312 946 8324
rect 962 8314 977 8318
rect 995 8315 1034 8334
rect 1053 8328 1060 8329
rect 1059 8321 1060 8328
rect 1043 8318 1044 8321
rect 1059 8318 1072 8321
rect 995 8314 1025 8315
rect 1034 8314 1040 8315
rect 1043 8314 1072 8318
rect 962 8313 1072 8314
rect 962 8312 1078 8313
rect 637 8304 688 8312
rect 637 8292 662 8304
rect 669 8292 688 8304
rect 719 8304 769 8312
rect 719 8296 735 8304
rect 742 8302 769 8304
rect 778 8302 999 8312
rect 742 8292 999 8302
rect 1028 8304 1078 8312
rect 1028 8295 1044 8304
rect 637 8284 688 8292
rect 735 8284 999 8292
rect 1025 8292 1044 8295
rect 1051 8292 1078 8304
rect 1025 8284 1078 8292
rect 653 8276 654 8284
rect 669 8276 682 8284
rect 653 8268 669 8276
rect 650 8261 669 8264
rect 650 8252 672 8261
rect 623 8242 672 8252
rect 623 8236 653 8242
rect 672 8237 677 8242
rect 595 8220 669 8236
rect 687 8228 717 8284
rect 752 8274 960 8284
rect 995 8280 1040 8284
rect 1043 8283 1044 8284
rect 1059 8283 1072 8284
rect 778 8244 967 8274
rect 793 8241 967 8244
rect 786 8238 967 8241
rect 595 8218 608 8220
rect 623 8218 657 8220
rect 595 8202 669 8218
rect 696 8214 709 8228
rect 724 8214 740 8230
rect 786 8225 797 8238
rect 579 8180 580 8196
rect 595 8180 608 8202
rect 623 8180 653 8202
rect 696 8198 758 8214
rect 786 8207 797 8223
rect 802 8218 812 8238
rect 822 8218 836 8238
rect 839 8225 848 8238
rect 864 8225 873 8238
rect 802 8207 836 8218
rect 839 8207 848 8223
rect 864 8207 873 8223
rect 880 8218 890 8238
rect 900 8218 914 8238
rect 915 8225 926 8238
rect 880 8207 914 8218
rect 915 8207 926 8223
rect 972 8214 988 8230
rect 995 8228 1025 8280
rect 1059 8276 1060 8283
rect 1044 8268 1060 8276
rect 1031 8236 1044 8255
rect 1059 8236 1089 8252
rect 1031 8220 1105 8236
rect 1031 8218 1044 8220
rect 1059 8218 1093 8220
rect 696 8196 709 8198
rect 724 8196 758 8198
rect 696 8180 758 8196
rect 802 8191 818 8194
rect 880 8191 910 8202
rect 958 8198 1004 8214
rect 1031 8202 1105 8218
rect 958 8196 992 8198
rect 957 8180 1004 8196
rect 1031 8180 1044 8202
rect 1059 8180 1089 8202
rect 1116 8180 1117 8196
rect 1132 8180 1145 8340
rect 1175 8236 1188 8340
rect 1233 8318 1234 8328
rect 1249 8318 1262 8328
rect 1233 8314 1262 8318
rect 1267 8314 1297 8340
rect 1315 8326 1331 8328
rect 1403 8326 1456 8340
rect 1404 8324 1468 8326
rect 1511 8324 1526 8340
rect 1575 8337 1605 8340
rect 1575 8334 1611 8337
rect 1541 8326 1557 8328
rect 1315 8314 1330 8318
rect 1233 8312 1330 8314
rect 1358 8312 1526 8324
rect 1542 8314 1557 8318
rect 1575 8315 1614 8334
rect 1633 8328 1640 8329
rect 1639 8321 1640 8328
rect 1623 8318 1624 8321
rect 1639 8318 1652 8321
rect 1575 8314 1605 8315
rect 1614 8314 1620 8315
rect 1623 8314 1652 8318
rect 1542 8313 1652 8314
rect 1542 8312 1658 8313
rect 1217 8304 1268 8312
rect 1217 8292 1242 8304
rect 1249 8292 1268 8304
rect 1299 8304 1349 8312
rect 1299 8296 1315 8304
rect 1322 8302 1349 8304
rect 1358 8302 1579 8312
rect 1322 8292 1579 8302
rect 1608 8304 1658 8312
rect 1608 8295 1624 8304
rect 1217 8284 1268 8292
rect 1315 8284 1579 8292
rect 1605 8292 1624 8295
rect 1631 8292 1658 8304
rect 1605 8284 1658 8292
rect 1233 8276 1234 8284
rect 1249 8276 1262 8284
rect 1233 8268 1249 8276
rect 1230 8261 1249 8264
rect 1230 8252 1252 8261
rect 1203 8242 1252 8252
rect 1203 8236 1233 8242
rect 1252 8237 1257 8242
rect 1175 8220 1249 8236
rect 1267 8228 1297 8284
rect 1332 8274 1540 8284
rect 1575 8280 1620 8284
rect 1623 8283 1624 8284
rect 1639 8283 1652 8284
rect 1358 8244 1547 8274
rect 1373 8241 1547 8244
rect 1366 8238 1547 8241
rect 1175 8218 1188 8220
rect 1203 8218 1237 8220
rect 1175 8202 1249 8218
rect 1276 8214 1289 8228
rect 1304 8214 1320 8230
rect 1366 8225 1377 8238
rect 1159 8180 1160 8196
rect 1175 8180 1188 8202
rect 1203 8180 1233 8202
rect 1276 8198 1338 8214
rect 1366 8207 1377 8223
rect 1382 8218 1392 8238
rect 1402 8218 1416 8238
rect 1419 8225 1428 8238
rect 1444 8225 1453 8238
rect 1382 8207 1416 8218
rect 1419 8207 1428 8223
rect 1444 8207 1453 8223
rect 1460 8218 1470 8238
rect 1480 8218 1494 8238
rect 1495 8225 1506 8238
rect 1460 8207 1494 8218
rect 1495 8207 1506 8223
rect 1552 8214 1568 8230
rect 1575 8228 1605 8280
rect 1639 8276 1640 8283
rect 1624 8268 1640 8276
rect 1611 8236 1624 8255
rect 1639 8236 1669 8252
rect 1611 8220 1685 8236
rect 1611 8218 1624 8220
rect 1639 8218 1673 8220
rect 1276 8196 1289 8198
rect 1304 8196 1338 8198
rect 1276 8180 1338 8196
rect 1382 8191 1398 8194
rect 1460 8191 1490 8202
rect 1538 8198 1584 8214
rect 1611 8202 1685 8218
rect 1538 8196 1572 8198
rect 1537 8180 1584 8196
rect 1611 8180 1624 8202
rect 1639 8180 1669 8202
rect 1696 8180 1697 8196
rect 1712 8180 1725 8340
rect 1755 8236 1768 8340
rect 1820 8336 1842 8340
rect 1813 8314 1842 8328
rect 1895 8314 1911 8328
rect 1949 8324 1955 8326
rect 1962 8324 2070 8340
rect 2077 8324 2083 8326
rect 2091 8324 2106 8340
rect 2172 8334 2191 8337
rect 1813 8312 1911 8314
rect 1938 8312 2106 8324
rect 2121 8314 2137 8328
rect 2172 8315 2194 8334
rect 2204 8328 2220 8329
rect 2203 8326 2220 8328
rect 2204 8321 2220 8326
rect 2194 8314 2200 8315
rect 2203 8314 2232 8321
rect 2121 8313 2232 8314
rect 2121 8312 2238 8313
rect 1797 8304 1848 8312
rect 1895 8304 1929 8312
rect 1797 8292 1822 8304
rect 1829 8292 1848 8304
rect 1902 8302 1929 8304
rect 1938 8302 2159 8312
rect 2194 8309 2200 8312
rect 1902 8298 2159 8302
rect 1797 8284 1848 8292
rect 1895 8284 2159 8298
rect 2203 8304 2238 8312
rect 1813 8276 1842 8284
rect 1813 8270 1830 8276
rect 1813 8268 1847 8270
rect 1895 8268 1911 8284
rect 1912 8274 2120 8284
rect 2121 8274 2137 8284
rect 2185 8280 2200 8295
rect 2203 8292 2204 8304
rect 2211 8292 2238 8304
rect 2203 8284 2238 8292
rect 2203 8283 2232 8284
rect 1923 8270 2137 8274
rect 1938 8268 2137 8270
rect 2172 8270 2185 8280
rect 2203 8270 2220 8283
rect 2172 8268 2220 8270
rect 1814 8264 1847 8268
rect 1810 8262 1847 8264
rect 1810 8261 1877 8262
rect 1810 8256 1841 8261
rect 1847 8256 1877 8261
rect 1810 8252 1877 8256
rect 1783 8249 1877 8252
rect 1783 8242 1832 8249
rect 1783 8236 1813 8242
rect 1832 8237 1837 8242
rect 1755 8220 1829 8236
rect 1841 8228 1877 8249
rect 1938 8244 2127 8268
rect 2172 8267 2219 8268
rect 2185 8262 2219 8267
rect 1953 8241 2127 8244
rect 1946 8238 2127 8241
rect 2155 8261 2219 8262
rect 1755 8218 1768 8220
rect 1783 8218 1817 8220
rect 1755 8202 1829 8218
rect 1739 8180 1740 8196
rect 1755 8180 1768 8202
rect 1783 8186 1813 8202
rect 1841 8180 1847 8228
rect 1850 8222 1869 8228
rect 1884 8222 1914 8230
rect 1850 8214 1914 8222
rect 1850 8198 1930 8214
rect 1946 8207 2008 8238
rect 2024 8207 2086 8238
rect 2155 8236 2204 8261
rect 2219 8236 2249 8252
rect 2118 8222 2148 8230
rect 2155 8228 2265 8236
rect 2118 8214 2163 8222
rect 1850 8196 1869 8198
rect 1884 8196 1930 8198
rect 1850 8180 1930 8196
rect 1957 8194 1992 8207
rect 2033 8204 2070 8207
rect 2033 8202 2075 8204
rect 1962 8191 1992 8194
rect 1971 8187 1978 8191
rect 1978 8186 1979 8187
rect 1937 8180 1947 8186
rect -7 8172 34 8180
rect -7 8146 8 8172
rect 15 8146 34 8172
rect 98 8168 160 8180
rect 172 8168 247 8180
rect 305 8168 380 8180
rect 392 8168 423 8180
rect 429 8168 464 8180
rect 98 8166 260 8168
rect -7 8138 34 8146
rect 116 8142 129 8166
rect 144 8164 159 8166
rect -1 8128 0 8138
rect 15 8128 28 8138
rect 43 8128 73 8142
rect 116 8128 159 8142
rect 183 8139 190 8146
rect 193 8142 260 8166
rect 292 8166 464 8168
rect 262 8144 290 8148
rect 292 8144 372 8166
rect 393 8164 408 8166
rect 262 8142 372 8144
rect 193 8138 372 8142
rect 166 8128 196 8138
rect 198 8128 351 8138
rect 359 8128 389 8138
rect 393 8128 423 8142
rect 451 8128 464 8166
rect 536 8172 571 8180
rect 536 8146 537 8172
rect 544 8146 571 8172
rect 479 8128 509 8142
rect 536 8138 571 8146
rect 573 8172 614 8180
rect 573 8146 588 8172
rect 595 8146 614 8172
rect 678 8168 740 8180
rect 752 8168 827 8180
rect 885 8168 960 8180
rect 972 8168 1003 8180
rect 1009 8168 1044 8180
rect 678 8166 840 8168
rect 573 8138 614 8146
rect 696 8142 709 8166
rect 724 8164 739 8166
rect 536 8128 537 8138
rect 552 8128 565 8138
rect 579 8128 580 8138
rect 595 8128 608 8138
rect 623 8128 653 8142
rect 696 8128 739 8142
rect 763 8139 770 8146
rect 773 8142 840 8166
rect 872 8166 1044 8168
rect 842 8144 870 8148
rect 872 8144 952 8166
rect 973 8164 988 8166
rect 842 8142 952 8144
rect 773 8138 952 8142
rect 746 8128 776 8138
rect 778 8128 931 8138
rect 939 8128 969 8138
rect 973 8128 1003 8142
rect 1031 8128 1044 8166
rect 1116 8172 1151 8180
rect 1116 8146 1117 8172
rect 1124 8146 1151 8172
rect 1059 8128 1089 8142
rect 1116 8138 1151 8146
rect 1153 8172 1194 8180
rect 1153 8146 1168 8172
rect 1175 8146 1194 8172
rect 1258 8168 1320 8180
rect 1332 8168 1407 8180
rect 1465 8168 1540 8180
rect 1552 8168 1583 8180
rect 1589 8168 1624 8180
rect 1258 8166 1420 8168
rect 1153 8138 1194 8146
rect 1276 8142 1289 8166
rect 1304 8164 1319 8166
rect 1116 8128 1117 8138
rect 1132 8128 1145 8138
rect 1159 8128 1160 8138
rect 1175 8128 1188 8138
rect 1203 8128 1233 8142
rect 1276 8128 1319 8142
rect 1343 8139 1350 8146
rect 1353 8142 1420 8166
rect 1452 8166 1624 8168
rect 1422 8144 1450 8148
rect 1452 8144 1532 8166
rect 1553 8164 1568 8166
rect 1422 8142 1532 8144
rect 1353 8138 1532 8142
rect 1326 8128 1356 8138
rect 1358 8128 1511 8138
rect 1519 8128 1549 8138
rect 1553 8128 1583 8142
rect 1611 8128 1624 8166
rect 1696 8172 1731 8180
rect 1696 8146 1697 8172
rect 1704 8146 1731 8172
rect 1639 8128 1669 8142
rect 1696 8138 1731 8146
rect 1733 8172 1774 8180
rect 1733 8146 1748 8172
rect 1755 8146 1774 8172
rect 1838 8168 1869 8180
rect 1884 8168 1987 8180
rect 1999 8170 2025 8196
rect 2040 8191 2070 8202
rect 2102 8198 2164 8214
rect 2102 8196 2148 8198
rect 2102 8180 2164 8196
rect 2176 8180 2182 8228
rect 2185 8220 2265 8228
rect 2185 8218 2204 8220
rect 2219 8218 2253 8220
rect 2185 8202 2265 8218
rect 2185 8180 2204 8202
rect 2219 8186 2249 8202
rect 2277 8196 2283 8270
rect 2286 8196 2305 8340
rect 2320 8196 2326 8340
rect 2335 8270 2348 8340
rect 2400 8336 2422 8340
rect 2393 8314 2422 8328
rect 2475 8314 2491 8328
rect 2529 8324 2535 8326
rect 2542 8324 2650 8340
rect 2657 8324 2663 8326
rect 2671 8324 2686 8340
rect 2752 8334 2771 8337
rect 2393 8312 2491 8314
rect 2518 8312 2686 8324
rect 2701 8314 2717 8328
rect 2752 8315 2774 8334
rect 2784 8328 2800 8329
rect 2783 8326 2800 8328
rect 2784 8321 2800 8326
rect 2774 8314 2780 8315
rect 2783 8314 2812 8321
rect 2701 8313 2812 8314
rect 2701 8312 2818 8313
rect 2377 8304 2428 8312
rect 2475 8304 2509 8312
rect 2377 8292 2402 8304
rect 2409 8292 2428 8304
rect 2482 8302 2509 8304
rect 2518 8302 2739 8312
rect 2774 8309 2780 8312
rect 2482 8298 2739 8302
rect 2377 8284 2428 8292
rect 2475 8284 2739 8298
rect 2783 8304 2818 8312
rect 2329 8236 2348 8270
rect 2393 8276 2422 8284
rect 2393 8270 2410 8276
rect 2393 8268 2427 8270
rect 2475 8268 2491 8284
rect 2492 8274 2700 8284
rect 2701 8274 2717 8284
rect 2765 8280 2780 8295
rect 2783 8292 2784 8304
rect 2791 8292 2818 8304
rect 2783 8284 2818 8292
rect 2783 8283 2812 8284
rect 2503 8270 2717 8274
rect 2518 8268 2717 8270
rect 2752 8270 2765 8280
rect 2783 8270 2800 8283
rect 2752 8268 2800 8270
rect 2394 8264 2427 8268
rect 2390 8262 2427 8264
rect 2390 8261 2457 8262
rect 2390 8256 2421 8261
rect 2427 8256 2457 8261
rect 2390 8252 2457 8256
rect 2363 8249 2457 8252
rect 2363 8242 2412 8249
rect 2363 8236 2393 8242
rect 2412 8237 2417 8242
rect 2329 8220 2409 8236
rect 2421 8228 2457 8249
rect 2518 8244 2707 8268
rect 2752 8267 2799 8268
rect 2765 8262 2799 8267
rect 2533 8241 2707 8244
rect 2526 8238 2707 8241
rect 2735 8261 2799 8262
rect 2329 8218 2348 8220
rect 2363 8218 2397 8220
rect 2329 8202 2409 8218
rect 2329 8196 2348 8202
rect 2045 8170 2148 8180
rect 1999 8168 2148 8170
rect 2169 8168 2204 8180
rect 1838 8166 2000 8168
rect 1850 8146 1869 8166
rect 1884 8164 1914 8166
rect 1733 8138 1774 8146
rect 1856 8142 1869 8146
rect 1921 8150 2000 8166
rect 2032 8166 2204 8168
rect 2032 8150 2111 8166
rect 2118 8164 2148 8166
rect 1696 8128 1697 8138
rect 1712 8128 1725 8138
rect 1739 8128 1740 8138
rect 1755 8128 1768 8138
rect 1783 8128 1813 8142
rect 1856 8128 1899 8142
rect 1921 8138 2111 8150
rect 2176 8146 2182 8166
rect 1906 8128 1936 8138
rect 1937 8128 2095 8138
rect 2099 8128 2129 8138
rect 2133 8128 2163 8142
rect 2191 8128 2204 8166
rect 2276 8180 2305 8196
rect 2319 8180 2348 8196
rect 2363 8186 2393 8202
rect 2421 8180 2427 8228
rect 2430 8222 2449 8228
rect 2464 8222 2494 8230
rect 2430 8214 2494 8222
rect 2430 8198 2510 8214
rect 2526 8207 2588 8238
rect 2604 8207 2666 8238
rect 2735 8236 2784 8261
rect 2799 8236 2829 8252
rect 2698 8222 2728 8230
rect 2735 8228 2845 8236
rect 2698 8214 2743 8222
rect 2430 8196 2449 8198
rect 2464 8196 2510 8198
rect 2430 8180 2510 8196
rect 2537 8194 2572 8207
rect 2613 8204 2650 8207
rect 2613 8202 2655 8204
rect 2542 8191 2572 8194
rect 2551 8187 2558 8191
rect 2558 8186 2559 8187
rect 2517 8180 2527 8186
rect 2276 8172 2311 8180
rect 2276 8146 2277 8172
rect 2284 8146 2311 8172
rect 2219 8128 2249 8142
rect 2276 8138 2311 8146
rect 2313 8172 2354 8180
rect 2313 8146 2328 8172
rect 2335 8146 2354 8172
rect 2418 8168 2449 8180
rect 2464 8168 2567 8180
rect 2579 8170 2605 8196
rect 2620 8191 2650 8202
rect 2682 8198 2744 8214
rect 2682 8196 2728 8198
rect 2682 8180 2744 8196
rect 2756 8180 2762 8228
rect 2765 8220 2845 8228
rect 2765 8218 2784 8220
rect 2799 8218 2833 8220
rect 2765 8202 2845 8218
rect 2765 8180 2784 8202
rect 2799 8186 2829 8202
rect 2857 8196 2863 8270
rect 2866 8196 2885 8340
rect 2900 8196 2906 8340
rect 2915 8270 2928 8340
rect 2980 8336 3002 8340
rect 2973 8314 3002 8328
rect 3055 8314 3071 8328
rect 3109 8324 3115 8326
rect 3122 8324 3230 8340
rect 3237 8324 3243 8326
rect 3251 8324 3266 8340
rect 3332 8334 3351 8337
rect 2973 8312 3071 8314
rect 3098 8312 3266 8324
rect 3281 8314 3297 8328
rect 3332 8315 3354 8334
rect 3364 8328 3380 8329
rect 3363 8326 3380 8328
rect 3364 8321 3380 8326
rect 3354 8314 3360 8315
rect 3363 8314 3392 8321
rect 3281 8313 3392 8314
rect 3281 8312 3398 8313
rect 2957 8304 3008 8312
rect 3055 8304 3089 8312
rect 2957 8292 2982 8304
rect 2989 8292 3008 8304
rect 3062 8302 3089 8304
rect 3098 8302 3319 8312
rect 3354 8309 3360 8312
rect 3062 8298 3319 8302
rect 2957 8284 3008 8292
rect 3055 8284 3319 8298
rect 3363 8304 3398 8312
rect 2909 8236 2928 8270
rect 2973 8276 3002 8284
rect 2973 8270 2990 8276
rect 2973 8268 3007 8270
rect 3055 8268 3071 8284
rect 3072 8274 3280 8284
rect 3281 8274 3297 8284
rect 3345 8280 3360 8295
rect 3363 8292 3364 8304
rect 3371 8292 3398 8304
rect 3363 8284 3398 8292
rect 3363 8283 3392 8284
rect 3083 8270 3297 8274
rect 3098 8268 3297 8270
rect 3332 8270 3345 8280
rect 3363 8270 3380 8283
rect 3332 8268 3380 8270
rect 2974 8264 3007 8268
rect 2970 8262 3007 8264
rect 2970 8261 3037 8262
rect 2970 8256 3001 8261
rect 3007 8256 3037 8261
rect 2970 8252 3037 8256
rect 2943 8249 3037 8252
rect 2943 8242 2992 8249
rect 2943 8236 2973 8242
rect 2992 8237 2997 8242
rect 2909 8220 2989 8236
rect 3001 8228 3037 8249
rect 3098 8244 3287 8268
rect 3332 8267 3379 8268
rect 3345 8262 3379 8267
rect 3113 8241 3287 8244
rect 3106 8238 3287 8241
rect 3315 8261 3379 8262
rect 2909 8218 2928 8220
rect 2943 8218 2977 8220
rect 2909 8202 2989 8218
rect 2909 8196 2928 8202
rect 2625 8170 2728 8180
rect 2579 8168 2728 8170
rect 2749 8168 2784 8180
rect 2418 8166 2580 8168
rect 2430 8146 2449 8166
rect 2464 8164 2494 8166
rect 2313 8138 2354 8146
rect 2436 8142 2449 8146
rect 2501 8150 2580 8166
rect 2612 8166 2784 8168
rect 2612 8150 2691 8166
rect 2698 8164 2728 8166
rect 2276 8128 2305 8138
rect 2319 8128 2348 8138
rect 2363 8128 2393 8142
rect 2436 8128 2479 8142
rect 2501 8138 2691 8150
rect 2756 8146 2762 8166
rect 2486 8128 2516 8138
rect 2517 8128 2675 8138
rect 2679 8128 2709 8138
rect 2713 8128 2743 8142
rect 2771 8128 2784 8166
rect 2856 8180 2885 8196
rect 2899 8180 2928 8196
rect 2943 8186 2973 8202
rect 3001 8180 3007 8228
rect 3010 8222 3029 8228
rect 3044 8222 3074 8230
rect 3010 8214 3074 8222
rect 3010 8198 3090 8214
rect 3106 8207 3168 8238
rect 3184 8207 3246 8238
rect 3315 8236 3364 8261
rect 3379 8236 3409 8252
rect 3278 8222 3308 8230
rect 3315 8228 3425 8236
rect 3278 8214 3323 8222
rect 3010 8196 3029 8198
rect 3044 8196 3090 8198
rect 3010 8180 3090 8196
rect 3117 8194 3152 8207
rect 3193 8204 3230 8207
rect 3193 8202 3235 8204
rect 3122 8191 3152 8194
rect 3131 8187 3138 8191
rect 3138 8186 3139 8187
rect 3097 8180 3107 8186
rect 2856 8172 2891 8180
rect 2856 8146 2857 8172
rect 2864 8146 2891 8172
rect 2799 8128 2829 8142
rect 2856 8138 2891 8146
rect 2893 8172 2934 8180
rect 2893 8146 2908 8172
rect 2915 8146 2934 8172
rect 2998 8168 3029 8180
rect 3044 8168 3147 8180
rect 3159 8170 3185 8196
rect 3200 8191 3230 8202
rect 3262 8198 3324 8214
rect 3262 8196 3308 8198
rect 3262 8180 3324 8196
rect 3336 8180 3342 8228
rect 3345 8220 3425 8228
rect 3345 8218 3364 8220
rect 3379 8218 3413 8220
rect 3345 8202 3425 8218
rect 3345 8180 3364 8202
rect 3379 8186 3409 8202
rect 3437 8196 3443 8270
rect 3446 8196 3465 8340
rect 3480 8196 3486 8340
rect 3495 8270 3508 8340
rect 3560 8336 3582 8340
rect 3553 8314 3582 8328
rect 3635 8314 3651 8328
rect 3689 8324 3695 8326
rect 3702 8324 3810 8340
rect 3817 8324 3823 8326
rect 3831 8324 3846 8340
rect 3912 8334 3931 8337
rect 3553 8312 3651 8314
rect 3678 8312 3846 8324
rect 3861 8314 3877 8328
rect 3912 8315 3934 8334
rect 3944 8328 3960 8329
rect 3943 8326 3960 8328
rect 3944 8321 3960 8326
rect 3934 8314 3940 8315
rect 3943 8314 3972 8321
rect 3861 8313 3972 8314
rect 3861 8312 3978 8313
rect 3537 8304 3588 8312
rect 3635 8304 3669 8312
rect 3537 8292 3562 8304
rect 3569 8292 3588 8304
rect 3642 8302 3669 8304
rect 3678 8302 3899 8312
rect 3934 8309 3940 8312
rect 3642 8298 3899 8302
rect 3537 8284 3588 8292
rect 3635 8284 3899 8298
rect 3943 8304 3978 8312
rect 3489 8236 3508 8270
rect 3553 8276 3582 8284
rect 3553 8270 3570 8276
rect 3553 8268 3587 8270
rect 3635 8268 3651 8284
rect 3652 8274 3860 8284
rect 3861 8274 3877 8284
rect 3925 8280 3940 8295
rect 3943 8292 3944 8304
rect 3951 8292 3978 8304
rect 3943 8284 3978 8292
rect 3943 8283 3972 8284
rect 3663 8270 3877 8274
rect 3678 8268 3877 8270
rect 3912 8270 3925 8280
rect 3943 8270 3960 8283
rect 3912 8268 3960 8270
rect 3554 8264 3587 8268
rect 3550 8262 3587 8264
rect 3550 8261 3617 8262
rect 3550 8256 3581 8261
rect 3587 8256 3617 8261
rect 3550 8252 3617 8256
rect 3523 8249 3617 8252
rect 3523 8242 3572 8249
rect 3523 8236 3553 8242
rect 3572 8237 3577 8242
rect 3489 8220 3569 8236
rect 3581 8228 3617 8249
rect 3678 8244 3867 8268
rect 3912 8267 3959 8268
rect 3925 8262 3959 8267
rect 3693 8241 3867 8244
rect 3686 8238 3867 8241
rect 3895 8261 3959 8262
rect 3489 8218 3508 8220
rect 3523 8218 3557 8220
rect 3489 8202 3569 8218
rect 3489 8196 3508 8202
rect 3205 8170 3308 8180
rect 3159 8168 3308 8170
rect 3329 8168 3364 8180
rect 2998 8166 3160 8168
rect 3010 8146 3029 8166
rect 3044 8164 3074 8166
rect 2893 8138 2934 8146
rect 3016 8142 3029 8146
rect 3081 8150 3160 8166
rect 3192 8166 3364 8168
rect 3192 8150 3271 8166
rect 3278 8164 3308 8166
rect 2856 8128 2885 8138
rect 2899 8128 2928 8138
rect 2943 8128 2973 8142
rect 3016 8128 3059 8142
rect 3081 8138 3271 8150
rect 3336 8146 3342 8166
rect 3066 8128 3096 8138
rect 3097 8128 3255 8138
rect 3259 8128 3289 8138
rect 3293 8128 3323 8142
rect 3351 8128 3364 8166
rect 3436 8180 3465 8196
rect 3479 8180 3508 8196
rect 3523 8186 3553 8202
rect 3581 8180 3587 8228
rect 3590 8222 3609 8228
rect 3624 8222 3654 8230
rect 3590 8214 3654 8222
rect 3590 8198 3670 8214
rect 3686 8207 3748 8238
rect 3764 8207 3826 8238
rect 3895 8236 3944 8261
rect 3959 8236 3989 8252
rect 3858 8222 3888 8230
rect 3895 8228 4005 8236
rect 3858 8214 3903 8222
rect 3590 8196 3609 8198
rect 3624 8196 3670 8198
rect 3590 8180 3670 8196
rect 3697 8194 3732 8207
rect 3773 8204 3810 8207
rect 3773 8202 3815 8204
rect 3702 8191 3732 8194
rect 3711 8187 3718 8191
rect 3718 8186 3719 8187
rect 3677 8180 3687 8186
rect 3436 8172 3471 8180
rect 3436 8146 3437 8172
rect 3444 8146 3471 8172
rect 3379 8128 3409 8142
rect 3436 8138 3471 8146
rect 3473 8172 3514 8180
rect 3473 8146 3488 8172
rect 3495 8146 3514 8172
rect 3578 8168 3609 8180
rect 3624 8168 3727 8180
rect 3739 8170 3765 8196
rect 3780 8191 3810 8202
rect 3842 8198 3904 8214
rect 3842 8196 3888 8198
rect 3842 8180 3904 8196
rect 3916 8180 3922 8228
rect 3925 8220 4005 8228
rect 3925 8218 3944 8220
rect 3959 8218 3993 8220
rect 3925 8202 4005 8218
rect 3925 8180 3944 8202
rect 3959 8186 3989 8202
rect 4017 8196 4023 8270
rect 4026 8196 4045 8340
rect 4060 8196 4066 8340
rect 4075 8270 4088 8340
rect 4140 8336 4162 8340
rect 4133 8314 4162 8328
rect 4215 8314 4231 8328
rect 4269 8324 4275 8326
rect 4282 8324 4390 8340
rect 4397 8324 4403 8326
rect 4411 8324 4426 8340
rect 4492 8334 4511 8337
rect 4133 8312 4231 8314
rect 4258 8312 4426 8324
rect 4441 8314 4457 8328
rect 4492 8315 4514 8334
rect 4524 8328 4540 8329
rect 4523 8326 4540 8328
rect 4524 8321 4540 8326
rect 4514 8314 4520 8315
rect 4523 8314 4552 8321
rect 4441 8313 4552 8314
rect 4441 8312 4558 8313
rect 4117 8304 4168 8312
rect 4215 8304 4249 8312
rect 4117 8292 4142 8304
rect 4149 8292 4168 8304
rect 4222 8302 4249 8304
rect 4258 8302 4479 8312
rect 4514 8309 4520 8312
rect 4222 8298 4479 8302
rect 4117 8284 4168 8292
rect 4215 8284 4479 8298
rect 4523 8304 4558 8312
rect 4069 8236 4088 8270
rect 4133 8276 4162 8284
rect 4133 8270 4150 8276
rect 4133 8268 4167 8270
rect 4215 8268 4231 8284
rect 4232 8274 4440 8284
rect 4441 8274 4457 8284
rect 4505 8280 4520 8295
rect 4523 8292 4524 8304
rect 4531 8292 4558 8304
rect 4523 8284 4558 8292
rect 4523 8283 4552 8284
rect 4243 8270 4457 8274
rect 4258 8268 4457 8270
rect 4492 8270 4505 8280
rect 4523 8270 4540 8283
rect 4492 8268 4540 8270
rect 4134 8264 4167 8268
rect 4130 8262 4167 8264
rect 4130 8261 4197 8262
rect 4130 8256 4161 8261
rect 4167 8256 4197 8261
rect 4130 8252 4197 8256
rect 4103 8249 4197 8252
rect 4103 8242 4152 8249
rect 4103 8236 4133 8242
rect 4152 8237 4157 8242
rect 4069 8220 4149 8236
rect 4161 8228 4197 8249
rect 4258 8244 4447 8268
rect 4492 8267 4539 8268
rect 4505 8262 4539 8267
rect 4273 8241 4447 8244
rect 4266 8238 4447 8241
rect 4475 8261 4539 8262
rect 4069 8218 4088 8220
rect 4103 8218 4137 8220
rect 4069 8202 4149 8218
rect 4069 8196 4088 8202
rect 3785 8170 3888 8180
rect 3739 8168 3888 8170
rect 3909 8168 3944 8180
rect 3578 8166 3740 8168
rect 3590 8146 3609 8166
rect 3624 8164 3654 8166
rect 3473 8138 3514 8146
rect 3596 8142 3609 8146
rect 3661 8150 3740 8166
rect 3772 8166 3944 8168
rect 3772 8150 3851 8166
rect 3858 8164 3888 8166
rect 3436 8128 3465 8138
rect 3479 8128 3508 8138
rect 3523 8128 3553 8142
rect 3596 8128 3639 8142
rect 3661 8138 3851 8150
rect 3916 8146 3922 8166
rect 3646 8128 3676 8138
rect 3677 8128 3835 8138
rect 3839 8128 3869 8138
rect 3873 8128 3903 8142
rect 3931 8128 3944 8166
rect 4016 8180 4045 8196
rect 4059 8180 4088 8196
rect 4103 8186 4133 8202
rect 4161 8180 4167 8228
rect 4170 8222 4189 8228
rect 4204 8222 4234 8230
rect 4170 8214 4234 8222
rect 4170 8198 4250 8214
rect 4266 8207 4328 8238
rect 4344 8207 4406 8238
rect 4475 8236 4524 8261
rect 4539 8236 4569 8252
rect 4438 8222 4468 8230
rect 4475 8228 4585 8236
rect 4438 8214 4483 8222
rect 4170 8196 4189 8198
rect 4204 8196 4250 8198
rect 4170 8180 4250 8196
rect 4277 8194 4312 8207
rect 4353 8204 4390 8207
rect 4353 8202 4395 8204
rect 4282 8191 4312 8194
rect 4291 8187 4298 8191
rect 4298 8186 4299 8187
rect 4257 8180 4267 8186
rect 4016 8172 4051 8180
rect 4016 8146 4017 8172
rect 4024 8146 4051 8172
rect 3959 8128 3989 8142
rect 4016 8138 4051 8146
rect 4053 8172 4094 8180
rect 4053 8146 4068 8172
rect 4075 8146 4094 8172
rect 4158 8168 4189 8180
rect 4204 8168 4307 8180
rect 4319 8170 4345 8196
rect 4360 8191 4390 8202
rect 4422 8198 4484 8214
rect 4422 8196 4468 8198
rect 4422 8180 4484 8196
rect 4496 8180 4502 8228
rect 4505 8220 4585 8228
rect 4505 8218 4524 8220
rect 4539 8218 4573 8220
rect 4505 8202 4585 8218
rect 4505 8180 4524 8202
rect 4539 8186 4569 8202
rect 4597 8196 4603 8270
rect 4606 8196 4625 8340
rect 4640 8196 4646 8340
rect 4655 8270 4668 8340
rect 4720 8336 4742 8340
rect 4713 8314 4742 8328
rect 4795 8314 4811 8328
rect 4849 8324 4855 8326
rect 4862 8324 4970 8340
rect 4977 8324 4983 8326
rect 4991 8324 5006 8340
rect 5072 8334 5091 8337
rect 4713 8312 4811 8314
rect 4838 8312 5006 8324
rect 5021 8314 5037 8328
rect 5072 8315 5094 8334
rect 5104 8328 5120 8329
rect 5103 8326 5120 8328
rect 5104 8321 5120 8326
rect 5094 8314 5100 8315
rect 5103 8314 5132 8321
rect 5021 8313 5132 8314
rect 5021 8312 5138 8313
rect 4697 8304 4748 8312
rect 4795 8304 4829 8312
rect 4697 8292 4722 8304
rect 4729 8292 4748 8304
rect 4802 8302 4829 8304
rect 4838 8302 5059 8312
rect 5094 8309 5100 8312
rect 4802 8298 5059 8302
rect 4697 8284 4748 8292
rect 4795 8284 5059 8298
rect 5103 8304 5138 8312
rect 4649 8236 4668 8270
rect 4713 8276 4742 8284
rect 4713 8270 4730 8276
rect 4713 8268 4747 8270
rect 4795 8268 4811 8284
rect 4812 8274 5020 8284
rect 5021 8274 5037 8284
rect 5085 8280 5100 8295
rect 5103 8292 5104 8304
rect 5111 8292 5138 8304
rect 5103 8284 5138 8292
rect 5103 8283 5132 8284
rect 4823 8270 5037 8274
rect 4838 8268 5037 8270
rect 5072 8270 5085 8280
rect 5103 8270 5120 8283
rect 5072 8268 5120 8270
rect 4714 8264 4747 8268
rect 4710 8262 4747 8264
rect 4710 8261 4777 8262
rect 4710 8256 4741 8261
rect 4747 8256 4777 8261
rect 4710 8252 4777 8256
rect 4683 8249 4777 8252
rect 4683 8242 4732 8249
rect 4683 8236 4713 8242
rect 4732 8237 4737 8242
rect 4649 8220 4729 8236
rect 4741 8228 4777 8249
rect 4838 8244 5027 8268
rect 5072 8267 5119 8268
rect 5085 8262 5119 8267
rect 4853 8241 5027 8244
rect 4846 8238 5027 8241
rect 5055 8261 5119 8262
rect 4649 8218 4668 8220
rect 4683 8218 4717 8220
rect 4649 8202 4729 8218
rect 4649 8196 4668 8202
rect 4365 8170 4468 8180
rect 4319 8168 4468 8170
rect 4489 8168 4524 8180
rect 4158 8166 4320 8168
rect 4170 8146 4189 8166
rect 4204 8164 4234 8166
rect 4053 8138 4094 8146
rect 4176 8142 4189 8146
rect 4241 8150 4320 8166
rect 4352 8166 4524 8168
rect 4352 8150 4431 8166
rect 4438 8164 4468 8166
rect 4016 8128 4045 8138
rect 4059 8128 4088 8138
rect 4103 8128 4133 8142
rect 4176 8128 4219 8142
rect 4241 8138 4431 8150
rect 4496 8146 4502 8166
rect 4226 8128 4256 8138
rect 4257 8128 4415 8138
rect 4419 8128 4449 8138
rect 4453 8128 4483 8142
rect 4511 8128 4524 8166
rect 4596 8180 4625 8196
rect 4639 8180 4668 8196
rect 4683 8186 4713 8202
rect 4741 8180 4747 8228
rect 4750 8222 4769 8228
rect 4784 8222 4814 8230
rect 4750 8214 4814 8222
rect 4750 8198 4830 8214
rect 4846 8207 4908 8238
rect 4924 8207 4986 8238
rect 5055 8236 5104 8261
rect 5119 8236 5149 8252
rect 5018 8222 5048 8230
rect 5055 8228 5165 8236
rect 5018 8214 5063 8222
rect 4750 8196 4769 8198
rect 4784 8196 4830 8198
rect 4750 8180 4830 8196
rect 4857 8194 4892 8207
rect 4933 8204 4970 8207
rect 4933 8202 4975 8204
rect 4862 8191 4892 8194
rect 4871 8187 4878 8191
rect 4878 8186 4879 8187
rect 4837 8180 4847 8186
rect 4596 8172 4631 8180
rect 4596 8146 4597 8172
rect 4604 8146 4631 8172
rect 4539 8128 4569 8142
rect 4596 8138 4631 8146
rect 4633 8172 4674 8180
rect 4633 8146 4648 8172
rect 4655 8146 4674 8172
rect 4738 8168 4769 8180
rect 4784 8168 4887 8180
rect 4899 8170 4925 8196
rect 4940 8191 4970 8202
rect 5002 8198 5064 8214
rect 5002 8196 5048 8198
rect 5002 8180 5064 8196
rect 5076 8180 5082 8228
rect 5085 8220 5165 8228
rect 5085 8218 5104 8220
rect 5119 8218 5153 8220
rect 5085 8202 5165 8218
rect 5085 8180 5104 8202
rect 5119 8186 5149 8202
rect 5177 8196 5183 8270
rect 5186 8196 5205 8340
rect 5220 8196 5226 8340
rect 5235 8270 5248 8340
rect 5300 8336 5322 8340
rect 5293 8314 5322 8328
rect 5375 8314 5391 8328
rect 5429 8324 5435 8326
rect 5442 8324 5550 8340
rect 5557 8324 5563 8326
rect 5571 8324 5586 8340
rect 5652 8334 5671 8337
rect 5293 8312 5391 8314
rect 5418 8312 5586 8324
rect 5601 8314 5617 8328
rect 5652 8315 5674 8334
rect 5684 8328 5700 8329
rect 5683 8326 5700 8328
rect 5684 8321 5700 8326
rect 5674 8314 5680 8315
rect 5683 8314 5712 8321
rect 5601 8313 5712 8314
rect 5601 8312 5718 8313
rect 5277 8304 5328 8312
rect 5375 8304 5409 8312
rect 5277 8292 5302 8304
rect 5309 8292 5328 8304
rect 5382 8302 5409 8304
rect 5418 8302 5639 8312
rect 5674 8309 5680 8312
rect 5382 8298 5639 8302
rect 5277 8284 5328 8292
rect 5375 8284 5639 8298
rect 5683 8304 5718 8312
rect 5229 8236 5248 8270
rect 5293 8276 5322 8284
rect 5293 8270 5310 8276
rect 5293 8268 5327 8270
rect 5375 8268 5391 8284
rect 5392 8274 5600 8284
rect 5601 8274 5617 8284
rect 5665 8280 5680 8295
rect 5683 8292 5684 8304
rect 5691 8292 5718 8304
rect 5683 8284 5718 8292
rect 5683 8283 5712 8284
rect 5403 8270 5617 8274
rect 5418 8268 5617 8270
rect 5652 8270 5665 8280
rect 5683 8270 5700 8283
rect 5652 8268 5700 8270
rect 5294 8264 5327 8268
rect 5290 8262 5327 8264
rect 5290 8261 5357 8262
rect 5290 8256 5321 8261
rect 5327 8256 5357 8261
rect 5290 8252 5357 8256
rect 5263 8249 5357 8252
rect 5263 8242 5312 8249
rect 5263 8236 5293 8242
rect 5312 8237 5317 8242
rect 5229 8220 5309 8236
rect 5321 8228 5357 8249
rect 5418 8244 5607 8268
rect 5652 8267 5699 8268
rect 5665 8262 5699 8267
rect 5433 8241 5607 8244
rect 5426 8238 5607 8241
rect 5635 8261 5699 8262
rect 5229 8218 5248 8220
rect 5263 8218 5297 8220
rect 5229 8202 5309 8218
rect 5229 8196 5248 8202
rect 4945 8170 5048 8180
rect 4899 8168 5048 8170
rect 5069 8168 5104 8180
rect 4738 8166 4900 8168
rect 4750 8146 4769 8166
rect 4784 8164 4814 8166
rect 4633 8138 4674 8146
rect 4756 8142 4769 8146
rect 4821 8150 4900 8166
rect 4932 8166 5104 8168
rect 4932 8150 5011 8166
rect 5018 8164 5048 8166
rect 4596 8128 4625 8138
rect 4639 8128 4668 8138
rect 4683 8128 4713 8142
rect 4756 8128 4799 8142
rect 4821 8138 5011 8150
rect 5076 8146 5082 8166
rect 4806 8128 4836 8138
rect 4837 8128 4995 8138
rect 4999 8128 5029 8138
rect 5033 8128 5063 8142
rect 5091 8128 5104 8166
rect 5176 8180 5205 8196
rect 5219 8180 5248 8196
rect 5263 8186 5293 8202
rect 5321 8180 5327 8228
rect 5330 8222 5349 8228
rect 5364 8222 5394 8230
rect 5330 8214 5394 8222
rect 5330 8198 5410 8214
rect 5426 8207 5488 8238
rect 5504 8207 5566 8238
rect 5635 8236 5684 8261
rect 5699 8236 5729 8252
rect 5598 8222 5628 8230
rect 5635 8228 5745 8236
rect 5598 8214 5643 8222
rect 5330 8196 5349 8198
rect 5364 8196 5410 8198
rect 5330 8180 5410 8196
rect 5437 8194 5472 8207
rect 5513 8204 5550 8207
rect 5513 8202 5555 8204
rect 5442 8191 5472 8194
rect 5451 8187 5458 8191
rect 5458 8186 5459 8187
rect 5417 8180 5427 8186
rect 5176 8172 5211 8180
rect 5176 8146 5177 8172
rect 5184 8146 5211 8172
rect 5119 8128 5149 8142
rect 5176 8138 5211 8146
rect 5213 8172 5254 8180
rect 5213 8146 5228 8172
rect 5235 8146 5254 8172
rect 5318 8168 5349 8180
rect 5364 8168 5467 8180
rect 5479 8170 5505 8196
rect 5520 8191 5550 8202
rect 5582 8198 5644 8214
rect 5582 8196 5628 8198
rect 5582 8180 5644 8196
rect 5656 8180 5662 8228
rect 5665 8220 5745 8228
rect 5665 8218 5684 8220
rect 5699 8218 5733 8220
rect 5665 8202 5745 8218
rect 5665 8180 5684 8202
rect 5699 8186 5729 8202
rect 5757 8196 5763 8270
rect 5766 8196 5785 8340
rect 5800 8196 5806 8340
rect 5815 8270 5828 8340
rect 5880 8336 5902 8340
rect 5873 8314 5902 8328
rect 5955 8314 5971 8328
rect 6009 8324 6015 8326
rect 6022 8324 6130 8340
rect 6137 8324 6143 8326
rect 6151 8324 6166 8340
rect 6232 8334 6251 8337
rect 5873 8312 5971 8314
rect 5998 8312 6166 8324
rect 6181 8314 6197 8328
rect 6232 8315 6254 8334
rect 6264 8328 6280 8329
rect 6263 8326 6280 8328
rect 6264 8321 6280 8326
rect 6254 8314 6260 8315
rect 6263 8314 6292 8321
rect 6181 8313 6292 8314
rect 6181 8312 6298 8313
rect 5857 8304 5908 8312
rect 5955 8304 5989 8312
rect 5857 8292 5882 8304
rect 5889 8292 5908 8304
rect 5962 8302 5989 8304
rect 5998 8302 6219 8312
rect 6254 8309 6260 8312
rect 5962 8298 6219 8302
rect 5857 8284 5908 8292
rect 5955 8284 6219 8298
rect 6263 8304 6298 8312
rect 5809 8236 5828 8270
rect 5873 8276 5902 8284
rect 5873 8270 5890 8276
rect 5873 8268 5907 8270
rect 5955 8268 5971 8284
rect 5972 8274 6180 8284
rect 6181 8274 6197 8284
rect 6245 8280 6260 8295
rect 6263 8292 6264 8304
rect 6271 8292 6298 8304
rect 6263 8284 6298 8292
rect 6263 8283 6292 8284
rect 5983 8270 6197 8274
rect 5998 8268 6197 8270
rect 6232 8270 6245 8280
rect 6263 8270 6280 8283
rect 6232 8268 6280 8270
rect 5874 8264 5907 8268
rect 5870 8262 5907 8264
rect 5870 8261 5937 8262
rect 5870 8256 5901 8261
rect 5907 8256 5937 8261
rect 5870 8252 5937 8256
rect 5843 8249 5937 8252
rect 5843 8242 5892 8249
rect 5843 8236 5873 8242
rect 5892 8237 5897 8242
rect 5809 8220 5889 8236
rect 5901 8228 5937 8249
rect 5998 8244 6187 8268
rect 6232 8267 6279 8268
rect 6245 8262 6279 8267
rect 6013 8241 6187 8244
rect 6006 8238 6187 8241
rect 6215 8261 6279 8262
rect 5809 8218 5828 8220
rect 5843 8218 5877 8220
rect 5809 8202 5889 8218
rect 5809 8196 5828 8202
rect 5525 8170 5628 8180
rect 5479 8168 5628 8170
rect 5649 8168 5684 8180
rect 5318 8166 5480 8168
rect 5330 8146 5349 8166
rect 5364 8164 5394 8166
rect 5213 8138 5254 8146
rect 5336 8142 5349 8146
rect 5401 8150 5480 8166
rect 5512 8166 5684 8168
rect 5512 8150 5591 8166
rect 5598 8164 5628 8166
rect 5176 8128 5205 8138
rect 5219 8128 5248 8138
rect 5263 8128 5293 8142
rect 5336 8128 5379 8142
rect 5401 8138 5591 8150
rect 5656 8146 5662 8166
rect 5386 8128 5416 8138
rect 5417 8128 5575 8138
rect 5579 8128 5609 8138
rect 5613 8128 5643 8142
rect 5671 8128 5684 8166
rect 5756 8180 5785 8196
rect 5799 8180 5828 8196
rect 5843 8186 5873 8202
rect 5901 8180 5907 8228
rect 5910 8222 5929 8228
rect 5944 8222 5974 8230
rect 5910 8214 5974 8222
rect 5910 8198 5990 8214
rect 6006 8207 6068 8238
rect 6084 8207 6146 8238
rect 6215 8236 6264 8261
rect 6279 8236 6309 8252
rect 6178 8222 6208 8230
rect 6215 8228 6325 8236
rect 6178 8214 6223 8222
rect 5910 8196 5929 8198
rect 5944 8196 5990 8198
rect 5910 8180 5990 8196
rect 6017 8194 6052 8207
rect 6093 8204 6130 8207
rect 6093 8202 6135 8204
rect 6022 8191 6052 8194
rect 6031 8187 6038 8191
rect 6038 8186 6039 8187
rect 5997 8180 6007 8186
rect 5756 8172 5791 8180
rect 5756 8146 5757 8172
rect 5764 8146 5791 8172
rect 5699 8128 5729 8142
rect 5756 8138 5791 8146
rect 5793 8172 5834 8180
rect 5793 8146 5808 8172
rect 5815 8146 5834 8172
rect 5898 8168 5929 8180
rect 5944 8168 6047 8180
rect 6059 8170 6085 8196
rect 6100 8191 6130 8202
rect 6162 8198 6224 8214
rect 6162 8196 6208 8198
rect 6162 8180 6224 8196
rect 6236 8180 6242 8228
rect 6245 8220 6325 8228
rect 6245 8218 6264 8220
rect 6279 8218 6313 8220
rect 6245 8202 6325 8218
rect 6245 8180 6264 8202
rect 6279 8186 6309 8202
rect 6337 8196 6343 8270
rect 6346 8196 6365 8340
rect 6380 8196 6386 8340
rect 6395 8270 6408 8340
rect 6460 8336 6482 8340
rect 6453 8314 6482 8328
rect 6535 8314 6551 8328
rect 6589 8324 6595 8326
rect 6602 8324 6710 8340
rect 6717 8324 6723 8326
rect 6731 8324 6746 8340
rect 6812 8334 6831 8337
rect 6453 8312 6551 8314
rect 6578 8312 6746 8324
rect 6761 8314 6777 8328
rect 6812 8315 6834 8334
rect 6844 8328 6860 8329
rect 6843 8326 6860 8328
rect 6844 8321 6860 8326
rect 6834 8314 6840 8315
rect 6843 8314 6872 8321
rect 6761 8313 6872 8314
rect 6761 8312 6878 8313
rect 6437 8304 6488 8312
rect 6535 8304 6569 8312
rect 6437 8292 6462 8304
rect 6469 8292 6488 8304
rect 6542 8302 6569 8304
rect 6578 8302 6799 8312
rect 6834 8309 6840 8312
rect 6542 8298 6799 8302
rect 6437 8284 6488 8292
rect 6535 8284 6799 8298
rect 6843 8304 6878 8312
rect 6389 8236 6408 8270
rect 6453 8276 6482 8284
rect 6453 8270 6470 8276
rect 6453 8268 6487 8270
rect 6535 8268 6551 8284
rect 6552 8274 6760 8284
rect 6761 8274 6777 8284
rect 6825 8280 6840 8295
rect 6843 8292 6844 8304
rect 6851 8292 6878 8304
rect 6843 8284 6878 8292
rect 6843 8283 6872 8284
rect 6563 8270 6777 8274
rect 6578 8268 6777 8270
rect 6812 8270 6825 8280
rect 6843 8270 6860 8283
rect 6812 8268 6860 8270
rect 6454 8264 6487 8268
rect 6450 8262 6487 8264
rect 6450 8261 6517 8262
rect 6450 8256 6481 8261
rect 6487 8256 6517 8261
rect 6450 8252 6517 8256
rect 6423 8249 6517 8252
rect 6423 8242 6472 8249
rect 6423 8236 6453 8242
rect 6472 8237 6477 8242
rect 6389 8220 6469 8236
rect 6481 8228 6517 8249
rect 6578 8244 6767 8268
rect 6812 8267 6859 8268
rect 6825 8262 6859 8267
rect 6593 8241 6767 8244
rect 6586 8238 6767 8241
rect 6795 8261 6859 8262
rect 6389 8218 6408 8220
rect 6423 8218 6457 8220
rect 6389 8202 6469 8218
rect 6389 8196 6408 8202
rect 6105 8170 6208 8180
rect 6059 8168 6208 8170
rect 6229 8168 6264 8180
rect 5898 8166 6060 8168
rect 5910 8146 5929 8166
rect 5944 8164 5974 8166
rect 5793 8138 5834 8146
rect 5916 8142 5929 8146
rect 5981 8150 6060 8166
rect 6092 8166 6264 8168
rect 6092 8150 6171 8166
rect 6178 8164 6208 8166
rect 5756 8128 5785 8138
rect 5799 8128 5828 8138
rect 5843 8128 5873 8142
rect 5916 8128 5959 8142
rect 5981 8138 6171 8150
rect 6236 8146 6242 8166
rect 5966 8128 5996 8138
rect 5997 8128 6155 8138
rect 6159 8128 6189 8138
rect 6193 8128 6223 8142
rect 6251 8128 6264 8166
rect 6336 8180 6365 8196
rect 6379 8180 6408 8196
rect 6423 8186 6453 8202
rect 6481 8180 6487 8228
rect 6490 8222 6509 8228
rect 6524 8222 6554 8230
rect 6490 8214 6554 8222
rect 6490 8198 6570 8214
rect 6586 8207 6648 8238
rect 6664 8207 6726 8238
rect 6795 8236 6844 8261
rect 6859 8236 6889 8252
rect 6758 8222 6788 8230
rect 6795 8228 6905 8236
rect 6758 8214 6803 8222
rect 6490 8196 6509 8198
rect 6524 8196 6570 8198
rect 6490 8180 6570 8196
rect 6597 8194 6632 8207
rect 6673 8204 6710 8207
rect 6673 8202 6715 8204
rect 6602 8191 6632 8194
rect 6611 8187 6618 8191
rect 6618 8186 6619 8187
rect 6577 8180 6587 8186
rect 6336 8172 6371 8180
rect 6336 8146 6337 8172
rect 6344 8146 6371 8172
rect 6279 8128 6309 8142
rect 6336 8138 6371 8146
rect 6373 8172 6414 8180
rect 6373 8146 6388 8172
rect 6395 8146 6414 8172
rect 6478 8168 6509 8180
rect 6524 8168 6627 8180
rect 6639 8170 6665 8196
rect 6680 8191 6710 8202
rect 6742 8198 6804 8214
rect 6742 8196 6788 8198
rect 6742 8180 6804 8196
rect 6816 8180 6822 8228
rect 6825 8220 6905 8228
rect 6825 8218 6844 8220
rect 6859 8218 6893 8220
rect 6825 8202 6905 8218
rect 6825 8180 6844 8202
rect 6859 8186 6889 8202
rect 6917 8196 6923 8270
rect 6926 8196 6945 8340
rect 6960 8196 6966 8340
rect 6975 8270 6988 8340
rect 7040 8336 7062 8340
rect 7033 8314 7062 8328
rect 7115 8314 7131 8328
rect 7169 8324 7175 8326
rect 7182 8324 7290 8340
rect 7297 8324 7303 8326
rect 7311 8324 7326 8340
rect 7392 8334 7411 8337
rect 7033 8312 7131 8314
rect 7158 8312 7326 8324
rect 7341 8314 7357 8328
rect 7392 8315 7414 8334
rect 7424 8328 7440 8329
rect 7423 8326 7440 8328
rect 7424 8321 7440 8326
rect 7414 8314 7420 8315
rect 7423 8314 7452 8321
rect 7341 8313 7452 8314
rect 7341 8312 7458 8313
rect 7017 8304 7068 8312
rect 7115 8304 7149 8312
rect 7017 8292 7042 8304
rect 7049 8292 7068 8304
rect 7122 8302 7149 8304
rect 7158 8302 7379 8312
rect 7414 8309 7420 8312
rect 7122 8298 7379 8302
rect 7017 8284 7068 8292
rect 7115 8284 7379 8298
rect 7423 8304 7458 8312
rect 6969 8236 6988 8270
rect 7033 8276 7062 8284
rect 7033 8270 7050 8276
rect 7033 8268 7067 8270
rect 7115 8268 7131 8284
rect 7132 8274 7340 8284
rect 7341 8274 7357 8284
rect 7405 8280 7420 8295
rect 7423 8292 7424 8304
rect 7431 8292 7458 8304
rect 7423 8284 7458 8292
rect 7423 8283 7452 8284
rect 7143 8270 7357 8274
rect 7158 8268 7357 8270
rect 7392 8270 7405 8280
rect 7423 8270 7440 8283
rect 7392 8268 7440 8270
rect 7034 8264 7067 8268
rect 7030 8262 7067 8264
rect 7030 8261 7097 8262
rect 7030 8256 7061 8261
rect 7067 8256 7097 8261
rect 7030 8252 7097 8256
rect 7003 8249 7097 8252
rect 7003 8242 7052 8249
rect 7003 8236 7033 8242
rect 7052 8237 7057 8242
rect 6969 8220 7049 8236
rect 7061 8228 7097 8249
rect 7158 8244 7347 8268
rect 7392 8267 7439 8268
rect 7405 8262 7439 8267
rect 7173 8241 7347 8244
rect 7166 8238 7347 8241
rect 7375 8261 7439 8262
rect 6969 8218 6988 8220
rect 7003 8218 7037 8220
rect 6969 8202 7049 8218
rect 6969 8196 6988 8202
rect 6685 8170 6788 8180
rect 6639 8168 6788 8170
rect 6809 8168 6844 8180
rect 6478 8166 6640 8168
rect 6490 8146 6509 8166
rect 6524 8164 6554 8166
rect 6373 8138 6414 8146
rect 6496 8142 6509 8146
rect 6561 8150 6640 8166
rect 6672 8166 6844 8168
rect 6672 8150 6751 8166
rect 6758 8164 6788 8166
rect 6336 8128 6365 8138
rect 6379 8128 6408 8138
rect 6423 8128 6453 8142
rect 6496 8128 6539 8142
rect 6561 8138 6751 8150
rect 6816 8146 6822 8166
rect 6546 8128 6576 8138
rect 6577 8128 6735 8138
rect 6739 8128 6769 8138
rect 6773 8128 6803 8142
rect 6831 8128 6844 8166
rect 6916 8180 6945 8196
rect 6959 8180 6988 8196
rect 7003 8186 7033 8202
rect 7061 8180 7067 8228
rect 7070 8222 7089 8228
rect 7104 8222 7134 8230
rect 7070 8214 7134 8222
rect 7070 8198 7150 8214
rect 7166 8207 7228 8238
rect 7244 8207 7306 8238
rect 7375 8236 7424 8261
rect 7439 8236 7469 8252
rect 7338 8222 7368 8230
rect 7375 8228 7485 8236
rect 7338 8214 7383 8222
rect 7070 8196 7089 8198
rect 7104 8196 7150 8198
rect 7070 8180 7150 8196
rect 7177 8194 7212 8207
rect 7253 8204 7290 8207
rect 7253 8202 7295 8204
rect 7182 8191 7212 8194
rect 7191 8187 7198 8191
rect 7198 8186 7199 8187
rect 7157 8180 7167 8186
rect 6916 8172 6951 8180
rect 6916 8146 6917 8172
rect 6924 8146 6951 8172
rect 6859 8128 6889 8142
rect 6916 8138 6951 8146
rect 6953 8172 6994 8180
rect 6953 8146 6968 8172
rect 6975 8146 6994 8172
rect 7058 8168 7089 8180
rect 7104 8168 7207 8180
rect 7219 8170 7245 8196
rect 7260 8191 7290 8202
rect 7322 8198 7384 8214
rect 7322 8196 7368 8198
rect 7322 8180 7384 8196
rect 7396 8180 7402 8228
rect 7405 8220 7485 8228
rect 7405 8218 7424 8220
rect 7439 8218 7473 8220
rect 7405 8202 7485 8218
rect 7405 8180 7424 8202
rect 7439 8186 7469 8202
rect 7497 8196 7503 8270
rect 7506 8196 7525 8340
rect 7540 8196 7546 8340
rect 7555 8270 7568 8340
rect 7613 8318 7614 8328
rect 7629 8318 7642 8328
rect 7613 8314 7642 8318
rect 7647 8314 7677 8340
rect 7695 8326 7711 8328
rect 7783 8326 7836 8340
rect 7784 8324 7848 8326
rect 7891 8324 7906 8340
rect 7955 8337 7985 8340
rect 7955 8334 7991 8337
rect 7921 8326 7937 8328
rect 7695 8314 7710 8318
rect 7613 8312 7710 8314
rect 7738 8312 7906 8324
rect 7922 8314 7937 8318
rect 7955 8315 7994 8334
rect 8013 8328 8020 8329
rect 8019 8321 8020 8328
rect 8003 8318 8004 8321
rect 8019 8318 8032 8321
rect 7955 8314 7985 8315
rect 7994 8314 8000 8315
rect 8003 8314 8032 8318
rect 7922 8313 8032 8314
rect 7922 8312 8038 8313
rect 7597 8304 7648 8312
rect 7597 8292 7622 8304
rect 7629 8292 7648 8304
rect 7679 8304 7729 8312
rect 7679 8296 7695 8304
rect 7702 8302 7729 8304
rect 7738 8302 7959 8312
rect 7702 8292 7959 8302
rect 7988 8304 8038 8312
rect 7988 8295 8004 8304
rect 7597 8284 7648 8292
rect 7695 8284 7959 8292
rect 7985 8292 8004 8295
rect 8011 8292 8038 8304
rect 7985 8284 8038 8292
rect 7549 8236 7568 8270
rect 7613 8276 7614 8284
rect 7629 8276 7642 8284
rect 7613 8268 7629 8276
rect 7610 8261 7629 8264
rect 7610 8252 7632 8261
rect 7583 8242 7632 8252
rect 7583 8236 7613 8242
rect 7632 8237 7637 8242
rect 7549 8220 7629 8236
rect 7647 8228 7677 8284
rect 7712 8274 7920 8284
rect 7955 8280 8000 8284
rect 8003 8283 8004 8284
rect 8019 8283 8032 8284
rect 7738 8244 7927 8274
rect 7753 8241 7927 8244
rect 7746 8238 7927 8241
rect 7549 8218 7568 8220
rect 7583 8218 7617 8220
rect 7549 8202 7629 8218
rect 7656 8214 7669 8228
rect 7684 8214 7700 8230
rect 7746 8225 7757 8238
rect 7549 8196 7568 8202
rect 7265 8170 7368 8180
rect 7219 8168 7368 8170
rect 7389 8168 7424 8180
rect 7058 8166 7220 8168
rect 7070 8146 7089 8166
rect 7104 8164 7134 8166
rect 6953 8138 6994 8146
rect 7076 8142 7089 8146
rect 7141 8150 7220 8166
rect 7252 8166 7424 8168
rect 7252 8150 7331 8166
rect 7338 8164 7368 8166
rect 6916 8128 6945 8138
rect 6959 8128 6988 8138
rect 7003 8128 7033 8142
rect 7076 8128 7119 8142
rect 7141 8138 7331 8150
rect 7396 8146 7402 8166
rect 7126 8128 7156 8138
rect 7157 8128 7315 8138
rect 7319 8128 7349 8138
rect 7353 8128 7383 8142
rect 7411 8128 7424 8166
rect 7496 8180 7525 8196
rect 7539 8180 7568 8196
rect 7583 8180 7613 8202
rect 7656 8198 7718 8214
rect 7746 8207 7757 8223
rect 7762 8218 7772 8238
rect 7782 8218 7796 8238
rect 7799 8225 7808 8238
rect 7824 8225 7833 8238
rect 7762 8207 7796 8218
rect 7799 8207 7808 8223
rect 7824 8207 7833 8223
rect 7840 8218 7850 8238
rect 7860 8218 7874 8238
rect 7875 8225 7886 8238
rect 7840 8207 7874 8218
rect 7875 8207 7886 8223
rect 7932 8214 7948 8230
rect 7955 8228 7985 8280
rect 8019 8276 8020 8283
rect 8004 8268 8020 8276
rect 7991 8236 8004 8255
rect 8019 8236 8049 8252
rect 7991 8220 8065 8236
rect 7991 8218 8004 8220
rect 8019 8218 8053 8220
rect 7656 8196 7669 8198
rect 7684 8196 7718 8198
rect 7656 8180 7718 8196
rect 7762 8191 7778 8194
rect 7840 8191 7870 8202
rect 7918 8198 7964 8214
rect 7991 8202 8065 8218
rect 7918 8196 7952 8198
rect 7917 8180 7964 8196
rect 7991 8180 8004 8202
rect 8019 8180 8049 8202
rect 8076 8180 8077 8196
rect 8092 8180 8105 8340
rect 8135 8236 8148 8340
rect 8193 8318 8194 8328
rect 8209 8318 8222 8328
rect 8193 8314 8222 8318
rect 8227 8314 8257 8340
rect 8275 8326 8291 8328
rect 8363 8326 8416 8340
rect 8364 8324 8428 8326
rect 8471 8324 8486 8340
rect 8535 8337 8565 8340
rect 8535 8334 8571 8337
rect 8501 8326 8517 8328
rect 8275 8314 8290 8318
rect 8193 8312 8290 8314
rect 8318 8312 8486 8324
rect 8502 8314 8517 8318
rect 8535 8315 8574 8334
rect 8593 8328 8600 8329
rect 8599 8321 8600 8328
rect 8583 8318 8584 8321
rect 8599 8318 8612 8321
rect 8535 8314 8565 8315
rect 8574 8314 8580 8315
rect 8583 8314 8612 8318
rect 8502 8313 8612 8314
rect 8502 8312 8618 8313
rect 8177 8304 8228 8312
rect 8177 8292 8202 8304
rect 8209 8292 8228 8304
rect 8259 8304 8309 8312
rect 8259 8296 8275 8304
rect 8282 8302 8309 8304
rect 8318 8302 8539 8312
rect 8282 8292 8539 8302
rect 8568 8304 8618 8312
rect 8568 8295 8584 8304
rect 8177 8284 8228 8292
rect 8275 8284 8539 8292
rect 8565 8292 8584 8295
rect 8591 8292 8618 8304
rect 8565 8284 8618 8292
rect 8193 8276 8194 8284
rect 8209 8276 8222 8284
rect 8193 8268 8209 8276
rect 8190 8261 8209 8264
rect 8190 8252 8212 8261
rect 8163 8242 8212 8252
rect 8163 8236 8193 8242
rect 8212 8237 8217 8242
rect 8135 8220 8209 8236
rect 8227 8228 8257 8284
rect 8292 8274 8500 8284
rect 8535 8280 8580 8284
rect 8583 8283 8584 8284
rect 8599 8283 8612 8284
rect 8318 8244 8507 8274
rect 8333 8241 8507 8244
rect 8326 8238 8507 8241
rect 8135 8218 8148 8220
rect 8163 8218 8197 8220
rect 8135 8202 8209 8218
rect 8236 8214 8249 8228
rect 8264 8214 8280 8230
rect 8326 8225 8337 8238
rect 8119 8180 8120 8196
rect 8135 8180 8148 8202
rect 8163 8180 8193 8202
rect 8236 8198 8298 8214
rect 8326 8207 8337 8223
rect 8342 8218 8352 8238
rect 8362 8218 8376 8238
rect 8379 8225 8388 8238
rect 8404 8225 8413 8238
rect 8342 8207 8376 8218
rect 8379 8207 8388 8223
rect 8404 8207 8413 8223
rect 8420 8218 8430 8238
rect 8440 8218 8454 8238
rect 8455 8225 8466 8238
rect 8420 8207 8454 8218
rect 8455 8207 8466 8223
rect 8512 8214 8528 8230
rect 8535 8228 8565 8280
rect 8599 8276 8600 8283
rect 8584 8268 8600 8276
rect 8571 8236 8584 8255
rect 8599 8236 8629 8252
rect 8571 8220 8645 8236
rect 8571 8218 8584 8220
rect 8599 8218 8633 8220
rect 8236 8196 8249 8198
rect 8264 8196 8298 8198
rect 8236 8180 8298 8196
rect 8342 8191 8358 8194
rect 8420 8191 8450 8202
rect 8498 8198 8544 8214
rect 8571 8202 8645 8218
rect 8498 8196 8532 8198
rect 8497 8180 8544 8196
rect 8571 8180 8584 8202
rect 8599 8180 8629 8202
rect 8656 8180 8657 8196
rect 8672 8180 8685 8340
rect 8715 8236 8728 8340
rect 8773 8318 8774 8328
rect 8789 8318 8802 8328
rect 8773 8314 8802 8318
rect 8807 8314 8837 8340
rect 8855 8326 8871 8328
rect 8943 8326 8996 8340
rect 8944 8324 9008 8326
rect 9051 8324 9066 8340
rect 9115 8337 9145 8340
rect 9115 8334 9151 8337
rect 9081 8326 9097 8328
rect 8855 8314 8870 8318
rect 8773 8312 8870 8314
rect 8898 8312 9066 8324
rect 9082 8314 9097 8318
rect 9115 8315 9154 8334
rect 9173 8328 9180 8329
rect 9179 8321 9180 8328
rect 9163 8318 9164 8321
rect 9179 8318 9192 8321
rect 9115 8314 9145 8315
rect 9154 8314 9160 8315
rect 9163 8314 9192 8318
rect 9082 8313 9192 8314
rect 9082 8312 9198 8313
rect 8757 8304 8808 8312
rect 8757 8292 8782 8304
rect 8789 8292 8808 8304
rect 8839 8304 8889 8312
rect 8839 8296 8855 8304
rect 8862 8302 8889 8304
rect 8898 8302 9119 8312
rect 8862 8292 9119 8302
rect 9148 8304 9198 8312
rect 9148 8295 9164 8304
rect 8757 8284 8808 8292
rect 8855 8284 9119 8292
rect 9145 8292 9164 8295
rect 9171 8292 9198 8304
rect 9145 8284 9198 8292
rect 8773 8276 8774 8284
rect 8789 8276 8802 8284
rect 8773 8268 8789 8276
rect 8770 8261 8789 8264
rect 8770 8252 8792 8261
rect 8743 8242 8792 8252
rect 8743 8236 8773 8242
rect 8792 8237 8797 8242
rect 8715 8220 8789 8236
rect 8807 8228 8837 8284
rect 8872 8274 9080 8284
rect 9115 8280 9160 8284
rect 9163 8283 9164 8284
rect 9179 8283 9192 8284
rect 8898 8244 9087 8274
rect 8913 8241 9087 8244
rect 8906 8238 9087 8241
rect 8715 8218 8728 8220
rect 8743 8218 8777 8220
rect 8715 8202 8789 8218
rect 8816 8214 8829 8228
rect 8844 8214 8860 8230
rect 8906 8225 8917 8238
rect 8699 8180 8700 8196
rect 8715 8180 8728 8202
rect 8743 8180 8773 8202
rect 8816 8198 8878 8214
rect 8906 8207 8917 8223
rect 8922 8218 8932 8238
rect 8942 8218 8956 8238
rect 8959 8225 8968 8238
rect 8984 8225 8993 8238
rect 8922 8207 8956 8218
rect 8959 8207 8968 8223
rect 8984 8207 8993 8223
rect 9000 8218 9010 8238
rect 9020 8218 9034 8238
rect 9035 8225 9046 8238
rect 9000 8207 9034 8218
rect 9035 8207 9046 8223
rect 9092 8214 9108 8230
rect 9115 8228 9145 8280
rect 9179 8276 9180 8283
rect 9164 8268 9180 8276
rect 9151 8236 9164 8255
rect 9179 8236 9209 8252
rect 9151 8220 9225 8236
rect 9151 8218 9164 8220
rect 9179 8218 9213 8220
rect 8816 8196 8829 8198
rect 8844 8196 8878 8198
rect 8816 8180 8878 8196
rect 8922 8191 8938 8194
rect 9000 8191 9030 8202
rect 9078 8198 9124 8214
rect 9151 8202 9225 8218
rect 9078 8196 9112 8198
rect 9077 8180 9124 8196
rect 9151 8180 9164 8202
rect 9179 8180 9209 8202
rect 9236 8180 9237 8196
rect 9252 8180 9265 8340
rect 7496 8172 7531 8180
rect 7496 8146 7497 8172
rect 7504 8146 7531 8172
rect 7439 8128 7469 8142
rect 7496 8138 7531 8146
rect 7533 8172 7574 8180
rect 7533 8146 7548 8172
rect 7555 8146 7574 8172
rect 7638 8168 7700 8180
rect 7712 8168 7787 8180
rect 7845 8168 7920 8180
rect 7932 8168 7963 8180
rect 7969 8168 8004 8180
rect 7638 8166 7800 8168
rect 7533 8138 7574 8146
rect 7656 8142 7669 8166
rect 7684 8164 7699 8166
rect 7496 8128 7525 8138
rect 7539 8128 7568 8138
rect 7583 8128 7613 8142
rect 7656 8128 7699 8142
rect 7723 8139 7730 8146
rect 7733 8142 7800 8166
rect 7832 8166 8004 8168
rect 7802 8144 7830 8148
rect 7832 8144 7912 8166
rect 7933 8164 7948 8166
rect 7802 8142 7912 8144
rect 7733 8138 7912 8142
rect 7706 8128 7736 8138
rect 7738 8128 7891 8138
rect 7899 8128 7929 8138
rect 7933 8128 7963 8142
rect 7991 8128 8004 8166
rect 8076 8172 8111 8180
rect 8076 8146 8077 8172
rect 8084 8146 8111 8172
rect 8019 8128 8049 8142
rect 8076 8138 8111 8146
rect 8113 8172 8154 8180
rect 8113 8146 8128 8172
rect 8135 8146 8154 8172
rect 8218 8168 8280 8180
rect 8292 8168 8367 8180
rect 8425 8168 8500 8180
rect 8512 8168 8543 8180
rect 8549 8168 8584 8180
rect 8218 8166 8380 8168
rect 8113 8138 8154 8146
rect 8236 8142 8249 8166
rect 8264 8164 8279 8166
rect 8076 8128 8077 8138
rect 8092 8128 8105 8138
rect 8119 8128 8120 8138
rect 8135 8128 8148 8138
rect 8163 8128 8193 8142
rect 8236 8128 8279 8142
rect 8303 8139 8310 8146
rect 8313 8142 8380 8166
rect 8412 8166 8584 8168
rect 8382 8144 8410 8148
rect 8412 8144 8492 8166
rect 8513 8164 8528 8166
rect 8382 8142 8492 8144
rect 8313 8138 8492 8142
rect 8286 8128 8316 8138
rect 8318 8128 8471 8138
rect 8479 8128 8509 8138
rect 8513 8128 8543 8142
rect 8571 8128 8584 8166
rect 8656 8172 8691 8180
rect 8656 8146 8657 8172
rect 8664 8146 8691 8172
rect 8599 8128 8629 8142
rect 8656 8138 8691 8146
rect 8693 8172 8734 8180
rect 8693 8146 8708 8172
rect 8715 8146 8734 8172
rect 8798 8168 8860 8180
rect 8872 8168 8947 8180
rect 9005 8168 9080 8180
rect 9092 8168 9123 8180
rect 9129 8168 9164 8180
rect 8798 8166 8960 8168
rect 8693 8138 8734 8146
rect 8816 8142 8829 8166
rect 8844 8164 8859 8166
rect 8656 8128 8657 8138
rect 8672 8128 8685 8138
rect 8699 8128 8700 8138
rect 8715 8128 8728 8138
rect 8743 8128 8773 8142
rect 8816 8128 8859 8142
rect 8883 8139 8890 8146
rect 8893 8142 8960 8166
rect 8992 8166 9164 8168
rect 8962 8144 8990 8148
rect 8992 8144 9072 8166
rect 9093 8164 9108 8166
rect 8962 8142 9072 8144
rect 8893 8138 9072 8142
rect 8866 8128 8896 8138
rect 8898 8128 9051 8138
rect 9059 8128 9089 8138
rect 9093 8128 9123 8142
rect 9151 8128 9164 8166
rect 9236 8172 9271 8180
rect 9236 8146 9237 8172
rect 9244 8146 9271 8172
rect 9179 8128 9209 8142
rect 9236 8138 9271 8146
rect 9236 8128 9237 8138
rect 9252 8128 9265 8138
rect -1 8122 9265 8128
rect 0 8114 9265 8122
rect 15 8084 28 8114
rect 43 8096 73 8114
rect 116 8100 130 8114
rect 166 8100 386 8114
rect 117 8098 130 8100
rect 83 8086 98 8098
rect 80 8084 102 8086
rect 107 8084 137 8098
rect 198 8096 351 8100
rect 180 8084 372 8096
rect 415 8084 445 8098
rect 451 8084 464 8114
rect 479 8096 509 8114
rect 552 8084 565 8114
rect 595 8084 608 8114
rect 623 8096 653 8114
rect 696 8100 710 8114
rect 746 8100 966 8114
rect 697 8098 710 8100
rect 663 8086 678 8098
rect 660 8084 682 8086
rect 687 8084 717 8098
rect 778 8096 931 8100
rect 760 8084 952 8096
rect 995 8084 1025 8098
rect 1031 8084 1044 8114
rect 1059 8096 1089 8114
rect 1132 8084 1145 8114
rect 1175 8084 1188 8114
rect 1203 8096 1233 8114
rect 1276 8100 1290 8114
rect 1326 8100 1546 8114
rect 1277 8098 1290 8100
rect 1243 8086 1258 8098
rect 1240 8084 1262 8086
rect 1267 8084 1297 8098
rect 1358 8096 1511 8100
rect 1340 8084 1532 8096
rect 1575 8084 1605 8098
rect 1611 8084 1624 8114
rect 1639 8096 1669 8114
rect 1712 8084 1725 8114
rect 1755 8084 1768 8114
rect 1783 8100 1813 8114
rect 1856 8100 1899 8114
rect 1906 8100 2126 8114
rect 2133 8100 2163 8114
rect 1823 8086 1838 8098
rect 1857 8086 1870 8100
rect 1938 8096 2091 8100
rect 1820 8084 1842 8086
rect 1920 8084 2112 8096
rect 2191 8084 2204 8114
rect 2219 8100 2249 8114
rect 2286 8084 2305 8114
rect 2320 8084 2326 8114
rect 2335 8084 2348 8114
rect 2363 8100 2393 8114
rect 2436 8100 2479 8114
rect 2486 8100 2706 8114
rect 2713 8100 2743 8114
rect 2403 8086 2418 8098
rect 2437 8086 2450 8100
rect 2518 8096 2671 8100
rect 2400 8084 2422 8086
rect 2500 8084 2692 8096
rect 2771 8084 2784 8114
rect 2799 8100 2829 8114
rect 2866 8084 2885 8114
rect 2900 8084 2906 8114
rect 2915 8084 2928 8114
rect 2943 8100 2973 8114
rect 3016 8100 3059 8114
rect 3066 8100 3286 8114
rect 3293 8100 3323 8114
rect 2983 8086 2998 8098
rect 3017 8086 3030 8100
rect 3098 8096 3251 8100
rect 2980 8084 3002 8086
rect 3080 8084 3272 8096
rect 3351 8084 3364 8114
rect 3379 8100 3409 8114
rect 3446 8084 3465 8114
rect 3480 8084 3486 8114
rect 3495 8084 3508 8114
rect 3523 8100 3553 8114
rect 3596 8100 3639 8114
rect 3646 8100 3866 8114
rect 3873 8100 3903 8114
rect 3563 8086 3578 8098
rect 3597 8086 3610 8100
rect 3678 8096 3831 8100
rect 3560 8084 3582 8086
rect 3660 8084 3852 8096
rect 3931 8084 3944 8114
rect 3959 8100 3989 8114
rect 4026 8084 4045 8114
rect 4060 8084 4066 8114
rect 4075 8084 4088 8114
rect 4103 8100 4133 8114
rect 4176 8100 4219 8114
rect 4226 8100 4446 8114
rect 4453 8100 4483 8114
rect 4143 8086 4158 8098
rect 4177 8086 4190 8100
rect 4258 8096 4411 8100
rect 4140 8084 4162 8086
rect 4240 8084 4432 8096
rect 4511 8084 4524 8114
rect 4539 8100 4569 8114
rect 4606 8084 4625 8114
rect 4640 8084 4646 8114
rect 4655 8084 4668 8114
rect 4683 8100 4713 8114
rect 4756 8100 4799 8114
rect 4806 8100 5026 8114
rect 5033 8100 5063 8114
rect 4723 8086 4738 8098
rect 4757 8086 4770 8100
rect 4838 8096 4991 8100
rect 4720 8084 4742 8086
rect 4820 8084 5012 8096
rect 5091 8084 5104 8114
rect 5119 8100 5149 8114
rect 5186 8084 5205 8114
rect 5220 8084 5226 8114
rect 5235 8084 5248 8114
rect 5263 8100 5293 8114
rect 5336 8100 5379 8114
rect 5386 8100 5606 8114
rect 5613 8100 5643 8114
rect 5303 8086 5318 8098
rect 5337 8086 5350 8100
rect 5418 8096 5571 8100
rect 5300 8084 5322 8086
rect 5400 8084 5592 8096
rect 5671 8084 5684 8114
rect 5699 8100 5729 8114
rect 5766 8084 5785 8114
rect 5800 8084 5806 8114
rect 5815 8084 5828 8114
rect 5843 8100 5873 8114
rect 5916 8100 5959 8114
rect 5966 8100 6186 8114
rect 6193 8100 6223 8114
rect 5883 8086 5898 8098
rect 5917 8086 5930 8100
rect 5998 8096 6151 8100
rect 5880 8084 5902 8086
rect 5980 8084 6172 8096
rect 6251 8084 6264 8114
rect 6279 8100 6309 8114
rect 6346 8084 6365 8114
rect 6380 8084 6386 8114
rect 6395 8084 6408 8114
rect 6423 8100 6453 8114
rect 6496 8100 6539 8114
rect 6546 8100 6766 8114
rect 6773 8100 6803 8114
rect 6463 8086 6478 8098
rect 6497 8086 6510 8100
rect 6578 8096 6731 8100
rect 6460 8084 6482 8086
rect 6560 8084 6752 8096
rect 6831 8084 6844 8114
rect 6859 8100 6889 8114
rect 6926 8084 6945 8114
rect 6960 8084 6966 8114
rect 6975 8084 6988 8114
rect 7003 8100 7033 8114
rect 7076 8100 7119 8114
rect 7126 8100 7346 8114
rect 7353 8100 7383 8114
rect 7043 8086 7058 8098
rect 7077 8086 7090 8100
rect 7158 8096 7311 8100
rect 7040 8084 7062 8086
rect 7140 8084 7332 8096
rect 7411 8084 7424 8114
rect 7439 8100 7469 8114
rect 7506 8084 7525 8114
rect 7540 8084 7546 8114
rect 7555 8084 7568 8114
rect 7583 8096 7613 8114
rect 7656 8100 7670 8114
rect 7706 8100 7926 8114
rect 7657 8098 7670 8100
rect 7623 8086 7638 8098
rect 7620 8084 7642 8086
rect 7647 8084 7677 8098
rect 7738 8096 7891 8100
rect 7720 8084 7912 8096
rect 7955 8084 7985 8098
rect 7991 8084 8004 8114
rect 8019 8096 8049 8114
rect 8092 8084 8105 8114
rect 8135 8084 8148 8114
rect 8163 8096 8193 8114
rect 8236 8100 8250 8114
rect 8286 8100 8506 8114
rect 8237 8098 8250 8100
rect 8203 8086 8218 8098
rect 8200 8084 8222 8086
rect 8227 8084 8257 8098
rect 8318 8096 8471 8100
rect 8300 8084 8492 8096
rect 8535 8084 8565 8098
rect 8571 8084 8584 8114
rect 8599 8096 8629 8114
rect 8672 8084 8685 8114
rect 8715 8084 8728 8114
rect 8743 8096 8773 8114
rect 8816 8100 8830 8114
rect 8866 8100 9086 8114
rect 8817 8098 8830 8100
rect 8783 8086 8798 8098
rect 8780 8084 8802 8086
rect 8807 8084 8837 8098
rect 8898 8096 9051 8100
rect 8880 8084 9072 8096
rect 9115 8084 9145 8098
rect 9151 8084 9164 8114
rect 9179 8096 9209 8114
rect 9252 8084 9265 8114
rect 0 8070 9265 8084
rect 15 7966 28 8070
rect 73 8048 74 8058
rect 89 8048 102 8058
rect 73 8044 102 8048
rect 107 8044 137 8070
rect 155 8056 171 8058
rect 243 8056 296 8070
rect 244 8054 308 8056
rect 351 8054 366 8070
rect 415 8067 445 8070
rect 415 8064 451 8067
rect 381 8056 397 8058
rect 155 8044 170 8048
rect 73 8042 170 8044
rect 198 8042 366 8054
rect 382 8044 397 8048
rect 415 8045 454 8064
rect 473 8058 480 8059
rect 479 8051 480 8058
rect 463 8048 464 8051
rect 479 8048 492 8051
rect 415 8044 445 8045
rect 454 8044 460 8045
rect 463 8044 492 8048
rect 382 8043 492 8044
rect 382 8042 498 8043
rect 57 8034 108 8042
rect 57 8022 82 8034
rect 89 8022 108 8034
rect 139 8034 189 8042
rect 139 8026 155 8034
rect 162 8032 189 8034
rect 198 8032 419 8042
rect 162 8022 419 8032
rect 448 8034 498 8042
rect 448 8025 464 8034
rect 57 8014 108 8022
rect 155 8014 419 8022
rect 445 8022 464 8025
rect 471 8022 498 8034
rect 445 8014 498 8022
rect 73 8006 74 8014
rect 89 8006 102 8014
rect 73 7998 89 8006
rect 70 7991 89 7994
rect 70 7982 92 7991
rect 43 7972 92 7982
rect 43 7966 73 7972
rect 92 7967 97 7972
rect 15 7950 89 7966
rect 107 7958 137 8014
rect 172 8004 380 8014
rect 415 8010 460 8014
rect 463 8013 464 8014
rect 479 8013 492 8014
rect 198 7974 387 8004
rect 213 7971 387 7974
rect 206 7968 387 7971
rect 15 7948 28 7950
rect 43 7948 77 7950
rect 15 7932 89 7948
rect 116 7944 129 7958
rect 144 7944 160 7960
rect 206 7955 217 7968
rect -1 7910 0 7926
rect 15 7910 28 7932
rect 43 7910 73 7932
rect 116 7928 178 7944
rect 206 7937 217 7953
rect 222 7948 232 7968
rect 242 7948 256 7968
rect 259 7955 268 7968
rect 284 7955 293 7968
rect 222 7937 256 7948
rect 259 7937 268 7953
rect 284 7937 293 7953
rect 300 7948 310 7968
rect 320 7948 334 7968
rect 335 7955 346 7968
rect 300 7937 334 7948
rect 335 7937 346 7953
rect 392 7944 408 7960
rect 415 7958 445 8010
rect 479 8006 480 8013
rect 464 7998 480 8006
rect 451 7966 464 7985
rect 479 7966 509 7982
rect 451 7950 525 7966
rect 451 7948 464 7950
rect 479 7948 513 7950
rect 116 7926 129 7928
rect 144 7926 178 7928
rect 116 7910 178 7926
rect 222 7921 238 7924
rect 300 7921 330 7932
rect 378 7928 424 7944
rect 451 7932 525 7948
rect 378 7926 412 7928
rect 377 7910 424 7926
rect 451 7910 464 7932
rect 479 7910 509 7932
rect 536 7910 537 7926
rect 552 7910 565 8070
rect 595 7966 608 8070
rect 653 8048 654 8058
rect 669 8048 682 8058
rect 653 8044 682 8048
rect 687 8044 717 8070
rect 735 8056 751 8058
rect 823 8056 876 8070
rect 824 8054 888 8056
rect 931 8054 946 8070
rect 995 8067 1025 8070
rect 995 8064 1031 8067
rect 961 8056 977 8058
rect 735 8044 750 8048
rect 653 8042 750 8044
rect 778 8042 946 8054
rect 962 8044 977 8048
rect 995 8045 1034 8064
rect 1053 8058 1060 8059
rect 1059 8051 1060 8058
rect 1043 8048 1044 8051
rect 1059 8048 1072 8051
rect 995 8044 1025 8045
rect 1034 8044 1040 8045
rect 1043 8044 1072 8048
rect 962 8043 1072 8044
rect 962 8042 1078 8043
rect 637 8034 688 8042
rect 637 8022 662 8034
rect 669 8022 688 8034
rect 719 8034 769 8042
rect 719 8026 735 8034
rect 742 8032 769 8034
rect 778 8032 999 8042
rect 742 8022 999 8032
rect 1028 8034 1078 8042
rect 1028 8025 1044 8034
rect 637 8014 688 8022
rect 735 8014 999 8022
rect 1025 8022 1044 8025
rect 1051 8022 1078 8034
rect 1025 8014 1078 8022
rect 653 8006 654 8014
rect 669 8006 682 8014
rect 653 7998 669 8006
rect 650 7991 669 7994
rect 650 7982 672 7991
rect 623 7972 672 7982
rect 623 7966 653 7972
rect 672 7967 677 7972
rect 595 7950 669 7966
rect 687 7958 717 8014
rect 752 8004 960 8014
rect 995 8010 1040 8014
rect 1043 8013 1044 8014
rect 1059 8013 1072 8014
rect 778 7974 967 8004
rect 793 7971 967 7974
rect 786 7968 967 7971
rect 595 7948 608 7950
rect 623 7948 657 7950
rect 595 7932 669 7948
rect 696 7944 709 7958
rect 724 7944 740 7960
rect 786 7955 797 7968
rect 579 7910 580 7926
rect 595 7910 608 7932
rect 623 7910 653 7932
rect 696 7928 758 7944
rect 786 7937 797 7953
rect 802 7948 812 7968
rect 822 7948 836 7968
rect 839 7955 848 7968
rect 864 7955 873 7968
rect 802 7937 836 7948
rect 839 7937 848 7953
rect 864 7937 873 7953
rect 880 7948 890 7968
rect 900 7948 914 7968
rect 915 7955 926 7968
rect 880 7937 914 7948
rect 915 7937 926 7953
rect 972 7944 988 7960
rect 995 7958 1025 8010
rect 1059 8006 1060 8013
rect 1044 7998 1060 8006
rect 1031 7966 1044 7985
rect 1059 7966 1089 7982
rect 1031 7950 1105 7966
rect 1031 7948 1044 7950
rect 1059 7948 1093 7950
rect 696 7926 709 7928
rect 724 7926 758 7928
rect 696 7910 758 7926
rect 802 7921 818 7924
rect 880 7921 910 7932
rect 958 7928 1004 7944
rect 1031 7932 1105 7948
rect 958 7926 992 7928
rect 957 7910 1004 7926
rect 1031 7910 1044 7932
rect 1059 7910 1089 7932
rect 1116 7910 1117 7926
rect 1132 7910 1145 8070
rect 1175 7966 1188 8070
rect 1233 8048 1234 8058
rect 1249 8048 1262 8058
rect 1233 8044 1262 8048
rect 1267 8044 1297 8070
rect 1315 8056 1331 8058
rect 1403 8056 1456 8070
rect 1404 8054 1468 8056
rect 1511 8054 1526 8070
rect 1575 8067 1605 8070
rect 1575 8064 1611 8067
rect 1541 8056 1557 8058
rect 1315 8044 1330 8048
rect 1233 8042 1330 8044
rect 1358 8042 1526 8054
rect 1542 8044 1557 8048
rect 1575 8045 1614 8064
rect 1633 8058 1640 8059
rect 1639 8051 1640 8058
rect 1623 8048 1624 8051
rect 1639 8048 1652 8051
rect 1575 8044 1605 8045
rect 1614 8044 1620 8045
rect 1623 8044 1652 8048
rect 1542 8043 1652 8044
rect 1542 8042 1658 8043
rect 1217 8034 1268 8042
rect 1217 8022 1242 8034
rect 1249 8022 1268 8034
rect 1299 8034 1349 8042
rect 1299 8026 1315 8034
rect 1322 8032 1349 8034
rect 1358 8032 1579 8042
rect 1322 8022 1579 8032
rect 1608 8034 1658 8042
rect 1608 8025 1624 8034
rect 1217 8014 1268 8022
rect 1315 8014 1579 8022
rect 1605 8022 1624 8025
rect 1631 8022 1658 8034
rect 1605 8014 1658 8022
rect 1233 8006 1234 8014
rect 1249 8006 1262 8014
rect 1233 7998 1249 8006
rect 1230 7991 1249 7994
rect 1230 7982 1252 7991
rect 1203 7972 1252 7982
rect 1203 7966 1233 7972
rect 1252 7967 1257 7972
rect 1175 7950 1249 7966
rect 1267 7958 1297 8014
rect 1332 8004 1540 8014
rect 1575 8010 1620 8014
rect 1623 8013 1624 8014
rect 1639 8013 1652 8014
rect 1358 7974 1547 8004
rect 1373 7971 1547 7974
rect 1366 7968 1547 7971
rect 1175 7948 1188 7950
rect 1203 7948 1237 7950
rect 1175 7932 1249 7948
rect 1276 7944 1289 7958
rect 1304 7944 1320 7960
rect 1366 7955 1377 7968
rect 1159 7910 1160 7926
rect 1175 7910 1188 7932
rect 1203 7910 1233 7932
rect 1276 7928 1338 7944
rect 1366 7937 1377 7953
rect 1382 7948 1392 7968
rect 1402 7948 1416 7968
rect 1419 7955 1428 7968
rect 1444 7955 1453 7968
rect 1382 7937 1416 7948
rect 1419 7937 1428 7953
rect 1444 7937 1453 7953
rect 1460 7948 1470 7968
rect 1480 7948 1494 7968
rect 1495 7955 1506 7968
rect 1460 7937 1494 7948
rect 1495 7937 1506 7953
rect 1552 7944 1568 7960
rect 1575 7958 1605 8010
rect 1639 8006 1640 8013
rect 1624 7998 1640 8006
rect 1611 7966 1624 7985
rect 1639 7966 1669 7982
rect 1611 7950 1685 7966
rect 1611 7948 1624 7950
rect 1639 7948 1673 7950
rect 1276 7926 1289 7928
rect 1304 7926 1338 7928
rect 1276 7910 1338 7926
rect 1382 7921 1398 7924
rect 1460 7921 1490 7932
rect 1538 7928 1584 7944
rect 1611 7932 1685 7948
rect 1538 7926 1572 7928
rect 1537 7910 1584 7926
rect 1611 7910 1624 7932
rect 1639 7910 1669 7932
rect 1696 7910 1697 7926
rect 1712 7910 1725 8070
rect 1755 7966 1768 8070
rect 1820 8066 1842 8070
rect 1813 8044 1842 8058
rect 1895 8044 1911 8058
rect 1949 8054 1955 8056
rect 1962 8054 2070 8070
rect 2077 8054 2083 8056
rect 2091 8054 2106 8070
rect 2172 8064 2191 8067
rect 1813 8042 1911 8044
rect 1938 8042 2106 8054
rect 2121 8044 2137 8058
rect 2172 8045 2194 8064
rect 2204 8058 2220 8059
rect 2203 8056 2220 8058
rect 2204 8051 2220 8056
rect 2194 8044 2200 8045
rect 2203 8044 2232 8051
rect 2121 8043 2232 8044
rect 2121 8042 2238 8043
rect 1797 8034 1848 8042
rect 1895 8034 1929 8042
rect 1797 8022 1822 8034
rect 1829 8022 1848 8034
rect 1902 8032 1929 8034
rect 1938 8032 2159 8042
rect 2194 8039 2200 8042
rect 1902 8028 2159 8032
rect 1797 8014 1848 8022
rect 1895 8014 2159 8028
rect 2203 8034 2238 8042
rect 1813 8006 1842 8014
rect 1813 8000 1830 8006
rect 1813 7998 1847 8000
rect 1895 7998 1911 8014
rect 1912 8004 2120 8014
rect 2121 8004 2137 8014
rect 2185 8010 2200 8025
rect 2203 8022 2204 8034
rect 2211 8022 2238 8034
rect 2203 8014 2238 8022
rect 2203 8013 2232 8014
rect 1923 8000 2137 8004
rect 1938 7998 2137 8000
rect 2172 8000 2185 8010
rect 2203 8000 2220 8013
rect 2172 7998 2220 8000
rect 1814 7994 1847 7998
rect 1810 7992 1847 7994
rect 1810 7991 1877 7992
rect 1810 7986 1841 7991
rect 1847 7986 1877 7991
rect 1810 7982 1877 7986
rect 1783 7979 1877 7982
rect 1783 7972 1832 7979
rect 1783 7966 1813 7972
rect 1832 7967 1837 7972
rect 1755 7950 1829 7966
rect 1841 7958 1877 7979
rect 1938 7974 2127 7998
rect 2172 7997 2219 7998
rect 2185 7992 2219 7997
rect 1953 7971 2127 7974
rect 1946 7968 2127 7971
rect 2155 7991 2219 7992
rect 1755 7948 1768 7950
rect 1783 7948 1817 7950
rect 1755 7932 1829 7948
rect 1739 7910 1740 7926
rect 1755 7910 1768 7932
rect 1783 7916 1813 7932
rect 1841 7910 1847 7958
rect 1850 7952 1869 7958
rect 1884 7952 1914 7960
rect 1850 7944 1914 7952
rect 1850 7928 1930 7944
rect 1946 7937 2008 7968
rect 2024 7937 2086 7968
rect 2155 7966 2204 7991
rect 2219 7966 2249 7982
rect 2118 7952 2148 7960
rect 2155 7958 2265 7966
rect 2118 7944 2163 7952
rect 1850 7926 1869 7928
rect 1884 7926 1930 7928
rect 1850 7910 1930 7926
rect 1957 7924 1992 7937
rect 2033 7934 2070 7937
rect 2033 7932 2075 7934
rect 1962 7921 1992 7924
rect 1971 7917 1978 7921
rect 1978 7916 1979 7917
rect 1937 7910 1947 7916
rect -7 7902 34 7910
rect -7 7876 8 7902
rect 15 7876 34 7902
rect 98 7898 160 7910
rect 172 7898 247 7910
rect 305 7898 380 7910
rect 392 7898 423 7910
rect 429 7898 464 7910
rect 98 7896 260 7898
rect -7 7868 34 7876
rect 116 7872 129 7896
rect 144 7894 159 7896
rect -1 7858 0 7868
rect 15 7858 28 7868
rect 43 7858 73 7872
rect 116 7858 159 7872
rect 183 7869 190 7876
rect 193 7872 260 7896
rect 292 7896 464 7898
rect 262 7874 290 7878
rect 292 7874 372 7896
rect 393 7894 408 7896
rect 262 7872 372 7874
rect 193 7868 372 7872
rect 166 7858 196 7868
rect 198 7858 351 7868
rect 359 7858 389 7868
rect 393 7858 423 7872
rect 451 7858 464 7896
rect 536 7902 571 7910
rect 536 7876 537 7902
rect 544 7876 571 7902
rect 479 7858 509 7872
rect 536 7868 571 7876
rect 573 7902 614 7910
rect 573 7876 588 7902
rect 595 7876 614 7902
rect 678 7898 740 7910
rect 752 7898 827 7910
rect 885 7898 960 7910
rect 972 7898 1003 7910
rect 1009 7898 1044 7910
rect 678 7896 840 7898
rect 573 7868 614 7876
rect 696 7872 709 7896
rect 724 7894 739 7896
rect 536 7858 537 7868
rect 552 7858 565 7868
rect 579 7858 580 7868
rect 595 7858 608 7868
rect 623 7858 653 7872
rect 696 7858 739 7872
rect 763 7869 770 7876
rect 773 7872 840 7896
rect 872 7896 1044 7898
rect 842 7874 870 7878
rect 872 7874 952 7896
rect 973 7894 988 7896
rect 842 7872 952 7874
rect 773 7868 952 7872
rect 746 7858 776 7868
rect 778 7858 931 7868
rect 939 7858 969 7868
rect 973 7858 1003 7872
rect 1031 7858 1044 7896
rect 1116 7902 1151 7910
rect 1116 7876 1117 7902
rect 1124 7876 1151 7902
rect 1059 7858 1089 7872
rect 1116 7868 1151 7876
rect 1153 7902 1194 7910
rect 1153 7876 1168 7902
rect 1175 7876 1194 7902
rect 1258 7898 1320 7910
rect 1332 7898 1407 7910
rect 1465 7898 1540 7910
rect 1552 7898 1583 7910
rect 1589 7898 1624 7910
rect 1258 7896 1420 7898
rect 1153 7868 1194 7876
rect 1276 7872 1289 7896
rect 1304 7894 1319 7896
rect 1116 7858 1117 7868
rect 1132 7858 1145 7868
rect 1159 7858 1160 7868
rect 1175 7858 1188 7868
rect 1203 7858 1233 7872
rect 1276 7858 1319 7872
rect 1343 7869 1350 7876
rect 1353 7872 1420 7896
rect 1452 7896 1624 7898
rect 1422 7874 1450 7878
rect 1452 7874 1532 7896
rect 1553 7894 1568 7896
rect 1422 7872 1532 7874
rect 1353 7868 1532 7872
rect 1326 7858 1356 7868
rect 1358 7858 1511 7868
rect 1519 7858 1549 7868
rect 1553 7858 1583 7872
rect 1611 7858 1624 7896
rect 1696 7902 1731 7910
rect 1696 7876 1697 7902
rect 1704 7876 1731 7902
rect 1639 7858 1669 7872
rect 1696 7868 1731 7876
rect 1733 7902 1774 7910
rect 1733 7876 1748 7902
rect 1755 7876 1774 7902
rect 1838 7898 1869 7910
rect 1884 7898 1987 7910
rect 1999 7900 2025 7926
rect 2040 7921 2070 7932
rect 2102 7928 2164 7944
rect 2102 7926 2148 7928
rect 2102 7910 2164 7926
rect 2176 7910 2182 7958
rect 2185 7950 2265 7958
rect 2185 7948 2204 7950
rect 2219 7948 2253 7950
rect 2185 7932 2265 7948
rect 2185 7910 2204 7932
rect 2219 7916 2249 7932
rect 2277 7926 2283 8000
rect 2286 7926 2305 8070
rect 2320 7926 2326 8070
rect 2335 8000 2348 8070
rect 2400 8066 2422 8070
rect 2393 8044 2422 8058
rect 2475 8044 2491 8058
rect 2529 8054 2535 8056
rect 2542 8054 2650 8070
rect 2657 8054 2663 8056
rect 2671 8054 2686 8070
rect 2752 8064 2771 8067
rect 2393 8042 2491 8044
rect 2518 8042 2686 8054
rect 2701 8044 2717 8058
rect 2752 8045 2774 8064
rect 2784 8058 2800 8059
rect 2783 8056 2800 8058
rect 2784 8051 2800 8056
rect 2774 8044 2780 8045
rect 2783 8044 2812 8051
rect 2701 8043 2812 8044
rect 2701 8042 2818 8043
rect 2377 8034 2428 8042
rect 2475 8034 2509 8042
rect 2377 8022 2402 8034
rect 2409 8022 2428 8034
rect 2482 8032 2509 8034
rect 2518 8032 2739 8042
rect 2774 8039 2780 8042
rect 2482 8028 2739 8032
rect 2377 8014 2428 8022
rect 2475 8014 2739 8028
rect 2783 8034 2818 8042
rect 2329 7966 2348 8000
rect 2393 8006 2422 8014
rect 2393 8000 2410 8006
rect 2393 7998 2427 8000
rect 2475 7998 2491 8014
rect 2492 8004 2700 8014
rect 2701 8004 2717 8014
rect 2765 8010 2780 8025
rect 2783 8022 2784 8034
rect 2791 8022 2818 8034
rect 2783 8014 2818 8022
rect 2783 8013 2812 8014
rect 2503 8000 2717 8004
rect 2518 7998 2717 8000
rect 2752 8000 2765 8010
rect 2783 8000 2800 8013
rect 2752 7998 2800 8000
rect 2394 7994 2427 7998
rect 2390 7992 2427 7994
rect 2390 7991 2457 7992
rect 2390 7986 2421 7991
rect 2427 7986 2457 7991
rect 2390 7982 2457 7986
rect 2363 7979 2457 7982
rect 2363 7972 2412 7979
rect 2363 7966 2393 7972
rect 2412 7967 2417 7972
rect 2329 7950 2409 7966
rect 2421 7958 2457 7979
rect 2518 7974 2707 7998
rect 2752 7997 2799 7998
rect 2765 7992 2799 7997
rect 2533 7971 2707 7974
rect 2526 7968 2707 7971
rect 2735 7991 2799 7992
rect 2329 7948 2348 7950
rect 2363 7948 2397 7950
rect 2329 7932 2409 7948
rect 2329 7926 2348 7932
rect 2045 7900 2148 7910
rect 1999 7898 2148 7900
rect 2169 7898 2204 7910
rect 1838 7896 2000 7898
rect 1850 7876 1869 7896
rect 1884 7894 1914 7896
rect 1733 7868 1774 7876
rect 1856 7872 1869 7876
rect 1921 7880 2000 7896
rect 2032 7896 2204 7898
rect 2032 7880 2111 7896
rect 2118 7894 2148 7896
rect 1696 7858 1697 7868
rect 1712 7858 1725 7868
rect 1739 7858 1740 7868
rect 1755 7858 1768 7868
rect 1783 7858 1813 7872
rect 1856 7858 1899 7872
rect 1921 7868 2111 7880
rect 2176 7876 2182 7896
rect 1906 7858 1936 7868
rect 1937 7858 2095 7868
rect 2099 7858 2129 7868
rect 2133 7858 2163 7872
rect 2191 7858 2204 7896
rect 2276 7910 2305 7926
rect 2319 7910 2348 7926
rect 2363 7916 2393 7932
rect 2421 7910 2427 7958
rect 2430 7952 2449 7958
rect 2464 7952 2494 7960
rect 2430 7944 2494 7952
rect 2430 7928 2510 7944
rect 2526 7937 2588 7968
rect 2604 7937 2666 7968
rect 2735 7966 2784 7991
rect 2799 7966 2829 7982
rect 2698 7952 2728 7960
rect 2735 7958 2845 7966
rect 2698 7944 2743 7952
rect 2430 7926 2449 7928
rect 2464 7926 2510 7928
rect 2430 7910 2510 7926
rect 2537 7924 2572 7937
rect 2613 7934 2650 7937
rect 2613 7932 2655 7934
rect 2542 7921 2572 7924
rect 2551 7917 2558 7921
rect 2558 7916 2559 7917
rect 2517 7910 2527 7916
rect 2276 7902 2311 7910
rect 2276 7876 2277 7902
rect 2284 7876 2311 7902
rect 2219 7858 2249 7872
rect 2276 7868 2311 7876
rect 2313 7902 2354 7910
rect 2313 7876 2328 7902
rect 2335 7876 2354 7902
rect 2418 7898 2449 7910
rect 2464 7898 2567 7910
rect 2579 7900 2605 7926
rect 2620 7921 2650 7932
rect 2682 7928 2744 7944
rect 2682 7926 2728 7928
rect 2682 7910 2744 7926
rect 2756 7910 2762 7958
rect 2765 7950 2845 7958
rect 2765 7948 2784 7950
rect 2799 7948 2833 7950
rect 2765 7932 2845 7948
rect 2765 7910 2784 7932
rect 2799 7916 2829 7932
rect 2857 7926 2863 8000
rect 2866 7926 2885 8070
rect 2900 7926 2906 8070
rect 2915 8000 2928 8070
rect 2980 8066 3002 8070
rect 2973 8044 3002 8058
rect 3055 8044 3071 8058
rect 3109 8054 3115 8056
rect 3122 8054 3230 8070
rect 3237 8054 3243 8056
rect 3251 8054 3266 8070
rect 3332 8064 3351 8067
rect 2973 8042 3071 8044
rect 3098 8042 3266 8054
rect 3281 8044 3297 8058
rect 3332 8045 3354 8064
rect 3364 8058 3380 8059
rect 3363 8056 3380 8058
rect 3364 8051 3380 8056
rect 3354 8044 3360 8045
rect 3363 8044 3392 8051
rect 3281 8043 3392 8044
rect 3281 8042 3398 8043
rect 2957 8034 3008 8042
rect 3055 8034 3089 8042
rect 2957 8022 2982 8034
rect 2989 8022 3008 8034
rect 3062 8032 3089 8034
rect 3098 8032 3319 8042
rect 3354 8039 3360 8042
rect 3062 8028 3319 8032
rect 2957 8014 3008 8022
rect 3055 8014 3319 8028
rect 3363 8034 3398 8042
rect 2909 7966 2928 8000
rect 2973 8006 3002 8014
rect 2973 8000 2990 8006
rect 2973 7998 3007 8000
rect 3055 7998 3071 8014
rect 3072 8004 3280 8014
rect 3281 8004 3297 8014
rect 3345 8010 3360 8025
rect 3363 8022 3364 8034
rect 3371 8022 3398 8034
rect 3363 8014 3398 8022
rect 3363 8013 3392 8014
rect 3083 8000 3297 8004
rect 3098 7998 3297 8000
rect 3332 8000 3345 8010
rect 3363 8000 3380 8013
rect 3332 7998 3380 8000
rect 2974 7994 3007 7998
rect 2970 7992 3007 7994
rect 2970 7991 3037 7992
rect 2970 7986 3001 7991
rect 3007 7986 3037 7991
rect 2970 7982 3037 7986
rect 2943 7979 3037 7982
rect 2943 7972 2992 7979
rect 2943 7966 2973 7972
rect 2992 7967 2997 7972
rect 2909 7950 2989 7966
rect 3001 7958 3037 7979
rect 3098 7974 3287 7998
rect 3332 7997 3379 7998
rect 3345 7992 3379 7997
rect 3113 7971 3287 7974
rect 3106 7968 3287 7971
rect 3315 7991 3379 7992
rect 2909 7948 2928 7950
rect 2943 7948 2977 7950
rect 2909 7932 2989 7948
rect 2909 7926 2928 7932
rect 2625 7900 2728 7910
rect 2579 7898 2728 7900
rect 2749 7898 2784 7910
rect 2418 7896 2580 7898
rect 2430 7876 2449 7896
rect 2464 7894 2494 7896
rect 2313 7868 2354 7876
rect 2436 7872 2449 7876
rect 2501 7880 2580 7896
rect 2612 7896 2784 7898
rect 2612 7880 2691 7896
rect 2698 7894 2728 7896
rect 2276 7858 2305 7868
rect 2319 7858 2348 7868
rect 2363 7858 2393 7872
rect 2436 7858 2479 7872
rect 2501 7868 2691 7880
rect 2756 7876 2762 7896
rect 2486 7858 2516 7868
rect 2517 7858 2675 7868
rect 2679 7858 2709 7868
rect 2713 7858 2743 7872
rect 2771 7858 2784 7896
rect 2856 7910 2885 7926
rect 2899 7910 2928 7926
rect 2943 7916 2973 7932
rect 3001 7910 3007 7958
rect 3010 7952 3029 7958
rect 3044 7952 3074 7960
rect 3010 7944 3074 7952
rect 3010 7928 3090 7944
rect 3106 7937 3168 7968
rect 3184 7937 3246 7968
rect 3315 7966 3364 7991
rect 3379 7966 3409 7982
rect 3278 7952 3308 7960
rect 3315 7958 3425 7966
rect 3278 7944 3323 7952
rect 3010 7926 3029 7928
rect 3044 7926 3090 7928
rect 3010 7910 3090 7926
rect 3117 7924 3152 7937
rect 3193 7934 3230 7937
rect 3193 7932 3235 7934
rect 3122 7921 3152 7924
rect 3131 7917 3138 7921
rect 3138 7916 3139 7917
rect 3097 7910 3107 7916
rect 2856 7902 2891 7910
rect 2856 7876 2857 7902
rect 2864 7876 2891 7902
rect 2799 7858 2829 7872
rect 2856 7868 2891 7876
rect 2893 7902 2934 7910
rect 2893 7876 2908 7902
rect 2915 7876 2934 7902
rect 2998 7898 3029 7910
rect 3044 7898 3147 7910
rect 3159 7900 3185 7926
rect 3200 7921 3230 7932
rect 3262 7928 3324 7944
rect 3262 7926 3308 7928
rect 3262 7910 3324 7926
rect 3336 7910 3342 7958
rect 3345 7950 3425 7958
rect 3345 7948 3364 7950
rect 3379 7948 3413 7950
rect 3345 7932 3425 7948
rect 3345 7910 3364 7932
rect 3379 7916 3409 7932
rect 3437 7926 3443 8000
rect 3446 7926 3465 8070
rect 3480 7926 3486 8070
rect 3495 8000 3508 8070
rect 3560 8066 3582 8070
rect 3553 8044 3582 8058
rect 3635 8044 3651 8058
rect 3689 8054 3695 8056
rect 3702 8054 3810 8070
rect 3817 8054 3823 8056
rect 3831 8054 3846 8070
rect 3912 8064 3931 8067
rect 3553 8042 3651 8044
rect 3678 8042 3846 8054
rect 3861 8044 3877 8058
rect 3912 8045 3934 8064
rect 3944 8058 3960 8059
rect 3943 8056 3960 8058
rect 3944 8051 3960 8056
rect 3934 8044 3940 8045
rect 3943 8044 3972 8051
rect 3861 8043 3972 8044
rect 3861 8042 3978 8043
rect 3537 8034 3588 8042
rect 3635 8034 3669 8042
rect 3537 8022 3562 8034
rect 3569 8022 3588 8034
rect 3642 8032 3669 8034
rect 3678 8032 3899 8042
rect 3934 8039 3940 8042
rect 3642 8028 3899 8032
rect 3537 8014 3588 8022
rect 3635 8014 3899 8028
rect 3943 8034 3978 8042
rect 3489 7966 3508 8000
rect 3553 8006 3582 8014
rect 3553 8000 3570 8006
rect 3553 7998 3587 8000
rect 3635 7998 3651 8014
rect 3652 8004 3860 8014
rect 3861 8004 3877 8014
rect 3925 8010 3940 8025
rect 3943 8022 3944 8034
rect 3951 8022 3978 8034
rect 3943 8014 3978 8022
rect 3943 8013 3972 8014
rect 3663 8000 3877 8004
rect 3678 7998 3877 8000
rect 3912 8000 3925 8010
rect 3943 8000 3960 8013
rect 3912 7998 3960 8000
rect 3554 7994 3587 7998
rect 3550 7992 3587 7994
rect 3550 7991 3617 7992
rect 3550 7986 3581 7991
rect 3587 7986 3617 7991
rect 3550 7982 3617 7986
rect 3523 7979 3617 7982
rect 3523 7972 3572 7979
rect 3523 7966 3553 7972
rect 3572 7967 3577 7972
rect 3489 7950 3569 7966
rect 3581 7958 3617 7979
rect 3678 7974 3867 7998
rect 3912 7997 3959 7998
rect 3925 7992 3959 7997
rect 3693 7971 3867 7974
rect 3686 7968 3867 7971
rect 3895 7991 3959 7992
rect 3489 7948 3508 7950
rect 3523 7948 3557 7950
rect 3489 7932 3569 7948
rect 3489 7926 3508 7932
rect 3205 7900 3308 7910
rect 3159 7898 3308 7900
rect 3329 7898 3364 7910
rect 2998 7896 3160 7898
rect 3010 7876 3029 7896
rect 3044 7894 3074 7896
rect 2893 7868 2934 7876
rect 3016 7872 3029 7876
rect 3081 7880 3160 7896
rect 3192 7896 3364 7898
rect 3192 7880 3271 7896
rect 3278 7894 3308 7896
rect 2856 7858 2885 7868
rect 2899 7858 2928 7868
rect 2943 7858 2973 7872
rect 3016 7858 3059 7872
rect 3081 7868 3271 7880
rect 3336 7876 3342 7896
rect 3066 7858 3096 7868
rect 3097 7858 3255 7868
rect 3259 7858 3289 7868
rect 3293 7858 3323 7872
rect 3351 7858 3364 7896
rect 3436 7910 3465 7926
rect 3479 7910 3508 7926
rect 3523 7916 3553 7932
rect 3581 7910 3587 7958
rect 3590 7952 3609 7958
rect 3624 7952 3654 7960
rect 3590 7944 3654 7952
rect 3590 7928 3670 7944
rect 3686 7937 3748 7968
rect 3764 7937 3826 7968
rect 3895 7966 3944 7991
rect 3959 7966 3989 7982
rect 3858 7952 3888 7960
rect 3895 7958 4005 7966
rect 3858 7944 3903 7952
rect 3590 7926 3609 7928
rect 3624 7926 3670 7928
rect 3590 7910 3670 7926
rect 3697 7924 3732 7937
rect 3773 7934 3810 7937
rect 3773 7932 3815 7934
rect 3702 7921 3732 7924
rect 3711 7917 3718 7921
rect 3718 7916 3719 7917
rect 3677 7910 3687 7916
rect 3436 7902 3471 7910
rect 3436 7876 3437 7902
rect 3444 7876 3471 7902
rect 3379 7858 3409 7872
rect 3436 7868 3471 7876
rect 3473 7902 3514 7910
rect 3473 7876 3488 7902
rect 3495 7876 3514 7902
rect 3578 7898 3609 7910
rect 3624 7898 3727 7910
rect 3739 7900 3765 7926
rect 3780 7921 3810 7932
rect 3842 7928 3904 7944
rect 3842 7926 3888 7928
rect 3842 7910 3904 7926
rect 3916 7910 3922 7958
rect 3925 7950 4005 7958
rect 3925 7948 3944 7950
rect 3959 7948 3993 7950
rect 3925 7932 4005 7948
rect 3925 7910 3944 7932
rect 3959 7916 3989 7932
rect 4017 7926 4023 8000
rect 4026 7926 4045 8070
rect 4060 7926 4066 8070
rect 4075 8000 4088 8070
rect 4140 8066 4162 8070
rect 4133 8044 4162 8058
rect 4215 8044 4231 8058
rect 4269 8054 4275 8056
rect 4282 8054 4390 8070
rect 4397 8054 4403 8056
rect 4411 8054 4426 8070
rect 4492 8064 4511 8067
rect 4133 8042 4231 8044
rect 4258 8042 4426 8054
rect 4441 8044 4457 8058
rect 4492 8045 4514 8064
rect 4524 8058 4540 8059
rect 4523 8056 4540 8058
rect 4524 8051 4540 8056
rect 4514 8044 4520 8045
rect 4523 8044 4552 8051
rect 4441 8043 4552 8044
rect 4441 8042 4558 8043
rect 4117 8034 4168 8042
rect 4215 8034 4249 8042
rect 4117 8022 4142 8034
rect 4149 8022 4168 8034
rect 4222 8032 4249 8034
rect 4258 8032 4479 8042
rect 4514 8039 4520 8042
rect 4222 8028 4479 8032
rect 4117 8014 4168 8022
rect 4215 8014 4479 8028
rect 4523 8034 4558 8042
rect 4069 7966 4088 8000
rect 4133 8006 4162 8014
rect 4133 8000 4150 8006
rect 4133 7998 4167 8000
rect 4215 7998 4231 8014
rect 4232 8004 4440 8014
rect 4441 8004 4457 8014
rect 4505 8010 4520 8025
rect 4523 8022 4524 8034
rect 4531 8022 4558 8034
rect 4523 8014 4558 8022
rect 4523 8013 4552 8014
rect 4243 8000 4457 8004
rect 4258 7998 4457 8000
rect 4492 8000 4505 8010
rect 4523 8000 4540 8013
rect 4492 7998 4540 8000
rect 4134 7994 4167 7998
rect 4130 7992 4167 7994
rect 4130 7991 4197 7992
rect 4130 7986 4161 7991
rect 4167 7986 4197 7991
rect 4130 7982 4197 7986
rect 4103 7979 4197 7982
rect 4103 7972 4152 7979
rect 4103 7966 4133 7972
rect 4152 7967 4157 7972
rect 4069 7950 4149 7966
rect 4161 7958 4197 7979
rect 4258 7974 4447 7998
rect 4492 7997 4539 7998
rect 4505 7992 4539 7997
rect 4273 7971 4447 7974
rect 4266 7968 4447 7971
rect 4475 7991 4539 7992
rect 4069 7948 4088 7950
rect 4103 7948 4137 7950
rect 4069 7932 4149 7948
rect 4069 7926 4088 7932
rect 3785 7900 3888 7910
rect 3739 7898 3888 7900
rect 3909 7898 3944 7910
rect 3578 7896 3740 7898
rect 3590 7876 3609 7896
rect 3624 7894 3654 7896
rect 3473 7868 3514 7876
rect 3596 7872 3609 7876
rect 3661 7880 3740 7896
rect 3772 7896 3944 7898
rect 3772 7880 3851 7896
rect 3858 7894 3888 7896
rect 3436 7858 3465 7868
rect 3479 7858 3508 7868
rect 3523 7858 3553 7872
rect 3596 7858 3639 7872
rect 3661 7868 3851 7880
rect 3916 7876 3922 7896
rect 3646 7858 3676 7868
rect 3677 7858 3835 7868
rect 3839 7858 3869 7868
rect 3873 7858 3903 7872
rect 3931 7858 3944 7896
rect 4016 7910 4045 7926
rect 4059 7910 4088 7926
rect 4103 7916 4133 7932
rect 4161 7910 4167 7958
rect 4170 7952 4189 7958
rect 4204 7952 4234 7960
rect 4170 7944 4234 7952
rect 4170 7928 4250 7944
rect 4266 7937 4328 7968
rect 4344 7937 4406 7968
rect 4475 7966 4524 7991
rect 4539 7966 4569 7982
rect 4438 7952 4468 7960
rect 4475 7958 4585 7966
rect 4438 7944 4483 7952
rect 4170 7926 4189 7928
rect 4204 7926 4250 7928
rect 4170 7910 4250 7926
rect 4277 7924 4312 7937
rect 4353 7934 4390 7937
rect 4353 7932 4395 7934
rect 4282 7921 4312 7924
rect 4291 7917 4298 7921
rect 4298 7916 4299 7917
rect 4257 7910 4267 7916
rect 4016 7902 4051 7910
rect 4016 7876 4017 7902
rect 4024 7876 4051 7902
rect 3959 7858 3989 7872
rect 4016 7868 4051 7876
rect 4053 7902 4094 7910
rect 4053 7876 4068 7902
rect 4075 7876 4094 7902
rect 4158 7898 4189 7910
rect 4204 7898 4307 7910
rect 4319 7900 4345 7926
rect 4360 7921 4390 7932
rect 4422 7928 4484 7944
rect 4422 7926 4468 7928
rect 4422 7910 4484 7926
rect 4496 7910 4502 7958
rect 4505 7950 4585 7958
rect 4505 7948 4524 7950
rect 4539 7948 4573 7950
rect 4505 7932 4585 7948
rect 4505 7910 4524 7932
rect 4539 7916 4569 7932
rect 4597 7926 4603 8000
rect 4606 7926 4625 8070
rect 4640 7926 4646 8070
rect 4655 8000 4668 8070
rect 4720 8066 4742 8070
rect 4713 8044 4742 8058
rect 4795 8044 4811 8058
rect 4849 8054 4855 8056
rect 4862 8054 4970 8070
rect 4977 8054 4983 8056
rect 4991 8054 5006 8070
rect 5072 8064 5091 8067
rect 4713 8042 4811 8044
rect 4838 8042 5006 8054
rect 5021 8044 5037 8058
rect 5072 8045 5094 8064
rect 5104 8058 5120 8059
rect 5103 8056 5120 8058
rect 5104 8051 5120 8056
rect 5094 8044 5100 8045
rect 5103 8044 5132 8051
rect 5021 8043 5132 8044
rect 5021 8042 5138 8043
rect 4697 8034 4748 8042
rect 4795 8034 4829 8042
rect 4697 8022 4722 8034
rect 4729 8022 4748 8034
rect 4802 8032 4829 8034
rect 4838 8032 5059 8042
rect 5094 8039 5100 8042
rect 4802 8028 5059 8032
rect 4697 8014 4748 8022
rect 4795 8014 5059 8028
rect 5103 8034 5138 8042
rect 4649 7966 4668 8000
rect 4713 8006 4742 8014
rect 4713 8000 4730 8006
rect 4713 7998 4747 8000
rect 4795 7998 4811 8014
rect 4812 8004 5020 8014
rect 5021 8004 5037 8014
rect 5085 8010 5100 8025
rect 5103 8022 5104 8034
rect 5111 8022 5138 8034
rect 5103 8014 5138 8022
rect 5103 8013 5132 8014
rect 4823 8000 5037 8004
rect 4838 7998 5037 8000
rect 5072 8000 5085 8010
rect 5103 8000 5120 8013
rect 5072 7998 5120 8000
rect 4714 7994 4747 7998
rect 4710 7992 4747 7994
rect 4710 7991 4777 7992
rect 4710 7986 4741 7991
rect 4747 7986 4777 7991
rect 4710 7982 4777 7986
rect 4683 7979 4777 7982
rect 4683 7972 4732 7979
rect 4683 7966 4713 7972
rect 4732 7967 4737 7972
rect 4649 7950 4729 7966
rect 4741 7958 4777 7979
rect 4838 7974 5027 7998
rect 5072 7997 5119 7998
rect 5085 7992 5119 7997
rect 4853 7971 5027 7974
rect 4846 7968 5027 7971
rect 5055 7991 5119 7992
rect 4649 7948 4668 7950
rect 4683 7948 4717 7950
rect 4649 7932 4729 7948
rect 4649 7926 4668 7932
rect 4365 7900 4468 7910
rect 4319 7898 4468 7900
rect 4489 7898 4524 7910
rect 4158 7896 4320 7898
rect 4170 7876 4189 7896
rect 4204 7894 4234 7896
rect 4053 7868 4094 7876
rect 4176 7872 4189 7876
rect 4241 7880 4320 7896
rect 4352 7896 4524 7898
rect 4352 7880 4431 7896
rect 4438 7894 4468 7896
rect 4016 7858 4045 7868
rect 4059 7858 4088 7868
rect 4103 7858 4133 7872
rect 4176 7858 4219 7872
rect 4241 7868 4431 7880
rect 4496 7876 4502 7896
rect 4226 7858 4256 7868
rect 4257 7858 4415 7868
rect 4419 7858 4449 7868
rect 4453 7858 4483 7872
rect 4511 7858 4524 7896
rect 4596 7910 4625 7926
rect 4639 7910 4668 7926
rect 4683 7916 4713 7932
rect 4741 7910 4747 7958
rect 4750 7952 4769 7958
rect 4784 7952 4814 7960
rect 4750 7944 4814 7952
rect 4750 7928 4830 7944
rect 4846 7937 4908 7968
rect 4924 7937 4986 7968
rect 5055 7966 5104 7991
rect 5119 7966 5149 7982
rect 5018 7952 5048 7960
rect 5055 7958 5165 7966
rect 5018 7944 5063 7952
rect 4750 7926 4769 7928
rect 4784 7926 4830 7928
rect 4750 7910 4830 7926
rect 4857 7924 4892 7937
rect 4933 7934 4970 7937
rect 4933 7932 4975 7934
rect 4862 7921 4892 7924
rect 4871 7917 4878 7921
rect 4878 7916 4879 7917
rect 4837 7910 4847 7916
rect 4596 7902 4631 7910
rect 4596 7876 4597 7902
rect 4604 7876 4631 7902
rect 4539 7858 4569 7872
rect 4596 7868 4631 7876
rect 4633 7902 4674 7910
rect 4633 7876 4648 7902
rect 4655 7876 4674 7902
rect 4738 7898 4769 7910
rect 4784 7898 4887 7910
rect 4899 7900 4925 7926
rect 4940 7921 4970 7932
rect 5002 7928 5064 7944
rect 5002 7926 5048 7928
rect 5002 7910 5064 7926
rect 5076 7910 5082 7958
rect 5085 7950 5165 7958
rect 5085 7948 5104 7950
rect 5119 7948 5153 7950
rect 5085 7932 5165 7948
rect 5085 7910 5104 7932
rect 5119 7916 5149 7932
rect 5177 7926 5183 8000
rect 5186 7926 5205 8070
rect 5220 7926 5226 8070
rect 5235 8000 5248 8070
rect 5300 8066 5322 8070
rect 5293 8044 5322 8058
rect 5375 8044 5391 8058
rect 5429 8054 5435 8056
rect 5442 8054 5550 8070
rect 5557 8054 5563 8056
rect 5571 8054 5586 8070
rect 5652 8064 5671 8067
rect 5293 8042 5391 8044
rect 5418 8042 5586 8054
rect 5601 8044 5617 8058
rect 5652 8045 5674 8064
rect 5684 8058 5700 8059
rect 5683 8056 5700 8058
rect 5684 8051 5700 8056
rect 5674 8044 5680 8045
rect 5683 8044 5712 8051
rect 5601 8043 5712 8044
rect 5601 8042 5718 8043
rect 5277 8034 5328 8042
rect 5375 8034 5409 8042
rect 5277 8022 5302 8034
rect 5309 8022 5328 8034
rect 5382 8032 5409 8034
rect 5418 8032 5639 8042
rect 5674 8039 5680 8042
rect 5382 8028 5639 8032
rect 5277 8014 5328 8022
rect 5375 8014 5639 8028
rect 5683 8034 5718 8042
rect 5229 7966 5248 8000
rect 5293 8006 5322 8014
rect 5293 8000 5310 8006
rect 5293 7998 5327 8000
rect 5375 7998 5391 8014
rect 5392 8004 5600 8014
rect 5601 8004 5617 8014
rect 5665 8010 5680 8025
rect 5683 8022 5684 8034
rect 5691 8022 5718 8034
rect 5683 8014 5718 8022
rect 5683 8013 5712 8014
rect 5403 8000 5617 8004
rect 5418 7998 5617 8000
rect 5652 8000 5665 8010
rect 5683 8000 5700 8013
rect 5652 7998 5700 8000
rect 5294 7994 5327 7998
rect 5290 7992 5327 7994
rect 5290 7991 5357 7992
rect 5290 7986 5321 7991
rect 5327 7986 5357 7991
rect 5290 7982 5357 7986
rect 5263 7979 5357 7982
rect 5263 7972 5312 7979
rect 5263 7966 5293 7972
rect 5312 7967 5317 7972
rect 5229 7950 5309 7966
rect 5321 7958 5357 7979
rect 5418 7974 5607 7998
rect 5652 7997 5699 7998
rect 5665 7992 5699 7997
rect 5433 7971 5607 7974
rect 5426 7968 5607 7971
rect 5635 7991 5699 7992
rect 5229 7948 5248 7950
rect 5263 7948 5297 7950
rect 5229 7932 5309 7948
rect 5229 7926 5248 7932
rect 4945 7900 5048 7910
rect 4899 7898 5048 7900
rect 5069 7898 5104 7910
rect 4738 7896 4900 7898
rect 4750 7876 4769 7896
rect 4784 7894 4814 7896
rect 4633 7868 4674 7876
rect 4756 7872 4769 7876
rect 4821 7880 4900 7896
rect 4932 7896 5104 7898
rect 4932 7880 5011 7896
rect 5018 7894 5048 7896
rect 4596 7858 4625 7868
rect 4639 7858 4668 7868
rect 4683 7858 4713 7872
rect 4756 7858 4799 7872
rect 4821 7868 5011 7880
rect 5076 7876 5082 7896
rect 4806 7858 4836 7868
rect 4837 7858 4995 7868
rect 4999 7858 5029 7868
rect 5033 7858 5063 7872
rect 5091 7858 5104 7896
rect 5176 7910 5205 7926
rect 5219 7910 5248 7926
rect 5263 7916 5293 7932
rect 5321 7910 5327 7958
rect 5330 7952 5349 7958
rect 5364 7952 5394 7960
rect 5330 7944 5394 7952
rect 5330 7928 5410 7944
rect 5426 7937 5488 7968
rect 5504 7937 5566 7968
rect 5635 7966 5684 7991
rect 5699 7966 5729 7982
rect 5598 7952 5628 7960
rect 5635 7958 5745 7966
rect 5598 7944 5643 7952
rect 5330 7926 5349 7928
rect 5364 7926 5410 7928
rect 5330 7910 5410 7926
rect 5437 7924 5472 7937
rect 5513 7934 5550 7937
rect 5513 7932 5555 7934
rect 5442 7921 5472 7924
rect 5451 7917 5458 7921
rect 5458 7916 5459 7917
rect 5417 7910 5427 7916
rect 5176 7902 5211 7910
rect 5176 7876 5177 7902
rect 5184 7876 5211 7902
rect 5119 7858 5149 7872
rect 5176 7868 5211 7876
rect 5213 7902 5254 7910
rect 5213 7876 5228 7902
rect 5235 7876 5254 7902
rect 5318 7898 5349 7910
rect 5364 7898 5467 7910
rect 5479 7900 5505 7926
rect 5520 7921 5550 7932
rect 5582 7928 5644 7944
rect 5582 7926 5628 7928
rect 5582 7910 5644 7926
rect 5656 7910 5662 7958
rect 5665 7950 5745 7958
rect 5665 7948 5684 7950
rect 5699 7948 5733 7950
rect 5665 7932 5745 7948
rect 5665 7910 5684 7932
rect 5699 7916 5729 7932
rect 5757 7926 5763 8000
rect 5766 7926 5785 8070
rect 5800 7926 5806 8070
rect 5815 8000 5828 8070
rect 5880 8066 5902 8070
rect 5873 8044 5902 8058
rect 5955 8044 5971 8058
rect 6009 8054 6015 8056
rect 6022 8054 6130 8070
rect 6137 8054 6143 8056
rect 6151 8054 6166 8070
rect 6232 8064 6251 8067
rect 5873 8042 5971 8044
rect 5998 8042 6166 8054
rect 6181 8044 6197 8058
rect 6232 8045 6254 8064
rect 6264 8058 6280 8059
rect 6263 8056 6280 8058
rect 6264 8051 6280 8056
rect 6254 8044 6260 8045
rect 6263 8044 6292 8051
rect 6181 8043 6292 8044
rect 6181 8042 6298 8043
rect 5857 8034 5908 8042
rect 5955 8034 5989 8042
rect 5857 8022 5882 8034
rect 5889 8022 5908 8034
rect 5962 8032 5989 8034
rect 5998 8032 6219 8042
rect 6254 8039 6260 8042
rect 5962 8028 6219 8032
rect 5857 8014 5908 8022
rect 5955 8014 6219 8028
rect 6263 8034 6298 8042
rect 5809 7966 5828 8000
rect 5873 8006 5902 8014
rect 5873 8000 5890 8006
rect 5873 7998 5907 8000
rect 5955 7998 5971 8014
rect 5972 8004 6180 8014
rect 6181 8004 6197 8014
rect 6245 8010 6260 8025
rect 6263 8022 6264 8034
rect 6271 8022 6298 8034
rect 6263 8014 6298 8022
rect 6263 8013 6292 8014
rect 5983 8000 6197 8004
rect 5998 7998 6197 8000
rect 6232 8000 6245 8010
rect 6263 8000 6280 8013
rect 6232 7998 6280 8000
rect 5874 7994 5907 7998
rect 5870 7992 5907 7994
rect 5870 7991 5937 7992
rect 5870 7986 5901 7991
rect 5907 7986 5937 7991
rect 5870 7982 5937 7986
rect 5843 7979 5937 7982
rect 5843 7972 5892 7979
rect 5843 7966 5873 7972
rect 5892 7967 5897 7972
rect 5809 7950 5889 7966
rect 5901 7958 5937 7979
rect 5998 7974 6187 7998
rect 6232 7997 6279 7998
rect 6245 7992 6279 7997
rect 6013 7971 6187 7974
rect 6006 7968 6187 7971
rect 6215 7991 6279 7992
rect 5809 7948 5828 7950
rect 5843 7948 5877 7950
rect 5809 7932 5889 7948
rect 5809 7926 5828 7932
rect 5525 7900 5628 7910
rect 5479 7898 5628 7900
rect 5649 7898 5684 7910
rect 5318 7896 5480 7898
rect 5330 7876 5349 7896
rect 5364 7894 5394 7896
rect 5213 7868 5254 7876
rect 5336 7872 5349 7876
rect 5401 7880 5480 7896
rect 5512 7896 5684 7898
rect 5512 7880 5591 7896
rect 5598 7894 5628 7896
rect 5176 7858 5205 7868
rect 5219 7858 5248 7868
rect 5263 7858 5293 7872
rect 5336 7858 5379 7872
rect 5401 7868 5591 7880
rect 5656 7876 5662 7896
rect 5386 7858 5416 7868
rect 5417 7858 5575 7868
rect 5579 7858 5609 7868
rect 5613 7858 5643 7872
rect 5671 7858 5684 7896
rect 5756 7910 5785 7926
rect 5799 7910 5828 7926
rect 5843 7916 5873 7932
rect 5901 7910 5907 7958
rect 5910 7952 5929 7958
rect 5944 7952 5974 7960
rect 5910 7944 5974 7952
rect 5910 7928 5990 7944
rect 6006 7937 6068 7968
rect 6084 7937 6146 7968
rect 6215 7966 6264 7991
rect 6279 7966 6309 7982
rect 6178 7952 6208 7960
rect 6215 7958 6325 7966
rect 6178 7944 6223 7952
rect 5910 7926 5929 7928
rect 5944 7926 5990 7928
rect 5910 7910 5990 7926
rect 6017 7924 6052 7937
rect 6093 7934 6130 7937
rect 6093 7932 6135 7934
rect 6022 7921 6052 7924
rect 6031 7917 6038 7921
rect 6038 7916 6039 7917
rect 5997 7910 6007 7916
rect 5756 7902 5791 7910
rect 5756 7876 5757 7902
rect 5764 7876 5791 7902
rect 5699 7858 5729 7872
rect 5756 7868 5791 7876
rect 5793 7902 5834 7910
rect 5793 7876 5808 7902
rect 5815 7876 5834 7902
rect 5898 7898 5929 7910
rect 5944 7898 6047 7910
rect 6059 7900 6085 7926
rect 6100 7921 6130 7932
rect 6162 7928 6224 7944
rect 6162 7926 6208 7928
rect 6162 7910 6224 7926
rect 6236 7910 6242 7958
rect 6245 7950 6325 7958
rect 6245 7948 6264 7950
rect 6279 7948 6313 7950
rect 6245 7932 6325 7948
rect 6245 7910 6264 7932
rect 6279 7916 6309 7932
rect 6337 7926 6343 8000
rect 6346 7926 6365 8070
rect 6380 7926 6386 8070
rect 6395 8000 6408 8070
rect 6460 8066 6482 8070
rect 6453 8044 6482 8058
rect 6535 8044 6551 8058
rect 6589 8054 6595 8056
rect 6602 8054 6710 8070
rect 6717 8054 6723 8056
rect 6731 8054 6746 8070
rect 6812 8064 6831 8067
rect 6453 8042 6551 8044
rect 6578 8042 6746 8054
rect 6761 8044 6777 8058
rect 6812 8045 6834 8064
rect 6844 8058 6860 8059
rect 6843 8056 6860 8058
rect 6844 8051 6860 8056
rect 6834 8044 6840 8045
rect 6843 8044 6872 8051
rect 6761 8043 6872 8044
rect 6761 8042 6878 8043
rect 6437 8034 6488 8042
rect 6535 8034 6569 8042
rect 6437 8022 6462 8034
rect 6469 8022 6488 8034
rect 6542 8032 6569 8034
rect 6578 8032 6799 8042
rect 6834 8039 6840 8042
rect 6542 8028 6799 8032
rect 6437 8014 6488 8022
rect 6535 8014 6799 8028
rect 6843 8034 6878 8042
rect 6389 7966 6408 8000
rect 6453 8006 6482 8014
rect 6453 8000 6470 8006
rect 6453 7998 6487 8000
rect 6535 7998 6551 8014
rect 6552 8004 6760 8014
rect 6761 8004 6777 8014
rect 6825 8010 6840 8025
rect 6843 8022 6844 8034
rect 6851 8022 6878 8034
rect 6843 8014 6878 8022
rect 6843 8013 6872 8014
rect 6563 8000 6777 8004
rect 6578 7998 6777 8000
rect 6812 8000 6825 8010
rect 6843 8000 6860 8013
rect 6812 7998 6860 8000
rect 6454 7994 6487 7998
rect 6450 7992 6487 7994
rect 6450 7991 6517 7992
rect 6450 7986 6481 7991
rect 6487 7986 6517 7991
rect 6450 7982 6517 7986
rect 6423 7979 6517 7982
rect 6423 7972 6472 7979
rect 6423 7966 6453 7972
rect 6472 7967 6477 7972
rect 6389 7950 6469 7966
rect 6481 7958 6517 7979
rect 6578 7974 6767 7998
rect 6812 7997 6859 7998
rect 6825 7992 6859 7997
rect 6593 7971 6767 7974
rect 6586 7968 6767 7971
rect 6795 7991 6859 7992
rect 6389 7948 6408 7950
rect 6423 7948 6457 7950
rect 6389 7932 6469 7948
rect 6389 7926 6408 7932
rect 6105 7900 6208 7910
rect 6059 7898 6208 7900
rect 6229 7898 6264 7910
rect 5898 7896 6060 7898
rect 5910 7876 5929 7896
rect 5944 7894 5974 7896
rect 5793 7868 5834 7876
rect 5916 7872 5929 7876
rect 5981 7880 6060 7896
rect 6092 7896 6264 7898
rect 6092 7880 6171 7896
rect 6178 7894 6208 7896
rect 5756 7858 5785 7868
rect 5799 7858 5828 7868
rect 5843 7858 5873 7872
rect 5916 7858 5959 7872
rect 5981 7868 6171 7880
rect 6236 7876 6242 7896
rect 5966 7858 5996 7868
rect 5997 7858 6155 7868
rect 6159 7858 6189 7868
rect 6193 7858 6223 7872
rect 6251 7858 6264 7896
rect 6336 7910 6365 7926
rect 6379 7910 6408 7926
rect 6423 7916 6453 7932
rect 6481 7910 6487 7958
rect 6490 7952 6509 7958
rect 6524 7952 6554 7960
rect 6490 7944 6554 7952
rect 6490 7928 6570 7944
rect 6586 7937 6648 7968
rect 6664 7937 6726 7968
rect 6795 7966 6844 7991
rect 6859 7966 6889 7982
rect 6758 7952 6788 7960
rect 6795 7958 6905 7966
rect 6758 7944 6803 7952
rect 6490 7926 6509 7928
rect 6524 7926 6570 7928
rect 6490 7910 6570 7926
rect 6597 7924 6632 7937
rect 6673 7934 6710 7937
rect 6673 7932 6715 7934
rect 6602 7921 6632 7924
rect 6611 7917 6618 7921
rect 6618 7916 6619 7917
rect 6577 7910 6587 7916
rect 6336 7902 6371 7910
rect 6336 7876 6337 7902
rect 6344 7876 6371 7902
rect 6279 7858 6309 7872
rect 6336 7868 6371 7876
rect 6373 7902 6414 7910
rect 6373 7876 6388 7902
rect 6395 7876 6414 7902
rect 6478 7898 6509 7910
rect 6524 7898 6627 7910
rect 6639 7900 6665 7926
rect 6680 7921 6710 7932
rect 6742 7928 6804 7944
rect 6742 7926 6788 7928
rect 6742 7910 6804 7926
rect 6816 7910 6822 7958
rect 6825 7950 6905 7958
rect 6825 7948 6844 7950
rect 6859 7948 6893 7950
rect 6825 7932 6905 7948
rect 6825 7910 6844 7932
rect 6859 7916 6889 7932
rect 6917 7926 6923 8000
rect 6926 7926 6945 8070
rect 6960 7926 6966 8070
rect 6975 8000 6988 8070
rect 7040 8066 7062 8070
rect 7033 8044 7062 8058
rect 7115 8044 7131 8058
rect 7169 8054 7175 8056
rect 7182 8054 7290 8070
rect 7297 8054 7303 8056
rect 7311 8054 7326 8070
rect 7392 8064 7411 8067
rect 7033 8042 7131 8044
rect 7158 8042 7326 8054
rect 7341 8044 7357 8058
rect 7392 8045 7414 8064
rect 7424 8058 7440 8059
rect 7423 8056 7440 8058
rect 7424 8051 7440 8056
rect 7414 8044 7420 8045
rect 7423 8044 7452 8051
rect 7341 8043 7452 8044
rect 7341 8042 7458 8043
rect 7017 8034 7068 8042
rect 7115 8034 7149 8042
rect 7017 8022 7042 8034
rect 7049 8022 7068 8034
rect 7122 8032 7149 8034
rect 7158 8032 7379 8042
rect 7414 8039 7420 8042
rect 7122 8028 7379 8032
rect 7017 8014 7068 8022
rect 7115 8014 7379 8028
rect 7423 8034 7458 8042
rect 6969 7966 6988 8000
rect 7033 8006 7062 8014
rect 7033 8000 7050 8006
rect 7033 7998 7067 8000
rect 7115 7998 7131 8014
rect 7132 8004 7340 8014
rect 7341 8004 7357 8014
rect 7405 8010 7420 8025
rect 7423 8022 7424 8034
rect 7431 8022 7458 8034
rect 7423 8014 7458 8022
rect 7423 8013 7452 8014
rect 7143 8000 7357 8004
rect 7158 7998 7357 8000
rect 7392 8000 7405 8010
rect 7423 8000 7440 8013
rect 7392 7998 7440 8000
rect 7034 7994 7067 7998
rect 7030 7992 7067 7994
rect 7030 7991 7097 7992
rect 7030 7986 7061 7991
rect 7067 7986 7097 7991
rect 7030 7982 7097 7986
rect 7003 7979 7097 7982
rect 7003 7972 7052 7979
rect 7003 7966 7033 7972
rect 7052 7967 7057 7972
rect 6969 7950 7049 7966
rect 7061 7958 7097 7979
rect 7158 7974 7347 7998
rect 7392 7997 7439 7998
rect 7405 7992 7439 7997
rect 7173 7971 7347 7974
rect 7166 7968 7347 7971
rect 7375 7991 7439 7992
rect 6969 7948 6988 7950
rect 7003 7948 7037 7950
rect 6969 7932 7049 7948
rect 6969 7926 6988 7932
rect 6685 7900 6788 7910
rect 6639 7898 6788 7900
rect 6809 7898 6844 7910
rect 6478 7896 6640 7898
rect 6490 7876 6509 7896
rect 6524 7894 6554 7896
rect 6373 7868 6414 7876
rect 6496 7872 6509 7876
rect 6561 7880 6640 7896
rect 6672 7896 6844 7898
rect 6672 7880 6751 7896
rect 6758 7894 6788 7896
rect 6336 7858 6365 7868
rect 6379 7858 6408 7868
rect 6423 7858 6453 7872
rect 6496 7858 6539 7872
rect 6561 7868 6751 7880
rect 6816 7876 6822 7896
rect 6546 7858 6576 7868
rect 6577 7858 6735 7868
rect 6739 7858 6769 7868
rect 6773 7858 6803 7872
rect 6831 7858 6844 7896
rect 6916 7910 6945 7926
rect 6959 7910 6988 7926
rect 7003 7916 7033 7932
rect 7061 7910 7067 7958
rect 7070 7952 7089 7958
rect 7104 7952 7134 7960
rect 7070 7944 7134 7952
rect 7070 7928 7150 7944
rect 7166 7937 7228 7968
rect 7244 7937 7306 7968
rect 7375 7966 7424 7991
rect 7439 7966 7469 7982
rect 7338 7952 7368 7960
rect 7375 7958 7485 7966
rect 7338 7944 7383 7952
rect 7070 7926 7089 7928
rect 7104 7926 7150 7928
rect 7070 7910 7150 7926
rect 7177 7924 7212 7937
rect 7253 7934 7290 7937
rect 7253 7932 7295 7934
rect 7182 7921 7212 7924
rect 7191 7917 7198 7921
rect 7198 7916 7199 7917
rect 7157 7910 7167 7916
rect 6916 7902 6951 7910
rect 6916 7876 6917 7902
rect 6924 7876 6951 7902
rect 6859 7858 6889 7872
rect 6916 7868 6951 7876
rect 6953 7902 6994 7910
rect 6953 7876 6968 7902
rect 6975 7876 6994 7902
rect 7058 7898 7089 7910
rect 7104 7898 7207 7910
rect 7219 7900 7245 7926
rect 7260 7921 7290 7932
rect 7322 7928 7384 7944
rect 7322 7926 7368 7928
rect 7322 7910 7384 7926
rect 7396 7910 7402 7958
rect 7405 7950 7485 7958
rect 7405 7948 7424 7950
rect 7439 7948 7473 7950
rect 7405 7932 7485 7948
rect 7405 7910 7424 7932
rect 7439 7916 7469 7932
rect 7497 7926 7503 8000
rect 7506 7926 7525 8070
rect 7540 7926 7546 8070
rect 7555 8000 7568 8070
rect 7613 8048 7614 8058
rect 7629 8048 7642 8058
rect 7613 8044 7642 8048
rect 7647 8044 7677 8070
rect 7695 8056 7711 8058
rect 7783 8056 7836 8070
rect 7784 8054 7848 8056
rect 7891 8054 7906 8070
rect 7955 8067 7985 8070
rect 7955 8064 7991 8067
rect 7921 8056 7937 8058
rect 7695 8044 7710 8048
rect 7613 8042 7710 8044
rect 7738 8042 7906 8054
rect 7922 8044 7937 8048
rect 7955 8045 7994 8064
rect 8013 8058 8020 8059
rect 8019 8051 8020 8058
rect 8003 8048 8004 8051
rect 8019 8048 8032 8051
rect 7955 8044 7985 8045
rect 7994 8044 8000 8045
rect 8003 8044 8032 8048
rect 7922 8043 8032 8044
rect 7922 8042 8038 8043
rect 7597 8034 7648 8042
rect 7597 8022 7622 8034
rect 7629 8022 7648 8034
rect 7679 8034 7729 8042
rect 7679 8026 7695 8034
rect 7702 8032 7729 8034
rect 7738 8032 7959 8042
rect 7702 8022 7959 8032
rect 7988 8034 8038 8042
rect 7988 8025 8004 8034
rect 7597 8014 7648 8022
rect 7695 8014 7959 8022
rect 7985 8022 8004 8025
rect 8011 8022 8038 8034
rect 7985 8014 8038 8022
rect 7549 7966 7568 8000
rect 7613 8006 7614 8014
rect 7629 8006 7642 8014
rect 7613 7998 7629 8006
rect 7610 7991 7629 7994
rect 7610 7982 7632 7991
rect 7583 7972 7632 7982
rect 7583 7966 7613 7972
rect 7632 7967 7637 7972
rect 7549 7950 7629 7966
rect 7647 7958 7677 8014
rect 7712 8004 7920 8014
rect 7955 8010 8000 8014
rect 8003 8013 8004 8014
rect 8019 8013 8032 8014
rect 7738 7974 7927 8004
rect 7753 7971 7927 7974
rect 7746 7968 7927 7971
rect 7549 7948 7568 7950
rect 7583 7948 7617 7950
rect 7549 7932 7629 7948
rect 7656 7944 7669 7958
rect 7684 7944 7700 7960
rect 7746 7955 7757 7968
rect 7549 7926 7568 7932
rect 7265 7900 7368 7910
rect 7219 7898 7368 7900
rect 7389 7898 7424 7910
rect 7058 7896 7220 7898
rect 7070 7876 7089 7896
rect 7104 7894 7134 7896
rect 6953 7868 6994 7876
rect 7076 7872 7089 7876
rect 7141 7880 7220 7896
rect 7252 7896 7424 7898
rect 7252 7880 7331 7896
rect 7338 7894 7368 7896
rect 6916 7858 6945 7868
rect 6959 7858 6988 7868
rect 7003 7858 7033 7872
rect 7076 7858 7119 7872
rect 7141 7868 7331 7880
rect 7396 7876 7402 7896
rect 7126 7858 7156 7868
rect 7157 7858 7315 7868
rect 7319 7858 7349 7868
rect 7353 7858 7383 7872
rect 7411 7858 7424 7896
rect 7496 7910 7525 7926
rect 7539 7910 7568 7926
rect 7583 7910 7613 7932
rect 7656 7928 7718 7944
rect 7746 7937 7757 7953
rect 7762 7948 7772 7968
rect 7782 7948 7796 7968
rect 7799 7955 7808 7968
rect 7824 7955 7833 7968
rect 7762 7937 7796 7948
rect 7799 7937 7808 7953
rect 7824 7937 7833 7953
rect 7840 7948 7850 7968
rect 7860 7948 7874 7968
rect 7875 7955 7886 7968
rect 7840 7937 7874 7948
rect 7875 7937 7886 7953
rect 7932 7944 7948 7960
rect 7955 7958 7985 8010
rect 8019 8006 8020 8013
rect 8004 7998 8020 8006
rect 7991 7966 8004 7985
rect 8019 7966 8049 7982
rect 7991 7950 8065 7966
rect 7991 7948 8004 7950
rect 8019 7948 8053 7950
rect 7656 7926 7669 7928
rect 7684 7926 7718 7928
rect 7656 7910 7718 7926
rect 7762 7921 7778 7924
rect 7840 7921 7870 7932
rect 7918 7928 7964 7944
rect 7991 7932 8065 7948
rect 7918 7926 7952 7928
rect 7917 7910 7964 7926
rect 7991 7910 8004 7932
rect 8019 7910 8049 7932
rect 8076 7910 8077 7926
rect 8092 7910 8105 8070
rect 8135 7966 8148 8070
rect 8193 8048 8194 8058
rect 8209 8048 8222 8058
rect 8193 8044 8222 8048
rect 8227 8044 8257 8070
rect 8275 8056 8291 8058
rect 8363 8056 8416 8070
rect 8364 8054 8428 8056
rect 8471 8054 8486 8070
rect 8535 8067 8565 8070
rect 8535 8064 8571 8067
rect 8501 8056 8517 8058
rect 8275 8044 8290 8048
rect 8193 8042 8290 8044
rect 8318 8042 8486 8054
rect 8502 8044 8517 8048
rect 8535 8045 8574 8064
rect 8593 8058 8600 8059
rect 8599 8051 8600 8058
rect 8583 8048 8584 8051
rect 8599 8048 8612 8051
rect 8535 8044 8565 8045
rect 8574 8044 8580 8045
rect 8583 8044 8612 8048
rect 8502 8043 8612 8044
rect 8502 8042 8618 8043
rect 8177 8034 8228 8042
rect 8177 8022 8202 8034
rect 8209 8022 8228 8034
rect 8259 8034 8309 8042
rect 8259 8026 8275 8034
rect 8282 8032 8309 8034
rect 8318 8032 8539 8042
rect 8282 8022 8539 8032
rect 8568 8034 8618 8042
rect 8568 8025 8584 8034
rect 8177 8014 8228 8022
rect 8275 8014 8539 8022
rect 8565 8022 8584 8025
rect 8591 8022 8618 8034
rect 8565 8014 8618 8022
rect 8193 8006 8194 8014
rect 8209 8006 8222 8014
rect 8193 7998 8209 8006
rect 8190 7991 8209 7994
rect 8190 7982 8212 7991
rect 8163 7972 8212 7982
rect 8163 7966 8193 7972
rect 8212 7967 8217 7972
rect 8135 7950 8209 7966
rect 8227 7958 8257 8014
rect 8292 8004 8500 8014
rect 8535 8010 8580 8014
rect 8583 8013 8584 8014
rect 8599 8013 8612 8014
rect 8318 7974 8507 8004
rect 8333 7971 8507 7974
rect 8326 7968 8507 7971
rect 8135 7948 8148 7950
rect 8163 7948 8197 7950
rect 8135 7932 8209 7948
rect 8236 7944 8249 7958
rect 8264 7944 8280 7960
rect 8326 7955 8337 7968
rect 8119 7910 8120 7926
rect 8135 7910 8148 7932
rect 8163 7910 8193 7932
rect 8236 7928 8298 7944
rect 8326 7937 8337 7953
rect 8342 7948 8352 7968
rect 8362 7948 8376 7968
rect 8379 7955 8388 7968
rect 8404 7955 8413 7968
rect 8342 7937 8376 7948
rect 8379 7937 8388 7953
rect 8404 7937 8413 7953
rect 8420 7948 8430 7968
rect 8440 7948 8454 7968
rect 8455 7955 8466 7968
rect 8420 7937 8454 7948
rect 8455 7937 8466 7953
rect 8512 7944 8528 7960
rect 8535 7958 8565 8010
rect 8599 8006 8600 8013
rect 8584 7998 8600 8006
rect 8571 7966 8584 7985
rect 8599 7966 8629 7982
rect 8571 7950 8645 7966
rect 8571 7948 8584 7950
rect 8599 7948 8633 7950
rect 8236 7926 8249 7928
rect 8264 7926 8298 7928
rect 8236 7910 8298 7926
rect 8342 7921 8358 7924
rect 8420 7921 8450 7932
rect 8498 7928 8544 7944
rect 8571 7932 8645 7948
rect 8498 7926 8532 7928
rect 8497 7910 8544 7926
rect 8571 7910 8584 7932
rect 8599 7910 8629 7932
rect 8656 7910 8657 7926
rect 8672 7910 8685 8070
rect 8715 7966 8728 8070
rect 8773 8048 8774 8058
rect 8789 8048 8802 8058
rect 8773 8044 8802 8048
rect 8807 8044 8837 8070
rect 8855 8056 8871 8058
rect 8943 8056 8996 8070
rect 8944 8054 9008 8056
rect 9051 8054 9066 8070
rect 9115 8067 9145 8070
rect 9115 8064 9151 8067
rect 9081 8056 9097 8058
rect 8855 8044 8870 8048
rect 8773 8042 8870 8044
rect 8898 8042 9066 8054
rect 9082 8044 9097 8048
rect 9115 8045 9154 8064
rect 9173 8058 9180 8059
rect 9179 8051 9180 8058
rect 9163 8048 9164 8051
rect 9179 8048 9192 8051
rect 9115 8044 9145 8045
rect 9154 8044 9160 8045
rect 9163 8044 9192 8048
rect 9082 8043 9192 8044
rect 9082 8042 9198 8043
rect 8757 8034 8808 8042
rect 8757 8022 8782 8034
rect 8789 8022 8808 8034
rect 8839 8034 8889 8042
rect 8839 8026 8855 8034
rect 8862 8032 8889 8034
rect 8898 8032 9119 8042
rect 8862 8022 9119 8032
rect 9148 8034 9198 8042
rect 9148 8025 9164 8034
rect 8757 8014 8808 8022
rect 8855 8014 9119 8022
rect 9145 8022 9164 8025
rect 9171 8022 9198 8034
rect 9145 8014 9198 8022
rect 8773 8006 8774 8014
rect 8789 8006 8802 8014
rect 8773 7998 8789 8006
rect 8770 7991 8789 7994
rect 8770 7982 8792 7991
rect 8743 7972 8792 7982
rect 8743 7966 8773 7972
rect 8792 7967 8797 7972
rect 8715 7950 8789 7966
rect 8807 7958 8837 8014
rect 8872 8004 9080 8014
rect 9115 8010 9160 8014
rect 9163 8013 9164 8014
rect 9179 8013 9192 8014
rect 8898 7974 9087 8004
rect 8913 7971 9087 7974
rect 8906 7968 9087 7971
rect 8715 7948 8728 7950
rect 8743 7948 8777 7950
rect 8715 7932 8789 7948
rect 8816 7944 8829 7958
rect 8844 7944 8860 7960
rect 8906 7955 8917 7968
rect 8699 7910 8700 7926
rect 8715 7910 8728 7932
rect 8743 7910 8773 7932
rect 8816 7928 8878 7944
rect 8906 7937 8917 7953
rect 8922 7948 8932 7968
rect 8942 7948 8956 7968
rect 8959 7955 8968 7968
rect 8984 7955 8993 7968
rect 8922 7937 8956 7948
rect 8959 7937 8968 7953
rect 8984 7937 8993 7953
rect 9000 7948 9010 7968
rect 9020 7948 9034 7968
rect 9035 7955 9046 7968
rect 9000 7937 9034 7948
rect 9035 7937 9046 7953
rect 9092 7944 9108 7960
rect 9115 7958 9145 8010
rect 9179 8006 9180 8013
rect 9164 7998 9180 8006
rect 9151 7966 9164 7985
rect 9179 7966 9209 7982
rect 9151 7950 9225 7966
rect 9151 7948 9164 7950
rect 9179 7948 9213 7950
rect 8816 7926 8829 7928
rect 8844 7926 8878 7928
rect 8816 7910 8878 7926
rect 8922 7921 8938 7924
rect 9000 7921 9030 7932
rect 9078 7928 9124 7944
rect 9151 7932 9225 7948
rect 9078 7926 9112 7928
rect 9077 7910 9124 7926
rect 9151 7910 9164 7932
rect 9179 7910 9209 7932
rect 9236 7910 9237 7926
rect 9252 7910 9265 8070
rect 7496 7902 7531 7910
rect 7496 7876 7497 7902
rect 7504 7876 7531 7902
rect 7439 7858 7469 7872
rect 7496 7868 7531 7876
rect 7533 7902 7574 7910
rect 7533 7876 7548 7902
rect 7555 7876 7574 7902
rect 7638 7898 7700 7910
rect 7712 7898 7787 7910
rect 7845 7898 7920 7910
rect 7932 7898 7963 7910
rect 7969 7898 8004 7910
rect 7638 7896 7800 7898
rect 7533 7868 7574 7876
rect 7656 7872 7669 7896
rect 7684 7894 7699 7896
rect 7496 7858 7525 7868
rect 7539 7858 7568 7868
rect 7583 7858 7613 7872
rect 7656 7858 7699 7872
rect 7723 7869 7730 7876
rect 7733 7872 7800 7896
rect 7832 7896 8004 7898
rect 7802 7874 7830 7878
rect 7832 7874 7912 7896
rect 7933 7894 7948 7896
rect 7802 7872 7912 7874
rect 7733 7868 7912 7872
rect 7706 7858 7736 7868
rect 7738 7858 7891 7868
rect 7899 7858 7929 7868
rect 7933 7858 7963 7872
rect 7991 7858 8004 7896
rect 8076 7902 8111 7910
rect 8076 7876 8077 7902
rect 8084 7876 8111 7902
rect 8019 7858 8049 7872
rect 8076 7868 8111 7876
rect 8113 7902 8154 7910
rect 8113 7876 8128 7902
rect 8135 7876 8154 7902
rect 8218 7898 8280 7910
rect 8292 7898 8367 7910
rect 8425 7898 8500 7910
rect 8512 7898 8543 7910
rect 8549 7898 8584 7910
rect 8218 7896 8380 7898
rect 8113 7868 8154 7876
rect 8236 7872 8249 7896
rect 8264 7894 8279 7896
rect 8076 7858 8077 7868
rect 8092 7858 8105 7868
rect 8119 7858 8120 7868
rect 8135 7858 8148 7868
rect 8163 7858 8193 7872
rect 8236 7858 8279 7872
rect 8303 7869 8310 7876
rect 8313 7872 8380 7896
rect 8412 7896 8584 7898
rect 8382 7874 8410 7878
rect 8412 7874 8492 7896
rect 8513 7894 8528 7896
rect 8382 7872 8492 7874
rect 8313 7868 8492 7872
rect 8286 7858 8316 7868
rect 8318 7858 8471 7868
rect 8479 7858 8509 7868
rect 8513 7858 8543 7872
rect 8571 7858 8584 7896
rect 8656 7902 8691 7910
rect 8656 7876 8657 7902
rect 8664 7876 8691 7902
rect 8599 7858 8629 7872
rect 8656 7868 8691 7876
rect 8693 7902 8734 7910
rect 8693 7876 8708 7902
rect 8715 7876 8734 7902
rect 8798 7898 8860 7910
rect 8872 7898 8947 7910
rect 9005 7898 9080 7910
rect 9092 7898 9123 7910
rect 9129 7898 9164 7910
rect 8798 7896 8960 7898
rect 8693 7868 8734 7876
rect 8816 7872 8829 7896
rect 8844 7894 8859 7896
rect 8656 7858 8657 7868
rect 8672 7858 8685 7868
rect 8699 7858 8700 7868
rect 8715 7858 8728 7868
rect 8743 7858 8773 7872
rect 8816 7858 8859 7872
rect 8883 7869 8890 7876
rect 8893 7872 8960 7896
rect 8992 7896 9164 7898
rect 8962 7874 8990 7878
rect 8992 7874 9072 7896
rect 9093 7894 9108 7896
rect 8962 7872 9072 7874
rect 8893 7868 9072 7872
rect 8866 7858 8896 7868
rect 8898 7858 9051 7868
rect 9059 7858 9089 7868
rect 9093 7858 9123 7872
rect 9151 7858 9164 7896
rect 9236 7902 9271 7910
rect 9236 7876 9237 7902
rect 9244 7876 9271 7902
rect 9179 7858 9209 7872
rect 9236 7868 9271 7876
rect 9236 7858 9237 7868
rect 9252 7858 9265 7868
rect -1 7852 9265 7858
rect 0 7844 9265 7852
rect 15 7814 28 7844
rect 43 7826 73 7844
rect 116 7830 130 7844
rect 166 7830 386 7844
rect 117 7828 130 7830
rect 83 7816 98 7828
rect 80 7814 102 7816
rect 107 7814 137 7828
rect 198 7826 351 7830
rect 180 7814 372 7826
rect 415 7814 445 7828
rect 451 7814 464 7844
rect 479 7826 509 7844
rect 552 7814 565 7844
rect 595 7814 608 7844
rect 623 7826 653 7844
rect 696 7830 710 7844
rect 746 7830 966 7844
rect 697 7828 710 7830
rect 663 7816 678 7828
rect 660 7814 682 7816
rect 687 7814 717 7828
rect 778 7826 931 7830
rect 760 7814 952 7826
rect 995 7814 1025 7828
rect 1031 7814 1044 7844
rect 1059 7826 1089 7844
rect 1132 7814 1145 7844
rect 1175 7814 1188 7844
rect 1203 7826 1233 7844
rect 1276 7830 1290 7844
rect 1326 7830 1546 7844
rect 1277 7828 1290 7830
rect 1243 7816 1258 7828
rect 1240 7814 1262 7816
rect 1267 7814 1297 7828
rect 1358 7826 1511 7830
rect 1340 7814 1532 7826
rect 1575 7814 1605 7828
rect 1611 7814 1624 7844
rect 1639 7826 1669 7844
rect 1712 7814 1725 7844
rect 1755 7814 1768 7844
rect 1783 7830 1813 7844
rect 1856 7830 1899 7844
rect 1906 7830 2126 7844
rect 2133 7830 2163 7844
rect 1823 7816 1838 7828
rect 1857 7816 1870 7830
rect 1938 7826 2091 7830
rect 1820 7814 1842 7816
rect 1920 7814 2112 7826
rect 2191 7814 2204 7844
rect 2219 7830 2249 7844
rect 2286 7814 2305 7844
rect 2320 7814 2326 7844
rect 2335 7814 2348 7844
rect 2363 7830 2393 7844
rect 2436 7830 2479 7844
rect 2486 7830 2706 7844
rect 2713 7830 2743 7844
rect 2403 7816 2418 7828
rect 2437 7816 2450 7830
rect 2518 7826 2671 7830
rect 2400 7814 2422 7816
rect 2500 7814 2692 7826
rect 2771 7814 2784 7844
rect 2799 7830 2829 7844
rect 2866 7814 2885 7844
rect 2900 7814 2906 7844
rect 2915 7814 2928 7844
rect 2943 7830 2973 7844
rect 3016 7830 3059 7844
rect 3066 7830 3286 7844
rect 3293 7830 3323 7844
rect 2983 7816 2998 7828
rect 3017 7816 3030 7830
rect 3098 7826 3251 7830
rect 2980 7814 3002 7816
rect 3080 7814 3272 7826
rect 3351 7814 3364 7844
rect 3379 7830 3409 7844
rect 3446 7814 3465 7844
rect 3480 7814 3486 7844
rect 3495 7814 3508 7844
rect 3523 7830 3553 7844
rect 3596 7830 3639 7844
rect 3646 7830 3866 7844
rect 3873 7830 3903 7844
rect 3563 7816 3578 7828
rect 3597 7816 3610 7830
rect 3678 7826 3831 7830
rect 3560 7814 3582 7816
rect 3660 7814 3852 7826
rect 3931 7814 3944 7844
rect 3959 7830 3989 7844
rect 4026 7814 4045 7844
rect 4060 7814 4066 7844
rect 4075 7814 4088 7844
rect 4103 7830 4133 7844
rect 4176 7830 4219 7844
rect 4226 7830 4446 7844
rect 4453 7830 4483 7844
rect 4143 7816 4158 7828
rect 4177 7816 4190 7830
rect 4258 7826 4411 7830
rect 4140 7814 4162 7816
rect 4240 7814 4432 7826
rect 4511 7814 4524 7844
rect 4539 7830 4569 7844
rect 4606 7814 4625 7844
rect 4640 7814 4646 7844
rect 4655 7814 4668 7844
rect 4683 7830 4713 7844
rect 4756 7830 4799 7844
rect 4806 7830 5026 7844
rect 5033 7830 5063 7844
rect 4723 7816 4738 7828
rect 4757 7816 4770 7830
rect 4838 7826 4991 7830
rect 4720 7814 4742 7816
rect 4820 7814 5012 7826
rect 5091 7814 5104 7844
rect 5119 7830 5149 7844
rect 5186 7814 5205 7844
rect 5220 7814 5226 7844
rect 5235 7814 5248 7844
rect 5263 7830 5293 7844
rect 5336 7830 5379 7844
rect 5386 7830 5606 7844
rect 5613 7830 5643 7844
rect 5303 7816 5318 7828
rect 5337 7816 5350 7830
rect 5418 7826 5571 7830
rect 5300 7814 5322 7816
rect 5400 7814 5592 7826
rect 5671 7814 5684 7844
rect 5699 7830 5729 7844
rect 5766 7814 5785 7844
rect 5800 7814 5806 7844
rect 5815 7814 5828 7844
rect 5843 7830 5873 7844
rect 5916 7830 5959 7844
rect 5966 7830 6186 7844
rect 6193 7830 6223 7844
rect 5883 7816 5898 7828
rect 5917 7816 5930 7830
rect 5998 7826 6151 7830
rect 5880 7814 5902 7816
rect 5980 7814 6172 7826
rect 6251 7814 6264 7844
rect 6279 7830 6309 7844
rect 6346 7814 6365 7844
rect 6380 7814 6386 7844
rect 6395 7814 6408 7844
rect 6423 7830 6453 7844
rect 6496 7830 6539 7844
rect 6546 7830 6766 7844
rect 6773 7830 6803 7844
rect 6463 7816 6478 7828
rect 6497 7816 6510 7830
rect 6578 7826 6731 7830
rect 6460 7814 6482 7816
rect 6560 7814 6752 7826
rect 6831 7814 6844 7844
rect 6859 7830 6889 7844
rect 6926 7814 6945 7844
rect 6960 7814 6966 7844
rect 6975 7814 6988 7844
rect 7003 7830 7033 7844
rect 7076 7830 7119 7844
rect 7126 7830 7346 7844
rect 7353 7830 7383 7844
rect 7043 7816 7058 7828
rect 7077 7816 7090 7830
rect 7158 7826 7311 7830
rect 7040 7814 7062 7816
rect 7140 7814 7332 7826
rect 7411 7814 7424 7844
rect 7439 7830 7469 7844
rect 7506 7814 7525 7844
rect 7540 7814 7546 7844
rect 7555 7814 7568 7844
rect 7583 7826 7613 7844
rect 7656 7830 7670 7844
rect 7706 7830 7926 7844
rect 7657 7828 7670 7830
rect 7623 7816 7638 7828
rect 7620 7814 7642 7816
rect 7647 7814 7677 7828
rect 7738 7826 7891 7830
rect 7720 7814 7912 7826
rect 7955 7814 7985 7828
rect 7991 7814 8004 7844
rect 8019 7826 8049 7844
rect 8092 7814 8105 7844
rect 8135 7814 8148 7844
rect 8163 7826 8193 7844
rect 8236 7830 8250 7844
rect 8286 7830 8506 7844
rect 8237 7828 8250 7830
rect 8203 7816 8218 7828
rect 8200 7814 8222 7816
rect 8227 7814 8257 7828
rect 8318 7826 8471 7830
rect 8300 7814 8492 7826
rect 8535 7814 8565 7828
rect 8571 7814 8584 7844
rect 8599 7826 8629 7844
rect 8672 7814 8685 7844
rect 8715 7814 8728 7844
rect 8743 7826 8773 7844
rect 8816 7830 8830 7844
rect 8866 7830 9086 7844
rect 8817 7828 8830 7830
rect 8783 7816 8798 7828
rect 8780 7814 8802 7816
rect 8807 7814 8837 7828
rect 8898 7826 9051 7830
rect 8880 7814 9072 7826
rect 9115 7814 9145 7828
rect 9151 7814 9164 7844
rect 9179 7826 9209 7844
rect 9252 7814 9265 7844
rect 0 7800 9265 7814
rect 15 7696 28 7800
rect 73 7778 74 7788
rect 89 7778 102 7788
rect 73 7774 102 7778
rect 107 7774 137 7800
rect 155 7786 171 7788
rect 243 7786 296 7800
rect 244 7784 308 7786
rect 351 7784 366 7800
rect 415 7797 445 7800
rect 415 7794 451 7797
rect 381 7786 397 7788
rect 155 7774 170 7778
rect 73 7772 170 7774
rect 198 7772 366 7784
rect 382 7774 397 7778
rect 415 7775 454 7794
rect 473 7788 480 7789
rect 479 7781 480 7788
rect 463 7778 464 7781
rect 479 7778 492 7781
rect 415 7774 445 7775
rect 454 7774 460 7775
rect 463 7774 492 7778
rect 382 7773 492 7774
rect 382 7772 498 7773
rect 57 7764 108 7772
rect 57 7752 82 7764
rect 89 7752 108 7764
rect 139 7764 189 7772
rect 139 7756 155 7764
rect 162 7762 189 7764
rect 198 7762 419 7772
rect 162 7752 419 7762
rect 448 7764 498 7772
rect 448 7755 464 7764
rect 57 7744 108 7752
rect 155 7744 419 7752
rect 445 7752 464 7755
rect 471 7752 498 7764
rect 445 7744 498 7752
rect 73 7736 74 7744
rect 89 7736 102 7744
rect 73 7728 89 7736
rect 70 7721 89 7724
rect 70 7712 92 7721
rect 43 7702 92 7712
rect 43 7696 73 7702
rect 92 7697 97 7702
rect 15 7680 89 7696
rect 107 7688 137 7744
rect 172 7734 380 7744
rect 415 7740 460 7744
rect 463 7743 464 7744
rect 479 7743 492 7744
rect 198 7704 387 7734
rect 213 7701 387 7704
rect 206 7698 387 7701
rect 15 7678 28 7680
rect 43 7678 77 7680
rect 15 7662 89 7678
rect 116 7674 129 7688
rect 144 7674 160 7690
rect 206 7685 217 7698
rect -1 7640 0 7656
rect 15 7640 28 7662
rect 43 7640 73 7662
rect 116 7658 178 7674
rect 206 7667 217 7683
rect 222 7678 232 7698
rect 242 7678 256 7698
rect 259 7685 268 7698
rect 284 7685 293 7698
rect 222 7667 256 7678
rect 259 7667 268 7683
rect 284 7667 293 7683
rect 300 7678 310 7698
rect 320 7678 334 7698
rect 335 7685 346 7698
rect 300 7667 334 7678
rect 335 7667 346 7683
rect 392 7674 408 7690
rect 415 7688 445 7740
rect 479 7736 480 7743
rect 464 7728 480 7736
rect 451 7696 464 7715
rect 479 7696 509 7712
rect 451 7680 525 7696
rect 451 7678 464 7680
rect 479 7678 513 7680
rect 116 7656 129 7658
rect 144 7656 178 7658
rect 116 7640 178 7656
rect 222 7651 238 7654
rect 300 7651 330 7662
rect 378 7658 424 7674
rect 451 7662 525 7678
rect 378 7656 412 7658
rect 377 7640 424 7656
rect 451 7640 464 7662
rect 479 7640 509 7662
rect 536 7640 537 7656
rect 552 7640 565 7800
rect 595 7696 608 7800
rect 653 7778 654 7788
rect 669 7778 682 7788
rect 653 7774 682 7778
rect 687 7774 717 7800
rect 735 7786 751 7788
rect 823 7786 876 7800
rect 824 7784 888 7786
rect 931 7784 946 7800
rect 995 7797 1025 7800
rect 995 7794 1031 7797
rect 961 7786 977 7788
rect 735 7774 750 7778
rect 653 7772 750 7774
rect 778 7772 946 7784
rect 962 7774 977 7778
rect 995 7775 1034 7794
rect 1053 7788 1060 7789
rect 1059 7781 1060 7788
rect 1043 7778 1044 7781
rect 1059 7778 1072 7781
rect 995 7774 1025 7775
rect 1034 7774 1040 7775
rect 1043 7774 1072 7778
rect 962 7773 1072 7774
rect 962 7772 1078 7773
rect 637 7764 688 7772
rect 637 7752 662 7764
rect 669 7752 688 7764
rect 719 7764 769 7772
rect 719 7756 735 7764
rect 742 7762 769 7764
rect 778 7762 999 7772
rect 742 7752 999 7762
rect 1028 7764 1078 7772
rect 1028 7755 1044 7764
rect 637 7744 688 7752
rect 735 7744 999 7752
rect 1025 7752 1044 7755
rect 1051 7752 1078 7764
rect 1025 7744 1078 7752
rect 653 7736 654 7744
rect 669 7736 682 7744
rect 653 7728 669 7736
rect 650 7721 669 7724
rect 650 7712 672 7721
rect 623 7702 672 7712
rect 623 7696 653 7702
rect 672 7697 677 7702
rect 595 7680 669 7696
rect 687 7688 717 7744
rect 752 7734 960 7744
rect 995 7740 1040 7744
rect 1043 7743 1044 7744
rect 1059 7743 1072 7744
rect 778 7704 967 7734
rect 793 7701 967 7704
rect 786 7698 967 7701
rect 595 7678 608 7680
rect 623 7678 657 7680
rect 595 7662 669 7678
rect 696 7674 709 7688
rect 724 7674 740 7690
rect 786 7685 797 7698
rect 579 7640 580 7656
rect 595 7640 608 7662
rect 623 7640 653 7662
rect 696 7658 758 7674
rect 786 7667 797 7683
rect 802 7678 812 7698
rect 822 7678 836 7698
rect 839 7685 848 7698
rect 864 7685 873 7698
rect 802 7667 836 7678
rect 839 7667 848 7683
rect 864 7667 873 7683
rect 880 7678 890 7698
rect 900 7678 914 7698
rect 915 7685 926 7698
rect 880 7667 914 7678
rect 915 7667 926 7683
rect 972 7674 988 7690
rect 995 7688 1025 7740
rect 1059 7736 1060 7743
rect 1044 7728 1060 7736
rect 1031 7696 1044 7715
rect 1059 7696 1089 7712
rect 1031 7680 1105 7696
rect 1031 7678 1044 7680
rect 1059 7678 1093 7680
rect 696 7656 709 7658
rect 724 7656 758 7658
rect 696 7640 758 7656
rect 802 7651 818 7654
rect 880 7651 910 7662
rect 958 7658 1004 7674
rect 1031 7662 1105 7678
rect 958 7656 992 7658
rect 957 7640 1004 7656
rect 1031 7640 1044 7662
rect 1059 7640 1089 7662
rect 1116 7640 1117 7656
rect 1132 7640 1145 7800
rect 1175 7696 1188 7800
rect 1233 7778 1234 7788
rect 1249 7778 1262 7788
rect 1233 7774 1262 7778
rect 1267 7774 1297 7800
rect 1315 7786 1331 7788
rect 1403 7786 1456 7800
rect 1404 7784 1468 7786
rect 1511 7784 1526 7800
rect 1575 7797 1605 7800
rect 1575 7794 1611 7797
rect 1541 7786 1557 7788
rect 1315 7774 1330 7778
rect 1233 7772 1330 7774
rect 1358 7772 1526 7784
rect 1542 7774 1557 7778
rect 1575 7775 1614 7794
rect 1633 7788 1640 7789
rect 1639 7781 1640 7788
rect 1623 7778 1624 7781
rect 1639 7778 1652 7781
rect 1575 7774 1605 7775
rect 1614 7774 1620 7775
rect 1623 7774 1652 7778
rect 1542 7773 1652 7774
rect 1542 7772 1658 7773
rect 1217 7764 1268 7772
rect 1217 7752 1242 7764
rect 1249 7752 1268 7764
rect 1299 7764 1349 7772
rect 1299 7756 1315 7764
rect 1322 7762 1349 7764
rect 1358 7762 1579 7772
rect 1322 7752 1579 7762
rect 1608 7764 1658 7772
rect 1608 7755 1624 7764
rect 1217 7744 1268 7752
rect 1315 7744 1579 7752
rect 1605 7752 1624 7755
rect 1631 7752 1658 7764
rect 1605 7744 1658 7752
rect 1233 7736 1234 7744
rect 1249 7736 1262 7744
rect 1233 7728 1249 7736
rect 1230 7721 1249 7724
rect 1230 7712 1252 7721
rect 1203 7702 1252 7712
rect 1203 7696 1233 7702
rect 1252 7697 1257 7702
rect 1175 7680 1249 7696
rect 1267 7688 1297 7744
rect 1332 7734 1540 7744
rect 1575 7740 1620 7744
rect 1623 7743 1624 7744
rect 1639 7743 1652 7744
rect 1358 7704 1547 7734
rect 1373 7701 1547 7704
rect 1366 7698 1547 7701
rect 1175 7678 1188 7680
rect 1203 7678 1237 7680
rect 1175 7662 1249 7678
rect 1276 7674 1289 7688
rect 1304 7674 1320 7690
rect 1366 7685 1377 7698
rect 1159 7640 1160 7656
rect 1175 7640 1188 7662
rect 1203 7640 1233 7662
rect 1276 7658 1338 7674
rect 1366 7667 1377 7683
rect 1382 7678 1392 7698
rect 1402 7678 1416 7698
rect 1419 7685 1428 7698
rect 1444 7685 1453 7698
rect 1382 7667 1416 7678
rect 1419 7667 1428 7683
rect 1444 7667 1453 7683
rect 1460 7678 1470 7698
rect 1480 7678 1494 7698
rect 1495 7685 1506 7698
rect 1460 7667 1494 7678
rect 1495 7667 1506 7683
rect 1552 7674 1568 7690
rect 1575 7688 1605 7740
rect 1639 7736 1640 7743
rect 1624 7728 1640 7736
rect 1611 7696 1624 7715
rect 1639 7696 1669 7712
rect 1611 7680 1685 7696
rect 1611 7678 1624 7680
rect 1639 7678 1673 7680
rect 1276 7656 1289 7658
rect 1304 7656 1338 7658
rect 1276 7640 1338 7656
rect 1382 7651 1398 7654
rect 1460 7651 1490 7662
rect 1538 7658 1584 7674
rect 1611 7662 1685 7678
rect 1538 7656 1572 7658
rect 1537 7640 1584 7656
rect 1611 7640 1624 7662
rect 1639 7640 1669 7662
rect 1696 7640 1697 7656
rect 1712 7640 1725 7800
rect 1755 7696 1768 7800
rect 1820 7796 1842 7800
rect 1813 7774 1842 7788
rect 1895 7774 1911 7788
rect 1949 7784 1955 7786
rect 1962 7784 2070 7800
rect 2077 7784 2083 7786
rect 2091 7784 2106 7800
rect 2172 7794 2191 7797
rect 1813 7772 1911 7774
rect 1938 7772 2106 7784
rect 2121 7774 2137 7788
rect 2172 7775 2194 7794
rect 2204 7788 2220 7789
rect 2203 7786 2220 7788
rect 2204 7781 2220 7786
rect 2194 7774 2200 7775
rect 2203 7774 2232 7781
rect 2121 7773 2232 7774
rect 2121 7772 2238 7773
rect 1797 7764 1848 7772
rect 1895 7764 1929 7772
rect 1797 7752 1822 7764
rect 1829 7752 1848 7764
rect 1902 7762 1929 7764
rect 1938 7762 2159 7772
rect 2194 7769 2200 7772
rect 1902 7758 2159 7762
rect 1797 7744 1848 7752
rect 1895 7744 2159 7758
rect 2203 7764 2238 7772
rect 1813 7736 1842 7744
rect 1813 7730 1830 7736
rect 1813 7728 1847 7730
rect 1895 7728 1911 7744
rect 1912 7734 2120 7744
rect 2121 7734 2137 7744
rect 2185 7740 2200 7755
rect 2203 7752 2204 7764
rect 2211 7752 2238 7764
rect 2203 7744 2238 7752
rect 2203 7743 2232 7744
rect 1923 7730 2137 7734
rect 1938 7728 2137 7730
rect 2172 7730 2185 7740
rect 2203 7730 2220 7743
rect 2172 7728 2220 7730
rect 1814 7724 1847 7728
rect 1810 7722 1847 7724
rect 1810 7721 1877 7722
rect 1810 7716 1841 7721
rect 1847 7716 1877 7721
rect 1810 7712 1877 7716
rect 1783 7709 1877 7712
rect 1783 7702 1832 7709
rect 1783 7696 1813 7702
rect 1832 7697 1837 7702
rect 1755 7680 1829 7696
rect 1841 7688 1877 7709
rect 1938 7704 2127 7728
rect 2172 7727 2219 7728
rect 2185 7722 2219 7727
rect 1953 7701 2127 7704
rect 1946 7698 2127 7701
rect 2155 7721 2219 7722
rect 1755 7678 1768 7680
rect 1783 7678 1817 7680
rect 1755 7662 1829 7678
rect 1739 7640 1740 7656
rect 1755 7640 1768 7662
rect 1783 7646 1813 7662
rect 1841 7640 1847 7688
rect 1850 7682 1869 7688
rect 1884 7682 1914 7690
rect 1850 7674 1914 7682
rect 1850 7658 1930 7674
rect 1946 7667 2008 7698
rect 2024 7667 2086 7698
rect 2155 7696 2204 7721
rect 2219 7696 2249 7712
rect 2118 7682 2148 7690
rect 2155 7688 2265 7696
rect 2118 7674 2163 7682
rect 1850 7656 1869 7658
rect 1884 7656 1930 7658
rect 1850 7640 1930 7656
rect 1957 7654 1992 7667
rect 2033 7664 2070 7667
rect 2033 7662 2075 7664
rect 1962 7651 1992 7654
rect 1971 7647 1978 7651
rect 1978 7646 1979 7647
rect 1937 7640 1947 7646
rect -7 7632 34 7640
rect -7 7606 8 7632
rect 15 7606 34 7632
rect 98 7628 160 7640
rect 172 7628 247 7640
rect 305 7628 380 7640
rect 392 7628 423 7640
rect 429 7628 464 7640
rect 98 7626 260 7628
rect -7 7598 34 7606
rect 116 7602 129 7626
rect 144 7624 159 7626
rect -1 7588 0 7598
rect 15 7588 28 7598
rect 43 7588 73 7602
rect 116 7588 159 7602
rect 183 7599 190 7606
rect 193 7602 260 7626
rect 292 7626 464 7628
rect 262 7604 290 7608
rect 292 7604 372 7626
rect 393 7624 408 7626
rect 262 7602 372 7604
rect 193 7598 372 7602
rect 166 7588 196 7598
rect 198 7588 351 7598
rect 359 7588 389 7598
rect 393 7588 423 7602
rect 451 7588 464 7626
rect 536 7632 571 7640
rect 536 7606 537 7632
rect 544 7606 571 7632
rect 479 7588 509 7602
rect 536 7598 571 7606
rect 573 7632 614 7640
rect 573 7606 588 7632
rect 595 7606 614 7632
rect 678 7628 740 7640
rect 752 7628 827 7640
rect 885 7628 960 7640
rect 972 7628 1003 7640
rect 1009 7628 1044 7640
rect 678 7626 840 7628
rect 573 7598 614 7606
rect 696 7602 709 7626
rect 724 7624 739 7626
rect 536 7588 537 7598
rect 552 7588 565 7598
rect 579 7588 580 7598
rect 595 7588 608 7598
rect 623 7588 653 7602
rect 696 7588 739 7602
rect 763 7599 770 7606
rect 773 7602 840 7626
rect 872 7626 1044 7628
rect 842 7604 870 7608
rect 872 7604 952 7626
rect 973 7624 988 7626
rect 842 7602 952 7604
rect 773 7598 952 7602
rect 746 7588 776 7598
rect 778 7588 931 7598
rect 939 7588 969 7598
rect 973 7588 1003 7602
rect 1031 7588 1044 7626
rect 1116 7632 1151 7640
rect 1116 7606 1117 7632
rect 1124 7606 1151 7632
rect 1059 7588 1089 7602
rect 1116 7598 1151 7606
rect 1153 7632 1194 7640
rect 1153 7606 1168 7632
rect 1175 7606 1194 7632
rect 1258 7628 1320 7640
rect 1332 7628 1407 7640
rect 1465 7628 1540 7640
rect 1552 7628 1583 7640
rect 1589 7628 1624 7640
rect 1258 7626 1420 7628
rect 1153 7598 1194 7606
rect 1276 7602 1289 7626
rect 1304 7624 1319 7626
rect 1116 7588 1117 7598
rect 1132 7588 1145 7598
rect 1159 7588 1160 7598
rect 1175 7588 1188 7598
rect 1203 7588 1233 7602
rect 1276 7588 1319 7602
rect 1343 7599 1350 7606
rect 1353 7602 1420 7626
rect 1452 7626 1624 7628
rect 1422 7604 1450 7608
rect 1452 7604 1532 7626
rect 1553 7624 1568 7626
rect 1422 7602 1532 7604
rect 1353 7598 1532 7602
rect 1326 7588 1356 7598
rect 1358 7588 1511 7598
rect 1519 7588 1549 7598
rect 1553 7588 1583 7602
rect 1611 7588 1624 7626
rect 1696 7632 1731 7640
rect 1696 7606 1697 7632
rect 1704 7606 1731 7632
rect 1639 7588 1669 7602
rect 1696 7598 1731 7606
rect 1733 7632 1774 7640
rect 1733 7606 1748 7632
rect 1755 7606 1774 7632
rect 1838 7628 1869 7640
rect 1884 7628 1987 7640
rect 1999 7630 2025 7656
rect 2040 7651 2070 7662
rect 2102 7658 2164 7674
rect 2102 7656 2148 7658
rect 2102 7640 2164 7656
rect 2176 7640 2182 7688
rect 2185 7680 2265 7688
rect 2185 7678 2204 7680
rect 2219 7678 2253 7680
rect 2185 7662 2265 7678
rect 2185 7640 2204 7662
rect 2219 7646 2249 7662
rect 2277 7656 2283 7730
rect 2286 7656 2305 7800
rect 2320 7656 2326 7800
rect 2335 7730 2348 7800
rect 2400 7796 2422 7800
rect 2393 7774 2422 7788
rect 2475 7774 2491 7788
rect 2529 7784 2535 7786
rect 2542 7784 2650 7800
rect 2657 7784 2663 7786
rect 2671 7784 2686 7800
rect 2752 7794 2771 7797
rect 2393 7772 2491 7774
rect 2518 7772 2686 7784
rect 2701 7774 2717 7788
rect 2752 7775 2774 7794
rect 2784 7788 2800 7789
rect 2783 7786 2800 7788
rect 2784 7781 2800 7786
rect 2774 7774 2780 7775
rect 2783 7774 2812 7781
rect 2701 7773 2812 7774
rect 2701 7772 2818 7773
rect 2377 7764 2428 7772
rect 2475 7764 2509 7772
rect 2377 7752 2402 7764
rect 2409 7752 2428 7764
rect 2482 7762 2509 7764
rect 2518 7762 2739 7772
rect 2774 7769 2780 7772
rect 2482 7758 2739 7762
rect 2377 7744 2428 7752
rect 2475 7744 2739 7758
rect 2783 7764 2818 7772
rect 2329 7696 2348 7730
rect 2393 7736 2422 7744
rect 2393 7730 2410 7736
rect 2393 7728 2427 7730
rect 2475 7728 2491 7744
rect 2492 7734 2700 7744
rect 2701 7734 2717 7744
rect 2765 7740 2780 7755
rect 2783 7752 2784 7764
rect 2791 7752 2818 7764
rect 2783 7744 2818 7752
rect 2783 7743 2812 7744
rect 2503 7730 2717 7734
rect 2518 7728 2717 7730
rect 2752 7730 2765 7740
rect 2783 7730 2800 7743
rect 2752 7728 2800 7730
rect 2394 7724 2427 7728
rect 2390 7722 2427 7724
rect 2390 7721 2457 7722
rect 2390 7716 2421 7721
rect 2427 7716 2457 7721
rect 2390 7712 2457 7716
rect 2363 7709 2457 7712
rect 2363 7702 2412 7709
rect 2363 7696 2393 7702
rect 2412 7697 2417 7702
rect 2329 7680 2409 7696
rect 2421 7688 2457 7709
rect 2518 7704 2707 7728
rect 2752 7727 2799 7728
rect 2765 7722 2799 7727
rect 2533 7701 2707 7704
rect 2526 7698 2707 7701
rect 2735 7721 2799 7722
rect 2329 7678 2348 7680
rect 2363 7678 2397 7680
rect 2329 7662 2409 7678
rect 2329 7656 2348 7662
rect 2045 7630 2148 7640
rect 1999 7628 2148 7630
rect 2169 7628 2204 7640
rect 1838 7626 2000 7628
rect 1850 7606 1869 7626
rect 1884 7624 1914 7626
rect 1733 7598 1774 7606
rect 1856 7602 1869 7606
rect 1921 7610 2000 7626
rect 2032 7626 2204 7628
rect 2032 7610 2111 7626
rect 2118 7624 2148 7626
rect 1696 7588 1697 7598
rect 1712 7588 1725 7598
rect 1739 7588 1740 7598
rect 1755 7588 1768 7598
rect 1783 7588 1813 7602
rect 1856 7588 1899 7602
rect 1921 7598 2111 7610
rect 2176 7606 2182 7626
rect 1906 7588 1936 7598
rect 1937 7588 2095 7598
rect 2099 7588 2129 7598
rect 2133 7588 2163 7602
rect 2191 7588 2204 7626
rect 2276 7640 2305 7656
rect 2319 7640 2348 7656
rect 2363 7646 2393 7662
rect 2421 7640 2427 7688
rect 2430 7682 2449 7688
rect 2464 7682 2494 7690
rect 2430 7674 2494 7682
rect 2430 7658 2510 7674
rect 2526 7667 2588 7698
rect 2604 7667 2666 7698
rect 2735 7696 2784 7721
rect 2799 7696 2829 7712
rect 2698 7682 2728 7690
rect 2735 7688 2845 7696
rect 2698 7674 2743 7682
rect 2430 7656 2449 7658
rect 2464 7656 2510 7658
rect 2430 7640 2510 7656
rect 2537 7654 2572 7667
rect 2613 7664 2650 7667
rect 2613 7662 2655 7664
rect 2542 7651 2572 7654
rect 2551 7647 2558 7651
rect 2558 7646 2559 7647
rect 2517 7640 2527 7646
rect 2276 7632 2311 7640
rect 2276 7606 2277 7632
rect 2284 7606 2311 7632
rect 2219 7588 2249 7602
rect 2276 7598 2311 7606
rect 2313 7632 2354 7640
rect 2313 7606 2328 7632
rect 2335 7606 2354 7632
rect 2418 7628 2449 7640
rect 2464 7628 2567 7640
rect 2579 7630 2605 7656
rect 2620 7651 2650 7662
rect 2682 7658 2744 7674
rect 2682 7656 2728 7658
rect 2682 7640 2744 7656
rect 2756 7640 2762 7688
rect 2765 7680 2845 7688
rect 2765 7678 2784 7680
rect 2799 7678 2833 7680
rect 2765 7662 2845 7678
rect 2765 7640 2784 7662
rect 2799 7646 2829 7662
rect 2857 7656 2863 7730
rect 2866 7656 2885 7800
rect 2900 7656 2906 7800
rect 2915 7730 2928 7800
rect 2980 7796 3002 7800
rect 2973 7774 3002 7788
rect 3055 7774 3071 7788
rect 3109 7784 3115 7786
rect 3122 7784 3230 7800
rect 3237 7784 3243 7786
rect 3251 7784 3266 7800
rect 3332 7794 3351 7797
rect 2973 7772 3071 7774
rect 3098 7772 3266 7784
rect 3281 7774 3297 7788
rect 3332 7775 3354 7794
rect 3364 7788 3380 7789
rect 3363 7786 3380 7788
rect 3364 7781 3380 7786
rect 3354 7774 3360 7775
rect 3363 7774 3392 7781
rect 3281 7773 3392 7774
rect 3281 7772 3398 7773
rect 2957 7764 3008 7772
rect 3055 7764 3089 7772
rect 2957 7752 2982 7764
rect 2989 7752 3008 7764
rect 3062 7762 3089 7764
rect 3098 7762 3319 7772
rect 3354 7769 3360 7772
rect 3062 7758 3319 7762
rect 2957 7744 3008 7752
rect 3055 7744 3319 7758
rect 3363 7764 3398 7772
rect 2909 7696 2928 7730
rect 2973 7736 3002 7744
rect 2973 7730 2990 7736
rect 2973 7728 3007 7730
rect 3055 7728 3071 7744
rect 3072 7734 3280 7744
rect 3281 7734 3297 7744
rect 3345 7740 3360 7755
rect 3363 7752 3364 7764
rect 3371 7752 3398 7764
rect 3363 7744 3398 7752
rect 3363 7743 3392 7744
rect 3083 7730 3297 7734
rect 3098 7728 3297 7730
rect 3332 7730 3345 7740
rect 3363 7730 3380 7743
rect 3332 7728 3380 7730
rect 2974 7724 3007 7728
rect 2970 7722 3007 7724
rect 2970 7721 3037 7722
rect 2970 7716 3001 7721
rect 3007 7716 3037 7721
rect 2970 7712 3037 7716
rect 2943 7709 3037 7712
rect 2943 7702 2992 7709
rect 2943 7696 2973 7702
rect 2992 7697 2997 7702
rect 2909 7680 2989 7696
rect 3001 7688 3037 7709
rect 3098 7704 3287 7728
rect 3332 7727 3379 7728
rect 3345 7722 3379 7727
rect 3113 7701 3287 7704
rect 3106 7698 3287 7701
rect 3315 7721 3379 7722
rect 2909 7678 2928 7680
rect 2943 7678 2977 7680
rect 2909 7662 2989 7678
rect 2909 7656 2928 7662
rect 2625 7630 2728 7640
rect 2579 7628 2728 7630
rect 2749 7628 2784 7640
rect 2418 7626 2580 7628
rect 2430 7606 2449 7626
rect 2464 7624 2494 7626
rect 2313 7598 2354 7606
rect 2436 7602 2449 7606
rect 2501 7610 2580 7626
rect 2612 7626 2784 7628
rect 2612 7610 2691 7626
rect 2698 7624 2728 7626
rect 2276 7588 2305 7598
rect 2319 7588 2348 7598
rect 2363 7588 2393 7602
rect 2436 7588 2479 7602
rect 2501 7598 2691 7610
rect 2756 7606 2762 7626
rect 2486 7588 2516 7598
rect 2517 7588 2675 7598
rect 2679 7588 2709 7598
rect 2713 7588 2743 7602
rect 2771 7588 2784 7626
rect 2856 7640 2885 7656
rect 2899 7640 2928 7656
rect 2943 7646 2973 7662
rect 3001 7640 3007 7688
rect 3010 7682 3029 7688
rect 3044 7682 3074 7690
rect 3010 7674 3074 7682
rect 3010 7658 3090 7674
rect 3106 7667 3168 7698
rect 3184 7667 3246 7698
rect 3315 7696 3364 7721
rect 3379 7696 3409 7712
rect 3278 7682 3308 7690
rect 3315 7688 3425 7696
rect 3278 7674 3323 7682
rect 3010 7656 3029 7658
rect 3044 7656 3090 7658
rect 3010 7640 3090 7656
rect 3117 7654 3152 7667
rect 3193 7664 3230 7667
rect 3193 7662 3235 7664
rect 3122 7651 3152 7654
rect 3131 7647 3138 7651
rect 3138 7646 3139 7647
rect 3097 7640 3107 7646
rect 2856 7632 2891 7640
rect 2856 7606 2857 7632
rect 2864 7606 2891 7632
rect 2799 7588 2829 7602
rect 2856 7598 2891 7606
rect 2893 7632 2934 7640
rect 2893 7606 2908 7632
rect 2915 7606 2934 7632
rect 2998 7628 3029 7640
rect 3044 7628 3147 7640
rect 3159 7630 3185 7656
rect 3200 7651 3230 7662
rect 3262 7658 3324 7674
rect 3262 7656 3308 7658
rect 3262 7640 3324 7656
rect 3336 7640 3342 7688
rect 3345 7680 3425 7688
rect 3345 7678 3364 7680
rect 3379 7678 3413 7680
rect 3345 7662 3425 7678
rect 3345 7640 3364 7662
rect 3379 7646 3409 7662
rect 3437 7656 3443 7730
rect 3446 7656 3465 7800
rect 3480 7656 3486 7800
rect 3495 7730 3508 7800
rect 3560 7796 3582 7800
rect 3553 7774 3582 7788
rect 3635 7774 3651 7788
rect 3689 7784 3695 7786
rect 3702 7784 3810 7800
rect 3817 7784 3823 7786
rect 3831 7784 3846 7800
rect 3912 7794 3931 7797
rect 3553 7772 3651 7774
rect 3678 7772 3846 7784
rect 3861 7774 3877 7788
rect 3912 7775 3934 7794
rect 3944 7788 3960 7789
rect 3943 7786 3960 7788
rect 3944 7781 3960 7786
rect 3934 7774 3940 7775
rect 3943 7774 3972 7781
rect 3861 7773 3972 7774
rect 3861 7772 3978 7773
rect 3537 7764 3588 7772
rect 3635 7764 3669 7772
rect 3537 7752 3562 7764
rect 3569 7752 3588 7764
rect 3642 7762 3669 7764
rect 3678 7762 3899 7772
rect 3934 7769 3940 7772
rect 3642 7758 3899 7762
rect 3537 7744 3588 7752
rect 3635 7744 3899 7758
rect 3943 7764 3978 7772
rect 3489 7696 3508 7730
rect 3553 7736 3582 7744
rect 3553 7730 3570 7736
rect 3553 7728 3587 7730
rect 3635 7728 3651 7744
rect 3652 7734 3860 7744
rect 3861 7734 3877 7744
rect 3925 7740 3940 7755
rect 3943 7752 3944 7764
rect 3951 7752 3978 7764
rect 3943 7744 3978 7752
rect 3943 7743 3972 7744
rect 3663 7730 3877 7734
rect 3678 7728 3877 7730
rect 3912 7730 3925 7740
rect 3943 7730 3960 7743
rect 3912 7728 3960 7730
rect 3554 7724 3587 7728
rect 3550 7722 3587 7724
rect 3550 7721 3617 7722
rect 3550 7716 3581 7721
rect 3587 7716 3617 7721
rect 3550 7712 3617 7716
rect 3523 7709 3617 7712
rect 3523 7702 3572 7709
rect 3523 7696 3553 7702
rect 3572 7697 3577 7702
rect 3489 7680 3569 7696
rect 3581 7688 3617 7709
rect 3678 7704 3867 7728
rect 3912 7727 3959 7728
rect 3925 7722 3959 7727
rect 3693 7701 3867 7704
rect 3686 7698 3867 7701
rect 3895 7721 3959 7722
rect 3489 7678 3508 7680
rect 3523 7678 3557 7680
rect 3489 7662 3569 7678
rect 3489 7656 3508 7662
rect 3205 7630 3308 7640
rect 3159 7628 3308 7630
rect 3329 7628 3364 7640
rect 2998 7626 3160 7628
rect 3010 7606 3029 7626
rect 3044 7624 3074 7626
rect 2893 7598 2934 7606
rect 3016 7602 3029 7606
rect 3081 7610 3160 7626
rect 3192 7626 3364 7628
rect 3192 7610 3271 7626
rect 3278 7624 3308 7626
rect 2856 7588 2885 7598
rect 2899 7588 2928 7598
rect 2943 7588 2973 7602
rect 3016 7588 3059 7602
rect 3081 7598 3271 7610
rect 3336 7606 3342 7626
rect 3066 7588 3096 7598
rect 3097 7588 3255 7598
rect 3259 7588 3289 7598
rect 3293 7588 3323 7602
rect 3351 7588 3364 7626
rect 3436 7640 3465 7656
rect 3479 7640 3508 7656
rect 3523 7646 3553 7662
rect 3581 7640 3587 7688
rect 3590 7682 3609 7688
rect 3624 7682 3654 7690
rect 3590 7674 3654 7682
rect 3590 7658 3670 7674
rect 3686 7667 3748 7698
rect 3764 7667 3826 7698
rect 3895 7696 3944 7721
rect 3959 7696 3989 7712
rect 3858 7682 3888 7690
rect 3895 7688 4005 7696
rect 3858 7674 3903 7682
rect 3590 7656 3609 7658
rect 3624 7656 3670 7658
rect 3590 7640 3670 7656
rect 3697 7654 3732 7667
rect 3773 7664 3810 7667
rect 3773 7662 3815 7664
rect 3702 7651 3732 7654
rect 3711 7647 3718 7651
rect 3718 7646 3719 7647
rect 3677 7640 3687 7646
rect 3436 7632 3471 7640
rect 3436 7606 3437 7632
rect 3444 7606 3471 7632
rect 3379 7588 3409 7602
rect 3436 7598 3471 7606
rect 3473 7632 3514 7640
rect 3473 7606 3488 7632
rect 3495 7606 3514 7632
rect 3578 7628 3609 7640
rect 3624 7628 3727 7640
rect 3739 7630 3765 7656
rect 3780 7651 3810 7662
rect 3842 7658 3904 7674
rect 3842 7656 3888 7658
rect 3842 7640 3904 7656
rect 3916 7640 3922 7688
rect 3925 7680 4005 7688
rect 3925 7678 3944 7680
rect 3959 7678 3993 7680
rect 3925 7662 4005 7678
rect 3925 7640 3944 7662
rect 3959 7646 3989 7662
rect 4017 7656 4023 7730
rect 4026 7656 4045 7800
rect 4060 7656 4066 7800
rect 4075 7730 4088 7800
rect 4140 7796 4162 7800
rect 4133 7774 4162 7788
rect 4215 7774 4231 7788
rect 4269 7784 4275 7786
rect 4282 7784 4390 7800
rect 4397 7784 4403 7786
rect 4411 7784 4426 7800
rect 4492 7794 4511 7797
rect 4133 7772 4231 7774
rect 4258 7772 4426 7784
rect 4441 7774 4457 7788
rect 4492 7775 4514 7794
rect 4524 7788 4540 7789
rect 4523 7786 4540 7788
rect 4524 7781 4540 7786
rect 4514 7774 4520 7775
rect 4523 7774 4552 7781
rect 4441 7773 4552 7774
rect 4441 7772 4558 7773
rect 4117 7764 4168 7772
rect 4215 7764 4249 7772
rect 4117 7752 4142 7764
rect 4149 7752 4168 7764
rect 4222 7762 4249 7764
rect 4258 7762 4479 7772
rect 4514 7769 4520 7772
rect 4222 7758 4479 7762
rect 4117 7744 4168 7752
rect 4215 7744 4479 7758
rect 4523 7764 4558 7772
rect 4069 7696 4088 7730
rect 4133 7736 4162 7744
rect 4133 7730 4150 7736
rect 4133 7728 4167 7730
rect 4215 7728 4231 7744
rect 4232 7734 4440 7744
rect 4441 7734 4457 7744
rect 4505 7740 4520 7755
rect 4523 7752 4524 7764
rect 4531 7752 4558 7764
rect 4523 7744 4558 7752
rect 4523 7743 4552 7744
rect 4243 7730 4457 7734
rect 4258 7728 4457 7730
rect 4492 7730 4505 7740
rect 4523 7730 4540 7743
rect 4492 7728 4540 7730
rect 4134 7724 4167 7728
rect 4130 7722 4167 7724
rect 4130 7721 4197 7722
rect 4130 7716 4161 7721
rect 4167 7716 4197 7721
rect 4130 7712 4197 7716
rect 4103 7709 4197 7712
rect 4103 7702 4152 7709
rect 4103 7696 4133 7702
rect 4152 7697 4157 7702
rect 4069 7680 4149 7696
rect 4161 7688 4197 7709
rect 4258 7704 4447 7728
rect 4492 7727 4539 7728
rect 4505 7722 4539 7727
rect 4273 7701 4447 7704
rect 4266 7698 4447 7701
rect 4475 7721 4539 7722
rect 4069 7678 4088 7680
rect 4103 7678 4137 7680
rect 4069 7662 4149 7678
rect 4069 7656 4088 7662
rect 3785 7630 3888 7640
rect 3739 7628 3888 7630
rect 3909 7628 3944 7640
rect 3578 7626 3740 7628
rect 3590 7606 3609 7626
rect 3624 7624 3654 7626
rect 3473 7598 3514 7606
rect 3596 7602 3609 7606
rect 3661 7610 3740 7626
rect 3772 7626 3944 7628
rect 3772 7610 3851 7626
rect 3858 7624 3888 7626
rect 3436 7588 3465 7598
rect 3479 7588 3508 7598
rect 3523 7588 3553 7602
rect 3596 7588 3639 7602
rect 3661 7598 3851 7610
rect 3916 7606 3922 7626
rect 3646 7588 3676 7598
rect 3677 7588 3835 7598
rect 3839 7588 3869 7598
rect 3873 7588 3903 7602
rect 3931 7588 3944 7626
rect 4016 7640 4045 7656
rect 4059 7640 4088 7656
rect 4103 7646 4133 7662
rect 4161 7640 4167 7688
rect 4170 7682 4189 7688
rect 4204 7682 4234 7690
rect 4170 7674 4234 7682
rect 4170 7658 4250 7674
rect 4266 7667 4328 7698
rect 4344 7667 4406 7698
rect 4475 7696 4524 7721
rect 4539 7696 4569 7712
rect 4438 7682 4468 7690
rect 4475 7688 4585 7696
rect 4438 7674 4483 7682
rect 4170 7656 4189 7658
rect 4204 7656 4250 7658
rect 4170 7640 4250 7656
rect 4277 7654 4312 7667
rect 4353 7664 4390 7667
rect 4353 7662 4395 7664
rect 4282 7651 4312 7654
rect 4291 7647 4298 7651
rect 4298 7646 4299 7647
rect 4257 7640 4267 7646
rect 4016 7632 4051 7640
rect 4016 7606 4017 7632
rect 4024 7606 4051 7632
rect 3959 7588 3989 7602
rect 4016 7598 4051 7606
rect 4053 7632 4094 7640
rect 4053 7606 4068 7632
rect 4075 7606 4094 7632
rect 4158 7628 4189 7640
rect 4204 7628 4307 7640
rect 4319 7630 4345 7656
rect 4360 7651 4390 7662
rect 4422 7658 4484 7674
rect 4422 7656 4468 7658
rect 4422 7640 4484 7656
rect 4496 7640 4502 7688
rect 4505 7680 4585 7688
rect 4505 7678 4524 7680
rect 4539 7678 4573 7680
rect 4505 7662 4585 7678
rect 4505 7640 4524 7662
rect 4539 7646 4569 7662
rect 4597 7656 4603 7730
rect 4606 7656 4625 7800
rect 4640 7656 4646 7800
rect 4655 7730 4668 7800
rect 4720 7796 4742 7800
rect 4713 7774 4742 7788
rect 4795 7774 4811 7788
rect 4849 7784 4855 7786
rect 4862 7784 4970 7800
rect 4977 7784 4983 7786
rect 4991 7784 5006 7800
rect 5072 7794 5091 7797
rect 4713 7772 4811 7774
rect 4838 7772 5006 7784
rect 5021 7774 5037 7788
rect 5072 7775 5094 7794
rect 5104 7788 5120 7789
rect 5103 7786 5120 7788
rect 5104 7781 5120 7786
rect 5094 7774 5100 7775
rect 5103 7774 5132 7781
rect 5021 7773 5132 7774
rect 5021 7772 5138 7773
rect 4697 7764 4748 7772
rect 4795 7764 4829 7772
rect 4697 7752 4722 7764
rect 4729 7752 4748 7764
rect 4802 7762 4829 7764
rect 4838 7762 5059 7772
rect 5094 7769 5100 7772
rect 4802 7758 5059 7762
rect 4697 7744 4748 7752
rect 4795 7744 5059 7758
rect 5103 7764 5138 7772
rect 4649 7696 4668 7730
rect 4713 7736 4742 7744
rect 4713 7730 4730 7736
rect 4713 7728 4747 7730
rect 4795 7728 4811 7744
rect 4812 7734 5020 7744
rect 5021 7734 5037 7744
rect 5085 7740 5100 7755
rect 5103 7752 5104 7764
rect 5111 7752 5138 7764
rect 5103 7744 5138 7752
rect 5103 7743 5132 7744
rect 4823 7730 5037 7734
rect 4838 7728 5037 7730
rect 5072 7730 5085 7740
rect 5103 7730 5120 7743
rect 5072 7728 5120 7730
rect 4714 7724 4747 7728
rect 4710 7722 4747 7724
rect 4710 7721 4777 7722
rect 4710 7716 4741 7721
rect 4747 7716 4777 7721
rect 4710 7712 4777 7716
rect 4683 7709 4777 7712
rect 4683 7702 4732 7709
rect 4683 7696 4713 7702
rect 4732 7697 4737 7702
rect 4649 7680 4729 7696
rect 4741 7688 4777 7709
rect 4838 7704 5027 7728
rect 5072 7727 5119 7728
rect 5085 7722 5119 7727
rect 4853 7701 5027 7704
rect 4846 7698 5027 7701
rect 5055 7721 5119 7722
rect 4649 7678 4668 7680
rect 4683 7678 4717 7680
rect 4649 7662 4729 7678
rect 4649 7656 4668 7662
rect 4365 7630 4468 7640
rect 4319 7628 4468 7630
rect 4489 7628 4524 7640
rect 4158 7626 4320 7628
rect 4170 7606 4189 7626
rect 4204 7624 4234 7626
rect 4053 7598 4094 7606
rect 4176 7602 4189 7606
rect 4241 7610 4320 7626
rect 4352 7626 4524 7628
rect 4352 7610 4431 7626
rect 4438 7624 4468 7626
rect 4016 7588 4045 7598
rect 4059 7588 4088 7598
rect 4103 7588 4133 7602
rect 4176 7588 4219 7602
rect 4241 7598 4431 7610
rect 4496 7606 4502 7626
rect 4226 7588 4256 7598
rect 4257 7588 4415 7598
rect 4419 7588 4449 7598
rect 4453 7588 4483 7602
rect 4511 7588 4524 7626
rect 4596 7640 4625 7656
rect 4639 7640 4668 7656
rect 4683 7646 4713 7662
rect 4741 7640 4747 7688
rect 4750 7682 4769 7688
rect 4784 7682 4814 7690
rect 4750 7674 4814 7682
rect 4750 7658 4830 7674
rect 4846 7667 4908 7698
rect 4924 7667 4986 7698
rect 5055 7696 5104 7721
rect 5119 7696 5149 7712
rect 5018 7682 5048 7690
rect 5055 7688 5165 7696
rect 5018 7674 5063 7682
rect 4750 7656 4769 7658
rect 4784 7656 4830 7658
rect 4750 7640 4830 7656
rect 4857 7654 4892 7667
rect 4933 7664 4970 7667
rect 4933 7662 4975 7664
rect 4862 7651 4892 7654
rect 4871 7647 4878 7651
rect 4878 7646 4879 7647
rect 4837 7640 4847 7646
rect 4596 7632 4631 7640
rect 4596 7606 4597 7632
rect 4604 7606 4631 7632
rect 4539 7588 4569 7602
rect 4596 7598 4631 7606
rect 4633 7632 4674 7640
rect 4633 7606 4648 7632
rect 4655 7606 4674 7632
rect 4738 7628 4769 7640
rect 4784 7628 4887 7640
rect 4899 7630 4925 7656
rect 4940 7651 4970 7662
rect 5002 7658 5064 7674
rect 5002 7656 5048 7658
rect 5002 7640 5064 7656
rect 5076 7640 5082 7688
rect 5085 7680 5165 7688
rect 5085 7678 5104 7680
rect 5119 7678 5153 7680
rect 5085 7662 5165 7678
rect 5085 7640 5104 7662
rect 5119 7646 5149 7662
rect 5177 7656 5183 7730
rect 5186 7656 5205 7800
rect 5220 7656 5226 7800
rect 5235 7730 5248 7800
rect 5300 7796 5322 7800
rect 5293 7774 5322 7788
rect 5375 7774 5391 7788
rect 5429 7784 5435 7786
rect 5442 7784 5550 7800
rect 5557 7784 5563 7786
rect 5571 7784 5586 7800
rect 5652 7794 5671 7797
rect 5293 7772 5391 7774
rect 5418 7772 5586 7784
rect 5601 7774 5617 7788
rect 5652 7775 5674 7794
rect 5684 7788 5700 7789
rect 5683 7786 5700 7788
rect 5684 7781 5700 7786
rect 5674 7774 5680 7775
rect 5683 7774 5712 7781
rect 5601 7773 5712 7774
rect 5601 7772 5718 7773
rect 5277 7764 5328 7772
rect 5375 7764 5409 7772
rect 5277 7752 5302 7764
rect 5309 7752 5328 7764
rect 5382 7762 5409 7764
rect 5418 7762 5639 7772
rect 5674 7769 5680 7772
rect 5382 7758 5639 7762
rect 5277 7744 5328 7752
rect 5375 7744 5639 7758
rect 5683 7764 5718 7772
rect 5229 7696 5248 7730
rect 5293 7736 5322 7744
rect 5293 7730 5310 7736
rect 5293 7728 5327 7730
rect 5375 7728 5391 7744
rect 5392 7734 5600 7744
rect 5601 7734 5617 7744
rect 5665 7740 5680 7755
rect 5683 7752 5684 7764
rect 5691 7752 5718 7764
rect 5683 7744 5718 7752
rect 5683 7743 5712 7744
rect 5403 7730 5617 7734
rect 5418 7728 5617 7730
rect 5652 7730 5665 7740
rect 5683 7730 5700 7743
rect 5652 7728 5700 7730
rect 5294 7724 5327 7728
rect 5290 7722 5327 7724
rect 5290 7721 5357 7722
rect 5290 7716 5321 7721
rect 5327 7716 5357 7721
rect 5290 7712 5357 7716
rect 5263 7709 5357 7712
rect 5263 7702 5312 7709
rect 5263 7696 5293 7702
rect 5312 7697 5317 7702
rect 5229 7680 5309 7696
rect 5321 7688 5357 7709
rect 5418 7704 5607 7728
rect 5652 7727 5699 7728
rect 5665 7722 5699 7727
rect 5433 7701 5607 7704
rect 5426 7698 5607 7701
rect 5635 7721 5699 7722
rect 5229 7678 5248 7680
rect 5263 7678 5297 7680
rect 5229 7662 5309 7678
rect 5229 7656 5248 7662
rect 4945 7630 5048 7640
rect 4899 7628 5048 7630
rect 5069 7628 5104 7640
rect 4738 7626 4900 7628
rect 4750 7606 4769 7626
rect 4784 7624 4814 7626
rect 4633 7598 4674 7606
rect 4756 7602 4769 7606
rect 4821 7610 4900 7626
rect 4932 7626 5104 7628
rect 4932 7610 5011 7626
rect 5018 7624 5048 7626
rect 4596 7588 4625 7598
rect 4639 7588 4668 7598
rect 4683 7588 4713 7602
rect 4756 7588 4799 7602
rect 4821 7598 5011 7610
rect 5076 7606 5082 7626
rect 4806 7588 4836 7598
rect 4837 7588 4995 7598
rect 4999 7588 5029 7598
rect 5033 7588 5063 7602
rect 5091 7588 5104 7626
rect 5176 7640 5205 7656
rect 5219 7640 5248 7656
rect 5263 7646 5293 7662
rect 5321 7640 5327 7688
rect 5330 7682 5349 7688
rect 5364 7682 5394 7690
rect 5330 7674 5394 7682
rect 5330 7658 5410 7674
rect 5426 7667 5488 7698
rect 5504 7667 5566 7698
rect 5635 7696 5684 7721
rect 5699 7696 5729 7712
rect 5598 7682 5628 7690
rect 5635 7688 5745 7696
rect 5598 7674 5643 7682
rect 5330 7656 5349 7658
rect 5364 7656 5410 7658
rect 5330 7640 5410 7656
rect 5437 7654 5472 7667
rect 5513 7664 5550 7667
rect 5513 7662 5555 7664
rect 5442 7651 5472 7654
rect 5451 7647 5458 7651
rect 5458 7646 5459 7647
rect 5417 7640 5427 7646
rect 5176 7632 5211 7640
rect 5176 7606 5177 7632
rect 5184 7606 5211 7632
rect 5119 7588 5149 7602
rect 5176 7598 5211 7606
rect 5213 7632 5254 7640
rect 5213 7606 5228 7632
rect 5235 7606 5254 7632
rect 5318 7628 5349 7640
rect 5364 7628 5467 7640
rect 5479 7630 5505 7656
rect 5520 7651 5550 7662
rect 5582 7658 5644 7674
rect 5582 7656 5628 7658
rect 5582 7640 5644 7656
rect 5656 7640 5662 7688
rect 5665 7680 5745 7688
rect 5665 7678 5684 7680
rect 5699 7678 5733 7680
rect 5665 7662 5745 7678
rect 5665 7640 5684 7662
rect 5699 7646 5729 7662
rect 5757 7656 5763 7730
rect 5766 7656 5785 7800
rect 5800 7656 5806 7800
rect 5815 7730 5828 7800
rect 5880 7796 5902 7800
rect 5873 7774 5902 7788
rect 5955 7774 5971 7788
rect 6009 7784 6015 7786
rect 6022 7784 6130 7800
rect 6137 7784 6143 7786
rect 6151 7784 6166 7800
rect 6232 7794 6251 7797
rect 5873 7772 5971 7774
rect 5998 7772 6166 7784
rect 6181 7774 6197 7788
rect 6232 7775 6254 7794
rect 6264 7788 6280 7789
rect 6263 7786 6280 7788
rect 6264 7781 6280 7786
rect 6254 7774 6260 7775
rect 6263 7774 6292 7781
rect 6181 7773 6292 7774
rect 6181 7772 6298 7773
rect 5857 7764 5908 7772
rect 5955 7764 5989 7772
rect 5857 7752 5882 7764
rect 5889 7752 5908 7764
rect 5962 7762 5989 7764
rect 5998 7762 6219 7772
rect 6254 7769 6260 7772
rect 5962 7758 6219 7762
rect 5857 7744 5908 7752
rect 5955 7744 6219 7758
rect 6263 7764 6298 7772
rect 5809 7696 5828 7730
rect 5873 7736 5902 7744
rect 5873 7730 5890 7736
rect 5873 7728 5907 7730
rect 5955 7728 5971 7744
rect 5972 7734 6180 7744
rect 6181 7734 6197 7744
rect 6245 7740 6260 7755
rect 6263 7752 6264 7764
rect 6271 7752 6298 7764
rect 6263 7744 6298 7752
rect 6263 7743 6292 7744
rect 5983 7730 6197 7734
rect 5998 7728 6197 7730
rect 6232 7730 6245 7740
rect 6263 7730 6280 7743
rect 6232 7728 6280 7730
rect 5874 7724 5907 7728
rect 5870 7722 5907 7724
rect 5870 7721 5937 7722
rect 5870 7716 5901 7721
rect 5907 7716 5937 7721
rect 5870 7712 5937 7716
rect 5843 7709 5937 7712
rect 5843 7702 5892 7709
rect 5843 7696 5873 7702
rect 5892 7697 5897 7702
rect 5809 7680 5889 7696
rect 5901 7688 5937 7709
rect 5998 7704 6187 7728
rect 6232 7727 6279 7728
rect 6245 7722 6279 7727
rect 6013 7701 6187 7704
rect 6006 7698 6187 7701
rect 6215 7721 6279 7722
rect 5809 7678 5828 7680
rect 5843 7678 5877 7680
rect 5809 7662 5889 7678
rect 5809 7656 5828 7662
rect 5525 7630 5628 7640
rect 5479 7628 5628 7630
rect 5649 7628 5684 7640
rect 5318 7626 5480 7628
rect 5330 7606 5349 7626
rect 5364 7624 5394 7626
rect 5213 7598 5254 7606
rect 5336 7602 5349 7606
rect 5401 7610 5480 7626
rect 5512 7626 5684 7628
rect 5512 7610 5591 7626
rect 5598 7624 5628 7626
rect 5176 7588 5205 7598
rect 5219 7588 5248 7598
rect 5263 7588 5293 7602
rect 5336 7588 5379 7602
rect 5401 7598 5591 7610
rect 5656 7606 5662 7626
rect 5386 7588 5416 7598
rect 5417 7588 5575 7598
rect 5579 7588 5609 7598
rect 5613 7588 5643 7602
rect 5671 7588 5684 7626
rect 5756 7640 5785 7656
rect 5799 7640 5828 7656
rect 5843 7646 5873 7662
rect 5901 7640 5907 7688
rect 5910 7682 5929 7688
rect 5944 7682 5974 7690
rect 5910 7674 5974 7682
rect 5910 7658 5990 7674
rect 6006 7667 6068 7698
rect 6084 7667 6146 7698
rect 6215 7696 6264 7721
rect 6279 7696 6309 7712
rect 6178 7682 6208 7690
rect 6215 7688 6325 7696
rect 6178 7674 6223 7682
rect 5910 7656 5929 7658
rect 5944 7656 5990 7658
rect 5910 7640 5990 7656
rect 6017 7654 6052 7667
rect 6093 7664 6130 7667
rect 6093 7662 6135 7664
rect 6022 7651 6052 7654
rect 6031 7647 6038 7651
rect 6038 7646 6039 7647
rect 5997 7640 6007 7646
rect 5756 7632 5791 7640
rect 5756 7606 5757 7632
rect 5764 7606 5791 7632
rect 5699 7588 5729 7602
rect 5756 7598 5791 7606
rect 5793 7632 5834 7640
rect 5793 7606 5808 7632
rect 5815 7606 5834 7632
rect 5898 7628 5929 7640
rect 5944 7628 6047 7640
rect 6059 7630 6085 7656
rect 6100 7651 6130 7662
rect 6162 7658 6224 7674
rect 6162 7656 6208 7658
rect 6162 7640 6224 7656
rect 6236 7640 6242 7688
rect 6245 7680 6325 7688
rect 6245 7678 6264 7680
rect 6279 7678 6313 7680
rect 6245 7662 6325 7678
rect 6245 7640 6264 7662
rect 6279 7646 6309 7662
rect 6337 7656 6343 7730
rect 6346 7656 6365 7800
rect 6380 7656 6386 7800
rect 6395 7730 6408 7800
rect 6460 7796 6482 7800
rect 6453 7774 6482 7788
rect 6535 7774 6551 7788
rect 6589 7784 6595 7786
rect 6602 7784 6710 7800
rect 6717 7784 6723 7786
rect 6731 7784 6746 7800
rect 6812 7794 6831 7797
rect 6453 7772 6551 7774
rect 6578 7772 6746 7784
rect 6761 7774 6777 7788
rect 6812 7775 6834 7794
rect 6844 7788 6860 7789
rect 6843 7786 6860 7788
rect 6844 7781 6860 7786
rect 6834 7774 6840 7775
rect 6843 7774 6872 7781
rect 6761 7773 6872 7774
rect 6761 7772 6878 7773
rect 6437 7764 6488 7772
rect 6535 7764 6569 7772
rect 6437 7752 6462 7764
rect 6469 7752 6488 7764
rect 6542 7762 6569 7764
rect 6578 7762 6799 7772
rect 6834 7769 6840 7772
rect 6542 7758 6799 7762
rect 6437 7744 6488 7752
rect 6535 7744 6799 7758
rect 6843 7764 6878 7772
rect 6389 7696 6408 7730
rect 6453 7736 6482 7744
rect 6453 7730 6470 7736
rect 6453 7728 6487 7730
rect 6535 7728 6551 7744
rect 6552 7734 6760 7744
rect 6761 7734 6777 7744
rect 6825 7740 6840 7755
rect 6843 7752 6844 7764
rect 6851 7752 6878 7764
rect 6843 7744 6878 7752
rect 6843 7743 6872 7744
rect 6563 7730 6777 7734
rect 6578 7728 6777 7730
rect 6812 7730 6825 7740
rect 6843 7730 6860 7743
rect 6812 7728 6860 7730
rect 6454 7724 6487 7728
rect 6450 7722 6487 7724
rect 6450 7721 6517 7722
rect 6450 7716 6481 7721
rect 6487 7716 6517 7721
rect 6450 7712 6517 7716
rect 6423 7709 6517 7712
rect 6423 7702 6472 7709
rect 6423 7696 6453 7702
rect 6472 7697 6477 7702
rect 6389 7680 6469 7696
rect 6481 7688 6517 7709
rect 6578 7704 6767 7728
rect 6812 7727 6859 7728
rect 6825 7722 6859 7727
rect 6593 7701 6767 7704
rect 6586 7698 6767 7701
rect 6795 7721 6859 7722
rect 6389 7678 6408 7680
rect 6423 7678 6457 7680
rect 6389 7662 6469 7678
rect 6389 7656 6408 7662
rect 6105 7630 6208 7640
rect 6059 7628 6208 7630
rect 6229 7628 6264 7640
rect 5898 7626 6060 7628
rect 5910 7606 5929 7626
rect 5944 7624 5974 7626
rect 5793 7598 5834 7606
rect 5916 7602 5929 7606
rect 5981 7610 6060 7626
rect 6092 7626 6264 7628
rect 6092 7610 6171 7626
rect 6178 7624 6208 7626
rect 5756 7588 5785 7598
rect 5799 7588 5828 7598
rect 5843 7588 5873 7602
rect 5916 7588 5959 7602
rect 5981 7598 6171 7610
rect 6236 7606 6242 7626
rect 5966 7588 5996 7598
rect 5997 7588 6155 7598
rect 6159 7588 6189 7598
rect 6193 7588 6223 7602
rect 6251 7588 6264 7626
rect 6336 7640 6365 7656
rect 6379 7640 6408 7656
rect 6423 7646 6453 7662
rect 6481 7640 6487 7688
rect 6490 7682 6509 7688
rect 6524 7682 6554 7690
rect 6490 7674 6554 7682
rect 6490 7658 6570 7674
rect 6586 7667 6648 7698
rect 6664 7667 6726 7698
rect 6795 7696 6844 7721
rect 6859 7696 6889 7712
rect 6758 7682 6788 7690
rect 6795 7688 6905 7696
rect 6758 7674 6803 7682
rect 6490 7656 6509 7658
rect 6524 7656 6570 7658
rect 6490 7640 6570 7656
rect 6597 7654 6632 7667
rect 6673 7664 6710 7667
rect 6673 7662 6715 7664
rect 6602 7651 6632 7654
rect 6611 7647 6618 7651
rect 6618 7646 6619 7647
rect 6577 7640 6587 7646
rect 6336 7632 6371 7640
rect 6336 7606 6337 7632
rect 6344 7606 6371 7632
rect 6279 7588 6309 7602
rect 6336 7598 6371 7606
rect 6373 7632 6414 7640
rect 6373 7606 6388 7632
rect 6395 7606 6414 7632
rect 6478 7628 6509 7640
rect 6524 7628 6627 7640
rect 6639 7630 6665 7656
rect 6680 7651 6710 7662
rect 6742 7658 6804 7674
rect 6742 7656 6788 7658
rect 6742 7640 6804 7656
rect 6816 7640 6822 7688
rect 6825 7680 6905 7688
rect 6825 7678 6844 7680
rect 6859 7678 6893 7680
rect 6825 7662 6905 7678
rect 6825 7640 6844 7662
rect 6859 7646 6889 7662
rect 6917 7656 6923 7730
rect 6926 7656 6945 7800
rect 6960 7656 6966 7800
rect 6975 7730 6988 7800
rect 7040 7796 7062 7800
rect 7033 7774 7062 7788
rect 7115 7774 7131 7788
rect 7169 7784 7175 7786
rect 7182 7784 7290 7800
rect 7297 7784 7303 7786
rect 7311 7784 7326 7800
rect 7392 7794 7411 7797
rect 7033 7772 7131 7774
rect 7158 7772 7326 7784
rect 7341 7774 7357 7788
rect 7392 7775 7414 7794
rect 7424 7788 7440 7789
rect 7423 7786 7440 7788
rect 7424 7781 7440 7786
rect 7414 7774 7420 7775
rect 7423 7774 7452 7781
rect 7341 7773 7452 7774
rect 7341 7772 7458 7773
rect 7017 7764 7068 7772
rect 7115 7764 7149 7772
rect 7017 7752 7042 7764
rect 7049 7752 7068 7764
rect 7122 7762 7149 7764
rect 7158 7762 7379 7772
rect 7414 7769 7420 7772
rect 7122 7758 7379 7762
rect 7017 7744 7068 7752
rect 7115 7744 7379 7758
rect 7423 7764 7458 7772
rect 6969 7696 6988 7730
rect 7033 7736 7062 7744
rect 7033 7730 7050 7736
rect 7033 7728 7067 7730
rect 7115 7728 7131 7744
rect 7132 7734 7340 7744
rect 7341 7734 7357 7744
rect 7405 7740 7420 7755
rect 7423 7752 7424 7764
rect 7431 7752 7458 7764
rect 7423 7744 7458 7752
rect 7423 7743 7452 7744
rect 7143 7730 7357 7734
rect 7158 7728 7357 7730
rect 7392 7730 7405 7740
rect 7423 7730 7440 7743
rect 7392 7728 7440 7730
rect 7034 7724 7067 7728
rect 7030 7722 7067 7724
rect 7030 7721 7097 7722
rect 7030 7716 7061 7721
rect 7067 7716 7097 7721
rect 7030 7712 7097 7716
rect 7003 7709 7097 7712
rect 7003 7702 7052 7709
rect 7003 7696 7033 7702
rect 7052 7697 7057 7702
rect 6969 7680 7049 7696
rect 7061 7688 7097 7709
rect 7158 7704 7347 7728
rect 7392 7727 7439 7728
rect 7405 7722 7439 7727
rect 7173 7701 7347 7704
rect 7166 7698 7347 7701
rect 7375 7721 7439 7722
rect 6969 7678 6988 7680
rect 7003 7678 7037 7680
rect 6969 7662 7049 7678
rect 6969 7656 6988 7662
rect 6685 7630 6788 7640
rect 6639 7628 6788 7630
rect 6809 7628 6844 7640
rect 6478 7626 6640 7628
rect 6490 7606 6509 7626
rect 6524 7624 6554 7626
rect 6373 7598 6414 7606
rect 6496 7602 6509 7606
rect 6561 7610 6640 7626
rect 6672 7626 6844 7628
rect 6672 7610 6751 7626
rect 6758 7624 6788 7626
rect 6336 7588 6365 7598
rect 6379 7588 6408 7598
rect 6423 7588 6453 7602
rect 6496 7588 6539 7602
rect 6561 7598 6751 7610
rect 6816 7606 6822 7626
rect 6546 7588 6576 7598
rect 6577 7588 6735 7598
rect 6739 7588 6769 7598
rect 6773 7588 6803 7602
rect 6831 7588 6844 7626
rect 6916 7640 6945 7656
rect 6959 7640 6988 7656
rect 7003 7646 7033 7662
rect 7061 7640 7067 7688
rect 7070 7682 7089 7688
rect 7104 7682 7134 7690
rect 7070 7674 7134 7682
rect 7070 7658 7150 7674
rect 7166 7667 7228 7698
rect 7244 7667 7306 7698
rect 7375 7696 7424 7721
rect 7439 7696 7469 7712
rect 7338 7682 7368 7690
rect 7375 7688 7485 7696
rect 7338 7674 7383 7682
rect 7070 7656 7089 7658
rect 7104 7656 7150 7658
rect 7070 7640 7150 7656
rect 7177 7654 7212 7667
rect 7253 7664 7290 7667
rect 7253 7662 7295 7664
rect 7182 7651 7212 7654
rect 7191 7647 7198 7651
rect 7198 7646 7199 7647
rect 7157 7640 7167 7646
rect 6916 7632 6951 7640
rect 6916 7606 6917 7632
rect 6924 7606 6951 7632
rect 6859 7588 6889 7602
rect 6916 7598 6951 7606
rect 6953 7632 6994 7640
rect 6953 7606 6968 7632
rect 6975 7606 6994 7632
rect 7058 7628 7089 7640
rect 7104 7628 7207 7640
rect 7219 7630 7245 7656
rect 7260 7651 7290 7662
rect 7322 7658 7384 7674
rect 7322 7656 7368 7658
rect 7322 7640 7384 7656
rect 7396 7640 7402 7688
rect 7405 7680 7485 7688
rect 7405 7678 7424 7680
rect 7439 7678 7473 7680
rect 7405 7662 7485 7678
rect 7405 7640 7424 7662
rect 7439 7646 7469 7662
rect 7497 7656 7503 7730
rect 7506 7656 7525 7800
rect 7540 7656 7546 7800
rect 7555 7730 7568 7800
rect 7613 7778 7614 7788
rect 7629 7778 7642 7788
rect 7613 7774 7642 7778
rect 7647 7774 7677 7800
rect 7695 7786 7711 7788
rect 7783 7786 7836 7800
rect 7784 7784 7848 7786
rect 7891 7784 7906 7800
rect 7955 7797 7985 7800
rect 7955 7794 7991 7797
rect 7921 7786 7937 7788
rect 7695 7774 7710 7778
rect 7613 7772 7710 7774
rect 7738 7772 7906 7784
rect 7922 7774 7937 7778
rect 7955 7775 7994 7794
rect 8013 7788 8020 7789
rect 8019 7781 8020 7788
rect 8003 7778 8004 7781
rect 8019 7778 8032 7781
rect 7955 7774 7985 7775
rect 7994 7774 8000 7775
rect 8003 7774 8032 7778
rect 7922 7773 8032 7774
rect 7922 7772 8038 7773
rect 7597 7764 7648 7772
rect 7597 7752 7622 7764
rect 7629 7752 7648 7764
rect 7679 7764 7729 7772
rect 7679 7756 7695 7764
rect 7702 7762 7729 7764
rect 7738 7762 7959 7772
rect 7702 7752 7959 7762
rect 7988 7764 8038 7772
rect 7988 7755 8004 7764
rect 7597 7744 7648 7752
rect 7695 7744 7959 7752
rect 7985 7752 8004 7755
rect 8011 7752 8038 7764
rect 7985 7744 8038 7752
rect 7549 7696 7568 7730
rect 7613 7736 7614 7744
rect 7629 7736 7642 7744
rect 7613 7728 7629 7736
rect 7610 7721 7629 7724
rect 7610 7712 7632 7721
rect 7583 7702 7632 7712
rect 7583 7696 7613 7702
rect 7632 7697 7637 7702
rect 7549 7680 7629 7696
rect 7647 7688 7677 7744
rect 7712 7734 7920 7744
rect 7955 7740 8000 7744
rect 8003 7743 8004 7744
rect 8019 7743 8032 7744
rect 7738 7704 7927 7734
rect 7753 7701 7927 7704
rect 7746 7698 7927 7701
rect 7549 7678 7568 7680
rect 7583 7678 7617 7680
rect 7549 7662 7629 7678
rect 7656 7674 7669 7688
rect 7684 7674 7700 7690
rect 7746 7685 7757 7698
rect 7549 7656 7568 7662
rect 7265 7630 7368 7640
rect 7219 7628 7368 7630
rect 7389 7628 7424 7640
rect 7058 7626 7220 7628
rect 7070 7606 7089 7626
rect 7104 7624 7134 7626
rect 6953 7598 6994 7606
rect 7076 7602 7089 7606
rect 7141 7610 7220 7626
rect 7252 7626 7424 7628
rect 7252 7610 7331 7626
rect 7338 7624 7368 7626
rect 6916 7588 6945 7598
rect 6959 7588 6988 7598
rect 7003 7588 7033 7602
rect 7076 7588 7119 7602
rect 7141 7598 7331 7610
rect 7396 7606 7402 7626
rect 7126 7588 7156 7598
rect 7157 7588 7315 7598
rect 7319 7588 7349 7598
rect 7353 7588 7383 7602
rect 7411 7588 7424 7626
rect 7496 7640 7525 7656
rect 7539 7640 7568 7656
rect 7583 7640 7613 7662
rect 7656 7658 7718 7674
rect 7746 7667 7757 7683
rect 7762 7678 7772 7698
rect 7782 7678 7796 7698
rect 7799 7685 7808 7698
rect 7824 7685 7833 7698
rect 7762 7667 7796 7678
rect 7799 7667 7808 7683
rect 7824 7667 7833 7683
rect 7840 7678 7850 7698
rect 7860 7678 7874 7698
rect 7875 7685 7886 7698
rect 7840 7667 7874 7678
rect 7875 7667 7886 7683
rect 7932 7674 7948 7690
rect 7955 7688 7985 7740
rect 8019 7736 8020 7743
rect 8004 7728 8020 7736
rect 7991 7696 8004 7715
rect 8019 7696 8049 7712
rect 7991 7680 8065 7696
rect 7991 7678 8004 7680
rect 8019 7678 8053 7680
rect 7656 7656 7669 7658
rect 7684 7656 7718 7658
rect 7656 7640 7718 7656
rect 7762 7651 7778 7654
rect 7840 7651 7870 7662
rect 7918 7658 7964 7674
rect 7991 7662 8065 7678
rect 7918 7656 7952 7658
rect 7917 7640 7964 7656
rect 7991 7640 8004 7662
rect 8019 7640 8049 7662
rect 8076 7640 8077 7656
rect 8092 7640 8105 7800
rect 8135 7696 8148 7800
rect 8193 7778 8194 7788
rect 8209 7778 8222 7788
rect 8193 7774 8222 7778
rect 8227 7774 8257 7800
rect 8275 7786 8291 7788
rect 8363 7786 8416 7800
rect 8364 7784 8428 7786
rect 8471 7784 8486 7800
rect 8535 7797 8565 7800
rect 8535 7794 8571 7797
rect 8501 7786 8517 7788
rect 8275 7774 8290 7778
rect 8193 7772 8290 7774
rect 8318 7772 8486 7784
rect 8502 7774 8517 7778
rect 8535 7775 8574 7794
rect 8593 7788 8600 7789
rect 8599 7781 8600 7788
rect 8583 7778 8584 7781
rect 8599 7778 8612 7781
rect 8535 7774 8565 7775
rect 8574 7774 8580 7775
rect 8583 7774 8612 7778
rect 8502 7773 8612 7774
rect 8502 7772 8618 7773
rect 8177 7764 8228 7772
rect 8177 7752 8202 7764
rect 8209 7752 8228 7764
rect 8259 7764 8309 7772
rect 8259 7756 8275 7764
rect 8282 7762 8309 7764
rect 8318 7762 8539 7772
rect 8282 7752 8539 7762
rect 8568 7764 8618 7772
rect 8568 7755 8584 7764
rect 8177 7744 8228 7752
rect 8275 7744 8539 7752
rect 8565 7752 8584 7755
rect 8591 7752 8618 7764
rect 8565 7744 8618 7752
rect 8193 7736 8194 7744
rect 8209 7736 8222 7744
rect 8193 7728 8209 7736
rect 8190 7721 8209 7724
rect 8190 7712 8212 7721
rect 8163 7702 8212 7712
rect 8163 7696 8193 7702
rect 8212 7697 8217 7702
rect 8135 7680 8209 7696
rect 8227 7688 8257 7744
rect 8292 7734 8500 7744
rect 8535 7740 8580 7744
rect 8583 7743 8584 7744
rect 8599 7743 8612 7744
rect 8318 7704 8507 7734
rect 8333 7701 8507 7704
rect 8326 7698 8507 7701
rect 8135 7678 8148 7680
rect 8163 7678 8197 7680
rect 8135 7662 8209 7678
rect 8236 7674 8249 7688
rect 8264 7674 8280 7690
rect 8326 7685 8337 7698
rect 8119 7640 8120 7656
rect 8135 7640 8148 7662
rect 8163 7640 8193 7662
rect 8236 7658 8298 7674
rect 8326 7667 8337 7683
rect 8342 7678 8352 7698
rect 8362 7678 8376 7698
rect 8379 7685 8388 7698
rect 8404 7685 8413 7698
rect 8342 7667 8376 7678
rect 8379 7667 8388 7683
rect 8404 7667 8413 7683
rect 8420 7678 8430 7698
rect 8440 7678 8454 7698
rect 8455 7685 8466 7698
rect 8420 7667 8454 7678
rect 8455 7667 8466 7683
rect 8512 7674 8528 7690
rect 8535 7688 8565 7740
rect 8599 7736 8600 7743
rect 8584 7728 8600 7736
rect 8571 7696 8584 7715
rect 8599 7696 8629 7712
rect 8571 7680 8645 7696
rect 8571 7678 8584 7680
rect 8599 7678 8633 7680
rect 8236 7656 8249 7658
rect 8264 7656 8298 7658
rect 8236 7640 8298 7656
rect 8342 7651 8358 7654
rect 8420 7651 8450 7662
rect 8498 7658 8544 7674
rect 8571 7662 8645 7678
rect 8498 7656 8532 7658
rect 8497 7640 8544 7656
rect 8571 7640 8584 7662
rect 8599 7640 8629 7662
rect 8656 7640 8657 7656
rect 8672 7640 8685 7800
rect 8715 7696 8728 7800
rect 8773 7778 8774 7788
rect 8789 7778 8802 7788
rect 8773 7774 8802 7778
rect 8807 7774 8837 7800
rect 8855 7786 8871 7788
rect 8943 7786 8996 7800
rect 8944 7784 9008 7786
rect 9051 7784 9066 7800
rect 9115 7797 9145 7800
rect 9115 7794 9151 7797
rect 9081 7786 9097 7788
rect 8855 7774 8870 7778
rect 8773 7772 8870 7774
rect 8898 7772 9066 7784
rect 9082 7774 9097 7778
rect 9115 7775 9154 7794
rect 9173 7788 9180 7789
rect 9179 7781 9180 7788
rect 9163 7778 9164 7781
rect 9179 7778 9192 7781
rect 9115 7774 9145 7775
rect 9154 7774 9160 7775
rect 9163 7774 9192 7778
rect 9082 7773 9192 7774
rect 9082 7772 9198 7773
rect 8757 7764 8808 7772
rect 8757 7752 8782 7764
rect 8789 7752 8808 7764
rect 8839 7764 8889 7772
rect 8839 7756 8855 7764
rect 8862 7762 8889 7764
rect 8898 7762 9119 7772
rect 8862 7752 9119 7762
rect 9148 7764 9198 7772
rect 9148 7755 9164 7764
rect 8757 7744 8808 7752
rect 8855 7744 9119 7752
rect 9145 7752 9164 7755
rect 9171 7752 9198 7764
rect 9145 7744 9198 7752
rect 8773 7736 8774 7744
rect 8789 7736 8802 7744
rect 8773 7728 8789 7736
rect 8770 7721 8789 7724
rect 8770 7712 8792 7721
rect 8743 7702 8792 7712
rect 8743 7696 8773 7702
rect 8792 7697 8797 7702
rect 8715 7680 8789 7696
rect 8807 7688 8837 7744
rect 8872 7734 9080 7744
rect 9115 7740 9160 7744
rect 9163 7743 9164 7744
rect 9179 7743 9192 7744
rect 8898 7704 9087 7734
rect 8913 7701 9087 7704
rect 8906 7698 9087 7701
rect 8715 7678 8728 7680
rect 8743 7678 8777 7680
rect 8715 7662 8789 7678
rect 8816 7674 8829 7688
rect 8844 7674 8860 7690
rect 8906 7685 8917 7698
rect 8699 7640 8700 7656
rect 8715 7640 8728 7662
rect 8743 7640 8773 7662
rect 8816 7658 8878 7674
rect 8906 7667 8917 7683
rect 8922 7678 8932 7698
rect 8942 7678 8956 7698
rect 8959 7685 8968 7698
rect 8984 7685 8993 7698
rect 8922 7667 8956 7678
rect 8959 7667 8968 7683
rect 8984 7667 8993 7683
rect 9000 7678 9010 7698
rect 9020 7678 9034 7698
rect 9035 7685 9046 7698
rect 9000 7667 9034 7678
rect 9035 7667 9046 7683
rect 9092 7674 9108 7690
rect 9115 7688 9145 7740
rect 9179 7736 9180 7743
rect 9164 7728 9180 7736
rect 9151 7696 9164 7715
rect 9179 7696 9209 7712
rect 9151 7680 9225 7696
rect 9151 7678 9164 7680
rect 9179 7678 9213 7680
rect 8816 7656 8829 7658
rect 8844 7656 8878 7658
rect 8816 7640 8878 7656
rect 8922 7651 8938 7654
rect 9000 7651 9030 7662
rect 9078 7658 9124 7674
rect 9151 7662 9225 7678
rect 9078 7656 9112 7658
rect 9077 7640 9124 7656
rect 9151 7640 9164 7662
rect 9179 7640 9209 7662
rect 9236 7640 9237 7656
rect 9252 7640 9265 7800
rect 7496 7632 7531 7640
rect 7496 7606 7497 7632
rect 7504 7606 7531 7632
rect 7439 7588 7469 7602
rect 7496 7598 7531 7606
rect 7533 7632 7574 7640
rect 7533 7606 7548 7632
rect 7555 7606 7574 7632
rect 7638 7628 7700 7640
rect 7712 7628 7787 7640
rect 7845 7628 7920 7640
rect 7932 7628 7963 7640
rect 7969 7628 8004 7640
rect 7638 7626 7800 7628
rect 7533 7598 7574 7606
rect 7656 7602 7669 7626
rect 7684 7624 7699 7626
rect 7496 7588 7525 7598
rect 7539 7588 7568 7598
rect 7583 7588 7613 7602
rect 7656 7588 7699 7602
rect 7723 7599 7730 7606
rect 7733 7602 7800 7626
rect 7832 7626 8004 7628
rect 7802 7604 7830 7608
rect 7832 7604 7912 7626
rect 7933 7624 7948 7626
rect 7802 7602 7912 7604
rect 7733 7598 7912 7602
rect 7706 7588 7736 7598
rect 7738 7588 7891 7598
rect 7899 7588 7929 7598
rect 7933 7588 7963 7602
rect 7991 7588 8004 7626
rect 8076 7632 8111 7640
rect 8076 7606 8077 7632
rect 8084 7606 8111 7632
rect 8019 7588 8049 7602
rect 8076 7598 8111 7606
rect 8113 7632 8154 7640
rect 8113 7606 8128 7632
rect 8135 7606 8154 7632
rect 8218 7628 8280 7640
rect 8292 7628 8367 7640
rect 8425 7628 8500 7640
rect 8512 7628 8543 7640
rect 8549 7628 8584 7640
rect 8218 7626 8380 7628
rect 8113 7598 8154 7606
rect 8236 7602 8249 7626
rect 8264 7624 8279 7626
rect 8076 7588 8077 7598
rect 8092 7588 8105 7598
rect 8119 7588 8120 7598
rect 8135 7588 8148 7598
rect 8163 7588 8193 7602
rect 8236 7588 8279 7602
rect 8303 7599 8310 7606
rect 8313 7602 8380 7626
rect 8412 7626 8584 7628
rect 8382 7604 8410 7608
rect 8412 7604 8492 7626
rect 8513 7624 8528 7626
rect 8382 7602 8492 7604
rect 8313 7598 8492 7602
rect 8286 7588 8316 7598
rect 8318 7588 8471 7598
rect 8479 7588 8509 7598
rect 8513 7588 8543 7602
rect 8571 7588 8584 7626
rect 8656 7632 8691 7640
rect 8656 7606 8657 7632
rect 8664 7606 8691 7632
rect 8599 7588 8629 7602
rect 8656 7598 8691 7606
rect 8693 7632 8734 7640
rect 8693 7606 8708 7632
rect 8715 7606 8734 7632
rect 8798 7628 8860 7640
rect 8872 7628 8947 7640
rect 9005 7628 9080 7640
rect 9092 7628 9123 7640
rect 9129 7628 9164 7640
rect 8798 7626 8960 7628
rect 8693 7598 8734 7606
rect 8816 7602 8829 7626
rect 8844 7624 8859 7626
rect 8656 7588 8657 7598
rect 8672 7588 8685 7598
rect 8699 7588 8700 7598
rect 8715 7588 8728 7598
rect 8743 7588 8773 7602
rect 8816 7588 8859 7602
rect 8883 7599 8890 7606
rect 8893 7602 8960 7626
rect 8992 7626 9164 7628
rect 8962 7604 8990 7608
rect 8992 7604 9072 7626
rect 9093 7624 9108 7626
rect 8962 7602 9072 7604
rect 8893 7598 9072 7602
rect 8866 7588 8896 7598
rect 8898 7588 9051 7598
rect 9059 7588 9089 7598
rect 9093 7588 9123 7602
rect 9151 7588 9164 7626
rect 9236 7632 9271 7640
rect 9236 7606 9237 7632
rect 9244 7606 9271 7632
rect 9179 7588 9209 7602
rect 9236 7598 9271 7606
rect 9236 7588 9237 7598
rect 9252 7588 9265 7598
rect -1 7582 9265 7588
rect 0 7574 9265 7582
rect 15 7544 28 7574
rect 43 7556 73 7574
rect 116 7560 130 7574
rect 166 7560 386 7574
rect 117 7558 130 7560
rect 83 7546 98 7558
rect 80 7544 102 7546
rect 107 7544 137 7558
rect 198 7556 351 7560
rect 180 7544 372 7556
rect 415 7544 445 7558
rect 451 7544 464 7574
rect 479 7556 509 7574
rect 552 7544 565 7574
rect 595 7544 608 7574
rect 623 7556 653 7574
rect 696 7560 710 7574
rect 746 7560 966 7574
rect 697 7558 710 7560
rect 663 7546 678 7558
rect 660 7544 682 7546
rect 687 7544 717 7558
rect 778 7556 931 7560
rect 760 7544 952 7556
rect 995 7544 1025 7558
rect 1031 7544 1044 7574
rect 1059 7556 1089 7574
rect 1132 7544 1145 7574
rect 1175 7544 1188 7574
rect 1203 7556 1233 7574
rect 1276 7560 1290 7574
rect 1326 7560 1546 7574
rect 1277 7558 1290 7560
rect 1243 7546 1258 7558
rect 1240 7544 1262 7546
rect 1267 7544 1297 7558
rect 1358 7556 1511 7560
rect 1340 7544 1532 7556
rect 1575 7544 1605 7558
rect 1611 7544 1624 7574
rect 1639 7556 1669 7574
rect 1712 7544 1725 7574
rect 1755 7544 1768 7574
rect 1783 7560 1813 7574
rect 1856 7560 1899 7574
rect 1906 7560 2126 7574
rect 2133 7560 2163 7574
rect 1823 7546 1838 7558
rect 1857 7546 1870 7560
rect 1938 7556 2091 7560
rect 1820 7544 1842 7546
rect 1920 7544 2112 7556
rect 2191 7544 2204 7574
rect 2219 7560 2249 7574
rect 2286 7544 2305 7574
rect 2320 7544 2326 7574
rect 2335 7544 2348 7574
rect 2363 7560 2393 7574
rect 2436 7560 2479 7574
rect 2486 7560 2706 7574
rect 2713 7560 2743 7574
rect 2403 7546 2418 7558
rect 2437 7546 2450 7560
rect 2518 7556 2671 7560
rect 2400 7544 2422 7546
rect 2500 7544 2692 7556
rect 2771 7544 2784 7574
rect 2799 7560 2829 7574
rect 2866 7544 2885 7574
rect 2900 7544 2906 7574
rect 2915 7544 2928 7574
rect 2943 7560 2973 7574
rect 3016 7560 3059 7574
rect 3066 7560 3286 7574
rect 3293 7560 3323 7574
rect 2983 7546 2998 7558
rect 3017 7546 3030 7560
rect 3098 7556 3251 7560
rect 2980 7544 3002 7546
rect 3080 7544 3272 7556
rect 3351 7544 3364 7574
rect 3379 7560 3409 7574
rect 3446 7544 3465 7574
rect 3480 7544 3486 7574
rect 3495 7544 3508 7574
rect 3523 7560 3553 7574
rect 3596 7560 3639 7574
rect 3646 7560 3866 7574
rect 3873 7560 3903 7574
rect 3563 7546 3578 7558
rect 3597 7546 3610 7560
rect 3678 7556 3831 7560
rect 3560 7544 3582 7546
rect 3660 7544 3852 7556
rect 3931 7544 3944 7574
rect 3959 7560 3989 7574
rect 4026 7544 4045 7574
rect 4060 7544 4066 7574
rect 4075 7544 4088 7574
rect 4103 7560 4133 7574
rect 4176 7560 4219 7574
rect 4226 7560 4446 7574
rect 4453 7560 4483 7574
rect 4143 7546 4158 7558
rect 4177 7546 4190 7560
rect 4258 7556 4411 7560
rect 4140 7544 4162 7546
rect 4240 7544 4432 7556
rect 4511 7544 4524 7574
rect 4539 7560 4569 7574
rect 4606 7544 4625 7574
rect 4640 7544 4646 7574
rect 4655 7544 4668 7574
rect 4683 7560 4713 7574
rect 4756 7560 4799 7574
rect 4806 7560 5026 7574
rect 5033 7560 5063 7574
rect 4723 7546 4738 7558
rect 4757 7546 4770 7560
rect 4838 7556 4991 7560
rect 4720 7544 4742 7546
rect 4820 7544 5012 7556
rect 5091 7544 5104 7574
rect 5119 7560 5149 7574
rect 5186 7544 5205 7574
rect 5220 7544 5226 7574
rect 5235 7544 5248 7574
rect 5263 7560 5293 7574
rect 5336 7560 5379 7574
rect 5386 7560 5606 7574
rect 5613 7560 5643 7574
rect 5303 7546 5318 7558
rect 5337 7546 5350 7560
rect 5418 7556 5571 7560
rect 5300 7544 5322 7546
rect 5400 7544 5592 7556
rect 5671 7544 5684 7574
rect 5699 7560 5729 7574
rect 5766 7544 5785 7574
rect 5800 7544 5806 7574
rect 5815 7544 5828 7574
rect 5843 7560 5873 7574
rect 5916 7560 5959 7574
rect 5966 7560 6186 7574
rect 6193 7560 6223 7574
rect 5883 7546 5898 7558
rect 5917 7546 5930 7560
rect 5998 7556 6151 7560
rect 5880 7544 5902 7546
rect 5980 7544 6172 7556
rect 6251 7544 6264 7574
rect 6279 7560 6309 7574
rect 6346 7544 6365 7574
rect 6380 7544 6386 7574
rect 6395 7544 6408 7574
rect 6423 7560 6453 7574
rect 6496 7560 6539 7574
rect 6546 7560 6766 7574
rect 6773 7560 6803 7574
rect 6463 7546 6478 7558
rect 6497 7546 6510 7560
rect 6578 7556 6731 7560
rect 6460 7544 6482 7546
rect 6560 7544 6752 7556
rect 6831 7544 6844 7574
rect 6859 7560 6889 7574
rect 6926 7544 6945 7574
rect 6960 7544 6966 7574
rect 6975 7544 6988 7574
rect 7003 7560 7033 7574
rect 7076 7560 7119 7574
rect 7126 7560 7346 7574
rect 7353 7560 7383 7574
rect 7043 7546 7058 7558
rect 7077 7546 7090 7560
rect 7158 7556 7311 7560
rect 7040 7544 7062 7546
rect 7140 7544 7332 7556
rect 7411 7544 7424 7574
rect 7439 7560 7469 7574
rect 7506 7544 7525 7574
rect 7540 7544 7546 7574
rect 7555 7544 7568 7574
rect 7583 7556 7613 7574
rect 7656 7560 7670 7574
rect 7706 7560 7926 7574
rect 7657 7558 7670 7560
rect 7623 7546 7638 7558
rect 7620 7544 7642 7546
rect 7647 7544 7677 7558
rect 7738 7556 7891 7560
rect 7720 7544 7912 7556
rect 7955 7544 7985 7558
rect 7991 7544 8004 7574
rect 8019 7556 8049 7574
rect 8092 7544 8105 7574
rect 8135 7544 8148 7574
rect 8163 7556 8193 7574
rect 8236 7560 8250 7574
rect 8286 7560 8506 7574
rect 8237 7558 8250 7560
rect 8203 7546 8218 7558
rect 8200 7544 8222 7546
rect 8227 7544 8257 7558
rect 8318 7556 8471 7560
rect 8300 7544 8492 7556
rect 8535 7544 8565 7558
rect 8571 7544 8584 7574
rect 8599 7556 8629 7574
rect 8672 7544 8685 7574
rect 8715 7544 8728 7574
rect 8743 7556 8773 7574
rect 8816 7560 8830 7574
rect 8866 7560 9086 7574
rect 8817 7558 8830 7560
rect 8783 7546 8798 7558
rect 8780 7544 8802 7546
rect 8807 7544 8837 7558
rect 8898 7556 9051 7560
rect 8880 7544 9072 7556
rect 9115 7544 9145 7558
rect 9151 7544 9164 7574
rect 9179 7556 9209 7574
rect 9252 7544 9265 7574
rect 0 7530 9265 7544
rect 15 7426 28 7530
rect 73 7508 74 7518
rect 89 7508 102 7518
rect 73 7504 102 7508
rect 107 7504 137 7530
rect 155 7516 171 7518
rect 243 7516 296 7530
rect 244 7514 308 7516
rect 351 7514 366 7530
rect 415 7527 445 7530
rect 415 7524 451 7527
rect 381 7516 397 7518
rect 155 7504 170 7508
rect 73 7502 170 7504
rect 198 7502 366 7514
rect 382 7504 397 7508
rect 415 7505 454 7524
rect 473 7518 480 7519
rect 479 7511 480 7518
rect 463 7508 464 7511
rect 479 7508 492 7511
rect 415 7504 445 7505
rect 454 7504 460 7505
rect 463 7504 492 7508
rect 382 7503 492 7504
rect 382 7502 498 7503
rect 57 7494 108 7502
rect 57 7482 82 7494
rect 89 7482 108 7494
rect 139 7494 189 7502
rect 139 7486 155 7494
rect 162 7492 189 7494
rect 198 7492 419 7502
rect 162 7482 419 7492
rect 448 7494 498 7502
rect 448 7485 464 7494
rect 57 7474 108 7482
rect 155 7474 419 7482
rect 445 7482 464 7485
rect 471 7482 498 7494
rect 445 7474 498 7482
rect 73 7466 74 7474
rect 89 7466 102 7474
rect 73 7458 89 7466
rect 70 7451 89 7454
rect 70 7442 92 7451
rect 43 7432 92 7442
rect 43 7426 73 7432
rect 92 7427 97 7432
rect 15 7410 89 7426
rect 107 7418 137 7474
rect 172 7464 380 7474
rect 415 7470 460 7474
rect 463 7473 464 7474
rect 479 7473 492 7474
rect 198 7434 387 7464
rect 213 7431 387 7434
rect 206 7428 387 7431
rect 15 7408 28 7410
rect 43 7408 77 7410
rect 15 7392 89 7408
rect 116 7404 129 7418
rect 144 7404 160 7420
rect 206 7415 217 7428
rect -1 7370 0 7386
rect 15 7370 28 7392
rect 43 7370 73 7392
rect 116 7388 178 7404
rect 206 7397 217 7413
rect 222 7408 232 7428
rect 242 7408 256 7428
rect 259 7415 268 7428
rect 284 7415 293 7428
rect 222 7397 256 7408
rect 259 7397 268 7413
rect 284 7397 293 7413
rect 300 7408 310 7428
rect 320 7408 334 7428
rect 335 7415 346 7428
rect 300 7397 334 7408
rect 335 7397 346 7413
rect 392 7404 408 7420
rect 415 7418 445 7470
rect 479 7466 480 7473
rect 464 7458 480 7466
rect 451 7426 464 7445
rect 479 7426 509 7442
rect 451 7410 525 7426
rect 451 7408 464 7410
rect 479 7408 513 7410
rect 116 7386 129 7388
rect 144 7386 178 7388
rect 116 7370 178 7386
rect 222 7381 238 7384
rect 300 7381 330 7392
rect 378 7388 424 7404
rect 451 7392 525 7408
rect 378 7386 412 7388
rect 377 7370 424 7386
rect 451 7370 464 7392
rect 479 7370 509 7392
rect 536 7370 537 7386
rect 552 7370 565 7530
rect 595 7426 608 7530
rect 653 7508 654 7518
rect 669 7508 682 7518
rect 653 7504 682 7508
rect 687 7504 717 7530
rect 735 7516 751 7518
rect 823 7516 876 7530
rect 824 7514 888 7516
rect 931 7514 946 7530
rect 995 7527 1025 7530
rect 995 7524 1031 7527
rect 961 7516 977 7518
rect 735 7504 750 7508
rect 653 7502 750 7504
rect 778 7502 946 7514
rect 962 7504 977 7508
rect 995 7505 1034 7524
rect 1053 7518 1060 7519
rect 1059 7511 1060 7518
rect 1043 7508 1044 7511
rect 1059 7508 1072 7511
rect 995 7504 1025 7505
rect 1034 7504 1040 7505
rect 1043 7504 1072 7508
rect 962 7503 1072 7504
rect 962 7502 1078 7503
rect 637 7494 688 7502
rect 637 7482 662 7494
rect 669 7482 688 7494
rect 719 7494 769 7502
rect 719 7486 735 7494
rect 742 7492 769 7494
rect 778 7492 999 7502
rect 742 7482 999 7492
rect 1028 7494 1078 7502
rect 1028 7485 1044 7494
rect 637 7474 688 7482
rect 735 7474 999 7482
rect 1025 7482 1044 7485
rect 1051 7482 1078 7494
rect 1025 7474 1078 7482
rect 653 7466 654 7474
rect 669 7466 682 7474
rect 653 7458 669 7466
rect 650 7451 669 7454
rect 650 7442 672 7451
rect 623 7432 672 7442
rect 623 7426 653 7432
rect 672 7427 677 7432
rect 595 7410 669 7426
rect 687 7418 717 7474
rect 752 7464 960 7474
rect 995 7470 1040 7474
rect 1043 7473 1044 7474
rect 1059 7473 1072 7474
rect 778 7434 967 7464
rect 793 7431 967 7434
rect 786 7428 967 7431
rect 595 7408 608 7410
rect 623 7408 657 7410
rect 595 7392 669 7408
rect 696 7404 709 7418
rect 724 7404 740 7420
rect 786 7415 797 7428
rect 579 7370 580 7386
rect 595 7370 608 7392
rect 623 7370 653 7392
rect 696 7388 758 7404
rect 786 7397 797 7413
rect 802 7408 812 7428
rect 822 7408 836 7428
rect 839 7415 848 7428
rect 864 7415 873 7428
rect 802 7397 836 7408
rect 839 7397 848 7413
rect 864 7397 873 7413
rect 880 7408 890 7428
rect 900 7408 914 7428
rect 915 7415 926 7428
rect 880 7397 914 7408
rect 915 7397 926 7413
rect 972 7404 988 7420
rect 995 7418 1025 7470
rect 1059 7466 1060 7473
rect 1044 7458 1060 7466
rect 1031 7426 1044 7445
rect 1059 7426 1089 7442
rect 1031 7410 1105 7426
rect 1031 7408 1044 7410
rect 1059 7408 1093 7410
rect 696 7386 709 7388
rect 724 7386 758 7388
rect 696 7370 758 7386
rect 802 7381 818 7384
rect 880 7381 910 7392
rect 958 7388 1004 7404
rect 1031 7392 1105 7408
rect 958 7386 992 7388
rect 957 7370 1004 7386
rect 1031 7370 1044 7392
rect 1059 7370 1089 7392
rect 1116 7370 1117 7386
rect 1132 7370 1145 7530
rect 1175 7426 1188 7530
rect 1233 7508 1234 7518
rect 1249 7508 1262 7518
rect 1233 7504 1262 7508
rect 1267 7504 1297 7530
rect 1315 7516 1331 7518
rect 1403 7516 1456 7530
rect 1404 7514 1468 7516
rect 1511 7514 1526 7530
rect 1575 7527 1605 7530
rect 1575 7524 1611 7527
rect 1541 7516 1557 7518
rect 1315 7504 1330 7508
rect 1233 7502 1330 7504
rect 1358 7502 1526 7514
rect 1542 7504 1557 7508
rect 1575 7505 1614 7524
rect 1633 7518 1640 7519
rect 1639 7511 1640 7518
rect 1623 7508 1624 7511
rect 1639 7508 1652 7511
rect 1575 7504 1605 7505
rect 1614 7504 1620 7505
rect 1623 7504 1652 7508
rect 1542 7503 1652 7504
rect 1542 7502 1658 7503
rect 1217 7494 1268 7502
rect 1217 7482 1242 7494
rect 1249 7482 1268 7494
rect 1299 7494 1349 7502
rect 1299 7486 1315 7494
rect 1322 7492 1349 7494
rect 1358 7492 1579 7502
rect 1322 7482 1579 7492
rect 1608 7494 1658 7502
rect 1608 7485 1624 7494
rect 1217 7474 1268 7482
rect 1315 7474 1579 7482
rect 1605 7482 1624 7485
rect 1631 7482 1658 7494
rect 1605 7474 1658 7482
rect 1233 7466 1234 7474
rect 1249 7466 1262 7474
rect 1233 7458 1249 7466
rect 1230 7451 1249 7454
rect 1230 7442 1252 7451
rect 1203 7432 1252 7442
rect 1203 7426 1233 7432
rect 1252 7427 1257 7432
rect 1175 7410 1249 7426
rect 1267 7418 1297 7474
rect 1332 7464 1540 7474
rect 1575 7470 1620 7474
rect 1623 7473 1624 7474
rect 1639 7473 1652 7474
rect 1358 7434 1547 7464
rect 1373 7431 1547 7434
rect 1366 7428 1547 7431
rect 1175 7408 1188 7410
rect 1203 7408 1237 7410
rect 1175 7392 1249 7408
rect 1276 7404 1289 7418
rect 1304 7404 1320 7420
rect 1366 7415 1377 7428
rect 1159 7370 1160 7386
rect 1175 7370 1188 7392
rect 1203 7370 1233 7392
rect 1276 7388 1338 7404
rect 1366 7397 1377 7413
rect 1382 7408 1392 7428
rect 1402 7408 1416 7428
rect 1419 7415 1428 7428
rect 1444 7415 1453 7428
rect 1382 7397 1416 7408
rect 1419 7397 1428 7413
rect 1444 7397 1453 7413
rect 1460 7408 1470 7428
rect 1480 7408 1494 7428
rect 1495 7415 1506 7428
rect 1460 7397 1494 7408
rect 1495 7397 1506 7413
rect 1552 7404 1568 7420
rect 1575 7418 1605 7470
rect 1639 7466 1640 7473
rect 1624 7458 1640 7466
rect 1611 7426 1624 7445
rect 1639 7426 1669 7442
rect 1611 7410 1685 7426
rect 1611 7408 1624 7410
rect 1639 7408 1673 7410
rect 1276 7386 1289 7388
rect 1304 7386 1338 7388
rect 1276 7370 1338 7386
rect 1382 7381 1398 7384
rect 1460 7381 1490 7392
rect 1538 7388 1584 7404
rect 1611 7392 1685 7408
rect 1538 7386 1572 7388
rect 1537 7370 1584 7386
rect 1611 7370 1624 7392
rect 1639 7370 1669 7392
rect 1696 7370 1697 7386
rect 1712 7370 1725 7530
rect 1755 7426 1768 7530
rect 1820 7526 1842 7530
rect 1813 7504 1842 7518
rect 1895 7504 1911 7518
rect 1949 7514 1955 7516
rect 1962 7514 2070 7530
rect 2077 7514 2083 7516
rect 2091 7514 2106 7530
rect 2172 7524 2191 7527
rect 1813 7502 1911 7504
rect 1938 7502 2106 7514
rect 2121 7504 2137 7518
rect 2172 7505 2194 7524
rect 2204 7518 2220 7519
rect 2203 7516 2220 7518
rect 2204 7511 2220 7516
rect 2194 7504 2200 7505
rect 2203 7504 2232 7511
rect 2121 7503 2232 7504
rect 2121 7502 2238 7503
rect 1797 7494 1848 7502
rect 1895 7494 1929 7502
rect 1797 7482 1822 7494
rect 1829 7482 1848 7494
rect 1902 7492 1929 7494
rect 1938 7492 2159 7502
rect 2194 7499 2200 7502
rect 1902 7488 2159 7492
rect 1797 7474 1848 7482
rect 1895 7474 2159 7488
rect 2203 7494 2238 7502
rect 1813 7466 1842 7474
rect 1813 7460 1830 7466
rect 1813 7458 1847 7460
rect 1895 7458 1911 7474
rect 1912 7464 2120 7474
rect 2121 7464 2137 7474
rect 2185 7470 2200 7485
rect 2203 7482 2204 7494
rect 2211 7482 2238 7494
rect 2203 7474 2238 7482
rect 2203 7473 2232 7474
rect 1923 7460 2137 7464
rect 1938 7458 2137 7460
rect 2172 7460 2185 7470
rect 2203 7460 2220 7473
rect 2172 7458 2220 7460
rect 1814 7454 1847 7458
rect 1810 7452 1847 7454
rect 1810 7451 1877 7452
rect 1810 7446 1841 7451
rect 1847 7446 1877 7451
rect 1810 7442 1877 7446
rect 1783 7439 1877 7442
rect 1783 7432 1832 7439
rect 1783 7426 1813 7432
rect 1832 7427 1837 7432
rect 1755 7410 1829 7426
rect 1841 7418 1877 7439
rect 1938 7434 2127 7458
rect 2172 7457 2219 7458
rect 2185 7452 2219 7457
rect 1953 7431 2127 7434
rect 1946 7428 2127 7431
rect 2155 7451 2219 7452
rect 1755 7408 1768 7410
rect 1783 7408 1817 7410
rect 1755 7392 1829 7408
rect 1739 7370 1740 7386
rect 1755 7370 1768 7392
rect 1783 7376 1813 7392
rect 1841 7370 1847 7418
rect 1850 7412 1869 7418
rect 1884 7412 1914 7420
rect 1850 7404 1914 7412
rect 1850 7388 1930 7404
rect 1946 7397 2008 7428
rect 2024 7397 2086 7428
rect 2155 7426 2204 7451
rect 2219 7426 2249 7442
rect 2118 7412 2148 7420
rect 2155 7418 2265 7426
rect 2118 7404 2163 7412
rect 1850 7386 1869 7388
rect 1884 7386 1930 7388
rect 1850 7370 1930 7386
rect 1957 7384 1992 7397
rect 2033 7394 2070 7397
rect 2033 7392 2075 7394
rect 1962 7381 1992 7384
rect 1971 7377 1978 7381
rect 1978 7376 1979 7377
rect 1937 7370 1947 7376
rect -7 7362 34 7370
rect -7 7336 8 7362
rect 15 7336 34 7362
rect 98 7358 160 7370
rect 172 7358 247 7370
rect 305 7358 380 7370
rect 392 7358 423 7370
rect 429 7358 464 7370
rect 98 7356 260 7358
rect -7 7328 34 7336
rect 116 7332 129 7356
rect 144 7354 159 7356
rect -1 7318 0 7328
rect 15 7318 28 7328
rect 43 7318 73 7332
rect 116 7318 159 7332
rect 183 7329 190 7336
rect 193 7332 260 7356
rect 292 7356 464 7358
rect 262 7334 290 7338
rect 292 7334 372 7356
rect 393 7354 408 7356
rect 262 7332 372 7334
rect 193 7328 372 7332
rect 166 7318 196 7328
rect 198 7318 351 7328
rect 359 7318 389 7328
rect 393 7318 423 7332
rect 451 7318 464 7356
rect 536 7362 571 7370
rect 536 7336 537 7362
rect 544 7336 571 7362
rect 479 7318 509 7332
rect 536 7328 571 7336
rect 573 7362 614 7370
rect 573 7336 588 7362
rect 595 7336 614 7362
rect 678 7358 740 7370
rect 752 7358 827 7370
rect 885 7358 960 7370
rect 972 7358 1003 7370
rect 1009 7358 1044 7370
rect 678 7356 840 7358
rect 573 7328 614 7336
rect 696 7332 709 7356
rect 724 7354 739 7356
rect 536 7318 537 7328
rect 552 7318 565 7328
rect 579 7318 580 7328
rect 595 7318 608 7328
rect 623 7318 653 7332
rect 696 7318 739 7332
rect 763 7329 770 7336
rect 773 7332 840 7356
rect 872 7356 1044 7358
rect 842 7334 870 7338
rect 872 7334 952 7356
rect 973 7354 988 7356
rect 842 7332 952 7334
rect 773 7328 952 7332
rect 746 7318 776 7328
rect 778 7318 931 7328
rect 939 7318 969 7328
rect 973 7318 1003 7332
rect 1031 7318 1044 7356
rect 1116 7362 1151 7370
rect 1116 7336 1117 7362
rect 1124 7336 1151 7362
rect 1059 7318 1089 7332
rect 1116 7328 1151 7336
rect 1153 7362 1194 7370
rect 1153 7336 1168 7362
rect 1175 7336 1194 7362
rect 1258 7358 1320 7370
rect 1332 7358 1407 7370
rect 1465 7358 1540 7370
rect 1552 7358 1583 7370
rect 1589 7358 1624 7370
rect 1258 7356 1420 7358
rect 1153 7328 1194 7336
rect 1276 7332 1289 7356
rect 1304 7354 1319 7356
rect 1116 7318 1117 7328
rect 1132 7318 1145 7328
rect 1159 7318 1160 7328
rect 1175 7318 1188 7328
rect 1203 7318 1233 7332
rect 1276 7318 1319 7332
rect 1343 7329 1350 7336
rect 1353 7332 1420 7356
rect 1452 7356 1624 7358
rect 1422 7334 1450 7338
rect 1452 7334 1532 7356
rect 1553 7354 1568 7356
rect 1422 7332 1532 7334
rect 1353 7328 1532 7332
rect 1326 7318 1356 7328
rect 1358 7318 1511 7328
rect 1519 7318 1549 7328
rect 1553 7318 1583 7332
rect 1611 7318 1624 7356
rect 1696 7362 1731 7370
rect 1696 7336 1697 7362
rect 1704 7336 1731 7362
rect 1639 7318 1669 7332
rect 1696 7328 1731 7336
rect 1733 7362 1774 7370
rect 1733 7336 1748 7362
rect 1755 7336 1774 7362
rect 1838 7358 1869 7370
rect 1884 7358 1987 7370
rect 1999 7360 2025 7386
rect 2040 7381 2070 7392
rect 2102 7388 2164 7404
rect 2102 7386 2148 7388
rect 2102 7370 2164 7386
rect 2176 7370 2182 7418
rect 2185 7410 2265 7418
rect 2185 7408 2204 7410
rect 2219 7408 2253 7410
rect 2185 7392 2265 7408
rect 2185 7370 2204 7392
rect 2219 7376 2249 7392
rect 2277 7386 2283 7460
rect 2286 7386 2305 7530
rect 2320 7386 2326 7530
rect 2335 7460 2348 7530
rect 2400 7526 2422 7530
rect 2393 7504 2422 7518
rect 2475 7504 2491 7518
rect 2529 7514 2535 7516
rect 2542 7514 2650 7530
rect 2657 7514 2663 7516
rect 2671 7514 2686 7530
rect 2752 7524 2771 7527
rect 2393 7502 2491 7504
rect 2518 7502 2686 7514
rect 2701 7504 2717 7518
rect 2752 7505 2774 7524
rect 2784 7518 2800 7519
rect 2783 7516 2800 7518
rect 2784 7511 2800 7516
rect 2774 7504 2780 7505
rect 2783 7504 2812 7511
rect 2701 7503 2812 7504
rect 2701 7502 2818 7503
rect 2377 7494 2428 7502
rect 2475 7494 2509 7502
rect 2377 7482 2402 7494
rect 2409 7482 2428 7494
rect 2482 7492 2509 7494
rect 2518 7492 2739 7502
rect 2774 7499 2780 7502
rect 2482 7488 2739 7492
rect 2377 7474 2428 7482
rect 2475 7474 2739 7488
rect 2783 7494 2818 7502
rect 2329 7426 2348 7460
rect 2393 7466 2422 7474
rect 2393 7460 2410 7466
rect 2393 7458 2427 7460
rect 2475 7458 2491 7474
rect 2492 7464 2700 7474
rect 2701 7464 2717 7474
rect 2765 7470 2780 7485
rect 2783 7482 2784 7494
rect 2791 7482 2818 7494
rect 2783 7474 2818 7482
rect 2783 7473 2812 7474
rect 2503 7460 2717 7464
rect 2518 7458 2717 7460
rect 2752 7460 2765 7470
rect 2783 7460 2800 7473
rect 2752 7458 2800 7460
rect 2394 7454 2427 7458
rect 2390 7452 2427 7454
rect 2390 7451 2457 7452
rect 2390 7446 2421 7451
rect 2427 7446 2457 7451
rect 2390 7442 2457 7446
rect 2363 7439 2457 7442
rect 2363 7432 2412 7439
rect 2363 7426 2393 7432
rect 2412 7427 2417 7432
rect 2329 7410 2409 7426
rect 2421 7418 2457 7439
rect 2518 7434 2707 7458
rect 2752 7457 2799 7458
rect 2765 7452 2799 7457
rect 2533 7431 2707 7434
rect 2526 7428 2707 7431
rect 2735 7451 2799 7452
rect 2329 7408 2348 7410
rect 2363 7408 2397 7410
rect 2329 7392 2409 7408
rect 2329 7386 2348 7392
rect 2045 7360 2148 7370
rect 1999 7358 2148 7360
rect 2169 7358 2204 7370
rect 1838 7356 2000 7358
rect 1850 7336 1869 7356
rect 1884 7354 1914 7356
rect 1733 7328 1774 7336
rect 1856 7332 1869 7336
rect 1921 7340 2000 7356
rect 2032 7356 2204 7358
rect 2032 7340 2111 7356
rect 2118 7354 2148 7356
rect 1696 7318 1697 7328
rect 1712 7318 1725 7328
rect 1739 7318 1740 7328
rect 1755 7318 1768 7328
rect 1783 7318 1813 7332
rect 1856 7318 1899 7332
rect 1921 7328 2111 7340
rect 2176 7336 2182 7356
rect 1906 7318 1936 7328
rect 1937 7318 2095 7328
rect 2099 7318 2129 7328
rect 2133 7318 2163 7332
rect 2191 7318 2204 7356
rect 2276 7370 2305 7386
rect 2319 7370 2348 7386
rect 2363 7376 2393 7392
rect 2421 7370 2427 7418
rect 2430 7412 2449 7418
rect 2464 7412 2494 7420
rect 2430 7404 2494 7412
rect 2430 7388 2510 7404
rect 2526 7397 2588 7428
rect 2604 7397 2666 7428
rect 2735 7426 2784 7451
rect 2799 7426 2829 7442
rect 2698 7412 2728 7420
rect 2735 7418 2845 7426
rect 2698 7404 2743 7412
rect 2430 7386 2449 7388
rect 2464 7386 2510 7388
rect 2430 7370 2510 7386
rect 2537 7384 2572 7397
rect 2613 7394 2650 7397
rect 2613 7392 2655 7394
rect 2542 7381 2572 7384
rect 2551 7377 2558 7381
rect 2558 7376 2559 7377
rect 2517 7370 2527 7376
rect 2276 7362 2311 7370
rect 2276 7336 2277 7362
rect 2284 7336 2311 7362
rect 2219 7318 2249 7332
rect 2276 7328 2311 7336
rect 2313 7362 2354 7370
rect 2313 7336 2328 7362
rect 2335 7336 2354 7362
rect 2418 7358 2449 7370
rect 2464 7358 2567 7370
rect 2579 7360 2605 7386
rect 2620 7381 2650 7392
rect 2682 7388 2744 7404
rect 2682 7386 2728 7388
rect 2682 7370 2744 7386
rect 2756 7370 2762 7418
rect 2765 7410 2845 7418
rect 2765 7408 2784 7410
rect 2799 7408 2833 7410
rect 2765 7392 2845 7408
rect 2765 7370 2784 7392
rect 2799 7376 2829 7392
rect 2857 7386 2863 7460
rect 2866 7386 2885 7530
rect 2900 7386 2906 7530
rect 2915 7460 2928 7530
rect 2980 7526 3002 7530
rect 2973 7504 3002 7518
rect 3055 7504 3071 7518
rect 3109 7514 3115 7516
rect 3122 7514 3230 7530
rect 3237 7514 3243 7516
rect 3251 7514 3266 7530
rect 3332 7524 3351 7527
rect 2973 7502 3071 7504
rect 3098 7502 3266 7514
rect 3281 7504 3297 7518
rect 3332 7505 3354 7524
rect 3364 7518 3380 7519
rect 3363 7516 3380 7518
rect 3364 7511 3380 7516
rect 3354 7504 3360 7505
rect 3363 7504 3392 7511
rect 3281 7503 3392 7504
rect 3281 7502 3398 7503
rect 2957 7494 3008 7502
rect 3055 7494 3089 7502
rect 2957 7482 2982 7494
rect 2989 7482 3008 7494
rect 3062 7492 3089 7494
rect 3098 7492 3319 7502
rect 3354 7499 3360 7502
rect 3062 7488 3319 7492
rect 2957 7474 3008 7482
rect 3055 7474 3319 7488
rect 3363 7494 3398 7502
rect 2909 7426 2928 7460
rect 2973 7466 3002 7474
rect 2973 7460 2990 7466
rect 2973 7458 3007 7460
rect 3055 7458 3071 7474
rect 3072 7464 3280 7474
rect 3281 7464 3297 7474
rect 3345 7470 3360 7485
rect 3363 7482 3364 7494
rect 3371 7482 3398 7494
rect 3363 7474 3398 7482
rect 3363 7473 3392 7474
rect 3083 7460 3297 7464
rect 3098 7458 3297 7460
rect 3332 7460 3345 7470
rect 3363 7460 3380 7473
rect 3332 7458 3380 7460
rect 2974 7454 3007 7458
rect 2970 7452 3007 7454
rect 2970 7451 3037 7452
rect 2970 7446 3001 7451
rect 3007 7446 3037 7451
rect 2970 7442 3037 7446
rect 2943 7439 3037 7442
rect 2943 7432 2992 7439
rect 2943 7426 2973 7432
rect 2992 7427 2997 7432
rect 2909 7410 2989 7426
rect 3001 7418 3037 7439
rect 3098 7434 3287 7458
rect 3332 7457 3379 7458
rect 3345 7452 3379 7457
rect 3113 7431 3287 7434
rect 3106 7428 3287 7431
rect 3315 7451 3379 7452
rect 2909 7408 2928 7410
rect 2943 7408 2977 7410
rect 2909 7392 2989 7408
rect 2909 7386 2928 7392
rect 2625 7360 2728 7370
rect 2579 7358 2728 7360
rect 2749 7358 2784 7370
rect 2418 7356 2580 7358
rect 2430 7336 2449 7356
rect 2464 7354 2494 7356
rect 2313 7328 2354 7336
rect 2436 7332 2449 7336
rect 2501 7340 2580 7356
rect 2612 7356 2784 7358
rect 2612 7340 2691 7356
rect 2698 7354 2728 7356
rect 2276 7318 2305 7328
rect 2319 7318 2348 7328
rect 2363 7318 2393 7332
rect 2436 7318 2479 7332
rect 2501 7328 2691 7340
rect 2756 7336 2762 7356
rect 2486 7318 2516 7328
rect 2517 7318 2675 7328
rect 2679 7318 2709 7328
rect 2713 7318 2743 7332
rect 2771 7318 2784 7356
rect 2856 7370 2885 7386
rect 2899 7370 2928 7386
rect 2943 7376 2973 7392
rect 3001 7370 3007 7418
rect 3010 7412 3029 7418
rect 3044 7412 3074 7420
rect 3010 7404 3074 7412
rect 3010 7388 3090 7404
rect 3106 7397 3168 7428
rect 3184 7397 3246 7428
rect 3315 7426 3364 7451
rect 3379 7426 3409 7442
rect 3278 7412 3308 7420
rect 3315 7418 3425 7426
rect 3278 7404 3323 7412
rect 3010 7386 3029 7388
rect 3044 7386 3090 7388
rect 3010 7370 3090 7386
rect 3117 7384 3152 7397
rect 3193 7394 3230 7397
rect 3193 7392 3235 7394
rect 3122 7381 3152 7384
rect 3131 7377 3138 7381
rect 3138 7376 3139 7377
rect 3097 7370 3107 7376
rect 2856 7362 2891 7370
rect 2856 7336 2857 7362
rect 2864 7336 2891 7362
rect 2799 7318 2829 7332
rect 2856 7328 2891 7336
rect 2893 7362 2934 7370
rect 2893 7336 2908 7362
rect 2915 7336 2934 7362
rect 2998 7358 3029 7370
rect 3044 7358 3147 7370
rect 3159 7360 3185 7386
rect 3200 7381 3230 7392
rect 3262 7388 3324 7404
rect 3262 7386 3308 7388
rect 3262 7370 3324 7386
rect 3336 7370 3342 7418
rect 3345 7410 3425 7418
rect 3345 7408 3364 7410
rect 3379 7408 3413 7410
rect 3345 7392 3425 7408
rect 3345 7370 3364 7392
rect 3379 7376 3409 7392
rect 3437 7386 3443 7460
rect 3446 7386 3465 7530
rect 3480 7386 3486 7530
rect 3495 7460 3508 7530
rect 3560 7526 3582 7530
rect 3553 7504 3582 7518
rect 3635 7504 3651 7518
rect 3689 7514 3695 7516
rect 3702 7514 3810 7530
rect 3817 7514 3823 7516
rect 3831 7514 3846 7530
rect 3912 7524 3931 7527
rect 3553 7502 3651 7504
rect 3678 7502 3846 7514
rect 3861 7504 3877 7518
rect 3912 7505 3934 7524
rect 3944 7518 3960 7519
rect 3943 7516 3960 7518
rect 3944 7511 3960 7516
rect 3934 7504 3940 7505
rect 3943 7504 3972 7511
rect 3861 7503 3972 7504
rect 3861 7502 3978 7503
rect 3537 7494 3588 7502
rect 3635 7494 3669 7502
rect 3537 7482 3562 7494
rect 3569 7482 3588 7494
rect 3642 7492 3669 7494
rect 3678 7492 3899 7502
rect 3934 7499 3940 7502
rect 3642 7488 3899 7492
rect 3537 7474 3588 7482
rect 3635 7474 3899 7488
rect 3943 7494 3978 7502
rect 3489 7426 3508 7460
rect 3553 7466 3582 7474
rect 3553 7460 3570 7466
rect 3553 7458 3587 7460
rect 3635 7458 3651 7474
rect 3652 7464 3860 7474
rect 3861 7464 3877 7474
rect 3925 7470 3940 7485
rect 3943 7482 3944 7494
rect 3951 7482 3978 7494
rect 3943 7474 3978 7482
rect 3943 7473 3972 7474
rect 3663 7460 3877 7464
rect 3678 7458 3877 7460
rect 3912 7460 3925 7470
rect 3943 7460 3960 7473
rect 3912 7458 3960 7460
rect 3554 7454 3587 7458
rect 3550 7452 3587 7454
rect 3550 7451 3617 7452
rect 3550 7446 3581 7451
rect 3587 7446 3617 7451
rect 3550 7442 3617 7446
rect 3523 7439 3617 7442
rect 3523 7432 3572 7439
rect 3523 7426 3553 7432
rect 3572 7427 3577 7432
rect 3489 7410 3569 7426
rect 3581 7418 3617 7439
rect 3678 7434 3867 7458
rect 3912 7457 3959 7458
rect 3925 7452 3959 7457
rect 3693 7431 3867 7434
rect 3686 7428 3867 7431
rect 3895 7451 3959 7452
rect 3489 7408 3508 7410
rect 3523 7408 3557 7410
rect 3489 7392 3569 7408
rect 3489 7386 3508 7392
rect 3205 7360 3308 7370
rect 3159 7358 3308 7360
rect 3329 7358 3364 7370
rect 2998 7356 3160 7358
rect 3010 7336 3029 7356
rect 3044 7354 3074 7356
rect 2893 7328 2934 7336
rect 3016 7332 3029 7336
rect 3081 7340 3160 7356
rect 3192 7356 3364 7358
rect 3192 7340 3271 7356
rect 3278 7354 3308 7356
rect 2856 7318 2885 7328
rect 2899 7318 2928 7328
rect 2943 7318 2973 7332
rect 3016 7318 3059 7332
rect 3081 7328 3271 7340
rect 3336 7336 3342 7356
rect 3066 7318 3096 7328
rect 3097 7318 3255 7328
rect 3259 7318 3289 7328
rect 3293 7318 3323 7332
rect 3351 7318 3364 7356
rect 3436 7370 3465 7386
rect 3479 7370 3508 7386
rect 3523 7376 3553 7392
rect 3581 7370 3587 7418
rect 3590 7412 3609 7418
rect 3624 7412 3654 7420
rect 3590 7404 3654 7412
rect 3590 7388 3670 7404
rect 3686 7397 3748 7428
rect 3764 7397 3826 7428
rect 3895 7426 3944 7451
rect 3959 7426 3989 7442
rect 3858 7412 3888 7420
rect 3895 7418 4005 7426
rect 3858 7404 3903 7412
rect 3590 7386 3609 7388
rect 3624 7386 3670 7388
rect 3590 7370 3670 7386
rect 3697 7384 3732 7397
rect 3773 7394 3810 7397
rect 3773 7392 3815 7394
rect 3702 7381 3732 7384
rect 3711 7377 3718 7381
rect 3718 7376 3719 7377
rect 3677 7370 3687 7376
rect 3436 7362 3471 7370
rect 3436 7336 3437 7362
rect 3444 7336 3471 7362
rect 3379 7318 3409 7332
rect 3436 7328 3471 7336
rect 3473 7362 3514 7370
rect 3473 7336 3488 7362
rect 3495 7336 3514 7362
rect 3578 7358 3609 7370
rect 3624 7358 3727 7370
rect 3739 7360 3765 7386
rect 3780 7381 3810 7392
rect 3842 7388 3904 7404
rect 3842 7386 3888 7388
rect 3842 7370 3904 7386
rect 3916 7370 3922 7418
rect 3925 7410 4005 7418
rect 3925 7408 3944 7410
rect 3959 7408 3993 7410
rect 3925 7392 4005 7408
rect 3925 7370 3944 7392
rect 3959 7376 3989 7392
rect 4017 7386 4023 7460
rect 4026 7386 4045 7530
rect 4060 7386 4066 7530
rect 4075 7460 4088 7530
rect 4140 7526 4162 7530
rect 4133 7504 4162 7518
rect 4215 7504 4231 7518
rect 4269 7514 4275 7516
rect 4282 7514 4390 7530
rect 4397 7514 4403 7516
rect 4411 7514 4426 7530
rect 4492 7524 4511 7527
rect 4133 7502 4231 7504
rect 4258 7502 4426 7514
rect 4441 7504 4457 7518
rect 4492 7505 4514 7524
rect 4524 7518 4540 7519
rect 4523 7516 4540 7518
rect 4524 7511 4540 7516
rect 4514 7504 4520 7505
rect 4523 7504 4552 7511
rect 4441 7503 4552 7504
rect 4441 7502 4558 7503
rect 4117 7494 4168 7502
rect 4215 7494 4249 7502
rect 4117 7482 4142 7494
rect 4149 7482 4168 7494
rect 4222 7492 4249 7494
rect 4258 7492 4479 7502
rect 4514 7499 4520 7502
rect 4222 7488 4479 7492
rect 4117 7474 4168 7482
rect 4215 7474 4479 7488
rect 4523 7494 4558 7502
rect 4069 7426 4088 7460
rect 4133 7466 4162 7474
rect 4133 7460 4150 7466
rect 4133 7458 4167 7460
rect 4215 7458 4231 7474
rect 4232 7464 4440 7474
rect 4441 7464 4457 7474
rect 4505 7470 4520 7485
rect 4523 7482 4524 7494
rect 4531 7482 4558 7494
rect 4523 7474 4558 7482
rect 4523 7473 4552 7474
rect 4243 7460 4457 7464
rect 4258 7458 4457 7460
rect 4492 7460 4505 7470
rect 4523 7460 4540 7473
rect 4492 7458 4540 7460
rect 4134 7454 4167 7458
rect 4130 7452 4167 7454
rect 4130 7451 4197 7452
rect 4130 7446 4161 7451
rect 4167 7446 4197 7451
rect 4130 7442 4197 7446
rect 4103 7439 4197 7442
rect 4103 7432 4152 7439
rect 4103 7426 4133 7432
rect 4152 7427 4157 7432
rect 4069 7410 4149 7426
rect 4161 7418 4197 7439
rect 4258 7434 4447 7458
rect 4492 7457 4539 7458
rect 4505 7452 4539 7457
rect 4273 7431 4447 7434
rect 4266 7428 4447 7431
rect 4475 7451 4539 7452
rect 4069 7408 4088 7410
rect 4103 7408 4137 7410
rect 4069 7392 4149 7408
rect 4069 7386 4088 7392
rect 3785 7360 3888 7370
rect 3739 7358 3888 7360
rect 3909 7358 3944 7370
rect 3578 7356 3740 7358
rect 3590 7336 3609 7356
rect 3624 7354 3654 7356
rect 3473 7328 3514 7336
rect 3596 7332 3609 7336
rect 3661 7340 3740 7356
rect 3772 7356 3944 7358
rect 3772 7340 3851 7356
rect 3858 7354 3888 7356
rect 3436 7318 3465 7328
rect 3479 7318 3508 7328
rect 3523 7318 3553 7332
rect 3596 7318 3639 7332
rect 3661 7328 3851 7340
rect 3916 7336 3922 7356
rect 3646 7318 3676 7328
rect 3677 7318 3835 7328
rect 3839 7318 3869 7328
rect 3873 7318 3903 7332
rect 3931 7318 3944 7356
rect 4016 7370 4045 7386
rect 4059 7370 4088 7386
rect 4103 7376 4133 7392
rect 4161 7370 4167 7418
rect 4170 7412 4189 7418
rect 4204 7412 4234 7420
rect 4170 7404 4234 7412
rect 4170 7388 4250 7404
rect 4266 7397 4328 7428
rect 4344 7397 4406 7428
rect 4475 7426 4524 7451
rect 4539 7426 4569 7442
rect 4438 7412 4468 7420
rect 4475 7418 4585 7426
rect 4438 7404 4483 7412
rect 4170 7386 4189 7388
rect 4204 7386 4250 7388
rect 4170 7370 4250 7386
rect 4277 7384 4312 7397
rect 4353 7394 4390 7397
rect 4353 7392 4395 7394
rect 4282 7381 4312 7384
rect 4291 7377 4298 7381
rect 4298 7376 4299 7377
rect 4257 7370 4267 7376
rect 4016 7362 4051 7370
rect 4016 7336 4017 7362
rect 4024 7336 4051 7362
rect 3959 7318 3989 7332
rect 4016 7328 4051 7336
rect 4053 7362 4094 7370
rect 4053 7336 4068 7362
rect 4075 7336 4094 7362
rect 4158 7358 4189 7370
rect 4204 7358 4307 7370
rect 4319 7360 4345 7386
rect 4360 7381 4390 7392
rect 4422 7388 4484 7404
rect 4422 7386 4468 7388
rect 4422 7370 4484 7386
rect 4496 7370 4502 7418
rect 4505 7410 4585 7418
rect 4505 7408 4524 7410
rect 4539 7408 4573 7410
rect 4505 7392 4585 7408
rect 4505 7370 4524 7392
rect 4539 7376 4569 7392
rect 4597 7386 4603 7460
rect 4606 7386 4625 7530
rect 4640 7386 4646 7530
rect 4655 7460 4668 7530
rect 4720 7526 4742 7530
rect 4713 7504 4742 7518
rect 4795 7504 4811 7518
rect 4849 7514 4855 7516
rect 4862 7514 4970 7530
rect 4977 7514 4983 7516
rect 4991 7514 5006 7530
rect 5072 7524 5091 7527
rect 4713 7502 4811 7504
rect 4838 7502 5006 7514
rect 5021 7504 5037 7518
rect 5072 7505 5094 7524
rect 5104 7518 5120 7519
rect 5103 7516 5120 7518
rect 5104 7511 5120 7516
rect 5094 7504 5100 7505
rect 5103 7504 5132 7511
rect 5021 7503 5132 7504
rect 5021 7502 5138 7503
rect 4697 7494 4748 7502
rect 4795 7494 4829 7502
rect 4697 7482 4722 7494
rect 4729 7482 4748 7494
rect 4802 7492 4829 7494
rect 4838 7492 5059 7502
rect 5094 7499 5100 7502
rect 4802 7488 5059 7492
rect 4697 7474 4748 7482
rect 4795 7474 5059 7488
rect 5103 7494 5138 7502
rect 4649 7426 4668 7460
rect 4713 7466 4742 7474
rect 4713 7460 4730 7466
rect 4713 7458 4747 7460
rect 4795 7458 4811 7474
rect 4812 7464 5020 7474
rect 5021 7464 5037 7474
rect 5085 7470 5100 7485
rect 5103 7482 5104 7494
rect 5111 7482 5138 7494
rect 5103 7474 5138 7482
rect 5103 7473 5132 7474
rect 4823 7460 5037 7464
rect 4838 7458 5037 7460
rect 5072 7460 5085 7470
rect 5103 7460 5120 7473
rect 5072 7458 5120 7460
rect 4714 7454 4747 7458
rect 4710 7452 4747 7454
rect 4710 7451 4777 7452
rect 4710 7446 4741 7451
rect 4747 7446 4777 7451
rect 4710 7442 4777 7446
rect 4683 7439 4777 7442
rect 4683 7432 4732 7439
rect 4683 7426 4713 7432
rect 4732 7427 4737 7432
rect 4649 7410 4729 7426
rect 4741 7418 4777 7439
rect 4838 7434 5027 7458
rect 5072 7457 5119 7458
rect 5085 7452 5119 7457
rect 4853 7431 5027 7434
rect 4846 7428 5027 7431
rect 5055 7451 5119 7452
rect 4649 7408 4668 7410
rect 4683 7408 4717 7410
rect 4649 7392 4729 7408
rect 4649 7386 4668 7392
rect 4365 7360 4468 7370
rect 4319 7358 4468 7360
rect 4489 7358 4524 7370
rect 4158 7356 4320 7358
rect 4170 7336 4189 7356
rect 4204 7354 4234 7356
rect 4053 7328 4094 7336
rect 4176 7332 4189 7336
rect 4241 7340 4320 7356
rect 4352 7356 4524 7358
rect 4352 7340 4431 7356
rect 4438 7354 4468 7356
rect 4016 7318 4045 7328
rect 4059 7318 4088 7328
rect 4103 7318 4133 7332
rect 4176 7318 4219 7332
rect 4241 7328 4431 7340
rect 4496 7336 4502 7356
rect 4226 7318 4256 7328
rect 4257 7318 4415 7328
rect 4419 7318 4449 7328
rect 4453 7318 4483 7332
rect 4511 7318 4524 7356
rect 4596 7370 4625 7386
rect 4639 7370 4668 7386
rect 4683 7376 4713 7392
rect 4741 7370 4747 7418
rect 4750 7412 4769 7418
rect 4784 7412 4814 7420
rect 4750 7404 4814 7412
rect 4750 7388 4830 7404
rect 4846 7397 4908 7428
rect 4924 7397 4986 7428
rect 5055 7426 5104 7451
rect 5119 7426 5149 7442
rect 5018 7412 5048 7420
rect 5055 7418 5165 7426
rect 5018 7404 5063 7412
rect 4750 7386 4769 7388
rect 4784 7386 4830 7388
rect 4750 7370 4830 7386
rect 4857 7384 4892 7397
rect 4933 7394 4970 7397
rect 4933 7392 4975 7394
rect 4862 7381 4892 7384
rect 4871 7377 4878 7381
rect 4878 7376 4879 7377
rect 4837 7370 4847 7376
rect 4596 7362 4631 7370
rect 4596 7336 4597 7362
rect 4604 7336 4631 7362
rect 4539 7318 4569 7332
rect 4596 7328 4631 7336
rect 4633 7362 4674 7370
rect 4633 7336 4648 7362
rect 4655 7336 4674 7362
rect 4738 7358 4769 7370
rect 4784 7358 4887 7370
rect 4899 7360 4925 7386
rect 4940 7381 4970 7392
rect 5002 7388 5064 7404
rect 5002 7386 5048 7388
rect 5002 7370 5064 7386
rect 5076 7370 5082 7418
rect 5085 7410 5165 7418
rect 5085 7408 5104 7410
rect 5119 7408 5153 7410
rect 5085 7392 5165 7408
rect 5085 7370 5104 7392
rect 5119 7376 5149 7392
rect 5177 7386 5183 7460
rect 5186 7386 5205 7530
rect 5220 7386 5226 7530
rect 5235 7460 5248 7530
rect 5300 7526 5322 7530
rect 5293 7504 5322 7518
rect 5375 7504 5391 7518
rect 5429 7514 5435 7516
rect 5442 7514 5550 7530
rect 5557 7514 5563 7516
rect 5571 7514 5586 7530
rect 5652 7524 5671 7527
rect 5293 7502 5391 7504
rect 5418 7502 5586 7514
rect 5601 7504 5617 7518
rect 5652 7505 5674 7524
rect 5684 7518 5700 7519
rect 5683 7516 5700 7518
rect 5684 7511 5700 7516
rect 5674 7504 5680 7505
rect 5683 7504 5712 7511
rect 5601 7503 5712 7504
rect 5601 7502 5718 7503
rect 5277 7494 5328 7502
rect 5375 7494 5409 7502
rect 5277 7482 5302 7494
rect 5309 7482 5328 7494
rect 5382 7492 5409 7494
rect 5418 7492 5639 7502
rect 5674 7499 5680 7502
rect 5382 7488 5639 7492
rect 5277 7474 5328 7482
rect 5375 7474 5639 7488
rect 5683 7494 5718 7502
rect 5229 7426 5248 7460
rect 5293 7466 5322 7474
rect 5293 7460 5310 7466
rect 5293 7458 5327 7460
rect 5375 7458 5391 7474
rect 5392 7464 5600 7474
rect 5601 7464 5617 7474
rect 5665 7470 5680 7485
rect 5683 7482 5684 7494
rect 5691 7482 5718 7494
rect 5683 7474 5718 7482
rect 5683 7473 5712 7474
rect 5403 7460 5617 7464
rect 5418 7458 5617 7460
rect 5652 7460 5665 7470
rect 5683 7460 5700 7473
rect 5652 7458 5700 7460
rect 5294 7454 5327 7458
rect 5290 7452 5327 7454
rect 5290 7451 5357 7452
rect 5290 7446 5321 7451
rect 5327 7446 5357 7451
rect 5290 7442 5357 7446
rect 5263 7439 5357 7442
rect 5263 7432 5312 7439
rect 5263 7426 5293 7432
rect 5312 7427 5317 7432
rect 5229 7410 5309 7426
rect 5321 7418 5357 7439
rect 5418 7434 5607 7458
rect 5652 7457 5699 7458
rect 5665 7452 5699 7457
rect 5433 7431 5607 7434
rect 5426 7428 5607 7431
rect 5635 7451 5699 7452
rect 5229 7408 5248 7410
rect 5263 7408 5297 7410
rect 5229 7392 5309 7408
rect 5229 7386 5248 7392
rect 4945 7360 5048 7370
rect 4899 7358 5048 7360
rect 5069 7358 5104 7370
rect 4738 7356 4900 7358
rect 4750 7336 4769 7356
rect 4784 7354 4814 7356
rect 4633 7328 4674 7336
rect 4756 7332 4769 7336
rect 4821 7340 4900 7356
rect 4932 7356 5104 7358
rect 4932 7340 5011 7356
rect 5018 7354 5048 7356
rect 4596 7318 4625 7328
rect 4639 7318 4668 7328
rect 4683 7318 4713 7332
rect 4756 7318 4799 7332
rect 4821 7328 5011 7340
rect 5076 7336 5082 7356
rect 4806 7318 4836 7328
rect 4837 7318 4995 7328
rect 4999 7318 5029 7328
rect 5033 7318 5063 7332
rect 5091 7318 5104 7356
rect 5176 7370 5205 7386
rect 5219 7370 5248 7386
rect 5263 7376 5293 7392
rect 5321 7370 5327 7418
rect 5330 7412 5349 7418
rect 5364 7412 5394 7420
rect 5330 7404 5394 7412
rect 5330 7388 5410 7404
rect 5426 7397 5488 7428
rect 5504 7397 5566 7428
rect 5635 7426 5684 7451
rect 5699 7426 5729 7442
rect 5598 7412 5628 7420
rect 5635 7418 5745 7426
rect 5598 7404 5643 7412
rect 5330 7386 5349 7388
rect 5364 7386 5410 7388
rect 5330 7370 5410 7386
rect 5437 7384 5472 7397
rect 5513 7394 5550 7397
rect 5513 7392 5555 7394
rect 5442 7381 5472 7384
rect 5451 7377 5458 7381
rect 5458 7376 5459 7377
rect 5417 7370 5427 7376
rect 5176 7362 5211 7370
rect 5176 7336 5177 7362
rect 5184 7336 5211 7362
rect 5119 7318 5149 7332
rect 5176 7328 5211 7336
rect 5213 7362 5254 7370
rect 5213 7336 5228 7362
rect 5235 7336 5254 7362
rect 5318 7358 5349 7370
rect 5364 7358 5467 7370
rect 5479 7360 5505 7386
rect 5520 7381 5550 7392
rect 5582 7388 5644 7404
rect 5582 7386 5628 7388
rect 5582 7370 5644 7386
rect 5656 7370 5662 7418
rect 5665 7410 5745 7418
rect 5665 7408 5684 7410
rect 5699 7408 5733 7410
rect 5665 7392 5745 7408
rect 5665 7370 5684 7392
rect 5699 7376 5729 7392
rect 5757 7386 5763 7460
rect 5766 7386 5785 7530
rect 5800 7386 5806 7530
rect 5815 7460 5828 7530
rect 5880 7526 5902 7530
rect 5873 7504 5902 7518
rect 5955 7504 5971 7518
rect 6009 7514 6015 7516
rect 6022 7514 6130 7530
rect 6137 7514 6143 7516
rect 6151 7514 6166 7530
rect 6232 7524 6251 7527
rect 5873 7502 5971 7504
rect 5998 7502 6166 7514
rect 6181 7504 6197 7518
rect 6232 7505 6254 7524
rect 6264 7518 6280 7519
rect 6263 7516 6280 7518
rect 6264 7511 6280 7516
rect 6254 7504 6260 7505
rect 6263 7504 6292 7511
rect 6181 7503 6292 7504
rect 6181 7502 6298 7503
rect 5857 7494 5908 7502
rect 5955 7494 5989 7502
rect 5857 7482 5882 7494
rect 5889 7482 5908 7494
rect 5962 7492 5989 7494
rect 5998 7492 6219 7502
rect 6254 7499 6260 7502
rect 5962 7488 6219 7492
rect 5857 7474 5908 7482
rect 5955 7474 6219 7488
rect 6263 7494 6298 7502
rect 5809 7426 5828 7460
rect 5873 7466 5902 7474
rect 5873 7460 5890 7466
rect 5873 7458 5907 7460
rect 5955 7458 5971 7474
rect 5972 7464 6180 7474
rect 6181 7464 6197 7474
rect 6245 7470 6260 7485
rect 6263 7482 6264 7494
rect 6271 7482 6298 7494
rect 6263 7474 6298 7482
rect 6263 7473 6292 7474
rect 5983 7460 6197 7464
rect 5998 7458 6197 7460
rect 6232 7460 6245 7470
rect 6263 7460 6280 7473
rect 6232 7458 6280 7460
rect 5874 7454 5907 7458
rect 5870 7452 5907 7454
rect 5870 7451 5937 7452
rect 5870 7446 5901 7451
rect 5907 7446 5937 7451
rect 5870 7442 5937 7446
rect 5843 7439 5937 7442
rect 5843 7432 5892 7439
rect 5843 7426 5873 7432
rect 5892 7427 5897 7432
rect 5809 7410 5889 7426
rect 5901 7418 5937 7439
rect 5998 7434 6187 7458
rect 6232 7457 6279 7458
rect 6245 7452 6279 7457
rect 6013 7431 6187 7434
rect 6006 7428 6187 7431
rect 6215 7451 6279 7452
rect 5809 7408 5828 7410
rect 5843 7408 5877 7410
rect 5809 7392 5889 7408
rect 5809 7386 5828 7392
rect 5525 7360 5628 7370
rect 5479 7358 5628 7360
rect 5649 7358 5684 7370
rect 5318 7356 5480 7358
rect 5330 7336 5349 7356
rect 5364 7354 5394 7356
rect 5213 7328 5254 7336
rect 5336 7332 5349 7336
rect 5401 7340 5480 7356
rect 5512 7356 5684 7358
rect 5512 7340 5591 7356
rect 5598 7354 5628 7356
rect 5176 7318 5205 7328
rect 5219 7318 5248 7328
rect 5263 7318 5293 7332
rect 5336 7318 5379 7332
rect 5401 7328 5591 7340
rect 5656 7336 5662 7356
rect 5386 7318 5416 7328
rect 5417 7318 5575 7328
rect 5579 7318 5609 7328
rect 5613 7318 5643 7332
rect 5671 7318 5684 7356
rect 5756 7370 5785 7386
rect 5799 7370 5828 7386
rect 5843 7376 5873 7392
rect 5901 7370 5907 7418
rect 5910 7412 5929 7418
rect 5944 7412 5974 7420
rect 5910 7404 5974 7412
rect 5910 7388 5990 7404
rect 6006 7397 6068 7428
rect 6084 7397 6146 7428
rect 6215 7426 6264 7451
rect 6279 7426 6309 7442
rect 6178 7412 6208 7420
rect 6215 7418 6325 7426
rect 6178 7404 6223 7412
rect 5910 7386 5929 7388
rect 5944 7386 5990 7388
rect 5910 7370 5990 7386
rect 6017 7384 6052 7397
rect 6093 7394 6130 7397
rect 6093 7392 6135 7394
rect 6022 7381 6052 7384
rect 6031 7377 6038 7381
rect 6038 7376 6039 7377
rect 5997 7370 6007 7376
rect 5756 7362 5791 7370
rect 5756 7336 5757 7362
rect 5764 7336 5791 7362
rect 5699 7318 5729 7332
rect 5756 7328 5791 7336
rect 5793 7362 5834 7370
rect 5793 7336 5808 7362
rect 5815 7336 5834 7362
rect 5898 7358 5929 7370
rect 5944 7358 6047 7370
rect 6059 7360 6085 7386
rect 6100 7381 6130 7392
rect 6162 7388 6224 7404
rect 6162 7386 6208 7388
rect 6162 7370 6224 7386
rect 6236 7370 6242 7418
rect 6245 7410 6325 7418
rect 6245 7408 6264 7410
rect 6279 7408 6313 7410
rect 6245 7392 6325 7408
rect 6245 7370 6264 7392
rect 6279 7376 6309 7392
rect 6337 7386 6343 7460
rect 6346 7386 6365 7530
rect 6380 7386 6386 7530
rect 6395 7460 6408 7530
rect 6460 7526 6482 7530
rect 6453 7504 6482 7518
rect 6535 7504 6551 7518
rect 6589 7514 6595 7516
rect 6602 7514 6710 7530
rect 6717 7514 6723 7516
rect 6731 7514 6746 7530
rect 6812 7524 6831 7527
rect 6453 7502 6551 7504
rect 6578 7502 6746 7514
rect 6761 7504 6777 7518
rect 6812 7505 6834 7524
rect 6844 7518 6860 7519
rect 6843 7516 6860 7518
rect 6844 7511 6860 7516
rect 6834 7504 6840 7505
rect 6843 7504 6872 7511
rect 6761 7503 6872 7504
rect 6761 7502 6878 7503
rect 6437 7494 6488 7502
rect 6535 7494 6569 7502
rect 6437 7482 6462 7494
rect 6469 7482 6488 7494
rect 6542 7492 6569 7494
rect 6578 7492 6799 7502
rect 6834 7499 6840 7502
rect 6542 7488 6799 7492
rect 6437 7474 6488 7482
rect 6535 7474 6799 7488
rect 6843 7494 6878 7502
rect 6389 7426 6408 7460
rect 6453 7466 6482 7474
rect 6453 7460 6470 7466
rect 6453 7458 6487 7460
rect 6535 7458 6551 7474
rect 6552 7464 6760 7474
rect 6761 7464 6777 7474
rect 6825 7470 6840 7485
rect 6843 7482 6844 7494
rect 6851 7482 6878 7494
rect 6843 7474 6878 7482
rect 6843 7473 6872 7474
rect 6563 7460 6777 7464
rect 6578 7458 6777 7460
rect 6812 7460 6825 7470
rect 6843 7460 6860 7473
rect 6812 7458 6860 7460
rect 6454 7454 6487 7458
rect 6450 7452 6487 7454
rect 6450 7451 6517 7452
rect 6450 7446 6481 7451
rect 6487 7446 6517 7451
rect 6450 7442 6517 7446
rect 6423 7439 6517 7442
rect 6423 7432 6472 7439
rect 6423 7426 6453 7432
rect 6472 7427 6477 7432
rect 6389 7410 6469 7426
rect 6481 7418 6517 7439
rect 6578 7434 6767 7458
rect 6812 7457 6859 7458
rect 6825 7452 6859 7457
rect 6593 7431 6767 7434
rect 6586 7428 6767 7431
rect 6795 7451 6859 7452
rect 6389 7408 6408 7410
rect 6423 7408 6457 7410
rect 6389 7392 6469 7408
rect 6389 7386 6408 7392
rect 6105 7360 6208 7370
rect 6059 7358 6208 7360
rect 6229 7358 6264 7370
rect 5898 7356 6060 7358
rect 5910 7336 5929 7356
rect 5944 7354 5974 7356
rect 5793 7328 5834 7336
rect 5916 7332 5929 7336
rect 5981 7340 6060 7356
rect 6092 7356 6264 7358
rect 6092 7340 6171 7356
rect 6178 7354 6208 7356
rect 5756 7318 5785 7328
rect 5799 7318 5828 7328
rect 5843 7318 5873 7332
rect 5916 7318 5959 7332
rect 5981 7328 6171 7340
rect 6236 7336 6242 7356
rect 5966 7318 5996 7328
rect 5997 7318 6155 7328
rect 6159 7318 6189 7328
rect 6193 7318 6223 7332
rect 6251 7318 6264 7356
rect 6336 7370 6365 7386
rect 6379 7370 6408 7386
rect 6423 7376 6453 7392
rect 6481 7370 6487 7418
rect 6490 7412 6509 7418
rect 6524 7412 6554 7420
rect 6490 7404 6554 7412
rect 6490 7388 6570 7404
rect 6586 7397 6648 7428
rect 6664 7397 6726 7428
rect 6795 7426 6844 7451
rect 6859 7426 6889 7442
rect 6758 7412 6788 7420
rect 6795 7418 6905 7426
rect 6758 7404 6803 7412
rect 6490 7386 6509 7388
rect 6524 7386 6570 7388
rect 6490 7370 6570 7386
rect 6597 7384 6632 7397
rect 6673 7394 6710 7397
rect 6673 7392 6715 7394
rect 6602 7381 6632 7384
rect 6611 7377 6618 7381
rect 6618 7376 6619 7377
rect 6577 7370 6587 7376
rect 6336 7362 6371 7370
rect 6336 7336 6337 7362
rect 6344 7336 6371 7362
rect 6279 7318 6309 7332
rect 6336 7328 6371 7336
rect 6373 7362 6414 7370
rect 6373 7336 6388 7362
rect 6395 7336 6414 7362
rect 6478 7358 6509 7370
rect 6524 7358 6627 7370
rect 6639 7360 6665 7386
rect 6680 7381 6710 7392
rect 6742 7388 6804 7404
rect 6742 7386 6788 7388
rect 6742 7370 6804 7386
rect 6816 7370 6822 7418
rect 6825 7410 6905 7418
rect 6825 7408 6844 7410
rect 6859 7408 6893 7410
rect 6825 7392 6905 7408
rect 6825 7370 6844 7392
rect 6859 7376 6889 7392
rect 6917 7386 6923 7460
rect 6926 7386 6945 7530
rect 6960 7386 6966 7530
rect 6975 7460 6988 7530
rect 7040 7526 7062 7530
rect 7033 7504 7062 7518
rect 7115 7504 7131 7518
rect 7169 7514 7175 7516
rect 7182 7514 7290 7530
rect 7297 7514 7303 7516
rect 7311 7514 7326 7530
rect 7392 7524 7411 7527
rect 7033 7502 7131 7504
rect 7158 7502 7326 7514
rect 7341 7504 7357 7518
rect 7392 7505 7414 7524
rect 7424 7518 7440 7519
rect 7423 7516 7440 7518
rect 7424 7511 7440 7516
rect 7414 7504 7420 7505
rect 7423 7504 7452 7511
rect 7341 7503 7452 7504
rect 7341 7502 7458 7503
rect 7017 7494 7068 7502
rect 7115 7494 7149 7502
rect 7017 7482 7042 7494
rect 7049 7482 7068 7494
rect 7122 7492 7149 7494
rect 7158 7492 7379 7502
rect 7414 7499 7420 7502
rect 7122 7488 7379 7492
rect 7017 7474 7068 7482
rect 7115 7474 7379 7488
rect 7423 7494 7458 7502
rect 6969 7426 6988 7460
rect 7033 7466 7062 7474
rect 7033 7460 7050 7466
rect 7033 7458 7067 7460
rect 7115 7458 7131 7474
rect 7132 7464 7340 7474
rect 7341 7464 7357 7474
rect 7405 7470 7420 7485
rect 7423 7482 7424 7494
rect 7431 7482 7458 7494
rect 7423 7474 7458 7482
rect 7423 7473 7452 7474
rect 7143 7460 7357 7464
rect 7158 7458 7357 7460
rect 7392 7460 7405 7470
rect 7423 7460 7440 7473
rect 7392 7458 7440 7460
rect 7034 7454 7067 7458
rect 7030 7452 7067 7454
rect 7030 7451 7097 7452
rect 7030 7446 7061 7451
rect 7067 7446 7097 7451
rect 7030 7442 7097 7446
rect 7003 7439 7097 7442
rect 7003 7432 7052 7439
rect 7003 7426 7033 7432
rect 7052 7427 7057 7432
rect 6969 7410 7049 7426
rect 7061 7418 7097 7439
rect 7158 7434 7347 7458
rect 7392 7457 7439 7458
rect 7405 7452 7439 7457
rect 7173 7431 7347 7434
rect 7166 7428 7347 7431
rect 7375 7451 7439 7452
rect 6969 7408 6988 7410
rect 7003 7408 7037 7410
rect 6969 7392 7049 7408
rect 6969 7386 6988 7392
rect 6685 7360 6788 7370
rect 6639 7358 6788 7360
rect 6809 7358 6844 7370
rect 6478 7356 6640 7358
rect 6490 7336 6509 7356
rect 6524 7354 6554 7356
rect 6373 7328 6414 7336
rect 6496 7332 6509 7336
rect 6561 7340 6640 7356
rect 6672 7356 6844 7358
rect 6672 7340 6751 7356
rect 6758 7354 6788 7356
rect 6336 7318 6365 7328
rect 6379 7318 6408 7328
rect 6423 7318 6453 7332
rect 6496 7318 6539 7332
rect 6561 7328 6751 7340
rect 6816 7336 6822 7356
rect 6546 7318 6576 7328
rect 6577 7318 6735 7328
rect 6739 7318 6769 7328
rect 6773 7318 6803 7332
rect 6831 7318 6844 7356
rect 6916 7370 6945 7386
rect 6959 7370 6988 7386
rect 7003 7376 7033 7392
rect 7061 7370 7067 7418
rect 7070 7412 7089 7418
rect 7104 7412 7134 7420
rect 7070 7404 7134 7412
rect 7070 7388 7150 7404
rect 7166 7397 7228 7428
rect 7244 7397 7306 7428
rect 7375 7426 7424 7451
rect 7439 7426 7469 7442
rect 7338 7412 7368 7420
rect 7375 7418 7485 7426
rect 7338 7404 7383 7412
rect 7070 7386 7089 7388
rect 7104 7386 7150 7388
rect 7070 7370 7150 7386
rect 7177 7384 7212 7397
rect 7253 7394 7290 7397
rect 7253 7392 7295 7394
rect 7182 7381 7212 7384
rect 7191 7377 7198 7381
rect 7198 7376 7199 7377
rect 7157 7370 7167 7376
rect 6916 7362 6951 7370
rect 6916 7336 6917 7362
rect 6924 7336 6951 7362
rect 6859 7318 6889 7332
rect 6916 7328 6951 7336
rect 6953 7362 6994 7370
rect 6953 7336 6968 7362
rect 6975 7336 6994 7362
rect 7058 7358 7089 7370
rect 7104 7358 7207 7370
rect 7219 7360 7245 7386
rect 7260 7381 7290 7392
rect 7322 7388 7384 7404
rect 7322 7386 7368 7388
rect 7322 7370 7384 7386
rect 7396 7370 7402 7418
rect 7405 7410 7485 7418
rect 7405 7408 7424 7410
rect 7439 7408 7473 7410
rect 7405 7392 7485 7408
rect 7405 7370 7424 7392
rect 7439 7376 7469 7392
rect 7497 7386 7503 7460
rect 7506 7386 7525 7530
rect 7540 7386 7546 7530
rect 7555 7460 7568 7530
rect 7613 7508 7614 7518
rect 7629 7508 7642 7518
rect 7613 7504 7642 7508
rect 7647 7504 7677 7530
rect 7695 7516 7711 7518
rect 7783 7516 7836 7530
rect 7784 7514 7848 7516
rect 7891 7514 7906 7530
rect 7955 7527 7985 7530
rect 7955 7524 7991 7527
rect 7921 7516 7937 7518
rect 7695 7504 7710 7508
rect 7613 7502 7710 7504
rect 7738 7502 7906 7514
rect 7922 7504 7937 7508
rect 7955 7505 7994 7524
rect 8013 7518 8020 7519
rect 8019 7511 8020 7518
rect 8003 7508 8004 7511
rect 8019 7508 8032 7511
rect 7955 7504 7985 7505
rect 7994 7504 8000 7505
rect 8003 7504 8032 7508
rect 7922 7503 8032 7504
rect 7922 7502 8038 7503
rect 7597 7494 7648 7502
rect 7597 7482 7622 7494
rect 7629 7482 7648 7494
rect 7679 7494 7729 7502
rect 7679 7486 7695 7494
rect 7702 7492 7729 7494
rect 7738 7492 7959 7502
rect 7702 7482 7959 7492
rect 7988 7494 8038 7502
rect 7988 7485 8004 7494
rect 7597 7474 7648 7482
rect 7695 7474 7959 7482
rect 7985 7482 8004 7485
rect 8011 7482 8038 7494
rect 7985 7474 8038 7482
rect 7549 7426 7568 7460
rect 7613 7466 7614 7474
rect 7629 7466 7642 7474
rect 7613 7458 7629 7466
rect 7610 7451 7629 7454
rect 7610 7442 7632 7451
rect 7583 7432 7632 7442
rect 7583 7426 7613 7432
rect 7632 7427 7637 7432
rect 7549 7410 7629 7426
rect 7647 7418 7677 7474
rect 7712 7464 7920 7474
rect 7955 7470 8000 7474
rect 8003 7473 8004 7474
rect 8019 7473 8032 7474
rect 7738 7434 7927 7464
rect 7753 7431 7927 7434
rect 7746 7428 7927 7431
rect 7549 7408 7568 7410
rect 7583 7408 7617 7410
rect 7549 7392 7629 7408
rect 7656 7404 7669 7418
rect 7684 7404 7700 7420
rect 7746 7415 7757 7428
rect 7549 7386 7568 7392
rect 7265 7360 7368 7370
rect 7219 7358 7368 7360
rect 7389 7358 7424 7370
rect 7058 7356 7220 7358
rect 7070 7336 7089 7356
rect 7104 7354 7134 7356
rect 6953 7328 6994 7336
rect 7076 7332 7089 7336
rect 7141 7340 7220 7356
rect 7252 7356 7424 7358
rect 7252 7340 7331 7356
rect 7338 7354 7368 7356
rect 6916 7318 6945 7328
rect 6959 7318 6988 7328
rect 7003 7318 7033 7332
rect 7076 7318 7119 7332
rect 7141 7328 7331 7340
rect 7396 7336 7402 7356
rect 7126 7318 7156 7328
rect 7157 7318 7315 7328
rect 7319 7318 7349 7328
rect 7353 7318 7383 7332
rect 7411 7318 7424 7356
rect 7496 7370 7525 7386
rect 7539 7370 7568 7386
rect 7583 7370 7613 7392
rect 7656 7388 7718 7404
rect 7746 7397 7757 7413
rect 7762 7408 7772 7428
rect 7782 7408 7796 7428
rect 7799 7415 7808 7428
rect 7824 7415 7833 7428
rect 7762 7397 7796 7408
rect 7799 7397 7808 7413
rect 7824 7397 7833 7413
rect 7840 7408 7850 7428
rect 7860 7408 7874 7428
rect 7875 7415 7886 7428
rect 7840 7397 7874 7408
rect 7875 7397 7886 7413
rect 7932 7404 7948 7420
rect 7955 7418 7985 7470
rect 8019 7466 8020 7473
rect 8004 7458 8020 7466
rect 7991 7426 8004 7445
rect 8019 7426 8049 7442
rect 7991 7410 8065 7426
rect 7991 7408 8004 7410
rect 8019 7408 8053 7410
rect 7656 7386 7669 7388
rect 7684 7386 7718 7388
rect 7656 7370 7718 7386
rect 7762 7381 7778 7384
rect 7840 7381 7870 7392
rect 7918 7388 7964 7404
rect 7991 7392 8065 7408
rect 7918 7386 7952 7388
rect 7917 7370 7964 7386
rect 7991 7370 8004 7392
rect 8019 7370 8049 7392
rect 8076 7370 8077 7386
rect 8092 7370 8105 7530
rect 8135 7426 8148 7530
rect 8193 7508 8194 7518
rect 8209 7508 8222 7518
rect 8193 7504 8222 7508
rect 8227 7504 8257 7530
rect 8275 7516 8291 7518
rect 8363 7516 8416 7530
rect 8364 7514 8428 7516
rect 8471 7514 8486 7530
rect 8535 7527 8565 7530
rect 8535 7524 8571 7527
rect 8501 7516 8517 7518
rect 8275 7504 8290 7508
rect 8193 7502 8290 7504
rect 8318 7502 8486 7514
rect 8502 7504 8517 7508
rect 8535 7505 8574 7524
rect 8593 7518 8600 7519
rect 8599 7511 8600 7518
rect 8583 7508 8584 7511
rect 8599 7508 8612 7511
rect 8535 7504 8565 7505
rect 8574 7504 8580 7505
rect 8583 7504 8612 7508
rect 8502 7503 8612 7504
rect 8502 7502 8618 7503
rect 8177 7494 8228 7502
rect 8177 7482 8202 7494
rect 8209 7482 8228 7494
rect 8259 7494 8309 7502
rect 8259 7486 8275 7494
rect 8282 7492 8309 7494
rect 8318 7492 8539 7502
rect 8282 7482 8539 7492
rect 8568 7494 8618 7502
rect 8568 7485 8584 7494
rect 8177 7474 8228 7482
rect 8275 7474 8539 7482
rect 8565 7482 8584 7485
rect 8591 7482 8618 7494
rect 8565 7474 8618 7482
rect 8193 7466 8194 7474
rect 8209 7466 8222 7474
rect 8193 7458 8209 7466
rect 8190 7451 8209 7454
rect 8190 7442 8212 7451
rect 8163 7432 8212 7442
rect 8163 7426 8193 7432
rect 8212 7427 8217 7432
rect 8135 7410 8209 7426
rect 8227 7418 8257 7474
rect 8292 7464 8500 7474
rect 8535 7470 8580 7474
rect 8583 7473 8584 7474
rect 8599 7473 8612 7474
rect 8318 7434 8507 7464
rect 8333 7431 8507 7434
rect 8326 7428 8507 7431
rect 8135 7408 8148 7410
rect 8163 7408 8197 7410
rect 8135 7392 8209 7408
rect 8236 7404 8249 7418
rect 8264 7404 8280 7420
rect 8326 7415 8337 7428
rect 8119 7370 8120 7386
rect 8135 7370 8148 7392
rect 8163 7370 8193 7392
rect 8236 7388 8298 7404
rect 8326 7397 8337 7413
rect 8342 7408 8352 7428
rect 8362 7408 8376 7428
rect 8379 7415 8388 7428
rect 8404 7415 8413 7428
rect 8342 7397 8376 7408
rect 8379 7397 8388 7413
rect 8404 7397 8413 7413
rect 8420 7408 8430 7428
rect 8440 7408 8454 7428
rect 8455 7415 8466 7428
rect 8420 7397 8454 7408
rect 8455 7397 8466 7413
rect 8512 7404 8528 7420
rect 8535 7418 8565 7470
rect 8599 7466 8600 7473
rect 8584 7458 8600 7466
rect 8571 7426 8584 7445
rect 8599 7426 8629 7442
rect 8571 7410 8645 7426
rect 8571 7408 8584 7410
rect 8599 7408 8633 7410
rect 8236 7386 8249 7388
rect 8264 7386 8298 7388
rect 8236 7370 8298 7386
rect 8342 7381 8358 7384
rect 8420 7381 8450 7392
rect 8498 7388 8544 7404
rect 8571 7392 8645 7408
rect 8498 7386 8532 7388
rect 8497 7370 8544 7386
rect 8571 7370 8584 7392
rect 8599 7370 8629 7392
rect 8656 7370 8657 7386
rect 8672 7370 8685 7530
rect 8715 7426 8728 7530
rect 8773 7508 8774 7518
rect 8789 7508 8802 7518
rect 8773 7504 8802 7508
rect 8807 7504 8837 7530
rect 8855 7516 8871 7518
rect 8943 7516 8996 7530
rect 8944 7514 9008 7516
rect 9051 7514 9066 7530
rect 9115 7527 9145 7530
rect 9115 7524 9151 7527
rect 9081 7516 9097 7518
rect 8855 7504 8870 7508
rect 8773 7502 8870 7504
rect 8898 7502 9066 7514
rect 9082 7504 9097 7508
rect 9115 7505 9154 7524
rect 9173 7518 9180 7519
rect 9179 7511 9180 7518
rect 9163 7508 9164 7511
rect 9179 7508 9192 7511
rect 9115 7504 9145 7505
rect 9154 7504 9160 7505
rect 9163 7504 9192 7508
rect 9082 7503 9192 7504
rect 9082 7502 9198 7503
rect 8757 7494 8808 7502
rect 8757 7482 8782 7494
rect 8789 7482 8808 7494
rect 8839 7494 8889 7502
rect 8839 7486 8855 7494
rect 8862 7492 8889 7494
rect 8898 7492 9119 7502
rect 8862 7482 9119 7492
rect 9148 7494 9198 7502
rect 9148 7485 9164 7494
rect 8757 7474 8808 7482
rect 8855 7474 9119 7482
rect 9145 7482 9164 7485
rect 9171 7482 9198 7494
rect 9145 7474 9198 7482
rect 8773 7466 8774 7474
rect 8789 7466 8802 7474
rect 8773 7458 8789 7466
rect 8770 7451 8789 7454
rect 8770 7442 8792 7451
rect 8743 7432 8792 7442
rect 8743 7426 8773 7432
rect 8792 7427 8797 7432
rect 8715 7410 8789 7426
rect 8807 7418 8837 7474
rect 8872 7464 9080 7474
rect 9115 7470 9160 7474
rect 9163 7473 9164 7474
rect 9179 7473 9192 7474
rect 8898 7434 9087 7464
rect 8913 7431 9087 7434
rect 8906 7428 9087 7431
rect 8715 7408 8728 7410
rect 8743 7408 8777 7410
rect 8715 7392 8789 7408
rect 8816 7404 8829 7418
rect 8844 7404 8860 7420
rect 8906 7415 8917 7428
rect 8699 7370 8700 7386
rect 8715 7370 8728 7392
rect 8743 7370 8773 7392
rect 8816 7388 8878 7404
rect 8906 7397 8917 7413
rect 8922 7408 8932 7428
rect 8942 7408 8956 7428
rect 8959 7415 8968 7428
rect 8984 7415 8993 7428
rect 8922 7397 8956 7408
rect 8959 7397 8968 7413
rect 8984 7397 8993 7413
rect 9000 7408 9010 7428
rect 9020 7408 9034 7428
rect 9035 7415 9046 7428
rect 9000 7397 9034 7408
rect 9035 7397 9046 7413
rect 9092 7404 9108 7420
rect 9115 7418 9145 7470
rect 9179 7466 9180 7473
rect 9164 7458 9180 7466
rect 9151 7426 9164 7445
rect 9179 7426 9209 7442
rect 9151 7410 9225 7426
rect 9151 7408 9164 7410
rect 9179 7408 9213 7410
rect 8816 7386 8829 7388
rect 8844 7386 8878 7388
rect 8816 7370 8878 7386
rect 8922 7381 8938 7384
rect 9000 7381 9030 7392
rect 9078 7388 9124 7404
rect 9151 7392 9225 7408
rect 9078 7386 9112 7388
rect 9077 7370 9124 7386
rect 9151 7370 9164 7392
rect 9179 7370 9209 7392
rect 9236 7370 9237 7386
rect 9252 7370 9265 7530
rect 7496 7362 7531 7370
rect 7496 7336 7497 7362
rect 7504 7336 7531 7362
rect 7439 7318 7469 7332
rect 7496 7328 7531 7336
rect 7533 7362 7574 7370
rect 7533 7336 7548 7362
rect 7555 7336 7574 7362
rect 7638 7358 7700 7370
rect 7712 7358 7787 7370
rect 7845 7358 7920 7370
rect 7932 7358 7963 7370
rect 7969 7358 8004 7370
rect 7638 7356 7800 7358
rect 7533 7328 7574 7336
rect 7656 7332 7669 7356
rect 7684 7354 7699 7356
rect 7496 7318 7525 7328
rect 7539 7318 7568 7328
rect 7583 7318 7613 7332
rect 7656 7318 7699 7332
rect 7723 7329 7730 7336
rect 7733 7332 7800 7356
rect 7832 7356 8004 7358
rect 7802 7334 7830 7338
rect 7832 7334 7912 7356
rect 7933 7354 7948 7356
rect 7802 7332 7912 7334
rect 7733 7328 7912 7332
rect 7706 7318 7736 7328
rect 7738 7318 7891 7328
rect 7899 7318 7929 7328
rect 7933 7318 7963 7332
rect 7991 7318 8004 7356
rect 8076 7362 8111 7370
rect 8076 7336 8077 7362
rect 8084 7336 8111 7362
rect 8019 7318 8049 7332
rect 8076 7328 8111 7336
rect 8113 7362 8154 7370
rect 8113 7336 8128 7362
rect 8135 7336 8154 7362
rect 8218 7358 8280 7370
rect 8292 7358 8367 7370
rect 8425 7358 8500 7370
rect 8512 7358 8543 7370
rect 8549 7358 8584 7370
rect 8218 7356 8380 7358
rect 8113 7328 8154 7336
rect 8236 7332 8249 7356
rect 8264 7354 8279 7356
rect 8076 7318 8077 7328
rect 8092 7318 8105 7328
rect 8119 7318 8120 7328
rect 8135 7318 8148 7328
rect 8163 7318 8193 7332
rect 8236 7318 8279 7332
rect 8303 7329 8310 7336
rect 8313 7332 8380 7356
rect 8412 7356 8584 7358
rect 8382 7334 8410 7338
rect 8412 7334 8492 7356
rect 8513 7354 8528 7356
rect 8382 7332 8492 7334
rect 8313 7328 8492 7332
rect 8286 7318 8316 7328
rect 8318 7318 8471 7328
rect 8479 7318 8509 7328
rect 8513 7318 8543 7332
rect 8571 7318 8584 7356
rect 8656 7362 8691 7370
rect 8656 7336 8657 7362
rect 8664 7336 8691 7362
rect 8599 7318 8629 7332
rect 8656 7328 8691 7336
rect 8693 7362 8734 7370
rect 8693 7336 8708 7362
rect 8715 7336 8734 7362
rect 8798 7358 8860 7370
rect 8872 7358 8947 7370
rect 9005 7358 9080 7370
rect 9092 7358 9123 7370
rect 9129 7358 9164 7370
rect 8798 7356 8960 7358
rect 8693 7328 8734 7336
rect 8816 7332 8829 7356
rect 8844 7354 8859 7356
rect 8656 7318 8657 7328
rect 8672 7318 8685 7328
rect 8699 7318 8700 7328
rect 8715 7318 8728 7328
rect 8743 7318 8773 7332
rect 8816 7318 8859 7332
rect 8883 7329 8890 7336
rect 8893 7332 8960 7356
rect 8992 7356 9164 7358
rect 8962 7334 8990 7338
rect 8992 7334 9072 7356
rect 9093 7354 9108 7356
rect 8962 7332 9072 7334
rect 8893 7328 9072 7332
rect 8866 7318 8896 7328
rect 8898 7318 9051 7328
rect 9059 7318 9089 7328
rect 9093 7318 9123 7332
rect 9151 7318 9164 7356
rect 9236 7362 9271 7370
rect 9236 7336 9237 7362
rect 9244 7336 9271 7362
rect 9179 7318 9209 7332
rect 9236 7328 9271 7336
rect 9236 7318 9237 7328
rect 9252 7318 9265 7328
rect -1 7312 9265 7318
rect 0 7304 9265 7312
rect 15 7274 28 7304
rect 43 7286 73 7304
rect 116 7290 130 7304
rect 166 7290 386 7304
rect 117 7288 130 7290
rect 83 7276 98 7288
rect 80 7274 102 7276
rect 107 7274 137 7288
rect 198 7286 351 7290
rect 180 7274 372 7286
rect 415 7274 445 7288
rect 451 7274 464 7304
rect 479 7286 509 7304
rect 552 7274 565 7304
rect 595 7274 608 7304
rect 623 7286 653 7304
rect 696 7290 710 7304
rect 746 7290 966 7304
rect 697 7288 710 7290
rect 663 7276 678 7288
rect 660 7274 682 7276
rect 687 7274 717 7288
rect 778 7286 931 7290
rect 760 7274 952 7286
rect 995 7274 1025 7288
rect 1031 7274 1044 7304
rect 1059 7286 1089 7304
rect 1132 7274 1145 7304
rect 1175 7274 1188 7304
rect 1203 7286 1233 7304
rect 1276 7290 1290 7304
rect 1326 7290 1546 7304
rect 1277 7288 1290 7290
rect 1243 7276 1258 7288
rect 1240 7274 1262 7276
rect 1267 7274 1297 7288
rect 1358 7286 1511 7290
rect 1340 7274 1532 7286
rect 1575 7274 1605 7288
rect 1611 7274 1624 7304
rect 1639 7286 1669 7304
rect 1712 7274 1725 7304
rect 1755 7274 1768 7304
rect 1783 7290 1813 7304
rect 1856 7290 1899 7304
rect 1906 7290 2126 7304
rect 2133 7290 2163 7304
rect 1823 7276 1838 7288
rect 1857 7276 1870 7290
rect 1938 7286 2091 7290
rect 1820 7274 1842 7276
rect 1920 7274 2112 7286
rect 2191 7274 2204 7304
rect 2219 7290 2249 7304
rect 2286 7274 2305 7304
rect 2320 7274 2326 7304
rect 2335 7274 2348 7304
rect 2363 7290 2393 7304
rect 2436 7290 2479 7304
rect 2486 7290 2706 7304
rect 2713 7290 2743 7304
rect 2403 7276 2418 7288
rect 2437 7276 2450 7290
rect 2518 7286 2671 7290
rect 2400 7274 2422 7276
rect 2500 7274 2692 7286
rect 2771 7274 2784 7304
rect 2799 7290 2829 7304
rect 2866 7274 2885 7304
rect 2900 7274 2906 7304
rect 2915 7274 2928 7304
rect 2943 7290 2973 7304
rect 3016 7290 3059 7304
rect 3066 7290 3286 7304
rect 3293 7290 3323 7304
rect 2983 7276 2998 7288
rect 3017 7276 3030 7290
rect 3098 7286 3251 7290
rect 2980 7274 3002 7276
rect 3080 7274 3272 7286
rect 3351 7274 3364 7304
rect 3379 7290 3409 7304
rect 3446 7274 3465 7304
rect 3480 7274 3486 7304
rect 3495 7274 3508 7304
rect 3523 7290 3553 7304
rect 3596 7290 3639 7304
rect 3646 7290 3866 7304
rect 3873 7290 3903 7304
rect 3563 7276 3578 7288
rect 3597 7276 3610 7290
rect 3678 7286 3831 7290
rect 3560 7274 3582 7276
rect 3660 7274 3852 7286
rect 3931 7274 3944 7304
rect 3959 7290 3989 7304
rect 4026 7274 4045 7304
rect 4060 7274 4066 7304
rect 4075 7274 4088 7304
rect 4103 7290 4133 7304
rect 4176 7290 4219 7304
rect 4226 7290 4446 7304
rect 4453 7290 4483 7304
rect 4143 7276 4158 7288
rect 4177 7276 4190 7290
rect 4258 7286 4411 7290
rect 4140 7274 4162 7276
rect 4240 7274 4432 7286
rect 4511 7274 4524 7304
rect 4539 7290 4569 7304
rect 4606 7274 4625 7304
rect 4640 7274 4646 7304
rect 4655 7274 4668 7304
rect 4683 7290 4713 7304
rect 4756 7290 4799 7304
rect 4806 7290 5026 7304
rect 5033 7290 5063 7304
rect 4723 7276 4738 7288
rect 4757 7276 4770 7290
rect 4838 7286 4991 7290
rect 4720 7274 4742 7276
rect 4820 7274 5012 7286
rect 5091 7274 5104 7304
rect 5119 7290 5149 7304
rect 5186 7274 5205 7304
rect 5220 7274 5226 7304
rect 5235 7274 5248 7304
rect 5263 7290 5293 7304
rect 5336 7290 5379 7304
rect 5386 7290 5606 7304
rect 5613 7290 5643 7304
rect 5303 7276 5318 7288
rect 5337 7276 5350 7290
rect 5418 7286 5571 7290
rect 5300 7274 5322 7276
rect 5400 7274 5592 7286
rect 5671 7274 5684 7304
rect 5699 7290 5729 7304
rect 5766 7274 5785 7304
rect 5800 7274 5806 7304
rect 5815 7274 5828 7304
rect 5843 7290 5873 7304
rect 5916 7290 5959 7304
rect 5966 7290 6186 7304
rect 6193 7290 6223 7304
rect 5883 7276 5898 7288
rect 5917 7276 5930 7290
rect 5998 7286 6151 7290
rect 5880 7274 5902 7276
rect 5980 7274 6172 7286
rect 6251 7274 6264 7304
rect 6279 7290 6309 7304
rect 6346 7274 6365 7304
rect 6380 7274 6386 7304
rect 6395 7274 6408 7304
rect 6423 7290 6453 7304
rect 6496 7290 6539 7304
rect 6546 7290 6766 7304
rect 6773 7290 6803 7304
rect 6463 7276 6478 7288
rect 6497 7276 6510 7290
rect 6578 7286 6731 7290
rect 6460 7274 6482 7276
rect 6560 7274 6752 7286
rect 6831 7274 6844 7304
rect 6859 7290 6889 7304
rect 6926 7274 6945 7304
rect 6960 7274 6966 7304
rect 6975 7274 6988 7304
rect 7003 7290 7033 7304
rect 7076 7290 7119 7304
rect 7126 7290 7346 7304
rect 7353 7290 7383 7304
rect 7043 7276 7058 7288
rect 7077 7276 7090 7290
rect 7158 7286 7311 7290
rect 7040 7274 7062 7276
rect 7140 7274 7332 7286
rect 7411 7274 7424 7304
rect 7439 7290 7469 7304
rect 7506 7274 7525 7304
rect 7540 7274 7546 7304
rect 7555 7274 7568 7304
rect 7583 7286 7613 7304
rect 7656 7290 7670 7304
rect 7706 7290 7926 7304
rect 7657 7288 7670 7290
rect 7623 7276 7638 7288
rect 7620 7274 7642 7276
rect 7647 7274 7677 7288
rect 7738 7286 7891 7290
rect 7720 7274 7912 7286
rect 7955 7274 7985 7288
rect 7991 7274 8004 7304
rect 8019 7286 8049 7304
rect 8092 7274 8105 7304
rect 8135 7274 8148 7304
rect 8163 7286 8193 7304
rect 8236 7290 8250 7304
rect 8286 7290 8506 7304
rect 8237 7288 8250 7290
rect 8203 7276 8218 7288
rect 8200 7274 8222 7276
rect 8227 7274 8257 7288
rect 8318 7286 8471 7290
rect 8300 7274 8492 7286
rect 8535 7274 8565 7288
rect 8571 7274 8584 7304
rect 8599 7286 8629 7304
rect 8672 7274 8685 7304
rect 8715 7274 8728 7304
rect 8743 7286 8773 7304
rect 8816 7290 8830 7304
rect 8866 7290 9086 7304
rect 8817 7288 8830 7290
rect 8783 7276 8798 7288
rect 8780 7274 8802 7276
rect 8807 7274 8837 7288
rect 8898 7286 9051 7290
rect 8880 7274 9072 7286
rect 9115 7274 9145 7288
rect 9151 7274 9164 7304
rect 9179 7286 9209 7304
rect 9252 7274 9265 7304
rect 0 7260 9265 7274
rect 15 7156 28 7260
rect 73 7238 74 7248
rect 89 7238 102 7248
rect 73 7234 102 7238
rect 107 7234 137 7260
rect 155 7246 171 7248
rect 243 7246 296 7260
rect 244 7244 308 7246
rect 351 7244 366 7260
rect 415 7257 445 7260
rect 415 7254 451 7257
rect 381 7246 397 7248
rect 155 7234 170 7238
rect 73 7232 170 7234
rect 198 7232 366 7244
rect 382 7234 397 7238
rect 415 7235 454 7254
rect 473 7248 480 7249
rect 479 7241 480 7248
rect 463 7238 464 7241
rect 479 7238 492 7241
rect 415 7234 445 7235
rect 454 7234 460 7235
rect 463 7234 492 7238
rect 382 7233 492 7234
rect 382 7232 498 7233
rect 57 7224 108 7232
rect 57 7212 82 7224
rect 89 7212 108 7224
rect 139 7224 189 7232
rect 139 7216 155 7224
rect 162 7222 189 7224
rect 198 7222 419 7232
rect 162 7212 419 7222
rect 448 7224 498 7232
rect 448 7215 464 7224
rect 57 7204 108 7212
rect 155 7204 419 7212
rect 445 7212 464 7215
rect 471 7212 498 7224
rect 445 7204 498 7212
rect 73 7196 74 7204
rect 89 7196 102 7204
rect 73 7188 89 7196
rect 70 7181 89 7184
rect 70 7172 92 7181
rect 43 7162 92 7172
rect 43 7156 73 7162
rect 92 7157 97 7162
rect 15 7140 89 7156
rect 107 7148 137 7204
rect 172 7194 380 7204
rect 415 7200 460 7204
rect 463 7203 464 7204
rect 479 7203 492 7204
rect 198 7164 387 7194
rect 213 7161 387 7164
rect 206 7158 387 7161
rect 15 7138 28 7140
rect 43 7138 77 7140
rect 15 7122 89 7138
rect 116 7134 129 7148
rect 144 7134 160 7150
rect 206 7145 217 7158
rect -1 7100 0 7116
rect 15 7100 28 7122
rect 43 7100 73 7122
rect 116 7118 178 7134
rect 206 7127 217 7143
rect 222 7138 232 7158
rect 242 7138 256 7158
rect 259 7145 268 7158
rect 284 7145 293 7158
rect 222 7127 256 7138
rect 259 7127 268 7143
rect 284 7127 293 7143
rect 300 7138 310 7158
rect 320 7138 334 7158
rect 335 7145 346 7158
rect 300 7127 334 7138
rect 335 7127 346 7143
rect 392 7134 408 7150
rect 415 7148 445 7200
rect 479 7196 480 7203
rect 464 7188 480 7196
rect 451 7156 464 7175
rect 479 7156 509 7172
rect 451 7140 525 7156
rect 451 7138 464 7140
rect 479 7138 513 7140
rect 116 7116 129 7118
rect 144 7116 178 7118
rect 116 7100 178 7116
rect 222 7111 238 7114
rect 300 7111 330 7122
rect 378 7118 424 7134
rect 451 7122 525 7138
rect 378 7116 412 7118
rect 377 7100 424 7116
rect 451 7100 464 7122
rect 479 7100 509 7122
rect 536 7100 537 7116
rect 552 7100 565 7260
rect 595 7156 608 7260
rect 653 7238 654 7248
rect 669 7238 682 7248
rect 653 7234 682 7238
rect 687 7234 717 7260
rect 735 7246 751 7248
rect 823 7246 876 7260
rect 824 7244 888 7246
rect 931 7244 946 7260
rect 995 7257 1025 7260
rect 995 7254 1031 7257
rect 961 7246 977 7248
rect 735 7234 750 7238
rect 653 7232 750 7234
rect 778 7232 946 7244
rect 962 7234 977 7238
rect 995 7235 1034 7254
rect 1053 7248 1060 7249
rect 1059 7241 1060 7248
rect 1043 7238 1044 7241
rect 1059 7238 1072 7241
rect 995 7234 1025 7235
rect 1034 7234 1040 7235
rect 1043 7234 1072 7238
rect 962 7233 1072 7234
rect 962 7232 1078 7233
rect 637 7224 688 7232
rect 637 7212 662 7224
rect 669 7212 688 7224
rect 719 7224 769 7232
rect 719 7216 735 7224
rect 742 7222 769 7224
rect 778 7222 999 7232
rect 742 7212 999 7222
rect 1028 7224 1078 7232
rect 1028 7215 1044 7224
rect 637 7204 688 7212
rect 735 7204 999 7212
rect 1025 7212 1044 7215
rect 1051 7212 1078 7224
rect 1025 7204 1078 7212
rect 653 7196 654 7204
rect 669 7196 682 7204
rect 653 7188 669 7196
rect 650 7181 669 7184
rect 650 7172 672 7181
rect 623 7162 672 7172
rect 623 7156 653 7162
rect 672 7157 677 7162
rect 595 7140 669 7156
rect 687 7148 717 7204
rect 752 7194 960 7204
rect 995 7200 1040 7204
rect 1043 7203 1044 7204
rect 1059 7203 1072 7204
rect 778 7164 967 7194
rect 793 7161 967 7164
rect 786 7158 967 7161
rect 595 7138 608 7140
rect 623 7138 657 7140
rect 595 7122 669 7138
rect 696 7134 709 7148
rect 724 7134 740 7150
rect 786 7145 797 7158
rect 579 7100 580 7116
rect 595 7100 608 7122
rect 623 7100 653 7122
rect 696 7118 758 7134
rect 786 7127 797 7143
rect 802 7138 812 7158
rect 822 7138 836 7158
rect 839 7145 848 7158
rect 864 7145 873 7158
rect 802 7127 836 7138
rect 839 7127 848 7143
rect 864 7127 873 7143
rect 880 7138 890 7158
rect 900 7138 914 7158
rect 915 7145 926 7158
rect 880 7127 914 7138
rect 915 7127 926 7143
rect 972 7134 988 7150
rect 995 7148 1025 7200
rect 1059 7196 1060 7203
rect 1044 7188 1060 7196
rect 1031 7156 1044 7175
rect 1059 7156 1089 7172
rect 1031 7140 1105 7156
rect 1031 7138 1044 7140
rect 1059 7138 1093 7140
rect 696 7116 709 7118
rect 724 7116 758 7118
rect 696 7100 758 7116
rect 802 7111 818 7114
rect 880 7111 910 7122
rect 958 7118 1004 7134
rect 1031 7122 1105 7138
rect 958 7116 992 7118
rect 957 7100 1004 7116
rect 1031 7100 1044 7122
rect 1059 7100 1089 7122
rect 1116 7100 1117 7116
rect 1132 7100 1145 7260
rect 1175 7156 1188 7260
rect 1233 7238 1234 7248
rect 1249 7238 1262 7248
rect 1233 7234 1262 7238
rect 1267 7234 1297 7260
rect 1315 7246 1331 7248
rect 1403 7246 1456 7260
rect 1404 7244 1468 7246
rect 1511 7244 1526 7260
rect 1575 7257 1605 7260
rect 1575 7254 1611 7257
rect 1541 7246 1557 7248
rect 1315 7234 1330 7238
rect 1233 7232 1330 7234
rect 1358 7232 1526 7244
rect 1542 7234 1557 7238
rect 1575 7235 1614 7254
rect 1633 7248 1640 7249
rect 1639 7241 1640 7248
rect 1623 7238 1624 7241
rect 1639 7238 1652 7241
rect 1575 7234 1605 7235
rect 1614 7234 1620 7235
rect 1623 7234 1652 7238
rect 1542 7233 1652 7234
rect 1542 7232 1658 7233
rect 1217 7224 1268 7232
rect 1217 7212 1242 7224
rect 1249 7212 1268 7224
rect 1299 7224 1349 7232
rect 1299 7216 1315 7224
rect 1322 7222 1349 7224
rect 1358 7222 1579 7232
rect 1322 7212 1579 7222
rect 1608 7224 1658 7232
rect 1608 7215 1624 7224
rect 1217 7204 1268 7212
rect 1315 7204 1579 7212
rect 1605 7212 1624 7215
rect 1631 7212 1658 7224
rect 1605 7204 1658 7212
rect 1233 7196 1234 7204
rect 1249 7196 1262 7204
rect 1233 7188 1249 7196
rect 1230 7181 1249 7184
rect 1230 7172 1252 7181
rect 1203 7162 1252 7172
rect 1203 7156 1233 7162
rect 1252 7157 1257 7162
rect 1175 7140 1249 7156
rect 1267 7148 1297 7204
rect 1332 7194 1540 7204
rect 1575 7200 1620 7204
rect 1623 7203 1624 7204
rect 1639 7203 1652 7204
rect 1358 7164 1547 7194
rect 1373 7161 1547 7164
rect 1366 7158 1547 7161
rect 1175 7138 1188 7140
rect 1203 7138 1237 7140
rect 1175 7122 1249 7138
rect 1276 7134 1289 7148
rect 1304 7134 1320 7150
rect 1366 7145 1377 7158
rect 1159 7100 1160 7116
rect 1175 7100 1188 7122
rect 1203 7100 1233 7122
rect 1276 7118 1338 7134
rect 1366 7127 1377 7143
rect 1382 7138 1392 7158
rect 1402 7138 1416 7158
rect 1419 7145 1428 7158
rect 1444 7145 1453 7158
rect 1382 7127 1416 7138
rect 1419 7127 1428 7143
rect 1444 7127 1453 7143
rect 1460 7138 1470 7158
rect 1480 7138 1494 7158
rect 1495 7145 1506 7158
rect 1460 7127 1494 7138
rect 1495 7127 1506 7143
rect 1552 7134 1568 7150
rect 1575 7148 1605 7200
rect 1639 7196 1640 7203
rect 1624 7188 1640 7196
rect 1611 7156 1624 7175
rect 1639 7156 1669 7172
rect 1611 7140 1685 7156
rect 1611 7138 1624 7140
rect 1639 7138 1673 7140
rect 1276 7116 1289 7118
rect 1304 7116 1338 7118
rect 1276 7100 1338 7116
rect 1382 7111 1398 7114
rect 1460 7111 1490 7122
rect 1538 7118 1584 7134
rect 1611 7122 1685 7138
rect 1538 7116 1572 7118
rect 1537 7100 1584 7116
rect 1611 7100 1624 7122
rect 1639 7100 1669 7122
rect 1696 7100 1697 7116
rect 1712 7100 1725 7260
rect 1755 7156 1768 7260
rect 1820 7256 1842 7260
rect 1813 7234 1842 7248
rect 1895 7234 1911 7248
rect 1949 7244 1955 7246
rect 1962 7244 2070 7260
rect 2077 7244 2083 7246
rect 2091 7244 2106 7260
rect 2172 7254 2191 7257
rect 1813 7232 1911 7234
rect 1938 7232 2106 7244
rect 2121 7234 2137 7248
rect 2172 7235 2194 7254
rect 2204 7248 2220 7249
rect 2203 7246 2220 7248
rect 2204 7241 2220 7246
rect 2194 7234 2200 7235
rect 2203 7234 2232 7241
rect 2121 7233 2232 7234
rect 2121 7232 2238 7233
rect 1797 7224 1848 7232
rect 1895 7224 1929 7232
rect 1797 7212 1822 7224
rect 1829 7212 1848 7224
rect 1902 7222 1929 7224
rect 1938 7222 2159 7232
rect 2194 7229 2200 7232
rect 1902 7218 2159 7222
rect 1797 7204 1848 7212
rect 1895 7204 2159 7218
rect 2203 7224 2238 7232
rect 1813 7196 1842 7204
rect 1813 7190 1830 7196
rect 1813 7188 1847 7190
rect 1895 7188 1911 7204
rect 1912 7194 2120 7204
rect 2121 7194 2137 7204
rect 2185 7200 2200 7215
rect 2203 7212 2204 7224
rect 2211 7212 2238 7224
rect 2203 7204 2238 7212
rect 2203 7203 2232 7204
rect 1923 7190 2137 7194
rect 1938 7188 2137 7190
rect 2172 7190 2185 7200
rect 2203 7190 2220 7203
rect 2172 7188 2220 7190
rect 1814 7184 1847 7188
rect 1810 7182 1847 7184
rect 1810 7181 1877 7182
rect 1810 7176 1841 7181
rect 1847 7176 1877 7181
rect 1810 7172 1877 7176
rect 1783 7169 1877 7172
rect 1783 7162 1832 7169
rect 1783 7156 1813 7162
rect 1832 7157 1837 7162
rect 1755 7140 1829 7156
rect 1841 7148 1877 7169
rect 1938 7164 2127 7188
rect 2172 7187 2219 7188
rect 2185 7182 2219 7187
rect 1953 7161 2127 7164
rect 1946 7158 2127 7161
rect 2155 7181 2219 7182
rect 1755 7138 1768 7140
rect 1783 7138 1817 7140
rect 1755 7122 1829 7138
rect 1739 7100 1740 7116
rect 1755 7100 1768 7122
rect 1783 7106 1813 7122
rect 1841 7100 1847 7148
rect 1850 7142 1869 7148
rect 1884 7142 1914 7150
rect 1850 7134 1914 7142
rect 1850 7118 1930 7134
rect 1946 7127 2008 7158
rect 2024 7127 2086 7158
rect 2155 7156 2204 7181
rect 2219 7156 2249 7172
rect 2118 7142 2148 7150
rect 2155 7148 2265 7156
rect 2118 7134 2163 7142
rect 1850 7116 1869 7118
rect 1884 7116 1930 7118
rect 1850 7100 1930 7116
rect 1957 7114 1992 7127
rect 2033 7124 2070 7127
rect 2033 7122 2075 7124
rect 1962 7111 1992 7114
rect 1971 7107 1978 7111
rect 1978 7106 1979 7107
rect 1937 7100 1947 7106
rect -7 7092 34 7100
rect -7 7066 8 7092
rect 15 7066 34 7092
rect 98 7088 160 7100
rect 172 7088 247 7100
rect 305 7088 380 7100
rect 392 7088 423 7100
rect 429 7088 464 7100
rect 98 7086 260 7088
rect -7 7058 34 7066
rect 116 7062 129 7086
rect 144 7084 159 7086
rect -1 7048 0 7058
rect 15 7048 28 7058
rect 43 7048 73 7062
rect 116 7048 159 7062
rect 183 7059 190 7066
rect 193 7062 260 7086
rect 292 7086 464 7088
rect 262 7064 290 7068
rect 292 7064 372 7086
rect 393 7084 408 7086
rect 262 7062 372 7064
rect 193 7058 372 7062
rect 166 7048 196 7058
rect 198 7048 351 7058
rect 359 7048 389 7058
rect 393 7048 423 7062
rect 451 7048 464 7086
rect 536 7092 571 7100
rect 536 7066 537 7092
rect 544 7066 571 7092
rect 479 7048 509 7062
rect 536 7058 571 7066
rect 573 7092 614 7100
rect 573 7066 588 7092
rect 595 7066 614 7092
rect 678 7088 740 7100
rect 752 7088 827 7100
rect 885 7088 960 7100
rect 972 7088 1003 7100
rect 1009 7088 1044 7100
rect 678 7086 840 7088
rect 573 7058 614 7066
rect 696 7062 709 7086
rect 724 7084 739 7086
rect 536 7048 537 7058
rect 552 7048 565 7058
rect 579 7048 580 7058
rect 595 7048 608 7058
rect 623 7048 653 7062
rect 696 7048 739 7062
rect 763 7059 770 7066
rect 773 7062 840 7086
rect 872 7086 1044 7088
rect 842 7064 870 7068
rect 872 7064 952 7086
rect 973 7084 988 7086
rect 842 7062 952 7064
rect 773 7058 952 7062
rect 746 7048 776 7058
rect 778 7048 931 7058
rect 939 7048 969 7058
rect 973 7048 1003 7062
rect 1031 7048 1044 7086
rect 1116 7092 1151 7100
rect 1116 7066 1117 7092
rect 1124 7066 1151 7092
rect 1059 7048 1089 7062
rect 1116 7058 1151 7066
rect 1153 7092 1194 7100
rect 1153 7066 1168 7092
rect 1175 7066 1194 7092
rect 1258 7088 1320 7100
rect 1332 7088 1407 7100
rect 1465 7088 1540 7100
rect 1552 7088 1583 7100
rect 1589 7088 1624 7100
rect 1258 7086 1420 7088
rect 1153 7058 1194 7066
rect 1276 7062 1289 7086
rect 1304 7084 1319 7086
rect 1116 7048 1117 7058
rect 1132 7048 1145 7058
rect 1159 7048 1160 7058
rect 1175 7048 1188 7058
rect 1203 7048 1233 7062
rect 1276 7048 1319 7062
rect 1343 7059 1350 7066
rect 1353 7062 1420 7086
rect 1452 7086 1624 7088
rect 1422 7064 1450 7068
rect 1452 7064 1532 7086
rect 1553 7084 1568 7086
rect 1422 7062 1532 7064
rect 1353 7058 1532 7062
rect 1326 7048 1356 7058
rect 1358 7048 1511 7058
rect 1519 7048 1549 7058
rect 1553 7048 1583 7062
rect 1611 7048 1624 7086
rect 1696 7092 1731 7100
rect 1696 7066 1697 7092
rect 1704 7066 1731 7092
rect 1639 7048 1669 7062
rect 1696 7058 1731 7066
rect 1733 7092 1774 7100
rect 1733 7066 1748 7092
rect 1755 7066 1774 7092
rect 1838 7088 1869 7100
rect 1884 7088 1987 7100
rect 1999 7090 2025 7116
rect 2040 7111 2070 7122
rect 2102 7118 2164 7134
rect 2102 7116 2148 7118
rect 2102 7100 2164 7116
rect 2176 7100 2182 7148
rect 2185 7140 2265 7148
rect 2185 7138 2204 7140
rect 2219 7138 2253 7140
rect 2185 7122 2265 7138
rect 2185 7100 2204 7122
rect 2219 7106 2249 7122
rect 2277 7116 2283 7190
rect 2286 7116 2305 7260
rect 2320 7116 2326 7260
rect 2335 7190 2348 7260
rect 2400 7256 2422 7260
rect 2393 7234 2422 7248
rect 2475 7234 2491 7248
rect 2529 7244 2535 7246
rect 2542 7244 2650 7260
rect 2657 7244 2663 7246
rect 2671 7244 2686 7260
rect 2752 7254 2771 7257
rect 2393 7232 2491 7234
rect 2518 7232 2686 7244
rect 2701 7234 2717 7248
rect 2752 7235 2774 7254
rect 2784 7248 2800 7249
rect 2783 7246 2800 7248
rect 2784 7241 2800 7246
rect 2774 7234 2780 7235
rect 2783 7234 2812 7241
rect 2701 7233 2812 7234
rect 2701 7232 2818 7233
rect 2377 7224 2428 7232
rect 2475 7224 2509 7232
rect 2377 7212 2402 7224
rect 2409 7212 2428 7224
rect 2482 7222 2509 7224
rect 2518 7222 2739 7232
rect 2774 7229 2780 7232
rect 2482 7218 2739 7222
rect 2377 7204 2428 7212
rect 2475 7204 2739 7218
rect 2783 7224 2818 7232
rect 2329 7156 2348 7190
rect 2393 7196 2422 7204
rect 2393 7190 2410 7196
rect 2393 7188 2427 7190
rect 2475 7188 2491 7204
rect 2492 7194 2700 7204
rect 2701 7194 2717 7204
rect 2765 7200 2780 7215
rect 2783 7212 2784 7224
rect 2791 7212 2818 7224
rect 2783 7204 2818 7212
rect 2783 7203 2812 7204
rect 2503 7190 2717 7194
rect 2518 7188 2717 7190
rect 2752 7190 2765 7200
rect 2783 7190 2800 7203
rect 2752 7188 2800 7190
rect 2394 7184 2427 7188
rect 2390 7182 2427 7184
rect 2390 7181 2457 7182
rect 2390 7176 2421 7181
rect 2427 7176 2457 7181
rect 2390 7172 2457 7176
rect 2363 7169 2457 7172
rect 2363 7162 2412 7169
rect 2363 7156 2393 7162
rect 2412 7157 2417 7162
rect 2329 7140 2409 7156
rect 2421 7148 2457 7169
rect 2518 7164 2707 7188
rect 2752 7187 2799 7188
rect 2765 7182 2799 7187
rect 2533 7161 2707 7164
rect 2526 7158 2707 7161
rect 2735 7181 2799 7182
rect 2329 7138 2348 7140
rect 2363 7138 2397 7140
rect 2329 7122 2409 7138
rect 2329 7116 2348 7122
rect 2045 7090 2148 7100
rect 1999 7088 2148 7090
rect 2169 7088 2204 7100
rect 1838 7086 2000 7088
rect 1850 7066 1869 7086
rect 1884 7084 1914 7086
rect 1733 7058 1774 7066
rect 1856 7062 1869 7066
rect 1921 7070 2000 7086
rect 2032 7086 2204 7088
rect 2032 7070 2111 7086
rect 2118 7084 2148 7086
rect 1696 7048 1697 7058
rect 1712 7048 1725 7058
rect 1739 7048 1740 7058
rect 1755 7048 1768 7058
rect 1783 7048 1813 7062
rect 1856 7048 1899 7062
rect 1921 7058 2111 7070
rect 2176 7066 2182 7086
rect 1906 7048 1936 7058
rect 1937 7048 2095 7058
rect 2099 7048 2129 7058
rect 2133 7048 2163 7062
rect 2191 7048 2204 7086
rect 2276 7100 2305 7116
rect 2319 7100 2348 7116
rect 2363 7106 2393 7122
rect 2421 7100 2427 7148
rect 2430 7142 2449 7148
rect 2464 7142 2494 7150
rect 2430 7134 2494 7142
rect 2430 7118 2510 7134
rect 2526 7127 2588 7158
rect 2604 7127 2666 7158
rect 2735 7156 2784 7181
rect 2799 7156 2829 7172
rect 2698 7142 2728 7150
rect 2735 7148 2845 7156
rect 2698 7134 2743 7142
rect 2430 7116 2449 7118
rect 2464 7116 2510 7118
rect 2430 7100 2510 7116
rect 2537 7114 2572 7127
rect 2613 7124 2650 7127
rect 2613 7122 2655 7124
rect 2542 7111 2572 7114
rect 2551 7107 2558 7111
rect 2558 7106 2559 7107
rect 2517 7100 2527 7106
rect 2276 7092 2311 7100
rect 2276 7066 2277 7092
rect 2284 7066 2311 7092
rect 2219 7048 2249 7062
rect 2276 7058 2311 7066
rect 2313 7092 2354 7100
rect 2313 7066 2328 7092
rect 2335 7066 2354 7092
rect 2418 7088 2449 7100
rect 2464 7088 2567 7100
rect 2579 7090 2605 7116
rect 2620 7111 2650 7122
rect 2682 7118 2744 7134
rect 2682 7116 2728 7118
rect 2682 7100 2744 7116
rect 2756 7100 2762 7148
rect 2765 7140 2845 7148
rect 2765 7138 2784 7140
rect 2799 7138 2833 7140
rect 2765 7122 2845 7138
rect 2765 7100 2784 7122
rect 2799 7106 2829 7122
rect 2857 7116 2863 7190
rect 2866 7116 2885 7260
rect 2900 7116 2906 7260
rect 2915 7190 2928 7260
rect 2980 7256 3002 7260
rect 2973 7234 3002 7248
rect 3055 7234 3071 7248
rect 3109 7244 3115 7246
rect 3122 7244 3230 7260
rect 3237 7244 3243 7246
rect 3251 7244 3266 7260
rect 3332 7254 3351 7257
rect 2973 7232 3071 7234
rect 3098 7232 3266 7244
rect 3281 7234 3297 7248
rect 3332 7235 3354 7254
rect 3364 7248 3380 7249
rect 3363 7246 3380 7248
rect 3364 7241 3380 7246
rect 3354 7234 3360 7235
rect 3363 7234 3392 7241
rect 3281 7233 3392 7234
rect 3281 7232 3398 7233
rect 2957 7224 3008 7232
rect 3055 7224 3089 7232
rect 2957 7212 2982 7224
rect 2989 7212 3008 7224
rect 3062 7222 3089 7224
rect 3098 7222 3319 7232
rect 3354 7229 3360 7232
rect 3062 7218 3319 7222
rect 2957 7204 3008 7212
rect 3055 7204 3319 7218
rect 3363 7224 3398 7232
rect 2909 7156 2928 7190
rect 2973 7196 3002 7204
rect 2973 7190 2990 7196
rect 2973 7188 3007 7190
rect 3055 7188 3071 7204
rect 3072 7194 3280 7204
rect 3281 7194 3297 7204
rect 3345 7200 3360 7215
rect 3363 7212 3364 7224
rect 3371 7212 3398 7224
rect 3363 7204 3398 7212
rect 3363 7203 3392 7204
rect 3083 7190 3297 7194
rect 3098 7188 3297 7190
rect 3332 7190 3345 7200
rect 3363 7190 3380 7203
rect 3332 7188 3380 7190
rect 2974 7184 3007 7188
rect 2970 7182 3007 7184
rect 2970 7181 3037 7182
rect 2970 7176 3001 7181
rect 3007 7176 3037 7181
rect 2970 7172 3037 7176
rect 2943 7169 3037 7172
rect 2943 7162 2992 7169
rect 2943 7156 2973 7162
rect 2992 7157 2997 7162
rect 2909 7140 2989 7156
rect 3001 7148 3037 7169
rect 3098 7164 3287 7188
rect 3332 7187 3379 7188
rect 3345 7182 3379 7187
rect 3113 7161 3287 7164
rect 3106 7158 3287 7161
rect 3315 7181 3379 7182
rect 2909 7138 2928 7140
rect 2943 7138 2977 7140
rect 2909 7122 2989 7138
rect 2909 7116 2928 7122
rect 2625 7090 2728 7100
rect 2579 7088 2728 7090
rect 2749 7088 2784 7100
rect 2418 7086 2580 7088
rect 2430 7066 2449 7086
rect 2464 7084 2494 7086
rect 2313 7058 2354 7066
rect 2436 7062 2449 7066
rect 2501 7070 2580 7086
rect 2612 7086 2784 7088
rect 2612 7070 2691 7086
rect 2698 7084 2728 7086
rect 2276 7048 2305 7058
rect 2319 7048 2348 7058
rect 2363 7048 2393 7062
rect 2436 7048 2479 7062
rect 2501 7058 2691 7070
rect 2756 7066 2762 7086
rect 2486 7048 2516 7058
rect 2517 7048 2675 7058
rect 2679 7048 2709 7058
rect 2713 7048 2743 7062
rect 2771 7048 2784 7086
rect 2856 7100 2885 7116
rect 2899 7100 2928 7116
rect 2943 7106 2973 7122
rect 3001 7100 3007 7148
rect 3010 7142 3029 7148
rect 3044 7142 3074 7150
rect 3010 7134 3074 7142
rect 3010 7118 3090 7134
rect 3106 7127 3168 7158
rect 3184 7127 3246 7158
rect 3315 7156 3364 7181
rect 3379 7156 3409 7172
rect 3278 7142 3308 7150
rect 3315 7148 3425 7156
rect 3278 7134 3323 7142
rect 3010 7116 3029 7118
rect 3044 7116 3090 7118
rect 3010 7100 3090 7116
rect 3117 7114 3152 7127
rect 3193 7124 3230 7127
rect 3193 7122 3235 7124
rect 3122 7111 3152 7114
rect 3131 7107 3138 7111
rect 3138 7106 3139 7107
rect 3097 7100 3107 7106
rect 2856 7092 2891 7100
rect 2856 7066 2857 7092
rect 2864 7066 2891 7092
rect 2799 7048 2829 7062
rect 2856 7058 2891 7066
rect 2893 7092 2934 7100
rect 2893 7066 2908 7092
rect 2915 7066 2934 7092
rect 2998 7088 3029 7100
rect 3044 7088 3147 7100
rect 3159 7090 3185 7116
rect 3200 7111 3230 7122
rect 3262 7118 3324 7134
rect 3262 7116 3308 7118
rect 3262 7100 3324 7116
rect 3336 7100 3342 7148
rect 3345 7140 3425 7148
rect 3345 7138 3364 7140
rect 3379 7138 3413 7140
rect 3345 7122 3425 7138
rect 3345 7100 3364 7122
rect 3379 7106 3409 7122
rect 3437 7116 3443 7190
rect 3446 7116 3465 7260
rect 3480 7116 3486 7260
rect 3495 7190 3508 7260
rect 3560 7256 3582 7260
rect 3553 7234 3582 7248
rect 3635 7234 3651 7248
rect 3689 7244 3695 7246
rect 3702 7244 3810 7260
rect 3817 7244 3823 7246
rect 3831 7244 3846 7260
rect 3912 7254 3931 7257
rect 3553 7232 3651 7234
rect 3678 7232 3846 7244
rect 3861 7234 3877 7248
rect 3912 7235 3934 7254
rect 3944 7248 3960 7249
rect 3943 7246 3960 7248
rect 3944 7241 3960 7246
rect 3934 7234 3940 7235
rect 3943 7234 3972 7241
rect 3861 7233 3972 7234
rect 3861 7232 3978 7233
rect 3537 7224 3588 7232
rect 3635 7224 3669 7232
rect 3537 7212 3562 7224
rect 3569 7212 3588 7224
rect 3642 7222 3669 7224
rect 3678 7222 3899 7232
rect 3934 7229 3940 7232
rect 3642 7218 3899 7222
rect 3537 7204 3588 7212
rect 3635 7204 3899 7218
rect 3943 7224 3978 7232
rect 3489 7156 3508 7190
rect 3553 7196 3582 7204
rect 3553 7190 3570 7196
rect 3553 7188 3587 7190
rect 3635 7188 3651 7204
rect 3652 7194 3860 7204
rect 3861 7194 3877 7204
rect 3925 7200 3940 7215
rect 3943 7212 3944 7224
rect 3951 7212 3978 7224
rect 3943 7204 3978 7212
rect 3943 7203 3972 7204
rect 3663 7190 3877 7194
rect 3678 7188 3877 7190
rect 3912 7190 3925 7200
rect 3943 7190 3960 7203
rect 3912 7188 3960 7190
rect 3554 7184 3587 7188
rect 3550 7182 3587 7184
rect 3550 7181 3617 7182
rect 3550 7176 3581 7181
rect 3587 7176 3617 7181
rect 3550 7172 3617 7176
rect 3523 7169 3617 7172
rect 3523 7162 3572 7169
rect 3523 7156 3553 7162
rect 3572 7157 3577 7162
rect 3489 7140 3569 7156
rect 3581 7148 3617 7169
rect 3678 7164 3867 7188
rect 3912 7187 3959 7188
rect 3925 7182 3959 7187
rect 3693 7161 3867 7164
rect 3686 7158 3867 7161
rect 3895 7181 3959 7182
rect 3489 7138 3508 7140
rect 3523 7138 3557 7140
rect 3489 7122 3569 7138
rect 3489 7116 3508 7122
rect 3205 7090 3308 7100
rect 3159 7088 3308 7090
rect 3329 7088 3364 7100
rect 2998 7086 3160 7088
rect 3010 7066 3029 7086
rect 3044 7084 3074 7086
rect 2893 7058 2934 7066
rect 3016 7062 3029 7066
rect 3081 7070 3160 7086
rect 3192 7086 3364 7088
rect 3192 7070 3271 7086
rect 3278 7084 3308 7086
rect 2856 7048 2885 7058
rect 2899 7048 2928 7058
rect 2943 7048 2973 7062
rect 3016 7048 3059 7062
rect 3081 7058 3271 7070
rect 3336 7066 3342 7086
rect 3066 7048 3096 7058
rect 3097 7048 3255 7058
rect 3259 7048 3289 7058
rect 3293 7048 3323 7062
rect 3351 7048 3364 7086
rect 3436 7100 3465 7116
rect 3479 7100 3508 7116
rect 3523 7106 3553 7122
rect 3581 7100 3587 7148
rect 3590 7142 3609 7148
rect 3624 7142 3654 7150
rect 3590 7134 3654 7142
rect 3590 7118 3670 7134
rect 3686 7127 3748 7158
rect 3764 7127 3826 7158
rect 3895 7156 3944 7181
rect 3959 7156 3989 7172
rect 3858 7142 3888 7150
rect 3895 7148 4005 7156
rect 3858 7134 3903 7142
rect 3590 7116 3609 7118
rect 3624 7116 3670 7118
rect 3590 7100 3670 7116
rect 3697 7114 3732 7127
rect 3773 7124 3810 7127
rect 3773 7122 3815 7124
rect 3702 7111 3732 7114
rect 3711 7107 3718 7111
rect 3718 7106 3719 7107
rect 3677 7100 3687 7106
rect 3436 7092 3471 7100
rect 3436 7066 3437 7092
rect 3444 7066 3471 7092
rect 3379 7048 3409 7062
rect 3436 7058 3471 7066
rect 3473 7092 3514 7100
rect 3473 7066 3488 7092
rect 3495 7066 3514 7092
rect 3578 7088 3609 7100
rect 3624 7088 3727 7100
rect 3739 7090 3765 7116
rect 3780 7111 3810 7122
rect 3842 7118 3904 7134
rect 3842 7116 3888 7118
rect 3842 7100 3904 7116
rect 3916 7100 3922 7148
rect 3925 7140 4005 7148
rect 3925 7138 3944 7140
rect 3959 7138 3993 7140
rect 3925 7122 4005 7138
rect 3925 7100 3944 7122
rect 3959 7106 3989 7122
rect 4017 7116 4023 7190
rect 4026 7116 4045 7260
rect 4060 7116 4066 7260
rect 4075 7190 4088 7260
rect 4140 7256 4162 7260
rect 4133 7234 4162 7248
rect 4215 7234 4231 7248
rect 4269 7244 4275 7246
rect 4282 7244 4390 7260
rect 4397 7244 4403 7246
rect 4411 7244 4426 7260
rect 4492 7254 4511 7257
rect 4133 7232 4231 7234
rect 4258 7232 4426 7244
rect 4441 7234 4457 7248
rect 4492 7235 4514 7254
rect 4524 7248 4540 7249
rect 4523 7246 4540 7248
rect 4524 7241 4540 7246
rect 4514 7234 4520 7235
rect 4523 7234 4552 7241
rect 4441 7233 4552 7234
rect 4441 7232 4558 7233
rect 4117 7224 4168 7232
rect 4215 7224 4249 7232
rect 4117 7212 4142 7224
rect 4149 7212 4168 7224
rect 4222 7222 4249 7224
rect 4258 7222 4479 7232
rect 4514 7229 4520 7232
rect 4222 7218 4479 7222
rect 4117 7204 4168 7212
rect 4215 7204 4479 7218
rect 4523 7224 4558 7232
rect 4069 7156 4088 7190
rect 4133 7196 4162 7204
rect 4133 7190 4150 7196
rect 4133 7188 4167 7190
rect 4215 7188 4231 7204
rect 4232 7194 4440 7204
rect 4441 7194 4457 7204
rect 4505 7200 4520 7215
rect 4523 7212 4524 7224
rect 4531 7212 4558 7224
rect 4523 7204 4558 7212
rect 4523 7203 4552 7204
rect 4243 7190 4457 7194
rect 4258 7188 4457 7190
rect 4492 7190 4505 7200
rect 4523 7190 4540 7203
rect 4492 7188 4540 7190
rect 4134 7184 4167 7188
rect 4130 7182 4167 7184
rect 4130 7181 4197 7182
rect 4130 7176 4161 7181
rect 4167 7176 4197 7181
rect 4130 7172 4197 7176
rect 4103 7169 4197 7172
rect 4103 7162 4152 7169
rect 4103 7156 4133 7162
rect 4152 7157 4157 7162
rect 4069 7140 4149 7156
rect 4161 7148 4197 7169
rect 4258 7164 4447 7188
rect 4492 7187 4539 7188
rect 4505 7182 4539 7187
rect 4273 7161 4447 7164
rect 4266 7158 4447 7161
rect 4475 7181 4539 7182
rect 4069 7138 4088 7140
rect 4103 7138 4137 7140
rect 4069 7122 4149 7138
rect 4069 7116 4088 7122
rect 3785 7090 3888 7100
rect 3739 7088 3888 7090
rect 3909 7088 3944 7100
rect 3578 7086 3740 7088
rect 3590 7066 3609 7086
rect 3624 7084 3654 7086
rect 3473 7058 3514 7066
rect 3596 7062 3609 7066
rect 3661 7070 3740 7086
rect 3772 7086 3944 7088
rect 3772 7070 3851 7086
rect 3858 7084 3888 7086
rect 3436 7048 3465 7058
rect 3479 7048 3508 7058
rect 3523 7048 3553 7062
rect 3596 7048 3639 7062
rect 3661 7058 3851 7070
rect 3916 7066 3922 7086
rect 3646 7048 3676 7058
rect 3677 7048 3835 7058
rect 3839 7048 3869 7058
rect 3873 7048 3903 7062
rect 3931 7048 3944 7086
rect 4016 7100 4045 7116
rect 4059 7100 4088 7116
rect 4103 7106 4133 7122
rect 4161 7100 4167 7148
rect 4170 7142 4189 7148
rect 4204 7142 4234 7150
rect 4170 7134 4234 7142
rect 4170 7118 4250 7134
rect 4266 7127 4328 7158
rect 4344 7127 4406 7158
rect 4475 7156 4524 7181
rect 4539 7156 4569 7172
rect 4438 7142 4468 7150
rect 4475 7148 4585 7156
rect 4438 7134 4483 7142
rect 4170 7116 4189 7118
rect 4204 7116 4250 7118
rect 4170 7100 4250 7116
rect 4277 7114 4312 7127
rect 4353 7124 4390 7127
rect 4353 7122 4395 7124
rect 4282 7111 4312 7114
rect 4291 7107 4298 7111
rect 4298 7106 4299 7107
rect 4257 7100 4267 7106
rect 4016 7092 4051 7100
rect 4016 7066 4017 7092
rect 4024 7066 4051 7092
rect 3959 7048 3989 7062
rect 4016 7058 4051 7066
rect 4053 7092 4094 7100
rect 4053 7066 4068 7092
rect 4075 7066 4094 7092
rect 4158 7088 4189 7100
rect 4204 7088 4307 7100
rect 4319 7090 4345 7116
rect 4360 7111 4390 7122
rect 4422 7118 4484 7134
rect 4422 7116 4468 7118
rect 4422 7100 4484 7116
rect 4496 7100 4502 7148
rect 4505 7140 4585 7148
rect 4505 7138 4524 7140
rect 4539 7138 4573 7140
rect 4505 7122 4585 7138
rect 4505 7100 4524 7122
rect 4539 7106 4569 7122
rect 4597 7116 4603 7190
rect 4606 7116 4625 7260
rect 4640 7116 4646 7260
rect 4655 7190 4668 7260
rect 4720 7256 4742 7260
rect 4713 7234 4742 7248
rect 4795 7234 4811 7248
rect 4849 7244 4855 7246
rect 4862 7244 4970 7260
rect 4977 7244 4983 7246
rect 4991 7244 5006 7260
rect 5072 7254 5091 7257
rect 4713 7232 4811 7234
rect 4838 7232 5006 7244
rect 5021 7234 5037 7248
rect 5072 7235 5094 7254
rect 5104 7248 5120 7249
rect 5103 7246 5120 7248
rect 5104 7241 5120 7246
rect 5094 7234 5100 7235
rect 5103 7234 5132 7241
rect 5021 7233 5132 7234
rect 5021 7232 5138 7233
rect 4697 7224 4748 7232
rect 4795 7224 4829 7232
rect 4697 7212 4722 7224
rect 4729 7212 4748 7224
rect 4802 7222 4829 7224
rect 4838 7222 5059 7232
rect 5094 7229 5100 7232
rect 4802 7218 5059 7222
rect 4697 7204 4748 7212
rect 4795 7204 5059 7218
rect 5103 7224 5138 7232
rect 4649 7156 4668 7190
rect 4713 7196 4742 7204
rect 4713 7190 4730 7196
rect 4713 7188 4747 7190
rect 4795 7188 4811 7204
rect 4812 7194 5020 7204
rect 5021 7194 5037 7204
rect 5085 7200 5100 7215
rect 5103 7212 5104 7224
rect 5111 7212 5138 7224
rect 5103 7204 5138 7212
rect 5103 7203 5132 7204
rect 4823 7190 5037 7194
rect 4838 7188 5037 7190
rect 5072 7190 5085 7200
rect 5103 7190 5120 7203
rect 5072 7188 5120 7190
rect 4714 7184 4747 7188
rect 4710 7182 4747 7184
rect 4710 7181 4777 7182
rect 4710 7176 4741 7181
rect 4747 7176 4777 7181
rect 4710 7172 4777 7176
rect 4683 7169 4777 7172
rect 4683 7162 4732 7169
rect 4683 7156 4713 7162
rect 4732 7157 4737 7162
rect 4649 7140 4729 7156
rect 4741 7148 4777 7169
rect 4838 7164 5027 7188
rect 5072 7187 5119 7188
rect 5085 7182 5119 7187
rect 4853 7161 5027 7164
rect 4846 7158 5027 7161
rect 5055 7181 5119 7182
rect 4649 7138 4668 7140
rect 4683 7138 4717 7140
rect 4649 7122 4729 7138
rect 4649 7116 4668 7122
rect 4365 7090 4468 7100
rect 4319 7088 4468 7090
rect 4489 7088 4524 7100
rect 4158 7086 4320 7088
rect 4170 7066 4189 7086
rect 4204 7084 4234 7086
rect 4053 7058 4094 7066
rect 4176 7062 4189 7066
rect 4241 7070 4320 7086
rect 4352 7086 4524 7088
rect 4352 7070 4431 7086
rect 4438 7084 4468 7086
rect 4016 7048 4045 7058
rect 4059 7048 4088 7058
rect 4103 7048 4133 7062
rect 4176 7048 4219 7062
rect 4241 7058 4431 7070
rect 4496 7066 4502 7086
rect 4226 7048 4256 7058
rect 4257 7048 4415 7058
rect 4419 7048 4449 7058
rect 4453 7048 4483 7062
rect 4511 7048 4524 7086
rect 4596 7100 4625 7116
rect 4639 7100 4668 7116
rect 4683 7106 4713 7122
rect 4741 7100 4747 7148
rect 4750 7142 4769 7148
rect 4784 7142 4814 7150
rect 4750 7134 4814 7142
rect 4750 7118 4830 7134
rect 4846 7127 4908 7158
rect 4924 7127 4986 7158
rect 5055 7156 5104 7181
rect 5119 7156 5149 7172
rect 5018 7142 5048 7150
rect 5055 7148 5165 7156
rect 5018 7134 5063 7142
rect 4750 7116 4769 7118
rect 4784 7116 4830 7118
rect 4750 7100 4830 7116
rect 4857 7114 4892 7127
rect 4933 7124 4970 7127
rect 4933 7122 4975 7124
rect 4862 7111 4892 7114
rect 4871 7107 4878 7111
rect 4878 7106 4879 7107
rect 4837 7100 4847 7106
rect 4596 7092 4631 7100
rect 4596 7066 4597 7092
rect 4604 7066 4631 7092
rect 4539 7048 4569 7062
rect 4596 7058 4631 7066
rect 4633 7092 4674 7100
rect 4633 7066 4648 7092
rect 4655 7066 4674 7092
rect 4738 7088 4769 7100
rect 4784 7088 4887 7100
rect 4899 7090 4925 7116
rect 4940 7111 4970 7122
rect 5002 7118 5064 7134
rect 5002 7116 5048 7118
rect 5002 7100 5064 7116
rect 5076 7100 5082 7148
rect 5085 7140 5165 7148
rect 5085 7138 5104 7140
rect 5119 7138 5153 7140
rect 5085 7122 5165 7138
rect 5085 7100 5104 7122
rect 5119 7106 5149 7122
rect 5177 7116 5183 7190
rect 5186 7116 5205 7260
rect 5220 7116 5226 7260
rect 5235 7190 5248 7260
rect 5300 7256 5322 7260
rect 5293 7234 5322 7248
rect 5375 7234 5391 7248
rect 5429 7244 5435 7246
rect 5442 7244 5550 7260
rect 5557 7244 5563 7246
rect 5571 7244 5586 7260
rect 5652 7254 5671 7257
rect 5293 7232 5391 7234
rect 5418 7232 5586 7244
rect 5601 7234 5617 7248
rect 5652 7235 5674 7254
rect 5684 7248 5700 7249
rect 5683 7246 5700 7248
rect 5684 7241 5700 7246
rect 5674 7234 5680 7235
rect 5683 7234 5712 7241
rect 5601 7233 5712 7234
rect 5601 7232 5718 7233
rect 5277 7224 5328 7232
rect 5375 7224 5409 7232
rect 5277 7212 5302 7224
rect 5309 7212 5328 7224
rect 5382 7222 5409 7224
rect 5418 7222 5639 7232
rect 5674 7229 5680 7232
rect 5382 7218 5639 7222
rect 5277 7204 5328 7212
rect 5375 7204 5639 7218
rect 5683 7224 5718 7232
rect 5229 7156 5248 7190
rect 5293 7196 5322 7204
rect 5293 7190 5310 7196
rect 5293 7188 5327 7190
rect 5375 7188 5391 7204
rect 5392 7194 5600 7204
rect 5601 7194 5617 7204
rect 5665 7200 5680 7215
rect 5683 7212 5684 7224
rect 5691 7212 5718 7224
rect 5683 7204 5718 7212
rect 5683 7203 5712 7204
rect 5403 7190 5617 7194
rect 5418 7188 5617 7190
rect 5652 7190 5665 7200
rect 5683 7190 5700 7203
rect 5652 7188 5700 7190
rect 5294 7184 5327 7188
rect 5290 7182 5327 7184
rect 5290 7181 5357 7182
rect 5290 7176 5321 7181
rect 5327 7176 5357 7181
rect 5290 7172 5357 7176
rect 5263 7169 5357 7172
rect 5263 7162 5312 7169
rect 5263 7156 5293 7162
rect 5312 7157 5317 7162
rect 5229 7140 5309 7156
rect 5321 7148 5357 7169
rect 5418 7164 5607 7188
rect 5652 7187 5699 7188
rect 5665 7182 5699 7187
rect 5433 7161 5607 7164
rect 5426 7158 5607 7161
rect 5635 7181 5699 7182
rect 5229 7138 5248 7140
rect 5263 7138 5297 7140
rect 5229 7122 5309 7138
rect 5229 7116 5248 7122
rect 4945 7090 5048 7100
rect 4899 7088 5048 7090
rect 5069 7088 5104 7100
rect 4738 7086 4900 7088
rect 4750 7066 4769 7086
rect 4784 7084 4814 7086
rect 4633 7058 4674 7066
rect 4756 7062 4769 7066
rect 4821 7070 4900 7086
rect 4932 7086 5104 7088
rect 4932 7070 5011 7086
rect 5018 7084 5048 7086
rect 4596 7048 4625 7058
rect 4639 7048 4668 7058
rect 4683 7048 4713 7062
rect 4756 7048 4799 7062
rect 4821 7058 5011 7070
rect 5076 7066 5082 7086
rect 4806 7048 4836 7058
rect 4837 7048 4995 7058
rect 4999 7048 5029 7058
rect 5033 7048 5063 7062
rect 5091 7048 5104 7086
rect 5176 7100 5205 7116
rect 5219 7100 5248 7116
rect 5263 7106 5293 7122
rect 5321 7100 5327 7148
rect 5330 7142 5349 7148
rect 5364 7142 5394 7150
rect 5330 7134 5394 7142
rect 5330 7118 5410 7134
rect 5426 7127 5488 7158
rect 5504 7127 5566 7158
rect 5635 7156 5684 7181
rect 5699 7156 5729 7172
rect 5598 7142 5628 7150
rect 5635 7148 5745 7156
rect 5598 7134 5643 7142
rect 5330 7116 5349 7118
rect 5364 7116 5410 7118
rect 5330 7100 5410 7116
rect 5437 7114 5472 7127
rect 5513 7124 5550 7127
rect 5513 7122 5555 7124
rect 5442 7111 5472 7114
rect 5451 7107 5458 7111
rect 5458 7106 5459 7107
rect 5417 7100 5427 7106
rect 5176 7092 5211 7100
rect 5176 7066 5177 7092
rect 5184 7066 5211 7092
rect 5119 7048 5149 7062
rect 5176 7058 5211 7066
rect 5213 7092 5254 7100
rect 5213 7066 5228 7092
rect 5235 7066 5254 7092
rect 5318 7088 5349 7100
rect 5364 7088 5467 7100
rect 5479 7090 5505 7116
rect 5520 7111 5550 7122
rect 5582 7118 5644 7134
rect 5582 7116 5628 7118
rect 5582 7100 5644 7116
rect 5656 7100 5662 7148
rect 5665 7140 5745 7148
rect 5665 7138 5684 7140
rect 5699 7138 5733 7140
rect 5665 7122 5745 7138
rect 5665 7100 5684 7122
rect 5699 7106 5729 7122
rect 5757 7116 5763 7190
rect 5766 7116 5785 7260
rect 5800 7116 5806 7260
rect 5815 7190 5828 7260
rect 5880 7256 5902 7260
rect 5873 7234 5902 7248
rect 5955 7234 5971 7248
rect 6009 7244 6015 7246
rect 6022 7244 6130 7260
rect 6137 7244 6143 7246
rect 6151 7244 6166 7260
rect 6232 7254 6251 7257
rect 5873 7232 5971 7234
rect 5998 7232 6166 7244
rect 6181 7234 6197 7248
rect 6232 7235 6254 7254
rect 6264 7248 6280 7249
rect 6263 7246 6280 7248
rect 6264 7241 6280 7246
rect 6254 7234 6260 7235
rect 6263 7234 6292 7241
rect 6181 7233 6292 7234
rect 6181 7232 6298 7233
rect 5857 7224 5908 7232
rect 5955 7224 5989 7232
rect 5857 7212 5882 7224
rect 5889 7212 5908 7224
rect 5962 7222 5989 7224
rect 5998 7222 6219 7232
rect 6254 7229 6260 7232
rect 5962 7218 6219 7222
rect 5857 7204 5908 7212
rect 5955 7204 6219 7218
rect 6263 7224 6298 7232
rect 5809 7156 5828 7190
rect 5873 7196 5902 7204
rect 5873 7190 5890 7196
rect 5873 7188 5907 7190
rect 5955 7188 5971 7204
rect 5972 7194 6180 7204
rect 6181 7194 6197 7204
rect 6245 7200 6260 7215
rect 6263 7212 6264 7224
rect 6271 7212 6298 7224
rect 6263 7204 6298 7212
rect 6263 7203 6292 7204
rect 5983 7190 6197 7194
rect 5998 7188 6197 7190
rect 6232 7190 6245 7200
rect 6263 7190 6280 7203
rect 6232 7188 6280 7190
rect 5874 7184 5907 7188
rect 5870 7182 5907 7184
rect 5870 7181 5937 7182
rect 5870 7176 5901 7181
rect 5907 7176 5937 7181
rect 5870 7172 5937 7176
rect 5843 7169 5937 7172
rect 5843 7162 5892 7169
rect 5843 7156 5873 7162
rect 5892 7157 5897 7162
rect 5809 7140 5889 7156
rect 5901 7148 5937 7169
rect 5998 7164 6187 7188
rect 6232 7187 6279 7188
rect 6245 7182 6279 7187
rect 6013 7161 6187 7164
rect 6006 7158 6187 7161
rect 6215 7181 6279 7182
rect 5809 7138 5828 7140
rect 5843 7138 5877 7140
rect 5809 7122 5889 7138
rect 5809 7116 5828 7122
rect 5525 7090 5628 7100
rect 5479 7088 5628 7090
rect 5649 7088 5684 7100
rect 5318 7086 5480 7088
rect 5330 7066 5349 7086
rect 5364 7084 5394 7086
rect 5213 7058 5254 7066
rect 5336 7062 5349 7066
rect 5401 7070 5480 7086
rect 5512 7086 5684 7088
rect 5512 7070 5591 7086
rect 5598 7084 5628 7086
rect 5176 7048 5205 7058
rect 5219 7048 5248 7058
rect 5263 7048 5293 7062
rect 5336 7048 5379 7062
rect 5401 7058 5591 7070
rect 5656 7066 5662 7086
rect 5386 7048 5416 7058
rect 5417 7048 5575 7058
rect 5579 7048 5609 7058
rect 5613 7048 5643 7062
rect 5671 7048 5684 7086
rect 5756 7100 5785 7116
rect 5799 7100 5828 7116
rect 5843 7106 5873 7122
rect 5901 7100 5907 7148
rect 5910 7142 5929 7148
rect 5944 7142 5974 7150
rect 5910 7134 5974 7142
rect 5910 7118 5990 7134
rect 6006 7127 6068 7158
rect 6084 7127 6146 7158
rect 6215 7156 6264 7181
rect 6279 7156 6309 7172
rect 6178 7142 6208 7150
rect 6215 7148 6325 7156
rect 6178 7134 6223 7142
rect 5910 7116 5929 7118
rect 5944 7116 5990 7118
rect 5910 7100 5990 7116
rect 6017 7114 6052 7127
rect 6093 7124 6130 7127
rect 6093 7122 6135 7124
rect 6022 7111 6052 7114
rect 6031 7107 6038 7111
rect 6038 7106 6039 7107
rect 5997 7100 6007 7106
rect 5756 7092 5791 7100
rect 5756 7066 5757 7092
rect 5764 7066 5791 7092
rect 5699 7048 5729 7062
rect 5756 7058 5791 7066
rect 5793 7092 5834 7100
rect 5793 7066 5808 7092
rect 5815 7066 5834 7092
rect 5898 7088 5929 7100
rect 5944 7088 6047 7100
rect 6059 7090 6085 7116
rect 6100 7111 6130 7122
rect 6162 7118 6224 7134
rect 6162 7116 6208 7118
rect 6162 7100 6224 7116
rect 6236 7100 6242 7148
rect 6245 7140 6325 7148
rect 6245 7138 6264 7140
rect 6279 7138 6313 7140
rect 6245 7122 6325 7138
rect 6245 7100 6264 7122
rect 6279 7106 6309 7122
rect 6337 7116 6343 7190
rect 6346 7116 6365 7260
rect 6380 7116 6386 7260
rect 6395 7190 6408 7260
rect 6460 7256 6482 7260
rect 6453 7234 6482 7248
rect 6535 7234 6551 7248
rect 6589 7244 6595 7246
rect 6602 7244 6710 7260
rect 6717 7244 6723 7246
rect 6731 7244 6746 7260
rect 6812 7254 6831 7257
rect 6453 7232 6551 7234
rect 6578 7232 6746 7244
rect 6761 7234 6777 7248
rect 6812 7235 6834 7254
rect 6844 7248 6860 7249
rect 6843 7246 6860 7248
rect 6844 7241 6860 7246
rect 6834 7234 6840 7235
rect 6843 7234 6872 7241
rect 6761 7233 6872 7234
rect 6761 7232 6878 7233
rect 6437 7224 6488 7232
rect 6535 7224 6569 7232
rect 6437 7212 6462 7224
rect 6469 7212 6488 7224
rect 6542 7222 6569 7224
rect 6578 7222 6799 7232
rect 6834 7229 6840 7232
rect 6542 7218 6799 7222
rect 6437 7204 6488 7212
rect 6535 7204 6799 7218
rect 6843 7224 6878 7232
rect 6389 7156 6408 7190
rect 6453 7196 6482 7204
rect 6453 7190 6470 7196
rect 6453 7188 6487 7190
rect 6535 7188 6551 7204
rect 6552 7194 6760 7204
rect 6761 7194 6777 7204
rect 6825 7200 6840 7215
rect 6843 7212 6844 7224
rect 6851 7212 6878 7224
rect 6843 7204 6878 7212
rect 6843 7203 6872 7204
rect 6563 7190 6777 7194
rect 6578 7188 6777 7190
rect 6812 7190 6825 7200
rect 6843 7190 6860 7203
rect 6812 7188 6860 7190
rect 6454 7184 6487 7188
rect 6450 7182 6487 7184
rect 6450 7181 6517 7182
rect 6450 7176 6481 7181
rect 6487 7176 6517 7181
rect 6450 7172 6517 7176
rect 6423 7169 6517 7172
rect 6423 7162 6472 7169
rect 6423 7156 6453 7162
rect 6472 7157 6477 7162
rect 6389 7140 6469 7156
rect 6481 7148 6517 7169
rect 6578 7164 6767 7188
rect 6812 7187 6859 7188
rect 6825 7182 6859 7187
rect 6593 7161 6767 7164
rect 6586 7158 6767 7161
rect 6795 7181 6859 7182
rect 6389 7138 6408 7140
rect 6423 7138 6457 7140
rect 6389 7122 6469 7138
rect 6389 7116 6408 7122
rect 6105 7090 6208 7100
rect 6059 7088 6208 7090
rect 6229 7088 6264 7100
rect 5898 7086 6060 7088
rect 5910 7066 5929 7086
rect 5944 7084 5974 7086
rect 5793 7058 5834 7066
rect 5916 7062 5929 7066
rect 5981 7070 6060 7086
rect 6092 7086 6264 7088
rect 6092 7070 6171 7086
rect 6178 7084 6208 7086
rect 5756 7048 5785 7058
rect 5799 7048 5828 7058
rect 5843 7048 5873 7062
rect 5916 7048 5959 7062
rect 5981 7058 6171 7070
rect 6236 7066 6242 7086
rect 5966 7048 5996 7058
rect 5997 7048 6155 7058
rect 6159 7048 6189 7058
rect 6193 7048 6223 7062
rect 6251 7048 6264 7086
rect 6336 7100 6365 7116
rect 6379 7100 6408 7116
rect 6423 7106 6453 7122
rect 6481 7100 6487 7148
rect 6490 7142 6509 7148
rect 6524 7142 6554 7150
rect 6490 7134 6554 7142
rect 6490 7118 6570 7134
rect 6586 7127 6648 7158
rect 6664 7127 6726 7158
rect 6795 7156 6844 7181
rect 6859 7156 6889 7172
rect 6758 7142 6788 7150
rect 6795 7148 6905 7156
rect 6758 7134 6803 7142
rect 6490 7116 6509 7118
rect 6524 7116 6570 7118
rect 6490 7100 6570 7116
rect 6597 7114 6632 7127
rect 6673 7124 6710 7127
rect 6673 7122 6715 7124
rect 6602 7111 6632 7114
rect 6611 7107 6618 7111
rect 6618 7106 6619 7107
rect 6577 7100 6587 7106
rect 6336 7092 6371 7100
rect 6336 7066 6337 7092
rect 6344 7066 6371 7092
rect 6279 7048 6309 7062
rect 6336 7058 6371 7066
rect 6373 7092 6414 7100
rect 6373 7066 6388 7092
rect 6395 7066 6414 7092
rect 6478 7088 6509 7100
rect 6524 7088 6627 7100
rect 6639 7090 6665 7116
rect 6680 7111 6710 7122
rect 6742 7118 6804 7134
rect 6742 7116 6788 7118
rect 6742 7100 6804 7116
rect 6816 7100 6822 7148
rect 6825 7140 6905 7148
rect 6825 7138 6844 7140
rect 6859 7138 6893 7140
rect 6825 7122 6905 7138
rect 6825 7100 6844 7122
rect 6859 7106 6889 7122
rect 6917 7116 6923 7190
rect 6926 7116 6945 7260
rect 6960 7116 6966 7260
rect 6975 7190 6988 7260
rect 7040 7256 7062 7260
rect 7033 7234 7062 7248
rect 7115 7234 7131 7248
rect 7169 7244 7175 7246
rect 7182 7244 7290 7260
rect 7297 7244 7303 7246
rect 7311 7244 7326 7260
rect 7392 7254 7411 7257
rect 7033 7232 7131 7234
rect 7158 7232 7326 7244
rect 7341 7234 7357 7248
rect 7392 7235 7414 7254
rect 7424 7248 7440 7249
rect 7423 7246 7440 7248
rect 7424 7241 7440 7246
rect 7414 7234 7420 7235
rect 7423 7234 7452 7241
rect 7341 7233 7452 7234
rect 7341 7232 7458 7233
rect 7017 7224 7068 7232
rect 7115 7224 7149 7232
rect 7017 7212 7042 7224
rect 7049 7212 7068 7224
rect 7122 7222 7149 7224
rect 7158 7222 7379 7232
rect 7414 7229 7420 7232
rect 7122 7218 7379 7222
rect 7017 7204 7068 7212
rect 7115 7204 7379 7218
rect 7423 7224 7458 7232
rect 6969 7156 6988 7190
rect 7033 7196 7062 7204
rect 7033 7190 7050 7196
rect 7033 7188 7067 7190
rect 7115 7188 7131 7204
rect 7132 7194 7340 7204
rect 7341 7194 7357 7204
rect 7405 7200 7420 7215
rect 7423 7212 7424 7224
rect 7431 7212 7458 7224
rect 7423 7204 7458 7212
rect 7423 7203 7452 7204
rect 7143 7190 7357 7194
rect 7158 7188 7357 7190
rect 7392 7190 7405 7200
rect 7423 7190 7440 7203
rect 7392 7188 7440 7190
rect 7034 7184 7067 7188
rect 7030 7182 7067 7184
rect 7030 7181 7097 7182
rect 7030 7176 7061 7181
rect 7067 7176 7097 7181
rect 7030 7172 7097 7176
rect 7003 7169 7097 7172
rect 7003 7162 7052 7169
rect 7003 7156 7033 7162
rect 7052 7157 7057 7162
rect 6969 7140 7049 7156
rect 7061 7148 7097 7169
rect 7158 7164 7347 7188
rect 7392 7187 7439 7188
rect 7405 7182 7439 7187
rect 7173 7161 7347 7164
rect 7166 7158 7347 7161
rect 7375 7181 7439 7182
rect 6969 7138 6988 7140
rect 7003 7138 7037 7140
rect 6969 7122 7049 7138
rect 6969 7116 6988 7122
rect 6685 7090 6788 7100
rect 6639 7088 6788 7090
rect 6809 7088 6844 7100
rect 6478 7086 6640 7088
rect 6490 7066 6509 7086
rect 6524 7084 6554 7086
rect 6373 7058 6414 7066
rect 6496 7062 6509 7066
rect 6561 7070 6640 7086
rect 6672 7086 6844 7088
rect 6672 7070 6751 7086
rect 6758 7084 6788 7086
rect 6336 7048 6365 7058
rect 6379 7048 6408 7058
rect 6423 7048 6453 7062
rect 6496 7048 6539 7062
rect 6561 7058 6751 7070
rect 6816 7066 6822 7086
rect 6546 7048 6576 7058
rect 6577 7048 6735 7058
rect 6739 7048 6769 7058
rect 6773 7048 6803 7062
rect 6831 7048 6844 7086
rect 6916 7100 6945 7116
rect 6959 7100 6988 7116
rect 7003 7106 7033 7122
rect 7061 7100 7067 7148
rect 7070 7142 7089 7148
rect 7104 7142 7134 7150
rect 7070 7134 7134 7142
rect 7070 7118 7150 7134
rect 7166 7127 7228 7158
rect 7244 7127 7306 7158
rect 7375 7156 7424 7181
rect 7439 7156 7469 7172
rect 7338 7142 7368 7150
rect 7375 7148 7485 7156
rect 7338 7134 7383 7142
rect 7070 7116 7089 7118
rect 7104 7116 7150 7118
rect 7070 7100 7150 7116
rect 7177 7114 7212 7127
rect 7253 7124 7290 7127
rect 7253 7122 7295 7124
rect 7182 7111 7212 7114
rect 7191 7107 7198 7111
rect 7198 7106 7199 7107
rect 7157 7100 7167 7106
rect 6916 7092 6951 7100
rect 6916 7066 6917 7092
rect 6924 7066 6951 7092
rect 6859 7048 6889 7062
rect 6916 7058 6951 7066
rect 6953 7092 6994 7100
rect 6953 7066 6968 7092
rect 6975 7066 6994 7092
rect 7058 7088 7089 7100
rect 7104 7088 7207 7100
rect 7219 7090 7245 7116
rect 7260 7111 7290 7122
rect 7322 7118 7384 7134
rect 7322 7116 7368 7118
rect 7322 7100 7384 7116
rect 7396 7100 7402 7148
rect 7405 7140 7485 7148
rect 7405 7138 7424 7140
rect 7439 7138 7473 7140
rect 7405 7122 7485 7138
rect 7405 7100 7424 7122
rect 7439 7106 7469 7122
rect 7497 7116 7503 7190
rect 7506 7116 7525 7260
rect 7540 7116 7546 7260
rect 7555 7190 7568 7260
rect 7613 7238 7614 7248
rect 7629 7238 7642 7248
rect 7613 7234 7642 7238
rect 7647 7234 7677 7260
rect 7695 7246 7711 7248
rect 7783 7246 7836 7260
rect 7784 7244 7848 7246
rect 7891 7244 7906 7260
rect 7955 7257 7985 7260
rect 7955 7254 7991 7257
rect 7921 7246 7937 7248
rect 7695 7234 7710 7238
rect 7613 7232 7710 7234
rect 7738 7232 7906 7244
rect 7922 7234 7937 7238
rect 7955 7235 7994 7254
rect 8013 7248 8020 7249
rect 8019 7241 8020 7248
rect 8003 7238 8004 7241
rect 8019 7238 8032 7241
rect 7955 7234 7985 7235
rect 7994 7234 8000 7235
rect 8003 7234 8032 7238
rect 7922 7233 8032 7234
rect 7922 7232 8038 7233
rect 7597 7224 7648 7232
rect 7597 7212 7622 7224
rect 7629 7212 7648 7224
rect 7679 7224 7729 7232
rect 7679 7216 7695 7224
rect 7702 7222 7729 7224
rect 7738 7222 7959 7232
rect 7702 7212 7959 7222
rect 7988 7224 8038 7232
rect 7988 7215 8004 7224
rect 7597 7204 7648 7212
rect 7695 7204 7959 7212
rect 7985 7212 8004 7215
rect 8011 7212 8038 7224
rect 7985 7204 8038 7212
rect 7549 7156 7568 7190
rect 7613 7196 7614 7204
rect 7629 7196 7642 7204
rect 7613 7188 7629 7196
rect 7610 7181 7629 7184
rect 7610 7172 7632 7181
rect 7583 7162 7632 7172
rect 7583 7156 7613 7162
rect 7632 7157 7637 7162
rect 7549 7140 7629 7156
rect 7647 7148 7677 7204
rect 7712 7194 7920 7204
rect 7955 7200 8000 7204
rect 8003 7203 8004 7204
rect 8019 7203 8032 7204
rect 7738 7164 7927 7194
rect 7753 7161 7927 7164
rect 7746 7158 7927 7161
rect 7549 7138 7568 7140
rect 7583 7138 7617 7140
rect 7549 7122 7629 7138
rect 7656 7134 7669 7148
rect 7684 7134 7700 7150
rect 7746 7145 7757 7158
rect 7549 7116 7568 7122
rect 7265 7090 7368 7100
rect 7219 7088 7368 7090
rect 7389 7088 7424 7100
rect 7058 7086 7220 7088
rect 7070 7066 7089 7086
rect 7104 7084 7134 7086
rect 6953 7058 6994 7066
rect 7076 7062 7089 7066
rect 7141 7070 7220 7086
rect 7252 7086 7424 7088
rect 7252 7070 7331 7086
rect 7338 7084 7368 7086
rect 6916 7048 6945 7058
rect 6959 7048 6988 7058
rect 7003 7048 7033 7062
rect 7076 7048 7119 7062
rect 7141 7058 7331 7070
rect 7396 7066 7402 7086
rect 7126 7048 7156 7058
rect 7157 7048 7315 7058
rect 7319 7048 7349 7058
rect 7353 7048 7383 7062
rect 7411 7048 7424 7086
rect 7496 7100 7525 7116
rect 7539 7100 7568 7116
rect 7583 7100 7613 7122
rect 7656 7118 7718 7134
rect 7746 7127 7757 7143
rect 7762 7138 7772 7158
rect 7782 7138 7796 7158
rect 7799 7145 7808 7158
rect 7824 7145 7833 7158
rect 7762 7127 7796 7138
rect 7799 7127 7808 7143
rect 7824 7127 7833 7143
rect 7840 7138 7850 7158
rect 7860 7138 7874 7158
rect 7875 7145 7886 7158
rect 7840 7127 7874 7138
rect 7875 7127 7886 7143
rect 7932 7134 7948 7150
rect 7955 7148 7985 7200
rect 8019 7196 8020 7203
rect 8004 7188 8020 7196
rect 7991 7156 8004 7175
rect 8019 7156 8049 7172
rect 7991 7140 8065 7156
rect 7991 7138 8004 7140
rect 8019 7138 8053 7140
rect 7656 7116 7669 7118
rect 7684 7116 7718 7118
rect 7656 7100 7718 7116
rect 7762 7111 7778 7114
rect 7840 7111 7870 7122
rect 7918 7118 7964 7134
rect 7991 7122 8065 7138
rect 7918 7116 7952 7118
rect 7917 7100 7964 7116
rect 7991 7100 8004 7122
rect 8019 7100 8049 7122
rect 8076 7100 8077 7116
rect 8092 7100 8105 7260
rect 8135 7156 8148 7260
rect 8193 7238 8194 7248
rect 8209 7238 8222 7248
rect 8193 7234 8222 7238
rect 8227 7234 8257 7260
rect 8275 7246 8291 7248
rect 8363 7246 8416 7260
rect 8364 7244 8428 7246
rect 8471 7244 8486 7260
rect 8535 7257 8565 7260
rect 8535 7254 8571 7257
rect 8501 7246 8517 7248
rect 8275 7234 8290 7238
rect 8193 7232 8290 7234
rect 8318 7232 8486 7244
rect 8502 7234 8517 7238
rect 8535 7235 8574 7254
rect 8593 7248 8600 7249
rect 8599 7241 8600 7248
rect 8583 7238 8584 7241
rect 8599 7238 8612 7241
rect 8535 7234 8565 7235
rect 8574 7234 8580 7235
rect 8583 7234 8612 7238
rect 8502 7233 8612 7234
rect 8502 7232 8618 7233
rect 8177 7224 8228 7232
rect 8177 7212 8202 7224
rect 8209 7212 8228 7224
rect 8259 7224 8309 7232
rect 8259 7216 8275 7224
rect 8282 7222 8309 7224
rect 8318 7222 8539 7232
rect 8282 7212 8539 7222
rect 8568 7224 8618 7232
rect 8568 7215 8584 7224
rect 8177 7204 8228 7212
rect 8275 7204 8539 7212
rect 8565 7212 8584 7215
rect 8591 7212 8618 7224
rect 8565 7204 8618 7212
rect 8193 7196 8194 7204
rect 8209 7196 8222 7204
rect 8193 7188 8209 7196
rect 8190 7181 8209 7184
rect 8190 7172 8212 7181
rect 8163 7162 8212 7172
rect 8163 7156 8193 7162
rect 8212 7157 8217 7162
rect 8135 7140 8209 7156
rect 8227 7148 8257 7204
rect 8292 7194 8500 7204
rect 8535 7200 8580 7204
rect 8583 7203 8584 7204
rect 8599 7203 8612 7204
rect 8318 7164 8507 7194
rect 8333 7161 8507 7164
rect 8326 7158 8507 7161
rect 8135 7138 8148 7140
rect 8163 7138 8197 7140
rect 8135 7122 8209 7138
rect 8236 7134 8249 7148
rect 8264 7134 8280 7150
rect 8326 7145 8337 7158
rect 8119 7100 8120 7116
rect 8135 7100 8148 7122
rect 8163 7100 8193 7122
rect 8236 7118 8298 7134
rect 8326 7127 8337 7143
rect 8342 7138 8352 7158
rect 8362 7138 8376 7158
rect 8379 7145 8388 7158
rect 8404 7145 8413 7158
rect 8342 7127 8376 7138
rect 8379 7127 8388 7143
rect 8404 7127 8413 7143
rect 8420 7138 8430 7158
rect 8440 7138 8454 7158
rect 8455 7145 8466 7158
rect 8420 7127 8454 7138
rect 8455 7127 8466 7143
rect 8512 7134 8528 7150
rect 8535 7148 8565 7200
rect 8599 7196 8600 7203
rect 8584 7188 8600 7196
rect 8571 7156 8584 7175
rect 8599 7156 8629 7172
rect 8571 7140 8645 7156
rect 8571 7138 8584 7140
rect 8599 7138 8633 7140
rect 8236 7116 8249 7118
rect 8264 7116 8298 7118
rect 8236 7100 8298 7116
rect 8342 7111 8358 7114
rect 8420 7111 8450 7122
rect 8498 7118 8544 7134
rect 8571 7122 8645 7138
rect 8498 7116 8532 7118
rect 8497 7100 8544 7116
rect 8571 7100 8584 7122
rect 8599 7100 8629 7122
rect 8656 7100 8657 7116
rect 8672 7100 8685 7260
rect 8715 7156 8728 7260
rect 8773 7238 8774 7248
rect 8789 7238 8802 7248
rect 8773 7234 8802 7238
rect 8807 7234 8837 7260
rect 8855 7246 8871 7248
rect 8943 7246 8996 7260
rect 8944 7244 9008 7246
rect 9051 7244 9066 7260
rect 9115 7257 9145 7260
rect 9115 7254 9151 7257
rect 9081 7246 9097 7248
rect 8855 7234 8870 7238
rect 8773 7232 8870 7234
rect 8898 7232 9066 7244
rect 9082 7234 9097 7238
rect 9115 7235 9154 7254
rect 9173 7248 9180 7249
rect 9179 7241 9180 7248
rect 9163 7238 9164 7241
rect 9179 7238 9192 7241
rect 9115 7234 9145 7235
rect 9154 7234 9160 7235
rect 9163 7234 9192 7238
rect 9082 7233 9192 7234
rect 9082 7232 9198 7233
rect 8757 7224 8808 7232
rect 8757 7212 8782 7224
rect 8789 7212 8808 7224
rect 8839 7224 8889 7232
rect 8839 7216 8855 7224
rect 8862 7222 8889 7224
rect 8898 7222 9119 7232
rect 8862 7212 9119 7222
rect 9148 7224 9198 7232
rect 9148 7215 9164 7224
rect 8757 7204 8808 7212
rect 8855 7204 9119 7212
rect 9145 7212 9164 7215
rect 9171 7212 9198 7224
rect 9145 7204 9198 7212
rect 8773 7196 8774 7204
rect 8789 7196 8802 7204
rect 8773 7188 8789 7196
rect 8770 7181 8789 7184
rect 8770 7172 8792 7181
rect 8743 7162 8792 7172
rect 8743 7156 8773 7162
rect 8792 7157 8797 7162
rect 8715 7140 8789 7156
rect 8807 7148 8837 7204
rect 8872 7194 9080 7204
rect 9115 7200 9160 7204
rect 9163 7203 9164 7204
rect 9179 7203 9192 7204
rect 8898 7164 9087 7194
rect 8913 7161 9087 7164
rect 8906 7158 9087 7161
rect 8715 7138 8728 7140
rect 8743 7138 8777 7140
rect 8715 7122 8789 7138
rect 8816 7134 8829 7148
rect 8844 7134 8860 7150
rect 8906 7145 8917 7158
rect 8699 7100 8700 7116
rect 8715 7100 8728 7122
rect 8743 7100 8773 7122
rect 8816 7118 8878 7134
rect 8906 7127 8917 7143
rect 8922 7138 8932 7158
rect 8942 7138 8956 7158
rect 8959 7145 8968 7158
rect 8984 7145 8993 7158
rect 8922 7127 8956 7138
rect 8959 7127 8968 7143
rect 8984 7127 8993 7143
rect 9000 7138 9010 7158
rect 9020 7138 9034 7158
rect 9035 7145 9046 7158
rect 9000 7127 9034 7138
rect 9035 7127 9046 7143
rect 9092 7134 9108 7150
rect 9115 7148 9145 7200
rect 9179 7196 9180 7203
rect 9164 7188 9180 7196
rect 9151 7156 9164 7175
rect 9179 7156 9209 7172
rect 9151 7140 9225 7156
rect 9151 7138 9164 7140
rect 9179 7138 9213 7140
rect 8816 7116 8829 7118
rect 8844 7116 8878 7118
rect 8816 7100 8878 7116
rect 8922 7111 8938 7114
rect 9000 7111 9030 7122
rect 9078 7118 9124 7134
rect 9151 7122 9225 7138
rect 9078 7116 9112 7118
rect 9077 7100 9124 7116
rect 9151 7100 9164 7122
rect 9179 7100 9209 7122
rect 9236 7100 9237 7116
rect 9252 7100 9265 7260
rect 7496 7092 7531 7100
rect 7496 7066 7497 7092
rect 7504 7066 7531 7092
rect 7439 7048 7469 7062
rect 7496 7058 7531 7066
rect 7533 7092 7574 7100
rect 7533 7066 7548 7092
rect 7555 7066 7574 7092
rect 7638 7088 7700 7100
rect 7712 7088 7787 7100
rect 7845 7088 7920 7100
rect 7932 7088 7963 7100
rect 7969 7088 8004 7100
rect 7638 7086 7800 7088
rect 7533 7058 7574 7066
rect 7656 7062 7669 7086
rect 7684 7084 7699 7086
rect 7496 7048 7525 7058
rect 7539 7048 7568 7058
rect 7583 7048 7613 7062
rect 7656 7048 7699 7062
rect 7723 7059 7730 7066
rect 7733 7062 7800 7086
rect 7832 7086 8004 7088
rect 7802 7064 7830 7068
rect 7832 7064 7912 7086
rect 7933 7084 7948 7086
rect 7802 7062 7912 7064
rect 7733 7058 7912 7062
rect 7706 7048 7736 7058
rect 7738 7048 7891 7058
rect 7899 7048 7929 7058
rect 7933 7048 7963 7062
rect 7991 7048 8004 7086
rect 8076 7092 8111 7100
rect 8076 7066 8077 7092
rect 8084 7066 8111 7092
rect 8019 7048 8049 7062
rect 8076 7058 8111 7066
rect 8113 7092 8154 7100
rect 8113 7066 8128 7092
rect 8135 7066 8154 7092
rect 8218 7088 8280 7100
rect 8292 7088 8367 7100
rect 8425 7088 8500 7100
rect 8512 7088 8543 7100
rect 8549 7088 8584 7100
rect 8218 7086 8380 7088
rect 8113 7058 8154 7066
rect 8236 7062 8249 7086
rect 8264 7084 8279 7086
rect 8076 7048 8077 7058
rect 8092 7048 8105 7058
rect 8119 7048 8120 7058
rect 8135 7048 8148 7058
rect 8163 7048 8193 7062
rect 8236 7048 8279 7062
rect 8303 7059 8310 7066
rect 8313 7062 8380 7086
rect 8412 7086 8584 7088
rect 8382 7064 8410 7068
rect 8412 7064 8492 7086
rect 8513 7084 8528 7086
rect 8382 7062 8492 7064
rect 8313 7058 8492 7062
rect 8286 7048 8316 7058
rect 8318 7048 8471 7058
rect 8479 7048 8509 7058
rect 8513 7048 8543 7062
rect 8571 7048 8584 7086
rect 8656 7092 8691 7100
rect 8656 7066 8657 7092
rect 8664 7066 8691 7092
rect 8599 7048 8629 7062
rect 8656 7058 8691 7066
rect 8693 7092 8734 7100
rect 8693 7066 8708 7092
rect 8715 7066 8734 7092
rect 8798 7088 8860 7100
rect 8872 7088 8947 7100
rect 9005 7088 9080 7100
rect 9092 7088 9123 7100
rect 9129 7088 9164 7100
rect 8798 7086 8960 7088
rect 8693 7058 8734 7066
rect 8816 7062 8829 7086
rect 8844 7084 8859 7086
rect 8656 7048 8657 7058
rect 8672 7048 8685 7058
rect 8699 7048 8700 7058
rect 8715 7048 8728 7058
rect 8743 7048 8773 7062
rect 8816 7048 8859 7062
rect 8883 7059 8890 7066
rect 8893 7062 8960 7086
rect 8992 7086 9164 7088
rect 8962 7064 8990 7068
rect 8992 7064 9072 7086
rect 9093 7084 9108 7086
rect 8962 7062 9072 7064
rect 8893 7058 9072 7062
rect 8866 7048 8896 7058
rect 8898 7048 9051 7058
rect 9059 7048 9089 7058
rect 9093 7048 9123 7062
rect 9151 7048 9164 7086
rect 9236 7092 9271 7100
rect 9236 7066 9237 7092
rect 9244 7066 9271 7092
rect 9179 7048 9209 7062
rect 9236 7058 9271 7066
rect 9236 7048 9237 7058
rect 9252 7048 9265 7058
rect -1 7042 9265 7048
rect 0 7034 9265 7042
rect 15 7004 28 7034
rect 43 7016 73 7034
rect 116 7020 130 7034
rect 166 7020 386 7034
rect 117 7018 130 7020
rect 83 7006 98 7018
rect 80 7004 102 7006
rect 107 7004 137 7018
rect 198 7016 351 7020
rect 180 7004 372 7016
rect 415 7004 445 7018
rect 451 7004 464 7034
rect 479 7016 509 7034
rect 552 7004 565 7034
rect 595 7004 608 7034
rect 623 7016 653 7034
rect 696 7020 710 7034
rect 746 7020 966 7034
rect 697 7018 710 7020
rect 663 7006 678 7018
rect 660 7004 682 7006
rect 687 7004 717 7018
rect 778 7016 931 7020
rect 760 7004 952 7016
rect 995 7004 1025 7018
rect 1031 7004 1044 7034
rect 1059 7016 1089 7034
rect 1132 7004 1145 7034
rect 1175 7004 1188 7034
rect 1203 7016 1233 7034
rect 1276 7020 1290 7034
rect 1326 7020 1546 7034
rect 1277 7018 1290 7020
rect 1243 7006 1258 7018
rect 1240 7004 1262 7006
rect 1267 7004 1297 7018
rect 1358 7016 1511 7020
rect 1340 7004 1532 7016
rect 1575 7004 1605 7018
rect 1611 7004 1624 7034
rect 1639 7016 1669 7034
rect 1712 7004 1725 7034
rect 1755 7004 1768 7034
rect 1783 7020 1813 7034
rect 1856 7020 1899 7034
rect 1906 7020 2126 7034
rect 2133 7020 2163 7034
rect 1823 7006 1838 7018
rect 1857 7006 1870 7020
rect 1938 7016 2091 7020
rect 1820 7004 1842 7006
rect 1920 7004 2112 7016
rect 2191 7004 2204 7034
rect 2219 7020 2249 7034
rect 2286 7004 2305 7034
rect 2320 7004 2326 7034
rect 2335 7004 2348 7034
rect 2363 7020 2393 7034
rect 2436 7020 2479 7034
rect 2486 7020 2706 7034
rect 2713 7020 2743 7034
rect 2403 7006 2418 7018
rect 2437 7006 2450 7020
rect 2518 7016 2671 7020
rect 2400 7004 2422 7006
rect 2500 7004 2692 7016
rect 2771 7004 2784 7034
rect 2799 7020 2829 7034
rect 2866 7004 2885 7034
rect 2900 7004 2906 7034
rect 2915 7004 2928 7034
rect 2943 7020 2973 7034
rect 3016 7020 3059 7034
rect 3066 7020 3286 7034
rect 3293 7020 3323 7034
rect 2983 7006 2998 7018
rect 3017 7006 3030 7020
rect 3098 7016 3251 7020
rect 2980 7004 3002 7006
rect 3080 7004 3272 7016
rect 3351 7004 3364 7034
rect 3379 7020 3409 7034
rect 3446 7004 3465 7034
rect 3480 7004 3486 7034
rect 3495 7004 3508 7034
rect 3523 7020 3553 7034
rect 3596 7020 3639 7034
rect 3646 7020 3866 7034
rect 3873 7020 3903 7034
rect 3563 7006 3578 7018
rect 3597 7006 3610 7020
rect 3678 7016 3831 7020
rect 3560 7004 3582 7006
rect 3660 7004 3852 7016
rect 3931 7004 3944 7034
rect 3959 7020 3989 7034
rect 4026 7004 4045 7034
rect 4060 7004 4066 7034
rect 4075 7004 4088 7034
rect 4103 7020 4133 7034
rect 4176 7020 4219 7034
rect 4226 7020 4446 7034
rect 4453 7020 4483 7034
rect 4143 7006 4158 7018
rect 4177 7006 4190 7020
rect 4258 7016 4411 7020
rect 4140 7004 4162 7006
rect 4240 7004 4432 7016
rect 4511 7004 4524 7034
rect 4539 7020 4569 7034
rect 4606 7004 4625 7034
rect 4640 7004 4646 7034
rect 4655 7004 4668 7034
rect 4683 7020 4713 7034
rect 4756 7020 4799 7034
rect 4806 7020 5026 7034
rect 5033 7020 5063 7034
rect 4723 7006 4738 7018
rect 4757 7006 4770 7020
rect 4838 7016 4991 7020
rect 4720 7004 4742 7006
rect 4820 7004 5012 7016
rect 5091 7004 5104 7034
rect 5119 7020 5149 7034
rect 5186 7004 5205 7034
rect 5220 7004 5226 7034
rect 5235 7004 5248 7034
rect 5263 7020 5293 7034
rect 5336 7020 5379 7034
rect 5386 7020 5606 7034
rect 5613 7020 5643 7034
rect 5303 7006 5318 7018
rect 5337 7006 5350 7020
rect 5418 7016 5571 7020
rect 5300 7004 5322 7006
rect 5400 7004 5592 7016
rect 5671 7004 5684 7034
rect 5699 7020 5729 7034
rect 5766 7004 5785 7034
rect 5800 7004 5806 7034
rect 5815 7004 5828 7034
rect 5843 7020 5873 7034
rect 5916 7020 5959 7034
rect 5966 7020 6186 7034
rect 6193 7020 6223 7034
rect 5883 7006 5898 7018
rect 5917 7006 5930 7020
rect 5998 7016 6151 7020
rect 5880 7004 5902 7006
rect 5980 7004 6172 7016
rect 6251 7004 6264 7034
rect 6279 7020 6309 7034
rect 6346 7004 6365 7034
rect 6380 7004 6386 7034
rect 6395 7004 6408 7034
rect 6423 7020 6453 7034
rect 6496 7020 6539 7034
rect 6546 7020 6766 7034
rect 6773 7020 6803 7034
rect 6463 7006 6478 7018
rect 6497 7006 6510 7020
rect 6578 7016 6731 7020
rect 6460 7004 6482 7006
rect 6560 7004 6752 7016
rect 6831 7004 6844 7034
rect 6859 7020 6889 7034
rect 6926 7004 6945 7034
rect 6960 7004 6966 7034
rect 6975 7004 6988 7034
rect 7003 7020 7033 7034
rect 7076 7020 7119 7034
rect 7126 7020 7346 7034
rect 7353 7020 7383 7034
rect 7043 7006 7058 7018
rect 7077 7006 7090 7020
rect 7158 7016 7311 7020
rect 7040 7004 7062 7006
rect 7140 7004 7332 7016
rect 7411 7004 7424 7034
rect 7439 7020 7469 7034
rect 7506 7004 7525 7034
rect 7540 7004 7546 7034
rect 7555 7004 7568 7034
rect 7583 7016 7613 7034
rect 7656 7020 7670 7034
rect 7706 7020 7926 7034
rect 7657 7018 7670 7020
rect 7623 7006 7638 7018
rect 7620 7004 7642 7006
rect 7647 7004 7677 7018
rect 7738 7016 7891 7020
rect 7720 7004 7912 7016
rect 7955 7004 7985 7018
rect 7991 7004 8004 7034
rect 8019 7016 8049 7034
rect 8092 7004 8105 7034
rect 8135 7004 8148 7034
rect 8163 7016 8193 7034
rect 8236 7020 8250 7034
rect 8286 7020 8506 7034
rect 8237 7018 8250 7020
rect 8203 7006 8218 7018
rect 8200 7004 8222 7006
rect 8227 7004 8257 7018
rect 8318 7016 8471 7020
rect 8300 7004 8492 7016
rect 8535 7004 8565 7018
rect 8571 7004 8584 7034
rect 8599 7016 8629 7034
rect 8672 7004 8685 7034
rect 8715 7004 8728 7034
rect 8743 7016 8773 7034
rect 8816 7020 8830 7034
rect 8866 7020 9086 7034
rect 8817 7018 8830 7020
rect 8783 7006 8798 7018
rect 8780 7004 8802 7006
rect 8807 7004 8837 7018
rect 8898 7016 9051 7020
rect 8880 7004 9072 7016
rect 9115 7004 9145 7018
rect 9151 7004 9164 7034
rect 9179 7016 9209 7034
rect 9252 7004 9265 7034
rect 0 6990 9265 7004
rect 15 6886 28 6990
rect 73 6968 74 6978
rect 89 6968 102 6978
rect 73 6964 102 6968
rect 107 6964 137 6990
rect 155 6976 171 6978
rect 243 6976 296 6990
rect 244 6974 308 6976
rect 351 6974 366 6990
rect 415 6987 445 6990
rect 415 6984 451 6987
rect 381 6976 397 6978
rect 155 6964 170 6968
rect 73 6962 170 6964
rect 198 6962 366 6974
rect 382 6964 397 6968
rect 415 6965 454 6984
rect 473 6978 480 6979
rect 479 6971 480 6978
rect 463 6968 464 6971
rect 479 6968 492 6971
rect 415 6964 445 6965
rect 454 6964 460 6965
rect 463 6964 492 6968
rect 382 6963 492 6964
rect 382 6962 498 6963
rect 57 6954 108 6962
rect 57 6942 82 6954
rect 89 6942 108 6954
rect 139 6954 189 6962
rect 139 6946 155 6954
rect 162 6952 189 6954
rect 198 6952 419 6962
rect 162 6942 419 6952
rect 448 6954 498 6962
rect 448 6945 464 6954
rect 57 6934 108 6942
rect 155 6934 419 6942
rect 445 6942 464 6945
rect 471 6942 498 6954
rect 445 6934 498 6942
rect 73 6926 74 6934
rect 89 6926 102 6934
rect 73 6918 89 6926
rect 70 6911 89 6914
rect 70 6902 92 6911
rect 43 6892 92 6902
rect 43 6886 73 6892
rect 92 6887 97 6892
rect 15 6882 89 6886
rect 107 6882 137 6934
rect 172 6924 380 6934
rect 415 6930 460 6934
rect 463 6933 464 6934
rect 479 6933 492 6934
rect 198 6894 387 6924
rect 213 6891 387 6894
rect 9 6870 89 6882
rect 101 6878 137 6882
rect 206 6888 387 6891
rect 206 6882 217 6888
rect 222 6882 232 6888
rect 242 6882 256 6888
rect 259 6882 268 6888
rect 9 6868 28 6870
rect 43 6868 77 6870
rect 9 6852 89 6868
rect 9 6846 28 6852
rect -1 6830 28 6846
rect 43 6836 73 6852
rect 101 6830 107 6878
rect 110 6872 129 6878
rect 144 6872 174 6880
rect 110 6864 174 6872
rect 110 6848 190 6864
rect 206 6857 268 6882
rect 284 6882 293 6888
rect 300 6882 310 6888
rect 320 6882 334 6888
rect 335 6882 346 6888
rect 284 6857 346 6882
rect 415 6882 445 6930
rect 479 6926 480 6933
rect 464 6918 480 6926
rect 451 6886 464 6905
rect 479 6886 509 6902
rect 451 6882 525 6886
rect 552 6882 565 6990
rect 595 6886 608 6990
rect 653 6968 654 6978
rect 669 6968 682 6978
rect 653 6964 682 6968
rect 687 6964 717 6990
rect 735 6976 751 6978
rect 823 6976 876 6990
rect 824 6974 888 6976
rect 931 6974 946 6990
rect 995 6987 1025 6990
rect 995 6984 1031 6987
rect 961 6976 977 6978
rect 735 6964 750 6968
rect 653 6962 750 6964
rect 778 6962 946 6974
rect 962 6964 977 6968
rect 995 6965 1034 6984
rect 1053 6978 1060 6979
rect 1059 6971 1060 6978
rect 1043 6968 1044 6971
rect 1059 6968 1072 6971
rect 995 6964 1025 6965
rect 1034 6964 1040 6965
rect 1043 6964 1072 6968
rect 962 6963 1072 6964
rect 962 6962 1078 6963
rect 637 6954 688 6962
rect 637 6942 662 6954
rect 669 6942 688 6954
rect 719 6954 769 6962
rect 719 6946 735 6954
rect 742 6952 769 6954
rect 778 6952 999 6962
rect 742 6942 999 6952
rect 1028 6954 1078 6962
rect 1028 6945 1044 6954
rect 637 6934 688 6942
rect 735 6934 999 6942
rect 1025 6942 1044 6945
rect 1051 6942 1078 6954
rect 1025 6934 1078 6942
rect 653 6926 654 6934
rect 669 6926 682 6934
rect 653 6918 669 6926
rect 650 6911 669 6914
rect 650 6902 672 6911
rect 623 6892 672 6902
rect 623 6886 653 6892
rect 672 6887 677 6892
rect 595 6882 669 6886
rect 687 6882 717 6934
rect 752 6924 960 6934
rect 995 6930 1040 6934
rect 1043 6933 1044 6934
rect 1059 6933 1072 6934
rect 778 6894 967 6924
rect 793 6891 967 6894
rect 378 6872 408 6880
rect 415 6878 525 6882
rect 378 6864 423 6872
rect 110 6846 129 6848
rect 144 6846 190 6848
rect 110 6830 190 6846
rect 217 6844 252 6857
rect 293 6854 330 6857
rect 293 6852 335 6854
rect 222 6841 252 6844
rect 231 6837 238 6841
rect 238 6836 239 6837
rect 197 6830 207 6836
rect -7 6822 34 6830
rect -7 6796 8 6822
rect 15 6796 34 6822
rect 98 6818 129 6830
rect 144 6818 247 6830
rect 259 6820 285 6846
rect 300 6841 330 6852
rect 362 6848 424 6864
rect 362 6846 408 6848
rect 362 6830 424 6846
rect 436 6830 442 6878
rect 445 6870 525 6878
rect 445 6868 464 6870
rect 479 6868 513 6870
rect 445 6852 525 6868
rect 445 6830 464 6852
rect 479 6836 509 6852
rect 537 6846 543 6882
rect 546 6846 565 6882
rect 580 6846 586 6882
rect 589 6870 669 6882
rect 681 6878 717 6882
rect 786 6888 967 6891
rect 786 6882 797 6888
rect 802 6882 812 6888
rect 822 6882 836 6888
rect 839 6882 848 6888
rect 589 6868 608 6870
rect 623 6868 657 6870
rect 589 6852 669 6868
rect 589 6846 608 6852
rect 305 6820 408 6830
rect 259 6818 408 6820
rect 429 6818 464 6830
rect 98 6816 260 6818
rect 110 6796 129 6816
rect 144 6814 174 6816
rect -7 6788 34 6796
rect 116 6792 129 6796
rect 181 6800 260 6816
rect 292 6816 464 6818
rect 292 6800 371 6816
rect 378 6814 408 6816
rect -1 6778 28 6788
rect 43 6778 73 6792
rect 116 6778 159 6792
rect 181 6788 371 6800
rect 436 6796 442 6816
rect 166 6778 196 6788
rect 197 6778 355 6788
rect 359 6778 389 6788
rect 393 6778 423 6792
rect 451 6778 464 6816
rect 536 6830 565 6846
rect 579 6830 608 6846
rect 623 6836 653 6852
rect 681 6830 687 6878
rect 690 6872 709 6878
rect 724 6872 754 6880
rect 690 6864 754 6872
rect 690 6848 770 6864
rect 786 6857 848 6882
rect 864 6882 873 6888
rect 880 6882 890 6888
rect 900 6882 914 6888
rect 915 6882 926 6888
rect 864 6857 926 6882
rect 995 6882 1025 6930
rect 1059 6926 1060 6933
rect 1044 6918 1060 6926
rect 1031 6886 1044 6905
rect 1059 6886 1089 6902
rect 1031 6882 1105 6886
rect 1132 6882 1145 6990
rect 1175 6886 1188 6990
rect 1233 6968 1234 6978
rect 1249 6968 1262 6978
rect 1233 6964 1262 6968
rect 1267 6964 1297 6990
rect 1315 6976 1331 6978
rect 1403 6976 1456 6990
rect 1404 6974 1468 6976
rect 1511 6974 1526 6990
rect 1575 6987 1605 6990
rect 1575 6984 1611 6987
rect 1541 6976 1557 6978
rect 1315 6964 1330 6968
rect 1233 6962 1330 6964
rect 1358 6962 1526 6974
rect 1542 6964 1557 6968
rect 1575 6965 1614 6984
rect 1633 6978 1640 6979
rect 1639 6971 1640 6978
rect 1623 6968 1624 6971
rect 1639 6968 1652 6971
rect 1575 6964 1605 6965
rect 1614 6964 1620 6965
rect 1623 6964 1652 6968
rect 1542 6963 1652 6964
rect 1542 6962 1658 6963
rect 1217 6954 1268 6962
rect 1217 6942 1242 6954
rect 1249 6942 1268 6954
rect 1299 6954 1349 6962
rect 1299 6946 1315 6954
rect 1322 6952 1349 6954
rect 1358 6952 1579 6962
rect 1322 6942 1579 6952
rect 1608 6954 1658 6962
rect 1608 6945 1624 6954
rect 1217 6934 1268 6942
rect 1315 6934 1579 6942
rect 1605 6942 1624 6945
rect 1631 6942 1658 6954
rect 1605 6934 1658 6942
rect 1233 6926 1234 6934
rect 1249 6926 1262 6934
rect 1233 6918 1249 6926
rect 1230 6911 1249 6914
rect 1230 6902 1252 6911
rect 1203 6892 1252 6902
rect 1203 6886 1233 6892
rect 1252 6887 1257 6892
rect 1175 6882 1249 6886
rect 1267 6882 1297 6934
rect 1332 6924 1540 6934
rect 1575 6930 1620 6934
rect 1623 6933 1624 6934
rect 1639 6933 1652 6934
rect 1358 6894 1547 6924
rect 1373 6891 1547 6894
rect 958 6872 988 6880
rect 995 6878 1105 6882
rect 958 6864 1003 6872
rect 690 6846 709 6848
rect 724 6846 770 6848
rect 690 6830 770 6846
rect 797 6844 832 6857
rect 873 6854 910 6857
rect 873 6852 915 6854
rect 802 6841 832 6844
rect 811 6837 818 6841
rect 818 6836 819 6837
rect 777 6830 787 6836
rect 536 6822 571 6830
rect 536 6796 537 6822
rect 544 6796 571 6822
rect 479 6778 509 6792
rect 536 6788 571 6796
rect 573 6822 614 6830
rect 573 6796 588 6822
rect 595 6796 614 6822
rect 678 6818 709 6830
rect 724 6818 827 6830
rect 839 6820 865 6846
rect 880 6841 910 6852
rect 942 6848 1004 6864
rect 942 6846 988 6848
rect 942 6830 1004 6846
rect 1016 6830 1022 6878
rect 1025 6870 1105 6878
rect 1025 6868 1044 6870
rect 1059 6868 1093 6870
rect 1025 6852 1105 6868
rect 1025 6830 1044 6852
rect 1059 6836 1089 6852
rect 1117 6846 1123 6882
rect 1126 6846 1145 6882
rect 1160 6846 1166 6882
rect 1169 6870 1249 6882
rect 1261 6878 1297 6882
rect 1366 6888 1547 6891
rect 1366 6882 1377 6888
rect 1382 6882 1392 6888
rect 1402 6882 1416 6888
rect 1419 6882 1428 6888
rect 1169 6868 1188 6870
rect 1203 6868 1237 6870
rect 1169 6852 1249 6868
rect 1169 6846 1188 6852
rect 885 6820 988 6830
rect 839 6818 988 6820
rect 1009 6818 1044 6830
rect 678 6816 840 6818
rect 690 6796 709 6816
rect 724 6814 754 6816
rect 573 6788 614 6796
rect 696 6792 709 6796
rect 761 6800 840 6816
rect 872 6816 1044 6818
rect 872 6800 951 6816
rect 958 6814 988 6816
rect 536 6778 565 6788
rect 579 6778 608 6788
rect 623 6778 653 6792
rect 696 6778 739 6792
rect 761 6788 951 6800
rect 1016 6796 1022 6816
rect 746 6778 776 6788
rect 777 6778 935 6788
rect 939 6778 969 6788
rect 973 6778 1003 6792
rect 1031 6778 1044 6816
rect 1116 6830 1145 6846
rect 1159 6830 1188 6846
rect 1203 6836 1233 6852
rect 1261 6830 1267 6878
rect 1270 6872 1289 6878
rect 1304 6872 1334 6880
rect 1270 6864 1334 6872
rect 1270 6848 1350 6864
rect 1366 6857 1428 6882
rect 1444 6882 1453 6888
rect 1460 6882 1470 6888
rect 1480 6882 1494 6888
rect 1495 6882 1506 6888
rect 1444 6857 1506 6882
rect 1575 6882 1605 6930
rect 1639 6926 1640 6933
rect 1624 6918 1640 6926
rect 1611 6886 1624 6905
rect 1639 6886 1669 6902
rect 1611 6882 1685 6886
rect 1712 6882 1725 6990
rect 1755 6886 1768 6990
rect 1820 6986 1842 6990
rect 1813 6964 1842 6978
rect 1895 6964 1911 6978
rect 1949 6974 1955 6976
rect 1962 6974 2070 6990
rect 2077 6974 2083 6976
rect 2091 6974 2106 6990
rect 2172 6984 2191 6987
rect 1813 6962 1911 6964
rect 1938 6962 2106 6974
rect 2121 6964 2137 6978
rect 2172 6965 2194 6984
rect 2204 6978 2220 6979
rect 2203 6976 2220 6978
rect 2204 6971 2220 6976
rect 2194 6964 2200 6965
rect 2203 6964 2232 6971
rect 2121 6963 2232 6964
rect 2121 6962 2238 6963
rect 1797 6954 1848 6962
rect 1895 6954 1929 6962
rect 1797 6942 1822 6954
rect 1829 6942 1848 6954
rect 1902 6952 1929 6954
rect 1938 6952 2159 6962
rect 2194 6959 2200 6962
rect 1902 6948 2159 6952
rect 1797 6934 1848 6942
rect 1895 6934 2159 6948
rect 2203 6954 2238 6962
rect 1813 6926 1842 6934
rect 1813 6920 1830 6926
rect 1813 6918 1847 6920
rect 1895 6918 1911 6934
rect 1912 6924 2120 6934
rect 2121 6924 2137 6934
rect 2185 6930 2200 6945
rect 2203 6942 2204 6954
rect 2211 6942 2238 6954
rect 2203 6934 2238 6942
rect 2203 6933 2232 6934
rect 1923 6920 2137 6924
rect 1938 6918 2137 6920
rect 2172 6920 2185 6930
rect 2203 6920 2220 6933
rect 2172 6918 2220 6920
rect 1814 6914 1847 6918
rect 1810 6912 1847 6914
rect 1810 6911 1877 6912
rect 1810 6906 1841 6911
rect 1847 6906 1877 6911
rect 1810 6902 1877 6906
rect 1783 6899 1877 6902
rect 1783 6892 1832 6899
rect 1783 6886 1813 6892
rect 1832 6887 1837 6892
rect 1755 6882 1829 6886
rect 1538 6872 1568 6880
rect 1575 6878 1685 6882
rect 1538 6864 1583 6872
rect 1270 6846 1289 6848
rect 1304 6846 1350 6848
rect 1270 6830 1350 6846
rect 1377 6844 1412 6857
rect 1453 6854 1490 6857
rect 1453 6852 1495 6854
rect 1382 6841 1412 6844
rect 1391 6837 1398 6841
rect 1398 6836 1399 6837
rect 1357 6830 1367 6836
rect 1116 6822 1151 6830
rect 1116 6796 1117 6822
rect 1124 6796 1151 6822
rect 1059 6778 1089 6792
rect 1116 6788 1151 6796
rect 1153 6822 1194 6830
rect 1153 6796 1168 6822
rect 1175 6796 1194 6822
rect 1258 6818 1289 6830
rect 1304 6818 1407 6830
rect 1419 6820 1445 6846
rect 1460 6841 1490 6852
rect 1522 6848 1584 6864
rect 1522 6846 1568 6848
rect 1522 6830 1584 6846
rect 1596 6830 1602 6878
rect 1605 6870 1685 6878
rect 1605 6868 1624 6870
rect 1639 6868 1673 6870
rect 1605 6852 1685 6868
rect 1605 6830 1624 6852
rect 1639 6836 1669 6852
rect 1697 6846 1703 6882
rect 1706 6846 1725 6882
rect 1740 6846 1746 6882
rect 1749 6870 1829 6882
rect 1841 6878 1877 6899
rect 1938 6894 2127 6918
rect 2172 6917 2219 6918
rect 2185 6912 2219 6917
rect 1953 6891 2127 6894
rect 1946 6888 2127 6891
rect 2155 6911 2219 6912
rect 1749 6868 1768 6870
rect 1783 6868 1817 6870
rect 1749 6852 1829 6868
rect 1749 6846 1768 6852
rect 1465 6820 1568 6830
rect 1419 6818 1568 6820
rect 1589 6818 1624 6830
rect 1258 6816 1420 6818
rect 1270 6796 1289 6816
rect 1304 6814 1334 6816
rect 1153 6788 1194 6796
rect 1276 6792 1289 6796
rect 1341 6800 1420 6816
rect 1452 6816 1624 6818
rect 1452 6800 1531 6816
rect 1538 6814 1568 6816
rect 1116 6778 1145 6788
rect 1159 6778 1188 6788
rect 1203 6778 1233 6792
rect 1276 6778 1319 6792
rect 1341 6788 1531 6800
rect 1596 6796 1602 6816
rect 1326 6778 1356 6788
rect 1357 6778 1515 6788
rect 1519 6778 1549 6788
rect 1553 6778 1583 6792
rect 1611 6778 1624 6816
rect 1696 6830 1725 6846
rect 1739 6830 1768 6846
rect 1783 6836 1813 6852
rect 1841 6830 1847 6878
rect 1850 6872 1869 6878
rect 1884 6872 1914 6880
rect 1850 6864 1914 6872
rect 1850 6848 1930 6864
rect 1946 6857 2008 6888
rect 2024 6857 2086 6888
rect 2155 6886 2204 6911
rect 2219 6886 2249 6902
rect 2118 6872 2148 6880
rect 2155 6878 2265 6886
rect 2118 6864 2163 6872
rect 1850 6846 1869 6848
rect 1884 6846 1930 6848
rect 1850 6830 1930 6846
rect 1957 6844 1992 6857
rect 2033 6854 2070 6857
rect 2033 6852 2075 6854
rect 1962 6841 1992 6844
rect 1971 6837 1978 6841
rect 1978 6836 1979 6837
rect 1937 6830 1947 6836
rect 1696 6822 1731 6830
rect 1696 6796 1697 6822
rect 1704 6796 1731 6822
rect 1639 6778 1669 6792
rect 1696 6788 1731 6796
rect 1733 6822 1774 6830
rect 1733 6796 1748 6822
rect 1755 6796 1774 6822
rect 1838 6818 1869 6830
rect 1884 6818 1987 6830
rect 1999 6820 2025 6846
rect 2040 6841 2070 6852
rect 2102 6848 2164 6864
rect 2102 6846 2148 6848
rect 2102 6830 2164 6846
rect 2176 6830 2182 6878
rect 2185 6870 2265 6878
rect 2185 6868 2204 6870
rect 2219 6868 2253 6870
rect 2185 6852 2265 6868
rect 2185 6830 2204 6852
rect 2219 6836 2249 6852
rect 2277 6846 2283 6920
rect 2286 6846 2305 6990
rect 2320 6846 2326 6990
rect 2335 6920 2348 6990
rect 2400 6986 2422 6990
rect 2393 6964 2422 6978
rect 2475 6964 2491 6978
rect 2529 6974 2535 6976
rect 2542 6974 2650 6990
rect 2657 6974 2663 6976
rect 2671 6974 2686 6990
rect 2752 6984 2771 6987
rect 2393 6962 2491 6964
rect 2518 6962 2686 6974
rect 2701 6964 2717 6978
rect 2752 6965 2774 6984
rect 2784 6978 2800 6979
rect 2783 6976 2800 6978
rect 2784 6971 2800 6976
rect 2774 6964 2780 6965
rect 2783 6964 2812 6971
rect 2701 6963 2812 6964
rect 2701 6962 2818 6963
rect 2377 6954 2428 6962
rect 2475 6954 2509 6962
rect 2377 6942 2402 6954
rect 2409 6942 2428 6954
rect 2482 6952 2509 6954
rect 2518 6952 2739 6962
rect 2774 6959 2780 6962
rect 2482 6948 2739 6952
rect 2377 6934 2428 6942
rect 2475 6934 2739 6948
rect 2783 6954 2818 6962
rect 2329 6886 2348 6920
rect 2393 6926 2422 6934
rect 2393 6920 2410 6926
rect 2393 6918 2427 6920
rect 2475 6918 2491 6934
rect 2492 6924 2700 6934
rect 2701 6924 2717 6934
rect 2765 6930 2780 6945
rect 2783 6942 2784 6954
rect 2791 6942 2818 6954
rect 2783 6934 2818 6942
rect 2783 6933 2812 6934
rect 2503 6920 2717 6924
rect 2518 6918 2717 6920
rect 2752 6920 2765 6930
rect 2783 6920 2800 6933
rect 2752 6918 2800 6920
rect 2394 6914 2427 6918
rect 2390 6912 2427 6914
rect 2390 6911 2457 6912
rect 2390 6906 2421 6911
rect 2427 6906 2457 6911
rect 2390 6902 2457 6906
rect 2363 6899 2457 6902
rect 2363 6892 2412 6899
rect 2363 6886 2393 6892
rect 2412 6887 2417 6892
rect 2329 6870 2409 6886
rect 2421 6878 2457 6899
rect 2518 6894 2707 6918
rect 2752 6917 2799 6918
rect 2765 6912 2799 6917
rect 2533 6891 2707 6894
rect 2526 6888 2707 6891
rect 2735 6911 2799 6912
rect 2329 6868 2348 6870
rect 2363 6868 2397 6870
rect 2329 6852 2409 6868
rect 2329 6846 2348 6852
rect 2045 6820 2148 6830
rect 1999 6818 2148 6820
rect 2169 6818 2204 6830
rect 1838 6816 2000 6818
rect 1850 6796 1869 6816
rect 1884 6814 1914 6816
rect 1733 6788 1774 6796
rect 1856 6792 1869 6796
rect 1921 6800 2000 6816
rect 2032 6816 2204 6818
rect 2032 6800 2111 6816
rect 2118 6814 2148 6816
rect 1696 6778 1725 6788
rect 1739 6778 1768 6788
rect 1783 6778 1813 6792
rect 1856 6778 1899 6792
rect 1921 6788 2111 6800
rect 2176 6796 2182 6816
rect 1906 6778 1936 6788
rect 1937 6778 2095 6788
rect 2099 6778 2129 6788
rect 2133 6778 2163 6792
rect 2191 6778 2204 6816
rect 2276 6830 2305 6846
rect 2319 6830 2348 6846
rect 2363 6836 2393 6852
rect 2421 6830 2427 6878
rect 2430 6872 2449 6878
rect 2464 6872 2494 6880
rect 2430 6864 2494 6872
rect 2430 6848 2510 6864
rect 2526 6857 2588 6888
rect 2604 6857 2666 6888
rect 2735 6886 2784 6911
rect 2799 6886 2829 6902
rect 2698 6872 2728 6880
rect 2735 6878 2845 6886
rect 2698 6864 2743 6872
rect 2430 6846 2449 6848
rect 2464 6846 2510 6848
rect 2430 6830 2510 6846
rect 2537 6844 2572 6857
rect 2613 6854 2650 6857
rect 2613 6852 2655 6854
rect 2542 6841 2572 6844
rect 2551 6837 2558 6841
rect 2558 6836 2559 6837
rect 2517 6830 2527 6836
rect 2276 6822 2311 6830
rect 2276 6796 2277 6822
rect 2284 6796 2311 6822
rect 2219 6778 2249 6792
rect 2276 6788 2311 6796
rect 2313 6822 2354 6830
rect 2313 6796 2328 6822
rect 2335 6796 2354 6822
rect 2418 6818 2449 6830
rect 2464 6818 2567 6830
rect 2579 6820 2605 6846
rect 2620 6841 2650 6852
rect 2682 6848 2744 6864
rect 2682 6846 2728 6848
rect 2682 6830 2744 6846
rect 2756 6830 2762 6878
rect 2765 6870 2845 6878
rect 2765 6868 2784 6870
rect 2799 6868 2833 6870
rect 2765 6852 2845 6868
rect 2765 6830 2784 6852
rect 2799 6836 2829 6852
rect 2857 6846 2863 6920
rect 2866 6846 2885 6990
rect 2900 6846 2906 6990
rect 2915 6920 2928 6990
rect 2980 6986 3002 6990
rect 2973 6964 3002 6978
rect 3055 6964 3071 6978
rect 3109 6974 3115 6976
rect 3122 6974 3230 6990
rect 3237 6974 3243 6976
rect 3251 6974 3266 6990
rect 3332 6984 3351 6987
rect 2973 6962 3071 6964
rect 3098 6962 3266 6974
rect 3281 6964 3297 6978
rect 3332 6965 3354 6984
rect 3364 6978 3380 6979
rect 3363 6976 3380 6978
rect 3364 6971 3380 6976
rect 3354 6964 3360 6965
rect 3363 6964 3392 6971
rect 3281 6963 3392 6964
rect 3281 6962 3398 6963
rect 2957 6954 3008 6962
rect 3055 6954 3089 6962
rect 2957 6942 2982 6954
rect 2989 6942 3008 6954
rect 3062 6952 3089 6954
rect 3098 6952 3319 6962
rect 3354 6959 3360 6962
rect 3062 6948 3319 6952
rect 2957 6934 3008 6942
rect 3055 6934 3319 6948
rect 3363 6954 3398 6962
rect 2909 6886 2928 6920
rect 2973 6926 3002 6934
rect 2973 6920 2990 6926
rect 2973 6918 3007 6920
rect 3055 6918 3071 6934
rect 3072 6924 3280 6934
rect 3281 6924 3297 6934
rect 3345 6930 3360 6945
rect 3363 6942 3364 6954
rect 3371 6942 3398 6954
rect 3363 6934 3398 6942
rect 3363 6933 3392 6934
rect 3083 6920 3297 6924
rect 3098 6918 3297 6920
rect 3332 6920 3345 6930
rect 3363 6920 3380 6933
rect 3332 6918 3380 6920
rect 2974 6914 3007 6918
rect 2970 6912 3007 6914
rect 2970 6911 3037 6912
rect 2970 6906 3001 6911
rect 3007 6906 3037 6911
rect 2970 6902 3037 6906
rect 2943 6899 3037 6902
rect 2943 6892 2992 6899
rect 2943 6886 2973 6892
rect 2992 6887 2997 6892
rect 2909 6870 2989 6886
rect 3001 6878 3037 6899
rect 3098 6894 3287 6918
rect 3332 6917 3379 6918
rect 3345 6912 3379 6917
rect 3113 6891 3287 6894
rect 3106 6888 3287 6891
rect 3315 6911 3379 6912
rect 2909 6868 2928 6870
rect 2943 6868 2977 6870
rect 2909 6852 2989 6868
rect 2909 6846 2928 6852
rect 2625 6820 2728 6830
rect 2579 6818 2728 6820
rect 2749 6818 2784 6830
rect 2418 6816 2580 6818
rect 2430 6796 2449 6816
rect 2464 6814 2494 6816
rect 2313 6788 2354 6796
rect 2436 6792 2449 6796
rect 2501 6800 2580 6816
rect 2612 6816 2784 6818
rect 2612 6800 2691 6816
rect 2698 6814 2728 6816
rect 2276 6778 2305 6788
rect 2319 6778 2348 6788
rect 2363 6778 2393 6792
rect 2436 6778 2479 6792
rect 2501 6788 2691 6800
rect 2756 6796 2762 6816
rect 2486 6778 2516 6788
rect 2517 6778 2675 6788
rect 2679 6778 2709 6788
rect 2713 6778 2743 6792
rect 2771 6778 2784 6816
rect 2856 6830 2885 6846
rect 2899 6830 2928 6846
rect 2943 6836 2973 6852
rect 3001 6830 3007 6878
rect 3010 6872 3029 6878
rect 3044 6872 3074 6880
rect 3010 6864 3074 6872
rect 3010 6848 3090 6864
rect 3106 6857 3168 6888
rect 3184 6857 3246 6888
rect 3315 6886 3364 6911
rect 3379 6886 3409 6902
rect 3278 6872 3308 6880
rect 3315 6878 3425 6886
rect 3278 6864 3323 6872
rect 3010 6846 3029 6848
rect 3044 6846 3090 6848
rect 3010 6830 3090 6846
rect 3117 6844 3152 6857
rect 3193 6854 3230 6857
rect 3193 6852 3235 6854
rect 3122 6841 3152 6844
rect 3131 6837 3138 6841
rect 3138 6836 3139 6837
rect 3097 6830 3107 6836
rect 2856 6822 2891 6830
rect 2856 6796 2857 6822
rect 2864 6796 2891 6822
rect 2799 6778 2829 6792
rect 2856 6788 2891 6796
rect 2893 6822 2934 6830
rect 2893 6796 2908 6822
rect 2915 6796 2934 6822
rect 2998 6818 3029 6830
rect 3044 6818 3147 6830
rect 3159 6820 3185 6846
rect 3200 6841 3230 6852
rect 3262 6848 3324 6864
rect 3262 6846 3308 6848
rect 3262 6830 3324 6846
rect 3336 6830 3342 6878
rect 3345 6870 3425 6878
rect 3345 6868 3364 6870
rect 3379 6868 3413 6870
rect 3345 6852 3425 6868
rect 3345 6830 3364 6852
rect 3379 6836 3409 6852
rect 3437 6846 3443 6920
rect 3446 6846 3465 6990
rect 3480 6846 3486 6990
rect 3495 6920 3508 6990
rect 3560 6986 3582 6990
rect 3553 6964 3582 6978
rect 3635 6964 3651 6978
rect 3689 6974 3695 6976
rect 3702 6974 3810 6990
rect 3817 6974 3823 6976
rect 3831 6974 3846 6990
rect 3912 6984 3931 6987
rect 3553 6962 3651 6964
rect 3678 6962 3846 6974
rect 3861 6964 3877 6978
rect 3912 6965 3934 6984
rect 3944 6978 3960 6979
rect 3943 6976 3960 6978
rect 3944 6971 3960 6976
rect 3934 6964 3940 6965
rect 3943 6964 3972 6971
rect 3861 6963 3972 6964
rect 3861 6962 3978 6963
rect 3537 6954 3588 6962
rect 3635 6954 3669 6962
rect 3537 6942 3562 6954
rect 3569 6942 3588 6954
rect 3642 6952 3669 6954
rect 3678 6952 3899 6962
rect 3934 6959 3940 6962
rect 3642 6948 3899 6952
rect 3537 6934 3588 6942
rect 3635 6934 3899 6948
rect 3943 6954 3978 6962
rect 3489 6886 3508 6920
rect 3553 6926 3582 6934
rect 3553 6920 3570 6926
rect 3553 6918 3587 6920
rect 3635 6918 3651 6934
rect 3652 6924 3860 6934
rect 3861 6924 3877 6934
rect 3925 6930 3940 6945
rect 3943 6942 3944 6954
rect 3951 6942 3978 6954
rect 3943 6934 3978 6942
rect 3943 6933 3972 6934
rect 3663 6920 3877 6924
rect 3678 6918 3877 6920
rect 3912 6920 3925 6930
rect 3943 6920 3960 6933
rect 3912 6918 3960 6920
rect 3554 6914 3587 6918
rect 3550 6912 3587 6914
rect 3550 6911 3617 6912
rect 3550 6906 3581 6911
rect 3587 6906 3617 6911
rect 3550 6902 3617 6906
rect 3523 6899 3617 6902
rect 3523 6892 3572 6899
rect 3523 6886 3553 6892
rect 3572 6887 3577 6892
rect 3489 6870 3569 6886
rect 3581 6878 3617 6899
rect 3678 6894 3867 6918
rect 3912 6917 3959 6918
rect 3925 6912 3959 6917
rect 3693 6891 3867 6894
rect 3686 6888 3867 6891
rect 3895 6911 3959 6912
rect 3489 6868 3508 6870
rect 3523 6868 3557 6870
rect 3489 6852 3569 6868
rect 3489 6846 3508 6852
rect 3205 6820 3308 6830
rect 3159 6818 3308 6820
rect 3329 6818 3364 6830
rect 2998 6816 3160 6818
rect 3010 6796 3029 6816
rect 3044 6814 3074 6816
rect 2893 6788 2934 6796
rect 3016 6792 3029 6796
rect 3081 6800 3160 6816
rect 3192 6816 3364 6818
rect 3192 6800 3271 6816
rect 3278 6814 3308 6816
rect 2856 6778 2885 6788
rect 2899 6778 2928 6788
rect 2943 6778 2973 6792
rect 3016 6778 3059 6792
rect 3081 6788 3271 6800
rect 3336 6796 3342 6816
rect 3066 6778 3096 6788
rect 3097 6778 3255 6788
rect 3259 6778 3289 6788
rect 3293 6778 3323 6792
rect 3351 6778 3364 6816
rect 3436 6830 3465 6846
rect 3479 6830 3508 6846
rect 3523 6836 3553 6852
rect 3581 6830 3587 6878
rect 3590 6872 3609 6878
rect 3624 6872 3654 6880
rect 3590 6864 3654 6872
rect 3590 6848 3670 6864
rect 3686 6857 3748 6888
rect 3764 6857 3826 6888
rect 3895 6886 3944 6911
rect 3959 6886 3989 6902
rect 3858 6872 3888 6880
rect 3895 6878 4005 6886
rect 3858 6864 3903 6872
rect 3590 6846 3609 6848
rect 3624 6846 3670 6848
rect 3590 6830 3670 6846
rect 3697 6844 3732 6857
rect 3773 6854 3810 6857
rect 3773 6852 3815 6854
rect 3702 6841 3732 6844
rect 3711 6837 3718 6841
rect 3718 6836 3719 6837
rect 3677 6830 3687 6836
rect 3436 6822 3471 6830
rect 3436 6796 3437 6822
rect 3444 6796 3471 6822
rect 3379 6778 3409 6792
rect 3436 6788 3471 6796
rect 3473 6822 3514 6830
rect 3473 6796 3488 6822
rect 3495 6796 3514 6822
rect 3578 6818 3609 6830
rect 3624 6818 3727 6830
rect 3739 6820 3765 6846
rect 3780 6841 3810 6852
rect 3842 6848 3904 6864
rect 3842 6846 3888 6848
rect 3842 6830 3904 6846
rect 3916 6830 3922 6878
rect 3925 6870 4005 6878
rect 3925 6868 3944 6870
rect 3959 6868 3993 6870
rect 3925 6852 4005 6868
rect 3925 6830 3944 6852
rect 3959 6836 3989 6852
rect 4017 6846 4023 6920
rect 4026 6846 4045 6990
rect 4060 6846 4066 6990
rect 4075 6920 4088 6990
rect 4140 6986 4162 6990
rect 4133 6964 4162 6978
rect 4215 6964 4231 6978
rect 4269 6974 4275 6976
rect 4282 6974 4390 6990
rect 4397 6974 4403 6976
rect 4411 6974 4426 6990
rect 4492 6984 4511 6987
rect 4133 6962 4231 6964
rect 4258 6962 4426 6974
rect 4441 6964 4457 6978
rect 4492 6965 4514 6984
rect 4524 6978 4540 6979
rect 4523 6976 4540 6978
rect 4524 6971 4540 6976
rect 4514 6964 4520 6965
rect 4523 6964 4552 6971
rect 4441 6963 4552 6964
rect 4441 6962 4558 6963
rect 4117 6954 4168 6962
rect 4215 6954 4249 6962
rect 4117 6942 4142 6954
rect 4149 6942 4168 6954
rect 4222 6952 4249 6954
rect 4258 6952 4479 6962
rect 4514 6959 4520 6962
rect 4222 6948 4479 6952
rect 4117 6934 4168 6942
rect 4215 6934 4479 6948
rect 4523 6954 4558 6962
rect 4069 6886 4088 6920
rect 4133 6926 4162 6934
rect 4133 6920 4150 6926
rect 4133 6918 4167 6920
rect 4215 6918 4231 6934
rect 4232 6924 4440 6934
rect 4441 6924 4457 6934
rect 4505 6930 4520 6945
rect 4523 6942 4524 6954
rect 4531 6942 4558 6954
rect 4523 6934 4558 6942
rect 4523 6933 4552 6934
rect 4243 6920 4457 6924
rect 4258 6918 4457 6920
rect 4492 6920 4505 6930
rect 4523 6920 4540 6933
rect 4492 6918 4540 6920
rect 4134 6914 4167 6918
rect 4130 6912 4167 6914
rect 4130 6911 4197 6912
rect 4130 6906 4161 6911
rect 4167 6906 4197 6911
rect 4130 6902 4197 6906
rect 4103 6899 4197 6902
rect 4103 6892 4152 6899
rect 4103 6886 4133 6892
rect 4152 6887 4157 6892
rect 4069 6870 4149 6886
rect 4161 6878 4197 6899
rect 4258 6894 4447 6918
rect 4492 6917 4539 6918
rect 4505 6912 4539 6917
rect 4273 6891 4447 6894
rect 4266 6888 4447 6891
rect 4475 6911 4539 6912
rect 4069 6868 4088 6870
rect 4103 6868 4137 6870
rect 4069 6852 4149 6868
rect 4069 6846 4088 6852
rect 3785 6820 3888 6830
rect 3739 6818 3888 6820
rect 3909 6818 3944 6830
rect 3578 6816 3740 6818
rect 3590 6796 3609 6816
rect 3624 6814 3654 6816
rect 3473 6788 3514 6796
rect 3596 6792 3609 6796
rect 3661 6800 3740 6816
rect 3772 6816 3944 6818
rect 3772 6800 3851 6816
rect 3858 6814 3888 6816
rect 3436 6778 3465 6788
rect 3479 6778 3508 6788
rect 3523 6778 3553 6792
rect 3596 6778 3639 6792
rect 3661 6788 3851 6800
rect 3916 6796 3922 6816
rect 3646 6778 3676 6788
rect 3677 6778 3835 6788
rect 3839 6778 3869 6788
rect 3873 6778 3903 6792
rect 3931 6778 3944 6816
rect 4016 6830 4045 6846
rect 4059 6830 4088 6846
rect 4103 6836 4133 6852
rect 4161 6830 4167 6878
rect 4170 6872 4189 6878
rect 4204 6872 4234 6880
rect 4170 6864 4234 6872
rect 4170 6848 4250 6864
rect 4266 6857 4328 6888
rect 4344 6857 4406 6888
rect 4475 6886 4524 6911
rect 4539 6886 4569 6902
rect 4438 6872 4468 6880
rect 4475 6878 4585 6886
rect 4438 6864 4483 6872
rect 4170 6846 4189 6848
rect 4204 6846 4250 6848
rect 4170 6830 4250 6846
rect 4277 6844 4312 6857
rect 4353 6854 4390 6857
rect 4353 6852 4395 6854
rect 4282 6841 4312 6844
rect 4291 6837 4298 6841
rect 4298 6836 4299 6837
rect 4257 6830 4267 6836
rect 4016 6822 4051 6830
rect 4016 6796 4017 6822
rect 4024 6796 4051 6822
rect 3959 6778 3989 6792
rect 4016 6788 4051 6796
rect 4053 6822 4094 6830
rect 4053 6796 4068 6822
rect 4075 6796 4094 6822
rect 4158 6818 4189 6830
rect 4204 6818 4307 6830
rect 4319 6820 4345 6846
rect 4360 6841 4390 6852
rect 4422 6848 4484 6864
rect 4422 6846 4468 6848
rect 4422 6830 4484 6846
rect 4496 6830 4502 6878
rect 4505 6870 4585 6878
rect 4505 6868 4524 6870
rect 4539 6868 4573 6870
rect 4505 6852 4585 6868
rect 4505 6830 4524 6852
rect 4539 6836 4569 6852
rect 4597 6846 4603 6920
rect 4606 6846 4625 6990
rect 4640 6846 4646 6990
rect 4655 6920 4668 6990
rect 4720 6986 4742 6990
rect 4713 6964 4742 6978
rect 4795 6964 4811 6978
rect 4849 6974 4855 6976
rect 4862 6974 4970 6990
rect 4977 6974 4983 6976
rect 4991 6974 5006 6990
rect 5072 6984 5091 6987
rect 4713 6962 4811 6964
rect 4838 6962 5006 6974
rect 5021 6964 5037 6978
rect 5072 6965 5094 6984
rect 5104 6978 5120 6979
rect 5103 6976 5120 6978
rect 5104 6971 5120 6976
rect 5094 6964 5100 6965
rect 5103 6964 5132 6971
rect 5021 6963 5132 6964
rect 5021 6962 5138 6963
rect 4697 6954 4748 6962
rect 4795 6954 4829 6962
rect 4697 6942 4722 6954
rect 4729 6942 4748 6954
rect 4802 6952 4829 6954
rect 4838 6952 5059 6962
rect 5094 6959 5100 6962
rect 4802 6948 5059 6952
rect 4697 6934 4748 6942
rect 4795 6934 5059 6948
rect 5103 6954 5138 6962
rect 4649 6886 4668 6920
rect 4713 6926 4742 6934
rect 4713 6920 4730 6926
rect 4713 6918 4747 6920
rect 4795 6918 4811 6934
rect 4812 6924 5020 6934
rect 5021 6924 5037 6934
rect 5085 6930 5100 6945
rect 5103 6942 5104 6954
rect 5111 6942 5138 6954
rect 5103 6934 5138 6942
rect 5103 6933 5132 6934
rect 4823 6920 5037 6924
rect 4838 6918 5037 6920
rect 5072 6920 5085 6930
rect 5103 6920 5120 6933
rect 5072 6918 5120 6920
rect 4714 6914 4747 6918
rect 4710 6912 4747 6914
rect 4710 6911 4777 6912
rect 4710 6906 4741 6911
rect 4747 6906 4777 6911
rect 4710 6902 4777 6906
rect 4683 6899 4777 6902
rect 4683 6892 4732 6899
rect 4683 6886 4713 6892
rect 4732 6887 4737 6892
rect 4649 6870 4729 6886
rect 4741 6878 4777 6899
rect 4838 6894 5027 6918
rect 5072 6917 5119 6918
rect 5085 6912 5119 6917
rect 4853 6891 5027 6894
rect 4846 6888 5027 6891
rect 5055 6911 5119 6912
rect 4649 6868 4668 6870
rect 4683 6868 4717 6870
rect 4649 6852 4729 6868
rect 4649 6846 4668 6852
rect 4365 6820 4468 6830
rect 4319 6818 4468 6820
rect 4489 6818 4524 6830
rect 4158 6816 4320 6818
rect 4170 6796 4189 6816
rect 4204 6814 4234 6816
rect 4053 6788 4094 6796
rect 4176 6792 4189 6796
rect 4241 6800 4320 6816
rect 4352 6816 4524 6818
rect 4352 6800 4431 6816
rect 4438 6814 4468 6816
rect 4016 6778 4045 6788
rect 4059 6778 4088 6788
rect 4103 6778 4133 6792
rect 4176 6778 4219 6792
rect 4241 6788 4431 6800
rect 4496 6796 4502 6816
rect 4226 6778 4256 6788
rect 4257 6778 4415 6788
rect 4419 6778 4449 6788
rect 4453 6778 4483 6792
rect 4511 6778 4524 6816
rect 4596 6830 4625 6846
rect 4639 6830 4668 6846
rect 4683 6836 4713 6852
rect 4741 6830 4747 6878
rect 4750 6872 4769 6878
rect 4784 6872 4814 6880
rect 4750 6864 4814 6872
rect 4750 6848 4830 6864
rect 4846 6857 4908 6888
rect 4924 6857 4986 6888
rect 5055 6886 5104 6911
rect 5119 6886 5149 6902
rect 5018 6872 5048 6880
rect 5055 6878 5165 6886
rect 5018 6864 5063 6872
rect 4750 6846 4769 6848
rect 4784 6846 4830 6848
rect 4750 6830 4830 6846
rect 4857 6844 4892 6857
rect 4933 6854 4970 6857
rect 4933 6852 4975 6854
rect 4862 6841 4892 6844
rect 4871 6837 4878 6841
rect 4878 6836 4879 6837
rect 4837 6830 4847 6836
rect 4596 6822 4631 6830
rect 4596 6796 4597 6822
rect 4604 6796 4631 6822
rect 4539 6778 4569 6792
rect 4596 6788 4631 6796
rect 4633 6822 4674 6830
rect 4633 6796 4648 6822
rect 4655 6796 4674 6822
rect 4738 6818 4769 6830
rect 4784 6818 4887 6830
rect 4899 6820 4925 6846
rect 4940 6841 4970 6852
rect 5002 6848 5064 6864
rect 5002 6846 5048 6848
rect 5002 6830 5064 6846
rect 5076 6830 5082 6878
rect 5085 6870 5165 6878
rect 5085 6868 5104 6870
rect 5119 6868 5153 6870
rect 5085 6852 5165 6868
rect 5085 6830 5104 6852
rect 5119 6836 5149 6852
rect 5177 6846 5183 6920
rect 5186 6846 5205 6990
rect 5220 6846 5226 6990
rect 5235 6920 5248 6990
rect 5300 6986 5322 6990
rect 5293 6964 5322 6978
rect 5375 6964 5391 6978
rect 5429 6974 5435 6976
rect 5442 6974 5550 6990
rect 5557 6974 5563 6976
rect 5571 6974 5586 6990
rect 5652 6984 5671 6987
rect 5293 6962 5391 6964
rect 5418 6962 5586 6974
rect 5601 6964 5617 6978
rect 5652 6965 5674 6984
rect 5684 6978 5700 6979
rect 5683 6976 5700 6978
rect 5684 6971 5700 6976
rect 5674 6964 5680 6965
rect 5683 6964 5712 6971
rect 5601 6963 5712 6964
rect 5601 6962 5718 6963
rect 5277 6954 5328 6962
rect 5375 6954 5409 6962
rect 5277 6942 5302 6954
rect 5309 6942 5328 6954
rect 5382 6952 5409 6954
rect 5418 6952 5639 6962
rect 5674 6959 5680 6962
rect 5382 6948 5639 6952
rect 5277 6934 5328 6942
rect 5375 6934 5639 6948
rect 5683 6954 5718 6962
rect 5229 6886 5248 6920
rect 5293 6926 5322 6934
rect 5293 6920 5310 6926
rect 5293 6918 5327 6920
rect 5375 6918 5391 6934
rect 5392 6924 5600 6934
rect 5601 6924 5617 6934
rect 5665 6930 5680 6945
rect 5683 6942 5684 6954
rect 5691 6942 5718 6954
rect 5683 6934 5718 6942
rect 5683 6933 5712 6934
rect 5403 6920 5617 6924
rect 5418 6918 5617 6920
rect 5652 6920 5665 6930
rect 5683 6920 5700 6933
rect 5652 6918 5700 6920
rect 5294 6914 5327 6918
rect 5290 6912 5327 6914
rect 5290 6911 5357 6912
rect 5290 6906 5321 6911
rect 5327 6906 5357 6911
rect 5290 6902 5357 6906
rect 5263 6899 5357 6902
rect 5263 6892 5312 6899
rect 5263 6886 5293 6892
rect 5312 6887 5317 6892
rect 5229 6870 5309 6886
rect 5321 6878 5357 6899
rect 5418 6894 5607 6918
rect 5652 6917 5699 6918
rect 5665 6912 5699 6917
rect 5433 6891 5607 6894
rect 5426 6888 5607 6891
rect 5635 6911 5699 6912
rect 5229 6868 5248 6870
rect 5263 6868 5297 6870
rect 5229 6852 5309 6868
rect 5229 6846 5248 6852
rect 4945 6820 5048 6830
rect 4899 6818 5048 6820
rect 5069 6818 5104 6830
rect 4738 6816 4900 6818
rect 4750 6796 4769 6816
rect 4784 6814 4814 6816
rect 4633 6788 4674 6796
rect 4756 6792 4769 6796
rect 4821 6800 4900 6816
rect 4932 6816 5104 6818
rect 4932 6800 5011 6816
rect 5018 6814 5048 6816
rect 4596 6778 4625 6788
rect 4639 6778 4668 6788
rect 4683 6778 4713 6792
rect 4756 6778 4799 6792
rect 4821 6788 5011 6800
rect 5076 6796 5082 6816
rect 4806 6778 4836 6788
rect 4837 6778 4995 6788
rect 4999 6778 5029 6788
rect 5033 6778 5063 6792
rect 5091 6778 5104 6816
rect 5176 6830 5205 6846
rect 5219 6830 5248 6846
rect 5263 6836 5293 6852
rect 5321 6830 5327 6878
rect 5330 6872 5349 6878
rect 5364 6872 5394 6880
rect 5330 6864 5394 6872
rect 5330 6848 5410 6864
rect 5426 6857 5488 6888
rect 5504 6857 5566 6888
rect 5635 6886 5684 6911
rect 5699 6886 5729 6902
rect 5598 6872 5628 6880
rect 5635 6878 5745 6886
rect 5598 6864 5643 6872
rect 5330 6846 5349 6848
rect 5364 6846 5410 6848
rect 5330 6830 5410 6846
rect 5437 6844 5472 6857
rect 5513 6854 5550 6857
rect 5513 6852 5555 6854
rect 5442 6841 5472 6844
rect 5451 6837 5458 6841
rect 5458 6836 5459 6837
rect 5417 6830 5427 6836
rect 5176 6822 5211 6830
rect 5176 6796 5177 6822
rect 5184 6796 5211 6822
rect 5119 6778 5149 6792
rect 5176 6788 5211 6796
rect 5213 6822 5254 6830
rect 5213 6796 5228 6822
rect 5235 6796 5254 6822
rect 5318 6818 5349 6830
rect 5364 6818 5467 6830
rect 5479 6820 5505 6846
rect 5520 6841 5550 6852
rect 5582 6848 5644 6864
rect 5582 6846 5628 6848
rect 5582 6830 5644 6846
rect 5656 6830 5662 6878
rect 5665 6870 5745 6878
rect 5665 6868 5684 6870
rect 5699 6868 5733 6870
rect 5665 6852 5745 6868
rect 5665 6830 5684 6852
rect 5699 6836 5729 6852
rect 5757 6846 5763 6920
rect 5766 6846 5785 6990
rect 5800 6846 5806 6990
rect 5815 6920 5828 6990
rect 5880 6986 5902 6990
rect 5873 6964 5902 6978
rect 5955 6964 5971 6978
rect 6009 6974 6015 6976
rect 6022 6974 6130 6990
rect 6137 6974 6143 6976
rect 6151 6974 6166 6990
rect 6232 6984 6251 6987
rect 5873 6962 5971 6964
rect 5998 6962 6166 6974
rect 6181 6964 6197 6978
rect 6232 6965 6254 6984
rect 6264 6978 6280 6979
rect 6263 6976 6280 6978
rect 6264 6971 6280 6976
rect 6254 6964 6260 6965
rect 6263 6964 6292 6971
rect 6181 6963 6292 6964
rect 6181 6962 6298 6963
rect 5857 6954 5908 6962
rect 5955 6954 5989 6962
rect 5857 6942 5882 6954
rect 5889 6942 5908 6954
rect 5962 6952 5989 6954
rect 5998 6952 6219 6962
rect 6254 6959 6260 6962
rect 5962 6948 6219 6952
rect 5857 6934 5908 6942
rect 5955 6934 6219 6948
rect 6263 6954 6298 6962
rect 5809 6886 5828 6920
rect 5873 6926 5902 6934
rect 5873 6920 5890 6926
rect 5873 6918 5907 6920
rect 5955 6918 5971 6934
rect 5972 6924 6180 6934
rect 6181 6924 6197 6934
rect 6245 6930 6260 6945
rect 6263 6942 6264 6954
rect 6271 6942 6298 6954
rect 6263 6934 6298 6942
rect 6263 6933 6292 6934
rect 5983 6920 6197 6924
rect 5998 6918 6197 6920
rect 6232 6920 6245 6930
rect 6263 6920 6280 6933
rect 6232 6918 6280 6920
rect 5874 6914 5907 6918
rect 5870 6912 5907 6914
rect 5870 6911 5937 6912
rect 5870 6906 5901 6911
rect 5907 6906 5937 6911
rect 5870 6902 5937 6906
rect 5843 6899 5937 6902
rect 5843 6892 5892 6899
rect 5843 6886 5873 6892
rect 5892 6887 5897 6892
rect 5809 6870 5889 6886
rect 5901 6878 5937 6899
rect 5998 6894 6187 6918
rect 6232 6917 6279 6918
rect 6245 6912 6279 6917
rect 6013 6891 6187 6894
rect 6006 6888 6187 6891
rect 6215 6911 6279 6912
rect 5809 6868 5828 6870
rect 5843 6868 5877 6870
rect 5809 6852 5889 6868
rect 5809 6846 5828 6852
rect 5525 6820 5628 6830
rect 5479 6818 5628 6820
rect 5649 6818 5684 6830
rect 5318 6816 5480 6818
rect 5330 6796 5349 6816
rect 5364 6814 5394 6816
rect 5213 6788 5254 6796
rect 5336 6792 5349 6796
rect 5401 6800 5480 6816
rect 5512 6816 5684 6818
rect 5512 6800 5591 6816
rect 5598 6814 5628 6816
rect 5176 6778 5205 6788
rect 5219 6778 5248 6788
rect 5263 6778 5293 6792
rect 5336 6778 5379 6792
rect 5401 6788 5591 6800
rect 5656 6796 5662 6816
rect 5386 6778 5416 6788
rect 5417 6778 5575 6788
rect 5579 6778 5609 6788
rect 5613 6778 5643 6792
rect 5671 6778 5684 6816
rect 5756 6830 5785 6846
rect 5799 6830 5828 6846
rect 5843 6836 5873 6852
rect 5901 6830 5907 6878
rect 5910 6872 5929 6878
rect 5944 6872 5974 6880
rect 5910 6864 5974 6872
rect 5910 6848 5990 6864
rect 6006 6857 6068 6888
rect 6084 6857 6146 6888
rect 6215 6886 6264 6911
rect 6279 6886 6309 6902
rect 6178 6872 6208 6880
rect 6215 6878 6325 6886
rect 6178 6864 6223 6872
rect 5910 6846 5929 6848
rect 5944 6846 5990 6848
rect 5910 6830 5990 6846
rect 6017 6844 6052 6857
rect 6093 6854 6130 6857
rect 6093 6852 6135 6854
rect 6022 6841 6052 6844
rect 6031 6837 6038 6841
rect 6038 6836 6039 6837
rect 5997 6830 6007 6836
rect 5756 6822 5791 6830
rect 5756 6796 5757 6822
rect 5764 6796 5791 6822
rect 5699 6778 5729 6792
rect 5756 6788 5791 6796
rect 5793 6822 5834 6830
rect 5793 6796 5808 6822
rect 5815 6796 5834 6822
rect 5898 6818 5929 6830
rect 5944 6818 6047 6830
rect 6059 6820 6085 6846
rect 6100 6841 6130 6852
rect 6162 6848 6224 6864
rect 6162 6846 6208 6848
rect 6162 6830 6224 6846
rect 6236 6830 6242 6878
rect 6245 6870 6325 6878
rect 6245 6868 6264 6870
rect 6279 6868 6313 6870
rect 6245 6852 6325 6868
rect 6245 6830 6264 6852
rect 6279 6836 6309 6852
rect 6337 6846 6343 6920
rect 6346 6846 6365 6990
rect 6380 6846 6386 6990
rect 6395 6920 6408 6990
rect 6460 6986 6482 6990
rect 6453 6964 6482 6978
rect 6535 6964 6551 6978
rect 6589 6974 6595 6976
rect 6602 6974 6710 6990
rect 6717 6974 6723 6976
rect 6731 6974 6746 6990
rect 6812 6984 6831 6987
rect 6453 6962 6551 6964
rect 6578 6962 6746 6974
rect 6761 6964 6777 6978
rect 6812 6965 6834 6984
rect 6844 6978 6860 6979
rect 6843 6976 6860 6978
rect 6844 6971 6860 6976
rect 6834 6964 6840 6965
rect 6843 6964 6872 6971
rect 6761 6963 6872 6964
rect 6761 6962 6878 6963
rect 6437 6954 6488 6962
rect 6535 6954 6569 6962
rect 6437 6942 6462 6954
rect 6469 6942 6488 6954
rect 6542 6952 6569 6954
rect 6578 6952 6799 6962
rect 6834 6959 6840 6962
rect 6542 6948 6799 6952
rect 6437 6934 6488 6942
rect 6535 6934 6799 6948
rect 6843 6954 6878 6962
rect 6389 6886 6408 6920
rect 6453 6926 6482 6934
rect 6453 6920 6470 6926
rect 6453 6918 6487 6920
rect 6535 6918 6551 6934
rect 6552 6924 6760 6934
rect 6761 6924 6777 6934
rect 6825 6930 6840 6945
rect 6843 6942 6844 6954
rect 6851 6942 6878 6954
rect 6843 6934 6878 6942
rect 6843 6933 6872 6934
rect 6563 6920 6777 6924
rect 6578 6918 6777 6920
rect 6812 6920 6825 6930
rect 6843 6920 6860 6933
rect 6812 6918 6860 6920
rect 6454 6914 6487 6918
rect 6450 6912 6487 6914
rect 6450 6911 6517 6912
rect 6450 6906 6481 6911
rect 6487 6906 6517 6911
rect 6450 6902 6517 6906
rect 6423 6899 6517 6902
rect 6423 6892 6472 6899
rect 6423 6886 6453 6892
rect 6472 6887 6477 6892
rect 6389 6870 6469 6886
rect 6481 6878 6517 6899
rect 6578 6894 6767 6918
rect 6812 6917 6859 6918
rect 6825 6912 6859 6917
rect 6593 6891 6767 6894
rect 6586 6888 6767 6891
rect 6795 6911 6859 6912
rect 6389 6868 6408 6870
rect 6423 6868 6457 6870
rect 6389 6852 6469 6868
rect 6389 6846 6408 6852
rect 6105 6820 6208 6830
rect 6059 6818 6208 6820
rect 6229 6818 6264 6830
rect 5898 6816 6060 6818
rect 5910 6796 5929 6816
rect 5944 6814 5974 6816
rect 5793 6788 5834 6796
rect 5916 6792 5929 6796
rect 5981 6800 6060 6816
rect 6092 6816 6264 6818
rect 6092 6800 6171 6816
rect 6178 6814 6208 6816
rect 5756 6778 5785 6788
rect 5799 6778 5828 6788
rect 5843 6778 5873 6792
rect 5916 6778 5959 6792
rect 5981 6788 6171 6800
rect 6236 6796 6242 6816
rect 5966 6778 5996 6788
rect 5997 6778 6155 6788
rect 6159 6778 6189 6788
rect 6193 6778 6223 6792
rect 6251 6778 6264 6816
rect 6336 6830 6365 6846
rect 6379 6830 6408 6846
rect 6423 6836 6453 6852
rect 6481 6830 6487 6878
rect 6490 6872 6509 6878
rect 6524 6872 6554 6880
rect 6490 6864 6554 6872
rect 6490 6848 6570 6864
rect 6586 6857 6648 6888
rect 6664 6857 6726 6888
rect 6795 6886 6844 6911
rect 6859 6886 6889 6902
rect 6758 6872 6788 6880
rect 6795 6878 6905 6886
rect 6758 6864 6803 6872
rect 6490 6846 6509 6848
rect 6524 6846 6570 6848
rect 6490 6830 6570 6846
rect 6597 6844 6632 6857
rect 6673 6854 6710 6857
rect 6673 6852 6715 6854
rect 6602 6841 6632 6844
rect 6611 6837 6618 6841
rect 6618 6836 6619 6837
rect 6577 6830 6587 6836
rect 6336 6822 6371 6830
rect 6336 6796 6337 6822
rect 6344 6796 6371 6822
rect 6279 6778 6309 6792
rect 6336 6788 6371 6796
rect 6373 6822 6414 6830
rect 6373 6796 6388 6822
rect 6395 6796 6414 6822
rect 6478 6818 6509 6830
rect 6524 6818 6627 6830
rect 6639 6820 6665 6846
rect 6680 6841 6710 6852
rect 6742 6848 6804 6864
rect 6742 6846 6788 6848
rect 6742 6830 6804 6846
rect 6816 6830 6822 6878
rect 6825 6870 6905 6878
rect 6825 6868 6844 6870
rect 6859 6868 6893 6870
rect 6825 6852 6905 6868
rect 6825 6830 6844 6852
rect 6859 6836 6889 6852
rect 6917 6846 6923 6920
rect 6926 6846 6945 6990
rect 6960 6846 6966 6990
rect 6975 6920 6988 6990
rect 7040 6986 7062 6990
rect 7033 6964 7062 6978
rect 7115 6964 7131 6978
rect 7169 6974 7175 6976
rect 7182 6974 7290 6990
rect 7297 6974 7303 6976
rect 7311 6974 7326 6990
rect 7392 6984 7411 6987
rect 7033 6962 7131 6964
rect 7158 6962 7326 6974
rect 7341 6964 7357 6978
rect 7392 6965 7414 6984
rect 7424 6978 7440 6979
rect 7423 6976 7440 6978
rect 7424 6971 7440 6976
rect 7414 6964 7420 6965
rect 7423 6964 7452 6971
rect 7341 6963 7452 6964
rect 7341 6962 7458 6963
rect 7017 6954 7068 6962
rect 7115 6954 7149 6962
rect 7017 6942 7042 6954
rect 7049 6942 7068 6954
rect 7122 6952 7149 6954
rect 7158 6952 7379 6962
rect 7414 6959 7420 6962
rect 7122 6948 7379 6952
rect 7017 6934 7068 6942
rect 7115 6934 7379 6948
rect 7423 6954 7458 6962
rect 6969 6886 6988 6920
rect 7033 6926 7062 6934
rect 7033 6920 7050 6926
rect 7033 6918 7067 6920
rect 7115 6918 7131 6934
rect 7132 6924 7340 6934
rect 7341 6924 7357 6934
rect 7405 6930 7420 6945
rect 7423 6942 7424 6954
rect 7431 6942 7458 6954
rect 7423 6934 7458 6942
rect 7423 6933 7452 6934
rect 7143 6920 7357 6924
rect 7158 6918 7357 6920
rect 7392 6920 7405 6930
rect 7423 6920 7440 6933
rect 7392 6918 7440 6920
rect 7034 6914 7067 6918
rect 7030 6912 7067 6914
rect 7030 6911 7097 6912
rect 7030 6906 7061 6911
rect 7067 6906 7097 6911
rect 7030 6902 7097 6906
rect 7003 6899 7097 6902
rect 7003 6892 7052 6899
rect 7003 6886 7033 6892
rect 7052 6887 7057 6892
rect 6969 6870 7049 6886
rect 7061 6878 7097 6899
rect 7158 6894 7347 6918
rect 7392 6917 7439 6918
rect 7405 6912 7439 6917
rect 7173 6891 7347 6894
rect 7166 6888 7347 6891
rect 7375 6911 7439 6912
rect 6969 6868 6988 6870
rect 7003 6868 7037 6870
rect 6969 6852 7049 6868
rect 6969 6846 6988 6852
rect 6685 6820 6788 6830
rect 6639 6818 6788 6820
rect 6809 6818 6844 6830
rect 6478 6816 6640 6818
rect 6490 6796 6509 6816
rect 6524 6814 6554 6816
rect 6373 6788 6414 6796
rect 6496 6792 6509 6796
rect 6561 6800 6640 6816
rect 6672 6816 6844 6818
rect 6672 6800 6751 6816
rect 6758 6814 6788 6816
rect 6336 6778 6365 6788
rect 6379 6778 6408 6788
rect 6423 6778 6453 6792
rect 6496 6778 6539 6792
rect 6561 6788 6751 6800
rect 6816 6796 6822 6816
rect 6546 6778 6576 6788
rect 6577 6778 6735 6788
rect 6739 6778 6769 6788
rect 6773 6778 6803 6792
rect 6831 6778 6844 6816
rect 6916 6830 6945 6846
rect 6959 6830 6988 6846
rect 7003 6836 7033 6852
rect 7061 6830 7067 6878
rect 7070 6872 7089 6878
rect 7104 6872 7134 6880
rect 7070 6864 7134 6872
rect 7070 6848 7150 6864
rect 7166 6857 7228 6888
rect 7244 6857 7306 6888
rect 7375 6886 7424 6911
rect 7439 6886 7469 6902
rect 7338 6872 7368 6880
rect 7375 6878 7485 6886
rect 7338 6864 7383 6872
rect 7070 6846 7089 6848
rect 7104 6846 7150 6848
rect 7070 6830 7150 6846
rect 7177 6844 7212 6857
rect 7253 6854 7290 6857
rect 7253 6852 7295 6854
rect 7182 6841 7212 6844
rect 7191 6837 7198 6841
rect 7198 6836 7199 6837
rect 7157 6830 7167 6836
rect 6916 6822 6951 6830
rect 6916 6796 6917 6822
rect 6924 6796 6951 6822
rect 6859 6778 6889 6792
rect 6916 6788 6951 6796
rect 6953 6822 6994 6830
rect 6953 6796 6968 6822
rect 6975 6796 6994 6822
rect 7058 6818 7089 6830
rect 7104 6818 7207 6830
rect 7219 6820 7245 6846
rect 7260 6841 7290 6852
rect 7322 6848 7384 6864
rect 7322 6846 7368 6848
rect 7322 6830 7384 6846
rect 7396 6830 7402 6878
rect 7405 6870 7485 6878
rect 7405 6868 7424 6870
rect 7439 6868 7473 6870
rect 7405 6852 7485 6868
rect 7405 6830 7424 6852
rect 7439 6836 7469 6852
rect 7497 6846 7503 6920
rect 7506 6846 7525 6990
rect 7540 6846 7546 6990
rect 7555 6920 7568 6990
rect 7613 6968 7614 6978
rect 7629 6968 7642 6978
rect 7613 6964 7642 6968
rect 7647 6964 7677 6990
rect 7695 6976 7711 6978
rect 7783 6976 7836 6990
rect 7784 6974 7848 6976
rect 7891 6974 7906 6990
rect 7955 6987 7985 6990
rect 7955 6984 7991 6987
rect 7921 6976 7937 6978
rect 7695 6964 7710 6968
rect 7613 6962 7710 6964
rect 7738 6962 7906 6974
rect 7922 6964 7937 6968
rect 7955 6965 7994 6984
rect 8013 6978 8020 6979
rect 8019 6971 8020 6978
rect 8003 6968 8004 6971
rect 8019 6968 8032 6971
rect 7955 6964 7985 6965
rect 7994 6964 8000 6965
rect 8003 6964 8032 6968
rect 7922 6963 8032 6964
rect 7922 6962 8038 6963
rect 7597 6954 7648 6962
rect 7597 6942 7622 6954
rect 7629 6942 7648 6954
rect 7679 6954 7729 6962
rect 7679 6946 7695 6954
rect 7702 6952 7729 6954
rect 7738 6952 7959 6962
rect 7702 6942 7959 6952
rect 7988 6954 8038 6962
rect 7988 6945 8004 6954
rect 7597 6934 7648 6942
rect 7695 6934 7959 6942
rect 7985 6942 8004 6945
rect 8011 6942 8038 6954
rect 7985 6934 8038 6942
rect 7549 6886 7568 6920
rect 7613 6926 7614 6934
rect 7629 6926 7642 6934
rect 7613 6918 7629 6926
rect 7610 6911 7629 6914
rect 7610 6902 7632 6911
rect 7583 6892 7632 6902
rect 7583 6886 7613 6892
rect 7632 6887 7637 6892
rect 7549 6870 7629 6886
rect 7647 6878 7677 6934
rect 7712 6924 7920 6934
rect 7955 6930 8000 6934
rect 8003 6933 8004 6934
rect 8019 6933 8032 6934
rect 7738 6894 7927 6924
rect 7753 6891 7927 6894
rect 7746 6888 7927 6891
rect 7549 6868 7568 6870
rect 7583 6868 7617 6870
rect 7549 6852 7629 6868
rect 7656 6864 7669 6878
rect 7684 6864 7700 6880
rect 7746 6875 7757 6888
rect 7549 6846 7568 6852
rect 7265 6820 7368 6830
rect 7219 6818 7368 6820
rect 7389 6818 7424 6830
rect 7058 6816 7220 6818
rect 7070 6796 7089 6816
rect 7104 6814 7134 6816
rect 6953 6788 6994 6796
rect 7076 6792 7089 6796
rect 7141 6800 7220 6816
rect 7252 6816 7424 6818
rect 7252 6800 7331 6816
rect 7338 6814 7368 6816
rect 6916 6778 6945 6788
rect 6959 6778 6988 6788
rect 7003 6778 7033 6792
rect 7076 6778 7119 6792
rect 7141 6788 7331 6800
rect 7396 6796 7402 6816
rect 7126 6778 7156 6788
rect 7157 6778 7315 6788
rect 7319 6778 7349 6788
rect 7353 6778 7383 6792
rect 7411 6778 7424 6816
rect 7496 6830 7525 6846
rect 7539 6830 7568 6846
rect 7583 6830 7613 6852
rect 7656 6848 7718 6864
rect 7746 6857 7757 6873
rect 7762 6868 7772 6888
rect 7782 6868 7796 6888
rect 7799 6875 7808 6888
rect 7824 6875 7833 6888
rect 7762 6857 7796 6868
rect 7799 6857 7808 6873
rect 7824 6857 7833 6873
rect 7840 6868 7850 6888
rect 7860 6868 7874 6888
rect 7875 6875 7886 6888
rect 7840 6857 7874 6868
rect 7875 6857 7886 6873
rect 7932 6864 7948 6880
rect 7955 6878 7985 6930
rect 8019 6926 8020 6933
rect 8004 6918 8020 6926
rect 7991 6886 8004 6905
rect 8019 6886 8049 6902
rect 7991 6870 8065 6886
rect 7991 6868 8004 6870
rect 8019 6868 8053 6870
rect 7656 6846 7669 6848
rect 7684 6846 7718 6848
rect 7656 6830 7718 6846
rect 7762 6841 7778 6844
rect 7840 6841 7870 6852
rect 7918 6848 7964 6864
rect 7991 6852 8065 6868
rect 7918 6846 7952 6848
rect 7917 6830 7964 6846
rect 7991 6830 8004 6852
rect 8019 6830 8049 6852
rect 8076 6830 8077 6846
rect 8092 6830 8105 6990
rect 8135 6886 8148 6990
rect 8193 6968 8194 6978
rect 8209 6968 8222 6978
rect 8193 6964 8222 6968
rect 8227 6964 8257 6990
rect 8275 6976 8291 6978
rect 8363 6976 8416 6990
rect 8364 6974 8428 6976
rect 8471 6974 8486 6990
rect 8535 6987 8565 6990
rect 8535 6984 8571 6987
rect 8501 6976 8517 6978
rect 8275 6964 8290 6968
rect 8193 6962 8290 6964
rect 8318 6962 8486 6974
rect 8502 6964 8517 6968
rect 8535 6965 8574 6984
rect 8593 6978 8600 6979
rect 8599 6971 8600 6978
rect 8583 6968 8584 6971
rect 8599 6968 8612 6971
rect 8535 6964 8565 6965
rect 8574 6964 8580 6965
rect 8583 6964 8612 6968
rect 8502 6963 8612 6964
rect 8502 6962 8618 6963
rect 8177 6954 8228 6962
rect 8177 6942 8202 6954
rect 8209 6942 8228 6954
rect 8259 6954 8309 6962
rect 8259 6946 8275 6954
rect 8282 6952 8309 6954
rect 8318 6952 8539 6962
rect 8282 6942 8539 6952
rect 8568 6954 8618 6962
rect 8568 6945 8584 6954
rect 8177 6934 8228 6942
rect 8275 6934 8539 6942
rect 8565 6942 8584 6945
rect 8591 6942 8618 6954
rect 8565 6934 8618 6942
rect 8193 6926 8194 6934
rect 8209 6926 8222 6934
rect 8193 6918 8209 6926
rect 8190 6911 8209 6914
rect 8190 6902 8212 6911
rect 8163 6892 8212 6902
rect 8163 6886 8193 6892
rect 8212 6887 8217 6892
rect 8135 6870 8209 6886
rect 8227 6878 8257 6934
rect 8292 6924 8500 6934
rect 8535 6930 8580 6934
rect 8583 6933 8584 6934
rect 8599 6933 8612 6934
rect 8318 6894 8507 6924
rect 8333 6891 8507 6894
rect 8326 6888 8507 6891
rect 8135 6868 8148 6870
rect 8163 6868 8197 6870
rect 8135 6852 8209 6868
rect 8236 6864 8249 6878
rect 8264 6864 8280 6880
rect 8326 6875 8337 6888
rect 8119 6830 8120 6846
rect 8135 6830 8148 6852
rect 8163 6830 8193 6852
rect 8236 6848 8298 6864
rect 8326 6857 8337 6873
rect 8342 6868 8352 6888
rect 8362 6868 8376 6888
rect 8379 6875 8388 6888
rect 8404 6875 8413 6888
rect 8342 6857 8376 6868
rect 8379 6857 8388 6873
rect 8404 6857 8413 6873
rect 8420 6868 8430 6888
rect 8440 6868 8454 6888
rect 8455 6875 8466 6888
rect 8420 6857 8454 6868
rect 8455 6857 8466 6873
rect 8512 6864 8528 6880
rect 8535 6878 8565 6930
rect 8599 6926 8600 6933
rect 8584 6918 8600 6926
rect 8571 6886 8584 6905
rect 8599 6886 8629 6902
rect 8571 6870 8645 6886
rect 8571 6868 8584 6870
rect 8599 6868 8633 6870
rect 8236 6846 8249 6848
rect 8264 6846 8298 6848
rect 8236 6830 8298 6846
rect 8342 6841 8358 6844
rect 8420 6841 8450 6852
rect 8498 6848 8544 6864
rect 8571 6852 8645 6868
rect 8498 6846 8532 6848
rect 8497 6830 8544 6846
rect 8571 6830 8584 6852
rect 8599 6830 8629 6852
rect 8656 6830 8657 6846
rect 8672 6830 8685 6990
rect 8715 6886 8728 6990
rect 8773 6968 8774 6978
rect 8789 6968 8802 6978
rect 8773 6964 8802 6968
rect 8807 6964 8837 6990
rect 8855 6976 8871 6978
rect 8943 6976 8996 6990
rect 8944 6974 9008 6976
rect 9051 6974 9066 6990
rect 9115 6987 9145 6990
rect 9115 6984 9151 6987
rect 9081 6976 9097 6978
rect 8855 6964 8870 6968
rect 8773 6962 8870 6964
rect 8898 6962 9066 6974
rect 9082 6964 9097 6968
rect 9115 6965 9154 6984
rect 9173 6978 9180 6979
rect 9179 6971 9180 6978
rect 9163 6968 9164 6971
rect 9179 6968 9192 6971
rect 9115 6964 9145 6965
rect 9154 6964 9160 6965
rect 9163 6964 9192 6968
rect 9082 6963 9192 6964
rect 9082 6962 9198 6963
rect 8757 6954 8808 6962
rect 8757 6942 8782 6954
rect 8789 6942 8808 6954
rect 8839 6954 8889 6962
rect 8839 6946 8855 6954
rect 8862 6952 8889 6954
rect 8898 6952 9119 6962
rect 8862 6942 9119 6952
rect 9148 6954 9198 6962
rect 9148 6945 9164 6954
rect 8757 6934 8808 6942
rect 8855 6934 9119 6942
rect 9145 6942 9164 6945
rect 9171 6942 9198 6954
rect 9145 6934 9198 6942
rect 8773 6926 8774 6934
rect 8789 6926 8802 6934
rect 8773 6918 8789 6926
rect 8770 6911 8789 6914
rect 8770 6902 8792 6911
rect 8743 6892 8792 6902
rect 8743 6886 8773 6892
rect 8792 6887 8797 6892
rect 8715 6870 8789 6886
rect 8807 6878 8837 6934
rect 8872 6924 9080 6934
rect 9115 6930 9160 6934
rect 9163 6933 9164 6934
rect 9179 6933 9192 6934
rect 8898 6894 9087 6924
rect 8913 6891 9087 6894
rect 8906 6888 9087 6891
rect 8715 6868 8728 6870
rect 8743 6868 8777 6870
rect 8715 6852 8789 6868
rect 8816 6864 8829 6878
rect 8844 6864 8860 6880
rect 8906 6875 8917 6888
rect 8699 6830 8700 6846
rect 8715 6830 8728 6852
rect 8743 6830 8773 6852
rect 8816 6848 8878 6864
rect 8906 6857 8917 6873
rect 8922 6868 8932 6888
rect 8942 6868 8956 6888
rect 8959 6875 8968 6888
rect 8984 6875 8993 6888
rect 8922 6857 8956 6868
rect 8959 6857 8968 6873
rect 8984 6857 8993 6873
rect 9000 6868 9010 6888
rect 9020 6868 9034 6888
rect 9035 6875 9046 6888
rect 9000 6857 9034 6868
rect 9035 6857 9046 6873
rect 9092 6864 9108 6880
rect 9115 6878 9145 6930
rect 9179 6926 9180 6933
rect 9164 6918 9180 6926
rect 9151 6886 9164 6905
rect 9179 6886 9209 6902
rect 9151 6870 9225 6886
rect 9151 6868 9164 6870
rect 9179 6868 9213 6870
rect 8816 6846 8829 6848
rect 8844 6846 8878 6848
rect 8816 6830 8878 6846
rect 8922 6841 8938 6844
rect 9000 6841 9030 6852
rect 9078 6848 9124 6864
rect 9151 6852 9225 6868
rect 9078 6846 9112 6848
rect 9077 6830 9124 6846
rect 9151 6830 9164 6852
rect 9179 6830 9209 6852
rect 9236 6830 9237 6846
rect 9252 6830 9265 6990
rect 7496 6822 7531 6830
rect 7496 6796 7497 6822
rect 7504 6796 7531 6822
rect 7439 6778 7469 6792
rect 7496 6788 7531 6796
rect 7533 6822 7574 6830
rect 7533 6796 7548 6822
rect 7555 6796 7574 6822
rect 7638 6818 7700 6830
rect 7712 6818 7787 6830
rect 7845 6818 7920 6830
rect 7932 6818 7963 6830
rect 7969 6818 8004 6830
rect 7638 6816 7800 6818
rect 7533 6788 7574 6796
rect 7656 6792 7669 6816
rect 7684 6814 7699 6816
rect 7496 6778 7525 6788
rect 7539 6778 7568 6788
rect 7583 6778 7613 6792
rect 7656 6778 7699 6792
rect 7723 6789 7730 6796
rect 7733 6792 7800 6816
rect 7832 6816 8004 6818
rect 7802 6794 7830 6798
rect 7832 6794 7912 6816
rect 7933 6814 7948 6816
rect 7802 6792 7912 6794
rect 7733 6788 7912 6792
rect 7706 6778 7736 6788
rect 7738 6778 7891 6788
rect 7899 6778 7929 6788
rect 7933 6778 7963 6792
rect 7991 6778 8004 6816
rect 8076 6822 8111 6830
rect 8076 6796 8077 6822
rect 8084 6796 8111 6822
rect 8019 6778 8049 6792
rect 8076 6788 8111 6796
rect 8113 6822 8154 6830
rect 8113 6796 8128 6822
rect 8135 6796 8154 6822
rect 8218 6818 8280 6830
rect 8292 6818 8367 6830
rect 8425 6818 8500 6830
rect 8512 6818 8543 6830
rect 8549 6818 8584 6830
rect 8218 6816 8380 6818
rect 8113 6788 8154 6796
rect 8236 6792 8249 6816
rect 8264 6814 8279 6816
rect 8076 6778 8077 6788
rect 8092 6778 8105 6788
rect 8119 6778 8120 6788
rect 8135 6778 8148 6788
rect 8163 6778 8193 6792
rect 8236 6778 8279 6792
rect 8303 6789 8310 6796
rect 8313 6792 8380 6816
rect 8412 6816 8584 6818
rect 8382 6794 8410 6798
rect 8412 6794 8492 6816
rect 8513 6814 8528 6816
rect 8382 6792 8492 6794
rect 8313 6788 8492 6792
rect 8286 6778 8316 6788
rect 8318 6778 8471 6788
rect 8479 6778 8509 6788
rect 8513 6778 8543 6792
rect 8571 6778 8584 6816
rect 8656 6822 8691 6830
rect 8656 6796 8657 6822
rect 8664 6796 8691 6822
rect 8599 6778 8629 6792
rect 8656 6788 8691 6796
rect 8693 6822 8734 6830
rect 8693 6796 8708 6822
rect 8715 6796 8734 6822
rect 8798 6818 8860 6830
rect 8872 6818 8947 6830
rect 9005 6818 9080 6830
rect 9092 6818 9123 6830
rect 9129 6818 9164 6830
rect 8798 6816 8960 6818
rect 8693 6788 8734 6796
rect 8816 6792 8829 6816
rect 8844 6814 8859 6816
rect 8656 6778 8657 6788
rect 8672 6778 8685 6788
rect 8699 6778 8700 6788
rect 8715 6778 8728 6788
rect 8743 6778 8773 6792
rect 8816 6778 8859 6792
rect 8883 6789 8890 6796
rect 8893 6792 8960 6816
rect 8992 6816 9164 6818
rect 8962 6794 8990 6798
rect 8992 6794 9072 6816
rect 9093 6814 9108 6816
rect 8962 6792 9072 6794
rect 8893 6788 9072 6792
rect 8866 6778 8896 6788
rect 8898 6778 9051 6788
rect 9059 6778 9089 6788
rect 9093 6778 9123 6792
rect 9151 6778 9164 6816
rect 9236 6822 9271 6830
rect 9236 6796 9237 6822
rect 9244 6796 9271 6822
rect 9179 6778 9209 6792
rect 9236 6788 9271 6796
rect 9236 6778 9237 6788
rect 9252 6778 9265 6788
rect -1 6772 9265 6778
rect 0 6764 9265 6772
rect 15 6734 28 6764
rect 43 6750 73 6764
rect 116 6750 159 6764
rect 166 6750 386 6764
rect 393 6750 423 6764
rect 83 6736 98 6748
rect 117 6736 130 6750
rect 198 6746 351 6750
rect 80 6734 102 6736
rect 180 6734 372 6746
rect 451 6734 464 6764
rect 479 6750 509 6764
rect 546 6734 565 6764
rect 580 6734 586 6764
rect 595 6734 608 6764
rect 623 6750 653 6764
rect 696 6750 739 6764
rect 746 6750 966 6764
rect 973 6750 1003 6764
rect 663 6736 678 6748
rect 697 6736 710 6750
rect 778 6746 931 6750
rect 660 6734 682 6736
rect 760 6734 952 6746
rect 1031 6734 1044 6764
rect 1059 6750 1089 6764
rect 1126 6734 1145 6764
rect 1160 6734 1166 6764
rect 1175 6734 1188 6764
rect 1203 6750 1233 6764
rect 1276 6750 1319 6764
rect 1326 6750 1546 6764
rect 1553 6750 1583 6764
rect 1243 6736 1258 6748
rect 1277 6736 1290 6750
rect 1358 6746 1511 6750
rect 1240 6734 1262 6736
rect 1340 6734 1532 6746
rect 1611 6734 1624 6764
rect 1639 6750 1669 6764
rect 1706 6734 1725 6764
rect 1740 6734 1746 6764
rect 1755 6734 1768 6764
rect 1783 6750 1813 6764
rect 1856 6750 1899 6764
rect 1906 6750 2126 6764
rect 2133 6750 2163 6764
rect 1823 6736 1838 6748
rect 1857 6736 1870 6750
rect 1938 6746 2091 6750
rect 1820 6734 1842 6736
rect 1920 6734 2112 6746
rect 2191 6734 2204 6764
rect 2219 6750 2249 6764
rect 2286 6734 2305 6764
rect 2320 6734 2326 6764
rect 2335 6734 2348 6764
rect 2363 6750 2393 6764
rect 2436 6750 2479 6764
rect 2486 6750 2706 6764
rect 2713 6750 2743 6764
rect 2403 6736 2418 6748
rect 2437 6736 2450 6750
rect 2518 6746 2671 6750
rect 2400 6734 2422 6736
rect 2500 6734 2692 6746
rect 2771 6734 2784 6764
rect 2799 6750 2829 6764
rect 2866 6734 2885 6764
rect 2900 6734 2906 6764
rect 2915 6734 2928 6764
rect 2943 6750 2973 6764
rect 3016 6750 3059 6764
rect 3066 6750 3286 6764
rect 3293 6750 3323 6764
rect 2983 6736 2998 6748
rect 3017 6736 3030 6750
rect 3098 6746 3251 6750
rect 2980 6734 3002 6736
rect 3080 6734 3272 6746
rect 3351 6734 3364 6764
rect 3379 6750 3409 6764
rect 3446 6734 3465 6764
rect 3480 6734 3486 6764
rect 3495 6734 3508 6764
rect 3523 6750 3553 6764
rect 3596 6750 3639 6764
rect 3646 6750 3866 6764
rect 3873 6750 3903 6764
rect 3563 6736 3578 6748
rect 3597 6736 3610 6750
rect 3678 6746 3831 6750
rect 3560 6734 3582 6736
rect 3660 6734 3852 6746
rect 3931 6734 3944 6764
rect 3959 6750 3989 6764
rect 4026 6734 4045 6764
rect 4060 6734 4066 6764
rect 4075 6734 4088 6764
rect 4103 6750 4133 6764
rect 4176 6750 4219 6764
rect 4226 6750 4446 6764
rect 4453 6750 4483 6764
rect 4143 6736 4158 6748
rect 4177 6736 4190 6750
rect 4258 6746 4411 6750
rect 4140 6734 4162 6736
rect 4240 6734 4432 6746
rect 4511 6734 4524 6764
rect 4539 6750 4569 6764
rect 4606 6734 4625 6764
rect 4640 6734 4646 6764
rect 4655 6734 4668 6764
rect 4683 6750 4713 6764
rect 4756 6750 4799 6764
rect 4806 6750 5026 6764
rect 5033 6750 5063 6764
rect 4723 6736 4738 6748
rect 4757 6736 4770 6750
rect 4838 6746 4991 6750
rect 4720 6734 4742 6736
rect 4820 6734 5012 6746
rect 5091 6734 5104 6764
rect 5119 6750 5149 6764
rect 5186 6734 5205 6764
rect 5220 6734 5226 6764
rect 5235 6734 5248 6764
rect 5263 6750 5293 6764
rect 5336 6750 5379 6764
rect 5386 6750 5606 6764
rect 5613 6750 5643 6764
rect 5303 6736 5318 6748
rect 5337 6736 5350 6750
rect 5418 6746 5571 6750
rect 5300 6734 5322 6736
rect 5400 6734 5592 6746
rect 5671 6734 5684 6764
rect 5699 6750 5729 6764
rect 5766 6734 5785 6764
rect 5800 6734 5806 6764
rect 5815 6734 5828 6764
rect 5843 6750 5873 6764
rect 5916 6750 5959 6764
rect 5966 6750 6186 6764
rect 6193 6750 6223 6764
rect 5883 6736 5898 6748
rect 5917 6736 5930 6750
rect 5998 6746 6151 6750
rect 5880 6734 5902 6736
rect 5980 6734 6172 6746
rect 6251 6734 6264 6764
rect 6279 6750 6309 6764
rect 6346 6734 6365 6764
rect 6380 6734 6386 6764
rect 6395 6734 6408 6764
rect 6423 6750 6453 6764
rect 6496 6750 6539 6764
rect 6546 6750 6766 6764
rect 6773 6750 6803 6764
rect 6463 6736 6478 6748
rect 6497 6736 6510 6750
rect 6578 6746 6731 6750
rect 6460 6734 6482 6736
rect 6560 6734 6752 6746
rect 6831 6734 6844 6764
rect 6859 6750 6889 6764
rect 6926 6734 6945 6764
rect 6960 6734 6966 6764
rect 6975 6734 6988 6764
rect 7003 6750 7033 6764
rect 7076 6750 7119 6764
rect 7126 6750 7346 6764
rect 7353 6750 7383 6764
rect 7043 6736 7058 6748
rect 7077 6736 7090 6750
rect 7158 6746 7311 6750
rect 7040 6734 7062 6736
rect 7140 6734 7332 6746
rect 7411 6734 7424 6764
rect 7439 6750 7469 6764
rect 7506 6734 7525 6764
rect 7540 6734 7546 6764
rect 7555 6734 7568 6764
rect 7583 6746 7613 6764
rect 7656 6750 7670 6764
rect 7706 6750 7926 6764
rect 7657 6748 7670 6750
rect 7623 6736 7638 6748
rect 7620 6734 7642 6736
rect 7647 6734 7677 6748
rect 7738 6746 7891 6750
rect 7720 6734 7912 6746
rect 7955 6734 7985 6748
rect 7991 6734 8004 6764
rect 8019 6746 8049 6764
rect 8092 6734 8105 6764
rect 8135 6734 8148 6764
rect 8163 6746 8193 6764
rect 8236 6750 8250 6764
rect 8286 6750 8506 6764
rect 8237 6748 8250 6750
rect 8203 6736 8218 6748
rect 8200 6734 8222 6736
rect 8227 6734 8257 6748
rect 8318 6746 8471 6750
rect 8300 6734 8492 6746
rect 8535 6734 8565 6748
rect 8571 6734 8584 6764
rect 8599 6746 8629 6764
rect 8672 6734 8685 6764
rect 8715 6734 8728 6764
rect 8743 6746 8773 6764
rect 8816 6750 8830 6764
rect 8866 6750 9086 6764
rect 8817 6748 8830 6750
rect 8783 6736 8798 6748
rect 8780 6734 8802 6736
rect 8807 6734 8837 6748
rect 8898 6746 9051 6750
rect 8880 6734 9072 6746
rect 9115 6734 9145 6748
rect 9151 6734 9164 6764
rect 9179 6746 9209 6764
rect 9252 6734 9265 6764
rect 0 6720 9265 6734
rect 15 6650 28 6720
rect 80 6716 102 6720
rect 73 6694 102 6708
rect 155 6694 171 6708
rect 209 6704 215 6706
rect 222 6704 330 6720
rect 337 6704 343 6706
rect 351 6704 366 6720
rect 432 6714 451 6717
rect 73 6692 171 6694
rect 198 6692 366 6704
rect 381 6694 397 6708
rect 432 6695 454 6714
rect 464 6708 480 6709
rect 463 6706 480 6708
rect 464 6701 480 6706
rect 454 6694 460 6695
rect 463 6694 492 6701
rect 381 6693 492 6694
rect 381 6692 498 6693
rect 57 6684 108 6692
rect 155 6684 189 6692
rect 57 6672 82 6684
rect 89 6672 108 6684
rect 162 6682 189 6684
rect 198 6682 419 6692
rect 454 6689 460 6692
rect 162 6678 419 6682
rect 57 6664 108 6672
rect 155 6664 419 6678
rect 463 6684 498 6692
rect 9 6616 28 6650
rect 73 6656 102 6664
rect 73 6650 90 6656
rect 73 6648 107 6650
rect 155 6648 171 6664
rect 172 6654 380 6664
rect 381 6654 397 6664
rect 445 6660 460 6675
rect 463 6672 464 6684
rect 471 6672 498 6684
rect 463 6664 498 6672
rect 463 6663 492 6664
rect 183 6650 397 6654
rect 198 6648 397 6650
rect 432 6650 445 6660
rect 463 6650 480 6663
rect 432 6648 480 6650
rect 74 6644 107 6648
rect 70 6642 107 6644
rect 70 6641 137 6642
rect 70 6636 101 6641
rect 107 6636 137 6641
rect 70 6632 137 6636
rect 43 6629 137 6632
rect 43 6622 92 6629
rect 43 6616 73 6622
rect 92 6617 97 6622
rect 9 6600 89 6616
rect 101 6608 137 6629
rect 198 6624 387 6648
rect 432 6647 479 6648
rect 445 6642 479 6647
rect 213 6621 387 6624
rect 206 6618 387 6621
rect 415 6641 479 6642
rect 9 6598 28 6600
rect 43 6598 77 6600
rect 9 6582 89 6598
rect 9 6576 28 6582
rect -1 6560 28 6576
rect 43 6566 73 6582
rect 101 6560 107 6608
rect 110 6602 129 6608
rect 144 6602 174 6610
rect 110 6594 174 6602
rect 110 6578 190 6594
rect 206 6587 268 6618
rect 284 6587 346 6618
rect 415 6616 464 6641
rect 479 6616 509 6632
rect 378 6602 408 6610
rect 415 6608 525 6616
rect 378 6594 423 6602
rect 110 6576 129 6578
rect 144 6576 190 6578
rect 110 6560 190 6576
rect 217 6574 252 6587
rect 293 6584 330 6587
rect 293 6582 335 6584
rect 222 6571 252 6574
rect 231 6567 238 6571
rect 238 6566 239 6567
rect 197 6560 207 6566
rect -7 6552 34 6560
rect -7 6526 8 6552
rect 15 6526 34 6552
rect 98 6548 129 6560
rect 144 6548 247 6560
rect 259 6550 285 6576
rect 300 6571 330 6582
rect 362 6578 424 6594
rect 362 6576 408 6578
rect 362 6560 424 6576
rect 436 6560 442 6608
rect 445 6600 525 6608
rect 445 6598 464 6600
rect 479 6598 513 6600
rect 445 6582 525 6598
rect 445 6560 464 6582
rect 479 6566 509 6582
rect 537 6576 543 6650
rect 546 6576 565 6720
rect 580 6576 586 6720
rect 595 6650 608 6720
rect 660 6716 682 6720
rect 653 6694 682 6708
rect 735 6694 751 6708
rect 789 6704 795 6706
rect 802 6704 910 6720
rect 917 6704 923 6706
rect 931 6704 946 6720
rect 1012 6714 1031 6717
rect 653 6692 751 6694
rect 778 6692 946 6704
rect 961 6694 977 6708
rect 1012 6695 1034 6714
rect 1044 6708 1060 6709
rect 1043 6706 1060 6708
rect 1044 6701 1060 6706
rect 1034 6694 1040 6695
rect 1043 6694 1072 6701
rect 961 6693 1072 6694
rect 961 6692 1078 6693
rect 637 6684 688 6692
rect 735 6684 769 6692
rect 637 6672 662 6684
rect 669 6672 688 6684
rect 742 6682 769 6684
rect 778 6682 999 6692
rect 1034 6689 1040 6692
rect 742 6678 999 6682
rect 637 6664 688 6672
rect 735 6664 999 6678
rect 1043 6684 1078 6692
rect 589 6616 608 6650
rect 653 6656 682 6664
rect 653 6650 670 6656
rect 653 6648 687 6650
rect 735 6648 751 6664
rect 752 6654 960 6664
rect 961 6654 977 6664
rect 1025 6660 1040 6675
rect 1043 6672 1044 6684
rect 1051 6672 1078 6684
rect 1043 6664 1078 6672
rect 1043 6663 1072 6664
rect 763 6650 977 6654
rect 778 6648 977 6650
rect 1012 6650 1025 6660
rect 1043 6650 1060 6663
rect 1012 6648 1060 6650
rect 654 6644 687 6648
rect 650 6642 687 6644
rect 650 6641 717 6642
rect 650 6636 681 6641
rect 687 6636 717 6641
rect 650 6632 717 6636
rect 623 6629 717 6632
rect 623 6622 672 6629
rect 623 6616 653 6622
rect 672 6617 677 6622
rect 589 6600 669 6616
rect 681 6608 717 6629
rect 778 6624 967 6648
rect 1012 6647 1059 6648
rect 1025 6642 1059 6647
rect 793 6621 967 6624
rect 786 6618 967 6621
rect 995 6641 1059 6642
rect 589 6598 608 6600
rect 623 6598 657 6600
rect 589 6582 669 6598
rect 589 6576 608 6582
rect 305 6550 408 6560
rect 259 6548 408 6550
rect 429 6548 464 6560
rect 98 6546 260 6548
rect 110 6526 129 6546
rect 144 6544 174 6546
rect -7 6518 34 6526
rect 116 6522 129 6526
rect 181 6530 260 6546
rect 292 6546 464 6548
rect 292 6530 371 6546
rect 378 6544 408 6546
rect -1 6508 28 6518
rect 43 6508 73 6522
rect 116 6508 159 6522
rect 181 6518 371 6530
rect 436 6526 442 6546
rect 166 6508 196 6518
rect 197 6508 355 6518
rect 359 6508 389 6518
rect 393 6508 423 6522
rect 451 6508 464 6546
rect 536 6560 565 6576
rect 579 6560 608 6576
rect 623 6566 653 6582
rect 681 6560 687 6608
rect 690 6602 709 6608
rect 724 6602 754 6610
rect 690 6594 754 6602
rect 690 6578 770 6594
rect 786 6587 848 6618
rect 864 6587 926 6618
rect 995 6616 1044 6641
rect 1059 6616 1089 6632
rect 958 6602 988 6610
rect 995 6608 1105 6616
rect 958 6594 1003 6602
rect 690 6576 709 6578
rect 724 6576 770 6578
rect 690 6560 770 6576
rect 797 6574 832 6587
rect 873 6584 910 6587
rect 873 6582 915 6584
rect 802 6571 832 6574
rect 811 6567 818 6571
rect 818 6566 819 6567
rect 777 6560 787 6566
rect 536 6552 571 6560
rect 536 6526 537 6552
rect 544 6526 571 6552
rect 479 6508 509 6522
rect 536 6518 571 6526
rect 573 6552 614 6560
rect 573 6526 588 6552
rect 595 6526 614 6552
rect 678 6548 709 6560
rect 724 6548 827 6560
rect 839 6550 865 6576
rect 880 6571 910 6582
rect 942 6578 1004 6594
rect 942 6576 988 6578
rect 942 6560 1004 6576
rect 1016 6560 1022 6608
rect 1025 6600 1105 6608
rect 1025 6598 1044 6600
rect 1059 6598 1093 6600
rect 1025 6582 1105 6598
rect 1025 6560 1044 6582
rect 1059 6566 1089 6582
rect 1117 6576 1123 6650
rect 1126 6576 1145 6720
rect 1160 6576 1166 6720
rect 1175 6650 1188 6720
rect 1240 6716 1262 6720
rect 1233 6694 1262 6708
rect 1315 6694 1331 6708
rect 1369 6704 1375 6706
rect 1382 6704 1490 6720
rect 1497 6704 1503 6706
rect 1511 6704 1526 6720
rect 1592 6714 1611 6717
rect 1233 6692 1331 6694
rect 1358 6692 1526 6704
rect 1541 6694 1557 6708
rect 1592 6695 1614 6714
rect 1624 6708 1640 6709
rect 1623 6706 1640 6708
rect 1624 6701 1640 6706
rect 1614 6694 1620 6695
rect 1623 6694 1652 6701
rect 1541 6693 1652 6694
rect 1541 6692 1658 6693
rect 1217 6684 1268 6692
rect 1315 6684 1349 6692
rect 1217 6672 1242 6684
rect 1249 6672 1268 6684
rect 1322 6682 1349 6684
rect 1358 6682 1579 6692
rect 1614 6689 1620 6692
rect 1322 6678 1579 6682
rect 1217 6664 1268 6672
rect 1315 6664 1579 6678
rect 1623 6684 1658 6692
rect 1169 6616 1188 6650
rect 1233 6656 1262 6664
rect 1233 6650 1250 6656
rect 1233 6648 1267 6650
rect 1315 6648 1331 6664
rect 1332 6654 1540 6664
rect 1541 6654 1557 6664
rect 1605 6660 1620 6675
rect 1623 6672 1624 6684
rect 1631 6672 1658 6684
rect 1623 6664 1658 6672
rect 1623 6663 1652 6664
rect 1343 6650 1557 6654
rect 1358 6648 1557 6650
rect 1592 6650 1605 6660
rect 1623 6650 1640 6663
rect 1592 6648 1640 6650
rect 1234 6644 1267 6648
rect 1230 6642 1267 6644
rect 1230 6641 1297 6642
rect 1230 6636 1261 6641
rect 1267 6636 1297 6641
rect 1230 6632 1297 6636
rect 1203 6629 1297 6632
rect 1203 6622 1252 6629
rect 1203 6616 1233 6622
rect 1252 6617 1257 6622
rect 1169 6600 1249 6616
rect 1261 6608 1297 6629
rect 1358 6624 1547 6648
rect 1592 6647 1639 6648
rect 1605 6642 1639 6647
rect 1373 6621 1547 6624
rect 1366 6618 1547 6621
rect 1575 6641 1639 6642
rect 1169 6598 1188 6600
rect 1203 6598 1237 6600
rect 1169 6582 1249 6598
rect 1169 6576 1188 6582
rect 885 6550 988 6560
rect 839 6548 988 6550
rect 1009 6548 1044 6560
rect 678 6546 840 6548
rect 690 6526 709 6546
rect 724 6544 754 6546
rect 573 6518 614 6526
rect 696 6522 709 6526
rect 761 6530 840 6546
rect 872 6546 1044 6548
rect 872 6530 951 6546
rect 958 6544 988 6546
rect 536 6508 565 6518
rect 579 6508 608 6518
rect 623 6508 653 6522
rect 696 6508 739 6522
rect 761 6518 951 6530
rect 1016 6526 1022 6546
rect 746 6508 776 6518
rect 777 6508 935 6518
rect 939 6508 969 6518
rect 973 6508 1003 6522
rect 1031 6508 1044 6546
rect 1116 6560 1145 6576
rect 1159 6560 1188 6576
rect 1203 6566 1233 6582
rect 1261 6560 1267 6608
rect 1270 6602 1289 6608
rect 1304 6602 1334 6610
rect 1270 6594 1334 6602
rect 1270 6578 1350 6594
rect 1366 6587 1428 6618
rect 1444 6587 1506 6618
rect 1575 6616 1624 6641
rect 1639 6616 1669 6632
rect 1538 6602 1568 6610
rect 1575 6608 1685 6616
rect 1538 6594 1583 6602
rect 1270 6576 1289 6578
rect 1304 6576 1350 6578
rect 1270 6560 1350 6576
rect 1377 6574 1412 6587
rect 1453 6584 1490 6587
rect 1453 6582 1495 6584
rect 1382 6571 1412 6574
rect 1391 6567 1398 6571
rect 1398 6566 1399 6567
rect 1357 6560 1367 6566
rect 1116 6552 1151 6560
rect 1116 6526 1117 6552
rect 1124 6526 1151 6552
rect 1059 6508 1089 6522
rect 1116 6518 1151 6526
rect 1153 6552 1194 6560
rect 1153 6526 1168 6552
rect 1175 6526 1194 6552
rect 1258 6548 1289 6560
rect 1304 6548 1407 6560
rect 1419 6550 1445 6576
rect 1460 6571 1490 6582
rect 1522 6578 1584 6594
rect 1522 6576 1568 6578
rect 1522 6560 1584 6576
rect 1596 6560 1602 6608
rect 1605 6600 1685 6608
rect 1605 6598 1624 6600
rect 1639 6598 1673 6600
rect 1605 6582 1685 6598
rect 1605 6560 1624 6582
rect 1639 6566 1669 6582
rect 1697 6576 1703 6650
rect 1706 6576 1725 6720
rect 1740 6576 1746 6720
rect 1755 6650 1768 6720
rect 1820 6716 1842 6720
rect 1813 6694 1842 6708
rect 1895 6694 1911 6708
rect 1949 6704 1955 6706
rect 1962 6704 2070 6720
rect 2077 6704 2083 6706
rect 2091 6704 2106 6720
rect 2172 6714 2191 6717
rect 1813 6692 1911 6694
rect 1938 6692 2106 6704
rect 2121 6694 2137 6708
rect 2172 6695 2194 6714
rect 2204 6708 2220 6709
rect 2203 6706 2220 6708
rect 2204 6701 2220 6706
rect 2194 6694 2200 6695
rect 2203 6694 2232 6701
rect 2121 6693 2232 6694
rect 2121 6692 2238 6693
rect 1797 6684 1848 6692
rect 1895 6684 1929 6692
rect 1797 6672 1822 6684
rect 1829 6672 1848 6684
rect 1902 6682 1929 6684
rect 1938 6682 2159 6692
rect 2194 6689 2200 6692
rect 1902 6678 2159 6682
rect 1797 6664 1848 6672
rect 1895 6664 2159 6678
rect 2203 6684 2238 6692
rect 1749 6616 1768 6650
rect 1813 6656 1842 6664
rect 1813 6650 1830 6656
rect 1813 6648 1847 6650
rect 1895 6648 1911 6664
rect 1912 6654 2120 6664
rect 2121 6654 2137 6664
rect 2185 6660 2200 6675
rect 2203 6672 2204 6684
rect 2211 6672 2238 6684
rect 2203 6664 2238 6672
rect 2203 6663 2232 6664
rect 1923 6650 2137 6654
rect 1938 6648 2137 6650
rect 2172 6650 2185 6660
rect 2203 6650 2220 6663
rect 2172 6648 2220 6650
rect 1814 6644 1847 6648
rect 1810 6642 1847 6644
rect 1810 6641 1877 6642
rect 1810 6636 1841 6641
rect 1847 6636 1877 6641
rect 1810 6632 1877 6636
rect 1783 6629 1877 6632
rect 1783 6622 1832 6629
rect 1783 6616 1813 6622
rect 1832 6617 1837 6622
rect 1749 6600 1829 6616
rect 1841 6608 1877 6629
rect 1938 6624 2127 6648
rect 2172 6647 2219 6648
rect 2185 6642 2219 6647
rect 1953 6621 2127 6624
rect 1946 6618 2127 6621
rect 2155 6641 2219 6642
rect 1749 6598 1768 6600
rect 1783 6598 1817 6600
rect 1749 6582 1829 6598
rect 1749 6576 1768 6582
rect 1465 6550 1568 6560
rect 1419 6548 1568 6550
rect 1589 6548 1624 6560
rect 1258 6546 1420 6548
rect 1270 6526 1289 6546
rect 1304 6544 1334 6546
rect 1153 6518 1194 6526
rect 1276 6522 1289 6526
rect 1341 6530 1420 6546
rect 1452 6546 1624 6548
rect 1452 6530 1531 6546
rect 1538 6544 1568 6546
rect 1116 6508 1145 6518
rect 1159 6508 1188 6518
rect 1203 6508 1233 6522
rect 1276 6508 1319 6522
rect 1341 6518 1531 6530
rect 1596 6526 1602 6546
rect 1326 6508 1356 6518
rect 1357 6508 1515 6518
rect 1519 6508 1549 6518
rect 1553 6508 1583 6522
rect 1611 6508 1624 6546
rect 1696 6560 1725 6576
rect 1739 6560 1768 6576
rect 1783 6566 1813 6582
rect 1841 6560 1847 6608
rect 1850 6602 1869 6608
rect 1884 6602 1914 6610
rect 1850 6594 1914 6602
rect 1850 6578 1930 6594
rect 1946 6587 2008 6618
rect 2024 6587 2086 6618
rect 2155 6616 2204 6641
rect 2219 6616 2249 6632
rect 2118 6602 2148 6610
rect 2155 6608 2265 6616
rect 2118 6594 2163 6602
rect 1850 6576 1869 6578
rect 1884 6576 1930 6578
rect 1850 6560 1930 6576
rect 1957 6574 1992 6587
rect 2033 6584 2070 6587
rect 2033 6582 2075 6584
rect 1962 6571 1992 6574
rect 1971 6567 1978 6571
rect 1978 6566 1979 6567
rect 1937 6560 1947 6566
rect 1696 6552 1731 6560
rect 1696 6526 1697 6552
rect 1704 6526 1731 6552
rect 1639 6508 1669 6522
rect 1696 6518 1731 6526
rect 1733 6552 1774 6560
rect 1733 6526 1748 6552
rect 1755 6526 1774 6552
rect 1838 6548 1869 6560
rect 1884 6548 1987 6560
rect 1999 6550 2025 6576
rect 2040 6571 2070 6582
rect 2102 6578 2164 6594
rect 2102 6576 2148 6578
rect 2102 6560 2164 6576
rect 2176 6560 2182 6608
rect 2185 6600 2265 6608
rect 2185 6598 2204 6600
rect 2219 6598 2253 6600
rect 2185 6582 2265 6598
rect 2185 6560 2204 6582
rect 2219 6566 2249 6582
rect 2277 6576 2283 6650
rect 2286 6576 2305 6720
rect 2320 6576 2326 6720
rect 2335 6650 2348 6720
rect 2400 6716 2422 6720
rect 2393 6694 2422 6708
rect 2475 6694 2491 6708
rect 2529 6704 2535 6706
rect 2542 6704 2650 6720
rect 2657 6704 2663 6706
rect 2671 6704 2686 6720
rect 2752 6714 2771 6717
rect 2393 6692 2491 6694
rect 2518 6692 2686 6704
rect 2701 6694 2717 6708
rect 2752 6695 2774 6714
rect 2784 6708 2800 6709
rect 2783 6706 2800 6708
rect 2784 6701 2800 6706
rect 2774 6694 2780 6695
rect 2783 6694 2812 6701
rect 2701 6693 2812 6694
rect 2701 6692 2818 6693
rect 2377 6684 2428 6692
rect 2475 6684 2509 6692
rect 2377 6672 2402 6684
rect 2409 6672 2428 6684
rect 2482 6682 2509 6684
rect 2518 6682 2739 6692
rect 2774 6689 2780 6692
rect 2482 6678 2739 6682
rect 2377 6664 2428 6672
rect 2475 6664 2739 6678
rect 2783 6684 2818 6692
rect 2329 6616 2348 6650
rect 2393 6656 2422 6664
rect 2393 6650 2410 6656
rect 2393 6648 2427 6650
rect 2475 6648 2491 6664
rect 2492 6654 2700 6664
rect 2701 6654 2717 6664
rect 2765 6660 2780 6675
rect 2783 6672 2784 6684
rect 2791 6672 2818 6684
rect 2783 6664 2818 6672
rect 2783 6663 2812 6664
rect 2503 6650 2717 6654
rect 2518 6648 2717 6650
rect 2752 6650 2765 6660
rect 2783 6650 2800 6663
rect 2752 6648 2800 6650
rect 2394 6644 2427 6648
rect 2390 6642 2427 6644
rect 2390 6641 2457 6642
rect 2390 6636 2421 6641
rect 2427 6636 2457 6641
rect 2390 6632 2457 6636
rect 2363 6629 2457 6632
rect 2363 6622 2412 6629
rect 2363 6616 2393 6622
rect 2412 6617 2417 6622
rect 2329 6600 2409 6616
rect 2421 6608 2457 6629
rect 2518 6624 2707 6648
rect 2752 6647 2799 6648
rect 2765 6642 2799 6647
rect 2533 6621 2707 6624
rect 2526 6618 2707 6621
rect 2735 6641 2799 6642
rect 2329 6598 2348 6600
rect 2363 6598 2397 6600
rect 2329 6582 2409 6598
rect 2329 6576 2348 6582
rect 2045 6550 2148 6560
rect 1999 6548 2148 6550
rect 2169 6548 2204 6560
rect 1838 6546 2000 6548
rect 1850 6526 1869 6546
rect 1884 6544 1914 6546
rect 1733 6518 1774 6526
rect 1856 6522 1869 6526
rect 1921 6530 2000 6546
rect 2032 6546 2204 6548
rect 2032 6530 2111 6546
rect 2118 6544 2148 6546
rect 1696 6508 1725 6518
rect 1739 6508 1768 6518
rect 1783 6508 1813 6522
rect 1856 6508 1899 6522
rect 1921 6518 2111 6530
rect 2176 6526 2182 6546
rect 1906 6508 1936 6518
rect 1937 6508 2095 6518
rect 2099 6508 2129 6518
rect 2133 6508 2163 6522
rect 2191 6508 2204 6546
rect 2276 6560 2305 6576
rect 2319 6560 2348 6576
rect 2363 6566 2393 6582
rect 2421 6560 2427 6608
rect 2430 6602 2449 6608
rect 2464 6602 2494 6610
rect 2430 6594 2494 6602
rect 2430 6578 2510 6594
rect 2526 6587 2588 6618
rect 2604 6587 2666 6618
rect 2735 6616 2784 6641
rect 2799 6616 2829 6632
rect 2698 6602 2728 6610
rect 2735 6608 2845 6616
rect 2698 6594 2743 6602
rect 2430 6576 2449 6578
rect 2464 6576 2510 6578
rect 2430 6560 2510 6576
rect 2537 6574 2572 6587
rect 2613 6584 2650 6587
rect 2613 6582 2655 6584
rect 2542 6571 2572 6574
rect 2551 6567 2558 6571
rect 2558 6566 2559 6567
rect 2517 6560 2527 6566
rect 2276 6552 2311 6560
rect 2276 6526 2277 6552
rect 2284 6526 2311 6552
rect 2219 6508 2249 6522
rect 2276 6518 2311 6526
rect 2313 6552 2354 6560
rect 2313 6526 2328 6552
rect 2335 6526 2354 6552
rect 2418 6548 2449 6560
rect 2464 6548 2567 6560
rect 2579 6550 2605 6576
rect 2620 6571 2650 6582
rect 2682 6578 2744 6594
rect 2682 6576 2728 6578
rect 2682 6560 2744 6576
rect 2756 6560 2762 6608
rect 2765 6600 2845 6608
rect 2765 6598 2784 6600
rect 2799 6598 2833 6600
rect 2765 6582 2845 6598
rect 2765 6560 2784 6582
rect 2799 6566 2829 6582
rect 2857 6576 2863 6650
rect 2866 6576 2885 6720
rect 2900 6576 2906 6720
rect 2915 6650 2928 6720
rect 2980 6716 3002 6720
rect 2973 6694 3002 6708
rect 3055 6694 3071 6708
rect 3109 6704 3115 6706
rect 3122 6704 3230 6720
rect 3237 6704 3243 6706
rect 3251 6704 3266 6720
rect 3332 6714 3351 6717
rect 2973 6692 3071 6694
rect 3098 6692 3266 6704
rect 3281 6694 3297 6708
rect 3332 6695 3354 6714
rect 3364 6708 3380 6709
rect 3363 6706 3380 6708
rect 3364 6701 3380 6706
rect 3354 6694 3360 6695
rect 3363 6694 3392 6701
rect 3281 6693 3392 6694
rect 3281 6692 3398 6693
rect 2957 6684 3008 6692
rect 3055 6684 3089 6692
rect 2957 6672 2982 6684
rect 2989 6672 3008 6684
rect 3062 6682 3089 6684
rect 3098 6682 3319 6692
rect 3354 6689 3360 6692
rect 3062 6678 3319 6682
rect 2957 6664 3008 6672
rect 3055 6664 3319 6678
rect 3363 6684 3398 6692
rect 2909 6616 2928 6650
rect 2973 6656 3002 6664
rect 2973 6650 2990 6656
rect 2973 6648 3007 6650
rect 3055 6648 3071 6664
rect 3072 6654 3280 6664
rect 3281 6654 3297 6664
rect 3345 6660 3360 6675
rect 3363 6672 3364 6684
rect 3371 6672 3398 6684
rect 3363 6664 3398 6672
rect 3363 6663 3392 6664
rect 3083 6650 3297 6654
rect 3098 6648 3297 6650
rect 3332 6650 3345 6660
rect 3363 6650 3380 6663
rect 3332 6648 3380 6650
rect 2974 6644 3007 6648
rect 2970 6642 3007 6644
rect 2970 6641 3037 6642
rect 2970 6636 3001 6641
rect 3007 6636 3037 6641
rect 2970 6632 3037 6636
rect 2943 6629 3037 6632
rect 2943 6622 2992 6629
rect 2943 6616 2973 6622
rect 2992 6617 2997 6622
rect 2909 6600 2989 6616
rect 3001 6608 3037 6629
rect 3098 6624 3287 6648
rect 3332 6647 3379 6648
rect 3345 6642 3379 6647
rect 3113 6621 3287 6624
rect 3106 6618 3287 6621
rect 3315 6641 3379 6642
rect 2909 6598 2928 6600
rect 2943 6598 2977 6600
rect 2909 6582 2989 6598
rect 2909 6576 2928 6582
rect 2625 6550 2728 6560
rect 2579 6548 2728 6550
rect 2749 6548 2784 6560
rect 2418 6546 2580 6548
rect 2430 6526 2449 6546
rect 2464 6544 2494 6546
rect 2313 6518 2354 6526
rect 2436 6522 2449 6526
rect 2501 6530 2580 6546
rect 2612 6546 2784 6548
rect 2612 6530 2691 6546
rect 2698 6544 2728 6546
rect 2276 6508 2305 6518
rect 2319 6508 2348 6518
rect 2363 6508 2393 6522
rect 2436 6508 2479 6522
rect 2501 6518 2691 6530
rect 2756 6526 2762 6546
rect 2486 6508 2516 6518
rect 2517 6508 2675 6518
rect 2679 6508 2709 6518
rect 2713 6508 2743 6522
rect 2771 6508 2784 6546
rect 2856 6560 2885 6576
rect 2899 6560 2928 6576
rect 2943 6566 2973 6582
rect 3001 6560 3007 6608
rect 3010 6602 3029 6608
rect 3044 6602 3074 6610
rect 3010 6594 3074 6602
rect 3010 6578 3090 6594
rect 3106 6587 3168 6618
rect 3184 6587 3246 6618
rect 3315 6616 3364 6641
rect 3379 6616 3409 6632
rect 3278 6602 3308 6610
rect 3315 6608 3425 6616
rect 3278 6594 3323 6602
rect 3010 6576 3029 6578
rect 3044 6576 3090 6578
rect 3010 6560 3090 6576
rect 3117 6574 3152 6587
rect 3193 6584 3230 6587
rect 3193 6582 3235 6584
rect 3122 6571 3152 6574
rect 3131 6567 3138 6571
rect 3138 6566 3139 6567
rect 3097 6560 3107 6566
rect 2856 6552 2891 6560
rect 2856 6526 2857 6552
rect 2864 6526 2891 6552
rect 2799 6508 2829 6522
rect 2856 6518 2891 6526
rect 2893 6552 2934 6560
rect 2893 6526 2908 6552
rect 2915 6526 2934 6552
rect 2998 6548 3029 6560
rect 3044 6548 3147 6560
rect 3159 6550 3185 6576
rect 3200 6571 3230 6582
rect 3262 6578 3324 6594
rect 3262 6576 3308 6578
rect 3262 6560 3324 6576
rect 3336 6560 3342 6608
rect 3345 6600 3425 6608
rect 3345 6598 3364 6600
rect 3379 6598 3413 6600
rect 3345 6582 3425 6598
rect 3345 6560 3364 6582
rect 3379 6566 3409 6582
rect 3437 6576 3443 6650
rect 3446 6576 3465 6720
rect 3480 6576 3486 6720
rect 3495 6650 3508 6720
rect 3560 6716 3582 6720
rect 3553 6694 3582 6708
rect 3635 6694 3651 6708
rect 3689 6704 3695 6706
rect 3702 6704 3810 6720
rect 3817 6704 3823 6706
rect 3831 6704 3846 6720
rect 3912 6714 3931 6717
rect 3553 6692 3651 6694
rect 3678 6692 3846 6704
rect 3861 6694 3877 6708
rect 3912 6695 3934 6714
rect 3944 6708 3960 6709
rect 3943 6706 3960 6708
rect 3944 6701 3960 6706
rect 3934 6694 3940 6695
rect 3943 6694 3972 6701
rect 3861 6693 3972 6694
rect 3861 6692 3978 6693
rect 3537 6684 3588 6692
rect 3635 6684 3669 6692
rect 3537 6672 3562 6684
rect 3569 6672 3588 6684
rect 3642 6682 3669 6684
rect 3678 6682 3899 6692
rect 3934 6689 3940 6692
rect 3642 6678 3899 6682
rect 3537 6664 3588 6672
rect 3635 6664 3899 6678
rect 3943 6684 3978 6692
rect 3489 6616 3508 6650
rect 3553 6656 3582 6664
rect 3553 6650 3570 6656
rect 3553 6648 3587 6650
rect 3635 6648 3651 6664
rect 3652 6654 3860 6664
rect 3861 6654 3877 6664
rect 3925 6660 3940 6675
rect 3943 6672 3944 6684
rect 3951 6672 3978 6684
rect 3943 6664 3978 6672
rect 3943 6663 3972 6664
rect 3663 6650 3877 6654
rect 3678 6648 3877 6650
rect 3912 6650 3925 6660
rect 3943 6650 3960 6663
rect 3912 6648 3960 6650
rect 3554 6644 3587 6648
rect 3550 6642 3587 6644
rect 3550 6641 3617 6642
rect 3550 6636 3581 6641
rect 3587 6636 3617 6641
rect 3550 6632 3617 6636
rect 3523 6629 3617 6632
rect 3523 6622 3572 6629
rect 3523 6616 3553 6622
rect 3572 6617 3577 6622
rect 3489 6600 3569 6616
rect 3581 6608 3617 6629
rect 3678 6624 3867 6648
rect 3912 6647 3959 6648
rect 3925 6642 3959 6647
rect 3693 6621 3867 6624
rect 3686 6618 3867 6621
rect 3895 6641 3959 6642
rect 3489 6598 3508 6600
rect 3523 6598 3557 6600
rect 3489 6582 3569 6598
rect 3489 6576 3508 6582
rect 3205 6550 3308 6560
rect 3159 6548 3308 6550
rect 3329 6548 3364 6560
rect 2998 6546 3160 6548
rect 3010 6526 3029 6546
rect 3044 6544 3074 6546
rect 2893 6518 2934 6526
rect 3016 6522 3029 6526
rect 3081 6530 3160 6546
rect 3192 6546 3364 6548
rect 3192 6530 3271 6546
rect 3278 6544 3308 6546
rect 2856 6508 2885 6518
rect 2899 6508 2928 6518
rect 2943 6508 2973 6522
rect 3016 6508 3059 6522
rect 3081 6518 3271 6530
rect 3336 6526 3342 6546
rect 3066 6508 3096 6518
rect 3097 6508 3255 6518
rect 3259 6508 3289 6518
rect 3293 6508 3323 6522
rect 3351 6508 3364 6546
rect 3436 6560 3465 6576
rect 3479 6560 3508 6576
rect 3523 6566 3553 6582
rect 3581 6560 3587 6608
rect 3590 6602 3609 6608
rect 3624 6602 3654 6610
rect 3590 6594 3654 6602
rect 3590 6578 3670 6594
rect 3686 6587 3748 6618
rect 3764 6587 3826 6618
rect 3895 6616 3944 6641
rect 3959 6616 3989 6632
rect 3858 6602 3888 6610
rect 3895 6608 4005 6616
rect 3858 6594 3903 6602
rect 3590 6576 3609 6578
rect 3624 6576 3670 6578
rect 3590 6560 3670 6576
rect 3697 6574 3732 6587
rect 3773 6584 3810 6587
rect 3773 6582 3815 6584
rect 3702 6571 3732 6574
rect 3711 6567 3718 6571
rect 3718 6566 3719 6567
rect 3677 6560 3687 6566
rect 3436 6552 3471 6560
rect 3436 6526 3437 6552
rect 3444 6526 3471 6552
rect 3379 6508 3409 6522
rect 3436 6518 3471 6526
rect 3473 6552 3514 6560
rect 3473 6526 3488 6552
rect 3495 6526 3514 6552
rect 3578 6548 3609 6560
rect 3624 6548 3727 6560
rect 3739 6550 3765 6576
rect 3780 6571 3810 6582
rect 3842 6578 3904 6594
rect 3842 6576 3888 6578
rect 3842 6560 3904 6576
rect 3916 6560 3922 6608
rect 3925 6600 4005 6608
rect 3925 6598 3944 6600
rect 3959 6598 3993 6600
rect 3925 6582 4005 6598
rect 3925 6560 3944 6582
rect 3959 6566 3989 6582
rect 4017 6576 4023 6650
rect 4026 6576 4045 6720
rect 4060 6576 4066 6720
rect 4075 6650 4088 6720
rect 4140 6716 4162 6720
rect 4133 6694 4162 6708
rect 4215 6694 4231 6708
rect 4269 6704 4275 6706
rect 4282 6704 4390 6720
rect 4397 6704 4403 6706
rect 4411 6704 4426 6720
rect 4492 6714 4511 6717
rect 4133 6692 4231 6694
rect 4258 6692 4426 6704
rect 4441 6694 4457 6708
rect 4492 6695 4514 6714
rect 4524 6708 4540 6709
rect 4523 6706 4540 6708
rect 4524 6701 4540 6706
rect 4514 6694 4520 6695
rect 4523 6694 4552 6701
rect 4441 6693 4552 6694
rect 4441 6692 4558 6693
rect 4117 6684 4168 6692
rect 4215 6684 4249 6692
rect 4117 6672 4142 6684
rect 4149 6672 4168 6684
rect 4222 6682 4249 6684
rect 4258 6682 4479 6692
rect 4514 6689 4520 6692
rect 4222 6678 4479 6682
rect 4117 6664 4168 6672
rect 4215 6664 4479 6678
rect 4523 6684 4558 6692
rect 4069 6616 4088 6650
rect 4133 6656 4162 6664
rect 4133 6650 4150 6656
rect 4133 6648 4167 6650
rect 4215 6648 4231 6664
rect 4232 6654 4440 6664
rect 4441 6654 4457 6664
rect 4505 6660 4520 6675
rect 4523 6672 4524 6684
rect 4531 6672 4558 6684
rect 4523 6664 4558 6672
rect 4523 6663 4552 6664
rect 4243 6650 4457 6654
rect 4258 6648 4457 6650
rect 4492 6650 4505 6660
rect 4523 6650 4540 6663
rect 4492 6648 4540 6650
rect 4134 6644 4167 6648
rect 4130 6642 4167 6644
rect 4130 6641 4197 6642
rect 4130 6636 4161 6641
rect 4167 6636 4197 6641
rect 4130 6632 4197 6636
rect 4103 6629 4197 6632
rect 4103 6622 4152 6629
rect 4103 6616 4133 6622
rect 4152 6617 4157 6622
rect 4069 6600 4149 6616
rect 4161 6608 4197 6629
rect 4258 6624 4447 6648
rect 4492 6647 4539 6648
rect 4505 6642 4539 6647
rect 4273 6621 4447 6624
rect 4266 6618 4447 6621
rect 4475 6641 4539 6642
rect 4069 6598 4088 6600
rect 4103 6598 4137 6600
rect 4069 6582 4149 6598
rect 4069 6576 4088 6582
rect 3785 6550 3888 6560
rect 3739 6548 3888 6550
rect 3909 6548 3944 6560
rect 3578 6546 3740 6548
rect 3590 6526 3609 6546
rect 3624 6544 3654 6546
rect 3473 6518 3514 6526
rect 3596 6522 3609 6526
rect 3661 6530 3740 6546
rect 3772 6546 3944 6548
rect 3772 6530 3851 6546
rect 3858 6544 3888 6546
rect 3436 6508 3465 6518
rect 3479 6508 3508 6518
rect 3523 6508 3553 6522
rect 3596 6508 3639 6522
rect 3661 6518 3851 6530
rect 3916 6526 3922 6546
rect 3646 6508 3676 6518
rect 3677 6508 3835 6518
rect 3839 6508 3869 6518
rect 3873 6508 3903 6522
rect 3931 6508 3944 6546
rect 4016 6560 4045 6576
rect 4059 6560 4088 6576
rect 4103 6566 4133 6582
rect 4161 6560 4167 6608
rect 4170 6602 4189 6608
rect 4204 6602 4234 6610
rect 4170 6594 4234 6602
rect 4170 6578 4250 6594
rect 4266 6587 4328 6618
rect 4344 6587 4406 6618
rect 4475 6616 4524 6641
rect 4539 6616 4569 6632
rect 4438 6602 4468 6610
rect 4475 6608 4585 6616
rect 4438 6594 4483 6602
rect 4170 6576 4189 6578
rect 4204 6576 4250 6578
rect 4170 6560 4250 6576
rect 4277 6574 4312 6587
rect 4353 6584 4390 6587
rect 4353 6582 4395 6584
rect 4282 6571 4312 6574
rect 4291 6567 4298 6571
rect 4298 6566 4299 6567
rect 4257 6560 4267 6566
rect 4016 6552 4051 6560
rect 4016 6526 4017 6552
rect 4024 6526 4051 6552
rect 3959 6508 3989 6522
rect 4016 6518 4051 6526
rect 4053 6552 4094 6560
rect 4053 6526 4068 6552
rect 4075 6526 4094 6552
rect 4158 6548 4189 6560
rect 4204 6548 4307 6560
rect 4319 6550 4345 6576
rect 4360 6571 4390 6582
rect 4422 6578 4484 6594
rect 4422 6576 4468 6578
rect 4422 6560 4484 6576
rect 4496 6560 4502 6608
rect 4505 6600 4585 6608
rect 4505 6598 4524 6600
rect 4539 6598 4573 6600
rect 4505 6582 4585 6598
rect 4505 6560 4524 6582
rect 4539 6566 4569 6582
rect 4597 6576 4603 6650
rect 4606 6576 4625 6720
rect 4640 6576 4646 6720
rect 4655 6650 4668 6720
rect 4720 6716 4742 6720
rect 4713 6694 4742 6708
rect 4795 6694 4811 6708
rect 4849 6704 4855 6706
rect 4862 6704 4970 6720
rect 4977 6704 4983 6706
rect 4991 6704 5006 6720
rect 5072 6714 5091 6717
rect 4713 6692 4811 6694
rect 4838 6692 5006 6704
rect 5021 6694 5037 6708
rect 5072 6695 5094 6714
rect 5104 6708 5120 6709
rect 5103 6706 5120 6708
rect 5104 6701 5120 6706
rect 5094 6694 5100 6695
rect 5103 6694 5132 6701
rect 5021 6693 5132 6694
rect 5021 6692 5138 6693
rect 4697 6684 4748 6692
rect 4795 6684 4829 6692
rect 4697 6672 4722 6684
rect 4729 6672 4748 6684
rect 4802 6682 4829 6684
rect 4838 6682 5059 6692
rect 5094 6689 5100 6692
rect 4802 6678 5059 6682
rect 4697 6664 4748 6672
rect 4795 6664 5059 6678
rect 5103 6684 5138 6692
rect 4649 6616 4668 6650
rect 4713 6656 4742 6664
rect 4713 6650 4730 6656
rect 4713 6648 4747 6650
rect 4795 6648 4811 6664
rect 4812 6654 5020 6664
rect 5021 6654 5037 6664
rect 5085 6660 5100 6675
rect 5103 6672 5104 6684
rect 5111 6672 5138 6684
rect 5103 6664 5138 6672
rect 5103 6663 5132 6664
rect 4823 6650 5037 6654
rect 4838 6648 5037 6650
rect 5072 6650 5085 6660
rect 5103 6650 5120 6663
rect 5072 6648 5120 6650
rect 4714 6644 4747 6648
rect 4710 6642 4747 6644
rect 4710 6641 4777 6642
rect 4710 6636 4741 6641
rect 4747 6636 4777 6641
rect 4710 6632 4777 6636
rect 4683 6629 4777 6632
rect 4683 6622 4732 6629
rect 4683 6616 4713 6622
rect 4732 6617 4737 6622
rect 4649 6600 4729 6616
rect 4741 6608 4777 6629
rect 4838 6624 5027 6648
rect 5072 6647 5119 6648
rect 5085 6642 5119 6647
rect 4853 6621 5027 6624
rect 4846 6618 5027 6621
rect 5055 6641 5119 6642
rect 4649 6598 4668 6600
rect 4683 6598 4717 6600
rect 4649 6582 4729 6598
rect 4649 6576 4668 6582
rect 4365 6550 4468 6560
rect 4319 6548 4468 6550
rect 4489 6548 4524 6560
rect 4158 6546 4320 6548
rect 4170 6526 4189 6546
rect 4204 6544 4234 6546
rect 4053 6518 4094 6526
rect 4176 6522 4189 6526
rect 4241 6530 4320 6546
rect 4352 6546 4524 6548
rect 4352 6530 4431 6546
rect 4438 6544 4468 6546
rect 4016 6508 4045 6518
rect 4059 6508 4088 6518
rect 4103 6508 4133 6522
rect 4176 6508 4219 6522
rect 4241 6518 4431 6530
rect 4496 6526 4502 6546
rect 4226 6508 4256 6518
rect 4257 6508 4415 6518
rect 4419 6508 4449 6518
rect 4453 6508 4483 6522
rect 4511 6508 4524 6546
rect 4596 6560 4625 6576
rect 4639 6560 4668 6576
rect 4683 6566 4713 6582
rect 4741 6560 4747 6608
rect 4750 6602 4769 6608
rect 4784 6602 4814 6610
rect 4750 6594 4814 6602
rect 4750 6578 4830 6594
rect 4846 6587 4908 6618
rect 4924 6587 4986 6618
rect 5055 6616 5104 6641
rect 5119 6616 5149 6632
rect 5018 6602 5048 6610
rect 5055 6608 5165 6616
rect 5018 6594 5063 6602
rect 4750 6576 4769 6578
rect 4784 6576 4830 6578
rect 4750 6560 4830 6576
rect 4857 6574 4892 6587
rect 4933 6584 4970 6587
rect 4933 6582 4975 6584
rect 4862 6571 4892 6574
rect 4871 6567 4878 6571
rect 4878 6566 4879 6567
rect 4837 6560 4847 6566
rect 4596 6552 4631 6560
rect 4596 6526 4597 6552
rect 4604 6526 4631 6552
rect 4539 6508 4569 6522
rect 4596 6518 4631 6526
rect 4633 6552 4674 6560
rect 4633 6526 4648 6552
rect 4655 6526 4674 6552
rect 4738 6548 4769 6560
rect 4784 6548 4887 6560
rect 4899 6550 4925 6576
rect 4940 6571 4970 6582
rect 5002 6578 5064 6594
rect 5002 6576 5048 6578
rect 5002 6560 5064 6576
rect 5076 6560 5082 6608
rect 5085 6600 5165 6608
rect 5085 6598 5104 6600
rect 5119 6598 5153 6600
rect 5085 6582 5165 6598
rect 5085 6560 5104 6582
rect 5119 6566 5149 6582
rect 5177 6576 5183 6650
rect 5186 6576 5205 6720
rect 5220 6576 5226 6720
rect 5235 6650 5248 6720
rect 5300 6716 5322 6720
rect 5293 6694 5322 6708
rect 5375 6694 5391 6708
rect 5429 6704 5435 6706
rect 5442 6704 5550 6720
rect 5557 6704 5563 6706
rect 5571 6704 5586 6720
rect 5652 6714 5671 6717
rect 5293 6692 5391 6694
rect 5418 6692 5586 6704
rect 5601 6694 5617 6708
rect 5652 6695 5674 6714
rect 5684 6708 5700 6709
rect 5683 6706 5700 6708
rect 5684 6701 5700 6706
rect 5674 6694 5680 6695
rect 5683 6694 5712 6701
rect 5601 6693 5712 6694
rect 5601 6692 5718 6693
rect 5277 6684 5328 6692
rect 5375 6684 5409 6692
rect 5277 6672 5302 6684
rect 5309 6672 5328 6684
rect 5382 6682 5409 6684
rect 5418 6682 5639 6692
rect 5674 6689 5680 6692
rect 5382 6678 5639 6682
rect 5277 6664 5328 6672
rect 5375 6664 5639 6678
rect 5683 6684 5718 6692
rect 5229 6616 5248 6650
rect 5293 6656 5322 6664
rect 5293 6650 5310 6656
rect 5293 6648 5327 6650
rect 5375 6648 5391 6664
rect 5392 6654 5600 6664
rect 5601 6654 5617 6664
rect 5665 6660 5680 6675
rect 5683 6672 5684 6684
rect 5691 6672 5718 6684
rect 5683 6664 5718 6672
rect 5683 6663 5712 6664
rect 5403 6650 5617 6654
rect 5418 6648 5617 6650
rect 5652 6650 5665 6660
rect 5683 6650 5700 6663
rect 5652 6648 5700 6650
rect 5294 6644 5327 6648
rect 5290 6642 5327 6644
rect 5290 6641 5357 6642
rect 5290 6636 5321 6641
rect 5327 6636 5357 6641
rect 5290 6632 5357 6636
rect 5263 6629 5357 6632
rect 5263 6622 5312 6629
rect 5263 6616 5293 6622
rect 5312 6617 5317 6622
rect 5229 6600 5309 6616
rect 5321 6608 5357 6629
rect 5418 6624 5607 6648
rect 5652 6647 5699 6648
rect 5665 6642 5699 6647
rect 5433 6621 5607 6624
rect 5426 6618 5607 6621
rect 5635 6641 5699 6642
rect 5229 6598 5248 6600
rect 5263 6598 5297 6600
rect 5229 6582 5309 6598
rect 5229 6576 5248 6582
rect 4945 6550 5048 6560
rect 4899 6548 5048 6550
rect 5069 6548 5104 6560
rect 4738 6546 4900 6548
rect 4750 6526 4769 6546
rect 4784 6544 4814 6546
rect 4633 6518 4674 6526
rect 4756 6522 4769 6526
rect 4821 6530 4900 6546
rect 4932 6546 5104 6548
rect 4932 6530 5011 6546
rect 5018 6544 5048 6546
rect 4596 6508 4625 6518
rect 4639 6508 4668 6518
rect 4683 6508 4713 6522
rect 4756 6508 4799 6522
rect 4821 6518 5011 6530
rect 5076 6526 5082 6546
rect 4806 6508 4836 6518
rect 4837 6508 4995 6518
rect 4999 6508 5029 6518
rect 5033 6508 5063 6522
rect 5091 6508 5104 6546
rect 5176 6560 5205 6576
rect 5219 6560 5248 6576
rect 5263 6566 5293 6582
rect 5321 6560 5327 6608
rect 5330 6602 5349 6608
rect 5364 6602 5394 6610
rect 5330 6594 5394 6602
rect 5330 6578 5410 6594
rect 5426 6587 5488 6618
rect 5504 6587 5566 6618
rect 5635 6616 5684 6641
rect 5699 6616 5729 6632
rect 5598 6602 5628 6610
rect 5635 6608 5745 6616
rect 5598 6594 5643 6602
rect 5330 6576 5349 6578
rect 5364 6576 5410 6578
rect 5330 6560 5410 6576
rect 5437 6574 5472 6587
rect 5513 6584 5550 6587
rect 5513 6582 5555 6584
rect 5442 6571 5472 6574
rect 5451 6567 5458 6571
rect 5458 6566 5459 6567
rect 5417 6560 5427 6566
rect 5176 6552 5211 6560
rect 5176 6526 5177 6552
rect 5184 6526 5211 6552
rect 5119 6508 5149 6522
rect 5176 6518 5211 6526
rect 5213 6552 5254 6560
rect 5213 6526 5228 6552
rect 5235 6526 5254 6552
rect 5318 6548 5349 6560
rect 5364 6548 5467 6560
rect 5479 6550 5505 6576
rect 5520 6571 5550 6582
rect 5582 6578 5644 6594
rect 5582 6576 5628 6578
rect 5582 6560 5644 6576
rect 5656 6560 5662 6608
rect 5665 6600 5745 6608
rect 5665 6598 5684 6600
rect 5699 6598 5733 6600
rect 5665 6582 5745 6598
rect 5665 6560 5684 6582
rect 5699 6566 5729 6582
rect 5757 6576 5763 6650
rect 5766 6576 5785 6720
rect 5800 6576 5806 6720
rect 5815 6650 5828 6720
rect 5880 6716 5902 6720
rect 5873 6694 5902 6708
rect 5955 6694 5971 6708
rect 6009 6704 6015 6706
rect 6022 6704 6130 6720
rect 6137 6704 6143 6706
rect 6151 6704 6166 6720
rect 6232 6714 6251 6717
rect 5873 6692 5971 6694
rect 5998 6692 6166 6704
rect 6181 6694 6197 6708
rect 6232 6695 6254 6714
rect 6264 6708 6280 6709
rect 6263 6706 6280 6708
rect 6264 6701 6280 6706
rect 6254 6694 6260 6695
rect 6263 6694 6292 6701
rect 6181 6693 6292 6694
rect 6181 6692 6298 6693
rect 5857 6684 5908 6692
rect 5955 6684 5989 6692
rect 5857 6672 5882 6684
rect 5889 6672 5908 6684
rect 5962 6682 5989 6684
rect 5998 6682 6219 6692
rect 6254 6689 6260 6692
rect 5962 6678 6219 6682
rect 5857 6664 5908 6672
rect 5955 6664 6219 6678
rect 6263 6684 6298 6692
rect 5809 6616 5828 6650
rect 5873 6656 5902 6664
rect 5873 6650 5890 6656
rect 5873 6648 5907 6650
rect 5955 6648 5971 6664
rect 5972 6654 6180 6664
rect 6181 6654 6197 6664
rect 6245 6660 6260 6675
rect 6263 6672 6264 6684
rect 6271 6672 6298 6684
rect 6263 6664 6298 6672
rect 6263 6663 6292 6664
rect 5983 6650 6197 6654
rect 5998 6648 6197 6650
rect 6232 6650 6245 6660
rect 6263 6650 6280 6663
rect 6232 6648 6280 6650
rect 5874 6644 5907 6648
rect 5870 6642 5907 6644
rect 5870 6641 5937 6642
rect 5870 6636 5901 6641
rect 5907 6636 5937 6641
rect 5870 6632 5937 6636
rect 5843 6629 5937 6632
rect 5843 6622 5892 6629
rect 5843 6616 5873 6622
rect 5892 6617 5897 6622
rect 5809 6600 5889 6616
rect 5901 6608 5937 6629
rect 5998 6624 6187 6648
rect 6232 6647 6279 6648
rect 6245 6642 6279 6647
rect 6013 6621 6187 6624
rect 6006 6618 6187 6621
rect 6215 6641 6279 6642
rect 5809 6598 5828 6600
rect 5843 6598 5877 6600
rect 5809 6582 5889 6598
rect 5809 6576 5828 6582
rect 5525 6550 5628 6560
rect 5479 6548 5628 6550
rect 5649 6548 5684 6560
rect 5318 6546 5480 6548
rect 5330 6526 5349 6546
rect 5364 6544 5394 6546
rect 5213 6518 5254 6526
rect 5336 6522 5349 6526
rect 5401 6530 5480 6546
rect 5512 6546 5684 6548
rect 5512 6530 5591 6546
rect 5598 6544 5628 6546
rect 5176 6508 5205 6518
rect 5219 6508 5248 6518
rect 5263 6508 5293 6522
rect 5336 6508 5379 6522
rect 5401 6518 5591 6530
rect 5656 6526 5662 6546
rect 5386 6508 5416 6518
rect 5417 6508 5575 6518
rect 5579 6508 5609 6518
rect 5613 6508 5643 6522
rect 5671 6508 5684 6546
rect 5756 6560 5785 6576
rect 5799 6560 5828 6576
rect 5843 6566 5873 6582
rect 5901 6560 5907 6608
rect 5910 6602 5929 6608
rect 5944 6602 5974 6610
rect 5910 6594 5974 6602
rect 5910 6578 5990 6594
rect 6006 6587 6068 6618
rect 6084 6587 6146 6618
rect 6215 6616 6264 6641
rect 6279 6616 6309 6632
rect 6178 6602 6208 6610
rect 6215 6608 6325 6616
rect 6178 6594 6223 6602
rect 5910 6576 5929 6578
rect 5944 6576 5990 6578
rect 5910 6560 5990 6576
rect 6017 6574 6052 6587
rect 6093 6584 6130 6587
rect 6093 6582 6135 6584
rect 6022 6571 6052 6574
rect 6031 6567 6038 6571
rect 6038 6566 6039 6567
rect 5997 6560 6007 6566
rect 5756 6552 5791 6560
rect 5756 6526 5757 6552
rect 5764 6526 5791 6552
rect 5699 6508 5729 6522
rect 5756 6518 5791 6526
rect 5793 6552 5834 6560
rect 5793 6526 5808 6552
rect 5815 6526 5834 6552
rect 5898 6548 5929 6560
rect 5944 6548 6047 6560
rect 6059 6550 6085 6576
rect 6100 6571 6130 6582
rect 6162 6578 6224 6594
rect 6162 6576 6208 6578
rect 6162 6560 6224 6576
rect 6236 6560 6242 6608
rect 6245 6600 6325 6608
rect 6245 6598 6264 6600
rect 6279 6598 6313 6600
rect 6245 6582 6325 6598
rect 6245 6560 6264 6582
rect 6279 6566 6309 6582
rect 6337 6576 6343 6650
rect 6346 6576 6365 6720
rect 6380 6576 6386 6720
rect 6395 6650 6408 6720
rect 6460 6716 6482 6720
rect 6453 6694 6482 6708
rect 6535 6694 6551 6708
rect 6589 6704 6595 6706
rect 6602 6704 6710 6720
rect 6717 6704 6723 6706
rect 6731 6704 6746 6720
rect 6812 6714 6831 6717
rect 6453 6692 6551 6694
rect 6578 6692 6746 6704
rect 6761 6694 6777 6708
rect 6812 6695 6834 6714
rect 6844 6708 6860 6709
rect 6843 6706 6860 6708
rect 6844 6701 6860 6706
rect 6834 6694 6840 6695
rect 6843 6694 6872 6701
rect 6761 6693 6872 6694
rect 6761 6692 6878 6693
rect 6437 6684 6488 6692
rect 6535 6684 6569 6692
rect 6437 6672 6462 6684
rect 6469 6672 6488 6684
rect 6542 6682 6569 6684
rect 6578 6682 6799 6692
rect 6834 6689 6840 6692
rect 6542 6678 6799 6682
rect 6437 6664 6488 6672
rect 6535 6664 6799 6678
rect 6843 6684 6878 6692
rect 6389 6616 6408 6650
rect 6453 6656 6482 6664
rect 6453 6650 6470 6656
rect 6453 6648 6487 6650
rect 6535 6648 6551 6664
rect 6552 6654 6760 6664
rect 6761 6654 6777 6664
rect 6825 6660 6840 6675
rect 6843 6672 6844 6684
rect 6851 6672 6878 6684
rect 6843 6664 6878 6672
rect 6843 6663 6872 6664
rect 6563 6650 6777 6654
rect 6578 6648 6777 6650
rect 6812 6650 6825 6660
rect 6843 6650 6860 6663
rect 6812 6648 6860 6650
rect 6454 6644 6487 6648
rect 6450 6642 6487 6644
rect 6450 6641 6517 6642
rect 6450 6636 6481 6641
rect 6487 6636 6517 6641
rect 6450 6632 6517 6636
rect 6423 6629 6517 6632
rect 6423 6622 6472 6629
rect 6423 6616 6453 6622
rect 6472 6617 6477 6622
rect 6389 6600 6469 6616
rect 6481 6608 6517 6629
rect 6578 6624 6767 6648
rect 6812 6647 6859 6648
rect 6825 6642 6859 6647
rect 6593 6621 6767 6624
rect 6586 6618 6767 6621
rect 6795 6641 6859 6642
rect 6389 6598 6408 6600
rect 6423 6598 6457 6600
rect 6389 6582 6469 6598
rect 6389 6576 6408 6582
rect 6105 6550 6208 6560
rect 6059 6548 6208 6550
rect 6229 6548 6264 6560
rect 5898 6546 6060 6548
rect 5910 6526 5929 6546
rect 5944 6544 5974 6546
rect 5793 6518 5834 6526
rect 5916 6522 5929 6526
rect 5981 6530 6060 6546
rect 6092 6546 6264 6548
rect 6092 6530 6171 6546
rect 6178 6544 6208 6546
rect 5756 6508 5785 6518
rect 5799 6508 5828 6518
rect 5843 6508 5873 6522
rect 5916 6508 5959 6522
rect 5981 6518 6171 6530
rect 6236 6526 6242 6546
rect 5966 6508 5996 6518
rect 5997 6508 6155 6518
rect 6159 6508 6189 6518
rect 6193 6508 6223 6522
rect 6251 6508 6264 6546
rect 6336 6560 6365 6576
rect 6379 6560 6408 6576
rect 6423 6566 6453 6582
rect 6481 6560 6487 6608
rect 6490 6602 6509 6608
rect 6524 6602 6554 6610
rect 6490 6594 6554 6602
rect 6490 6578 6570 6594
rect 6586 6587 6648 6618
rect 6664 6587 6726 6618
rect 6795 6616 6844 6641
rect 6859 6616 6889 6632
rect 6758 6602 6788 6610
rect 6795 6608 6905 6616
rect 6758 6594 6803 6602
rect 6490 6576 6509 6578
rect 6524 6576 6570 6578
rect 6490 6560 6570 6576
rect 6597 6574 6632 6587
rect 6673 6584 6710 6587
rect 6673 6582 6715 6584
rect 6602 6571 6632 6574
rect 6611 6567 6618 6571
rect 6618 6566 6619 6567
rect 6577 6560 6587 6566
rect 6336 6552 6371 6560
rect 6336 6526 6337 6552
rect 6344 6526 6371 6552
rect 6279 6508 6309 6522
rect 6336 6518 6371 6526
rect 6373 6552 6414 6560
rect 6373 6526 6388 6552
rect 6395 6526 6414 6552
rect 6478 6548 6509 6560
rect 6524 6548 6627 6560
rect 6639 6550 6665 6576
rect 6680 6571 6710 6582
rect 6742 6578 6804 6594
rect 6742 6576 6788 6578
rect 6742 6560 6804 6576
rect 6816 6560 6822 6608
rect 6825 6600 6905 6608
rect 6825 6598 6844 6600
rect 6859 6598 6893 6600
rect 6825 6582 6905 6598
rect 6825 6560 6844 6582
rect 6859 6566 6889 6582
rect 6917 6576 6923 6650
rect 6926 6576 6945 6720
rect 6960 6576 6966 6720
rect 6975 6650 6988 6720
rect 7040 6716 7062 6720
rect 7033 6694 7062 6708
rect 7115 6694 7131 6708
rect 7169 6704 7175 6706
rect 7182 6704 7290 6720
rect 7297 6704 7303 6706
rect 7311 6704 7326 6720
rect 7392 6714 7411 6717
rect 7033 6692 7131 6694
rect 7158 6692 7326 6704
rect 7341 6694 7357 6708
rect 7392 6695 7414 6714
rect 7424 6708 7440 6709
rect 7423 6706 7440 6708
rect 7424 6701 7440 6706
rect 7414 6694 7420 6695
rect 7423 6694 7452 6701
rect 7341 6693 7452 6694
rect 7341 6692 7458 6693
rect 7017 6684 7068 6692
rect 7115 6684 7149 6692
rect 7017 6672 7042 6684
rect 7049 6672 7068 6684
rect 7122 6682 7149 6684
rect 7158 6682 7379 6692
rect 7414 6689 7420 6692
rect 7122 6678 7379 6682
rect 7017 6664 7068 6672
rect 7115 6664 7379 6678
rect 7423 6684 7458 6692
rect 6969 6616 6988 6650
rect 7033 6656 7062 6664
rect 7033 6650 7050 6656
rect 7033 6648 7067 6650
rect 7115 6648 7131 6664
rect 7132 6654 7340 6664
rect 7341 6654 7357 6664
rect 7405 6660 7420 6675
rect 7423 6672 7424 6684
rect 7431 6672 7458 6684
rect 7423 6664 7458 6672
rect 7423 6663 7452 6664
rect 7143 6650 7357 6654
rect 7158 6648 7357 6650
rect 7392 6650 7405 6660
rect 7423 6650 7440 6663
rect 7392 6648 7440 6650
rect 7034 6644 7067 6648
rect 7030 6642 7067 6644
rect 7030 6641 7097 6642
rect 7030 6636 7061 6641
rect 7067 6636 7097 6641
rect 7030 6632 7097 6636
rect 7003 6629 7097 6632
rect 7003 6622 7052 6629
rect 7003 6616 7033 6622
rect 7052 6617 7057 6622
rect 6969 6600 7049 6616
rect 7061 6608 7097 6629
rect 7158 6624 7347 6648
rect 7392 6647 7439 6648
rect 7405 6642 7439 6647
rect 7173 6621 7347 6624
rect 7166 6618 7347 6621
rect 7375 6641 7439 6642
rect 6969 6598 6988 6600
rect 7003 6598 7037 6600
rect 6969 6582 7049 6598
rect 6969 6576 6988 6582
rect 6685 6550 6788 6560
rect 6639 6548 6788 6550
rect 6809 6548 6844 6560
rect 6478 6546 6640 6548
rect 6490 6526 6509 6546
rect 6524 6544 6554 6546
rect 6373 6518 6414 6526
rect 6496 6522 6509 6526
rect 6561 6530 6640 6546
rect 6672 6546 6844 6548
rect 6672 6530 6751 6546
rect 6758 6544 6788 6546
rect 6336 6508 6365 6518
rect 6379 6508 6408 6518
rect 6423 6508 6453 6522
rect 6496 6508 6539 6522
rect 6561 6518 6751 6530
rect 6816 6526 6822 6546
rect 6546 6508 6576 6518
rect 6577 6508 6735 6518
rect 6739 6508 6769 6518
rect 6773 6508 6803 6522
rect 6831 6508 6844 6546
rect 6916 6560 6945 6576
rect 6959 6560 6988 6576
rect 7003 6566 7033 6582
rect 7061 6560 7067 6608
rect 7070 6602 7089 6608
rect 7104 6602 7134 6610
rect 7070 6594 7134 6602
rect 7070 6578 7150 6594
rect 7166 6587 7228 6618
rect 7244 6587 7306 6618
rect 7375 6616 7424 6641
rect 7439 6616 7469 6632
rect 7338 6602 7368 6610
rect 7375 6608 7485 6616
rect 7338 6594 7383 6602
rect 7070 6576 7089 6578
rect 7104 6576 7150 6578
rect 7070 6560 7150 6576
rect 7177 6574 7212 6587
rect 7253 6584 7290 6587
rect 7253 6582 7295 6584
rect 7182 6571 7212 6574
rect 7191 6567 7198 6571
rect 7198 6566 7199 6567
rect 7157 6560 7167 6566
rect 6916 6552 6951 6560
rect 6916 6526 6917 6552
rect 6924 6526 6951 6552
rect 6859 6508 6889 6522
rect 6916 6518 6951 6526
rect 6953 6552 6994 6560
rect 6953 6526 6968 6552
rect 6975 6526 6994 6552
rect 7058 6548 7089 6560
rect 7104 6548 7207 6560
rect 7219 6550 7245 6576
rect 7260 6571 7290 6582
rect 7322 6578 7384 6594
rect 7322 6576 7368 6578
rect 7322 6560 7384 6576
rect 7396 6560 7402 6608
rect 7405 6600 7485 6608
rect 7405 6598 7424 6600
rect 7439 6598 7473 6600
rect 7405 6582 7485 6598
rect 7405 6560 7424 6582
rect 7439 6566 7469 6582
rect 7497 6576 7503 6650
rect 7506 6576 7525 6720
rect 7540 6576 7546 6720
rect 7555 6650 7568 6720
rect 7613 6698 7614 6708
rect 7629 6698 7642 6708
rect 7613 6694 7642 6698
rect 7647 6694 7677 6720
rect 7695 6706 7711 6708
rect 7783 6706 7836 6720
rect 7784 6704 7848 6706
rect 7891 6704 7906 6720
rect 7955 6717 7985 6720
rect 7955 6714 7991 6717
rect 7921 6706 7937 6708
rect 7695 6694 7710 6698
rect 7613 6692 7710 6694
rect 7738 6692 7906 6704
rect 7922 6694 7937 6698
rect 7955 6695 7994 6714
rect 8013 6708 8020 6709
rect 8019 6701 8020 6708
rect 8003 6698 8004 6701
rect 8019 6698 8032 6701
rect 7955 6694 7985 6695
rect 7994 6694 8000 6695
rect 8003 6694 8032 6698
rect 7922 6693 8032 6694
rect 7922 6692 8038 6693
rect 7597 6684 7648 6692
rect 7597 6672 7622 6684
rect 7629 6672 7648 6684
rect 7679 6684 7729 6692
rect 7679 6676 7695 6684
rect 7702 6682 7729 6684
rect 7738 6682 7959 6692
rect 7702 6672 7959 6682
rect 7988 6684 8038 6692
rect 7988 6675 8004 6684
rect 7597 6664 7648 6672
rect 7695 6664 7959 6672
rect 7985 6672 8004 6675
rect 8011 6672 8038 6684
rect 7985 6664 8038 6672
rect 7549 6616 7568 6650
rect 7613 6656 7614 6664
rect 7629 6656 7642 6664
rect 7613 6648 7629 6656
rect 7610 6641 7629 6644
rect 7610 6632 7632 6641
rect 7583 6622 7632 6632
rect 7583 6616 7613 6622
rect 7632 6617 7637 6622
rect 7549 6600 7629 6616
rect 7647 6608 7677 6664
rect 7712 6654 7920 6664
rect 7955 6660 8000 6664
rect 8003 6663 8004 6664
rect 8019 6663 8032 6664
rect 7738 6624 7927 6654
rect 7753 6621 7927 6624
rect 7746 6618 7927 6621
rect 7549 6598 7568 6600
rect 7583 6598 7617 6600
rect 7549 6582 7629 6598
rect 7656 6594 7669 6608
rect 7684 6594 7700 6610
rect 7746 6605 7757 6618
rect 7549 6576 7568 6582
rect 7265 6550 7368 6560
rect 7219 6548 7368 6550
rect 7389 6548 7424 6560
rect 7058 6546 7220 6548
rect 7070 6526 7089 6546
rect 7104 6544 7134 6546
rect 6953 6518 6994 6526
rect 7076 6522 7089 6526
rect 7141 6530 7220 6546
rect 7252 6546 7424 6548
rect 7252 6530 7331 6546
rect 7338 6544 7368 6546
rect 6916 6508 6945 6518
rect 6959 6508 6988 6518
rect 7003 6508 7033 6522
rect 7076 6508 7119 6522
rect 7141 6518 7331 6530
rect 7396 6526 7402 6546
rect 7126 6508 7156 6518
rect 7157 6508 7315 6518
rect 7319 6508 7349 6518
rect 7353 6508 7383 6522
rect 7411 6508 7424 6546
rect 7496 6560 7525 6576
rect 7539 6560 7568 6576
rect 7583 6560 7613 6582
rect 7656 6578 7718 6594
rect 7746 6587 7757 6603
rect 7762 6598 7772 6618
rect 7782 6598 7796 6618
rect 7799 6605 7808 6618
rect 7824 6605 7833 6618
rect 7762 6587 7796 6598
rect 7799 6587 7808 6603
rect 7824 6587 7833 6603
rect 7840 6598 7850 6618
rect 7860 6598 7874 6618
rect 7875 6605 7886 6618
rect 7840 6587 7874 6598
rect 7875 6587 7886 6603
rect 7932 6594 7948 6610
rect 7955 6608 7985 6660
rect 8019 6656 8020 6663
rect 8004 6648 8020 6656
rect 7991 6616 8004 6635
rect 8019 6616 8049 6632
rect 7991 6600 8065 6616
rect 7991 6598 8004 6600
rect 8019 6598 8053 6600
rect 7656 6576 7669 6578
rect 7684 6576 7718 6578
rect 7656 6560 7718 6576
rect 7762 6571 7778 6574
rect 7840 6571 7870 6582
rect 7918 6578 7964 6594
rect 7991 6582 8065 6598
rect 7918 6576 7952 6578
rect 7917 6560 7964 6576
rect 7991 6560 8004 6582
rect 8019 6560 8049 6582
rect 8076 6560 8077 6576
rect 8092 6560 8105 6720
rect 8135 6616 8148 6720
rect 8193 6698 8194 6708
rect 8209 6698 8222 6708
rect 8193 6694 8222 6698
rect 8227 6694 8257 6720
rect 8275 6706 8291 6708
rect 8363 6706 8416 6720
rect 8364 6704 8428 6706
rect 8471 6704 8486 6720
rect 8535 6717 8565 6720
rect 8535 6714 8571 6717
rect 8501 6706 8517 6708
rect 8275 6694 8290 6698
rect 8193 6692 8290 6694
rect 8318 6692 8486 6704
rect 8502 6694 8517 6698
rect 8535 6695 8574 6714
rect 8593 6708 8600 6709
rect 8599 6701 8600 6708
rect 8583 6698 8584 6701
rect 8599 6698 8612 6701
rect 8535 6694 8565 6695
rect 8574 6694 8580 6695
rect 8583 6694 8612 6698
rect 8502 6693 8612 6694
rect 8502 6692 8618 6693
rect 8177 6684 8228 6692
rect 8177 6672 8202 6684
rect 8209 6672 8228 6684
rect 8259 6684 8309 6692
rect 8259 6676 8275 6684
rect 8282 6682 8309 6684
rect 8318 6682 8539 6692
rect 8282 6672 8539 6682
rect 8568 6684 8618 6692
rect 8568 6675 8584 6684
rect 8177 6664 8228 6672
rect 8275 6664 8539 6672
rect 8565 6672 8584 6675
rect 8591 6672 8618 6684
rect 8565 6664 8618 6672
rect 8193 6656 8194 6664
rect 8209 6656 8222 6664
rect 8193 6648 8209 6656
rect 8190 6641 8209 6644
rect 8190 6632 8212 6641
rect 8163 6622 8212 6632
rect 8163 6616 8193 6622
rect 8212 6617 8217 6622
rect 8135 6600 8209 6616
rect 8227 6608 8257 6664
rect 8292 6654 8500 6664
rect 8535 6660 8580 6664
rect 8583 6663 8584 6664
rect 8599 6663 8612 6664
rect 8318 6624 8507 6654
rect 8333 6621 8507 6624
rect 8326 6618 8507 6621
rect 8135 6598 8148 6600
rect 8163 6598 8197 6600
rect 8135 6582 8209 6598
rect 8236 6594 8249 6608
rect 8264 6594 8280 6610
rect 8326 6605 8337 6618
rect 8119 6560 8120 6576
rect 8135 6560 8148 6582
rect 8163 6560 8193 6582
rect 8236 6578 8298 6594
rect 8326 6587 8337 6603
rect 8342 6598 8352 6618
rect 8362 6598 8376 6618
rect 8379 6605 8388 6618
rect 8404 6605 8413 6618
rect 8342 6587 8376 6598
rect 8379 6587 8388 6603
rect 8404 6587 8413 6603
rect 8420 6598 8430 6618
rect 8440 6598 8454 6618
rect 8455 6605 8466 6618
rect 8420 6587 8454 6598
rect 8455 6587 8466 6603
rect 8512 6594 8528 6610
rect 8535 6608 8565 6660
rect 8599 6656 8600 6663
rect 8584 6648 8600 6656
rect 8571 6616 8584 6635
rect 8599 6616 8629 6632
rect 8571 6600 8645 6616
rect 8571 6598 8584 6600
rect 8599 6598 8633 6600
rect 8236 6576 8249 6578
rect 8264 6576 8298 6578
rect 8236 6560 8298 6576
rect 8342 6571 8358 6574
rect 8420 6571 8450 6582
rect 8498 6578 8544 6594
rect 8571 6582 8645 6598
rect 8498 6576 8532 6578
rect 8497 6560 8544 6576
rect 8571 6560 8584 6582
rect 8599 6560 8629 6582
rect 8656 6560 8657 6576
rect 8672 6560 8685 6720
rect 8715 6616 8728 6720
rect 8773 6698 8774 6708
rect 8789 6698 8802 6708
rect 8773 6694 8802 6698
rect 8807 6694 8837 6720
rect 8855 6706 8871 6708
rect 8943 6706 8996 6720
rect 8944 6704 9008 6706
rect 9051 6704 9066 6720
rect 9115 6717 9145 6720
rect 9115 6714 9151 6717
rect 9081 6706 9097 6708
rect 8855 6694 8870 6698
rect 8773 6692 8870 6694
rect 8898 6692 9066 6704
rect 9082 6694 9097 6698
rect 9115 6695 9154 6714
rect 9173 6708 9180 6709
rect 9179 6701 9180 6708
rect 9163 6698 9164 6701
rect 9179 6698 9192 6701
rect 9115 6694 9145 6695
rect 9154 6694 9160 6695
rect 9163 6694 9192 6698
rect 9082 6693 9192 6694
rect 9082 6692 9198 6693
rect 8757 6684 8808 6692
rect 8757 6672 8782 6684
rect 8789 6672 8808 6684
rect 8839 6684 8889 6692
rect 8839 6676 8855 6684
rect 8862 6682 8889 6684
rect 8898 6682 9119 6692
rect 8862 6672 9119 6682
rect 9148 6684 9198 6692
rect 9148 6675 9164 6684
rect 8757 6664 8808 6672
rect 8855 6664 9119 6672
rect 9145 6672 9164 6675
rect 9171 6672 9198 6684
rect 9145 6664 9198 6672
rect 8773 6656 8774 6664
rect 8789 6656 8802 6664
rect 8773 6648 8789 6656
rect 8770 6641 8789 6644
rect 8770 6632 8792 6641
rect 8743 6622 8792 6632
rect 8743 6616 8773 6622
rect 8792 6617 8797 6622
rect 8715 6600 8789 6616
rect 8807 6608 8837 6664
rect 8872 6654 9080 6664
rect 9115 6660 9160 6664
rect 9163 6663 9164 6664
rect 9179 6663 9192 6664
rect 8898 6624 9087 6654
rect 8913 6621 9087 6624
rect 8906 6618 9087 6621
rect 8715 6598 8728 6600
rect 8743 6598 8777 6600
rect 8715 6582 8789 6598
rect 8816 6594 8829 6608
rect 8844 6594 8860 6610
rect 8906 6605 8917 6618
rect 8699 6560 8700 6576
rect 8715 6560 8728 6582
rect 8743 6560 8773 6582
rect 8816 6578 8878 6594
rect 8906 6587 8917 6603
rect 8922 6598 8932 6618
rect 8942 6598 8956 6618
rect 8959 6605 8968 6618
rect 8984 6605 8993 6618
rect 8922 6587 8956 6598
rect 8959 6587 8968 6603
rect 8984 6587 8993 6603
rect 9000 6598 9010 6618
rect 9020 6598 9034 6618
rect 9035 6605 9046 6618
rect 9000 6587 9034 6598
rect 9035 6587 9046 6603
rect 9092 6594 9108 6610
rect 9115 6608 9145 6660
rect 9179 6656 9180 6663
rect 9164 6648 9180 6656
rect 9151 6616 9164 6635
rect 9179 6616 9209 6632
rect 9151 6600 9225 6616
rect 9151 6598 9164 6600
rect 9179 6598 9213 6600
rect 8816 6576 8829 6578
rect 8844 6576 8878 6578
rect 8816 6560 8878 6576
rect 8922 6571 8938 6574
rect 9000 6571 9030 6582
rect 9078 6578 9124 6594
rect 9151 6582 9225 6598
rect 9078 6576 9112 6578
rect 9077 6560 9124 6576
rect 9151 6560 9164 6582
rect 9179 6560 9209 6582
rect 9236 6560 9237 6576
rect 9252 6560 9265 6720
rect 7496 6552 7531 6560
rect 7496 6526 7497 6552
rect 7504 6526 7531 6552
rect 7439 6508 7469 6522
rect 7496 6518 7531 6526
rect 7533 6552 7574 6560
rect 7533 6526 7548 6552
rect 7555 6526 7574 6552
rect 7638 6548 7700 6560
rect 7712 6548 7787 6560
rect 7845 6548 7920 6560
rect 7932 6548 7963 6560
rect 7969 6548 8004 6560
rect 7638 6546 7800 6548
rect 7533 6518 7574 6526
rect 7656 6522 7669 6546
rect 7684 6544 7699 6546
rect 7496 6508 7525 6518
rect 7539 6508 7568 6518
rect 7583 6508 7613 6522
rect 7656 6508 7699 6522
rect 7723 6519 7730 6526
rect 7733 6522 7800 6546
rect 7832 6546 8004 6548
rect 7802 6524 7830 6528
rect 7832 6524 7912 6546
rect 7933 6544 7948 6546
rect 7802 6522 7912 6524
rect 7733 6518 7912 6522
rect 7706 6508 7736 6518
rect 7738 6508 7891 6518
rect 7899 6508 7929 6518
rect 7933 6508 7963 6522
rect 7991 6508 8004 6546
rect 8076 6552 8111 6560
rect 8076 6526 8077 6552
rect 8084 6526 8111 6552
rect 8019 6508 8049 6522
rect 8076 6518 8111 6526
rect 8113 6552 8154 6560
rect 8113 6526 8128 6552
rect 8135 6526 8154 6552
rect 8218 6548 8280 6560
rect 8292 6548 8367 6560
rect 8425 6548 8500 6560
rect 8512 6548 8543 6560
rect 8549 6548 8584 6560
rect 8218 6546 8380 6548
rect 8113 6518 8154 6526
rect 8236 6522 8249 6546
rect 8264 6544 8279 6546
rect 8076 6508 8077 6518
rect 8092 6508 8105 6518
rect 8119 6508 8120 6518
rect 8135 6508 8148 6518
rect 8163 6508 8193 6522
rect 8236 6508 8279 6522
rect 8303 6519 8310 6526
rect 8313 6522 8380 6546
rect 8412 6546 8584 6548
rect 8382 6524 8410 6528
rect 8412 6524 8492 6546
rect 8513 6544 8528 6546
rect 8382 6522 8492 6524
rect 8313 6518 8492 6522
rect 8286 6508 8316 6518
rect 8318 6508 8471 6518
rect 8479 6508 8509 6518
rect 8513 6508 8543 6522
rect 8571 6508 8584 6546
rect 8656 6552 8691 6560
rect 8656 6526 8657 6552
rect 8664 6526 8691 6552
rect 8599 6508 8629 6522
rect 8656 6518 8691 6526
rect 8693 6552 8734 6560
rect 8693 6526 8708 6552
rect 8715 6526 8734 6552
rect 8798 6548 8860 6560
rect 8872 6548 8947 6560
rect 9005 6548 9080 6560
rect 9092 6548 9123 6560
rect 9129 6548 9164 6560
rect 8798 6546 8960 6548
rect 8693 6518 8734 6526
rect 8816 6522 8829 6546
rect 8844 6544 8859 6546
rect 8656 6508 8657 6518
rect 8672 6508 8685 6518
rect 8699 6508 8700 6518
rect 8715 6508 8728 6518
rect 8743 6508 8773 6522
rect 8816 6508 8859 6522
rect 8883 6519 8890 6526
rect 8893 6522 8960 6546
rect 8992 6546 9164 6548
rect 8962 6524 8990 6528
rect 8992 6524 9072 6546
rect 9093 6544 9108 6546
rect 8962 6522 9072 6524
rect 8893 6518 9072 6522
rect 8866 6508 8896 6518
rect 8898 6508 9051 6518
rect 9059 6508 9089 6518
rect 9093 6508 9123 6522
rect 9151 6508 9164 6546
rect 9236 6552 9271 6560
rect 9236 6526 9237 6552
rect 9244 6526 9271 6552
rect 9179 6508 9209 6522
rect 9236 6518 9271 6526
rect 9236 6508 9237 6518
rect 9252 6508 9265 6518
rect -1 6502 9265 6508
rect 0 6494 9265 6502
rect 15 6464 28 6494
rect 43 6480 73 6494
rect 116 6480 159 6494
rect 166 6480 386 6494
rect 393 6480 423 6494
rect 83 6466 98 6478
rect 117 6466 130 6480
rect 198 6476 351 6480
rect 80 6464 102 6466
rect 180 6464 372 6476
rect 451 6464 464 6494
rect 479 6480 509 6494
rect 546 6464 565 6494
rect 580 6464 586 6494
rect 595 6464 608 6494
rect 623 6480 653 6494
rect 696 6480 739 6494
rect 746 6480 966 6494
rect 973 6480 1003 6494
rect 663 6466 678 6478
rect 697 6466 710 6480
rect 778 6476 931 6480
rect 660 6464 682 6466
rect 760 6464 952 6476
rect 1031 6464 1044 6494
rect 1059 6480 1089 6494
rect 1126 6464 1145 6494
rect 1160 6464 1166 6494
rect 1175 6464 1188 6494
rect 1203 6480 1233 6494
rect 1276 6480 1319 6494
rect 1326 6480 1546 6494
rect 1553 6480 1583 6494
rect 1243 6466 1258 6478
rect 1277 6466 1290 6480
rect 1358 6476 1511 6480
rect 1240 6464 1262 6466
rect 1340 6464 1532 6476
rect 1611 6464 1624 6494
rect 1639 6480 1669 6494
rect 1706 6464 1725 6494
rect 1740 6464 1746 6494
rect 1755 6464 1768 6494
rect 1783 6480 1813 6494
rect 1856 6480 1899 6494
rect 1906 6480 2126 6494
rect 2133 6480 2163 6494
rect 1823 6466 1838 6478
rect 1857 6466 1870 6480
rect 1938 6476 2091 6480
rect 1820 6464 1842 6466
rect 1920 6464 2112 6476
rect 2191 6464 2204 6494
rect 2219 6480 2249 6494
rect 2286 6464 2305 6494
rect 2320 6464 2326 6494
rect 2335 6464 2348 6494
rect 2363 6480 2393 6494
rect 2436 6480 2479 6494
rect 2486 6480 2706 6494
rect 2713 6480 2743 6494
rect 2403 6466 2418 6478
rect 2437 6466 2450 6480
rect 2518 6476 2671 6480
rect 2400 6464 2422 6466
rect 2500 6464 2692 6476
rect 2771 6464 2784 6494
rect 2799 6480 2829 6494
rect 2866 6464 2885 6494
rect 2900 6464 2906 6494
rect 2915 6464 2928 6494
rect 2943 6480 2973 6494
rect 3016 6480 3059 6494
rect 3066 6480 3286 6494
rect 3293 6480 3323 6494
rect 2983 6466 2998 6478
rect 3017 6466 3030 6480
rect 3098 6476 3251 6480
rect 2980 6464 3002 6466
rect 3080 6464 3272 6476
rect 3351 6464 3364 6494
rect 3379 6480 3409 6494
rect 3446 6464 3465 6494
rect 3480 6464 3486 6494
rect 3495 6464 3508 6494
rect 3523 6480 3553 6494
rect 3596 6480 3639 6494
rect 3646 6480 3866 6494
rect 3873 6480 3903 6494
rect 3563 6466 3578 6478
rect 3597 6466 3610 6480
rect 3678 6476 3831 6480
rect 3560 6464 3582 6466
rect 3660 6464 3852 6476
rect 3931 6464 3944 6494
rect 3959 6480 3989 6494
rect 4026 6464 4045 6494
rect 4060 6464 4066 6494
rect 4075 6464 4088 6494
rect 4103 6480 4133 6494
rect 4176 6480 4219 6494
rect 4226 6480 4446 6494
rect 4453 6480 4483 6494
rect 4143 6466 4158 6478
rect 4177 6466 4190 6480
rect 4258 6476 4411 6480
rect 4140 6464 4162 6466
rect 4240 6464 4432 6476
rect 4511 6464 4524 6494
rect 4539 6480 4569 6494
rect 4606 6464 4625 6494
rect 4640 6464 4646 6494
rect 4655 6464 4668 6494
rect 4683 6480 4713 6494
rect 4756 6480 4799 6494
rect 4806 6480 5026 6494
rect 5033 6480 5063 6494
rect 4723 6466 4738 6478
rect 4757 6466 4770 6480
rect 4838 6476 4991 6480
rect 4720 6464 4742 6466
rect 4820 6464 5012 6476
rect 5091 6464 5104 6494
rect 5119 6480 5149 6494
rect 5186 6464 5205 6494
rect 5220 6464 5226 6494
rect 5235 6464 5248 6494
rect 5263 6480 5293 6494
rect 5336 6480 5379 6494
rect 5386 6480 5606 6494
rect 5613 6480 5643 6494
rect 5303 6466 5318 6478
rect 5337 6466 5350 6480
rect 5418 6476 5571 6480
rect 5300 6464 5322 6466
rect 5400 6464 5592 6476
rect 5671 6464 5684 6494
rect 5699 6480 5729 6494
rect 5766 6464 5785 6494
rect 5800 6464 5806 6494
rect 5815 6464 5828 6494
rect 5843 6480 5873 6494
rect 5916 6480 5959 6494
rect 5966 6480 6186 6494
rect 6193 6480 6223 6494
rect 5883 6466 5898 6478
rect 5917 6466 5930 6480
rect 5998 6476 6151 6480
rect 5880 6464 5902 6466
rect 5980 6464 6172 6476
rect 6251 6464 6264 6494
rect 6279 6480 6309 6494
rect 6346 6464 6365 6494
rect 6380 6464 6386 6494
rect 6395 6464 6408 6494
rect 6423 6480 6453 6494
rect 6496 6480 6539 6494
rect 6546 6480 6766 6494
rect 6773 6480 6803 6494
rect 6463 6466 6478 6478
rect 6497 6466 6510 6480
rect 6578 6476 6731 6480
rect 6460 6464 6482 6466
rect 6560 6464 6752 6476
rect 6831 6464 6844 6494
rect 6859 6480 6889 6494
rect 6926 6464 6945 6494
rect 6960 6464 6966 6494
rect 6975 6464 6988 6494
rect 7003 6480 7033 6494
rect 7076 6480 7119 6494
rect 7126 6480 7346 6494
rect 7353 6480 7383 6494
rect 7043 6466 7058 6478
rect 7077 6466 7090 6480
rect 7158 6476 7311 6480
rect 7040 6464 7062 6466
rect 7140 6464 7332 6476
rect 7411 6464 7424 6494
rect 7439 6480 7469 6494
rect 7506 6464 7525 6494
rect 7540 6464 7546 6494
rect 7555 6464 7568 6494
rect 7583 6476 7613 6494
rect 7656 6480 7670 6494
rect 7706 6480 7926 6494
rect 7657 6478 7670 6480
rect 7623 6466 7638 6478
rect 7620 6464 7642 6466
rect 7647 6464 7677 6478
rect 7738 6476 7891 6480
rect 7720 6464 7912 6476
rect 7955 6464 7985 6478
rect 7991 6464 8004 6494
rect 8019 6476 8049 6494
rect 8092 6464 8105 6494
rect 8135 6464 8148 6494
rect 8163 6476 8193 6494
rect 8236 6480 8250 6494
rect 8286 6480 8506 6494
rect 8237 6478 8250 6480
rect 8203 6466 8218 6478
rect 8200 6464 8222 6466
rect 8227 6464 8257 6478
rect 8318 6476 8471 6480
rect 8300 6464 8492 6476
rect 8535 6464 8565 6478
rect 8571 6464 8584 6494
rect 8599 6476 8629 6494
rect 8672 6464 8685 6494
rect 8715 6464 8728 6494
rect 8743 6476 8773 6494
rect 8816 6480 8830 6494
rect 8866 6480 9086 6494
rect 8817 6478 8830 6480
rect 8783 6466 8798 6478
rect 8780 6464 8802 6466
rect 8807 6464 8837 6478
rect 8898 6476 9051 6480
rect 8880 6464 9072 6476
rect 9115 6464 9145 6478
rect 9151 6464 9164 6494
rect 9179 6476 9209 6494
rect 9252 6464 9265 6494
rect 0 6450 9265 6464
rect 15 6380 28 6450
rect 80 6446 102 6450
rect 73 6424 102 6438
rect 155 6424 171 6438
rect 209 6434 215 6436
rect 222 6434 330 6450
rect 337 6434 343 6436
rect 351 6434 366 6450
rect 432 6444 451 6447
rect 73 6422 171 6424
rect 198 6422 366 6434
rect 381 6424 397 6438
rect 432 6425 454 6444
rect 464 6438 480 6439
rect 463 6436 480 6438
rect 464 6431 480 6436
rect 454 6424 460 6425
rect 463 6424 492 6431
rect 381 6423 492 6424
rect 381 6422 498 6423
rect 57 6414 108 6422
rect 155 6414 189 6422
rect 57 6402 82 6414
rect 89 6402 108 6414
rect 162 6412 189 6414
rect 198 6412 419 6422
rect 454 6419 460 6422
rect 162 6408 419 6412
rect 57 6394 108 6402
rect 155 6394 419 6408
rect 463 6414 498 6422
rect 9 6346 28 6380
rect 73 6386 102 6394
rect 73 6380 90 6386
rect 73 6378 107 6380
rect 155 6378 171 6394
rect 172 6384 380 6394
rect 381 6384 397 6394
rect 445 6390 460 6405
rect 463 6402 464 6414
rect 471 6402 498 6414
rect 463 6394 498 6402
rect 463 6393 492 6394
rect 183 6380 397 6384
rect 198 6378 397 6380
rect 432 6380 445 6390
rect 463 6380 480 6393
rect 432 6378 480 6380
rect 74 6374 107 6378
rect 70 6372 107 6374
rect 70 6371 137 6372
rect 70 6366 101 6371
rect 107 6366 137 6371
rect 70 6362 137 6366
rect 43 6359 137 6362
rect 43 6352 92 6359
rect 43 6346 73 6352
rect 92 6347 97 6352
rect 9 6330 89 6346
rect 101 6338 137 6359
rect 198 6354 387 6378
rect 432 6377 479 6378
rect 445 6372 479 6377
rect 213 6351 387 6354
rect 206 6348 387 6351
rect 415 6371 479 6372
rect 9 6328 28 6330
rect 43 6328 77 6330
rect 9 6312 89 6328
rect 9 6306 28 6312
rect -1 6290 28 6306
rect 43 6296 73 6312
rect 101 6290 107 6338
rect 110 6332 129 6338
rect 144 6332 174 6340
rect 110 6324 174 6332
rect 110 6308 190 6324
rect 206 6317 268 6348
rect 284 6317 346 6348
rect 415 6346 464 6371
rect 479 6346 509 6362
rect 378 6332 408 6340
rect 415 6338 525 6346
rect 378 6324 423 6332
rect 110 6306 129 6308
rect 144 6306 190 6308
rect 110 6290 190 6306
rect 217 6304 252 6317
rect 293 6314 330 6317
rect 293 6312 335 6314
rect 222 6301 252 6304
rect 231 6297 238 6301
rect 238 6296 239 6297
rect 197 6290 207 6296
rect -7 6282 34 6290
rect -7 6256 8 6282
rect 15 6256 34 6282
rect 98 6278 129 6290
rect 144 6278 247 6290
rect 259 6280 285 6306
rect 300 6301 330 6312
rect 362 6308 424 6324
rect 362 6306 408 6308
rect 362 6290 424 6306
rect 436 6290 442 6338
rect 445 6330 525 6338
rect 445 6328 464 6330
rect 479 6328 513 6330
rect 445 6312 525 6328
rect 445 6290 464 6312
rect 479 6296 509 6312
rect 537 6306 543 6380
rect 546 6306 565 6450
rect 580 6306 586 6450
rect 595 6380 608 6450
rect 660 6446 682 6450
rect 653 6424 682 6438
rect 735 6424 751 6438
rect 789 6434 795 6436
rect 802 6434 910 6450
rect 917 6434 923 6436
rect 931 6434 946 6450
rect 1012 6444 1031 6447
rect 653 6422 751 6424
rect 778 6422 946 6434
rect 961 6424 977 6438
rect 1012 6425 1034 6444
rect 1044 6438 1060 6439
rect 1043 6436 1060 6438
rect 1044 6431 1060 6436
rect 1034 6424 1040 6425
rect 1043 6424 1072 6431
rect 961 6423 1072 6424
rect 961 6422 1078 6423
rect 637 6414 688 6422
rect 735 6414 769 6422
rect 637 6402 662 6414
rect 669 6402 688 6414
rect 742 6412 769 6414
rect 778 6412 999 6422
rect 1034 6419 1040 6422
rect 742 6408 999 6412
rect 637 6394 688 6402
rect 735 6394 999 6408
rect 1043 6414 1078 6422
rect 589 6346 608 6380
rect 653 6386 682 6394
rect 653 6380 670 6386
rect 653 6378 687 6380
rect 735 6378 751 6394
rect 752 6384 960 6394
rect 961 6384 977 6394
rect 1025 6390 1040 6405
rect 1043 6402 1044 6414
rect 1051 6402 1078 6414
rect 1043 6394 1078 6402
rect 1043 6393 1072 6394
rect 763 6380 977 6384
rect 778 6378 977 6380
rect 1012 6380 1025 6390
rect 1043 6380 1060 6393
rect 1012 6378 1060 6380
rect 654 6374 687 6378
rect 650 6372 687 6374
rect 650 6371 717 6372
rect 650 6366 681 6371
rect 687 6366 717 6371
rect 650 6362 717 6366
rect 623 6359 717 6362
rect 623 6352 672 6359
rect 623 6346 653 6352
rect 672 6347 677 6352
rect 589 6330 669 6346
rect 681 6338 717 6359
rect 778 6354 967 6378
rect 1012 6377 1059 6378
rect 1025 6372 1059 6377
rect 793 6351 967 6354
rect 786 6348 967 6351
rect 995 6371 1059 6372
rect 589 6328 608 6330
rect 623 6328 657 6330
rect 589 6312 669 6328
rect 589 6306 608 6312
rect 305 6280 408 6290
rect 259 6278 408 6280
rect 429 6278 464 6290
rect 98 6276 260 6278
rect 110 6256 129 6276
rect 144 6274 174 6276
rect -7 6248 34 6256
rect 116 6252 129 6256
rect 181 6260 260 6276
rect 292 6276 464 6278
rect 292 6260 371 6276
rect 378 6274 408 6276
rect -1 6238 28 6248
rect 43 6238 73 6252
rect 116 6238 159 6252
rect 181 6248 371 6260
rect 436 6256 442 6276
rect 166 6238 196 6248
rect 197 6238 355 6248
rect 359 6238 389 6248
rect 393 6238 423 6252
rect 451 6238 464 6276
rect 536 6290 565 6306
rect 579 6290 608 6306
rect 623 6296 653 6312
rect 681 6290 687 6338
rect 690 6332 709 6338
rect 724 6332 754 6340
rect 690 6324 754 6332
rect 690 6308 770 6324
rect 786 6317 848 6348
rect 864 6317 926 6348
rect 995 6346 1044 6371
rect 1059 6346 1089 6362
rect 958 6332 988 6340
rect 995 6338 1105 6346
rect 958 6324 1003 6332
rect 690 6306 709 6308
rect 724 6306 770 6308
rect 690 6290 770 6306
rect 797 6304 832 6317
rect 873 6314 910 6317
rect 873 6312 915 6314
rect 802 6301 832 6304
rect 811 6297 818 6301
rect 818 6296 819 6297
rect 777 6290 787 6296
rect 536 6282 571 6290
rect 536 6256 537 6282
rect 544 6256 571 6282
rect 479 6238 509 6252
rect 536 6248 571 6256
rect 573 6282 614 6290
rect 573 6256 588 6282
rect 595 6256 614 6282
rect 678 6278 709 6290
rect 724 6278 827 6290
rect 839 6280 865 6306
rect 880 6301 910 6312
rect 942 6308 1004 6324
rect 942 6306 988 6308
rect 942 6290 1004 6306
rect 1016 6290 1022 6338
rect 1025 6330 1105 6338
rect 1025 6328 1044 6330
rect 1059 6328 1093 6330
rect 1025 6312 1105 6328
rect 1025 6290 1044 6312
rect 1059 6296 1089 6312
rect 1117 6306 1123 6380
rect 1126 6306 1145 6450
rect 1160 6306 1166 6450
rect 1175 6380 1188 6450
rect 1240 6446 1262 6450
rect 1233 6424 1262 6438
rect 1315 6424 1331 6438
rect 1369 6434 1375 6436
rect 1382 6434 1490 6450
rect 1497 6434 1503 6436
rect 1511 6434 1526 6450
rect 1592 6444 1611 6447
rect 1233 6422 1331 6424
rect 1358 6422 1526 6434
rect 1541 6424 1557 6438
rect 1592 6425 1614 6444
rect 1624 6438 1640 6439
rect 1623 6436 1640 6438
rect 1624 6431 1640 6436
rect 1614 6424 1620 6425
rect 1623 6424 1652 6431
rect 1541 6423 1652 6424
rect 1541 6422 1658 6423
rect 1217 6414 1268 6422
rect 1315 6414 1349 6422
rect 1217 6402 1242 6414
rect 1249 6402 1268 6414
rect 1322 6412 1349 6414
rect 1358 6412 1579 6422
rect 1614 6419 1620 6422
rect 1322 6408 1579 6412
rect 1217 6394 1268 6402
rect 1315 6394 1579 6408
rect 1623 6414 1658 6422
rect 1169 6346 1188 6380
rect 1233 6386 1262 6394
rect 1233 6380 1250 6386
rect 1233 6378 1267 6380
rect 1315 6378 1331 6394
rect 1332 6384 1540 6394
rect 1541 6384 1557 6394
rect 1605 6390 1620 6405
rect 1623 6402 1624 6414
rect 1631 6402 1658 6414
rect 1623 6394 1658 6402
rect 1623 6393 1652 6394
rect 1343 6380 1557 6384
rect 1358 6378 1557 6380
rect 1592 6380 1605 6390
rect 1623 6380 1640 6393
rect 1592 6378 1640 6380
rect 1234 6374 1267 6378
rect 1230 6372 1267 6374
rect 1230 6371 1297 6372
rect 1230 6366 1261 6371
rect 1267 6366 1297 6371
rect 1230 6362 1297 6366
rect 1203 6359 1297 6362
rect 1203 6352 1252 6359
rect 1203 6346 1233 6352
rect 1252 6347 1257 6352
rect 1169 6330 1249 6346
rect 1261 6338 1297 6359
rect 1358 6354 1547 6378
rect 1592 6377 1639 6378
rect 1605 6372 1639 6377
rect 1373 6351 1547 6354
rect 1366 6348 1547 6351
rect 1575 6371 1639 6372
rect 1169 6328 1188 6330
rect 1203 6328 1237 6330
rect 1169 6312 1249 6328
rect 1169 6306 1188 6312
rect 885 6280 988 6290
rect 839 6278 988 6280
rect 1009 6278 1044 6290
rect 678 6276 840 6278
rect 690 6256 709 6276
rect 724 6274 754 6276
rect 573 6248 614 6256
rect 696 6252 709 6256
rect 761 6260 840 6276
rect 872 6276 1044 6278
rect 872 6260 951 6276
rect 958 6274 988 6276
rect 536 6238 565 6248
rect 579 6238 608 6248
rect 623 6238 653 6252
rect 696 6238 739 6252
rect 761 6248 951 6260
rect 1016 6256 1022 6276
rect 746 6238 776 6248
rect 777 6238 935 6248
rect 939 6238 969 6248
rect 973 6238 1003 6252
rect 1031 6238 1044 6276
rect 1116 6290 1145 6306
rect 1159 6290 1188 6306
rect 1203 6296 1233 6312
rect 1261 6290 1267 6338
rect 1270 6332 1289 6338
rect 1304 6332 1334 6340
rect 1270 6324 1334 6332
rect 1270 6308 1350 6324
rect 1366 6317 1428 6348
rect 1444 6317 1506 6348
rect 1575 6346 1624 6371
rect 1639 6346 1669 6362
rect 1538 6332 1568 6340
rect 1575 6338 1685 6346
rect 1538 6324 1583 6332
rect 1270 6306 1289 6308
rect 1304 6306 1350 6308
rect 1270 6290 1350 6306
rect 1377 6304 1412 6317
rect 1453 6314 1490 6317
rect 1453 6312 1495 6314
rect 1382 6301 1412 6304
rect 1391 6297 1398 6301
rect 1398 6296 1399 6297
rect 1357 6290 1367 6296
rect 1116 6282 1151 6290
rect 1116 6256 1117 6282
rect 1124 6256 1151 6282
rect 1059 6238 1089 6252
rect 1116 6248 1151 6256
rect 1153 6282 1194 6290
rect 1153 6256 1168 6282
rect 1175 6256 1194 6282
rect 1258 6278 1289 6290
rect 1304 6278 1407 6290
rect 1419 6280 1445 6306
rect 1460 6301 1490 6312
rect 1522 6308 1584 6324
rect 1522 6306 1568 6308
rect 1522 6290 1584 6306
rect 1596 6290 1602 6338
rect 1605 6330 1685 6338
rect 1605 6328 1624 6330
rect 1639 6328 1673 6330
rect 1605 6312 1685 6328
rect 1605 6290 1624 6312
rect 1639 6296 1669 6312
rect 1697 6306 1703 6380
rect 1706 6306 1725 6450
rect 1740 6306 1746 6450
rect 1755 6380 1768 6450
rect 1820 6446 1842 6450
rect 1813 6424 1842 6438
rect 1895 6424 1911 6438
rect 1949 6434 1955 6436
rect 1962 6434 2070 6450
rect 2077 6434 2083 6436
rect 2091 6434 2106 6450
rect 2172 6444 2191 6447
rect 1813 6422 1911 6424
rect 1938 6422 2106 6434
rect 2121 6424 2137 6438
rect 2172 6425 2194 6444
rect 2204 6438 2220 6439
rect 2203 6436 2220 6438
rect 2204 6431 2220 6436
rect 2194 6424 2200 6425
rect 2203 6424 2232 6431
rect 2121 6423 2232 6424
rect 2121 6422 2238 6423
rect 1797 6414 1848 6422
rect 1895 6414 1929 6422
rect 1797 6402 1822 6414
rect 1829 6402 1848 6414
rect 1902 6412 1929 6414
rect 1938 6412 2159 6422
rect 2194 6419 2200 6422
rect 1902 6408 2159 6412
rect 1797 6394 1848 6402
rect 1895 6394 2159 6408
rect 2203 6414 2238 6422
rect 1749 6346 1768 6380
rect 1813 6386 1842 6394
rect 1813 6380 1830 6386
rect 1813 6378 1847 6380
rect 1895 6378 1911 6394
rect 1912 6384 2120 6394
rect 2121 6384 2137 6394
rect 2185 6390 2200 6405
rect 2203 6402 2204 6414
rect 2211 6402 2238 6414
rect 2203 6394 2238 6402
rect 2203 6393 2232 6394
rect 1923 6380 2137 6384
rect 1938 6378 2137 6380
rect 2172 6380 2185 6390
rect 2203 6380 2220 6393
rect 2172 6378 2220 6380
rect 1814 6374 1847 6378
rect 1810 6372 1847 6374
rect 1810 6371 1877 6372
rect 1810 6366 1841 6371
rect 1847 6366 1877 6371
rect 1810 6362 1877 6366
rect 1783 6359 1877 6362
rect 1783 6352 1832 6359
rect 1783 6346 1813 6352
rect 1832 6347 1837 6352
rect 1749 6330 1829 6346
rect 1841 6338 1877 6359
rect 1938 6354 2127 6378
rect 2172 6377 2219 6378
rect 2185 6372 2219 6377
rect 1953 6351 2127 6354
rect 1946 6348 2127 6351
rect 2155 6371 2219 6372
rect 1749 6328 1768 6330
rect 1783 6328 1817 6330
rect 1749 6312 1829 6328
rect 1749 6306 1768 6312
rect 1465 6280 1568 6290
rect 1419 6278 1568 6280
rect 1589 6278 1624 6290
rect 1258 6276 1420 6278
rect 1270 6256 1289 6276
rect 1304 6274 1334 6276
rect 1153 6248 1194 6256
rect 1276 6252 1289 6256
rect 1341 6260 1420 6276
rect 1452 6276 1624 6278
rect 1452 6260 1531 6276
rect 1538 6274 1568 6276
rect 1116 6238 1145 6248
rect 1159 6238 1188 6248
rect 1203 6238 1233 6252
rect 1276 6238 1319 6252
rect 1341 6248 1531 6260
rect 1596 6256 1602 6276
rect 1326 6238 1356 6248
rect 1357 6238 1515 6248
rect 1519 6238 1549 6248
rect 1553 6238 1583 6252
rect 1611 6238 1624 6276
rect 1696 6290 1725 6306
rect 1739 6290 1768 6306
rect 1783 6296 1813 6312
rect 1841 6290 1847 6338
rect 1850 6332 1869 6338
rect 1884 6332 1914 6340
rect 1850 6324 1914 6332
rect 1850 6308 1930 6324
rect 1946 6317 2008 6348
rect 2024 6317 2086 6348
rect 2155 6346 2204 6371
rect 2219 6346 2249 6362
rect 2118 6332 2148 6340
rect 2155 6338 2265 6346
rect 2118 6324 2163 6332
rect 1850 6306 1869 6308
rect 1884 6306 1930 6308
rect 1850 6290 1930 6306
rect 1957 6304 1992 6317
rect 2033 6314 2070 6317
rect 2033 6312 2075 6314
rect 1962 6301 1992 6304
rect 1971 6297 1978 6301
rect 1978 6296 1979 6297
rect 1937 6290 1947 6296
rect 1696 6282 1731 6290
rect 1696 6256 1697 6282
rect 1704 6256 1731 6282
rect 1639 6238 1669 6252
rect 1696 6248 1731 6256
rect 1733 6282 1774 6290
rect 1733 6256 1748 6282
rect 1755 6256 1774 6282
rect 1838 6278 1869 6290
rect 1884 6278 1987 6290
rect 1999 6280 2025 6306
rect 2040 6301 2070 6312
rect 2102 6308 2164 6324
rect 2102 6306 2148 6308
rect 2102 6290 2164 6306
rect 2176 6290 2182 6338
rect 2185 6330 2265 6338
rect 2185 6328 2204 6330
rect 2219 6328 2253 6330
rect 2185 6312 2265 6328
rect 2185 6290 2204 6312
rect 2219 6296 2249 6312
rect 2277 6306 2283 6380
rect 2286 6306 2305 6450
rect 2320 6306 2326 6450
rect 2335 6380 2348 6450
rect 2400 6446 2422 6450
rect 2393 6424 2422 6438
rect 2475 6424 2491 6438
rect 2529 6434 2535 6436
rect 2542 6434 2650 6450
rect 2657 6434 2663 6436
rect 2671 6434 2686 6450
rect 2752 6444 2771 6447
rect 2393 6422 2491 6424
rect 2518 6422 2686 6434
rect 2701 6424 2717 6438
rect 2752 6425 2774 6444
rect 2784 6438 2800 6439
rect 2783 6436 2800 6438
rect 2784 6431 2800 6436
rect 2774 6424 2780 6425
rect 2783 6424 2812 6431
rect 2701 6423 2812 6424
rect 2701 6422 2818 6423
rect 2377 6414 2428 6422
rect 2475 6414 2509 6422
rect 2377 6402 2402 6414
rect 2409 6402 2428 6414
rect 2482 6412 2509 6414
rect 2518 6412 2739 6422
rect 2774 6419 2780 6422
rect 2482 6408 2739 6412
rect 2377 6394 2428 6402
rect 2475 6394 2739 6408
rect 2783 6414 2818 6422
rect 2329 6346 2348 6380
rect 2393 6386 2422 6394
rect 2393 6380 2410 6386
rect 2393 6378 2427 6380
rect 2475 6378 2491 6394
rect 2492 6384 2700 6394
rect 2701 6384 2717 6394
rect 2765 6390 2780 6405
rect 2783 6402 2784 6414
rect 2791 6402 2818 6414
rect 2783 6394 2818 6402
rect 2783 6393 2812 6394
rect 2503 6380 2717 6384
rect 2518 6378 2717 6380
rect 2752 6380 2765 6390
rect 2783 6380 2800 6393
rect 2752 6378 2800 6380
rect 2394 6374 2427 6378
rect 2390 6372 2427 6374
rect 2390 6371 2457 6372
rect 2390 6366 2421 6371
rect 2427 6366 2457 6371
rect 2390 6362 2457 6366
rect 2363 6359 2457 6362
rect 2363 6352 2412 6359
rect 2363 6346 2393 6352
rect 2412 6347 2417 6352
rect 2329 6330 2409 6346
rect 2421 6338 2457 6359
rect 2518 6354 2707 6378
rect 2752 6377 2799 6378
rect 2765 6372 2799 6377
rect 2533 6351 2707 6354
rect 2526 6348 2707 6351
rect 2735 6371 2799 6372
rect 2329 6328 2348 6330
rect 2363 6328 2397 6330
rect 2329 6312 2409 6328
rect 2329 6306 2348 6312
rect 2045 6280 2148 6290
rect 1999 6278 2148 6280
rect 2169 6278 2204 6290
rect 1838 6276 2000 6278
rect 1850 6256 1869 6276
rect 1884 6274 1914 6276
rect 1733 6248 1774 6256
rect 1856 6252 1869 6256
rect 1921 6260 2000 6276
rect 2032 6276 2204 6278
rect 2032 6260 2111 6276
rect 2118 6274 2148 6276
rect 1696 6238 1725 6248
rect 1739 6238 1768 6248
rect 1783 6238 1813 6252
rect 1856 6238 1899 6252
rect 1921 6248 2111 6260
rect 2176 6256 2182 6276
rect 1906 6238 1936 6248
rect 1937 6238 2095 6248
rect 2099 6238 2129 6248
rect 2133 6238 2163 6252
rect 2191 6238 2204 6276
rect 2276 6290 2305 6306
rect 2319 6290 2348 6306
rect 2363 6296 2393 6312
rect 2421 6290 2427 6338
rect 2430 6332 2449 6338
rect 2464 6332 2494 6340
rect 2430 6324 2494 6332
rect 2430 6308 2510 6324
rect 2526 6317 2588 6348
rect 2604 6317 2666 6348
rect 2735 6346 2784 6371
rect 2799 6346 2829 6362
rect 2698 6332 2728 6340
rect 2735 6338 2845 6346
rect 2698 6324 2743 6332
rect 2430 6306 2449 6308
rect 2464 6306 2510 6308
rect 2430 6290 2510 6306
rect 2537 6304 2572 6317
rect 2613 6314 2650 6317
rect 2613 6312 2655 6314
rect 2542 6301 2572 6304
rect 2551 6297 2558 6301
rect 2558 6296 2559 6297
rect 2517 6290 2527 6296
rect 2276 6282 2311 6290
rect 2276 6256 2277 6282
rect 2284 6256 2311 6282
rect 2219 6238 2249 6252
rect 2276 6248 2311 6256
rect 2313 6282 2354 6290
rect 2313 6256 2328 6282
rect 2335 6256 2354 6282
rect 2418 6278 2449 6290
rect 2464 6278 2567 6290
rect 2579 6280 2605 6306
rect 2620 6301 2650 6312
rect 2682 6308 2744 6324
rect 2682 6306 2728 6308
rect 2682 6290 2744 6306
rect 2756 6290 2762 6338
rect 2765 6330 2845 6338
rect 2765 6328 2784 6330
rect 2799 6328 2833 6330
rect 2765 6312 2845 6328
rect 2765 6290 2784 6312
rect 2799 6296 2829 6312
rect 2857 6306 2863 6380
rect 2866 6306 2885 6450
rect 2900 6306 2906 6450
rect 2915 6380 2928 6450
rect 2980 6446 3002 6450
rect 2973 6424 3002 6438
rect 3055 6424 3071 6438
rect 3109 6434 3115 6436
rect 3122 6434 3230 6450
rect 3237 6434 3243 6436
rect 3251 6434 3266 6450
rect 3332 6444 3351 6447
rect 2973 6422 3071 6424
rect 3098 6422 3266 6434
rect 3281 6424 3297 6438
rect 3332 6425 3354 6444
rect 3364 6438 3380 6439
rect 3363 6436 3380 6438
rect 3364 6431 3380 6436
rect 3354 6424 3360 6425
rect 3363 6424 3392 6431
rect 3281 6423 3392 6424
rect 3281 6422 3398 6423
rect 2957 6414 3008 6422
rect 3055 6414 3089 6422
rect 2957 6402 2982 6414
rect 2989 6402 3008 6414
rect 3062 6412 3089 6414
rect 3098 6412 3319 6422
rect 3354 6419 3360 6422
rect 3062 6408 3319 6412
rect 2957 6394 3008 6402
rect 3055 6394 3319 6408
rect 3363 6414 3398 6422
rect 2909 6346 2928 6380
rect 2973 6386 3002 6394
rect 2973 6380 2990 6386
rect 2973 6378 3007 6380
rect 3055 6378 3071 6394
rect 3072 6384 3280 6394
rect 3281 6384 3297 6394
rect 3345 6390 3360 6405
rect 3363 6402 3364 6414
rect 3371 6402 3398 6414
rect 3363 6394 3398 6402
rect 3363 6393 3392 6394
rect 3083 6380 3297 6384
rect 3098 6378 3297 6380
rect 3332 6380 3345 6390
rect 3363 6380 3380 6393
rect 3332 6378 3380 6380
rect 2974 6374 3007 6378
rect 2970 6372 3007 6374
rect 2970 6371 3037 6372
rect 2970 6366 3001 6371
rect 3007 6366 3037 6371
rect 2970 6362 3037 6366
rect 2943 6359 3037 6362
rect 2943 6352 2992 6359
rect 2943 6346 2973 6352
rect 2992 6347 2997 6352
rect 2909 6330 2989 6346
rect 3001 6338 3037 6359
rect 3098 6354 3287 6378
rect 3332 6377 3379 6378
rect 3345 6372 3379 6377
rect 3113 6351 3287 6354
rect 3106 6348 3287 6351
rect 3315 6371 3379 6372
rect 2909 6328 2928 6330
rect 2943 6328 2977 6330
rect 2909 6312 2989 6328
rect 2909 6306 2928 6312
rect 2625 6280 2728 6290
rect 2579 6278 2728 6280
rect 2749 6278 2784 6290
rect 2418 6276 2580 6278
rect 2430 6256 2449 6276
rect 2464 6274 2494 6276
rect 2313 6248 2354 6256
rect 2436 6252 2449 6256
rect 2501 6260 2580 6276
rect 2612 6276 2784 6278
rect 2612 6260 2691 6276
rect 2698 6274 2728 6276
rect 2276 6238 2305 6248
rect 2319 6238 2348 6248
rect 2363 6238 2393 6252
rect 2436 6238 2479 6252
rect 2501 6248 2691 6260
rect 2756 6256 2762 6276
rect 2486 6238 2516 6248
rect 2517 6238 2675 6248
rect 2679 6238 2709 6248
rect 2713 6238 2743 6252
rect 2771 6238 2784 6276
rect 2856 6290 2885 6306
rect 2899 6290 2928 6306
rect 2943 6296 2973 6312
rect 3001 6290 3007 6338
rect 3010 6332 3029 6338
rect 3044 6332 3074 6340
rect 3010 6324 3074 6332
rect 3010 6308 3090 6324
rect 3106 6317 3168 6348
rect 3184 6317 3246 6348
rect 3315 6346 3364 6371
rect 3379 6346 3409 6362
rect 3278 6332 3308 6340
rect 3315 6338 3425 6346
rect 3278 6324 3323 6332
rect 3010 6306 3029 6308
rect 3044 6306 3090 6308
rect 3010 6290 3090 6306
rect 3117 6304 3152 6317
rect 3193 6314 3230 6317
rect 3193 6312 3235 6314
rect 3122 6301 3152 6304
rect 3131 6297 3138 6301
rect 3138 6296 3139 6297
rect 3097 6290 3107 6296
rect 2856 6282 2891 6290
rect 2856 6256 2857 6282
rect 2864 6256 2891 6282
rect 2799 6238 2829 6252
rect 2856 6248 2891 6256
rect 2893 6282 2934 6290
rect 2893 6256 2908 6282
rect 2915 6256 2934 6282
rect 2998 6278 3029 6290
rect 3044 6278 3147 6290
rect 3159 6280 3185 6306
rect 3200 6301 3230 6312
rect 3262 6308 3324 6324
rect 3262 6306 3308 6308
rect 3262 6290 3324 6306
rect 3336 6290 3342 6338
rect 3345 6330 3425 6338
rect 3345 6328 3364 6330
rect 3379 6328 3413 6330
rect 3345 6312 3425 6328
rect 3345 6290 3364 6312
rect 3379 6296 3409 6312
rect 3437 6306 3443 6380
rect 3446 6306 3465 6450
rect 3480 6306 3486 6450
rect 3495 6380 3508 6450
rect 3560 6446 3582 6450
rect 3553 6424 3582 6438
rect 3635 6424 3651 6438
rect 3689 6434 3695 6436
rect 3702 6434 3810 6450
rect 3817 6434 3823 6436
rect 3831 6434 3846 6450
rect 3912 6444 3931 6447
rect 3553 6422 3651 6424
rect 3678 6422 3846 6434
rect 3861 6424 3877 6438
rect 3912 6425 3934 6444
rect 3944 6438 3960 6439
rect 3943 6436 3960 6438
rect 3944 6431 3960 6436
rect 3934 6424 3940 6425
rect 3943 6424 3972 6431
rect 3861 6423 3972 6424
rect 3861 6422 3978 6423
rect 3537 6414 3588 6422
rect 3635 6414 3669 6422
rect 3537 6402 3562 6414
rect 3569 6402 3588 6414
rect 3642 6412 3669 6414
rect 3678 6412 3899 6422
rect 3934 6419 3940 6422
rect 3642 6408 3899 6412
rect 3537 6394 3588 6402
rect 3635 6394 3899 6408
rect 3943 6414 3978 6422
rect 3489 6346 3508 6380
rect 3553 6386 3582 6394
rect 3553 6380 3570 6386
rect 3553 6378 3587 6380
rect 3635 6378 3651 6394
rect 3652 6384 3860 6394
rect 3861 6384 3877 6394
rect 3925 6390 3940 6405
rect 3943 6402 3944 6414
rect 3951 6402 3978 6414
rect 3943 6394 3978 6402
rect 3943 6393 3972 6394
rect 3663 6380 3877 6384
rect 3678 6378 3877 6380
rect 3912 6380 3925 6390
rect 3943 6380 3960 6393
rect 3912 6378 3960 6380
rect 3554 6374 3587 6378
rect 3550 6372 3587 6374
rect 3550 6371 3617 6372
rect 3550 6366 3581 6371
rect 3587 6366 3617 6371
rect 3550 6362 3617 6366
rect 3523 6359 3617 6362
rect 3523 6352 3572 6359
rect 3523 6346 3553 6352
rect 3572 6347 3577 6352
rect 3489 6330 3569 6346
rect 3581 6338 3617 6359
rect 3678 6354 3867 6378
rect 3912 6377 3959 6378
rect 3925 6372 3959 6377
rect 3693 6351 3867 6354
rect 3686 6348 3867 6351
rect 3895 6371 3959 6372
rect 3489 6328 3508 6330
rect 3523 6328 3557 6330
rect 3489 6312 3569 6328
rect 3489 6306 3508 6312
rect 3205 6280 3308 6290
rect 3159 6278 3308 6280
rect 3329 6278 3364 6290
rect 2998 6276 3160 6278
rect 3010 6256 3029 6276
rect 3044 6274 3074 6276
rect 2893 6248 2934 6256
rect 3016 6252 3029 6256
rect 3081 6260 3160 6276
rect 3192 6276 3364 6278
rect 3192 6260 3271 6276
rect 3278 6274 3308 6276
rect 2856 6238 2885 6248
rect 2899 6238 2928 6248
rect 2943 6238 2973 6252
rect 3016 6238 3059 6252
rect 3081 6248 3271 6260
rect 3336 6256 3342 6276
rect 3066 6238 3096 6248
rect 3097 6238 3255 6248
rect 3259 6238 3289 6248
rect 3293 6238 3323 6252
rect 3351 6238 3364 6276
rect 3436 6290 3465 6306
rect 3479 6290 3508 6306
rect 3523 6296 3553 6312
rect 3581 6290 3587 6338
rect 3590 6332 3609 6338
rect 3624 6332 3654 6340
rect 3590 6324 3654 6332
rect 3590 6308 3670 6324
rect 3686 6317 3748 6348
rect 3764 6317 3826 6348
rect 3895 6346 3944 6371
rect 3959 6346 3989 6362
rect 3858 6332 3888 6340
rect 3895 6338 4005 6346
rect 3858 6324 3903 6332
rect 3590 6306 3609 6308
rect 3624 6306 3670 6308
rect 3590 6290 3670 6306
rect 3697 6304 3732 6317
rect 3773 6314 3810 6317
rect 3773 6312 3815 6314
rect 3702 6301 3732 6304
rect 3711 6297 3718 6301
rect 3718 6296 3719 6297
rect 3677 6290 3687 6296
rect 3436 6282 3471 6290
rect 3436 6256 3437 6282
rect 3444 6256 3471 6282
rect 3379 6238 3409 6252
rect 3436 6248 3471 6256
rect 3473 6282 3514 6290
rect 3473 6256 3488 6282
rect 3495 6256 3514 6282
rect 3578 6278 3609 6290
rect 3624 6278 3727 6290
rect 3739 6280 3765 6306
rect 3780 6301 3810 6312
rect 3842 6308 3904 6324
rect 3842 6306 3888 6308
rect 3842 6290 3904 6306
rect 3916 6290 3922 6338
rect 3925 6330 4005 6338
rect 3925 6328 3944 6330
rect 3959 6328 3993 6330
rect 3925 6312 4005 6328
rect 3925 6290 3944 6312
rect 3959 6296 3989 6312
rect 4017 6306 4023 6380
rect 4026 6306 4045 6450
rect 4060 6306 4066 6450
rect 4075 6380 4088 6450
rect 4140 6446 4162 6450
rect 4133 6424 4162 6438
rect 4215 6424 4231 6438
rect 4269 6434 4275 6436
rect 4282 6434 4390 6450
rect 4397 6434 4403 6436
rect 4411 6434 4426 6450
rect 4492 6444 4511 6447
rect 4133 6422 4231 6424
rect 4258 6422 4426 6434
rect 4441 6424 4457 6438
rect 4492 6425 4514 6444
rect 4524 6438 4540 6439
rect 4523 6436 4540 6438
rect 4524 6431 4540 6436
rect 4514 6424 4520 6425
rect 4523 6424 4552 6431
rect 4441 6423 4552 6424
rect 4441 6422 4558 6423
rect 4117 6414 4168 6422
rect 4215 6414 4249 6422
rect 4117 6402 4142 6414
rect 4149 6402 4168 6414
rect 4222 6412 4249 6414
rect 4258 6412 4479 6422
rect 4514 6419 4520 6422
rect 4222 6408 4479 6412
rect 4117 6394 4168 6402
rect 4215 6394 4479 6408
rect 4523 6414 4558 6422
rect 4069 6346 4088 6380
rect 4133 6386 4162 6394
rect 4133 6380 4150 6386
rect 4133 6378 4167 6380
rect 4215 6378 4231 6394
rect 4232 6384 4440 6394
rect 4441 6384 4457 6394
rect 4505 6390 4520 6405
rect 4523 6402 4524 6414
rect 4531 6402 4558 6414
rect 4523 6394 4558 6402
rect 4523 6393 4552 6394
rect 4243 6380 4457 6384
rect 4258 6378 4457 6380
rect 4492 6380 4505 6390
rect 4523 6380 4540 6393
rect 4492 6378 4540 6380
rect 4134 6374 4167 6378
rect 4130 6372 4167 6374
rect 4130 6371 4197 6372
rect 4130 6366 4161 6371
rect 4167 6366 4197 6371
rect 4130 6362 4197 6366
rect 4103 6359 4197 6362
rect 4103 6352 4152 6359
rect 4103 6346 4133 6352
rect 4152 6347 4157 6352
rect 4069 6330 4149 6346
rect 4161 6338 4197 6359
rect 4258 6354 4447 6378
rect 4492 6377 4539 6378
rect 4505 6372 4539 6377
rect 4273 6351 4447 6354
rect 4266 6348 4447 6351
rect 4475 6371 4539 6372
rect 4069 6328 4088 6330
rect 4103 6328 4137 6330
rect 4069 6312 4149 6328
rect 4069 6306 4088 6312
rect 3785 6280 3888 6290
rect 3739 6278 3888 6280
rect 3909 6278 3944 6290
rect 3578 6276 3740 6278
rect 3590 6256 3609 6276
rect 3624 6274 3654 6276
rect 3473 6248 3514 6256
rect 3596 6252 3609 6256
rect 3661 6260 3740 6276
rect 3772 6276 3944 6278
rect 3772 6260 3851 6276
rect 3858 6274 3888 6276
rect 3436 6238 3465 6248
rect 3479 6238 3508 6248
rect 3523 6238 3553 6252
rect 3596 6238 3639 6252
rect 3661 6248 3851 6260
rect 3916 6256 3922 6276
rect 3646 6238 3676 6248
rect 3677 6238 3835 6248
rect 3839 6238 3869 6248
rect 3873 6238 3903 6252
rect 3931 6238 3944 6276
rect 4016 6290 4045 6306
rect 4059 6290 4088 6306
rect 4103 6296 4133 6312
rect 4161 6290 4167 6338
rect 4170 6332 4189 6338
rect 4204 6332 4234 6340
rect 4170 6324 4234 6332
rect 4170 6308 4250 6324
rect 4266 6317 4328 6348
rect 4344 6317 4406 6348
rect 4475 6346 4524 6371
rect 4539 6346 4569 6362
rect 4438 6332 4468 6340
rect 4475 6338 4585 6346
rect 4438 6324 4483 6332
rect 4170 6306 4189 6308
rect 4204 6306 4250 6308
rect 4170 6290 4250 6306
rect 4277 6304 4312 6317
rect 4353 6314 4390 6317
rect 4353 6312 4395 6314
rect 4282 6301 4312 6304
rect 4291 6297 4298 6301
rect 4298 6296 4299 6297
rect 4257 6290 4267 6296
rect 4016 6282 4051 6290
rect 4016 6256 4017 6282
rect 4024 6256 4051 6282
rect 3959 6238 3989 6252
rect 4016 6248 4051 6256
rect 4053 6282 4094 6290
rect 4053 6256 4068 6282
rect 4075 6256 4094 6282
rect 4158 6278 4189 6290
rect 4204 6278 4307 6290
rect 4319 6280 4345 6306
rect 4360 6301 4390 6312
rect 4422 6308 4484 6324
rect 4422 6306 4468 6308
rect 4422 6290 4484 6306
rect 4496 6290 4502 6338
rect 4505 6330 4585 6338
rect 4505 6328 4524 6330
rect 4539 6328 4573 6330
rect 4505 6312 4585 6328
rect 4505 6290 4524 6312
rect 4539 6296 4569 6312
rect 4597 6306 4603 6380
rect 4606 6306 4625 6450
rect 4640 6306 4646 6450
rect 4655 6380 4668 6450
rect 4720 6446 4742 6450
rect 4713 6424 4742 6438
rect 4795 6424 4811 6438
rect 4849 6434 4855 6436
rect 4862 6434 4970 6450
rect 4977 6434 4983 6436
rect 4991 6434 5006 6450
rect 5072 6444 5091 6447
rect 4713 6422 4811 6424
rect 4838 6422 5006 6434
rect 5021 6424 5037 6438
rect 5072 6425 5094 6444
rect 5104 6438 5120 6439
rect 5103 6436 5120 6438
rect 5104 6431 5120 6436
rect 5094 6424 5100 6425
rect 5103 6424 5132 6431
rect 5021 6423 5132 6424
rect 5021 6422 5138 6423
rect 4697 6414 4748 6422
rect 4795 6414 4829 6422
rect 4697 6402 4722 6414
rect 4729 6402 4748 6414
rect 4802 6412 4829 6414
rect 4838 6412 5059 6422
rect 5094 6419 5100 6422
rect 4802 6408 5059 6412
rect 4697 6394 4748 6402
rect 4795 6394 5059 6408
rect 5103 6414 5138 6422
rect 4649 6346 4668 6380
rect 4713 6386 4742 6394
rect 4713 6380 4730 6386
rect 4713 6378 4747 6380
rect 4795 6378 4811 6394
rect 4812 6384 5020 6394
rect 5021 6384 5037 6394
rect 5085 6390 5100 6405
rect 5103 6402 5104 6414
rect 5111 6402 5138 6414
rect 5103 6394 5138 6402
rect 5103 6393 5132 6394
rect 4823 6380 5037 6384
rect 4838 6378 5037 6380
rect 5072 6380 5085 6390
rect 5103 6380 5120 6393
rect 5072 6378 5120 6380
rect 4714 6374 4747 6378
rect 4710 6372 4747 6374
rect 4710 6371 4777 6372
rect 4710 6366 4741 6371
rect 4747 6366 4777 6371
rect 4710 6362 4777 6366
rect 4683 6359 4777 6362
rect 4683 6352 4732 6359
rect 4683 6346 4713 6352
rect 4732 6347 4737 6352
rect 4649 6330 4729 6346
rect 4741 6338 4777 6359
rect 4838 6354 5027 6378
rect 5072 6377 5119 6378
rect 5085 6372 5119 6377
rect 4853 6351 5027 6354
rect 4846 6348 5027 6351
rect 5055 6371 5119 6372
rect 4649 6328 4668 6330
rect 4683 6328 4717 6330
rect 4649 6312 4729 6328
rect 4649 6306 4668 6312
rect 4365 6280 4468 6290
rect 4319 6278 4468 6280
rect 4489 6278 4524 6290
rect 4158 6276 4320 6278
rect 4170 6256 4189 6276
rect 4204 6274 4234 6276
rect 4053 6248 4094 6256
rect 4176 6252 4189 6256
rect 4241 6260 4320 6276
rect 4352 6276 4524 6278
rect 4352 6260 4431 6276
rect 4438 6274 4468 6276
rect 4016 6238 4045 6248
rect 4059 6238 4088 6248
rect 4103 6238 4133 6252
rect 4176 6238 4219 6252
rect 4241 6248 4431 6260
rect 4496 6256 4502 6276
rect 4226 6238 4256 6248
rect 4257 6238 4415 6248
rect 4419 6238 4449 6248
rect 4453 6238 4483 6252
rect 4511 6238 4524 6276
rect 4596 6290 4625 6306
rect 4639 6290 4668 6306
rect 4683 6296 4713 6312
rect 4741 6290 4747 6338
rect 4750 6332 4769 6338
rect 4784 6332 4814 6340
rect 4750 6324 4814 6332
rect 4750 6308 4830 6324
rect 4846 6317 4908 6348
rect 4924 6317 4986 6348
rect 5055 6346 5104 6371
rect 5119 6346 5149 6362
rect 5018 6332 5048 6340
rect 5055 6338 5165 6346
rect 5018 6324 5063 6332
rect 4750 6306 4769 6308
rect 4784 6306 4830 6308
rect 4750 6290 4830 6306
rect 4857 6304 4892 6317
rect 4933 6314 4970 6317
rect 4933 6312 4975 6314
rect 4862 6301 4892 6304
rect 4871 6297 4878 6301
rect 4878 6296 4879 6297
rect 4837 6290 4847 6296
rect 4596 6282 4631 6290
rect 4596 6256 4597 6282
rect 4604 6256 4631 6282
rect 4539 6238 4569 6252
rect 4596 6248 4631 6256
rect 4633 6282 4674 6290
rect 4633 6256 4648 6282
rect 4655 6256 4674 6282
rect 4738 6278 4769 6290
rect 4784 6278 4887 6290
rect 4899 6280 4925 6306
rect 4940 6301 4970 6312
rect 5002 6308 5064 6324
rect 5002 6306 5048 6308
rect 5002 6290 5064 6306
rect 5076 6290 5082 6338
rect 5085 6330 5165 6338
rect 5085 6328 5104 6330
rect 5119 6328 5153 6330
rect 5085 6312 5165 6328
rect 5085 6290 5104 6312
rect 5119 6296 5149 6312
rect 5177 6306 5183 6380
rect 5186 6306 5205 6450
rect 5220 6306 5226 6450
rect 5235 6380 5248 6450
rect 5300 6446 5322 6450
rect 5293 6424 5322 6438
rect 5375 6424 5391 6438
rect 5429 6434 5435 6436
rect 5442 6434 5550 6450
rect 5557 6434 5563 6436
rect 5571 6434 5586 6450
rect 5652 6444 5671 6447
rect 5293 6422 5391 6424
rect 5418 6422 5586 6434
rect 5601 6424 5617 6438
rect 5652 6425 5674 6444
rect 5684 6438 5700 6439
rect 5683 6436 5700 6438
rect 5684 6431 5700 6436
rect 5674 6424 5680 6425
rect 5683 6424 5712 6431
rect 5601 6423 5712 6424
rect 5601 6422 5718 6423
rect 5277 6414 5328 6422
rect 5375 6414 5409 6422
rect 5277 6402 5302 6414
rect 5309 6402 5328 6414
rect 5382 6412 5409 6414
rect 5418 6412 5639 6422
rect 5674 6419 5680 6422
rect 5382 6408 5639 6412
rect 5277 6394 5328 6402
rect 5375 6394 5639 6408
rect 5683 6414 5718 6422
rect 5229 6346 5248 6380
rect 5293 6386 5322 6394
rect 5293 6380 5310 6386
rect 5293 6378 5327 6380
rect 5375 6378 5391 6394
rect 5392 6384 5600 6394
rect 5601 6384 5617 6394
rect 5665 6390 5680 6405
rect 5683 6402 5684 6414
rect 5691 6402 5718 6414
rect 5683 6394 5718 6402
rect 5683 6393 5712 6394
rect 5403 6380 5617 6384
rect 5418 6378 5617 6380
rect 5652 6380 5665 6390
rect 5683 6380 5700 6393
rect 5652 6378 5700 6380
rect 5294 6374 5327 6378
rect 5290 6372 5327 6374
rect 5290 6371 5357 6372
rect 5290 6366 5321 6371
rect 5327 6366 5357 6371
rect 5290 6362 5357 6366
rect 5263 6359 5357 6362
rect 5263 6352 5312 6359
rect 5263 6346 5293 6352
rect 5312 6347 5317 6352
rect 5229 6330 5309 6346
rect 5321 6338 5357 6359
rect 5418 6354 5607 6378
rect 5652 6377 5699 6378
rect 5665 6372 5699 6377
rect 5433 6351 5607 6354
rect 5426 6348 5607 6351
rect 5635 6371 5699 6372
rect 5229 6328 5248 6330
rect 5263 6328 5297 6330
rect 5229 6312 5309 6328
rect 5229 6306 5248 6312
rect 4945 6280 5048 6290
rect 4899 6278 5048 6280
rect 5069 6278 5104 6290
rect 4738 6276 4900 6278
rect 4750 6256 4769 6276
rect 4784 6274 4814 6276
rect 4633 6248 4674 6256
rect 4756 6252 4769 6256
rect 4821 6260 4900 6276
rect 4932 6276 5104 6278
rect 4932 6260 5011 6276
rect 5018 6274 5048 6276
rect 4596 6238 4625 6248
rect 4639 6238 4668 6248
rect 4683 6238 4713 6252
rect 4756 6238 4799 6252
rect 4821 6248 5011 6260
rect 5076 6256 5082 6276
rect 4806 6238 4836 6248
rect 4837 6238 4995 6248
rect 4999 6238 5029 6248
rect 5033 6238 5063 6252
rect 5091 6238 5104 6276
rect 5176 6290 5205 6306
rect 5219 6290 5248 6306
rect 5263 6296 5293 6312
rect 5321 6290 5327 6338
rect 5330 6332 5349 6338
rect 5364 6332 5394 6340
rect 5330 6324 5394 6332
rect 5330 6308 5410 6324
rect 5426 6317 5488 6348
rect 5504 6317 5566 6348
rect 5635 6346 5684 6371
rect 5699 6346 5729 6362
rect 5598 6332 5628 6340
rect 5635 6338 5745 6346
rect 5598 6324 5643 6332
rect 5330 6306 5349 6308
rect 5364 6306 5410 6308
rect 5330 6290 5410 6306
rect 5437 6304 5472 6317
rect 5513 6314 5550 6317
rect 5513 6312 5555 6314
rect 5442 6301 5472 6304
rect 5451 6297 5458 6301
rect 5458 6296 5459 6297
rect 5417 6290 5427 6296
rect 5176 6282 5211 6290
rect 5176 6256 5177 6282
rect 5184 6256 5211 6282
rect 5119 6238 5149 6252
rect 5176 6248 5211 6256
rect 5213 6282 5254 6290
rect 5213 6256 5228 6282
rect 5235 6256 5254 6282
rect 5318 6278 5349 6290
rect 5364 6278 5467 6290
rect 5479 6280 5505 6306
rect 5520 6301 5550 6312
rect 5582 6308 5644 6324
rect 5582 6306 5628 6308
rect 5582 6290 5644 6306
rect 5656 6290 5662 6338
rect 5665 6330 5745 6338
rect 5665 6328 5684 6330
rect 5699 6328 5733 6330
rect 5665 6312 5745 6328
rect 5665 6290 5684 6312
rect 5699 6296 5729 6312
rect 5757 6306 5763 6380
rect 5766 6306 5785 6450
rect 5800 6306 5806 6450
rect 5815 6380 5828 6450
rect 5880 6446 5902 6450
rect 5873 6424 5902 6438
rect 5955 6424 5971 6438
rect 6009 6434 6015 6436
rect 6022 6434 6130 6450
rect 6137 6434 6143 6436
rect 6151 6434 6166 6450
rect 6232 6444 6251 6447
rect 5873 6422 5971 6424
rect 5998 6422 6166 6434
rect 6181 6424 6197 6438
rect 6232 6425 6254 6444
rect 6264 6438 6280 6439
rect 6263 6436 6280 6438
rect 6264 6431 6280 6436
rect 6254 6424 6260 6425
rect 6263 6424 6292 6431
rect 6181 6423 6292 6424
rect 6181 6422 6298 6423
rect 5857 6414 5908 6422
rect 5955 6414 5989 6422
rect 5857 6402 5882 6414
rect 5889 6402 5908 6414
rect 5962 6412 5989 6414
rect 5998 6412 6219 6422
rect 6254 6419 6260 6422
rect 5962 6408 6219 6412
rect 5857 6394 5908 6402
rect 5955 6394 6219 6408
rect 6263 6414 6298 6422
rect 5809 6346 5828 6380
rect 5873 6386 5902 6394
rect 5873 6380 5890 6386
rect 5873 6378 5907 6380
rect 5955 6378 5971 6394
rect 5972 6384 6180 6394
rect 6181 6384 6197 6394
rect 6245 6390 6260 6405
rect 6263 6402 6264 6414
rect 6271 6402 6298 6414
rect 6263 6394 6298 6402
rect 6263 6393 6292 6394
rect 5983 6380 6197 6384
rect 5998 6378 6197 6380
rect 6232 6380 6245 6390
rect 6263 6380 6280 6393
rect 6232 6378 6280 6380
rect 5874 6374 5907 6378
rect 5870 6372 5907 6374
rect 5870 6371 5937 6372
rect 5870 6366 5901 6371
rect 5907 6366 5937 6371
rect 5870 6362 5937 6366
rect 5843 6359 5937 6362
rect 5843 6352 5892 6359
rect 5843 6346 5873 6352
rect 5892 6347 5897 6352
rect 5809 6330 5889 6346
rect 5901 6338 5937 6359
rect 5998 6354 6187 6378
rect 6232 6377 6279 6378
rect 6245 6372 6279 6377
rect 6013 6351 6187 6354
rect 6006 6348 6187 6351
rect 6215 6371 6279 6372
rect 5809 6328 5828 6330
rect 5843 6328 5877 6330
rect 5809 6312 5889 6328
rect 5809 6306 5828 6312
rect 5525 6280 5628 6290
rect 5479 6278 5628 6280
rect 5649 6278 5684 6290
rect 5318 6276 5480 6278
rect 5330 6256 5349 6276
rect 5364 6274 5394 6276
rect 5213 6248 5254 6256
rect 5336 6252 5349 6256
rect 5401 6260 5480 6276
rect 5512 6276 5684 6278
rect 5512 6260 5591 6276
rect 5598 6274 5628 6276
rect 5176 6238 5205 6248
rect 5219 6238 5248 6248
rect 5263 6238 5293 6252
rect 5336 6238 5379 6252
rect 5401 6248 5591 6260
rect 5656 6256 5662 6276
rect 5386 6238 5416 6248
rect 5417 6238 5575 6248
rect 5579 6238 5609 6248
rect 5613 6238 5643 6252
rect 5671 6238 5684 6276
rect 5756 6290 5785 6306
rect 5799 6290 5828 6306
rect 5843 6296 5873 6312
rect 5901 6290 5907 6338
rect 5910 6332 5929 6338
rect 5944 6332 5974 6340
rect 5910 6324 5974 6332
rect 5910 6308 5990 6324
rect 6006 6317 6068 6348
rect 6084 6317 6146 6348
rect 6215 6346 6264 6371
rect 6279 6346 6309 6362
rect 6178 6332 6208 6340
rect 6215 6338 6325 6346
rect 6178 6324 6223 6332
rect 5910 6306 5929 6308
rect 5944 6306 5990 6308
rect 5910 6290 5990 6306
rect 6017 6304 6052 6317
rect 6093 6314 6130 6317
rect 6093 6312 6135 6314
rect 6022 6301 6052 6304
rect 6031 6297 6038 6301
rect 6038 6296 6039 6297
rect 5997 6290 6007 6296
rect 5756 6282 5791 6290
rect 5756 6256 5757 6282
rect 5764 6256 5791 6282
rect 5699 6238 5729 6252
rect 5756 6248 5791 6256
rect 5793 6282 5834 6290
rect 5793 6256 5808 6282
rect 5815 6256 5834 6282
rect 5898 6278 5929 6290
rect 5944 6278 6047 6290
rect 6059 6280 6085 6306
rect 6100 6301 6130 6312
rect 6162 6308 6224 6324
rect 6162 6306 6208 6308
rect 6162 6290 6224 6306
rect 6236 6290 6242 6338
rect 6245 6330 6325 6338
rect 6245 6328 6264 6330
rect 6279 6328 6313 6330
rect 6245 6312 6325 6328
rect 6245 6290 6264 6312
rect 6279 6296 6309 6312
rect 6337 6306 6343 6380
rect 6346 6306 6365 6450
rect 6380 6306 6386 6450
rect 6395 6380 6408 6450
rect 6460 6446 6482 6450
rect 6453 6424 6482 6438
rect 6535 6424 6551 6438
rect 6589 6434 6595 6436
rect 6602 6434 6710 6450
rect 6717 6434 6723 6436
rect 6731 6434 6746 6450
rect 6812 6444 6831 6447
rect 6453 6422 6551 6424
rect 6578 6422 6746 6434
rect 6761 6424 6777 6438
rect 6812 6425 6834 6444
rect 6844 6438 6860 6439
rect 6843 6436 6860 6438
rect 6844 6431 6860 6436
rect 6834 6424 6840 6425
rect 6843 6424 6872 6431
rect 6761 6423 6872 6424
rect 6761 6422 6878 6423
rect 6437 6414 6488 6422
rect 6535 6414 6569 6422
rect 6437 6402 6462 6414
rect 6469 6402 6488 6414
rect 6542 6412 6569 6414
rect 6578 6412 6799 6422
rect 6834 6419 6840 6422
rect 6542 6408 6799 6412
rect 6437 6394 6488 6402
rect 6535 6394 6799 6408
rect 6843 6414 6878 6422
rect 6389 6346 6408 6380
rect 6453 6386 6482 6394
rect 6453 6380 6470 6386
rect 6453 6378 6487 6380
rect 6535 6378 6551 6394
rect 6552 6384 6760 6394
rect 6761 6384 6777 6394
rect 6825 6390 6840 6405
rect 6843 6402 6844 6414
rect 6851 6402 6878 6414
rect 6843 6394 6878 6402
rect 6843 6393 6872 6394
rect 6563 6380 6777 6384
rect 6578 6378 6777 6380
rect 6812 6380 6825 6390
rect 6843 6380 6860 6393
rect 6812 6378 6860 6380
rect 6454 6374 6487 6378
rect 6450 6372 6487 6374
rect 6450 6371 6517 6372
rect 6450 6366 6481 6371
rect 6487 6366 6517 6371
rect 6450 6362 6517 6366
rect 6423 6359 6517 6362
rect 6423 6352 6472 6359
rect 6423 6346 6453 6352
rect 6472 6347 6477 6352
rect 6389 6330 6469 6346
rect 6481 6338 6517 6359
rect 6578 6354 6767 6378
rect 6812 6377 6859 6378
rect 6825 6372 6859 6377
rect 6593 6351 6767 6354
rect 6586 6348 6767 6351
rect 6795 6371 6859 6372
rect 6389 6328 6408 6330
rect 6423 6328 6457 6330
rect 6389 6312 6469 6328
rect 6389 6306 6408 6312
rect 6105 6280 6208 6290
rect 6059 6278 6208 6280
rect 6229 6278 6264 6290
rect 5898 6276 6060 6278
rect 5910 6256 5929 6276
rect 5944 6274 5974 6276
rect 5793 6248 5834 6256
rect 5916 6252 5929 6256
rect 5981 6260 6060 6276
rect 6092 6276 6264 6278
rect 6092 6260 6171 6276
rect 6178 6274 6208 6276
rect 5756 6238 5785 6248
rect 5799 6238 5828 6248
rect 5843 6238 5873 6252
rect 5916 6238 5959 6252
rect 5981 6248 6171 6260
rect 6236 6256 6242 6276
rect 5966 6238 5996 6248
rect 5997 6238 6155 6248
rect 6159 6238 6189 6248
rect 6193 6238 6223 6252
rect 6251 6238 6264 6276
rect 6336 6290 6365 6306
rect 6379 6290 6408 6306
rect 6423 6296 6453 6312
rect 6481 6290 6487 6338
rect 6490 6332 6509 6338
rect 6524 6332 6554 6340
rect 6490 6324 6554 6332
rect 6490 6308 6570 6324
rect 6586 6317 6648 6348
rect 6664 6317 6726 6348
rect 6795 6346 6844 6371
rect 6859 6346 6889 6362
rect 6758 6332 6788 6340
rect 6795 6338 6905 6346
rect 6758 6324 6803 6332
rect 6490 6306 6509 6308
rect 6524 6306 6570 6308
rect 6490 6290 6570 6306
rect 6597 6304 6632 6317
rect 6673 6314 6710 6317
rect 6673 6312 6715 6314
rect 6602 6301 6632 6304
rect 6611 6297 6618 6301
rect 6618 6296 6619 6297
rect 6577 6290 6587 6296
rect 6336 6282 6371 6290
rect 6336 6256 6337 6282
rect 6344 6256 6371 6282
rect 6279 6238 6309 6252
rect 6336 6248 6371 6256
rect 6373 6282 6414 6290
rect 6373 6256 6388 6282
rect 6395 6256 6414 6282
rect 6478 6278 6509 6290
rect 6524 6278 6627 6290
rect 6639 6280 6665 6306
rect 6680 6301 6710 6312
rect 6742 6308 6804 6324
rect 6742 6306 6788 6308
rect 6742 6290 6804 6306
rect 6816 6290 6822 6338
rect 6825 6330 6905 6338
rect 6825 6328 6844 6330
rect 6859 6328 6893 6330
rect 6825 6312 6905 6328
rect 6825 6290 6844 6312
rect 6859 6296 6889 6312
rect 6917 6306 6923 6380
rect 6926 6306 6945 6450
rect 6960 6306 6966 6450
rect 6975 6380 6988 6450
rect 7040 6446 7062 6450
rect 7033 6424 7062 6438
rect 7115 6424 7131 6438
rect 7169 6434 7175 6436
rect 7182 6434 7290 6450
rect 7297 6434 7303 6436
rect 7311 6434 7326 6450
rect 7392 6444 7411 6447
rect 7033 6422 7131 6424
rect 7158 6422 7326 6434
rect 7341 6424 7357 6438
rect 7392 6425 7414 6444
rect 7424 6438 7440 6439
rect 7423 6436 7440 6438
rect 7424 6431 7440 6436
rect 7414 6424 7420 6425
rect 7423 6424 7452 6431
rect 7341 6423 7452 6424
rect 7341 6422 7458 6423
rect 7017 6414 7068 6422
rect 7115 6414 7149 6422
rect 7017 6402 7042 6414
rect 7049 6402 7068 6414
rect 7122 6412 7149 6414
rect 7158 6412 7379 6422
rect 7414 6419 7420 6422
rect 7122 6408 7379 6412
rect 7017 6394 7068 6402
rect 7115 6394 7379 6408
rect 7423 6414 7458 6422
rect 6969 6346 6988 6380
rect 7033 6386 7062 6394
rect 7033 6380 7050 6386
rect 7033 6378 7067 6380
rect 7115 6378 7131 6394
rect 7132 6384 7340 6394
rect 7341 6384 7357 6394
rect 7405 6390 7420 6405
rect 7423 6402 7424 6414
rect 7431 6402 7458 6414
rect 7423 6394 7458 6402
rect 7423 6393 7452 6394
rect 7143 6380 7357 6384
rect 7158 6378 7357 6380
rect 7392 6380 7405 6390
rect 7423 6380 7440 6393
rect 7392 6378 7440 6380
rect 7034 6374 7067 6378
rect 7030 6372 7067 6374
rect 7030 6371 7097 6372
rect 7030 6366 7061 6371
rect 7067 6366 7097 6371
rect 7030 6362 7097 6366
rect 7003 6359 7097 6362
rect 7003 6352 7052 6359
rect 7003 6346 7033 6352
rect 7052 6347 7057 6352
rect 6969 6330 7049 6346
rect 7061 6338 7097 6359
rect 7158 6354 7347 6378
rect 7392 6377 7439 6378
rect 7405 6372 7439 6377
rect 7173 6351 7347 6354
rect 7166 6348 7347 6351
rect 7375 6371 7439 6372
rect 6969 6328 6988 6330
rect 7003 6328 7037 6330
rect 6969 6312 7049 6328
rect 6969 6306 6988 6312
rect 6685 6280 6788 6290
rect 6639 6278 6788 6280
rect 6809 6278 6844 6290
rect 6478 6276 6640 6278
rect 6490 6256 6509 6276
rect 6524 6274 6554 6276
rect 6373 6248 6414 6256
rect 6496 6252 6509 6256
rect 6561 6260 6640 6276
rect 6672 6276 6844 6278
rect 6672 6260 6751 6276
rect 6758 6274 6788 6276
rect 6336 6238 6365 6248
rect 6379 6238 6408 6248
rect 6423 6238 6453 6252
rect 6496 6238 6539 6252
rect 6561 6248 6751 6260
rect 6816 6256 6822 6276
rect 6546 6238 6576 6248
rect 6577 6238 6735 6248
rect 6739 6238 6769 6248
rect 6773 6238 6803 6252
rect 6831 6238 6844 6276
rect 6916 6290 6945 6306
rect 6959 6290 6988 6306
rect 7003 6296 7033 6312
rect 7061 6290 7067 6338
rect 7070 6332 7089 6338
rect 7104 6332 7134 6340
rect 7070 6324 7134 6332
rect 7070 6308 7150 6324
rect 7166 6317 7228 6348
rect 7244 6317 7306 6348
rect 7375 6346 7424 6371
rect 7439 6346 7469 6362
rect 7338 6332 7368 6340
rect 7375 6338 7485 6346
rect 7338 6324 7383 6332
rect 7070 6306 7089 6308
rect 7104 6306 7150 6308
rect 7070 6290 7150 6306
rect 7177 6304 7212 6317
rect 7253 6314 7290 6317
rect 7253 6312 7295 6314
rect 7182 6301 7212 6304
rect 7191 6297 7198 6301
rect 7198 6296 7199 6297
rect 7157 6290 7167 6296
rect 6916 6282 6951 6290
rect 6916 6256 6917 6282
rect 6924 6256 6951 6282
rect 6859 6238 6889 6252
rect 6916 6248 6951 6256
rect 6953 6282 6994 6290
rect 6953 6256 6968 6282
rect 6975 6256 6994 6282
rect 7058 6278 7089 6290
rect 7104 6278 7207 6290
rect 7219 6280 7245 6306
rect 7260 6301 7290 6312
rect 7322 6308 7384 6324
rect 7322 6306 7368 6308
rect 7322 6290 7384 6306
rect 7396 6290 7402 6338
rect 7405 6330 7485 6338
rect 7405 6328 7424 6330
rect 7439 6328 7473 6330
rect 7405 6312 7485 6328
rect 7405 6290 7424 6312
rect 7439 6296 7469 6312
rect 7497 6306 7503 6380
rect 7506 6306 7525 6450
rect 7540 6306 7546 6450
rect 7555 6380 7568 6450
rect 7613 6428 7614 6438
rect 7629 6428 7642 6438
rect 7613 6424 7642 6428
rect 7647 6424 7677 6450
rect 7695 6436 7711 6438
rect 7783 6436 7836 6450
rect 7784 6434 7848 6436
rect 7891 6434 7906 6450
rect 7955 6447 7985 6450
rect 7955 6444 7991 6447
rect 7921 6436 7937 6438
rect 7695 6424 7710 6428
rect 7613 6422 7710 6424
rect 7738 6422 7906 6434
rect 7922 6424 7937 6428
rect 7955 6425 7994 6444
rect 8013 6438 8020 6439
rect 8019 6431 8020 6438
rect 8003 6428 8004 6431
rect 8019 6428 8032 6431
rect 7955 6424 7985 6425
rect 7994 6424 8000 6425
rect 8003 6424 8032 6428
rect 7922 6423 8032 6424
rect 7922 6422 8038 6423
rect 7597 6414 7648 6422
rect 7597 6402 7622 6414
rect 7629 6402 7648 6414
rect 7679 6414 7729 6422
rect 7679 6406 7695 6414
rect 7702 6412 7729 6414
rect 7738 6412 7959 6422
rect 7702 6402 7959 6412
rect 7988 6414 8038 6422
rect 7988 6405 8004 6414
rect 7597 6394 7648 6402
rect 7695 6394 7959 6402
rect 7985 6402 8004 6405
rect 8011 6402 8038 6414
rect 7985 6394 8038 6402
rect 7549 6346 7568 6380
rect 7613 6386 7614 6394
rect 7629 6386 7642 6394
rect 7613 6378 7629 6386
rect 7610 6371 7629 6374
rect 7610 6362 7632 6371
rect 7583 6352 7632 6362
rect 7583 6346 7613 6352
rect 7632 6347 7637 6352
rect 7549 6330 7629 6346
rect 7647 6338 7677 6394
rect 7712 6384 7920 6394
rect 7955 6390 8000 6394
rect 8003 6393 8004 6394
rect 8019 6393 8032 6394
rect 7738 6354 7927 6384
rect 7753 6351 7927 6354
rect 7746 6348 7927 6351
rect 7549 6328 7568 6330
rect 7583 6328 7617 6330
rect 7549 6312 7629 6328
rect 7656 6324 7669 6338
rect 7684 6324 7700 6340
rect 7746 6335 7757 6348
rect 7549 6306 7568 6312
rect 7265 6280 7368 6290
rect 7219 6278 7368 6280
rect 7389 6278 7424 6290
rect 7058 6276 7220 6278
rect 7070 6256 7089 6276
rect 7104 6274 7134 6276
rect 6953 6248 6994 6256
rect 7076 6252 7089 6256
rect 7141 6260 7220 6276
rect 7252 6276 7424 6278
rect 7252 6260 7331 6276
rect 7338 6274 7368 6276
rect 6916 6238 6945 6248
rect 6959 6238 6988 6248
rect 7003 6238 7033 6252
rect 7076 6238 7119 6252
rect 7141 6248 7331 6260
rect 7396 6256 7402 6276
rect 7126 6238 7156 6248
rect 7157 6238 7315 6248
rect 7319 6238 7349 6248
rect 7353 6238 7383 6252
rect 7411 6238 7424 6276
rect 7496 6290 7525 6306
rect 7539 6290 7568 6306
rect 7583 6290 7613 6312
rect 7656 6308 7718 6324
rect 7746 6317 7757 6333
rect 7762 6328 7772 6348
rect 7782 6328 7796 6348
rect 7799 6335 7808 6348
rect 7824 6335 7833 6348
rect 7762 6317 7796 6328
rect 7799 6317 7808 6333
rect 7824 6317 7833 6333
rect 7840 6328 7850 6348
rect 7860 6328 7874 6348
rect 7875 6335 7886 6348
rect 7840 6317 7874 6328
rect 7875 6317 7886 6333
rect 7932 6324 7948 6340
rect 7955 6338 7985 6390
rect 8019 6386 8020 6393
rect 8004 6378 8020 6386
rect 7991 6346 8004 6365
rect 8019 6346 8049 6362
rect 7991 6330 8065 6346
rect 7991 6328 8004 6330
rect 8019 6328 8053 6330
rect 7656 6306 7669 6308
rect 7684 6306 7718 6308
rect 7656 6290 7718 6306
rect 7762 6301 7778 6304
rect 7840 6301 7870 6312
rect 7918 6308 7964 6324
rect 7991 6312 8065 6328
rect 7918 6306 7952 6308
rect 7917 6290 7964 6306
rect 7991 6290 8004 6312
rect 8019 6290 8049 6312
rect 8076 6290 8077 6306
rect 8092 6290 8105 6450
rect 8135 6346 8148 6450
rect 8193 6428 8194 6438
rect 8209 6428 8222 6438
rect 8193 6424 8222 6428
rect 8227 6424 8257 6450
rect 8275 6436 8291 6438
rect 8363 6436 8416 6450
rect 8364 6434 8428 6436
rect 8471 6434 8486 6450
rect 8535 6447 8565 6450
rect 8535 6444 8571 6447
rect 8501 6436 8517 6438
rect 8275 6424 8290 6428
rect 8193 6422 8290 6424
rect 8318 6422 8486 6434
rect 8502 6424 8517 6428
rect 8535 6425 8574 6444
rect 8593 6438 8600 6439
rect 8599 6431 8600 6438
rect 8583 6428 8584 6431
rect 8599 6428 8612 6431
rect 8535 6424 8565 6425
rect 8574 6424 8580 6425
rect 8583 6424 8612 6428
rect 8502 6423 8612 6424
rect 8502 6422 8618 6423
rect 8177 6414 8228 6422
rect 8177 6402 8202 6414
rect 8209 6402 8228 6414
rect 8259 6414 8309 6422
rect 8259 6406 8275 6414
rect 8282 6412 8309 6414
rect 8318 6412 8539 6422
rect 8282 6402 8539 6412
rect 8568 6414 8618 6422
rect 8568 6405 8584 6414
rect 8177 6394 8228 6402
rect 8275 6394 8539 6402
rect 8565 6402 8584 6405
rect 8591 6402 8618 6414
rect 8565 6394 8618 6402
rect 8193 6386 8194 6394
rect 8209 6386 8222 6394
rect 8193 6378 8209 6386
rect 8190 6371 8209 6374
rect 8190 6362 8212 6371
rect 8163 6352 8212 6362
rect 8163 6346 8193 6352
rect 8212 6347 8217 6352
rect 8135 6330 8209 6346
rect 8227 6338 8257 6394
rect 8292 6384 8500 6394
rect 8535 6390 8580 6394
rect 8583 6393 8584 6394
rect 8599 6393 8612 6394
rect 8318 6354 8507 6384
rect 8333 6351 8507 6354
rect 8326 6348 8507 6351
rect 8135 6328 8148 6330
rect 8163 6328 8197 6330
rect 8135 6312 8209 6328
rect 8236 6324 8249 6338
rect 8264 6324 8280 6340
rect 8326 6335 8337 6348
rect 8119 6290 8120 6306
rect 8135 6290 8148 6312
rect 8163 6290 8193 6312
rect 8236 6308 8298 6324
rect 8326 6317 8337 6333
rect 8342 6328 8352 6348
rect 8362 6328 8376 6348
rect 8379 6335 8388 6348
rect 8404 6335 8413 6348
rect 8342 6317 8376 6328
rect 8379 6317 8388 6333
rect 8404 6317 8413 6333
rect 8420 6328 8430 6348
rect 8440 6328 8454 6348
rect 8455 6335 8466 6348
rect 8420 6317 8454 6328
rect 8455 6317 8466 6333
rect 8512 6324 8528 6340
rect 8535 6338 8565 6390
rect 8599 6386 8600 6393
rect 8584 6378 8600 6386
rect 8571 6346 8584 6365
rect 8599 6346 8629 6362
rect 8571 6330 8645 6346
rect 8571 6328 8584 6330
rect 8599 6328 8633 6330
rect 8236 6306 8249 6308
rect 8264 6306 8298 6308
rect 8236 6290 8298 6306
rect 8342 6301 8358 6304
rect 8420 6301 8450 6312
rect 8498 6308 8544 6324
rect 8571 6312 8645 6328
rect 8498 6306 8532 6308
rect 8497 6290 8544 6306
rect 8571 6290 8584 6312
rect 8599 6290 8629 6312
rect 8656 6290 8657 6306
rect 8672 6290 8685 6450
rect 8715 6346 8728 6450
rect 8773 6428 8774 6438
rect 8789 6428 8802 6438
rect 8773 6424 8802 6428
rect 8807 6424 8837 6450
rect 8855 6436 8871 6438
rect 8943 6436 8996 6450
rect 8944 6434 9008 6436
rect 9051 6434 9066 6450
rect 9115 6447 9145 6450
rect 9115 6444 9151 6447
rect 9081 6436 9097 6438
rect 8855 6424 8870 6428
rect 8773 6422 8870 6424
rect 8898 6422 9066 6434
rect 9082 6424 9097 6428
rect 9115 6425 9154 6444
rect 9173 6438 9180 6439
rect 9179 6431 9180 6438
rect 9163 6428 9164 6431
rect 9179 6428 9192 6431
rect 9115 6424 9145 6425
rect 9154 6424 9160 6425
rect 9163 6424 9192 6428
rect 9082 6423 9192 6424
rect 9082 6422 9198 6423
rect 8757 6414 8808 6422
rect 8757 6402 8782 6414
rect 8789 6402 8808 6414
rect 8839 6414 8889 6422
rect 8839 6406 8855 6414
rect 8862 6412 8889 6414
rect 8898 6412 9119 6422
rect 8862 6402 9119 6412
rect 9148 6414 9198 6422
rect 9148 6405 9164 6414
rect 8757 6394 8808 6402
rect 8855 6394 9119 6402
rect 9145 6402 9164 6405
rect 9171 6402 9198 6414
rect 9145 6394 9198 6402
rect 8773 6386 8774 6394
rect 8789 6386 8802 6394
rect 8773 6378 8789 6386
rect 8770 6371 8789 6374
rect 8770 6362 8792 6371
rect 8743 6352 8792 6362
rect 8743 6346 8773 6352
rect 8792 6347 8797 6352
rect 8715 6330 8789 6346
rect 8807 6338 8837 6394
rect 8872 6384 9080 6394
rect 9115 6390 9160 6394
rect 9163 6393 9164 6394
rect 9179 6393 9192 6394
rect 8898 6354 9087 6384
rect 8913 6351 9087 6354
rect 8906 6348 9087 6351
rect 8715 6328 8728 6330
rect 8743 6328 8777 6330
rect 8715 6312 8789 6328
rect 8816 6324 8829 6338
rect 8844 6324 8860 6340
rect 8906 6335 8917 6348
rect 8699 6290 8700 6306
rect 8715 6290 8728 6312
rect 8743 6290 8773 6312
rect 8816 6308 8878 6324
rect 8906 6317 8917 6333
rect 8922 6328 8932 6348
rect 8942 6328 8956 6348
rect 8959 6335 8968 6348
rect 8984 6335 8993 6348
rect 8922 6317 8956 6328
rect 8959 6317 8968 6333
rect 8984 6317 8993 6333
rect 9000 6328 9010 6348
rect 9020 6328 9034 6348
rect 9035 6335 9046 6348
rect 9000 6317 9034 6328
rect 9035 6317 9046 6333
rect 9092 6324 9108 6340
rect 9115 6338 9145 6390
rect 9179 6386 9180 6393
rect 9164 6378 9180 6386
rect 9151 6346 9164 6365
rect 9179 6346 9209 6362
rect 9151 6330 9225 6346
rect 9151 6328 9164 6330
rect 9179 6328 9213 6330
rect 8816 6306 8829 6308
rect 8844 6306 8878 6308
rect 8816 6290 8878 6306
rect 8922 6301 8938 6304
rect 9000 6301 9030 6312
rect 9078 6308 9124 6324
rect 9151 6312 9225 6328
rect 9078 6306 9112 6308
rect 9077 6290 9124 6306
rect 9151 6290 9164 6312
rect 9179 6290 9209 6312
rect 9236 6290 9237 6306
rect 9252 6290 9265 6450
rect 7496 6282 7531 6290
rect 7496 6256 7497 6282
rect 7504 6256 7531 6282
rect 7439 6238 7469 6252
rect 7496 6248 7531 6256
rect 7533 6282 7574 6290
rect 7533 6256 7548 6282
rect 7555 6256 7574 6282
rect 7638 6278 7700 6290
rect 7712 6278 7787 6290
rect 7845 6278 7920 6290
rect 7932 6278 7963 6290
rect 7969 6278 8004 6290
rect 7638 6276 7800 6278
rect 7533 6248 7574 6256
rect 7656 6252 7669 6276
rect 7684 6274 7699 6276
rect 7496 6238 7525 6248
rect 7539 6238 7568 6248
rect 7583 6238 7613 6252
rect 7656 6238 7699 6252
rect 7723 6249 7730 6256
rect 7733 6252 7800 6276
rect 7832 6276 8004 6278
rect 7802 6254 7830 6258
rect 7832 6254 7912 6276
rect 7933 6274 7948 6276
rect 7802 6252 7912 6254
rect 7733 6248 7912 6252
rect 7706 6238 7736 6248
rect 7738 6238 7891 6248
rect 7899 6238 7929 6248
rect 7933 6238 7963 6252
rect 7991 6238 8004 6276
rect 8076 6282 8111 6290
rect 8076 6256 8077 6282
rect 8084 6256 8111 6282
rect 8019 6238 8049 6252
rect 8076 6248 8111 6256
rect 8113 6282 8154 6290
rect 8113 6256 8128 6282
rect 8135 6256 8154 6282
rect 8218 6278 8280 6290
rect 8292 6278 8367 6290
rect 8425 6278 8500 6290
rect 8512 6278 8543 6290
rect 8549 6278 8584 6290
rect 8218 6276 8380 6278
rect 8113 6248 8154 6256
rect 8236 6252 8249 6276
rect 8264 6274 8279 6276
rect 8076 6238 8077 6248
rect 8092 6238 8105 6248
rect 8119 6238 8120 6248
rect 8135 6238 8148 6248
rect 8163 6238 8193 6252
rect 8236 6238 8279 6252
rect 8303 6249 8310 6256
rect 8313 6252 8380 6276
rect 8412 6276 8584 6278
rect 8382 6254 8410 6258
rect 8412 6254 8492 6276
rect 8513 6274 8528 6276
rect 8382 6252 8492 6254
rect 8313 6248 8492 6252
rect 8286 6238 8316 6248
rect 8318 6238 8471 6248
rect 8479 6238 8509 6248
rect 8513 6238 8543 6252
rect 8571 6238 8584 6276
rect 8656 6282 8691 6290
rect 8656 6256 8657 6282
rect 8664 6256 8691 6282
rect 8599 6238 8629 6252
rect 8656 6248 8691 6256
rect 8693 6282 8734 6290
rect 8693 6256 8708 6282
rect 8715 6256 8734 6282
rect 8798 6278 8860 6290
rect 8872 6278 8947 6290
rect 9005 6278 9080 6290
rect 9092 6278 9123 6290
rect 9129 6278 9164 6290
rect 8798 6276 8960 6278
rect 8693 6248 8734 6256
rect 8816 6252 8829 6276
rect 8844 6274 8859 6276
rect 8656 6238 8657 6248
rect 8672 6238 8685 6248
rect 8699 6238 8700 6248
rect 8715 6238 8728 6248
rect 8743 6238 8773 6252
rect 8816 6238 8859 6252
rect 8883 6249 8890 6256
rect 8893 6252 8960 6276
rect 8992 6276 9164 6278
rect 8962 6254 8990 6258
rect 8992 6254 9072 6276
rect 9093 6274 9108 6276
rect 8962 6252 9072 6254
rect 8893 6248 9072 6252
rect 8866 6238 8896 6248
rect 8898 6238 9051 6248
rect 9059 6238 9089 6248
rect 9093 6238 9123 6252
rect 9151 6238 9164 6276
rect 9236 6282 9271 6290
rect 9236 6256 9237 6282
rect 9244 6256 9271 6282
rect 9179 6238 9209 6252
rect 9236 6248 9271 6256
rect 9236 6238 9237 6248
rect 9252 6238 9265 6248
rect -1 6232 9265 6238
rect 0 6224 9265 6232
rect 15 6194 28 6224
rect 43 6210 73 6224
rect 116 6210 159 6224
rect 166 6210 386 6224
rect 393 6210 423 6224
rect 83 6196 98 6208
rect 117 6196 130 6210
rect 198 6206 351 6210
rect 80 6194 102 6196
rect 180 6194 372 6206
rect 451 6194 464 6224
rect 479 6210 509 6224
rect 546 6194 565 6224
rect 580 6194 586 6224
rect 595 6194 608 6224
rect 623 6210 653 6224
rect 696 6210 739 6224
rect 746 6210 966 6224
rect 973 6210 1003 6224
rect 663 6196 678 6208
rect 697 6196 710 6210
rect 778 6206 931 6210
rect 660 6194 682 6196
rect 760 6194 952 6206
rect 1031 6194 1044 6224
rect 1059 6210 1089 6224
rect 1126 6194 1145 6224
rect 1160 6194 1166 6224
rect 1175 6194 1188 6224
rect 1203 6210 1233 6224
rect 1276 6210 1319 6224
rect 1326 6210 1546 6224
rect 1553 6210 1583 6224
rect 1243 6196 1258 6208
rect 1277 6196 1290 6210
rect 1358 6206 1511 6210
rect 1240 6194 1262 6196
rect 1340 6194 1532 6206
rect 1611 6194 1624 6224
rect 1639 6210 1669 6224
rect 1706 6194 1725 6224
rect 1740 6194 1746 6224
rect 1755 6194 1768 6224
rect 1783 6210 1813 6224
rect 1856 6210 1899 6224
rect 1906 6210 2126 6224
rect 2133 6210 2163 6224
rect 1823 6196 1838 6208
rect 1857 6196 1870 6210
rect 1938 6206 2091 6210
rect 1820 6194 1842 6196
rect 1920 6194 2112 6206
rect 2191 6194 2204 6224
rect 2219 6210 2249 6224
rect 2286 6194 2305 6224
rect 2320 6194 2326 6224
rect 2335 6194 2348 6224
rect 2363 6210 2393 6224
rect 2436 6210 2479 6224
rect 2486 6210 2706 6224
rect 2713 6210 2743 6224
rect 2403 6196 2418 6208
rect 2437 6196 2450 6210
rect 2518 6206 2671 6210
rect 2400 6194 2422 6196
rect 2500 6194 2692 6206
rect 2771 6194 2784 6224
rect 2799 6210 2829 6224
rect 2866 6194 2885 6224
rect 2900 6194 2906 6224
rect 2915 6194 2928 6224
rect 2943 6210 2973 6224
rect 3016 6210 3059 6224
rect 3066 6210 3286 6224
rect 3293 6210 3323 6224
rect 2983 6196 2998 6208
rect 3017 6196 3030 6210
rect 3098 6206 3251 6210
rect 2980 6194 3002 6196
rect 3080 6194 3272 6206
rect 3351 6194 3364 6224
rect 3379 6210 3409 6224
rect 3446 6194 3465 6224
rect 3480 6194 3486 6224
rect 3495 6194 3508 6224
rect 3523 6210 3553 6224
rect 3596 6210 3639 6224
rect 3646 6210 3866 6224
rect 3873 6210 3903 6224
rect 3563 6196 3578 6208
rect 3597 6196 3610 6210
rect 3678 6206 3831 6210
rect 3560 6194 3582 6196
rect 3660 6194 3852 6206
rect 3931 6194 3944 6224
rect 3959 6210 3989 6224
rect 4026 6194 4045 6224
rect 4060 6194 4066 6224
rect 4075 6194 4088 6224
rect 4103 6210 4133 6224
rect 4176 6210 4219 6224
rect 4226 6210 4446 6224
rect 4453 6210 4483 6224
rect 4143 6196 4158 6208
rect 4177 6196 4190 6210
rect 4258 6206 4411 6210
rect 4140 6194 4162 6196
rect 4240 6194 4432 6206
rect 4511 6194 4524 6224
rect 4539 6210 4569 6224
rect 4606 6194 4625 6224
rect 4640 6194 4646 6224
rect 4655 6194 4668 6224
rect 4683 6210 4713 6224
rect 4756 6210 4799 6224
rect 4806 6210 5026 6224
rect 5033 6210 5063 6224
rect 4723 6196 4738 6208
rect 4757 6196 4770 6210
rect 4838 6206 4991 6210
rect 4720 6194 4742 6196
rect 4820 6194 5012 6206
rect 5091 6194 5104 6224
rect 5119 6210 5149 6224
rect 5186 6194 5205 6224
rect 5220 6194 5226 6224
rect 5235 6194 5248 6224
rect 5263 6210 5293 6224
rect 5336 6210 5379 6224
rect 5386 6210 5606 6224
rect 5613 6210 5643 6224
rect 5303 6196 5318 6208
rect 5337 6196 5350 6210
rect 5418 6206 5571 6210
rect 5300 6194 5322 6196
rect 5400 6194 5592 6206
rect 5671 6194 5684 6224
rect 5699 6210 5729 6224
rect 5766 6194 5785 6224
rect 5800 6194 5806 6224
rect 5815 6194 5828 6224
rect 5843 6210 5873 6224
rect 5916 6210 5959 6224
rect 5966 6210 6186 6224
rect 6193 6210 6223 6224
rect 5883 6196 5898 6208
rect 5917 6196 5930 6210
rect 5998 6206 6151 6210
rect 5880 6194 5902 6196
rect 5980 6194 6172 6206
rect 6251 6194 6264 6224
rect 6279 6210 6309 6224
rect 6346 6194 6365 6224
rect 6380 6194 6386 6224
rect 6395 6194 6408 6224
rect 6423 6210 6453 6224
rect 6496 6210 6539 6224
rect 6546 6210 6766 6224
rect 6773 6210 6803 6224
rect 6463 6196 6478 6208
rect 6497 6196 6510 6210
rect 6578 6206 6731 6210
rect 6460 6194 6482 6196
rect 6560 6194 6752 6206
rect 6831 6194 6844 6224
rect 6859 6210 6889 6224
rect 6926 6194 6945 6224
rect 6960 6194 6966 6224
rect 6975 6194 6988 6224
rect 7003 6210 7033 6224
rect 7076 6210 7119 6224
rect 7126 6210 7346 6224
rect 7353 6210 7383 6224
rect 7043 6196 7058 6208
rect 7077 6196 7090 6210
rect 7158 6206 7311 6210
rect 7040 6194 7062 6196
rect 7140 6194 7332 6206
rect 7411 6194 7424 6224
rect 7439 6210 7469 6224
rect 7506 6194 7525 6224
rect 7540 6194 7546 6224
rect 7555 6194 7568 6224
rect 7583 6206 7613 6224
rect 7656 6210 7670 6224
rect 7706 6210 7926 6224
rect 7657 6208 7670 6210
rect 7623 6196 7638 6208
rect 7620 6194 7642 6196
rect 7647 6194 7677 6208
rect 7738 6206 7891 6210
rect 7720 6194 7912 6206
rect 7955 6194 7985 6208
rect 7991 6194 8004 6224
rect 8019 6206 8049 6224
rect 8092 6194 8105 6224
rect 8135 6194 8148 6224
rect 8163 6206 8193 6224
rect 8236 6210 8250 6224
rect 8286 6210 8506 6224
rect 8237 6208 8250 6210
rect 8203 6196 8218 6208
rect 8200 6194 8222 6196
rect 8227 6194 8257 6208
rect 8318 6206 8471 6210
rect 8300 6194 8492 6206
rect 8535 6194 8565 6208
rect 8571 6194 8584 6224
rect 8599 6206 8629 6224
rect 8672 6194 8685 6224
rect 8715 6194 8728 6224
rect 8743 6206 8773 6224
rect 8816 6210 8830 6224
rect 8866 6210 9086 6224
rect 8817 6208 8830 6210
rect 8783 6196 8798 6208
rect 8780 6194 8802 6196
rect 8807 6194 8837 6208
rect 8898 6206 9051 6210
rect 8880 6194 9072 6206
rect 9115 6194 9145 6208
rect 9151 6194 9164 6224
rect 9179 6206 9209 6224
rect 9252 6194 9265 6224
rect 0 6180 9265 6194
rect 15 6110 28 6180
rect 80 6176 102 6180
rect 73 6154 102 6168
rect 155 6154 171 6168
rect 209 6164 215 6166
rect 222 6164 330 6180
rect 337 6164 343 6166
rect 351 6164 366 6180
rect 432 6174 451 6177
rect 73 6152 171 6154
rect 198 6152 366 6164
rect 381 6154 397 6168
rect 432 6155 454 6174
rect 464 6168 480 6169
rect 463 6166 480 6168
rect 464 6161 480 6166
rect 454 6154 460 6155
rect 463 6154 492 6161
rect 381 6153 492 6154
rect 381 6152 498 6153
rect 57 6144 108 6152
rect 155 6144 189 6152
rect 57 6132 82 6144
rect 89 6132 108 6144
rect 162 6142 189 6144
rect 198 6142 419 6152
rect 454 6149 460 6152
rect 162 6138 419 6142
rect 57 6124 108 6132
rect 155 6124 419 6138
rect 463 6144 498 6152
rect 9 6076 28 6110
rect 73 6116 102 6124
rect 73 6110 90 6116
rect 73 6108 107 6110
rect 155 6108 171 6124
rect 172 6114 380 6124
rect 381 6114 397 6124
rect 445 6120 460 6135
rect 463 6132 464 6144
rect 471 6132 498 6144
rect 463 6124 498 6132
rect 463 6123 492 6124
rect 183 6110 397 6114
rect 198 6108 397 6110
rect 432 6110 445 6120
rect 463 6110 480 6123
rect 432 6108 480 6110
rect 74 6104 107 6108
rect 70 6102 107 6104
rect 70 6101 137 6102
rect 70 6096 101 6101
rect 107 6096 137 6101
rect 70 6092 137 6096
rect 43 6089 137 6092
rect 43 6082 92 6089
rect 43 6076 73 6082
rect 92 6077 97 6082
rect 9 6060 89 6076
rect 101 6068 137 6089
rect 198 6084 387 6108
rect 432 6107 479 6108
rect 445 6102 479 6107
rect 213 6081 387 6084
rect 206 6078 387 6081
rect 415 6101 479 6102
rect 9 6058 28 6060
rect 43 6058 77 6060
rect 9 6042 89 6058
rect 9 6036 28 6042
rect -1 6020 28 6036
rect 43 6026 73 6042
rect 101 6020 107 6068
rect 110 6062 129 6068
rect 144 6062 174 6070
rect 110 6054 174 6062
rect 110 6038 190 6054
rect 206 6047 268 6078
rect 284 6047 346 6078
rect 415 6076 464 6101
rect 479 6076 509 6092
rect 378 6062 408 6070
rect 415 6068 525 6076
rect 378 6054 423 6062
rect 110 6036 129 6038
rect 144 6036 190 6038
rect 110 6020 190 6036
rect 217 6034 252 6047
rect 293 6044 330 6047
rect 293 6042 335 6044
rect 222 6031 252 6034
rect 231 6027 238 6031
rect 238 6026 239 6027
rect 197 6020 207 6026
rect -7 6012 34 6020
rect -7 5986 8 6012
rect 15 5986 34 6012
rect 98 6008 129 6020
rect 144 6008 247 6020
rect 259 6010 285 6036
rect 300 6031 330 6042
rect 362 6038 424 6054
rect 362 6036 408 6038
rect 362 6020 424 6036
rect 436 6020 442 6068
rect 445 6060 525 6068
rect 445 6058 464 6060
rect 479 6058 513 6060
rect 445 6042 525 6058
rect 445 6020 464 6042
rect 479 6026 509 6042
rect 537 6036 543 6110
rect 546 6036 565 6180
rect 580 6036 586 6180
rect 595 6110 608 6180
rect 660 6176 682 6180
rect 653 6154 682 6168
rect 735 6154 751 6168
rect 789 6164 795 6166
rect 802 6164 910 6180
rect 917 6164 923 6166
rect 931 6164 946 6180
rect 1012 6174 1031 6177
rect 653 6152 751 6154
rect 778 6152 946 6164
rect 961 6154 977 6168
rect 1012 6155 1034 6174
rect 1044 6168 1060 6169
rect 1043 6166 1060 6168
rect 1044 6161 1060 6166
rect 1034 6154 1040 6155
rect 1043 6154 1072 6161
rect 961 6153 1072 6154
rect 961 6152 1078 6153
rect 637 6144 688 6152
rect 735 6144 769 6152
rect 637 6132 662 6144
rect 669 6132 688 6144
rect 742 6142 769 6144
rect 778 6142 999 6152
rect 1034 6149 1040 6152
rect 742 6138 999 6142
rect 637 6124 688 6132
rect 735 6124 999 6138
rect 1043 6144 1078 6152
rect 589 6076 608 6110
rect 653 6116 682 6124
rect 653 6110 670 6116
rect 653 6108 687 6110
rect 735 6108 751 6124
rect 752 6114 960 6124
rect 961 6114 977 6124
rect 1025 6120 1040 6135
rect 1043 6132 1044 6144
rect 1051 6132 1078 6144
rect 1043 6124 1078 6132
rect 1043 6123 1072 6124
rect 763 6110 977 6114
rect 778 6108 977 6110
rect 1012 6110 1025 6120
rect 1043 6110 1060 6123
rect 1012 6108 1060 6110
rect 654 6104 687 6108
rect 650 6102 687 6104
rect 650 6101 717 6102
rect 650 6096 681 6101
rect 687 6096 717 6101
rect 650 6092 717 6096
rect 623 6089 717 6092
rect 623 6082 672 6089
rect 623 6076 653 6082
rect 672 6077 677 6082
rect 589 6060 669 6076
rect 681 6068 717 6089
rect 778 6084 967 6108
rect 1012 6107 1059 6108
rect 1025 6102 1059 6107
rect 793 6081 967 6084
rect 786 6078 967 6081
rect 995 6101 1059 6102
rect 589 6058 608 6060
rect 623 6058 657 6060
rect 589 6042 669 6058
rect 589 6036 608 6042
rect 305 6010 408 6020
rect 259 6008 408 6010
rect 429 6008 464 6020
rect 98 6006 260 6008
rect 110 5986 129 6006
rect 144 6004 174 6006
rect -7 5978 34 5986
rect 116 5982 129 5986
rect 181 5990 260 6006
rect 292 6006 464 6008
rect 292 5990 371 6006
rect 378 6004 408 6006
rect -1 5968 28 5978
rect 43 5968 73 5982
rect 116 5968 159 5982
rect 181 5978 371 5990
rect 436 5986 442 6006
rect 166 5968 196 5978
rect 197 5968 355 5978
rect 359 5968 389 5978
rect 393 5968 423 5982
rect 451 5968 464 6006
rect 536 6020 565 6036
rect 579 6020 608 6036
rect 623 6026 653 6042
rect 681 6020 687 6068
rect 690 6062 709 6068
rect 724 6062 754 6070
rect 690 6054 754 6062
rect 690 6038 770 6054
rect 786 6047 848 6078
rect 864 6047 926 6078
rect 995 6076 1044 6101
rect 1059 6076 1089 6092
rect 958 6062 988 6070
rect 995 6068 1105 6076
rect 958 6054 1003 6062
rect 690 6036 709 6038
rect 724 6036 770 6038
rect 690 6020 770 6036
rect 797 6034 832 6047
rect 873 6044 910 6047
rect 873 6042 915 6044
rect 802 6031 832 6034
rect 811 6027 818 6031
rect 818 6026 819 6027
rect 777 6020 787 6026
rect 536 6012 571 6020
rect 536 5986 537 6012
rect 544 5986 571 6012
rect 479 5968 509 5982
rect 536 5978 571 5986
rect 573 6012 614 6020
rect 573 5986 588 6012
rect 595 5986 614 6012
rect 678 6008 709 6020
rect 724 6008 827 6020
rect 839 6010 865 6036
rect 880 6031 910 6042
rect 942 6038 1004 6054
rect 942 6036 988 6038
rect 942 6020 1004 6036
rect 1016 6020 1022 6068
rect 1025 6060 1105 6068
rect 1025 6058 1044 6060
rect 1059 6058 1093 6060
rect 1025 6042 1105 6058
rect 1025 6020 1044 6042
rect 1059 6026 1089 6042
rect 1117 6036 1123 6110
rect 1126 6036 1145 6180
rect 1160 6036 1166 6180
rect 1175 6110 1188 6180
rect 1240 6176 1262 6180
rect 1233 6154 1262 6168
rect 1315 6154 1331 6168
rect 1369 6164 1375 6166
rect 1382 6164 1490 6180
rect 1497 6164 1503 6166
rect 1511 6164 1526 6180
rect 1592 6174 1611 6177
rect 1233 6152 1331 6154
rect 1358 6152 1526 6164
rect 1541 6154 1557 6168
rect 1592 6155 1614 6174
rect 1624 6168 1640 6169
rect 1623 6166 1640 6168
rect 1624 6161 1640 6166
rect 1614 6154 1620 6155
rect 1623 6154 1652 6161
rect 1541 6153 1652 6154
rect 1541 6152 1658 6153
rect 1217 6144 1268 6152
rect 1315 6144 1349 6152
rect 1217 6132 1242 6144
rect 1249 6132 1268 6144
rect 1322 6142 1349 6144
rect 1358 6142 1579 6152
rect 1614 6149 1620 6152
rect 1322 6138 1579 6142
rect 1217 6124 1268 6132
rect 1315 6124 1579 6138
rect 1623 6144 1658 6152
rect 1169 6076 1188 6110
rect 1233 6116 1262 6124
rect 1233 6110 1250 6116
rect 1233 6108 1267 6110
rect 1315 6108 1331 6124
rect 1332 6114 1540 6124
rect 1541 6114 1557 6124
rect 1605 6120 1620 6135
rect 1623 6132 1624 6144
rect 1631 6132 1658 6144
rect 1623 6124 1658 6132
rect 1623 6123 1652 6124
rect 1343 6110 1557 6114
rect 1358 6108 1557 6110
rect 1592 6110 1605 6120
rect 1623 6110 1640 6123
rect 1592 6108 1640 6110
rect 1234 6104 1267 6108
rect 1230 6102 1267 6104
rect 1230 6101 1297 6102
rect 1230 6096 1261 6101
rect 1267 6096 1297 6101
rect 1230 6092 1297 6096
rect 1203 6089 1297 6092
rect 1203 6082 1252 6089
rect 1203 6076 1233 6082
rect 1252 6077 1257 6082
rect 1169 6060 1249 6076
rect 1261 6068 1297 6089
rect 1358 6084 1547 6108
rect 1592 6107 1639 6108
rect 1605 6102 1639 6107
rect 1373 6081 1547 6084
rect 1366 6078 1547 6081
rect 1575 6101 1639 6102
rect 1169 6058 1188 6060
rect 1203 6058 1237 6060
rect 1169 6042 1249 6058
rect 1169 6036 1188 6042
rect 885 6010 988 6020
rect 839 6008 988 6010
rect 1009 6008 1044 6020
rect 678 6006 840 6008
rect 690 5986 709 6006
rect 724 6004 754 6006
rect 573 5978 614 5986
rect 696 5982 709 5986
rect 761 5990 840 6006
rect 872 6006 1044 6008
rect 872 5990 951 6006
rect 958 6004 988 6006
rect 536 5968 565 5978
rect 579 5968 608 5978
rect 623 5968 653 5982
rect 696 5968 739 5982
rect 761 5978 951 5990
rect 1016 5986 1022 6006
rect 746 5968 776 5978
rect 777 5968 935 5978
rect 939 5968 969 5978
rect 973 5968 1003 5982
rect 1031 5968 1044 6006
rect 1116 6020 1145 6036
rect 1159 6020 1188 6036
rect 1203 6026 1233 6042
rect 1261 6020 1267 6068
rect 1270 6062 1289 6068
rect 1304 6062 1334 6070
rect 1270 6054 1334 6062
rect 1270 6038 1350 6054
rect 1366 6047 1428 6078
rect 1444 6047 1506 6078
rect 1575 6076 1624 6101
rect 1639 6076 1669 6092
rect 1538 6062 1568 6070
rect 1575 6068 1685 6076
rect 1538 6054 1583 6062
rect 1270 6036 1289 6038
rect 1304 6036 1350 6038
rect 1270 6020 1350 6036
rect 1377 6034 1412 6047
rect 1453 6044 1490 6047
rect 1453 6042 1495 6044
rect 1382 6031 1412 6034
rect 1391 6027 1398 6031
rect 1398 6026 1399 6027
rect 1357 6020 1367 6026
rect 1116 6012 1151 6020
rect 1116 5986 1117 6012
rect 1124 5986 1151 6012
rect 1059 5968 1089 5982
rect 1116 5978 1151 5986
rect 1153 6012 1194 6020
rect 1153 5986 1168 6012
rect 1175 5986 1194 6012
rect 1258 6008 1289 6020
rect 1304 6008 1407 6020
rect 1419 6010 1445 6036
rect 1460 6031 1490 6042
rect 1522 6038 1584 6054
rect 1522 6036 1568 6038
rect 1522 6020 1584 6036
rect 1596 6020 1602 6068
rect 1605 6060 1685 6068
rect 1605 6058 1624 6060
rect 1639 6058 1673 6060
rect 1605 6042 1685 6058
rect 1605 6020 1624 6042
rect 1639 6026 1669 6042
rect 1697 6036 1703 6110
rect 1706 6036 1725 6180
rect 1740 6036 1746 6180
rect 1755 6110 1768 6180
rect 1820 6176 1842 6180
rect 1813 6154 1842 6168
rect 1895 6154 1911 6168
rect 1949 6164 1955 6166
rect 1962 6164 2070 6180
rect 2077 6164 2083 6166
rect 2091 6164 2106 6180
rect 2172 6174 2191 6177
rect 1813 6152 1911 6154
rect 1938 6152 2106 6164
rect 2121 6154 2137 6168
rect 2172 6155 2194 6174
rect 2204 6168 2220 6169
rect 2203 6166 2220 6168
rect 2204 6161 2220 6166
rect 2194 6154 2200 6155
rect 2203 6154 2232 6161
rect 2121 6153 2232 6154
rect 2121 6152 2238 6153
rect 1797 6144 1848 6152
rect 1895 6144 1929 6152
rect 1797 6132 1822 6144
rect 1829 6132 1848 6144
rect 1902 6142 1929 6144
rect 1938 6142 2159 6152
rect 2194 6149 2200 6152
rect 1902 6138 2159 6142
rect 1797 6124 1848 6132
rect 1895 6124 2159 6138
rect 2203 6144 2238 6152
rect 1749 6076 1768 6110
rect 1813 6116 1842 6124
rect 1813 6110 1830 6116
rect 1813 6108 1847 6110
rect 1895 6108 1911 6124
rect 1912 6114 2120 6124
rect 2121 6114 2137 6124
rect 2185 6120 2200 6135
rect 2203 6132 2204 6144
rect 2211 6132 2238 6144
rect 2203 6124 2238 6132
rect 2203 6123 2232 6124
rect 1923 6110 2137 6114
rect 1938 6108 2137 6110
rect 2172 6110 2185 6120
rect 2203 6110 2220 6123
rect 2172 6108 2220 6110
rect 1814 6104 1847 6108
rect 1810 6102 1847 6104
rect 1810 6101 1877 6102
rect 1810 6096 1841 6101
rect 1847 6096 1877 6101
rect 1810 6092 1877 6096
rect 1783 6089 1877 6092
rect 1783 6082 1832 6089
rect 1783 6076 1813 6082
rect 1832 6077 1837 6082
rect 1749 6060 1829 6076
rect 1841 6068 1877 6089
rect 1938 6084 2127 6108
rect 2172 6107 2219 6108
rect 2185 6102 2219 6107
rect 1953 6081 2127 6084
rect 1946 6078 2127 6081
rect 2155 6101 2219 6102
rect 1749 6058 1768 6060
rect 1783 6058 1817 6060
rect 1749 6042 1829 6058
rect 1749 6036 1768 6042
rect 1465 6010 1568 6020
rect 1419 6008 1568 6010
rect 1589 6008 1624 6020
rect 1258 6006 1420 6008
rect 1270 5986 1289 6006
rect 1304 6004 1334 6006
rect 1153 5978 1194 5986
rect 1276 5982 1289 5986
rect 1341 5990 1420 6006
rect 1452 6006 1624 6008
rect 1452 5990 1531 6006
rect 1538 6004 1568 6006
rect 1116 5968 1145 5978
rect 1159 5968 1188 5978
rect 1203 5968 1233 5982
rect 1276 5968 1319 5982
rect 1341 5978 1531 5990
rect 1596 5986 1602 6006
rect 1326 5968 1356 5978
rect 1357 5968 1515 5978
rect 1519 5968 1549 5978
rect 1553 5968 1583 5982
rect 1611 5968 1624 6006
rect 1696 6020 1725 6036
rect 1739 6020 1768 6036
rect 1783 6026 1813 6042
rect 1841 6020 1847 6068
rect 1850 6062 1869 6068
rect 1884 6062 1914 6070
rect 1850 6054 1914 6062
rect 1850 6038 1930 6054
rect 1946 6047 2008 6078
rect 2024 6047 2086 6078
rect 2155 6076 2204 6101
rect 2219 6076 2249 6092
rect 2118 6062 2148 6070
rect 2155 6068 2265 6076
rect 2118 6054 2163 6062
rect 1850 6036 1869 6038
rect 1884 6036 1930 6038
rect 1850 6020 1930 6036
rect 1957 6034 1992 6047
rect 2033 6044 2070 6047
rect 2033 6042 2075 6044
rect 1962 6031 1992 6034
rect 1971 6027 1978 6031
rect 1978 6026 1979 6027
rect 1937 6020 1947 6026
rect 1696 6012 1731 6020
rect 1696 5986 1697 6012
rect 1704 5986 1731 6012
rect 1639 5968 1669 5982
rect 1696 5978 1731 5986
rect 1733 6012 1774 6020
rect 1733 5986 1748 6012
rect 1755 5986 1774 6012
rect 1838 6008 1869 6020
rect 1884 6008 1987 6020
rect 1999 6010 2025 6036
rect 2040 6031 2070 6042
rect 2102 6038 2164 6054
rect 2102 6036 2148 6038
rect 2102 6020 2164 6036
rect 2176 6020 2182 6068
rect 2185 6060 2265 6068
rect 2185 6058 2204 6060
rect 2219 6058 2253 6060
rect 2185 6042 2265 6058
rect 2185 6020 2204 6042
rect 2219 6026 2249 6042
rect 2277 6036 2283 6110
rect 2286 6036 2305 6180
rect 2320 6036 2326 6180
rect 2335 6110 2348 6180
rect 2400 6176 2422 6180
rect 2393 6154 2422 6168
rect 2475 6154 2491 6168
rect 2529 6164 2535 6166
rect 2542 6164 2650 6180
rect 2657 6164 2663 6166
rect 2671 6164 2686 6180
rect 2752 6174 2771 6177
rect 2393 6152 2491 6154
rect 2518 6152 2686 6164
rect 2701 6154 2717 6168
rect 2752 6155 2774 6174
rect 2784 6168 2800 6169
rect 2783 6166 2800 6168
rect 2784 6161 2800 6166
rect 2774 6154 2780 6155
rect 2783 6154 2812 6161
rect 2701 6153 2812 6154
rect 2701 6152 2818 6153
rect 2377 6144 2428 6152
rect 2475 6144 2509 6152
rect 2377 6132 2402 6144
rect 2409 6132 2428 6144
rect 2482 6142 2509 6144
rect 2518 6142 2739 6152
rect 2774 6149 2780 6152
rect 2482 6138 2739 6142
rect 2377 6124 2428 6132
rect 2475 6124 2739 6138
rect 2783 6144 2818 6152
rect 2329 6076 2348 6110
rect 2393 6116 2422 6124
rect 2393 6110 2410 6116
rect 2393 6108 2427 6110
rect 2475 6108 2491 6124
rect 2492 6114 2700 6124
rect 2701 6114 2717 6124
rect 2765 6120 2780 6135
rect 2783 6132 2784 6144
rect 2791 6132 2818 6144
rect 2783 6124 2818 6132
rect 2783 6123 2812 6124
rect 2503 6110 2717 6114
rect 2518 6108 2717 6110
rect 2752 6110 2765 6120
rect 2783 6110 2800 6123
rect 2752 6108 2800 6110
rect 2394 6104 2427 6108
rect 2390 6102 2427 6104
rect 2390 6101 2457 6102
rect 2390 6096 2421 6101
rect 2427 6096 2457 6101
rect 2390 6092 2457 6096
rect 2363 6089 2457 6092
rect 2363 6082 2412 6089
rect 2363 6076 2393 6082
rect 2412 6077 2417 6082
rect 2329 6060 2409 6076
rect 2421 6068 2457 6089
rect 2518 6084 2707 6108
rect 2752 6107 2799 6108
rect 2765 6102 2799 6107
rect 2533 6081 2707 6084
rect 2526 6078 2707 6081
rect 2735 6101 2799 6102
rect 2329 6058 2348 6060
rect 2363 6058 2397 6060
rect 2329 6042 2409 6058
rect 2329 6036 2348 6042
rect 2045 6010 2148 6020
rect 1999 6008 2148 6010
rect 2169 6008 2204 6020
rect 1838 6006 2000 6008
rect 1850 5986 1869 6006
rect 1884 6004 1914 6006
rect 1733 5978 1774 5986
rect 1856 5982 1869 5986
rect 1921 5990 2000 6006
rect 2032 6006 2204 6008
rect 2032 5990 2111 6006
rect 2118 6004 2148 6006
rect 1696 5968 1725 5978
rect 1739 5968 1768 5978
rect 1783 5968 1813 5982
rect 1856 5968 1899 5982
rect 1921 5978 2111 5990
rect 2176 5986 2182 6006
rect 1906 5968 1936 5978
rect 1937 5968 2095 5978
rect 2099 5968 2129 5978
rect 2133 5968 2163 5982
rect 2191 5968 2204 6006
rect 2276 6020 2305 6036
rect 2319 6020 2348 6036
rect 2363 6026 2393 6042
rect 2421 6020 2427 6068
rect 2430 6062 2449 6068
rect 2464 6062 2494 6070
rect 2430 6054 2494 6062
rect 2430 6038 2510 6054
rect 2526 6047 2588 6078
rect 2604 6047 2666 6078
rect 2735 6076 2784 6101
rect 2799 6076 2829 6092
rect 2698 6062 2728 6070
rect 2735 6068 2845 6076
rect 2698 6054 2743 6062
rect 2430 6036 2449 6038
rect 2464 6036 2510 6038
rect 2430 6020 2510 6036
rect 2537 6034 2572 6047
rect 2613 6044 2650 6047
rect 2613 6042 2655 6044
rect 2542 6031 2572 6034
rect 2551 6027 2558 6031
rect 2558 6026 2559 6027
rect 2517 6020 2527 6026
rect 2276 6012 2311 6020
rect 2276 5986 2277 6012
rect 2284 5986 2311 6012
rect 2219 5968 2249 5982
rect 2276 5978 2311 5986
rect 2313 6012 2354 6020
rect 2313 5986 2328 6012
rect 2335 5986 2354 6012
rect 2418 6008 2449 6020
rect 2464 6008 2567 6020
rect 2579 6010 2605 6036
rect 2620 6031 2650 6042
rect 2682 6038 2744 6054
rect 2682 6036 2728 6038
rect 2682 6020 2744 6036
rect 2756 6020 2762 6068
rect 2765 6060 2845 6068
rect 2765 6058 2784 6060
rect 2799 6058 2833 6060
rect 2765 6042 2845 6058
rect 2765 6020 2784 6042
rect 2799 6026 2829 6042
rect 2857 6036 2863 6110
rect 2866 6036 2885 6180
rect 2900 6036 2906 6180
rect 2915 6110 2928 6180
rect 2980 6176 3002 6180
rect 2973 6154 3002 6168
rect 3055 6154 3071 6168
rect 3109 6164 3115 6166
rect 3122 6164 3230 6180
rect 3237 6164 3243 6166
rect 3251 6164 3266 6180
rect 3332 6174 3351 6177
rect 2973 6152 3071 6154
rect 3098 6152 3266 6164
rect 3281 6154 3297 6168
rect 3332 6155 3354 6174
rect 3364 6168 3380 6169
rect 3363 6166 3380 6168
rect 3364 6161 3380 6166
rect 3354 6154 3360 6155
rect 3363 6154 3392 6161
rect 3281 6153 3392 6154
rect 3281 6152 3398 6153
rect 2957 6144 3008 6152
rect 3055 6144 3089 6152
rect 2957 6132 2982 6144
rect 2989 6132 3008 6144
rect 3062 6142 3089 6144
rect 3098 6142 3319 6152
rect 3354 6149 3360 6152
rect 3062 6138 3319 6142
rect 2957 6124 3008 6132
rect 3055 6124 3319 6138
rect 3363 6144 3398 6152
rect 2909 6076 2928 6110
rect 2973 6116 3002 6124
rect 2973 6110 2990 6116
rect 2973 6108 3007 6110
rect 3055 6108 3071 6124
rect 3072 6114 3280 6124
rect 3281 6114 3297 6124
rect 3345 6120 3360 6135
rect 3363 6132 3364 6144
rect 3371 6132 3398 6144
rect 3363 6124 3398 6132
rect 3363 6123 3392 6124
rect 3083 6110 3297 6114
rect 3098 6108 3297 6110
rect 3332 6110 3345 6120
rect 3363 6110 3380 6123
rect 3332 6108 3380 6110
rect 2974 6104 3007 6108
rect 2970 6102 3007 6104
rect 2970 6101 3037 6102
rect 2970 6096 3001 6101
rect 3007 6096 3037 6101
rect 2970 6092 3037 6096
rect 2943 6089 3037 6092
rect 2943 6082 2992 6089
rect 2943 6076 2973 6082
rect 2992 6077 2997 6082
rect 2909 6060 2989 6076
rect 3001 6068 3037 6089
rect 3098 6084 3287 6108
rect 3332 6107 3379 6108
rect 3345 6102 3379 6107
rect 3113 6081 3287 6084
rect 3106 6078 3287 6081
rect 3315 6101 3379 6102
rect 2909 6058 2928 6060
rect 2943 6058 2977 6060
rect 2909 6042 2989 6058
rect 2909 6036 2928 6042
rect 2625 6010 2728 6020
rect 2579 6008 2728 6010
rect 2749 6008 2784 6020
rect 2418 6006 2580 6008
rect 2430 5986 2449 6006
rect 2464 6004 2494 6006
rect 2313 5978 2354 5986
rect 2436 5982 2449 5986
rect 2501 5990 2580 6006
rect 2612 6006 2784 6008
rect 2612 5990 2691 6006
rect 2698 6004 2728 6006
rect 2276 5968 2305 5978
rect 2319 5968 2348 5978
rect 2363 5968 2393 5982
rect 2436 5968 2479 5982
rect 2501 5978 2691 5990
rect 2756 5986 2762 6006
rect 2486 5968 2516 5978
rect 2517 5968 2675 5978
rect 2679 5968 2709 5978
rect 2713 5968 2743 5982
rect 2771 5968 2784 6006
rect 2856 6020 2885 6036
rect 2899 6020 2928 6036
rect 2943 6026 2973 6042
rect 3001 6020 3007 6068
rect 3010 6062 3029 6068
rect 3044 6062 3074 6070
rect 3010 6054 3074 6062
rect 3010 6038 3090 6054
rect 3106 6047 3168 6078
rect 3184 6047 3246 6078
rect 3315 6076 3364 6101
rect 3379 6076 3409 6092
rect 3278 6062 3308 6070
rect 3315 6068 3425 6076
rect 3278 6054 3323 6062
rect 3010 6036 3029 6038
rect 3044 6036 3090 6038
rect 3010 6020 3090 6036
rect 3117 6034 3152 6047
rect 3193 6044 3230 6047
rect 3193 6042 3235 6044
rect 3122 6031 3152 6034
rect 3131 6027 3138 6031
rect 3138 6026 3139 6027
rect 3097 6020 3107 6026
rect 2856 6012 2891 6020
rect 2856 5986 2857 6012
rect 2864 5986 2891 6012
rect 2799 5968 2829 5982
rect 2856 5978 2891 5986
rect 2893 6012 2934 6020
rect 2893 5986 2908 6012
rect 2915 5986 2934 6012
rect 2998 6008 3029 6020
rect 3044 6008 3147 6020
rect 3159 6010 3185 6036
rect 3200 6031 3230 6042
rect 3262 6038 3324 6054
rect 3262 6036 3308 6038
rect 3262 6020 3324 6036
rect 3336 6020 3342 6068
rect 3345 6060 3425 6068
rect 3345 6058 3364 6060
rect 3379 6058 3413 6060
rect 3345 6042 3425 6058
rect 3345 6020 3364 6042
rect 3379 6026 3409 6042
rect 3437 6036 3443 6110
rect 3446 6036 3465 6180
rect 3480 6036 3486 6180
rect 3495 6110 3508 6180
rect 3560 6176 3582 6180
rect 3553 6154 3582 6168
rect 3635 6154 3651 6168
rect 3689 6164 3695 6166
rect 3702 6164 3810 6180
rect 3817 6164 3823 6166
rect 3831 6164 3846 6180
rect 3912 6174 3931 6177
rect 3553 6152 3651 6154
rect 3678 6152 3846 6164
rect 3861 6154 3877 6168
rect 3912 6155 3934 6174
rect 3944 6168 3960 6169
rect 3943 6166 3960 6168
rect 3944 6161 3960 6166
rect 3934 6154 3940 6155
rect 3943 6154 3972 6161
rect 3861 6153 3972 6154
rect 3861 6152 3978 6153
rect 3537 6144 3588 6152
rect 3635 6144 3669 6152
rect 3537 6132 3562 6144
rect 3569 6132 3588 6144
rect 3642 6142 3669 6144
rect 3678 6142 3899 6152
rect 3934 6149 3940 6152
rect 3642 6138 3899 6142
rect 3537 6124 3588 6132
rect 3635 6124 3899 6138
rect 3943 6144 3978 6152
rect 3489 6076 3508 6110
rect 3553 6116 3582 6124
rect 3553 6110 3570 6116
rect 3553 6108 3587 6110
rect 3635 6108 3651 6124
rect 3652 6114 3860 6124
rect 3861 6114 3877 6124
rect 3925 6120 3940 6135
rect 3943 6132 3944 6144
rect 3951 6132 3978 6144
rect 3943 6124 3978 6132
rect 3943 6123 3972 6124
rect 3663 6110 3877 6114
rect 3678 6108 3877 6110
rect 3912 6110 3925 6120
rect 3943 6110 3960 6123
rect 3912 6108 3960 6110
rect 3554 6104 3587 6108
rect 3550 6102 3587 6104
rect 3550 6101 3617 6102
rect 3550 6096 3581 6101
rect 3587 6096 3617 6101
rect 3550 6092 3617 6096
rect 3523 6089 3617 6092
rect 3523 6082 3572 6089
rect 3523 6076 3553 6082
rect 3572 6077 3577 6082
rect 3489 6060 3569 6076
rect 3581 6068 3617 6089
rect 3678 6084 3867 6108
rect 3912 6107 3959 6108
rect 3925 6102 3959 6107
rect 3693 6081 3867 6084
rect 3686 6078 3867 6081
rect 3895 6101 3959 6102
rect 3489 6058 3508 6060
rect 3523 6058 3557 6060
rect 3489 6042 3569 6058
rect 3489 6036 3508 6042
rect 3205 6010 3308 6020
rect 3159 6008 3308 6010
rect 3329 6008 3364 6020
rect 2998 6006 3160 6008
rect 3010 5986 3029 6006
rect 3044 6004 3074 6006
rect 2893 5978 2934 5986
rect 3016 5982 3029 5986
rect 3081 5990 3160 6006
rect 3192 6006 3364 6008
rect 3192 5990 3271 6006
rect 3278 6004 3308 6006
rect 2856 5968 2885 5978
rect 2899 5968 2928 5978
rect 2943 5968 2973 5982
rect 3016 5968 3059 5982
rect 3081 5978 3271 5990
rect 3336 5986 3342 6006
rect 3066 5968 3096 5978
rect 3097 5968 3255 5978
rect 3259 5968 3289 5978
rect 3293 5968 3323 5982
rect 3351 5968 3364 6006
rect 3436 6020 3465 6036
rect 3479 6020 3508 6036
rect 3523 6026 3553 6042
rect 3581 6020 3587 6068
rect 3590 6062 3609 6068
rect 3624 6062 3654 6070
rect 3590 6054 3654 6062
rect 3590 6038 3670 6054
rect 3686 6047 3748 6078
rect 3764 6047 3826 6078
rect 3895 6076 3944 6101
rect 3959 6076 3989 6092
rect 3858 6062 3888 6070
rect 3895 6068 4005 6076
rect 3858 6054 3903 6062
rect 3590 6036 3609 6038
rect 3624 6036 3670 6038
rect 3590 6020 3670 6036
rect 3697 6034 3732 6047
rect 3773 6044 3810 6047
rect 3773 6042 3815 6044
rect 3702 6031 3732 6034
rect 3711 6027 3718 6031
rect 3718 6026 3719 6027
rect 3677 6020 3687 6026
rect 3436 6012 3471 6020
rect 3436 5986 3437 6012
rect 3444 5986 3471 6012
rect 3379 5968 3409 5982
rect 3436 5978 3471 5986
rect 3473 6012 3514 6020
rect 3473 5986 3488 6012
rect 3495 5986 3514 6012
rect 3578 6008 3609 6020
rect 3624 6008 3727 6020
rect 3739 6010 3765 6036
rect 3780 6031 3810 6042
rect 3842 6038 3904 6054
rect 3842 6036 3888 6038
rect 3842 6020 3904 6036
rect 3916 6020 3922 6068
rect 3925 6060 4005 6068
rect 3925 6058 3944 6060
rect 3959 6058 3993 6060
rect 3925 6042 4005 6058
rect 3925 6020 3944 6042
rect 3959 6026 3989 6042
rect 4017 6036 4023 6110
rect 4026 6036 4045 6180
rect 4060 6036 4066 6180
rect 4075 6110 4088 6180
rect 4140 6176 4162 6180
rect 4133 6154 4162 6168
rect 4215 6154 4231 6168
rect 4269 6164 4275 6166
rect 4282 6164 4390 6180
rect 4397 6164 4403 6166
rect 4411 6164 4426 6180
rect 4492 6174 4511 6177
rect 4133 6152 4231 6154
rect 4258 6152 4426 6164
rect 4441 6154 4457 6168
rect 4492 6155 4514 6174
rect 4524 6168 4540 6169
rect 4523 6166 4540 6168
rect 4524 6161 4540 6166
rect 4514 6154 4520 6155
rect 4523 6154 4552 6161
rect 4441 6153 4552 6154
rect 4441 6152 4558 6153
rect 4117 6144 4168 6152
rect 4215 6144 4249 6152
rect 4117 6132 4142 6144
rect 4149 6132 4168 6144
rect 4222 6142 4249 6144
rect 4258 6142 4479 6152
rect 4514 6149 4520 6152
rect 4222 6138 4479 6142
rect 4117 6124 4168 6132
rect 4215 6124 4479 6138
rect 4523 6144 4558 6152
rect 4069 6076 4088 6110
rect 4133 6116 4162 6124
rect 4133 6110 4150 6116
rect 4133 6108 4167 6110
rect 4215 6108 4231 6124
rect 4232 6114 4440 6124
rect 4441 6114 4457 6124
rect 4505 6120 4520 6135
rect 4523 6132 4524 6144
rect 4531 6132 4558 6144
rect 4523 6124 4558 6132
rect 4523 6123 4552 6124
rect 4243 6110 4457 6114
rect 4258 6108 4457 6110
rect 4492 6110 4505 6120
rect 4523 6110 4540 6123
rect 4492 6108 4540 6110
rect 4134 6104 4167 6108
rect 4130 6102 4167 6104
rect 4130 6101 4197 6102
rect 4130 6096 4161 6101
rect 4167 6096 4197 6101
rect 4130 6092 4197 6096
rect 4103 6089 4197 6092
rect 4103 6082 4152 6089
rect 4103 6076 4133 6082
rect 4152 6077 4157 6082
rect 4069 6060 4149 6076
rect 4161 6068 4197 6089
rect 4258 6084 4447 6108
rect 4492 6107 4539 6108
rect 4505 6102 4539 6107
rect 4273 6081 4447 6084
rect 4266 6078 4447 6081
rect 4475 6101 4539 6102
rect 4069 6058 4088 6060
rect 4103 6058 4137 6060
rect 4069 6042 4149 6058
rect 4069 6036 4088 6042
rect 3785 6010 3888 6020
rect 3739 6008 3888 6010
rect 3909 6008 3944 6020
rect 3578 6006 3740 6008
rect 3590 5986 3609 6006
rect 3624 6004 3654 6006
rect 3473 5978 3514 5986
rect 3596 5982 3609 5986
rect 3661 5990 3740 6006
rect 3772 6006 3944 6008
rect 3772 5990 3851 6006
rect 3858 6004 3888 6006
rect 3436 5968 3465 5978
rect 3479 5968 3508 5978
rect 3523 5968 3553 5982
rect 3596 5968 3639 5982
rect 3661 5978 3851 5990
rect 3916 5986 3922 6006
rect 3646 5968 3676 5978
rect 3677 5968 3835 5978
rect 3839 5968 3869 5978
rect 3873 5968 3903 5982
rect 3931 5968 3944 6006
rect 4016 6020 4045 6036
rect 4059 6020 4088 6036
rect 4103 6026 4133 6042
rect 4161 6020 4167 6068
rect 4170 6062 4189 6068
rect 4204 6062 4234 6070
rect 4170 6054 4234 6062
rect 4170 6038 4250 6054
rect 4266 6047 4328 6078
rect 4344 6047 4406 6078
rect 4475 6076 4524 6101
rect 4539 6076 4569 6092
rect 4438 6062 4468 6070
rect 4475 6068 4585 6076
rect 4438 6054 4483 6062
rect 4170 6036 4189 6038
rect 4204 6036 4250 6038
rect 4170 6020 4250 6036
rect 4277 6034 4312 6047
rect 4353 6044 4390 6047
rect 4353 6042 4395 6044
rect 4282 6031 4312 6034
rect 4291 6027 4298 6031
rect 4298 6026 4299 6027
rect 4257 6020 4267 6026
rect 4016 6012 4051 6020
rect 4016 5986 4017 6012
rect 4024 5986 4051 6012
rect 3959 5968 3989 5982
rect 4016 5978 4051 5986
rect 4053 6012 4094 6020
rect 4053 5986 4068 6012
rect 4075 5986 4094 6012
rect 4158 6008 4189 6020
rect 4204 6008 4307 6020
rect 4319 6010 4345 6036
rect 4360 6031 4390 6042
rect 4422 6038 4484 6054
rect 4422 6036 4468 6038
rect 4422 6020 4484 6036
rect 4496 6020 4502 6068
rect 4505 6060 4585 6068
rect 4505 6058 4524 6060
rect 4539 6058 4573 6060
rect 4505 6042 4585 6058
rect 4505 6020 4524 6042
rect 4539 6026 4569 6042
rect 4597 6036 4603 6110
rect 4606 6036 4625 6180
rect 4640 6036 4646 6180
rect 4655 6110 4668 6180
rect 4720 6176 4742 6180
rect 4713 6154 4742 6168
rect 4795 6154 4811 6168
rect 4849 6164 4855 6166
rect 4862 6164 4970 6180
rect 4977 6164 4983 6166
rect 4991 6164 5006 6180
rect 5072 6174 5091 6177
rect 4713 6152 4811 6154
rect 4838 6152 5006 6164
rect 5021 6154 5037 6168
rect 5072 6155 5094 6174
rect 5104 6168 5120 6169
rect 5103 6166 5120 6168
rect 5104 6161 5120 6166
rect 5094 6154 5100 6155
rect 5103 6154 5132 6161
rect 5021 6153 5132 6154
rect 5021 6152 5138 6153
rect 4697 6144 4748 6152
rect 4795 6144 4829 6152
rect 4697 6132 4722 6144
rect 4729 6132 4748 6144
rect 4802 6142 4829 6144
rect 4838 6142 5059 6152
rect 5094 6149 5100 6152
rect 4802 6138 5059 6142
rect 4697 6124 4748 6132
rect 4795 6124 5059 6138
rect 5103 6144 5138 6152
rect 4649 6076 4668 6110
rect 4713 6116 4742 6124
rect 4713 6110 4730 6116
rect 4713 6108 4747 6110
rect 4795 6108 4811 6124
rect 4812 6114 5020 6124
rect 5021 6114 5037 6124
rect 5085 6120 5100 6135
rect 5103 6132 5104 6144
rect 5111 6132 5138 6144
rect 5103 6124 5138 6132
rect 5103 6123 5132 6124
rect 4823 6110 5037 6114
rect 4838 6108 5037 6110
rect 5072 6110 5085 6120
rect 5103 6110 5120 6123
rect 5072 6108 5120 6110
rect 4714 6104 4747 6108
rect 4710 6102 4747 6104
rect 4710 6101 4777 6102
rect 4710 6096 4741 6101
rect 4747 6096 4777 6101
rect 4710 6092 4777 6096
rect 4683 6089 4777 6092
rect 4683 6082 4732 6089
rect 4683 6076 4713 6082
rect 4732 6077 4737 6082
rect 4649 6060 4729 6076
rect 4741 6068 4777 6089
rect 4838 6084 5027 6108
rect 5072 6107 5119 6108
rect 5085 6102 5119 6107
rect 4853 6081 5027 6084
rect 4846 6078 5027 6081
rect 5055 6101 5119 6102
rect 4649 6058 4668 6060
rect 4683 6058 4717 6060
rect 4649 6042 4729 6058
rect 4649 6036 4668 6042
rect 4365 6010 4468 6020
rect 4319 6008 4468 6010
rect 4489 6008 4524 6020
rect 4158 6006 4320 6008
rect 4170 5986 4189 6006
rect 4204 6004 4234 6006
rect 4053 5978 4094 5986
rect 4176 5982 4189 5986
rect 4241 5990 4320 6006
rect 4352 6006 4524 6008
rect 4352 5990 4431 6006
rect 4438 6004 4468 6006
rect 4016 5968 4045 5978
rect 4059 5968 4088 5978
rect 4103 5968 4133 5982
rect 4176 5968 4219 5982
rect 4241 5978 4431 5990
rect 4496 5986 4502 6006
rect 4226 5968 4256 5978
rect 4257 5968 4415 5978
rect 4419 5968 4449 5978
rect 4453 5968 4483 5982
rect 4511 5968 4524 6006
rect 4596 6020 4625 6036
rect 4639 6020 4668 6036
rect 4683 6026 4713 6042
rect 4741 6020 4747 6068
rect 4750 6062 4769 6068
rect 4784 6062 4814 6070
rect 4750 6054 4814 6062
rect 4750 6038 4830 6054
rect 4846 6047 4908 6078
rect 4924 6047 4986 6078
rect 5055 6076 5104 6101
rect 5119 6076 5149 6092
rect 5018 6062 5048 6070
rect 5055 6068 5165 6076
rect 5018 6054 5063 6062
rect 4750 6036 4769 6038
rect 4784 6036 4830 6038
rect 4750 6020 4830 6036
rect 4857 6034 4892 6047
rect 4933 6044 4970 6047
rect 4933 6042 4975 6044
rect 4862 6031 4892 6034
rect 4871 6027 4878 6031
rect 4878 6026 4879 6027
rect 4837 6020 4847 6026
rect 4596 6012 4631 6020
rect 4596 5986 4597 6012
rect 4604 5986 4631 6012
rect 4539 5968 4569 5982
rect 4596 5978 4631 5986
rect 4633 6012 4674 6020
rect 4633 5986 4648 6012
rect 4655 5986 4674 6012
rect 4738 6008 4769 6020
rect 4784 6008 4887 6020
rect 4899 6010 4925 6036
rect 4940 6031 4970 6042
rect 5002 6038 5064 6054
rect 5002 6036 5048 6038
rect 5002 6020 5064 6036
rect 5076 6020 5082 6068
rect 5085 6060 5165 6068
rect 5085 6058 5104 6060
rect 5119 6058 5153 6060
rect 5085 6042 5165 6058
rect 5085 6020 5104 6042
rect 5119 6026 5149 6042
rect 5177 6036 5183 6110
rect 5186 6036 5205 6180
rect 5220 6036 5226 6180
rect 5235 6110 5248 6180
rect 5300 6176 5322 6180
rect 5293 6154 5322 6168
rect 5375 6154 5391 6168
rect 5429 6164 5435 6166
rect 5442 6164 5550 6180
rect 5557 6164 5563 6166
rect 5571 6164 5586 6180
rect 5652 6174 5671 6177
rect 5293 6152 5391 6154
rect 5418 6152 5586 6164
rect 5601 6154 5617 6168
rect 5652 6155 5674 6174
rect 5684 6168 5700 6169
rect 5683 6166 5700 6168
rect 5684 6161 5700 6166
rect 5674 6154 5680 6155
rect 5683 6154 5712 6161
rect 5601 6153 5712 6154
rect 5601 6152 5718 6153
rect 5277 6144 5328 6152
rect 5375 6144 5409 6152
rect 5277 6132 5302 6144
rect 5309 6132 5328 6144
rect 5382 6142 5409 6144
rect 5418 6142 5639 6152
rect 5674 6149 5680 6152
rect 5382 6138 5639 6142
rect 5277 6124 5328 6132
rect 5375 6124 5639 6138
rect 5683 6144 5718 6152
rect 5229 6076 5248 6110
rect 5293 6116 5322 6124
rect 5293 6110 5310 6116
rect 5293 6108 5327 6110
rect 5375 6108 5391 6124
rect 5392 6114 5600 6124
rect 5601 6114 5617 6124
rect 5665 6120 5680 6135
rect 5683 6132 5684 6144
rect 5691 6132 5718 6144
rect 5683 6124 5718 6132
rect 5683 6123 5712 6124
rect 5403 6110 5617 6114
rect 5418 6108 5617 6110
rect 5652 6110 5665 6120
rect 5683 6110 5700 6123
rect 5652 6108 5700 6110
rect 5294 6104 5327 6108
rect 5290 6102 5327 6104
rect 5290 6101 5357 6102
rect 5290 6096 5321 6101
rect 5327 6096 5357 6101
rect 5290 6092 5357 6096
rect 5263 6089 5357 6092
rect 5263 6082 5312 6089
rect 5263 6076 5293 6082
rect 5312 6077 5317 6082
rect 5229 6060 5309 6076
rect 5321 6068 5357 6089
rect 5418 6084 5607 6108
rect 5652 6107 5699 6108
rect 5665 6102 5699 6107
rect 5433 6081 5607 6084
rect 5426 6078 5607 6081
rect 5635 6101 5699 6102
rect 5229 6058 5248 6060
rect 5263 6058 5297 6060
rect 5229 6042 5309 6058
rect 5229 6036 5248 6042
rect 4945 6010 5048 6020
rect 4899 6008 5048 6010
rect 5069 6008 5104 6020
rect 4738 6006 4900 6008
rect 4750 5986 4769 6006
rect 4784 6004 4814 6006
rect 4633 5978 4674 5986
rect 4756 5982 4769 5986
rect 4821 5990 4900 6006
rect 4932 6006 5104 6008
rect 4932 5990 5011 6006
rect 5018 6004 5048 6006
rect 4596 5968 4625 5978
rect 4639 5968 4668 5978
rect 4683 5968 4713 5982
rect 4756 5968 4799 5982
rect 4821 5978 5011 5990
rect 5076 5986 5082 6006
rect 4806 5968 4836 5978
rect 4837 5968 4995 5978
rect 4999 5968 5029 5978
rect 5033 5968 5063 5982
rect 5091 5968 5104 6006
rect 5176 6020 5205 6036
rect 5219 6020 5248 6036
rect 5263 6026 5293 6042
rect 5321 6020 5327 6068
rect 5330 6062 5349 6068
rect 5364 6062 5394 6070
rect 5330 6054 5394 6062
rect 5330 6038 5410 6054
rect 5426 6047 5488 6078
rect 5504 6047 5566 6078
rect 5635 6076 5684 6101
rect 5699 6076 5729 6092
rect 5598 6062 5628 6070
rect 5635 6068 5745 6076
rect 5598 6054 5643 6062
rect 5330 6036 5349 6038
rect 5364 6036 5410 6038
rect 5330 6020 5410 6036
rect 5437 6034 5472 6047
rect 5513 6044 5550 6047
rect 5513 6042 5555 6044
rect 5442 6031 5472 6034
rect 5451 6027 5458 6031
rect 5458 6026 5459 6027
rect 5417 6020 5427 6026
rect 5176 6012 5211 6020
rect 5176 5986 5177 6012
rect 5184 5986 5211 6012
rect 5119 5968 5149 5982
rect 5176 5978 5211 5986
rect 5213 6012 5254 6020
rect 5213 5986 5228 6012
rect 5235 5986 5254 6012
rect 5318 6008 5349 6020
rect 5364 6008 5467 6020
rect 5479 6010 5505 6036
rect 5520 6031 5550 6042
rect 5582 6038 5644 6054
rect 5582 6036 5628 6038
rect 5582 6020 5644 6036
rect 5656 6020 5662 6068
rect 5665 6060 5745 6068
rect 5665 6058 5684 6060
rect 5699 6058 5733 6060
rect 5665 6042 5745 6058
rect 5665 6020 5684 6042
rect 5699 6026 5729 6042
rect 5757 6036 5763 6110
rect 5766 6036 5785 6180
rect 5800 6036 5806 6180
rect 5815 6110 5828 6180
rect 5880 6176 5902 6180
rect 5873 6154 5902 6168
rect 5955 6154 5971 6168
rect 6009 6164 6015 6166
rect 6022 6164 6130 6180
rect 6137 6164 6143 6166
rect 6151 6164 6166 6180
rect 6232 6174 6251 6177
rect 5873 6152 5971 6154
rect 5998 6152 6166 6164
rect 6181 6154 6197 6168
rect 6232 6155 6254 6174
rect 6264 6168 6280 6169
rect 6263 6166 6280 6168
rect 6264 6161 6280 6166
rect 6254 6154 6260 6155
rect 6263 6154 6292 6161
rect 6181 6153 6292 6154
rect 6181 6152 6298 6153
rect 5857 6144 5908 6152
rect 5955 6144 5989 6152
rect 5857 6132 5882 6144
rect 5889 6132 5908 6144
rect 5962 6142 5989 6144
rect 5998 6142 6219 6152
rect 6254 6149 6260 6152
rect 5962 6138 6219 6142
rect 5857 6124 5908 6132
rect 5955 6124 6219 6138
rect 6263 6144 6298 6152
rect 5809 6076 5828 6110
rect 5873 6116 5902 6124
rect 5873 6110 5890 6116
rect 5873 6108 5907 6110
rect 5955 6108 5971 6124
rect 5972 6114 6180 6124
rect 6181 6114 6197 6124
rect 6245 6120 6260 6135
rect 6263 6132 6264 6144
rect 6271 6132 6298 6144
rect 6263 6124 6298 6132
rect 6263 6123 6292 6124
rect 5983 6110 6197 6114
rect 5998 6108 6197 6110
rect 6232 6110 6245 6120
rect 6263 6110 6280 6123
rect 6232 6108 6280 6110
rect 5874 6104 5907 6108
rect 5870 6102 5907 6104
rect 5870 6101 5937 6102
rect 5870 6096 5901 6101
rect 5907 6096 5937 6101
rect 5870 6092 5937 6096
rect 5843 6089 5937 6092
rect 5843 6082 5892 6089
rect 5843 6076 5873 6082
rect 5892 6077 5897 6082
rect 5809 6060 5889 6076
rect 5901 6068 5937 6089
rect 5998 6084 6187 6108
rect 6232 6107 6279 6108
rect 6245 6102 6279 6107
rect 6013 6081 6187 6084
rect 6006 6078 6187 6081
rect 6215 6101 6279 6102
rect 5809 6058 5828 6060
rect 5843 6058 5877 6060
rect 5809 6042 5889 6058
rect 5809 6036 5828 6042
rect 5525 6010 5628 6020
rect 5479 6008 5628 6010
rect 5649 6008 5684 6020
rect 5318 6006 5480 6008
rect 5330 5986 5349 6006
rect 5364 6004 5394 6006
rect 5213 5978 5254 5986
rect 5336 5982 5349 5986
rect 5401 5990 5480 6006
rect 5512 6006 5684 6008
rect 5512 5990 5591 6006
rect 5598 6004 5628 6006
rect 5176 5968 5205 5978
rect 5219 5968 5248 5978
rect 5263 5968 5293 5982
rect 5336 5968 5379 5982
rect 5401 5978 5591 5990
rect 5656 5986 5662 6006
rect 5386 5968 5416 5978
rect 5417 5968 5575 5978
rect 5579 5968 5609 5978
rect 5613 5968 5643 5982
rect 5671 5968 5684 6006
rect 5756 6020 5785 6036
rect 5799 6020 5828 6036
rect 5843 6026 5873 6042
rect 5901 6020 5907 6068
rect 5910 6062 5929 6068
rect 5944 6062 5974 6070
rect 5910 6054 5974 6062
rect 5910 6038 5990 6054
rect 6006 6047 6068 6078
rect 6084 6047 6146 6078
rect 6215 6076 6264 6101
rect 6279 6076 6309 6092
rect 6178 6062 6208 6070
rect 6215 6068 6325 6076
rect 6178 6054 6223 6062
rect 5910 6036 5929 6038
rect 5944 6036 5990 6038
rect 5910 6020 5990 6036
rect 6017 6034 6052 6047
rect 6093 6044 6130 6047
rect 6093 6042 6135 6044
rect 6022 6031 6052 6034
rect 6031 6027 6038 6031
rect 6038 6026 6039 6027
rect 5997 6020 6007 6026
rect 5756 6012 5791 6020
rect 5756 5986 5757 6012
rect 5764 5986 5791 6012
rect 5699 5968 5729 5982
rect 5756 5978 5791 5986
rect 5793 6012 5834 6020
rect 5793 5986 5808 6012
rect 5815 5986 5834 6012
rect 5898 6008 5929 6020
rect 5944 6008 6047 6020
rect 6059 6010 6085 6036
rect 6100 6031 6130 6042
rect 6162 6038 6224 6054
rect 6162 6036 6208 6038
rect 6162 6020 6224 6036
rect 6236 6020 6242 6068
rect 6245 6060 6325 6068
rect 6245 6058 6264 6060
rect 6279 6058 6313 6060
rect 6245 6042 6325 6058
rect 6245 6020 6264 6042
rect 6279 6026 6309 6042
rect 6337 6036 6343 6110
rect 6346 6036 6365 6180
rect 6380 6036 6386 6180
rect 6395 6110 6408 6180
rect 6460 6176 6482 6180
rect 6453 6154 6482 6168
rect 6535 6154 6551 6168
rect 6589 6164 6595 6166
rect 6602 6164 6710 6180
rect 6717 6164 6723 6166
rect 6731 6164 6746 6180
rect 6812 6174 6831 6177
rect 6453 6152 6551 6154
rect 6578 6152 6746 6164
rect 6761 6154 6777 6168
rect 6812 6155 6834 6174
rect 6844 6168 6860 6169
rect 6843 6166 6860 6168
rect 6844 6161 6860 6166
rect 6834 6154 6840 6155
rect 6843 6154 6872 6161
rect 6761 6153 6872 6154
rect 6761 6152 6878 6153
rect 6437 6144 6488 6152
rect 6535 6144 6569 6152
rect 6437 6132 6462 6144
rect 6469 6132 6488 6144
rect 6542 6142 6569 6144
rect 6578 6142 6799 6152
rect 6834 6149 6840 6152
rect 6542 6138 6799 6142
rect 6437 6124 6488 6132
rect 6535 6124 6799 6138
rect 6843 6144 6878 6152
rect 6389 6076 6408 6110
rect 6453 6116 6482 6124
rect 6453 6110 6470 6116
rect 6453 6108 6487 6110
rect 6535 6108 6551 6124
rect 6552 6114 6760 6124
rect 6761 6114 6777 6124
rect 6825 6120 6840 6135
rect 6843 6132 6844 6144
rect 6851 6132 6878 6144
rect 6843 6124 6878 6132
rect 6843 6123 6872 6124
rect 6563 6110 6777 6114
rect 6578 6108 6777 6110
rect 6812 6110 6825 6120
rect 6843 6110 6860 6123
rect 6812 6108 6860 6110
rect 6454 6104 6487 6108
rect 6450 6102 6487 6104
rect 6450 6101 6517 6102
rect 6450 6096 6481 6101
rect 6487 6096 6517 6101
rect 6450 6092 6517 6096
rect 6423 6089 6517 6092
rect 6423 6082 6472 6089
rect 6423 6076 6453 6082
rect 6472 6077 6477 6082
rect 6389 6060 6469 6076
rect 6481 6068 6517 6089
rect 6578 6084 6767 6108
rect 6812 6107 6859 6108
rect 6825 6102 6859 6107
rect 6593 6081 6767 6084
rect 6586 6078 6767 6081
rect 6795 6101 6859 6102
rect 6389 6058 6408 6060
rect 6423 6058 6457 6060
rect 6389 6042 6469 6058
rect 6389 6036 6408 6042
rect 6105 6010 6208 6020
rect 6059 6008 6208 6010
rect 6229 6008 6264 6020
rect 5898 6006 6060 6008
rect 5910 5986 5929 6006
rect 5944 6004 5974 6006
rect 5793 5978 5834 5986
rect 5916 5982 5929 5986
rect 5981 5990 6060 6006
rect 6092 6006 6264 6008
rect 6092 5990 6171 6006
rect 6178 6004 6208 6006
rect 5756 5968 5785 5978
rect 5799 5968 5828 5978
rect 5843 5968 5873 5982
rect 5916 5968 5959 5982
rect 5981 5978 6171 5990
rect 6236 5986 6242 6006
rect 5966 5968 5996 5978
rect 5997 5968 6155 5978
rect 6159 5968 6189 5978
rect 6193 5968 6223 5982
rect 6251 5968 6264 6006
rect 6336 6020 6365 6036
rect 6379 6020 6408 6036
rect 6423 6026 6453 6042
rect 6481 6020 6487 6068
rect 6490 6062 6509 6068
rect 6524 6062 6554 6070
rect 6490 6054 6554 6062
rect 6490 6038 6570 6054
rect 6586 6047 6648 6078
rect 6664 6047 6726 6078
rect 6795 6076 6844 6101
rect 6859 6076 6889 6092
rect 6758 6062 6788 6070
rect 6795 6068 6905 6076
rect 6758 6054 6803 6062
rect 6490 6036 6509 6038
rect 6524 6036 6570 6038
rect 6490 6020 6570 6036
rect 6597 6034 6632 6047
rect 6673 6044 6710 6047
rect 6673 6042 6715 6044
rect 6602 6031 6632 6034
rect 6611 6027 6618 6031
rect 6618 6026 6619 6027
rect 6577 6020 6587 6026
rect 6336 6012 6371 6020
rect 6336 5986 6337 6012
rect 6344 5986 6371 6012
rect 6279 5968 6309 5982
rect 6336 5978 6371 5986
rect 6373 6012 6414 6020
rect 6373 5986 6388 6012
rect 6395 5986 6414 6012
rect 6478 6008 6509 6020
rect 6524 6008 6627 6020
rect 6639 6010 6665 6036
rect 6680 6031 6710 6042
rect 6742 6038 6804 6054
rect 6742 6036 6788 6038
rect 6742 6020 6804 6036
rect 6816 6020 6822 6068
rect 6825 6060 6905 6068
rect 6825 6058 6844 6060
rect 6859 6058 6893 6060
rect 6825 6042 6905 6058
rect 6825 6020 6844 6042
rect 6859 6026 6889 6042
rect 6917 6036 6923 6110
rect 6926 6036 6945 6180
rect 6960 6036 6966 6180
rect 6975 6110 6988 6180
rect 7040 6176 7062 6180
rect 7033 6154 7062 6168
rect 7115 6154 7131 6168
rect 7169 6164 7175 6166
rect 7182 6164 7290 6180
rect 7297 6164 7303 6166
rect 7311 6164 7326 6180
rect 7392 6174 7411 6177
rect 7033 6152 7131 6154
rect 7158 6152 7326 6164
rect 7341 6154 7357 6168
rect 7392 6155 7414 6174
rect 7424 6168 7440 6169
rect 7423 6166 7440 6168
rect 7424 6161 7440 6166
rect 7414 6154 7420 6155
rect 7423 6154 7452 6161
rect 7341 6153 7452 6154
rect 7341 6152 7458 6153
rect 7017 6144 7068 6152
rect 7115 6144 7149 6152
rect 7017 6132 7042 6144
rect 7049 6132 7068 6144
rect 7122 6142 7149 6144
rect 7158 6142 7379 6152
rect 7414 6149 7420 6152
rect 7122 6138 7379 6142
rect 7017 6124 7068 6132
rect 7115 6124 7379 6138
rect 7423 6144 7458 6152
rect 6969 6076 6988 6110
rect 7033 6116 7062 6124
rect 7033 6110 7050 6116
rect 7033 6108 7067 6110
rect 7115 6108 7131 6124
rect 7132 6114 7340 6124
rect 7341 6114 7357 6124
rect 7405 6120 7420 6135
rect 7423 6132 7424 6144
rect 7431 6132 7458 6144
rect 7423 6124 7458 6132
rect 7423 6123 7452 6124
rect 7143 6110 7357 6114
rect 7158 6108 7357 6110
rect 7392 6110 7405 6120
rect 7423 6110 7440 6123
rect 7392 6108 7440 6110
rect 7034 6104 7067 6108
rect 7030 6102 7067 6104
rect 7030 6101 7097 6102
rect 7030 6096 7061 6101
rect 7067 6096 7097 6101
rect 7030 6092 7097 6096
rect 7003 6089 7097 6092
rect 7003 6082 7052 6089
rect 7003 6076 7033 6082
rect 7052 6077 7057 6082
rect 6969 6060 7049 6076
rect 7061 6068 7097 6089
rect 7158 6084 7347 6108
rect 7392 6107 7439 6108
rect 7405 6102 7439 6107
rect 7173 6081 7347 6084
rect 7166 6078 7347 6081
rect 7375 6101 7439 6102
rect 6969 6058 6988 6060
rect 7003 6058 7037 6060
rect 6969 6042 7049 6058
rect 6969 6036 6988 6042
rect 6685 6010 6788 6020
rect 6639 6008 6788 6010
rect 6809 6008 6844 6020
rect 6478 6006 6640 6008
rect 6490 5986 6509 6006
rect 6524 6004 6554 6006
rect 6373 5978 6414 5986
rect 6496 5982 6509 5986
rect 6561 5990 6640 6006
rect 6672 6006 6844 6008
rect 6672 5990 6751 6006
rect 6758 6004 6788 6006
rect 6336 5968 6365 5978
rect 6379 5968 6408 5978
rect 6423 5968 6453 5982
rect 6496 5968 6539 5982
rect 6561 5978 6751 5990
rect 6816 5986 6822 6006
rect 6546 5968 6576 5978
rect 6577 5968 6735 5978
rect 6739 5968 6769 5978
rect 6773 5968 6803 5982
rect 6831 5968 6844 6006
rect 6916 6020 6945 6036
rect 6959 6020 6988 6036
rect 7003 6026 7033 6042
rect 7061 6020 7067 6068
rect 7070 6062 7089 6068
rect 7104 6062 7134 6070
rect 7070 6054 7134 6062
rect 7070 6038 7150 6054
rect 7166 6047 7228 6078
rect 7244 6047 7306 6078
rect 7375 6076 7424 6101
rect 7439 6076 7469 6092
rect 7338 6062 7368 6070
rect 7375 6068 7485 6076
rect 7338 6054 7383 6062
rect 7070 6036 7089 6038
rect 7104 6036 7150 6038
rect 7070 6020 7150 6036
rect 7177 6034 7212 6047
rect 7253 6044 7290 6047
rect 7253 6042 7295 6044
rect 7182 6031 7212 6034
rect 7191 6027 7198 6031
rect 7198 6026 7199 6027
rect 7157 6020 7167 6026
rect 6916 6012 6951 6020
rect 6916 5986 6917 6012
rect 6924 5986 6951 6012
rect 6859 5968 6889 5982
rect 6916 5978 6951 5986
rect 6953 6012 6994 6020
rect 6953 5986 6968 6012
rect 6975 5986 6994 6012
rect 7058 6008 7089 6020
rect 7104 6008 7207 6020
rect 7219 6010 7245 6036
rect 7260 6031 7290 6042
rect 7322 6038 7384 6054
rect 7322 6036 7368 6038
rect 7322 6020 7384 6036
rect 7396 6020 7402 6068
rect 7405 6060 7485 6068
rect 7405 6058 7424 6060
rect 7439 6058 7473 6060
rect 7405 6042 7485 6058
rect 7405 6020 7424 6042
rect 7439 6026 7469 6042
rect 7497 6036 7503 6110
rect 7506 6036 7525 6180
rect 7540 6036 7546 6180
rect 7555 6110 7568 6180
rect 7613 6158 7614 6168
rect 7629 6158 7642 6168
rect 7613 6154 7642 6158
rect 7647 6154 7677 6180
rect 7695 6166 7711 6168
rect 7783 6166 7836 6180
rect 7784 6164 7848 6166
rect 7891 6164 7906 6180
rect 7955 6177 7985 6180
rect 7955 6174 7991 6177
rect 7921 6166 7937 6168
rect 7695 6154 7710 6158
rect 7613 6152 7710 6154
rect 7738 6152 7906 6164
rect 7922 6154 7937 6158
rect 7955 6155 7994 6174
rect 8013 6168 8020 6169
rect 8019 6161 8020 6168
rect 8003 6158 8004 6161
rect 8019 6158 8032 6161
rect 7955 6154 7985 6155
rect 7994 6154 8000 6155
rect 8003 6154 8032 6158
rect 7922 6153 8032 6154
rect 7922 6152 8038 6153
rect 7597 6144 7648 6152
rect 7597 6132 7622 6144
rect 7629 6132 7648 6144
rect 7679 6144 7729 6152
rect 7679 6136 7695 6144
rect 7702 6142 7729 6144
rect 7738 6142 7959 6152
rect 7702 6132 7959 6142
rect 7988 6144 8038 6152
rect 7988 6135 8004 6144
rect 7597 6124 7648 6132
rect 7695 6124 7959 6132
rect 7985 6132 8004 6135
rect 8011 6132 8038 6144
rect 7985 6124 8038 6132
rect 7549 6076 7568 6110
rect 7613 6116 7614 6124
rect 7629 6116 7642 6124
rect 7613 6108 7629 6116
rect 7610 6101 7629 6104
rect 7610 6092 7632 6101
rect 7583 6082 7632 6092
rect 7583 6076 7613 6082
rect 7632 6077 7637 6082
rect 7549 6060 7629 6076
rect 7647 6068 7677 6124
rect 7712 6114 7920 6124
rect 7955 6120 8000 6124
rect 8003 6123 8004 6124
rect 8019 6123 8032 6124
rect 7738 6084 7927 6114
rect 7753 6081 7927 6084
rect 7746 6078 7927 6081
rect 7549 6058 7568 6060
rect 7583 6058 7617 6060
rect 7549 6042 7629 6058
rect 7656 6054 7669 6068
rect 7684 6054 7700 6070
rect 7746 6065 7757 6078
rect 7549 6036 7568 6042
rect 7265 6010 7368 6020
rect 7219 6008 7368 6010
rect 7389 6008 7424 6020
rect 7058 6006 7220 6008
rect 7070 5986 7089 6006
rect 7104 6004 7134 6006
rect 6953 5978 6994 5986
rect 7076 5982 7089 5986
rect 7141 5990 7220 6006
rect 7252 6006 7424 6008
rect 7252 5990 7331 6006
rect 7338 6004 7368 6006
rect 6916 5968 6945 5978
rect 6959 5968 6988 5978
rect 7003 5968 7033 5982
rect 7076 5968 7119 5982
rect 7141 5978 7331 5990
rect 7396 5986 7402 6006
rect 7126 5968 7156 5978
rect 7157 5968 7315 5978
rect 7319 5968 7349 5978
rect 7353 5968 7383 5982
rect 7411 5968 7424 6006
rect 7496 6020 7525 6036
rect 7539 6020 7568 6036
rect 7583 6020 7613 6042
rect 7656 6038 7718 6054
rect 7746 6047 7757 6063
rect 7762 6058 7772 6078
rect 7782 6058 7796 6078
rect 7799 6065 7808 6078
rect 7824 6065 7833 6078
rect 7762 6047 7796 6058
rect 7799 6047 7808 6063
rect 7824 6047 7833 6063
rect 7840 6058 7850 6078
rect 7860 6058 7874 6078
rect 7875 6065 7886 6078
rect 7840 6047 7874 6058
rect 7875 6047 7886 6063
rect 7932 6054 7948 6070
rect 7955 6068 7985 6120
rect 8019 6116 8020 6123
rect 8004 6108 8020 6116
rect 7991 6076 8004 6095
rect 8019 6076 8049 6092
rect 7991 6060 8065 6076
rect 7991 6058 8004 6060
rect 8019 6058 8053 6060
rect 7656 6036 7669 6038
rect 7684 6036 7718 6038
rect 7656 6020 7718 6036
rect 7762 6031 7778 6034
rect 7840 6031 7870 6042
rect 7918 6038 7964 6054
rect 7991 6042 8065 6058
rect 7918 6036 7952 6038
rect 7917 6020 7964 6036
rect 7991 6020 8004 6042
rect 8019 6020 8049 6042
rect 8076 6020 8077 6036
rect 8092 6020 8105 6180
rect 8135 6076 8148 6180
rect 8193 6158 8194 6168
rect 8209 6158 8222 6168
rect 8193 6154 8222 6158
rect 8227 6154 8257 6180
rect 8275 6166 8291 6168
rect 8363 6166 8416 6180
rect 8364 6164 8428 6166
rect 8471 6164 8486 6180
rect 8535 6177 8565 6180
rect 8535 6174 8571 6177
rect 8501 6166 8517 6168
rect 8275 6154 8290 6158
rect 8193 6152 8290 6154
rect 8318 6152 8486 6164
rect 8502 6154 8517 6158
rect 8535 6155 8574 6174
rect 8593 6168 8600 6169
rect 8599 6161 8600 6168
rect 8583 6158 8584 6161
rect 8599 6158 8612 6161
rect 8535 6154 8565 6155
rect 8574 6154 8580 6155
rect 8583 6154 8612 6158
rect 8502 6153 8612 6154
rect 8502 6152 8618 6153
rect 8177 6144 8228 6152
rect 8177 6132 8202 6144
rect 8209 6132 8228 6144
rect 8259 6144 8309 6152
rect 8259 6136 8275 6144
rect 8282 6142 8309 6144
rect 8318 6142 8539 6152
rect 8282 6132 8539 6142
rect 8568 6144 8618 6152
rect 8568 6135 8584 6144
rect 8177 6124 8228 6132
rect 8275 6124 8539 6132
rect 8565 6132 8584 6135
rect 8591 6132 8618 6144
rect 8565 6124 8618 6132
rect 8193 6116 8194 6124
rect 8209 6116 8222 6124
rect 8193 6108 8209 6116
rect 8190 6101 8209 6104
rect 8190 6092 8212 6101
rect 8163 6082 8212 6092
rect 8163 6076 8193 6082
rect 8212 6077 8217 6082
rect 8135 6060 8209 6076
rect 8227 6068 8257 6124
rect 8292 6114 8500 6124
rect 8535 6120 8580 6124
rect 8583 6123 8584 6124
rect 8599 6123 8612 6124
rect 8318 6084 8507 6114
rect 8333 6081 8507 6084
rect 8326 6078 8507 6081
rect 8135 6058 8148 6060
rect 8163 6058 8197 6060
rect 8135 6042 8209 6058
rect 8236 6054 8249 6068
rect 8264 6054 8280 6070
rect 8326 6065 8337 6078
rect 8119 6020 8120 6036
rect 8135 6020 8148 6042
rect 8163 6020 8193 6042
rect 8236 6038 8298 6054
rect 8326 6047 8337 6063
rect 8342 6058 8352 6078
rect 8362 6058 8376 6078
rect 8379 6065 8388 6078
rect 8404 6065 8413 6078
rect 8342 6047 8376 6058
rect 8379 6047 8388 6063
rect 8404 6047 8413 6063
rect 8420 6058 8430 6078
rect 8440 6058 8454 6078
rect 8455 6065 8466 6078
rect 8420 6047 8454 6058
rect 8455 6047 8466 6063
rect 8512 6054 8528 6070
rect 8535 6068 8565 6120
rect 8599 6116 8600 6123
rect 8584 6108 8600 6116
rect 8571 6076 8584 6095
rect 8599 6076 8629 6092
rect 8571 6060 8645 6076
rect 8571 6058 8584 6060
rect 8599 6058 8633 6060
rect 8236 6036 8249 6038
rect 8264 6036 8298 6038
rect 8236 6020 8298 6036
rect 8342 6031 8358 6034
rect 8420 6031 8450 6042
rect 8498 6038 8544 6054
rect 8571 6042 8645 6058
rect 8498 6036 8532 6038
rect 8497 6020 8544 6036
rect 8571 6020 8584 6042
rect 8599 6020 8629 6042
rect 8656 6020 8657 6036
rect 8672 6020 8685 6180
rect 8715 6076 8728 6180
rect 8773 6158 8774 6168
rect 8789 6158 8802 6168
rect 8773 6154 8802 6158
rect 8807 6154 8837 6180
rect 8855 6166 8871 6168
rect 8943 6166 8996 6180
rect 8944 6164 9008 6166
rect 9051 6164 9066 6180
rect 9115 6177 9145 6180
rect 9115 6174 9151 6177
rect 9081 6166 9097 6168
rect 8855 6154 8870 6158
rect 8773 6152 8870 6154
rect 8898 6152 9066 6164
rect 9082 6154 9097 6158
rect 9115 6155 9154 6174
rect 9173 6168 9180 6169
rect 9179 6161 9180 6168
rect 9163 6158 9164 6161
rect 9179 6158 9192 6161
rect 9115 6154 9145 6155
rect 9154 6154 9160 6155
rect 9163 6154 9192 6158
rect 9082 6153 9192 6154
rect 9082 6152 9198 6153
rect 8757 6144 8808 6152
rect 8757 6132 8782 6144
rect 8789 6132 8808 6144
rect 8839 6144 8889 6152
rect 8839 6136 8855 6144
rect 8862 6142 8889 6144
rect 8898 6142 9119 6152
rect 8862 6132 9119 6142
rect 9148 6144 9198 6152
rect 9148 6135 9164 6144
rect 8757 6124 8808 6132
rect 8855 6124 9119 6132
rect 9145 6132 9164 6135
rect 9171 6132 9198 6144
rect 9145 6124 9198 6132
rect 8773 6116 8774 6124
rect 8789 6116 8802 6124
rect 8773 6108 8789 6116
rect 8770 6101 8789 6104
rect 8770 6092 8792 6101
rect 8743 6082 8792 6092
rect 8743 6076 8773 6082
rect 8792 6077 8797 6082
rect 8715 6060 8789 6076
rect 8807 6068 8837 6124
rect 8872 6114 9080 6124
rect 9115 6120 9160 6124
rect 9163 6123 9164 6124
rect 9179 6123 9192 6124
rect 8898 6084 9087 6114
rect 8913 6081 9087 6084
rect 8906 6078 9087 6081
rect 8715 6058 8728 6060
rect 8743 6058 8777 6060
rect 8715 6042 8789 6058
rect 8816 6054 8829 6068
rect 8844 6054 8860 6070
rect 8906 6065 8917 6078
rect 8699 6020 8700 6036
rect 8715 6020 8728 6042
rect 8743 6020 8773 6042
rect 8816 6038 8878 6054
rect 8906 6047 8917 6063
rect 8922 6058 8932 6078
rect 8942 6058 8956 6078
rect 8959 6065 8968 6078
rect 8984 6065 8993 6078
rect 8922 6047 8956 6058
rect 8959 6047 8968 6063
rect 8984 6047 8993 6063
rect 9000 6058 9010 6078
rect 9020 6058 9034 6078
rect 9035 6065 9046 6078
rect 9000 6047 9034 6058
rect 9035 6047 9046 6063
rect 9092 6054 9108 6070
rect 9115 6068 9145 6120
rect 9179 6116 9180 6123
rect 9164 6108 9180 6116
rect 9151 6076 9164 6095
rect 9179 6076 9209 6092
rect 9151 6060 9225 6076
rect 9151 6058 9164 6060
rect 9179 6058 9213 6060
rect 8816 6036 8829 6038
rect 8844 6036 8878 6038
rect 8816 6020 8878 6036
rect 8922 6031 8938 6034
rect 9000 6031 9030 6042
rect 9078 6038 9124 6054
rect 9151 6042 9225 6058
rect 9078 6036 9112 6038
rect 9077 6020 9124 6036
rect 9151 6020 9164 6042
rect 9179 6020 9209 6042
rect 9236 6020 9237 6036
rect 9252 6020 9265 6180
rect 7496 6012 7531 6020
rect 7496 5986 7497 6012
rect 7504 5986 7531 6012
rect 7439 5968 7469 5982
rect 7496 5978 7531 5986
rect 7533 6012 7574 6020
rect 7533 5986 7548 6012
rect 7555 5986 7574 6012
rect 7638 6008 7700 6020
rect 7712 6008 7787 6020
rect 7845 6008 7920 6020
rect 7932 6008 7963 6020
rect 7969 6008 8004 6020
rect 7638 6006 7800 6008
rect 7533 5978 7574 5986
rect 7656 5982 7669 6006
rect 7684 6004 7699 6006
rect 7496 5968 7525 5978
rect 7539 5968 7568 5978
rect 7583 5968 7613 5982
rect 7656 5968 7699 5982
rect 7723 5979 7730 5986
rect 7733 5982 7800 6006
rect 7832 6006 8004 6008
rect 7802 5984 7830 5988
rect 7832 5984 7912 6006
rect 7933 6004 7948 6006
rect 7802 5982 7912 5984
rect 7733 5978 7912 5982
rect 7706 5968 7736 5978
rect 7738 5968 7891 5978
rect 7899 5968 7929 5978
rect 7933 5968 7963 5982
rect 7991 5968 8004 6006
rect 8076 6012 8111 6020
rect 8076 5986 8077 6012
rect 8084 5986 8111 6012
rect 8019 5968 8049 5982
rect 8076 5978 8111 5986
rect 8113 6012 8154 6020
rect 8113 5986 8128 6012
rect 8135 5986 8154 6012
rect 8218 6008 8280 6020
rect 8292 6008 8367 6020
rect 8425 6008 8500 6020
rect 8512 6008 8543 6020
rect 8549 6008 8584 6020
rect 8218 6006 8380 6008
rect 8113 5978 8154 5986
rect 8236 5982 8249 6006
rect 8264 6004 8279 6006
rect 8076 5968 8077 5978
rect 8092 5968 8105 5978
rect 8119 5968 8120 5978
rect 8135 5968 8148 5978
rect 8163 5968 8193 5982
rect 8236 5968 8279 5982
rect 8303 5979 8310 5986
rect 8313 5982 8380 6006
rect 8412 6006 8584 6008
rect 8382 5984 8410 5988
rect 8412 5984 8492 6006
rect 8513 6004 8528 6006
rect 8382 5982 8492 5984
rect 8313 5978 8492 5982
rect 8286 5968 8316 5978
rect 8318 5968 8471 5978
rect 8479 5968 8509 5978
rect 8513 5968 8543 5982
rect 8571 5968 8584 6006
rect 8656 6012 8691 6020
rect 8656 5986 8657 6012
rect 8664 5986 8691 6012
rect 8599 5968 8629 5982
rect 8656 5978 8691 5986
rect 8693 6012 8734 6020
rect 8693 5986 8708 6012
rect 8715 5986 8734 6012
rect 8798 6008 8860 6020
rect 8872 6008 8947 6020
rect 9005 6008 9080 6020
rect 9092 6008 9123 6020
rect 9129 6008 9164 6020
rect 8798 6006 8960 6008
rect 8693 5978 8734 5986
rect 8816 5982 8829 6006
rect 8844 6004 8859 6006
rect 8656 5968 8657 5978
rect 8672 5968 8685 5978
rect 8699 5968 8700 5978
rect 8715 5968 8728 5978
rect 8743 5968 8773 5982
rect 8816 5968 8859 5982
rect 8883 5979 8890 5986
rect 8893 5982 8960 6006
rect 8992 6006 9164 6008
rect 8962 5984 8990 5988
rect 8992 5984 9072 6006
rect 9093 6004 9108 6006
rect 8962 5982 9072 5984
rect 8893 5978 9072 5982
rect 8866 5968 8896 5978
rect 8898 5968 9051 5978
rect 9059 5968 9089 5978
rect 9093 5968 9123 5982
rect 9151 5968 9164 6006
rect 9236 6012 9271 6020
rect 9236 5986 9237 6012
rect 9244 5986 9271 6012
rect 9179 5968 9209 5982
rect 9236 5978 9271 5986
rect 9236 5968 9237 5978
rect 9252 5968 9265 5978
rect -1 5962 9265 5968
rect 0 5954 9265 5962
rect 15 5924 28 5954
rect 43 5940 73 5954
rect 116 5940 159 5954
rect 166 5940 386 5954
rect 393 5940 423 5954
rect 83 5926 98 5938
rect 117 5926 130 5940
rect 198 5936 351 5940
rect 80 5924 102 5926
rect 180 5924 372 5936
rect 451 5924 464 5954
rect 479 5940 509 5954
rect 546 5924 565 5954
rect 580 5924 586 5954
rect 595 5924 608 5954
rect 623 5940 653 5954
rect 696 5940 739 5954
rect 746 5940 966 5954
rect 973 5940 1003 5954
rect 663 5926 678 5938
rect 697 5926 710 5940
rect 778 5936 931 5940
rect 660 5924 682 5926
rect 760 5924 952 5936
rect 1031 5924 1044 5954
rect 1059 5940 1089 5954
rect 1126 5924 1145 5954
rect 1160 5924 1166 5954
rect 1175 5924 1188 5954
rect 1203 5940 1233 5954
rect 1276 5940 1319 5954
rect 1326 5940 1546 5954
rect 1553 5940 1583 5954
rect 1243 5926 1258 5938
rect 1277 5926 1290 5940
rect 1358 5936 1511 5940
rect 1240 5924 1262 5926
rect 1340 5924 1532 5936
rect 1611 5924 1624 5954
rect 1639 5940 1669 5954
rect 1706 5924 1725 5954
rect 1740 5924 1746 5954
rect 1755 5924 1768 5954
rect 1783 5940 1813 5954
rect 1856 5940 1899 5954
rect 1906 5940 2126 5954
rect 2133 5940 2163 5954
rect 1823 5926 1838 5938
rect 1857 5926 1870 5940
rect 1938 5936 2091 5940
rect 1820 5924 1842 5926
rect 1920 5924 2112 5936
rect 2191 5924 2204 5954
rect 2219 5940 2249 5954
rect 2286 5924 2305 5954
rect 2320 5924 2326 5954
rect 2335 5924 2348 5954
rect 2363 5940 2393 5954
rect 2436 5940 2479 5954
rect 2486 5940 2706 5954
rect 2713 5940 2743 5954
rect 2403 5926 2418 5938
rect 2437 5926 2450 5940
rect 2518 5936 2671 5940
rect 2400 5924 2422 5926
rect 2500 5924 2692 5936
rect 2771 5924 2784 5954
rect 2799 5940 2829 5954
rect 2866 5924 2885 5954
rect 2900 5924 2906 5954
rect 2915 5924 2928 5954
rect 2943 5940 2973 5954
rect 3016 5940 3059 5954
rect 3066 5940 3286 5954
rect 3293 5940 3323 5954
rect 2983 5926 2998 5938
rect 3017 5926 3030 5940
rect 3098 5936 3251 5940
rect 2980 5924 3002 5926
rect 3080 5924 3272 5936
rect 3351 5924 3364 5954
rect 3379 5940 3409 5954
rect 3446 5924 3465 5954
rect 3480 5924 3486 5954
rect 3495 5924 3508 5954
rect 3523 5940 3553 5954
rect 3596 5940 3639 5954
rect 3646 5940 3866 5954
rect 3873 5940 3903 5954
rect 3563 5926 3578 5938
rect 3597 5926 3610 5940
rect 3678 5936 3831 5940
rect 3560 5924 3582 5926
rect 3660 5924 3852 5936
rect 3931 5924 3944 5954
rect 3959 5940 3989 5954
rect 4026 5924 4045 5954
rect 4060 5924 4066 5954
rect 4075 5924 4088 5954
rect 4103 5940 4133 5954
rect 4176 5940 4219 5954
rect 4226 5940 4446 5954
rect 4453 5940 4483 5954
rect 4143 5926 4158 5938
rect 4177 5926 4190 5940
rect 4258 5936 4411 5940
rect 4140 5924 4162 5926
rect 4240 5924 4432 5936
rect 4511 5924 4524 5954
rect 4539 5940 4569 5954
rect 4606 5924 4625 5954
rect 4640 5924 4646 5954
rect 4655 5924 4668 5954
rect 4683 5940 4713 5954
rect 4756 5940 4799 5954
rect 4806 5940 5026 5954
rect 5033 5940 5063 5954
rect 4723 5926 4738 5938
rect 4757 5926 4770 5940
rect 4838 5936 4991 5940
rect 4720 5924 4742 5926
rect 4820 5924 5012 5936
rect 5091 5924 5104 5954
rect 5119 5940 5149 5954
rect 5186 5924 5205 5954
rect 5220 5924 5226 5954
rect 5235 5924 5248 5954
rect 5263 5940 5293 5954
rect 5336 5940 5379 5954
rect 5386 5940 5606 5954
rect 5613 5940 5643 5954
rect 5303 5926 5318 5938
rect 5337 5926 5350 5940
rect 5418 5936 5571 5940
rect 5300 5924 5322 5926
rect 5400 5924 5592 5936
rect 5671 5924 5684 5954
rect 5699 5940 5729 5954
rect 5766 5924 5785 5954
rect 5800 5924 5806 5954
rect 5815 5924 5828 5954
rect 5843 5940 5873 5954
rect 5916 5940 5959 5954
rect 5966 5940 6186 5954
rect 6193 5940 6223 5954
rect 5883 5926 5898 5938
rect 5917 5926 5930 5940
rect 5998 5936 6151 5940
rect 5880 5924 5902 5926
rect 5980 5924 6172 5936
rect 6251 5924 6264 5954
rect 6279 5940 6309 5954
rect 6346 5924 6365 5954
rect 6380 5924 6386 5954
rect 6395 5924 6408 5954
rect 6423 5940 6453 5954
rect 6496 5940 6539 5954
rect 6546 5940 6766 5954
rect 6773 5940 6803 5954
rect 6463 5926 6478 5938
rect 6497 5926 6510 5940
rect 6578 5936 6731 5940
rect 6460 5924 6482 5926
rect 6560 5924 6752 5936
rect 6831 5924 6844 5954
rect 6859 5940 6889 5954
rect 6926 5924 6945 5954
rect 6960 5924 6966 5954
rect 6975 5924 6988 5954
rect 7003 5940 7033 5954
rect 7076 5940 7119 5954
rect 7126 5940 7346 5954
rect 7353 5940 7383 5954
rect 7043 5926 7058 5938
rect 7077 5926 7090 5940
rect 7158 5936 7311 5940
rect 7040 5924 7062 5926
rect 7140 5924 7332 5936
rect 7411 5924 7424 5954
rect 7439 5940 7469 5954
rect 7506 5924 7525 5954
rect 7540 5924 7546 5954
rect 7555 5924 7568 5954
rect 7583 5936 7613 5954
rect 7656 5940 7670 5954
rect 7706 5940 7926 5954
rect 7657 5938 7670 5940
rect 7623 5926 7638 5938
rect 7620 5924 7642 5926
rect 7647 5924 7677 5938
rect 7738 5936 7891 5940
rect 7720 5924 7912 5936
rect 7955 5924 7985 5938
rect 7991 5924 8004 5954
rect 8019 5936 8049 5954
rect 8092 5924 8105 5954
rect 8135 5924 8148 5954
rect 8163 5936 8193 5954
rect 8236 5940 8250 5954
rect 8286 5940 8506 5954
rect 8237 5938 8250 5940
rect 8203 5926 8218 5938
rect 8200 5924 8222 5926
rect 8227 5924 8257 5938
rect 8318 5936 8471 5940
rect 8300 5924 8492 5936
rect 8535 5924 8565 5938
rect 8571 5924 8584 5954
rect 8599 5936 8629 5954
rect 8672 5924 8685 5954
rect 8715 5924 8728 5954
rect 8743 5936 8773 5954
rect 8816 5940 8830 5954
rect 8866 5940 9086 5954
rect 8817 5938 8830 5940
rect 8783 5926 8798 5938
rect 8780 5924 8802 5926
rect 8807 5924 8837 5938
rect 8898 5936 9051 5940
rect 8880 5924 9072 5936
rect 9115 5924 9145 5938
rect 9151 5924 9164 5954
rect 9179 5936 9209 5954
rect 9252 5924 9265 5954
rect 0 5910 9265 5924
rect 15 5840 28 5910
rect 80 5906 102 5910
rect 73 5884 102 5898
rect 155 5884 171 5898
rect 209 5894 215 5896
rect 222 5894 330 5910
rect 337 5894 343 5896
rect 351 5894 366 5910
rect 432 5904 451 5907
rect 73 5882 171 5884
rect 198 5882 366 5894
rect 381 5884 397 5898
rect 432 5885 454 5904
rect 464 5898 480 5899
rect 463 5896 480 5898
rect 464 5891 480 5896
rect 454 5884 460 5885
rect 463 5884 492 5891
rect 381 5883 492 5884
rect 381 5882 498 5883
rect 57 5874 108 5882
rect 155 5874 189 5882
rect 57 5862 82 5874
rect 89 5862 108 5874
rect 162 5872 189 5874
rect 198 5872 419 5882
rect 454 5879 460 5882
rect 162 5868 419 5872
rect 57 5854 108 5862
rect 155 5854 419 5868
rect 463 5874 498 5882
rect 9 5806 28 5840
rect 73 5846 102 5854
rect 73 5840 90 5846
rect 73 5838 107 5840
rect 155 5838 171 5854
rect 172 5844 380 5854
rect 381 5844 397 5854
rect 445 5850 460 5865
rect 463 5862 464 5874
rect 471 5862 498 5874
rect 463 5854 498 5862
rect 463 5853 492 5854
rect 183 5840 397 5844
rect 198 5838 397 5840
rect 432 5840 445 5850
rect 463 5840 480 5853
rect 432 5838 480 5840
rect 74 5834 107 5838
rect 70 5832 107 5834
rect 70 5831 137 5832
rect 70 5826 101 5831
rect 107 5826 137 5831
rect 70 5822 137 5826
rect 43 5819 137 5822
rect 43 5812 92 5819
rect 43 5806 73 5812
rect 92 5807 97 5812
rect 9 5790 89 5806
rect 101 5798 137 5819
rect 198 5814 387 5838
rect 432 5837 479 5838
rect 445 5832 479 5837
rect 213 5811 387 5814
rect 206 5808 387 5811
rect 415 5831 479 5832
rect 9 5788 28 5790
rect 43 5788 77 5790
rect 9 5772 89 5788
rect 9 5766 28 5772
rect -1 5750 28 5766
rect 43 5756 73 5772
rect 101 5750 107 5798
rect 110 5792 129 5798
rect 144 5792 174 5800
rect 110 5784 174 5792
rect 110 5768 190 5784
rect 206 5777 268 5808
rect 284 5777 346 5808
rect 415 5806 464 5831
rect 479 5806 509 5822
rect 378 5792 408 5800
rect 415 5798 525 5806
rect 378 5784 423 5792
rect 110 5766 129 5768
rect 144 5766 190 5768
rect 110 5750 190 5766
rect 217 5764 252 5777
rect 293 5774 330 5777
rect 293 5772 335 5774
rect 222 5761 252 5764
rect 231 5757 238 5761
rect 238 5756 239 5757
rect 197 5750 207 5756
rect -7 5742 34 5750
rect -7 5716 8 5742
rect 15 5716 34 5742
rect 98 5738 129 5750
rect 144 5738 247 5750
rect 259 5740 285 5766
rect 300 5761 330 5772
rect 362 5768 424 5784
rect 362 5766 408 5768
rect 362 5750 424 5766
rect 436 5750 442 5798
rect 445 5790 525 5798
rect 445 5788 464 5790
rect 479 5788 513 5790
rect 445 5772 525 5788
rect 445 5750 464 5772
rect 479 5756 509 5772
rect 537 5766 543 5840
rect 546 5766 565 5910
rect 580 5766 586 5910
rect 595 5840 608 5910
rect 660 5906 682 5910
rect 653 5884 682 5898
rect 735 5884 751 5898
rect 789 5894 795 5896
rect 802 5894 910 5910
rect 917 5894 923 5896
rect 931 5894 946 5910
rect 1012 5904 1031 5907
rect 653 5882 751 5884
rect 778 5882 946 5894
rect 961 5884 977 5898
rect 1012 5885 1034 5904
rect 1044 5898 1060 5899
rect 1043 5896 1060 5898
rect 1044 5891 1060 5896
rect 1034 5884 1040 5885
rect 1043 5884 1072 5891
rect 961 5883 1072 5884
rect 961 5882 1078 5883
rect 637 5874 688 5882
rect 735 5874 769 5882
rect 637 5862 662 5874
rect 669 5862 688 5874
rect 742 5872 769 5874
rect 778 5872 999 5882
rect 1034 5879 1040 5882
rect 742 5868 999 5872
rect 637 5854 688 5862
rect 735 5854 999 5868
rect 1043 5874 1078 5882
rect 589 5806 608 5840
rect 653 5846 682 5854
rect 653 5840 670 5846
rect 653 5838 687 5840
rect 735 5838 751 5854
rect 752 5844 960 5854
rect 961 5844 977 5854
rect 1025 5850 1040 5865
rect 1043 5862 1044 5874
rect 1051 5862 1078 5874
rect 1043 5854 1078 5862
rect 1043 5853 1072 5854
rect 763 5840 977 5844
rect 778 5838 977 5840
rect 1012 5840 1025 5850
rect 1043 5840 1060 5853
rect 1012 5838 1060 5840
rect 654 5834 687 5838
rect 650 5832 687 5834
rect 650 5831 717 5832
rect 650 5826 681 5831
rect 687 5826 717 5831
rect 650 5822 717 5826
rect 623 5819 717 5822
rect 623 5812 672 5819
rect 623 5806 653 5812
rect 672 5807 677 5812
rect 589 5790 669 5806
rect 681 5798 717 5819
rect 778 5814 967 5838
rect 1012 5837 1059 5838
rect 1025 5832 1059 5837
rect 793 5811 967 5814
rect 786 5808 967 5811
rect 995 5831 1059 5832
rect 589 5788 608 5790
rect 623 5788 657 5790
rect 589 5772 669 5788
rect 589 5766 608 5772
rect 305 5740 408 5750
rect 259 5738 408 5740
rect 429 5738 464 5750
rect 98 5736 260 5738
rect 110 5716 129 5736
rect 144 5734 174 5736
rect -7 5708 34 5716
rect 116 5712 129 5716
rect 181 5720 260 5736
rect 292 5736 464 5738
rect 292 5720 371 5736
rect 378 5734 408 5736
rect -1 5698 28 5708
rect 43 5698 73 5712
rect 116 5698 159 5712
rect 181 5708 371 5720
rect 436 5716 442 5736
rect 166 5698 196 5708
rect 197 5698 355 5708
rect 359 5698 389 5708
rect 393 5698 423 5712
rect 451 5698 464 5736
rect 536 5750 565 5766
rect 579 5750 608 5766
rect 623 5756 653 5772
rect 681 5750 687 5798
rect 690 5792 709 5798
rect 724 5792 754 5800
rect 690 5784 754 5792
rect 690 5768 770 5784
rect 786 5777 848 5808
rect 864 5777 926 5808
rect 995 5806 1044 5831
rect 1059 5806 1089 5822
rect 958 5792 988 5800
rect 995 5798 1105 5806
rect 958 5784 1003 5792
rect 690 5766 709 5768
rect 724 5766 770 5768
rect 690 5750 770 5766
rect 797 5764 832 5777
rect 873 5774 910 5777
rect 873 5772 915 5774
rect 802 5761 832 5764
rect 811 5757 818 5761
rect 818 5756 819 5757
rect 777 5750 787 5756
rect 536 5742 571 5750
rect 536 5716 537 5742
rect 544 5716 571 5742
rect 479 5698 509 5712
rect 536 5708 571 5716
rect 573 5742 614 5750
rect 573 5716 588 5742
rect 595 5716 614 5742
rect 678 5738 709 5750
rect 724 5738 827 5750
rect 839 5740 865 5766
rect 880 5761 910 5772
rect 942 5768 1004 5784
rect 942 5766 988 5768
rect 942 5750 1004 5766
rect 1016 5750 1022 5798
rect 1025 5790 1105 5798
rect 1025 5788 1044 5790
rect 1059 5788 1093 5790
rect 1025 5772 1105 5788
rect 1025 5750 1044 5772
rect 1059 5756 1089 5772
rect 1117 5766 1123 5840
rect 1126 5766 1145 5910
rect 1160 5766 1166 5910
rect 1175 5840 1188 5910
rect 1240 5906 1262 5910
rect 1233 5884 1262 5898
rect 1315 5884 1331 5898
rect 1369 5894 1375 5896
rect 1382 5894 1490 5910
rect 1497 5894 1503 5896
rect 1511 5894 1526 5910
rect 1592 5904 1611 5907
rect 1233 5882 1331 5884
rect 1358 5882 1526 5894
rect 1541 5884 1557 5898
rect 1592 5885 1614 5904
rect 1624 5898 1640 5899
rect 1623 5896 1640 5898
rect 1624 5891 1640 5896
rect 1614 5884 1620 5885
rect 1623 5884 1652 5891
rect 1541 5883 1652 5884
rect 1541 5882 1658 5883
rect 1217 5874 1268 5882
rect 1315 5874 1349 5882
rect 1217 5862 1242 5874
rect 1249 5862 1268 5874
rect 1322 5872 1349 5874
rect 1358 5872 1579 5882
rect 1614 5879 1620 5882
rect 1322 5868 1579 5872
rect 1217 5854 1268 5862
rect 1315 5854 1579 5868
rect 1623 5874 1658 5882
rect 1169 5806 1188 5840
rect 1233 5846 1262 5854
rect 1233 5840 1250 5846
rect 1233 5838 1267 5840
rect 1315 5838 1331 5854
rect 1332 5844 1540 5854
rect 1541 5844 1557 5854
rect 1605 5850 1620 5865
rect 1623 5862 1624 5874
rect 1631 5862 1658 5874
rect 1623 5854 1658 5862
rect 1623 5853 1652 5854
rect 1343 5840 1557 5844
rect 1358 5838 1557 5840
rect 1592 5840 1605 5850
rect 1623 5840 1640 5853
rect 1592 5838 1640 5840
rect 1234 5834 1267 5838
rect 1230 5832 1267 5834
rect 1230 5831 1297 5832
rect 1230 5826 1261 5831
rect 1267 5826 1297 5831
rect 1230 5822 1297 5826
rect 1203 5819 1297 5822
rect 1203 5812 1252 5819
rect 1203 5806 1233 5812
rect 1252 5807 1257 5812
rect 1169 5790 1249 5806
rect 1261 5798 1297 5819
rect 1358 5814 1547 5838
rect 1592 5837 1639 5838
rect 1605 5832 1639 5837
rect 1373 5811 1547 5814
rect 1366 5808 1547 5811
rect 1575 5831 1639 5832
rect 1169 5788 1188 5790
rect 1203 5788 1237 5790
rect 1169 5772 1249 5788
rect 1169 5766 1188 5772
rect 885 5740 988 5750
rect 839 5738 988 5740
rect 1009 5738 1044 5750
rect 678 5736 840 5738
rect 690 5716 709 5736
rect 724 5734 754 5736
rect 573 5708 614 5716
rect 696 5712 709 5716
rect 761 5720 840 5736
rect 872 5736 1044 5738
rect 872 5720 951 5736
rect 958 5734 988 5736
rect 536 5698 565 5708
rect 579 5698 608 5708
rect 623 5698 653 5712
rect 696 5698 739 5712
rect 761 5708 951 5720
rect 1016 5716 1022 5736
rect 746 5698 776 5708
rect 777 5698 935 5708
rect 939 5698 969 5708
rect 973 5698 1003 5712
rect 1031 5698 1044 5736
rect 1116 5750 1145 5766
rect 1159 5750 1188 5766
rect 1203 5756 1233 5772
rect 1261 5750 1267 5798
rect 1270 5792 1289 5798
rect 1304 5792 1334 5800
rect 1270 5784 1334 5792
rect 1270 5768 1350 5784
rect 1366 5777 1428 5808
rect 1444 5777 1506 5808
rect 1575 5806 1624 5831
rect 1639 5806 1669 5822
rect 1538 5792 1568 5800
rect 1575 5798 1685 5806
rect 1538 5784 1583 5792
rect 1270 5766 1289 5768
rect 1304 5766 1350 5768
rect 1270 5750 1350 5766
rect 1377 5764 1412 5777
rect 1453 5774 1490 5777
rect 1453 5772 1495 5774
rect 1382 5761 1412 5764
rect 1391 5757 1398 5761
rect 1398 5756 1399 5757
rect 1357 5750 1367 5756
rect 1116 5742 1151 5750
rect 1116 5716 1117 5742
rect 1124 5716 1151 5742
rect 1059 5698 1089 5712
rect 1116 5708 1151 5716
rect 1153 5742 1194 5750
rect 1153 5716 1168 5742
rect 1175 5716 1194 5742
rect 1258 5738 1289 5750
rect 1304 5738 1407 5750
rect 1419 5740 1445 5766
rect 1460 5761 1490 5772
rect 1522 5768 1584 5784
rect 1522 5766 1568 5768
rect 1522 5750 1584 5766
rect 1596 5750 1602 5798
rect 1605 5790 1685 5798
rect 1605 5788 1624 5790
rect 1639 5788 1673 5790
rect 1605 5772 1685 5788
rect 1605 5750 1624 5772
rect 1639 5756 1669 5772
rect 1697 5766 1703 5840
rect 1706 5766 1725 5910
rect 1740 5766 1746 5910
rect 1755 5840 1768 5910
rect 1820 5906 1842 5910
rect 1813 5884 1842 5898
rect 1895 5884 1911 5898
rect 1949 5894 1955 5896
rect 1962 5894 2070 5910
rect 2077 5894 2083 5896
rect 2091 5894 2106 5910
rect 2172 5904 2191 5907
rect 1813 5882 1911 5884
rect 1938 5882 2106 5894
rect 2121 5884 2137 5898
rect 2172 5885 2194 5904
rect 2204 5898 2220 5899
rect 2203 5896 2220 5898
rect 2204 5891 2220 5896
rect 2194 5884 2200 5885
rect 2203 5884 2232 5891
rect 2121 5883 2232 5884
rect 2121 5882 2238 5883
rect 1797 5874 1848 5882
rect 1895 5874 1929 5882
rect 1797 5862 1822 5874
rect 1829 5862 1848 5874
rect 1902 5872 1929 5874
rect 1938 5872 2159 5882
rect 2194 5879 2200 5882
rect 1902 5868 2159 5872
rect 1797 5854 1848 5862
rect 1895 5854 2159 5868
rect 2203 5874 2238 5882
rect 1749 5806 1768 5840
rect 1813 5846 1842 5854
rect 1813 5840 1830 5846
rect 1813 5838 1847 5840
rect 1895 5838 1911 5854
rect 1912 5844 2120 5854
rect 2121 5844 2137 5854
rect 2185 5850 2200 5865
rect 2203 5862 2204 5874
rect 2211 5862 2238 5874
rect 2203 5854 2238 5862
rect 2203 5853 2232 5854
rect 1923 5840 2137 5844
rect 1938 5838 2137 5840
rect 2172 5840 2185 5850
rect 2203 5840 2220 5853
rect 2172 5838 2220 5840
rect 1814 5834 1847 5838
rect 1810 5832 1847 5834
rect 1810 5831 1877 5832
rect 1810 5826 1841 5831
rect 1847 5826 1877 5831
rect 1810 5822 1877 5826
rect 1783 5819 1877 5822
rect 1783 5812 1832 5819
rect 1783 5806 1813 5812
rect 1832 5807 1837 5812
rect 1749 5790 1829 5806
rect 1841 5798 1877 5819
rect 1938 5814 2127 5838
rect 2172 5837 2219 5838
rect 2185 5832 2219 5837
rect 1953 5811 2127 5814
rect 1946 5808 2127 5811
rect 2155 5831 2219 5832
rect 1749 5788 1768 5790
rect 1783 5788 1817 5790
rect 1749 5772 1829 5788
rect 1749 5766 1768 5772
rect 1465 5740 1568 5750
rect 1419 5738 1568 5740
rect 1589 5738 1624 5750
rect 1258 5736 1420 5738
rect 1270 5716 1289 5736
rect 1304 5734 1334 5736
rect 1153 5708 1194 5716
rect 1276 5712 1289 5716
rect 1341 5720 1420 5736
rect 1452 5736 1624 5738
rect 1452 5720 1531 5736
rect 1538 5734 1568 5736
rect 1116 5698 1145 5708
rect 1159 5698 1188 5708
rect 1203 5698 1233 5712
rect 1276 5698 1319 5712
rect 1341 5708 1531 5720
rect 1596 5716 1602 5736
rect 1326 5698 1356 5708
rect 1357 5698 1515 5708
rect 1519 5698 1549 5708
rect 1553 5698 1583 5712
rect 1611 5698 1624 5736
rect 1696 5750 1725 5766
rect 1739 5750 1768 5766
rect 1783 5756 1813 5772
rect 1841 5750 1847 5798
rect 1850 5792 1869 5798
rect 1884 5792 1914 5800
rect 1850 5784 1914 5792
rect 1850 5768 1930 5784
rect 1946 5777 2008 5808
rect 2024 5777 2086 5808
rect 2155 5806 2204 5831
rect 2219 5806 2249 5822
rect 2118 5792 2148 5800
rect 2155 5798 2265 5806
rect 2118 5784 2163 5792
rect 1850 5766 1869 5768
rect 1884 5766 1930 5768
rect 1850 5750 1930 5766
rect 1957 5764 1992 5777
rect 2033 5774 2070 5777
rect 2033 5772 2075 5774
rect 1962 5761 1992 5764
rect 1971 5757 1978 5761
rect 1978 5756 1979 5757
rect 1937 5750 1947 5756
rect 1696 5742 1731 5750
rect 1696 5716 1697 5742
rect 1704 5716 1731 5742
rect 1639 5698 1669 5712
rect 1696 5708 1731 5716
rect 1733 5742 1774 5750
rect 1733 5716 1748 5742
rect 1755 5716 1774 5742
rect 1838 5738 1869 5750
rect 1884 5738 1987 5750
rect 1999 5740 2025 5766
rect 2040 5761 2070 5772
rect 2102 5768 2164 5784
rect 2102 5766 2148 5768
rect 2102 5750 2164 5766
rect 2176 5750 2182 5798
rect 2185 5790 2265 5798
rect 2185 5788 2204 5790
rect 2219 5788 2253 5790
rect 2185 5772 2265 5788
rect 2185 5750 2204 5772
rect 2219 5756 2249 5772
rect 2277 5766 2283 5840
rect 2286 5766 2305 5910
rect 2320 5766 2326 5910
rect 2335 5840 2348 5910
rect 2400 5906 2422 5910
rect 2393 5884 2422 5898
rect 2475 5884 2491 5898
rect 2529 5894 2535 5896
rect 2542 5894 2650 5910
rect 2657 5894 2663 5896
rect 2671 5894 2686 5910
rect 2752 5904 2771 5907
rect 2393 5882 2491 5884
rect 2518 5882 2686 5894
rect 2701 5884 2717 5898
rect 2752 5885 2774 5904
rect 2784 5898 2800 5899
rect 2783 5896 2800 5898
rect 2784 5891 2800 5896
rect 2774 5884 2780 5885
rect 2783 5884 2812 5891
rect 2701 5883 2812 5884
rect 2701 5882 2818 5883
rect 2377 5874 2428 5882
rect 2475 5874 2509 5882
rect 2377 5862 2402 5874
rect 2409 5862 2428 5874
rect 2482 5872 2509 5874
rect 2518 5872 2739 5882
rect 2774 5879 2780 5882
rect 2482 5868 2739 5872
rect 2377 5854 2428 5862
rect 2475 5854 2739 5868
rect 2783 5874 2818 5882
rect 2329 5806 2348 5840
rect 2393 5846 2422 5854
rect 2393 5840 2410 5846
rect 2393 5838 2427 5840
rect 2475 5838 2491 5854
rect 2492 5844 2700 5854
rect 2701 5844 2717 5854
rect 2765 5850 2780 5865
rect 2783 5862 2784 5874
rect 2791 5862 2818 5874
rect 2783 5854 2818 5862
rect 2783 5853 2812 5854
rect 2503 5840 2717 5844
rect 2518 5838 2717 5840
rect 2752 5840 2765 5850
rect 2783 5840 2800 5853
rect 2752 5838 2800 5840
rect 2394 5834 2427 5838
rect 2390 5832 2427 5834
rect 2390 5831 2457 5832
rect 2390 5826 2421 5831
rect 2427 5826 2457 5831
rect 2390 5822 2457 5826
rect 2363 5819 2457 5822
rect 2363 5812 2412 5819
rect 2363 5806 2393 5812
rect 2412 5807 2417 5812
rect 2329 5790 2409 5806
rect 2421 5798 2457 5819
rect 2518 5814 2707 5838
rect 2752 5837 2799 5838
rect 2765 5832 2799 5837
rect 2533 5811 2707 5814
rect 2526 5808 2707 5811
rect 2735 5831 2799 5832
rect 2329 5788 2348 5790
rect 2363 5788 2397 5790
rect 2329 5772 2409 5788
rect 2329 5766 2348 5772
rect 2045 5740 2148 5750
rect 1999 5738 2148 5740
rect 2169 5738 2204 5750
rect 1838 5736 2000 5738
rect 1850 5716 1869 5736
rect 1884 5734 1914 5736
rect 1733 5708 1774 5716
rect 1856 5712 1869 5716
rect 1921 5720 2000 5736
rect 2032 5736 2204 5738
rect 2032 5720 2111 5736
rect 2118 5734 2148 5736
rect 1696 5698 1725 5708
rect 1739 5698 1768 5708
rect 1783 5698 1813 5712
rect 1856 5698 1899 5712
rect 1921 5708 2111 5720
rect 2176 5716 2182 5736
rect 1906 5698 1936 5708
rect 1937 5698 2095 5708
rect 2099 5698 2129 5708
rect 2133 5698 2163 5712
rect 2191 5698 2204 5736
rect 2276 5750 2305 5766
rect 2319 5750 2348 5766
rect 2363 5756 2393 5772
rect 2421 5750 2427 5798
rect 2430 5792 2449 5798
rect 2464 5792 2494 5800
rect 2430 5784 2494 5792
rect 2430 5768 2510 5784
rect 2526 5777 2588 5808
rect 2604 5777 2666 5808
rect 2735 5806 2784 5831
rect 2799 5806 2829 5822
rect 2698 5792 2728 5800
rect 2735 5798 2845 5806
rect 2698 5784 2743 5792
rect 2430 5766 2449 5768
rect 2464 5766 2510 5768
rect 2430 5750 2510 5766
rect 2537 5764 2572 5777
rect 2613 5774 2650 5777
rect 2613 5772 2655 5774
rect 2542 5761 2572 5764
rect 2551 5757 2558 5761
rect 2558 5756 2559 5757
rect 2517 5750 2527 5756
rect 2276 5742 2311 5750
rect 2276 5716 2277 5742
rect 2284 5716 2311 5742
rect 2219 5698 2249 5712
rect 2276 5708 2311 5716
rect 2313 5742 2354 5750
rect 2313 5716 2328 5742
rect 2335 5716 2354 5742
rect 2418 5738 2449 5750
rect 2464 5738 2567 5750
rect 2579 5740 2605 5766
rect 2620 5761 2650 5772
rect 2682 5768 2744 5784
rect 2682 5766 2728 5768
rect 2682 5750 2744 5766
rect 2756 5750 2762 5798
rect 2765 5790 2845 5798
rect 2765 5788 2784 5790
rect 2799 5788 2833 5790
rect 2765 5772 2845 5788
rect 2765 5750 2784 5772
rect 2799 5756 2829 5772
rect 2857 5766 2863 5840
rect 2866 5766 2885 5910
rect 2900 5766 2906 5910
rect 2915 5840 2928 5910
rect 2980 5906 3002 5910
rect 2973 5884 3002 5898
rect 3055 5884 3071 5898
rect 3109 5894 3115 5896
rect 3122 5894 3230 5910
rect 3237 5894 3243 5896
rect 3251 5894 3266 5910
rect 3332 5904 3351 5907
rect 2973 5882 3071 5884
rect 3098 5882 3266 5894
rect 3281 5884 3297 5898
rect 3332 5885 3354 5904
rect 3364 5898 3380 5899
rect 3363 5896 3380 5898
rect 3364 5891 3380 5896
rect 3354 5884 3360 5885
rect 3363 5884 3392 5891
rect 3281 5883 3392 5884
rect 3281 5882 3398 5883
rect 2957 5874 3008 5882
rect 3055 5874 3089 5882
rect 2957 5862 2982 5874
rect 2989 5862 3008 5874
rect 3062 5872 3089 5874
rect 3098 5872 3319 5882
rect 3354 5879 3360 5882
rect 3062 5868 3319 5872
rect 2957 5854 3008 5862
rect 3055 5854 3319 5868
rect 3363 5874 3398 5882
rect 2909 5806 2928 5840
rect 2973 5846 3002 5854
rect 2973 5840 2990 5846
rect 2973 5838 3007 5840
rect 3055 5838 3071 5854
rect 3072 5844 3280 5854
rect 3281 5844 3297 5854
rect 3345 5850 3360 5865
rect 3363 5862 3364 5874
rect 3371 5862 3398 5874
rect 3363 5854 3398 5862
rect 3363 5853 3392 5854
rect 3083 5840 3297 5844
rect 3098 5838 3297 5840
rect 3332 5840 3345 5850
rect 3363 5840 3380 5853
rect 3332 5838 3380 5840
rect 2974 5834 3007 5838
rect 2970 5832 3007 5834
rect 2970 5831 3037 5832
rect 2970 5826 3001 5831
rect 3007 5826 3037 5831
rect 2970 5822 3037 5826
rect 2943 5819 3037 5822
rect 2943 5812 2992 5819
rect 2943 5806 2973 5812
rect 2992 5807 2997 5812
rect 2909 5790 2989 5806
rect 3001 5798 3037 5819
rect 3098 5814 3287 5838
rect 3332 5837 3379 5838
rect 3345 5832 3379 5837
rect 3113 5811 3287 5814
rect 3106 5808 3287 5811
rect 3315 5831 3379 5832
rect 2909 5788 2928 5790
rect 2943 5788 2977 5790
rect 2909 5772 2989 5788
rect 2909 5766 2928 5772
rect 2625 5740 2728 5750
rect 2579 5738 2728 5740
rect 2749 5738 2784 5750
rect 2418 5736 2580 5738
rect 2430 5716 2449 5736
rect 2464 5734 2494 5736
rect 2313 5708 2354 5716
rect 2436 5712 2449 5716
rect 2501 5720 2580 5736
rect 2612 5736 2784 5738
rect 2612 5720 2691 5736
rect 2698 5734 2728 5736
rect 2276 5698 2305 5708
rect 2319 5698 2348 5708
rect 2363 5698 2393 5712
rect 2436 5698 2479 5712
rect 2501 5708 2691 5720
rect 2756 5716 2762 5736
rect 2486 5698 2516 5708
rect 2517 5698 2675 5708
rect 2679 5698 2709 5708
rect 2713 5698 2743 5712
rect 2771 5698 2784 5736
rect 2856 5750 2885 5766
rect 2899 5750 2928 5766
rect 2943 5756 2973 5772
rect 3001 5750 3007 5798
rect 3010 5792 3029 5798
rect 3044 5792 3074 5800
rect 3010 5784 3074 5792
rect 3010 5768 3090 5784
rect 3106 5777 3168 5808
rect 3184 5777 3246 5808
rect 3315 5806 3364 5831
rect 3379 5806 3409 5822
rect 3278 5792 3308 5800
rect 3315 5798 3425 5806
rect 3278 5784 3323 5792
rect 3010 5766 3029 5768
rect 3044 5766 3090 5768
rect 3010 5750 3090 5766
rect 3117 5764 3152 5777
rect 3193 5774 3230 5777
rect 3193 5772 3235 5774
rect 3122 5761 3152 5764
rect 3131 5757 3138 5761
rect 3138 5756 3139 5757
rect 3097 5750 3107 5756
rect 2856 5742 2891 5750
rect 2856 5716 2857 5742
rect 2864 5716 2891 5742
rect 2799 5698 2829 5712
rect 2856 5708 2891 5716
rect 2893 5742 2934 5750
rect 2893 5716 2908 5742
rect 2915 5716 2934 5742
rect 2998 5738 3029 5750
rect 3044 5738 3147 5750
rect 3159 5740 3185 5766
rect 3200 5761 3230 5772
rect 3262 5768 3324 5784
rect 3262 5766 3308 5768
rect 3262 5750 3324 5766
rect 3336 5750 3342 5798
rect 3345 5790 3425 5798
rect 3345 5788 3364 5790
rect 3379 5788 3413 5790
rect 3345 5772 3425 5788
rect 3345 5750 3364 5772
rect 3379 5756 3409 5772
rect 3437 5766 3443 5840
rect 3446 5766 3465 5910
rect 3480 5766 3486 5910
rect 3495 5840 3508 5910
rect 3560 5906 3582 5910
rect 3553 5884 3582 5898
rect 3635 5884 3651 5898
rect 3689 5894 3695 5896
rect 3702 5894 3810 5910
rect 3817 5894 3823 5896
rect 3831 5894 3846 5910
rect 3912 5904 3931 5907
rect 3553 5882 3651 5884
rect 3678 5882 3846 5894
rect 3861 5884 3877 5898
rect 3912 5885 3934 5904
rect 3944 5898 3960 5899
rect 3943 5896 3960 5898
rect 3944 5891 3960 5896
rect 3934 5884 3940 5885
rect 3943 5884 3972 5891
rect 3861 5883 3972 5884
rect 3861 5882 3978 5883
rect 3537 5874 3588 5882
rect 3635 5874 3669 5882
rect 3537 5862 3562 5874
rect 3569 5862 3588 5874
rect 3642 5872 3669 5874
rect 3678 5872 3899 5882
rect 3934 5879 3940 5882
rect 3642 5868 3899 5872
rect 3537 5854 3588 5862
rect 3635 5854 3899 5868
rect 3943 5874 3978 5882
rect 3489 5806 3508 5840
rect 3553 5846 3582 5854
rect 3553 5840 3570 5846
rect 3553 5838 3587 5840
rect 3635 5838 3651 5854
rect 3652 5844 3860 5854
rect 3861 5844 3877 5854
rect 3925 5850 3940 5865
rect 3943 5862 3944 5874
rect 3951 5862 3978 5874
rect 3943 5854 3978 5862
rect 3943 5853 3972 5854
rect 3663 5840 3877 5844
rect 3678 5838 3877 5840
rect 3912 5840 3925 5850
rect 3943 5840 3960 5853
rect 3912 5838 3960 5840
rect 3554 5834 3587 5838
rect 3550 5832 3587 5834
rect 3550 5831 3617 5832
rect 3550 5826 3581 5831
rect 3587 5826 3617 5831
rect 3550 5822 3617 5826
rect 3523 5819 3617 5822
rect 3523 5812 3572 5819
rect 3523 5806 3553 5812
rect 3572 5807 3577 5812
rect 3489 5790 3569 5806
rect 3581 5798 3617 5819
rect 3678 5814 3867 5838
rect 3912 5837 3959 5838
rect 3925 5832 3959 5837
rect 3693 5811 3867 5814
rect 3686 5808 3867 5811
rect 3895 5831 3959 5832
rect 3489 5788 3508 5790
rect 3523 5788 3557 5790
rect 3489 5772 3569 5788
rect 3489 5766 3508 5772
rect 3205 5740 3308 5750
rect 3159 5738 3308 5740
rect 3329 5738 3364 5750
rect 2998 5736 3160 5738
rect 3010 5716 3029 5736
rect 3044 5734 3074 5736
rect 2893 5708 2934 5716
rect 3016 5712 3029 5716
rect 3081 5720 3160 5736
rect 3192 5736 3364 5738
rect 3192 5720 3271 5736
rect 3278 5734 3308 5736
rect 2856 5698 2885 5708
rect 2899 5698 2928 5708
rect 2943 5698 2973 5712
rect 3016 5698 3059 5712
rect 3081 5708 3271 5720
rect 3336 5716 3342 5736
rect 3066 5698 3096 5708
rect 3097 5698 3255 5708
rect 3259 5698 3289 5708
rect 3293 5698 3323 5712
rect 3351 5698 3364 5736
rect 3436 5750 3465 5766
rect 3479 5750 3508 5766
rect 3523 5756 3553 5772
rect 3581 5750 3587 5798
rect 3590 5792 3609 5798
rect 3624 5792 3654 5800
rect 3590 5784 3654 5792
rect 3590 5768 3670 5784
rect 3686 5777 3748 5808
rect 3764 5777 3826 5808
rect 3895 5806 3944 5831
rect 3959 5806 3989 5822
rect 3858 5792 3888 5800
rect 3895 5798 4005 5806
rect 3858 5784 3903 5792
rect 3590 5766 3609 5768
rect 3624 5766 3670 5768
rect 3590 5750 3670 5766
rect 3697 5764 3732 5777
rect 3773 5774 3810 5777
rect 3773 5772 3815 5774
rect 3702 5761 3732 5764
rect 3711 5757 3718 5761
rect 3718 5756 3719 5757
rect 3677 5750 3687 5756
rect 3436 5742 3471 5750
rect 3436 5716 3437 5742
rect 3444 5716 3471 5742
rect 3379 5698 3409 5712
rect 3436 5708 3471 5716
rect 3473 5742 3514 5750
rect 3473 5716 3488 5742
rect 3495 5716 3514 5742
rect 3578 5738 3609 5750
rect 3624 5738 3727 5750
rect 3739 5740 3765 5766
rect 3780 5761 3810 5772
rect 3842 5768 3904 5784
rect 3842 5766 3888 5768
rect 3842 5750 3904 5766
rect 3916 5750 3922 5798
rect 3925 5790 4005 5798
rect 3925 5788 3944 5790
rect 3959 5788 3993 5790
rect 3925 5772 4005 5788
rect 3925 5750 3944 5772
rect 3959 5756 3989 5772
rect 4017 5766 4023 5840
rect 4026 5766 4045 5910
rect 4060 5766 4066 5910
rect 4075 5840 4088 5910
rect 4140 5906 4162 5910
rect 4133 5884 4162 5898
rect 4215 5884 4231 5898
rect 4269 5894 4275 5896
rect 4282 5894 4390 5910
rect 4397 5894 4403 5896
rect 4411 5894 4426 5910
rect 4492 5904 4511 5907
rect 4133 5882 4231 5884
rect 4258 5882 4426 5894
rect 4441 5884 4457 5898
rect 4492 5885 4514 5904
rect 4524 5898 4540 5899
rect 4523 5896 4540 5898
rect 4524 5891 4540 5896
rect 4514 5884 4520 5885
rect 4523 5884 4552 5891
rect 4441 5883 4552 5884
rect 4441 5882 4558 5883
rect 4117 5874 4168 5882
rect 4215 5874 4249 5882
rect 4117 5862 4142 5874
rect 4149 5862 4168 5874
rect 4222 5872 4249 5874
rect 4258 5872 4479 5882
rect 4514 5879 4520 5882
rect 4222 5868 4479 5872
rect 4117 5854 4168 5862
rect 4215 5854 4479 5868
rect 4523 5874 4558 5882
rect 4069 5806 4088 5840
rect 4133 5846 4162 5854
rect 4133 5840 4150 5846
rect 4133 5838 4167 5840
rect 4215 5838 4231 5854
rect 4232 5844 4440 5854
rect 4441 5844 4457 5854
rect 4505 5850 4520 5865
rect 4523 5862 4524 5874
rect 4531 5862 4558 5874
rect 4523 5854 4558 5862
rect 4523 5853 4552 5854
rect 4243 5840 4457 5844
rect 4258 5838 4457 5840
rect 4492 5840 4505 5850
rect 4523 5840 4540 5853
rect 4492 5838 4540 5840
rect 4134 5834 4167 5838
rect 4130 5832 4167 5834
rect 4130 5831 4197 5832
rect 4130 5826 4161 5831
rect 4167 5826 4197 5831
rect 4130 5822 4197 5826
rect 4103 5819 4197 5822
rect 4103 5812 4152 5819
rect 4103 5806 4133 5812
rect 4152 5807 4157 5812
rect 4069 5790 4149 5806
rect 4161 5798 4197 5819
rect 4258 5814 4447 5838
rect 4492 5837 4539 5838
rect 4505 5832 4539 5837
rect 4273 5811 4447 5814
rect 4266 5808 4447 5811
rect 4475 5831 4539 5832
rect 4069 5788 4088 5790
rect 4103 5788 4137 5790
rect 4069 5772 4149 5788
rect 4069 5766 4088 5772
rect 3785 5740 3888 5750
rect 3739 5738 3888 5740
rect 3909 5738 3944 5750
rect 3578 5736 3740 5738
rect 3590 5716 3609 5736
rect 3624 5734 3654 5736
rect 3473 5708 3514 5716
rect 3596 5712 3609 5716
rect 3661 5720 3740 5736
rect 3772 5736 3944 5738
rect 3772 5720 3851 5736
rect 3858 5734 3888 5736
rect 3436 5698 3465 5708
rect 3479 5698 3508 5708
rect 3523 5698 3553 5712
rect 3596 5698 3639 5712
rect 3661 5708 3851 5720
rect 3916 5716 3922 5736
rect 3646 5698 3676 5708
rect 3677 5698 3835 5708
rect 3839 5698 3869 5708
rect 3873 5698 3903 5712
rect 3931 5698 3944 5736
rect 4016 5750 4045 5766
rect 4059 5750 4088 5766
rect 4103 5756 4133 5772
rect 4161 5750 4167 5798
rect 4170 5792 4189 5798
rect 4204 5792 4234 5800
rect 4170 5784 4234 5792
rect 4170 5768 4250 5784
rect 4266 5777 4328 5808
rect 4344 5777 4406 5808
rect 4475 5806 4524 5831
rect 4539 5806 4569 5822
rect 4438 5792 4468 5800
rect 4475 5798 4585 5806
rect 4438 5784 4483 5792
rect 4170 5766 4189 5768
rect 4204 5766 4250 5768
rect 4170 5750 4250 5766
rect 4277 5764 4312 5777
rect 4353 5774 4390 5777
rect 4353 5772 4395 5774
rect 4282 5761 4312 5764
rect 4291 5757 4298 5761
rect 4298 5756 4299 5757
rect 4257 5750 4267 5756
rect 4016 5742 4051 5750
rect 4016 5716 4017 5742
rect 4024 5716 4051 5742
rect 3959 5698 3989 5712
rect 4016 5708 4051 5716
rect 4053 5742 4094 5750
rect 4053 5716 4068 5742
rect 4075 5716 4094 5742
rect 4158 5738 4189 5750
rect 4204 5738 4307 5750
rect 4319 5740 4345 5766
rect 4360 5761 4390 5772
rect 4422 5768 4484 5784
rect 4422 5766 4468 5768
rect 4422 5750 4484 5766
rect 4496 5750 4502 5798
rect 4505 5790 4585 5798
rect 4505 5788 4524 5790
rect 4539 5788 4573 5790
rect 4505 5772 4585 5788
rect 4505 5750 4524 5772
rect 4539 5756 4569 5772
rect 4597 5766 4603 5840
rect 4606 5766 4625 5910
rect 4640 5766 4646 5910
rect 4655 5840 4668 5910
rect 4720 5906 4742 5910
rect 4713 5884 4742 5898
rect 4795 5884 4811 5898
rect 4849 5894 4855 5896
rect 4862 5894 4970 5910
rect 4977 5894 4983 5896
rect 4991 5894 5006 5910
rect 5072 5904 5091 5907
rect 4713 5882 4811 5884
rect 4838 5882 5006 5894
rect 5021 5884 5037 5898
rect 5072 5885 5094 5904
rect 5104 5898 5120 5899
rect 5103 5896 5120 5898
rect 5104 5891 5120 5896
rect 5094 5884 5100 5885
rect 5103 5884 5132 5891
rect 5021 5883 5132 5884
rect 5021 5882 5138 5883
rect 4697 5874 4748 5882
rect 4795 5874 4829 5882
rect 4697 5862 4722 5874
rect 4729 5862 4748 5874
rect 4802 5872 4829 5874
rect 4838 5872 5059 5882
rect 5094 5879 5100 5882
rect 4802 5868 5059 5872
rect 4697 5854 4748 5862
rect 4795 5854 5059 5868
rect 5103 5874 5138 5882
rect 4649 5806 4668 5840
rect 4713 5846 4742 5854
rect 4713 5840 4730 5846
rect 4713 5838 4747 5840
rect 4795 5838 4811 5854
rect 4812 5844 5020 5854
rect 5021 5844 5037 5854
rect 5085 5850 5100 5865
rect 5103 5862 5104 5874
rect 5111 5862 5138 5874
rect 5103 5854 5138 5862
rect 5103 5853 5132 5854
rect 4823 5840 5037 5844
rect 4838 5838 5037 5840
rect 5072 5840 5085 5850
rect 5103 5840 5120 5853
rect 5072 5838 5120 5840
rect 4714 5834 4747 5838
rect 4710 5832 4747 5834
rect 4710 5831 4777 5832
rect 4710 5826 4741 5831
rect 4747 5826 4777 5831
rect 4710 5822 4777 5826
rect 4683 5819 4777 5822
rect 4683 5812 4732 5819
rect 4683 5806 4713 5812
rect 4732 5807 4737 5812
rect 4649 5790 4729 5806
rect 4741 5798 4777 5819
rect 4838 5814 5027 5838
rect 5072 5837 5119 5838
rect 5085 5832 5119 5837
rect 4853 5811 5027 5814
rect 4846 5808 5027 5811
rect 5055 5831 5119 5832
rect 4649 5788 4668 5790
rect 4683 5788 4717 5790
rect 4649 5772 4729 5788
rect 4649 5766 4668 5772
rect 4365 5740 4468 5750
rect 4319 5738 4468 5740
rect 4489 5738 4524 5750
rect 4158 5736 4320 5738
rect 4170 5716 4189 5736
rect 4204 5734 4234 5736
rect 4053 5708 4094 5716
rect 4176 5712 4189 5716
rect 4241 5720 4320 5736
rect 4352 5736 4524 5738
rect 4352 5720 4431 5736
rect 4438 5734 4468 5736
rect 4016 5698 4045 5708
rect 4059 5698 4088 5708
rect 4103 5698 4133 5712
rect 4176 5698 4219 5712
rect 4241 5708 4431 5720
rect 4496 5716 4502 5736
rect 4226 5698 4256 5708
rect 4257 5698 4415 5708
rect 4419 5698 4449 5708
rect 4453 5698 4483 5712
rect 4511 5698 4524 5736
rect 4596 5750 4625 5766
rect 4639 5750 4668 5766
rect 4683 5756 4713 5772
rect 4741 5750 4747 5798
rect 4750 5792 4769 5798
rect 4784 5792 4814 5800
rect 4750 5784 4814 5792
rect 4750 5768 4830 5784
rect 4846 5777 4908 5808
rect 4924 5777 4986 5808
rect 5055 5806 5104 5831
rect 5119 5806 5149 5822
rect 5018 5792 5048 5800
rect 5055 5798 5165 5806
rect 5018 5784 5063 5792
rect 4750 5766 4769 5768
rect 4784 5766 4830 5768
rect 4750 5750 4830 5766
rect 4857 5764 4892 5777
rect 4933 5774 4970 5777
rect 4933 5772 4975 5774
rect 4862 5761 4892 5764
rect 4871 5757 4878 5761
rect 4878 5756 4879 5757
rect 4837 5750 4847 5756
rect 4596 5742 4631 5750
rect 4596 5716 4597 5742
rect 4604 5716 4631 5742
rect 4539 5698 4569 5712
rect 4596 5708 4631 5716
rect 4633 5742 4674 5750
rect 4633 5716 4648 5742
rect 4655 5716 4674 5742
rect 4738 5738 4769 5750
rect 4784 5738 4887 5750
rect 4899 5740 4925 5766
rect 4940 5761 4970 5772
rect 5002 5768 5064 5784
rect 5002 5766 5048 5768
rect 5002 5750 5064 5766
rect 5076 5750 5082 5798
rect 5085 5790 5165 5798
rect 5085 5788 5104 5790
rect 5119 5788 5153 5790
rect 5085 5772 5165 5788
rect 5085 5750 5104 5772
rect 5119 5756 5149 5772
rect 5177 5766 5183 5840
rect 5186 5766 5205 5910
rect 5220 5766 5226 5910
rect 5235 5840 5248 5910
rect 5300 5906 5322 5910
rect 5293 5884 5322 5898
rect 5375 5884 5391 5898
rect 5429 5894 5435 5896
rect 5442 5894 5550 5910
rect 5557 5894 5563 5896
rect 5571 5894 5586 5910
rect 5652 5904 5671 5907
rect 5293 5882 5391 5884
rect 5418 5882 5586 5894
rect 5601 5884 5617 5898
rect 5652 5885 5674 5904
rect 5684 5898 5700 5899
rect 5683 5896 5700 5898
rect 5684 5891 5700 5896
rect 5674 5884 5680 5885
rect 5683 5884 5712 5891
rect 5601 5883 5712 5884
rect 5601 5882 5718 5883
rect 5277 5874 5328 5882
rect 5375 5874 5409 5882
rect 5277 5862 5302 5874
rect 5309 5862 5328 5874
rect 5382 5872 5409 5874
rect 5418 5872 5639 5882
rect 5674 5879 5680 5882
rect 5382 5868 5639 5872
rect 5277 5854 5328 5862
rect 5375 5854 5639 5868
rect 5683 5874 5718 5882
rect 5229 5806 5248 5840
rect 5293 5846 5322 5854
rect 5293 5840 5310 5846
rect 5293 5838 5327 5840
rect 5375 5838 5391 5854
rect 5392 5844 5600 5854
rect 5601 5844 5617 5854
rect 5665 5850 5680 5865
rect 5683 5862 5684 5874
rect 5691 5862 5718 5874
rect 5683 5854 5718 5862
rect 5683 5853 5712 5854
rect 5403 5840 5617 5844
rect 5418 5838 5617 5840
rect 5652 5840 5665 5850
rect 5683 5840 5700 5853
rect 5652 5838 5700 5840
rect 5294 5834 5327 5838
rect 5290 5832 5327 5834
rect 5290 5831 5357 5832
rect 5290 5826 5321 5831
rect 5327 5826 5357 5831
rect 5290 5822 5357 5826
rect 5263 5819 5357 5822
rect 5263 5812 5312 5819
rect 5263 5806 5293 5812
rect 5312 5807 5317 5812
rect 5229 5790 5309 5806
rect 5321 5798 5357 5819
rect 5418 5814 5607 5838
rect 5652 5837 5699 5838
rect 5665 5832 5699 5837
rect 5433 5811 5607 5814
rect 5426 5808 5607 5811
rect 5635 5831 5699 5832
rect 5229 5788 5248 5790
rect 5263 5788 5297 5790
rect 5229 5772 5309 5788
rect 5229 5766 5248 5772
rect 4945 5740 5048 5750
rect 4899 5738 5048 5740
rect 5069 5738 5104 5750
rect 4738 5736 4900 5738
rect 4750 5716 4769 5736
rect 4784 5734 4814 5736
rect 4633 5708 4674 5716
rect 4756 5712 4769 5716
rect 4821 5720 4900 5736
rect 4932 5736 5104 5738
rect 4932 5720 5011 5736
rect 5018 5734 5048 5736
rect 4596 5698 4625 5708
rect 4639 5698 4668 5708
rect 4683 5698 4713 5712
rect 4756 5698 4799 5712
rect 4821 5708 5011 5720
rect 5076 5716 5082 5736
rect 4806 5698 4836 5708
rect 4837 5698 4995 5708
rect 4999 5698 5029 5708
rect 5033 5698 5063 5712
rect 5091 5698 5104 5736
rect 5176 5750 5205 5766
rect 5219 5750 5248 5766
rect 5263 5756 5293 5772
rect 5321 5750 5327 5798
rect 5330 5792 5349 5798
rect 5364 5792 5394 5800
rect 5330 5784 5394 5792
rect 5330 5768 5410 5784
rect 5426 5777 5488 5808
rect 5504 5777 5566 5808
rect 5635 5806 5684 5831
rect 5699 5806 5729 5822
rect 5598 5792 5628 5800
rect 5635 5798 5745 5806
rect 5598 5784 5643 5792
rect 5330 5766 5349 5768
rect 5364 5766 5410 5768
rect 5330 5750 5410 5766
rect 5437 5764 5472 5777
rect 5513 5774 5550 5777
rect 5513 5772 5555 5774
rect 5442 5761 5472 5764
rect 5451 5757 5458 5761
rect 5458 5756 5459 5757
rect 5417 5750 5427 5756
rect 5176 5742 5211 5750
rect 5176 5716 5177 5742
rect 5184 5716 5211 5742
rect 5119 5698 5149 5712
rect 5176 5708 5211 5716
rect 5213 5742 5254 5750
rect 5213 5716 5228 5742
rect 5235 5716 5254 5742
rect 5318 5738 5349 5750
rect 5364 5738 5467 5750
rect 5479 5740 5505 5766
rect 5520 5761 5550 5772
rect 5582 5768 5644 5784
rect 5582 5766 5628 5768
rect 5582 5750 5644 5766
rect 5656 5750 5662 5798
rect 5665 5790 5745 5798
rect 5665 5788 5684 5790
rect 5699 5788 5733 5790
rect 5665 5772 5745 5788
rect 5665 5750 5684 5772
rect 5699 5756 5729 5772
rect 5757 5766 5763 5840
rect 5766 5766 5785 5910
rect 5800 5766 5806 5910
rect 5815 5840 5828 5910
rect 5880 5906 5902 5910
rect 5873 5884 5902 5898
rect 5955 5884 5971 5898
rect 6009 5894 6015 5896
rect 6022 5894 6130 5910
rect 6137 5894 6143 5896
rect 6151 5894 6166 5910
rect 6232 5904 6251 5907
rect 5873 5882 5971 5884
rect 5998 5882 6166 5894
rect 6181 5884 6197 5898
rect 6232 5885 6254 5904
rect 6264 5898 6280 5899
rect 6263 5896 6280 5898
rect 6264 5891 6280 5896
rect 6254 5884 6260 5885
rect 6263 5884 6292 5891
rect 6181 5883 6292 5884
rect 6181 5882 6298 5883
rect 5857 5874 5908 5882
rect 5955 5874 5989 5882
rect 5857 5862 5882 5874
rect 5889 5862 5908 5874
rect 5962 5872 5989 5874
rect 5998 5872 6219 5882
rect 6254 5879 6260 5882
rect 5962 5868 6219 5872
rect 5857 5854 5908 5862
rect 5955 5854 6219 5868
rect 6263 5874 6298 5882
rect 5809 5806 5828 5840
rect 5873 5846 5902 5854
rect 5873 5840 5890 5846
rect 5873 5838 5907 5840
rect 5955 5838 5971 5854
rect 5972 5844 6180 5854
rect 6181 5844 6197 5854
rect 6245 5850 6260 5865
rect 6263 5862 6264 5874
rect 6271 5862 6298 5874
rect 6263 5854 6298 5862
rect 6263 5853 6292 5854
rect 5983 5840 6197 5844
rect 5998 5838 6197 5840
rect 6232 5840 6245 5850
rect 6263 5840 6280 5853
rect 6232 5838 6280 5840
rect 5874 5834 5907 5838
rect 5870 5832 5907 5834
rect 5870 5831 5937 5832
rect 5870 5826 5901 5831
rect 5907 5826 5937 5831
rect 5870 5822 5937 5826
rect 5843 5819 5937 5822
rect 5843 5812 5892 5819
rect 5843 5806 5873 5812
rect 5892 5807 5897 5812
rect 5809 5790 5889 5806
rect 5901 5798 5937 5819
rect 5998 5814 6187 5838
rect 6232 5837 6279 5838
rect 6245 5832 6279 5837
rect 6013 5811 6187 5814
rect 6006 5808 6187 5811
rect 6215 5831 6279 5832
rect 5809 5788 5828 5790
rect 5843 5788 5877 5790
rect 5809 5772 5889 5788
rect 5809 5766 5828 5772
rect 5525 5740 5628 5750
rect 5479 5738 5628 5740
rect 5649 5738 5684 5750
rect 5318 5736 5480 5738
rect 5330 5716 5349 5736
rect 5364 5734 5394 5736
rect 5213 5708 5254 5716
rect 5336 5712 5349 5716
rect 5401 5720 5480 5736
rect 5512 5736 5684 5738
rect 5512 5720 5591 5736
rect 5598 5734 5628 5736
rect 5176 5698 5205 5708
rect 5219 5698 5248 5708
rect 5263 5698 5293 5712
rect 5336 5698 5379 5712
rect 5401 5708 5591 5720
rect 5656 5716 5662 5736
rect 5386 5698 5416 5708
rect 5417 5698 5575 5708
rect 5579 5698 5609 5708
rect 5613 5698 5643 5712
rect 5671 5698 5684 5736
rect 5756 5750 5785 5766
rect 5799 5750 5828 5766
rect 5843 5756 5873 5772
rect 5901 5750 5907 5798
rect 5910 5792 5929 5798
rect 5944 5792 5974 5800
rect 5910 5784 5974 5792
rect 5910 5768 5990 5784
rect 6006 5777 6068 5808
rect 6084 5777 6146 5808
rect 6215 5806 6264 5831
rect 6279 5806 6309 5822
rect 6178 5792 6208 5800
rect 6215 5798 6325 5806
rect 6178 5784 6223 5792
rect 5910 5766 5929 5768
rect 5944 5766 5990 5768
rect 5910 5750 5990 5766
rect 6017 5764 6052 5777
rect 6093 5774 6130 5777
rect 6093 5772 6135 5774
rect 6022 5761 6052 5764
rect 6031 5757 6038 5761
rect 6038 5756 6039 5757
rect 5997 5750 6007 5756
rect 5756 5742 5791 5750
rect 5756 5716 5757 5742
rect 5764 5716 5791 5742
rect 5699 5698 5729 5712
rect 5756 5708 5791 5716
rect 5793 5742 5834 5750
rect 5793 5716 5808 5742
rect 5815 5716 5834 5742
rect 5898 5738 5929 5750
rect 5944 5738 6047 5750
rect 6059 5740 6085 5766
rect 6100 5761 6130 5772
rect 6162 5768 6224 5784
rect 6162 5766 6208 5768
rect 6162 5750 6224 5766
rect 6236 5750 6242 5798
rect 6245 5790 6325 5798
rect 6245 5788 6264 5790
rect 6279 5788 6313 5790
rect 6245 5772 6325 5788
rect 6245 5750 6264 5772
rect 6279 5756 6309 5772
rect 6337 5766 6343 5840
rect 6346 5766 6365 5910
rect 6380 5766 6386 5910
rect 6395 5840 6408 5910
rect 6460 5906 6482 5910
rect 6453 5884 6482 5898
rect 6535 5884 6551 5898
rect 6589 5894 6595 5896
rect 6602 5894 6710 5910
rect 6717 5894 6723 5896
rect 6731 5894 6746 5910
rect 6812 5904 6831 5907
rect 6453 5882 6551 5884
rect 6578 5882 6746 5894
rect 6761 5884 6777 5898
rect 6812 5885 6834 5904
rect 6844 5898 6860 5899
rect 6843 5896 6860 5898
rect 6844 5891 6860 5896
rect 6834 5884 6840 5885
rect 6843 5884 6872 5891
rect 6761 5883 6872 5884
rect 6761 5882 6878 5883
rect 6437 5874 6488 5882
rect 6535 5874 6569 5882
rect 6437 5862 6462 5874
rect 6469 5862 6488 5874
rect 6542 5872 6569 5874
rect 6578 5872 6799 5882
rect 6834 5879 6840 5882
rect 6542 5868 6799 5872
rect 6437 5854 6488 5862
rect 6535 5854 6799 5868
rect 6843 5874 6878 5882
rect 6389 5806 6408 5840
rect 6453 5846 6482 5854
rect 6453 5840 6470 5846
rect 6453 5838 6487 5840
rect 6535 5838 6551 5854
rect 6552 5844 6760 5854
rect 6761 5844 6777 5854
rect 6825 5850 6840 5865
rect 6843 5862 6844 5874
rect 6851 5862 6878 5874
rect 6843 5854 6878 5862
rect 6843 5853 6872 5854
rect 6563 5840 6777 5844
rect 6578 5838 6777 5840
rect 6812 5840 6825 5850
rect 6843 5840 6860 5853
rect 6812 5838 6860 5840
rect 6454 5834 6487 5838
rect 6450 5832 6487 5834
rect 6450 5831 6517 5832
rect 6450 5826 6481 5831
rect 6487 5826 6517 5831
rect 6450 5822 6517 5826
rect 6423 5819 6517 5822
rect 6423 5812 6472 5819
rect 6423 5806 6453 5812
rect 6472 5807 6477 5812
rect 6389 5790 6469 5806
rect 6481 5798 6517 5819
rect 6578 5814 6767 5838
rect 6812 5837 6859 5838
rect 6825 5832 6859 5837
rect 6593 5811 6767 5814
rect 6586 5808 6767 5811
rect 6795 5831 6859 5832
rect 6389 5788 6408 5790
rect 6423 5788 6457 5790
rect 6389 5772 6469 5788
rect 6389 5766 6408 5772
rect 6105 5740 6208 5750
rect 6059 5738 6208 5740
rect 6229 5738 6264 5750
rect 5898 5736 6060 5738
rect 5910 5716 5929 5736
rect 5944 5734 5974 5736
rect 5793 5708 5834 5716
rect 5916 5712 5929 5716
rect 5981 5720 6060 5736
rect 6092 5736 6264 5738
rect 6092 5720 6171 5736
rect 6178 5734 6208 5736
rect 5756 5698 5785 5708
rect 5799 5698 5828 5708
rect 5843 5698 5873 5712
rect 5916 5698 5959 5712
rect 5981 5708 6171 5720
rect 6236 5716 6242 5736
rect 5966 5698 5996 5708
rect 5997 5698 6155 5708
rect 6159 5698 6189 5708
rect 6193 5698 6223 5712
rect 6251 5698 6264 5736
rect 6336 5750 6365 5766
rect 6379 5750 6408 5766
rect 6423 5756 6453 5772
rect 6481 5750 6487 5798
rect 6490 5792 6509 5798
rect 6524 5792 6554 5800
rect 6490 5784 6554 5792
rect 6490 5768 6570 5784
rect 6586 5777 6648 5808
rect 6664 5777 6726 5808
rect 6795 5806 6844 5831
rect 6859 5806 6889 5822
rect 6758 5792 6788 5800
rect 6795 5798 6905 5806
rect 6758 5784 6803 5792
rect 6490 5766 6509 5768
rect 6524 5766 6570 5768
rect 6490 5750 6570 5766
rect 6597 5764 6632 5777
rect 6673 5774 6710 5777
rect 6673 5772 6715 5774
rect 6602 5761 6632 5764
rect 6611 5757 6618 5761
rect 6618 5756 6619 5757
rect 6577 5750 6587 5756
rect 6336 5742 6371 5750
rect 6336 5716 6337 5742
rect 6344 5716 6371 5742
rect 6279 5698 6309 5712
rect 6336 5708 6371 5716
rect 6373 5742 6414 5750
rect 6373 5716 6388 5742
rect 6395 5716 6414 5742
rect 6478 5738 6509 5750
rect 6524 5738 6627 5750
rect 6639 5740 6665 5766
rect 6680 5761 6710 5772
rect 6742 5768 6804 5784
rect 6742 5766 6788 5768
rect 6742 5750 6804 5766
rect 6816 5750 6822 5798
rect 6825 5790 6905 5798
rect 6825 5788 6844 5790
rect 6859 5788 6893 5790
rect 6825 5772 6905 5788
rect 6825 5750 6844 5772
rect 6859 5756 6889 5772
rect 6917 5766 6923 5840
rect 6926 5766 6945 5910
rect 6960 5766 6966 5910
rect 6975 5840 6988 5910
rect 7040 5906 7062 5910
rect 7033 5884 7062 5898
rect 7115 5884 7131 5898
rect 7169 5894 7175 5896
rect 7182 5894 7290 5910
rect 7297 5894 7303 5896
rect 7311 5894 7326 5910
rect 7392 5904 7411 5907
rect 7033 5882 7131 5884
rect 7158 5882 7326 5894
rect 7341 5884 7357 5898
rect 7392 5885 7414 5904
rect 7424 5898 7440 5899
rect 7423 5896 7440 5898
rect 7424 5891 7440 5896
rect 7414 5884 7420 5885
rect 7423 5884 7452 5891
rect 7341 5883 7452 5884
rect 7341 5882 7458 5883
rect 7017 5874 7068 5882
rect 7115 5874 7149 5882
rect 7017 5862 7042 5874
rect 7049 5862 7068 5874
rect 7122 5872 7149 5874
rect 7158 5872 7379 5882
rect 7414 5879 7420 5882
rect 7122 5868 7379 5872
rect 7017 5854 7068 5862
rect 7115 5854 7379 5868
rect 7423 5874 7458 5882
rect 6969 5806 6988 5840
rect 7033 5846 7062 5854
rect 7033 5840 7050 5846
rect 7033 5838 7067 5840
rect 7115 5838 7131 5854
rect 7132 5844 7340 5854
rect 7341 5844 7357 5854
rect 7405 5850 7420 5865
rect 7423 5862 7424 5874
rect 7431 5862 7458 5874
rect 7423 5854 7458 5862
rect 7423 5853 7452 5854
rect 7143 5840 7357 5844
rect 7158 5838 7357 5840
rect 7392 5840 7405 5850
rect 7423 5840 7440 5853
rect 7392 5838 7440 5840
rect 7034 5834 7067 5838
rect 7030 5832 7067 5834
rect 7030 5831 7097 5832
rect 7030 5826 7061 5831
rect 7067 5826 7097 5831
rect 7030 5822 7097 5826
rect 7003 5819 7097 5822
rect 7003 5812 7052 5819
rect 7003 5806 7033 5812
rect 7052 5807 7057 5812
rect 6969 5790 7049 5806
rect 7061 5798 7097 5819
rect 7158 5814 7347 5838
rect 7392 5837 7439 5838
rect 7405 5832 7439 5837
rect 7173 5811 7347 5814
rect 7166 5808 7347 5811
rect 7375 5831 7439 5832
rect 6969 5788 6988 5790
rect 7003 5788 7037 5790
rect 6969 5772 7049 5788
rect 6969 5766 6988 5772
rect 6685 5740 6788 5750
rect 6639 5738 6788 5740
rect 6809 5738 6844 5750
rect 6478 5736 6640 5738
rect 6490 5716 6509 5736
rect 6524 5734 6554 5736
rect 6373 5708 6414 5716
rect 6496 5712 6509 5716
rect 6561 5720 6640 5736
rect 6672 5736 6844 5738
rect 6672 5720 6751 5736
rect 6758 5734 6788 5736
rect 6336 5698 6365 5708
rect 6379 5698 6408 5708
rect 6423 5698 6453 5712
rect 6496 5698 6539 5712
rect 6561 5708 6751 5720
rect 6816 5716 6822 5736
rect 6546 5698 6576 5708
rect 6577 5698 6735 5708
rect 6739 5698 6769 5708
rect 6773 5698 6803 5712
rect 6831 5698 6844 5736
rect 6916 5750 6945 5766
rect 6959 5750 6988 5766
rect 7003 5756 7033 5772
rect 7061 5750 7067 5798
rect 7070 5792 7089 5798
rect 7104 5792 7134 5800
rect 7070 5784 7134 5792
rect 7070 5768 7150 5784
rect 7166 5777 7228 5808
rect 7244 5777 7306 5808
rect 7375 5806 7424 5831
rect 7439 5806 7469 5822
rect 7338 5792 7368 5800
rect 7375 5798 7485 5806
rect 7338 5784 7383 5792
rect 7070 5766 7089 5768
rect 7104 5766 7150 5768
rect 7070 5750 7150 5766
rect 7177 5764 7212 5777
rect 7253 5774 7290 5777
rect 7253 5772 7295 5774
rect 7182 5761 7212 5764
rect 7191 5757 7198 5761
rect 7198 5756 7199 5757
rect 7157 5750 7167 5756
rect 6916 5742 6951 5750
rect 6916 5716 6917 5742
rect 6924 5716 6951 5742
rect 6859 5698 6889 5712
rect 6916 5708 6951 5716
rect 6953 5742 6994 5750
rect 6953 5716 6968 5742
rect 6975 5716 6994 5742
rect 7058 5738 7089 5750
rect 7104 5738 7207 5750
rect 7219 5740 7245 5766
rect 7260 5761 7290 5772
rect 7322 5768 7384 5784
rect 7322 5766 7368 5768
rect 7322 5750 7384 5766
rect 7396 5750 7402 5798
rect 7405 5790 7485 5798
rect 7405 5788 7424 5790
rect 7439 5788 7473 5790
rect 7405 5772 7485 5788
rect 7405 5750 7424 5772
rect 7439 5756 7469 5772
rect 7497 5766 7503 5840
rect 7506 5766 7525 5910
rect 7540 5766 7546 5910
rect 7555 5840 7568 5910
rect 7613 5888 7614 5898
rect 7629 5888 7642 5898
rect 7613 5884 7642 5888
rect 7647 5884 7677 5910
rect 7695 5896 7711 5898
rect 7783 5896 7836 5910
rect 7784 5894 7848 5896
rect 7891 5894 7906 5910
rect 7955 5907 7985 5910
rect 7955 5904 7991 5907
rect 7921 5896 7937 5898
rect 7695 5884 7710 5888
rect 7613 5882 7710 5884
rect 7738 5882 7906 5894
rect 7922 5884 7937 5888
rect 7955 5885 7994 5904
rect 8013 5898 8020 5899
rect 8019 5891 8020 5898
rect 8003 5888 8004 5891
rect 8019 5888 8032 5891
rect 7955 5884 7985 5885
rect 7994 5884 8000 5885
rect 8003 5884 8032 5888
rect 7922 5883 8032 5884
rect 7922 5882 8038 5883
rect 7597 5874 7648 5882
rect 7597 5862 7622 5874
rect 7629 5862 7648 5874
rect 7679 5874 7729 5882
rect 7679 5866 7695 5874
rect 7702 5872 7729 5874
rect 7738 5872 7959 5882
rect 7702 5862 7959 5872
rect 7988 5874 8038 5882
rect 7988 5865 8004 5874
rect 7597 5854 7648 5862
rect 7695 5854 7959 5862
rect 7985 5862 8004 5865
rect 8011 5862 8038 5874
rect 7985 5854 8038 5862
rect 7549 5806 7568 5840
rect 7613 5846 7614 5854
rect 7629 5846 7642 5854
rect 7613 5838 7629 5846
rect 7610 5831 7629 5834
rect 7610 5822 7632 5831
rect 7583 5812 7632 5822
rect 7583 5806 7613 5812
rect 7632 5807 7637 5812
rect 7549 5790 7629 5806
rect 7647 5798 7677 5854
rect 7712 5844 7920 5854
rect 7955 5850 8000 5854
rect 8003 5853 8004 5854
rect 8019 5853 8032 5854
rect 7738 5814 7927 5844
rect 7753 5811 7927 5814
rect 7746 5808 7927 5811
rect 7549 5788 7568 5790
rect 7583 5788 7617 5790
rect 7549 5772 7629 5788
rect 7656 5784 7669 5798
rect 7684 5784 7700 5800
rect 7746 5795 7757 5808
rect 7549 5766 7568 5772
rect 7265 5740 7368 5750
rect 7219 5738 7368 5740
rect 7389 5738 7424 5750
rect 7058 5736 7220 5738
rect 7070 5716 7089 5736
rect 7104 5734 7134 5736
rect 6953 5708 6994 5716
rect 7076 5712 7089 5716
rect 7141 5720 7220 5736
rect 7252 5736 7424 5738
rect 7252 5720 7331 5736
rect 7338 5734 7368 5736
rect 6916 5698 6945 5708
rect 6959 5698 6988 5708
rect 7003 5698 7033 5712
rect 7076 5698 7119 5712
rect 7141 5708 7331 5720
rect 7396 5716 7402 5736
rect 7126 5698 7156 5708
rect 7157 5698 7315 5708
rect 7319 5698 7349 5708
rect 7353 5698 7383 5712
rect 7411 5698 7424 5736
rect 7496 5750 7525 5766
rect 7539 5750 7568 5766
rect 7583 5750 7613 5772
rect 7656 5768 7718 5784
rect 7746 5777 7757 5793
rect 7762 5788 7772 5808
rect 7782 5788 7796 5808
rect 7799 5795 7808 5808
rect 7824 5795 7833 5808
rect 7762 5777 7796 5788
rect 7799 5777 7808 5793
rect 7824 5777 7833 5793
rect 7840 5788 7850 5808
rect 7860 5788 7874 5808
rect 7875 5795 7886 5808
rect 7840 5777 7874 5788
rect 7875 5777 7886 5793
rect 7932 5784 7948 5800
rect 7955 5798 7985 5850
rect 8019 5846 8020 5853
rect 8004 5838 8020 5846
rect 7991 5806 8004 5825
rect 8019 5806 8049 5822
rect 7991 5790 8065 5806
rect 7991 5788 8004 5790
rect 8019 5788 8053 5790
rect 7656 5766 7669 5768
rect 7684 5766 7718 5768
rect 7656 5750 7718 5766
rect 7762 5761 7778 5764
rect 7840 5761 7870 5772
rect 7918 5768 7964 5784
rect 7991 5772 8065 5788
rect 7918 5766 7952 5768
rect 7917 5750 7964 5766
rect 7991 5750 8004 5772
rect 8019 5750 8049 5772
rect 8076 5750 8077 5766
rect 8092 5750 8105 5910
rect 8135 5806 8148 5910
rect 8193 5888 8194 5898
rect 8209 5888 8222 5898
rect 8193 5884 8222 5888
rect 8227 5884 8257 5910
rect 8275 5896 8291 5898
rect 8363 5896 8416 5910
rect 8364 5894 8428 5896
rect 8471 5894 8486 5910
rect 8535 5907 8565 5910
rect 8535 5904 8571 5907
rect 8501 5896 8517 5898
rect 8275 5884 8290 5888
rect 8193 5882 8290 5884
rect 8318 5882 8486 5894
rect 8502 5884 8517 5888
rect 8535 5885 8574 5904
rect 8593 5898 8600 5899
rect 8599 5891 8600 5898
rect 8583 5888 8584 5891
rect 8599 5888 8612 5891
rect 8535 5884 8565 5885
rect 8574 5884 8580 5885
rect 8583 5884 8612 5888
rect 8502 5883 8612 5884
rect 8502 5882 8618 5883
rect 8177 5874 8228 5882
rect 8177 5862 8202 5874
rect 8209 5862 8228 5874
rect 8259 5874 8309 5882
rect 8259 5866 8275 5874
rect 8282 5872 8309 5874
rect 8318 5872 8539 5882
rect 8282 5862 8539 5872
rect 8568 5874 8618 5882
rect 8568 5865 8584 5874
rect 8177 5854 8228 5862
rect 8275 5854 8539 5862
rect 8565 5862 8584 5865
rect 8591 5862 8618 5874
rect 8565 5854 8618 5862
rect 8193 5846 8194 5854
rect 8209 5846 8222 5854
rect 8193 5838 8209 5846
rect 8190 5831 8209 5834
rect 8190 5822 8212 5831
rect 8163 5812 8212 5822
rect 8163 5806 8193 5812
rect 8212 5807 8217 5812
rect 8135 5790 8209 5806
rect 8227 5798 8257 5854
rect 8292 5844 8500 5854
rect 8535 5850 8580 5854
rect 8583 5853 8584 5854
rect 8599 5853 8612 5854
rect 8318 5814 8507 5844
rect 8333 5811 8507 5814
rect 8326 5808 8507 5811
rect 8135 5788 8148 5790
rect 8163 5788 8197 5790
rect 8135 5772 8209 5788
rect 8236 5784 8249 5798
rect 8264 5784 8280 5800
rect 8326 5795 8337 5808
rect 8119 5750 8120 5766
rect 8135 5750 8148 5772
rect 8163 5750 8193 5772
rect 8236 5768 8298 5784
rect 8326 5777 8337 5793
rect 8342 5788 8352 5808
rect 8362 5788 8376 5808
rect 8379 5795 8388 5808
rect 8404 5795 8413 5808
rect 8342 5777 8376 5788
rect 8379 5777 8388 5793
rect 8404 5777 8413 5793
rect 8420 5788 8430 5808
rect 8440 5788 8454 5808
rect 8455 5795 8466 5808
rect 8420 5777 8454 5788
rect 8455 5777 8466 5793
rect 8512 5784 8528 5800
rect 8535 5798 8565 5850
rect 8599 5846 8600 5853
rect 8584 5838 8600 5846
rect 8571 5806 8584 5825
rect 8599 5806 8629 5822
rect 8571 5790 8645 5806
rect 8571 5788 8584 5790
rect 8599 5788 8633 5790
rect 8236 5766 8249 5768
rect 8264 5766 8298 5768
rect 8236 5750 8298 5766
rect 8342 5761 8358 5764
rect 8420 5761 8450 5772
rect 8498 5768 8544 5784
rect 8571 5772 8645 5788
rect 8498 5766 8532 5768
rect 8497 5750 8544 5766
rect 8571 5750 8584 5772
rect 8599 5750 8629 5772
rect 8656 5750 8657 5766
rect 8672 5750 8685 5910
rect 8715 5806 8728 5910
rect 8773 5888 8774 5898
rect 8789 5888 8802 5898
rect 8773 5884 8802 5888
rect 8807 5884 8837 5910
rect 8855 5896 8871 5898
rect 8943 5896 8996 5910
rect 8944 5894 9008 5896
rect 9051 5894 9066 5910
rect 9115 5907 9145 5910
rect 9115 5904 9151 5907
rect 9081 5896 9097 5898
rect 8855 5884 8870 5888
rect 8773 5882 8870 5884
rect 8898 5882 9066 5894
rect 9082 5884 9097 5888
rect 9115 5885 9154 5904
rect 9173 5898 9180 5899
rect 9179 5891 9180 5898
rect 9163 5888 9164 5891
rect 9179 5888 9192 5891
rect 9115 5884 9145 5885
rect 9154 5884 9160 5885
rect 9163 5884 9192 5888
rect 9082 5883 9192 5884
rect 9082 5882 9198 5883
rect 8757 5874 8808 5882
rect 8757 5862 8782 5874
rect 8789 5862 8808 5874
rect 8839 5874 8889 5882
rect 8839 5866 8855 5874
rect 8862 5872 8889 5874
rect 8898 5872 9119 5882
rect 8862 5862 9119 5872
rect 9148 5874 9198 5882
rect 9148 5865 9164 5874
rect 8757 5854 8808 5862
rect 8855 5854 9119 5862
rect 9145 5862 9164 5865
rect 9171 5862 9198 5874
rect 9145 5854 9198 5862
rect 8773 5846 8774 5854
rect 8789 5846 8802 5854
rect 8773 5838 8789 5846
rect 8770 5831 8789 5834
rect 8770 5822 8792 5831
rect 8743 5812 8792 5822
rect 8743 5806 8773 5812
rect 8792 5807 8797 5812
rect 8715 5790 8789 5806
rect 8807 5798 8837 5854
rect 8872 5844 9080 5854
rect 9115 5850 9160 5854
rect 9163 5853 9164 5854
rect 9179 5853 9192 5854
rect 8898 5814 9087 5844
rect 8913 5811 9087 5814
rect 8906 5808 9087 5811
rect 8715 5788 8728 5790
rect 8743 5788 8777 5790
rect 8715 5772 8789 5788
rect 8816 5784 8829 5798
rect 8844 5784 8860 5800
rect 8906 5795 8917 5808
rect 8699 5750 8700 5766
rect 8715 5750 8728 5772
rect 8743 5750 8773 5772
rect 8816 5768 8878 5784
rect 8906 5777 8917 5793
rect 8922 5788 8932 5808
rect 8942 5788 8956 5808
rect 8959 5795 8968 5808
rect 8984 5795 8993 5808
rect 8922 5777 8956 5788
rect 8959 5777 8968 5793
rect 8984 5777 8993 5793
rect 9000 5788 9010 5808
rect 9020 5788 9034 5808
rect 9035 5795 9046 5808
rect 9000 5777 9034 5788
rect 9035 5777 9046 5793
rect 9092 5784 9108 5800
rect 9115 5798 9145 5850
rect 9179 5846 9180 5853
rect 9164 5838 9180 5846
rect 9151 5806 9164 5825
rect 9179 5806 9209 5822
rect 9151 5790 9225 5806
rect 9151 5788 9164 5790
rect 9179 5788 9213 5790
rect 8816 5766 8829 5768
rect 8844 5766 8878 5768
rect 8816 5750 8878 5766
rect 8922 5761 8938 5764
rect 9000 5761 9030 5772
rect 9078 5768 9124 5784
rect 9151 5772 9225 5788
rect 9078 5766 9112 5768
rect 9077 5750 9124 5766
rect 9151 5750 9164 5772
rect 9179 5750 9209 5772
rect 9236 5750 9237 5766
rect 9252 5750 9265 5910
rect 7496 5742 7531 5750
rect 7496 5716 7497 5742
rect 7504 5716 7531 5742
rect 7439 5698 7469 5712
rect 7496 5708 7531 5716
rect 7533 5742 7574 5750
rect 7533 5716 7548 5742
rect 7555 5716 7574 5742
rect 7638 5738 7700 5750
rect 7712 5738 7787 5750
rect 7845 5738 7920 5750
rect 7932 5738 7963 5750
rect 7969 5738 8004 5750
rect 7638 5736 7800 5738
rect 7533 5708 7574 5716
rect 7656 5712 7669 5736
rect 7684 5734 7699 5736
rect 7496 5698 7525 5708
rect 7539 5698 7568 5708
rect 7583 5698 7613 5712
rect 7656 5698 7699 5712
rect 7723 5709 7730 5716
rect 7733 5712 7800 5736
rect 7832 5736 8004 5738
rect 7802 5714 7830 5718
rect 7832 5714 7912 5736
rect 7933 5734 7948 5736
rect 7802 5712 7912 5714
rect 7733 5708 7912 5712
rect 7706 5698 7736 5708
rect 7738 5698 7891 5708
rect 7899 5698 7929 5708
rect 7933 5698 7963 5712
rect 7991 5698 8004 5736
rect 8076 5742 8111 5750
rect 8076 5716 8077 5742
rect 8084 5716 8111 5742
rect 8019 5698 8049 5712
rect 8076 5708 8111 5716
rect 8113 5742 8154 5750
rect 8113 5716 8128 5742
rect 8135 5716 8154 5742
rect 8218 5738 8280 5750
rect 8292 5738 8367 5750
rect 8425 5738 8500 5750
rect 8512 5738 8543 5750
rect 8549 5738 8584 5750
rect 8218 5736 8380 5738
rect 8113 5708 8154 5716
rect 8236 5712 8249 5736
rect 8264 5734 8279 5736
rect 8076 5698 8077 5708
rect 8092 5698 8105 5708
rect 8119 5698 8120 5708
rect 8135 5698 8148 5708
rect 8163 5698 8193 5712
rect 8236 5698 8279 5712
rect 8303 5709 8310 5716
rect 8313 5712 8380 5736
rect 8412 5736 8584 5738
rect 8382 5714 8410 5718
rect 8412 5714 8492 5736
rect 8513 5734 8528 5736
rect 8382 5712 8492 5714
rect 8313 5708 8492 5712
rect 8286 5698 8316 5708
rect 8318 5698 8471 5708
rect 8479 5698 8509 5708
rect 8513 5698 8543 5712
rect 8571 5698 8584 5736
rect 8656 5742 8691 5750
rect 8656 5716 8657 5742
rect 8664 5716 8691 5742
rect 8599 5698 8629 5712
rect 8656 5708 8691 5716
rect 8693 5742 8734 5750
rect 8693 5716 8708 5742
rect 8715 5716 8734 5742
rect 8798 5738 8860 5750
rect 8872 5738 8947 5750
rect 9005 5738 9080 5750
rect 9092 5738 9123 5750
rect 9129 5738 9164 5750
rect 8798 5736 8960 5738
rect 8693 5708 8734 5716
rect 8816 5712 8829 5736
rect 8844 5734 8859 5736
rect 8656 5698 8657 5708
rect 8672 5698 8685 5708
rect 8699 5698 8700 5708
rect 8715 5698 8728 5708
rect 8743 5698 8773 5712
rect 8816 5698 8859 5712
rect 8883 5709 8890 5716
rect 8893 5712 8960 5736
rect 8992 5736 9164 5738
rect 8962 5714 8990 5718
rect 8992 5714 9072 5736
rect 9093 5734 9108 5736
rect 8962 5712 9072 5714
rect 8893 5708 9072 5712
rect 8866 5698 8896 5708
rect 8898 5698 9051 5708
rect 9059 5698 9089 5708
rect 9093 5698 9123 5712
rect 9151 5698 9164 5736
rect 9236 5742 9271 5750
rect 9236 5716 9237 5742
rect 9244 5716 9271 5742
rect 9179 5698 9209 5712
rect 9236 5708 9271 5716
rect 9236 5698 9237 5708
rect 9252 5698 9265 5708
rect -1 5692 9265 5698
rect 0 5684 9265 5692
rect 15 5654 28 5684
rect 43 5670 73 5684
rect 116 5670 159 5684
rect 166 5670 386 5684
rect 393 5670 423 5684
rect 83 5656 98 5668
rect 117 5656 130 5670
rect 198 5666 351 5670
rect 80 5654 102 5656
rect 180 5654 372 5666
rect 451 5654 464 5684
rect 479 5670 509 5684
rect 546 5654 565 5684
rect 580 5654 586 5684
rect 595 5654 608 5684
rect 623 5670 653 5684
rect 696 5670 739 5684
rect 746 5670 966 5684
rect 973 5670 1003 5684
rect 663 5656 678 5668
rect 697 5656 710 5670
rect 778 5666 931 5670
rect 660 5654 682 5656
rect 760 5654 952 5666
rect 1031 5654 1044 5684
rect 1059 5670 1089 5684
rect 1126 5654 1145 5684
rect 1160 5654 1166 5684
rect 1175 5654 1188 5684
rect 1203 5670 1233 5684
rect 1276 5670 1319 5684
rect 1326 5670 1546 5684
rect 1553 5670 1583 5684
rect 1243 5656 1258 5668
rect 1277 5656 1290 5670
rect 1358 5666 1511 5670
rect 1240 5654 1262 5656
rect 1340 5654 1532 5666
rect 1611 5654 1624 5684
rect 1639 5670 1669 5684
rect 1706 5654 1725 5684
rect 1740 5654 1746 5684
rect 1755 5654 1768 5684
rect 1783 5670 1813 5684
rect 1856 5670 1899 5684
rect 1906 5670 2126 5684
rect 2133 5670 2163 5684
rect 1823 5656 1838 5668
rect 1857 5656 1870 5670
rect 1938 5666 2091 5670
rect 1820 5654 1842 5656
rect 1920 5654 2112 5666
rect 2191 5654 2204 5684
rect 2219 5670 2249 5684
rect 2286 5654 2305 5684
rect 2320 5654 2326 5684
rect 2335 5654 2348 5684
rect 2363 5670 2393 5684
rect 2436 5670 2479 5684
rect 2486 5670 2706 5684
rect 2713 5670 2743 5684
rect 2403 5656 2418 5668
rect 2437 5656 2450 5670
rect 2518 5666 2671 5670
rect 2400 5654 2422 5656
rect 2500 5654 2692 5666
rect 2771 5654 2784 5684
rect 2799 5670 2829 5684
rect 2866 5654 2885 5684
rect 2900 5654 2906 5684
rect 2915 5654 2928 5684
rect 2943 5670 2973 5684
rect 3016 5670 3059 5684
rect 3066 5670 3286 5684
rect 3293 5670 3323 5684
rect 2983 5656 2998 5668
rect 3017 5656 3030 5670
rect 3098 5666 3251 5670
rect 2980 5654 3002 5656
rect 3080 5654 3272 5666
rect 3351 5654 3364 5684
rect 3379 5670 3409 5684
rect 3446 5654 3465 5684
rect 3480 5654 3486 5684
rect 3495 5654 3508 5684
rect 3523 5670 3553 5684
rect 3596 5670 3639 5684
rect 3646 5670 3866 5684
rect 3873 5670 3903 5684
rect 3563 5656 3578 5668
rect 3597 5656 3610 5670
rect 3678 5666 3831 5670
rect 3560 5654 3582 5656
rect 3660 5654 3852 5666
rect 3931 5654 3944 5684
rect 3959 5670 3989 5684
rect 4026 5654 4045 5684
rect 4060 5654 4066 5684
rect 4075 5654 4088 5684
rect 4103 5670 4133 5684
rect 4176 5670 4219 5684
rect 4226 5670 4446 5684
rect 4453 5670 4483 5684
rect 4143 5656 4158 5668
rect 4177 5656 4190 5670
rect 4258 5666 4411 5670
rect 4140 5654 4162 5656
rect 4240 5654 4432 5666
rect 4511 5654 4524 5684
rect 4539 5670 4569 5684
rect 4606 5654 4625 5684
rect 4640 5654 4646 5684
rect 4655 5654 4668 5684
rect 4683 5670 4713 5684
rect 4756 5670 4799 5684
rect 4806 5670 5026 5684
rect 5033 5670 5063 5684
rect 4723 5656 4738 5668
rect 4757 5656 4770 5670
rect 4838 5666 4991 5670
rect 4720 5654 4742 5656
rect 4820 5654 5012 5666
rect 5091 5654 5104 5684
rect 5119 5670 5149 5684
rect 5186 5654 5205 5684
rect 5220 5654 5226 5684
rect 5235 5654 5248 5684
rect 5263 5670 5293 5684
rect 5336 5670 5379 5684
rect 5386 5670 5606 5684
rect 5613 5670 5643 5684
rect 5303 5656 5318 5668
rect 5337 5656 5350 5670
rect 5418 5666 5571 5670
rect 5300 5654 5322 5656
rect 5400 5654 5592 5666
rect 5671 5654 5684 5684
rect 5699 5670 5729 5684
rect 5766 5654 5785 5684
rect 5800 5654 5806 5684
rect 5815 5654 5828 5684
rect 5843 5670 5873 5684
rect 5916 5670 5959 5684
rect 5966 5670 6186 5684
rect 6193 5670 6223 5684
rect 5883 5656 5898 5668
rect 5917 5656 5930 5670
rect 5998 5666 6151 5670
rect 5880 5654 5902 5656
rect 5980 5654 6172 5666
rect 6251 5654 6264 5684
rect 6279 5670 6309 5684
rect 6346 5654 6365 5684
rect 6380 5654 6386 5684
rect 6395 5654 6408 5684
rect 6423 5670 6453 5684
rect 6496 5670 6539 5684
rect 6546 5670 6766 5684
rect 6773 5670 6803 5684
rect 6463 5656 6478 5668
rect 6497 5656 6510 5670
rect 6578 5666 6731 5670
rect 6460 5654 6482 5656
rect 6560 5654 6752 5666
rect 6831 5654 6844 5684
rect 6859 5670 6889 5684
rect 6926 5654 6945 5684
rect 6960 5654 6966 5684
rect 6975 5654 6988 5684
rect 7003 5670 7033 5684
rect 7076 5670 7119 5684
rect 7126 5670 7346 5684
rect 7353 5670 7383 5684
rect 7043 5656 7058 5668
rect 7077 5656 7090 5670
rect 7158 5666 7311 5670
rect 7040 5654 7062 5656
rect 7140 5654 7332 5666
rect 7411 5654 7424 5684
rect 7439 5670 7469 5684
rect 7506 5654 7525 5684
rect 7540 5654 7546 5684
rect 7555 5654 7568 5684
rect 7583 5666 7613 5684
rect 7656 5670 7670 5684
rect 7706 5670 7926 5684
rect 7657 5668 7670 5670
rect 7623 5656 7638 5668
rect 7620 5654 7642 5656
rect 7647 5654 7677 5668
rect 7738 5666 7891 5670
rect 7720 5654 7912 5666
rect 7955 5654 7985 5668
rect 7991 5654 8004 5684
rect 8019 5666 8049 5684
rect 8092 5654 8105 5684
rect 8135 5654 8148 5684
rect 8163 5666 8193 5684
rect 8236 5670 8250 5684
rect 8286 5670 8506 5684
rect 8237 5668 8250 5670
rect 8203 5656 8218 5668
rect 8200 5654 8222 5656
rect 8227 5654 8257 5668
rect 8318 5666 8471 5670
rect 8300 5654 8492 5666
rect 8535 5654 8565 5668
rect 8571 5654 8584 5684
rect 8599 5666 8629 5684
rect 8672 5654 8685 5684
rect 8715 5654 8728 5684
rect 8743 5666 8773 5684
rect 8816 5670 8830 5684
rect 8866 5670 9086 5684
rect 8817 5668 8830 5670
rect 8783 5656 8798 5668
rect 8780 5654 8802 5656
rect 8807 5654 8837 5668
rect 8898 5666 9051 5670
rect 8880 5654 9072 5666
rect 9115 5654 9145 5668
rect 9151 5654 9164 5684
rect 9179 5666 9209 5684
rect 9252 5654 9265 5684
rect 0 5640 9265 5654
rect 15 5570 28 5640
rect 80 5636 102 5640
rect 73 5614 102 5628
rect 155 5614 171 5628
rect 209 5624 215 5626
rect 222 5624 330 5640
rect 337 5624 343 5626
rect 351 5624 366 5640
rect 432 5634 451 5637
rect 73 5612 171 5614
rect 198 5612 366 5624
rect 381 5614 397 5628
rect 432 5615 454 5634
rect 464 5628 480 5629
rect 463 5626 480 5628
rect 464 5621 480 5626
rect 454 5614 460 5615
rect 463 5614 492 5621
rect 381 5613 492 5614
rect 381 5612 498 5613
rect 57 5604 108 5612
rect 155 5604 189 5612
rect 57 5592 82 5604
rect 89 5592 108 5604
rect 162 5602 189 5604
rect 198 5602 419 5612
rect 454 5609 460 5612
rect 162 5598 419 5602
rect 57 5584 108 5592
rect 155 5584 419 5598
rect 463 5604 498 5612
rect 9 5536 28 5570
rect 73 5576 102 5584
rect 73 5570 90 5576
rect 73 5568 107 5570
rect 155 5568 171 5584
rect 172 5574 380 5584
rect 381 5574 397 5584
rect 445 5580 460 5595
rect 463 5592 464 5604
rect 471 5592 498 5604
rect 463 5584 498 5592
rect 463 5583 492 5584
rect 183 5570 397 5574
rect 198 5568 397 5570
rect 432 5570 445 5580
rect 463 5570 480 5583
rect 432 5568 480 5570
rect 74 5564 107 5568
rect 70 5562 107 5564
rect 70 5561 137 5562
rect 70 5556 101 5561
rect 107 5556 137 5561
rect 70 5552 137 5556
rect 43 5549 137 5552
rect 43 5542 92 5549
rect 43 5536 73 5542
rect 92 5537 97 5542
rect 9 5520 89 5536
rect 101 5528 137 5549
rect 198 5544 387 5568
rect 432 5567 479 5568
rect 445 5562 479 5567
rect 213 5541 387 5544
rect 206 5538 387 5541
rect 415 5561 479 5562
rect 9 5518 28 5520
rect 43 5518 77 5520
rect 9 5502 89 5518
rect 9 5496 28 5502
rect -1 5480 28 5496
rect 43 5486 73 5502
rect 101 5480 107 5528
rect 110 5522 129 5528
rect 144 5522 174 5530
rect 110 5514 174 5522
rect 110 5498 190 5514
rect 206 5507 268 5538
rect 284 5507 346 5538
rect 415 5536 464 5561
rect 479 5536 509 5552
rect 378 5522 408 5530
rect 415 5528 525 5536
rect 378 5514 423 5522
rect 110 5496 129 5498
rect 144 5496 190 5498
rect 110 5480 190 5496
rect 217 5494 252 5507
rect 293 5504 330 5507
rect 293 5502 335 5504
rect 222 5491 252 5494
rect 231 5487 238 5491
rect 238 5486 239 5487
rect 197 5480 207 5486
rect -7 5472 34 5480
rect -7 5446 8 5472
rect 15 5446 34 5472
rect 98 5468 129 5480
rect 144 5468 247 5480
rect 259 5470 285 5496
rect 300 5491 330 5502
rect 362 5498 424 5514
rect 362 5496 408 5498
rect 362 5480 424 5496
rect 436 5480 442 5528
rect 445 5520 525 5528
rect 445 5518 464 5520
rect 479 5518 513 5520
rect 445 5502 525 5518
rect 445 5480 464 5502
rect 479 5486 509 5502
rect 537 5496 543 5570
rect 546 5496 565 5640
rect 580 5496 586 5640
rect 595 5570 608 5640
rect 660 5636 682 5640
rect 653 5614 682 5628
rect 735 5614 751 5628
rect 789 5624 795 5626
rect 802 5624 910 5640
rect 917 5624 923 5626
rect 931 5624 946 5640
rect 1012 5634 1031 5637
rect 653 5612 751 5614
rect 778 5612 946 5624
rect 961 5614 977 5628
rect 1012 5615 1034 5634
rect 1044 5628 1060 5629
rect 1043 5626 1060 5628
rect 1044 5621 1060 5626
rect 1034 5614 1040 5615
rect 1043 5614 1072 5621
rect 961 5613 1072 5614
rect 961 5612 1078 5613
rect 637 5604 688 5612
rect 735 5604 769 5612
rect 637 5592 662 5604
rect 669 5592 688 5604
rect 742 5602 769 5604
rect 778 5602 999 5612
rect 1034 5609 1040 5612
rect 742 5598 999 5602
rect 637 5584 688 5592
rect 735 5584 999 5598
rect 1043 5604 1078 5612
rect 589 5536 608 5570
rect 653 5576 682 5584
rect 653 5570 670 5576
rect 653 5568 687 5570
rect 735 5568 751 5584
rect 752 5574 960 5584
rect 961 5574 977 5584
rect 1025 5580 1040 5595
rect 1043 5592 1044 5604
rect 1051 5592 1078 5604
rect 1043 5584 1078 5592
rect 1043 5583 1072 5584
rect 763 5570 977 5574
rect 778 5568 977 5570
rect 1012 5570 1025 5580
rect 1043 5570 1060 5583
rect 1012 5568 1060 5570
rect 654 5564 687 5568
rect 650 5562 687 5564
rect 650 5561 717 5562
rect 650 5556 681 5561
rect 687 5556 717 5561
rect 650 5552 717 5556
rect 623 5549 717 5552
rect 623 5542 672 5549
rect 623 5536 653 5542
rect 672 5537 677 5542
rect 589 5520 669 5536
rect 681 5528 717 5549
rect 778 5544 967 5568
rect 1012 5567 1059 5568
rect 1025 5562 1059 5567
rect 793 5541 967 5544
rect 786 5538 967 5541
rect 995 5561 1059 5562
rect 589 5518 608 5520
rect 623 5518 657 5520
rect 589 5502 669 5518
rect 589 5496 608 5502
rect 305 5470 408 5480
rect 259 5468 408 5470
rect 429 5468 464 5480
rect 98 5466 260 5468
rect 110 5446 129 5466
rect 144 5464 174 5466
rect -7 5438 34 5446
rect 116 5442 129 5446
rect 181 5450 260 5466
rect 292 5466 464 5468
rect 292 5450 371 5466
rect 378 5464 408 5466
rect -1 5428 28 5438
rect 43 5428 73 5442
rect 116 5428 159 5442
rect 181 5438 371 5450
rect 436 5446 442 5466
rect 166 5428 196 5438
rect 197 5428 355 5438
rect 359 5428 389 5438
rect 393 5428 423 5442
rect 451 5428 464 5466
rect 536 5480 565 5496
rect 579 5480 608 5496
rect 623 5486 653 5502
rect 681 5480 687 5528
rect 690 5522 709 5528
rect 724 5522 754 5530
rect 690 5514 754 5522
rect 690 5498 770 5514
rect 786 5507 848 5538
rect 864 5507 926 5538
rect 995 5536 1044 5561
rect 1059 5536 1089 5552
rect 958 5522 988 5530
rect 995 5528 1105 5536
rect 958 5514 1003 5522
rect 690 5496 709 5498
rect 724 5496 770 5498
rect 690 5480 770 5496
rect 797 5494 832 5507
rect 873 5504 910 5507
rect 873 5502 915 5504
rect 802 5491 832 5494
rect 811 5487 818 5491
rect 818 5486 819 5487
rect 777 5480 787 5486
rect 536 5472 571 5480
rect 536 5446 537 5472
rect 544 5446 571 5472
rect 479 5428 509 5442
rect 536 5438 571 5446
rect 573 5472 614 5480
rect 573 5446 588 5472
rect 595 5446 614 5472
rect 678 5468 709 5480
rect 724 5468 827 5480
rect 839 5470 865 5496
rect 880 5491 910 5502
rect 942 5498 1004 5514
rect 942 5496 988 5498
rect 942 5480 1004 5496
rect 1016 5480 1022 5528
rect 1025 5520 1105 5528
rect 1025 5518 1044 5520
rect 1059 5518 1093 5520
rect 1025 5502 1105 5518
rect 1025 5480 1044 5502
rect 1059 5486 1089 5502
rect 1117 5496 1123 5570
rect 1126 5496 1145 5640
rect 1160 5496 1166 5640
rect 1175 5570 1188 5640
rect 1240 5636 1262 5640
rect 1233 5614 1262 5628
rect 1315 5614 1331 5628
rect 1369 5624 1375 5626
rect 1382 5624 1490 5640
rect 1497 5624 1503 5626
rect 1511 5624 1526 5640
rect 1592 5634 1611 5637
rect 1233 5612 1331 5614
rect 1358 5612 1526 5624
rect 1541 5614 1557 5628
rect 1592 5615 1614 5634
rect 1624 5628 1640 5629
rect 1623 5626 1640 5628
rect 1624 5621 1640 5626
rect 1614 5614 1620 5615
rect 1623 5614 1652 5621
rect 1541 5613 1652 5614
rect 1541 5612 1658 5613
rect 1217 5604 1268 5612
rect 1315 5604 1349 5612
rect 1217 5592 1242 5604
rect 1249 5592 1268 5604
rect 1322 5602 1349 5604
rect 1358 5602 1579 5612
rect 1614 5609 1620 5612
rect 1322 5598 1579 5602
rect 1217 5584 1268 5592
rect 1315 5584 1579 5598
rect 1623 5604 1658 5612
rect 1169 5536 1188 5570
rect 1233 5576 1262 5584
rect 1233 5570 1250 5576
rect 1233 5568 1267 5570
rect 1315 5568 1331 5584
rect 1332 5574 1540 5584
rect 1541 5574 1557 5584
rect 1605 5580 1620 5595
rect 1623 5592 1624 5604
rect 1631 5592 1658 5604
rect 1623 5584 1658 5592
rect 1623 5583 1652 5584
rect 1343 5570 1557 5574
rect 1358 5568 1557 5570
rect 1592 5570 1605 5580
rect 1623 5570 1640 5583
rect 1592 5568 1640 5570
rect 1234 5564 1267 5568
rect 1230 5562 1267 5564
rect 1230 5561 1297 5562
rect 1230 5556 1261 5561
rect 1267 5556 1297 5561
rect 1230 5552 1297 5556
rect 1203 5549 1297 5552
rect 1203 5542 1252 5549
rect 1203 5536 1233 5542
rect 1252 5537 1257 5542
rect 1169 5520 1249 5536
rect 1261 5528 1297 5549
rect 1358 5544 1547 5568
rect 1592 5567 1639 5568
rect 1605 5562 1639 5567
rect 1373 5541 1547 5544
rect 1366 5538 1547 5541
rect 1575 5561 1639 5562
rect 1169 5518 1188 5520
rect 1203 5518 1237 5520
rect 1169 5502 1249 5518
rect 1169 5496 1188 5502
rect 885 5470 988 5480
rect 839 5468 988 5470
rect 1009 5468 1044 5480
rect 678 5466 840 5468
rect 690 5446 709 5466
rect 724 5464 754 5466
rect 573 5438 614 5446
rect 696 5442 709 5446
rect 761 5450 840 5466
rect 872 5466 1044 5468
rect 872 5450 951 5466
rect 958 5464 988 5466
rect 536 5428 565 5438
rect 579 5428 608 5438
rect 623 5428 653 5442
rect 696 5428 739 5442
rect 761 5438 951 5450
rect 1016 5446 1022 5466
rect 746 5428 776 5438
rect 777 5428 935 5438
rect 939 5428 969 5438
rect 973 5428 1003 5442
rect 1031 5428 1044 5466
rect 1116 5480 1145 5496
rect 1159 5480 1188 5496
rect 1203 5486 1233 5502
rect 1261 5480 1267 5528
rect 1270 5522 1289 5528
rect 1304 5522 1334 5530
rect 1270 5514 1334 5522
rect 1270 5498 1350 5514
rect 1366 5507 1428 5538
rect 1444 5507 1506 5538
rect 1575 5536 1624 5561
rect 1639 5536 1669 5552
rect 1538 5522 1568 5530
rect 1575 5528 1685 5536
rect 1538 5514 1583 5522
rect 1270 5496 1289 5498
rect 1304 5496 1350 5498
rect 1270 5480 1350 5496
rect 1377 5494 1412 5507
rect 1453 5504 1490 5507
rect 1453 5502 1495 5504
rect 1382 5491 1412 5494
rect 1391 5487 1398 5491
rect 1398 5486 1399 5487
rect 1357 5480 1367 5486
rect 1116 5472 1151 5480
rect 1116 5446 1117 5472
rect 1124 5446 1151 5472
rect 1059 5428 1089 5442
rect 1116 5438 1151 5446
rect 1153 5472 1194 5480
rect 1153 5446 1168 5472
rect 1175 5446 1194 5472
rect 1258 5468 1289 5480
rect 1304 5468 1407 5480
rect 1419 5470 1445 5496
rect 1460 5491 1490 5502
rect 1522 5498 1584 5514
rect 1522 5496 1568 5498
rect 1522 5480 1584 5496
rect 1596 5480 1602 5528
rect 1605 5520 1685 5528
rect 1605 5518 1624 5520
rect 1639 5518 1673 5520
rect 1605 5502 1685 5518
rect 1605 5480 1624 5502
rect 1639 5486 1669 5502
rect 1697 5496 1703 5570
rect 1706 5496 1725 5640
rect 1740 5496 1746 5640
rect 1755 5570 1768 5640
rect 1820 5636 1842 5640
rect 1813 5614 1842 5628
rect 1895 5614 1911 5628
rect 1949 5624 1955 5626
rect 1962 5624 2070 5640
rect 2077 5624 2083 5626
rect 2091 5624 2106 5640
rect 2172 5634 2191 5637
rect 1813 5612 1911 5614
rect 1938 5612 2106 5624
rect 2121 5614 2137 5628
rect 2172 5615 2194 5634
rect 2204 5628 2220 5629
rect 2203 5626 2220 5628
rect 2204 5621 2220 5626
rect 2194 5614 2200 5615
rect 2203 5614 2232 5621
rect 2121 5613 2232 5614
rect 2121 5612 2238 5613
rect 1797 5604 1848 5612
rect 1895 5604 1929 5612
rect 1797 5592 1822 5604
rect 1829 5592 1848 5604
rect 1902 5602 1929 5604
rect 1938 5602 2159 5612
rect 2194 5609 2200 5612
rect 1902 5598 2159 5602
rect 1797 5584 1848 5592
rect 1895 5584 2159 5598
rect 2203 5604 2238 5612
rect 1749 5536 1768 5570
rect 1813 5576 1842 5584
rect 1813 5570 1830 5576
rect 1813 5568 1847 5570
rect 1895 5568 1911 5584
rect 1912 5574 2120 5584
rect 2121 5574 2137 5584
rect 2185 5580 2200 5595
rect 2203 5592 2204 5604
rect 2211 5592 2238 5604
rect 2203 5584 2238 5592
rect 2203 5583 2232 5584
rect 1923 5570 2137 5574
rect 1938 5568 2137 5570
rect 2172 5570 2185 5580
rect 2203 5570 2220 5583
rect 2172 5568 2220 5570
rect 1814 5564 1847 5568
rect 1810 5562 1847 5564
rect 1810 5561 1877 5562
rect 1810 5556 1841 5561
rect 1847 5556 1877 5561
rect 1810 5552 1877 5556
rect 1783 5549 1877 5552
rect 1783 5542 1832 5549
rect 1783 5536 1813 5542
rect 1832 5537 1837 5542
rect 1749 5520 1829 5536
rect 1841 5528 1877 5549
rect 1938 5544 2127 5568
rect 2172 5567 2219 5568
rect 2185 5562 2219 5567
rect 1953 5541 2127 5544
rect 1946 5538 2127 5541
rect 2155 5561 2219 5562
rect 1749 5518 1768 5520
rect 1783 5518 1817 5520
rect 1749 5502 1829 5518
rect 1749 5496 1768 5502
rect 1465 5470 1568 5480
rect 1419 5468 1568 5470
rect 1589 5468 1624 5480
rect 1258 5466 1420 5468
rect 1270 5446 1289 5466
rect 1304 5464 1334 5466
rect 1153 5438 1194 5446
rect 1276 5442 1289 5446
rect 1341 5450 1420 5466
rect 1452 5466 1624 5468
rect 1452 5450 1531 5466
rect 1538 5464 1568 5466
rect 1116 5428 1145 5438
rect 1159 5428 1188 5438
rect 1203 5428 1233 5442
rect 1276 5428 1319 5442
rect 1341 5438 1531 5450
rect 1596 5446 1602 5466
rect 1326 5428 1356 5438
rect 1357 5428 1515 5438
rect 1519 5428 1549 5438
rect 1553 5428 1583 5442
rect 1611 5428 1624 5466
rect 1696 5480 1725 5496
rect 1739 5480 1768 5496
rect 1783 5486 1813 5502
rect 1841 5480 1847 5528
rect 1850 5522 1869 5528
rect 1884 5522 1914 5530
rect 1850 5514 1914 5522
rect 1850 5498 1930 5514
rect 1946 5507 2008 5538
rect 2024 5507 2086 5538
rect 2155 5536 2204 5561
rect 2219 5536 2249 5552
rect 2118 5522 2148 5530
rect 2155 5528 2265 5536
rect 2118 5514 2163 5522
rect 1850 5496 1869 5498
rect 1884 5496 1930 5498
rect 1850 5480 1930 5496
rect 1957 5494 1992 5507
rect 2033 5504 2070 5507
rect 2033 5502 2075 5504
rect 1962 5491 1992 5494
rect 1971 5487 1978 5491
rect 1978 5486 1979 5487
rect 1937 5480 1947 5486
rect 1696 5472 1731 5480
rect 1696 5446 1697 5472
rect 1704 5446 1731 5472
rect 1639 5428 1669 5442
rect 1696 5438 1731 5446
rect 1733 5472 1774 5480
rect 1733 5446 1748 5472
rect 1755 5446 1774 5472
rect 1838 5468 1869 5480
rect 1884 5468 1987 5480
rect 1999 5470 2025 5496
rect 2040 5491 2070 5502
rect 2102 5498 2164 5514
rect 2102 5496 2148 5498
rect 2102 5480 2164 5496
rect 2176 5480 2182 5528
rect 2185 5520 2265 5528
rect 2185 5518 2204 5520
rect 2219 5518 2253 5520
rect 2185 5502 2265 5518
rect 2185 5480 2204 5502
rect 2219 5486 2249 5502
rect 2277 5496 2283 5570
rect 2286 5496 2305 5640
rect 2320 5496 2326 5640
rect 2335 5570 2348 5640
rect 2400 5636 2422 5640
rect 2393 5614 2422 5628
rect 2475 5614 2491 5628
rect 2529 5624 2535 5626
rect 2542 5624 2650 5640
rect 2657 5624 2663 5626
rect 2671 5624 2686 5640
rect 2752 5634 2771 5637
rect 2393 5612 2491 5614
rect 2518 5612 2686 5624
rect 2701 5614 2717 5628
rect 2752 5615 2774 5634
rect 2784 5628 2800 5629
rect 2783 5626 2800 5628
rect 2784 5621 2800 5626
rect 2774 5614 2780 5615
rect 2783 5614 2812 5621
rect 2701 5613 2812 5614
rect 2701 5612 2818 5613
rect 2377 5604 2428 5612
rect 2475 5604 2509 5612
rect 2377 5592 2402 5604
rect 2409 5592 2428 5604
rect 2482 5602 2509 5604
rect 2518 5602 2739 5612
rect 2774 5609 2780 5612
rect 2482 5598 2739 5602
rect 2377 5584 2428 5592
rect 2475 5584 2739 5598
rect 2783 5604 2818 5612
rect 2329 5536 2348 5570
rect 2393 5576 2422 5584
rect 2393 5570 2410 5576
rect 2393 5568 2427 5570
rect 2475 5568 2491 5584
rect 2492 5574 2700 5584
rect 2701 5574 2717 5584
rect 2765 5580 2780 5595
rect 2783 5592 2784 5604
rect 2791 5592 2818 5604
rect 2783 5584 2818 5592
rect 2783 5583 2812 5584
rect 2503 5570 2717 5574
rect 2518 5568 2717 5570
rect 2752 5570 2765 5580
rect 2783 5570 2800 5583
rect 2752 5568 2800 5570
rect 2394 5564 2427 5568
rect 2390 5562 2427 5564
rect 2390 5561 2457 5562
rect 2390 5556 2421 5561
rect 2427 5556 2457 5561
rect 2390 5552 2457 5556
rect 2363 5549 2457 5552
rect 2363 5542 2412 5549
rect 2363 5536 2393 5542
rect 2412 5537 2417 5542
rect 2329 5520 2409 5536
rect 2421 5528 2457 5549
rect 2518 5544 2707 5568
rect 2752 5567 2799 5568
rect 2765 5562 2799 5567
rect 2533 5541 2707 5544
rect 2526 5538 2707 5541
rect 2735 5561 2799 5562
rect 2329 5518 2348 5520
rect 2363 5518 2397 5520
rect 2329 5502 2409 5518
rect 2329 5496 2348 5502
rect 2045 5470 2148 5480
rect 1999 5468 2148 5470
rect 2169 5468 2204 5480
rect 1838 5466 2000 5468
rect 1850 5446 1869 5466
rect 1884 5464 1914 5466
rect 1733 5438 1774 5446
rect 1856 5442 1869 5446
rect 1921 5450 2000 5466
rect 2032 5466 2204 5468
rect 2032 5450 2111 5466
rect 2118 5464 2148 5466
rect 1696 5428 1725 5438
rect 1739 5428 1768 5438
rect 1783 5428 1813 5442
rect 1856 5428 1899 5442
rect 1921 5438 2111 5450
rect 2176 5446 2182 5466
rect 1906 5428 1936 5438
rect 1937 5428 2095 5438
rect 2099 5428 2129 5438
rect 2133 5428 2163 5442
rect 2191 5428 2204 5466
rect 2276 5480 2305 5496
rect 2319 5480 2348 5496
rect 2363 5486 2393 5502
rect 2421 5480 2427 5528
rect 2430 5522 2449 5528
rect 2464 5522 2494 5530
rect 2430 5514 2494 5522
rect 2430 5498 2510 5514
rect 2526 5507 2588 5538
rect 2604 5507 2666 5538
rect 2735 5536 2784 5561
rect 2799 5536 2829 5552
rect 2698 5522 2728 5530
rect 2735 5528 2845 5536
rect 2698 5514 2743 5522
rect 2430 5496 2449 5498
rect 2464 5496 2510 5498
rect 2430 5480 2510 5496
rect 2537 5494 2572 5507
rect 2613 5504 2650 5507
rect 2613 5502 2655 5504
rect 2542 5491 2572 5494
rect 2551 5487 2558 5491
rect 2558 5486 2559 5487
rect 2517 5480 2527 5486
rect 2276 5472 2311 5480
rect 2276 5446 2277 5472
rect 2284 5446 2311 5472
rect 2219 5428 2249 5442
rect 2276 5438 2311 5446
rect 2313 5472 2354 5480
rect 2313 5446 2328 5472
rect 2335 5446 2354 5472
rect 2418 5468 2449 5480
rect 2464 5468 2567 5480
rect 2579 5470 2605 5496
rect 2620 5491 2650 5502
rect 2682 5498 2744 5514
rect 2682 5496 2728 5498
rect 2682 5480 2744 5496
rect 2756 5480 2762 5528
rect 2765 5520 2845 5528
rect 2765 5518 2784 5520
rect 2799 5518 2833 5520
rect 2765 5502 2845 5518
rect 2765 5480 2784 5502
rect 2799 5486 2829 5502
rect 2857 5496 2863 5570
rect 2866 5496 2885 5640
rect 2900 5496 2906 5640
rect 2915 5570 2928 5640
rect 2980 5636 3002 5640
rect 2973 5614 3002 5628
rect 3055 5614 3071 5628
rect 3109 5624 3115 5626
rect 3122 5624 3230 5640
rect 3237 5624 3243 5626
rect 3251 5624 3266 5640
rect 3332 5634 3351 5637
rect 2973 5612 3071 5614
rect 3098 5612 3266 5624
rect 3281 5614 3297 5628
rect 3332 5615 3354 5634
rect 3364 5628 3380 5629
rect 3363 5626 3380 5628
rect 3364 5621 3380 5626
rect 3354 5614 3360 5615
rect 3363 5614 3392 5621
rect 3281 5613 3392 5614
rect 3281 5612 3398 5613
rect 2957 5604 3008 5612
rect 3055 5604 3089 5612
rect 2957 5592 2982 5604
rect 2989 5592 3008 5604
rect 3062 5602 3089 5604
rect 3098 5602 3319 5612
rect 3354 5609 3360 5612
rect 3062 5598 3319 5602
rect 2957 5584 3008 5592
rect 3055 5584 3319 5598
rect 3363 5604 3398 5612
rect 2909 5536 2928 5570
rect 2973 5576 3002 5584
rect 2973 5570 2990 5576
rect 2973 5568 3007 5570
rect 3055 5568 3071 5584
rect 3072 5574 3280 5584
rect 3281 5574 3297 5584
rect 3345 5580 3360 5595
rect 3363 5592 3364 5604
rect 3371 5592 3398 5604
rect 3363 5584 3398 5592
rect 3363 5583 3392 5584
rect 3083 5570 3297 5574
rect 3098 5568 3297 5570
rect 3332 5570 3345 5580
rect 3363 5570 3380 5583
rect 3332 5568 3380 5570
rect 2974 5564 3007 5568
rect 2970 5562 3007 5564
rect 2970 5561 3037 5562
rect 2970 5556 3001 5561
rect 3007 5556 3037 5561
rect 2970 5552 3037 5556
rect 2943 5549 3037 5552
rect 2943 5542 2992 5549
rect 2943 5536 2973 5542
rect 2992 5537 2997 5542
rect 2909 5520 2989 5536
rect 3001 5528 3037 5549
rect 3098 5544 3287 5568
rect 3332 5567 3379 5568
rect 3345 5562 3379 5567
rect 3113 5541 3287 5544
rect 3106 5538 3287 5541
rect 3315 5561 3379 5562
rect 2909 5518 2928 5520
rect 2943 5518 2977 5520
rect 2909 5502 2989 5518
rect 2909 5496 2928 5502
rect 2625 5470 2728 5480
rect 2579 5468 2728 5470
rect 2749 5468 2784 5480
rect 2418 5466 2580 5468
rect 2430 5446 2449 5466
rect 2464 5464 2494 5466
rect 2313 5438 2354 5446
rect 2436 5442 2449 5446
rect 2501 5450 2580 5466
rect 2612 5466 2784 5468
rect 2612 5450 2691 5466
rect 2698 5464 2728 5466
rect 2276 5428 2305 5438
rect 2319 5428 2348 5438
rect 2363 5428 2393 5442
rect 2436 5428 2479 5442
rect 2501 5438 2691 5450
rect 2756 5446 2762 5466
rect 2486 5428 2516 5438
rect 2517 5428 2675 5438
rect 2679 5428 2709 5438
rect 2713 5428 2743 5442
rect 2771 5428 2784 5466
rect 2856 5480 2885 5496
rect 2899 5480 2928 5496
rect 2943 5486 2973 5502
rect 3001 5480 3007 5528
rect 3010 5522 3029 5528
rect 3044 5522 3074 5530
rect 3010 5514 3074 5522
rect 3010 5498 3090 5514
rect 3106 5507 3168 5538
rect 3184 5507 3246 5538
rect 3315 5536 3364 5561
rect 3379 5536 3409 5552
rect 3278 5522 3308 5530
rect 3315 5528 3425 5536
rect 3278 5514 3323 5522
rect 3010 5496 3029 5498
rect 3044 5496 3090 5498
rect 3010 5480 3090 5496
rect 3117 5494 3152 5507
rect 3193 5504 3230 5507
rect 3193 5502 3235 5504
rect 3122 5491 3152 5494
rect 3131 5487 3138 5491
rect 3138 5486 3139 5487
rect 3097 5480 3107 5486
rect 2856 5472 2891 5480
rect 2856 5446 2857 5472
rect 2864 5446 2891 5472
rect 2799 5428 2829 5442
rect 2856 5438 2891 5446
rect 2893 5472 2934 5480
rect 2893 5446 2908 5472
rect 2915 5446 2934 5472
rect 2998 5468 3029 5480
rect 3044 5468 3147 5480
rect 3159 5470 3185 5496
rect 3200 5491 3230 5502
rect 3262 5498 3324 5514
rect 3262 5496 3308 5498
rect 3262 5480 3324 5496
rect 3336 5480 3342 5528
rect 3345 5520 3425 5528
rect 3345 5518 3364 5520
rect 3379 5518 3413 5520
rect 3345 5502 3425 5518
rect 3345 5480 3364 5502
rect 3379 5486 3409 5502
rect 3437 5496 3443 5570
rect 3446 5496 3465 5640
rect 3480 5496 3486 5640
rect 3495 5570 3508 5640
rect 3560 5636 3582 5640
rect 3553 5614 3582 5628
rect 3635 5614 3651 5628
rect 3689 5624 3695 5626
rect 3702 5624 3810 5640
rect 3817 5624 3823 5626
rect 3831 5624 3846 5640
rect 3912 5634 3931 5637
rect 3553 5612 3651 5614
rect 3678 5612 3846 5624
rect 3861 5614 3877 5628
rect 3912 5615 3934 5634
rect 3944 5628 3960 5629
rect 3943 5626 3960 5628
rect 3944 5621 3960 5626
rect 3934 5614 3940 5615
rect 3943 5614 3972 5621
rect 3861 5613 3972 5614
rect 3861 5612 3978 5613
rect 3537 5604 3588 5612
rect 3635 5604 3669 5612
rect 3537 5592 3562 5604
rect 3569 5592 3588 5604
rect 3642 5602 3669 5604
rect 3678 5602 3899 5612
rect 3934 5609 3940 5612
rect 3642 5598 3899 5602
rect 3537 5584 3588 5592
rect 3635 5584 3899 5598
rect 3943 5604 3978 5612
rect 3489 5536 3508 5570
rect 3553 5576 3582 5584
rect 3553 5570 3570 5576
rect 3553 5568 3587 5570
rect 3635 5568 3651 5584
rect 3652 5574 3860 5584
rect 3861 5574 3877 5584
rect 3925 5580 3940 5595
rect 3943 5592 3944 5604
rect 3951 5592 3978 5604
rect 3943 5584 3978 5592
rect 3943 5583 3972 5584
rect 3663 5570 3877 5574
rect 3678 5568 3877 5570
rect 3912 5570 3925 5580
rect 3943 5570 3960 5583
rect 3912 5568 3960 5570
rect 3554 5564 3587 5568
rect 3550 5562 3587 5564
rect 3550 5561 3617 5562
rect 3550 5556 3581 5561
rect 3587 5556 3617 5561
rect 3550 5552 3617 5556
rect 3523 5549 3617 5552
rect 3523 5542 3572 5549
rect 3523 5536 3553 5542
rect 3572 5537 3577 5542
rect 3489 5520 3569 5536
rect 3581 5528 3617 5549
rect 3678 5544 3867 5568
rect 3912 5567 3959 5568
rect 3925 5562 3959 5567
rect 3693 5541 3867 5544
rect 3686 5538 3867 5541
rect 3895 5561 3959 5562
rect 3489 5518 3508 5520
rect 3523 5518 3557 5520
rect 3489 5502 3569 5518
rect 3489 5496 3508 5502
rect 3205 5470 3308 5480
rect 3159 5468 3308 5470
rect 3329 5468 3364 5480
rect 2998 5466 3160 5468
rect 3010 5446 3029 5466
rect 3044 5464 3074 5466
rect 2893 5438 2934 5446
rect 3016 5442 3029 5446
rect 3081 5450 3160 5466
rect 3192 5466 3364 5468
rect 3192 5450 3271 5466
rect 3278 5464 3308 5466
rect 2856 5428 2885 5438
rect 2899 5428 2928 5438
rect 2943 5428 2973 5442
rect 3016 5428 3059 5442
rect 3081 5438 3271 5450
rect 3336 5446 3342 5466
rect 3066 5428 3096 5438
rect 3097 5428 3255 5438
rect 3259 5428 3289 5438
rect 3293 5428 3323 5442
rect 3351 5428 3364 5466
rect 3436 5480 3465 5496
rect 3479 5480 3508 5496
rect 3523 5486 3553 5502
rect 3581 5480 3587 5528
rect 3590 5522 3609 5528
rect 3624 5522 3654 5530
rect 3590 5514 3654 5522
rect 3590 5498 3670 5514
rect 3686 5507 3748 5538
rect 3764 5507 3826 5538
rect 3895 5536 3944 5561
rect 3959 5536 3989 5552
rect 3858 5522 3888 5530
rect 3895 5528 4005 5536
rect 3858 5514 3903 5522
rect 3590 5496 3609 5498
rect 3624 5496 3670 5498
rect 3590 5480 3670 5496
rect 3697 5494 3732 5507
rect 3773 5504 3810 5507
rect 3773 5502 3815 5504
rect 3702 5491 3732 5494
rect 3711 5487 3718 5491
rect 3718 5486 3719 5487
rect 3677 5480 3687 5486
rect 3436 5472 3471 5480
rect 3436 5446 3437 5472
rect 3444 5446 3471 5472
rect 3379 5428 3409 5442
rect 3436 5438 3471 5446
rect 3473 5472 3514 5480
rect 3473 5446 3488 5472
rect 3495 5446 3514 5472
rect 3578 5468 3609 5480
rect 3624 5468 3727 5480
rect 3739 5470 3765 5496
rect 3780 5491 3810 5502
rect 3842 5498 3904 5514
rect 3842 5496 3888 5498
rect 3842 5480 3904 5496
rect 3916 5480 3922 5528
rect 3925 5520 4005 5528
rect 3925 5518 3944 5520
rect 3959 5518 3993 5520
rect 3925 5502 4005 5518
rect 3925 5480 3944 5502
rect 3959 5486 3989 5502
rect 4017 5496 4023 5570
rect 4026 5496 4045 5640
rect 4060 5496 4066 5640
rect 4075 5570 4088 5640
rect 4140 5636 4162 5640
rect 4133 5614 4162 5628
rect 4215 5614 4231 5628
rect 4269 5624 4275 5626
rect 4282 5624 4390 5640
rect 4397 5624 4403 5626
rect 4411 5624 4426 5640
rect 4492 5634 4511 5637
rect 4133 5612 4231 5614
rect 4258 5612 4426 5624
rect 4441 5614 4457 5628
rect 4492 5615 4514 5634
rect 4524 5628 4540 5629
rect 4523 5626 4540 5628
rect 4524 5621 4540 5626
rect 4514 5614 4520 5615
rect 4523 5614 4552 5621
rect 4441 5613 4552 5614
rect 4441 5612 4558 5613
rect 4117 5604 4168 5612
rect 4215 5604 4249 5612
rect 4117 5592 4142 5604
rect 4149 5592 4168 5604
rect 4222 5602 4249 5604
rect 4258 5602 4479 5612
rect 4514 5609 4520 5612
rect 4222 5598 4479 5602
rect 4117 5584 4168 5592
rect 4215 5584 4479 5598
rect 4523 5604 4558 5612
rect 4069 5536 4088 5570
rect 4133 5576 4162 5584
rect 4133 5570 4150 5576
rect 4133 5568 4167 5570
rect 4215 5568 4231 5584
rect 4232 5574 4440 5584
rect 4441 5574 4457 5584
rect 4505 5580 4520 5595
rect 4523 5592 4524 5604
rect 4531 5592 4558 5604
rect 4523 5584 4558 5592
rect 4523 5583 4552 5584
rect 4243 5570 4457 5574
rect 4258 5568 4457 5570
rect 4492 5570 4505 5580
rect 4523 5570 4540 5583
rect 4492 5568 4540 5570
rect 4134 5564 4167 5568
rect 4130 5562 4167 5564
rect 4130 5561 4197 5562
rect 4130 5556 4161 5561
rect 4167 5556 4197 5561
rect 4130 5552 4197 5556
rect 4103 5549 4197 5552
rect 4103 5542 4152 5549
rect 4103 5536 4133 5542
rect 4152 5537 4157 5542
rect 4069 5520 4149 5536
rect 4161 5528 4197 5549
rect 4258 5544 4447 5568
rect 4492 5567 4539 5568
rect 4505 5562 4539 5567
rect 4273 5541 4447 5544
rect 4266 5538 4447 5541
rect 4475 5561 4539 5562
rect 4069 5518 4088 5520
rect 4103 5518 4137 5520
rect 4069 5502 4149 5518
rect 4069 5496 4088 5502
rect 3785 5470 3888 5480
rect 3739 5468 3888 5470
rect 3909 5468 3944 5480
rect 3578 5466 3740 5468
rect 3590 5446 3609 5466
rect 3624 5464 3654 5466
rect 3473 5438 3514 5446
rect 3596 5442 3609 5446
rect 3661 5450 3740 5466
rect 3772 5466 3944 5468
rect 3772 5450 3851 5466
rect 3858 5464 3888 5466
rect 3436 5428 3465 5438
rect 3479 5428 3508 5438
rect 3523 5428 3553 5442
rect 3596 5428 3639 5442
rect 3661 5438 3851 5450
rect 3916 5446 3922 5466
rect 3646 5428 3676 5438
rect 3677 5428 3835 5438
rect 3839 5428 3869 5438
rect 3873 5428 3903 5442
rect 3931 5428 3944 5466
rect 4016 5480 4045 5496
rect 4059 5480 4088 5496
rect 4103 5486 4133 5502
rect 4161 5480 4167 5528
rect 4170 5522 4189 5528
rect 4204 5522 4234 5530
rect 4170 5514 4234 5522
rect 4170 5498 4250 5514
rect 4266 5507 4328 5538
rect 4344 5507 4406 5538
rect 4475 5536 4524 5561
rect 4539 5536 4569 5552
rect 4438 5522 4468 5530
rect 4475 5528 4585 5536
rect 4438 5514 4483 5522
rect 4170 5496 4189 5498
rect 4204 5496 4250 5498
rect 4170 5480 4250 5496
rect 4277 5494 4312 5507
rect 4353 5504 4390 5507
rect 4353 5502 4395 5504
rect 4282 5491 4312 5494
rect 4291 5487 4298 5491
rect 4298 5486 4299 5487
rect 4257 5480 4267 5486
rect 4016 5472 4051 5480
rect 4016 5446 4017 5472
rect 4024 5446 4051 5472
rect 3959 5428 3989 5442
rect 4016 5438 4051 5446
rect 4053 5472 4094 5480
rect 4053 5446 4068 5472
rect 4075 5446 4094 5472
rect 4158 5468 4189 5480
rect 4204 5468 4307 5480
rect 4319 5470 4345 5496
rect 4360 5491 4390 5502
rect 4422 5498 4484 5514
rect 4422 5496 4468 5498
rect 4422 5480 4484 5496
rect 4496 5480 4502 5528
rect 4505 5520 4585 5528
rect 4505 5518 4524 5520
rect 4539 5518 4573 5520
rect 4505 5502 4585 5518
rect 4505 5480 4524 5502
rect 4539 5486 4569 5502
rect 4597 5496 4603 5570
rect 4606 5496 4625 5640
rect 4640 5496 4646 5640
rect 4655 5570 4668 5640
rect 4720 5636 4742 5640
rect 4713 5614 4742 5628
rect 4795 5614 4811 5628
rect 4849 5624 4855 5626
rect 4862 5624 4970 5640
rect 4977 5624 4983 5626
rect 4991 5624 5006 5640
rect 5072 5634 5091 5637
rect 4713 5612 4811 5614
rect 4838 5612 5006 5624
rect 5021 5614 5037 5628
rect 5072 5615 5094 5634
rect 5104 5628 5120 5629
rect 5103 5626 5120 5628
rect 5104 5621 5120 5626
rect 5094 5614 5100 5615
rect 5103 5614 5132 5621
rect 5021 5613 5132 5614
rect 5021 5612 5138 5613
rect 4697 5604 4748 5612
rect 4795 5604 4829 5612
rect 4697 5592 4722 5604
rect 4729 5592 4748 5604
rect 4802 5602 4829 5604
rect 4838 5602 5059 5612
rect 5094 5609 5100 5612
rect 4802 5598 5059 5602
rect 4697 5584 4748 5592
rect 4795 5584 5059 5598
rect 5103 5604 5138 5612
rect 4649 5536 4668 5570
rect 4713 5576 4742 5584
rect 4713 5570 4730 5576
rect 4713 5568 4747 5570
rect 4795 5568 4811 5584
rect 4812 5574 5020 5584
rect 5021 5574 5037 5584
rect 5085 5580 5100 5595
rect 5103 5592 5104 5604
rect 5111 5592 5138 5604
rect 5103 5584 5138 5592
rect 5103 5583 5132 5584
rect 4823 5570 5037 5574
rect 4838 5568 5037 5570
rect 5072 5570 5085 5580
rect 5103 5570 5120 5583
rect 5072 5568 5120 5570
rect 4714 5564 4747 5568
rect 4710 5562 4747 5564
rect 4710 5561 4777 5562
rect 4710 5556 4741 5561
rect 4747 5556 4777 5561
rect 4710 5552 4777 5556
rect 4683 5549 4777 5552
rect 4683 5542 4732 5549
rect 4683 5536 4713 5542
rect 4732 5537 4737 5542
rect 4649 5520 4729 5536
rect 4741 5528 4777 5549
rect 4838 5544 5027 5568
rect 5072 5567 5119 5568
rect 5085 5562 5119 5567
rect 4853 5541 5027 5544
rect 4846 5538 5027 5541
rect 5055 5561 5119 5562
rect 4649 5518 4668 5520
rect 4683 5518 4717 5520
rect 4649 5502 4729 5518
rect 4649 5496 4668 5502
rect 4365 5470 4468 5480
rect 4319 5468 4468 5470
rect 4489 5468 4524 5480
rect 4158 5466 4320 5468
rect 4170 5446 4189 5466
rect 4204 5464 4234 5466
rect 4053 5438 4094 5446
rect 4176 5442 4189 5446
rect 4241 5450 4320 5466
rect 4352 5466 4524 5468
rect 4352 5450 4431 5466
rect 4438 5464 4468 5466
rect 4016 5428 4045 5438
rect 4059 5428 4088 5438
rect 4103 5428 4133 5442
rect 4176 5428 4219 5442
rect 4241 5438 4431 5450
rect 4496 5446 4502 5466
rect 4226 5428 4256 5438
rect 4257 5428 4415 5438
rect 4419 5428 4449 5438
rect 4453 5428 4483 5442
rect 4511 5428 4524 5466
rect 4596 5480 4625 5496
rect 4639 5480 4668 5496
rect 4683 5486 4713 5502
rect 4741 5480 4747 5528
rect 4750 5522 4769 5528
rect 4784 5522 4814 5530
rect 4750 5514 4814 5522
rect 4750 5498 4830 5514
rect 4846 5507 4908 5538
rect 4924 5507 4986 5538
rect 5055 5536 5104 5561
rect 5119 5536 5149 5552
rect 5018 5522 5048 5530
rect 5055 5528 5165 5536
rect 5018 5514 5063 5522
rect 4750 5496 4769 5498
rect 4784 5496 4830 5498
rect 4750 5480 4830 5496
rect 4857 5494 4892 5507
rect 4933 5504 4970 5507
rect 4933 5502 4975 5504
rect 4862 5491 4892 5494
rect 4871 5487 4878 5491
rect 4878 5486 4879 5487
rect 4837 5480 4847 5486
rect 4596 5472 4631 5480
rect 4596 5446 4597 5472
rect 4604 5446 4631 5472
rect 4539 5428 4569 5442
rect 4596 5438 4631 5446
rect 4633 5472 4674 5480
rect 4633 5446 4648 5472
rect 4655 5446 4674 5472
rect 4738 5468 4769 5480
rect 4784 5468 4887 5480
rect 4899 5470 4925 5496
rect 4940 5491 4970 5502
rect 5002 5498 5064 5514
rect 5002 5496 5048 5498
rect 5002 5480 5064 5496
rect 5076 5480 5082 5528
rect 5085 5520 5165 5528
rect 5085 5518 5104 5520
rect 5119 5518 5153 5520
rect 5085 5502 5165 5518
rect 5085 5480 5104 5502
rect 5119 5486 5149 5502
rect 5177 5496 5183 5570
rect 5186 5496 5205 5640
rect 5220 5496 5226 5640
rect 5235 5570 5248 5640
rect 5300 5636 5322 5640
rect 5293 5614 5322 5628
rect 5375 5614 5391 5628
rect 5429 5624 5435 5626
rect 5442 5624 5550 5640
rect 5557 5624 5563 5626
rect 5571 5624 5586 5640
rect 5652 5634 5671 5637
rect 5293 5612 5391 5614
rect 5418 5612 5586 5624
rect 5601 5614 5617 5628
rect 5652 5615 5674 5634
rect 5684 5628 5700 5629
rect 5683 5626 5700 5628
rect 5684 5621 5700 5626
rect 5674 5614 5680 5615
rect 5683 5614 5712 5621
rect 5601 5613 5712 5614
rect 5601 5612 5718 5613
rect 5277 5604 5328 5612
rect 5375 5604 5409 5612
rect 5277 5592 5302 5604
rect 5309 5592 5328 5604
rect 5382 5602 5409 5604
rect 5418 5602 5639 5612
rect 5674 5609 5680 5612
rect 5382 5598 5639 5602
rect 5277 5584 5328 5592
rect 5375 5584 5639 5598
rect 5683 5604 5718 5612
rect 5229 5536 5248 5570
rect 5293 5576 5322 5584
rect 5293 5570 5310 5576
rect 5293 5568 5327 5570
rect 5375 5568 5391 5584
rect 5392 5574 5600 5584
rect 5601 5574 5617 5584
rect 5665 5580 5680 5595
rect 5683 5592 5684 5604
rect 5691 5592 5718 5604
rect 5683 5584 5718 5592
rect 5683 5583 5712 5584
rect 5403 5570 5617 5574
rect 5418 5568 5617 5570
rect 5652 5570 5665 5580
rect 5683 5570 5700 5583
rect 5652 5568 5700 5570
rect 5294 5564 5327 5568
rect 5290 5562 5327 5564
rect 5290 5561 5357 5562
rect 5290 5556 5321 5561
rect 5327 5556 5357 5561
rect 5290 5552 5357 5556
rect 5263 5549 5357 5552
rect 5263 5542 5312 5549
rect 5263 5536 5293 5542
rect 5312 5537 5317 5542
rect 5229 5520 5309 5536
rect 5321 5528 5357 5549
rect 5418 5544 5607 5568
rect 5652 5567 5699 5568
rect 5665 5562 5699 5567
rect 5433 5541 5607 5544
rect 5426 5538 5607 5541
rect 5635 5561 5699 5562
rect 5229 5518 5248 5520
rect 5263 5518 5297 5520
rect 5229 5502 5309 5518
rect 5229 5496 5248 5502
rect 4945 5470 5048 5480
rect 4899 5468 5048 5470
rect 5069 5468 5104 5480
rect 4738 5466 4900 5468
rect 4750 5446 4769 5466
rect 4784 5464 4814 5466
rect 4633 5438 4674 5446
rect 4756 5442 4769 5446
rect 4821 5450 4900 5466
rect 4932 5466 5104 5468
rect 4932 5450 5011 5466
rect 5018 5464 5048 5466
rect 4596 5428 4625 5438
rect 4639 5428 4668 5438
rect 4683 5428 4713 5442
rect 4756 5428 4799 5442
rect 4821 5438 5011 5450
rect 5076 5446 5082 5466
rect 4806 5428 4836 5438
rect 4837 5428 4995 5438
rect 4999 5428 5029 5438
rect 5033 5428 5063 5442
rect 5091 5428 5104 5466
rect 5176 5480 5205 5496
rect 5219 5480 5248 5496
rect 5263 5486 5293 5502
rect 5321 5480 5327 5528
rect 5330 5522 5349 5528
rect 5364 5522 5394 5530
rect 5330 5514 5394 5522
rect 5330 5498 5410 5514
rect 5426 5507 5488 5538
rect 5504 5507 5566 5538
rect 5635 5536 5684 5561
rect 5699 5536 5729 5552
rect 5598 5522 5628 5530
rect 5635 5528 5745 5536
rect 5598 5514 5643 5522
rect 5330 5496 5349 5498
rect 5364 5496 5410 5498
rect 5330 5480 5410 5496
rect 5437 5494 5472 5507
rect 5513 5504 5550 5507
rect 5513 5502 5555 5504
rect 5442 5491 5472 5494
rect 5451 5487 5458 5491
rect 5458 5486 5459 5487
rect 5417 5480 5427 5486
rect 5176 5472 5211 5480
rect 5176 5446 5177 5472
rect 5184 5446 5211 5472
rect 5119 5428 5149 5442
rect 5176 5438 5211 5446
rect 5213 5472 5254 5480
rect 5213 5446 5228 5472
rect 5235 5446 5254 5472
rect 5318 5468 5349 5480
rect 5364 5468 5467 5480
rect 5479 5470 5505 5496
rect 5520 5491 5550 5502
rect 5582 5498 5644 5514
rect 5582 5496 5628 5498
rect 5582 5480 5644 5496
rect 5656 5480 5662 5528
rect 5665 5520 5745 5528
rect 5665 5518 5684 5520
rect 5699 5518 5733 5520
rect 5665 5502 5745 5518
rect 5665 5480 5684 5502
rect 5699 5486 5729 5502
rect 5757 5496 5763 5570
rect 5766 5496 5785 5640
rect 5800 5496 5806 5640
rect 5815 5570 5828 5640
rect 5880 5636 5902 5640
rect 5873 5614 5902 5628
rect 5955 5614 5971 5628
rect 6009 5624 6015 5626
rect 6022 5624 6130 5640
rect 6137 5624 6143 5626
rect 6151 5624 6166 5640
rect 6232 5634 6251 5637
rect 5873 5612 5971 5614
rect 5998 5612 6166 5624
rect 6181 5614 6197 5628
rect 6232 5615 6254 5634
rect 6264 5628 6280 5629
rect 6263 5626 6280 5628
rect 6264 5621 6280 5626
rect 6254 5614 6260 5615
rect 6263 5614 6292 5621
rect 6181 5613 6292 5614
rect 6181 5612 6298 5613
rect 5857 5604 5908 5612
rect 5955 5604 5989 5612
rect 5857 5592 5882 5604
rect 5889 5592 5908 5604
rect 5962 5602 5989 5604
rect 5998 5602 6219 5612
rect 6254 5609 6260 5612
rect 5962 5598 6219 5602
rect 5857 5584 5908 5592
rect 5955 5584 6219 5598
rect 6263 5604 6298 5612
rect 5809 5536 5828 5570
rect 5873 5576 5902 5584
rect 5873 5570 5890 5576
rect 5873 5568 5907 5570
rect 5955 5568 5971 5584
rect 5972 5574 6180 5584
rect 6181 5574 6197 5584
rect 6245 5580 6260 5595
rect 6263 5592 6264 5604
rect 6271 5592 6298 5604
rect 6263 5584 6298 5592
rect 6263 5583 6292 5584
rect 5983 5570 6197 5574
rect 5998 5568 6197 5570
rect 6232 5570 6245 5580
rect 6263 5570 6280 5583
rect 6232 5568 6280 5570
rect 5874 5564 5907 5568
rect 5870 5562 5907 5564
rect 5870 5561 5937 5562
rect 5870 5556 5901 5561
rect 5907 5556 5937 5561
rect 5870 5552 5937 5556
rect 5843 5549 5937 5552
rect 5843 5542 5892 5549
rect 5843 5536 5873 5542
rect 5892 5537 5897 5542
rect 5809 5520 5889 5536
rect 5901 5528 5937 5549
rect 5998 5544 6187 5568
rect 6232 5567 6279 5568
rect 6245 5562 6279 5567
rect 6013 5541 6187 5544
rect 6006 5538 6187 5541
rect 6215 5561 6279 5562
rect 5809 5518 5828 5520
rect 5843 5518 5877 5520
rect 5809 5502 5889 5518
rect 5809 5496 5828 5502
rect 5525 5470 5628 5480
rect 5479 5468 5628 5470
rect 5649 5468 5684 5480
rect 5318 5466 5480 5468
rect 5330 5446 5349 5466
rect 5364 5464 5394 5466
rect 5213 5438 5254 5446
rect 5336 5442 5349 5446
rect 5401 5450 5480 5466
rect 5512 5466 5684 5468
rect 5512 5450 5591 5466
rect 5598 5464 5628 5466
rect 5176 5428 5205 5438
rect 5219 5428 5248 5438
rect 5263 5428 5293 5442
rect 5336 5428 5379 5442
rect 5401 5438 5591 5450
rect 5656 5446 5662 5466
rect 5386 5428 5416 5438
rect 5417 5428 5575 5438
rect 5579 5428 5609 5438
rect 5613 5428 5643 5442
rect 5671 5428 5684 5466
rect 5756 5480 5785 5496
rect 5799 5480 5828 5496
rect 5843 5486 5873 5502
rect 5901 5480 5907 5528
rect 5910 5522 5929 5528
rect 5944 5522 5974 5530
rect 5910 5514 5974 5522
rect 5910 5498 5990 5514
rect 6006 5507 6068 5538
rect 6084 5507 6146 5538
rect 6215 5536 6264 5561
rect 6279 5536 6309 5552
rect 6178 5522 6208 5530
rect 6215 5528 6325 5536
rect 6178 5514 6223 5522
rect 5910 5496 5929 5498
rect 5944 5496 5990 5498
rect 5910 5480 5990 5496
rect 6017 5494 6052 5507
rect 6093 5504 6130 5507
rect 6093 5502 6135 5504
rect 6022 5491 6052 5494
rect 6031 5487 6038 5491
rect 6038 5486 6039 5487
rect 5997 5480 6007 5486
rect 5756 5472 5791 5480
rect 5756 5446 5757 5472
rect 5764 5446 5791 5472
rect 5699 5428 5729 5442
rect 5756 5438 5791 5446
rect 5793 5472 5834 5480
rect 5793 5446 5808 5472
rect 5815 5446 5834 5472
rect 5898 5468 5929 5480
rect 5944 5468 6047 5480
rect 6059 5470 6085 5496
rect 6100 5491 6130 5502
rect 6162 5498 6224 5514
rect 6162 5496 6208 5498
rect 6162 5480 6224 5496
rect 6236 5480 6242 5528
rect 6245 5520 6325 5528
rect 6245 5518 6264 5520
rect 6279 5518 6313 5520
rect 6245 5502 6325 5518
rect 6245 5480 6264 5502
rect 6279 5486 6309 5502
rect 6337 5496 6343 5570
rect 6346 5496 6365 5640
rect 6380 5496 6386 5640
rect 6395 5570 6408 5640
rect 6460 5636 6482 5640
rect 6453 5614 6482 5628
rect 6535 5614 6551 5628
rect 6589 5624 6595 5626
rect 6602 5624 6710 5640
rect 6717 5624 6723 5626
rect 6731 5624 6746 5640
rect 6812 5634 6831 5637
rect 6453 5612 6551 5614
rect 6578 5612 6746 5624
rect 6761 5614 6777 5628
rect 6812 5615 6834 5634
rect 6844 5628 6860 5629
rect 6843 5626 6860 5628
rect 6844 5621 6860 5626
rect 6834 5614 6840 5615
rect 6843 5614 6872 5621
rect 6761 5613 6872 5614
rect 6761 5612 6878 5613
rect 6437 5604 6488 5612
rect 6535 5604 6569 5612
rect 6437 5592 6462 5604
rect 6469 5592 6488 5604
rect 6542 5602 6569 5604
rect 6578 5602 6799 5612
rect 6834 5609 6840 5612
rect 6542 5598 6799 5602
rect 6437 5584 6488 5592
rect 6535 5584 6799 5598
rect 6843 5604 6878 5612
rect 6389 5536 6408 5570
rect 6453 5576 6482 5584
rect 6453 5570 6470 5576
rect 6453 5568 6487 5570
rect 6535 5568 6551 5584
rect 6552 5574 6760 5584
rect 6761 5574 6777 5584
rect 6825 5580 6840 5595
rect 6843 5592 6844 5604
rect 6851 5592 6878 5604
rect 6843 5584 6878 5592
rect 6843 5583 6872 5584
rect 6563 5570 6777 5574
rect 6578 5568 6777 5570
rect 6812 5570 6825 5580
rect 6843 5570 6860 5583
rect 6812 5568 6860 5570
rect 6454 5564 6487 5568
rect 6450 5562 6487 5564
rect 6450 5561 6517 5562
rect 6450 5556 6481 5561
rect 6487 5556 6517 5561
rect 6450 5552 6517 5556
rect 6423 5549 6517 5552
rect 6423 5542 6472 5549
rect 6423 5536 6453 5542
rect 6472 5537 6477 5542
rect 6389 5520 6469 5536
rect 6481 5528 6517 5549
rect 6578 5544 6767 5568
rect 6812 5567 6859 5568
rect 6825 5562 6859 5567
rect 6593 5541 6767 5544
rect 6586 5538 6767 5541
rect 6795 5561 6859 5562
rect 6389 5518 6408 5520
rect 6423 5518 6457 5520
rect 6389 5502 6469 5518
rect 6389 5496 6408 5502
rect 6105 5470 6208 5480
rect 6059 5468 6208 5470
rect 6229 5468 6264 5480
rect 5898 5466 6060 5468
rect 5910 5446 5929 5466
rect 5944 5464 5974 5466
rect 5793 5438 5834 5446
rect 5916 5442 5929 5446
rect 5981 5450 6060 5466
rect 6092 5466 6264 5468
rect 6092 5450 6171 5466
rect 6178 5464 6208 5466
rect 5756 5428 5785 5438
rect 5799 5428 5828 5438
rect 5843 5428 5873 5442
rect 5916 5428 5959 5442
rect 5981 5438 6171 5450
rect 6236 5446 6242 5466
rect 5966 5428 5996 5438
rect 5997 5428 6155 5438
rect 6159 5428 6189 5438
rect 6193 5428 6223 5442
rect 6251 5428 6264 5466
rect 6336 5480 6365 5496
rect 6379 5480 6408 5496
rect 6423 5486 6453 5502
rect 6481 5480 6487 5528
rect 6490 5522 6509 5528
rect 6524 5522 6554 5530
rect 6490 5514 6554 5522
rect 6490 5498 6570 5514
rect 6586 5507 6648 5538
rect 6664 5507 6726 5538
rect 6795 5536 6844 5561
rect 6859 5536 6889 5552
rect 6758 5522 6788 5530
rect 6795 5528 6905 5536
rect 6758 5514 6803 5522
rect 6490 5496 6509 5498
rect 6524 5496 6570 5498
rect 6490 5480 6570 5496
rect 6597 5494 6632 5507
rect 6673 5504 6710 5507
rect 6673 5502 6715 5504
rect 6602 5491 6632 5494
rect 6611 5487 6618 5491
rect 6618 5486 6619 5487
rect 6577 5480 6587 5486
rect 6336 5472 6371 5480
rect 6336 5446 6337 5472
rect 6344 5446 6371 5472
rect 6279 5428 6309 5442
rect 6336 5438 6371 5446
rect 6373 5472 6414 5480
rect 6373 5446 6388 5472
rect 6395 5446 6414 5472
rect 6478 5468 6509 5480
rect 6524 5468 6627 5480
rect 6639 5470 6665 5496
rect 6680 5491 6710 5502
rect 6742 5498 6804 5514
rect 6742 5496 6788 5498
rect 6742 5480 6804 5496
rect 6816 5480 6822 5528
rect 6825 5520 6905 5528
rect 6825 5518 6844 5520
rect 6859 5518 6893 5520
rect 6825 5502 6905 5518
rect 6825 5480 6844 5502
rect 6859 5486 6889 5502
rect 6917 5496 6923 5570
rect 6926 5496 6945 5640
rect 6960 5496 6966 5640
rect 6975 5570 6988 5640
rect 7040 5636 7062 5640
rect 7033 5614 7062 5628
rect 7115 5614 7131 5628
rect 7169 5624 7175 5626
rect 7182 5624 7290 5640
rect 7297 5624 7303 5626
rect 7311 5624 7326 5640
rect 7392 5634 7411 5637
rect 7033 5612 7131 5614
rect 7158 5612 7326 5624
rect 7341 5614 7357 5628
rect 7392 5615 7414 5634
rect 7424 5628 7440 5629
rect 7423 5626 7440 5628
rect 7424 5621 7440 5626
rect 7414 5614 7420 5615
rect 7423 5614 7452 5621
rect 7341 5613 7452 5614
rect 7341 5612 7458 5613
rect 7017 5604 7068 5612
rect 7115 5604 7149 5612
rect 7017 5592 7042 5604
rect 7049 5592 7068 5604
rect 7122 5602 7149 5604
rect 7158 5602 7379 5612
rect 7414 5609 7420 5612
rect 7122 5598 7379 5602
rect 7017 5584 7068 5592
rect 7115 5584 7379 5598
rect 7423 5604 7458 5612
rect 6969 5536 6988 5570
rect 7033 5576 7062 5584
rect 7033 5570 7050 5576
rect 7033 5568 7067 5570
rect 7115 5568 7131 5584
rect 7132 5574 7340 5584
rect 7341 5574 7357 5584
rect 7405 5580 7420 5595
rect 7423 5592 7424 5604
rect 7431 5592 7458 5604
rect 7423 5584 7458 5592
rect 7423 5583 7452 5584
rect 7143 5570 7357 5574
rect 7158 5568 7357 5570
rect 7392 5570 7405 5580
rect 7423 5570 7440 5583
rect 7392 5568 7440 5570
rect 7034 5564 7067 5568
rect 7030 5562 7067 5564
rect 7030 5561 7097 5562
rect 7030 5556 7061 5561
rect 7067 5556 7097 5561
rect 7030 5552 7097 5556
rect 7003 5549 7097 5552
rect 7003 5542 7052 5549
rect 7003 5536 7033 5542
rect 7052 5537 7057 5542
rect 6969 5520 7049 5536
rect 7061 5528 7097 5549
rect 7158 5544 7347 5568
rect 7392 5567 7439 5568
rect 7405 5562 7439 5567
rect 7173 5541 7347 5544
rect 7166 5538 7347 5541
rect 7375 5561 7439 5562
rect 6969 5518 6988 5520
rect 7003 5518 7037 5520
rect 6969 5502 7049 5518
rect 6969 5496 6988 5502
rect 6685 5470 6788 5480
rect 6639 5468 6788 5470
rect 6809 5468 6844 5480
rect 6478 5466 6640 5468
rect 6490 5446 6509 5466
rect 6524 5464 6554 5466
rect 6373 5438 6414 5446
rect 6496 5442 6509 5446
rect 6561 5450 6640 5466
rect 6672 5466 6844 5468
rect 6672 5450 6751 5466
rect 6758 5464 6788 5466
rect 6336 5428 6365 5438
rect 6379 5428 6408 5438
rect 6423 5428 6453 5442
rect 6496 5428 6539 5442
rect 6561 5438 6751 5450
rect 6816 5446 6822 5466
rect 6546 5428 6576 5438
rect 6577 5428 6735 5438
rect 6739 5428 6769 5438
rect 6773 5428 6803 5442
rect 6831 5428 6844 5466
rect 6916 5480 6945 5496
rect 6959 5480 6988 5496
rect 7003 5486 7033 5502
rect 7061 5480 7067 5528
rect 7070 5522 7089 5528
rect 7104 5522 7134 5530
rect 7070 5514 7134 5522
rect 7070 5498 7150 5514
rect 7166 5507 7228 5538
rect 7244 5507 7306 5538
rect 7375 5536 7424 5561
rect 7439 5536 7469 5552
rect 7338 5522 7368 5530
rect 7375 5528 7485 5536
rect 7338 5514 7383 5522
rect 7070 5496 7089 5498
rect 7104 5496 7150 5498
rect 7070 5480 7150 5496
rect 7177 5494 7212 5507
rect 7253 5504 7290 5507
rect 7253 5502 7295 5504
rect 7182 5491 7212 5494
rect 7191 5487 7198 5491
rect 7198 5486 7199 5487
rect 7157 5480 7167 5486
rect 6916 5472 6951 5480
rect 6916 5446 6917 5472
rect 6924 5446 6951 5472
rect 6859 5428 6889 5442
rect 6916 5438 6951 5446
rect 6953 5472 6994 5480
rect 6953 5446 6968 5472
rect 6975 5446 6994 5472
rect 7058 5468 7089 5480
rect 7104 5468 7207 5480
rect 7219 5470 7245 5496
rect 7260 5491 7290 5502
rect 7322 5498 7384 5514
rect 7322 5496 7368 5498
rect 7322 5480 7384 5496
rect 7396 5480 7402 5528
rect 7405 5520 7485 5528
rect 7405 5518 7424 5520
rect 7439 5518 7473 5520
rect 7405 5502 7485 5518
rect 7405 5480 7424 5502
rect 7439 5486 7469 5502
rect 7497 5496 7503 5570
rect 7506 5496 7525 5640
rect 7540 5496 7546 5640
rect 7555 5570 7568 5640
rect 7613 5618 7614 5628
rect 7629 5618 7642 5628
rect 7613 5614 7642 5618
rect 7647 5614 7677 5640
rect 7695 5626 7711 5628
rect 7783 5626 7836 5640
rect 7784 5624 7848 5626
rect 7891 5624 7906 5640
rect 7955 5637 7985 5640
rect 7955 5634 7991 5637
rect 7921 5626 7937 5628
rect 7695 5614 7710 5618
rect 7613 5612 7710 5614
rect 7738 5612 7906 5624
rect 7922 5614 7937 5618
rect 7955 5615 7994 5634
rect 8013 5628 8020 5629
rect 8019 5621 8020 5628
rect 8003 5618 8004 5621
rect 8019 5618 8032 5621
rect 7955 5614 7985 5615
rect 7994 5614 8000 5615
rect 8003 5614 8032 5618
rect 7922 5613 8032 5614
rect 7922 5612 8038 5613
rect 7597 5604 7648 5612
rect 7597 5592 7622 5604
rect 7629 5592 7648 5604
rect 7679 5604 7729 5612
rect 7679 5596 7695 5604
rect 7702 5602 7729 5604
rect 7738 5602 7959 5612
rect 7702 5592 7959 5602
rect 7988 5604 8038 5612
rect 7988 5595 8004 5604
rect 7597 5584 7648 5592
rect 7695 5584 7959 5592
rect 7985 5592 8004 5595
rect 8011 5592 8038 5604
rect 7985 5584 8038 5592
rect 7549 5536 7568 5570
rect 7613 5576 7614 5584
rect 7629 5576 7642 5584
rect 7613 5568 7629 5576
rect 7610 5561 7629 5564
rect 7610 5552 7632 5561
rect 7583 5542 7632 5552
rect 7583 5536 7613 5542
rect 7632 5537 7637 5542
rect 7549 5520 7629 5536
rect 7647 5528 7677 5584
rect 7712 5574 7920 5584
rect 7955 5580 8000 5584
rect 8003 5583 8004 5584
rect 8019 5583 8032 5584
rect 7738 5544 7927 5574
rect 7753 5541 7927 5544
rect 7746 5538 7927 5541
rect 7549 5518 7568 5520
rect 7583 5518 7617 5520
rect 7549 5502 7629 5518
rect 7656 5514 7669 5528
rect 7684 5514 7700 5530
rect 7746 5525 7757 5538
rect 7549 5496 7568 5502
rect 7265 5470 7368 5480
rect 7219 5468 7368 5470
rect 7389 5468 7424 5480
rect 7058 5466 7220 5468
rect 7070 5446 7089 5466
rect 7104 5464 7134 5466
rect 6953 5438 6994 5446
rect 7076 5442 7089 5446
rect 7141 5450 7220 5466
rect 7252 5466 7424 5468
rect 7252 5450 7331 5466
rect 7338 5464 7368 5466
rect 6916 5428 6945 5438
rect 6959 5428 6988 5438
rect 7003 5428 7033 5442
rect 7076 5428 7119 5442
rect 7141 5438 7331 5450
rect 7396 5446 7402 5466
rect 7126 5428 7156 5438
rect 7157 5428 7315 5438
rect 7319 5428 7349 5438
rect 7353 5428 7383 5442
rect 7411 5428 7424 5466
rect 7496 5480 7525 5496
rect 7539 5480 7568 5496
rect 7583 5480 7613 5502
rect 7656 5498 7718 5514
rect 7746 5507 7757 5523
rect 7762 5518 7772 5538
rect 7782 5518 7796 5538
rect 7799 5525 7808 5538
rect 7824 5525 7833 5538
rect 7762 5507 7796 5518
rect 7799 5507 7808 5523
rect 7824 5507 7833 5523
rect 7840 5518 7850 5538
rect 7860 5518 7874 5538
rect 7875 5525 7886 5538
rect 7840 5507 7874 5518
rect 7875 5507 7886 5523
rect 7932 5514 7948 5530
rect 7955 5528 7985 5580
rect 8019 5576 8020 5583
rect 8004 5568 8020 5576
rect 7991 5536 8004 5555
rect 8019 5536 8049 5552
rect 7991 5520 8065 5536
rect 7991 5518 8004 5520
rect 8019 5518 8053 5520
rect 7656 5496 7669 5498
rect 7684 5496 7718 5498
rect 7656 5480 7718 5496
rect 7762 5491 7778 5494
rect 7840 5491 7870 5502
rect 7918 5498 7964 5514
rect 7991 5502 8065 5518
rect 7918 5496 7952 5498
rect 7917 5480 7964 5496
rect 7991 5480 8004 5502
rect 8019 5480 8049 5502
rect 8076 5480 8077 5496
rect 8092 5480 8105 5640
rect 8135 5536 8148 5640
rect 8193 5618 8194 5628
rect 8209 5618 8222 5628
rect 8193 5614 8222 5618
rect 8227 5614 8257 5640
rect 8275 5626 8291 5628
rect 8363 5626 8416 5640
rect 8364 5624 8428 5626
rect 8471 5624 8486 5640
rect 8535 5637 8565 5640
rect 8535 5634 8571 5637
rect 8501 5626 8517 5628
rect 8275 5614 8290 5618
rect 8193 5612 8290 5614
rect 8318 5612 8486 5624
rect 8502 5614 8517 5618
rect 8535 5615 8574 5634
rect 8593 5628 8600 5629
rect 8599 5621 8600 5628
rect 8583 5618 8584 5621
rect 8599 5618 8612 5621
rect 8535 5614 8565 5615
rect 8574 5614 8580 5615
rect 8583 5614 8612 5618
rect 8502 5613 8612 5614
rect 8502 5612 8618 5613
rect 8177 5604 8228 5612
rect 8177 5592 8202 5604
rect 8209 5592 8228 5604
rect 8259 5604 8309 5612
rect 8259 5596 8275 5604
rect 8282 5602 8309 5604
rect 8318 5602 8539 5612
rect 8282 5592 8539 5602
rect 8568 5604 8618 5612
rect 8568 5595 8584 5604
rect 8177 5584 8228 5592
rect 8275 5584 8539 5592
rect 8565 5592 8584 5595
rect 8591 5592 8618 5604
rect 8565 5584 8618 5592
rect 8193 5576 8194 5584
rect 8209 5576 8222 5584
rect 8193 5568 8209 5576
rect 8190 5561 8209 5564
rect 8190 5552 8212 5561
rect 8163 5542 8212 5552
rect 8163 5536 8193 5542
rect 8212 5537 8217 5542
rect 8135 5520 8209 5536
rect 8227 5528 8257 5584
rect 8292 5574 8500 5584
rect 8535 5580 8580 5584
rect 8583 5583 8584 5584
rect 8599 5583 8612 5584
rect 8318 5544 8507 5574
rect 8333 5541 8507 5544
rect 8326 5538 8507 5541
rect 8135 5518 8148 5520
rect 8163 5518 8197 5520
rect 8135 5502 8209 5518
rect 8236 5514 8249 5528
rect 8264 5514 8280 5530
rect 8326 5525 8337 5538
rect 8119 5480 8120 5496
rect 8135 5480 8148 5502
rect 8163 5480 8193 5502
rect 8236 5498 8298 5514
rect 8326 5507 8337 5523
rect 8342 5518 8352 5538
rect 8362 5518 8376 5538
rect 8379 5525 8388 5538
rect 8404 5525 8413 5538
rect 8342 5507 8376 5518
rect 8379 5507 8388 5523
rect 8404 5507 8413 5523
rect 8420 5518 8430 5538
rect 8440 5518 8454 5538
rect 8455 5525 8466 5538
rect 8420 5507 8454 5518
rect 8455 5507 8466 5523
rect 8512 5514 8528 5530
rect 8535 5528 8565 5580
rect 8599 5576 8600 5583
rect 8584 5568 8600 5576
rect 8571 5536 8584 5555
rect 8599 5536 8629 5552
rect 8571 5520 8645 5536
rect 8571 5518 8584 5520
rect 8599 5518 8633 5520
rect 8236 5496 8249 5498
rect 8264 5496 8298 5498
rect 8236 5480 8298 5496
rect 8342 5491 8358 5494
rect 8420 5491 8450 5502
rect 8498 5498 8544 5514
rect 8571 5502 8645 5518
rect 8498 5496 8532 5498
rect 8497 5480 8544 5496
rect 8571 5480 8584 5502
rect 8599 5480 8629 5502
rect 8656 5480 8657 5496
rect 8672 5480 8685 5640
rect 8715 5536 8728 5640
rect 8773 5618 8774 5628
rect 8789 5618 8802 5628
rect 8773 5614 8802 5618
rect 8807 5614 8837 5640
rect 8855 5626 8871 5628
rect 8943 5626 8996 5640
rect 8944 5624 9008 5626
rect 9051 5624 9066 5640
rect 9115 5637 9145 5640
rect 9115 5634 9151 5637
rect 9081 5626 9097 5628
rect 8855 5614 8870 5618
rect 8773 5612 8870 5614
rect 8898 5612 9066 5624
rect 9082 5614 9097 5618
rect 9115 5615 9154 5634
rect 9173 5628 9180 5629
rect 9179 5621 9180 5628
rect 9163 5618 9164 5621
rect 9179 5618 9192 5621
rect 9115 5614 9145 5615
rect 9154 5614 9160 5615
rect 9163 5614 9192 5618
rect 9082 5613 9192 5614
rect 9082 5612 9198 5613
rect 8757 5604 8808 5612
rect 8757 5592 8782 5604
rect 8789 5592 8808 5604
rect 8839 5604 8889 5612
rect 8839 5596 8855 5604
rect 8862 5602 8889 5604
rect 8898 5602 9119 5612
rect 8862 5592 9119 5602
rect 9148 5604 9198 5612
rect 9148 5595 9164 5604
rect 8757 5584 8808 5592
rect 8855 5584 9119 5592
rect 9145 5592 9164 5595
rect 9171 5592 9198 5604
rect 9145 5584 9198 5592
rect 8773 5576 8774 5584
rect 8789 5576 8802 5584
rect 8773 5568 8789 5576
rect 8770 5561 8789 5564
rect 8770 5552 8792 5561
rect 8743 5542 8792 5552
rect 8743 5536 8773 5542
rect 8792 5537 8797 5542
rect 8715 5520 8789 5536
rect 8807 5528 8837 5584
rect 8872 5574 9080 5584
rect 9115 5580 9160 5584
rect 9163 5583 9164 5584
rect 9179 5583 9192 5584
rect 8898 5544 9087 5574
rect 8913 5541 9087 5544
rect 8906 5538 9087 5541
rect 8715 5518 8728 5520
rect 8743 5518 8777 5520
rect 8715 5502 8789 5518
rect 8816 5514 8829 5528
rect 8844 5514 8860 5530
rect 8906 5525 8917 5538
rect 8699 5480 8700 5496
rect 8715 5480 8728 5502
rect 8743 5480 8773 5502
rect 8816 5498 8878 5514
rect 8906 5507 8917 5523
rect 8922 5518 8932 5538
rect 8942 5518 8956 5538
rect 8959 5525 8968 5538
rect 8984 5525 8993 5538
rect 8922 5507 8956 5518
rect 8959 5507 8968 5523
rect 8984 5507 8993 5523
rect 9000 5518 9010 5538
rect 9020 5518 9034 5538
rect 9035 5525 9046 5538
rect 9000 5507 9034 5518
rect 9035 5507 9046 5523
rect 9092 5514 9108 5530
rect 9115 5528 9145 5580
rect 9179 5576 9180 5583
rect 9164 5568 9180 5576
rect 9151 5536 9164 5555
rect 9179 5536 9209 5552
rect 9151 5520 9225 5536
rect 9151 5518 9164 5520
rect 9179 5518 9213 5520
rect 8816 5496 8829 5498
rect 8844 5496 8878 5498
rect 8816 5480 8878 5496
rect 8922 5491 8938 5494
rect 9000 5491 9030 5502
rect 9078 5498 9124 5514
rect 9151 5502 9225 5518
rect 9078 5496 9112 5498
rect 9077 5480 9124 5496
rect 9151 5480 9164 5502
rect 9179 5480 9209 5502
rect 9236 5480 9237 5496
rect 9252 5480 9265 5640
rect 7496 5472 7531 5480
rect 7496 5446 7497 5472
rect 7504 5446 7531 5472
rect 7439 5428 7469 5442
rect 7496 5438 7531 5446
rect 7533 5472 7574 5480
rect 7533 5446 7548 5472
rect 7555 5446 7574 5472
rect 7638 5468 7700 5480
rect 7712 5468 7787 5480
rect 7845 5468 7920 5480
rect 7932 5468 7963 5480
rect 7969 5468 8004 5480
rect 7638 5466 7800 5468
rect 7533 5438 7574 5446
rect 7656 5442 7669 5466
rect 7684 5464 7699 5466
rect 7496 5428 7525 5438
rect 7539 5428 7568 5438
rect 7583 5428 7613 5442
rect 7656 5428 7699 5442
rect 7723 5439 7730 5446
rect 7733 5442 7800 5466
rect 7832 5466 8004 5468
rect 7802 5444 7830 5448
rect 7832 5444 7912 5466
rect 7933 5464 7948 5466
rect 7802 5442 7912 5444
rect 7733 5438 7912 5442
rect 7706 5428 7736 5438
rect 7738 5428 7891 5438
rect 7899 5428 7929 5438
rect 7933 5428 7963 5442
rect 7991 5428 8004 5466
rect 8076 5472 8111 5480
rect 8076 5446 8077 5472
rect 8084 5446 8111 5472
rect 8019 5428 8049 5442
rect 8076 5438 8111 5446
rect 8113 5472 8154 5480
rect 8113 5446 8128 5472
rect 8135 5446 8154 5472
rect 8218 5468 8280 5480
rect 8292 5468 8367 5480
rect 8425 5468 8500 5480
rect 8512 5468 8543 5480
rect 8549 5468 8584 5480
rect 8218 5466 8380 5468
rect 8113 5438 8154 5446
rect 8236 5442 8249 5466
rect 8264 5464 8279 5466
rect 8076 5428 8077 5438
rect 8092 5428 8105 5438
rect 8119 5428 8120 5438
rect 8135 5428 8148 5438
rect 8163 5428 8193 5442
rect 8236 5428 8279 5442
rect 8303 5439 8310 5446
rect 8313 5442 8380 5466
rect 8412 5466 8584 5468
rect 8382 5444 8410 5448
rect 8412 5444 8492 5466
rect 8513 5464 8528 5466
rect 8382 5442 8492 5444
rect 8313 5438 8492 5442
rect 8286 5428 8316 5438
rect 8318 5428 8471 5438
rect 8479 5428 8509 5438
rect 8513 5428 8543 5442
rect 8571 5428 8584 5466
rect 8656 5472 8691 5480
rect 8656 5446 8657 5472
rect 8664 5446 8691 5472
rect 8599 5428 8629 5442
rect 8656 5438 8691 5446
rect 8693 5472 8734 5480
rect 8693 5446 8708 5472
rect 8715 5446 8734 5472
rect 8798 5468 8860 5480
rect 8872 5468 8947 5480
rect 9005 5468 9080 5480
rect 9092 5468 9123 5480
rect 9129 5468 9164 5480
rect 8798 5466 8960 5468
rect 8693 5438 8734 5446
rect 8816 5442 8829 5466
rect 8844 5464 8859 5466
rect 8656 5428 8657 5438
rect 8672 5428 8685 5438
rect 8699 5428 8700 5438
rect 8715 5428 8728 5438
rect 8743 5428 8773 5442
rect 8816 5428 8859 5442
rect 8883 5439 8890 5446
rect 8893 5442 8960 5466
rect 8992 5466 9164 5468
rect 8962 5444 8990 5448
rect 8992 5444 9072 5466
rect 9093 5464 9108 5466
rect 8962 5442 9072 5444
rect 8893 5438 9072 5442
rect 8866 5428 8896 5438
rect 8898 5428 9051 5438
rect 9059 5428 9089 5438
rect 9093 5428 9123 5442
rect 9151 5428 9164 5466
rect 9236 5472 9271 5480
rect 9236 5446 9237 5472
rect 9244 5446 9271 5472
rect 9179 5428 9209 5442
rect 9236 5438 9271 5446
rect 9236 5428 9237 5438
rect 9252 5428 9265 5438
rect -1 5422 9265 5428
rect 0 5414 9265 5422
rect 15 5384 28 5414
rect 43 5400 73 5414
rect 116 5400 159 5414
rect 166 5400 386 5414
rect 393 5400 423 5414
rect 83 5386 98 5398
rect 117 5386 130 5400
rect 198 5396 351 5400
rect 80 5384 102 5386
rect 180 5384 372 5396
rect 451 5384 464 5414
rect 479 5400 509 5414
rect 546 5384 565 5414
rect 580 5384 586 5414
rect 595 5384 608 5414
rect 623 5400 653 5414
rect 696 5400 739 5414
rect 746 5400 966 5414
rect 973 5400 1003 5414
rect 663 5386 678 5398
rect 697 5386 710 5400
rect 778 5396 931 5400
rect 660 5384 682 5386
rect 760 5384 952 5396
rect 1031 5384 1044 5414
rect 1059 5400 1089 5414
rect 1126 5384 1145 5414
rect 1160 5384 1166 5414
rect 1175 5384 1188 5414
rect 1203 5400 1233 5414
rect 1276 5400 1319 5414
rect 1326 5400 1546 5414
rect 1553 5400 1583 5414
rect 1243 5386 1258 5398
rect 1277 5386 1290 5400
rect 1358 5396 1511 5400
rect 1240 5384 1262 5386
rect 1340 5384 1532 5396
rect 1611 5384 1624 5414
rect 1639 5400 1669 5414
rect 1706 5384 1725 5414
rect 1740 5384 1746 5414
rect 1755 5384 1768 5414
rect 1783 5400 1813 5414
rect 1856 5400 1899 5414
rect 1906 5400 2126 5414
rect 2133 5400 2163 5414
rect 1823 5386 1838 5398
rect 1857 5386 1870 5400
rect 1938 5396 2091 5400
rect 1820 5384 1842 5386
rect 1920 5384 2112 5396
rect 2191 5384 2204 5414
rect 2219 5400 2249 5414
rect 2286 5384 2305 5414
rect 2320 5384 2326 5414
rect 2335 5384 2348 5414
rect 2363 5400 2393 5414
rect 2436 5400 2479 5414
rect 2486 5400 2706 5414
rect 2713 5400 2743 5414
rect 2403 5386 2418 5398
rect 2437 5386 2450 5400
rect 2518 5396 2671 5400
rect 2400 5384 2422 5386
rect 2500 5384 2692 5396
rect 2771 5384 2784 5414
rect 2799 5400 2829 5414
rect 2866 5384 2885 5414
rect 2900 5384 2906 5414
rect 2915 5384 2928 5414
rect 2943 5400 2973 5414
rect 3016 5400 3059 5414
rect 3066 5400 3286 5414
rect 3293 5400 3323 5414
rect 2983 5386 2998 5398
rect 3017 5386 3030 5400
rect 3098 5396 3251 5400
rect 2980 5384 3002 5386
rect 3080 5384 3272 5396
rect 3351 5384 3364 5414
rect 3379 5400 3409 5414
rect 3446 5384 3465 5414
rect 3480 5384 3486 5414
rect 3495 5384 3508 5414
rect 3523 5400 3553 5414
rect 3596 5400 3639 5414
rect 3646 5400 3866 5414
rect 3873 5400 3903 5414
rect 3563 5386 3578 5398
rect 3597 5386 3610 5400
rect 3678 5396 3831 5400
rect 3560 5384 3582 5386
rect 3660 5384 3852 5396
rect 3931 5384 3944 5414
rect 3959 5400 3989 5414
rect 4026 5384 4045 5414
rect 4060 5384 4066 5414
rect 4075 5384 4088 5414
rect 4103 5400 4133 5414
rect 4176 5400 4219 5414
rect 4226 5400 4446 5414
rect 4453 5400 4483 5414
rect 4143 5386 4158 5398
rect 4177 5386 4190 5400
rect 4258 5396 4411 5400
rect 4140 5384 4162 5386
rect 4240 5384 4432 5396
rect 4511 5384 4524 5414
rect 4539 5400 4569 5414
rect 4606 5384 4625 5414
rect 4640 5384 4646 5414
rect 4655 5384 4668 5414
rect 4683 5400 4713 5414
rect 4756 5400 4799 5414
rect 4806 5400 5026 5414
rect 5033 5400 5063 5414
rect 4723 5386 4738 5398
rect 4757 5386 4770 5400
rect 4838 5396 4991 5400
rect 4720 5384 4742 5386
rect 4820 5384 5012 5396
rect 5091 5384 5104 5414
rect 5119 5400 5149 5414
rect 5186 5384 5205 5414
rect 5220 5384 5226 5414
rect 5235 5384 5248 5414
rect 5263 5400 5293 5414
rect 5336 5400 5379 5414
rect 5386 5400 5606 5414
rect 5613 5400 5643 5414
rect 5303 5386 5318 5398
rect 5337 5386 5350 5400
rect 5418 5396 5571 5400
rect 5300 5384 5322 5386
rect 5400 5384 5592 5396
rect 5671 5384 5684 5414
rect 5699 5400 5729 5414
rect 5766 5384 5785 5414
rect 5800 5384 5806 5414
rect 5815 5384 5828 5414
rect 5843 5400 5873 5414
rect 5916 5400 5959 5414
rect 5966 5400 6186 5414
rect 6193 5400 6223 5414
rect 5883 5386 5898 5398
rect 5917 5386 5930 5400
rect 5998 5396 6151 5400
rect 5880 5384 5902 5386
rect 5980 5384 6172 5396
rect 6251 5384 6264 5414
rect 6279 5400 6309 5414
rect 6346 5384 6365 5414
rect 6380 5384 6386 5414
rect 6395 5384 6408 5414
rect 6423 5400 6453 5414
rect 6496 5400 6539 5414
rect 6546 5400 6766 5414
rect 6773 5400 6803 5414
rect 6463 5386 6478 5398
rect 6497 5386 6510 5400
rect 6578 5396 6731 5400
rect 6460 5384 6482 5386
rect 6560 5384 6752 5396
rect 6831 5384 6844 5414
rect 6859 5400 6889 5414
rect 6926 5384 6945 5414
rect 6960 5384 6966 5414
rect 6975 5384 6988 5414
rect 7003 5400 7033 5414
rect 7076 5400 7119 5414
rect 7126 5400 7346 5414
rect 7353 5400 7383 5414
rect 7043 5386 7058 5398
rect 7077 5386 7090 5400
rect 7158 5396 7311 5400
rect 7040 5384 7062 5386
rect 7140 5384 7332 5396
rect 7411 5384 7424 5414
rect 7439 5400 7469 5414
rect 7506 5384 7525 5414
rect 7540 5384 7546 5414
rect 7555 5384 7568 5414
rect 7583 5396 7613 5414
rect 7656 5400 7670 5414
rect 7706 5400 7926 5414
rect 7657 5398 7670 5400
rect 7623 5386 7638 5398
rect 7620 5384 7642 5386
rect 7647 5384 7677 5398
rect 7738 5396 7891 5400
rect 7720 5384 7912 5396
rect 7955 5384 7985 5398
rect 7991 5384 8004 5414
rect 8019 5396 8049 5414
rect 8092 5384 8105 5414
rect 8135 5384 8148 5414
rect 8163 5396 8193 5414
rect 8236 5400 8250 5414
rect 8286 5400 8506 5414
rect 8237 5398 8250 5400
rect 8203 5386 8218 5398
rect 8200 5384 8222 5386
rect 8227 5384 8257 5398
rect 8318 5396 8471 5400
rect 8300 5384 8492 5396
rect 8535 5384 8565 5398
rect 8571 5384 8584 5414
rect 8599 5396 8629 5414
rect 8672 5384 8685 5414
rect 8715 5384 8728 5414
rect 8743 5396 8773 5414
rect 8816 5400 8830 5414
rect 8866 5400 9086 5414
rect 8817 5398 8830 5400
rect 8783 5386 8798 5398
rect 8780 5384 8802 5386
rect 8807 5384 8837 5398
rect 8898 5396 9051 5400
rect 8880 5384 9072 5396
rect 9115 5384 9145 5398
rect 9151 5384 9164 5414
rect 9179 5396 9209 5414
rect 9252 5384 9265 5414
rect 0 5370 9265 5384
rect 15 5300 28 5370
rect 80 5366 102 5370
rect 73 5344 102 5358
rect 155 5344 171 5358
rect 209 5354 215 5356
rect 222 5354 330 5370
rect 337 5354 343 5356
rect 351 5354 366 5370
rect 432 5364 451 5367
rect 73 5342 171 5344
rect 198 5342 366 5354
rect 381 5344 397 5358
rect 432 5345 454 5364
rect 464 5358 480 5359
rect 463 5356 480 5358
rect 464 5351 480 5356
rect 454 5344 460 5345
rect 463 5344 492 5351
rect 381 5343 492 5344
rect 381 5342 498 5343
rect 57 5334 108 5342
rect 155 5334 189 5342
rect 57 5322 82 5334
rect 89 5322 108 5334
rect 162 5332 189 5334
rect 198 5332 419 5342
rect 454 5339 460 5342
rect 162 5328 419 5332
rect 57 5314 108 5322
rect 155 5314 419 5328
rect 463 5334 498 5342
rect 9 5266 28 5300
rect 73 5306 102 5314
rect 73 5300 90 5306
rect 73 5298 107 5300
rect 155 5298 171 5314
rect 172 5304 380 5314
rect 381 5304 397 5314
rect 445 5310 460 5325
rect 463 5322 464 5334
rect 471 5322 498 5334
rect 463 5314 498 5322
rect 463 5313 492 5314
rect 183 5300 397 5304
rect 198 5298 397 5300
rect 432 5300 445 5310
rect 463 5300 480 5313
rect 432 5298 480 5300
rect 74 5294 107 5298
rect 70 5292 107 5294
rect 70 5291 137 5292
rect 70 5286 101 5291
rect 107 5286 137 5291
rect 70 5282 137 5286
rect 43 5279 137 5282
rect 43 5272 92 5279
rect 43 5266 73 5272
rect 92 5267 97 5272
rect 9 5250 89 5266
rect 101 5258 137 5279
rect 198 5274 387 5298
rect 432 5297 479 5298
rect 445 5292 479 5297
rect 213 5271 387 5274
rect 206 5268 387 5271
rect 415 5291 479 5292
rect 9 5248 28 5250
rect 43 5248 77 5250
rect 9 5232 89 5248
rect 9 5226 28 5232
rect -1 5210 28 5226
rect 43 5216 73 5232
rect 101 5210 107 5258
rect 110 5252 129 5258
rect 144 5252 174 5260
rect 110 5244 174 5252
rect 110 5228 190 5244
rect 206 5237 268 5268
rect 284 5237 346 5268
rect 415 5266 464 5291
rect 479 5266 509 5282
rect 378 5252 408 5260
rect 415 5258 525 5266
rect 378 5244 423 5252
rect 110 5226 129 5228
rect 144 5226 190 5228
rect 110 5210 190 5226
rect 217 5224 252 5237
rect 293 5234 330 5237
rect 293 5232 335 5234
rect 222 5221 252 5224
rect 231 5217 238 5221
rect 238 5216 239 5217
rect 197 5210 207 5216
rect -7 5202 34 5210
rect -7 5176 8 5202
rect 15 5176 34 5202
rect 98 5198 129 5210
rect 144 5198 247 5210
rect 259 5200 285 5226
rect 300 5221 330 5232
rect 362 5228 424 5244
rect 362 5226 408 5228
rect 362 5210 424 5226
rect 436 5210 442 5258
rect 445 5250 525 5258
rect 445 5248 464 5250
rect 479 5248 513 5250
rect 445 5232 525 5248
rect 445 5210 464 5232
rect 479 5216 509 5232
rect 537 5226 543 5300
rect 546 5226 565 5370
rect 580 5226 586 5370
rect 595 5300 608 5370
rect 660 5366 682 5370
rect 653 5344 682 5358
rect 735 5344 751 5358
rect 789 5354 795 5356
rect 802 5354 910 5370
rect 917 5354 923 5356
rect 931 5354 946 5370
rect 1012 5364 1031 5367
rect 653 5342 751 5344
rect 778 5342 946 5354
rect 961 5344 977 5358
rect 1012 5345 1034 5364
rect 1044 5358 1060 5359
rect 1043 5356 1060 5358
rect 1044 5351 1060 5356
rect 1034 5344 1040 5345
rect 1043 5344 1072 5351
rect 961 5343 1072 5344
rect 961 5342 1078 5343
rect 637 5334 688 5342
rect 735 5334 769 5342
rect 637 5322 662 5334
rect 669 5322 688 5334
rect 742 5332 769 5334
rect 778 5332 999 5342
rect 1034 5339 1040 5342
rect 742 5328 999 5332
rect 637 5314 688 5322
rect 735 5314 999 5328
rect 1043 5334 1078 5342
rect 589 5266 608 5300
rect 653 5306 682 5314
rect 653 5300 670 5306
rect 653 5298 687 5300
rect 735 5298 751 5314
rect 752 5304 960 5314
rect 961 5304 977 5314
rect 1025 5310 1040 5325
rect 1043 5322 1044 5334
rect 1051 5322 1078 5334
rect 1043 5314 1078 5322
rect 1043 5313 1072 5314
rect 763 5300 977 5304
rect 778 5298 977 5300
rect 1012 5300 1025 5310
rect 1043 5300 1060 5313
rect 1012 5298 1060 5300
rect 654 5294 687 5298
rect 650 5292 687 5294
rect 650 5291 717 5292
rect 650 5286 681 5291
rect 687 5286 717 5291
rect 650 5282 717 5286
rect 623 5279 717 5282
rect 623 5272 672 5279
rect 623 5266 653 5272
rect 672 5267 677 5272
rect 589 5250 669 5266
rect 681 5258 717 5279
rect 778 5274 967 5298
rect 1012 5297 1059 5298
rect 1025 5292 1059 5297
rect 793 5271 967 5274
rect 786 5268 967 5271
rect 995 5291 1059 5292
rect 589 5248 608 5250
rect 623 5248 657 5250
rect 589 5232 669 5248
rect 589 5226 608 5232
rect 305 5200 408 5210
rect 259 5198 408 5200
rect 429 5198 464 5210
rect 98 5196 260 5198
rect 110 5176 129 5196
rect 144 5194 174 5196
rect -7 5168 34 5176
rect 116 5172 129 5176
rect 181 5180 260 5196
rect 292 5196 464 5198
rect 292 5180 371 5196
rect 378 5194 408 5196
rect -1 5158 28 5168
rect 43 5158 73 5172
rect 116 5158 159 5172
rect 181 5168 371 5180
rect 436 5176 442 5196
rect 166 5158 196 5168
rect 197 5158 355 5168
rect 359 5158 389 5168
rect 393 5158 423 5172
rect 451 5158 464 5196
rect 536 5210 565 5226
rect 579 5210 608 5226
rect 623 5216 653 5232
rect 681 5210 687 5258
rect 690 5252 709 5258
rect 724 5252 754 5260
rect 690 5244 754 5252
rect 690 5228 770 5244
rect 786 5237 848 5268
rect 864 5237 926 5268
rect 995 5266 1044 5291
rect 1059 5266 1089 5282
rect 958 5252 988 5260
rect 995 5258 1105 5266
rect 958 5244 1003 5252
rect 690 5226 709 5228
rect 724 5226 770 5228
rect 690 5210 770 5226
rect 797 5224 832 5237
rect 873 5234 910 5237
rect 873 5232 915 5234
rect 802 5221 832 5224
rect 811 5217 818 5221
rect 818 5216 819 5217
rect 777 5210 787 5216
rect 536 5202 571 5210
rect 536 5176 537 5202
rect 544 5176 571 5202
rect 479 5158 509 5172
rect 536 5168 571 5176
rect 573 5202 614 5210
rect 573 5176 588 5202
rect 595 5176 614 5202
rect 678 5198 709 5210
rect 724 5198 827 5210
rect 839 5200 865 5226
rect 880 5221 910 5232
rect 942 5228 1004 5244
rect 942 5226 988 5228
rect 942 5210 1004 5226
rect 1016 5210 1022 5258
rect 1025 5250 1105 5258
rect 1025 5248 1044 5250
rect 1059 5248 1093 5250
rect 1025 5232 1105 5248
rect 1025 5210 1044 5232
rect 1059 5216 1089 5232
rect 1117 5226 1123 5300
rect 1126 5226 1145 5370
rect 1160 5226 1166 5370
rect 1175 5300 1188 5370
rect 1240 5366 1262 5370
rect 1233 5344 1262 5358
rect 1315 5344 1331 5358
rect 1369 5354 1375 5356
rect 1382 5354 1490 5370
rect 1497 5354 1503 5356
rect 1511 5354 1526 5370
rect 1592 5364 1611 5367
rect 1233 5342 1331 5344
rect 1358 5342 1526 5354
rect 1541 5344 1557 5358
rect 1592 5345 1614 5364
rect 1624 5358 1640 5359
rect 1623 5356 1640 5358
rect 1624 5351 1640 5356
rect 1614 5344 1620 5345
rect 1623 5344 1652 5351
rect 1541 5343 1652 5344
rect 1541 5342 1658 5343
rect 1217 5334 1268 5342
rect 1315 5334 1349 5342
rect 1217 5322 1242 5334
rect 1249 5322 1268 5334
rect 1322 5332 1349 5334
rect 1358 5332 1579 5342
rect 1614 5339 1620 5342
rect 1322 5328 1579 5332
rect 1217 5314 1268 5322
rect 1315 5314 1579 5328
rect 1623 5334 1658 5342
rect 1169 5266 1188 5300
rect 1233 5306 1262 5314
rect 1233 5300 1250 5306
rect 1233 5298 1267 5300
rect 1315 5298 1331 5314
rect 1332 5304 1540 5314
rect 1541 5304 1557 5314
rect 1605 5310 1620 5325
rect 1623 5322 1624 5334
rect 1631 5322 1658 5334
rect 1623 5314 1658 5322
rect 1623 5313 1652 5314
rect 1343 5300 1557 5304
rect 1358 5298 1557 5300
rect 1592 5300 1605 5310
rect 1623 5300 1640 5313
rect 1592 5298 1640 5300
rect 1234 5294 1267 5298
rect 1230 5292 1267 5294
rect 1230 5291 1297 5292
rect 1230 5286 1261 5291
rect 1267 5286 1297 5291
rect 1230 5282 1297 5286
rect 1203 5279 1297 5282
rect 1203 5272 1252 5279
rect 1203 5266 1233 5272
rect 1252 5267 1257 5272
rect 1169 5250 1249 5266
rect 1261 5258 1297 5279
rect 1358 5274 1547 5298
rect 1592 5297 1639 5298
rect 1605 5292 1639 5297
rect 1373 5271 1547 5274
rect 1366 5268 1547 5271
rect 1575 5291 1639 5292
rect 1169 5248 1188 5250
rect 1203 5248 1237 5250
rect 1169 5232 1249 5248
rect 1169 5226 1188 5232
rect 885 5200 988 5210
rect 839 5198 988 5200
rect 1009 5198 1044 5210
rect 678 5196 840 5198
rect 690 5176 709 5196
rect 724 5194 754 5196
rect 573 5168 614 5176
rect 696 5172 709 5176
rect 761 5180 840 5196
rect 872 5196 1044 5198
rect 872 5180 951 5196
rect 958 5194 988 5196
rect 536 5158 565 5168
rect 579 5158 608 5168
rect 623 5158 653 5172
rect 696 5158 739 5172
rect 761 5168 951 5180
rect 1016 5176 1022 5196
rect 746 5158 776 5168
rect 777 5158 935 5168
rect 939 5158 969 5168
rect 973 5158 1003 5172
rect 1031 5158 1044 5196
rect 1116 5210 1145 5226
rect 1159 5210 1188 5226
rect 1203 5216 1233 5232
rect 1261 5210 1267 5258
rect 1270 5252 1289 5258
rect 1304 5252 1334 5260
rect 1270 5244 1334 5252
rect 1270 5228 1350 5244
rect 1366 5237 1428 5268
rect 1444 5237 1506 5268
rect 1575 5266 1624 5291
rect 1639 5266 1669 5282
rect 1538 5252 1568 5260
rect 1575 5258 1685 5266
rect 1538 5244 1583 5252
rect 1270 5226 1289 5228
rect 1304 5226 1350 5228
rect 1270 5210 1350 5226
rect 1377 5224 1412 5237
rect 1453 5234 1490 5237
rect 1453 5232 1495 5234
rect 1382 5221 1412 5224
rect 1391 5217 1398 5221
rect 1398 5216 1399 5217
rect 1357 5210 1367 5216
rect 1116 5202 1151 5210
rect 1116 5176 1117 5202
rect 1124 5176 1151 5202
rect 1059 5158 1089 5172
rect 1116 5168 1151 5176
rect 1153 5202 1194 5210
rect 1153 5176 1168 5202
rect 1175 5176 1194 5202
rect 1258 5198 1289 5210
rect 1304 5198 1407 5210
rect 1419 5200 1445 5226
rect 1460 5221 1490 5232
rect 1522 5228 1584 5244
rect 1522 5226 1568 5228
rect 1522 5210 1584 5226
rect 1596 5210 1602 5258
rect 1605 5250 1685 5258
rect 1605 5248 1624 5250
rect 1639 5248 1673 5250
rect 1605 5232 1685 5248
rect 1605 5210 1624 5232
rect 1639 5216 1669 5232
rect 1697 5226 1703 5300
rect 1706 5226 1725 5370
rect 1740 5226 1746 5370
rect 1755 5300 1768 5370
rect 1820 5366 1842 5370
rect 1813 5344 1842 5358
rect 1895 5344 1911 5358
rect 1949 5354 1955 5356
rect 1962 5354 2070 5370
rect 2077 5354 2083 5356
rect 2091 5354 2106 5370
rect 2172 5364 2191 5367
rect 1813 5342 1911 5344
rect 1938 5342 2106 5354
rect 2121 5344 2137 5358
rect 2172 5345 2194 5364
rect 2204 5358 2220 5359
rect 2203 5356 2220 5358
rect 2204 5351 2220 5356
rect 2194 5344 2200 5345
rect 2203 5344 2232 5351
rect 2121 5343 2232 5344
rect 2121 5342 2238 5343
rect 1797 5334 1848 5342
rect 1895 5334 1929 5342
rect 1797 5322 1822 5334
rect 1829 5322 1848 5334
rect 1902 5332 1929 5334
rect 1938 5332 2159 5342
rect 2194 5339 2200 5342
rect 1902 5328 2159 5332
rect 1797 5314 1848 5322
rect 1895 5314 2159 5328
rect 2203 5334 2238 5342
rect 1749 5266 1768 5300
rect 1813 5306 1842 5314
rect 1813 5300 1830 5306
rect 1813 5298 1847 5300
rect 1895 5298 1911 5314
rect 1912 5304 2120 5314
rect 2121 5304 2137 5314
rect 2185 5310 2200 5325
rect 2203 5322 2204 5334
rect 2211 5322 2238 5334
rect 2203 5314 2238 5322
rect 2203 5313 2232 5314
rect 1923 5300 2137 5304
rect 1938 5298 2137 5300
rect 2172 5300 2185 5310
rect 2203 5300 2220 5313
rect 2172 5298 2220 5300
rect 1814 5294 1847 5298
rect 1810 5292 1847 5294
rect 1810 5291 1877 5292
rect 1810 5286 1841 5291
rect 1847 5286 1877 5291
rect 1810 5282 1877 5286
rect 1783 5279 1877 5282
rect 1783 5272 1832 5279
rect 1783 5266 1813 5272
rect 1832 5267 1837 5272
rect 1749 5250 1829 5266
rect 1841 5258 1877 5279
rect 1938 5274 2127 5298
rect 2172 5297 2219 5298
rect 2185 5292 2219 5297
rect 1953 5271 2127 5274
rect 1946 5268 2127 5271
rect 2155 5291 2219 5292
rect 1749 5248 1768 5250
rect 1783 5248 1817 5250
rect 1749 5232 1829 5248
rect 1749 5226 1768 5232
rect 1465 5200 1568 5210
rect 1419 5198 1568 5200
rect 1589 5198 1624 5210
rect 1258 5196 1420 5198
rect 1270 5176 1289 5196
rect 1304 5194 1334 5196
rect 1153 5168 1194 5176
rect 1276 5172 1289 5176
rect 1341 5180 1420 5196
rect 1452 5196 1624 5198
rect 1452 5180 1531 5196
rect 1538 5194 1568 5196
rect 1116 5158 1145 5168
rect 1159 5158 1188 5168
rect 1203 5158 1233 5172
rect 1276 5158 1319 5172
rect 1341 5168 1531 5180
rect 1596 5176 1602 5196
rect 1326 5158 1356 5168
rect 1357 5158 1515 5168
rect 1519 5158 1549 5168
rect 1553 5158 1583 5172
rect 1611 5158 1624 5196
rect 1696 5210 1725 5226
rect 1739 5210 1768 5226
rect 1783 5216 1813 5232
rect 1841 5210 1847 5258
rect 1850 5252 1869 5258
rect 1884 5252 1914 5260
rect 1850 5244 1914 5252
rect 1850 5228 1930 5244
rect 1946 5237 2008 5268
rect 2024 5237 2086 5268
rect 2155 5266 2204 5291
rect 2219 5266 2249 5282
rect 2118 5252 2148 5260
rect 2155 5258 2265 5266
rect 2118 5244 2163 5252
rect 1850 5226 1869 5228
rect 1884 5226 1930 5228
rect 1850 5210 1930 5226
rect 1957 5224 1992 5237
rect 2033 5234 2070 5237
rect 2033 5232 2075 5234
rect 1962 5221 1992 5224
rect 1971 5217 1978 5221
rect 1978 5216 1979 5217
rect 1937 5210 1947 5216
rect 1696 5202 1731 5210
rect 1696 5176 1697 5202
rect 1704 5176 1731 5202
rect 1639 5158 1669 5172
rect 1696 5168 1731 5176
rect 1733 5202 1774 5210
rect 1733 5176 1748 5202
rect 1755 5176 1774 5202
rect 1838 5198 1869 5210
rect 1884 5198 1987 5210
rect 1999 5200 2025 5226
rect 2040 5221 2070 5232
rect 2102 5228 2164 5244
rect 2102 5226 2148 5228
rect 2102 5210 2164 5226
rect 2176 5210 2182 5258
rect 2185 5250 2265 5258
rect 2185 5248 2204 5250
rect 2219 5248 2253 5250
rect 2185 5232 2265 5248
rect 2185 5210 2204 5232
rect 2219 5216 2249 5232
rect 2277 5226 2283 5300
rect 2286 5226 2305 5370
rect 2320 5226 2326 5370
rect 2335 5300 2348 5370
rect 2400 5366 2422 5370
rect 2393 5344 2422 5358
rect 2475 5344 2491 5358
rect 2529 5354 2535 5356
rect 2542 5354 2650 5370
rect 2657 5354 2663 5356
rect 2671 5354 2686 5370
rect 2752 5364 2771 5367
rect 2393 5342 2491 5344
rect 2518 5342 2686 5354
rect 2701 5344 2717 5358
rect 2752 5345 2774 5364
rect 2784 5358 2800 5359
rect 2783 5356 2800 5358
rect 2784 5351 2800 5356
rect 2774 5344 2780 5345
rect 2783 5344 2812 5351
rect 2701 5343 2812 5344
rect 2701 5342 2818 5343
rect 2377 5334 2428 5342
rect 2475 5334 2509 5342
rect 2377 5322 2402 5334
rect 2409 5322 2428 5334
rect 2482 5332 2509 5334
rect 2518 5332 2739 5342
rect 2774 5339 2780 5342
rect 2482 5328 2739 5332
rect 2377 5314 2428 5322
rect 2475 5314 2739 5328
rect 2783 5334 2818 5342
rect 2329 5266 2348 5300
rect 2393 5306 2422 5314
rect 2393 5300 2410 5306
rect 2393 5298 2427 5300
rect 2475 5298 2491 5314
rect 2492 5304 2700 5314
rect 2701 5304 2717 5314
rect 2765 5310 2780 5325
rect 2783 5322 2784 5334
rect 2791 5322 2818 5334
rect 2783 5314 2818 5322
rect 2783 5313 2812 5314
rect 2503 5300 2717 5304
rect 2518 5298 2717 5300
rect 2752 5300 2765 5310
rect 2783 5300 2800 5313
rect 2752 5298 2800 5300
rect 2394 5294 2427 5298
rect 2390 5292 2427 5294
rect 2390 5291 2457 5292
rect 2390 5286 2421 5291
rect 2427 5286 2457 5291
rect 2390 5282 2457 5286
rect 2363 5279 2457 5282
rect 2363 5272 2412 5279
rect 2363 5266 2393 5272
rect 2412 5267 2417 5272
rect 2329 5250 2409 5266
rect 2421 5258 2457 5279
rect 2518 5274 2707 5298
rect 2752 5297 2799 5298
rect 2765 5292 2799 5297
rect 2533 5271 2707 5274
rect 2526 5268 2707 5271
rect 2735 5291 2799 5292
rect 2329 5248 2348 5250
rect 2363 5248 2397 5250
rect 2329 5232 2409 5248
rect 2329 5226 2348 5232
rect 2045 5200 2148 5210
rect 1999 5198 2148 5200
rect 2169 5198 2204 5210
rect 1838 5196 2000 5198
rect 1850 5176 1869 5196
rect 1884 5194 1914 5196
rect 1733 5168 1774 5176
rect 1856 5172 1869 5176
rect 1921 5180 2000 5196
rect 2032 5196 2204 5198
rect 2032 5180 2111 5196
rect 2118 5194 2148 5196
rect 1696 5158 1725 5168
rect 1739 5158 1768 5168
rect 1783 5158 1813 5172
rect 1856 5158 1899 5172
rect 1921 5168 2111 5180
rect 2176 5176 2182 5196
rect 1906 5158 1936 5168
rect 1937 5158 2095 5168
rect 2099 5158 2129 5168
rect 2133 5158 2163 5172
rect 2191 5158 2204 5196
rect 2276 5210 2305 5226
rect 2319 5210 2348 5226
rect 2363 5216 2393 5232
rect 2421 5210 2427 5258
rect 2430 5252 2449 5258
rect 2464 5252 2494 5260
rect 2430 5244 2494 5252
rect 2430 5228 2510 5244
rect 2526 5237 2588 5268
rect 2604 5237 2666 5268
rect 2735 5266 2784 5291
rect 2799 5266 2829 5282
rect 2698 5252 2728 5260
rect 2735 5258 2845 5266
rect 2698 5244 2743 5252
rect 2430 5226 2449 5228
rect 2464 5226 2510 5228
rect 2430 5210 2510 5226
rect 2537 5224 2572 5237
rect 2613 5234 2650 5237
rect 2613 5232 2655 5234
rect 2542 5221 2572 5224
rect 2551 5217 2558 5221
rect 2558 5216 2559 5217
rect 2517 5210 2527 5216
rect 2276 5202 2311 5210
rect 2276 5176 2277 5202
rect 2284 5176 2311 5202
rect 2219 5158 2249 5172
rect 2276 5168 2311 5176
rect 2313 5202 2354 5210
rect 2313 5176 2328 5202
rect 2335 5176 2354 5202
rect 2418 5198 2449 5210
rect 2464 5198 2567 5210
rect 2579 5200 2605 5226
rect 2620 5221 2650 5232
rect 2682 5228 2744 5244
rect 2682 5226 2728 5228
rect 2682 5210 2744 5226
rect 2756 5210 2762 5258
rect 2765 5250 2845 5258
rect 2765 5248 2784 5250
rect 2799 5248 2833 5250
rect 2765 5232 2845 5248
rect 2765 5210 2784 5232
rect 2799 5216 2829 5232
rect 2857 5226 2863 5300
rect 2866 5226 2885 5370
rect 2900 5226 2906 5370
rect 2915 5300 2928 5370
rect 2980 5366 3002 5370
rect 2973 5344 3002 5358
rect 3055 5344 3071 5358
rect 3109 5354 3115 5356
rect 3122 5354 3230 5370
rect 3237 5354 3243 5356
rect 3251 5354 3266 5370
rect 3332 5364 3351 5367
rect 2973 5342 3071 5344
rect 3098 5342 3266 5354
rect 3281 5344 3297 5358
rect 3332 5345 3354 5364
rect 3364 5358 3380 5359
rect 3363 5356 3380 5358
rect 3364 5351 3380 5356
rect 3354 5344 3360 5345
rect 3363 5344 3392 5351
rect 3281 5343 3392 5344
rect 3281 5342 3398 5343
rect 2957 5334 3008 5342
rect 3055 5334 3089 5342
rect 2957 5322 2982 5334
rect 2989 5322 3008 5334
rect 3062 5332 3089 5334
rect 3098 5332 3319 5342
rect 3354 5339 3360 5342
rect 3062 5328 3319 5332
rect 2957 5314 3008 5322
rect 3055 5314 3319 5328
rect 3363 5334 3398 5342
rect 2909 5266 2928 5300
rect 2973 5306 3002 5314
rect 2973 5300 2990 5306
rect 2973 5298 3007 5300
rect 3055 5298 3071 5314
rect 3072 5304 3280 5314
rect 3281 5304 3297 5314
rect 3345 5310 3360 5325
rect 3363 5322 3364 5334
rect 3371 5322 3398 5334
rect 3363 5314 3398 5322
rect 3363 5313 3392 5314
rect 3083 5300 3297 5304
rect 3098 5298 3297 5300
rect 3332 5300 3345 5310
rect 3363 5300 3380 5313
rect 3332 5298 3380 5300
rect 2974 5294 3007 5298
rect 2970 5292 3007 5294
rect 2970 5291 3037 5292
rect 2970 5286 3001 5291
rect 3007 5286 3037 5291
rect 2970 5282 3037 5286
rect 2943 5279 3037 5282
rect 2943 5272 2992 5279
rect 2943 5266 2973 5272
rect 2992 5267 2997 5272
rect 2909 5250 2989 5266
rect 3001 5258 3037 5279
rect 3098 5274 3287 5298
rect 3332 5297 3379 5298
rect 3345 5292 3379 5297
rect 3113 5271 3287 5274
rect 3106 5268 3287 5271
rect 3315 5291 3379 5292
rect 2909 5248 2928 5250
rect 2943 5248 2977 5250
rect 2909 5232 2989 5248
rect 2909 5226 2928 5232
rect 2625 5200 2728 5210
rect 2579 5198 2728 5200
rect 2749 5198 2784 5210
rect 2418 5196 2580 5198
rect 2430 5176 2449 5196
rect 2464 5194 2494 5196
rect 2313 5168 2354 5176
rect 2436 5172 2449 5176
rect 2501 5180 2580 5196
rect 2612 5196 2784 5198
rect 2612 5180 2691 5196
rect 2698 5194 2728 5196
rect 2276 5158 2305 5168
rect 2319 5158 2348 5168
rect 2363 5158 2393 5172
rect 2436 5158 2479 5172
rect 2501 5168 2691 5180
rect 2756 5176 2762 5196
rect 2486 5158 2516 5168
rect 2517 5158 2675 5168
rect 2679 5158 2709 5168
rect 2713 5158 2743 5172
rect 2771 5158 2784 5196
rect 2856 5210 2885 5226
rect 2899 5210 2928 5226
rect 2943 5216 2973 5232
rect 3001 5210 3007 5258
rect 3010 5252 3029 5258
rect 3044 5252 3074 5260
rect 3010 5244 3074 5252
rect 3010 5228 3090 5244
rect 3106 5237 3168 5268
rect 3184 5237 3246 5268
rect 3315 5266 3364 5291
rect 3379 5266 3409 5282
rect 3278 5252 3308 5260
rect 3315 5258 3425 5266
rect 3278 5244 3323 5252
rect 3010 5226 3029 5228
rect 3044 5226 3090 5228
rect 3010 5210 3090 5226
rect 3117 5224 3152 5237
rect 3193 5234 3230 5237
rect 3193 5232 3235 5234
rect 3122 5221 3152 5224
rect 3131 5217 3138 5221
rect 3138 5216 3139 5217
rect 3097 5210 3107 5216
rect 2856 5202 2891 5210
rect 2856 5176 2857 5202
rect 2864 5176 2891 5202
rect 2799 5158 2829 5172
rect 2856 5168 2891 5176
rect 2893 5202 2934 5210
rect 2893 5176 2908 5202
rect 2915 5176 2934 5202
rect 2998 5198 3029 5210
rect 3044 5198 3147 5210
rect 3159 5200 3185 5226
rect 3200 5221 3230 5232
rect 3262 5228 3324 5244
rect 3262 5226 3308 5228
rect 3262 5210 3324 5226
rect 3336 5210 3342 5258
rect 3345 5250 3425 5258
rect 3345 5248 3364 5250
rect 3379 5248 3413 5250
rect 3345 5232 3425 5248
rect 3345 5210 3364 5232
rect 3379 5216 3409 5232
rect 3437 5226 3443 5300
rect 3446 5226 3465 5370
rect 3480 5226 3486 5370
rect 3495 5300 3508 5370
rect 3560 5366 3582 5370
rect 3553 5344 3582 5358
rect 3635 5344 3651 5358
rect 3689 5354 3695 5356
rect 3702 5354 3810 5370
rect 3817 5354 3823 5356
rect 3831 5354 3846 5370
rect 3912 5364 3931 5367
rect 3553 5342 3651 5344
rect 3678 5342 3846 5354
rect 3861 5344 3877 5358
rect 3912 5345 3934 5364
rect 3944 5358 3960 5359
rect 3943 5356 3960 5358
rect 3944 5351 3960 5356
rect 3934 5344 3940 5345
rect 3943 5344 3972 5351
rect 3861 5343 3972 5344
rect 3861 5342 3978 5343
rect 3537 5334 3588 5342
rect 3635 5334 3669 5342
rect 3537 5322 3562 5334
rect 3569 5322 3588 5334
rect 3642 5332 3669 5334
rect 3678 5332 3899 5342
rect 3934 5339 3940 5342
rect 3642 5328 3899 5332
rect 3537 5314 3588 5322
rect 3635 5314 3899 5328
rect 3943 5334 3978 5342
rect 3489 5266 3508 5300
rect 3553 5306 3582 5314
rect 3553 5300 3570 5306
rect 3553 5298 3587 5300
rect 3635 5298 3651 5314
rect 3652 5304 3860 5314
rect 3861 5304 3877 5314
rect 3925 5310 3940 5325
rect 3943 5322 3944 5334
rect 3951 5322 3978 5334
rect 3943 5314 3978 5322
rect 3943 5313 3972 5314
rect 3663 5300 3877 5304
rect 3678 5298 3877 5300
rect 3912 5300 3925 5310
rect 3943 5300 3960 5313
rect 3912 5298 3960 5300
rect 3554 5294 3587 5298
rect 3550 5292 3587 5294
rect 3550 5291 3617 5292
rect 3550 5286 3581 5291
rect 3587 5286 3617 5291
rect 3550 5282 3617 5286
rect 3523 5279 3617 5282
rect 3523 5272 3572 5279
rect 3523 5266 3553 5272
rect 3572 5267 3577 5272
rect 3489 5250 3569 5266
rect 3581 5258 3617 5279
rect 3678 5274 3867 5298
rect 3912 5297 3959 5298
rect 3925 5292 3959 5297
rect 3693 5271 3867 5274
rect 3686 5268 3867 5271
rect 3895 5291 3959 5292
rect 3489 5248 3508 5250
rect 3523 5248 3557 5250
rect 3489 5232 3569 5248
rect 3489 5226 3508 5232
rect 3205 5200 3308 5210
rect 3159 5198 3308 5200
rect 3329 5198 3364 5210
rect 2998 5196 3160 5198
rect 3010 5176 3029 5196
rect 3044 5194 3074 5196
rect 2893 5168 2934 5176
rect 3016 5172 3029 5176
rect 3081 5180 3160 5196
rect 3192 5196 3364 5198
rect 3192 5180 3271 5196
rect 3278 5194 3308 5196
rect 2856 5158 2885 5168
rect 2899 5158 2928 5168
rect 2943 5158 2973 5172
rect 3016 5158 3059 5172
rect 3081 5168 3271 5180
rect 3336 5176 3342 5196
rect 3066 5158 3096 5168
rect 3097 5158 3255 5168
rect 3259 5158 3289 5168
rect 3293 5158 3323 5172
rect 3351 5158 3364 5196
rect 3436 5210 3465 5226
rect 3479 5210 3508 5226
rect 3523 5216 3553 5232
rect 3581 5210 3587 5258
rect 3590 5252 3609 5258
rect 3624 5252 3654 5260
rect 3590 5244 3654 5252
rect 3590 5228 3670 5244
rect 3686 5237 3748 5268
rect 3764 5237 3826 5268
rect 3895 5266 3944 5291
rect 3959 5266 3989 5282
rect 3858 5252 3888 5260
rect 3895 5258 4005 5266
rect 3858 5244 3903 5252
rect 3590 5226 3609 5228
rect 3624 5226 3670 5228
rect 3590 5210 3670 5226
rect 3697 5224 3732 5237
rect 3773 5234 3810 5237
rect 3773 5232 3815 5234
rect 3702 5221 3732 5224
rect 3711 5217 3718 5221
rect 3718 5216 3719 5217
rect 3677 5210 3687 5216
rect 3436 5202 3471 5210
rect 3436 5176 3437 5202
rect 3444 5176 3471 5202
rect 3379 5158 3409 5172
rect 3436 5168 3471 5176
rect 3473 5202 3514 5210
rect 3473 5176 3488 5202
rect 3495 5176 3514 5202
rect 3578 5198 3609 5210
rect 3624 5198 3727 5210
rect 3739 5200 3765 5226
rect 3780 5221 3810 5232
rect 3842 5228 3904 5244
rect 3842 5226 3888 5228
rect 3842 5210 3904 5226
rect 3916 5210 3922 5258
rect 3925 5250 4005 5258
rect 3925 5248 3944 5250
rect 3959 5248 3993 5250
rect 3925 5232 4005 5248
rect 3925 5210 3944 5232
rect 3959 5216 3989 5232
rect 4017 5226 4023 5300
rect 4026 5226 4045 5370
rect 4060 5226 4066 5370
rect 4075 5300 4088 5370
rect 4140 5366 4162 5370
rect 4133 5344 4162 5358
rect 4215 5344 4231 5358
rect 4269 5354 4275 5356
rect 4282 5354 4390 5370
rect 4397 5354 4403 5356
rect 4411 5354 4426 5370
rect 4492 5364 4511 5367
rect 4133 5342 4231 5344
rect 4258 5342 4426 5354
rect 4441 5344 4457 5358
rect 4492 5345 4514 5364
rect 4524 5358 4540 5359
rect 4523 5356 4540 5358
rect 4524 5351 4540 5356
rect 4514 5344 4520 5345
rect 4523 5344 4552 5351
rect 4441 5343 4552 5344
rect 4441 5342 4558 5343
rect 4117 5334 4168 5342
rect 4215 5334 4249 5342
rect 4117 5322 4142 5334
rect 4149 5322 4168 5334
rect 4222 5332 4249 5334
rect 4258 5332 4479 5342
rect 4514 5339 4520 5342
rect 4222 5328 4479 5332
rect 4117 5314 4168 5322
rect 4215 5314 4479 5328
rect 4523 5334 4558 5342
rect 4069 5266 4088 5300
rect 4133 5306 4162 5314
rect 4133 5300 4150 5306
rect 4133 5298 4167 5300
rect 4215 5298 4231 5314
rect 4232 5304 4440 5314
rect 4441 5304 4457 5314
rect 4505 5310 4520 5325
rect 4523 5322 4524 5334
rect 4531 5322 4558 5334
rect 4523 5314 4558 5322
rect 4523 5313 4552 5314
rect 4243 5300 4457 5304
rect 4258 5298 4457 5300
rect 4492 5300 4505 5310
rect 4523 5300 4540 5313
rect 4492 5298 4540 5300
rect 4134 5294 4167 5298
rect 4130 5292 4167 5294
rect 4130 5291 4197 5292
rect 4130 5286 4161 5291
rect 4167 5286 4197 5291
rect 4130 5282 4197 5286
rect 4103 5279 4197 5282
rect 4103 5272 4152 5279
rect 4103 5266 4133 5272
rect 4152 5267 4157 5272
rect 4069 5250 4149 5266
rect 4161 5258 4197 5279
rect 4258 5274 4447 5298
rect 4492 5297 4539 5298
rect 4505 5292 4539 5297
rect 4273 5271 4447 5274
rect 4266 5268 4447 5271
rect 4475 5291 4539 5292
rect 4069 5248 4088 5250
rect 4103 5248 4137 5250
rect 4069 5232 4149 5248
rect 4069 5226 4088 5232
rect 3785 5200 3888 5210
rect 3739 5198 3888 5200
rect 3909 5198 3944 5210
rect 3578 5196 3740 5198
rect 3590 5176 3609 5196
rect 3624 5194 3654 5196
rect 3473 5168 3514 5176
rect 3596 5172 3609 5176
rect 3661 5180 3740 5196
rect 3772 5196 3944 5198
rect 3772 5180 3851 5196
rect 3858 5194 3888 5196
rect 3436 5158 3465 5168
rect 3479 5158 3508 5168
rect 3523 5158 3553 5172
rect 3596 5158 3639 5172
rect 3661 5168 3851 5180
rect 3916 5176 3922 5196
rect 3646 5158 3676 5168
rect 3677 5158 3835 5168
rect 3839 5158 3869 5168
rect 3873 5158 3903 5172
rect 3931 5158 3944 5196
rect 4016 5210 4045 5226
rect 4059 5210 4088 5226
rect 4103 5216 4133 5232
rect 4161 5210 4167 5258
rect 4170 5252 4189 5258
rect 4204 5252 4234 5260
rect 4170 5244 4234 5252
rect 4170 5228 4250 5244
rect 4266 5237 4328 5268
rect 4344 5237 4406 5268
rect 4475 5266 4524 5291
rect 4539 5266 4569 5282
rect 4438 5252 4468 5260
rect 4475 5258 4585 5266
rect 4438 5244 4483 5252
rect 4170 5226 4189 5228
rect 4204 5226 4250 5228
rect 4170 5210 4250 5226
rect 4277 5224 4312 5237
rect 4353 5234 4390 5237
rect 4353 5232 4395 5234
rect 4282 5221 4312 5224
rect 4291 5217 4298 5221
rect 4298 5216 4299 5217
rect 4257 5210 4267 5216
rect 4016 5202 4051 5210
rect 4016 5176 4017 5202
rect 4024 5176 4051 5202
rect 3959 5158 3989 5172
rect 4016 5168 4051 5176
rect 4053 5202 4094 5210
rect 4053 5176 4068 5202
rect 4075 5176 4094 5202
rect 4158 5198 4189 5210
rect 4204 5198 4307 5210
rect 4319 5200 4345 5226
rect 4360 5221 4390 5232
rect 4422 5228 4484 5244
rect 4422 5226 4468 5228
rect 4422 5210 4484 5226
rect 4496 5210 4502 5258
rect 4505 5250 4585 5258
rect 4505 5248 4524 5250
rect 4539 5248 4573 5250
rect 4505 5232 4585 5248
rect 4505 5210 4524 5232
rect 4539 5216 4569 5232
rect 4597 5226 4603 5300
rect 4606 5226 4625 5370
rect 4640 5226 4646 5370
rect 4655 5300 4668 5370
rect 4720 5366 4742 5370
rect 4713 5344 4742 5358
rect 4795 5344 4811 5358
rect 4849 5354 4855 5356
rect 4862 5354 4970 5370
rect 4977 5354 4983 5356
rect 4991 5354 5006 5370
rect 5072 5364 5091 5367
rect 4713 5342 4811 5344
rect 4838 5342 5006 5354
rect 5021 5344 5037 5358
rect 5072 5345 5094 5364
rect 5104 5358 5120 5359
rect 5103 5356 5120 5358
rect 5104 5351 5120 5356
rect 5094 5344 5100 5345
rect 5103 5344 5132 5351
rect 5021 5343 5132 5344
rect 5021 5342 5138 5343
rect 4697 5334 4748 5342
rect 4795 5334 4829 5342
rect 4697 5322 4722 5334
rect 4729 5322 4748 5334
rect 4802 5332 4829 5334
rect 4838 5332 5059 5342
rect 5094 5339 5100 5342
rect 4802 5328 5059 5332
rect 4697 5314 4748 5322
rect 4795 5314 5059 5328
rect 5103 5334 5138 5342
rect 4649 5266 4668 5300
rect 4713 5306 4742 5314
rect 4713 5300 4730 5306
rect 4713 5298 4747 5300
rect 4795 5298 4811 5314
rect 4812 5304 5020 5314
rect 5021 5304 5037 5314
rect 5085 5310 5100 5325
rect 5103 5322 5104 5334
rect 5111 5322 5138 5334
rect 5103 5314 5138 5322
rect 5103 5313 5132 5314
rect 4823 5300 5037 5304
rect 4838 5298 5037 5300
rect 5072 5300 5085 5310
rect 5103 5300 5120 5313
rect 5072 5298 5120 5300
rect 4714 5294 4747 5298
rect 4710 5292 4747 5294
rect 4710 5291 4777 5292
rect 4710 5286 4741 5291
rect 4747 5286 4777 5291
rect 4710 5282 4777 5286
rect 4683 5279 4777 5282
rect 4683 5272 4732 5279
rect 4683 5266 4713 5272
rect 4732 5267 4737 5272
rect 4649 5250 4729 5266
rect 4741 5258 4777 5279
rect 4838 5274 5027 5298
rect 5072 5297 5119 5298
rect 5085 5292 5119 5297
rect 4853 5271 5027 5274
rect 4846 5268 5027 5271
rect 5055 5291 5119 5292
rect 4649 5248 4668 5250
rect 4683 5248 4717 5250
rect 4649 5232 4729 5248
rect 4649 5226 4668 5232
rect 4365 5200 4468 5210
rect 4319 5198 4468 5200
rect 4489 5198 4524 5210
rect 4158 5196 4320 5198
rect 4170 5176 4189 5196
rect 4204 5194 4234 5196
rect 4053 5168 4094 5176
rect 4176 5172 4189 5176
rect 4241 5180 4320 5196
rect 4352 5196 4524 5198
rect 4352 5180 4431 5196
rect 4438 5194 4468 5196
rect 4016 5158 4045 5168
rect 4059 5158 4088 5168
rect 4103 5158 4133 5172
rect 4176 5158 4219 5172
rect 4241 5168 4431 5180
rect 4496 5176 4502 5196
rect 4226 5158 4256 5168
rect 4257 5158 4415 5168
rect 4419 5158 4449 5168
rect 4453 5158 4483 5172
rect 4511 5158 4524 5196
rect 4596 5210 4625 5226
rect 4639 5210 4668 5226
rect 4683 5216 4713 5232
rect 4741 5210 4747 5258
rect 4750 5252 4769 5258
rect 4784 5252 4814 5260
rect 4750 5244 4814 5252
rect 4750 5228 4830 5244
rect 4846 5237 4908 5268
rect 4924 5237 4986 5268
rect 5055 5266 5104 5291
rect 5119 5266 5149 5282
rect 5018 5252 5048 5260
rect 5055 5258 5165 5266
rect 5018 5244 5063 5252
rect 4750 5226 4769 5228
rect 4784 5226 4830 5228
rect 4750 5210 4830 5226
rect 4857 5224 4892 5237
rect 4933 5234 4970 5237
rect 4933 5232 4975 5234
rect 4862 5221 4892 5224
rect 4871 5217 4878 5221
rect 4878 5216 4879 5217
rect 4837 5210 4847 5216
rect 4596 5202 4631 5210
rect 4596 5176 4597 5202
rect 4604 5176 4631 5202
rect 4539 5158 4569 5172
rect 4596 5168 4631 5176
rect 4633 5202 4674 5210
rect 4633 5176 4648 5202
rect 4655 5176 4674 5202
rect 4738 5198 4769 5210
rect 4784 5198 4887 5210
rect 4899 5200 4925 5226
rect 4940 5221 4970 5232
rect 5002 5228 5064 5244
rect 5002 5226 5048 5228
rect 5002 5210 5064 5226
rect 5076 5210 5082 5258
rect 5085 5250 5165 5258
rect 5085 5248 5104 5250
rect 5119 5248 5153 5250
rect 5085 5232 5165 5248
rect 5085 5210 5104 5232
rect 5119 5216 5149 5232
rect 5177 5226 5183 5300
rect 5186 5226 5205 5370
rect 5220 5226 5226 5370
rect 5235 5300 5248 5370
rect 5300 5366 5322 5370
rect 5293 5344 5322 5358
rect 5375 5344 5391 5358
rect 5429 5354 5435 5356
rect 5442 5354 5550 5370
rect 5557 5354 5563 5356
rect 5571 5354 5586 5370
rect 5652 5364 5671 5367
rect 5293 5342 5391 5344
rect 5418 5342 5586 5354
rect 5601 5344 5617 5358
rect 5652 5345 5674 5364
rect 5684 5358 5700 5359
rect 5683 5356 5700 5358
rect 5684 5351 5700 5356
rect 5674 5344 5680 5345
rect 5683 5344 5712 5351
rect 5601 5343 5712 5344
rect 5601 5342 5718 5343
rect 5277 5334 5328 5342
rect 5375 5334 5409 5342
rect 5277 5322 5302 5334
rect 5309 5322 5328 5334
rect 5382 5332 5409 5334
rect 5418 5332 5639 5342
rect 5674 5339 5680 5342
rect 5382 5328 5639 5332
rect 5277 5314 5328 5322
rect 5375 5314 5639 5328
rect 5683 5334 5718 5342
rect 5229 5266 5248 5300
rect 5293 5306 5322 5314
rect 5293 5300 5310 5306
rect 5293 5298 5327 5300
rect 5375 5298 5391 5314
rect 5392 5304 5600 5314
rect 5601 5304 5617 5314
rect 5665 5310 5680 5325
rect 5683 5322 5684 5334
rect 5691 5322 5718 5334
rect 5683 5314 5718 5322
rect 5683 5313 5712 5314
rect 5403 5300 5617 5304
rect 5418 5298 5617 5300
rect 5652 5300 5665 5310
rect 5683 5300 5700 5313
rect 5652 5298 5700 5300
rect 5294 5294 5327 5298
rect 5290 5292 5327 5294
rect 5290 5291 5357 5292
rect 5290 5286 5321 5291
rect 5327 5286 5357 5291
rect 5290 5282 5357 5286
rect 5263 5279 5357 5282
rect 5263 5272 5312 5279
rect 5263 5266 5293 5272
rect 5312 5267 5317 5272
rect 5229 5250 5309 5266
rect 5321 5258 5357 5279
rect 5418 5274 5607 5298
rect 5652 5297 5699 5298
rect 5665 5292 5699 5297
rect 5433 5271 5607 5274
rect 5426 5268 5607 5271
rect 5635 5291 5699 5292
rect 5229 5248 5248 5250
rect 5263 5248 5297 5250
rect 5229 5232 5309 5248
rect 5229 5226 5248 5232
rect 4945 5200 5048 5210
rect 4899 5198 5048 5200
rect 5069 5198 5104 5210
rect 4738 5196 4900 5198
rect 4750 5176 4769 5196
rect 4784 5194 4814 5196
rect 4633 5168 4674 5176
rect 4756 5172 4769 5176
rect 4821 5180 4900 5196
rect 4932 5196 5104 5198
rect 4932 5180 5011 5196
rect 5018 5194 5048 5196
rect 4596 5158 4625 5168
rect 4639 5158 4668 5168
rect 4683 5158 4713 5172
rect 4756 5158 4799 5172
rect 4821 5168 5011 5180
rect 5076 5176 5082 5196
rect 4806 5158 4836 5168
rect 4837 5158 4995 5168
rect 4999 5158 5029 5168
rect 5033 5158 5063 5172
rect 5091 5158 5104 5196
rect 5176 5210 5205 5226
rect 5219 5210 5248 5226
rect 5263 5216 5293 5232
rect 5321 5210 5327 5258
rect 5330 5252 5349 5258
rect 5364 5252 5394 5260
rect 5330 5244 5394 5252
rect 5330 5228 5410 5244
rect 5426 5237 5488 5268
rect 5504 5237 5566 5268
rect 5635 5266 5684 5291
rect 5699 5266 5729 5282
rect 5598 5252 5628 5260
rect 5635 5258 5745 5266
rect 5598 5244 5643 5252
rect 5330 5226 5349 5228
rect 5364 5226 5410 5228
rect 5330 5210 5410 5226
rect 5437 5224 5472 5237
rect 5513 5234 5550 5237
rect 5513 5232 5555 5234
rect 5442 5221 5472 5224
rect 5451 5217 5458 5221
rect 5458 5216 5459 5217
rect 5417 5210 5427 5216
rect 5176 5202 5211 5210
rect 5176 5176 5177 5202
rect 5184 5176 5211 5202
rect 5119 5158 5149 5172
rect 5176 5168 5211 5176
rect 5213 5202 5254 5210
rect 5213 5176 5228 5202
rect 5235 5176 5254 5202
rect 5318 5198 5349 5210
rect 5364 5198 5467 5210
rect 5479 5200 5505 5226
rect 5520 5221 5550 5232
rect 5582 5228 5644 5244
rect 5582 5226 5628 5228
rect 5582 5210 5644 5226
rect 5656 5210 5662 5258
rect 5665 5250 5745 5258
rect 5665 5248 5684 5250
rect 5699 5248 5733 5250
rect 5665 5232 5745 5248
rect 5665 5210 5684 5232
rect 5699 5216 5729 5232
rect 5757 5226 5763 5300
rect 5766 5226 5785 5370
rect 5800 5226 5806 5370
rect 5815 5300 5828 5370
rect 5880 5366 5902 5370
rect 5873 5344 5902 5358
rect 5955 5344 5971 5358
rect 6009 5354 6015 5356
rect 6022 5354 6130 5370
rect 6137 5354 6143 5356
rect 6151 5354 6166 5370
rect 6232 5364 6251 5367
rect 5873 5342 5971 5344
rect 5998 5342 6166 5354
rect 6181 5344 6197 5358
rect 6232 5345 6254 5364
rect 6264 5358 6280 5359
rect 6263 5356 6280 5358
rect 6264 5351 6280 5356
rect 6254 5344 6260 5345
rect 6263 5344 6292 5351
rect 6181 5343 6292 5344
rect 6181 5342 6298 5343
rect 5857 5334 5908 5342
rect 5955 5334 5989 5342
rect 5857 5322 5882 5334
rect 5889 5322 5908 5334
rect 5962 5332 5989 5334
rect 5998 5332 6219 5342
rect 6254 5339 6260 5342
rect 5962 5328 6219 5332
rect 5857 5314 5908 5322
rect 5955 5314 6219 5328
rect 6263 5334 6298 5342
rect 5809 5266 5828 5300
rect 5873 5306 5902 5314
rect 5873 5300 5890 5306
rect 5873 5298 5907 5300
rect 5955 5298 5971 5314
rect 5972 5304 6180 5314
rect 6181 5304 6197 5314
rect 6245 5310 6260 5325
rect 6263 5322 6264 5334
rect 6271 5322 6298 5334
rect 6263 5314 6298 5322
rect 6263 5313 6292 5314
rect 5983 5300 6197 5304
rect 5998 5298 6197 5300
rect 6232 5300 6245 5310
rect 6263 5300 6280 5313
rect 6232 5298 6280 5300
rect 5874 5294 5907 5298
rect 5870 5292 5907 5294
rect 5870 5291 5937 5292
rect 5870 5286 5901 5291
rect 5907 5286 5937 5291
rect 5870 5282 5937 5286
rect 5843 5279 5937 5282
rect 5843 5272 5892 5279
rect 5843 5266 5873 5272
rect 5892 5267 5897 5272
rect 5809 5250 5889 5266
rect 5901 5258 5937 5279
rect 5998 5274 6187 5298
rect 6232 5297 6279 5298
rect 6245 5292 6279 5297
rect 6013 5271 6187 5274
rect 6006 5268 6187 5271
rect 6215 5291 6279 5292
rect 5809 5248 5828 5250
rect 5843 5248 5877 5250
rect 5809 5232 5889 5248
rect 5809 5226 5828 5232
rect 5525 5200 5628 5210
rect 5479 5198 5628 5200
rect 5649 5198 5684 5210
rect 5318 5196 5480 5198
rect 5330 5176 5349 5196
rect 5364 5194 5394 5196
rect 5213 5168 5254 5176
rect 5336 5172 5349 5176
rect 5401 5180 5480 5196
rect 5512 5196 5684 5198
rect 5512 5180 5591 5196
rect 5598 5194 5628 5196
rect 5176 5158 5205 5168
rect 5219 5158 5248 5168
rect 5263 5158 5293 5172
rect 5336 5158 5379 5172
rect 5401 5168 5591 5180
rect 5656 5176 5662 5196
rect 5386 5158 5416 5168
rect 5417 5158 5575 5168
rect 5579 5158 5609 5168
rect 5613 5158 5643 5172
rect 5671 5158 5684 5196
rect 5756 5210 5785 5226
rect 5799 5210 5828 5226
rect 5843 5216 5873 5232
rect 5901 5210 5907 5258
rect 5910 5252 5929 5258
rect 5944 5252 5974 5260
rect 5910 5244 5974 5252
rect 5910 5228 5990 5244
rect 6006 5237 6068 5268
rect 6084 5237 6146 5268
rect 6215 5266 6264 5291
rect 6279 5266 6309 5282
rect 6178 5252 6208 5260
rect 6215 5258 6325 5266
rect 6178 5244 6223 5252
rect 5910 5226 5929 5228
rect 5944 5226 5990 5228
rect 5910 5210 5990 5226
rect 6017 5224 6052 5237
rect 6093 5234 6130 5237
rect 6093 5232 6135 5234
rect 6022 5221 6052 5224
rect 6031 5217 6038 5221
rect 6038 5216 6039 5217
rect 5997 5210 6007 5216
rect 5756 5202 5791 5210
rect 5756 5176 5757 5202
rect 5764 5176 5791 5202
rect 5699 5158 5729 5172
rect 5756 5168 5791 5176
rect 5793 5202 5834 5210
rect 5793 5176 5808 5202
rect 5815 5176 5834 5202
rect 5898 5198 5929 5210
rect 5944 5198 6047 5210
rect 6059 5200 6085 5226
rect 6100 5221 6130 5232
rect 6162 5228 6224 5244
rect 6162 5226 6208 5228
rect 6162 5210 6224 5226
rect 6236 5210 6242 5258
rect 6245 5250 6325 5258
rect 6245 5248 6264 5250
rect 6279 5248 6313 5250
rect 6245 5232 6325 5248
rect 6245 5210 6264 5232
rect 6279 5216 6309 5232
rect 6337 5226 6343 5300
rect 6346 5226 6365 5370
rect 6380 5226 6386 5370
rect 6395 5300 6408 5370
rect 6460 5366 6482 5370
rect 6453 5344 6482 5358
rect 6535 5344 6551 5358
rect 6589 5354 6595 5356
rect 6602 5354 6710 5370
rect 6717 5354 6723 5356
rect 6731 5354 6746 5370
rect 6812 5364 6831 5367
rect 6453 5342 6551 5344
rect 6578 5342 6746 5354
rect 6761 5344 6777 5358
rect 6812 5345 6834 5364
rect 6844 5358 6860 5359
rect 6843 5356 6860 5358
rect 6844 5351 6860 5356
rect 6834 5344 6840 5345
rect 6843 5344 6872 5351
rect 6761 5343 6872 5344
rect 6761 5342 6878 5343
rect 6437 5334 6488 5342
rect 6535 5334 6569 5342
rect 6437 5322 6462 5334
rect 6469 5322 6488 5334
rect 6542 5332 6569 5334
rect 6578 5332 6799 5342
rect 6834 5339 6840 5342
rect 6542 5328 6799 5332
rect 6437 5314 6488 5322
rect 6535 5314 6799 5328
rect 6843 5334 6878 5342
rect 6389 5266 6408 5300
rect 6453 5306 6482 5314
rect 6453 5300 6470 5306
rect 6453 5298 6487 5300
rect 6535 5298 6551 5314
rect 6552 5304 6760 5314
rect 6761 5304 6777 5314
rect 6825 5310 6840 5325
rect 6843 5322 6844 5334
rect 6851 5322 6878 5334
rect 6843 5314 6878 5322
rect 6843 5313 6872 5314
rect 6563 5300 6777 5304
rect 6578 5298 6777 5300
rect 6812 5300 6825 5310
rect 6843 5300 6860 5313
rect 6812 5298 6860 5300
rect 6454 5294 6487 5298
rect 6450 5292 6487 5294
rect 6450 5291 6517 5292
rect 6450 5286 6481 5291
rect 6487 5286 6517 5291
rect 6450 5282 6517 5286
rect 6423 5279 6517 5282
rect 6423 5272 6472 5279
rect 6423 5266 6453 5272
rect 6472 5267 6477 5272
rect 6389 5250 6469 5266
rect 6481 5258 6517 5279
rect 6578 5274 6767 5298
rect 6812 5297 6859 5298
rect 6825 5292 6859 5297
rect 6593 5271 6767 5274
rect 6586 5268 6767 5271
rect 6795 5291 6859 5292
rect 6389 5248 6408 5250
rect 6423 5248 6457 5250
rect 6389 5232 6469 5248
rect 6389 5226 6408 5232
rect 6105 5200 6208 5210
rect 6059 5198 6208 5200
rect 6229 5198 6264 5210
rect 5898 5196 6060 5198
rect 5910 5176 5929 5196
rect 5944 5194 5974 5196
rect 5793 5168 5834 5176
rect 5916 5172 5929 5176
rect 5981 5180 6060 5196
rect 6092 5196 6264 5198
rect 6092 5180 6171 5196
rect 6178 5194 6208 5196
rect 5756 5158 5785 5168
rect 5799 5158 5828 5168
rect 5843 5158 5873 5172
rect 5916 5158 5959 5172
rect 5981 5168 6171 5180
rect 6236 5176 6242 5196
rect 5966 5158 5996 5168
rect 5997 5158 6155 5168
rect 6159 5158 6189 5168
rect 6193 5158 6223 5172
rect 6251 5158 6264 5196
rect 6336 5210 6365 5226
rect 6379 5210 6408 5226
rect 6423 5216 6453 5232
rect 6481 5210 6487 5258
rect 6490 5252 6509 5258
rect 6524 5252 6554 5260
rect 6490 5244 6554 5252
rect 6490 5228 6570 5244
rect 6586 5237 6648 5268
rect 6664 5237 6726 5268
rect 6795 5266 6844 5291
rect 6859 5266 6889 5282
rect 6758 5252 6788 5260
rect 6795 5258 6905 5266
rect 6758 5244 6803 5252
rect 6490 5226 6509 5228
rect 6524 5226 6570 5228
rect 6490 5210 6570 5226
rect 6597 5224 6632 5237
rect 6673 5234 6710 5237
rect 6673 5232 6715 5234
rect 6602 5221 6632 5224
rect 6611 5217 6618 5221
rect 6618 5216 6619 5217
rect 6577 5210 6587 5216
rect 6336 5202 6371 5210
rect 6336 5176 6337 5202
rect 6344 5176 6371 5202
rect 6279 5158 6309 5172
rect 6336 5168 6371 5176
rect 6373 5202 6414 5210
rect 6373 5176 6388 5202
rect 6395 5176 6414 5202
rect 6478 5198 6509 5210
rect 6524 5198 6627 5210
rect 6639 5200 6665 5226
rect 6680 5221 6710 5232
rect 6742 5228 6804 5244
rect 6742 5226 6788 5228
rect 6742 5210 6804 5226
rect 6816 5210 6822 5258
rect 6825 5250 6905 5258
rect 6825 5248 6844 5250
rect 6859 5248 6893 5250
rect 6825 5232 6905 5248
rect 6825 5210 6844 5232
rect 6859 5216 6889 5232
rect 6917 5226 6923 5300
rect 6926 5226 6945 5370
rect 6960 5226 6966 5370
rect 6975 5300 6988 5370
rect 7040 5366 7062 5370
rect 7033 5344 7062 5358
rect 7115 5344 7131 5358
rect 7169 5354 7175 5356
rect 7182 5354 7290 5370
rect 7297 5354 7303 5356
rect 7311 5354 7326 5370
rect 7392 5364 7411 5367
rect 7033 5342 7131 5344
rect 7158 5342 7326 5354
rect 7341 5344 7357 5358
rect 7392 5345 7414 5364
rect 7424 5358 7440 5359
rect 7423 5356 7440 5358
rect 7424 5351 7440 5356
rect 7414 5344 7420 5345
rect 7423 5344 7452 5351
rect 7341 5343 7452 5344
rect 7341 5342 7458 5343
rect 7017 5334 7068 5342
rect 7115 5334 7149 5342
rect 7017 5322 7042 5334
rect 7049 5322 7068 5334
rect 7122 5332 7149 5334
rect 7158 5332 7379 5342
rect 7414 5339 7420 5342
rect 7122 5328 7379 5332
rect 7017 5314 7068 5322
rect 7115 5314 7379 5328
rect 7423 5334 7458 5342
rect 6969 5266 6988 5300
rect 7033 5306 7062 5314
rect 7033 5300 7050 5306
rect 7033 5298 7067 5300
rect 7115 5298 7131 5314
rect 7132 5304 7340 5314
rect 7341 5304 7357 5314
rect 7405 5310 7420 5325
rect 7423 5322 7424 5334
rect 7431 5322 7458 5334
rect 7423 5314 7458 5322
rect 7423 5313 7452 5314
rect 7143 5300 7357 5304
rect 7158 5298 7357 5300
rect 7392 5300 7405 5310
rect 7423 5300 7440 5313
rect 7392 5298 7440 5300
rect 7034 5294 7067 5298
rect 7030 5292 7067 5294
rect 7030 5291 7097 5292
rect 7030 5286 7061 5291
rect 7067 5286 7097 5291
rect 7030 5282 7097 5286
rect 7003 5279 7097 5282
rect 7003 5272 7052 5279
rect 7003 5266 7033 5272
rect 7052 5267 7057 5272
rect 6969 5250 7049 5266
rect 7061 5258 7097 5279
rect 7158 5274 7347 5298
rect 7392 5297 7439 5298
rect 7405 5292 7439 5297
rect 7173 5271 7347 5274
rect 7166 5268 7347 5271
rect 7375 5291 7439 5292
rect 6969 5248 6988 5250
rect 7003 5248 7037 5250
rect 6969 5232 7049 5248
rect 6969 5226 6988 5232
rect 6685 5200 6788 5210
rect 6639 5198 6788 5200
rect 6809 5198 6844 5210
rect 6478 5196 6640 5198
rect 6490 5176 6509 5196
rect 6524 5194 6554 5196
rect 6373 5168 6414 5176
rect 6496 5172 6509 5176
rect 6561 5180 6640 5196
rect 6672 5196 6844 5198
rect 6672 5180 6751 5196
rect 6758 5194 6788 5196
rect 6336 5158 6365 5168
rect 6379 5158 6408 5168
rect 6423 5158 6453 5172
rect 6496 5158 6539 5172
rect 6561 5168 6751 5180
rect 6816 5176 6822 5196
rect 6546 5158 6576 5168
rect 6577 5158 6735 5168
rect 6739 5158 6769 5168
rect 6773 5158 6803 5172
rect 6831 5158 6844 5196
rect 6916 5210 6945 5226
rect 6959 5210 6988 5226
rect 7003 5216 7033 5232
rect 7061 5210 7067 5258
rect 7070 5252 7089 5258
rect 7104 5252 7134 5260
rect 7070 5244 7134 5252
rect 7070 5228 7150 5244
rect 7166 5237 7228 5268
rect 7244 5237 7306 5268
rect 7375 5266 7424 5291
rect 7439 5266 7469 5282
rect 7338 5252 7368 5260
rect 7375 5258 7485 5266
rect 7338 5244 7383 5252
rect 7070 5226 7089 5228
rect 7104 5226 7150 5228
rect 7070 5210 7150 5226
rect 7177 5224 7212 5237
rect 7253 5234 7290 5237
rect 7253 5232 7295 5234
rect 7182 5221 7212 5224
rect 7191 5217 7198 5221
rect 7198 5216 7199 5217
rect 7157 5210 7167 5216
rect 6916 5202 6951 5210
rect 6916 5176 6917 5202
rect 6924 5176 6951 5202
rect 6859 5158 6889 5172
rect 6916 5168 6951 5176
rect 6953 5202 6994 5210
rect 6953 5176 6968 5202
rect 6975 5176 6994 5202
rect 7058 5198 7089 5210
rect 7104 5198 7207 5210
rect 7219 5200 7245 5226
rect 7260 5221 7290 5232
rect 7322 5228 7384 5244
rect 7322 5226 7368 5228
rect 7322 5210 7384 5226
rect 7396 5210 7402 5258
rect 7405 5250 7485 5258
rect 7405 5248 7424 5250
rect 7439 5248 7473 5250
rect 7405 5232 7485 5248
rect 7405 5210 7424 5232
rect 7439 5216 7469 5232
rect 7497 5226 7503 5300
rect 7506 5226 7525 5370
rect 7540 5226 7546 5370
rect 7555 5300 7568 5370
rect 7613 5348 7614 5358
rect 7629 5348 7642 5358
rect 7613 5344 7642 5348
rect 7647 5344 7677 5370
rect 7695 5356 7711 5358
rect 7783 5356 7836 5370
rect 7784 5354 7848 5356
rect 7891 5354 7906 5370
rect 7955 5367 7985 5370
rect 7955 5364 7991 5367
rect 7921 5356 7937 5358
rect 7695 5344 7710 5348
rect 7613 5342 7710 5344
rect 7738 5342 7906 5354
rect 7922 5344 7937 5348
rect 7955 5345 7994 5364
rect 8013 5358 8020 5359
rect 8019 5351 8020 5358
rect 8003 5348 8004 5351
rect 8019 5348 8032 5351
rect 7955 5344 7985 5345
rect 7994 5344 8000 5345
rect 8003 5344 8032 5348
rect 7922 5343 8032 5344
rect 7922 5342 8038 5343
rect 7597 5334 7648 5342
rect 7597 5322 7622 5334
rect 7629 5322 7648 5334
rect 7679 5334 7729 5342
rect 7679 5326 7695 5334
rect 7702 5332 7729 5334
rect 7738 5332 7959 5342
rect 7702 5322 7959 5332
rect 7988 5334 8038 5342
rect 7988 5325 8004 5334
rect 7597 5314 7648 5322
rect 7695 5314 7959 5322
rect 7985 5322 8004 5325
rect 8011 5322 8038 5334
rect 7985 5314 8038 5322
rect 7549 5266 7568 5300
rect 7613 5306 7614 5314
rect 7629 5306 7642 5314
rect 7613 5298 7629 5306
rect 7610 5291 7629 5294
rect 7610 5282 7632 5291
rect 7583 5272 7632 5282
rect 7583 5266 7613 5272
rect 7632 5267 7637 5272
rect 7549 5250 7629 5266
rect 7647 5258 7677 5314
rect 7712 5304 7920 5314
rect 7955 5310 8000 5314
rect 8003 5313 8004 5314
rect 8019 5313 8032 5314
rect 7738 5274 7927 5304
rect 7753 5271 7927 5274
rect 7746 5268 7927 5271
rect 7549 5248 7568 5250
rect 7583 5248 7617 5250
rect 7549 5232 7629 5248
rect 7656 5244 7669 5258
rect 7684 5244 7700 5260
rect 7746 5255 7757 5268
rect 7549 5226 7568 5232
rect 7265 5200 7368 5210
rect 7219 5198 7368 5200
rect 7389 5198 7424 5210
rect 7058 5196 7220 5198
rect 7070 5176 7089 5196
rect 7104 5194 7134 5196
rect 6953 5168 6994 5176
rect 7076 5172 7089 5176
rect 7141 5180 7220 5196
rect 7252 5196 7424 5198
rect 7252 5180 7331 5196
rect 7338 5194 7368 5196
rect 6916 5158 6945 5168
rect 6959 5158 6988 5168
rect 7003 5158 7033 5172
rect 7076 5158 7119 5172
rect 7141 5168 7331 5180
rect 7396 5176 7402 5196
rect 7126 5158 7156 5168
rect 7157 5158 7315 5168
rect 7319 5158 7349 5168
rect 7353 5158 7383 5172
rect 7411 5158 7424 5196
rect 7496 5210 7525 5226
rect 7539 5210 7568 5226
rect 7583 5210 7613 5232
rect 7656 5228 7718 5244
rect 7746 5237 7757 5253
rect 7762 5248 7772 5268
rect 7782 5248 7796 5268
rect 7799 5255 7808 5268
rect 7824 5255 7833 5268
rect 7762 5237 7796 5248
rect 7799 5237 7808 5253
rect 7824 5237 7833 5253
rect 7840 5248 7850 5268
rect 7860 5248 7874 5268
rect 7875 5255 7886 5268
rect 7840 5237 7874 5248
rect 7875 5237 7886 5253
rect 7932 5244 7948 5260
rect 7955 5258 7985 5310
rect 8019 5306 8020 5313
rect 8004 5298 8020 5306
rect 7991 5266 8004 5285
rect 8019 5266 8049 5282
rect 7991 5250 8065 5266
rect 7991 5248 8004 5250
rect 8019 5248 8053 5250
rect 7656 5226 7669 5228
rect 7684 5226 7718 5228
rect 7656 5210 7718 5226
rect 7762 5221 7778 5224
rect 7840 5221 7870 5232
rect 7918 5228 7964 5244
rect 7991 5232 8065 5248
rect 7918 5226 7952 5228
rect 7917 5210 7964 5226
rect 7991 5210 8004 5232
rect 8019 5210 8049 5232
rect 8076 5210 8077 5226
rect 8092 5210 8105 5370
rect 8135 5266 8148 5370
rect 8193 5348 8194 5358
rect 8209 5348 8222 5358
rect 8193 5344 8222 5348
rect 8227 5344 8257 5370
rect 8275 5356 8291 5358
rect 8363 5356 8416 5370
rect 8364 5354 8428 5356
rect 8471 5354 8486 5370
rect 8535 5367 8565 5370
rect 8535 5364 8571 5367
rect 8501 5356 8517 5358
rect 8275 5344 8290 5348
rect 8193 5342 8290 5344
rect 8318 5342 8486 5354
rect 8502 5344 8517 5348
rect 8535 5345 8574 5364
rect 8593 5358 8600 5359
rect 8599 5351 8600 5358
rect 8583 5348 8584 5351
rect 8599 5348 8612 5351
rect 8535 5344 8565 5345
rect 8574 5344 8580 5345
rect 8583 5344 8612 5348
rect 8502 5343 8612 5344
rect 8502 5342 8618 5343
rect 8177 5334 8228 5342
rect 8177 5322 8202 5334
rect 8209 5322 8228 5334
rect 8259 5334 8309 5342
rect 8259 5326 8275 5334
rect 8282 5332 8309 5334
rect 8318 5332 8539 5342
rect 8282 5322 8539 5332
rect 8568 5334 8618 5342
rect 8568 5325 8584 5334
rect 8177 5314 8228 5322
rect 8275 5314 8539 5322
rect 8565 5322 8584 5325
rect 8591 5322 8618 5334
rect 8565 5314 8618 5322
rect 8193 5306 8194 5314
rect 8209 5306 8222 5314
rect 8193 5298 8209 5306
rect 8190 5291 8209 5294
rect 8190 5282 8212 5291
rect 8163 5272 8212 5282
rect 8163 5266 8193 5272
rect 8212 5267 8217 5272
rect 8135 5250 8209 5266
rect 8227 5258 8257 5314
rect 8292 5304 8500 5314
rect 8535 5310 8580 5314
rect 8583 5313 8584 5314
rect 8599 5313 8612 5314
rect 8318 5274 8507 5304
rect 8333 5271 8507 5274
rect 8326 5268 8507 5271
rect 8135 5248 8148 5250
rect 8163 5248 8197 5250
rect 8135 5232 8209 5248
rect 8236 5244 8249 5258
rect 8264 5244 8280 5260
rect 8326 5255 8337 5268
rect 8119 5210 8120 5226
rect 8135 5210 8148 5232
rect 8163 5210 8193 5232
rect 8236 5228 8298 5244
rect 8326 5237 8337 5253
rect 8342 5248 8352 5268
rect 8362 5248 8376 5268
rect 8379 5255 8388 5268
rect 8404 5255 8413 5268
rect 8342 5237 8376 5248
rect 8379 5237 8388 5253
rect 8404 5237 8413 5253
rect 8420 5248 8430 5268
rect 8440 5248 8454 5268
rect 8455 5255 8466 5268
rect 8420 5237 8454 5248
rect 8455 5237 8466 5253
rect 8512 5244 8528 5260
rect 8535 5258 8565 5310
rect 8599 5306 8600 5313
rect 8584 5298 8600 5306
rect 8571 5266 8584 5285
rect 8599 5266 8629 5282
rect 8571 5250 8645 5266
rect 8571 5248 8584 5250
rect 8599 5248 8633 5250
rect 8236 5226 8249 5228
rect 8264 5226 8298 5228
rect 8236 5210 8298 5226
rect 8342 5221 8358 5224
rect 8420 5221 8450 5232
rect 8498 5228 8544 5244
rect 8571 5232 8645 5248
rect 8498 5226 8532 5228
rect 8497 5210 8544 5226
rect 8571 5210 8584 5232
rect 8599 5210 8629 5232
rect 8656 5210 8657 5226
rect 8672 5210 8685 5370
rect 8715 5266 8728 5370
rect 8773 5348 8774 5358
rect 8789 5348 8802 5358
rect 8773 5344 8802 5348
rect 8807 5344 8837 5370
rect 8855 5356 8871 5358
rect 8943 5356 8996 5370
rect 8944 5354 9008 5356
rect 9051 5354 9066 5370
rect 9115 5367 9145 5370
rect 9115 5364 9151 5367
rect 9081 5356 9097 5358
rect 8855 5344 8870 5348
rect 8773 5342 8870 5344
rect 8898 5342 9066 5354
rect 9082 5344 9097 5348
rect 9115 5345 9154 5364
rect 9173 5358 9180 5359
rect 9179 5351 9180 5358
rect 9163 5348 9164 5351
rect 9179 5348 9192 5351
rect 9115 5344 9145 5345
rect 9154 5344 9160 5345
rect 9163 5344 9192 5348
rect 9082 5343 9192 5344
rect 9082 5342 9198 5343
rect 8757 5334 8808 5342
rect 8757 5322 8782 5334
rect 8789 5322 8808 5334
rect 8839 5334 8889 5342
rect 8839 5326 8855 5334
rect 8862 5332 8889 5334
rect 8898 5332 9119 5342
rect 8862 5322 9119 5332
rect 9148 5334 9198 5342
rect 9148 5325 9164 5334
rect 8757 5314 8808 5322
rect 8855 5314 9119 5322
rect 9145 5322 9164 5325
rect 9171 5322 9198 5334
rect 9145 5314 9198 5322
rect 8773 5306 8774 5314
rect 8789 5306 8802 5314
rect 8773 5298 8789 5306
rect 8770 5291 8789 5294
rect 8770 5282 8792 5291
rect 8743 5272 8792 5282
rect 8743 5266 8773 5272
rect 8792 5267 8797 5272
rect 8715 5250 8789 5266
rect 8807 5258 8837 5314
rect 8872 5304 9080 5314
rect 9115 5310 9160 5314
rect 9163 5313 9164 5314
rect 9179 5313 9192 5314
rect 8898 5274 9087 5304
rect 8913 5271 9087 5274
rect 8906 5268 9087 5271
rect 8715 5248 8728 5250
rect 8743 5248 8777 5250
rect 8715 5232 8789 5248
rect 8816 5244 8829 5258
rect 8844 5244 8860 5260
rect 8906 5255 8917 5268
rect 8699 5210 8700 5226
rect 8715 5210 8728 5232
rect 8743 5210 8773 5232
rect 8816 5228 8878 5244
rect 8906 5237 8917 5253
rect 8922 5248 8932 5268
rect 8942 5248 8956 5268
rect 8959 5255 8968 5268
rect 8984 5255 8993 5268
rect 8922 5237 8956 5248
rect 8959 5237 8968 5253
rect 8984 5237 8993 5253
rect 9000 5248 9010 5268
rect 9020 5248 9034 5268
rect 9035 5255 9046 5268
rect 9000 5237 9034 5248
rect 9035 5237 9046 5253
rect 9092 5244 9108 5260
rect 9115 5258 9145 5310
rect 9179 5306 9180 5313
rect 9164 5298 9180 5306
rect 9151 5266 9164 5285
rect 9179 5266 9209 5282
rect 9151 5250 9225 5266
rect 9151 5248 9164 5250
rect 9179 5248 9213 5250
rect 8816 5226 8829 5228
rect 8844 5226 8878 5228
rect 8816 5210 8878 5226
rect 8922 5221 8938 5224
rect 9000 5221 9030 5232
rect 9078 5228 9124 5244
rect 9151 5232 9225 5248
rect 9078 5226 9112 5228
rect 9077 5210 9124 5226
rect 9151 5210 9164 5232
rect 9179 5210 9209 5232
rect 9236 5210 9237 5226
rect 9252 5210 9265 5370
rect 7496 5202 7531 5210
rect 7496 5176 7497 5202
rect 7504 5176 7531 5202
rect 7439 5158 7469 5172
rect 7496 5168 7531 5176
rect 7533 5202 7574 5210
rect 7533 5176 7548 5202
rect 7555 5176 7574 5202
rect 7638 5198 7700 5210
rect 7712 5198 7787 5210
rect 7845 5198 7920 5210
rect 7932 5198 7963 5210
rect 7969 5198 8004 5210
rect 7638 5196 7800 5198
rect 7533 5168 7574 5176
rect 7656 5172 7669 5196
rect 7684 5194 7699 5196
rect 7496 5158 7525 5168
rect 7539 5158 7568 5168
rect 7583 5158 7613 5172
rect 7656 5158 7699 5172
rect 7723 5169 7730 5176
rect 7733 5172 7800 5196
rect 7832 5196 8004 5198
rect 7802 5174 7830 5178
rect 7832 5174 7912 5196
rect 7933 5194 7948 5196
rect 7802 5172 7912 5174
rect 7733 5168 7912 5172
rect 7706 5158 7736 5168
rect 7738 5158 7891 5168
rect 7899 5158 7929 5168
rect 7933 5158 7963 5172
rect 7991 5158 8004 5196
rect 8076 5202 8111 5210
rect 8076 5176 8077 5202
rect 8084 5176 8111 5202
rect 8019 5158 8049 5172
rect 8076 5168 8111 5176
rect 8113 5202 8154 5210
rect 8113 5176 8128 5202
rect 8135 5176 8154 5202
rect 8218 5198 8280 5210
rect 8292 5198 8367 5210
rect 8425 5198 8500 5210
rect 8512 5198 8543 5210
rect 8549 5198 8584 5210
rect 8218 5196 8380 5198
rect 8113 5168 8154 5176
rect 8236 5172 8249 5196
rect 8264 5194 8279 5196
rect 8076 5158 8077 5168
rect 8092 5158 8105 5168
rect 8119 5158 8120 5168
rect 8135 5158 8148 5168
rect 8163 5158 8193 5172
rect 8236 5158 8279 5172
rect 8303 5169 8310 5176
rect 8313 5172 8380 5196
rect 8412 5196 8584 5198
rect 8382 5174 8410 5178
rect 8412 5174 8492 5196
rect 8513 5194 8528 5196
rect 8382 5172 8492 5174
rect 8313 5168 8492 5172
rect 8286 5158 8316 5168
rect 8318 5158 8471 5168
rect 8479 5158 8509 5168
rect 8513 5158 8543 5172
rect 8571 5158 8584 5196
rect 8656 5202 8691 5210
rect 8656 5176 8657 5202
rect 8664 5176 8691 5202
rect 8599 5158 8629 5172
rect 8656 5168 8691 5176
rect 8693 5202 8734 5210
rect 8693 5176 8708 5202
rect 8715 5176 8734 5202
rect 8798 5198 8860 5210
rect 8872 5198 8947 5210
rect 9005 5198 9080 5210
rect 9092 5198 9123 5210
rect 9129 5198 9164 5210
rect 8798 5196 8960 5198
rect 8693 5168 8734 5176
rect 8816 5172 8829 5196
rect 8844 5194 8859 5196
rect 8656 5158 8657 5168
rect 8672 5158 8685 5168
rect 8699 5158 8700 5168
rect 8715 5158 8728 5168
rect 8743 5158 8773 5172
rect 8816 5158 8859 5172
rect 8883 5169 8890 5176
rect 8893 5172 8960 5196
rect 8992 5196 9164 5198
rect 8962 5174 8990 5178
rect 8992 5174 9072 5196
rect 9093 5194 9108 5196
rect 8962 5172 9072 5174
rect 8893 5168 9072 5172
rect 8866 5158 8896 5168
rect 8898 5158 9051 5168
rect 9059 5158 9089 5168
rect 9093 5158 9123 5172
rect 9151 5158 9164 5196
rect 9236 5202 9271 5210
rect 9236 5176 9237 5202
rect 9244 5176 9271 5202
rect 9179 5158 9209 5172
rect 9236 5168 9271 5176
rect 9236 5158 9237 5168
rect 9252 5158 9265 5168
rect -1 5152 9265 5158
rect 0 5144 9265 5152
rect 15 5114 28 5144
rect 43 5130 73 5144
rect 116 5130 159 5144
rect 166 5130 386 5144
rect 393 5130 423 5144
rect 83 5116 98 5128
rect 117 5116 130 5130
rect 198 5126 351 5130
rect 80 5114 102 5116
rect 180 5114 372 5126
rect 451 5114 464 5144
rect 479 5130 509 5144
rect 546 5114 565 5144
rect 580 5114 586 5144
rect 595 5114 608 5144
rect 623 5130 653 5144
rect 696 5130 739 5144
rect 746 5130 966 5144
rect 973 5130 1003 5144
rect 663 5116 678 5128
rect 697 5116 710 5130
rect 778 5126 931 5130
rect 660 5114 682 5116
rect 760 5114 952 5126
rect 1031 5114 1044 5144
rect 1059 5130 1089 5144
rect 1126 5114 1145 5144
rect 1160 5114 1166 5144
rect 1175 5114 1188 5144
rect 1203 5130 1233 5144
rect 1276 5130 1319 5144
rect 1326 5130 1546 5144
rect 1553 5130 1583 5144
rect 1243 5116 1258 5128
rect 1277 5116 1290 5130
rect 1358 5126 1511 5130
rect 1240 5114 1262 5116
rect 1340 5114 1532 5126
rect 1611 5114 1624 5144
rect 1639 5130 1669 5144
rect 1706 5114 1725 5144
rect 1740 5114 1746 5144
rect 1755 5114 1768 5144
rect 1783 5130 1813 5144
rect 1856 5130 1899 5144
rect 1906 5130 2126 5144
rect 2133 5130 2163 5144
rect 1823 5116 1838 5128
rect 1857 5116 1870 5130
rect 1938 5126 2091 5130
rect 1820 5114 1842 5116
rect 1920 5114 2112 5126
rect 2191 5114 2204 5144
rect 2219 5130 2249 5144
rect 2286 5114 2305 5144
rect 2320 5114 2326 5144
rect 2335 5114 2348 5144
rect 2363 5130 2393 5144
rect 2436 5130 2479 5144
rect 2486 5130 2706 5144
rect 2713 5130 2743 5144
rect 2403 5116 2418 5128
rect 2437 5116 2450 5130
rect 2518 5126 2671 5130
rect 2400 5114 2422 5116
rect 2500 5114 2692 5126
rect 2771 5114 2784 5144
rect 2799 5130 2829 5144
rect 2866 5114 2885 5144
rect 2900 5114 2906 5144
rect 2915 5114 2928 5144
rect 2943 5130 2973 5144
rect 3016 5130 3059 5144
rect 3066 5130 3286 5144
rect 3293 5130 3323 5144
rect 2983 5116 2998 5128
rect 3017 5116 3030 5130
rect 3098 5126 3251 5130
rect 2980 5114 3002 5116
rect 3080 5114 3272 5126
rect 3351 5114 3364 5144
rect 3379 5130 3409 5144
rect 3446 5114 3465 5144
rect 3480 5114 3486 5144
rect 3495 5114 3508 5144
rect 3523 5130 3553 5144
rect 3596 5130 3639 5144
rect 3646 5130 3866 5144
rect 3873 5130 3903 5144
rect 3563 5116 3578 5128
rect 3597 5116 3610 5130
rect 3678 5126 3831 5130
rect 3560 5114 3582 5116
rect 3660 5114 3852 5126
rect 3931 5114 3944 5144
rect 3959 5130 3989 5144
rect 4026 5114 4045 5144
rect 4060 5114 4066 5144
rect 4075 5114 4088 5144
rect 4103 5130 4133 5144
rect 4176 5130 4219 5144
rect 4226 5130 4446 5144
rect 4453 5130 4483 5144
rect 4143 5116 4158 5128
rect 4177 5116 4190 5130
rect 4258 5126 4411 5130
rect 4140 5114 4162 5116
rect 4240 5114 4432 5126
rect 4511 5114 4524 5144
rect 4539 5130 4569 5144
rect 4606 5114 4625 5144
rect 4640 5114 4646 5144
rect 4655 5114 4668 5144
rect 4683 5130 4713 5144
rect 4756 5130 4799 5144
rect 4806 5130 5026 5144
rect 5033 5130 5063 5144
rect 4723 5116 4738 5128
rect 4757 5116 4770 5130
rect 4838 5126 4991 5130
rect 4720 5114 4742 5116
rect 4820 5114 5012 5126
rect 5091 5114 5104 5144
rect 5119 5130 5149 5144
rect 5186 5114 5205 5144
rect 5220 5114 5226 5144
rect 5235 5114 5248 5144
rect 5263 5130 5293 5144
rect 5336 5130 5379 5144
rect 5386 5130 5606 5144
rect 5613 5130 5643 5144
rect 5303 5116 5318 5128
rect 5337 5116 5350 5130
rect 5418 5126 5571 5130
rect 5300 5114 5322 5116
rect 5400 5114 5592 5126
rect 5671 5114 5684 5144
rect 5699 5130 5729 5144
rect 5766 5114 5785 5144
rect 5800 5114 5806 5144
rect 5815 5114 5828 5144
rect 5843 5130 5873 5144
rect 5916 5130 5959 5144
rect 5966 5130 6186 5144
rect 6193 5130 6223 5144
rect 5883 5116 5898 5128
rect 5917 5116 5930 5130
rect 5998 5126 6151 5130
rect 5880 5114 5902 5116
rect 5980 5114 6172 5126
rect 6251 5114 6264 5144
rect 6279 5130 6309 5144
rect 6346 5114 6365 5144
rect 6380 5114 6386 5144
rect 6395 5114 6408 5144
rect 6423 5130 6453 5144
rect 6496 5130 6539 5144
rect 6546 5130 6766 5144
rect 6773 5130 6803 5144
rect 6463 5116 6478 5128
rect 6497 5116 6510 5130
rect 6578 5126 6731 5130
rect 6460 5114 6482 5116
rect 6560 5114 6752 5126
rect 6831 5114 6844 5144
rect 6859 5130 6889 5144
rect 6926 5114 6945 5144
rect 6960 5114 6966 5144
rect 6975 5114 6988 5144
rect 7003 5130 7033 5144
rect 7076 5130 7119 5144
rect 7126 5130 7346 5144
rect 7353 5130 7383 5144
rect 7043 5116 7058 5128
rect 7077 5116 7090 5130
rect 7158 5126 7311 5130
rect 7040 5114 7062 5116
rect 7140 5114 7332 5126
rect 7411 5114 7424 5144
rect 7439 5130 7469 5144
rect 7506 5114 7525 5144
rect 7540 5114 7546 5144
rect 7555 5114 7568 5144
rect 7583 5126 7613 5144
rect 7656 5130 7670 5144
rect 7706 5130 7926 5144
rect 7657 5128 7670 5130
rect 7623 5116 7638 5128
rect 7620 5114 7642 5116
rect 7647 5114 7677 5128
rect 7738 5126 7891 5130
rect 7720 5114 7912 5126
rect 7955 5114 7985 5128
rect 7991 5114 8004 5144
rect 8019 5126 8049 5144
rect 8092 5114 8105 5144
rect 8135 5114 8148 5144
rect 8163 5126 8193 5144
rect 8236 5130 8250 5144
rect 8286 5130 8506 5144
rect 8237 5128 8250 5130
rect 8203 5116 8218 5128
rect 8200 5114 8222 5116
rect 8227 5114 8257 5128
rect 8318 5126 8471 5130
rect 8300 5114 8492 5126
rect 8535 5114 8565 5128
rect 8571 5114 8584 5144
rect 8599 5126 8629 5144
rect 8672 5114 8685 5144
rect 8715 5114 8728 5144
rect 8743 5126 8773 5144
rect 8816 5130 8830 5144
rect 8866 5130 9086 5144
rect 8817 5128 8830 5130
rect 8783 5116 8798 5128
rect 8780 5114 8802 5116
rect 8807 5114 8837 5128
rect 8898 5126 9051 5130
rect 8880 5114 9072 5126
rect 9115 5114 9145 5128
rect 9151 5114 9164 5144
rect 9179 5126 9209 5144
rect 9252 5114 9265 5144
rect 0 5100 9265 5114
rect 15 5030 28 5100
rect 80 5096 102 5100
rect 73 5074 102 5088
rect 155 5074 171 5088
rect 209 5084 215 5086
rect 222 5084 330 5100
rect 337 5084 343 5086
rect 351 5084 366 5100
rect 432 5094 451 5097
rect 73 5072 171 5074
rect 198 5072 366 5084
rect 381 5074 397 5088
rect 432 5075 454 5094
rect 464 5088 480 5089
rect 463 5086 480 5088
rect 464 5081 480 5086
rect 454 5074 460 5075
rect 463 5074 492 5081
rect 381 5073 492 5074
rect 381 5072 498 5073
rect 57 5064 108 5072
rect 155 5064 189 5072
rect 57 5052 82 5064
rect 89 5052 108 5064
rect 162 5062 189 5064
rect 198 5062 419 5072
rect 454 5069 460 5072
rect 162 5058 419 5062
rect 57 5044 108 5052
rect 155 5044 419 5058
rect 463 5064 498 5072
rect 9 4996 28 5030
rect 73 5036 102 5044
rect 73 5030 90 5036
rect 73 5028 107 5030
rect 155 5028 171 5044
rect 172 5034 380 5044
rect 381 5034 397 5044
rect 445 5040 460 5055
rect 463 5052 464 5064
rect 471 5052 498 5064
rect 463 5044 498 5052
rect 463 5043 492 5044
rect 183 5030 397 5034
rect 198 5028 397 5030
rect 432 5030 445 5040
rect 463 5030 480 5043
rect 432 5028 480 5030
rect 74 5024 107 5028
rect 70 5022 107 5024
rect 70 5021 137 5022
rect 70 5016 101 5021
rect 107 5016 137 5021
rect 70 5012 137 5016
rect 43 5009 137 5012
rect 43 5002 92 5009
rect 43 4996 73 5002
rect 92 4997 97 5002
rect 9 4980 89 4996
rect 101 4988 137 5009
rect 198 5004 387 5028
rect 432 5027 479 5028
rect 445 5022 479 5027
rect 213 5001 387 5004
rect 206 4998 387 5001
rect 415 5021 479 5022
rect 9 4978 28 4980
rect 43 4978 77 4980
rect 9 4962 89 4978
rect 9 4956 28 4962
rect -1 4940 28 4956
rect 43 4946 73 4962
rect 101 4940 107 4988
rect 110 4982 129 4988
rect 144 4982 174 4990
rect 110 4974 174 4982
rect 110 4958 190 4974
rect 206 4967 268 4998
rect 284 4967 346 4998
rect 415 4996 464 5021
rect 479 4996 509 5012
rect 378 4982 408 4990
rect 415 4988 525 4996
rect 378 4974 423 4982
rect 110 4956 129 4958
rect 144 4956 190 4958
rect 110 4940 190 4956
rect 217 4954 252 4967
rect 293 4964 330 4967
rect 293 4962 335 4964
rect 222 4951 252 4954
rect 231 4947 238 4951
rect 238 4946 239 4947
rect 197 4940 207 4946
rect -7 4932 34 4940
rect -7 4906 8 4932
rect 15 4906 34 4932
rect 98 4928 129 4940
rect 144 4928 247 4940
rect 259 4930 285 4956
rect 300 4951 330 4962
rect 362 4958 424 4974
rect 362 4956 408 4958
rect 362 4940 424 4956
rect 436 4940 442 4988
rect 445 4980 525 4988
rect 445 4978 464 4980
rect 479 4978 513 4980
rect 445 4962 525 4978
rect 445 4940 464 4962
rect 479 4946 509 4962
rect 537 4956 543 5030
rect 546 4956 565 5100
rect 580 4956 586 5100
rect 595 5030 608 5100
rect 660 5096 682 5100
rect 653 5074 682 5088
rect 735 5074 751 5088
rect 789 5084 795 5086
rect 802 5084 910 5100
rect 917 5084 923 5086
rect 931 5084 946 5100
rect 1012 5094 1031 5097
rect 653 5072 751 5074
rect 778 5072 946 5084
rect 961 5074 977 5088
rect 1012 5075 1034 5094
rect 1044 5088 1060 5089
rect 1043 5086 1060 5088
rect 1044 5081 1060 5086
rect 1034 5074 1040 5075
rect 1043 5074 1072 5081
rect 961 5073 1072 5074
rect 961 5072 1078 5073
rect 637 5064 688 5072
rect 735 5064 769 5072
rect 637 5052 662 5064
rect 669 5052 688 5064
rect 742 5062 769 5064
rect 778 5062 999 5072
rect 1034 5069 1040 5072
rect 742 5058 999 5062
rect 637 5044 688 5052
rect 735 5044 999 5058
rect 1043 5064 1078 5072
rect 589 4996 608 5030
rect 653 5036 682 5044
rect 653 5030 670 5036
rect 653 5028 687 5030
rect 735 5028 751 5044
rect 752 5034 960 5044
rect 961 5034 977 5044
rect 1025 5040 1040 5055
rect 1043 5052 1044 5064
rect 1051 5052 1078 5064
rect 1043 5044 1078 5052
rect 1043 5043 1072 5044
rect 763 5030 977 5034
rect 778 5028 977 5030
rect 1012 5030 1025 5040
rect 1043 5030 1060 5043
rect 1012 5028 1060 5030
rect 654 5024 687 5028
rect 650 5022 687 5024
rect 650 5021 717 5022
rect 650 5016 681 5021
rect 687 5016 717 5021
rect 650 5012 717 5016
rect 623 5009 717 5012
rect 623 5002 672 5009
rect 623 4996 653 5002
rect 672 4997 677 5002
rect 589 4980 669 4996
rect 681 4988 717 5009
rect 778 5004 967 5028
rect 1012 5027 1059 5028
rect 1025 5022 1059 5027
rect 793 5001 967 5004
rect 786 4998 967 5001
rect 995 5021 1059 5022
rect 589 4978 608 4980
rect 623 4978 657 4980
rect 589 4962 669 4978
rect 589 4956 608 4962
rect 305 4930 408 4940
rect 259 4928 408 4930
rect 429 4928 464 4940
rect 98 4926 260 4928
rect 110 4906 129 4926
rect 144 4924 174 4926
rect -7 4898 34 4906
rect 116 4902 129 4906
rect 181 4910 260 4926
rect 292 4926 464 4928
rect 292 4910 371 4926
rect 378 4924 408 4926
rect -1 4888 28 4898
rect 43 4888 73 4902
rect 116 4888 159 4902
rect 181 4898 371 4910
rect 436 4906 442 4926
rect 166 4888 196 4898
rect 197 4888 355 4898
rect 359 4888 389 4898
rect 393 4888 423 4902
rect 451 4888 464 4926
rect 536 4940 565 4956
rect 579 4940 608 4956
rect 623 4946 653 4962
rect 681 4940 687 4988
rect 690 4982 709 4988
rect 724 4982 754 4990
rect 690 4974 754 4982
rect 690 4958 770 4974
rect 786 4967 848 4998
rect 864 4967 926 4998
rect 995 4996 1044 5021
rect 1059 4996 1089 5012
rect 958 4982 988 4990
rect 995 4988 1105 4996
rect 958 4974 1003 4982
rect 690 4956 709 4958
rect 724 4956 770 4958
rect 690 4940 770 4956
rect 797 4954 832 4967
rect 873 4964 910 4967
rect 873 4962 915 4964
rect 802 4951 832 4954
rect 811 4947 818 4951
rect 818 4946 819 4947
rect 777 4940 787 4946
rect 536 4932 571 4940
rect 536 4906 537 4932
rect 544 4906 571 4932
rect 479 4888 509 4902
rect 536 4898 571 4906
rect 573 4932 614 4940
rect 573 4906 588 4932
rect 595 4906 614 4932
rect 678 4928 709 4940
rect 724 4928 827 4940
rect 839 4930 865 4956
rect 880 4951 910 4962
rect 942 4958 1004 4974
rect 942 4956 988 4958
rect 942 4940 1004 4956
rect 1016 4940 1022 4988
rect 1025 4980 1105 4988
rect 1025 4978 1044 4980
rect 1059 4978 1093 4980
rect 1025 4962 1105 4978
rect 1025 4940 1044 4962
rect 1059 4946 1089 4962
rect 1117 4956 1123 5030
rect 1126 4956 1145 5100
rect 1160 4956 1166 5100
rect 1175 5030 1188 5100
rect 1240 5096 1262 5100
rect 1233 5074 1262 5088
rect 1315 5074 1331 5088
rect 1369 5084 1375 5086
rect 1382 5084 1490 5100
rect 1497 5084 1503 5086
rect 1511 5084 1526 5100
rect 1592 5094 1611 5097
rect 1233 5072 1331 5074
rect 1358 5072 1526 5084
rect 1541 5074 1557 5088
rect 1592 5075 1614 5094
rect 1624 5088 1640 5089
rect 1623 5086 1640 5088
rect 1624 5081 1640 5086
rect 1614 5074 1620 5075
rect 1623 5074 1652 5081
rect 1541 5073 1652 5074
rect 1541 5072 1658 5073
rect 1217 5064 1268 5072
rect 1315 5064 1349 5072
rect 1217 5052 1242 5064
rect 1249 5052 1268 5064
rect 1322 5062 1349 5064
rect 1358 5062 1579 5072
rect 1614 5069 1620 5072
rect 1322 5058 1579 5062
rect 1217 5044 1268 5052
rect 1315 5044 1579 5058
rect 1623 5064 1658 5072
rect 1169 4996 1188 5030
rect 1233 5036 1262 5044
rect 1233 5030 1250 5036
rect 1233 5028 1267 5030
rect 1315 5028 1331 5044
rect 1332 5034 1540 5044
rect 1541 5034 1557 5044
rect 1605 5040 1620 5055
rect 1623 5052 1624 5064
rect 1631 5052 1658 5064
rect 1623 5044 1658 5052
rect 1623 5043 1652 5044
rect 1343 5030 1557 5034
rect 1358 5028 1557 5030
rect 1592 5030 1605 5040
rect 1623 5030 1640 5043
rect 1592 5028 1640 5030
rect 1234 5024 1267 5028
rect 1230 5022 1267 5024
rect 1230 5021 1297 5022
rect 1230 5016 1261 5021
rect 1267 5016 1297 5021
rect 1230 5012 1297 5016
rect 1203 5009 1297 5012
rect 1203 5002 1252 5009
rect 1203 4996 1233 5002
rect 1252 4997 1257 5002
rect 1169 4980 1249 4996
rect 1261 4988 1297 5009
rect 1358 5004 1547 5028
rect 1592 5027 1639 5028
rect 1605 5022 1639 5027
rect 1373 5001 1547 5004
rect 1366 4998 1547 5001
rect 1575 5021 1639 5022
rect 1169 4978 1188 4980
rect 1203 4978 1237 4980
rect 1169 4962 1249 4978
rect 1169 4956 1188 4962
rect 885 4930 988 4940
rect 839 4928 988 4930
rect 1009 4928 1044 4940
rect 678 4926 840 4928
rect 690 4906 709 4926
rect 724 4924 754 4926
rect 573 4898 614 4906
rect 696 4902 709 4906
rect 761 4910 840 4926
rect 872 4926 1044 4928
rect 872 4910 951 4926
rect 958 4924 988 4926
rect 536 4888 565 4898
rect 579 4888 608 4898
rect 623 4888 653 4902
rect 696 4888 739 4902
rect 761 4898 951 4910
rect 1016 4906 1022 4926
rect 746 4888 776 4898
rect 777 4888 935 4898
rect 939 4888 969 4898
rect 973 4888 1003 4902
rect 1031 4888 1044 4926
rect 1116 4940 1145 4956
rect 1159 4940 1188 4956
rect 1203 4946 1233 4962
rect 1261 4940 1267 4988
rect 1270 4982 1289 4988
rect 1304 4982 1334 4990
rect 1270 4974 1334 4982
rect 1270 4958 1350 4974
rect 1366 4967 1428 4998
rect 1444 4967 1506 4998
rect 1575 4996 1624 5021
rect 1639 4996 1669 5012
rect 1538 4982 1568 4990
rect 1575 4988 1685 4996
rect 1538 4974 1583 4982
rect 1270 4956 1289 4958
rect 1304 4956 1350 4958
rect 1270 4940 1350 4956
rect 1377 4954 1412 4967
rect 1453 4964 1490 4967
rect 1453 4962 1495 4964
rect 1382 4951 1412 4954
rect 1391 4947 1398 4951
rect 1398 4946 1399 4947
rect 1357 4940 1367 4946
rect 1116 4932 1151 4940
rect 1116 4906 1117 4932
rect 1124 4906 1151 4932
rect 1059 4888 1089 4902
rect 1116 4898 1151 4906
rect 1153 4932 1194 4940
rect 1153 4906 1168 4932
rect 1175 4906 1194 4932
rect 1258 4928 1289 4940
rect 1304 4928 1407 4940
rect 1419 4930 1445 4956
rect 1460 4951 1490 4962
rect 1522 4958 1584 4974
rect 1522 4956 1568 4958
rect 1522 4940 1584 4956
rect 1596 4940 1602 4988
rect 1605 4980 1685 4988
rect 1605 4978 1624 4980
rect 1639 4978 1673 4980
rect 1605 4962 1685 4978
rect 1605 4940 1624 4962
rect 1639 4946 1669 4962
rect 1697 4956 1703 5030
rect 1706 4956 1725 5100
rect 1740 4956 1746 5100
rect 1755 5030 1768 5100
rect 1820 5096 1842 5100
rect 1813 5074 1842 5088
rect 1895 5074 1911 5088
rect 1949 5084 1955 5086
rect 1962 5084 2070 5100
rect 2077 5084 2083 5086
rect 2091 5084 2106 5100
rect 2172 5094 2191 5097
rect 1813 5072 1911 5074
rect 1938 5072 2106 5084
rect 2121 5074 2137 5088
rect 2172 5075 2194 5094
rect 2204 5088 2220 5089
rect 2203 5086 2220 5088
rect 2204 5081 2220 5086
rect 2194 5074 2200 5075
rect 2203 5074 2232 5081
rect 2121 5073 2232 5074
rect 2121 5072 2238 5073
rect 1797 5064 1848 5072
rect 1895 5064 1929 5072
rect 1797 5052 1822 5064
rect 1829 5052 1848 5064
rect 1902 5062 1929 5064
rect 1938 5062 2159 5072
rect 2194 5069 2200 5072
rect 1902 5058 2159 5062
rect 1797 5044 1848 5052
rect 1895 5044 2159 5058
rect 2203 5064 2238 5072
rect 1749 4996 1768 5030
rect 1813 5036 1842 5044
rect 1813 5030 1830 5036
rect 1813 5028 1847 5030
rect 1895 5028 1911 5044
rect 1912 5034 2120 5044
rect 2121 5034 2137 5044
rect 2185 5040 2200 5055
rect 2203 5052 2204 5064
rect 2211 5052 2238 5064
rect 2203 5044 2238 5052
rect 2203 5043 2232 5044
rect 1923 5030 2137 5034
rect 1938 5028 2137 5030
rect 2172 5030 2185 5040
rect 2203 5030 2220 5043
rect 2172 5028 2220 5030
rect 1814 5024 1847 5028
rect 1810 5022 1847 5024
rect 1810 5021 1877 5022
rect 1810 5016 1841 5021
rect 1847 5016 1877 5021
rect 1810 5012 1877 5016
rect 1783 5009 1877 5012
rect 1783 5002 1832 5009
rect 1783 4996 1813 5002
rect 1832 4997 1837 5002
rect 1749 4980 1829 4996
rect 1841 4988 1877 5009
rect 1938 5004 2127 5028
rect 2172 5027 2219 5028
rect 2185 5022 2219 5027
rect 1953 5001 2127 5004
rect 1946 4998 2127 5001
rect 2155 5021 2219 5022
rect 1749 4978 1768 4980
rect 1783 4978 1817 4980
rect 1749 4962 1829 4978
rect 1749 4956 1768 4962
rect 1465 4930 1568 4940
rect 1419 4928 1568 4930
rect 1589 4928 1624 4940
rect 1258 4926 1420 4928
rect 1270 4906 1289 4926
rect 1304 4924 1334 4926
rect 1153 4898 1194 4906
rect 1276 4902 1289 4906
rect 1341 4910 1420 4926
rect 1452 4926 1624 4928
rect 1452 4910 1531 4926
rect 1538 4924 1568 4926
rect 1116 4888 1145 4898
rect 1159 4888 1188 4898
rect 1203 4888 1233 4902
rect 1276 4888 1319 4902
rect 1341 4898 1531 4910
rect 1596 4906 1602 4926
rect 1326 4888 1356 4898
rect 1357 4888 1515 4898
rect 1519 4888 1549 4898
rect 1553 4888 1583 4902
rect 1611 4888 1624 4926
rect 1696 4940 1725 4956
rect 1739 4940 1768 4956
rect 1783 4946 1813 4962
rect 1841 4940 1847 4988
rect 1850 4982 1869 4988
rect 1884 4982 1914 4990
rect 1850 4974 1914 4982
rect 1850 4958 1930 4974
rect 1946 4967 2008 4998
rect 2024 4967 2086 4998
rect 2155 4996 2204 5021
rect 2219 4996 2249 5012
rect 2118 4982 2148 4990
rect 2155 4988 2265 4996
rect 2118 4974 2163 4982
rect 1850 4956 1869 4958
rect 1884 4956 1930 4958
rect 1850 4940 1930 4956
rect 1957 4954 1992 4967
rect 2033 4964 2070 4967
rect 2033 4962 2075 4964
rect 1962 4951 1992 4954
rect 1971 4947 1978 4951
rect 1978 4946 1979 4947
rect 1937 4940 1947 4946
rect 1696 4932 1731 4940
rect 1696 4906 1697 4932
rect 1704 4906 1731 4932
rect 1639 4888 1669 4902
rect 1696 4898 1731 4906
rect 1733 4932 1774 4940
rect 1733 4906 1748 4932
rect 1755 4906 1774 4932
rect 1838 4928 1869 4940
rect 1884 4928 1987 4940
rect 1999 4930 2025 4956
rect 2040 4951 2070 4962
rect 2102 4958 2164 4974
rect 2102 4956 2148 4958
rect 2102 4940 2164 4956
rect 2176 4940 2182 4988
rect 2185 4980 2265 4988
rect 2185 4978 2204 4980
rect 2219 4978 2253 4980
rect 2185 4962 2265 4978
rect 2185 4940 2204 4962
rect 2219 4946 2249 4962
rect 2277 4956 2283 5030
rect 2286 4956 2305 5100
rect 2320 4956 2326 5100
rect 2335 5030 2348 5100
rect 2400 5096 2422 5100
rect 2393 5074 2422 5088
rect 2475 5074 2491 5088
rect 2529 5084 2535 5086
rect 2542 5084 2650 5100
rect 2657 5084 2663 5086
rect 2671 5084 2686 5100
rect 2752 5094 2771 5097
rect 2393 5072 2491 5074
rect 2518 5072 2686 5084
rect 2701 5074 2717 5088
rect 2752 5075 2774 5094
rect 2784 5088 2800 5089
rect 2783 5086 2800 5088
rect 2784 5081 2800 5086
rect 2774 5074 2780 5075
rect 2783 5074 2812 5081
rect 2701 5073 2812 5074
rect 2701 5072 2818 5073
rect 2377 5064 2428 5072
rect 2475 5064 2509 5072
rect 2377 5052 2402 5064
rect 2409 5052 2428 5064
rect 2482 5062 2509 5064
rect 2518 5062 2739 5072
rect 2774 5069 2780 5072
rect 2482 5058 2739 5062
rect 2377 5044 2428 5052
rect 2475 5044 2739 5058
rect 2783 5064 2818 5072
rect 2329 4996 2348 5030
rect 2393 5036 2422 5044
rect 2393 5030 2410 5036
rect 2393 5028 2427 5030
rect 2475 5028 2491 5044
rect 2492 5034 2700 5044
rect 2701 5034 2717 5044
rect 2765 5040 2780 5055
rect 2783 5052 2784 5064
rect 2791 5052 2818 5064
rect 2783 5044 2818 5052
rect 2783 5043 2812 5044
rect 2503 5030 2717 5034
rect 2518 5028 2717 5030
rect 2752 5030 2765 5040
rect 2783 5030 2800 5043
rect 2752 5028 2800 5030
rect 2394 5024 2427 5028
rect 2390 5022 2427 5024
rect 2390 5021 2457 5022
rect 2390 5016 2421 5021
rect 2427 5016 2457 5021
rect 2390 5012 2457 5016
rect 2363 5009 2457 5012
rect 2363 5002 2412 5009
rect 2363 4996 2393 5002
rect 2412 4997 2417 5002
rect 2329 4980 2409 4996
rect 2421 4988 2457 5009
rect 2518 5004 2707 5028
rect 2752 5027 2799 5028
rect 2765 5022 2799 5027
rect 2533 5001 2707 5004
rect 2526 4998 2707 5001
rect 2735 5021 2799 5022
rect 2329 4978 2348 4980
rect 2363 4978 2397 4980
rect 2329 4962 2409 4978
rect 2329 4956 2348 4962
rect 2045 4930 2148 4940
rect 1999 4928 2148 4930
rect 2169 4928 2204 4940
rect 1838 4926 2000 4928
rect 1850 4906 1869 4926
rect 1884 4924 1914 4926
rect 1733 4898 1774 4906
rect 1856 4902 1869 4906
rect 1921 4910 2000 4926
rect 2032 4926 2204 4928
rect 2032 4910 2111 4926
rect 2118 4924 2148 4926
rect 1696 4888 1725 4898
rect 1739 4888 1768 4898
rect 1783 4888 1813 4902
rect 1856 4888 1899 4902
rect 1921 4898 2111 4910
rect 2176 4906 2182 4926
rect 1906 4888 1936 4898
rect 1937 4888 2095 4898
rect 2099 4888 2129 4898
rect 2133 4888 2163 4902
rect 2191 4888 2204 4926
rect 2276 4940 2305 4956
rect 2319 4940 2348 4956
rect 2363 4946 2393 4962
rect 2421 4940 2427 4988
rect 2430 4982 2449 4988
rect 2464 4982 2494 4990
rect 2430 4974 2494 4982
rect 2430 4958 2510 4974
rect 2526 4967 2588 4998
rect 2604 4967 2666 4998
rect 2735 4996 2784 5021
rect 2799 4996 2829 5012
rect 2698 4982 2728 4990
rect 2735 4988 2845 4996
rect 2698 4974 2743 4982
rect 2430 4956 2449 4958
rect 2464 4956 2510 4958
rect 2430 4940 2510 4956
rect 2537 4954 2572 4967
rect 2613 4964 2650 4967
rect 2613 4962 2655 4964
rect 2542 4951 2572 4954
rect 2551 4947 2558 4951
rect 2558 4946 2559 4947
rect 2517 4940 2527 4946
rect 2276 4932 2311 4940
rect 2276 4906 2277 4932
rect 2284 4906 2311 4932
rect 2219 4888 2249 4902
rect 2276 4898 2311 4906
rect 2313 4932 2354 4940
rect 2313 4906 2328 4932
rect 2335 4906 2354 4932
rect 2418 4928 2449 4940
rect 2464 4928 2567 4940
rect 2579 4930 2605 4956
rect 2620 4951 2650 4962
rect 2682 4958 2744 4974
rect 2682 4956 2728 4958
rect 2682 4940 2744 4956
rect 2756 4940 2762 4988
rect 2765 4980 2845 4988
rect 2765 4978 2784 4980
rect 2799 4978 2833 4980
rect 2765 4962 2845 4978
rect 2765 4940 2784 4962
rect 2799 4946 2829 4962
rect 2857 4956 2863 5030
rect 2866 4956 2885 5100
rect 2900 4956 2906 5100
rect 2915 5030 2928 5100
rect 2980 5096 3002 5100
rect 2973 5074 3002 5088
rect 3055 5074 3071 5088
rect 3109 5084 3115 5086
rect 3122 5084 3230 5100
rect 3237 5084 3243 5086
rect 3251 5084 3266 5100
rect 3332 5094 3351 5097
rect 2973 5072 3071 5074
rect 3098 5072 3266 5084
rect 3281 5074 3297 5088
rect 3332 5075 3354 5094
rect 3364 5088 3380 5089
rect 3363 5086 3380 5088
rect 3364 5081 3380 5086
rect 3354 5074 3360 5075
rect 3363 5074 3392 5081
rect 3281 5073 3392 5074
rect 3281 5072 3398 5073
rect 2957 5064 3008 5072
rect 3055 5064 3089 5072
rect 2957 5052 2982 5064
rect 2989 5052 3008 5064
rect 3062 5062 3089 5064
rect 3098 5062 3319 5072
rect 3354 5069 3360 5072
rect 3062 5058 3319 5062
rect 2957 5044 3008 5052
rect 3055 5044 3319 5058
rect 3363 5064 3398 5072
rect 2909 4996 2928 5030
rect 2973 5036 3002 5044
rect 2973 5030 2990 5036
rect 2973 5028 3007 5030
rect 3055 5028 3071 5044
rect 3072 5034 3280 5044
rect 3281 5034 3297 5044
rect 3345 5040 3360 5055
rect 3363 5052 3364 5064
rect 3371 5052 3398 5064
rect 3363 5044 3398 5052
rect 3363 5043 3392 5044
rect 3083 5030 3297 5034
rect 3098 5028 3297 5030
rect 3332 5030 3345 5040
rect 3363 5030 3380 5043
rect 3332 5028 3380 5030
rect 2974 5024 3007 5028
rect 2970 5022 3007 5024
rect 2970 5021 3037 5022
rect 2970 5016 3001 5021
rect 3007 5016 3037 5021
rect 2970 5012 3037 5016
rect 2943 5009 3037 5012
rect 2943 5002 2992 5009
rect 2943 4996 2973 5002
rect 2992 4997 2997 5002
rect 2909 4980 2989 4996
rect 3001 4988 3037 5009
rect 3098 5004 3287 5028
rect 3332 5027 3379 5028
rect 3345 5022 3379 5027
rect 3113 5001 3287 5004
rect 3106 4998 3287 5001
rect 3315 5021 3379 5022
rect 2909 4978 2928 4980
rect 2943 4978 2977 4980
rect 2909 4962 2989 4978
rect 2909 4956 2928 4962
rect 2625 4930 2728 4940
rect 2579 4928 2728 4930
rect 2749 4928 2784 4940
rect 2418 4926 2580 4928
rect 2430 4906 2449 4926
rect 2464 4924 2494 4926
rect 2313 4898 2354 4906
rect 2436 4902 2449 4906
rect 2501 4910 2580 4926
rect 2612 4926 2784 4928
rect 2612 4910 2691 4926
rect 2698 4924 2728 4926
rect 2276 4888 2305 4898
rect 2319 4888 2348 4898
rect 2363 4888 2393 4902
rect 2436 4888 2479 4902
rect 2501 4898 2691 4910
rect 2756 4906 2762 4926
rect 2486 4888 2516 4898
rect 2517 4888 2675 4898
rect 2679 4888 2709 4898
rect 2713 4888 2743 4902
rect 2771 4888 2784 4926
rect 2856 4940 2885 4956
rect 2899 4940 2928 4956
rect 2943 4946 2973 4962
rect 3001 4940 3007 4988
rect 3010 4982 3029 4988
rect 3044 4982 3074 4990
rect 3010 4974 3074 4982
rect 3010 4958 3090 4974
rect 3106 4967 3168 4998
rect 3184 4967 3246 4998
rect 3315 4996 3364 5021
rect 3379 4996 3409 5012
rect 3278 4982 3308 4990
rect 3315 4988 3425 4996
rect 3278 4974 3323 4982
rect 3010 4956 3029 4958
rect 3044 4956 3090 4958
rect 3010 4940 3090 4956
rect 3117 4954 3152 4967
rect 3193 4964 3230 4967
rect 3193 4962 3235 4964
rect 3122 4951 3152 4954
rect 3131 4947 3138 4951
rect 3138 4946 3139 4947
rect 3097 4940 3107 4946
rect 2856 4932 2891 4940
rect 2856 4906 2857 4932
rect 2864 4906 2891 4932
rect 2799 4888 2829 4902
rect 2856 4898 2891 4906
rect 2893 4932 2934 4940
rect 2893 4906 2908 4932
rect 2915 4906 2934 4932
rect 2998 4928 3029 4940
rect 3044 4928 3147 4940
rect 3159 4930 3185 4956
rect 3200 4951 3230 4962
rect 3262 4958 3324 4974
rect 3262 4956 3308 4958
rect 3262 4940 3324 4956
rect 3336 4940 3342 4988
rect 3345 4980 3425 4988
rect 3345 4978 3364 4980
rect 3379 4978 3413 4980
rect 3345 4962 3425 4978
rect 3345 4940 3364 4962
rect 3379 4946 3409 4962
rect 3437 4956 3443 5030
rect 3446 4956 3465 5100
rect 3480 4956 3486 5100
rect 3495 5030 3508 5100
rect 3560 5096 3582 5100
rect 3553 5074 3582 5088
rect 3635 5074 3651 5088
rect 3689 5084 3695 5086
rect 3702 5084 3810 5100
rect 3817 5084 3823 5086
rect 3831 5084 3846 5100
rect 3912 5094 3931 5097
rect 3553 5072 3651 5074
rect 3678 5072 3846 5084
rect 3861 5074 3877 5088
rect 3912 5075 3934 5094
rect 3944 5088 3960 5089
rect 3943 5086 3960 5088
rect 3944 5081 3960 5086
rect 3934 5074 3940 5075
rect 3943 5074 3972 5081
rect 3861 5073 3972 5074
rect 3861 5072 3978 5073
rect 3537 5064 3588 5072
rect 3635 5064 3669 5072
rect 3537 5052 3562 5064
rect 3569 5052 3588 5064
rect 3642 5062 3669 5064
rect 3678 5062 3899 5072
rect 3934 5069 3940 5072
rect 3642 5058 3899 5062
rect 3537 5044 3588 5052
rect 3635 5044 3899 5058
rect 3943 5064 3978 5072
rect 3489 4996 3508 5030
rect 3553 5036 3582 5044
rect 3553 5030 3570 5036
rect 3553 5028 3587 5030
rect 3635 5028 3651 5044
rect 3652 5034 3860 5044
rect 3861 5034 3877 5044
rect 3925 5040 3940 5055
rect 3943 5052 3944 5064
rect 3951 5052 3978 5064
rect 3943 5044 3978 5052
rect 3943 5043 3972 5044
rect 3663 5030 3877 5034
rect 3678 5028 3877 5030
rect 3912 5030 3925 5040
rect 3943 5030 3960 5043
rect 3912 5028 3960 5030
rect 3554 5024 3587 5028
rect 3550 5022 3587 5024
rect 3550 5021 3617 5022
rect 3550 5016 3581 5021
rect 3587 5016 3617 5021
rect 3550 5012 3617 5016
rect 3523 5009 3617 5012
rect 3523 5002 3572 5009
rect 3523 4996 3553 5002
rect 3572 4997 3577 5002
rect 3489 4980 3569 4996
rect 3581 4988 3617 5009
rect 3678 5004 3867 5028
rect 3912 5027 3959 5028
rect 3925 5022 3959 5027
rect 3693 5001 3867 5004
rect 3686 4998 3867 5001
rect 3895 5021 3959 5022
rect 3489 4978 3508 4980
rect 3523 4978 3557 4980
rect 3489 4962 3569 4978
rect 3489 4956 3508 4962
rect 3205 4930 3308 4940
rect 3159 4928 3308 4930
rect 3329 4928 3364 4940
rect 2998 4926 3160 4928
rect 3010 4906 3029 4926
rect 3044 4924 3074 4926
rect 2893 4898 2934 4906
rect 3016 4902 3029 4906
rect 3081 4910 3160 4926
rect 3192 4926 3364 4928
rect 3192 4910 3271 4926
rect 3278 4924 3308 4926
rect 2856 4888 2885 4898
rect 2899 4888 2928 4898
rect 2943 4888 2973 4902
rect 3016 4888 3059 4902
rect 3081 4898 3271 4910
rect 3336 4906 3342 4926
rect 3066 4888 3096 4898
rect 3097 4888 3255 4898
rect 3259 4888 3289 4898
rect 3293 4888 3323 4902
rect 3351 4888 3364 4926
rect 3436 4940 3465 4956
rect 3479 4940 3508 4956
rect 3523 4946 3553 4962
rect 3581 4940 3587 4988
rect 3590 4982 3609 4988
rect 3624 4982 3654 4990
rect 3590 4974 3654 4982
rect 3590 4958 3670 4974
rect 3686 4967 3748 4998
rect 3764 4967 3826 4998
rect 3895 4996 3944 5021
rect 3959 4996 3989 5012
rect 3858 4982 3888 4990
rect 3895 4988 4005 4996
rect 3858 4974 3903 4982
rect 3590 4956 3609 4958
rect 3624 4956 3670 4958
rect 3590 4940 3670 4956
rect 3697 4954 3732 4967
rect 3773 4964 3810 4967
rect 3773 4962 3815 4964
rect 3702 4951 3732 4954
rect 3711 4947 3718 4951
rect 3718 4946 3719 4947
rect 3677 4940 3687 4946
rect 3436 4932 3471 4940
rect 3436 4906 3437 4932
rect 3444 4906 3471 4932
rect 3379 4888 3409 4902
rect 3436 4898 3471 4906
rect 3473 4932 3514 4940
rect 3473 4906 3488 4932
rect 3495 4906 3514 4932
rect 3578 4928 3609 4940
rect 3624 4928 3727 4940
rect 3739 4930 3765 4956
rect 3780 4951 3810 4962
rect 3842 4958 3904 4974
rect 3842 4956 3888 4958
rect 3842 4940 3904 4956
rect 3916 4940 3922 4988
rect 3925 4980 4005 4988
rect 3925 4978 3944 4980
rect 3959 4978 3993 4980
rect 3925 4962 4005 4978
rect 3925 4940 3944 4962
rect 3959 4946 3989 4962
rect 4017 4956 4023 5030
rect 4026 4956 4045 5100
rect 4060 4956 4066 5100
rect 4075 5030 4088 5100
rect 4140 5096 4162 5100
rect 4133 5074 4162 5088
rect 4215 5074 4231 5088
rect 4269 5084 4275 5086
rect 4282 5084 4390 5100
rect 4397 5084 4403 5086
rect 4411 5084 4426 5100
rect 4492 5094 4511 5097
rect 4133 5072 4231 5074
rect 4258 5072 4426 5084
rect 4441 5074 4457 5088
rect 4492 5075 4514 5094
rect 4524 5088 4540 5089
rect 4523 5086 4540 5088
rect 4524 5081 4540 5086
rect 4514 5074 4520 5075
rect 4523 5074 4552 5081
rect 4441 5073 4552 5074
rect 4441 5072 4558 5073
rect 4117 5064 4168 5072
rect 4215 5064 4249 5072
rect 4117 5052 4142 5064
rect 4149 5052 4168 5064
rect 4222 5062 4249 5064
rect 4258 5062 4479 5072
rect 4514 5069 4520 5072
rect 4222 5058 4479 5062
rect 4117 5044 4168 5052
rect 4215 5044 4479 5058
rect 4523 5064 4558 5072
rect 4069 4996 4088 5030
rect 4133 5036 4162 5044
rect 4133 5030 4150 5036
rect 4133 5028 4167 5030
rect 4215 5028 4231 5044
rect 4232 5034 4440 5044
rect 4441 5034 4457 5044
rect 4505 5040 4520 5055
rect 4523 5052 4524 5064
rect 4531 5052 4558 5064
rect 4523 5044 4558 5052
rect 4523 5043 4552 5044
rect 4243 5030 4457 5034
rect 4258 5028 4457 5030
rect 4492 5030 4505 5040
rect 4523 5030 4540 5043
rect 4492 5028 4540 5030
rect 4134 5024 4167 5028
rect 4130 5022 4167 5024
rect 4130 5021 4197 5022
rect 4130 5016 4161 5021
rect 4167 5016 4197 5021
rect 4130 5012 4197 5016
rect 4103 5009 4197 5012
rect 4103 5002 4152 5009
rect 4103 4996 4133 5002
rect 4152 4997 4157 5002
rect 4069 4980 4149 4996
rect 4161 4988 4197 5009
rect 4258 5004 4447 5028
rect 4492 5027 4539 5028
rect 4505 5022 4539 5027
rect 4273 5001 4447 5004
rect 4266 4998 4447 5001
rect 4475 5021 4539 5022
rect 4069 4978 4088 4980
rect 4103 4978 4137 4980
rect 4069 4962 4149 4978
rect 4069 4956 4088 4962
rect 3785 4930 3888 4940
rect 3739 4928 3888 4930
rect 3909 4928 3944 4940
rect 3578 4926 3740 4928
rect 3590 4906 3609 4926
rect 3624 4924 3654 4926
rect 3473 4898 3514 4906
rect 3596 4902 3609 4906
rect 3661 4910 3740 4926
rect 3772 4926 3944 4928
rect 3772 4910 3851 4926
rect 3858 4924 3888 4926
rect 3436 4888 3465 4898
rect 3479 4888 3508 4898
rect 3523 4888 3553 4902
rect 3596 4888 3639 4902
rect 3661 4898 3851 4910
rect 3916 4906 3922 4926
rect 3646 4888 3676 4898
rect 3677 4888 3835 4898
rect 3839 4888 3869 4898
rect 3873 4888 3903 4902
rect 3931 4888 3944 4926
rect 4016 4940 4045 4956
rect 4059 4940 4088 4956
rect 4103 4946 4133 4962
rect 4161 4940 4167 4988
rect 4170 4982 4189 4988
rect 4204 4982 4234 4990
rect 4170 4974 4234 4982
rect 4170 4958 4250 4974
rect 4266 4967 4328 4998
rect 4344 4967 4406 4998
rect 4475 4996 4524 5021
rect 4539 4996 4569 5012
rect 4438 4982 4468 4990
rect 4475 4988 4585 4996
rect 4438 4974 4483 4982
rect 4170 4956 4189 4958
rect 4204 4956 4250 4958
rect 4170 4940 4250 4956
rect 4277 4954 4312 4967
rect 4353 4964 4390 4967
rect 4353 4962 4395 4964
rect 4282 4951 4312 4954
rect 4291 4947 4298 4951
rect 4298 4946 4299 4947
rect 4257 4940 4267 4946
rect 4016 4932 4051 4940
rect 4016 4906 4017 4932
rect 4024 4906 4051 4932
rect 3959 4888 3989 4902
rect 4016 4898 4051 4906
rect 4053 4932 4094 4940
rect 4053 4906 4068 4932
rect 4075 4906 4094 4932
rect 4158 4928 4189 4940
rect 4204 4928 4307 4940
rect 4319 4930 4345 4956
rect 4360 4951 4390 4962
rect 4422 4958 4484 4974
rect 4422 4956 4468 4958
rect 4422 4940 4484 4956
rect 4496 4940 4502 4988
rect 4505 4980 4585 4988
rect 4505 4978 4524 4980
rect 4539 4978 4573 4980
rect 4505 4962 4585 4978
rect 4505 4940 4524 4962
rect 4539 4946 4569 4962
rect 4597 4956 4603 5030
rect 4606 4956 4625 5100
rect 4640 4956 4646 5100
rect 4655 5030 4668 5100
rect 4720 5096 4742 5100
rect 4713 5074 4742 5088
rect 4795 5074 4811 5088
rect 4849 5084 4855 5086
rect 4862 5084 4970 5100
rect 4977 5084 4983 5086
rect 4991 5084 5006 5100
rect 5072 5094 5091 5097
rect 4713 5072 4811 5074
rect 4838 5072 5006 5084
rect 5021 5074 5037 5088
rect 5072 5075 5094 5094
rect 5104 5088 5120 5089
rect 5103 5086 5120 5088
rect 5104 5081 5120 5086
rect 5094 5074 5100 5075
rect 5103 5074 5132 5081
rect 5021 5073 5132 5074
rect 5021 5072 5138 5073
rect 4697 5064 4748 5072
rect 4795 5064 4829 5072
rect 4697 5052 4722 5064
rect 4729 5052 4748 5064
rect 4802 5062 4829 5064
rect 4838 5062 5059 5072
rect 5094 5069 5100 5072
rect 4802 5058 5059 5062
rect 4697 5044 4748 5052
rect 4795 5044 5059 5058
rect 5103 5064 5138 5072
rect 4649 4996 4668 5030
rect 4713 5036 4742 5044
rect 4713 5030 4730 5036
rect 4713 5028 4747 5030
rect 4795 5028 4811 5044
rect 4812 5034 5020 5044
rect 5021 5034 5037 5044
rect 5085 5040 5100 5055
rect 5103 5052 5104 5064
rect 5111 5052 5138 5064
rect 5103 5044 5138 5052
rect 5103 5043 5132 5044
rect 4823 5030 5037 5034
rect 4838 5028 5037 5030
rect 5072 5030 5085 5040
rect 5103 5030 5120 5043
rect 5072 5028 5120 5030
rect 4714 5024 4747 5028
rect 4710 5022 4747 5024
rect 4710 5021 4777 5022
rect 4710 5016 4741 5021
rect 4747 5016 4777 5021
rect 4710 5012 4777 5016
rect 4683 5009 4777 5012
rect 4683 5002 4732 5009
rect 4683 4996 4713 5002
rect 4732 4997 4737 5002
rect 4649 4980 4729 4996
rect 4741 4988 4777 5009
rect 4838 5004 5027 5028
rect 5072 5027 5119 5028
rect 5085 5022 5119 5027
rect 4853 5001 5027 5004
rect 4846 4998 5027 5001
rect 5055 5021 5119 5022
rect 4649 4978 4668 4980
rect 4683 4978 4717 4980
rect 4649 4962 4729 4978
rect 4649 4956 4668 4962
rect 4365 4930 4468 4940
rect 4319 4928 4468 4930
rect 4489 4928 4524 4940
rect 4158 4926 4320 4928
rect 4170 4906 4189 4926
rect 4204 4924 4234 4926
rect 4053 4898 4094 4906
rect 4176 4902 4189 4906
rect 4241 4910 4320 4926
rect 4352 4926 4524 4928
rect 4352 4910 4431 4926
rect 4438 4924 4468 4926
rect 4016 4888 4045 4898
rect 4059 4888 4088 4898
rect 4103 4888 4133 4902
rect 4176 4888 4219 4902
rect 4241 4898 4431 4910
rect 4496 4906 4502 4926
rect 4226 4888 4256 4898
rect 4257 4888 4415 4898
rect 4419 4888 4449 4898
rect 4453 4888 4483 4902
rect 4511 4888 4524 4926
rect 4596 4940 4625 4956
rect 4639 4940 4668 4956
rect 4683 4946 4713 4962
rect 4741 4940 4747 4988
rect 4750 4982 4769 4988
rect 4784 4982 4814 4990
rect 4750 4974 4814 4982
rect 4750 4958 4830 4974
rect 4846 4967 4908 4998
rect 4924 4967 4986 4998
rect 5055 4996 5104 5021
rect 5119 4996 5149 5012
rect 5018 4982 5048 4990
rect 5055 4988 5165 4996
rect 5018 4974 5063 4982
rect 4750 4956 4769 4958
rect 4784 4956 4830 4958
rect 4750 4940 4830 4956
rect 4857 4954 4892 4967
rect 4933 4964 4970 4967
rect 4933 4962 4975 4964
rect 4862 4951 4892 4954
rect 4871 4947 4878 4951
rect 4878 4946 4879 4947
rect 4837 4940 4847 4946
rect 4596 4932 4631 4940
rect 4596 4906 4597 4932
rect 4604 4906 4631 4932
rect 4539 4888 4569 4902
rect 4596 4898 4631 4906
rect 4633 4932 4674 4940
rect 4633 4906 4648 4932
rect 4655 4906 4674 4932
rect 4738 4928 4769 4940
rect 4784 4928 4887 4940
rect 4899 4930 4925 4956
rect 4940 4951 4970 4962
rect 5002 4958 5064 4974
rect 5002 4956 5048 4958
rect 5002 4940 5064 4956
rect 5076 4940 5082 4988
rect 5085 4980 5165 4988
rect 5085 4978 5104 4980
rect 5119 4978 5153 4980
rect 5085 4962 5165 4978
rect 5085 4940 5104 4962
rect 5119 4946 5149 4962
rect 5177 4956 5183 5030
rect 5186 4956 5205 5100
rect 5220 4956 5226 5100
rect 5235 5030 5248 5100
rect 5300 5096 5322 5100
rect 5293 5074 5322 5088
rect 5375 5074 5391 5088
rect 5429 5084 5435 5086
rect 5442 5084 5550 5100
rect 5557 5084 5563 5086
rect 5571 5084 5586 5100
rect 5652 5094 5671 5097
rect 5293 5072 5391 5074
rect 5418 5072 5586 5084
rect 5601 5074 5617 5088
rect 5652 5075 5674 5094
rect 5684 5088 5700 5089
rect 5683 5086 5700 5088
rect 5684 5081 5700 5086
rect 5674 5074 5680 5075
rect 5683 5074 5712 5081
rect 5601 5073 5712 5074
rect 5601 5072 5718 5073
rect 5277 5064 5328 5072
rect 5375 5064 5409 5072
rect 5277 5052 5302 5064
rect 5309 5052 5328 5064
rect 5382 5062 5409 5064
rect 5418 5062 5639 5072
rect 5674 5069 5680 5072
rect 5382 5058 5639 5062
rect 5277 5044 5328 5052
rect 5375 5044 5639 5058
rect 5683 5064 5718 5072
rect 5229 4996 5248 5030
rect 5293 5036 5322 5044
rect 5293 5030 5310 5036
rect 5293 5028 5327 5030
rect 5375 5028 5391 5044
rect 5392 5034 5600 5044
rect 5601 5034 5617 5044
rect 5665 5040 5680 5055
rect 5683 5052 5684 5064
rect 5691 5052 5718 5064
rect 5683 5044 5718 5052
rect 5683 5043 5712 5044
rect 5403 5030 5617 5034
rect 5418 5028 5617 5030
rect 5652 5030 5665 5040
rect 5683 5030 5700 5043
rect 5652 5028 5700 5030
rect 5294 5024 5327 5028
rect 5290 5022 5327 5024
rect 5290 5021 5357 5022
rect 5290 5016 5321 5021
rect 5327 5016 5357 5021
rect 5290 5012 5357 5016
rect 5263 5009 5357 5012
rect 5263 5002 5312 5009
rect 5263 4996 5293 5002
rect 5312 4997 5317 5002
rect 5229 4980 5309 4996
rect 5321 4988 5357 5009
rect 5418 5004 5607 5028
rect 5652 5027 5699 5028
rect 5665 5022 5699 5027
rect 5433 5001 5607 5004
rect 5426 4998 5607 5001
rect 5635 5021 5699 5022
rect 5229 4978 5248 4980
rect 5263 4978 5297 4980
rect 5229 4962 5309 4978
rect 5229 4956 5248 4962
rect 4945 4930 5048 4940
rect 4899 4928 5048 4930
rect 5069 4928 5104 4940
rect 4738 4926 4900 4928
rect 4750 4906 4769 4926
rect 4784 4924 4814 4926
rect 4633 4898 4674 4906
rect 4756 4902 4769 4906
rect 4821 4910 4900 4926
rect 4932 4926 5104 4928
rect 4932 4910 5011 4926
rect 5018 4924 5048 4926
rect 4596 4888 4625 4898
rect 4639 4888 4668 4898
rect 4683 4888 4713 4902
rect 4756 4888 4799 4902
rect 4821 4898 5011 4910
rect 5076 4906 5082 4926
rect 4806 4888 4836 4898
rect 4837 4888 4995 4898
rect 4999 4888 5029 4898
rect 5033 4888 5063 4902
rect 5091 4888 5104 4926
rect 5176 4940 5205 4956
rect 5219 4940 5248 4956
rect 5263 4946 5293 4962
rect 5321 4940 5327 4988
rect 5330 4982 5349 4988
rect 5364 4982 5394 4990
rect 5330 4974 5394 4982
rect 5330 4958 5410 4974
rect 5426 4967 5488 4998
rect 5504 4967 5566 4998
rect 5635 4996 5684 5021
rect 5699 4996 5729 5012
rect 5598 4982 5628 4990
rect 5635 4988 5745 4996
rect 5598 4974 5643 4982
rect 5330 4956 5349 4958
rect 5364 4956 5410 4958
rect 5330 4940 5410 4956
rect 5437 4954 5472 4967
rect 5513 4964 5550 4967
rect 5513 4962 5555 4964
rect 5442 4951 5472 4954
rect 5451 4947 5458 4951
rect 5458 4946 5459 4947
rect 5417 4940 5427 4946
rect 5176 4932 5211 4940
rect 5176 4906 5177 4932
rect 5184 4906 5211 4932
rect 5119 4888 5149 4902
rect 5176 4898 5211 4906
rect 5213 4932 5254 4940
rect 5213 4906 5228 4932
rect 5235 4906 5254 4932
rect 5318 4928 5349 4940
rect 5364 4928 5467 4940
rect 5479 4930 5505 4956
rect 5520 4951 5550 4962
rect 5582 4958 5644 4974
rect 5582 4956 5628 4958
rect 5582 4940 5644 4956
rect 5656 4940 5662 4988
rect 5665 4980 5745 4988
rect 5665 4978 5684 4980
rect 5699 4978 5733 4980
rect 5665 4962 5745 4978
rect 5665 4940 5684 4962
rect 5699 4946 5729 4962
rect 5757 4956 5763 5030
rect 5766 4956 5785 5100
rect 5800 4956 5806 5100
rect 5815 5030 5828 5100
rect 5880 5096 5902 5100
rect 5873 5074 5902 5088
rect 5955 5074 5971 5088
rect 6009 5084 6015 5086
rect 6022 5084 6130 5100
rect 6137 5084 6143 5086
rect 6151 5084 6166 5100
rect 6232 5094 6251 5097
rect 5873 5072 5971 5074
rect 5998 5072 6166 5084
rect 6181 5074 6197 5088
rect 6232 5075 6254 5094
rect 6264 5088 6280 5089
rect 6263 5086 6280 5088
rect 6264 5081 6280 5086
rect 6254 5074 6260 5075
rect 6263 5074 6292 5081
rect 6181 5073 6292 5074
rect 6181 5072 6298 5073
rect 5857 5064 5908 5072
rect 5955 5064 5989 5072
rect 5857 5052 5882 5064
rect 5889 5052 5908 5064
rect 5962 5062 5989 5064
rect 5998 5062 6219 5072
rect 6254 5069 6260 5072
rect 5962 5058 6219 5062
rect 5857 5044 5908 5052
rect 5955 5044 6219 5058
rect 6263 5064 6298 5072
rect 5809 4996 5828 5030
rect 5873 5036 5902 5044
rect 5873 5030 5890 5036
rect 5873 5028 5907 5030
rect 5955 5028 5971 5044
rect 5972 5034 6180 5044
rect 6181 5034 6197 5044
rect 6245 5040 6260 5055
rect 6263 5052 6264 5064
rect 6271 5052 6298 5064
rect 6263 5044 6298 5052
rect 6263 5043 6292 5044
rect 5983 5030 6197 5034
rect 5998 5028 6197 5030
rect 6232 5030 6245 5040
rect 6263 5030 6280 5043
rect 6232 5028 6280 5030
rect 5874 5024 5907 5028
rect 5870 5022 5907 5024
rect 5870 5021 5937 5022
rect 5870 5016 5901 5021
rect 5907 5016 5937 5021
rect 5870 5012 5937 5016
rect 5843 5009 5937 5012
rect 5843 5002 5892 5009
rect 5843 4996 5873 5002
rect 5892 4997 5897 5002
rect 5809 4980 5889 4996
rect 5901 4988 5937 5009
rect 5998 5004 6187 5028
rect 6232 5027 6279 5028
rect 6245 5022 6279 5027
rect 6013 5001 6187 5004
rect 6006 4998 6187 5001
rect 6215 5021 6279 5022
rect 5809 4978 5828 4980
rect 5843 4978 5877 4980
rect 5809 4962 5889 4978
rect 5809 4956 5828 4962
rect 5525 4930 5628 4940
rect 5479 4928 5628 4930
rect 5649 4928 5684 4940
rect 5318 4926 5480 4928
rect 5330 4906 5349 4926
rect 5364 4924 5394 4926
rect 5213 4898 5254 4906
rect 5336 4902 5349 4906
rect 5401 4910 5480 4926
rect 5512 4926 5684 4928
rect 5512 4910 5591 4926
rect 5598 4924 5628 4926
rect 5176 4888 5205 4898
rect 5219 4888 5248 4898
rect 5263 4888 5293 4902
rect 5336 4888 5379 4902
rect 5401 4898 5591 4910
rect 5656 4906 5662 4926
rect 5386 4888 5416 4898
rect 5417 4888 5575 4898
rect 5579 4888 5609 4898
rect 5613 4888 5643 4902
rect 5671 4888 5684 4926
rect 5756 4940 5785 4956
rect 5799 4940 5828 4956
rect 5843 4946 5873 4962
rect 5901 4940 5907 4988
rect 5910 4982 5929 4988
rect 5944 4982 5974 4990
rect 5910 4974 5974 4982
rect 5910 4958 5990 4974
rect 6006 4967 6068 4998
rect 6084 4967 6146 4998
rect 6215 4996 6264 5021
rect 6279 4996 6309 5012
rect 6178 4982 6208 4990
rect 6215 4988 6325 4996
rect 6178 4974 6223 4982
rect 5910 4956 5929 4958
rect 5944 4956 5990 4958
rect 5910 4940 5990 4956
rect 6017 4954 6052 4967
rect 6093 4964 6130 4967
rect 6093 4962 6135 4964
rect 6022 4951 6052 4954
rect 6031 4947 6038 4951
rect 6038 4946 6039 4947
rect 5997 4940 6007 4946
rect 5756 4932 5791 4940
rect 5756 4906 5757 4932
rect 5764 4906 5791 4932
rect 5699 4888 5729 4902
rect 5756 4898 5791 4906
rect 5793 4932 5834 4940
rect 5793 4906 5808 4932
rect 5815 4906 5834 4932
rect 5898 4928 5929 4940
rect 5944 4928 6047 4940
rect 6059 4930 6085 4956
rect 6100 4951 6130 4962
rect 6162 4958 6224 4974
rect 6162 4956 6208 4958
rect 6162 4940 6224 4956
rect 6236 4940 6242 4988
rect 6245 4980 6325 4988
rect 6245 4978 6264 4980
rect 6279 4978 6313 4980
rect 6245 4962 6325 4978
rect 6245 4940 6264 4962
rect 6279 4946 6309 4962
rect 6337 4956 6343 5030
rect 6346 4956 6365 5100
rect 6380 4956 6386 5100
rect 6395 5030 6408 5100
rect 6460 5096 6482 5100
rect 6453 5074 6482 5088
rect 6535 5074 6551 5088
rect 6589 5084 6595 5086
rect 6602 5084 6710 5100
rect 6717 5084 6723 5086
rect 6731 5084 6746 5100
rect 6812 5094 6831 5097
rect 6453 5072 6551 5074
rect 6578 5072 6746 5084
rect 6761 5074 6777 5088
rect 6812 5075 6834 5094
rect 6844 5088 6860 5089
rect 6843 5086 6860 5088
rect 6844 5081 6860 5086
rect 6834 5074 6840 5075
rect 6843 5074 6872 5081
rect 6761 5073 6872 5074
rect 6761 5072 6878 5073
rect 6437 5064 6488 5072
rect 6535 5064 6569 5072
rect 6437 5052 6462 5064
rect 6469 5052 6488 5064
rect 6542 5062 6569 5064
rect 6578 5062 6799 5072
rect 6834 5069 6840 5072
rect 6542 5058 6799 5062
rect 6437 5044 6488 5052
rect 6535 5044 6799 5058
rect 6843 5064 6878 5072
rect 6389 4996 6408 5030
rect 6453 5036 6482 5044
rect 6453 5030 6470 5036
rect 6453 5028 6487 5030
rect 6535 5028 6551 5044
rect 6552 5034 6760 5044
rect 6761 5034 6777 5044
rect 6825 5040 6840 5055
rect 6843 5052 6844 5064
rect 6851 5052 6878 5064
rect 6843 5044 6878 5052
rect 6843 5043 6872 5044
rect 6563 5030 6777 5034
rect 6578 5028 6777 5030
rect 6812 5030 6825 5040
rect 6843 5030 6860 5043
rect 6812 5028 6860 5030
rect 6454 5024 6487 5028
rect 6450 5022 6487 5024
rect 6450 5021 6517 5022
rect 6450 5016 6481 5021
rect 6487 5016 6517 5021
rect 6450 5012 6517 5016
rect 6423 5009 6517 5012
rect 6423 5002 6472 5009
rect 6423 4996 6453 5002
rect 6472 4997 6477 5002
rect 6389 4980 6469 4996
rect 6481 4988 6517 5009
rect 6578 5004 6767 5028
rect 6812 5027 6859 5028
rect 6825 5022 6859 5027
rect 6593 5001 6767 5004
rect 6586 4998 6767 5001
rect 6795 5021 6859 5022
rect 6389 4978 6408 4980
rect 6423 4978 6457 4980
rect 6389 4962 6469 4978
rect 6389 4956 6408 4962
rect 6105 4930 6208 4940
rect 6059 4928 6208 4930
rect 6229 4928 6264 4940
rect 5898 4926 6060 4928
rect 5910 4906 5929 4926
rect 5944 4924 5974 4926
rect 5793 4898 5834 4906
rect 5916 4902 5929 4906
rect 5981 4910 6060 4926
rect 6092 4926 6264 4928
rect 6092 4910 6171 4926
rect 6178 4924 6208 4926
rect 5756 4888 5785 4898
rect 5799 4888 5828 4898
rect 5843 4888 5873 4902
rect 5916 4888 5959 4902
rect 5981 4898 6171 4910
rect 6236 4906 6242 4926
rect 5966 4888 5996 4898
rect 5997 4888 6155 4898
rect 6159 4888 6189 4898
rect 6193 4888 6223 4902
rect 6251 4888 6264 4926
rect 6336 4940 6365 4956
rect 6379 4940 6408 4956
rect 6423 4946 6453 4962
rect 6481 4940 6487 4988
rect 6490 4982 6509 4988
rect 6524 4982 6554 4990
rect 6490 4974 6554 4982
rect 6490 4958 6570 4974
rect 6586 4967 6648 4998
rect 6664 4967 6726 4998
rect 6795 4996 6844 5021
rect 6859 4996 6889 5012
rect 6758 4982 6788 4990
rect 6795 4988 6905 4996
rect 6758 4974 6803 4982
rect 6490 4956 6509 4958
rect 6524 4956 6570 4958
rect 6490 4940 6570 4956
rect 6597 4954 6632 4967
rect 6673 4964 6710 4967
rect 6673 4962 6715 4964
rect 6602 4951 6632 4954
rect 6611 4947 6618 4951
rect 6618 4946 6619 4947
rect 6577 4940 6587 4946
rect 6336 4932 6371 4940
rect 6336 4906 6337 4932
rect 6344 4906 6371 4932
rect 6279 4888 6309 4902
rect 6336 4898 6371 4906
rect 6373 4932 6414 4940
rect 6373 4906 6388 4932
rect 6395 4906 6414 4932
rect 6478 4928 6509 4940
rect 6524 4928 6627 4940
rect 6639 4930 6665 4956
rect 6680 4951 6710 4962
rect 6742 4958 6804 4974
rect 6742 4956 6788 4958
rect 6742 4940 6804 4956
rect 6816 4940 6822 4988
rect 6825 4980 6905 4988
rect 6825 4978 6844 4980
rect 6859 4978 6893 4980
rect 6825 4962 6905 4978
rect 6825 4940 6844 4962
rect 6859 4946 6889 4962
rect 6917 4956 6923 5030
rect 6926 4956 6945 5100
rect 6960 4956 6966 5100
rect 6975 5030 6988 5100
rect 7040 5096 7062 5100
rect 7033 5074 7062 5088
rect 7115 5074 7131 5088
rect 7169 5084 7175 5086
rect 7182 5084 7290 5100
rect 7297 5084 7303 5086
rect 7311 5084 7326 5100
rect 7392 5094 7411 5097
rect 7033 5072 7131 5074
rect 7158 5072 7326 5084
rect 7341 5074 7357 5088
rect 7392 5075 7414 5094
rect 7424 5088 7440 5089
rect 7423 5086 7440 5088
rect 7424 5081 7440 5086
rect 7414 5074 7420 5075
rect 7423 5074 7452 5081
rect 7341 5073 7452 5074
rect 7341 5072 7458 5073
rect 7017 5064 7068 5072
rect 7115 5064 7149 5072
rect 7017 5052 7042 5064
rect 7049 5052 7068 5064
rect 7122 5062 7149 5064
rect 7158 5062 7379 5072
rect 7414 5069 7420 5072
rect 7122 5058 7379 5062
rect 7017 5044 7068 5052
rect 7115 5044 7379 5058
rect 7423 5064 7458 5072
rect 6969 4996 6988 5030
rect 7033 5036 7062 5044
rect 7033 5030 7050 5036
rect 7033 5028 7067 5030
rect 7115 5028 7131 5044
rect 7132 5034 7340 5044
rect 7341 5034 7357 5044
rect 7405 5040 7420 5055
rect 7423 5052 7424 5064
rect 7431 5052 7458 5064
rect 7423 5044 7458 5052
rect 7423 5043 7452 5044
rect 7143 5030 7357 5034
rect 7158 5028 7357 5030
rect 7392 5030 7405 5040
rect 7423 5030 7440 5043
rect 7392 5028 7440 5030
rect 7034 5024 7067 5028
rect 7030 5022 7067 5024
rect 7030 5021 7097 5022
rect 7030 5016 7061 5021
rect 7067 5016 7097 5021
rect 7030 5012 7097 5016
rect 7003 5009 7097 5012
rect 7003 5002 7052 5009
rect 7003 4996 7033 5002
rect 7052 4997 7057 5002
rect 6969 4980 7049 4996
rect 7061 4988 7097 5009
rect 7158 5004 7347 5028
rect 7392 5027 7439 5028
rect 7405 5022 7439 5027
rect 7173 5001 7347 5004
rect 7166 4998 7347 5001
rect 7375 5021 7439 5022
rect 6969 4978 6988 4980
rect 7003 4978 7037 4980
rect 6969 4962 7049 4978
rect 6969 4956 6988 4962
rect 6685 4930 6788 4940
rect 6639 4928 6788 4930
rect 6809 4928 6844 4940
rect 6478 4926 6640 4928
rect 6490 4906 6509 4926
rect 6524 4924 6554 4926
rect 6373 4898 6414 4906
rect 6496 4902 6509 4906
rect 6561 4910 6640 4926
rect 6672 4926 6844 4928
rect 6672 4910 6751 4926
rect 6758 4924 6788 4926
rect 6336 4888 6365 4898
rect 6379 4888 6408 4898
rect 6423 4888 6453 4902
rect 6496 4888 6539 4902
rect 6561 4898 6751 4910
rect 6816 4906 6822 4926
rect 6546 4888 6576 4898
rect 6577 4888 6735 4898
rect 6739 4888 6769 4898
rect 6773 4888 6803 4902
rect 6831 4888 6844 4926
rect 6916 4940 6945 4956
rect 6959 4940 6988 4956
rect 7003 4946 7033 4962
rect 7061 4940 7067 4988
rect 7070 4982 7089 4988
rect 7104 4982 7134 4990
rect 7070 4974 7134 4982
rect 7070 4958 7150 4974
rect 7166 4967 7228 4998
rect 7244 4967 7306 4998
rect 7375 4996 7424 5021
rect 7439 4996 7469 5012
rect 7338 4982 7368 4990
rect 7375 4988 7485 4996
rect 7338 4974 7383 4982
rect 7070 4956 7089 4958
rect 7104 4956 7150 4958
rect 7070 4940 7150 4956
rect 7177 4954 7212 4967
rect 7253 4964 7290 4967
rect 7253 4962 7295 4964
rect 7182 4951 7212 4954
rect 7191 4947 7198 4951
rect 7198 4946 7199 4947
rect 7157 4940 7167 4946
rect 6916 4932 6951 4940
rect 6916 4906 6917 4932
rect 6924 4906 6951 4932
rect 6859 4888 6889 4902
rect 6916 4898 6951 4906
rect 6953 4932 6994 4940
rect 6953 4906 6968 4932
rect 6975 4906 6994 4932
rect 7058 4928 7089 4940
rect 7104 4928 7207 4940
rect 7219 4930 7245 4956
rect 7260 4951 7290 4962
rect 7322 4958 7384 4974
rect 7322 4956 7368 4958
rect 7322 4940 7384 4956
rect 7396 4940 7402 4988
rect 7405 4980 7485 4988
rect 7405 4978 7424 4980
rect 7439 4978 7473 4980
rect 7405 4962 7485 4978
rect 7405 4940 7424 4962
rect 7439 4946 7469 4962
rect 7497 4956 7503 5030
rect 7506 4956 7525 5100
rect 7540 4956 7546 5100
rect 7555 5030 7568 5100
rect 7613 5078 7614 5088
rect 7629 5078 7642 5088
rect 7613 5074 7642 5078
rect 7647 5074 7677 5100
rect 7695 5086 7711 5088
rect 7783 5086 7836 5100
rect 7784 5084 7848 5086
rect 7891 5084 7906 5100
rect 7955 5097 7985 5100
rect 7955 5094 7991 5097
rect 7921 5086 7937 5088
rect 7695 5074 7710 5078
rect 7613 5072 7710 5074
rect 7738 5072 7906 5084
rect 7922 5074 7937 5078
rect 7955 5075 7994 5094
rect 8013 5088 8020 5089
rect 8019 5081 8020 5088
rect 8003 5078 8004 5081
rect 8019 5078 8032 5081
rect 7955 5074 7985 5075
rect 7994 5074 8000 5075
rect 8003 5074 8032 5078
rect 7922 5073 8032 5074
rect 7922 5072 8038 5073
rect 7597 5064 7648 5072
rect 7597 5052 7622 5064
rect 7629 5052 7648 5064
rect 7679 5064 7729 5072
rect 7679 5056 7695 5064
rect 7702 5062 7729 5064
rect 7738 5062 7959 5072
rect 7702 5052 7959 5062
rect 7988 5064 8038 5072
rect 7988 5055 8004 5064
rect 7597 5044 7648 5052
rect 7695 5044 7959 5052
rect 7985 5052 8004 5055
rect 8011 5052 8038 5064
rect 7985 5044 8038 5052
rect 7549 4996 7568 5030
rect 7613 5036 7614 5044
rect 7629 5036 7642 5044
rect 7613 5028 7629 5036
rect 7610 5021 7629 5024
rect 7610 5012 7632 5021
rect 7583 5002 7632 5012
rect 7583 4996 7613 5002
rect 7632 4997 7637 5002
rect 7549 4980 7629 4996
rect 7647 4988 7677 5044
rect 7712 5034 7920 5044
rect 7955 5040 8000 5044
rect 8003 5043 8004 5044
rect 8019 5043 8032 5044
rect 7738 5004 7927 5034
rect 7753 5001 7927 5004
rect 7746 4998 7927 5001
rect 7549 4978 7568 4980
rect 7583 4978 7617 4980
rect 7549 4962 7629 4978
rect 7656 4974 7669 4988
rect 7684 4974 7700 4990
rect 7746 4985 7757 4998
rect 7549 4956 7568 4962
rect 7265 4930 7368 4940
rect 7219 4928 7368 4930
rect 7389 4928 7424 4940
rect 7058 4926 7220 4928
rect 7070 4906 7089 4926
rect 7104 4924 7134 4926
rect 6953 4898 6994 4906
rect 7076 4902 7089 4906
rect 7141 4910 7220 4926
rect 7252 4926 7424 4928
rect 7252 4910 7331 4926
rect 7338 4924 7368 4926
rect 6916 4888 6945 4898
rect 6959 4888 6988 4898
rect 7003 4888 7033 4902
rect 7076 4888 7119 4902
rect 7141 4898 7331 4910
rect 7396 4906 7402 4926
rect 7126 4888 7156 4898
rect 7157 4888 7315 4898
rect 7319 4888 7349 4898
rect 7353 4888 7383 4902
rect 7411 4888 7424 4926
rect 7496 4940 7525 4956
rect 7539 4940 7568 4956
rect 7583 4940 7613 4962
rect 7656 4958 7718 4974
rect 7746 4967 7757 4983
rect 7762 4978 7772 4998
rect 7782 4978 7796 4998
rect 7799 4985 7808 4998
rect 7824 4985 7833 4998
rect 7762 4967 7796 4978
rect 7799 4967 7808 4983
rect 7824 4967 7833 4983
rect 7840 4978 7850 4998
rect 7860 4978 7874 4998
rect 7875 4985 7886 4998
rect 7840 4967 7874 4978
rect 7875 4967 7886 4983
rect 7932 4974 7948 4990
rect 7955 4988 7985 5040
rect 8019 5036 8020 5043
rect 8004 5028 8020 5036
rect 7991 4996 8004 5015
rect 8019 4996 8049 5012
rect 7991 4980 8065 4996
rect 7991 4978 8004 4980
rect 8019 4978 8053 4980
rect 7656 4956 7669 4958
rect 7684 4956 7718 4958
rect 7656 4940 7718 4956
rect 7762 4951 7778 4954
rect 7840 4951 7870 4962
rect 7918 4958 7964 4974
rect 7991 4962 8065 4978
rect 7918 4956 7952 4958
rect 7917 4940 7964 4956
rect 7991 4940 8004 4962
rect 8019 4940 8049 4962
rect 8076 4940 8077 4956
rect 8092 4940 8105 5100
rect 8135 4996 8148 5100
rect 8193 5078 8194 5088
rect 8209 5078 8222 5088
rect 8193 5074 8222 5078
rect 8227 5074 8257 5100
rect 8275 5086 8291 5088
rect 8363 5086 8416 5100
rect 8364 5084 8428 5086
rect 8471 5084 8486 5100
rect 8535 5097 8565 5100
rect 8535 5094 8571 5097
rect 8501 5086 8517 5088
rect 8275 5074 8290 5078
rect 8193 5072 8290 5074
rect 8318 5072 8486 5084
rect 8502 5074 8517 5078
rect 8535 5075 8574 5094
rect 8593 5088 8600 5089
rect 8599 5081 8600 5088
rect 8583 5078 8584 5081
rect 8599 5078 8612 5081
rect 8535 5074 8565 5075
rect 8574 5074 8580 5075
rect 8583 5074 8612 5078
rect 8502 5073 8612 5074
rect 8502 5072 8618 5073
rect 8177 5064 8228 5072
rect 8177 5052 8202 5064
rect 8209 5052 8228 5064
rect 8259 5064 8309 5072
rect 8259 5056 8275 5064
rect 8282 5062 8309 5064
rect 8318 5062 8539 5072
rect 8282 5052 8539 5062
rect 8568 5064 8618 5072
rect 8568 5055 8584 5064
rect 8177 5044 8228 5052
rect 8275 5044 8539 5052
rect 8565 5052 8584 5055
rect 8591 5052 8618 5064
rect 8565 5044 8618 5052
rect 8193 5036 8194 5044
rect 8209 5036 8222 5044
rect 8193 5028 8209 5036
rect 8190 5021 8209 5024
rect 8190 5012 8212 5021
rect 8163 5002 8212 5012
rect 8163 4996 8193 5002
rect 8212 4997 8217 5002
rect 8135 4980 8209 4996
rect 8227 4988 8257 5044
rect 8292 5034 8500 5044
rect 8535 5040 8580 5044
rect 8583 5043 8584 5044
rect 8599 5043 8612 5044
rect 8318 5004 8507 5034
rect 8333 5001 8507 5004
rect 8326 4998 8507 5001
rect 8135 4978 8148 4980
rect 8163 4978 8197 4980
rect 8135 4962 8209 4978
rect 8236 4974 8249 4988
rect 8264 4974 8280 4990
rect 8326 4985 8337 4998
rect 8119 4940 8120 4956
rect 8135 4940 8148 4962
rect 8163 4940 8193 4962
rect 8236 4958 8298 4974
rect 8326 4967 8337 4983
rect 8342 4978 8352 4998
rect 8362 4978 8376 4998
rect 8379 4985 8388 4998
rect 8404 4985 8413 4998
rect 8342 4967 8376 4978
rect 8379 4967 8388 4983
rect 8404 4967 8413 4983
rect 8420 4978 8430 4998
rect 8440 4978 8454 4998
rect 8455 4985 8466 4998
rect 8420 4967 8454 4978
rect 8455 4967 8466 4983
rect 8512 4974 8528 4990
rect 8535 4988 8565 5040
rect 8599 5036 8600 5043
rect 8584 5028 8600 5036
rect 8571 4996 8584 5015
rect 8599 4996 8629 5012
rect 8571 4980 8645 4996
rect 8571 4978 8584 4980
rect 8599 4978 8633 4980
rect 8236 4956 8249 4958
rect 8264 4956 8298 4958
rect 8236 4940 8298 4956
rect 8342 4951 8358 4954
rect 8420 4951 8450 4962
rect 8498 4958 8544 4974
rect 8571 4962 8645 4978
rect 8498 4956 8532 4958
rect 8497 4940 8544 4956
rect 8571 4940 8584 4962
rect 8599 4940 8629 4962
rect 8656 4940 8657 4956
rect 8672 4940 8685 5100
rect 8715 4996 8728 5100
rect 8773 5078 8774 5088
rect 8789 5078 8802 5088
rect 8773 5074 8802 5078
rect 8807 5074 8837 5100
rect 8855 5086 8871 5088
rect 8943 5086 8996 5100
rect 8944 5084 9008 5086
rect 9051 5084 9066 5100
rect 9115 5097 9145 5100
rect 9115 5094 9151 5097
rect 9081 5086 9097 5088
rect 8855 5074 8870 5078
rect 8773 5072 8870 5074
rect 8898 5072 9066 5084
rect 9082 5074 9097 5078
rect 9115 5075 9154 5094
rect 9173 5088 9180 5089
rect 9179 5081 9180 5088
rect 9163 5078 9164 5081
rect 9179 5078 9192 5081
rect 9115 5074 9145 5075
rect 9154 5074 9160 5075
rect 9163 5074 9192 5078
rect 9082 5073 9192 5074
rect 9082 5072 9198 5073
rect 8757 5064 8808 5072
rect 8757 5052 8782 5064
rect 8789 5052 8808 5064
rect 8839 5064 8889 5072
rect 8839 5056 8855 5064
rect 8862 5062 8889 5064
rect 8898 5062 9119 5072
rect 8862 5052 9119 5062
rect 9148 5064 9198 5072
rect 9148 5055 9164 5064
rect 8757 5044 8808 5052
rect 8855 5044 9119 5052
rect 9145 5052 9164 5055
rect 9171 5052 9198 5064
rect 9145 5044 9198 5052
rect 8773 5036 8774 5044
rect 8789 5036 8802 5044
rect 8773 5028 8789 5036
rect 8770 5021 8789 5024
rect 8770 5012 8792 5021
rect 8743 5002 8792 5012
rect 8743 4996 8773 5002
rect 8792 4997 8797 5002
rect 8715 4980 8789 4996
rect 8807 4988 8837 5044
rect 8872 5034 9080 5044
rect 9115 5040 9160 5044
rect 9163 5043 9164 5044
rect 9179 5043 9192 5044
rect 8898 5004 9087 5034
rect 8913 5001 9087 5004
rect 8906 4998 9087 5001
rect 8715 4978 8728 4980
rect 8743 4978 8777 4980
rect 8715 4962 8789 4978
rect 8816 4974 8829 4988
rect 8844 4974 8860 4990
rect 8906 4985 8917 4998
rect 8699 4940 8700 4956
rect 8715 4940 8728 4962
rect 8743 4940 8773 4962
rect 8816 4958 8878 4974
rect 8906 4967 8917 4983
rect 8922 4978 8932 4998
rect 8942 4978 8956 4998
rect 8959 4985 8968 4998
rect 8984 4985 8993 4998
rect 8922 4967 8956 4978
rect 8959 4967 8968 4983
rect 8984 4967 8993 4983
rect 9000 4978 9010 4998
rect 9020 4978 9034 4998
rect 9035 4985 9046 4998
rect 9000 4967 9034 4978
rect 9035 4967 9046 4983
rect 9092 4974 9108 4990
rect 9115 4988 9145 5040
rect 9179 5036 9180 5043
rect 9164 5028 9180 5036
rect 9151 4996 9164 5015
rect 9179 4996 9209 5012
rect 9151 4980 9225 4996
rect 9151 4978 9164 4980
rect 9179 4978 9213 4980
rect 8816 4956 8829 4958
rect 8844 4956 8878 4958
rect 8816 4940 8878 4956
rect 8922 4951 8938 4954
rect 9000 4951 9030 4962
rect 9078 4958 9124 4974
rect 9151 4962 9225 4978
rect 9078 4956 9112 4958
rect 9077 4940 9124 4956
rect 9151 4940 9164 4962
rect 9179 4940 9209 4962
rect 9236 4940 9237 4956
rect 9252 4940 9265 5100
rect 7496 4932 7531 4940
rect 7496 4906 7497 4932
rect 7504 4906 7531 4932
rect 7439 4888 7469 4902
rect 7496 4898 7531 4906
rect 7533 4932 7574 4940
rect 7533 4906 7548 4932
rect 7555 4906 7574 4932
rect 7638 4928 7700 4940
rect 7712 4928 7787 4940
rect 7845 4928 7920 4940
rect 7932 4928 7963 4940
rect 7969 4928 8004 4940
rect 7638 4926 7800 4928
rect 7533 4898 7574 4906
rect 7656 4902 7669 4926
rect 7684 4924 7699 4926
rect 7496 4888 7525 4898
rect 7539 4888 7568 4898
rect 7583 4888 7613 4902
rect 7656 4888 7699 4902
rect 7723 4899 7730 4906
rect 7733 4902 7800 4926
rect 7832 4926 8004 4928
rect 7802 4904 7830 4908
rect 7832 4904 7912 4926
rect 7933 4924 7948 4926
rect 7802 4902 7912 4904
rect 7733 4898 7912 4902
rect 7706 4888 7736 4898
rect 7738 4888 7891 4898
rect 7899 4888 7929 4898
rect 7933 4888 7963 4902
rect 7991 4888 8004 4926
rect 8076 4932 8111 4940
rect 8076 4906 8077 4932
rect 8084 4906 8111 4932
rect 8019 4888 8049 4902
rect 8076 4898 8111 4906
rect 8113 4932 8154 4940
rect 8113 4906 8128 4932
rect 8135 4906 8154 4932
rect 8218 4928 8280 4940
rect 8292 4928 8367 4940
rect 8425 4928 8500 4940
rect 8512 4928 8543 4940
rect 8549 4928 8584 4940
rect 8218 4926 8380 4928
rect 8113 4898 8154 4906
rect 8236 4902 8249 4926
rect 8264 4924 8279 4926
rect 8076 4888 8077 4898
rect 8092 4888 8105 4898
rect 8119 4888 8120 4898
rect 8135 4888 8148 4898
rect 8163 4888 8193 4902
rect 8236 4888 8279 4902
rect 8303 4899 8310 4906
rect 8313 4902 8380 4926
rect 8412 4926 8584 4928
rect 8382 4904 8410 4908
rect 8412 4904 8492 4926
rect 8513 4924 8528 4926
rect 8382 4902 8492 4904
rect 8313 4898 8492 4902
rect 8286 4888 8316 4898
rect 8318 4888 8471 4898
rect 8479 4888 8509 4898
rect 8513 4888 8543 4902
rect 8571 4888 8584 4926
rect 8656 4932 8691 4940
rect 8656 4906 8657 4932
rect 8664 4906 8691 4932
rect 8599 4888 8629 4902
rect 8656 4898 8691 4906
rect 8693 4932 8734 4940
rect 8693 4906 8708 4932
rect 8715 4906 8734 4932
rect 8798 4928 8860 4940
rect 8872 4928 8947 4940
rect 9005 4928 9080 4940
rect 9092 4928 9123 4940
rect 9129 4928 9164 4940
rect 8798 4926 8960 4928
rect 8693 4898 8734 4906
rect 8816 4902 8829 4926
rect 8844 4924 8859 4926
rect 8656 4888 8657 4898
rect 8672 4888 8685 4898
rect 8699 4888 8700 4898
rect 8715 4888 8728 4898
rect 8743 4888 8773 4902
rect 8816 4888 8859 4902
rect 8883 4899 8890 4906
rect 8893 4902 8960 4926
rect 8992 4926 9164 4928
rect 8962 4904 8990 4908
rect 8992 4904 9072 4926
rect 9093 4924 9108 4926
rect 8962 4902 9072 4904
rect 8893 4898 9072 4902
rect 8866 4888 8896 4898
rect 8898 4888 9051 4898
rect 9059 4888 9089 4898
rect 9093 4888 9123 4902
rect 9151 4888 9164 4926
rect 9236 4932 9271 4940
rect 9236 4906 9237 4932
rect 9244 4906 9271 4932
rect 9179 4888 9209 4902
rect 9236 4898 9271 4906
rect 9236 4888 9237 4898
rect 9252 4888 9265 4898
rect -1 4882 9265 4888
rect 0 4874 9265 4882
rect 15 4844 28 4874
rect 43 4860 73 4874
rect 116 4860 159 4874
rect 166 4860 386 4874
rect 393 4860 423 4874
rect 83 4846 98 4858
rect 117 4846 130 4860
rect 198 4856 351 4860
rect 80 4844 102 4846
rect 180 4844 372 4856
rect 451 4844 464 4874
rect 479 4860 509 4874
rect 546 4844 565 4874
rect 580 4844 586 4874
rect 595 4844 608 4874
rect 623 4860 653 4874
rect 696 4860 739 4874
rect 746 4860 966 4874
rect 973 4860 1003 4874
rect 663 4846 678 4858
rect 697 4846 710 4860
rect 778 4856 931 4860
rect 660 4844 682 4846
rect 760 4844 952 4856
rect 1031 4844 1044 4874
rect 1059 4860 1089 4874
rect 1126 4844 1145 4874
rect 1160 4844 1166 4874
rect 1175 4844 1188 4874
rect 1203 4860 1233 4874
rect 1276 4860 1319 4874
rect 1326 4860 1546 4874
rect 1553 4860 1583 4874
rect 1243 4846 1258 4858
rect 1277 4846 1290 4860
rect 1358 4856 1511 4860
rect 1240 4844 1262 4846
rect 1340 4844 1532 4856
rect 1611 4844 1624 4874
rect 1639 4860 1669 4874
rect 1706 4844 1725 4874
rect 1740 4844 1746 4874
rect 1755 4844 1768 4874
rect 1783 4860 1813 4874
rect 1856 4860 1899 4874
rect 1906 4860 2126 4874
rect 2133 4860 2163 4874
rect 1823 4846 1838 4858
rect 1857 4846 1870 4860
rect 1938 4856 2091 4860
rect 1820 4844 1842 4846
rect 1920 4844 2112 4856
rect 2191 4844 2204 4874
rect 2219 4860 2249 4874
rect 2286 4844 2305 4874
rect 2320 4844 2326 4874
rect 2335 4844 2348 4874
rect 2363 4860 2393 4874
rect 2436 4860 2479 4874
rect 2486 4860 2706 4874
rect 2713 4860 2743 4874
rect 2403 4846 2418 4858
rect 2437 4846 2450 4860
rect 2518 4856 2671 4860
rect 2400 4844 2422 4846
rect 2500 4844 2692 4856
rect 2771 4844 2784 4874
rect 2799 4860 2829 4874
rect 2866 4844 2885 4874
rect 2900 4844 2906 4874
rect 2915 4844 2928 4874
rect 2943 4860 2973 4874
rect 3016 4860 3059 4874
rect 3066 4860 3286 4874
rect 3293 4860 3323 4874
rect 2983 4846 2998 4858
rect 3017 4846 3030 4860
rect 3098 4856 3251 4860
rect 2980 4844 3002 4846
rect 3080 4844 3272 4856
rect 3351 4844 3364 4874
rect 3379 4860 3409 4874
rect 3446 4844 3465 4874
rect 3480 4844 3486 4874
rect 3495 4844 3508 4874
rect 3523 4860 3553 4874
rect 3596 4860 3639 4874
rect 3646 4860 3866 4874
rect 3873 4860 3903 4874
rect 3563 4846 3578 4858
rect 3597 4846 3610 4860
rect 3678 4856 3831 4860
rect 3560 4844 3582 4846
rect 3660 4844 3852 4856
rect 3931 4844 3944 4874
rect 3959 4860 3989 4874
rect 4026 4844 4045 4874
rect 4060 4844 4066 4874
rect 4075 4844 4088 4874
rect 4103 4860 4133 4874
rect 4176 4860 4219 4874
rect 4226 4860 4446 4874
rect 4453 4860 4483 4874
rect 4143 4846 4158 4858
rect 4177 4846 4190 4860
rect 4258 4856 4411 4860
rect 4140 4844 4162 4846
rect 4240 4844 4432 4856
rect 4511 4844 4524 4874
rect 4539 4860 4569 4874
rect 4606 4844 4625 4874
rect 4640 4844 4646 4874
rect 4655 4844 4668 4874
rect 4683 4860 4713 4874
rect 4756 4860 4799 4874
rect 4806 4860 5026 4874
rect 5033 4860 5063 4874
rect 4723 4846 4738 4858
rect 4757 4846 4770 4860
rect 4838 4856 4991 4860
rect 4720 4844 4742 4846
rect 4820 4844 5012 4856
rect 5091 4844 5104 4874
rect 5119 4860 5149 4874
rect 5186 4844 5205 4874
rect 5220 4844 5226 4874
rect 5235 4844 5248 4874
rect 5263 4860 5293 4874
rect 5336 4860 5379 4874
rect 5386 4860 5606 4874
rect 5613 4860 5643 4874
rect 5303 4846 5318 4858
rect 5337 4846 5350 4860
rect 5418 4856 5571 4860
rect 5300 4844 5322 4846
rect 5400 4844 5592 4856
rect 5671 4844 5684 4874
rect 5699 4860 5729 4874
rect 5766 4844 5785 4874
rect 5800 4844 5806 4874
rect 5815 4844 5828 4874
rect 5843 4860 5873 4874
rect 5916 4860 5959 4874
rect 5966 4860 6186 4874
rect 6193 4860 6223 4874
rect 5883 4846 5898 4858
rect 5917 4846 5930 4860
rect 5998 4856 6151 4860
rect 5880 4844 5902 4846
rect 5980 4844 6172 4856
rect 6251 4844 6264 4874
rect 6279 4860 6309 4874
rect 6346 4844 6365 4874
rect 6380 4844 6386 4874
rect 6395 4844 6408 4874
rect 6423 4860 6453 4874
rect 6496 4860 6539 4874
rect 6546 4860 6766 4874
rect 6773 4860 6803 4874
rect 6463 4846 6478 4858
rect 6497 4846 6510 4860
rect 6578 4856 6731 4860
rect 6460 4844 6482 4846
rect 6560 4844 6752 4856
rect 6831 4844 6844 4874
rect 6859 4860 6889 4874
rect 6926 4844 6945 4874
rect 6960 4844 6966 4874
rect 6975 4844 6988 4874
rect 7003 4860 7033 4874
rect 7076 4860 7119 4874
rect 7126 4860 7346 4874
rect 7353 4860 7383 4874
rect 7043 4846 7058 4858
rect 7077 4846 7090 4860
rect 7158 4856 7311 4860
rect 7040 4844 7062 4846
rect 7140 4844 7332 4856
rect 7411 4844 7424 4874
rect 7439 4860 7469 4874
rect 7506 4844 7525 4874
rect 7540 4844 7546 4874
rect 7555 4844 7568 4874
rect 7583 4856 7613 4874
rect 7656 4860 7670 4874
rect 7706 4860 7926 4874
rect 7657 4858 7670 4860
rect 7623 4846 7638 4858
rect 7620 4844 7642 4846
rect 7647 4844 7677 4858
rect 7738 4856 7891 4860
rect 7720 4844 7912 4856
rect 7955 4844 7985 4858
rect 7991 4844 8004 4874
rect 8019 4856 8049 4874
rect 8092 4844 8105 4874
rect 8135 4844 8148 4874
rect 8163 4856 8193 4874
rect 8236 4860 8250 4874
rect 8286 4860 8506 4874
rect 8237 4858 8250 4860
rect 8203 4846 8218 4858
rect 8200 4844 8222 4846
rect 8227 4844 8257 4858
rect 8318 4856 8471 4860
rect 8300 4844 8492 4856
rect 8535 4844 8565 4858
rect 8571 4844 8584 4874
rect 8599 4856 8629 4874
rect 8672 4844 8685 4874
rect 8715 4844 8728 4874
rect 8743 4856 8773 4874
rect 8816 4860 8830 4874
rect 8866 4860 9086 4874
rect 8817 4858 8830 4860
rect 8783 4846 8798 4858
rect 8780 4844 8802 4846
rect 8807 4844 8837 4858
rect 8898 4856 9051 4860
rect 8880 4844 9072 4856
rect 9115 4844 9145 4858
rect 9151 4844 9164 4874
rect 9179 4856 9209 4874
rect 9252 4844 9265 4874
rect 0 4830 9265 4844
rect 15 4760 28 4830
rect 80 4826 102 4830
rect 73 4804 102 4818
rect 155 4804 171 4818
rect 209 4814 215 4816
rect 222 4814 330 4830
rect 337 4814 343 4816
rect 351 4814 366 4830
rect 432 4824 451 4827
rect 73 4802 171 4804
rect 198 4802 366 4814
rect 381 4804 397 4818
rect 432 4805 454 4824
rect 464 4818 480 4819
rect 463 4816 480 4818
rect 464 4811 480 4816
rect 454 4804 460 4805
rect 463 4804 492 4811
rect 381 4803 492 4804
rect 381 4802 498 4803
rect 57 4794 108 4802
rect 155 4794 189 4802
rect 57 4782 82 4794
rect 89 4782 108 4794
rect 162 4792 189 4794
rect 198 4792 419 4802
rect 454 4799 460 4802
rect 162 4788 419 4792
rect 57 4774 108 4782
rect 155 4774 419 4788
rect 463 4794 498 4802
rect 9 4726 28 4760
rect 73 4766 102 4774
rect 73 4760 90 4766
rect 73 4758 107 4760
rect 155 4758 171 4774
rect 172 4764 380 4774
rect 381 4764 397 4774
rect 445 4770 460 4785
rect 463 4782 464 4794
rect 471 4782 498 4794
rect 463 4774 498 4782
rect 463 4773 492 4774
rect 183 4760 397 4764
rect 198 4758 397 4760
rect 432 4760 445 4770
rect 463 4760 480 4773
rect 432 4758 480 4760
rect 74 4754 107 4758
rect 70 4752 107 4754
rect 70 4751 137 4752
rect 70 4746 101 4751
rect 107 4746 137 4751
rect 70 4742 137 4746
rect 43 4739 137 4742
rect 43 4732 92 4739
rect 43 4726 73 4732
rect 92 4727 97 4732
rect 9 4710 89 4726
rect 101 4718 137 4739
rect 198 4734 387 4758
rect 432 4757 479 4758
rect 445 4752 479 4757
rect 213 4731 387 4734
rect 206 4728 387 4731
rect 415 4751 479 4752
rect 9 4708 28 4710
rect 43 4708 77 4710
rect 9 4692 89 4708
rect 9 4686 28 4692
rect -1 4670 28 4686
rect 43 4676 73 4692
rect 101 4670 107 4718
rect 110 4712 129 4718
rect 144 4712 174 4720
rect 110 4704 174 4712
rect 110 4688 190 4704
rect 206 4697 268 4728
rect 284 4697 346 4728
rect 415 4726 464 4751
rect 479 4726 509 4742
rect 378 4712 408 4720
rect 415 4718 525 4726
rect 378 4704 423 4712
rect 110 4686 129 4688
rect 144 4686 190 4688
rect 110 4670 190 4686
rect 217 4684 252 4697
rect 293 4694 330 4697
rect 293 4692 335 4694
rect 222 4681 252 4684
rect 231 4677 238 4681
rect 238 4676 239 4677
rect 197 4670 207 4676
rect -7 4662 34 4670
rect -7 4636 8 4662
rect 15 4636 34 4662
rect 98 4658 129 4670
rect 144 4658 247 4670
rect 259 4660 285 4686
rect 300 4681 330 4692
rect 362 4688 424 4704
rect 362 4686 408 4688
rect 362 4670 424 4686
rect 436 4670 442 4718
rect 445 4710 525 4718
rect 445 4708 464 4710
rect 479 4708 513 4710
rect 445 4692 525 4708
rect 445 4670 464 4692
rect 479 4676 509 4692
rect 537 4686 543 4760
rect 546 4686 565 4830
rect 580 4686 586 4830
rect 595 4760 608 4830
rect 660 4826 682 4830
rect 653 4804 682 4818
rect 735 4804 751 4818
rect 789 4814 795 4816
rect 802 4814 910 4830
rect 917 4814 923 4816
rect 931 4814 946 4830
rect 1012 4824 1031 4827
rect 653 4802 751 4804
rect 778 4802 946 4814
rect 961 4804 977 4818
rect 1012 4805 1034 4824
rect 1044 4818 1060 4819
rect 1043 4816 1060 4818
rect 1044 4811 1060 4816
rect 1034 4804 1040 4805
rect 1043 4804 1072 4811
rect 961 4803 1072 4804
rect 961 4802 1078 4803
rect 637 4794 688 4802
rect 735 4794 769 4802
rect 637 4782 662 4794
rect 669 4782 688 4794
rect 742 4792 769 4794
rect 778 4792 999 4802
rect 1034 4799 1040 4802
rect 742 4788 999 4792
rect 637 4774 688 4782
rect 735 4774 999 4788
rect 1043 4794 1078 4802
rect 589 4726 608 4760
rect 653 4766 682 4774
rect 653 4760 670 4766
rect 653 4758 687 4760
rect 735 4758 751 4774
rect 752 4764 960 4774
rect 961 4764 977 4774
rect 1025 4770 1040 4785
rect 1043 4782 1044 4794
rect 1051 4782 1078 4794
rect 1043 4774 1078 4782
rect 1043 4773 1072 4774
rect 763 4760 977 4764
rect 778 4758 977 4760
rect 1012 4760 1025 4770
rect 1043 4760 1060 4773
rect 1012 4758 1060 4760
rect 654 4754 687 4758
rect 650 4752 687 4754
rect 650 4751 717 4752
rect 650 4746 681 4751
rect 687 4746 717 4751
rect 650 4742 717 4746
rect 623 4739 717 4742
rect 623 4732 672 4739
rect 623 4726 653 4732
rect 672 4727 677 4732
rect 589 4710 669 4726
rect 681 4718 717 4739
rect 778 4734 967 4758
rect 1012 4757 1059 4758
rect 1025 4752 1059 4757
rect 793 4731 967 4734
rect 786 4728 967 4731
rect 995 4751 1059 4752
rect 589 4708 608 4710
rect 623 4708 657 4710
rect 589 4692 669 4708
rect 589 4686 608 4692
rect 305 4660 408 4670
rect 259 4658 408 4660
rect 429 4658 464 4670
rect 98 4656 260 4658
rect 110 4636 129 4656
rect 144 4654 174 4656
rect -7 4628 34 4636
rect 116 4632 129 4636
rect 181 4640 260 4656
rect 292 4656 464 4658
rect 292 4640 371 4656
rect 378 4654 408 4656
rect -1 4618 28 4628
rect 43 4618 73 4632
rect 116 4618 159 4632
rect 181 4628 371 4640
rect 436 4636 442 4656
rect 166 4618 196 4628
rect 197 4618 355 4628
rect 359 4618 389 4628
rect 393 4618 423 4632
rect 451 4618 464 4656
rect 536 4670 565 4686
rect 579 4670 608 4686
rect 623 4676 653 4692
rect 681 4670 687 4718
rect 690 4712 709 4718
rect 724 4712 754 4720
rect 690 4704 754 4712
rect 690 4688 770 4704
rect 786 4697 848 4728
rect 864 4697 926 4728
rect 995 4726 1044 4751
rect 1059 4726 1089 4742
rect 958 4712 988 4720
rect 995 4718 1105 4726
rect 958 4704 1003 4712
rect 690 4686 709 4688
rect 724 4686 770 4688
rect 690 4670 770 4686
rect 797 4684 832 4697
rect 873 4694 910 4697
rect 873 4692 915 4694
rect 802 4681 832 4684
rect 811 4677 818 4681
rect 818 4676 819 4677
rect 777 4670 787 4676
rect 536 4662 571 4670
rect 536 4636 537 4662
rect 544 4636 571 4662
rect 479 4618 509 4632
rect 536 4628 571 4636
rect 573 4662 614 4670
rect 573 4636 588 4662
rect 595 4636 614 4662
rect 678 4658 709 4670
rect 724 4658 827 4670
rect 839 4660 865 4686
rect 880 4681 910 4692
rect 942 4688 1004 4704
rect 942 4686 988 4688
rect 942 4670 1004 4686
rect 1016 4670 1022 4718
rect 1025 4710 1105 4718
rect 1025 4708 1044 4710
rect 1059 4708 1093 4710
rect 1025 4692 1105 4708
rect 1025 4670 1044 4692
rect 1059 4676 1089 4692
rect 1117 4686 1123 4760
rect 1126 4686 1145 4830
rect 1160 4686 1166 4830
rect 1175 4760 1188 4830
rect 1240 4826 1262 4830
rect 1233 4804 1262 4818
rect 1315 4804 1331 4818
rect 1369 4814 1375 4816
rect 1382 4814 1490 4830
rect 1497 4814 1503 4816
rect 1511 4814 1526 4830
rect 1592 4824 1611 4827
rect 1233 4802 1331 4804
rect 1358 4802 1526 4814
rect 1541 4804 1557 4818
rect 1592 4805 1614 4824
rect 1624 4818 1640 4819
rect 1623 4816 1640 4818
rect 1624 4811 1640 4816
rect 1614 4804 1620 4805
rect 1623 4804 1652 4811
rect 1541 4803 1652 4804
rect 1541 4802 1658 4803
rect 1217 4794 1268 4802
rect 1315 4794 1349 4802
rect 1217 4782 1242 4794
rect 1249 4782 1268 4794
rect 1322 4792 1349 4794
rect 1358 4792 1579 4802
rect 1614 4799 1620 4802
rect 1322 4788 1579 4792
rect 1217 4774 1268 4782
rect 1315 4774 1579 4788
rect 1623 4794 1658 4802
rect 1169 4726 1188 4760
rect 1233 4766 1262 4774
rect 1233 4760 1250 4766
rect 1233 4758 1267 4760
rect 1315 4758 1331 4774
rect 1332 4764 1540 4774
rect 1541 4764 1557 4774
rect 1605 4770 1620 4785
rect 1623 4782 1624 4794
rect 1631 4782 1658 4794
rect 1623 4774 1658 4782
rect 1623 4773 1652 4774
rect 1343 4760 1557 4764
rect 1358 4758 1557 4760
rect 1592 4760 1605 4770
rect 1623 4760 1640 4773
rect 1592 4758 1640 4760
rect 1234 4754 1267 4758
rect 1230 4752 1267 4754
rect 1230 4751 1297 4752
rect 1230 4746 1261 4751
rect 1267 4746 1297 4751
rect 1230 4742 1297 4746
rect 1203 4739 1297 4742
rect 1203 4732 1252 4739
rect 1203 4726 1233 4732
rect 1252 4727 1257 4732
rect 1169 4710 1249 4726
rect 1261 4718 1297 4739
rect 1358 4734 1547 4758
rect 1592 4757 1639 4758
rect 1605 4752 1639 4757
rect 1373 4731 1547 4734
rect 1366 4728 1547 4731
rect 1575 4751 1639 4752
rect 1169 4708 1188 4710
rect 1203 4708 1237 4710
rect 1169 4692 1249 4708
rect 1169 4686 1188 4692
rect 885 4660 988 4670
rect 839 4658 988 4660
rect 1009 4658 1044 4670
rect 678 4656 840 4658
rect 690 4636 709 4656
rect 724 4654 754 4656
rect 573 4628 614 4636
rect 696 4632 709 4636
rect 761 4640 840 4656
rect 872 4656 1044 4658
rect 872 4640 951 4656
rect 958 4654 988 4656
rect 536 4618 565 4628
rect 579 4618 608 4628
rect 623 4618 653 4632
rect 696 4618 739 4632
rect 761 4628 951 4640
rect 1016 4636 1022 4656
rect 746 4618 776 4628
rect 777 4618 935 4628
rect 939 4618 969 4628
rect 973 4618 1003 4632
rect 1031 4618 1044 4656
rect 1116 4670 1145 4686
rect 1159 4670 1188 4686
rect 1203 4676 1233 4692
rect 1261 4670 1267 4718
rect 1270 4712 1289 4718
rect 1304 4712 1334 4720
rect 1270 4704 1334 4712
rect 1270 4688 1350 4704
rect 1366 4697 1428 4728
rect 1444 4697 1506 4728
rect 1575 4726 1624 4751
rect 1639 4726 1669 4742
rect 1538 4712 1568 4720
rect 1575 4718 1685 4726
rect 1538 4704 1583 4712
rect 1270 4686 1289 4688
rect 1304 4686 1350 4688
rect 1270 4670 1350 4686
rect 1377 4684 1412 4697
rect 1453 4694 1490 4697
rect 1453 4692 1495 4694
rect 1382 4681 1412 4684
rect 1391 4677 1398 4681
rect 1398 4676 1399 4677
rect 1357 4670 1367 4676
rect 1116 4662 1151 4670
rect 1116 4636 1117 4662
rect 1124 4636 1151 4662
rect 1059 4618 1089 4632
rect 1116 4628 1151 4636
rect 1153 4662 1194 4670
rect 1153 4636 1168 4662
rect 1175 4636 1194 4662
rect 1258 4658 1289 4670
rect 1304 4658 1407 4670
rect 1419 4660 1445 4686
rect 1460 4681 1490 4692
rect 1522 4688 1584 4704
rect 1522 4686 1568 4688
rect 1522 4670 1584 4686
rect 1596 4670 1602 4718
rect 1605 4710 1685 4718
rect 1605 4708 1624 4710
rect 1639 4708 1673 4710
rect 1605 4692 1685 4708
rect 1605 4670 1624 4692
rect 1639 4676 1669 4692
rect 1697 4686 1703 4760
rect 1706 4686 1725 4830
rect 1740 4686 1746 4830
rect 1755 4760 1768 4830
rect 1820 4826 1842 4830
rect 1813 4804 1842 4818
rect 1895 4804 1911 4818
rect 1949 4814 1955 4816
rect 1962 4814 2070 4830
rect 2077 4814 2083 4816
rect 2091 4814 2106 4830
rect 2172 4824 2191 4827
rect 1813 4802 1911 4804
rect 1938 4802 2106 4814
rect 2121 4804 2137 4818
rect 2172 4805 2194 4824
rect 2204 4818 2220 4819
rect 2203 4816 2220 4818
rect 2204 4811 2220 4816
rect 2194 4804 2200 4805
rect 2203 4804 2232 4811
rect 2121 4803 2232 4804
rect 2121 4802 2238 4803
rect 1797 4794 1848 4802
rect 1895 4794 1929 4802
rect 1797 4782 1822 4794
rect 1829 4782 1848 4794
rect 1902 4792 1929 4794
rect 1938 4792 2159 4802
rect 2194 4799 2200 4802
rect 1902 4788 2159 4792
rect 1797 4774 1848 4782
rect 1895 4774 2159 4788
rect 2203 4794 2238 4802
rect 1749 4726 1768 4760
rect 1813 4766 1842 4774
rect 1813 4760 1830 4766
rect 1813 4758 1847 4760
rect 1895 4758 1911 4774
rect 1912 4764 2120 4774
rect 2121 4764 2137 4774
rect 2185 4770 2200 4785
rect 2203 4782 2204 4794
rect 2211 4782 2238 4794
rect 2203 4774 2238 4782
rect 2203 4773 2232 4774
rect 1923 4760 2137 4764
rect 1938 4758 2137 4760
rect 2172 4760 2185 4770
rect 2203 4760 2220 4773
rect 2172 4758 2220 4760
rect 1814 4754 1847 4758
rect 1810 4752 1847 4754
rect 1810 4751 1877 4752
rect 1810 4746 1841 4751
rect 1847 4746 1877 4751
rect 1810 4742 1877 4746
rect 1783 4739 1877 4742
rect 1783 4732 1832 4739
rect 1783 4726 1813 4732
rect 1832 4727 1837 4732
rect 1749 4710 1829 4726
rect 1841 4718 1877 4739
rect 1938 4734 2127 4758
rect 2172 4757 2219 4758
rect 2185 4752 2219 4757
rect 1953 4731 2127 4734
rect 1946 4728 2127 4731
rect 2155 4751 2219 4752
rect 1749 4708 1768 4710
rect 1783 4708 1817 4710
rect 1749 4692 1829 4708
rect 1749 4686 1768 4692
rect 1465 4660 1568 4670
rect 1419 4658 1568 4660
rect 1589 4658 1624 4670
rect 1258 4656 1420 4658
rect 1270 4636 1289 4656
rect 1304 4654 1334 4656
rect 1153 4628 1194 4636
rect 1276 4632 1289 4636
rect 1341 4640 1420 4656
rect 1452 4656 1624 4658
rect 1452 4640 1531 4656
rect 1538 4654 1568 4656
rect 1116 4618 1145 4628
rect 1159 4618 1188 4628
rect 1203 4618 1233 4632
rect 1276 4618 1319 4632
rect 1341 4628 1531 4640
rect 1596 4636 1602 4656
rect 1326 4618 1356 4628
rect 1357 4618 1515 4628
rect 1519 4618 1549 4628
rect 1553 4618 1583 4632
rect 1611 4618 1624 4656
rect 1696 4670 1725 4686
rect 1739 4670 1768 4686
rect 1783 4676 1813 4692
rect 1841 4670 1847 4718
rect 1850 4712 1869 4718
rect 1884 4712 1914 4720
rect 1850 4704 1914 4712
rect 1850 4688 1930 4704
rect 1946 4697 2008 4728
rect 2024 4697 2086 4728
rect 2155 4726 2204 4751
rect 2219 4726 2249 4742
rect 2118 4712 2148 4720
rect 2155 4718 2265 4726
rect 2118 4704 2163 4712
rect 1850 4686 1869 4688
rect 1884 4686 1930 4688
rect 1850 4670 1930 4686
rect 1957 4684 1992 4697
rect 2033 4694 2070 4697
rect 2033 4692 2075 4694
rect 1962 4681 1992 4684
rect 1971 4677 1978 4681
rect 1978 4676 1979 4677
rect 1937 4670 1947 4676
rect 1696 4662 1731 4670
rect 1696 4636 1697 4662
rect 1704 4636 1731 4662
rect 1639 4618 1669 4632
rect 1696 4628 1731 4636
rect 1733 4662 1774 4670
rect 1733 4636 1748 4662
rect 1755 4636 1774 4662
rect 1838 4658 1869 4670
rect 1884 4658 1987 4670
rect 1999 4660 2025 4686
rect 2040 4681 2070 4692
rect 2102 4688 2164 4704
rect 2102 4686 2148 4688
rect 2102 4670 2164 4686
rect 2176 4670 2182 4718
rect 2185 4710 2265 4718
rect 2185 4708 2204 4710
rect 2219 4708 2253 4710
rect 2185 4692 2265 4708
rect 2185 4670 2204 4692
rect 2219 4676 2249 4692
rect 2277 4686 2283 4760
rect 2286 4686 2305 4830
rect 2320 4686 2326 4830
rect 2335 4760 2348 4830
rect 2400 4826 2422 4830
rect 2393 4804 2422 4818
rect 2475 4804 2491 4818
rect 2529 4814 2535 4816
rect 2542 4814 2650 4830
rect 2657 4814 2663 4816
rect 2671 4814 2686 4830
rect 2752 4824 2771 4827
rect 2393 4802 2491 4804
rect 2518 4802 2686 4814
rect 2701 4804 2717 4818
rect 2752 4805 2774 4824
rect 2784 4818 2800 4819
rect 2783 4816 2800 4818
rect 2784 4811 2800 4816
rect 2774 4804 2780 4805
rect 2783 4804 2812 4811
rect 2701 4803 2812 4804
rect 2701 4802 2818 4803
rect 2377 4794 2428 4802
rect 2475 4794 2509 4802
rect 2377 4782 2402 4794
rect 2409 4782 2428 4794
rect 2482 4792 2509 4794
rect 2518 4792 2739 4802
rect 2774 4799 2780 4802
rect 2482 4788 2739 4792
rect 2377 4774 2428 4782
rect 2475 4774 2739 4788
rect 2783 4794 2818 4802
rect 2329 4726 2348 4760
rect 2393 4766 2422 4774
rect 2393 4760 2410 4766
rect 2393 4758 2427 4760
rect 2475 4758 2491 4774
rect 2492 4764 2700 4774
rect 2701 4764 2717 4774
rect 2765 4770 2780 4785
rect 2783 4782 2784 4794
rect 2791 4782 2818 4794
rect 2783 4774 2818 4782
rect 2783 4773 2812 4774
rect 2503 4760 2717 4764
rect 2518 4758 2717 4760
rect 2752 4760 2765 4770
rect 2783 4760 2800 4773
rect 2752 4758 2800 4760
rect 2394 4754 2427 4758
rect 2390 4752 2427 4754
rect 2390 4751 2457 4752
rect 2390 4746 2421 4751
rect 2427 4746 2457 4751
rect 2390 4742 2457 4746
rect 2363 4739 2457 4742
rect 2363 4732 2412 4739
rect 2363 4726 2393 4732
rect 2412 4727 2417 4732
rect 2329 4710 2409 4726
rect 2421 4718 2457 4739
rect 2518 4734 2707 4758
rect 2752 4757 2799 4758
rect 2765 4752 2799 4757
rect 2533 4731 2707 4734
rect 2526 4728 2707 4731
rect 2735 4751 2799 4752
rect 2329 4708 2348 4710
rect 2363 4708 2397 4710
rect 2329 4692 2409 4708
rect 2329 4686 2348 4692
rect 2045 4660 2148 4670
rect 1999 4658 2148 4660
rect 2169 4658 2204 4670
rect 1838 4656 2000 4658
rect 1850 4636 1869 4656
rect 1884 4654 1914 4656
rect 1733 4628 1774 4636
rect 1856 4632 1869 4636
rect 1921 4640 2000 4656
rect 2032 4656 2204 4658
rect 2032 4640 2111 4656
rect 2118 4654 2148 4656
rect 1696 4618 1725 4628
rect 1739 4618 1768 4628
rect 1783 4618 1813 4632
rect 1856 4618 1899 4632
rect 1921 4628 2111 4640
rect 2176 4636 2182 4656
rect 1906 4618 1936 4628
rect 1937 4618 2095 4628
rect 2099 4618 2129 4628
rect 2133 4618 2163 4632
rect 2191 4618 2204 4656
rect 2276 4670 2305 4686
rect 2319 4670 2348 4686
rect 2363 4676 2393 4692
rect 2421 4670 2427 4718
rect 2430 4712 2449 4718
rect 2464 4712 2494 4720
rect 2430 4704 2494 4712
rect 2430 4688 2510 4704
rect 2526 4697 2588 4728
rect 2604 4697 2666 4728
rect 2735 4726 2784 4751
rect 2799 4726 2829 4742
rect 2698 4712 2728 4720
rect 2735 4718 2845 4726
rect 2698 4704 2743 4712
rect 2430 4686 2449 4688
rect 2464 4686 2510 4688
rect 2430 4670 2510 4686
rect 2537 4684 2572 4697
rect 2613 4694 2650 4697
rect 2613 4692 2655 4694
rect 2542 4681 2572 4684
rect 2551 4677 2558 4681
rect 2558 4676 2559 4677
rect 2517 4670 2527 4676
rect 2276 4662 2311 4670
rect 2276 4636 2277 4662
rect 2284 4636 2311 4662
rect 2219 4618 2249 4632
rect 2276 4628 2311 4636
rect 2313 4662 2354 4670
rect 2313 4636 2328 4662
rect 2335 4636 2354 4662
rect 2418 4658 2449 4670
rect 2464 4658 2567 4670
rect 2579 4660 2605 4686
rect 2620 4681 2650 4692
rect 2682 4688 2744 4704
rect 2682 4686 2728 4688
rect 2682 4670 2744 4686
rect 2756 4670 2762 4718
rect 2765 4710 2845 4718
rect 2765 4708 2784 4710
rect 2799 4708 2833 4710
rect 2765 4692 2845 4708
rect 2765 4670 2784 4692
rect 2799 4676 2829 4692
rect 2857 4686 2863 4760
rect 2866 4686 2885 4830
rect 2900 4686 2906 4830
rect 2915 4760 2928 4830
rect 2980 4826 3002 4830
rect 2973 4804 3002 4818
rect 3055 4804 3071 4818
rect 3109 4814 3115 4816
rect 3122 4814 3230 4830
rect 3237 4814 3243 4816
rect 3251 4814 3266 4830
rect 3332 4824 3351 4827
rect 2973 4802 3071 4804
rect 3098 4802 3266 4814
rect 3281 4804 3297 4818
rect 3332 4805 3354 4824
rect 3364 4818 3380 4819
rect 3363 4816 3380 4818
rect 3364 4811 3380 4816
rect 3354 4804 3360 4805
rect 3363 4804 3392 4811
rect 3281 4803 3392 4804
rect 3281 4802 3398 4803
rect 2957 4794 3008 4802
rect 3055 4794 3089 4802
rect 2957 4782 2982 4794
rect 2989 4782 3008 4794
rect 3062 4792 3089 4794
rect 3098 4792 3319 4802
rect 3354 4799 3360 4802
rect 3062 4788 3319 4792
rect 2957 4774 3008 4782
rect 3055 4774 3319 4788
rect 3363 4794 3398 4802
rect 2909 4726 2928 4760
rect 2973 4766 3002 4774
rect 2973 4760 2990 4766
rect 2973 4758 3007 4760
rect 3055 4758 3071 4774
rect 3072 4764 3280 4774
rect 3281 4764 3297 4774
rect 3345 4770 3360 4785
rect 3363 4782 3364 4794
rect 3371 4782 3398 4794
rect 3363 4774 3398 4782
rect 3363 4773 3392 4774
rect 3083 4760 3297 4764
rect 3098 4758 3297 4760
rect 3332 4760 3345 4770
rect 3363 4760 3380 4773
rect 3332 4758 3380 4760
rect 2974 4754 3007 4758
rect 2970 4752 3007 4754
rect 2970 4751 3037 4752
rect 2970 4746 3001 4751
rect 3007 4746 3037 4751
rect 2970 4742 3037 4746
rect 2943 4739 3037 4742
rect 2943 4732 2992 4739
rect 2943 4726 2973 4732
rect 2992 4727 2997 4732
rect 2909 4710 2989 4726
rect 3001 4718 3037 4739
rect 3098 4734 3287 4758
rect 3332 4757 3379 4758
rect 3345 4752 3379 4757
rect 3113 4731 3287 4734
rect 3106 4728 3287 4731
rect 3315 4751 3379 4752
rect 2909 4708 2928 4710
rect 2943 4708 2977 4710
rect 2909 4692 2989 4708
rect 2909 4686 2928 4692
rect 2625 4660 2728 4670
rect 2579 4658 2728 4660
rect 2749 4658 2784 4670
rect 2418 4656 2580 4658
rect 2430 4636 2449 4656
rect 2464 4654 2494 4656
rect 2313 4628 2354 4636
rect 2436 4632 2449 4636
rect 2501 4640 2580 4656
rect 2612 4656 2784 4658
rect 2612 4640 2691 4656
rect 2698 4654 2728 4656
rect 2276 4618 2305 4628
rect 2319 4618 2348 4628
rect 2363 4618 2393 4632
rect 2436 4618 2479 4632
rect 2501 4628 2691 4640
rect 2756 4636 2762 4656
rect 2486 4618 2516 4628
rect 2517 4618 2675 4628
rect 2679 4618 2709 4628
rect 2713 4618 2743 4632
rect 2771 4618 2784 4656
rect 2856 4670 2885 4686
rect 2899 4670 2928 4686
rect 2943 4676 2973 4692
rect 3001 4670 3007 4718
rect 3010 4712 3029 4718
rect 3044 4712 3074 4720
rect 3010 4704 3074 4712
rect 3010 4688 3090 4704
rect 3106 4697 3168 4728
rect 3184 4697 3246 4728
rect 3315 4726 3364 4751
rect 3379 4726 3409 4742
rect 3278 4712 3308 4720
rect 3315 4718 3425 4726
rect 3278 4704 3323 4712
rect 3010 4686 3029 4688
rect 3044 4686 3090 4688
rect 3010 4670 3090 4686
rect 3117 4684 3152 4697
rect 3193 4694 3230 4697
rect 3193 4692 3235 4694
rect 3122 4681 3152 4684
rect 3131 4677 3138 4681
rect 3138 4676 3139 4677
rect 3097 4670 3107 4676
rect 2856 4662 2891 4670
rect 2856 4636 2857 4662
rect 2864 4636 2891 4662
rect 2799 4618 2829 4632
rect 2856 4628 2891 4636
rect 2893 4662 2934 4670
rect 2893 4636 2908 4662
rect 2915 4636 2934 4662
rect 2998 4658 3029 4670
rect 3044 4658 3147 4670
rect 3159 4660 3185 4686
rect 3200 4681 3230 4692
rect 3262 4688 3324 4704
rect 3262 4686 3308 4688
rect 3262 4670 3324 4686
rect 3336 4670 3342 4718
rect 3345 4710 3425 4718
rect 3345 4708 3364 4710
rect 3379 4708 3413 4710
rect 3345 4692 3425 4708
rect 3345 4670 3364 4692
rect 3379 4676 3409 4692
rect 3437 4686 3443 4760
rect 3446 4686 3465 4830
rect 3480 4686 3486 4830
rect 3495 4760 3508 4830
rect 3560 4826 3582 4830
rect 3553 4804 3582 4818
rect 3635 4804 3651 4818
rect 3689 4814 3695 4816
rect 3702 4814 3810 4830
rect 3817 4814 3823 4816
rect 3831 4814 3846 4830
rect 3912 4824 3931 4827
rect 3553 4802 3651 4804
rect 3678 4802 3846 4814
rect 3861 4804 3877 4818
rect 3912 4805 3934 4824
rect 3944 4818 3960 4819
rect 3943 4816 3960 4818
rect 3944 4811 3960 4816
rect 3934 4804 3940 4805
rect 3943 4804 3972 4811
rect 3861 4803 3972 4804
rect 3861 4802 3978 4803
rect 3537 4794 3588 4802
rect 3635 4794 3669 4802
rect 3537 4782 3562 4794
rect 3569 4782 3588 4794
rect 3642 4792 3669 4794
rect 3678 4792 3899 4802
rect 3934 4799 3940 4802
rect 3642 4788 3899 4792
rect 3537 4774 3588 4782
rect 3635 4774 3899 4788
rect 3943 4794 3978 4802
rect 3489 4726 3508 4760
rect 3553 4766 3582 4774
rect 3553 4760 3570 4766
rect 3553 4758 3587 4760
rect 3635 4758 3651 4774
rect 3652 4764 3860 4774
rect 3861 4764 3877 4774
rect 3925 4770 3940 4785
rect 3943 4782 3944 4794
rect 3951 4782 3978 4794
rect 3943 4774 3978 4782
rect 3943 4773 3972 4774
rect 3663 4760 3877 4764
rect 3678 4758 3877 4760
rect 3912 4760 3925 4770
rect 3943 4760 3960 4773
rect 3912 4758 3960 4760
rect 3554 4754 3587 4758
rect 3550 4752 3587 4754
rect 3550 4751 3617 4752
rect 3550 4746 3581 4751
rect 3587 4746 3617 4751
rect 3550 4742 3617 4746
rect 3523 4739 3617 4742
rect 3523 4732 3572 4739
rect 3523 4726 3553 4732
rect 3572 4727 3577 4732
rect 3489 4710 3569 4726
rect 3581 4718 3617 4739
rect 3678 4734 3867 4758
rect 3912 4757 3959 4758
rect 3925 4752 3959 4757
rect 3693 4731 3867 4734
rect 3686 4728 3867 4731
rect 3895 4751 3959 4752
rect 3489 4708 3508 4710
rect 3523 4708 3557 4710
rect 3489 4692 3569 4708
rect 3489 4686 3508 4692
rect 3205 4660 3308 4670
rect 3159 4658 3308 4660
rect 3329 4658 3364 4670
rect 2998 4656 3160 4658
rect 3010 4636 3029 4656
rect 3044 4654 3074 4656
rect 2893 4628 2934 4636
rect 3016 4632 3029 4636
rect 3081 4640 3160 4656
rect 3192 4656 3364 4658
rect 3192 4640 3271 4656
rect 3278 4654 3308 4656
rect 2856 4618 2885 4628
rect 2899 4618 2928 4628
rect 2943 4618 2973 4632
rect 3016 4618 3059 4632
rect 3081 4628 3271 4640
rect 3336 4636 3342 4656
rect 3066 4618 3096 4628
rect 3097 4618 3255 4628
rect 3259 4618 3289 4628
rect 3293 4618 3323 4632
rect 3351 4618 3364 4656
rect 3436 4670 3465 4686
rect 3479 4670 3508 4686
rect 3523 4676 3553 4692
rect 3581 4670 3587 4718
rect 3590 4712 3609 4718
rect 3624 4712 3654 4720
rect 3590 4704 3654 4712
rect 3590 4688 3670 4704
rect 3686 4697 3748 4728
rect 3764 4697 3826 4728
rect 3895 4726 3944 4751
rect 3959 4726 3989 4742
rect 3858 4712 3888 4720
rect 3895 4718 4005 4726
rect 3858 4704 3903 4712
rect 3590 4686 3609 4688
rect 3624 4686 3670 4688
rect 3590 4670 3670 4686
rect 3697 4684 3732 4697
rect 3773 4694 3810 4697
rect 3773 4692 3815 4694
rect 3702 4681 3732 4684
rect 3711 4677 3718 4681
rect 3718 4676 3719 4677
rect 3677 4670 3687 4676
rect 3436 4662 3471 4670
rect 3436 4636 3437 4662
rect 3444 4636 3471 4662
rect 3379 4618 3409 4632
rect 3436 4628 3471 4636
rect 3473 4662 3514 4670
rect 3473 4636 3488 4662
rect 3495 4636 3514 4662
rect 3578 4658 3609 4670
rect 3624 4658 3727 4670
rect 3739 4660 3765 4686
rect 3780 4681 3810 4692
rect 3842 4688 3904 4704
rect 3842 4686 3888 4688
rect 3842 4670 3904 4686
rect 3916 4670 3922 4718
rect 3925 4710 4005 4718
rect 3925 4708 3944 4710
rect 3959 4708 3993 4710
rect 3925 4692 4005 4708
rect 3925 4670 3944 4692
rect 3959 4676 3989 4692
rect 4017 4686 4023 4760
rect 4026 4686 4045 4830
rect 4060 4686 4066 4830
rect 4075 4760 4088 4830
rect 4140 4826 4162 4830
rect 4133 4804 4162 4818
rect 4215 4804 4231 4818
rect 4269 4814 4275 4816
rect 4282 4814 4390 4830
rect 4397 4814 4403 4816
rect 4411 4814 4426 4830
rect 4492 4824 4511 4827
rect 4133 4802 4231 4804
rect 4258 4802 4426 4814
rect 4441 4804 4457 4818
rect 4492 4805 4514 4824
rect 4524 4818 4540 4819
rect 4523 4816 4540 4818
rect 4524 4811 4540 4816
rect 4514 4804 4520 4805
rect 4523 4804 4552 4811
rect 4441 4803 4552 4804
rect 4441 4802 4558 4803
rect 4117 4794 4168 4802
rect 4215 4794 4249 4802
rect 4117 4782 4142 4794
rect 4149 4782 4168 4794
rect 4222 4792 4249 4794
rect 4258 4792 4479 4802
rect 4514 4799 4520 4802
rect 4222 4788 4479 4792
rect 4117 4774 4168 4782
rect 4215 4774 4479 4788
rect 4523 4794 4558 4802
rect 4069 4726 4088 4760
rect 4133 4766 4162 4774
rect 4133 4760 4150 4766
rect 4133 4758 4167 4760
rect 4215 4758 4231 4774
rect 4232 4764 4440 4774
rect 4441 4764 4457 4774
rect 4505 4770 4520 4785
rect 4523 4782 4524 4794
rect 4531 4782 4558 4794
rect 4523 4774 4558 4782
rect 4523 4773 4552 4774
rect 4243 4760 4457 4764
rect 4258 4758 4457 4760
rect 4492 4760 4505 4770
rect 4523 4760 4540 4773
rect 4492 4758 4540 4760
rect 4134 4754 4167 4758
rect 4130 4752 4167 4754
rect 4130 4751 4197 4752
rect 4130 4746 4161 4751
rect 4167 4746 4197 4751
rect 4130 4742 4197 4746
rect 4103 4739 4197 4742
rect 4103 4732 4152 4739
rect 4103 4726 4133 4732
rect 4152 4727 4157 4732
rect 4069 4710 4149 4726
rect 4161 4718 4197 4739
rect 4258 4734 4447 4758
rect 4492 4757 4539 4758
rect 4505 4752 4539 4757
rect 4273 4731 4447 4734
rect 4266 4728 4447 4731
rect 4475 4751 4539 4752
rect 4069 4708 4088 4710
rect 4103 4708 4137 4710
rect 4069 4692 4149 4708
rect 4069 4686 4088 4692
rect 3785 4660 3888 4670
rect 3739 4658 3888 4660
rect 3909 4658 3944 4670
rect 3578 4656 3740 4658
rect 3590 4636 3609 4656
rect 3624 4654 3654 4656
rect 3473 4628 3514 4636
rect 3596 4632 3609 4636
rect 3661 4640 3740 4656
rect 3772 4656 3944 4658
rect 3772 4640 3851 4656
rect 3858 4654 3888 4656
rect 3436 4618 3465 4628
rect 3479 4618 3508 4628
rect 3523 4618 3553 4632
rect 3596 4618 3639 4632
rect 3661 4628 3851 4640
rect 3916 4636 3922 4656
rect 3646 4618 3676 4628
rect 3677 4618 3835 4628
rect 3839 4618 3869 4628
rect 3873 4618 3903 4632
rect 3931 4618 3944 4656
rect 4016 4670 4045 4686
rect 4059 4670 4088 4686
rect 4103 4676 4133 4692
rect 4161 4670 4167 4718
rect 4170 4712 4189 4718
rect 4204 4712 4234 4720
rect 4170 4704 4234 4712
rect 4170 4688 4250 4704
rect 4266 4697 4328 4728
rect 4344 4697 4406 4728
rect 4475 4726 4524 4751
rect 4539 4726 4569 4742
rect 4438 4712 4468 4720
rect 4475 4718 4585 4726
rect 4438 4704 4483 4712
rect 4170 4686 4189 4688
rect 4204 4686 4250 4688
rect 4170 4670 4250 4686
rect 4277 4684 4312 4697
rect 4353 4694 4390 4697
rect 4353 4692 4395 4694
rect 4282 4681 4312 4684
rect 4291 4677 4298 4681
rect 4298 4676 4299 4677
rect 4257 4670 4267 4676
rect 4016 4662 4051 4670
rect 4016 4636 4017 4662
rect 4024 4636 4051 4662
rect 3959 4618 3989 4632
rect 4016 4628 4051 4636
rect 4053 4662 4094 4670
rect 4053 4636 4068 4662
rect 4075 4636 4094 4662
rect 4158 4658 4189 4670
rect 4204 4658 4307 4670
rect 4319 4660 4345 4686
rect 4360 4681 4390 4692
rect 4422 4688 4484 4704
rect 4422 4686 4468 4688
rect 4422 4670 4484 4686
rect 4496 4670 4502 4718
rect 4505 4710 4585 4718
rect 4505 4708 4524 4710
rect 4539 4708 4573 4710
rect 4505 4692 4585 4708
rect 4505 4670 4524 4692
rect 4539 4676 4569 4692
rect 4597 4686 4603 4760
rect 4606 4686 4625 4830
rect 4640 4686 4646 4830
rect 4655 4760 4668 4830
rect 4720 4826 4742 4830
rect 4713 4804 4742 4818
rect 4795 4804 4811 4818
rect 4849 4814 4855 4816
rect 4862 4814 4970 4830
rect 4977 4814 4983 4816
rect 4991 4814 5006 4830
rect 5072 4824 5091 4827
rect 4713 4802 4811 4804
rect 4838 4802 5006 4814
rect 5021 4804 5037 4818
rect 5072 4805 5094 4824
rect 5104 4818 5120 4819
rect 5103 4816 5120 4818
rect 5104 4811 5120 4816
rect 5094 4804 5100 4805
rect 5103 4804 5132 4811
rect 5021 4803 5132 4804
rect 5021 4802 5138 4803
rect 4697 4794 4748 4802
rect 4795 4794 4829 4802
rect 4697 4782 4722 4794
rect 4729 4782 4748 4794
rect 4802 4792 4829 4794
rect 4838 4792 5059 4802
rect 5094 4799 5100 4802
rect 4802 4788 5059 4792
rect 4697 4774 4748 4782
rect 4795 4774 5059 4788
rect 5103 4794 5138 4802
rect 4649 4726 4668 4760
rect 4713 4766 4742 4774
rect 4713 4760 4730 4766
rect 4713 4758 4747 4760
rect 4795 4758 4811 4774
rect 4812 4764 5020 4774
rect 5021 4764 5037 4774
rect 5085 4770 5100 4785
rect 5103 4782 5104 4794
rect 5111 4782 5138 4794
rect 5103 4774 5138 4782
rect 5103 4773 5132 4774
rect 4823 4760 5037 4764
rect 4838 4758 5037 4760
rect 5072 4760 5085 4770
rect 5103 4760 5120 4773
rect 5072 4758 5120 4760
rect 4714 4754 4747 4758
rect 4710 4752 4747 4754
rect 4710 4751 4777 4752
rect 4710 4746 4741 4751
rect 4747 4746 4777 4751
rect 4710 4742 4777 4746
rect 4683 4739 4777 4742
rect 4683 4732 4732 4739
rect 4683 4726 4713 4732
rect 4732 4727 4737 4732
rect 4649 4710 4729 4726
rect 4741 4718 4777 4739
rect 4838 4734 5027 4758
rect 5072 4757 5119 4758
rect 5085 4752 5119 4757
rect 4853 4731 5027 4734
rect 4846 4728 5027 4731
rect 5055 4751 5119 4752
rect 4649 4708 4668 4710
rect 4683 4708 4717 4710
rect 4649 4692 4729 4708
rect 4649 4686 4668 4692
rect 4365 4660 4468 4670
rect 4319 4658 4468 4660
rect 4489 4658 4524 4670
rect 4158 4656 4320 4658
rect 4170 4636 4189 4656
rect 4204 4654 4234 4656
rect 4053 4628 4094 4636
rect 4176 4632 4189 4636
rect 4241 4640 4320 4656
rect 4352 4656 4524 4658
rect 4352 4640 4431 4656
rect 4438 4654 4468 4656
rect 4016 4618 4045 4628
rect 4059 4618 4088 4628
rect 4103 4618 4133 4632
rect 4176 4618 4219 4632
rect 4241 4628 4431 4640
rect 4496 4636 4502 4656
rect 4226 4618 4256 4628
rect 4257 4618 4415 4628
rect 4419 4618 4449 4628
rect 4453 4618 4483 4632
rect 4511 4618 4524 4656
rect 4596 4670 4625 4686
rect 4639 4670 4668 4686
rect 4683 4676 4713 4692
rect 4741 4670 4747 4718
rect 4750 4712 4769 4718
rect 4784 4712 4814 4720
rect 4750 4704 4814 4712
rect 4750 4688 4830 4704
rect 4846 4697 4908 4728
rect 4924 4697 4986 4728
rect 5055 4726 5104 4751
rect 5119 4726 5149 4742
rect 5018 4712 5048 4720
rect 5055 4718 5165 4726
rect 5018 4704 5063 4712
rect 4750 4686 4769 4688
rect 4784 4686 4830 4688
rect 4750 4670 4830 4686
rect 4857 4684 4892 4697
rect 4933 4694 4970 4697
rect 4933 4692 4975 4694
rect 4862 4681 4892 4684
rect 4871 4677 4878 4681
rect 4878 4676 4879 4677
rect 4837 4670 4847 4676
rect 4596 4662 4631 4670
rect 4596 4636 4597 4662
rect 4604 4636 4631 4662
rect 4539 4618 4569 4632
rect 4596 4628 4631 4636
rect 4633 4662 4674 4670
rect 4633 4636 4648 4662
rect 4655 4636 4674 4662
rect 4738 4658 4769 4670
rect 4784 4658 4887 4670
rect 4899 4660 4925 4686
rect 4940 4681 4970 4692
rect 5002 4688 5064 4704
rect 5002 4686 5048 4688
rect 5002 4670 5064 4686
rect 5076 4670 5082 4718
rect 5085 4710 5165 4718
rect 5085 4708 5104 4710
rect 5119 4708 5153 4710
rect 5085 4692 5165 4708
rect 5085 4670 5104 4692
rect 5119 4676 5149 4692
rect 5177 4686 5183 4760
rect 5186 4686 5205 4830
rect 5220 4686 5226 4830
rect 5235 4760 5248 4830
rect 5300 4826 5322 4830
rect 5293 4804 5322 4818
rect 5375 4804 5391 4818
rect 5429 4814 5435 4816
rect 5442 4814 5550 4830
rect 5557 4814 5563 4816
rect 5571 4814 5586 4830
rect 5652 4824 5671 4827
rect 5293 4802 5391 4804
rect 5418 4802 5586 4814
rect 5601 4804 5617 4818
rect 5652 4805 5674 4824
rect 5684 4818 5700 4819
rect 5683 4816 5700 4818
rect 5684 4811 5700 4816
rect 5674 4804 5680 4805
rect 5683 4804 5712 4811
rect 5601 4803 5712 4804
rect 5601 4802 5718 4803
rect 5277 4794 5328 4802
rect 5375 4794 5409 4802
rect 5277 4782 5302 4794
rect 5309 4782 5328 4794
rect 5382 4792 5409 4794
rect 5418 4792 5639 4802
rect 5674 4799 5680 4802
rect 5382 4788 5639 4792
rect 5277 4774 5328 4782
rect 5375 4774 5639 4788
rect 5683 4794 5718 4802
rect 5229 4726 5248 4760
rect 5293 4766 5322 4774
rect 5293 4760 5310 4766
rect 5293 4758 5327 4760
rect 5375 4758 5391 4774
rect 5392 4764 5600 4774
rect 5601 4764 5617 4774
rect 5665 4770 5680 4785
rect 5683 4782 5684 4794
rect 5691 4782 5718 4794
rect 5683 4774 5718 4782
rect 5683 4773 5712 4774
rect 5403 4760 5617 4764
rect 5418 4758 5617 4760
rect 5652 4760 5665 4770
rect 5683 4760 5700 4773
rect 5652 4758 5700 4760
rect 5294 4754 5327 4758
rect 5290 4752 5327 4754
rect 5290 4751 5357 4752
rect 5290 4746 5321 4751
rect 5327 4746 5357 4751
rect 5290 4742 5357 4746
rect 5263 4739 5357 4742
rect 5263 4732 5312 4739
rect 5263 4726 5293 4732
rect 5312 4727 5317 4732
rect 5229 4710 5309 4726
rect 5321 4718 5357 4739
rect 5418 4734 5607 4758
rect 5652 4757 5699 4758
rect 5665 4752 5699 4757
rect 5433 4731 5607 4734
rect 5426 4728 5607 4731
rect 5635 4751 5699 4752
rect 5229 4708 5248 4710
rect 5263 4708 5297 4710
rect 5229 4692 5309 4708
rect 5229 4686 5248 4692
rect 4945 4660 5048 4670
rect 4899 4658 5048 4660
rect 5069 4658 5104 4670
rect 4738 4656 4900 4658
rect 4750 4636 4769 4656
rect 4784 4654 4814 4656
rect 4633 4628 4674 4636
rect 4756 4632 4769 4636
rect 4821 4640 4900 4656
rect 4932 4656 5104 4658
rect 4932 4640 5011 4656
rect 5018 4654 5048 4656
rect 4596 4618 4625 4628
rect 4639 4618 4668 4628
rect 4683 4618 4713 4632
rect 4756 4618 4799 4632
rect 4821 4628 5011 4640
rect 5076 4636 5082 4656
rect 4806 4618 4836 4628
rect 4837 4618 4995 4628
rect 4999 4618 5029 4628
rect 5033 4618 5063 4632
rect 5091 4618 5104 4656
rect 5176 4670 5205 4686
rect 5219 4670 5248 4686
rect 5263 4676 5293 4692
rect 5321 4670 5327 4718
rect 5330 4712 5349 4718
rect 5364 4712 5394 4720
rect 5330 4704 5394 4712
rect 5330 4688 5410 4704
rect 5426 4697 5488 4728
rect 5504 4697 5566 4728
rect 5635 4726 5684 4751
rect 5699 4726 5729 4742
rect 5598 4712 5628 4720
rect 5635 4718 5745 4726
rect 5598 4704 5643 4712
rect 5330 4686 5349 4688
rect 5364 4686 5410 4688
rect 5330 4670 5410 4686
rect 5437 4684 5472 4697
rect 5513 4694 5550 4697
rect 5513 4692 5555 4694
rect 5442 4681 5472 4684
rect 5451 4677 5458 4681
rect 5458 4676 5459 4677
rect 5417 4670 5427 4676
rect 5176 4662 5211 4670
rect 5176 4636 5177 4662
rect 5184 4636 5211 4662
rect 5119 4618 5149 4632
rect 5176 4628 5211 4636
rect 5213 4662 5254 4670
rect 5213 4636 5228 4662
rect 5235 4636 5254 4662
rect 5318 4658 5349 4670
rect 5364 4658 5467 4670
rect 5479 4660 5505 4686
rect 5520 4681 5550 4692
rect 5582 4688 5644 4704
rect 5582 4686 5628 4688
rect 5582 4670 5644 4686
rect 5656 4670 5662 4718
rect 5665 4710 5745 4718
rect 5665 4708 5684 4710
rect 5699 4708 5733 4710
rect 5665 4692 5745 4708
rect 5665 4670 5684 4692
rect 5699 4676 5729 4692
rect 5757 4686 5763 4760
rect 5766 4686 5785 4830
rect 5800 4686 5806 4830
rect 5815 4760 5828 4830
rect 5880 4826 5902 4830
rect 5873 4804 5902 4818
rect 5955 4804 5971 4818
rect 6009 4814 6015 4816
rect 6022 4814 6130 4830
rect 6137 4814 6143 4816
rect 6151 4814 6166 4830
rect 6232 4824 6251 4827
rect 5873 4802 5971 4804
rect 5998 4802 6166 4814
rect 6181 4804 6197 4818
rect 6232 4805 6254 4824
rect 6264 4818 6280 4819
rect 6263 4816 6280 4818
rect 6264 4811 6280 4816
rect 6254 4804 6260 4805
rect 6263 4804 6292 4811
rect 6181 4803 6292 4804
rect 6181 4802 6298 4803
rect 5857 4794 5908 4802
rect 5955 4794 5989 4802
rect 5857 4782 5882 4794
rect 5889 4782 5908 4794
rect 5962 4792 5989 4794
rect 5998 4792 6219 4802
rect 6254 4799 6260 4802
rect 5962 4788 6219 4792
rect 5857 4774 5908 4782
rect 5955 4774 6219 4788
rect 6263 4794 6298 4802
rect 5809 4726 5828 4760
rect 5873 4766 5902 4774
rect 5873 4760 5890 4766
rect 5873 4758 5907 4760
rect 5955 4758 5971 4774
rect 5972 4764 6180 4774
rect 6181 4764 6197 4774
rect 6245 4770 6260 4785
rect 6263 4782 6264 4794
rect 6271 4782 6298 4794
rect 6263 4774 6298 4782
rect 6263 4773 6292 4774
rect 5983 4760 6197 4764
rect 5998 4758 6197 4760
rect 6232 4760 6245 4770
rect 6263 4760 6280 4773
rect 6232 4758 6280 4760
rect 5874 4754 5907 4758
rect 5870 4752 5907 4754
rect 5870 4751 5937 4752
rect 5870 4746 5901 4751
rect 5907 4746 5937 4751
rect 5870 4742 5937 4746
rect 5843 4739 5937 4742
rect 5843 4732 5892 4739
rect 5843 4726 5873 4732
rect 5892 4727 5897 4732
rect 5809 4710 5889 4726
rect 5901 4718 5937 4739
rect 5998 4734 6187 4758
rect 6232 4757 6279 4758
rect 6245 4752 6279 4757
rect 6013 4731 6187 4734
rect 6006 4728 6187 4731
rect 6215 4751 6279 4752
rect 5809 4708 5828 4710
rect 5843 4708 5877 4710
rect 5809 4692 5889 4708
rect 5809 4686 5828 4692
rect 5525 4660 5628 4670
rect 5479 4658 5628 4660
rect 5649 4658 5684 4670
rect 5318 4656 5480 4658
rect 5330 4636 5349 4656
rect 5364 4654 5394 4656
rect 5213 4628 5254 4636
rect 5336 4632 5349 4636
rect 5401 4640 5480 4656
rect 5512 4656 5684 4658
rect 5512 4640 5591 4656
rect 5598 4654 5628 4656
rect 5176 4618 5205 4628
rect 5219 4618 5248 4628
rect 5263 4618 5293 4632
rect 5336 4618 5379 4632
rect 5401 4628 5591 4640
rect 5656 4636 5662 4656
rect 5386 4618 5416 4628
rect 5417 4618 5575 4628
rect 5579 4618 5609 4628
rect 5613 4618 5643 4632
rect 5671 4618 5684 4656
rect 5756 4670 5785 4686
rect 5799 4670 5828 4686
rect 5843 4676 5873 4692
rect 5901 4670 5907 4718
rect 5910 4712 5929 4718
rect 5944 4712 5974 4720
rect 5910 4704 5974 4712
rect 5910 4688 5990 4704
rect 6006 4697 6068 4728
rect 6084 4697 6146 4728
rect 6215 4726 6264 4751
rect 6279 4726 6309 4742
rect 6178 4712 6208 4720
rect 6215 4718 6325 4726
rect 6178 4704 6223 4712
rect 5910 4686 5929 4688
rect 5944 4686 5990 4688
rect 5910 4670 5990 4686
rect 6017 4684 6052 4697
rect 6093 4694 6130 4697
rect 6093 4692 6135 4694
rect 6022 4681 6052 4684
rect 6031 4677 6038 4681
rect 6038 4676 6039 4677
rect 5997 4670 6007 4676
rect 5756 4662 5791 4670
rect 5756 4636 5757 4662
rect 5764 4636 5791 4662
rect 5699 4618 5729 4632
rect 5756 4628 5791 4636
rect 5793 4662 5834 4670
rect 5793 4636 5808 4662
rect 5815 4636 5834 4662
rect 5898 4658 5929 4670
rect 5944 4658 6047 4670
rect 6059 4660 6085 4686
rect 6100 4681 6130 4692
rect 6162 4688 6224 4704
rect 6162 4686 6208 4688
rect 6162 4670 6224 4686
rect 6236 4670 6242 4718
rect 6245 4710 6325 4718
rect 6245 4708 6264 4710
rect 6279 4708 6313 4710
rect 6245 4692 6325 4708
rect 6245 4670 6264 4692
rect 6279 4676 6309 4692
rect 6337 4686 6343 4760
rect 6346 4686 6365 4830
rect 6380 4686 6386 4830
rect 6395 4760 6408 4830
rect 6460 4826 6482 4830
rect 6453 4804 6482 4818
rect 6535 4804 6551 4818
rect 6589 4814 6595 4816
rect 6602 4814 6710 4830
rect 6717 4814 6723 4816
rect 6731 4814 6746 4830
rect 6812 4824 6831 4827
rect 6453 4802 6551 4804
rect 6578 4802 6746 4814
rect 6761 4804 6777 4818
rect 6812 4805 6834 4824
rect 6844 4818 6860 4819
rect 6843 4816 6860 4818
rect 6844 4811 6860 4816
rect 6834 4804 6840 4805
rect 6843 4804 6872 4811
rect 6761 4803 6872 4804
rect 6761 4802 6878 4803
rect 6437 4794 6488 4802
rect 6535 4794 6569 4802
rect 6437 4782 6462 4794
rect 6469 4782 6488 4794
rect 6542 4792 6569 4794
rect 6578 4792 6799 4802
rect 6834 4799 6840 4802
rect 6542 4788 6799 4792
rect 6437 4774 6488 4782
rect 6535 4774 6799 4788
rect 6843 4794 6878 4802
rect 6389 4726 6408 4760
rect 6453 4766 6482 4774
rect 6453 4760 6470 4766
rect 6453 4758 6487 4760
rect 6535 4758 6551 4774
rect 6552 4764 6760 4774
rect 6761 4764 6777 4774
rect 6825 4770 6840 4785
rect 6843 4782 6844 4794
rect 6851 4782 6878 4794
rect 6843 4774 6878 4782
rect 6843 4773 6872 4774
rect 6563 4760 6777 4764
rect 6578 4758 6777 4760
rect 6812 4760 6825 4770
rect 6843 4760 6860 4773
rect 6812 4758 6860 4760
rect 6454 4754 6487 4758
rect 6450 4752 6487 4754
rect 6450 4751 6517 4752
rect 6450 4746 6481 4751
rect 6487 4746 6517 4751
rect 6450 4742 6517 4746
rect 6423 4739 6517 4742
rect 6423 4732 6472 4739
rect 6423 4726 6453 4732
rect 6472 4727 6477 4732
rect 6389 4710 6469 4726
rect 6481 4718 6517 4739
rect 6578 4734 6767 4758
rect 6812 4757 6859 4758
rect 6825 4752 6859 4757
rect 6593 4731 6767 4734
rect 6586 4728 6767 4731
rect 6795 4751 6859 4752
rect 6389 4708 6408 4710
rect 6423 4708 6457 4710
rect 6389 4692 6469 4708
rect 6389 4686 6408 4692
rect 6105 4660 6208 4670
rect 6059 4658 6208 4660
rect 6229 4658 6264 4670
rect 5898 4656 6060 4658
rect 5910 4636 5929 4656
rect 5944 4654 5974 4656
rect 5793 4628 5834 4636
rect 5916 4632 5929 4636
rect 5981 4640 6060 4656
rect 6092 4656 6264 4658
rect 6092 4640 6171 4656
rect 6178 4654 6208 4656
rect 5756 4618 5785 4628
rect 5799 4618 5828 4628
rect 5843 4618 5873 4632
rect 5916 4618 5959 4632
rect 5981 4628 6171 4640
rect 6236 4636 6242 4656
rect 5966 4618 5996 4628
rect 5997 4618 6155 4628
rect 6159 4618 6189 4628
rect 6193 4618 6223 4632
rect 6251 4618 6264 4656
rect 6336 4670 6365 4686
rect 6379 4670 6408 4686
rect 6423 4676 6453 4692
rect 6481 4670 6487 4718
rect 6490 4712 6509 4718
rect 6524 4712 6554 4720
rect 6490 4704 6554 4712
rect 6490 4688 6570 4704
rect 6586 4697 6648 4728
rect 6664 4697 6726 4728
rect 6795 4726 6844 4751
rect 6859 4726 6889 4742
rect 6758 4712 6788 4720
rect 6795 4718 6905 4726
rect 6758 4704 6803 4712
rect 6490 4686 6509 4688
rect 6524 4686 6570 4688
rect 6490 4670 6570 4686
rect 6597 4684 6632 4697
rect 6673 4694 6710 4697
rect 6673 4692 6715 4694
rect 6602 4681 6632 4684
rect 6611 4677 6618 4681
rect 6618 4676 6619 4677
rect 6577 4670 6587 4676
rect 6336 4662 6371 4670
rect 6336 4636 6337 4662
rect 6344 4636 6371 4662
rect 6279 4618 6309 4632
rect 6336 4628 6371 4636
rect 6373 4662 6414 4670
rect 6373 4636 6388 4662
rect 6395 4636 6414 4662
rect 6478 4658 6509 4670
rect 6524 4658 6627 4670
rect 6639 4660 6665 4686
rect 6680 4681 6710 4692
rect 6742 4688 6804 4704
rect 6742 4686 6788 4688
rect 6742 4670 6804 4686
rect 6816 4670 6822 4718
rect 6825 4710 6905 4718
rect 6825 4708 6844 4710
rect 6859 4708 6893 4710
rect 6825 4692 6905 4708
rect 6825 4670 6844 4692
rect 6859 4676 6889 4692
rect 6917 4686 6923 4760
rect 6926 4686 6945 4830
rect 6960 4686 6966 4830
rect 6975 4760 6988 4830
rect 7040 4826 7062 4830
rect 7033 4804 7062 4818
rect 7115 4804 7131 4818
rect 7169 4814 7175 4816
rect 7182 4814 7290 4830
rect 7297 4814 7303 4816
rect 7311 4814 7326 4830
rect 7392 4824 7411 4827
rect 7033 4802 7131 4804
rect 7158 4802 7326 4814
rect 7341 4804 7357 4818
rect 7392 4805 7414 4824
rect 7424 4818 7440 4819
rect 7423 4816 7440 4818
rect 7424 4811 7440 4816
rect 7414 4804 7420 4805
rect 7423 4804 7452 4811
rect 7341 4803 7452 4804
rect 7341 4802 7458 4803
rect 7017 4794 7068 4802
rect 7115 4794 7149 4802
rect 7017 4782 7042 4794
rect 7049 4782 7068 4794
rect 7122 4792 7149 4794
rect 7158 4792 7379 4802
rect 7414 4799 7420 4802
rect 7122 4788 7379 4792
rect 7017 4774 7068 4782
rect 7115 4774 7379 4788
rect 7423 4794 7458 4802
rect 6969 4726 6988 4760
rect 7033 4766 7062 4774
rect 7033 4760 7050 4766
rect 7033 4758 7067 4760
rect 7115 4758 7131 4774
rect 7132 4764 7340 4774
rect 7341 4764 7357 4774
rect 7405 4770 7420 4785
rect 7423 4782 7424 4794
rect 7431 4782 7458 4794
rect 7423 4774 7458 4782
rect 7423 4773 7452 4774
rect 7143 4760 7357 4764
rect 7158 4758 7357 4760
rect 7392 4760 7405 4770
rect 7423 4760 7440 4773
rect 7392 4758 7440 4760
rect 7034 4754 7067 4758
rect 7030 4752 7067 4754
rect 7030 4751 7097 4752
rect 7030 4746 7061 4751
rect 7067 4746 7097 4751
rect 7030 4742 7097 4746
rect 7003 4739 7097 4742
rect 7003 4732 7052 4739
rect 7003 4726 7033 4732
rect 7052 4727 7057 4732
rect 6969 4710 7049 4726
rect 7061 4718 7097 4739
rect 7158 4734 7347 4758
rect 7392 4757 7439 4758
rect 7405 4752 7439 4757
rect 7173 4731 7347 4734
rect 7166 4728 7347 4731
rect 7375 4751 7439 4752
rect 6969 4708 6988 4710
rect 7003 4708 7037 4710
rect 6969 4692 7049 4708
rect 6969 4686 6988 4692
rect 6685 4660 6788 4670
rect 6639 4658 6788 4660
rect 6809 4658 6844 4670
rect 6478 4656 6640 4658
rect 6490 4636 6509 4656
rect 6524 4654 6554 4656
rect 6373 4628 6414 4636
rect 6496 4632 6509 4636
rect 6561 4640 6640 4656
rect 6672 4656 6844 4658
rect 6672 4640 6751 4656
rect 6758 4654 6788 4656
rect 6336 4618 6365 4628
rect 6379 4618 6408 4628
rect 6423 4618 6453 4632
rect 6496 4618 6539 4632
rect 6561 4628 6751 4640
rect 6816 4636 6822 4656
rect 6546 4618 6576 4628
rect 6577 4618 6735 4628
rect 6739 4618 6769 4628
rect 6773 4618 6803 4632
rect 6831 4618 6844 4656
rect 6916 4670 6945 4686
rect 6959 4670 6988 4686
rect 7003 4676 7033 4692
rect 7061 4670 7067 4718
rect 7070 4712 7089 4718
rect 7104 4712 7134 4720
rect 7070 4704 7134 4712
rect 7070 4688 7150 4704
rect 7166 4697 7228 4728
rect 7244 4697 7306 4728
rect 7375 4726 7424 4751
rect 7439 4726 7469 4742
rect 7338 4712 7368 4720
rect 7375 4718 7485 4726
rect 7338 4704 7383 4712
rect 7070 4686 7089 4688
rect 7104 4686 7150 4688
rect 7070 4670 7150 4686
rect 7177 4684 7212 4697
rect 7253 4694 7290 4697
rect 7253 4692 7295 4694
rect 7182 4681 7212 4684
rect 7191 4677 7198 4681
rect 7198 4676 7199 4677
rect 7157 4670 7167 4676
rect 6916 4662 6951 4670
rect 6916 4636 6917 4662
rect 6924 4636 6951 4662
rect 6859 4618 6889 4632
rect 6916 4628 6951 4636
rect 6953 4662 6994 4670
rect 6953 4636 6968 4662
rect 6975 4636 6994 4662
rect 7058 4658 7089 4670
rect 7104 4658 7207 4670
rect 7219 4660 7245 4686
rect 7260 4681 7290 4692
rect 7322 4688 7384 4704
rect 7322 4686 7368 4688
rect 7322 4670 7384 4686
rect 7396 4670 7402 4718
rect 7405 4710 7485 4718
rect 7405 4708 7424 4710
rect 7439 4708 7473 4710
rect 7405 4692 7485 4708
rect 7405 4670 7424 4692
rect 7439 4676 7469 4692
rect 7497 4686 7503 4760
rect 7506 4686 7525 4830
rect 7540 4686 7546 4830
rect 7555 4760 7568 4830
rect 7613 4808 7614 4818
rect 7629 4808 7642 4818
rect 7613 4804 7642 4808
rect 7647 4804 7677 4830
rect 7695 4816 7711 4818
rect 7783 4816 7836 4830
rect 7784 4814 7848 4816
rect 7891 4814 7906 4830
rect 7955 4827 7985 4830
rect 7955 4824 7991 4827
rect 7921 4816 7937 4818
rect 7695 4804 7710 4808
rect 7613 4802 7710 4804
rect 7738 4802 7906 4814
rect 7922 4804 7937 4808
rect 7955 4805 7994 4824
rect 8013 4818 8020 4819
rect 8019 4811 8020 4818
rect 8003 4808 8004 4811
rect 8019 4808 8032 4811
rect 7955 4804 7985 4805
rect 7994 4804 8000 4805
rect 8003 4804 8032 4808
rect 7922 4803 8032 4804
rect 7922 4802 8038 4803
rect 7597 4794 7648 4802
rect 7597 4782 7622 4794
rect 7629 4782 7648 4794
rect 7679 4794 7729 4802
rect 7679 4786 7695 4794
rect 7702 4792 7729 4794
rect 7738 4792 7959 4802
rect 7702 4782 7959 4792
rect 7988 4794 8038 4802
rect 7988 4785 8004 4794
rect 7597 4774 7648 4782
rect 7695 4774 7959 4782
rect 7985 4782 8004 4785
rect 8011 4782 8038 4794
rect 7985 4774 8038 4782
rect 7549 4726 7568 4760
rect 7613 4766 7614 4774
rect 7629 4766 7642 4774
rect 7613 4758 7629 4766
rect 7610 4751 7629 4754
rect 7610 4742 7632 4751
rect 7583 4732 7632 4742
rect 7583 4726 7613 4732
rect 7632 4727 7637 4732
rect 7549 4710 7629 4726
rect 7647 4718 7677 4774
rect 7712 4764 7920 4774
rect 7955 4770 8000 4774
rect 8003 4773 8004 4774
rect 8019 4773 8032 4774
rect 7738 4734 7927 4764
rect 7753 4731 7927 4734
rect 7746 4728 7927 4731
rect 7549 4708 7568 4710
rect 7583 4708 7617 4710
rect 7549 4692 7629 4708
rect 7656 4704 7669 4718
rect 7684 4704 7700 4720
rect 7746 4715 7757 4728
rect 7549 4686 7568 4692
rect 7265 4660 7368 4670
rect 7219 4658 7368 4660
rect 7389 4658 7424 4670
rect 7058 4656 7220 4658
rect 7070 4636 7089 4656
rect 7104 4654 7134 4656
rect 6953 4628 6994 4636
rect 7076 4632 7089 4636
rect 7141 4640 7220 4656
rect 7252 4656 7424 4658
rect 7252 4640 7331 4656
rect 7338 4654 7368 4656
rect 6916 4618 6945 4628
rect 6959 4618 6988 4628
rect 7003 4618 7033 4632
rect 7076 4618 7119 4632
rect 7141 4628 7331 4640
rect 7396 4636 7402 4656
rect 7126 4618 7156 4628
rect 7157 4618 7315 4628
rect 7319 4618 7349 4628
rect 7353 4618 7383 4632
rect 7411 4618 7424 4656
rect 7496 4670 7525 4686
rect 7539 4670 7568 4686
rect 7583 4670 7613 4692
rect 7656 4688 7718 4704
rect 7746 4697 7757 4713
rect 7762 4708 7772 4728
rect 7782 4708 7796 4728
rect 7799 4715 7808 4728
rect 7824 4715 7833 4728
rect 7762 4697 7796 4708
rect 7799 4697 7808 4713
rect 7824 4697 7833 4713
rect 7840 4708 7850 4728
rect 7860 4708 7874 4728
rect 7875 4715 7886 4728
rect 7840 4697 7874 4708
rect 7875 4697 7886 4713
rect 7932 4704 7948 4720
rect 7955 4718 7985 4770
rect 8019 4766 8020 4773
rect 8004 4758 8020 4766
rect 7991 4726 8004 4745
rect 8019 4726 8049 4742
rect 7991 4710 8065 4726
rect 7991 4708 8004 4710
rect 8019 4708 8053 4710
rect 7656 4686 7669 4688
rect 7684 4686 7718 4688
rect 7656 4670 7718 4686
rect 7762 4681 7778 4684
rect 7840 4681 7870 4692
rect 7918 4688 7964 4704
rect 7991 4692 8065 4708
rect 7918 4686 7952 4688
rect 7917 4670 7964 4686
rect 7991 4670 8004 4692
rect 8019 4670 8049 4692
rect 8076 4670 8077 4686
rect 8092 4670 8105 4830
rect 8135 4726 8148 4830
rect 8193 4808 8194 4818
rect 8209 4808 8222 4818
rect 8193 4804 8222 4808
rect 8227 4804 8257 4830
rect 8275 4816 8291 4818
rect 8363 4816 8416 4830
rect 8364 4814 8428 4816
rect 8471 4814 8486 4830
rect 8535 4827 8565 4830
rect 8535 4824 8571 4827
rect 8501 4816 8517 4818
rect 8275 4804 8290 4808
rect 8193 4802 8290 4804
rect 8318 4802 8486 4814
rect 8502 4804 8517 4808
rect 8535 4805 8574 4824
rect 8593 4818 8600 4819
rect 8599 4811 8600 4818
rect 8583 4808 8584 4811
rect 8599 4808 8612 4811
rect 8535 4804 8565 4805
rect 8574 4804 8580 4805
rect 8583 4804 8612 4808
rect 8502 4803 8612 4804
rect 8502 4802 8618 4803
rect 8177 4794 8228 4802
rect 8177 4782 8202 4794
rect 8209 4782 8228 4794
rect 8259 4794 8309 4802
rect 8259 4786 8275 4794
rect 8282 4792 8309 4794
rect 8318 4792 8539 4802
rect 8282 4782 8539 4792
rect 8568 4794 8618 4802
rect 8568 4785 8584 4794
rect 8177 4774 8228 4782
rect 8275 4774 8539 4782
rect 8565 4782 8584 4785
rect 8591 4782 8618 4794
rect 8565 4774 8618 4782
rect 8193 4766 8194 4774
rect 8209 4766 8222 4774
rect 8193 4758 8209 4766
rect 8190 4751 8209 4754
rect 8190 4742 8212 4751
rect 8163 4732 8212 4742
rect 8163 4726 8193 4732
rect 8212 4727 8217 4732
rect 8135 4710 8209 4726
rect 8227 4718 8257 4774
rect 8292 4764 8500 4774
rect 8535 4770 8580 4774
rect 8583 4773 8584 4774
rect 8599 4773 8612 4774
rect 8318 4734 8507 4764
rect 8333 4731 8507 4734
rect 8326 4728 8507 4731
rect 8135 4708 8148 4710
rect 8163 4708 8197 4710
rect 8135 4692 8209 4708
rect 8236 4704 8249 4718
rect 8264 4704 8280 4720
rect 8326 4715 8337 4728
rect 8119 4670 8120 4686
rect 8135 4670 8148 4692
rect 8163 4670 8193 4692
rect 8236 4688 8298 4704
rect 8326 4697 8337 4713
rect 8342 4708 8352 4728
rect 8362 4708 8376 4728
rect 8379 4715 8388 4728
rect 8404 4715 8413 4728
rect 8342 4697 8376 4708
rect 8379 4697 8388 4713
rect 8404 4697 8413 4713
rect 8420 4708 8430 4728
rect 8440 4708 8454 4728
rect 8455 4715 8466 4728
rect 8420 4697 8454 4708
rect 8455 4697 8466 4713
rect 8512 4704 8528 4720
rect 8535 4718 8565 4770
rect 8599 4766 8600 4773
rect 8584 4758 8600 4766
rect 8571 4726 8584 4745
rect 8599 4726 8629 4742
rect 8571 4710 8645 4726
rect 8571 4708 8584 4710
rect 8599 4708 8633 4710
rect 8236 4686 8249 4688
rect 8264 4686 8298 4688
rect 8236 4670 8298 4686
rect 8342 4681 8358 4684
rect 8420 4681 8450 4692
rect 8498 4688 8544 4704
rect 8571 4692 8645 4708
rect 8498 4686 8532 4688
rect 8497 4670 8544 4686
rect 8571 4670 8584 4692
rect 8599 4670 8629 4692
rect 8656 4670 8657 4686
rect 8672 4670 8685 4830
rect 8715 4726 8728 4830
rect 8773 4808 8774 4818
rect 8789 4808 8802 4818
rect 8773 4804 8802 4808
rect 8807 4804 8837 4830
rect 8855 4816 8871 4818
rect 8943 4816 8996 4830
rect 8944 4814 9008 4816
rect 9051 4814 9066 4830
rect 9115 4827 9145 4830
rect 9115 4824 9151 4827
rect 9081 4816 9097 4818
rect 8855 4804 8870 4808
rect 8773 4802 8870 4804
rect 8898 4802 9066 4814
rect 9082 4804 9097 4808
rect 9115 4805 9154 4824
rect 9173 4818 9180 4819
rect 9179 4811 9180 4818
rect 9163 4808 9164 4811
rect 9179 4808 9192 4811
rect 9115 4804 9145 4805
rect 9154 4804 9160 4805
rect 9163 4804 9192 4808
rect 9082 4803 9192 4804
rect 9082 4802 9198 4803
rect 8757 4794 8808 4802
rect 8757 4782 8782 4794
rect 8789 4782 8808 4794
rect 8839 4794 8889 4802
rect 8839 4786 8855 4794
rect 8862 4792 8889 4794
rect 8898 4792 9119 4802
rect 8862 4782 9119 4792
rect 9148 4794 9198 4802
rect 9148 4785 9164 4794
rect 8757 4774 8808 4782
rect 8855 4774 9119 4782
rect 9145 4782 9164 4785
rect 9171 4782 9198 4794
rect 9145 4774 9198 4782
rect 8773 4766 8774 4774
rect 8789 4766 8802 4774
rect 8773 4758 8789 4766
rect 8770 4751 8789 4754
rect 8770 4742 8792 4751
rect 8743 4732 8792 4742
rect 8743 4726 8773 4732
rect 8792 4727 8797 4732
rect 8715 4710 8789 4726
rect 8807 4718 8837 4774
rect 8872 4764 9080 4774
rect 9115 4770 9160 4774
rect 9163 4773 9164 4774
rect 9179 4773 9192 4774
rect 8898 4734 9087 4764
rect 8913 4731 9087 4734
rect 8906 4728 9087 4731
rect 8715 4708 8728 4710
rect 8743 4708 8777 4710
rect 8715 4692 8789 4708
rect 8816 4704 8829 4718
rect 8844 4704 8860 4720
rect 8906 4715 8917 4728
rect 8699 4670 8700 4686
rect 8715 4670 8728 4692
rect 8743 4670 8773 4692
rect 8816 4688 8878 4704
rect 8906 4697 8917 4713
rect 8922 4708 8932 4728
rect 8942 4708 8956 4728
rect 8959 4715 8968 4728
rect 8984 4715 8993 4728
rect 8922 4697 8956 4708
rect 8959 4697 8968 4713
rect 8984 4697 8993 4713
rect 9000 4708 9010 4728
rect 9020 4708 9034 4728
rect 9035 4715 9046 4728
rect 9000 4697 9034 4708
rect 9035 4697 9046 4713
rect 9092 4704 9108 4720
rect 9115 4718 9145 4770
rect 9179 4766 9180 4773
rect 9164 4758 9180 4766
rect 9151 4726 9164 4745
rect 9179 4726 9209 4742
rect 9151 4710 9225 4726
rect 9151 4708 9164 4710
rect 9179 4708 9213 4710
rect 8816 4686 8829 4688
rect 8844 4686 8878 4688
rect 8816 4670 8878 4686
rect 8922 4681 8938 4684
rect 9000 4681 9030 4692
rect 9078 4688 9124 4704
rect 9151 4692 9225 4708
rect 9078 4686 9112 4688
rect 9077 4670 9124 4686
rect 9151 4670 9164 4692
rect 9179 4670 9209 4692
rect 9236 4670 9237 4686
rect 9252 4670 9265 4830
rect 7496 4662 7531 4670
rect 7496 4636 7497 4662
rect 7504 4636 7531 4662
rect 7439 4618 7469 4632
rect 7496 4628 7531 4636
rect 7533 4662 7574 4670
rect 7533 4636 7548 4662
rect 7555 4636 7574 4662
rect 7638 4658 7700 4670
rect 7712 4658 7787 4670
rect 7845 4658 7920 4670
rect 7932 4658 7963 4670
rect 7969 4658 8004 4670
rect 7638 4656 7800 4658
rect 7533 4628 7574 4636
rect 7656 4632 7669 4656
rect 7684 4654 7699 4656
rect 7496 4618 7525 4628
rect 7539 4618 7568 4628
rect 7583 4618 7613 4632
rect 7656 4618 7699 4632
rect 7723 4629 7730 4636
rect 7733 4632 7800 4656
rect 7832 4656 8004 4658
rect 7802 4634 7830 4638
rect 7832 4634 7912 4656
rect 7933 4654 7948 4656
rect 7802 4632 7912 4634
rect 7733 4628 7912 4632
rect 7706 4618 7736 4628
rect 7738 4618 7891 4628
rect 7899 4618 7929 4628
rect 7933 4618 7963 4632
rect 7991 4618 8004 4656
rect 8076 4662 8111 4670
rect 8076 4636 8077 4662
rect 8084 4636 8111 4662
rect 8019 4618 8049 4632
rect 8076 4628 8111 4636
rect 8113 4662 8154 4670
rect 8113 4636 8128 4662
rect 8135 4636 8154 4662
rect 8218 4658 8280 4670
rect 8292 4658 8367 4670
rect 8425 4658 8500 4670
rect 8512 4658 8543 4670
rect 8549 4658 8584 4670
rect 8218 4656 8380 4658
rect 8113 4628 8154 4636
rect 8236 4632 8249 4656
rect 8264 4654 8279 4656
rect 8076 4618 8077 4628
rect 8092 4618 8105 4628
rect 8119 4618 8120 4628
rect 8135 4618 8148 4628
rect 8163 4618 8193 4632
rect 8236 4618 8279 4632
rect 8303 4629 8310 4636
rect 8313 4632 8380 4656
rect 8412 4656 8584 4658
rect 8382 4634 8410 4638
rect 8412 4634 8492 4656
rect 8513 4654 8528 4656
rect 8382 4632 8492 4634
rect 8313 4628 8492 4632
rect 8286 4618 8316 4628
rect 8318 4618 8471 4628
rect 8479 4618 8509 4628
rect 8513 4618 8543 4632
rect 8571 4618 8584 4656
rect 8656 4662 8691 4670
rect 8656 4636 8657 4662
rect 8664 4636 8691 4662
rect 8599 4618 8629 4632
rect 8656 4628 8691 4636
rect 8693 4662 8734 4670
rect 8693 4636 8708 4662
rect 8715 4636 8734 4662
rect 8798 4658 8860 4670
rect 8872 4658 8947 4670
rect 9005 4658 9080 4670
rect 9092 4658 9123 4670
rect 9129 4658 9164 4670
rect 8798 4656 8960 4658
rect 8693 4628 8734 4636
rect 8816 4632 8829 4656
rect 8844 4654 8859 4656
rect 8656 4618 8657 4628
rect 8672 4618 8685 4628
rect 8699 4618 8700 4628
rect 8715 4618 8728 4628
rect 8743 4618 8773 4632
rect 8816 4618 8859 4632
rect 8883 4629 8890 4636
rect 8893 4632 8960 4656
rect 8992 4656 9164 4658
rect 8962 4634 8990 4638
rect 8992 4634 9072 4656
rect 9093 4654 9108 4656
rect 8962 4632 9072 4634
rect 8893 4628 9072 4632
rect 8866 4618 8896 4628
rect 8898 4618 9051 4628
rect 9059 4618 9089 4628
rect 9093 4618 9123 4632
rect 9151 4618 9164 4656
rect 9236 4662 9271 4670
rect 9236 4636 9237 4662
rect 9244 4636 9271 4662
rect 9179 4618 9209 4632
rect 9236 4628 9271 4636
rect 9236 4618 9237 4628
rect 9252 4618 9265 4628
rect -1 4612 9265 4618
rect 0 4604 9265 4612
rect 15 4574 28 4604
rect 43 4590 73 4604
rect 116 4590 159 4604
rect 166 4590 386 4604
rect 393 4590 423 4604
rect 83 4576 98 4588
rect 117 4576 130 4590
rect 198 4586 351 4590
rect 80 4574 102 4576
rect 180 4574 372 4586
rect 451 4574 464 4604
rect 479 4590 509 4604
rect 546 4574 565 4604
rect 580 4574 586 4604
rect 595 4574 608 4604
rect 623 4590 653 4604
rect 696 4590 739 4604
rect 746 4590 966 4604
rect 973 4590 1003 4604
rect 663 4576 678 4588
rect 697 4576 710 4590
rect 778 4586 931 4590
rect 660 4574 682 4576
rect 760 4574 952 4586
rect 1031 4574 1044 4604
rect 1059 4590 1089 4604
rect 1126 4574 1145 4604
rect 1160 4574 1166 4604
rect 1175 4574 1188 4604
rect 1203 4590 1233 4604
rect 1276 4590 1319 4604
rect 1326 4590 1546 4604
rect 1553 4590 1583 4604
rect 1243 4576 1258 4588
rect 1277 4576 1290 4590
rect 1358 4586 1511 4590
rect 1240 4574 1262 4576
rect 1340 4574 1532 4586
rect 1611 4574 1624 4604
rect 1639 4590 1669 4604
rect 1706 4574 1725 4604
rect 1740 4574 1746 4604
rect 1755 4574 1768 4604
rect 1783 4590 1813 4604
rect 1856 4590 1899 4604
rect 1906 4590 2126 4604
rect 2133 4590 2163 4604
rect 1823 4576 1838 4588
rect 1857 4576 1870 4590
rect 1938 4586 2091 4590
rect 1820 4574 1842 4576
rect 1920 4574 2112 4586
rect 2191 4574 2204 4604
rect 2219 4590 2249 4604
rect 2286 4574 2305 4604
rect 2320 4574 2326 4604
rect 2335 4574 2348 4604
rect 2363 4590 2393 4604
rect 2436 4590 2479 4604
rect 2486 4590 2706 4604
rect 2713 4590 2743 4604
rect 2403 4576 2418 4588
rect 2437 4576 2450 4590
rect 2518 4586 2671 4590
rect 2400 4574 2422 4576
rect 2500 4574 2692 4586
rect 2771 4574 2784 4604
rect 2799 4590 2829 4604
rect 2866 4574 2885 4604
rect 2900 4574 2906 4604
rect 2915 4574 2928 4604
rect 2943 4590 2973 4604
rect 3016 4590 3059 4604
rect 3066 4590 3286 4604
rect 3293 4590 3323 4604
rect 2983 4576 2998 4588
rect 3017 4576 3030 4590
rect 3098 4586 3251 4590
rect 2980 4574 3002 4576
rect 3080 4574 3272 4586
rect 3351 4574 3364 4604
rect 3379 4590 3409 4604
rect 3446 4574 3465 4604
rect 3480 4574 3486 4604
rect 3495 4574 3508 4604
rect 3523 4590 3553 4604
rect 3596 4590 3639 4604
rect 3646 4590 3866 4604
rect 3873 4590 3903 4604
rect 3563 4576 3578 4588
rect 3597 4576 3610 4590
rect 3678 4586 3831 4590
rect 3560 4574 3582 4576
rect 3660 4574 3852 4586
rect 3931 4574 3944 4604
rect 3959 4590 3989 4604
rect 4026 4574 4045 4604
rect 4060 4574 4066 4604
rect 4075 4574 4088 4604
rect 4103 4590 4133 4604
rect 4176 4590 4219 4604
rect 4226 4590 4446 4604
rect 4453 4590 4483 4604
rect 4143 4576 4158 4588
rect 4177 4576 4190 4590
rect 4258 4586 4411 4590
rect 4140 4574 4162 4576
rect 4240 4574 4432 4586
rect 4511 4574 4524 4604
rect 4539 4590 4569 4604
rect 4606 4574 4625 4604
rect 4640 4574 4646 4604
rect 4655 4574 4668 4604
rect 4683 4590 4713 4604
rect 4756 4590 4799 4604
rect 4806 4590 5026 4604
rect 5033 4590 5063 4604
rect 4723 4576 4738 4588
rect 4757 4576 4770 4590
rect 4838 4586 4991 4590
rect 4720 4574 4742 4576
rect 4820 4574 5012 4586
rect 5091 4574 5104 4604
rect 5119 4590 5149 4604
rect 5186 4574 5205 4604
rect 5220 4574 5226 4604
rect 5235 4574 5248 4604
rect 5263 4590 5293 4604
rect 5336 4590 5379 4604
rect 5386 4590 5606 4604
rect 5613 4590 5643 4604
rect 5303 4576 5318 4588
rect 5337 4576 5350 4590
rect 5418 4586 5571 4590
rect 5300 4574 5322 4576
rect 5400 4574 5592 4586
rect 5671 4574 5684 4604
rect 5699 4590 5729 4604
rect 5766 4574 5785 4604
rect 5800 4574 5806 4604
rect 5815 4574 5828 4604
rect 5843 4590 5873 4604
rect 5916 4590 5959 4604
rect 5966 4590 6186 4604
rect 6193 4590 6223 4604
rect 5883 4576 5898 4588
rect 5917 4576 5930 4590
rect 5998 4586 6151 4590
rect 5880 4574 5902 4576
rect 5980 4574 6172 4586
rect 6251 4574 6264 4604
rect 6279 4590 6309 4604
rect 6346 4574 6365 4604
rect 6380 4574 6386 4604
rect 6395 4574 6408 4604
rect 6423 4590 6453 4604
rect 6496 4590 6539 4604
rect 6546 4590 6766 4604
rect 6773 4590 6803 4604
rect 6463 4576 6478 4588
rect 6497 4576 6510 4590
rect 6578 4586 6731 4590
rect 6460 4574 6482 4576
rect 6560 4574 6752 4586
rect 6831 4574 6844 4604
rect 6859 4590 6889 4604
rect 6926 4574 6945 4604
rect 6960 4574 6966 4604
rect 6975 4574 6988 4604
rect 7003 4590 7033 4604
rect 7076 4590 7119 4604
rect 7126 4590 7346 4604
rect 7353 4590 7383 4604
rect 7043 4576 7058 4588
rect 7077 4576 7090 4590
rect 7158 4586 7311 4590
rect 7040 4574 7062 4576
rect 7140 4574 7332 4586
rect 7411 4574 7424 4604
rect 7439 4590 7469 4604
rect 7506 4574 7525 4604
rect 7540 4574 7546 4604
rect 7555 4574 7568 4604
rect 7583 4586 7613 4604
rect 7656 4590 7670 4604
rect 7706 4590 7926 4604
rect 7657 4588 7670 4590
rect 7623 4576 7638 4588
rect 7620 4574 7642 4576
rect 7647 4574 7677 4588
rect 7738 4586 7891 4590
rect 7720 4574 7912 4586
rect 7955 4574 7985 4588
rect 7991 4574 8004 4604
rect 8019 4586 8049 4604
rect 8092 4574 8105 4604
rect 8135 4574 8148 4604
rect 8163 4586 8193 4604
rect 8236 4590 8250 4604
rect 8286 4590 8506 4604
rect 8237 4588 8250 4590
rect 8203 4576 8218 4588
rect 8200 4574 8222 4576
rect 8227 4574 8257 4588
rect 8318 4586 8471 4590
rect 8300 4574 8492 4586
rect 8535 4574 8565 4588
rect 8571 4574 8584 4604
rect 8599 4586 8629 4604
rect 8672 4574 8685 4604
rect 8715 4574 8728 4604
rect 8743 4586 8773 4604
rect 8816 4590 8830 4604
rect 8866 4590 9086 4604
rect 8817 4588 8830 4590
rect 8783 4576 8798 4588
rect 8780 4574 8802 4576
rect 8807 4574 8837 4588
rect 8898 4586 9051 4590
rect 8880 4574 9072 4586
rect 9115 4574 9145 4588
rect 9151 4574 9164 4604
rect 9179 4586 9209 4604
rect 9252 4574 9265 4604
rect 0 4560 9265 4574
rect 15 4490 28 4560
rect 80 4556 102 4560
rect 73 4534 102 4548
rect 155 4534 171 4548
rect 209 4544 215 4546
rect 222 4544 330 4560
rect 337 4544 343 4546
rect 351 4544 366 4560
rect 432 4554 451 4557
rect 73 4532 171 4534
rect 198 4532 366 4544
rect 381 4534 397 4548
rect 432 4535 454 4554
rect 464 4548 480 4549
rect 463 4546 480 4548
rect 464 4541 480 4546
rect 454 4534 460 4535
rect 463 4534 492 4541
rect 381 4533 492 4534
rect 381 4532 498 4533
rect 57 4524 108 4532
rect 155 4524 189 4532
rect 57 4512 82 4524
rect 89 4512 108 4524
rect 162 4522 189 4524
rect 198 4522 419 4532
rect 454 4529 460 4532
rect 162 4518 419 4522
rect 57 4504 108 4512
rect 155 4504 419 4518
rect 463 4524 498 4532
rect 9 4456 28 4490
rect 73 4496 102 4504
rect 73 4490 90 4496
rect 73 4488 107 4490
rect 155 4488 171 4504
rect 172 4494 380 4504
rect 381 4494 397 4504
rect 445 4500 460 4515
rect 463 4512 464 4524
rect 471 4512 498 4524
rect 463 4504 498 4512
rect 463 4503 492 4504
rect 183 4490 397 4494
rect 198 4488 397 4490
rect 432 4490 445 4500
rect 463 4490 480 4503
rect 432 4488 480 4490
rect 74 4484 107 4488
rect 70 4482 107 4484
rect 70 4481 137 4482
rect 70 4476 101 4481
rect 107 4476 137 4481
rect 70 4472 137 4476
rect 43 4469 137 4472
rect 43 4462 92 4469
rect 43 4456 73 4462
rect 92 4457 97 4462
rect 9 4440 89 4456
rect 101 4448 137 4469
rect 198 4464 387 4488
rect 432 4487 479 4488
rect 445 4482 479 4487
rect 213 4461 387 4464
rect 206 4458 387 4461
rect 415 4481 479 4482
rect 9 4438 28 4440
rect 43 4438 77 4440
rect 9 4422 89 4438
rect 9 4416 28 4422
rect -1 4400 28 4416
rect 43 4406 73 4422
rect 101 4400 107 4448
rect 110 4442 129 4448
rect 144 4442 174 4450
rect 110 4434 174 4442
rect 110 4418 190 4434
rect 206 4427 268 4458
rect 284 4427 346 4458
rect 415 4456 464 4481
rect 479 4456 509 4472
rect 378 4442 408 4450
rect 415 4448 525 4456
rect 378 4434 423 4442
rect 110 4416 129 4418
rect 144 4416 190 4418
rect 110 4400 190 4416
rect 217 4414 252 4427
rect 293 4424 330 4427
rect 293 4422 335 4424
rect 222 4411 252 4414
rect 231 4407 238 4411
rect 238 4406 239 4407
rect 197 4400 207 4406
rect -7 4392 34 4400
rect -7 4366 8 4392
rect 15 4366 34 4392
rect 98 4388 129 4400
rect 144 4388 247 4400
rect 259 4390 285 4416
rect 300 4411 330 4422
rect 362 4418 424 4434
rect 362 4416 408 4418
rect 362 4400 424 4416
rect 436 4400 442 4448
rect 445 4440 525 4448
rect 445 4438 464 4440
rect 479 4438 513 4440
rect 445 4422 525 4438
rect 445 4400 464 4422
rect 479 4406 509 4422
rect 537 4416 543 4490
rect 546 4416 565 4560
rect 580 4416 586 4560
rect 595 4490 608 4560
rect 660 4556 682 4560
rect 653 4534 682 4548
rect 735 4534 751 4548
rect 789 4544 795 4546
rect 802 4544 910 4560
rect 917 4544 923 4546
rect 931 4544 946 4560
rect 1012 4554 1031 4557
rect 653 4532 751 4534
rect 778 4532 946 4544
rect 961 4534 977 4548
rect 1012 4535 1034 4554
rect 1044 4548 1060 4549
rect 1043 4546 1060 4548
rect 1044 4541 1060 4546
rect 1034 4534 1040 4535
rect 1043 4534 1072 4541
rect 961 4533 1072 4534
rect 961 4532 1078 4533
rect 637 4524 688 4532
rect 735 4524 769 4532
rect 637 4512 662 4524
rect 669 4512 688 4524
rect 742 4522 769 4524
rect 778 4522 999 4532
rect 1034 4529 1040 4532
rect 742 4518 999 4522
rect 637 4504 688 4512
rect 735 4504 999 4518
rect 1043 4524 1078 4532
rect 589 4456 608 4490
rect 653 4496 682 4504
rect 653 4490 670 4496
rect 653 4488 687 4490
rect 735 4488 751 4504
rect 752 4494 960 4504
rect 961 4494 977 4504
rect 1025 4500 1040 4515
rect 1043 4512 1044 4524
rect 1051 4512 1078 4524
rect 1043 4504 1078 4512
rect 1043 4503 1072 4504
rect 763 4490 977 4494
rect 778 4488 977 4490
rect 1012 4490 1025 4500
rect 1043 4490 1060 4503
rect 1012 4488 1060 4490
rect 654 4484 687 4488
rect 650 4482 687 4484
rect 650 4481 717 4482
rect 650 4476 681 4481
rect 687 4476 717 4481
rect 650 4472 717 4476
rect 623 4469 717 4472
rect 623 4462 672 4469
rect 623 4456 653 4462
rect 672 4457 677 4462
rect 589 4440 669 4456
rect 681 4448 717 4469
rect 778 4464 967 4488
rect 1012 4487 1059 4488
rect 1025 4482 1059 4487
rect 793 4461 967 4464
rect 786 4458 967 4461
rect 995 4481 1059 4482
rect 589 4438 608 4440
rect 623 4438 657 4440
rect 589 4422 669 4438
rect 589 4416 608 4422
rect 305 4390 408 4400
rect 259 4388 408 4390
rect 429 4388 464 4400
rect 98 4386 260 4388
rect 110 4366 129 4386
rect 144 4384 174 4386
rect -7 4358 34 4366
rect 116 4362 129 4366
rect 181 4370 260 4386
rect 292 4386 464 4388
rect 292 4370 371 4386
rect 378 4384 408 4386
rect -1 4348 28 4358
rect 43 4348 73 4362
rect 116 4348 159 4362
rect 181 4358 371 4370
rect 436 4366 442 4386
rect 166 4348 196 4358
rect 197 4348 355 4358
rect 359 4348 389 4358
rect 393 4348 423 4362
rect 451 4348 464 4386
rect 536 4400 565 4416
rect 579 4400 608 4416
rect 623 4406 653 4422
rect 681 4400 687 4448
rect 690 4442 709 4448
rect 724 4442 754 4450
rect 690 4434 754 4442
rect 690 4418 770 4434
rect 786 4427 848 4458
rect 864 4427 926 4458
rect 995 4456 1044 4481
rect 1059 4456 1089 4472
rect 958 4442 988 4450
rect 995 4448 1105 4456
rect 958 4434 1003 4442
rect 690 4416 709 4418
rect 724 4416 770 4418
rect 690 4400 770 4416
rect 797 4414 832 4427
rect 873 4424 910 4427
rect 873 4422 915 4424
rect 802 4411 832 4414
rect 811 4407 818 4411
rect 818 4406 819 4407
rect 777 4400 787 4406
rect 536 4392 571 4400
rect 536 4366 537 4392
rect 544 4366 571 4392
rect 479 4348 509 4362
rect 536 4358 571 4366
rect 573 4392 614 4400
rect 573 4366 588 4392
rect 595 4366 614 4392
rect 678 4388 709 4400
rect 724 4388 827 4400
rect 839 4390 865 4416
rect 880 4411 910 4422
rect 942 4418 1004 4434
rect 942 4416 988 4418
rect 942 4400 1004 4416
rect 1016 4400 1022 4448
rect 1025 4440 1105 4448
rect 1025 4438 1044 4440
rect 1059 4438 1093 4440
rect 1025 4422 1105 4438
rect 1025 4400 1044 4422
rect 1059 4406 1089 4422
rect 1117 4416 1123 4490
rect 1126 4416 1145 4560
rect 1160 4416 1166 4560
rect 1175 4490 1188 4560
rect 1240 4556 1262 4560
rect 1233 4534 1262 4548
rect 1315 4534 1331 4548
rect 1369 4544 1375 4546
rect 1382 4544 1490 4560
rect 1497 4544 1503 4546
rect 1511 4544 1526 4560
rect 1592 4554 1611 4557
rect 1233 4532 1331 4534
rect 1358 4532 1526 4544
rect 1541 4534 1557 4548
rect 1592 4535 1614 4554
rect 1624 4548 1640 4549
rect 1623 4546 1640 4548
rect 1624 4541 1640 4546
rect 1614 4534 1620 4535
rect 1623 4534 1652 4541
rect 1541 4533 1652 4534
rect 1541 4532 1658 4533
rect 1217 4524 1268 4532
rect 1315 4524 1349 4532
rect 1217 4512 1242 4524
rect 1249 4512 1268 4524
rect 1322 4522 1349 4524
rect 1358 4522 1579 4532
rect 1614 4529 1620 4532
rect 1322 4518 1579 4522
rect 1217 4504 1268 4512
rect 1315 4504 1579 4518
rect 1623 4524 1658 4532
rect 1169 4456 1188 4490
rect 1233 4496 1262 4504
rect 1233 4490 1250 4496
rect 1233 4488 1267 4490
rect 1315 4488 1331 4504
rect 1332 4494 1540 4504
rect 1541 4494 1557 4504
rect 1605 4500 1620 4515
rect 1623 4512 1624 4524
rect 1631 4512 1658 4524
rect 1623 4504 1658 4512
rect 1623 4503 1652 4504
rect 1343 4490 1557 4494
rect 1358 4488 1557 4490
rect 1592 4490 1605 4500
rect 1623 4490 1640 4503
rect 1592 4488 1640 4490
rect 1234 4484 1267 4488
rect 1230 4482 1267 4484
rect 1230 4481 1297 4482
rect 1230 4476 1261 4481
rect 1267 4476 1297 4481
rect 1230 4472 1297 4476
rect 1203 4469 1297 4472
rect 1203 4462 1252 4469
rect 1203 4456 1233 4462
rect 1252 4457 1257 4462
rect 1169 4440 1249 4456
rect 1261 4448 1297 4469
rect 1358 4464 1547 4488
rect 1592 4487 1639 4488
rect 1605 4482 1639 4487
rect 1373 4461 1547 4464
rect 1366 4458 1547 4461
rect 1575 4481 1639 4482
rect 1169 4438 1188 4440
rect 1203 4438 1237 4440
rect 1169 4422 1249 4438
rect 1169 4416 1188 4422
rect 885 4390 988 4400
rect 839 4388 988 4390
rect 1009 4388 1044 4400
rect 678 4386 840 4388
rect 690 4366 709 4386
rect 724 4384 754 4386
rect 573 4358 614 4366
rect 696 4362 709 4366
rect 761 4370 840 4386
rect 872 4386 1044 4388
rect 872 4370 951 4386
rect 958 4384 988 4386
rect 536 4348 565 4358
rect 579 4348 608 4358
rect 623 4348 653 4362
rect 696 4348 739 4362
rect 761 4358 951 4370
rect 1016 4366 1022 4386
rect 746 4348 776 4358
rect 777 4348 935 4358
rect 939 4348 969 4358
rect 973 4348 1003 4362
rect 1031 4348 1044 4386
rect 1116 4400 1145 4416
rect 1159 4400 1188 4416
rect 1203 4406 1233 4422
rect 1261 4400 1267 4448
rect 1270 4442 1289 4448
rect 1304 4442 1334 4450
rect 1270 4434 1334 4442
rect 1270 4418 1350 4434
rect 1366 4427 1428 4458
rect 1444 4427 1506 4458
rect 1575 4456 1624 4481
rect 1639 4456 1669 4472
rect 1538 4442 1568 4450
rect 1575 4448 1685 4456
rect 1538 4434 1583 4442
rect 1270 4416 1289 4418
rect 1304 4416 1350 4418
rect 1270 4400 1350 4416
rect 1377 4414 1412 4427
rect 1453 4424 1490 4427
rect 1453 4422 1495 4424
rect 1382 4411 1412 4414
rect 1391 4407 1398 4411
rect 1398 4406 1399 4407
rect 1357 4400 1367 4406
rect 1116 4392 1151 4400
rect 1116 4366 1117 4392
rect 1124 4366 1151 4392
rect 1059 4348 1089 4362
rect 1116 4358 1151 4366
rect 1153 4392 1194 4400
rect 1153 4366 1168 4392
rect 1175 4366 1194 4392
rect 1258 4388 1289 4400
rect 1304 4388 1407 4400
rect 1419 4390 1445 4416
rect 1460 4411 1490 4422
rect 1522 4418 1584 4434
rect 1522 4416 1568 4418
rect 1522 4400 1584 4416
rect 1596 4400 1602 4448
rect 1605 4440 1685 4448
rect 1605 4438 1624 4440
rect 1639 4438 1673 4440
rect 1605 4422 1685 4438
rect 1605 4400 1624 4422
rect 1639 4406 1669 4422
rect 1697 4416 1703 4490
rect 1706 4416 1725 4560
rect 1740 4416 1746 4560
rect 1755 4490 1768 4560
rect 1820 4556 1842 4560
rect 1813 4534 1842 4548
rect 1895 4534 1911 4548
rect 1949 4544 1955 4546
rect 1962 4544 2070 4560
rect 2077 4544 2083 4546
rect 2091 4544 2106 4560
rect 2172 4554 2191 4557
rect 1813 4532 1911 4534
rect 1938 4532 2106 4544
rect 2121 4534 2137 4548
rect 2172 4535 2194 4554
rect 2204 4548 2220 4549
rect 2203 4546 2220 4548
rect 2204 4541 2220 4546
rect 2194 4534 2200 4535
rect 2203 4534 2232 4541
rect 2121 4533 2232 4534
rect 2121 4532 2238 4533
rect 1797 4524 1848 4532
rect 1895 4524 1929 4532
rect 1797 4512 1822 4524
rect 1829 4512 1848 4524
rect 1902 4522 1929 4524
rect 1938 4522 2159 4532
rect 2194 4529 2200 4532
rect 1902 4518 2159 4522
rect 1797 4504 1848 4512
rect 1895 4504 2159 4518
rect 2203 4524 2238 4532
rect 1749 4456 1768 4490
rect 1813 4496 1842 4504
rect 1813 4490 1830 4496
rect 1813 4488 1847 4490
rect 1895 4488 1911 4504
rect 1912 4494 2120 4504
rect 2121 4494 2137 4504
rect 2185 4500 2200 4515
rect 2203 4512 2204 4524
rect 2211 4512 2238 4524
rect 2203 4504 2238 4512
rect 2203 4503 2232 4504
rect 1923 4490 2137 4494
rect 1938 4488 2137 4490
rect 2172 4490 2185 4500
rect 2203 4490 2220 4503
rect 2172 4488 2220 4490
rect 1814 4484 1847 4488
rect 1810 4482 1847 4484
rect 1810 4481 1877 4482
rect 1810 4476 1841 4481
rect 1847 4476 1877 4481
rect 1810 4472 1877 4476
rect 1783 4469 1877 4472
rect 1783 4462 1832 4469
rect 1783 4456 1813 4462
rect 1832 4457 1837 4462
rect 1749 4440 1829 4456
rect 1841 4448 1877 4469
rect 1938 4464 2127 4488
rect 2172 4487 2219 4488
rect 2185 4482 2219 4487
rect 1953 4461 2127 4464
rect 1946 4458 2127 4461
rect 2155 4481 2219 4482
rect 1749 4438 1768 4440
rect 1783 4438 1817 4440
rect 1749 4422 1829 4438
rect 1749 4416 1768 4422
rect 1465 4390 1568 4400
rect 1419 4388 1568 4390
rect 1589 4388 1624 4400
rect 1258 4386 1420 4388
rect 1270 4366 1289 4386
rect 1304 4384 1334 4386
rect 1153 4358 1194 4366
rect 1276 4362 1289 4366
rect 1341 4370 1420 4386
rect 1452 4386 1624 4388
rect 1452 4370 1531 4386
rect 1538 4384 1568 4386
rect 1116 4348 1145 4358
rect 1159 4348 1188 4358
rect 1203 4348 1233 4362
rect 1276 4348 1319 4362
rect 1341 4358 1531 4370
rect 1596 4366 1602 4386
rect 1326 4348 1356 4358
rect 1357 4348 1515 4358
rect 1519 4348 1549 4358
rect 1553 4348 1583 4362
rect 1611 4348 1624 4386
rect 1696 4400 1725 4416
rect 1739 4400 1768 4416
rect 1783 4406 1813 4422
rect 1841 4400 1847 4448
rect 1850 4442 1869 4448
rect 1884 4442 1914 4450
rect 1850 4434 1914 4442
rect 1850 4418 1930 4434
rect 1946 4427 2008 4458
rect 2024 4427 2086 4458
rect 2155 4456 2204 4481
rect 2219 4456 2249 4472
rect 2118 4442 2148 4450
rect 2155 4448 2265 4456
rect 2118 4434 2163 4442
rect 1850 4416 1869 4418
rect 1884 4416 1930 4418
rect 1850 4400 1930 4416
rect 1957 4414 1992 4427
rect 2033 4424 2070 4427
rect 2033 4422 2075 4424
rect 1962 4411 1992 4414
rect 1971 4407 1978 4411
rect 1978 4406 1979 4407
rect 1937 4400 1947 4406
rect 1696 4392 1731 4400
rect 1696 4366 1697 4392
rect 1704 4366 1731 4392
rect 1639 4348 1669 4362
rect 1696 4358 1731 4366
rect 1733 4392 1774 4400
rect 1733 4366 1748 4392
rect 1755 4366 1774 4392
rect 1838 4388 1869 4400
rect 1884 4388 1987 4400
rect 1999 4390 2025 4416
rect 2040 4411 2070 4422
rect 2102 4418 2164 4434
rect 2102 4416 2148 4418
rect 2102 4400 2164 4416
rect 2176 4400 2182 4448
rect 2185 4440 2265 4448
rect 2185 4438 2204 4440
rect 2219 4438 2253 4440
rect 2185 4422 2265 4438
rect 2185 4400 2204 4422
rect 2219 4406 2249 4422
rect 2277 4416 2283 4490
rect 2286 4416 2305 4560
rect 2320 4416 2326 4560
rect 2335 4490 2348 4560
rect 2400 4556 2422 4560
rect 2393 4534 2422 4548
rect 2475 4534 2491 4548
rect 2529 4544 2535 4546
rect 2542 4544 2650 4560
rect 2657 4544 2663 4546
rect 2671 4544 2686 4560
rect 2752 4554 2771 4557
rect 2393 4532 2491 4534
rect 2518 4532 2686 4544
rect 2701 4534 2717 4548
rect 2752 4535 2774 4554
rect 2784 4548 2800 4549
rect 2783 4546 2800 4548
rect 2784 4541 2800 4546
rect 2774 4534 2780 4535
rect 2783 4534 2812 4541
rect 2701 4533 2812 4534
rect 2701 4532 2818 4533
rect 2377 4524 2428 4532
rect 2475 4524 2509 4532
rect 2377 4512 2402 4524
rect 2409 4512 2428 4524
rect 2482 4522 2509 4524
rect 2518 4522 2739 4532
rect 2774 4529 2780 4532
rect 2482 4518 2739 4522
rect 2377 4504 2428 4512
rect 2475 4504 2739 4518
rect 2783 4524 2818 4532
rect 2329 4456 2348 4490
rect 2393 4496 2422 4504
rect 2393 4490 2410 4496
rect 2393 4488 2427 4490
rect 2475 4488 2491 4504
rect 2492 4494 2700 4504
rect 2701 4494 2717 4504
rect 2765 4500 2780 4515
rect 2783 4512 2784 4524
rect 2791 4512 2818 4524
rect 2783 4504 2818 4512
rect 2783 4503 2812 4504
rect 2503 4490 2717 4494
rect 2518 4488 2717 4490
rect 2752 4490 2765 4500
rect 2783 4490 2800 4503
rect 2752 4488 2800 4490
rect 2394 4484 2427 4488
rect 2390 4482 2427 4484
rect 2390 4481 2457 4482
rect 2390 4476 2421 4481
rect 2427 4476 2457 4481
rect 2390 4472 2457 4476
rect 2363 4469 2457 4472
rect 2363 4462 2412 4469
rect 2363 4456 2393 4462
rect 2412 4457 2417 4462
rect 2329 4440 2409 4456
rect 2421 4448 2457 4469
rect 2518 4464 2707 4488
rect 2752 4487 2799 4488
rect 2765 4482 2799 4487
rect 2533 4461 2707 4464
rect 2526 4458 2707 4461
rect 2735 4481 2799 4482
rect 2329 4438 2348 4440
rect 2363 4438 2397 4440
rect 2329 4422 2409 4438
rect 2329 4416 2348 4422
rect 2045 4390 2148 4400
rect 1999 4388 2148 4390
rect 2169 4388 2204 4400
rect 1838 4386 2000 4388
rect 1850 4366 1869 4386
rect 1884 4384 1914 4386
rect 1733 4358 1774 4366
rect 1856 4362 1869 4366
rect 1921 4370 2000 4386
rect 2032 4386 2204 4388
rect 2032 4370 2111 4386
rect 2118 4384 2148 4386
rect 1696 4348 1725 4358
rect 1739 4348 1768 4358
rect 1783 4348 1813 4362
rect 1856 4348 1899 4362
rect 1921 4358 2111 4370
rect 2176 4366 2182 4386
rect 1906 4348 1936 4358
rect 1937 4348 2095 4358
rect 2099 4348 2129 4358
rect 2133 4348 2163 4362
rect 2191 4348 2204 4386
rect 2276 4400 2305 4416
rect 2319 4400 2348 4416
rect 2363 4406 2393 4422
rect 2421 4400 2427 4448
rect 2430 4442 2449 4448
rect 2464 4442 2494 4450
rect 2430 4434 2494 4442
rect 2430 4418 2510 4434
rect 2526 4427 2588 4458
rect 2604 4427 2666 4458
rect 2735 4456 2784 4481
rect 2799 4456 2829 4472
rect 2698 4442 2728 4450
rect 2735 4448 2845 4456
rect 2698 4434 2743 4442
rect 2430 4416 2449 4418
rect 2464 4416 2510 4418
rect 2430 4400 2510 4416
rect 2537 4414 2572 4427
rect 2613 4424 2650 4427
rect 2613 4422 2655 4424
rect 2542 4411 2572 4414
rect 2551 4407 2558 4411
rect 2558 4406 2559 4407
rect 2517 4400 2527 4406
rect 2276 4392 2311 4400
rect 2276 4366 2277 4392
rect 2284 4366 2311 4392
rect 2219 4348 2249 4362
rect 2276 4358 2311 4366
rect 2313 4392 2354 4400
rect 2313 4366 2328 4392
rect 2335 4366 2354 4392
rect 2418 4388 2449 4400
rect 2464 4388 2567 4400
rect 2579 4390 2605 4416
rect 2620 4411 2650 4422
rect 2682 4418 2744 4434
rect 2682 4416 2728 4418
rect 2682 4400 2744 4416
rect 2756 4400 2762 4448
rect 2765 4440 2845 4448
rect 2765 4438 2784 4440
rect 2799 4438 2833 4440
rect 2765 4422 2845 4438
rect 2765 4400 2784 4422
rect 2799 4406 2829 4422
rect 2857 4416 2863 4490
rect 2866 4416 2885 4560
rect 2900 4416 2906 4560
rect 2915 4490 2928 4560
rect 2980 4556 3002 4560
rect 2973 4534 3002 4548
rect 3055 4534 3071 4548
rect 3109 4544 3115 4546
rect 3122 4544 3230 4560
rect 3237 4544 3243 4546
rect 3251 4544 3266 4560
rect 3332 4554 3351 4557
rect 2973 4532 3071 4534
rect 3098 4532 3266 4544
rect 3281 4534 3297 4548
rect 3332 4535 3354 4554
rect 3364 4548 3380 4549
rect 3363 4546 3380 4548
rect 3364 4541 3380 4546
rect 3354 4534 3360 4535
rect 3363 4534 3392 4541
rect 3281 4533 3392 4534
rect 3281 4532 3398 4533
rect 2957 4524 3008 4532
rect 3055 4524 3089 4532
rect 2957 4512 2982 4524
rect 2989 4512 3008 4524
rect 3062 4522 3089 4524
rect 3098 4522 3319 4532
rect 3354 4529 3360 4532
rect 3062 4518 3319 4522
rect 2957 4504 3008 4512
rect 3055 4504 3319 4518
rect 3363 4524 3398 4532
rect 2909 4456 2928 4490
rect 2973 4496 3002 4504
rect 2973 4490 2990 4496
rect 2973 4488 3007 4490
rect 3055 4488 3071 4504
rect 3072 4494 3280 4504
rect 3281 4494 3297 4504
rect 3345 4500 3360 4515
rect 3363 4512 3364 4524
rect 3371 4512 3398 4524
rect 3363 4504 3398 4512
rect 3363 4503 3392 4504
rect 3083 4490 3297 4494
rect 3098 4488 3297 4490
rect 3332 4490 3345 4500
rect 3363 4490 3380 4503
rect 3332 4488 3380 4490
rect 2974 4484 3007 4488
rect 2970 4482 3007 4484
rect 2970 4481 3037 4482
rect 2970 4476 3001 4481
rect 3007 4476 3037 4481
rect 2970 4472 3037 4476
rect 2943 4469 3037 4472
rect 2943 4462 2992 4469
rect 2943 4456 2973 4462
rect 2992 4457 2997 4462
rect 2909 4440 2989 4456
rect 3001 4448 3037 4469
rect 3098 4464 3287 4488
rect 3332 4487 3379 4488
rect 3345 4482 3379 4487
rect 3113 4461 3287 4464
rect 3106 4458 3287 4461
rect 3315 4481 3379 4482
rect 2909 4438 2928 4440
rect 2943 4438 2977 4440
rect 2909 4422 2989 4438
rect 2909 4416 2928 4422
rect 2625 4390 2728 4400
rect 2579 4388 2728 4390
rect 2749 4388 2784 4400
rect 2418 4386 2580 4388
rect 2430 4366 2449 4386
rect 2464 4384 2494 4386
rect 2313 4358 2354 4366
rect 2436 4362 2449 4366
rect 2501 4370 2580 4386
rect 2612 4386 2784 4388
rect 2612 4370 2691 4386
rect 2698 4384 2728 4386
rect 2276 4348 2305 4358
rect 2319 4348 2348 4358
rect 2363 4348 2393 4362
rect 2436 4348 2479 4362
rect 2501 4358 2691 4370
rect 2756 4366 2762 4386
rect 2486 4348 2516 4358
rect 2517 4348 2675 4358
rect 2679 4348 2709 4358
rect 2713 4348 2743 4362
rect 2771 4348 2784 4386
rect 2856 4400 2885 4416
rect 2899 4400 2928 4416
rect 2943 4406 2973 4422
rect 3001 4400 3007 4448
rect 3010 4442 3029 4448
rect 3044 4442 3074 4450
rect 3010 4434 3074 4442
rect 3010 4418 3090 4434
rect 3106 4427 3168 4458
rect 3184 4427 3246 4458
rect 3315 4456 3364 4481
rect 3379 4456 3409 4472
rect 3278 4442 3308 4450
rect 3315 4448 3425 4456
rect 3278 4434 3323 4442
rect 3010 4416 3029 4418
rect 3044 4416 3090 4418
rect 3010 4400 3090 4416
rect 3117 4414 3152 4427
rect 3193 4424 3230 4427
rect 3193 4422 3235 4424
rect 3122 4411 3152 4414
rect 3131 4407 3138 4411
rect 3138 4406 3139 4407
rect 3097 4400 3107 4406
rect 2856 4392 2891 4400
rect 2856 4366 2857 4392
rect 2864 4366 2891 4392
rect 2799 4348 2829 4362
rect 2856 4358 2891 4366
rect 2893 4392 2934 4400
rect 2893 4366 2908 4392
rect 2915 4366 2934 4392
rect 2998 4388 3029 4400
rect 3044 4388 3147 4400
rect 3159 4390 3185 4416
rect 3200 4411 3230 4422
rect 3262 4418 3324 4434
rect 3262 4416 3308 4418
rect 3262 4400 3324 4416
rect 3336 4400 3342 4448
rect 3345 4440 3425 4448
rect 3345 4438 3364 4440
rect 3379 4438 3413 4440
rect 3345 4422 3425 4438
rect 3345 4400 3364 4422
rect 3379 4406 3409 4422
rect 3437 4416 3443 4490
rect 3446 4416 3465 4560
rect 3480 4416 3486 4560
rect 3495 4490 3508 4560
rect 3560 4556 3582 4560
rect 3553 4534 3582 4548
rect 3635 4534 3651 4548
rect 3689 4544 3695 4546
rect 3702 4544 3810 4560
rect 3817 4544 3823 4546
rect 3831 4544 3846 4560
rect 3912 4554 3931 4557
rect 3553 4532 3651 4534
rect 3678 4532 3846 4544
rect 3861 4534 3877 4548
rect 3912 4535 3934 4554
rect 3944 4548 3960 4549
rect 3943 4546 3960 4548
rect 3944 4541 3960 4546
rect 3934 4534 3940 4535
rect 3943 4534 3972 4541
rect 3861 4533 3972 4534
rect 3861 4532 3978 4533
rect 3537 4524 3588 4532
rect 3635 4524 3669 4532
rect 3537 4512 3562 4524
rect 3569 4512 3588 4524
rect 3642 4522 3669 4524
rect 3678 4522 3899 4532
rect 3934 4529 3940 4532
rect 3642 4518 3899 4522
rect 3537 4504 3588 4512
rect 3635 4504 3899 4518
rect 3943 4524 3978 4532
rect 3489 4456 3508 4490
rect 3553 4496 3582 4504
rect 3553 4490 3570 4496
rect 3553 4488 3587 4490
rect 3635 4488 3651 4504
rect 3652 4494 3860 4504
rect 3861 4494 3877 4504
rect 3925 4500 3940 4515
rect 3943 4512 3944 4524
rect 3951 4512 3978 4524
rect 3943 4504 3978 4512
rect 3943 4503 3972 4504
rect 3663 4490 3877 4494
rect 3678 4488 3877 4490
rect 3912 4490 3925 4500
rect 3943 4490 3960 4503
rect 3912 4488 3960 4490
rect 3554 4484 3587 4488
rect 3550 4482 3587 4484
rect 3550 4481 3617 4482
rect 3550 4476 3581 4481
rect 3587 4476 3617 4481
rect 3550 4472 3617 4476
rect 3523 4469 3617 4472
rect 3523 4462 3572 4469
rect 3523 4456 3553 4462
rect 3572 4457 3577 4462
rect 3489 4440 3569 4456
rect 3581 4448 3617 4469
rect 3678 4464 3867 4488
rect 3912 4487 3959 4488
rect 3925 4482 3959 4487
rect 3693 4461 3867 4464
rect 3686 4458 3867 4461
rect 3895 4481 3959 4482
rect 3489 4438 3508 4440
rect 3523 4438 3557 4440
rect 3489 4422 3569 4438
rect 3489 4416 3508 4422
rect 3205 4390 3308 4400
rect 3159 4388 3308 4390
rect 3329 4388 3364 4400
rect 2998 4386 3160 4388
rect 3010 4366 3029 4386
rect 3044 4384 3074 4386
rect 2893 4358 2934 4366
rect 3016 4362 3029 4366
rect 3081 4370 3160 4386
rect 3192 4386 3364 4388
rect 3192 4370 3271 4386
rect 3278 4384 3308 4386
rect 2856 4348 2885 4358
rect 2899 4348 2928 4358
rect 2943 4348 2973 4362
rect 3016 4348 3059 4362
rect 3081 4358 3271 4370
rect 3336 4366 3342 4386
rect 3066 4348 3096 4358
rect 3097 4348 3255 4358
rect 3259 4348 3289 4358
rect 3293 4348 3323 4362
rect 3351 4348 3364 4386
rect 3436 4400 3465 4416
rect 3479 4400 3508 4416
rect 3523 4406 3553 4422
rect 3581 4400 3587 4448
rect 3590 4442 3609 4448
rect 3624 4442 3654 4450
rect 3590 4434 3654 4442
rect 3590 4418 3670 4434
rect 3686 4427 3748 4458
rect 3764 4427 3826 4458
rect 3895 4456 3944 4481
rect 3959 4456 3989 4472
rect 3858 4442 3888 4450
rect 3895 4448 4005 4456
rect 3858 4434 3903 4442
rect 3590 4416 3609 4418
rect 3624 4416 3670 4418
rect 3590 4400 3670 4416
rect 3697 4414 3732 4427
rect 3773 4424 3810 4427
rect 3773 4422 3815 4424
rect 3702 4411 3732 4414
rect 3711 4407 3718 4411
rect 3718 4406 3719 4407
rect 3677 4400 3687 4406
rect 3436 4392 3471 4400
rect 3436 4366 3437 4392
rect 3444 4366 3471 4392
rect 3379 4348 3409 4362
rect 3436 4358 3471 4366
rect 3473 4392 3514 4400
rect 3473 4366 3488 4392
rect 3495 4366 3514 4392
rect 3578 4388 3609 4400
rect 3624 4388 3727 4400
rect 3739 4390 3765 4416
rect 3780 4411 3810 4422
rect 3842 4418 3904 4434
rect 3842 4416 3888 4418
rect 3842 4400 3904 4416
rect 3916 4400 3922 4448
rect 3925 4440 4005 4448
rect 3925 4438 3944 4440
rect 3959 4438 3993 4440
rect 3925 4422 4005 4438
rect 3925 4400 3944 4422
rect 3959 4406 3989 4422
rect 4017 4416 4023 4490
rect 4026 4416 4045 4560
rect 4060 4416 4066 4560
rect 4075 4490 4088 4560
rect 4140 4556 4162 4560
rect 4133 4534 4162 4548
rect 4215 4534 4231 4548
rect 4269 4544 4275 4546
rect 4282 4544 4390 4560
rect 4397 4544 4403 4546
rect 4411 4544 4426 4560
rect 4492 4554 4511 4557
rect 4133 4532 4231 4534
rect 4258 4532 4426 4544
rect 4441 4534 4457 4548
rect 4492 4535 4514 4554
rect 4524 4548 4540 4549
rect 4523 4546 4540 4548
rect 4524 4541 4540 4546
rect 4514 4534 4520 4535
rect 4523 4534 4552 4541
rect 4441 4533 4552 4534
rect 4441 4532 4558 4533
rect 4117 4524 4168 4532
rect 4215 4524 4249 4532
rect 4117 4512 4142 4524
rect 4149 4512 4168 4524
rect 4222 4522 4249 4524
rect 4258 4522 4479 4532
rect 4514 4529 4520 4532
rect 4222 4518 4479 4522
rect 4117 4504 4168 4512
rect 4215 4504 4479 4518
rect 4523 4524 4558 4532
rect 4069 4456 4088 4490
rect 4133 4496 4162 4504
rect 4133 4490 4150 4496
rect 4133 4488 4167 4490
rect 4215 4488 4231 4504
rect 4232 4494 4440 4504
rect 4441 4494 4457 4504
rect 4505 4500 4520 4515
rect 4523 4512 4524 4524
rect 4531 4512 4558 4524
rect 4523 4504 4558 4512
rect 4523 4503 4552 4504
rect 4243 4490 4457 4494
rect 4258 4488 4457 4490
rect 4492 4490 4505 4500
rect 4523 4490 4540 4503
rect 4492 4488 4540 4490
rect 4134 4484 4167 4488
rect 4130 4482 4167 4484
rect 4130 4481 4197 4482
rect 4130 4476 4161 4481
rect 4167 4476 4197 4481
rect 4130 4472 4197 4476
rect 4103 4469 4197 4472
rect 4103 4462 4152 4469
rect 4103 4456 4133 4462
rect 4152 4457 4157 4462
rect 4069 4440 4149 4456
rect 4161 4448 4197 4469
rect 4258 4464 4447 4488
rect 4492 4487 4539 4488
rect 4505 4482 4539 4487
rect 4273 4461 4447 4464
rect 4266 4458 4447 4461
rect 4475 4481 4539 4482
rect 4069 4438 4088 4440
rect 4103 4438 4137 4440
rect 4069 4422 4149 4438
rect 4069 4416 4088 4422
rect 3785 4390 3888 4400
rect 3739 4388 3888 4390
rect 3909 4388 3944 4400
rect 3578 4386 3740 4388
rect 3590 4366 3609 4386
rect 3624 4384 3654 4386
rect 3473 4358 3514 4366
rect 3596 4362 3609 4366
rect 3661 4370 3740 4386
rect 3772 4386 3944 4388
rect 3772 4370 3851 4386
rect 3858 4384 3888 4386
rect 3436 4348 3465 4358
rect 3479 4348 3508 4358
rect 3523 4348 3553 4362
rect 3596 4348 3639 4362
rect 3661 4358 3851 4370
rect 3916 4366 3922 4386
rect 3646 4348 3676 4358
rect 3677 4348 3835 4358
rect 3839 4348 3869 4358
rect 3873 4348 3903 4362
rect 3931 4348 3944 4386
rect 4016 4400 4045 4416
rect 4059 4400 4088 4416
rect 4103 4406 4133 4422
rect 4161 4400 4167 4448
rect 4170 4442 4189 4448
rect 4204 4442 4234 4450
rect 4170 4434 4234 4442
rect 4170 4418 4250 4434
rect 4266 4427 4328 4458
rect 4344 4427 4406 4458
rect 4475 4456 4524 4481
rect 4539 4456 4569 4472
rect 4438 4442 4468 4450
rect 4475 4448 4585 4456
rect 4438 4434 4483 4442
rect 4170 4416 4189 4418
rect 4204 4416 4250 4418
rect 4170 4400 4250 4416
rect 4277 4414 4312 4427
rect 4353 4424 4390 4427
rect 4353 4422 4395 4424
rect 4282 4411 4312 4414
rect 4291 4407 4298 4411
rect 4298 4406 4299 4407
rect 4257 4400 4267 4406
rect 4016 4392 4051 4400
rect 4016 4366 4017 4392
rect 4024 4366 4051 4392
rect 3959 4348 3989 4362
rect 4016 4358 4051 4366
rect 4053 4392 4094 4400
rect 4053 4366 4068 4392
rect 4075 4366 4094 4392
rect 4158 4388 4189 4400
rect 4204 4388 4307 4400
rect 4319 4390 4345 4416
rect 4360 4411 4390 4422
rect 4422 4418 4484 4434
rect 4422 4416 4468 4418
rect 4422 4400 4484 4416
rect 4496 4400 4502 4448
rect 4505 4440 4585 4448
rect 4505 4438 4524 4440
rect 4539 4438 4573 4440
rect 4505 4422 4585 4438
rect 4505 4400 4524 4422
rect 4539 4406 4569 4422
rect 4597 4416 4603 4490
rect 4606 4416 4625 4560
rect 4640 4416 4646 4560
rect 4655 4490 4668 4560
rect 4720 4556 4742 4560
rect 4713 4534 4742 4548
rect 4795 4534 4811 4548
rect 4849 4544 4855 4546
rect 4862 4544 4970 4560
rect 4977 4544 4983 4546
rect 4991 4544 5006 4560
rect 5072 4554 5091 4557
rect 4713 4532 4811 4534
rect 4838 4532 5006 4544
rect 5021 4534 5037 4548
rect 5072 4535 5094 4554
rect 5104 4548 5120 4549
rect 5103 4546 5120 4548
rect 5104 4541 5120 4546
rect 5094 4534 5100 4535
rect 5103 4534 5132 4541
rect 5021 4533 5132 4534
rect 5021 4532 5138 4533
rect 4697 4524 4748 4532
rect 4795 4524 4829 4532
rect 4697 4512 4722 4524
rect 4729 4512 4748 4524
rect 4802 4522 4829 4524
rect 4838 4522 5059 4532
rect 5094 4529 5100 4532
rect 4802 4518 5059 4522
rect 4697 4504 4748 4512
rect 4795 4504 5059 4518
rect 5103 4524 5138 4532
rect 4649 4456 4668 4490
rect 4713 4496 4742 4504
rect 4713 4490 4730 4496
rect 4713 4488 4747 4490
rect 4795 4488 4811 4504
rect 4812 4494 5020 4504
rect 5021 4494 5037 4504
rect 5085 4500 5100 4515
rect 5103 4512 5104 4524
rect 5111 4512 5138 4524
rect 5103 4504 5138 4512
rect 5103 4503 5132 4504
rect 4823 4490 5037 4494
rect 4838 4488 5037 4490
rect 5072 4490 5085 4500
rect 5103 4490 5120 4503
rect 5072 4488 5120 4490
rect 4714 4484 4747 4488
rect 4710 4482 4747 4484
rect 4710 4481 4777 4482
rect 4710 4476 4741 4481
rect 4747 4476 4777 4481
rect 4710 4472 4777 4476
rect 4683 4469 4777 4472
rect 4683 4462 4732 4469
rect 4683 4456 4713 4462
rect 4732 4457 4737 4462
rect 4649 4440 4729 4456
rect 4741 4448 4777 4469
rect 4838 4464 5027 4488
rect 5072 4487 5119 4488
rect 5085 4482 5119 4487
rect 4853 4461 5027 4464
rect 4846 4458 5027 4461
rect 5055 4481 5119 4482
rect 4649 4438 4668 4440
rect 4683 4438 4717 4440
rect 4649 4422 4729 4438
rect 4649 4416 4668 4422
rect 4365 4390 4468 4400
rect 4319 4388 4468 4390
rect 4489 4388 4524 4400
rect 4158 4386 4320 4388
rect 4170 4366 4189 4386
rect 4204 4384 4234 4386
rect 4053 4358 4094 4366
rect 4176 4362 4189 4366
rect 4241 4370 4320 4386
rect 4352 4386 4524 4388
rect 4352 4370 4431 4386
rect 4438 4384 4468 4386
rect 4016 4348 4045 4358
rect 4059 4348 4088 4358
rect 4103 4348 4133 4362
rect 4176 4348 4219 4362
rect 4241 4358 4431 4370
rect 4496 4366 4502 4386
rect 4226 4348 4256 4358
rect 4257 4348 4415 4358
rect 4419 4348 4449 4358
rect 4453 4348 4483 4362
rect 4511 4348 4524 4386
rect 4596 4400 4625 4416
rect 4639 4400 4668 4416
rect 4683 4406 4713 4422
rect 4741 4400 4747 4448
rect 4750 4442 4769 4448
rect 4784 4442 4814 4450
rect 4750 4434 4814 4442
rect 4750 4418 4830 4434
rect 4846 4427 4908 4458
rect 4924 4427 4986 4458
rect 5055 4456 5104 4481
rect 5119 4456 5149 4472
rect 5018 4442 5048 4450
rect 5055 4448 5165 4456
rect 5018 4434 5063 4442
rect 4750 4416 4769 4418
rect 4784 4416 4830 4418
rect 4750 4400 4830 4416
rect 4857 4414 4892 4427
rect 4933 4424 4970 4427
rect 4933 4422 4975 4424
rect 4862 4411 4892 4414
rect 4871 4407 4878 4411
rect 4878 4406 4879 4407
rect 4837 4400 4847 4406
rect 4596 4392 4631 4400
rect 4596 4366 4597 4392
rect 4604 4366 4631 4392
rect 4539 4348 4569 4362
rect 4596 4358 4631 4366
rect 4633 4392 4674 4400
rect 4633 4366 4648 4392
rect 4655 4366 4674 4392
rect 4738 4388 4769 4400
rect 4784 4388 4887 4400
rect 4899 4390 4925 4416
rect 4940 4411 4970 4422
rect 5002 4418 5064 4434
rect 5002 4416 5048 4418
rect 5002 4400 5064 4416
rect 5076 4400 5082 4448
rect 5085 4440 5165 4448
rect 5085 4438 5104 4440
rect 5119 4438 5153 4440
rect 5085 4422 5165 4438
rect 5085 4400 5104 4422
rect 5119 4406 5149 4422
rect 5177 4416 5183 4490
rect 5186 4416 5205 4560
rect 5220 4416 5226 4560
rect 5235 4490 5248 4560
rect 5300 4556 5322 4560
rect 5293 4534 5322 4548
rect 5375 4534 5391 4548
rect 5429 4544 5435 4546
rect 5442 4544 5550 4560
rect 5557 4544 5563 4546
rect 5571 4544 5586 4560
rect 5652 4554 5671 4557
rect 5293 4532 5391 4534
rect 5418 4532 5586 4544
rect 5601 4534 5617 4548
rect 5652 4535 5674 4554
rect 5684 4548 5700 4549
rect 5683 4546 5700 4548
rect 5684 4541 5700 4546
rect 5674 4534 5680 4535
rect 5683 4534 5712 4541
rect 5601 4533 5712 4534
rect 5601 4532 5718 4533
rect 5277 4524 5328 4532
rect 5375 4524 5409 4532
rect 5277 4512 5302 4524
rect 5309 4512 5328 4524
rect 5382 4522 5409 4524
rect 5418 4522 5639 4532
rect 5674 4529 5680 4532
rect 5382 4518 5639 4522
rect 5277 4504 5328 4512
rect 5375 4504 5639 4518
rect 5683 4524 5718 4532
rect 5229 4456 5248 4490
rect 5293 4496 5322 4504
rect 5293 4490 5310 4496
rect 5293 4488 5327 4490
rect 5375 4488 5391 4504
rect 5392 4494 5600 4504
rect 5601 4494 5617 4504
rect 5665 4500 5680 4515
rect 5683 4512 5684 4524
rect 5691 4512 5718 4524
rect 5683 4504 5718 4512
rect 5683 4503 5712 4504
rect 5403 4490 5617 4494
rect 5418 4488 5617 4490
rect 5652 4490 5665 4500
rect 5683 4490 5700 4503
rect 5652 4488 5700 4490
rect 5294 4484 5327 4488
rect 5290 4482 5327 4484
rect 5290 4481 5357 4482
rect 5290 4476 5321 4481
rect 5327 4476 5357 4481
rect 5290 4472 5357 4476
rect 5263 4469 5357 4472
rect 5263 4462 5312 4469
rect 5263 4456 5293 4462
rect 5312 4457 5317 4462
rect 5229 4440 5309 4456
rect 5321 4448 5357 4469
rect 5418 4464 5607 4488
rect 5652 4487 5699 4488
rect 5665 4482 5699 4487
rect 5433 4461 5607 4464
rect 5426 4458 5607 4461
rect 5635 4481 5699 4482
rect 5229 4438 5248 4440
rect 5263 4438 5297 4440
rect 5229 4422 5309 4438
rect 5229 4416 5248 4422
rect 4945 4390 5048 4400
rect 4899 4388 5048 4390
rect 5069 4388 5104 4400
rect 4738 4386 4900 4388
rect 4750 4366 4769 4386
rect 4784 4384 4814 4386
rect 4633 4358 4674 4366
rect 4756 4362 4769 4366
rect 4821 4370 4900 4386
rect 4932 4386 5104 4388
rect 4932 4370 5011 4386
rect 5018 4384 5048 4386
rect 4596 4348 4625 4358
rect 4639 4348 4668 4358
rect 4683 4348 4713 4362
rect 4756 4348 4799 4362
rect 4821 4358 5011 4370
rect 5076 4366 5082 4386
rect 4806 4348 4836 4358
rect 4837 4348 4995 4358
rect 4999 4348 5029 4358
rect 5033 4348 5063 4362
rect 5091 4348 5104 4386
rect 5176 4400 5205 4416
rect 5219 4400 5248 4416
rect 5263 4406 5293 4422
rect 5321 4400 5327 4448
rect 5330 4442 5349 4448
rect 5364 4442 5394 4450
rect 5330 4434 5394 4442
rect 5330 4418 5410 4434
rect 5426 4427 5488 4458
rect 5504 4427 5566 4458
rect 5635 4456 5684 4481
rect 5699 4456 5729 4472
rect 5598 4442 5628 4450
rect 5635 4448 5745 4456
rect 5598 4434 5643 4442
rect 5330 4416 5349 4418
rect 5364 4416 5410 4418
rect 5330 4400 5410 4416
rect 5437 4414 5472 4427
rect 5513 4424 5550 4427
rect 5513 4422 5555 4424
rect 5442 4411 5472 4414
rect 5451 4407 5458 4411
rect 5458 4406 5459 4407
rect 5417 4400 5427 4406
rect 5176 4392 5211 4400
rect 5176 4366 5177 4392
rect 5184 4366 5211 4392
rect 5119 4348 5149 4362
rect 5176 4358 5211 4366
rect 5213 4392 5254 4400
rect 5213 4366 5228 4392
rect 5235 4366 5254 4392
rect 5318 4388 5349 4400
rect 5364 4388 5467 4400
rect 5479 4390 5505 4416
rect 5520 4411 5550 4422
rect 5582 4418 5644 4434
rect 5582 4416 5628 4418
rect 5582 4400 5644 4416
rect 5656 4400 5662 4448
rect 5665 4440 5745 4448
rect 5665 4438 5684 4440
rect 5699 4438 5733 4440
rect 5665 4422 5745 4438
rect 5665 4400 5684 4422
rect 5699 4406 5729 4422
rect 5757 4416 5763 4490
rect 5766 4416 5785 4560
rect 5800 4416 5806 4560
rect 5815 4490 5828 4560
rect 5880 4556 5902 4560
rect 5873 4534 5902 4548
rect 5955 4534 5971 4548
rect 6009 4544 6015 4546
rect 6022 4544 6130 4560
rect 6137 4544 6143 4546
rect 6151 4544 6166 4560
rect 6232 4554 6251 4557
rect 5873 4532 5971 4534
rect 5998 4532 6166 4544
rect 6181 4534 6197 4548
rect 6232 4535 6254 4554
rect 6264 4548 6280 4549
rect 6263 4546 6280 4548
rect 6264 4541 6280 4546
rect 6254 4534 6260 4535
rect 6263 4534 6292 4541
rect 6181 4533 6292 4534
rect 6181 4532 6298 4533
rect 5857 4524 5908 4532
rect 5955 4524 5989 4532
rect 5857 4512 5882 4524
rect 5889 4512 5908 4524
rect 5962 4522 5989 4524
rect 5998 4522 6219 4532
rect 6254 4529 6260 4532
rect 5962 4518 6219 4522
rect 5857 4504 5908 4512
rect 5955 4504 6219 4518
rect 6263 4524 6298 4532
rect 5809 4456 5828 4490
rect 5873 4496 5902 4504
rect 5873 4490 5890 4496
rect 5873 4488 5907 4490
rect 5955 4488 5971 4504
rect 5972 4494 6180 4504
rect 6181 4494 6197 4504
rect 6245 4500 6260 4515
rect 6263 4512 6264 4524
rect 6271 4512 6298 4524
rect 6263 4504 6298 4512
rect 6263 4503 6292 4504
rect 5983 4490 6197 4494
rect 5998 4488 6197 4490
rect 6232 4490 6245 4500
rect 6263 4490 6280 4503
rect 6232 4488 6280 4490
rect 5874 4484 5907 4488
rect 5870 4482 5907 4484
rect 5870 4481 5937 4482
rect 5870 4476 5901 4481
rect 5907 4476 5937 4481
rect 5870 4472 5937 4476
rect 5843 4469 5937 4472
rect 5843 4462 5892 4469
rect 5843 4456 5873 4462
rect 5892 4457 5897 4462
rect 5809 4440 5889 4456
rect 5901 4448 5937 4469
rect 5998 4464 6187 4488
rect 6232 4487 6279 4488
rect 6245 4482 6279 4487
rect 6013 4461 6187 4464
rect 6006 4458 6187 4461
rect 6215 4481 6279 4482
rect 5809 4438 5828 4440
rect 5843 4438 5877 4440
rect 5809 4422 5889 4438
rect 5809 4416 5828 4422
rect 5525 4390 5628 4400
rect 5479 4388 5628 4390
rect 5649 4388 5684 4400
rect 5318 4386 5480 4388
rect 5330 4366 5349 4386
rect 5364 4384 5394 4386
rect 5213 4358 5254 4366
rect 5336 4362 5349 4366
rect 5401 4370 5480 4386
rect 5512 4386 5684 4388
rect 5512 4370 5591 4386
rect 5598 4384 5628 4386
rect 5176 4348 5205 4358
rect 5219 4348 5248 4358
rect 5263 4348 5293 4362
rect 5336 4348 5379 4362
rect 5401 4358 5591 4370
rect 5656 4366 5662 4386
rect 5386 4348 5416 4358
rect 5417 4348 5575 4358
rect 5579 4348 5609 4358
rect 5613 4348 5643 4362
rect 5671 4348 5684 4386
rect 5756 4400 5785 4416
rect 5799 4400 5828 4416
rect 5843 4406 5873 4422
rect 5901 4400 5907 4448
rect 5910 4442 5929 4448
rect 5944 4442 5974 4450
rect 5910 4434 5974 4442
rect 5910 4418 5990 4434
rect 6006 4427 6068 4458
rect 6084 4427 6146 4458
rect 6215 4456 6264 4481
rect 6279 4456 6309 4472
rect 6178 4442 6208 4450
rect 6215 4448 6325 4456
rect 6178 4434 6223 4442
rect 5910 4416 5929 4418
rect 5944 4416 5990 4418
rect 5910 4400 5990 4416
rect 6017 4414 6052 4427
rect 6093 4424 6130 4427
rect 6093 4422 6135 4424
rect 6022 4411 6052 4414
rect 6031 4407 6038 4411
rect 6038 4406 6039 4407
rect 5997 4400 6007 4406
rect 5756 4392 5791 4400
rect 5756 4366 5757 4392
rect 5764 4366 5791 4392
rect 5699 4348 5729 4362
rect 5756 4358 5791 4366
rect 5793 4392 5834 4400
rect 5793 4366 5808 4392
rect 5815 4366 5834 4392
rect 5898 4388 5929 4400
rect 5944 4388 6047 4400
rect 6059 4390 6085 4416
rect 6100 4411 6130 4422
rect 6162 4418 6224 4434
rect 6162 4416 6208 4418
rect 6162 4400 6224 4416
rect 6236 4400 6242 4448
rect 6245 4440 6325 4448
rect 6245 4438 6264 4440
rect 6279 4438 6313 4440
rect 6245 4422 6325 4438
rect 6245 4400 6264 4422
rect 6279 4406 6309 4422
rect 6337 4416 6343 4490
rect 6346 4416 6365 4560
rect 6380 4416 6386 4560
rect 6395 4490 6408 4560
rect 6460 4556 6482 4560
rect 6453 4534 6482 4548
rect 6535 4534 6551 4548
rect 6589 4544 6595 4546
rect 6602 4544 6710 4560
rect 6717 4544 6723 4546
rect 6731 4544 6746 4560
rect 6812 4554 6831 4557
rect 6453 4532 6551 4534
rect 6578 4532 6746 4544
rect 6761 4534 6777 4548
rect 6812 4535 6834 4554
rect 6844 4548 6860 4549
rect 6843 4546 6860 4548
rect 6844 4541 6860 4546
rect 6834 4534 6840 4535
rect 6843 4534 6872 4541
rect 6761 4533 6872 4534
rect 6761 4532 6878 4533
rect 6437 4524 6488 4532
rect 6535 4524 6569 4532
rect 6437 4512 6462 4524
rect 6469 4512 6488 4524
rect 6542 4522 6569 4524
rect 6578 4522 6799 4532
rect 6834 4529 6840 4532
rect 6542 4518 6799 4522
rect 6437 4504 6488 4512
rect 6535 4504 6799 4518
rect 6843 4524 6878 4532
rect 6389 4456 6408 4490
rect 6453 4496 6482 4504
rect 6453 4490 6470 4496
rect 6453 4488 6487 4490
rect 6535 4488 6551 4504
rect 6552 4494 6760 4504
rect 6761 4494 6777 4504
rect 6825 4500 6840 4515
rect 6843 4512 6844 4524
rect 6851 4512 6878 4524
rect 6843 4504 6878 4512
rect 6843 4503 6872 4504
rect 6563 4490 6777 4494
rect 6578 4488 6777 4490
rect 6812 4490 6825 4500
rect 6843 4490 6860 4503
rect 6812 4488 6860 4490
rect 6454 4484 6487 4488
rect 6450 4482 6487 4484
rect 6450 4481 6517 4482
rect 6450 4476 6481 4481
rect 6487 4476 6517 4481
rect 6450 4472 6517 4476
rect 6423 4469 6517 4472
rect 6423 4462 6472 4469
rect 6423 4456 6453 4462
rect 6472 4457 6477 4462
rect 6389 4440 6469 4456
rect 6481 4448 6517 4469
rect 6578 4464 6767 4488
rect 6812 4487 6859 4488
rect 6825 4482 6859 4487
rect 6593 4461 6767 4464
rect 6586 4458 6767 4461
rect 6795 4481 6859 4482
rect 6389 4438 6408 4440
rect 6423 4438 6457 4440
rect 6389 4422 6469 4438
rect 6389 4416 6408 4422
rect 6105 4390 6208 4400
rect 6059 4388 6208 4390
rect 6229 4388 6264 4400
rect 5898 4386 6060 4388
rect 5910 4366 5929 4386
rect 5944 4384 5974 4386
rect 5793 4358 5834 4366
rect 5916 4362 5929 4366
rect 5981 4370 6060 4386
rect 6092 4386 6264 4388
rect 6092 4370 6171 4386
rect 6178 4384 6208 4386
rect 5756 4348 5785 4358
rect 5799 4348 5828 4358
rect 5843 4348 5873 4362
rect 5916 4348 5959 4362
rect 5981 4358 6171 4370
rect 6236 4366 6242 4386
rect 5966 4348 5996 4358
rect 5997 4348 6155 4358
rect 6159 4348 6189 4358
rect 6193 4348 6223 4362
rect 6251 4348 6264 4386
rect 6336 4400 6365 4416
rect 6379 4400 6408 4416
rect 6423 4406 6453 4422
rect 6481 4400 6487 4448
rect 6490 4442 6509 4448
rect 6524 4442 6554 4450
rect 6490 4434 6554 4442
rect 6490 4418 6570 4434
rect 6586 4427 6648 4458
rect 6664 4427 6726 4458
rect 6795 4456 6844 4481
rect 6859 4456 6889 4472
rect 6758 4442 6788 4450
rect 6795 4448 6905 4456
rect 6758 4434 6803 4442
rect 6490 4416 6509 4418
rect 6524 4416 6570 4418
rect 6490 4400 6570 4416
rect 6597 4414 6632 4427
rect 6673 4424 6710 4427
rect 6673 4422 6715 4424
rect 6602 4411 6632 4414
rect 6611 4407 6618 4411
rect 6618 4406 6619 4407
rect 6577 4400 6587 4406
rect 6336 4392 6371 4400
rect 6336 4366 6337 4392
rect 6344 4366 6371 4392
rect 6279 4348 6309 4362
rect 6336 4358 6371 4366
rect 6373 4392 6414 4400
rect 6373 4366 6388 4392
rect 6395 4366 6414 4392
rect 6478 4388 6509 4400
rect 6524 4388 6627 4400
rect 6639 4390 6665 4416
rect 6680 4411 6710 4422
rect 6742 4418 6804 4434
rect 6742 4416 6788 4418
rect 6742 4400 6804 4416
rect 6816 4400 6822 4448
rect 6825 4440 6905 4448
rect 6825 4438 6844 4440
rect 6859 4438 6893 4440
rect 6825 4422 6905 4438
rect 6825 4400 6844 4422
rect 6859 4406 6889 4422
rect 6917 4416 6923 4490
rect 6926 4416 6945 4560
rect 6960 4416 6966 4560
rect 6975 4490 6988 4560
rect 7040 4556 7062 4560
rect 7033 4534 7062 4548
rect 7115 4534 7131 4548
rect 7169 4544 7175 4546
rect 7182 4544 7290 4560
rect 7297 4544 7303 4546
rect 7311 4544 7326 4560
rect 7392 4554 7411 4557
rect 7033 4532 7131 4534
rect 7158 4532 7326 4544
rect 7341 4534 7357 4548
rect 7392 4535 7414 4554
rect 7424 4548 7440 4549
rect 7423 4546 7440 4548
rect 7424 4541 7440 4546
rect 7414 4534 7420 4535
rect 7423 4534 7452 4541
rect 7341 4533 7452 4534
rect 7341 4532 7458 4533
rect 7017 4524 7068 4532
rect 7115 4524 7149 4532
rect 7017 4512 7042 4524
rect 7049 4512 7068 4524
rect 7122 4522 7149 4524
rect 7158 4522 7379 4532
rect 7414 4529 7420 4532
rect 7122 4518 7379 4522
rect 7017 4504 7068 4512
rect 7115 4504 7379 4518
rect 7423 4524 7458 4532
rect 6969 4456 6988 4490
rect 7033 4496 7062 4504
rect 7033 4490 7050 4496
rect 7033 4488 7067 4490
rect 7115 4488 7131 4504
rect 7132 4494 7340 4504
rect 7341 4494 7357 4504
rect 7405 4500 7420 4515
rect 7423 4512 7424 4524
rect 7431 4512 7458 4524
rect 7423 4504 7458 4512
rect 7423 4503 7452 4504
rect 7143 4490 7357 4494
rect 7158 4488 7357 4490
rect 7392 4490 7405 4500
rect 7423 4490 7440 4503
rect 7392 4488 7440 4490
rect 7034 4484 7067 4488
rect 7030 4482 7067 4484
rect 7030 4481 7097 4482
rect 7030 4476 7061 4481
rect 7067 4476 7097 4481
rect 7030 4472 7097 4476
rect 7003 4469 7097 4472
rect 7003 4462 7052 4469
rect 7003 4456 7033 4462
rect 7052 4457 7057 4462
rect 6969 4440 7049 4456
rect 7061 4448 7097 4469
rect 7158 4464 7347 4488
rect 7392 4487 7439 4488
rect 7405 4482 7439 4487
rect 7173 4461 7347 4464
rect 7166 4458 7347 4461
rect 7375 4481 7439 4482
rect 6969 4438 6988 4440
rect 7003 4438 7037 4440
rect 6969 4422 7049 4438
rect 6969 4416 6988 4422
rect 6685 4390 6788 4400
rect 6639 4388 6788 4390
rect 6809 4388 6844 4400
rect 6478 4386 6640 4388
rect 6490 4366 6509 4386
rect 6524 4384 6554 4386
rect 6373 4358 6414 4366
rect 6496 4362 6509 4366
rect 6561 4370 6640 4386
rect 6672 4386 6844 4388
rect 6672 4370 6751 4386
rect 6758 4384 6788 4386
rect 6336 4348 6365 4358
rect 6379 4348 6408 4358
rect 6423 4348 6453 4362
rect 6496 4348 6539 4362
rect 6561 4358 6751 4370
rect 6816 4366 6822 4386
rect 6546 4348 6576 4358
rect 6577 4348 6735 4358
rect 6739 4348 6769 4358
rect 6773 4348 6803 4362
rect 6831 4348 6844 4386
rect 6916 4400 6945 4416
rect 6959 4400 6988 4416
rect 7003 4406 7033 4422
rect 7061 4400 7067 4448
rect 7070 4442 7089 4448
rect 7104 4442 7134 4450
rect 7070 4434 7134 4442
rect 7070 4418 7150 4434
rect 7166 4427 7228 4458
rect 7244 4427 7306 4458
rect 7375 4456 7424 4481
rect 7439 4456 7469 4472
rect 7338 4442 7368 4450
rect 7375 4448 7485 4456
rect 7338 4434 7383 4442
rect 7070 4416 7089 4418
rect 7104 4416 7150 4418
rect 7070 4400 7150 4416
rect 7177 4414 7212 4427
rect 7253 4424 7290 4427
rect 7253 4422 7295 4424
rect 7182 4411 7212 4414
rect 7191 4407 7198 4411
rect 7198 4406 7199 4407
rect 7157 4400 7167 4406
rect 6916 4392 6951 4400
rect 6916 4366 6917 4392
rect 6924 4366 6951 4392
rect 6859 4348 6889 4362
rect 6916 4358 6951 4366
rect 6953 4392 6994 4400
rect 6953 4366 6968 4392
rect 6975 4366 6994 4392
rect 7058 4388 7089 4400
rect 7104 4388 7207 4400
rect 7219 4390 7245 4416
rect 7260 4411 7290 4422
rect 7322 4418 7384 4434
rect 7322 4416 7368 4418
rect 7322 4400 7384 4416
rect 7396 4400 7402 4448
rect 7405 4440 7485 4448
rect 7405 4438 7424 4440
rect 7439 4438 7473 4440
rect 7405 4422 7485 4438
rect 7405 4400 7424 4422
rect 7439 4406 7469 4422
rect 7497 4416 7503 4490
rect 7506 4416 7525 4560
rect 7540 4416 7546 4560
rect 7555 4490 7568 4560
rect 7613 4538 7614 4548
rect 7629 4538 7642 4548
rect 7613 4534 7642 4538
rect 7647 4534 7677 4560
rect 7695 4546 7711 4548
rect 7783 4546 7836 4560
rect 7784 4544 7848 4546
rect 7891 4544 7906 4560
rect 7955 4557 7985 4560
rect 7955 4554 7991 4557
rect 7921 4546 7937 4548
rect 7695 4534 7710 4538
rect 7613 4532 7710 4534
rect 7738 4532 7906 4544
rect 7922 4534 7937 4538
rect 7955 4535 7994 4554
rect 8013 4548 8020 4549
rect 8019 4541 8020 4548
rect 8003 4538 8004 4541
rect 8019 4538 8032 4541
rect 7955 4534 7985 4535
rect 7994 4534 8000 4535
rect 8003 4534 8032 4538
rect 7922 4533 8032 4534
rect 7922 4532 8038 4533
rect 7597 4524 7648 4532
rect 7597 4512 7622 4524
rect 7629 4512 7648 4524
rect 7679 4524 7729 4532
rect 7679 4516 7695 4524
rect 7702 4522 7729 4524
rect 7738 4522 7959 4532
rect 7702 4512 7959 4522
rect 7988 4524 8038 4532
rect 7988 4515 8004 4524
rect 7597 4504 7648 4512
rect 7695 4504 7959 4512
rect 7985 4512 8004 4515
rect 8011 4512 8038 4524
rect 7985 4504 8038 4512
rect 7549 4456 7568 4490
rect 7613 4496 7614 4504
rect 7629 4496 7642 4504
rect 7613 4488 7629 4496
rect 7610 4481 7629 4484
rect 7610 4472 7632 4481
rect 7583 4462 7632 4472
rect 7583 4456 7613 4462
rect 7632 4457 7637 4462
rect 7549 4440 7629 4456
rect 7647 4448 7677 4504
rect 7712 4494 7920 4504
rect 7955 4500 8000 4504
rect 8003 4503 8004 4504
rect 8019 4503 8032 4504
rect 7738 4464 7927 4494
rect 7753 4461 7927 4464
rect 7746 4458 7927 4461
rect 7549 4438 7568 4440
rect 7583 4438 7617 4440
rect 7549 4422 7629 4438
rect 7656 4434 7669 4448
rect 7684 4434 7700 4450
rect 7746 4445 7757 4458
rect 7549 4416 7568 4422
rect 7265 4390 7368 4400
rect 7219 4388 7368 4390
rect 7389 4388 7424 4400
rect 7058 4386 7220 4388
rect 7070 4366 7089 4386
rect 7104 4384 7134 4386
rect 6953 4358 6994 4366
rect 7076 4362 7089 4366
rect 7141 4370 7220 4386
rect 7252 4386 7424 4388
rect 7252 4370 7331 4386
rect 7338 4384 7368 4386
rect 6916 4348 6945 4358
rect 6959 4348 6988 4358
rect 7003 4348 7033 4362
rect 7076 4348 7119 4362
rect 7141 4358 7331 4370
rect 7396 4366 7402 4386
rect 7126 4348 7156 4358
rect 7157 4348 7315 4358
rect 7319 4348 7349 4358
rect 7353 4348 7383 4362
rect 7411 4348 7424 4386
rect 7496 4400 7525 4416
rect 7539 4400 7568 4416
rect 7583 4400 7613 4422
rect 7656 4418 7718 4434
rect 7746 4427 7757 4443
rect 7762 4438 7772 4458
rect 7782 4438 7796 4458
rect 7799 4445 7808 4458
rect 7824 4445 7833 4458
rect 7762 4427 7796 4438
rect 7799 4427 7808 4443
rect 7824 4427 7833 4443
rect 7840 4438 7850 4458
rect 7860 4438 7874 4458
rect 7875 4445 7886 4458
rect 7840 4427 7874 4438
rect 7875 4427 7886 4443
rect 7932 4434 7948 4450
rect 7955 4448 7985 4500
rect 8019 4496 8020 4503
rect 8004 4488 8020 4496
rect 7991 4456 8004 4475
rect 8019 4456 8049 4472
rect 7991 4440 8065 4456
rect 7991 4438 8004 4440
rect 8019 4438 8053 4440
rect 7656 4416 7669 4418
rect 7684 4416 7718 4418
rect 7656 4400 7718 4416
rect 7762 4411 7778 4414
rect 7840 4411 7870 4422
rect 7918 4418 7964 4434
rect 7991 4422 8065 4438
rect 7918 4416 7952 4418
rect 7917 4400 7964 4416
rect 7991 4400 8004 4422
rect 8019 4400 8049 4422
rect 8076 4400 8077 4416
rect 8092 4400 8105 4560
rect 8135 4456 8148 4560
rect 8193 4538 8194 4548
rect 8209 4538 8222 4548
rect 8193 4534 8222 4538
rect 8227 4534 8257 4560
rect 8275 4546 8291 4548
rect 8363 4546 8416 4560
rect 8364 4544 8428 4546
rect 8471 4544 8486 4560
rect 8535 4557 8565 4560
rect 8535 4554 8571 4557
rect 8501 4546 8517 4548
rect 8275 4534 8290 4538
rect 8193 4532 8290 4534
rect 8318 4532 8486 4544
rect 8502 4534 8517 4538
rect 8535 4535 8574 4554
rect 8593 4548 8600 4549
rect 8599 4541 8600 4548
rect 8583 4538 8584 4541
rect 8599 4538 8612 4541
rect 8535 4534 8565 4535
rect 8574 4534 8580 4535
rect 8583 4534 8612 4538
rect 8502 4533 8612 4534
rect 8502 4532 8618 4533
rect 8177 4524 8228 4532
rect 8177 4512 8202 4524
rect 8209 4512 8228 4524
rect 8259 4524 8309 4532
rect 8259 4516 8275 4524
rect 8282 4522 8309 4524
rect 8318 4522 8539 4532
rect 8282 4512 8539 4522
rect 8568 4524 8618 4532
rect 8568 4515 8584 4524
rect 8177 4504 8228 4512
rect 8275 4504 8539 4512
rect 8565 4512 8584 4515
rect 8591 4512 8618 4524
rect 8565 4504 8618 4512
rect 8193 4496 8194 4504
rect 8209 4496 8222 4504
rect 8193 4488 8209 4496
rect 8190 4481 8209 4484
rect 8190 4472 8212 4481
rect 8163 4462 8212 4472
rect 8163 4456 8193 4462
rect 8212 4457 8217 4462
rect 8135 4440 8209 4456
rect 8227 4448 8257 4504
rect 8292 4494 8500 4504
rect 8535 4500 8580 4504
rect 8583 4503 8584 4504
rect 8599 4503 8612 4504
rect 8318 4464 8507 4494
rect 8333 4461 8507 4464
rect 8326 4458 8507 4461
rect 8135 4438 8148 4440
rect 8163 4438 8197 4440
rect 8135 4422 8209 4438
rect 8236 4434 8249 4448
rect 8264 4434 8280 4450
rect 8326 4445 8337 4458
rect 8119 4400 8120 4416
rect 8135 4400 8148 4422
rect 8163 4400 8193 4422
rect 8236 4418 8298 4434
rect 8326 4427 8337 4443
rect 8342 4438 8352 4458
rect 8362 4438 8376 4458
rect 8379 4445 8388 4458
rect 8404 4445 8413 4458
rect 8342 4427 8376 4438
rect 8379 4427 8388 4443
rect 8404 4427 8413 4443
rect 8420 4438 8430 4458
rect 8440 4438 8454 4458
rect 8455 4445 8466 4458
rect 8420 4427 8454 4438
rect 8455 4427 8466 4443
rect 8512 4434 8528 4450
rect 8535 4448 8565 4500
rect 8599 4496 8600 4503
rect 8584 4488 8600 4496
rect 8571 4456 8584 4475
rect 8599 4456 8629 4472
rect 8571 4440 8645 4456
rect 8571 4438 8584 4440
rect 8599 4438 8633 4440
rect 8236 4416 8249 4418
rect 8264 4416 8298 4418
rect 8236 4400 8298 4416
rect 8342 4411 8358 4414
rect 8420 4411 8450 4422
rect 8498 4418 8544 4434
rect 8571 4422 8645 4438
rect 8498 4416 8532 4418
rect 8497 4400 8544 4416
rect 8571 4400 8584 4422
rect 8599 4400 8629 4422
rect 8656 4400 8657 4416
rect 8672 4400 8685 4560
rect 8715 4456 8728 4560
rect 8773 4538 8774 4548
rect 8789 4538 8802 4548
rect 8773 4534 8802 4538
rect 8807 4534 8837 4560
rect 8855 4546 8871 4548
rect 8943 4546 8996 4560
rect 8944 4544 9008 4546
rect 9051 4544 9066 4560
rect 9115 4557 9145 4560
rect 9115 4554 9151 4557
rect 9081 4546 9097 4548
rect 8855 4534 8870 4538
rect 8773 4532 8870 4534
rect 8898 4532 9066 4544
rect 9082 4534 9097 4538
rect 9115 4535 9154 4554
rect 9173 4548 9180 4549
rect 9179 4541 9180 4548
rect 9163 4538 9164 4541
rect 9179 4538 9192 4541
rect 9115 4534 9145 4535
rect 9154 4534 9160 4535
rect 9163 4534 9192 4538
rect 9082 4533 9192 4534
rect 9082 4532 9198 4533
rect 8757 4524 8808 4532
rect 8757 4512 8782 4524
rect 8789 4512 8808 4524
rect 8839 4524 8889 4532
rect 8839 4516 8855 4524
rect 8862 4522 8889 4524
rect 8898 4522 9119 4532
rect 8862 4512 9119 4522
rect 9148 4524 9198 4532
rect 9148 4515 9164 4524
rect 8757 4504 8808 4512
rect 8855 4504 9119 4512
rect 9145 4512 9164 4515
rect 9171 4512 9198 4524
rect 9145 4504 9198 4512
rect 8773 4496 8774 4504
rect 8789 4496 8802 4504
rect 8773 4488 8789 4496
rect 8770 4481 8789 4484
rect 8770 4472 8792 4481
rect 8743 4462 8792 4472
rect 8743 4456 8773 4462
rect 8792 4457 8797 4462
rect 8715 4440 8789 4456
rect 8807 4448 8837 4504
rect 8872 4494 9080 4504
rect 9115 4500 9160 4504
rect 9163 4503 9164 4504
rect 9179 4503 9192 4504
rect 8898 4464 9087 4494
rect 8913 4461 9087 4464
rect 8906 4458 9087 4461
rect 8715 4438 8728 4440
rect 8743 4438 8777 4440
rect 8715 4422 8789 4438
rect 8816 4434 8829 4448
rect 8844 4434 8860 4450
rect 8906 4445 8917 4458
rect 8699 4400 8700 4416
rect 8715 4400 8728 4422
rect 8743 4400 8773 4422
rect 8816 4418 8878 4434
rect 8906 4427 8917 4443
rect 8922 4438 8932 4458
rect 8942 4438 8956 4458
rect 8959 4445 8968 4458
rect 8984 4445 8993 4458
rect 8922 4427 8956 4438
rect 8959 4427 8968 4443
rect 8984 4427 8993 4443
rect 9000 4438 9010 4458
rect 9020 4438 9034 4458
rect 9035 4445 9046 4458
rect 9000 4427 9034 4438
rect 9035 4427 9046 4443
rect 9092 4434 9108 4450
rect 9115 4448 9145 4500
rect 9179 4496 9180 4503
rect 9164 4488 9180 4496
rect 9151 4456 9164 4475
rect 9179 4456 9209 4472
rect 9151 4440 9225 4456
rect 9151 4438 9164 4440
rect 9179 4438 9213 4440
rect 8816 4416 8829 4418
rect 8844 4416 8878 4418
rect 8816 4400 8878 4416
rect 8922 4411 8938 4414
rect 9000 4411 9030 4422
rect 9078 4418 9124 4434
rect 9151 4422 9225 4438
rect 9078 4416 9112 4418
rect 9077 4400 9124 4416
rect 9151 4400 9164 4422
rect 9179 4400 9209 4422
rect 9236 4400 9237 4416
rect 9252 4400 9265 4560
rect 7496 4392 7531 4400
rect 7496 4366 7497 4392
rect 7504 4366 7531 4392
rect 7439 4348 7469 4362
rect 7496 4358 7531 4366
rect 7533 4392 7574 4400
rect 7533 4366 7548 4392
rect 7555 4366 7574 4392
rect 7638 4388 7700 4400
rect 7712 4388 7787 4400
rect 7845 4388 7920 4400
rect 7932 4388 7963 4400
rect 7969 4388 8004 4400
rect 7638 4386 7800 4388
rect 7533 4358 7574 4366
rect 7656 4362 7669 4386
rect 7684 4384 7699 4386
rect 7496 4348 7525 4358
rect 7539 4348 7568 4358
rect 7583 4348 7613 4362
rect 7656 4348 7699 4362
rect 7723 4359 7730 4366
rect 7733 4362 7800 4386
rect 7832 4386 8004 4388
rect 7802 4364 7830 4368
rect 7832 4364 7912 4386
rect 7933 4384 7948 4386
rect 7802 4362 7912 4364
rect 7733 4358 7912 4362
rect 7706 4348 7736 4358
rect 7738 4348 7891 4358
rect 7899 4348 7929 4358
rect 7933 4348 7963 4362
rect 7991 4348 8004 4386
rect 8076 4392 8111 4400
rect 8076 4366 8077 4392
rect 8084 4366 8111 4392
rect 8019 4348 8049 4362
rect 8076 4358 8111 4366
rect 8113 4392 8154 4400
rect 8113 4366 8128 4392
rect 8135 4366 8154 4392
rect 8218 4388 8280 4400
rect 8292 4388 8367 4400
rect 8425 4388 8500 4400
rect 8512 4388 8543 4400
rect 8549 4388 8584 4400
rect 8218 4386 8380 4388
rect 8113 4358 8154 4366
rect 8236 4362 8249 4386
rect 8264 4384 8279 4386
rect 8076 4348 8077 4358
rect 8092 4348 8105 4358
rect 8119 4348 8120 4358
rect 8135 4348 8148 4358
rect 8163 4348 8193 4362
rect 8236 4348 8279 4362
rect 8303 4359 8310 4366
rect 8313 4362 8380 4386
rect 8412 4386 8584 4388
rect 8382 4364 8410 4368
rect 8412 4364 8492 4386
rect 8513 4384 8528 4386
rect 8382 4362 8492 4364
rect 8313 4358 8492 4362
rect 8286 4348 8316 4358
rect 8318 4348 8471 4358
rect 8479 4348 8509 4358
rect 8513 4348 8543 4362
rect 8571 4348 8584 4386
rect 8656 4392 8691 4400
rect 8656 4366 8657 4392
rect 8664 4366 8691 4392
rect 8599 4348 8629 4362
rect 8656 4358 8691 4366
rect 8693 4392 8734 4400
rect 8693 4366 8708 4392
rect 8715 4366 8734 4392
rect 8798 4388 8860 4400
rect 8872 4388 8947 4400
rect 9005 4388 9080 4400
rect 9092 4388 9123 4400
rect 9129 4388 9164 4400
rect 8798 4386 8960 4388
rect 8693 4358 8734 4366
rect 8816 4362 8829 4386
rect 8844 4384 8859 4386
rect 8656 4348 8657 4358
rect 8672 4348 8685 4358
rect 8699 4348 8700 4358
rect 8715 4348 8728 4358
rect 8743 4348 8773 4362
rect 8816 4348 8859 4362
rect 8883 4359 8890 4366
rect 8893 4362 8960 4386
rect 8992 4386 9164 4388
rect 8962 4364 8990 4368
rect 8992 4364 9072 4386
rect 9093 4384 9108 4386
rect 8962 4362 9072 4364
rect 8893 4358 9072 4362
rect 8866 4348 8896 4358
rect 8898 4348 9051 4358
rect 9059 4348 9089 4358
rect 9093 4348 9123 4362
rect 9151 4348 9164 4386
rect 9236 4392 9271 4400
rect 9236 4366 9237 4392
rect 9244 4366 9271 4392
rect 9179 4348 9209 4362
rect 9236 4358 9271 4366
rect 9236 4348 9237 4358
rect 9252 4348 9265 4358
rect -1 4342 9265 4348
rect 0 4334 9265 4342
rect 15 4304 28 4334
rect 43 4320 73 4334
rect 116 4320 159 4334
rect 166 4320 386 4334
rect 393 4320 423 4334
rect 83 4306 98 4318
rect 117 4306 130 4320
rect 198 4316 351 4320
rect 80 4304 102 4306
rect 180 4304 372 4316
rect 451 4304 464 4334
rect 479 4320 509 4334
rect 546 4304 565 4334
rect 580 4304 586 4334
rect 595 4304 608 4334
rect 623 4320 653 4334
rect 696 4320 739 4334
rect 746 4320 966 4334
rect 973 4320 1003 4334
rect 663 4306 678 4318
rect 697 4306 710 4320
rect 778 4316 931 4320
rect 660 4304 682 4306
rect 760 4304 952 4316
rect 1031 4304 1044 4334
rect 1059 4320 1089 4334
rect 1126 4304 1145 4334
rect 1160 4304 1166 4334
rect 1175 4304 1188 4334
rect 1203 4320 1233 4334
rect 1276 4320 1319 4334
rect 1326 4320 1546 4334
rect 1553 4320 1583 4334
rect 1243 4306 1258 4318
rect 1277 4306 1290 4320
rect 1358 4316 1511 4320
rect 1240 4304 1262 4306
rect 1340 4304 1532 4316
rect 1611 4304 1624 4334
rect 1639 4320 1669 4334
rect 1706 4304 1725 4334
rect 1740 4304 1746 4334
rect 1755 4304 1768 4334
rect 1783 4320 1813 4334
rect 1856 4320 1899 4334
rect 1906 4320 2126 4334
rect 2133 4320 2163 4334
rect 1823 4306 1838 4318
rect 1857 4306 1870 4320
rect 1938 4316 2091 4320
rect 1820 4304 1842 4306
rect 1920 4304 2112 4316
rect 2191 4304 2204 4334
rect 2219 4320 2249 4334
rect 2286 4304 2305 4334
rect 2320 4304 2326 4334
rect 2335 4304 2348 4334
rect 2363 4320 2393 4334
rect 2436 4320 2479 4334
rect 2486 4320 2706 4334
rect 2713 4320 2743 4334
rect 2403 4306 2418 4318
rect 2437 4306 2450 4320
rect 2518 4316 2671 4320
rect 2400 4304 2422 4306
rect 2500 4304 2692 4316
rect 2771 4304 2784 4334
rect 2799 4320 2829 4334
rect 2866 4304 2885 4334
rect 2900 4304 2906 4334
rect 2915 4304 2928 4334
rect 2943 4320 2973 4334
rect 3016 4320 3059 4334
rect 3066 4320 3286 4334
rect 3293 4320 3323 4334
rect 2983 4306 2998 4318
rect 3017 4306 3030 4320
rect 3098 4316 3251 4320
rect 2980 4304 3002 4306
rect 3080 4304 3272 4316
rect 3351 4304 3364 4334
rect 3379 4320 3409 4334
rect 3446 4304 3465 4334
rect 3480 4304 3486 4334
rect 3495 4304 3508 4334
rect 3523 4320 3553 4334
rect 3596 4320 3639 4334
rect 3646 4320 3866 4334
rect 3873 4320 3903 4334
rect 3563 4306 3578 4318
rect 3597 4306 3610 4320
rect 3678 4316 3831 4320
rect 3560 4304 3582 4306
rect 3660 4304 3852 4316
rect 3931 4304 3944 4334
rect 3959 4320 3989 4334
rect 4026 4304 4045 4334
rect 4060 4304 4066 4334
rect 4075 4304 4088 4334
rect 4103 4320 4133 4334
rect 4176 4320 4219 4334
rect 4226 4320 4446 4334
rect 4453 4320 4483 4334
rect 4143 4306 4158 4318
rect 4177 4306 4190 4320
rect 4258 4316 4411 4320
rect 4140 4304 4162 4306
rect 4240 4304 4432 4316
rect 4511 4304 4524 4334
rect 4539 4320 4569 4334
rect 4606 4304 4625 4334
rect 4640 4304 4646 4334
rect 4655 4304 4668 4334
rect 4683 4320 4713 4334
rect 4756 4320 4799 4334
rect 4806 4320 5026 4334
rect 5033 4320 5063 4334
rect 4723 4306 4738 4318
rect 4757 4306 4770 4320
rect 4838 4316 4991 4320
rect 4720 4304 4742 4306
rect 4820 4304 5012 4316
rect 5091 4304 5104 4334
rect 5119 4320 5149 4334
rect 5186 4304 5205 4334
rect 5220 4304 5226 4334
rect 5235 4304 5248 4334
rect 5263 4320 5293 4334
rect 5336 4320 5379 4334
rect 5386 4320 5606 4334
rect 5613 4320 5643 4334
rect 5303 4306 5318 4318
rect 5337 4306 5350 4320
rect 5418 4316 5571 4320
rect 5300 4304 5322 4306
rect 5400 4304 5592 4316
rect 5671 4304 5684 4334
rect 5699 4320 5729 4334
rect 5766 4304 5785 4334
rect 5800 4304 5806 4334
rect 5815 4304 5828 4334
rect 5843 4320 5873 4334
rect 5916 4320 5959 4334
rect 5966 4320 6186 4334
rect 6193 4320 6223 4334
rect 5883 4306 5898 4318
rect 5917 4306 5930 4320
rect 5998 4316 6151 4320
rect 5880 4304 5902 4306
rect 5980 4304 6172 4316
rect 6251 4304 6264 4334
rect 6279 4320 6309 4334
rect 6346 4304 6365 4334
rect 6380 4304 6386 4334
rect 6395 4304 6408 4334
rect 6423 4320 6453 4334
rect 6496 4320 6539 4334
rect 6546 4320 6766 4334
rect 6773 4320 6803 4334
rect 6463 4306 6478 4318
rect 6497 4306 6510 4320
rect 6578 4316 6731 4320
rect 6460 4304 6482 4306
rect 6560 4304 6752 4316
rect 6831 4304 6844 4334
rect 6859 4320 6889 4334
rect 6926 4304 6945 4334
rect 6960 4304 6966 4334
rect 6975 4304 6988 4334
rect 7003 4320 7033 4334
rect 7076 4320 7119 4334
rect 7126 4320 7346 4334
rect 7353 4320 7383 4334
rect 7043 4306 7058 4318
rect 7077 4306 7090 4320
rect 7158 4316 7311 4320
rect 7040 4304 7062 4306
rect 7140 4304 7332 4316
rect 7411 4304 7424 4334
rect 7439 4320 7469 4334
rect 7506 4304 7525 4334
rect 7540 4304 7546 4334
rect 7555 4304 7568 4334
rect 7583 4316 7613 4334
rect 7656 4320 7670 4334
rect 7706 4320 7926 4334
rect 7657 4318 7670 4320
rect 7623 4306 7638 4318
rect 7620 4304 7642 4306
rect 7647 4304 7677 4318
rect 7738 4316 7891 4320
rect 7720 4304 7912 4316
rect 7955 4304 7985 4318
rect 7991 4304 8004 4334
rect 8019 4316 8049 4334
rect 8092 4304 8105 4334
rect 8135 4304 8148 4334
rect 8163 4316 8193 4334
rect 8236 4320 8250 4334
rect 8286 4320 8506 4334
rect 8237 4318 8250 4320
rect 8203 4306 8218 4318
rect 8200 4304 8222 4306
rect 8227 4304 8257 4318
rect 8318 4316 8471 4320
rect 8300 4304 8492 4316
rect 8535 4304 8565 4318
rect 8571 4304 8584 4334
rect 8599 4316 8629 4334
rect 8672 4304 8685 4334
rect 8715 4304 8728 4334
rect 8743 4316 8773 4334
rect 8816 4320 8830 4334
rect 8866 4320 9086 4334
rect 8817 4318 8830 4320
rect 8783 4306 8798 4318
rect 8780 4304 8802 4306
rect 8807 4304 8837 4318
rect 8898 4316 9051 4320
rect 8880 4304 9072 4316
rect 9115 4304 9145 4318
rect 9151 4304 9164 4334
rect 9179 4316 9209 4334
rect 9252 4304 9265 4334
rect 0 4290 9265 4304
rect 15 4220 28 4290
rect 80 4286 102 4290
rect 73 4264 102 4278
rect 155 4264 171 4278
rect 209 4274 215 4276
rect 222 4274 330 4290
rect 337 4274 343 4276
rect 351 4274 366 4290
rect 432 4284 451 4287
rect 73 4262 171 4264
rect 198 4262 366 4274
rect 381 4264 397 4278
rect 432 4265 454 4284
rect 464 4278 480 4279
rect 463 4276 480 4278
rect 464 4271 480 4276
rect 454 4264 460 4265
rect 463 4264 492 4271
rect 381 4263 492 4264
rect 381 4262 498 4263
rect 57 4254 108 4262
rect 155 4254 189 4262
rect 57 4242 82 4254
rect 89 4242 108 4254
rect 162 4252 189 4254
rect 198 4252 419 4262
rect 454 4259 460 4262
rect 162 4248 419 4252
rect 57 4234 108 4242
rect 155 4234 419 4248
rect 463 4254 498 4262
rect 9 4186 28 4220
rect 73 4226 102 4234
rect 73 4220 90 4226
rect 73 4218 107 4220
rect 155 4218 171 4234
rect 172 4224 380 4234
rect 381 4224 397 4234
rect 445 4230 460 4245
rect 463 4242 464 4254
rect 471 4242 498 4254
rect 463 4234 498 4242
rect 463 4233 492 4234
rect 183 4220 397 4224
rect 198 4218 397 4220
rect 432 4220 445 4230
rect 463 4220 480 4233
rect 432 4218 480 4220
rect 74 4214 107 4218
rect 70 4212 107 4214
rect 70 4211 137 4212
rect 70 4206 101 4211
rect 107 4206 137 4211
rect 70 4202 137 4206
rect 43 4199 137 4202
rect 43 4192 92 4199
rect 43 4186 73 4192
rect 92 4187 97 4192
rect 9 4170 89 4186
rect 101 4178 137 4199
rect 198 4194 387 4218
rect 432 4217 479 4218
rect 445 4212 479 4217
rect 213 4191 387 4194
rect 206 4188 387 4191
rect 415 4211 479 4212
rect 9 4168 28 4170
rect 43 4168 77 4170
rect 9 4152 89 4168
rect 9 4146 28 4152
rect -1 4130 28 4146
rect 43 4136 73 4152
rect 101 4130 107 4178
rect 110 4172 129 4178
rect 144 4172 174 4180
rect 110 4164 174 4172
rect 110 4148 190 4164
rect 206 4157 268 4188
rect 284 4157 346 4188
rect 415 4186 464 4211
rect 479 4186 509 4202
rect 378 4172 408 4180
rect 415 4178 525 4186
rect 378 4164 423 4172
rect 110 4146 129 4148
rect 144 4146 190 4148
rect 110 4130 190 4146
rect 217 4144 252 4157
rect 293 4154 330 4157
rect 293 4152 335 4154
rect 222 4141 252 4144
rect 231 4137 238 4141
rect 238 4136 239 4137
rect 197 4130 207 4136
rect -7 4122 34 4130
rect -7 4096 8 4122
rect 15 4096 34 4122
rect 98 4118 129 4130
rect 144 4118 247 4130
rect 259 4120 285 4146
rect 300 4141 330 4152
rect 362 4148 424 4164
rect 362 4146 408 4148
rect 362 4130 424 4146
rect 436 4130 442 4178
rect 445 4170 525 4178
rect 445 4168 464 4170
rect 479 4168 513 4170
rect 445 4152 525 4168
rect 445 4130 464 4152
rect 479 4136 509 4152
rect 537 4146 543 4220
rect 546 4146 565 4290
rect 580 4146 586 4290
rect 595 4220 608 4290
rect 660 4286 682 4290
rect 653 4264 682 4278
rect 735 4264 751 4278
rect 789 4274 795 4276
rect 802 4274 910 4290
rect 917 4274 923 4276
rect 931 4274 946 4290
rect 1012 4284 1031 4287
rect 653 4262 751 4264
rect 778 4262 946 4274
rect 961 4264 977 4278
rect 1012 4265 1034 4284
rect 1044 4278 1060 4279
rect 1043 4276 1060 4278
rect 1044 4271 1060 4276
rect 1034 4264 1040 4265
rect 1043 4264 1072 4271
rect 961 4263 1072 4264
rect 961 4262 1078 4263
rect 637 4254 688 4262
rect 735 4254 769 4262
rect 637 4242 662 4254
rect 669 4242 688 4254
rect 742 4252 769 4254
rect 778 4252 999 4262
rect 1034 4259 1040 4262
rect 742 4248 999 4252
rect 637 4234 688 4242
rect 735 4234 999 4248
rect 1043 4254 1078 4262
rect 589 4186 608 4220
rect 653 4226 682 4234
rect 653 4220 670 4226
rect 653 4218 687 4220
rect 735 4218 751 4234
rect 752 4224 960 4234
rect 961 4224 977 4234
rect 1025 4230 1040 4245
rect 1043 4242 1044 4254
rect 1051 4242 1078 4254
rect 1043 4234 1078 4242
rect 1043 4233 1072 4234
rect 763 4220 977 4224
rect 778 4218 977 4220
rect 1012 4220 1025 4230
rect 1043 4220 1060 4233
rect 1012 4218 1060 4220
rect 654 4214 687 4218
rect 650 4212 687 4214
rect 650 4211 717 4212
rect 650 4206 681 4211
rect 687 4206 717 4211
rect 650 4202 717 4206
rect 623 4199 717 4202
rect 623 4192 672 4199
rect 623 4186 653 4192
rect 672 4187 677 4192
rect 589 4170 669 4186
rect 681 4178 717 4199
rect 778 4194 967 4218
rect 1012 4217 1059 4218
rect 1025 4212 1059 4217
rect 793 4191 967 4194
rect 786 4188 967 4191
rect 995 4211 1059 4212
rect 589 4168 608 4170
rect 623 4168 657 4170
rect 589 4152 669 4168
rect 589 4146 608 4152
rect 305 4120 408 4130
rect 259 4118 408 4120
rect 429 4118 464 4130
rect 98 4116 260 4118
rect 110 4096 129 4116
rect 144 4114 174 4116
rect -7 4088 34 4096
rect 116 4092 129 4096
rect 181 4100 260 4116
rect 292 4116 464 4118
rect 292 4100 371 4116
rect 378 4114 408 4116
rect -1 4078 28 4088
rect 43 4078 73 4092
rect 116 4078 159 4092
rect 181 4088 371 4100
rect 436 4096 442 4116
rect 166 4078 196 4088
rect 197 4078 355 4088
rect 359 4078 389 4088
rect 393 4078 423 4092
rect 451 4078 464 4116
rect 536 4130 565 4146
rect 579 4130 608 4146
rect 623 4136 653 4152
rect 681 4130 687 4178
rect 690 4172 709 4178
rect 724 4172 754 4180
rect 690 4164 754 4172
rect 690 4148 770 4164
rect 786 4157 848 4188
rect 864 4157 926 4188
rect 995 4186 1044 4211
rect 1059 4186 1089 4202
rect 958 4172 988 4180
rect 995 4178 1105 4186
rect 958 4164 1003 4172
rect 690 4146 709 4148
rect 724 4146 770 4148
rect 690 4130 770 4146
rect 797 4144 832 4157
rect 873 4154 910 4157
rect 873 4152 915 4154
rect 802 4141 832 4144
rect 811 4137 818 4141
rect 818 4136 819 4137
rect 777 4130 787 4136
rect 536 4122 571 4130
rect 536 4096 537 4122
rect 544 4096 571 4122
rect 479 4078 509 4092
rect 536 4088 571 4096
rect 573 4122 614 4130
rect 573 4096 588 4122
rect 595 4096 614 4122
rect 678 4118 709 4130
rect 724 4118 827 4130
rect 839 4120 865 4146
rect 880 4141 910 4152
rect 942 4148 1004 4164
rect 942 4146 988 4148
rect 942 4130 1004 4146
rect 1016 4130 1022 4178
rect 1025 4170 1105 4178
rect 1025 4168 1044 4170
rect 1059 4168 1093 4170
rect 1025 4152 1105 4168
rect 1025 4130 1044 4152
rect 1059 4136 1089 4152
rect 1117 4146 1123 4220
rect 1126 4146 1145 4290
rect 1160 4146 1166 4290
rect 1175 4220 1188 4290
rect 1240 4286 1262 4290
rect 1233 4264 1262 4278
rect 1315 4264 1331 4278
rect 1369 4274 1375 4276
rect 1382 4274 1490 4290
rect 1497 4274 1503 4276
rect 1511 4274 1526 4290
rect 1592 4284 1611 4287
rect 1233 4262 1331 4264
rect 1358 4262 1526 4274
rect 1541 4264 1557 4278
rect 1592 4265 1614 4284
rect 1624 4278 1640 4279
rect 1623 4276 1640 4278
rect 1624 4271 1640 4276
rect 1614 4264 1620 4265
rect 1623 4264 1652 4271
rect 1541 4263 1652 4264
rect 1541 4262 1658 4263
rect 1217 4254 1268 4262
rect 1315 4254 1349 4262
rect 1217 4242 1242 4254
rect 1249 4242 1268 4254
rect 1322 4252 1349 4254
rect 1358 4252 1579 4262
rect 1614 4259 1620 4262
rect 1322 4248 1579 4252
rect 1217 4234 1268 4242
rect 1315 4234 1579 4248
rect 1623 4254 1658 4262
rect 1169 4186 1188 4220
rect 1233 4226 1262 4234
rect 1233 4220 1250 4226
rect 1233 4218 1267 4220
rect 1315 4218 1331 4234
rect 1332 4224 1540 4234
rect 1541 4224 1557 4234
rect 1605 4230 1620 4245
rect 1623 4242 1624 4254
rect 1631 4242 1658 4254
rect 1623 4234 1658 4242
rect 1623 4233 1652 4234
rect 1343 4220 1557 4224
rect 1358 4218 1557 4220
rect 1592 4220 1605 4230
rect 1623 4220 1640 4233
rect 1592 4218 1640 4220
rect 1234 4214 1267 4218
rect 1230 4212 1267 4214
rect 1230 4211 1297 4212
rect 1230 4206 1261 4211
rect 1267 4206 1297 4211
rect 1230 4202 1297 4206
rect 1203 4199 1297 4202
rect 1203 4192 1252 4199
rect 1203 4186 1233 4192
rect 1252 4187 1257 4192
rect 1169 4170 1249 4186
rect 1261 4178 1297 4199
rect 1358 4194 1547 4218
rect 1592 4217 1639 4218
rect 1605 4212 1639 4217
rect 1373 4191 1547 4194
rect 1366 4188 1547 4191
rect 1575 4211 1639 4212
rect 1169 4168 1188 4170
rect 1203 4168 1237 4170
rect 1169 4152 1249 4168
rect 1169 4146 1188 4152
rect 885 4120 988 4130
rect 839 4118 988 4120
rect 1009 4118 1044 4130
rect 678 4116 840 4118
rect 690 4096 709 4116
rect 724 4114 754 4116
rect 573 4088 614 4096
rect 696 4092 709 4096
rect 761 4100 840 4116
rect 872 4116 1044 4118
rect 872 4100 951 4116
rect 958 4114 988 4116
rect 536 4078 565 4088
rect 579 4078 608 4088
rect 623 4078 653 4092
rect 696 4078 739 4092
rect 761 4088 951 4100
rect 1016 4096 1022 4116
rect 746 4078 776 4088
rect 777 4078 935 4088
rect 939 4078 969 4088
rect 973 4078 1003 4092
rect 1031 4078 1044 4116
rect 1116 4130 1145 4146
rect 1159 4130 1188 4146
rect 1203 4136 1233 4152
rect 1261 4130 1267 4178
rect 1270 4172 1289 4178
rect 1304 4172 1334 4180
rect 1270 4164 1334 4172
rect 1270 4148 1350 4164
rect 1366 4157 1428 4188
rect 1444 4157 1506 4188
rect 1575 4186 1624 4211
rect 1639 4186 1669 4202
rect 1538 4172 1568 4180
rect 1575 4178 1685 4186
rect 1538 4164 1583 4172
rect 1270 4146 1289 4148
rect 1304 4146 1350 4148
rect 1270 4130 1350 4146
rect 1377 4144 1412 4157
rect 1453 4154 1490 4157
rect 1453 4152 1495 4154
rect 1382 4141 1412 4144
rect 1391 4137 1398 4141
rect 1398 4136 1399 4137
rect 1357 4130 1367 4136
rect 1116 4122 1151 4130
rect 1116 4096 1117 4122
rect 1124 4096 1151 4122
rect 1059 4078 1089 4092
rect 1116 4088 1151 4096
rect 1153 4122 1194 4130
rect 1153 4096 1168 4122
rect 1175 4096 1194 4122
rect 1258 4118 1289 4130
rect 1304 4118 1407 4130
rect 1419 4120 1445 4146
rect 1460 4141 1490 4152
rect 1522 4148 1584 4164
rect 1522 4146 1568 4148
rect 1522 4130 1584 4146
rect 1596 4130 1602 4178
rect 1605 4170 1685 4178
rect 1605 4168 1624 4170
rect 1639 4168 1673 4170
rect 1605 4152 1685 4168
rect 1605 4130 1624 4152
rect 1639 4136 1669 4152
rect 1697 4146 1703 4220
rect 1706 4146 1725 4290
rect 1740 4146 1746 4290
rect 1755 4220 1768 4290
rect 1820 4286 1842 4290
rect 1813 4264 1842 4278
rect 1895 4264 1911 4278
rect 1949 4274 1955 4276
rect 1962 4274 2070 4290
rect 2077 4274 2083 4276
rect 2091 4274 2106 4290
rect 2172 4284 2191 4287
rect 1813 4262 1911 4264
rect 1938 4262 2106 4274
rect 2121 4264 2137 4278
rect 2172 4265 2194 4284
rect 2204 4278 2220 4279
rect 2203 4276 2220 4278
rect 2204 4271 2220 4276
rect 2194 4264 2200 4265
rect 2203 4264 2232 4271
rect 2121 4263 2232 4264
rect 2121 4262 2238 4263
rect 1797 4254 1848 4262
rect 1895 4254 1929 4262
rect 1797 4242 1822 4254
rect 1829 4242 1848 4254
rect 1902 4252 1929 4254
rect 1938 4252 2159 4262
rect 2194 4259 2200 4262
rect 1902 4248 2159 4252
rect 1797 4234 1848 4242
rect 1895 4234 2159 4248
rect 2203 4254 2238 4262
rect 1749 4186 1768 4220
rect 1813 4226 1842 4234
rect 1813 4220 1830 4226
rect 1813 4218 1847 4220
rect 1895 4218 1911 4234
rect 1912 4224 2120 4234
rect 2121 4224 2137 4234
rect 2185 4230 2200 4245
rect 2203 4242 2204 4254
rect 2211 4242 2238 4254
rect 2203 4234 2238 4242
rect 2203 4233 2232 4234
rect 1923 4220 2137 4224
rect 1938 4218 2137 4220
rect 2172 4220 2185 4230
rect 2203 4220 2220 4233
rect 2172 4218 2220 4220
rect 1814 4214 1847 4218
rect 1810 4212 1847 4214
rect 1810 4211 1877 4212
rect 1810 4206 1841 4211
rect 1847 4206 1877 4211
rect 1810 4202 1877 4206
rect 1783 4199 1877 4202
rect 1783 4192 1832 4199
rect 1783 4186 1813 4192
rect 1832 4187 1837 4192
rect 1749 4170 1829 4186
rect 1841 4178 1877 4199
rect 1938 4194 2127 4218
rect 2172 4217 2219 4218
rect 2185 4212 2219 4217
rect 1953 4191 2127 4194
rect 1946 4188 2127 4191
rect 2155 4211 2219 4212
rect 1749 4168 1768 4170
rect 1783 4168 1817 4170
rect 1749 4152 1829 4168
rect 1749 4146 1768 4152
rect 1465 4120 1568 4130
rect 1419 4118 1568 4120
rect 1589 4118 1624 4130
rect 1258 4116 1420 4118
rect 1270 4096 1289 4116
rect 1304 4114 1334 4116
rect 1153 4088 1194 4096
rect 1276 4092 1289 4096
rect 1341 4100 1420 4116
rect 1452 4116 1624 4118
rect 1452 4100 1531 4116
rect 1538 4114 1568 4116
rect 1116 4078 1145 4088
rect 1159 4078 1188 4088
rect 1203 4078 1233 4092
rect 1276 4078 1319 4092
rect 1341 4088 1531 4100
rect 1596 4096 1602 4116
rect 1326 4078 1356 4088
rect 1357 4078 1515 4088
rect 1519 4078 1549 4088
rect 1553 4078 1583 4092
rect 1611 4078 1624 4116
rect 1696 4130 1725 4146
rect 1739 4130 1768 4146
rect 1783 4136 1813 4152
rect 1841 4130 1847 4178
rect 1850 4172 1869 4178
rect 1884 4172 1914 4180
rect 1850 4164 1914 4172
rect 1850 4148 1930 4164
rect 1946 4157 2008 4188
rect 2024 4157 2086 4188
rect 2155 4186 2204 4211
rect 2219 4186 2249 4202
rect 2118 4172 2148 4180
rect 2155 4178 2265 4186
rect 2118 4164 2163 4172
rect 1850 4146 1869 4148
rect 1884 4146 1930 4148
rect 1850 4130 1930 4146
rect 1957 4144 1992 4157
rect 2033 4154 2070 4157
rect 2033 4152 2075 4154
rect 1962 4141 1992 4144
rect 1971 4137 1978 4141
rect 1978 4136 1979 4137
rect 1937 4130 1947 4136
rect 1696 4122 1731 4130
rect 1696 4096 1697 4122
rect 1704 4096 1731 4122
rect 1639 4078 1669 4092
rect 1696 4088 1731 4096
rect 1733 4122 1774 4130
rect 1733 4096 1748 4122
rect 1755 4096 1774 4122
rect 1838 4118 1869 4130
rect 1884 4118 1987 4130
rect 1999 4120 2025 4146
rect 2040 4141 2070 4152
rect 2102 4148 2164 4164
rect 2102 4146 2148 4148
rect 2102 4130 2164 4146
rect 2176 4130 2182 4178
rect 2185 4170 2265 4178
rect 2185 4168 2204 4170
rect 2219 4168 2253 4170
rect 2185 4152 2265 4168
rect 2185 4130 2204 4152
rect 2219 4136 2249 4152
rect 2277 4146 2283 4220
rect 2286 4146 2305 4290
rect 2320 4146 2326 4290
rect 2335 4220 2348 4290
rect 2400 4286 2422 4290
rect 2393 4264 2422 4278
rect 2475 4264 2491 4278
rect 2529 4274 2535 4276
rect 2542 4274 2650 4290
rect 2657 4274 2663 4276
rect 2671 4274 2686 4290
rect 2752 4284 2771 4287
rect 2393 4262 2491 4264
rect 2518 4262 2686 4274
rect 2701 4264 2717 4278
rect 2752 4265 2774 4284
rect 2784 4278 2800 4279
rect 2783 4276 2800 4278
rect 2784 4271 2800 4276
rect 2774 4264 2780 4265
rect 2783 4264 2812 4271
rect 2701 4263 2812 4264
rect 2701 4262 2818 4263
rect 2377 4254 2428 4262
rect 2475 4254 2509 4262
rect 2377 4242 2402 4254
rect 2409 4242 2428 4254
rect 2482 4252 2509 4254
rect 2518 4252 2739 4262
rect 2774 4259 2780 4262
rect 2482 4248 2739 4252
rect 2377 4234 2428 4242
rect 2475 4234 2739 4248
rect 2783 4254 2818 4262
rect 2329 4186 2348 4220
rect 2393 4226 2422 4234
rect 2393 4220 2410 4226
rect 2393 4218 2427 4220
rect 2475 4218 2491 4234
rect 2492 4224 2700 4234
rect 2701 4224 2717 4234
rect 2765 4230 2780 4245
rect 2783 4242 2784 4254
rect 2791 4242 2818 4254
rect 2783 4234 2818 4242
rect 2783 4233 2812 4234
rect 2503 4220 2717 4224
rect 2518 4218 2717 4220
rect 2752 4220 2765 4230
rect 2783 4220 2800 4233
rect 2752 4218 2800 4220
rect 2394 4214 2427 4218
rect 2390 4212 2427 4214
rect 2390 4211 2457 4212
rect 2390 4206 2421 4211
rect 2427 4206 2457 4211
rect 2390 4202 2457 4206
rect 2363 4199 2457 4202
rect 2363 4192 2412 4199
rect 2363 4186 2393 4192
rect 2412 4187 2417 4192
rect 2329 4170 2409 4186
rect 2421 4178 2457 4199
rect 2518 4194 2707 4218
rect 2752 4217 2799 4218
rect 2765 4212 2799 4217
rect 2533 4191 2707 4194
rect 2526 4188 2707 4191
rect 2735 4211 2799 4212
rect 2329 4168 2348 4170
rect 2363 4168 2397 4170
rect 2329 4152 2409 4168
rect 2329 4146 2348 4152
rect 2045 4120 2148 4130
rect 1999 4118 2148 4120
rect 2169 4118 2204 4130
rect 1838 4116 2000 4118
rect 1850 4096 1869 4116
rect 1884 4114 1914 4116
rect 1733 4088 1774 4096
rect 1856 4092 1869 4096
rect 1921 4100 2000 4116
rect 2032 4116 2204 4118
rect 2032 4100 2111 4116
rect 2118 4114 2148 4116
rect 1696 4078 1725 4088
rect 1739 4078 1768 4088
rect 1783 4078 1813 4092
rect 1856 4078 1899 4092
rect 1921 4088 2111 4100
rect 2176 4096 2182 4116
rect 1906 4078 1936 4088
rect 1937 4078 2095 4088
rect 2099 4078 2129 4088
rect 2133 4078 2163 4092
rect 2191 4078 2204 4116
rect 2276 4130 2305 4146
rect 2319 4130 2348 4146
rect 2363 4136 2393 4152
rect 2421 4130 2427 4178
rect 2430 4172 2449 4178
rect 2464 4172 2494 4180
rect 2430 4164 2494 4172
rect 2430 4148 2510 4164
rect 2526 4157 2588 4188
rect 2604 4157 2666 4188
rect 2735 4186 2784 4211
rect 2799 4186 2829 4202
rect 2698 4172 2728 4180
rect 2735 4178 2845 4186
rect 2698 4164 2743 4172
rect 2430 4146 2449 4148
rect 2464 4146 2510 4148
rect 2430 4130 2510 4146
rect 2537 4144 2572 4157
rect 2613 4154 2650 4157
rect 2613 4152 2655 4154
rect 2542 4141 2572 4144
rect 2551 4137 2558 4141
rect 2558 4136 2559 4137
rect 2517 4130 2527 4136
rect 2276 4122 2311 4130
rect 2276 4096 2277 4122
rect 2284 4096 2311 4122
rect 2219 4078 2249 4092
rect 2276 4088 2311 4096
rect 2313 4122 2354 4130
rect 2313 4096 2328 4122
rect 2335 4096 2354 4122
rect 2418 4118 2449 4130
rect 2464 4118 2567 4130
rect 2579 4120 2605 4146
rect 2620 4141 2650 4152
rect 2682 4148 2744 4164
rect 2682 4146 2728 4148
rect 2682 4130 2744 4146
rect 2756 4130 2762 4178
rect 2765 4170 2845 4178
rect 2765 4168 2784 4170
rect 2799 4168 2833 4170
rect 2765 4152 2845 4168
rect 2765 4130 2784 4152
rect 2799 4136 2829 4152
rect 2857 4146 2863 4220
rect 2866 4146 2885 4290
rect 2900 4146 2906 4290
rect 2915 4220 2928 4290
rect 2980 4286 3002 4290
rect 2973 4264 3002 4278
rect 3055 4264 3071 4278
rect 3109 4274 3115 4276
rect 3122 4274 3230 4290
rect 3237 4274 3243 4276
rect 3251 4274 3266 4290
rect 3332 4284 3351 4287
rect 2973 4262 3071 4264
rect 3098 4262 3266 4274
rect 3281 4264 3297 4278
rect 3332 4265 3354 4284
rect 3364 4278 3380 4279
rect 3363 4276 3380 4278
rect 3364 4271 3380 4276
rect 3354 4264 3360 4265
rect 3363 4264 3392 4271
rect 3281 4263 3392 4264
rect 3281 4262 3398 4263
rect 2957 4254 3008 4262
rect 3055 4254 3089 4262
rect 2957 4242 2982 4254
rect 2989 4242 3008 4254
rect 3062 4252 3089 4254
rect 3098 4252 3319 4262
rect 3354 4259 3360 4262
rect 3062 4248 3319 4252
rect 2957 4234 3008 4242
rect 3055 4234 3319 4248
rect 3363 4254 3398 4262
rect 2909 4186 2928 4220
rect 2973 4226 3002 4234
rect 2973 4220 2990 4226
rect 2973 4218 3007 4220
rect 3055 4218 3071 4234
rect 3072 4224 3280 4234
rect 3281 4224 3297 4234
rect 3345 4230 3360 4245
rect 3363 4242 3364 4254
rect 3371 4242 3398 4254
rect 3363 4234 3398 4242
rect 3363 4233 3392 4234
rect 3083 4220 3297 4224
rect 3098 4218 3297 4220
rect 3332 4220 3345 4230
rect 3363 4220 3380 4233
rect 3332 4218 3380 4220
rect 2974 4214 3007 4218
rect 2970 4212 3007 4214
rect 2970 4211 3037 4212
rect 2970 4206 3001 4211
rect 3007 4206 3037 4211
rect 2970 4202 3037 4206
rect 2943 4199 3037 4202
rect 2943 4192 2992 4199
rect 2943 4186 2973 4192
rect 2992 4187 2997 4192
rect 2909 4170 2989 4186
rect 3001 4178 3037 4199
rect 3098 4194 3287 4218
rect 3332 4217 3379 4218
rect 3345 4212 3379 4217
rect 3113 4191 3287 4194
rect 3106 4188 3287 4191
rect 3315 4211 3379 4212
rect 2909 4168 2928 4170
rect 2943 4168 2977 4170
rect 2909 4152 2989 4168
rect 2909 4146 2928 4152
rect 2625 4120 2728 4130
rect 2579 4118 2728 4120
rect 2749 4118 2784 4130
rect 2418 4116 2580 4118
rect 2430 4096 2449 4116
rect 2464 4114 2494 4116
rect 2313 4088 2354 4096
rect 2436 4092 2449 4096
rect 2501 4100 2580 4116
rect 2612 4116 2784 4118
rect 2612 4100 2691 4116
rect 2698 4114 2728 4116
rect 2276 4078 2305 4088
rect 2319 4078 2348 4088
rect 2363 4078 2393 4092
rect 2436 4078 2479 4092
rect 2501 4088 2691 4100
rect 2756 4096 2762 4116
rect 2486 4078 2516 4088
rect 2517 4078 2675 4088
rect 2679 4078 2709 4088
rect 2713 4078 2743 4092
rect 2771 4078 2784 4116
rect 2856 4130 2885 4146
rect 2899 4130 2928 4146
rect 2943 4136 2973 4152
rect 3001 4130 3007 4178
rect 3010 4172 3029 4178
rect 3044 4172 3074 4180
rect 3010 4164 3074 4172
rect 3010 4148 3090 4164
rect 3106 4157 3168 4188
rect 3184 4157 3246 4188
rect 3315 4186 3364 4211
rect 3379 4186 3409 4202
rect 3278 4172 3308 4180
rect 3315 4178 3425 4186
rect 3278 4164 3323 4172
rect 3010 4146 3029 4148
rect 3044 4146 3090 4148
rect 3010 4130 3090 4146
rect 3117 4144 3152 4157
rect 3193 4154 3230 4157
rect 3193 4152 3235 4154
rect 3122 4141 3152 4144
rect 3131 4137 3138 4141
rect 3138 4136 3139 4137
rect 3097 4130 3107 4136
rect 2856 4122 2891 4130
rect 2856 4096 2857 4122
rect 2864 4096 2891 4122
rect 2799 4078 2829 4092
rect 2856 4088 2891 4096
rect 2893 4122 2934 4130
rect 2893 4096 2908 4122
rect 2915 4096 2934 4122
rect 2998 4118 3029 4130
rect 3044 4118 3147 4130
rect 3159 4120 3185 4146
rect 3200 4141 3230 4152
rect 3262 4148 3324 4164
rect 3262 4146 3308 4148
rect 3262 4130 3324 4146
rect 3336 4130 3342 4178
rect 3345 4170 3425 4178
rect 3345 4168 3364 4170
rect 3379 4168 3413 4170
rect 3345 4152 3425 4168
rect 3345 4130 3364 4152
rect 3379 4136 3409 4152
rect 3437 4146 3443 4220
rect 3446 4146 3465 4290
rect 3480 4146 3486 4290
rect 3495 4220 3508 4290
rect 3560 4286 3582 4290
rect 3553 4264 3582 4278
rect 3635 4264 3651 4278
rect 3689 4274 3695 4276
rect 3702 4274 3810 4290
rect 3817 4274 3823 4276
rect 3831 4274 3846 4290
rect 3912 4284 3931 4287
rect 3553 4262 3651 4264
rect 3678 4262 3846 4274
rect 3861 4264 3877 4278
rect 3912 4265 3934 4284
rect 3944 4278 3960 4279
rect 3943 4276 3960 4278
rect 3944 4271 3960 4276
rect 3934 4264 3940 4265
rect 3943 4264 3972 4271
rect 3861 4263 3972 4264
rect 3861 4262 3978 4263
rect 3537 4254 3588 4262
rect 3635 4254 3669 4262
rect 3537 4242 3562 4254
rect 3569 4242 3588 4254
rect 3642 4252 3669 4254
rect 3678 4252 3899 4262
rect 3934 4259 3940 4262
rect 3642 4248 3899 4252
rect 3537 4234 3588 4242
rect 3635 4234 3899 4248
rect 3943 4254 3978 4262
rect 3489 4186 3508 4220
rect 3553 4226 3582 4234
rect 3553 4220 3570 4226
rect 3553 4218 3587 4220
rect 3635 4218 3651 4234
rect 3652 4224 3860 4234
rect 3861 4224 3877 4234
rect 3925 4230 3940 4245
rect 3943 4242 3944 4254
rect 3951 4242 3978 4254
rect 3943 4234 3978 4242
rect 3943 4233 3972 4234
rect 3663 4220 3877 4224
rect 3678 4218 3877 4220
rect 3912 4220 3925 4230
rect 3943 4220 3960 4233
rect 3912 4218 3960 4220
rect 3554 4214 3587 4218
rect 3550 4212 3587 4214
rect 3550 4211 3617 4212
rect 3550 4206 3581 4211
rect 3587 4206 3617 4211
rect 3550 4202 3617 4206
rect 3523 4199 3617 4202
rect 3523 4192 3572 4199
rect 3523 4186 3553 4192
rect 3572 4187 3577 4192
rect 3489 4170 3569 4186
rect 3581 4178 3617 4199
rect 3678 4194 3867 4218
rect 3912 4217 3959 4218
rect 3925 4212 3959 4217
rect 3693 4191 3867 4194
rect 3686 4188 3867 4191
rect 3895 4211 3959 4212
rect 3489 4168 3508 4170
rect 3523 4168 3557 4170
rect 3489 4152 3569 4168
rect 3489 4146 3508 4152
rect 3205 4120 3308 4130
rect 3159 4118 3308 4120
rect 3329 4118 3364 4130
rect 2998 4116 3160 4118
rect 3010 4096 3029 4116
rect 3044 4114 3074 4116
rect 2893 4088 2934 4096
rect 3016 4092 3029 4096
rect 3081 4100 3160 4116
rect 3192 4116 3364 4118
rect 3192 4100 3271 4116
rect 3278 4114 3308 4116
rect 2856 4078 2885 4088
rect 2899 4078 2928 4088
rect 2943 4078 2973 4092
rect 3016 4078 3059 4092
rect 3081 4088 3271 4100
rect 3336 4096 3342 4116
rect 3066 4078 3096 4088
rect 3097 4078 3255 4088
rect 3259 4078 3289 4088
rect 3293 4078 3323 4092
rect 3351 4078 3364 4116
rect 3436 4130 3465 4146
rect 3479 4130 3508 4146
rect 3523 4136 3553 4152
rect 3581 4130 3587 4178
rect 3590 4172 3609 4178
rect 3624 4172 3654 4180
rect 3590 4164 3654 4172
rect 3590 4148 3670 4164
rect 3686 4157 3748 4188
rect 3764 4157 3826 4188
rect 3895 4186 3944 4211
rect 3959 4186 3989 4202
rect 3858 4172 3888 4180
rect 3895 4178 4005 4186
rect 3858 4164 3903 4172
rect 3590 4146 3609 4148
rect 3624 4146 3670 4148
rect 3590 4130 3670 4146
rect 3697 4144 3732 4157
rect 3773 4154 3810 4157
rect 3773 4152 3815 4154
rect 3702 4141 3732 4144
rect 3711 4137 3718 4141
rect 3718 4136 3719 4137
rect 3677 4130 3687 4136
rect 3436 4122 3471 4130
rect 3436 4096 3437 4122
rect 3444 4096 3471 4122
rect 3379 4078 3409 4092
rect 3436 4088 3471 4096
rect 3473 4122 3514 4130
rect 3473 4096 3488 4122
rect 3495 4096 3514 4122
rect 3578 4118 3609 4130
rect 3624 4118 3727 4130
rect 3739 4120 3765 4146
rect 3780 4141 3810 4152
rect 3842 4148 3904 4164
rect 3842 4146 3888 4148
rect 3842 4130 3904 4146
rect 3916 4130 3922 4178
rect 3925 4170 4005 4178
rect 3925 4168 3944 4170
rect 3959 4168 3993 4170
rect 3925 4152 4005 4168
rect 3925 4130 3944 4152
rect 3959 4136 3989 4152
rect 4017 4146 4023 4220
rect 4026 4146 4045 4290
rect 4060 4146 4066 4290
rect 4075 4220 4088 4290
rect 4140 4286 4162 4290
rect 4133 4264 4162 4278
rect 4215 4264 4231 4278
rect 4269 4274 4275 4276
rect 4282 4274 4390 4290
rect 4397 4274 4403 4276
rect 4411 4274 4426 4290
rect 4492 4284 4511 4287
rect 4133 4262 4231 4264
rect 4258 4262 4426 4274
rect 4441 4264 4457 4278
rect 4492 4265 4514 4284
rect 4524 4278 4540 4279
rect 4523 4276 4540 4278
rect 4524 4271 4540 4276
rect 4514 4264 4520 4265
rect 4523 4264 4552 4271
rect 4441 4263 4552 4264
rect 4441 4262 4558 4263
rect 4117 4254 4168 4262
rect 4215 4254 4249 4262
rect 4117 4242 4142 4254
rect 4149 4242 4168 4254
rect 4222 4252 4249 4254
rect 4258 4252 4479 4262
rect 4514 4259 4520 4262
rect 4222 4248 4479 4252
rect 4117 4234 4168 4242
rect 4215 4234 4479 4248
rect 4523 4254 4558 4262
rect 4069 4186 4088 4220
rect 4133 4226 4162 4234
rect 4133 4220 4150 4226
rect 4133 4218 4167 4220
rect 4215 4218 4231 4234
rect 4232 4224 4440 4234
rect 4441 4224 4457 4234
rect 4505 4230 4520 4245
rect 4523 4242 4524 4254
rect 4531 4242 4558 4254
rect 4523 4234 4558 4242
rect 4523 4233 4552 4234
rect 4243 4220 4457 4224
rect 4258 4218 4457 4220
rect 4492 4220 4505 4230
rect 4523 4220 4540 4233
rect 4492 4218 4540 4220
rect 4134 4214 4167 4218
rect 4130 4212 4167 4214
rect 4130 4211 4197 4212
rect 4130 4206 4161 4211
rect 4167 4206 4197 4211
rect 4130 4202 4197 4206
rect 4103 4199 4197 4202
rect 4103 4192 4152 4199
rect 4103 4186 4133 4192
rect 4152 4187 4157 4192
rect 4069 4170 4149 4186
rect 4161 4178 4197 4199
rect 4258 4194 4447 4218
rect 4492 4217 4539 4218
rect 4505 4212 4539 4217
rect 4273 4191 4447 4194
rect 4266 4188 4447 4191
rect 4475 4211 4539 4212
rect 4069 4168 4088 4170
rect 4103 4168 4137 4170
rect 4069 4152 4149 4168
rect 4069 4146 4088 4152
rect 3785 4120 3888 4130
rect 3739 4118 3888 4120
rect 3909 4118 3944 4130
rect 3578 4116 3740 4118
rect 3590 4096 3609 4116
rect 3624 4114 3654 4116
rect 3473 4088 3514 4096
rect 3596 4092 3609 4096
rect 3661 4100 3740 4116
rect 3772 4116 3944 4118
rect 3772 4100 3851 4116
rect 3858 4114 3888 4116
rect 3436 4078 3465 4088
rect 3479 4078 3508 4088
rect 3523 4078 3553 4092
rect 3596 4078 3639 4092
rect 3661 4088 3851 4100
rect 3916 4096 3922 4116
rect 3646 4078 3676 4088
rect 3677 4078 3835 4088
rect 3839 4078 3869 4088
rect 3873 4078 3903 4092
rect 3931 4078 3944 4116
rect 4016 4130 4045 4146
rect 4059 4130 4088 4146
rect 4103 4136 4133 4152
rect 4161 4130 4167 4178
rect 4170 4172 4189 4178
rect 4204 4172 4234 4180
rect 4170 4164 4234 4172
rect 4170 4148 4250 4164
rect 4266 4157 4328 4188
rect 4344 4157 4406 4188
rect 4475 4186 4524 4211
rect 4539 4186 4569 4202
rect 4438 4172 4468 4180
rect 4475 4178 4585 4186
rect 4438 4164 4483 4172
rect 4170 4146 4189 4148
rect 4204 4146 4250 4148
rect 4170 4130 4250 4146
rect 4277 4144 4312 4157
rect 4353 4154 4390 4157
rect 4353 4152 4395 4154
rect 4282 4141 4312 4144
rect 4291 4137 4298 4141
rect 4298 4136 4299 4137
rect 4257 4130 4267 4136
rect 4016 4122 4051 4130
rect 4016 4096 4017 4122
rect 4024 4096 4051 4122
rect 3959 4078 3989 4092
rect 4016 4088 4051 4096
rect 4053 4122 4094 4130
rect 4053 4096 4068 4122
rect 4075 4096 4094 4122
rect 4158 4118 4189 4130
rect 4204 4118 4307 4130
rect 4319 4120 4345 4146
rect 4360 4141 4390 4152
rect 4422 4148 4484 4164
rect 4422 4146 4468 4148
rect 4422 4130 4484 4146
rect 4496 4130 4502 4178
rect 4505 4170 4585 4178
rect 4505 4168 4524 4170
rect 4539 4168 4573 4170
rect 4505 4152 4585 4168
rect 4505 4130 4524 4152
rect 4539 4136 4569 4152
rect 4597 4146 4603 4220
rect 4606 4146 4625 4290
rect 4640 4146 4646 4290
rect 4655 4220 4668 4290
rect 4720 4286 4742 4290
rect 4713 4264 4742 4278
rect 4795 4264 4811 4278
rect 4849 4274 4855 4276
rect 4862 4274 4970 4290
rect 4977 4274 4983 4276
rect 4991 4274 5006 4290
rect 5072 4284 5091 4287
rect 4713 4262 4811 4264
rect 4838 4262 5006 4274
rect 5021 4264 5037 4278
rect 5072 4265 5094 4284
rect 5104 4278 5120 4279
rect 5103 4276 5120 4278
rect 5104 4271 5120 4276
rect 5094 4264 5100 4265
rect 5103 4264 5132 4271
rect 5021 4263 5132 4264
rect 5021 4262 5138 4263
rect 4697 4254 4748 4262
rect 4795 4254 4829 4262
rect 4697 4242 4722 4254
rect 4729 4242 4748 4254
rect 4802 4252 4829 4254
rect 4838 4252 5059 4262
rect 5094 4259 5100 4262
rect 4802 4248 5059 4252
rect 4697 4234 4748 4242
rect 4795 4234 5059 4248
rect 5103 4254 5138 4262
rect 4649 4186 4668 4220
rect 4713 4226 4742 4234
rect 4713 4220 4730 4226
rect 4713 4218 4747 4220
rect 4795 4218 4811 4234
rect 4812 4224 5020 4234
rect 5021 4224 5037 4234
rect 5085 4230 5100 4245
rect 5103 4242 5104 4254
rect 5111 4242 5138 4254
rect 5103 4234 5138 4242
rect 5103 4233 5132 4234
rect 4823 4220 5037 4224
rect 4838 4218 5037 4220
rect 5072 4220 5085 4230
rect 5103 4220 5120 4233
rect 5072 4218 5120 4220
rect 4714 4214 4747 4218
rect 4710 4212 4747 4214
rect 4710 4211 4777 4212
rect 4710 4206 4741 4211
rect 4747 4206 4777 4211
rect 4710 4202 4777 4206
rect 4683 4199 4777 4202
rect 4683 4192 4732 4199
rect 4683 4186 4713 4192
rect 4732 4187 4737 4192
rect 4649 4170 4729 4186
rect 4741 4178 4777 4199
rect 4838 4194 5027 4218
rect 5072 4217 5119 4218
rect 5085 4212 5119 4217
rect 4853 4191 5027 4194
rect 4846 4188 5027 4191
rect 5055 4211 5119 4212
rect 4649 4168 4668 4170
rect 4683 4168 4717 4170
rect 4649 4152 4729 4168
rect 4649 4146 4668 4152
rect 4365 4120 4468 4130
rect 4319 4118 4468 4120
rect 4489 4118 4524 4130
rect 4158 4116 4320 4118
rect 4170 4096 4189 4116
rect 4204 4114 4234 4116
rect 4053 4088 4094 4096
rect 4176 4092 4189 4096
rect 4241 4100 4320 4116
rect 4352 4116 4524 4118
rect 4352 4100 4431 4116
rect 4438 4114 4468 4116
rect 4016 4078 4045 4088
rect 4059 4078 4088 4088
rect 4103 4078 4133 4092
rect 4176 4078 4219 4092
rect 4241 4088 4431 4100
rect 4496 4096 4502 4116
rect 4226 4078 4256 4088
rect 4257 4078 4415 4088
rect 4419 4078 4449 4088
rect 4453 4078 4483 4092
rect 4511 4078 4524 4116
rect 4596 4130 4625 4146
rect 4639 4130 4668 4146
rect 4683 4136 4713 4152
rect 4741 4130 4747 4178
rect 4750 4172 4769 4178
rect 4784 4172 4814 4180
rect 4750 4164 4814 4172
rect 4750 4148 4830 4164
rect 4846 4157 4908 4188
rect 4924 4157 4986 4188
rect 5055 4186 5104 4211
rect 5119 4186 5149 4202
rect 5018 4172 5048 4180
rect 5055 4178 5165 4186
rect 5018 4164 5063 4172
rect 4750 4146 4769 4148
rect 4784 4146 4830 4148
rect 4750 4130 4830 4146
rect 4857 4144 4892 4157
rect 4933 4154 4970 4157
rect 4933 4152 4975 4154
rect 4862 4141 4892 4144
rect 4871 4137 4878 4141
rect 4878 4136 4879 4137
rect 4837 4130 4847 4136
rect 4596 4122 4631 4130
rect 4596 4096 4597 4122
rect 4604 4096 4631 4122
rect 4539 4078 4569 4092
rect 4596 4088 4631 4096
rect 4633 4122 4674 4130
rect 4633 4096 4648 4122
rect 4655 4096 4674 4122
rect 4738 4118 4769 4130
rect 4784 4118 4887 4130
rect 4899 4120 4925 4146
rect 4940 4141 4970 4152
rect 5002 4148 5064 4164
rect 5002 4146 5048 4148
rect 5002 4130 5064 4146
rect 5076 4130 5082 4178
rect 5085 4170 5165 4178
rect 5085 4168 5104 4170
rect 5119 4168 5153 4170
rect 5085 4152 5165 4168
rect 5085 4130 5104 4152
rect 5119 4136 5149 4152
rect 5177 4146 5183 4220
rect 5186 4146 5205 4290
rect 5220 4146 5226 4290
rect 5235 4220 5248 4290
rect 5300 4286 5322 4290
rect 5293 4264 5322 4278
rect 5375 4264 5391 4278
rect 5429 4274 5435 4276
rect 5442 4274 5550 4290
rect 5557 4274 5563 4276
rect 5571 4274 5586 4290
rect 5652 4284 5671 4287
rect 5293 4262 5391 4264
rect 5418 4262 5586 4274
rect 5601 4264 5617 4278
rect 5652 4265 5674 4284
rect 5684 4278 5700 4279
rect 5683 4276 5700 4278
rect 5684 4271 5700 4276
rect 5674 4264 5680 4265
rect 5683 4264 5712 4271
rect 5601 4263 5712 4264
rect 5601 4262 5718 4263
rect 5277 4254 5328 4262
rect 5375 4254 5409 4262
rect 5277 4242 5302 4254
rect 5309 4242 5328 4254
rect 5382 4252 5409 4254
rect 5418 4252 5639 4262
rect 5674 4259 5680 4262
rect 5382 4248 5639 4252
rect 5277 4234 5328 4242
rect 5375 4234 5639 4248
rect 5683 4254 5718 4262
rect 5229 4186 5248 4220
rect 5293 4226 5322 4234
rect 5293 4220 5310 4226
rect 5293 4218 5327 4220
rect 5375 4218 5391 4234
rect 5392 4224 5600 4234
rect 5601 4224 5617 4234
rect 5665 4230 5680 4245
rect 5683 4242 5684 4254
rect 5691 4242 5718 4254
rect 5683 4234 5718 4242
rect 5683 4233 5712 4234
rect 5403 4220 5617 4224
rect 5418 4218 5617 4220
rect 5652 4220 5665 4230
rect 5683 4220 5700 4233
rect 5652 4218 5700 4220
rect 5294 4214 5327 4218
rect 5290 4212 5327 4214
rect 5290 4211 5357 4212
rect 5290 4206 5321 4211
rect 5327 4206 5357 4211
rect 5290 4202 5357 4206
rect 5263 4199 5357 4202
rect 5263 4192 5312 4199
rect 5263 4186 5293 4192
rect 5312 4187 5317 4192
rect 5229 4170 5309 4186
rect 5321 4178 5357 4199
rect 5418 4194 5607 4218
rect 5652 4217 5699 4218
rect 5665 4212 5699 4217
rect 5433 4191 5607 4194
rect 5426 4188 5607 4191
rect 5635 4211 5699 4212
rect 5229 4168 5248 4170
rect 5263 4168 5297 4170
rect 5229 4152 5309 4168
rect 5229 4146 5248 4152
rect 4945 4120 5048 4130
rect 4899 4118 5048 4120
rect 5069 4118 5104 4130
rect 4738 4116 4900 4118
rect 4750 4096 4769 4116
rect 4784 4114 4814 4116
rect 4633 4088 4674 4096
rect 4756 4092 4769 4096
rect 4821 4100 4900 4116
rect 4932 4116 5104 4118
rect 4932 4100 5011 4116
rect 5018 4114 5048 4116
rect 4596 4078 4625 4088
rect 4639 4078 4668 4088
rect 4683 4078 4713 4092
rect 4756 4078 4799 4092
rect 4821 4088 5011 4100
rect 5076 4096 5082 4116
rect 4806 4078 4836 4088
rect 4837 4078 4995 4088
rect 4999 4078 5029 4088
rect 5033 4078 5063 4092
rect 5091 4078 5104 4116
rect 5176 4130 5205 4146
rect 5219 4130 5248 4146
rect 5263 4136 5293 4152
rect 5321 4130 5327 4178
rect 5330 4172 5349 4178
rect 5364 4172 5394 4180
rect 5330 4164 5394 4172
rect 5330 4148 5410 4164
rect 5426 4157 5488 4188
rect 5504 4157 5566 4188
rect 5635 4186 5684 4211
rect 5699 4186 5729 4202
rect 5598 4172 5628 4180
rect 5635 4178 5745 4186
rect 5598 4164 5643 4172
rect 5330 4146 5349 4148
rect 5364 4146 5410 4148
rect 5330 4130 5410 4146
rect 5437 4144 5472 4157
rect 5513 4154 5550 4157
rect 5513 4152 5555 4154
rect 5442 4141 5472 4144
rect 5451 4137 5458 4141
rect 5458 4136 5459 4137
rect 5417 4130 5427 4136
rect 5176 4122 5211 4130
rect 5176 4096 5177 4122
rect 5184 4096 5211 4122
rect 5119 4078 5149 4092
rect 5176 4088 5211 4096
rect 5213 4122 5254 4130
rect 5213 4096 5228 4122
rect 5235 4096 5254 4122
rect 5318 4118 5349 4130
rect 5364 4118 5467 4130
rect 5479 4120 5505 4146
rect 5520 4141 5550 4152
rect 5582 4148 5644 4164
rect 5582 4146 5628 4148
rect 5582 4130 5644 4146
rect 5656 4130 5662 4178
rect 5665 4170 5745 4178
rect 5665 4168 5684 4170
rect 5699 4168 5733 4170
rect 5665 4152 5745 4168
rect 5665 4130 5684 4152
rect 5699 4136 5729 4152
rect 5757 4146 5763 4220
rect 5766 4146 5785 4290
rect 5800 4146 5806 4290
rect 5815 4220 5828 4290
rect 5880 4286 5902 4290
rect 5873 4264 5902 4278
rect 5955 4264 5971 4278
rect 6009 4274 6015 4276
rect 6022 4274 6130 4290
rect 6137 4274 6143 4276
rect 6151 4274 6166 4290
rect 6232 4284 6251 4287
rect 5873 4262 5971 4264
rect 5998 4262 6166 4274
rect 6181 4264 6197 4278
rect 6232 4265 6254 4284
rect 6264 4278 6280 4279
rect 6263 4276 6280 4278
rect 6264 4271 6280 4276
rect 6254 4264 6260 4265
rect 6263 4264 6292 4271
rect 6181 4263 6292 4264
rect 6181 4262 6298 4263
rect 5857 4254 5908 4262
rect 5955 4254 5989 4262
rect 5857 4242 5882 4254
rect 5889 4242 5908 4254
rect 5962 4252 5989 4254
rect 5998 4252 6219 4262
rect 6254 4259 6260 4262
rect 5962 4248 6219 4252
rect 5857 4234 5908 4242
rect 5955 4234 6219 4248
rect 6263 4254 6298 4262
rect 5809 4186 5828 4220
rect 5873 4226 5902 4234
rect 5873 4220 5890 4226
rect 5873 4218 5907 4220
rect 5955 4218 5971 4234
rect 5972 4224 6180 4234
rect 6181 4224 6197 4234
rect 6245 4230 6260 4245
rect 6263 4242 6264 4254
rect 6271 4242 6298 4254
rect 6263 4234 6298 4242
rect 6263 4233 6292 4234
rect 5983 4220 6197 4224
rect 5998 4218 6197 4220
rect 6232 4220 6245 4230
rect 6263 4220 6280 4233
rect 6232 4218 6280 4220
rect 5874 4214 5907 4218
rect 5870 4212 5907 4214
rect 5870 4211 5937 4212
rect 5870 4206 5901 4211
rect 5907 4206 5937 4211
rect 5870 4202 5937 4206
rect 5843 4199 5937 4202
rect 5843 4192 5892 4199
rect 5843 4186 5873 4192
rect 5892 4187 5897 4192
rect 5809 4170 5889 4186
rect 5901 4178 5937 4199
rect 5998 4194 6187 4218
rect 6232 4217 6279 4218
rect 6245 4212 6279 4217
rect 6013 4191 6187 4194
rect 6006 4188 6187 4191
rect 6215 4211 6279 4212
rect 5809 4168 5828 4170
rect 5843 4168 5877 4170
rect 5809 4152 5889 4168
rect 5809 4146 5828 4152
rect 5525 4120 5628 4130
rect 5479 4118 5628 4120
rect 5649 4118 5684 4130
rect 5318 4116 5480 4118
rect 5330 4096 5349 4116
rect 5364 4114 5394 4116
rect 5213 4088 5254 4096
rect 5336 4092 5349 4096
rect 5401 4100 5480 4116
rect 5512 4116 5684 4118
rect 5512 4100 5591 4116
rect 5598 4114 5628 4116
rect 5176 4078 5205 4088
rect 5219 4078 5248 4088
rect 5263 4078 5293 4092
rect 5336 4078 5379 4092
rect 5401 4088 5591 4100
rect 5656 4096 5662 4116
rect 5386 4078 5416 4088
rect 5417 4078 5575 4088
rect 5579 4078 5609 4088
rect 5613 4078 5643 4092
rect 5671 4078 5684 4116
rect 5756 4130 5785 4146
rect 5799 4130 5828 4146
rect 5843 4136 5873 4152
rect 5901 4130 5907 4178
rect 5910 4172 5929 4178
rect 5944 4172 5974 4180
rect 5910 4164 5974 4172
rect 5910 4148 5990 4164
rect 6006 4157 6068 4188
rect 6084 4157 6146 4188
rect 6215 4186 6264 4211
rect 6279 4186 6309 4202
rect 6178 4172 6208 4180
rect 6215 4178 6325 4186
rect 6178 4164 6223 4172
rect 5910 4146 5929 4148
rect 5944 4146 5990 4148
rect 5910 4130 5990 4146
rect 6017 4144 6052 4157
rect 6093 4154 6130 4157
rect 6093 4152 6135 4154
rect 6022 4141 6052 4144
rect 6031 4137 6038 4141
rect 6038 4136 6039 4137
rect 5997 4130 6007 4136
rect 5756 4122 5791 4130
rect 5756 4096 5757 4122
rect 5764 4096 5791 4122
rect 5699 4078 5729 4092
rect 5756 4088 5791 4096
rect 5793 4122 5834 4130
rect 5793 4096 5808 4122
rect 5815 4096 5834 4122
rect 5898 4118 5929 4130
rect 5944 4118 6047 4130
rect 6059 4120 6085 4146
rect 6100 4141 6130 4152
rect 6162 4148 6224 4164
rect 6162 4146 6208 4148
rect 6162 4130 6224 4146
rect 6236 4130 6242 4178
rect 6245 4170 6325 4178
rect 6245 4168 6264 4170
rect 6279 4168 6313 4170
rect 6245 4152 6325 4168
rect 6245 4130 6264 4152
rect 6279 4136 6309 4152
rect 6337 4146 6343 4220
rect 6346 4146 6365 4290
rect 6380 4146 6386 4290
rect 6395 4220 6408 4290
rect 6460 4286 6482 4290
rect 6453 4264 6482 4278
rect 6535 4264 6551 4278
rect 6589 4274 6595 4276
rect 6602 4274 6710 4290
rect 6717 4274 6723 4276
rect 6731 4274 6746 4290
rect 6812 4284 6831 4287
rect 6453 4262 6551 4264
rect 6578 4262 6746 4274
rect 6761 4264 6777 4278
rect 6812 4265 6834 4284
rect 6844 4278 6860 4279
rect 6843 4276 6860 4278
rect 6844 4271 6860 4276
rect 6834 4264 6840 4265
rect 6843 4264 6872 4271
rect 6761 4263 6872 4264
rect 6761 4262 6878 4263
rect 6437 4254 6488 4262
rect 6535 4254 6569 4262
rect 6437 4242 6462 4254
rect 6469 4242 6488 4254
rect 6542 4252 6569 4254
rect 6578 4252 6799 4262
rect 6834 4259 6840 4262
rect 6542 4248 6799 4252
rect 6437 4234 6488 4242
rect 6535 4234 6799 4248
rect 6843 4254 6878 4262
rect 6389 4186 6408 4220
rect 6453 4226 6482 4234
rect 6453 4220 6470 4226
rect 6453 4218 6487 4220
rect 6535 4218 6551 4234
rect 6552 4224 6760 4234
rect 6761 4224 6777 4234
rect 6825 4230 6840 4245
rect 6843 4242 6844 4254
rect 6851 4242 6878 4254
rect 6843 4234 6878 4242
rect 6843 4233 6872 4234
rect 6563 4220 6777 4224
rect 6578 4218 6777 4220
rect 6812 4220 6825 4230
rect 6843 4220 6860 4233
rect 6812 4218 6860 4220
rect 6454 4214 6487 4218
rect 6450 4212 6487 4214
rect 6450 4211 6517 4212
rect 6450 4206 6481 4211
rect 6487 4206 6517 4211
rect 6450 4202 6517 4206
rect 6423 4199 6517 4202
rect 6423 4192 6472 4199
rect 6423 4186 6453 4192
rect 6472 4187 6477 4192
rect 6389 4170 6469 4186
rect 6481 4178 6517 4199
rect 6578 4194 6767 4218
rect 6812 4217 6859 4218
rect 6825 4212 6859 4217
rect 6593 4191 6767 4194
rect 6586 4188 6767 4191
rect 6795 4211 6859 4212
rect 6389 4168 6408 4170
rect 6423 4168 6457 4170
rect 6389 4152 6469 4168
rect 6389 4146 6408 4152
rect 6105 4120 6208 4130
rect 6059 4118 6208 4120
rect 6229 4118 6264 4130
rect 5898 4116 6060 4118
rect 5910 4096 5929 4116
rect 5944 4114 5974 4116
rect 5793 4088 5834 4096
rect 5916 4092 5929 4096
rect 5981 4100 6060 4116
rect 6092 4116 6264 4118
rect 6092 4100 6171 4116
rect 6178 4114 6208 4116
rect 5756 4078 5785 4088
rect 5799 4078 5828 4088
rect 5843 4078 5873 4092
rect 5916 4078 5959 4092
rect 5981 4088 6171 4100
rect 6236 4096 6242 4116
rect 5966 4078 5996 4088
rect 5997 4078 6155 4088
rect 6159 4078 6189 4088
rect 6193 4078 6223 4092
rect 6251 4078 6264 4116
rect 6336 4130 6365 4146
rect 6379 4130 6408 4146
rect 6423 4136 6453 4152
rect 6481 4130 6487 4178
rect 6490 4172 6509 4178
rect 6524 4172 6554 4180
rect 6490 4164 6554 4172
rect 6490 4148 6570 4164
rect 6586 4157 6648 4188
rect 6664 4157 6726 4188
rect 6795 4186 6844 4211
rect 6859 4186 6889 4202
rect 6758 4172 6788 4180
rect 6795 4178 6905 4186
rect 6758 4164 6803 4172
rect 6490 4146 6509 4148
rect 6524 4146 6570 4148
rect 6490 4130 6570 4146
rect 6597 4144 6632 4157
rect 6673 4154 6710 4157
rect 6673 4152 6715 4154
rect 6602 4141 6632 4144
rect 6611 4137 6618 4141
rect 6618 4136 6619 4137
rect 6577 4130 6587 4136
rect 6336 4122 6371 4130
rect 6336 4096 6337 4122
rect 6344 4096 6371 4122
rect 6279 4078 6309 4092
rect 6336 4088 6371 4096
rect 6373 4122 6414 4130
rect 6373 4096 6388 4122
rect 6395 4096 6414 4122
rect 6478 4118 6509 4130
rect 6524 4118 6627 4130
rect 6639 4120 6665 4146
rect 6680 4141 6710 4152
rect 6742 4148 6804 4164
rect 6742 4146 6788 4148
rect 6742 4130 6804 4146
rect 6816 4130 6822 4178
rect 6825 4170 6905 4178
rect 6825 4168 6844 4170
rect 6859 4168 6893 4170
rect 6825 4152 6905 4168
rect 6825 4130 6844 4152
rect 6859 4136 6889 4152
rect 6917 4146 6923 4220
rect 6926 4146 6945 4290
rect 6960 4146 6966 4290
rect 6975 4220 6988 4290
rect 7040 4286 7062 4290
rect 7033 4264 7062 4278
rect 7115 4264 7131 4278
rect 7169 4274 7175 4276
rect 7182 4274 7290 4290
rect 7297 4274 7303 4276
rect 7311 4274 7326 4290
rect 7392 4284 7411 4287
rect 7033 4262 7131 4264
rect 7158 4262 7326 4274
rect 7341 4264 7357 4278
rect 7392 4265 7414 4284
rect 7424 4278 7440 4279
rect 7423 4276 7440 4278
rect 7424 4271 7440 4276
rect 7414 4264 7420 4265
rect 7423 4264 7452 4271
rect 7341 4263 7452 4264
rect 7341 4262 7458 4263
rect 7017 4254 7068 4262
rect 7115 4254 7149 4262
rect 7017 4242 7042 4254
rect 7049 4242 7068 4254
rect 7122 4252 7149 4254
rect 7158 4252 7379 4262
rect 7414 4259 7420 4262
rect 7122 4248 7379 4252
rect 7017 4234 7068 4242
rect 7115 4234 7379 4248
rect 7423 4254 7458 4262
rect 6969 4186 6988 4220
rect 7033 4226 7062 4234
rect 7033 4220 7050 4226
rect 7033 4218 7067 4220
rect 7115 4218 7131 4234
rect 7132 4224 7340 4234
rect 7341 4224 7357 4234
rect 7405 4230 7420 4245
rect 7423 4242 7424 4254
rect 7431 4242 7458 4254
rect 7423 4234 7458 4242
rect 7423 4233 7452 4234
rect 7143 4220 7357 4224
rect 7158 4218 7357 4220
rect 7392 4220 7405 4230
rect 7423 4220 7440 4233
rect 7392 4218 7440 4220
rect 7034 4214 7067 4218
rect 7030 4212 7067 4214
rect 7030 4211 7097 4212
rect 7030 4206 7061 4211
rect 7067 4206 7097 4211
rect 7030 4202 7097 4206
rect 7003 4199 7097 4202
rect 7003 4192 7052 4199
rect 7003 4186 7033 4192
rect 7052 4187 7057 4192
rect 6969 4170 7049 4186
rect 7061 4178 7097 4199
rect 7158 4194 7347 4218
rect 7392 4217 7439 4218
rect 7405 4212 7439 4217
rect 7173 4191 7347 4194
rect 7166 4188 7347 4191
rect 7375 4211 7439 4212
rect 6969 4168 6988 4170
rect 7003 4168 7037 4170
rect 6969 4152 7049 4168
rect 6969 4146 6988 4152
rect 6685 4120 6788 4130
rect 6639 4118 6788 4120
rect 6809 4118 6844 4130
rect 6478 4116 6640 4118
rect 6490 4096 6509 4116
rect 6524 4114 6554 4116
rect 6373 4088 6414 4096
rect 6496 4092 6509 4096
rect 6561 4100 6640 4116
rect 6672 4116 6844 4118
rect 6672 4100 6751 4116
rect 6758 4114 6788 4116
rect 6336 4078 6365 4088
rect 6379 4078 6408 4088
rect 6423 4078 6453 4092
rect 6496 4078 6539 4092
rect 6561 4088 6751 4100
rect 6816 4096 6822 4116
rect 6546 4078 6576 4088
rect 6577 4078 6735 4088
rect 6739 4078 6769 4088
rect 6773 4078 6803 4092
rect 6831 4078 6844 4116
rect 6916 4130 6945 4146
rect 6959 4130 6988 4146
rect 7003 4136 7033 4152
rect 7061 4130 7067 4178
rect 7070 4172 7089 4178
rect 7104 4172 7134 4180
rect 7070 4164 7134 4172
rect 7070 4148 7150 4164
rect 7166 4157 7228 4188
rect 7244 4157 7306 4188
rect 7375 4186 7424 4211
rect 7439 4186 7469 4202
rect 7338 4172 7368 4180
rect 7375 4178 7485 4186
rect 7338 4164 7383 4172
rect 7070 4146 7089 4148
rect 7104 4146 7150 4148
rect 7070 4130 7150 4146
rect 7177 4144 7212 4157
rect 7253 4154 7290 4157
rect 7253 4152 7295 4154
rect 7182 4141 7212 4144
rect 7191 4137 7198 4141
rect 7198 4136 7199 4137
rect 7157 4130 7167 4136
rect 6916 4122 6951 4130
rect 6916 4096 6917 4122
rect 6924 4096 6951 4122
rect 6859 4078 6889 4092
rect 6916 4088 6951 4096
rect 6953 4122 6994 4130
rect 6953 4096 6968 4122
rect 6975 4096 6994 4122
rect 7058 4118 7089 4130
rect 7104 4118 7207 4130
rect 7219 4120 7245 4146
rect 7260 4141 7290 4152
rect 7322 4148 7384 4164
rect 7322 4146 7368 4148
rect 7322 4130 7384 4146
rect 7396 4130 7402 4178
rect 7405 4170 7485 4178
rect 7405 4168 7424 4170
rect 7439 4168 7473 4170
rect 7405 4152 7485 4168
rect 7405 4130 7424 4152
rect 7439 4136 7469 4152
rect 7497 4146 7503 4220
rect 7506 4146 7525 4290
rect 7540 4146 7546 4290
rect 7555 4220 7568 4290
rect 7613 4268 7614 4278
rect 7629 4268 7642 4278
rect 7613 4264 7642 4268
rect 7647 4264 7677 4290
rect 7695 4276 7711 4278
rect 7783 4276 7836 4290
rect 7784 4274 7848 4276
rect 7891 4274 7906 4290
rect 7955 4287 7985 4290
rect 7955 4284 7991 4287
rect 7921 4276 7937 4278
rect 7695 4264 7710 4268
rect 7613 4262 7710 4264
rect 7738 4262 7906 4274
rect 7922 4264 7937 4268
rect 7955 4265 7994 4284
rect 8013 4278 8020 4279
rect 8019 4271 8020 4278
rect 8003 4268 8004 4271
rect 8019 4268 8032 4271
rect 7955 4264 7985 4265
rect 7994 4264 8000 4265
rect 8003 4264 8032 4268
rect 7922 4263 8032 4264
rect 7922 4262 8038 4263
rect 7597 4254 7648 4262
rect 7597 4242 7622 4254
rect 7629 4242 7648 4254
rect 7679 4254 7729 4262
rect 7679 4246 7695 4254
rect 7702 4252 7729 4254
rect 7738 4252 7959 4262
rect 7702 4242 7959 4252
rect 7988 4254 8038 4262
rect 7988 4245 8004 4254
rect 7597 4234 7648 4242
rect 7695 4234 7959 4242
rect 7985 4242 8004 4245
rect 8011 4242 8038 4254
rect 7985 4234 8038 4242
rect 7549 4186 7568 4220
rect 7613 4226 7614 4234
rect 7629 4226 7642 4234
rect 7613 4218 7629 4226
rect 7610 4211 7629 4214
rect 7610 4202 7632 4211
rect 7583 4192 7632 4202
rect 7583 4186 7613 4192
rect 7632 4187 7637 4192
rect 7549 4170 7629 4186
rect 7647 4178 7677 4234
rect 7712 4224 7920 4234
rect 7955 4230 8000 4234
rect 8003 4233 8004 4234
rect 8019 4233 8032 4234
rect 7738 4194 7927 4224
rect 7753 4191 7927 4194
rect 7746 4188 7927 4191
rect 7549 4168 7568 4170
rect 7583 4168 7617 4170
rect 7549 4152 7629 4168
rect 7656 4164 7669 4178
rect 7684 4164 7700 4180
rect 7746 4175 7757 4188
rect 7549 4146 7568 4152
rect 7265 4120 7368 4130
rect 7219 4118 7368 4120
rect 7389 4118 7424 4130
rect 7058 4116 7220 4118
rect 7070 4096 7089 4116
rect 7104 4114 7134 4116
rect 6953 4088 6994 4096
rect 7076 4092 7089 4096
rect 7141 4100 7220 4116
rect 7252 4116 7424 4118
rect 7252 4100 7331 4116
rect 7338 4114 7368 4116
rect 6916 4078 6945 4088
rect 6959 4078 6988 4088
rect 7003 4078 7033 4092
rect 7076 4078 7119 4092
rect 7141 4088 7331 4100
rect 7396 4096 7402 4116
rect 7126 4078 7156 4088
rect 7157 4078 7315 4088
rect 7319 4078 7349 4088
rect 7353 4078 7383 4092
rect 7411 4078 7424 4116
rect 7496 4130 7525 4146
rect 7539 4130 7568 4146
rect 7583 4130 7613 4152
rect 7656 4148 7718 4164
rect 7746 4157 7757 4173
rect 7762 4168 7772 4188
rect 7782 4168 7796 4188
rect 7799 4175 7808 4188
rect 7824 4175 7833 4188
rect 7762 4157 7796 4168
rect 7799 4157 7808 4173
rect 7824 4157 7833 4173
rect 7840 4168 7850 4188
rect 7860 4168 7874 4188
rect 7875 4175 7886 4188
rect 7840 4157 7874 4168
rect 7875 4157 7886 4173
rect 7932 4164 7948 4180
rect 7955 4178 7985 4230
rect 8019 4226 8020 4233
rect 8004 4218 8020 4226
rect 7991 4186 8004 4205
rect 8019 4186 8049 4202
rect 7991 4170 8065 4186
rect 7991 4168 8004 4170
rect 8019 4168 8053 4170
rect 7656 4146 7669 4148
rect 7684 4146 7718 4148
rect 7656 4130 7718 4146
rect 7762 4141 7778 4144
rect 7840 4141 7870 4152
rect 7918 4148 7964 4164
rect 7991 4152 8065 4168
rect 7918 4146 7952 4148
rect 7917 4130 7964 4146
rect 7991 4130 8004 4152
rect 8019 4130 8049 4152
rect 8076 4130 8077 4146
rect 8092 4130 8105 4290
rect 8135 4186 8148 4290
rect 8193 4268 8194 4278
rect 8209 4268 8222 4278
rect 8193 4264 8222 4268
rect 8227 4264 8257 4290
rect 8275 4276 8291 4278
rect 8363 4276 8416 4290
rect 8364 4274 8428 4276
rect 8471 4274 8486 4290
rect 8535 4287 8565 4290
rect 8535 4284 8571 4287
rect 8501 4276 8517 4278
rect 8275 4264 8290 4268
rect 8193 4262 8290 4264
rect 8318 4262 8486 4274
rect 8502 4264 8517 4268
rect 8535 4265 8574 4284
rect 8593 4278 8600 4279
rect 8599 4271 8600 4278
rect 8583 4268 8584 4271
rect 8599 4268 8612 4271
rect 8535 4264 8565 4265
rect 8574 4264 8580 4265
rect 8583 4264 8612 4268
rect 8502 4263 8612 4264
rect 8502 4262 8618 4263
rect 8177 4254 8228 4262
rect 8177 4242 8202 4254
rect 8209 4242 8228 4254
rect 8259 4254 8309 4262
rect 8259 4246 8275 4254
rect 8282 4252 8309 4254
rect 8318 4252 8539 4262
rect 8282 4242 8539 4252
rect 8568 4254 8618 4262
rect 8568 4245 8584 4254
rect 8177 4234 8228 4242
rect 8275 4234 8539 4242
rect 8565 4242 8584 4245
rect 8591 4242 8618 4254
rect 8565 4234 8618 4242
rect 8193 4226 8194 4234
rect 8209 4226 8222 4234
rect 8193 4218 8209 4226
rect 8190 4211 8209 4214
rect 8190 4202 8212 4211
rect 8163 4192 8212 4202
rect 8163 4186 8193 4192
rect 8212 4187 8217 4192
rect 8135 4170 8209 4186
rect 8227 4178 8257 4234
rect 8292 4224 8500 4234
rect 8535 4230 8580 4234
rect 8583 4233 8584 4234
rect 8599 4233 8612 4234
rect 8318 4194 8507 4224
rect 8333 4191 8507 4194
rect 8326 4188 8507 4191
rect 8135 4168 8148 4170
rect 8163 4168 8197 4170
rect 8135 4152 8209 4168
rect 8236 4164 8249 4178
rect 8264 4164 8280 4180
rect 8326 4175 8337 4188
rect 8119 4130 8120 4146
rect 8135 4130 8148 4152
rect 8163 4130 8193 4152
rect 8236 4148 8298 4164
rect 8326 4157 8337 4173
rect 8342 4168 8352 4188
rect 8362 4168 8376 4188
rect 8379 4175 8388 4188
rect 8404 4175 8413 4188
rect 8342 4157 8376 4168
rect 8379 4157 8388 4173
rect 8404 4157 8413 4173
rect 8420 4168 8430 4188
rect 8440 4168 8454 4188
rect 8455 4175 8466 4188
rect 8420 4157 8454 4168
rect 8455 4157 8466 4173
rect 8512 4164 8528 4180
rect 8535 4178 8565 4230
rect 8599 4226 8600 4233
rect 8584 4218 8600 4226
rect 8571 4186 8584 4205
rect 8599 4186 8629 4202
rect 8571 4170 8645 4186
rect 8571 4168 8584 4170
rect 8599 4168 8633 4170
rect 8236 4146 8249 4148
rect 8264 4146 8298 4148
rect 8236 4130 8298 4146
rect 8342 4141 8358 4144
rect 8420 4141 8450 4152
rect 8498 4148 8544 4164
rect 8571 4152 8645 4168
rect 8498 4146 8532 4148
rect 8497 4130 8544 4146
rect 8571 4130 8584 4152
rect 8599 4130 8629 4152
rect 8656 4130 8657 4146
rect 8672 4130 8685 4290
rect 8715 4186 8728 4290
rect 8773 4268 8774 4278
rect 8789 4268 8802 4278
rect 8773 4264 8802 4268
rect 8807 4264 8837 4290
rect 8855 4276 8871 4278
rect 8943 4276 8996 4290
rect 8944 4274 9008 4276
rect 9051 4274 9066 4290
rect 9115 4287 9145 4290
rect 9115 4284 9151 4287
rect 9081 4276 9097 4278
rect 8855 4264 8870 4268
rect 8773 4262 8870 4264
rect 8898 4262 9066 4274
rect 9082 4264 9097 4268
rect 9115 4265 9154 4284
rect 9173 4278 9180 4279
rect 9179 4271 9180 4278
rect 9163 4268 9164 4271
rect 9179 4268 9192 4271
rect 9115 4264 9145 4265
rect 9154 4264 9160 4265
rect 9163 4264 9192 4268
rect 9082 4263 9192 4264
rect 9082 4262 9198 4263
rect 8757 4254 8808 4262
rect 8757 4242 8782 4254
rect 8789 4242 8808 4254
rect 8839 4254 8889 4262
rect 8839 4246 8855 4254
rect 8862 4252 8889 4254
rect 8898 4252 9119 4262
rect 8862 4242 9119 4252
rect 9148 4254 9198 4262
rect 9148 4245 9164 4254
rect 8757 4234 8808 4242
rect 8855 4234 9119 4242
rect 9145 4242 9164 4245
rect 9171 4242 9198 4254
rect 9145 4234 9198 4242
rect 8773 4226 8774 4234
rect 8789 4226 8802 4234
rect 8773 4218 8789 4226
rect 8770 4211 8789 4214
rect 8770 4202 8792 4211
rect 8743 4192 8792 4202
rect 8743 4186 8773 4192
rect 8792 4187 8797 4192
rect 8715 4170 8789 4186
rect 8807 4178 8837 4234
rect 8872 4224 9080 4234
rect 9115 4230 9160 4234
rect 9163 4233 9164 4234
rect 9179 4233 9192 4234
rect 8898 4194 9087 4224
rect 8913 4191 9087 4194
rect 8906 4188 9087 4191
rect 8715 4168 8728 4170
rect 8743 4168 8777 4170
rect 8715 4152 8789 4168
rect 8816 4164 8829 4178
rect 8844 4164 8860 4180
rect 8906 4175 8917 4188
rect 8699 4130 8700 4146
rect 8715 4130 8728 4152
rect 8743 4130 8773 4152
rect 8816 4148 8878 4164
rect 8906 4157 8917 4173
rect 8922 4168 8932 4188
rect 8942 4168 8956 4188
rect 8959 4175 8968 4188
rect 8984 4175 8993 4188
rect 8922 4157 8956 4168
rect 8959 4157 8968 4173
rect 8984 4157 8993 4173
rect 9000 4168 9010 4188
rect 9020 4168 9034 4188
rect 9035 4175 9046 4188
rect 9000 4157 9034 4168
rect 9035 4157 9046 4173
rect 9092 4164 9108 4180
rect 9115 4178 9145 4230
rect 9179 4226 9180 4233
rect 9164 4218 9180 4226
rect 9151 4186 9164 4205
rect 9179 4186 9209 4202
rect 9151 4170 9225 4186
rect 9151 4168 9164 4170
rect 9179 4168 9213 4170
rect 8816 4146 8829 4148
rect 8844 4146 8878 4148
rect 8816 4130 8878 4146
rect 8922 4141 8938 4144
rect 9000 4141 9030 4152
rect 9078 4148 9124 4164
rect 9151 4152 9225 4168
rect 9078 4146 9112 4148
rect 9077 4130 9124 4146
rect 9151 4130 9164 4152
rect 9179 4130 9209 4152
rect 9236 4130 9237 4146
rect 9252 4130 9265 4290
rect 7496 4122 7531 4130
rect 7496 4096 7497 4122
rect 7504 4096 7531 4122
rect 7439 4078 7469 4092
rect 7496 4088 7531 4096
rect 7533 4122 7574 4130
rect 7533 4096 7548 4122
rect 7555 4096 7574 4122
rect 7638 4118 7700 4130
rect 7712 4118 7787 4130
rect 7845 4118 7920 4130
rect 7932 4118 7963 4130
rect 7969 4118 8004 4130
rect 7638 4116 7800 4118
rect 7533 4088 7574 4096
rect 7656 4092 7669 4116
rect 7684 4114 7699 4116
rect 7496 4078 7525 4088
rect 7539 4078 7568 4088
rect 7583 4078 7613 4092
rect 7656 4078 7699 4092
rect 7723 4089 7730 4096
rect 7733 4092 7800 4116
rect 7832 4116 8004 4118
rect 7802 4094 7830 4098
rect 7832 4094 7912 4116
rect 7933 4114 7948 4116
rect 7802 4092 7912 4094
rect 7733 4088 7912 4092
rect 7706 4078 7736 4088
rect 7738 4078 7891 4088
rect 7899 4078 7929 4088
rect 7933 4078 7963 4092
rect 7991 4078 8004 4116
rect 8076 4122 8111 4130
rect 8076 4096 8077 4122
rect 8084 4096 8111 4122
rect 8019 4078 8049 4092
rect 8076 4088 8111 4096
rect 8113 4122 8154 4130
rect 8113 4096 8128 4122
rect 8135 4096 8154 4122
rect 8218 4118 8280 4130
rect 8292 4118 8367 4130
rect 8425 4118 8500 4130
rect 8512 4118 8543 4130
rect 8549 4118 8584 4130
rect 8218 4116 8380 4118
rect 8113 4088 8154 4096
rect 8236 4092 8249 4116
rect 8264 4114 8279 4116
rect 8076 4078 8077 4088
rect 8092 4078 8105 4088
rect 8119 4078 8120 4088
rect 8135 4078 8148 4088
rect 8163 4078 8193 4092
rect 8236 4078 8279 4092
rect 8303 4089 8310 4096
rect 8313 4092 8380 4116
rect 8412 4116 8584 4118
rect 8382 4094 8410 4098
rect 8412 4094 8492 4116
rect 8513 4114 8528 4116
rect 8382 4092 8492 4094
rect 8313 4088 8492 4092
rect 8286 4078 8316 4088
rect 8318 4078 8471 4088
rect 8479 4078 8509 4088
rect 8513 4078 8543 4092
rect 8571 4078 8584 4116
rect 8656 4122 8691 4130
rect 8656 4096 8657 4122
rect 8664 4096 8691 4122
rect 8599 4078 8629 4092
rect 8656 4088 8691 4096
rect 8693 4122 8734 4130
rect 8693 4096 8708 4122
rect 8715 4096 8734 4122
rect 8798 4118 8860 4130
rect 8872 4118 8947 4130
rect 9005 4118 9080 4130
rect 9092 4118 9123 4130
rect 9129 4118 9164 4130
rect 8798 4116 8960 4118
rect 8693 4088 8734 4096
rect 8816 4092 8829 4116
rect 8844 4114 8859 4116
rect 8656 4078 8657 4088
rect 8672 4078 8685 4088
rect 8699 4078 8700 4088
rect 8715 4078 8728 4088
rect 8743 4078 8773 4092
rect 8816 4078 8859 4092
rect 8883 4089 8890 4096
rect 8893 4092 8960 4116
rect 8992 4116 9164 4118
rect 8962 4094 8990 4098
rect 8992 4094 9072 4116
rect 9093 4114 9108 4116
rect 8962 4092 9072 4094
rect 8893 4088 9072 4092
rect 8866 4078 8896 4088
rect 8898 4078 9051 4088
rect 9059 4078 9089 4088
rect 9093 4078 9123 4092
rect 9151 4078 9164 4116
rect 9236 4122 9271 4130
rect 9236 4096 9237 4122
rect 9244 4096 9271 4122
rect 9179 4078 9209 4092
rect 9236 4088 9271 4096
rect 9236 4078 9237 4088
rect 9252 4078 9265 4088
rect -1 4072 9265 4078
rect 0 4064 9265 4072
rect 15 4034 28 4064
rect 43 4050 73 4064
rect 116 4050 159 4064
rect 166 4050 386 4064
rect 393 4050 423 4064
rect 83 4036 98 4048
rect 117 4036 130 4050
rect 198 4046 351 4050
rect 80 4034 102 4036
rect 180 4034 372 4046
rect 451 4034 464 4064
rect 479 4050 509 4064
rect 546 4034 565 4064
rect 580 4034 586 4064
rect 595 4034 608 4064
rect 623 4050 653 4064
rect 696 4050 739 4064
rect 746 4050 966 4064
rect 973 4050 1003 4064
rect 663 4036 678 4048
rect 697 4036 710 4050
rect 778 4046 931 4050
rect 660 4034 682 4036
rect 760 4034 952 4046
rect 1031 4034 1044 4064
rect 1059 4050 1089 4064
rect 1126 4034 1145 4064
rect 1160 4034 1166 4064
rect 1175 4034 1188 4064
rect 1203 4050 1233 4064
rect 1276 4050 1319 4064
rect 1326 4050 1546 4064
rect 1553 4050 1583 4064
rect 1243 4036 1258 4048
rect 1277 4036 1290 4050
rect 1358 4046 1511 4050
rect 1240 4034 1262 4036
rect 1340 4034 1532 4046
rect 1611 4034 1624 4064
rect 1639 4050 1669 4064
rect 1706 4034 1725 4064
rect 1740 4034 1746 4064
rect 1755 4034 1768 4064
rect 1783 4050 1813 4064
rect 1856 4050 1899 4064
rect 1906 4050 2126 4064
rect 2133 4050 2163 4064
rect 1823 4036 1838 4048
rect 1857 4036 1870 4050
rect 1938 4046 2091 4050
rect 1820 4034 1842 4036
rect 1920 4034 2112 4046
rect 2191 4034 2204 4064
rect 2219 4050 2249 4064
rect 2286 4034 2305 4064
rect 2320 4034 2326 4064
rect 2335 4034 2348 4064
rect 2363 4050 2393 4064
rect 2436 4050 2479 4064
rect 2486 4050 2706 4064
rect 2713 4050 2743 4064
rect 2403 4036 2418 4048
rect 2437 4036 2450 4050
rect 2518 4046 2671 4050
rect 2400 4034 2422 4036
rect 2500 4034 2692 4046
rect 2771 4034 2784 4064
rect 2799 4050 2829 4064
rect 2866 4034 2885 4064
rect 2900 4034 2906 4064
rect 2915 4034 2928 4064
rect 2943 4050 2973 4064
rect 3016 4050 3059 4064
rect 3066 4050 3286 4064
rect 3293 4050 3323 4064
rect 2983 4036 2998 4048
rect 3017 4036 3030 4050
rect 3098 4046 3251 4050
rect 2980 4034 3002 4036
rect 3080 4034 3272 4046
rect 3351 4034 3364 4064
rect 3379 4050 3409 4064
rect 3446 4034 3465 4064
rect 3480 4034 3486 4064
rect 3495 4034 3508 4064
rect 3523 4050 3553 4064
rect 3596 4050 3639 4064
rect 3646 4050 3866 4064
rect 3873 4050 3903 4064
rect 3563 4036 3578 4048
rect 3597 4036 3610 4050
rect 3678 4046 3831 4050
rect 3560 4034 3582 4036
rect 3660 4034 3852 4046
rect 3931 4034 3944 4064
rect 3959 4050 3989 4064
rect 4026 4034 4045 4064
rect 4060 4034 4066 4064
rect 4075 4034 4088 4064
rect 4103 4050 4133 4064
rect 4176 4050 4219 4064
rect 4226 4050 4446 4064
rect 4453 4050 4483 4064
rect 4143 4036 4158 4048
rect 4177 4036 4190 4050
rect 4258 4046 4411 4050
rect 4140 4034 4162 4036
rect 4240 4034 4432 4046
rect 4511 4034 4524 4064
rect 4539 4050 4569 4064
rect 4606 4034 4625 4064
rect 4640 4034 4646 4064
rect 4655 4034 4668 4064
rect 4683 4050 4713 4064
rect 4756 4050 4799 4064
rect 4806 4050 5026 4064
rect 5033 4050 5063 4064
rect 4723 4036 4738 4048
rect 4757 4036 4770 4050
rect 4838 4046 4991 4050
rect 4720 4034 4742 4036
rect 4820 4034 5012 4046
rect 5091 4034 5104 4064
rect 5119 4050 5149 4064
rect 5186 4034 5205 4064
rect 5220 4034 5226 4064
rect 5235 4034 5248 4064
rect 5263 4050 5293 4064
rect 5336 4050 5379 4064
rect 5386 4050 5606 4064
rect 5613 4050 5643 4064
rect 5303 4036 5318 4048
rect 5337 4036 5350 4050
rect 5418 4046 5571 4050
rect 5300 4034 5322 4036
rect 5400 4034 5592 4046
rect 5671 4034 5684 4064
rect 5699 4050 5729 4064
rect 5766 4034 5785 4064
rect 5800 4034 5806 4064
rect 5815 4034 5828 4064
rect 5843 4050 5873 4064
rect 5916 4050 5959 4064
rect 5966 4050 6186 4064
rect 6193 4050 6223 4064
rect 5883 4036 5898 4048
rect 5917 4036 5930 4050
rect 5998 4046 6151 4050
rect 5880 4034 5902 4036
rect 5980 4034 6172 4046
rect 6251 4034 6264 4064
rect 6279 4050 6309 4064
rect 6346 4034 6365 4064
rect 6380 4034 6386 4064
rect 6395 4034 6408 4064
rect 6423 4050 6453 4064
rect 6496 4050 6539 4064
rect 6546 4050 6766 4064
rect 6773 4050 6803 4064
rect 6463 4036 6478 4048
rect 6497 4036 6510 4050
rect 6578 4046 6731 4050
rect 6460 4034 6482 4036
rect 6560 4034 6752 4046
rect 6831 4034 6844 4064
rect 6859 4050 6889 4064
rect 6926 4034 6945 4064
rect 6960 4034 6966 4064
rect 6975 4034 6988 4064
rect 7003 4050 7033 4064
rect 7076 4050 7119 4064
rect 7126 4050 7346 4064
rect 7353 4050 7383 4064
rect 7043 4036 7058 4048
rect 7077 4036 7090 4050
rect 7158 4046 7311 4050
rect 7040 4034 7062 4036
rect 7140 4034 7332 4046
rect 7411 4034 7424 4064
rect 7439 4050 7469 4064
rect 7506 4034 7525 4064
rect 7540 4034 7546 4064
rect 7555 4034 7568 4064
rect 7583 4046 7613 4064
rect 7656 4050 7670 4064
rect 7706 4050 7926 4064
rect 7657 4048 7670 4050
rect 7623 4036 7638 4048
rect 7620 4034 7642 4036
rect 7647 4034 7677 4048
rect 7738 4046 7891 4050
rect 7720 4034 7912 4046
rect 7955 4034 7985 4048
rect 7991 4034 8004 4064
rect 8019 4046 8049 4064
rect 8092 4034 8105 4064
rect 8135 4034 8148 4064
rect 8163 4046 8193 4064
rect 8236 4050 8250 4064
rect 8286 4050 8506 4064
rect 8237 4048 8250 4050
rect 8203 4036 8218 4048
rect 8200 4034 8222 4036
rect 8227 4034 8257 4048
rect 8318 4046 8471 4050
rect 8300 4034 8492 4046
rect 8535 4034 8565 4048
rect 8571 4034 8584 4064
rect 8599 4046 8629 4064
rect 8672 4034 8685 4064
rect 8715 4034 8728 4064
rect 8743 4046 8773 4064
rect 8816 4050 8830 4064
rect 8866 4050 9086 4064
rect 8817 4048 8830 4050
rect 8783 4036 8798 4048
rect 8780 4034 8802 4036
rect 8807 4034 8837 4048
rect 8898 4046 9051 4050
rect 8880 4034 9072 4046
rect 9115 4034 9145 4048
rect 9151 4034 9164 4064
rect 9179 4046 9209 4064
rect 9252 4034 9265 4064
rect 0 4020 9265 4034
rect 15 3950 28 4020
rect 80 4016 102 4020
rect 73 3994 102 4008
rect 155 3994 171 4008
rect 209 4004 215 4006
rect 222 4004 330 4020
rect 337 4004 343 4006
rect 351 4004 366 4020
rect 432 4014 451 4017
rect 73 3992 171 3994
rect 198 3992 366 4004
rect 381 3994 397 4008
rect 432 3995 454 4014
rect 464 4008 480 4009
rect 463 4006 480 4008
rect 464 4001 480 4006
rect 454 3994 460 3995
rect 463 3994 492 4001
rect 381 3993 492 3994
rect 381 3992 498 3993
rect 57 3984 108 3992
rect 155 3984 189 3992
rect 57 3972 82 3984
rect 89 3972 108 3984
rect 162 3982 189 3984
rect 198 3982 419 3992
rect 454 3989 460 3992
rect 162 3978 419 3982
rect 57 3964 108 3972
rect 155 3964 419 3978
rect 463 3984 498 3992
rect 9 3916 28 3950
rect 73 3956 102 3964
rect 73 3950 90 3956
rect 73 3948 107 3950
rect 155 3948 171 3964
rect 172 3954 380 3964
rect 381 3954 397 3964
rect 445 3960 460 3975
rect 463 3972 464 3984
rect 471 3972 498 3984
rect 463 3964 498 3972
rect 463 3963 492 3964
rect 183 3950 397 3954
rect 198 3948 397 3950
rect 432 3950 445 3960
rect 463 3950 480 3963
rect 432 3948 480 3950
rect 74 3944 107 3948
rect 70 3942 107 3944
rect 70 3941 137 3942
rect 70 3936 101 3941
rect 107 3936 137 3941
rect 70 3932 137 3936
rect 43 3929 137 3932
rect 43 3922 92 3929
rect 43 3916 73 3922
rect 92 3917 97 3922
rect 9 3900 89 3916
rect 101 3908 137 3929
rect 198 3924 387 3948
rect 432 3947 479 3948
rect 445 3942 479 3947
rect 213 3921 387 3924
rect 206 3918 387 3921
rect 415 3941 479 3942
rect 9 3898 28 3900
rect 43 3898 77 3900
rect 9 3882 89 3898
rect 9 3876 28 3882
rect -1 3860 28 3876
rect 43 3866 73 3882
rect 101 3860 107 3908
rect 110 3902 129 3908
rect 144 3902 174 3910
rect 110 3894 174 3902
rect 110 3878 190 3894
rect 206 3887 268 3918
rect 284 3887 346 3918
rect 415 3916 464 3941
rect 479 3916 509 3932
rect 378 3902 408 3910
rect 415 3908 525 3916
rect 378 3894 423 3902
rect 110 3876 129 3878
rect 144 3876 190 3878
rect 110 3860 190 3876
rect 217 3874 252 3887
rect 293 3884 330 3887
rect 293 3882 335 3884
rect 222 3871 252 3874
rect 231 3867 238 3871
rect 238 3866 239 3867
rect 197 3860 207 3866
rect -7 3852 34 3860
rect -7 3826 8 3852
rect 15 3826 34 3852
rect 98 3848 129 3860
rect 144 3848 247 3860
rect 259 3850 285 3876
rect 300 3871 330 3882
rect 362 3878 424 3894
rect 362 3876 408 3878
rect 362 3860 424 3876
rect 436 3860 442 3908
rect 445 3900 525 3908
rect 445 3898 464 3900
rect 479 3898 513 3900
rect 445 3882 525 3898
rect 445 3860 464 3882
rect 479 3866 509 3882
rect 537 3876 543 3950
rect 546 3876 565 4020
rect 580 3876 586 4020
rect 595 3950 608 4020
rect 660 4016 682 4020
rect 653 3994 682 4008
rect 735 3994 751 4008
rect 789 4004 795 4006
rect 802 4004 910 4020
rect 917 4004 923 4006
rect 931 4004 946 4020
rect 1012 4014 1031 4017
rect 653 3992 751 3994
rect 778 3992 946 4004
rect 961 3994 977 4008
rect 1012 3995 1034 4014
rect 1044 4008 1060 4009
rect 1043 4006 1060 4008
rect 1044 4001 1060 4006
rect 1034 3994 1040 3995
rect 1043 3994 1072 4001
rect 961 3993 1072 3994
rect 961 3992 1078 3993
rect 637 3984 688 3992
rect 735 3984 769 3992
rect 637 3972 662 3984
rect 669 3972 688 3984
rect 742 3982 769 3984
rect 778 3982 999 3992
rect 1034 3989 1040 3992
rect 742 3978 999 3982
rect 637 3964 688 3972
rect 735 3964 999 3978
rect 1043 3984 1078 3992
rect 589 3916 608 3950
rect 653 3956 682 3964
rect 653 3950 670 3956
rect 653 3948 687 3950
rect 735 3948 751 3964
rect 752 3954 960 3964
rect 961 3954 977 3964
rect 1025 3960 1040 3975
rect 1043 3972 1044 3984
rect 1051 3972 1078 3984
rect 1043 3964 1078 3972
rect 1043 3963 1072 3964
rect 763 3950 977 3954
rect 778 3948 977 3950
rect 1012 3950 1025 3960
rect 1043 3950 1060 3963
rect 1012 3948 1060 3950
rect 654 3944 687 3948
rect 650 3942 687 3944
rect 650 3941 717 3942
rect 650 3936 681 3941
rect 687 3936 717 3941
rect 650 3932 717 3936
rect 623 3929 717 3932
rect 623 3922 672 3929
rect 623 3916 653 3922
rect 672 3917 677 3922
rect 589 3900 669 3916
rect 681 3908 717 3929
rect 778 3924 967 3948
rect 1012 3947 1059 3948
rect 1025 3942 1059 3947
rect 793 3921 967 3924
rect 786 3918 967 3921
rect 995 3941 1059 3942
rect 589 3898 608 3900
rect 623 3898 657 3900
rect 589 3882 669 3898
rect 589 3876 608 3882
rect 305 3850 408 3860
rect 259 3848 408 3850
rect 429 3848 464 3860
rect 98 3846 260 3848
rect 110 3826 129 3846
rect 144 3844 174 3846
rect -7 3818 34 3826
rect 116 3822 129 3826
rect 181 3830 260 3846
rect 292 3846 464 3848
rect 292 3830 371 3846
rect 378 3844 408 3846
rect -1 3808 28 3818
rect 43 3808 73 3822
rect 116 3808 159 3822
rect 181 3818 371 3830
rect 436 3826 442 3846
rect 166 3808 196 3818
rect 197 3808 355 3818
rect 359 3808 389 3818
rect 393 3808 423 3822
rect 451 3808 464 3846
rect 536 3860 565 3876
rect 579 3860 608 3876
rect 623 3866 653 3882
rect 681 3860 687 3908
rect 690 3902 709 3908
rect 724 3902 754 3910
rect 690 3894 754 3902
rect 690 3878 770 3894
rect 786 3887 848 3918
rect 864 3887 926 3918
rect 995 3916 1044 3941
rect 1059 3916 1089 3932
rect 958 3902 988 3910
rect 995 3908 1105 3916
rect 958 3894 1003 3902
rect 690 3876 709 3878
rect 724 3876 770 3878
rect 690 3860 770 3876
rect 797 3874 832 3887
rect 873 3884 910 3887
rect 873 3882 915 3884
rect 802 3871 832 3874
rect 811 3867 818 3871
rect 818 3866 819 3867
rect 777 3860 787 3866
rect 536 3852 571 3860
rect 536 3826 537 3852
rect 544 3826 571 3852
rect 479 3808 509 3822
rect 536 3818 571 3826
rect 573 3852 614 3860
rect 573 3826 588 3852
rect 595 3826 614 3852
rect 678 3848 709 3860
rect 724 3848 827 3860
rect 839 3850 865 3876
rect 880 3871 910 3882
rect 942 3878 1004 3894
rect 942 3876 988 3878
rect 942 3860 1004 3876
rect 1016 3860 1022 3908
rect 1025 3900 1105 3908
rect 1025 3898 1044 3900
rect 1059 3898 1093 3900
rect 1025 3882 1105 3898
rect 1025 3860 1044 3882
rect 1059 3866 1089 3882
rect 1117 3876 1123 3950
rect 1126 3876 1145 4020
rect 1160 3876 1166 4020
rect 1175 3950 1188 4020
rect 1240 4016 1262 4020
rect 1233 3994 1262 4008
rect 1315 3994 1331 4008
rect 1369 4004 1375 4006
rect 1382 4004 1490 4020
rect 1497 4004 1503 4006
rect 1511 4004 1526 4020
rect 1592 4014 1611 4017
rect 1233 3992 1331 3994
rect 1358 3992 1526 4004
rect 1541 3994 1557 4008
rect 1592 3995 1614 4014
rect 1624 4008 1640 4009
rect 1623 4006 1640 4008
rect 1624 4001 1640 4006
rect 1614 3994 1620 3995
rect 1623 3994 1652 4001
rect 1541 3993 1652 3994
rect 1541 3992 1658 3993
rect 1217 3984 1268 3992
rect 1315 3984 1349 3992
rect 1217 3972 1242 3984
rect 1249 3972 1268 3984
rect 1322 3982 1349 3984
rect 1358 3982 1579 3992
rect 1614 3989 1620 3992
rect 1322 3978 1579 3982
rect 1217 3964 1268 3972
rect 1315 3964 1579 3978
rect 1623 3984 1658 3992
rect 1169 3916 1188 3950
rect 1233 3956 1262 3964
rect 1233 3950 1250 3956
rect 1233 3948 1267 3950
rect 1315 3948 1331 3964
rect 1332 3954 1540 3964
rect 1541 3954 1557 3964
rect 1605 3960 1620 3975
rect 1623 3972 1624 3984
rect 1631 3972 1658 3984
rect 1623 3964 1658 3972
rect 1623 3963 1652 3964
rect 1343 3950 1557 3954
rect 1358 3948 1557 3950
rect 1592 3950 1605 3960
rect 1623 3950 1640 3963
rect 1592 3948 1640 3950
rect 1234 3944 1267 3948
rect 1230 3942 1267 3944
rect 1230 3941 1297 3942
rect 1230 3936 1261 3941
rect 1267 3936 1297 3941
rect 1230 3932 1297 3936
rect 1203 3929 1297 3932
rect 1203 3922 1252 3929
rect 1203 3916 1233 3922
rect 1252 3917 1257 3922
rect 1169 3900 1249 3916
rect 1261 3908 1297 3929
rect 1358 3924 1547 3948
rect 1592 3947 1639 3948
rect 1605 3942 1639 3947
rect 1373 3921 1547 3924
rect 1366 3918 1547 3921
rect 1575 3941 1639 3942
rect 1169 3898 1188 3900
rect 1203 3898 1237 3900
rect 1169 3882 1249 3898
rect 1169 3876 1188 3882
rect 885 3850 988 3860
rect 839 3848 988 3850
rect 1009 3848 1044 3860
rect 678 3846 840 3848
rect 690 3826 709 3846
rect 724 3844 754 3846
rect 573 3818 614 3826
rect 696 3822 709 3826
rect 761 3830 840 3846
rect 872 3846 1044 3848
rect 872 3830 951 3846
rect 958 3844 988 3846
rect 536 3808 565 3818
rect 579 3808 608 3818
rect 623 3808 653 3822
rect 696 3808 739 3822
rect 761 3818 951 3830
rect 1016 3826 1022 3846
rect 746 3808 776 3818
rect 777 3808 935 3818
rect 939 3808 969 3818
rect 973 3808 1003 3822
rect 1031 3808 1044 3846
rect 1116 3860 1145 3876
rect 1159 3860 1188 3876
rect 1203 3866 1233 3882
rect 1261 3860 1267 3908
rect 1270 3902 1289 3908
rect 1304 3902 1334 3910
rect 1270 3894 1334 3902
rect 1270 3878 1350 3894
rect 1366 3887 1428 3918
rect 1444 3887 1506 3918
rect 1575 3916 1624 3941
rect 1639 3916 1669 3932
rect 1538 3902 1568 3910
rect 1575 3908 1685 3916
rect 1538 3894 1583 3902
rect 1270 3876 1289 3878
rect 1304 3876 1350 3878
rect 1270 3860 1350 3876
rect 1377 3874 1412 3887
rect 1453 3884 1490 3887
rect 1453 3882 1495 3884
rect 1382 3871 1412 3874
rect 1391 3867 1398 3871
rect 1398 3866 1399 3867
rect 1357 3860 1367 3866
rect 1116 3852 1151 3860
rect 1116 3826 1117 3852
rect 1124 3826 1151 3852
rect 1059 3808 1089 3822
rect 1116 3818 1151 3826
rect 1153 3852 1194 3860
rect 1153 3826 1168 3852
rect 1175 3826 1194 3852
rect 1258 3848 1289 3860
rect 1304 3848 1407 3860
rect 1419 3850 1445 3876
rect 1460 3871 1490 3882
rect 1522 3878 1584 3894
rect 1522 3876 1568 3878
rect 1522 3860 1584 3876
rect 1596 3860 1602 3908
rect 1605 3900 1685 3908
rect 1605 3898 1624 3900
rect 1639 3898 1673 3900
rect 1605 3882 1685 3898
rect 1605 3860 1624 3882
rect 1639 3866 1669 3882
rect 1697 3876 1703 3950
rect 1706 3876 1725 4020
rect 1740 3876 1746 4020
rect 1755 3950 1768 4020
rect 1820 4016 1842 4020
rect 1813 3994 1842 4008
rect 1895 3994 1911 4008
rect 1949 4004 1955 4006
rect 1962 4004 2070 4020
rect 2077 4004 2083 4006
rect 2091 4004 2106 4020
rect 2172 4014 2191 4017
rect 1813 3992 1911 3994
rect 1938 3992 2106 4004
rect 2121 3994 2137 4008
rect 2172 3995 2194 4014
rect 2204 4008 2220 4009
rect 2203 4006 2220 4008
rect 2204 4001 2220 4006
rect 2194 3994 2200 3995
rect 2203 3994 2232 4001
rect 2121 3993 2232 3994
rect 2121 3992 2238 3993
rect 1797 3984 1848 3992
rect 1895 3984 1929 3992
rect 1797 3972 1822 3984
rect 1829 3972 1848 3984
rect 1902 3982 1929 3984
rect 1938 3982 2159 3992
rect 2194 3989 2200 3992
rect 1902 3978 2159 3982
rect 1797 3964 1848 3972
rect 1895 3964 2159 3978
rect 2203 3984 2238 3992
rect 1749 3916 1768 3950
rect 1813 3956 1842 3964
rect 1813 3950 1830 3956
rect 1813 3948 1847 3950
rect 1895 3948 1911 3964
rect 1912 3954 2120 3964
rect 2121 3954 2137 3964
rect 2185 3960 2200 3975
rect 2203 3972 2204 3984
rect 2211 3972 2238 3984
rect 2203 3964 2238 3972
rect 2203 3963 2232 3964
rect 1923 3950 2137 3954
rect 1938 3948 2137 3950
rect 2172 3950 2185 3960
rect 2203 3950 2220 3963
rect 2172 3948 2220 3950
rect 1814 3944 1847 3948
rect 1810 3942 1847 3944
rect 1810 3941 1877 3942
rect 1810 3936 1841 3941
rect 1847 3936 1877 3941
rect 1810 3932 1877 3936
rect 1783 3929 1877 3932
rect 1783 3922 1832 3929
rect 1783 3916 1813 3922
rect 1832 3917 1837 3922
rect 1749 3900 1829 3916
rect 1841 3908 1877 3929
rect 1938 3924 2127 3948
rect 2172 3947 2219 3948
rect 2185 3942 2219 3947
rect 1953 3921 2127 3924
rect 1946 3918 2127 3921
rect 2155 3941 2219 3942
rect 1749 3898 1768 3900
rect 1783 3898 1817 3900
rect 1749 3882 1829 3898
rect 1749 3876 1768 3882
rect 1465 3850 1568 3860
rect 1419 3848 1568 3850
rect 1589 3848 1624 3860
rect 1258 3846 1420 3848
rect 1270 3826 1289 3846
rect 1304 3844 1334 3846
rect 1153 3818 1194 3826
rect 1276 3822 1289 3826
rect 1341 3830 1420 3846
rect 1452 3846 1624 3848
rect 1452 3830 1531 3846
rect 1538 3844 1568 3846
rect 1116 3808 1145 3818
rect 1159 3808 1188 3818
rect 1203 3808 1233 3822
rect 1276 3808 1319 3822
rect 1341 3818 1531 3830
rect 1596 3826 1602 3846
rect 1326 3808 1356 3818
rect 1357 3808 1515 3818
rect 1519 3808 1549 3818
rect 1553 3808 1583 3822
rect 1611 3808 1624 3846
rect 1696 3860 1725 3876
rect 1739 3860 1768 3876
rect 1783 3866 1813 3882
rect 1841 3860 1847 3908
rect 1850 3902 1869 3908
rect 1884 3902 1914 3910
rect 1850 3894 1914 3902
rect 1850 3878 1930 3894
rect 1946 3887 2008 3918
rect 2024 3887 2086 3918
rect 2155 3916 2204 3941
rect 2219 3916 2249 3932
rect 2118 3902 2148 3910
rect 2155 3908 2265 3916
rect 2118 3894 2163 3902
rect 1850 3876 1869 3878
rect 1884 3876 1930 3878
rect 1850 3860 1930 3876
rect 1957 3874 1992 3887
rect 2033 3884 2070 3887
rect 2033 3882 2075 3884
rect 1962 3871 1992 3874
rect 1971 3867 1978 3871
rect 1978 3866 1979 3867
rect 1937 3860 1947 3866
rect 1696 3852 1731 3860
rect 1696 3826 1697 3852
rect 1704 3826 1731 3852
rect 1639 3808 1669 3822
rect 1696 3818 1731 3826
rect 1733 3852 1774 3860
rect 1733 3826 1748 3852
rect 1755 3826 1774 3852
rect 1838 3848 1869 3860
rect 1884 3848 1987 3860
rect 1999 3850 2025 3876
rect 2040 3871 2070 3882
rect 2102 3878 2164 3894
rect 2102 3876 2148 3878
rect 2102 3860 2164 3876
rect 2176 3860 2182 3908
rect 2185 3900 2265 3908
rect 2185 3898 2204 3900
rect 2219 3898 2253 3900
rect 2185 3882 2265 3898
rect 2185 3860 2204 3882
rect 2219 3866 2249 3882
rect 2277 3876 2283 3950
rect 2286 3876 2305 4020
rect 2320 3876 2326 4020
rect 2335 3950 2348 4020
rect 2400 4016 2422 4020
rect 2393 3994 2422 4008
rect 2475 3994 2491 4008
rect 2529 4004 2535 4006
rect 2542 4004 2650 4020
rect 2657 4004 2663 4006
rect 2671 4004 2686 4020
rect 2752 4014 2771 4017
rect 2393 3992 2491 3994
rect 2518 3992 2686 4004
rect 2701 3994 2717 4008
rect 2752 3995 2774 4014
rect 2784 4008 2800 4009
rect 2783 4006 2800 4008
rect 2784 4001 2800 4006
rect 2774 3994 2780 3995
rect 2783 3994 2812 4001
rect 2701 3993 2812 3994
rect 2701 3992 2818 3993
rect 2377 3984 2428 3992
rect 2475 3984 2509 3992
rect 2377 3972 2402 3984
rect 2409 3972 2428 3984
rect 2482 3982 2509 3984
rect 2518 3982 2739 3992
rect 2774 3989 2780 3992
rect 2482 3978 2739 3982
rect 2377 3964 2428 3972
rect 2475 3964 2739 3978
rect 2783 3984 2818 3992
rect 2329 3916 2348 3950
rect 2393 3956 2422 3964
rect 2393 3950 2410 3956
rect 2393 3948 2427 3950
rect 2475 3948 2491 3964
rect 2492 3954 2700 3964
rect 2701 3954 2717 3964
rect 2765 3960 2780 3975
rect 2783 3972 2784 3984
rect 2791 3972 2818 3984
rect 2783 3964 2818 3972
rect 2783 3963 2812 3964
rect 2503 3950 2717 3954
rect 2518 3948 2717 3950
rect 2752 3950 2765 3960
rect 2783 3950 2800 3963
rect 2752 3948 2800 3950
rect 2394 3944 2427 3948
rect 2390 3942 2427 3944
rect 2390 3941 2457 3942
rect 2390 3936 2421 3941
rect 2427 3936 2457 3941
rect 2390 3932 2457 3936
rect 2363 3929 2457 3932
rect 2363 3922 2412 3929
rect 2363 3916 2393 3922
rect 2412 3917 2417 3922
rect 2329 3900 2409 3916
rect 2421 3908 2457 3929
rect 2518 3924 2707 3948
rect 2752 3947 2799 3948
rect 2765 3942 2799 3947
rect 2533 3921 2707 3924
rect 2526 3918 2707 3921
rect 2735 3941 2799 3942
rect 2329 3898 2348 3900
rect 2363 3898 2397 3900
rect 2329 3882 2409 3898
rect 2329 3876 2348 3882
rect 2045 3850 2148 3860
rect 1999 3848 2148 3850
rect 2169 3848 2204 3860
rect 1838 3846 2000 3848
rect 1850 3826 1869 3846
rect 1884 3844 1914 3846
rect 1733 3818 1774 3826
rect 1856 3822 1869 3826
rect 1921 3830 2000 3846
rect 2032 3846 2204 3848
rect 2032 3830 2111 3846
rect 2118 3844 2148 3846
rect 1696 3808 1725 3818
rect 1739 3808 1768 3818
rect 1783 3808 1813 3822
rect 1856 3808 1899 3822
rect 1921 3818 2111 3830
rect 2176 3826 2182 3846
rect 1906 3808 1936 3818
rect 1937 3808 2095 3818
rect 2099 3808 2129 3818
rect 2133 3808 2163 3822
rect 2191 3808 2204 3846
rect 2276 3860 2305 3876
rect 2319 3860 2348 3876
rect 2363 3866 2393 3882
rect 2421 3860 2427 3908
rect 2430 3902 2449 3908
rect 2464 3902 2494 3910
rect 2430 3894 2494 3902
rect 2430 3878 2510 3894
rect 2526 3887 2588 3918
rect 2604 3887 2666 3918
rect 2735 3916 2784 3941
rect 2799 3916 2829 3932
rect 2698 3902 2728 3910
rect 2735 3908 2845 3916
rect 2698 3894 2743 3902
rect 2430 3876 2449 3878
rect 2464 3876 2510 3878
rect 2430 3860 2510 3876
rect 2537 3874 2572 3887
rect 2613 3884 2650 3887
rect 2613 3882 2655 3884
rect 2542 3871 2572 3874
rect 2551 3867 2558 3871
rect 2558 3866 2559 3867
rect 2517 3860 2527 3866
rect 2276 3852 2311 3860
rect 2276 3826 2277 3852
rect 2284 3826 2311 3852
rect 2219 3808 2249 3822
rect 2276 3818 2311 3826
rect 2313 3852 2354 3860
rect 2313 3826 2328 3852
rect 2335 3826 2354 3852
rect 2418 3848 2449 3860
rect 2464 3848 2567 3860
rect 2579 3850 2605 3876
rect 2620 3871 2650 3882
rect 2682 3878 2744 3894
rect 2682 3876 2728 3878
rect 2682 3860 2744 3876
rect 2756 3860 2762 3908
rect 2765 3900 2845 3908
rect 2765 3898 2784 3900
rect 2799 3898 2833 3900
rect 2765 3882 2845 3898
rect 2765 3860 2784 3882
rect 2799 3866 2829 3882
rect 2857 3876 2863 3950
rect 2866 3876 2885 4020
rect 2900 3876 2906 4020
rect 2915 3950 2928 4020
rect 2980 4016 3002 4020
rect 2973 3994 3002 4008
rect 3055 3994 3071 4008
rect 3109 4004 3115 4006
rect 3122 4004 3230 4020
rect 3237 4004 3243 4006
rect 3251 4004 3266 4020
rect 3332 4014 3351 4017
rect 2973 3992 3071 3994
rect 3098 3992 3266 4004
rect 3281 3994 3297 4008
rect 3332 3995 3354 4014
rect 3364 4008 3380 4009
rect 3363 4006 3380 4008
rect 3364 4001 3380 4006
rect 3354 3994 3360 3995
rect 3363 3994 3392 4001
rect 3281 3993 3392 3994
rect 3281 3992 3398 3993
rect 2957 3984 3008 3992
rect 3055 3984 3089 3992
rect 2957 3972 2982 3984
rect 2989 3972 3008 3984
rect 3062 3982 3089 3984
rect 3098 3982 3319 3992
rect 3354 3989 3360 3992
rect 3062 3978 3319 3982
rect 2957 3964 3008 3972
rect 3055 3964 3319 3978
rect 3363 3984 3398 3992
rect 2909 3916 2928 3950
rect 2973 3956 3002 3964
rect 2973 3950 2990 3956
rect 2973 3948 3007 3950
rect 3055 3948 3071 3964
rect 3072 3954 3280 3964
rect 3281 3954 3297 3964
rect 3345 3960 3360 3975
rect 3363 3972 3364 3984
rect 3371 3972 3398 3984
rect 3363 3964 3398 3972
rect 3363 3963 3392 3964
rect 3083 3950 3297 3954
rect 3098 3948 3297 3950
rect 3332 3950 3345 3960
rect 3363 3950 3380 3963
rect 3332 3948 3380 3950
rect 2974 3944 3007 3948
rect 2970 3942 3007 3944
rect 2970 3941 3037 3942
rect 2970 3936 3001 3941
rect 3007 3936 3037 3941
rect 2970 3932 3037 3936
rect 2943 3929 3037 3932
rect 2943 3922 2992 3929
rect 2943 3916 2973 3922
rect 2992 3917 2997 3922
rect 2909 3900 2989 3916
rect 3001 3908 3037 3929
rect 3098 3924 3287 3948
rect 3332 3947 3379 3948
rect 3345 3942 3379 3947
rect 3113 3921 3287 3924
rect 3106 3918 3287 3921
rect 3315 3941 3379 3942
rect 2909 3898 2928 3900
rect 2943 3898 2977 3900
rect 2909 3882 2989 3898
rect 2909 3876 2928 3882
rect 2625 3850 2728 3860
rect 2579 3848 2728 3850
rect 2749 3848 2784 3860
rect 2418 3846 2580 3848
rect 2430 3826 2449 3846
rect 2464 3844 2494 3846
rect 2313 3818 2354 3826
rect 2436 3822 2449 3826
rect 2501 3830 2580 3846
rect 2612 3846 2784 3848
rect 2612 3830 2691 3846
rect 2698 3844 2728 3846
rect 2276 3808 2305 3818
rect 2319 3808 2348 3818
rect 2363 3808 2393 3822
rect 2436 3808 2479 3822
rect 2501 3818 2691 3830
rect 2756 3826 2762 3846
rect 2486 3808 2516 3818
rect 2517 3808 2675 3818
rect 2679 3808 2709 3818
rect 2713 3808 2743 3822
rect 2771 3808 2784 3846
rect 2856 3860 2885 3876
rect 2899 3860 2928 3876
rect 2943 3866 2973 3882
rect 3001 3860 3007 3908
rect 3010 3902 3029 3908
rect 3044 3902 3074 3910
rect 3010 3894 3074 3902
rect 3010 3878 3090 3894
rect 3106 3887 3168 3918
rect 3184 3887 3246 3918
rect 3315 3916 3364 3941
rect 3379 3916 3409 3932
rect 3278 3902 3308 3910
rect 3315 3908 3425 3916
rect 3278 3894 3323 3902
rect 3010 3876 3029 3878
rect 3044 3876 3090 3878
rect 3010 3860 3090 3876
rect 3117 3874 3152 3887
rect 3193 3884 3230 3887
rect 3193 3882 3235 3884
rect 3122 3871 3152 3874
rect 3131 3867 3138 3871
rect 3138 3866 3139 3867
rect 3097 3860 3107 3866
rect 2856 3852 2891 3860
rect 2856 3826 2857 3852
rect 2864 3826 2891 3852
rect 2799 3808 2829 3822
rect 2856 3818 2891 3826
rect 2893 3852 2934 3860
rect 2893 3826 2908 3852
rect 2915 3826 2934 3852
rect 2998 3848 3029 3860
rect 3044 3848 3147 3860
rect 3159 3850 3185 3876
rect 3200 3871 3230 3882
rect 3262 3878 3324 3894
rect 3262 3876 3308 3878
rect 3262 3860 3324 3876
rect 3336 3860 3342 3908
rect 3345 3900 3425 3908
rect 3345 3898 3364 3900
rect 3379 3898 3413 3900
rect 3345 3882 3425 3898
rect 3345 3860 3364 3882
rect 3379 3866 3409 3882
rect 3437 3876 3443 3950
rect 3446 3876 3465 4020
rect 3480 3876 3486 4020
rect 3495 3950 3508 4020
rect 3560 4016 3582 4020
rect 3553 3994 3582 4008
rect 3635 3994 3651 4008
rect 3689 4004 3695 4006
rect 3702 4004 3810 4020
rect 3817 4004 3823 4006
rect 3831 4004 3846 4020
rect 3912 4014 3931 4017
rect 3553 3992 3651 3994
rect 3678 3992 3846 4004
rect 3861 3994 3877 4008
rect 3912 3995 3934 4014
rect 3944 4008 3960 4009
rect 3943 4006 3960 4008
rect 3944 4001 3960 4006
rect 3934 3994 3940 3995
rect 3943 3994 3972 4001
rect 3861 3993 3972 3994
rect 3861 3992 3978 3993
rect 3537 3984 3588 3992
rect 3635 3984 3669 3992
rect 3537 3972 3562 3984
rect 3569 3972 3588 3984
rect 3642 3982 3669 3984
rect 3678 3982 3899 3992
rect 3934 3989 3940 3992
rect 3642 3978 3899 3982
rect 3537 3964 3588 3972
rect 3635 3964 3899 3978
rect 3943 3984 3978 3992
rect 3489 3916 3508 3950
rect 3553 3956 3582 3964
rect 3553 3950 3570 3956
rect 3553 3948 3587 3950
rect 3635 3948 3651 3964
rect 3652 3954 3860 3964
rect 3861 3954 3877 3964
rect 3925 3960 3940 3975
rect 3943 3972 3944 3984
rect 3951 3972 3978 3984
rect 3943 3964 3978 3972
rect 3943 3963 3972 3964
rect 3663 3950 3877 3954
rect 3678 3948 3877 3950
rect 3912 3950 3925 3960
rect 3943 3950 3960 3963
rect 3912 3948 3960 3950
rect 3554 3944 3587 3948
rect 3550 3942 3587 3944
rect 3550 3941 3617 3942
rect 3550 3936 3581 3941
rect 3587 3936 3617 3941
rect 3550 3932 3617 3936
rect 3523 3929 3617 3932
rect 3523 3922 3572 3929
rect 3523 3916 3553 3922
rect 3572 3917 3577 3922
rect 3489 3900 3569 3916
rect 3581 3908 3617 3929
rect 3678 3924 3867 3948
rect 3912 3947 3959 3948
rect 3925 3942 3959 3947
rect 3693 3921 3867 3924
rect 3686 3918 3867 3921
rect 3895 3941 3959 3942
rect 3489 3898 3508 3900
rect 3523 3898 3557 3900
rect 3489 3882 3569 3898
rect 3489 3876 3508 3882
rect 3205 3850 3308 3860
rect 3159 3848 3308 3850
rect 3329 3848 3364 3860
rect 2998 3846 3160 3848
rect 3010 3826 3029 3846
rect 3044 3844 3074 3846
rect 2893 3818 2934 3826
rect 3016 3822 3029 3826
rect 3081 3830 3160 3846
rect 3192 3846 3364 3848
rect 3192 3830 3271 3846
rect 3278 3844 3308 3846
rect 2856 3808 2885 3818
rect 2899 3808 2928 3818
rect 2943 3808 2973 3822
rect 3016 3808 3059 3822
rect 3081 3818 3271 3830
rect 3336 3826 3342 3846
rect 3066 3808 3096 3818
rect 3097 3808 3255 3818
rect 3259 3808 3289 3818
rect 3293 3808 3323 3822
rect 3351 3808 3364 3846
rect 3436 3860 3465 3876
rect 3479 3860 3508 3876
rect 3523 3866 3553 3882
rect 3581 3860 3587 3908
rect 3590 3902 3609 3908
rect 3624 3902 3654 3910
rect 3590 3894 3654 3902
rect 3590 3878 3670 3894
rect 3686 3887 3748 3918
rect 3764 3887 3826 3918
rect 3895 3916 3944 3941
rect 3959 3916 3989 3932
rect 3858 3902 3888 3910
rect 3895 3908 4005 3916
rect 3858 3894 3903 3902
rect 3590 3876 3609 3878
rect 3624 3876 3670 3878
rect 3590 3860 3670 3876
rect 3697 3874 3732 3887
rect 3773 3884 3810 3887
rect 3773 3882 3815 3884
rect 3702 3871 3732 3874
rect 3711 3867 3718 3871
rect 3718 3866 3719 3867
rect 3677 3860 3687 3866
rect 3436 3852 3471 3860
rect 3436 3826 3437 3852
rect 3444 3826 3471 3852
rect 3379 3808 3409 3822
rect 3436 3818 3471 3826
rect 3473 3852 3514 3860
rect 3473 3826 3488 3852
rect 3495 3826 3514 3852
rect 3578 3848 3609 3860
rect 3624 3848 3727 3860
rect 3739 3850 3765 3876
rect 3780 3871 3810 3882
rect 3842 3878 3904 3894
rect 3842 3876 3888 3878
rect 3842 3860 3904 3876
rect 3916 3860 3922 3908
rect 3925 3900 4005 3908
rect 3925 3898 3944 3900
rect 3959 3898 3993 3900
rect 3925 3882 4005 3898
rect 3925 3860 3944 3882
rect 3959 3866 3989 3882
rect 4017 3876 4023 3950
rect 4026 3876 4045 4020
rect 4060 3876 4066 4020
rect 4075 3950 4088 4020
rect 4140 4016 4162 4020
rect 4133 3994 4162 4008
rect 4215 3994 4231 4008
rect 4269 4004 4275 4006
rect 4282 4004 4390 4020
rect 4397 4004 4403 4006
rect 4411 4004 4426 4020
rect 4492 4014 4511 4017
rect 4133 3992 4231 3994
rect 4258 3992 4426 4004
rect 4441 3994 4457 4008
rect 4492 3995 4514 4014
rect 4524 4008 4540 4009
rect 4523 4006 4540 4008
rect 4524 4001 4540 4006
rect 4514 3994 4520 3995
rect 4523 3994 4552 4001
rect 4441 3993 4552 3994
rect 4441 3992 4558 3993
rect 4117 3984 4168 3992
rect 4215 3984 4249 3992
rect 4117 3972 4142 3984
rect 4149 3972 4168 3984
rect 4222 3982 4249 3984
rect 4258 3982 4479 3992
rect 4514 3989 4520 3992
rect 4222 3978 4479 3982
rect 4117 3964 4168 3972
rect 4215 3964 4479 3978
rect 4523 3984 4558 3992
rect 4069 3916 4088 3950
rect 4133 3956 4162 3964
rect 4133 3950 4150 3956
rect 4133 3948 4167 3950
rect 4215 3948 4231 3964
rect 4232 3954 4440 3964
rect 4441 3954 4457 3964
rect 4505 3960 4520 3975
rect 4523 3972 4524 3984
rect 4531 3972 4558 3984
rect 4523 3964 4558 3972
rect 4523 3963 4552 3964
rect 4243 3950 4457 3954
rect 4258 3948 4457 3950
rect 4492 3950 4505 3960
rect 4523 3950 4540 3963
rect 4492 3948 4540 3950
rect 4134 3944 4167 3948
rect 4130 3942 4167 3944
rect 4130 3941 4197 3942
rect 4130 3936 4161 3941
rect 4167 3936 4197 3941
rect 4130 3932 4197 3936
rect 4103 3929 4197 3932
rect 4103 3922 4152 3929
rect 4103 3916 4133 3922
rect 4152 3917 4157 3922
rect 4069 3900 4149 3916
rect 4161 3908 4197 3929
rect 4258 3924 4447 3948
rect 4492 3947 4539 3948
rect 4505 3942 4539 3947
rect 4273 3921 4447 3924
rect 4266 3918 4447 3921
rect 4475 3941 4539 3942
rect 4069 3898 4088 3900
rect 4103 3898 4137 3900
rect 4069 3882 4149 3898
rect 4069 3876 4088 3882
rect 3785 3850 3888 3860
rect 3739 3848 3888 3850
rect 3909 3848 3944 3860
rect 3578 3846 3740 3848
rect 3590 3826 3609 3846
rect 3624 3844 3654 3846
rect 3473 3818 3514 3826
rect 3596 3822 3609 3826
rect 3661 3830 3740 3846
rect 3772 3846 3944 3848
rect 3772 3830 3851 3846
rect 3858 3844 3888 3846
rect 3436 3808 3465 3818
rect 3479 3808 3508 3818
rect 3523 3808 3553 3822
rect 3596 3808 3639 3822
rect 3661 3818 3851 3830
rect 3916 3826 3922 3846
rect 3646 3808 3676 3818
rect 3677 3808 3835 3818
rect 3839 3808 3869 3818
rect 3873 3808 3903 3822
rect 3931 3808 3944 3846
rect 4016 3860 4045 3876
rect 4059 3860 4088 3876
rect 4103 3866 4133 3882
rect 4161 3860 4167 3908
rect 4170 3902 4189 3908
rect 4204 3902 4234 3910
rect 4170 3894 4234 3902
rect 4170 3878 4250 3894
rect 4266 3887 4328 3918
rect 4344 3887 4406 3918
rect 4475 3916 4524 3941
rect 4539 3916 4569 3932
rect 4438 3902 4468 3910
rect 4475 3908 4585 3916
rect 4438 3894 4483 3902
rect 4170 3876 4189 3878
rect 4204 3876 4250 3878
rect 4170 3860 4250 3876
rect 4277 3874 4312 3887
rect 4353 3884 4390 3887
rect 4353 3882 4395 3884
rect 4282 3871 4312 3874
rect 4291 3867 4298 3871
rect 4298 3866 4299 3867
rect 4257 3860 4267 3866
rect 4016 3852 4051 3860
rect 4016 3826 4017 3852
rect 4024 3826 4051 3852
rect 3959 3808 3989 3822
rect 4016 3818 4051 3826
rect 4053 3852 4094 3860
rect 4053 3826 4068 3852
rect 4075 3826 4094 3852
rect 4158 3848 4189 3860
rect 4204 3848 4307 3860
rect 4319 3850 4345 3876
rect 4360 3871 4390 3882
rect 4422 3878 4484 3894
rect 4422 3876 4468 3878
rect 4422 3860 4484 3876
rect 4496 3860 4502 3908
rect 4505 3900 4585 3908
rect 4505 3898 4524 3900
rect 4539 3898 4573 3900
rect 4505 3882 4585 3898
rect 4505 3860 4524 3882
rect 4539 3866 4569 3882
rect 4597 3876 4603 3950
rect 4606 3876 4625 4020
rect 4640 3876 4646 4020
rect 4655 3950 4668 4020
rect 4720 4016 4742 4020
rect 4713 3994 4742 4008
rect 4795 3994 4811 4008
rect 4849 4004 4855 4006
rect 4862 4004 4970 4020
rect 4977 4004 4983 4006
rect 4991 4004 5006 4020
rect 5072 4014 5091 4017
rect 4713 3992 4811 3994
rect 4838 3992 5006 4004
rect 5021 3994 5037 4008
rect 5072 3995 5094 4014
rect 5104 4008 5120 4009
rect 5103 4006 5120 4008
rect 5104 4001 5120 4006
rect 5094 3994 5100 3995
rect 5103 3994 5132 4001
rect 5021 3993 5132 3994
rect 5021 3992 5138 3993
rect 4697 3984 4748 3992
rect 4795 3984 4829 3992
rect 4697 3972 4722 3984
rect 4729 3972 4748 3984
rect 4802 3982 4829 3984
rect 4838 3982 5059 3992
rect 5094 3989 5100 3992
rect 4802 3978 5059 3982
rect 4697 3964 4748 3972
rect 4795 3964 5059 3978
rect 5103 3984 5138 3992
rect 4649 3916 4668 3950
rect 4713 3956 4742 3964
rect 4713 3950 4730 3956
rect 4713 3948 4747 3950
rect 4795 3948 4811 3964
rect 4812 3954 5020 3964
rect 5021 3954 5037 3964
rect 5085 3960 5100 3975
rect 5103 3972 5104 3984
rect 5111 3972 5138 3984
rect 5103 3964 5138 3972
rect 5103 3963 5132 3964
rect 4823 3950 5037 3954
rect 4838 3948 5037 3950
rect 5072 3950 5085 3960
rect 5103 3950 5120 3963
rect 5072 3948 5120 3950
rect 4714 3944 4747 3948
rect 4710 3942 4747 3944
rect 4710 3941 4777 3942
rect 4710 3936 4741 3941
rect 4747 3936 4777 3941
rect 4710 3932 4777 3936
rect 4683 3929 4777 3932
rect 4683 3922 4732 3929
rect 4683 3916 4713 3922
rect 4732 3917 4737 3922
rect 4649 3900 4729 3916
rect 4741 3908 4777 3929
rect 4838 3924 5027 3948
rect 5072 3947 5119 3948
rect 5085 3942 5119 3947
rect 4853 3921 5027 3924
rect 4846 3918 5027 3921
rect 5055 3941 5119 3942
rect 4649 3898 4668 3900
rect 4683 3898 4717 3900
rect 4649 3882 4729 3898
rect 4649 3876 4668 3882
rect 4365 3850 4468 3860
rect 4319 3848 4468 3850
rect 4489 3848 4524 3860
rect 4158 3846 4320 3848
rect 4170 3826 4189 3846
rect 4204 3844 4234 3846
rect 4053 3818 4094 3826
rect 4176 3822 4189 3826
rect 4241 3830 4320 3846
rect 4352 3846 4524 3848
rect 4352 3830 4431 3846
rect 4438 3844 4468 3846
rect 4016 3808 4045 3818
rect 4059 3808 4088 3818
rect 4103 3808 4133 3822
rect 4176 3808 4219 3822
rect 4241 3818 4431 3830
rect 4496 3826 4502 3846
rect 4226 3808 4256 3818
rect 4257 3808 4415 3818
rect 4419 3808 4449 3818
rect 4453 3808 4483 3822
rect 4511 3808 4524 3846
rect 4596 3860 4625 3876
rect 4639 3860 4668 3876
rect 4683 3866 4713 3882
rect 4741 3860 4747 3908
rect 4750 3902 4769 3908
rect 4784 3902 4814 3910
rect 4750 3894 4814 3902
rect 4750 3878 4830 3894
rect 4846 3887 4908 3918
rect 4924 3887 4986 3918
rect 5055 3916 5104 3941
rect 5119 3916 5149 3932
rect 5018 3902 5048 3910
rect 5055 3908 5165 3916
rect 5018 3894 5063 3902
rect 4750 3876 4769 3878
rect 4784 3876 4830 3878
rect 4750 3860 4830 3876
rect 4857 3874 4892 3887
rect 4933 3884 4970 3887
rect 4933 3882 4975 3884
rect 4862 3871 4892 3874
rect 4871 3867 4878 3871
rect 4878 3866 4879 3867
rect 4837 3860 4847 3866
rect 4596 3852 4631 3860
rect 4596 3826 4597 3852
rect 4604 3826 4631 3852
rect 4539 3808 4569 3822
rect 4596 3818 4631 3826
rect 4633 3852 4674 3860
rect 4633 3826 4648 3852
rect 4655 3826 4674 3852
rect 4738 3848 4769 3860
rect 4784 3848 4887 3860
rect 4899 3850 4925 3876
rect 4940 3871 4970 3882
rect 5002 3878 5064 3894
rect 5002 3876 5048 3878
rect 5002 3860 5064 3876
rect 5076 3860 5082 3908
rect 5085 3900 5165 3908
rect 5085 3898 5104 3900
rect 5119 3898 5153 3900
rect 5085 3882 5165 3898
rect 5085 3860 5104 3882
rect 5119 3866 5149 3882
rect 5177 3876 5183 3950
rect 5186 3876 5205 4020
rect 5220 3876 5226 4020
rect 5235 3950 5248 4020
rect 5300 4016 5322 4020
rect 5293 3994 5322 4008
rect 5375 3994 5391 4008
rect 5429 4004 5435 4006
rect 5442 4004 5550 4020
rect 5557 4004 5563 4006
rect 5571 4004 5586 4020
rect 5652 4014 5671 4017
rect 5293 3992 5391 3994
rect 5418 3992 5586 4004
rect 5601 3994 5617 4008
rect 5652 3995 5674 4014
rect 5684 4008 5700 4009
rect 5683 4006 5700 4008
rect 5684 4001 5700 4006
rect 5674 3994 5680 3995
rect 5683 3994 5712 4001
rect 5601 3993 5712 3994
rect 5601 3992 5718 3993
rect 5277 3984 5328 3992
rect 5375 3984 5409 3992
rect 5277 3972 5302 3984
rect 5309 3972 5328 3984
rect 5382 3982 5409 3984
rect 5418 3982 5639 3992
rect 5674 3989 5680 3992
rect 5382 3978 5639 3982
rect 5277 3964 5328 3972
rect 5375 3964 5639 3978
rect 5683 3984 5718 3992
rect 5229 3916 5248 3950
rect 5293 3956 5322 3964
rect 5293 3950 5310 3956
rect 5293 3948 5327 3950
rect 5375 3948 5391 3964
rect 5392 3954 5600 3964
rect 5601 3954 5617 3964
rect 5665 3960 5680 3975
rect 5683 3972 5684 3984
rect 5691 3972 5718 3984
rect 5683 3964 5718 3972
rect 5683 3963 5712 3964
rect 5403 3950 5617 3954
rect 5418 3948 5617 3950
rect 5652 3950 5665 3960
rect 5683 3950 5700 3963
rect 5652 3948 5700 3950
rect 5294 3944 5327 3948
rect 5290 3942 5327 3944
rect 5290 3941 5357 3942
rect 5290 3936 5321 3941
rect 5327 3936 5357 3941
rect 5290 3932 5357 3936
rect 5263 3929 5357 3932
rect 5263 3922 5312 3929
rect 5263 3916 5293 3922
rect 5312 3917 5317 3922
rect 5229 3900 5309 3916
rect 5321 3908 5357 3929
rect 5418 3924 5607 3948
rect 5652 3947 5699 3948
rect 5665 3942 5699 3947
rect 5433 3921 5607 3924
rect 5426 3918 5607 3921
rect 5635 3941 5699 3942
rect 5229 3898 5248 3900
rect 5263 3898 5297 3900
rect 5229 3882 5309 3898
rect 5229 3876 5248 3882
rect 4945 3850 5048 3860
rect 4899 3848 5048 3850
rect 5069 3848 5104 3860
rect 4738 3846 4900 3848
rect 4750 3826 4769 3846
rect 4784 3844 4814 3846
rect 4633 3818 4674 3826
rect 4756 3822 4769 3826
rect 4821 3830 4900 3846
rect 4932 3846 5104 3848
rect 4932 3830 5011 3846
rect 5018 3844 5048 3846
rect 4596 3808 4625 3818
rect 4639 3808 4668 3818
rect 4683 3808 4713 3822
rect 4756 3808 4799 3822
rect 4821 3818 5011 3830
rect 5076 3826 5082 3846
rect 4806 3808 4836 3818
rect 4837 3808 4995 3818
rect 4999 3808 5029 3818
rect 5033 3808 5063 3822
rect 5091 3808 5104 3846
rect 5176 3860 5205 3876
rect 5219 3860 5248 3876
rect 5263 3866 5293 3882
rect 5321 3860 5327 3908
rect 5330 3902 5349 3908
rect 5364 3902 5394 3910
rect 5330 3894 5394 3902
rect 5330 3878 5410 3894
rect 5426 3887 5488 3918
rect 5504 3887 5566 3918
rect 5635 3916 5684 3941
rect 5699 3916 5729 3932
rect 5598 3902 5628 3910
rect 5635 3908 5745 3916
rect 5598 3894 5643 3902
rect 5330 3876 5349 3878
rect 5364 3876 5410 3878
rect 5330 3860 5410 3876
rect 5437 3874 5472 3887
rect 5513 3884 5550 3887
rect 5513 3882 5555 3884
rect 5442 3871 5472 3874
rect 5451 3867 5458 3871
rect 5458 3866 5459 3867
rect 5417 3860 5427 3866
rect 5176 3852 5211 3860
rect 5176 3826 5177 3852
rect 5184 3826 5211 3852
rect 5119 3808 5149 3822
rect 5176 3818 5211 3826
rect 5213 3852 5254 3860
rect 5213 3826 5228 3852
rect 5235 3826 5254 3852
rect 5318 3848 5349 3860
rect 5364 3848 5467 3860
rect 5479 3850 5505 3876
rect 5520 3871 5550 3882
rect 5582 3878 5644 3894
rect 5582 3876 5628 3878
rect 5582 3860 5644 3876
rect 5656 3860 5662 3908
rect 5665 3900 5745 3908
rect 5665 3898 5684 3900
rect 5699 3898 5733 3900
rect 5665 3882 5745 3898
rect 5665 3860 5684 3882
rect 5699 3866 5729 3882
rect 5757 3876 5763 3950
rect 5766 3876 5785 4020
rect 5800 3876 5806 4020
rect 5815 3950 5828 4020
rect 5880 4016 5902 4020
rect 5873 3994 5902 4008
rect 5955 3994 5971 4008
rect 6009 4004 6015 4006
rect 6022 4004 6130 4020
rect 6137 4004 6143 4006
rect 6151 4004 6166 4020
rect 6232 4014 6251 4017
rect 5873 3992 5971 3994
rect 5998 3992 6166 4004
rect 6181 3994 6197 4008
rect 6232 3995 6254 4014
rect 6264 4008 6280 4009
rect 6263 4006 6280 4008
rect 6264 4001 6280 4006
rect 6254 3994 6260 3995
rect 6263 3994 6292 4001
rect 6181 3993 6292 3994
rect 6181 3992 6298 3993
rect 5857 3984 5908 3992
rect 5955 3984 5989 3992
rect 5857 3972 5882 3984
rect 5889 3972 5908 3984
rect 5962 3982 5989 3984
rect 5998 3982 6219 3992
rect 6254 3989 6260 3992
rect 5962 3978 6219 3982
rect 5857 3964 5908 3972
rect 5955 3964 6219 3978
rect 6263 3984 6298 3992
rect 5809 3916 5828 3950
rect 5873 3956 5902 3964
rect 5873 3950 5890 3956
rect 5873 3948 5907 3950
rect 5955 3948 5971 3964
rect 5972 3954 6180 3964
rect 6181 3954 6197 3964
rect 6245 3960 6260 3975
rect 6263 3972 6264 3984
rect 6271 3972 6298 3984
rect 6263 3964 6298 3972
rect 6263 3963 6292 3964
rect 5983 3950 6197 3954
rect 5998 3948 6197 3950
rect 6232 3950 6245 3960
rect 6263 3950 6280 3963
rect 6232 3948 6280 3950
rect 5874 3944 5907 3948
rect 5870 3942 5907 3944
rect 5870 3941 5937 3942
rect 5870 3936 5901 3941
rect 5907 3936 5937 3941
rect 5870 3932 5937 3936
rect 5843 3929 5937 3932
rect 5843 3922 5892 3929
rect 5843 3916 5873 3922
rect 5892 3917 5897 3922
rect 5809 3900 5889 3916
rect 5901 3908 5937 3929
rect 5998 3924 6187 3948
rect 6232 3947 6279 3948
rect 6245 3942 6279 3947
rect 6013 3921 6187 3924
rect 6006 3918 6187 3921
rect 6215 3941 6279 3942
rect 5809 3898 5828 3900
rect 5843 3898 5877 3900
rect 5809 3882 5889 3898
rect 5809 3876 5828 3882
rect 5525 3850 5628 3860
rect 5479 3848 5628 3850
rect 5649 3848 5684 3860
rect 5318 3846 5480 3848
rect 5330 3826 5349 3846
rect 5364 3844 5394 3846
rect 5213 3818 5254 3826
rect 5336 3822 5349 3826
rect 5401 3830 5480 3846
rect 5512 3846 5684 3848
rect 5512 3830 5591 3846
rect 5598 3844 5628 3846
rect 5176 3808 5205 3818
rect 5219 3808 5248 3818
rect 5263 3808 5293 3822
rect 5336 3808 5379 3822
rect 5401 3818 5591 3830
rect 5656 3826 5662 3846
rect 5386 3808 5416 3818
rect 5417 3808 5575 3818
rect 5579 3808 5609 3818
rect 5613 3808 5643 3822
rect 5671 3808 5684 3846
rect 5756 3860 5785 3876
rect 5799 3860 5828 3876
rect 5843 3866 5873 3882
rect 5901 3860 5907 3908
rect 5910 3902 5929 3908
rect 5944 3902 5974 3910
rect 5910 3894 5974 3902
rect 5910 3878 5990 3894
rect 6006 3887 6068 3918
rect 6084 3887 6146 3918
rect 6215 3916 6264 3941
rect 6279 3916 6309 3932
rect 6178 3902 6208 3910
rect 6215 3908 6325 3916
rect 6178 3894 6223 3902
rect 5910 3876 5929 3878
rect 5944 3876 5990 3878
rect 5910 3860 5990 3876
rect 6017 3874 6052 3887
rect 6093 3884 6130 3887
rect 6093 3882 6135 3884
rect 6022 3871 6052 3874
rect 6031 3867 6038 3871
rect 6038 3866 6039 3867
rect 5997 3860 6007 3866
rect 5756 3852 5791 3860
rect 5756 3826 5757 3852
rect 5764 3826 5791 3852
rect 5699 3808 5729 3822
rect 5756 3818 5791 3826
rect 5793 3852 5834 3860
rect 5793 3826 5808 3852
rect 5815 3826 5834 3852
rect 5898 3848 5929 3860
rect 5944 3848 6047 3860
rect 6059 3850 6085 3876
rect 6100 3871 6130 3882
rect 6162 3878 6224 3894
rect 6162 3876 6208 3878
rect 6162 3860 6224 3876
rect 6236 3860 6242 3908
rect 6245 3900 6325 3908
rect 6245 3898 6264 3900
rect 6279 3898 6313 3900
rect 6245 3882 6325 3898
rect 6245 3860 6264 3882
rect 6279 3866 6309 3882
rect 6337 3876 6343 3950
rect 6346 3876 6365 4020
rect 6380 3876 6386 4020
rect 6395 3950 6408 4020
rect 6460 4016 6482 4020
rect 6453 3994 6482 4008
rect 6535 3994 6551 4008
rect 6589 4004 6595 4006
rect 6602 4004 6710 4020
rect 6717 4004 6723 4006
rect 6731 4004 6746 4020
rect 6812 4014 6831 4017
rect 6453 3992 6551 3994
rect 6578 3992 6746 4004
rect 6761 3994 6777 4008
rect 6812 3995 6834 4014
rect 6844 4008 6860 4009
rect 6843 4006 6860 4008
rect 6844 4001 6860 4006
rect 6834 3994 6840 3995
rect 6843 3994 6872 4001
rect 6761 3993 6872 3994
rect 6761 3992 6878 3993
rect 6437 3984 6488 3992
rect 6535 3984 6569 3992
rect 6437 3972 6462 3984
rect 6469 3972 6488 3984
rect 6542 3982 6569 3984
rect 6578 3982 6799 3992
rect 6834 3989 6840 3992
rect 6542 3978 6799 3982
rect 6437 3964 6488 3972
rect 6535 3964 6799 3978
rect 6843 3984 6878 3992
rect 6389 3916 6408 3950
rect 6453 3956 6482 3964
rect 6453 3950 6470 3956
rect 6453 3948 6487 3950
rect 6535 3948 6551 3964
rect 6552 3954 6760 3964
rect 6761 3954 6777 3964
rect 6825 3960 6840 3975
rect 6843 3972 6844 3984
rect 6851 3972 6878 3984
rect 6843 3964 6878 3972
rect 6843 3963 6872 3964
rect 6563 3950 6777 3954
rect 6578 3948 6777 3950
rect 6812 3950 6825 3960
rect 6843 3950 6860 3963
rect 6812 3948 6860 3950
rect 6454 3944 6487 3948
rect 6450 3942 6487 3944
rect 6450 3941 6517 3942
rect 6450 3936 6481 3941
rect 6487 3936 6517 3941
rect 6450 3932 6517 3936
rect 6423 3929 6517 3932
rect 6423 3922 6472 3929
rect 6423 3916 6453 3922
rect 6472 3917 6477 3922
rect 6389 3900 6469 3916
rect 6481 3908 6517 3929
rect 6578 3924 6767 3948
rect 6812 3947 6859 3948
rect 6825 3942 6859 3947
rect 6593 3921 6767 3924
rect 6586 3918 6767 3921
rect 6795 3941 6859 3942
rect 6389 3898 6408 3900
rect 6423 3898 6457 3900
rect 6389 3882 6469 3898
rect 6389 3876 6408 3882
rect 6105 3850 6208 3860
rect 6059 3848 6208 3850
rect 6229 3848 6264 3860
rect 5898 3846 6060 3848
rect 5910 3826 5929 3846
rect 5944 3844 5974 3846
rect 5793 3818 5834 3826
rect 5916 3822 5929 3826
rect 5981 3830 6060 3846
rect 6092 3846 6264 3848
rect 6092 3830 6171 3846
rect 6178 3844 6208 3846
rect 5756 3808 5785 3818
rect 5799 3808 5828 3818
rect 5843 3808 5873 3822
rect 5916 3808 5959 3822
rect 5981 3818 6171 3830
rect 6236 3826 6242 3846
rect 5966 3808 5996 3818
rect 5997 3808 6155 3818
rect 6159 3808 6189 3818
rect 6193 3808 6223 3822
rect 6251 3808 6264 3846
rect 6336 3860 6365 3876
rect 6379 3860 6408 3876
rect 6423 3866 6453 3882
rect 6481 3860 6487 3908
rect 6490 3902 6509 3908
rect 6524 3902 6554 3910
rect 6490 3894 6554 3902
rect 6490 3878 6570 3894
rect 6586 3887 6648 3918
rect 6664 3887 6726 3918
rect 6795 3916 6844 3941
rect 6859 3916 6889 3932
rect 6758 3902 6788 3910
rect 6795 3908 6905 3916
rect 6758 3894 6803 3902
rect 6490 3876 6509 3878
rect 6524 3876 6570 3878
rect 6490 3860 6570 3876
rect 6597 3874 6632 3887
rect 6673 3884 6710 3887
rect 6673 3882 6715 3884
rect 6602 3871 6632 3874
rect 6611 3867 6618 3871
rect 6618 3866 6619 3867
rect 6577 3860 6587 3866
rect 6336 3852 6371 3860
rect 6336 3826 6337 3852
rect 6344 3826 6371 3852
rect 6279 3808 6309 3822
rect 6336 3818 6371 3826
rect 6373 3852 6414 3860
rect 6373 3826 6388 3852
rect 6395 3826 6414 3852
rect 6478 3848 6509 3860
rect 6524 3848 6627 3860
rect 6639 3850 6665 3876
rect 6680 3871 6710 3882
rect 6742 3878 6804 3894
rect 6742 3876 6788 3878
rect 6742 3860 6804 3876
rect 6816 3860 6822 3908
rect 6825 3900 6905 3908
rect 6825 3898 6844 3900
rect 6859 3898 6893 3900
rect 6825 3882 6905 3898
rect 6825 3860 6844 3882
rect 6859 3866 6889 3882
rect 6917 3876 6923 3950
rect 6926 3876 6945 4020
rect 6960 3876 6966 4020
rect 6975 3950 6988 4020
rect 7040 4016 7062 4020
rect 7033 3994 7062 4008
rect 7115 3994 7131 4008
rect 7169 4004 7175 4006
rect 7182 4004 7290 4020
rect 7297 4004 7303 4006
rect 7311 4004 7326 4020
rect 7392 4014 7411 4017
rect 7033 3992 7131 3994
rect 7158 3992 7326 4004
rect 7341 3994 7357 4008
rect 7392 3995 7414 4014
rect 7424 4008 7440 4009
rect 7423 4006 7440 4008
rect 7424 4001 7440 4006
rect 7414 3994 7420 3995
rect 7423 3994 7452 4001
rect 7341 3993 7452 3994
rect 7341 3992 7458 3993
rect 7017 3984 7068 3992
rect 7115 3984 7149 3992
rect 7017 3972 7042 3984
rect 7049 3972 7068 3984
rect 7122 3982 7149 3984
rect 7158 3982 7379 3992
rect 7414 3989 7420 3992
rect 7122 3978 7379 3982
rect 7017 3964 7068 3972
rect 7115 3964 7379 3978
rect 7423 3984 7458 3992
rect 6969 3916 6988 3950
rect 7033 3956 7062 3964
rect 7033 3950 7050 3956
rect 7033 3948 7067 3950
rect 7115 3948 7131 3964
rect 7132 3954 7340 3964
rect 7341 3954 7357 3964
rect 7405 3960 7420 3975
rect 7423 3972 7424 3984
rect 7431 3972 7458 3984
rect 7423 3964 7458 3972
rect 7423 3963 7452 3964
rect 7143 3950 7357 3954
rect 7158 3948 7357 3950
rect 7392 3950 7405 3960
rect 7423 3950 7440 3963
rect 7392 3948 7440 3950
rect 7034 3944 7067 3948
rect 7030 3942 7067 3944
rect 7030 3941 7097 3942
rect 7030 3936 7061 3941
rect 7067 3936 7097 3941
rect 7030 3932 7097 3936
rect 7003 3929 7097 3932
rect 7003 3922 7052 3929
rect 7003 3916 7033 3922
rect 7052 3917 7057 3922
rect 6969 3900 7049 3916
rect 7061 3908 7097 3929
rect 7158 3924 7347 3948
rect 7392 3947 7439 3948
rect 7405 3942 7439 3947
rect 7173 3921 7347 3924
rect 7166 3918 7347 3921
rect 7375 3941 7439 3942
rect 6969 3898 6988 3900
rect 7003 3898 7037 3900
rect 6969 3882 7049 3898
rect 6969 3876 6988 3882
rect 6685 3850 6788 3860
rect 6639 3848 6788 3850
rect 6809 3848 6844 3860
rect 6478 3846 6640 3848
rect 6490 3826 6509 3846
rect 6524 3844 6554 3846
rect 6373 3818 6414 3826
rect 6496 3822 6509 3826
rect 6561 3830 6640 3846
rect 6672 3846 6844 3848
rect 6672 3830 6751 3846
rect 6758 3844 6788 3846
rect 6336 3808 6365 3818
rect 6379 3808 6408 3818
rect 6423 3808 6453 3822
rect 6496 3808 6539 3822
rect 6561 3818 6751 3830
rect 6816 3826 6822 3846
rect 6546 3808 6576 3818
rect 6577 3808 6735 3818
rect 6739 3808 6769 3818
rect 6773 3808 6803 3822
rect 6831 3808 6844 3846
rect 6916 3860 6945 3876
rect 6959 3860 6988 3876
rect 7003 3866 7033 3882
rect 7061 3860 7067 3908
rect 7070 3902 7089 3908
rect 7104 3902 7134 3910
rect 7070 3894 7134 3902
rect 7070 3878 7150 3894
rect 7166 3887 7228 3918
rect 7244 3887 7306 3918
rect 7375 3916 7424 3941
rect 7439 3916 7469 3932
rect 7338 3902 7368 3910
rect 7375 3908 7485 3916
rect 7338 3894 7383 3902
rect 7070 3876 7089 3878
rect 7104 3876 7150 3878
rect 7070 3860 7150 3876
rect 7177 3874 7212 3887
rect 7253 3884 7290 3887
rect 7253 3882 7295 3884
rect 7182 3871 7212 3874
rect 7191 3867 7198 3871
rect 7198 3866 7199 3867
rect 7157 3860 7167 3866
rect 6916 3852 6951 3860
rect 6916 3826 6917 3852
rect 6924 3826 6951 3852
rect 6859 3808 6889 3822
rect 6916 3818 6951 3826
rect 6953 3852 6994 3860
rect 6953 3826 6968 3852
rect 6975 3826 6994 3852
rect 7058 3848 7089 3860
rect 7104 3848 7207 3860
rect 7219 3850 7245 3876
rect 7260 3871 7290 3882
rect 7322 3878 7384 3894
rect 7322 3876 7368 3878
rect 7322 3860 7384 3876
rect 7396 3860 7402 3908
rect 7405 3900 7485 3908
rect 7405 3898 7424 3900
rect 7439 3898 7473 3900
rect 7405 3882 7485 3898
rect 7405 3860 7424 3882
rect 7439 3866 7469 3882
rect 7497 3876 7503 3950
rect 7506 3876 7525 4020
rect 7540 3876 7546 4020
rect 7555 3950 7568 4020
rect 7613 3998 7614 4008
rect 7629 3998 7642 4008
rect 7613 3994 7642 3998
rect 7647 3994 7677 4020
rect 7695 4006 7711 4008
rect 7783 4006 7836 4020
rect 7784 4004 7848 4006
rect 7891 4004 7906 4020
rect 7955 4017 7985 4020
rect 7955 4014 7991 4017
rect 7921 4006 7937 4008
rect 7695 3994 7710 3998
rect 7613 3992 7710 3994
rect 7738 3992 7906 4004
rect 7922 3994 7937 3998
rect 7955 3995 7994 4014
rect 8013 4008 8020 4009
rect 8019 4001 8020 4008
rect 8003 3998 8004 4001
rect 8019 3998 8032 4001
rect 7955 3994 7985 3995
rect 7994 3994 8000 3995
rect 8003 3994 8032 3998
rect 7922 3993 8032 3994
rect 7922 3992 8038 3993
rect 7597 3984 7648 3992
rect 7597 3972 7622 3984
rect 7629 3972 7648 3984
rect 7679 3984 7729 3992
rect 7679 3976 7695 3984
rect 7702 3982 7729 3984
rect 7738 3982 7959 3992
rect 7702 3972 7959 3982
rect 7988 3984 8038 3992
rect 7988 3975 8004 3984
rect 7597 3964 7648 3972
rect 7695 3964 7959 3972
rect 7985 3972 8004 3975
rect 8011 3972 8038 3984
rect 7985 3964 8038 3972
rect 7549 3916 7568 3950
rect 7613 3956 7614 3964
rect 7629 3956 7642 3964
rect 7613 3948 7629 3956
rect 7610 3941 7629 3944
rect 7610 3932 7632 3941
rect 7583 3922 7632 3932
rect 7583 3916 7613 3922
rect 7632 3917 7637 3922
rect 7549 3900 7629 3916
rect 7647 3908 7677 3964
rect 7712 3954 7920 3964
rect 7955 3960 8000 3964
rect 8003 3963 8004 3964
rect 8019 3963 8032 3964
rect 7738 3924 7927 3954
rect 7753 3921 7927 3924
rect 7746 3918 7927 3921
rect 7549 3898 7568 3900
rect 7583 3898 7617 3900
rect 7549 3882 7629 3898
rect 7656 3894 7669 3908
rect 7684 3894 7700 3910
rect 7746 3905 7757 3918
rect 7549 3876 7568 3882
rect 7265 3850 7368 3860
rect 7219 3848 7368 3850
rect 7389 3848 7424 3860
rect 7058 3846 7220 3848
rect 7070 3826 7089 3846
rect 7104 3844 7134 3846
rect 6953 3818 6994 3826
rect 7076 3822 7089 3826
rect 7141 3830 7220 3846
rect 7252 3846 7424 3848
rect 7252 3830 7331 3846
rect 7338 3844 7368 3846
rect 6916 3808 6945 3818
rect 6959 3808 6988 3818
rect 7003 3808 7033 3822
rect 7076 3808 7119 3822
rect 7141 3818 7331 3830
rect 7396 3826 7402 3846
rect 7126 3808 7156 3818
rect 7157 3808 7315 3818
rect 7319 3808 7349 3818
rect 7353 3808 7383 3822
rect 7411 3808 7424 3846
rect 7496 3860 7525 3876
rect 7539 3860 7568 3876
rect 7583 3860 7613 3882
rect 7656 3878 7718 3894
rect 7746 3887 7757 3903
rect 7762 3898 7772 3918
rect 7782 3898 7796 3918
rect 7799 3905 7808 3918
rect 7824 3905 7833 3918
rect 7762 3887 7796 3898
rect 7799 3887 7808 3903
rect 7824 3887 7833 3903
rect 7840 3898 7850 3918
rect 7860 3898 7874 3918
rect 7875 3905 7886 3918
rect 7840 3887 7874 3898
rect 7875 3887 7886 3903
rect 7932 3894 7948 3910
rect 7955 3908 7985 3960
rect 8019 3956 8020 3963
rect 8004 3948 8020 3956
rect 7991 3916 8004 3935
rect 8019 3916 8049 3932
rect 7991 3900 8065 3916
rect 7991 3898 8004 3900
rect 8019 3898 8053 3900
rect 7656 3876 7669 3878
rect 7684 3876 7718 3878
rect 7656 3860 7718 3876
rect 7762 3871 7778 3874
rect 7840 3871 7870 3882
rect 7918 3878 7964 3894
rect 7991 3882 8065 3898
rect 7918 3876 7952 3878
rect 7917 3860 7964 3876
rect 7991 3860 8004 3882
rect 8019 3860 8049 3882
rect 8076 3860 8077 3876
rect 8092 3860 8105 4020
rect 8135 3916 8148 4020
rect 8193 3998 8194 4008
rect 8209 3998 8222 4008
rect 8193 3994 8222 3998
rect 8227 3994 8257 4020
rect 8275 4006 8291 4008
rect 8363 4006 8416 4020
rect 8364 4004 8428 4006
rect 8471 4004 8486 4020
rect 8535 4017 8565 4020
rect 8535 4014 8571 4017
rect 8501 4006 8517 4008
rect 8275 3994 8290 3998
rect 8193 3992 8290 3994
rect 8318 3992 8486 4004
rect 8502 3994 8517 3998
rect 8535 3995 8574 4014
rect 8593 4008 8600 4009
rect 8599 4001 8600 4008
rect 8583 3998 8584 4001
rect 8599 3998 8612 4001
rect 8535 3994 8565 3995
rect 8574 3994 8580 3995
rect 8583 3994 8612 3998
rect 8502 3993 8612 3994
rect 8502 3992 8618 3993
rect 8177 3984 8228 3992
rect 8177 3972 8202 3984
rect 8209 3972 8228 3984
rect 8259 3984 8309 3992
rect 8259 3976 8275 3984
rect 8282 3982 8309 3984
rect 8318 3982 8539 3992
rect 8282 3972 8539 3982
rect 8568 3984 8618 3992
rect 8568 3975 8584 3984
rect 8177 3964 8228 3972
rect 8275 3964 8539 3972
rect 8565 3972 8584 3975
rect 8591 3972 8618 3984
rect 8565 3964 8618 3972
rect 8193 3956 8194 3964
rect 8209 3956 8222 3964
rect 8193 3948 8209 3956
rect 8190 3941 8209 3944
rect 8190 3932 8212 3941
rect 8163 3922 8212 3932
rect 8163 3916 8193 3922
rect 8212 3917 8217 3922
rect 8135 3900 8209 3916
rect 8227 3908 8257 3964
rect 8292 3954 8500 3964
rect 8535 3960 8580 3964
rect 8583 3963 8584 3964
rect 8599 3963 8612 3964
rect 8318 3924 8507 3954
rect 8333 3921 8507 3924
rect 8326 3918 8507 3921
rect 8135 3898 8148 3900
rect 8163 3898 8197 3900
rect 8135 3882 8209 3898
rect 8236 3894 8249 3908
rect 8264 3894 8280 3910
rect 8326 3905 8337 3918
rect 8119 3860 8120 3876
rect 8135 3860 8148 3882
rect 8163 3860 8193 3882
rect 8236 3878 8298 3894
rect 8326 3887 8337 3903
rect 8342 3898 8352 3918
rect 8362 3898 8376 3918
rect 8379 3905 8388 3918
rect 8404 3905 8413 3918
rect 8342 3887 8376 3898
rect 8379 3887 8388 3903
rect 8404 3887 8413 3903
rect 8420 3898 8430 3918
rect 8440 3898 8454 3918
rect 8455 3905 8466 3918
rect 8420 3887 8454 3898
rect 8455 3887 8466 3903
rect 8512 3894 8528 3910
rect 8535 3908 8565 3960
rect 8599 3956 8600 3963
rect 8584 3948 8600 3956
rect 8571 3916 8584 3935
rect 8599 3916 8629 3932
rect 8571 3900 8645 3916
rect 8571 3898 8584 3900
rect 8599 3898 8633 3900
rect 8236 3876 8249 3878
rect 8264 3876 8298 3878
rect 8236 3860 8298 3876
rect 8342 3871 8358 3874
rect 8420 3871 8450 3882
rect 8498 3878 8544 3894
rect 8571 3882 8645 3898
rect 8498 3876 8532 3878
rect 8497 3860 8544 3876
rect 8571 3860 8584 3882
rect 8599 3860 8629 3882
rect 8656 3860 8657 3876
rect 8672 3860 8685 4020
rect 8715 3916 8728 4020
rect 8773 3998 8774 4008
rect 8789 3998 8802 4008
rect 8773 3994 8802 3998
rect 8807 3994 8837 4020
rect 8855 4006 8871 4008
rect 8943 4006 8996 4020
rect 8944 4004 9008 4006
rect 9051 4004 9066 4020
rect 9115 4017 9145 4020
rect 9115 4014 9151 4017
rect 9081 4006 9097 4008
rect 8855 3994 8870 3998
rect 8773 3992 8870 3994
rect 8898 3992 9066 4004
rect 9082 3994 9097 3998
rect 9115 3995 9154 4014
rect 9173 4008 9180 4009
rect 9179 4001 9180 4008
rect 9163 3998 9164 4001
rect 9179 3998 9192 4001
rect 9115 3994 9145 3995
rect 9154 3994 9160 3995
rect 9163 3994 9192 3998
rect 9082 3993 9192 3994
rect 9082 3992 9198 3993
rect 8757 3984 8808 3992
rect 8757 3972 8782 3984
rect 8789 3972 8808 3984
rect 8839 3984 8889 3992
rect 8839 3976 8855 3984
rect 8862 3982 8889 3984
rect 8898 3982 9119 3992
rect 8862 3972 9119 3982
rect 9148 3984 9198 3992
rect 9148 3975 9164 3984
rect 8757 3964 8808 3972
rect 8855 3964 9119 3972
rect 9145 3972 9164 3975
rect 9171 3972 9198 3984
rect 9145 3964 9198 3972
rect 8773 3956 8774 3964
rect 8789 3956 8802 3964
rect 8773 3948 8789 3956
rect 8770 3941 8789 3944
rect 8770 3932 8792 3941
rect 8743 3922 8792 3932
rect 8743 3916 8773 3922
rect 8792 3917 8797 3922
rect 8715 3900 8789 3916
rect 8807 3908 8837 3964
rect 8872 3954 9080 3964
rect 9115 3960 9160 3964
rect 9163 3963 9164 3964
rect 9179 3963 9192 3964
rect 8898 3924 9087 3954
rect 8913 3921 9087 3924
rect 8906 3918 9087 3921
rect 8715 3898 8728 3900
rect 8743 3898 8777 3900
rect 8715 3882 8789 3898
rect 8816 3894 8829 3908
rect 8844 3894 8860 3910
rect 8906 3905 8917 3918
rect 8699 3860 8700 3876
rect 8715 3860 8728 3882
rect 8743 3860 8773 3882
rect 8816 3878 8878 3894
rect 8906 3887 8917 3903
rect 8922 3898 8932 3918
rect 8942 3898 8956 3918
rect 8959 3905 8968 3918
rect 8984 3905 8993 3918
rect 8922 3887 8956 3898
rect 8959 3887 8968 3903
rect 8984 3887 8993 3903
rect 9000 3898 9010 3918
rect 9020 3898 9034 3918
rect 9035 3905 9046 3918
rect 9000 3887 9034 3898
rect 9035 3887 9046 3903
rect 9092 3894 9108 3910
rect 9115 3908 9145 3960
rect 9179 3956 9180 3963
rect 9164 3948 9180 3956
rect 9151 3916 9164 3935
rect 9179 3916 9209 3932
rect 9151 3900 9225 3916
rect 9151 3898 9164 3900
rect 9179 3898 9213 3900
rect 8816 3876 8829 3878
rect 8844 3876 8878 3878
rect 8816 3860 8878 3876
rect 8922 3871 8938 3874
rect 9000 3871 9030 3882
rect 9078 3878 9124 3894
rect 9151 3882 9225 3898
rect 9078 3876 9112 3878
rect 9077 3860 9124 3876
rect 9151 3860 9164 3882
rect 9179 3860 9209 3882
rect 9236 3860 9237 3876
rect 9252 3860 9265 4020
rect 7496 3852 7531 3860
rect 7496 3826 7497 3852
rect 7504 3826 7531 3852
rect 7439 3808 7469 3822
rect 7496 3818 7531 3826
rect 7533 3852 7574 3860
rect 7533 3826 7548 3852
rect 7555 3826 7574 3852
rect 7638 3848 7700 3860
rect 7712 3848 7787 3860
rect 7845 3848 7920 3860
rect 7932 3848 7963 3860
rect 7969 3848 8004 3860
rect 7638 3846 7800 3848
rect 7533 3818 7574 3826
rect 7656 3822 7669 3846
rect 7684 3844 7699 3846
rect 7496 3808 7525 3818
rect 7539 3808 7568 3818
rect 7583 3808 7613 3822
rect 7656 3808 7699 3822
rect 7723 3819 7730 3826
rect 7733 3822 7800 3846
rect 7832 3846 8004 3848
rect 7802 3824 7830 3828
rect 7832 3824 7912 3846
rect 7933 3844 7948 3846
rect 7802 3822 7912 3824
rect 7733 3818 7912 3822
rect 7706 3808 7736 3818
rect 7738 3808 7891 3818
rect 7899 3808 7929 3818
rect 7933 3808 7963 3822
rect 7991 3808 8004 3846
rect 8076 3852 8111 3860
rect 8076 3826 8077 3852
rect 8084 3826 8111 3852
rect 8019 3808 8049 3822
rect 8076 3818 8111 3826
rect 8113 3852 8154 3860
rect 8113 3826 8128 3852
rect 8135 3826 8154 3852
rect 8218 3848 8280 3860
rect 8292 3848 8367 3860
rect 8425 3848 8500 3860
rect 8512 3848 8543 3860
rect 8549 3848 8584 3860
rect 8218 3846 8380 3848
rect 8113 3818 8154 3826
rect 8236 3822 8249 3846
rect 8264 3844 8279 3846
rect 8076 3808 8077 3818
rect 8092 3808 8105 3818
rect 8119 3808 8120 3818
rect 8135 3808 8148 3818
rect 8163 3808 8193 3822
rect 8236 3808 8279 3822
rect 8303 3819 8310 3826
rect 8313 3822 8380 3846
rect 8412 3846 8584 3848
rect 8382 3824 8410 3828
rect 8412 3824 8492 3846
rect 8513 3844 8528 3846
rect 8382 3822 8492 3824
rect 8313 3818 8492 3822
rect 8286 3808 8316 3818
rect 8318 3808 8471 3818
rect 8479 3808 8509 3818
rect 8513 3808 8543 3822
rect 8571 3808 8584 3846
rect 8656 3852 8691 3860
rect 8656 3826 8657 3852
rect 8664 3826 8691 3852
rect 8599 3808 8629 3822
rect 8656 3818 8691 3826
rect 8693 3852 8734 3860
rect 8693 3826 8708 3852
rect 8715 3826 8734 3852
rect 8798 3848 8860 3860
rect 8872 3848 8947 3860
rect 9005 3848 9080 3860
rect 9092 3848 9123 3860
rect 9129 3848 9164 3860
rect 8798 3846 8960 3848
rect 8693 3818 8734 3826
rect 8816 3822 8829 3846
rect 8844 3844 8859 3846
rect 8656 3808 8657 3818
rect 8672 3808 8685 3818
rect 8699 3808 8700 3818
rect 8715 3808 8728 3818
rect 8743 3808 8773 3822
rect 8816 3808 8859 3822
rect 8883 3819 8890 3826
rect 8893 3822 8960 3846
rect 8992 3846 9164 3848
rect 8962 3824 8990 3828
rect 8992 3824 9072 3846
rect 9093 3844 9108 3846
rect 8962 3822 9072 3824
rect 8893 3818 9072 3822
rect 8866 3808 8896 3818
rect 8898 3808 9051 3818
rect 9059 3808 9089 3818
rect 9093 3808 9123 3822
rect 9151 3808 9164 3846
rect 9236 3852 9271 3860
rect 9236 3826 9237 3852
rect 9244 3826 9271 3852
rect 9179 3808 9209 3822
rect 9236 3818 9271 3826
rect 9236 3808 9237 3818
rect 9252 3808 9265 3818
rect -1 3802 9265 3808
rect 0 3794 9265 3802
rect 15 3764 28 3794
rect 43 3780 73 3794
rect 116 3780 159 3794
rect 166 3780 386 3794
rect 393 3780 423 3794
rect 83 3766 98 3778
rect 117 3766 130 3780
rect 198 3776 351 3780
rect 80 3764 102 3766
rect 180 3764 372 3776
rect 451 3764 464 3794
rect 479 3780 509 3794
rect 546 3764 565 3794
rect 580 3764 586 3794
rect 595 3764 608 3794
rect 623 3780 653 3794
rect 696 3780 739 3794
rect 746 3780 966 3794
rect 973 3780 1003 3794
rect 663 3766 678 3778
rect 697 3766 710 3780
rect 778 3776 931 3780
rect 660 3764 682 3766
rect 760 3764 952 3776
rect 1031 3764 1044 3794
rect 1059 3780 1089 3794
rect 1126 3764 1145 3794
rect 1160 3764 1166 3794
rect 1175 3764 1188 3794
rect 1203 3780 1233 3794
rect 1276 3780 1319 3794
rect 1326 3780 1546 3794
rect 1553 3780 1583 3794
rect 1243 3766 1258 3778
rect 1277 3766 1290 3780
rect 1358 3776 1511 3780
rect 1240 3764 1262 3766
rect 1340 3764 1532 3776
rect 1611 3764 1624 3794
rect 1639 3780 1669 3794
rect 1706 3764 1725 3794
rect 1740 3764 1746 3794
rect 1755 3764 1768 3794
rect 1783 3780 1813 3794
rect 1856 3780 1899 3794
rect 1906 3780 2126 3794
rect 2133 3780 2163 3794
rect 1823 3766 1838 3778
rect 1857 3766 1870 3780
rect 1938 3776 2091 3780
rect 1820 3764 1842 3766
rect 1920 3764 2112 3776
rect 2191 3764 2204 3794
rect 2219 3780 2249 3794
rect 2286 3764 2305 3794
rect 2320 3764 2326 3794
rect 2335 3764 2348 3794
rect 2363 3780 2393 3794
rect 2436 3780 2479 3794
rect 2486 3780 2706 3794
rect 2713 3780 2743 3794
rect 2403 3766 2418 3778
rect 2437 3766 2450 3780
rect 2518 3776 2671 3780
rect 2400 3764 2422 3766
rect 2500 3764 2692 3776
rect 2771 3764 2784 3794
rect 2799 3780 2829 3794
rect 2866 3764 2885 3794
rect 2900 3764 2906 3794
rect 2915 3764 2928 3794
rect 2943 3780 2973 3794
rect 3016 3780 3059 3794
rect 3066 3780 3286 3794
rect 3293 3780 3323 3794
rect 2983 3766 2998 3778
rect 3017 3766 3030 3780
rect 3098 3776 3251 3780
rect 2980 3764 3002 3766
rect 3080 3764 3272 3776
rect 3351 3764 3364 3794
rect 3379 3780 3409 3794
rect 3446 3764 3465 3794
rect 3480 3764 3486 3794
rect 3495 3764 3508 3794
rect 3523 3780 3553 3794
rect 3596 3780 3639 3794
rect 3646 3780 3866 3794
rect 3873 3780 3903 3794
rect 3563 3766 3578 3778
rect 3597 3766 3610 3780
rect 3678 3776 3831 3780
rect 3560 3764 3582 3766
rect 3660 3764 3852 3776
rect 3931 3764 3944 3794
rect 3959 3780 3989 3794
rect 4026 3764 4045 3794
rect 4060 3764 4066 3794
rect 4075 3764 4088 3794
rect 4103 3780 4133 3794
rect 4176 3780 4219 3794
rect 4226 3780 4446 3794
rect 4453 3780 4483 3794
rect 4143 3766 4158 3778
rect 4177 3766 4190 3780
rect 4258 3776 4411 3780
rect 4140 3764 4162 3766
rect 4240 3764 4432 3776
rect 4511 3764 4524 3794
rect 4539 3780 4569 3794
rect 4606 3764 4625 3794
rect 4640 3764 4646 3794
rect 4655 3764 4668 3794
rect 4683 3780 4713 3794
rect 4756 3780 4799 3794
rect 4806 3780 5026 3794
rect 5033 3780 5063 3794
rect 4723 3766 4738 3778
rect 4757 3766 4770 3780
rect 4838 3776 4991 3780
rect 4720 3764 4742 3766
rect 4820 3764 5012 3776
rect 5091 3764 5104 3794
rect 5119 3780 5149 3794
rect 5186 3764 5205 3794
rect 5220 3764 5226 3794
rect 5235 3764 5248 3794
rect 5263 3780 5293 3794
rect 5336 3780 5379 3794
rect 5386 3780 5606 3794
rect 5613 3780 5643 3794
rect 5303 3766 5318 3778
rect 5337 3766 5350 3780
rect 5418 3776 5571 3780
rect 5300 3764 5322 3766
rect 5400 3764 5592 3776
rect 5671 3764 5684 3794
rect 5699 3780 5729 3794
rect 5766 3764 5785 3794
rect 5800 3764 5806 3794
rect 5815 3764 5828 3794
rect 5843 3780 5873 3794
rect 5916 3780 5959 3794
rect 5966 3780 6186 3794
rect 6193 3780 6223 3794
rect 5883 3766 5898 3778
rect 5917 3766 5930 3780
rect 5998 3776 6151 3780
rect 5880 3764 5902 3766
rect 5980 3764 6172 3776
rect 6251 3764 6264 3794
rect 6279 3780 6309 3794
rect 6346 3764 6365 3794
rect 6380 3764 6386 3794
rect 6395 3764 6408 3794
rect 6423 3780 6453 3794
rect 6496 3780 6539 3794
rect 6546 3780 6766 3794
rect 6773 3780 6803 3794
rect 6463 3766 6478 3778
rect 6497 3766 6510 3780
rect 6578 3776 6731 3780
rect 6460 3764 6482 3766
rect 6560 3764 6752 3776
rect 6831 3764 6844 3794
rect 6859 3780 6889 3794
rect 6926 3764 6945 3794
rect 6960 3764 6966 3794
rect 6975 3764 6988 3794
rect 7003 3780 7033 3794
rect 7076 3780 7119 3794
rect 7126 3780 7346 3794
rect 7353 3780 7383 3794
rect 7043 3766 7058 3778
rect 7077 3766 7090 3780
rect 7158 3776 7311 3780
rect 7040 3764 7062 3766
rect 7140 3764 7332 3776
rect 7411 3764 7424 3794
rect 7439 3780 7469 3794
rect 7506 3764 7525 3794
rect 7540 3764 7546 3794
rect 7555 3764 7568 3794
rect 7583 3776 7613 3794
rect 7656 3780 7670 3794
rect 7706 3780 7926 3794
rect 7657 3778 7670 3780
rect 7623 3766 7638 3778
rect 7620 3764 7642 3766
rect 7647 3764 7677 3778
rect 7738 3776 7891 3780
rect 7720 3764 7912 3776
rect 7955 3764 7985 3778
rect 7991 3764 8004 3794
rect 8019 3776 8049 3794
rect 8092 3764 8105 3794
rect 8135 3764 8148 3794
rect 8163 3776 8193 3794
rect 8236 3780 8250 3794
rect 8286 3780 8506 3794
rect 8237 3778 8250 3780
rect 8203 3766 8218 3778
rect 8200 3764 8222 3766
rect 8227 3764 8257 3778
rect 8318 3776 8471 3780
rect 8300 3764 8492 3776
rect 8535 3764 8565 3778
rect 8571 3764 8584 3794
rect 8599 3776 8629 3794
rect 8672 3764 8685 3794
rect 8715 3764 8728 3794
rect 8743 3776 8773 3794
rect 8816 3780 8830 3794
rect 8866 3780 9086 3794
rect 8817 3778 8830 3780
rect 8783 3766 8798 3778
rect 8780 3764 8802 3766
rect 8807 3764 8837 3778
rect 8898 3776 9051 3780
rect 8880 3764 9072 3776
rect 9115 3764 9145 3778
rect 9151 3764 9164 3794
rect 9179 3776 9209 3794
rect 9252 3764 9265 3794
rect 0 3750 9265 3764
rect 15 3680 28 3750
rect 80 3746 102 3750
rect 73 3724 102 3738
rect 155 3724 171 3738
rect 209 3734 215 3736
rect 222 3734 330 3750
rect 337 3734 343 3736
rect 351 3734 366 3750
rect 432 3744 451 3747
rect 73 3722 171 3724
rect 198 3722 366 3734
rect 381 3724 397 3738
rect 432 3725 454 3744
rect 464 3738 480 3739
rect 463 3736 480 3738
rect 464 3731 480 3736
rect 454 3724 460 3725
rect 463 3724 492 3731
rect 381 3723 492 3724
rect 381 3722 498 3723
rect 57 3714 108 3722
rect 155 3714 189 3722
rect 57 3702 82 3714
rect 89 3702 108 3714
rect 162 3712 189 3714
rect 198 3712 419 3722
rect 454 3719 460 3722
rect 162 3708 419 3712
rect 57 3694 108 3702
rect 155 3694 419 3708
rect 463 3714 498 3722
rect 9 3646 28 3680
rect 73 3686 102 3694
rect 73 3680 90 3686
rect 73 3678 107 3680
rect 155 3678 171 3694
rect 172 3684 380 3694
rect 381 3684 397 3694
rect 445 3690 460 3705
rect 463 3702 464 3714
rect 471 3702 498 3714
rect 463 3694 498 3702
rect 463 3693 492 3694
rect 183 3680 397 3684
rect 198 3678 397 3680
rect 432 3680 445 3690
rect 463 3680 480 3693
rect 432 3678 480 3680
rect 74 3674 107 3678
rect 70 3672 107 3674
rect 70 3671 137 3672
rect 70 3666 101 3671
rect 107 3666 137 3671
rect 70 3662 137 3666
rect 43 3659 137 3662
rect 43 3652 92 3659
rect 43 3646 73 3652
rect 92 3647 97 3652
rect 9 3630 89 3646
rect 101 3638 137 3659
rect 198 3654 387 3678
rect 432 3677 479 3678
rect 445 3672 479 3677
rect 213 3651 387 3654
rect 206 3648 387 3651
rect 415 3671 479 3672
rect 9 3628 28 3630
rect 43 3628 77 3630
rect 9 3612 89 3628
rect 9 3606 28 3612
rect -1 3590 28 3606
rect 43 3596 73 3612
rect 101 3590 107 3638
rect 110 3632 129 3638
rect 144 3632 174 3640
rect 110 3624 174 3632
rect 110 3608 190 3624
rect 206 3617 268 3648
rect 284 3617 346 3648
rect 415 3646 464 3671
rect 479 3646 509 3662
rect 378 3632 408 3640
rect 415 3638 525 3646
rect 378 3624 423 3632
rect 110 3606 129 3608
rect 144 3606 190 3608
rect 110 3590 190 3606
rect 217 3604 252 3617
rect 293 3614 330 3617
rect 293 3612 335 3614
rect 222 3601 252 3604
rect 231 3597 238 3601
rect 238 3596 239 3597
rect 197 3590 207 3596
rect -7 3582 34 3590
rect -7 3556 8 3582
rect 15 3556 34 3582
rect 98 3578 129 3590
rect 144 3578 247 3590
rect 259 3580 285 3606
rect 300 3601 330 3612
rect 362 3608 424 3624
rect 362 3606 408 3608
rect 362 3590 424 3606
rect 436 3590 442 3638
rect 445 3630 525 3638
rect 445 3628 464 3630
rect 479 3628 513 3630
rect 445 3612 525 3628
rect 445 3590 464 3612
rect 479 3596 509 3612
rect 537 3606 543 3680
rect 546 3606 565 3750
rect 580 3606 586 3750
rect 595 3680 608 3750
rect 660 3746 682 3750
rect 653 3724 682 3738
rect 735 3724 751 3738
rect 789 3734 795 3736
rect 802 3734 910 3750
rect 917 3734 923 3736
rect 931 3734 946 3750
rect 1012 3744 1031 3747
rect 653 3722 751 3724
rect 778 3722 946 3734
rect 961 3724 977 3738
rect 1012 3725 1034 3744
rect 1044 3738 1060 3739
rect 1043 3736 1060 3738
rect 1044 3731 1060 3736
rect 1034 3724 1040 3725
rect 1043 3724 1072 3731
rect 961 3723 1072 3724
rect 961 3722 1078 3723
rect 637 3714 688 3722
rect 735 3714 769 3722
rect 637 3702 662 3714
rect 669 3702 688 3714
rect 742 3712 769 3714
rect 778 3712 999 3722
rect 1034 3719 1040 3722
rect 742 3708 999 3712
rect 637 3694 688 3702
rect 735 3694 999 3708
rect 1043 3714 1078 3722
rect 589 3646 608 3680
rect 653 3686 682 3694
rect 653 3680 670 3686
rect 653 3678 687 3680
rect 735 3678 751 3694
rect 752 3684 960 3694
rect 961 3684 977 3694
rect 1025 3690 1040 3705
rect 1043 3702 1044 3714
rect 1051 3702 1078 3714
rect 1043 3694 1078 3702
rect 1043 3693 1072 3694
rect 763 3680 977 3684
rect 778 3678 977 3680
rect 1012 3680 1025 3690
rect 1043 3680 1060 3693
rect 1012 3678 1060 3680
rect 654 3674 687 3678
rect 650 3672 687 3674
rect 650 3671 717 3672
rect 650 3666 681 3671
rect 687 3666 717 3671
rect 650 3662 717 3666
rect 623 3659 717 3662
rect 623 3652 672 3659
rect 623 3646 653 3652
rect 672 3647 677 3652
rect 589 3630 669 3646
rect 681 3638 717 3659
rect 778 3654 967 3678
rect 1012 3677 1059 3678
rect 1025 3672 1059 3677
rect 793 3651 967 3654
rect 786 3648 967 3651
rect 995 3671 1059 3672
rect 589 3628 608 3630
rect 623 3628 657 3630
rect 589 3612 669 3628
rect 589 3606 608 3612
rect 305 3580 408 3590
rect 259 3578 408 3580
rect 429 3578 464 3590
rect 98 3576 260 3578
rect 110 3556 129 3576
rect 144 3574 174 3576
rect -7 3548 34 3556
rect 116 3552 129 3556
rect 181 3560 260 3576
rect 292 3576 464 3578
rect 292 3560 371 3576
rect 378 3574 408 3576
rect -1 3538 28 3548
rect 43 3538 73 3552
rect 116 3538 159 3552
rect 181 3548 371 3560
rect 436 3556 442 3576
rect 166 3538 196 3548
rect 197 3538 355 3548
rect 359 3538 389 3548
rect 393 3538 423 3552
rect 451 3538 464 3576
rect 536 3590 565 3606
rect 579 3590 608 3606
rect 623 3596 653 3612
rect 681 3590 687 3638
rect 690 3632 709 3638
rect 724 3632 754 3640
rect 690 3624 754 3632
rect 690 3608 770 3624
rect 786 3617 848 3648
rect 864 3617 926 3648
rect 995 3646 1044 3671
rect 1059 3646 1089 3662
rect 958 3632 988 3640
rect 995 3638 1105 3646
rect 958 3624 1003 3632
rect 690 3606 709 3608
rect 724 3606 770 3608
rect 690 3590 770 3606
rect 797 3604 832 3617
rect 873 3614 910 3617
rect 873 3612 915 3614
rect 802 3601 832 3604
rect 811 3597 818 3601
rect 818 3596 819 3597
rect 777 3590 787 3596
rect 536 3582 571 3590
rect 536 3556 537 3582
rect 544 3556 571 3582
rect 479 3538 509 3552
rect 536 3548 571 3556
rect 573 3582 614 3590
rect 573 3556 588 3582
rect 595 3556 614 3582
rect 678 3578 709 3590
rect 724 3578 827 3590
rect 839 3580 865 3606
rect 880 3601 910 3612
rect 942 3608 1004 3624
rect 942 3606 988 3608
rect 942 3590 1004 3606
rect 1016 3590 1022 3638
rect 1025 3630 1105 3638
rect 1025 3628 1044 3630
rect 1059 3628 1093 3630
rect 1025 3612 1105 3628
rect 1025 3590 1044 3612
rect 1059 3596 1089 3612
rect 1117 3606 1123 3680
rect 1126 3606 1145 3750
rect 1160 3606 1166 3750
rect 1175 3680 1188 3750
rect 1240 3746 1262 3750
rect 1233 3724 1262 3738
rect 1315 3724 1331 3738
rect 1369 3734 1375 3736
rect 1382 3734 1490 3750
rect 1497 3734 1503 3736
rect 1511 3734 1526 3750
rect 1592 3744 1611 3747
rect 1233 3722 1331 3724
rect 1358 3722 1526 3734
rect 1541 3724 1557 3738
rect 1592 3725 1614 3744
rect 1624 3738 1640 3739
rect 1623 3736 1640 3738
rect 1624 3731 1640 3736
rect 1614 3724 1620 3725
rect 1623 3724 1652 3731
rect 1541 3723 1652 3724
rect 1541 3722 1658 3723
rect 1217 3714 1268 3722
rect 1315 3714 1349 3722
rect 1217 3702 1242 3714
rect 1249 3702 1268 3714
rect 1322 3712 1349 3714
rect 1358 3712 1579 3722
rect 1614 3719 1620 3722
rect 1322 3708 1579 3712
rect 1217 3694 1268 3702
rect 1315 3694 1579 3708
rect 1623 3714 1658 3722
rect 1169 3646 1188 3680
rect 1233 3686 1262 3694
rect 1233 3680 1250 3686
rect 1233 3678 1267 3680
rect 1315 3678 1331 3694
rect 1332 3684 1540 3694
rect 1541 3684 1557 3694
rect 1605 3690 1620 3705
rect 1623 3702 1624 3714
rect 1631 3702 1658 3714
rect 1623 3694 1658 3702
rect 1623 3693 1652 3694
rect 1343 3680 1557 3684
rect 1358 3678 1557 3680
rect 1592 3680 1605 3690
rect 1623 3680 1640 3693
rect 1592 3678 1640 3680
rect 1234 3674 1267 3678
rect 1230 3672 1267 3674
rect 1230 3671 1297 3672
rect 1230 3666 1261 3671
rect 1267 3666 1297 3671
rect 1230 3662 1297 3666
rect 1203 3659 1297 3662
rect 1203 3652 1252 3659
rect 1203 3646 1233 3652
rect 1252 3647 1257 3652
rect 1169 3630 1249 3646
rect 1261 3638 1297 3659
rect 1358 3654 1547 3678
rect 1592 3677 1639 3678
rect 1605 3672 1639 3677
rect 1373 3651 1547 3654
rect 1366 3648 1547 3651
rect 1575 3671 1639 3672
rect 1169 3628 1188 3630
rect 1203 3628 1237 3630
rect 1169 3612 1249 3628
rect 1169 3606 1188 3612
rect 885 3580 988 3590
rect 839 3578 988 3580
rect 1009 3578 1044 3590
rect 678 3576 840 3578
rect 690 3556 709 3576
rect 724 3574 754 3576
rect 573 3548 614 3556
rect 696 3552 709 3556
rect 761 3560 840 3576
rect 872 3576 1044 3578
rect 872 3560 951 3576
rect 958 3574 988 3576
rect 536 3538 565 3548
rect 579 3538 608 3548
rect 623 3538 653 3552
rect 696 3538 739 3552
rect 761 3548 951 3560
rect 1016 3556 1022 3576
rect 746 3538 776 3548
rect 777 3538 935 3548
rect 939 3538 969 3548
rect 973 3538 1003 3552
rect 1031 3538 1044 3576
rect 1116 3590 1145 3606
rect 1159 3590 1188 3606
rect 1203 3596 1233 3612
rect 1261 3590 1267 3638
rect 1270 3632 1289 3638
rect 1304 3632 1334 3640
rect 1270 3624 1334 3632
rect 1270 3608 1350 3624
rect 1366 3617 1428 3648
rect 1444 3617 1506 3648
rect 1575 3646 1624 3671
rect 1639 3646 1669 3662
rect 1538 3632 1568 3640
rect 1575 3638 1685 3646
rect 1538 3624 1583 3632
rect 1270 3606 1289 3608
rect 1304 3606 1350 3608
rect 1270 3590 1350 3606
rect 1377 3604 1412 3617
rect 1453 3614 1490 3617
rect 1453 3612 1495 3614
rect 1382 3601 1412 3604
rect 1391 3597 1398 3601
rect 1398 3596 1399 3597
rect 1357 3590 1367 3596
rect 1116 3582 1151 3590
rect 1116 3556 1117 3582
rect 1124 3556 1151 3582
rect 1059 3538 1089 3552
rect 1116 3548 1151 3556
rect 1153 3582 1194 3590
rect 1153 3556 1168 3582
rect 1175 3556 1194 3582
rect 1258 3578 1289 3590
rect 1304 3578 1407 3590
rect 1419 3580 1445 3606
rect 1460 3601 1490 3612
rect 1522 3608 1584 3624
rect 1522 3606 1568 3608
rect 1522 3590 1584 3606
rect 1596 3590 1602 3638
rect 1605 3630 1685 3638
rect 1605 3628 1624 3630
rect 1639 3628 1673 3630
rect 1605 3612 1685 3628
rect 1605 3590 1624 3612
rect 1639 3596 1669 3612
rect 1697 3606 1703 3680
rect 1706 3606 1725 3750
rect 1740 3606 1746 3750
rect 1755 3680 1768 3750
rect 1820 3746 1842 3750
rect 1813 3724 1842 3738
rect 1895 3724 1911 3738
rect 1949 3734 1955 3736
rect 1962 3734 2070 3750
rect 2077 3734 2083 3736
rect 2091 3734 2106 3750
rect 2172 3744 2191 3747
rect 1813 3722 1911 3724
rect 1938 3722 2106 3734
rect 2121 3724 2137 3738
rect 2172 3725 2194 3744
rect 2204 3738 2220 3739
rect 2203 3736 2220 3738
rect 2204 3731 2220 3736
rect 2194 3724 2200 3725
rect 2203 3724 2232 3731
rect 2121 3723 2232 3724
rect 2121 3722 2238 3723
rect 1797 3714 1848 3722
rect 1895 3714 1929 3722
rect 1797 3702 1822 3714
rect 1829 3702 1848 3714
rect 1902 3712 1929 3714
rect 1938 3712 2159 3722
rect 2194 3719 2200 3722
rect 1902 3708 2159 3712
rect 1797 3694 1848 3702
rect 1895 3694 2159 3708
rect 2203 3714 2238 3722
rect 1749 3646 1768 3680
rect 1813 3686 1842 3694
rect 1813 3680 1830 3686
rect 1813 3678 1847 3680
rect 1895 3678 1911 3694
rect 1912 3684 2120 3694
rect 2121 3684 2137 3694
rect 2185 3690 2200 3705
rect 2203 3702 2204 3714
rect 2211 3702 2238 3714
rect 2203 3694 2238 3702
rect 2203 3693 2232 3694
rect 1923 3680 2137 3684
rect 1938 3678 2137 3680
rect 2172 3680 2185 3690
rect 2203 3680 2220 3693
rect 2172 3678 2220 3680
rect 1814 3674 1847 3678
rect 1810 3672 1847 3674
rect 1810 3671 1877 3672
rect 1810 3666 1841 3671
rect 1847 3666 1877 3671
rect 1810 3662 1877 3666
rect 1783 3659 1877 3662
rect 1783 3652 1832 3659
rect 1783 3646 1813 3652
rect 1832 3647 1837 3652
rect 1749 3630 1829 3646
rect 1841 3638 1877 3659
rect 1938 3654 2127 3678
rect 2172 3677 2219 3678
rect 2185 3672 2219 3677
rect 1953 3651 2127 3654
rect 1946 3648 2127 3651
rect 2155 3671 2219 3672
rect 1749 3628 1768 3630
rect 1783 3628 1817 3630
rect 1749 3612 1829 3628
rect 1749 3606 1768 3612
rect 1465 3580 1568 3590
rect 1419 3578 1568 3580
rect 1589 3578 1624 3590
rect 1258 3576 1420 3578
rect 1270 3556 1289 3576
rect 1304 3574 1334 3576
rect 1153 3548 1194 3556
rect 1276 3552 1289 3556
rect 1341 3560 1420 3576
rect 1452 3576 1624 3578
rect 1452 3560 1531 3576
rect 1538 3574 1568 3576
rect 1116 3538 1145 3548
rect 1159 3538 1188 3548
rect 1203 3538 1233 3552
rect 1276 3538 1319 3552
rect 1341 3548 1531 3560
rect 1596 3556 1602 3576
rect 1326 3538 1356 3548
rect 1357 3538 1515 3548
rect 1519 3538 1549 3548
rect 1553 3538 1583 3552
rect 1611 3538 1624 3576
rect 1696 3590 1725 3606
rect 1739 3590 1768 3606
rect 1783 3596 1813 3612
rect 1841 3590 1847 3638
rect 1850 3632 1869 3638
rect 1884 3632 1914 3640
rect 1850 3624 1914 3632
rect 1850 3608 1930 3624
rect 1946 3617 2008 3648
rect 2024 3617 2086 3648
rect 2155 3646 2204 3671
rect 2219 3646 2249 3662
rect 2118 3632 2148 3640
rect 2155 3638 2265 3646
rect 2118 3624 2163 3632
rect 1850 3606 1869 3608
rect 1884 3606 1930 3608
rect 1850 3590 1930 3606
rect 1957 3604 1992 3617
rect 2033 3614 2070 3617
rect 2033 3612 2075 3614
rect 1962 3601 1992 3604
rect 1971 3597 1978 3601
rect 1978 3596 1979 3597
rect 1937 3590 1947 3596
rect 1696 3582 1731 3590
rect 1696 3556 1697 3582
rect 1704 3556 1731 3582
rect 1639 3538 1669 3552
rect 1696 3548 1731 3556
rect 1733 3582 1774 3590
rect 1733 3556 1748 3582
rect 1755 3556 1774 3582
rect 1838 3578 1869 3590
rect 1884 3578 1987 3590
rect 1999 3580 2025 3606
rect 2040 3601 2070 3612
rect 2102 3608 2164 3624
rect 2102 3606 2148 3608
rect 2102 3590 2164 3606
rect 2176 3590 2182 3638
rect 2185 3630 2265 3638
rect 2185 3628 2204 3630
rect 2219 3628 2253 3630
rect 2185 3612 2265 3628
rect 2185 3590 2204 3612
rect 2219 3596 2249 3612
rect 2277 3606 2283 3680
rect 2286 3606 2305 3750
rect 2320 3606 2326 3750
rect 2335 3680 2348 3750
rect 2400 3746 2422 3750
rect 2393 3724 2422 3738
rect 2475 3724 2491 3738
rect 2529 3734 2535 3736
rect 2542 3734 2650 3750
rect 2657 3734 2663 3736
rect 2671 3734 2686 3750
rect 2752 3744 2771 3747
rect 2393 3722 2491 3724
rect 2518 3722 2686 3734
rect 2701 3724 2717 3738
rect 2752 3725 2774 3744
rect 2784 3738 2800 3739
rect 2783 3736 2800 3738
rect 2784 3731 2800 3736
rect 2774 3724 2780 3725
rect 2783 3724 2812 3731
rect 2701 3723 2812 3724
rect 2701 3722 2818 3723
rect 2377 3714 2428 3722
rect 2475 3714 2509 3722
rect 2377 3702 2402 3714
rect 2409 3702 2428 3714
rect 2482 3712 2509 3714
rect 2518 3712 2739 3722
rect 2774 3719 2780 3722
rect 2482 3708 2739 3712
rect 2377 3694 2428 3702
rect 2475 3694 2739 3708
rect 2783 3714 2818 3722
rect 2329 3646 2348 3680
rect 2393 3686 2422 3694
rect 2393 3680 2410 3686
rect 2393 3678 2427 3680
rect 2475 3678 2491 3694
rect 2492 3684 2700 3694
rect 2701 3684 2717 3694
rect 2765 3690 2780 3705
rect 2783 3702 2784 3714
rect 2791 3702 2818 3714
rect 2783 3694 2818 3702
rect 2783 3693 2812 3694
rect 2503 3680 2717 3684
rect 2518 3678 2717 3680
rect 2752 3680 2765 3690
rect 2783 3680 2800 3693
rect 2752 3678 2800 3680
rect 2394 3674 2427 3678
rect 2390 3672 2427 3674
rect 2390 3671 2457 3672
rect 2390 3666 2421 3671
rect 2427 3666 2457 3671
rect 2390 3662 2457 3666
rect 2363 3659 2457 3662
rect 2363 3652 2412 3659
rect 2363 3646 2393 3652
rect 2412 3647 2417 3652
rect 2329 3630 2409 3646
rect 2421 3638 2457 3659
rect 2518 3654 2707 3678
rect 2752 3677 2799 3678
rect 2765 3672 2799 3677
rect 2533 3651 2707 3654
rect 2526 3648 2707 3651
rect 2735 3671 2799 3672
rect 2329 3628 2348 3630
rect 2363 3628 2397 3630
rect 2329 3612 2409 3628
rect 2329 3606 2348 3612
rect 2045 3580 2148 3590
rect 1999 3578 2148 3580
rect 2169 3578 2204 3590
rect 1838 3576 2000 3578
rect 1850 3556 1869 3576
rect 1884 3574 1914 3576
rect 1733 3548 1774 3556
rect 1856 3552 1869 3556
rect 1921 3560 2000 3576
rect 2032 3576 2204 3578
rect 2032 3560 2111 3576
rect 2118 3574 2148 3576
rect 1696 3538 1725 3548
rect 1739 3538 1768 3548
rect 1783 3538 1813 3552
rect 1856 3538 1899 3552
rect 1921 3548 2111 3560
rect 2176 3556 2182 3576
rect 1906 3538 1936 3548
rect 1937 3538 2095 3548
rect 2099 3538 2129 3548
rect 2133 3538 2163 3552
rect 2191 3538 2204 3576
rect 2276 3590 2305 3606
rect 2319 3590 2348 3606
rect 2363 3596 2393 3612
rect 2421 3590 2427 3638
rect 2430 3632 2449 3638
rect 2464 3632 2494 3640
rect 2430 3624 2494 3632
rect 2430 3608 2510 3624
rect 2526 3617 2588 3648
rect 2604 3617 2666 3648
rect 2735 3646 2784 3671
rect 2799 3646 2829 3662
rect 2698 3632 2728 3640
rect 2735 3638 2845 3646
rect 2698 3624 2743 3632
rect 2430 3606 2449 3608
rect 2464 3606 2510 3608
rect 2430 3590 2510 3606
rect 2537 3604 2572 3617
rect 2613 3614 2650 3617
rect 2613 3612 2655 3614
rect 2542 3601 2572 3604
rect 2551 3597 2558 3601
rect 2558 3596 2559 3597
rect 2517 3590 2527 3596
rect 2276 3582 2311 3590
rect 2276 3556 2277 3582
rect 2284 3556 2311 3582
rect 2219 3538 2249 3552
rect 2276 3548 2311 3556
rect 2313 3582 2354 3590
rect 2313 3556 2328 3582
rect 2335 3556 2354 3582
rect 2418 3578 2449 3590
rect 2464 3578 2567 3590
rect 2579 3580 2605 3606
rect 2620 3601 2650 3612
rect 2682 3608 2744 3624
rect 2682 3606 2728 3608
rect 2682 3590 2744 3606
rect 2756 3590 2762 3638
rect 2765 3630 2845 3638
rect 2765 3628 2784 3630
rect 2799 3628 2833 3630
rect 2765 3612 2845 3628
rect 2765 3590 2784 3612
rect 2799 3596 2829 3612
rect 2857 3606 2863 3680
rect 2866 3606 2885 3750
rect 2900 3606 2906 3750
rect 2915 3680 2928 3750
rect 2980 3746 3002 3750
rect 2973 3724 3002 3738
rect 3055 3724 3071 3738
rect 3109 3734 3115 3736
rect 3122 3734 3230 3750
rect 3237 3734 3243 3736
rect 3251 3734 3266 3750
rect 3332 3744 3351 3747
rect 2973 3722 3071 3724
rect 3098 3722 3266 3734
rect 3281 3724 3297 3738
rect 3332 3725 3354 3744
rect 3364 3738 3380 3739
rect 3363 3736 3380 3738
rect 3364 3731 3380 3736
rect 3354 3724 3360 3725
rect 3363 3724 3392 3731
rect 3281 3723 3392 3724
rect 3281 3722 3398 3723
rect 2957 3714 3008 3722
rect 3055 3714 3089 3722
rect 2957 3702 2982 3714
rect 2989 3702 3008 3714
rect 3062 3712 3089 3714
rect 3098 3712 3319 3722
rect 3354 3719 3360 3722
rect 3062 3708 3319 3712
rect 2957 3694 3008 3702
rect 3055 3694 3319 3708
rect 3363 3714 3398 3722
rect 2909 3646 2928 3680
rect 2973 3686 3002 3694
rect 2973 3680 2990 3686
rect 2973 3678 3007 3680
rect 3055 3678 3071 3694
rect 3072 3684 3280 3694
rect 3281 3684 3297 3694
rect 3345 3690 3360 3705
rect 3363 3702 3364 3714
rect 3371 3702 3398 3714
rect 3363 3694 3398 3702
rect 3363 3693 3392 3694
rect 3083 3680 3297 3684
rect 3098 3678 3297 3680
rect 3332 3680 3345 3690
rect 3363 3680 3380 3693
rect 3332 3678 3380 3680
rect 2974 3674 3007 3678
rect 2970 3672 3007 3674
rect 2970 3671 3037 3672
rect 2970 3666 3001 3671
rect 3007 3666 3037 3671
rect 2970 3662 3037 3666
rect 2943 3659 3037 3662
rect 2943 3652 2992 3659
rect 2943 3646 2973 3652
rect 2992 3647 2997 3652
rect 2909 3630 2989 3646
rect 3001 3638 3037 3659
rect 3098 3654 3287 3678
rect 3332 3677 3379 3678
rect 3345 3672 3379 3677
rect 3113 3651 3287 3654
rect 3106 3648 3287 3651
rect 3315 3671 3379 3672
rect 2909 3628 2928 3630
rect 2943 3628 2977 3630
rect 2909 3612 2989 3628
rect 2909 3606 2928 3612
rect 2625 3580 2728 3590
rect 2579 3578 2728 3580
rect 2749 3578 2784 3590
rect 2418 3576 2580 3578
rect 2430 3556 2449 3576
rect 2464 3574 2494 3576
rect 2313 3548 2354 3556
rect 2436 3552 2449 3556
rect 2501 3560 2580 3576
rect 2612 3576 2784 3578
rect 2612 3560 2691 3576
rect 2698 3574 2728 3576
rect 2276 3538 2305 3548
rect 2319 3538 2348 3548
rect 2363 3538 2393 3552
rect 2436 3538 2479 3552
rect 2501 3548 2691 3560
rect 2756 3556 2762 3576
rect 2486 3538 2516 3548
rect 2517 3538 2675 3548
rect 2679 3538 2709 3548
rect 2713 3538 2743 3552
rect 2771 3538 2784 3576
rect 2856 3590 2885 3606
rect 2899 3590 2928 3606
rect 2943 3596 2973 3612
rect 3001 3590 3007 3638
rect 3010 3632 3029 3638
rect 3044 3632 3074 3640
rect 3010 3624 3074 3632
rect 3010 3608 3090 3624
rect 3106 3617 3168 3648
rect 3184 3617 3246 3648
rect 3315 3646 3364 3671
rect 3379 3646 3409 3662
rect 3278 3632 3308 3640
rect 3315 3638 3425 3646
rect 3278 3624 3323 3632
rect 3010 3606 3029 3608
rect 3044 3606 3090 3608
rect 3010 3590 3090 3606
rect 3117 3604 3152 3617
rect 3193 3614 3230 3617
rect 3193 3612 3235 3614
rect 3122 3601 3152 3604
rect 3131 3597 3138 3601
rect 3138 3596 3139 3597
rect 3097 3590 3107 3596
rect 2856 3582 2891 3590
rect 2856 3556 2857 3582
rect 2864 3556 2891 3582
rect 2799 3538 2829 3552
rect 2856 3548 2891 3556
rect 2893 3582 2934 3590
rect 2893 3556 2908 3582
rect 2915 3556 2934 3582
rect 2998 3578 3029 3590
rect 3044 3578 3147 3590
rect 3159 3580 3185 3606
rect 3200 3601 3230 3612
rect 3262 3608 3324 3624
rect 3262 3606 3308 3608
rect 3262 3590 3324 3606
rect 3336 3590 3342 3638
rect 3345 3630 3425 3638
rect 3345 3628 3364 3630
rect 3379 3628 3413 3630
rect 3345 3612 3425 3628
rect 3345 3590 3364 3612
rect 3379 3596 3409 3612
rect 3437 3606 3443 3680
rect 3446 3606 3465 3750
rect 3480 3606 3486 3750
rect 3495 3680 3508 3750
rect 3560 3746 3582 3750
rect 3553 3724 3582 3738
rect 3635 3724 3651 3738
rect 3689 3734 3695 3736
rect 3702 3734 3810 3750
rect 3817 3734 3823 3736
rect 3831 3734 3846 3750
rect 3912 3744 3931 3747
rect 3553 3722 3651 3724
rect 3678 3722 3846 3734
rect 3861 3724 3877 3738
rect 3912 3725 3934 3744
rect 3944 3738 3960 3739
rect 3943 3736 3960 3738
rect 3944 3731 3960 3736
rect 3934 3724 3940 3725
rect 3943 3724 3972 3731
rect 3861 3723 3972 3724
rect 3861 3722 3978 3723
rect 3537 3714 3588 3722
rect 3635 3714 3669 3722
rect 3537 3702 3562 3714
rect 3569 3702 3588 3714
rect 3642 3712 3669 3714
rect 3678 3712 3899 3722
rect 3934 3719 3940 3722
rect 3642 3708 3899 3712
rect 3537 3694 3588 3702
rect 3635 3694 3899 3708
rect 3943 3714 3978 3722
rect 3489 3646 3508 3680
rect 3553 3686 3582 3694
rect 3553 3680 3570 3686
rect 3553 3678 3587 3680
rect 3635 3678 3651 3694
rect 3652 3684 3860 3694
rect 3861 3684 3877 3694
rect 3925 3690 3940 3705
rect 3943 3702 3944 3714
rect 3951 3702 3978 3714
rect 3943 3694 3978 3702
rect 3943 3693 3972 3694
rect 3663 3680 3877 3684
rect 3678 3678 3877 3680
rect 3912 3680 3925 3690
rect 3943 3680 3960 3693
rect 3912 3678 3960 3680
rect 3554 3674 3587 3678
rect 3550 3672 3587 3674
rect 3550 3671 3617 3672
rect 3550 3666 3581 3671
rect 3587 3666 3617 3671
rect 3550 3662 3617 3666
rect 3523 3659 3617 3662
rect 3523 3652 3572 3659
rect 3523 3646 3553 3652
rect 3572 3647 3577 3652
rect 3489 3630 3569 3646
rect 3581 3638 3617 3659
rect 3678 3654 3867 3678
rect 3912 3677 3959 3678
rect 3925 3672 3959 3677
rect 3693 3651 3867 3654
rect 3686 3648 3867 3651
rect 3895 3671 3959 3672
rect 3489 3628 3508 3630
rect 3523 3628 3557 3630
rect 3489 3612 3569 3628
rect 3489 3606 3508 3612
rect 3205 3580 3308 3590
rect 3159 3578 3308 3580
rect 3329 3578 3364 3590
rect 2998 3576 3160 3578
rect 3010 3556 3029 3576
rect 3044 3574 3074 3576
rect 2893 3548 2934 3556
rect 3016 3552 3029 3556
rect 3081 3560 3160 3576
rect 3192 3576 3364 3578
rect 3192 3560 3271 3576
rect 3278 3574 3308 3576
rect 2856 3538 2885 3548
rect 2899 3538 2928 3548
rect 2943 3538 2973 3552
rect 3016 3538 3059 3552
rect 3081 3548 3271 3560
rect 3336 3556 3342 3576
rect 3066 3538 3096 3548
rect 3097 3538 3255 3548
rect 3259 3538 3289 3548
rect 3293 3538 3323 3552
rect 3351 3538 3364 3576
rect 3436 3590 3465 3606
rect 3479 3590 3508 3606
rect 3523 3596 3553 3612
rect 3581 3590 3587 3638
rect 3590 3632 3609 3638
rect 3624 3632 3654 3640
rect 3590 3624 3654 3632
rect 3590 3608 3670 3624
rect 3686 3617 3748 3648
rect 3764 3617 3826 3648
rect 3895 3646 3944 3671
rect 3959 3646 3989 3662
rect 3858 3632 3888 3640
rect 3895 3638 4005 3646
rect 3858 3624 3903 3632
rect 3590 3606 3609 3608
rect 3624 3606 3670 3608
rect 3590 3590 3670 3606
rect 3697 3604 3732 3617
rect 3773 3614 3810 3617
rect 3773 3612 3815 3614
rect 3702 3601 3732 3604
rect 3711 3597 3718 3601
rect 3718 3596 3719 3597
rect 3677 3590 3687 3596
rect 3436 3582 3471 3590
rect 3436 3556 3437 3582
rect 3444 3556 3471 3582
rect 3379 3538 3409 3552
rect 3436 3548 3471 3556
rect 3473 3582 3514 3590
rect 3473 3556 3488 3582
rect 3495 3556 3514 3582
rect 3578 3578 3609 3590
rect 3624 3578 3727 3590
rect 3739 3580 3765 3606
rect 3780 3601 3810 3612
rect 3842 3608 3904 3624
rect 3842 3606 3888 3608
rect 3842 3590 3904 3606
rect 3916 3590 3922 3638
rect 3925 3630 4005 3638
rect 3925 3628 3944 3630
rect 3959 3628 3993 3630
rect 3925 3612 4005 3628
rect 3925 3590 3944 3612
rect 3959 3596 3989 3612
rect 4017 3606 4023 3680
rect 4026 3606 4045 3750
rect 4060 3606 4066 3750
rect 4075 3680 4088 3750
rect 4140 3746 4162 3750
rect 4133 3724 4162 3738
rect 4215 3724 4231 3738
rect 4269 3734 4275 3736
rect 4282 3734 4390 3750
rect 4397 3734 4403 3736
rect 4411 3734 4426 3750
rect 4492 3744 4511 3747
rect 4133 3722 4231 3724
rect 4258 3722 4426 3734
rect 4441 3724 4457 3738
rect 4492 3725 4514 3744
rect 4524 3738 4540 3739
rect 4523 3736 4540 3738
rect 4524 3731 4540 3736
rect 4514 3724 4520 3725
rect 4523 3724 4552 3731
rect 4441 3723 4552 3724
rect 4441 3722 4558 3723
rect 4117 3714 4168 3722
rect 4215 3714 4249 3722
rect 4117 3702 4142 3714
rect 4149 3702 4168 3714
rect 4222 3712 4249 3714
rect 4258 3712 4479 3722
rect 4514 3719 4520 3722
rect 4222 3708 4479 3712
rect 4117 3694 4168 3702
rect 4215 3694 4479 3708
rect 4523 3714 4558 3722
rect 4069 3646 4088 3680
rect 4133 3686 4162 3694
rect 4133 3680 4150 3686
rect 4133 3678 4167 3680
rect 4215 3678 4231 3694
rect 4232 3684 4440 3694
rect 4441 3684 4457 3694
rect 4505 3690 4520 3705
rect 4523 3702 4524 3714
rect 4531 3702 4558 3714
rect 4523 3694 4558 3702
rect 4523 3693 4552 3694
rect 4243 3680 4457 3684
rect 4258 3678 4457 3680
rect 4492 3680 4505 3690
rect 4523 3680 4540 3693
rect 4492 3678 4540 3680
rect 4134 3674 4167 3678
rect 4130 3672 4167 3674
rect 4130 3671 4197 3672
rect 4130 3666 4161 3671
rect 4167 3666 4197 3671
rect 4130 3662 4197 3666
rect 4103 3659 4197 3662
rect 4103 3652 4152 3659
rect 4103 3646 4133 3652
rect 4152 3647 4157 3652
rect 4069 3630 4149 3646
rect 4161 3638 4197 3659
rect 4258 3654 4447 3678
rect 4492 3677 4539 3678
rect 4505 3672 4539 3677
rect 4273 3651 4447 3654
rect 4266 3648 4447 3651
rect 4475 3671 4539 3672
rect 4069 3628 4088 3630
rect 4103 3628 4137 3630
rect 4069 3612 4149 3628
rect 4069 3606 4088 3612
rect 3785 3580 3888 3590
rect 3739 3578 3888 3580
rect 3909 3578 3944 3590
rect 3578 3576 3740 3578
rect 3590 3556 3609 3576
rect 3624 3574 3654 3576
rect 3473 3548 3514 3556
rect 3596 3552 3609 3556
rect 3661 3560 3740 3576
rect 3772 3576 3944 3578
rect 3772 3560 3851 3576
rect 3858 3574 3888 3576
rect 3436 3538 3465 3548
rect 3479 3538 3508 3548
rect 3523 3538 3553 3552
rect 3596 3538 3639 3552
rect 3661 3548 3851 3560
rect 3916 3556 3922 3576
rect 3646 3538 3676 3548
rect 3677 3538 3835 3548
rect 3839 3538 3869 3548
rect 3873 3538 3903 3552
rect 3931 3538 3944 3576
rect 4016 3590 4045 3606
rect 4059 3590 4088 3606
rect 4103 3596 4133 3612
rect 4161 3590 4167 3638
rect 4170 3632 4189 3638
rect 4204 3632 4234 3640
rect 4170 3624 4234 3632
rect 4170 3608 4250 3624
rect 4266 3617 4328 3648
rect 4344 3617 4406 3648
rect 4475 3646 4524 3671
rect 4539 3646 4569 3662
rect 4438 3632 4468 3640
rect 4475 3638 4585 3646
rect 4438 3624 4483 3632
rect 4170 3606 4189 3608
rect 4204 3606 4250 3608
rect 4170 3590 4250 3606
rect 4277 3604 4312 3617
rect 4353 3614 4390 3617
rect 4353 3612 4395 3614
rect 4282 3601 4312 3604
rect 4291 3597 4298 3601
rect 4298 3596 4299 3597
rect 4257 3590 4267 3596
rect 4016 3582 4051 3590
rect 4016 3556 4017 3582
rect 4024 3556 4051 3582
rect 3959 3538 3989 3552
rect 4016 3548 4051 3556
rect 4053 3582 4094 3590
rect 4053 3556 4068 3582
rect 4075 3556 4094 3582
rect 4158 3578 4189 3590
rect 4204 3578 4307 3590
rect 4319 3580 4345 3606
rect 4360 3601 4390 3612
rect 4422 3608 4484 3624
rect 4422 3606 4468 3608
rect 4422 3590 4484 3606
rect 4496 3590 4502 3638
rect 4505 3630 4585 3638
rect 4505 3628 4524 3630
rect 4539 3628 4573 3630
rect 4505 3612 4585 3628
rect 4505 3590 4524 3612
rect 4539 3596 4569 3612
rect 4597 3606 4603 3680
rect 4606 3606 4625 3750
rect 4640 3606 4646 3750
rect 4655 3680 4668 3750
rect 4720 3746 4742 3750
rect 4713 3724 4742 3738
rect 4795 3724 4811 3738
rect 4849 3734 4855 3736
rect 4862 3734 4970 3750
rect 4977 3734 4983 3736
rect 4991 3734 5006 3750
rect 5072 3744 5091 3747
rect 4713 3722 4811 3724
rect 4838 3722 5006 3734
rect 5021 3724 5037 3738
rect 5072 3725 5094 3744
rect 5104 3738 5120 3739
rect 5103 3736 5120 3738
rect 5104 3731 5120 3736
rect 5094 3724 5100 3725
rect 5103 3724 5132 3731
rect 5021 3723 5132 3724
rect 5021 3722 5138 3723
rect 4697 3714 4748 3722
rect 4795 3714 4829 3722
rect 4697 3702 4722 3714
rect 4729 3702 4748 3714
rect 4802 3712 4829 3714
rect 4838 3712 5059 3722
rect 5094 3719 5100 3722
rect 4802 3708 5059 3712
rect 4697 3694 4748 3702
rect 4795 3694 5059 3708
rect 5103 3714 5138 3722
rect 4649 3646 4668 3680
rect 4713 3686 4742 3694
rect 4713 3680 4730 3686
rect 4713 3678 4747 3680
rect 4795 3678 4811 3694
rect 4812 3684 5020 3694
rect 5021 3684 5037 3694
rect 5085 3690 5100 3705
rect 5103 3702 5104 3714
rect 5111 3702 5138 3714
rect 5103 3694 5138 3702
rect 5103 3693 5132 3694
rect 4823 3680 5037 3684
rect 4838 3678 5037 3680
rect 5072 3680 5085 3690
rect 5103 3680 5120 3693
rect 5072 3678 5120 3680
rect 4714 3674 4747 3678
rect 4710 3672 4747 3674
rect 4710 3671 4777 3672
rect 4710 3666 4741 3671
rect 4747 3666 4777 3671
rect 4710 3662 4777 3666
rect 4683 3659 4777 3662
rect 4683 3652 4732 3659
rect 4683 3646 4713 3652
rect 4732 3647 4737 3652
rect 4649 3630 4729 3646
rect 4741 3638 4777 3659
rect 4838 3654 5027 3678
rect 5072 3677 5119 3678
rect 5085 3672 5119 3677
rect 4853 3651 5027 3654
rect 4846 3648 5027 3651
rect 5055 3671 5119 3672
rect 4649 3628 4668 3630
rect 4683 3628 4717 3630
rect 4649 3612 4729 3628
rect 4649 3606 4668 3612
rect 4365 3580 4468 3590
rect 4319 3578 4468 3580
rect 4489 3578 4524 3590
rect 4158 3576 4320 3578
rect 4170 3556 4189 3576
rect 4204 3574 4234 3576
rect 4053 3548 4094 3556
rect 4176 3552 4189 3556
rect 4241 3560 4320 3576
rect 4352 3576 4524 3578
rect 4352 3560 4431 3576
rect 4438 3574 4468 3576
rect 4016 3538 4045 3548
rect 4059 3538 4088 3548
rect 4103 3538 4133 3552
rect 4176 3538 4219 3552
rect 4241 3548 4431 3560
rect 4496 3556 4502 3576
rect 4226 3538 4256 3548
rect 4257 3538 4415 3548
rect 4419 3538 4449 3548
rect 4453 3538 4483 3552
rect 4511 3538 4524 3576
rect 4596 3590 4625 3606
rect 4639 3590 4668 3606
rect 4683 3596 4713 3612
rect 4741 3590 4747 3638
rect 4750 3632 4769 3638
rect 4784 3632 4814 3640
rect 4750 3624 4814 3632
rect 4750 3608 4830 3624
rect 4846 3617 4908 3648
rect 4924 3617 4986 3648
rect 5055 3646 5104 3671
rect 5119 3646 5149 3662
rect 5018 3632 5048 3640
rect 5055 3638 5165 3646
rect 5018 3624 5063 3632
rect 4750 3606 4769 3608
rect 4784 3606 4830 3608
rect 4750 3590 4830 3606
rect 4857 3604 4892 3617
rect 4933 3614 4970 3617
rect 4933 3612 4975 3614
rect 4862 3601 4892 3604
rect 4871 3597 4878 3601
rect 4878 3596 4879 3597
rect 4837 3590 4847 3596
rect 4596 3582 4631 3590
rect 4596 3556 4597 3582
rect 4604 3556 4631 3582
rect 4539 3538 4569 3552
rect 4596 3548 4631 3556
rect 4633 3582 4674 3590
rect 4633 3556 4648 3582
rect 4655 3556 4674 3582
rect 4738 3578 4769 3590
rect 4784 3578 4887 3590
rect 4899 3580 4925 3606
rect 4940 3601 4970 3612
rect 5002 3608 5064 3624
rect 5002 3606 5048 3608
rect 5002 3590 5064 3606
rect 5076 3590 5082 3638
rect 5085 3630 5165 3638
rect 5085 3628 5104 3630
rect 5119 3628 5153 3630
rect 5085 3612 5165 3628
rect 5085 3590 5104 3612
rect 5119 3596 5149 3612
rect 5177 3606 5183 3680
rect 5186 3606 5205 3750
rect 5220 3606 5226 3750
rect 5235 3680 5248 3750
rect 5300 3746 5322 3750
rect 5293 3724 5322 3738
rect 5375 3724 5391 3738
rect 5429 3734 5435 3736
rect 5442 3734 5550 3750
rect 5557 3734 5563 3736
rect 5571 3734 5586 3750
rect 5652 3744 5671 3747
rect 5293 3722 5391 3724
rect 5418 3722 5586 3734
rect 5601 3724 5617 3738
rect 5652 3725 5674 3744
rect 5684 3738 5700 3739
rect 5683 3736 5700 3738
rect 5684 3731 5700 3736
rect 5674 3724 5680 3725
rect 5683 3724 5712 3731
rect 5601 3723 5712 3724
rect 5601 3722 5718 3723
rect 5277 3714 5328 3722
rect 5375 3714 5409 3722
rect 5277 3702 5302 3714
rect 5309 3702 5328 3714
rect 5382 3712 5409 3714
rect 5418 3712 5639 3722
rect 5674 3719 5680 3722
rect 5382 3708 5639 3712
rect 5277 3694 5328 3702
rect 5375 3694 5639 3708
rect 5683 3714 5718 3722
rect 5229 3646 5248 3680
rect 5293 3686 5322 3694
rect 5293 3680 5310 3686
rect 5293 3678 5327 3680
rect 5375 3678 5391 3694
rect 5392 3684 5600 3694
rect 5601 3684 5617 3694
rect 5665 3690 5680 3705
rect 5683 3702 5684 3714
rect 5691 3702 5718 3714
rect 5683 3694 5718 3702
rect 5683 3693 5712 3694
rect 5403 3680 5617 3684
rect 5418 3678 5617 3680
rect 5652 3680 5665 3690
rect 5683 3680 5700 3693
rect 5652 3678 5700 3680
rect 5294 3674 5327 3678
rect 5290 3672 5327 3674
rect 5290 3671 5357 3672
rect 5290 3666 5321 3671
rect 5327 3666 5357 3671
rect 5290 3662 5357 3666
rect 5263 3659 5357 3662
rect 5263 3652 5312 3659
rect 5263 3646 5293 3652
rect 5312 3647 5317 3652
rect 5229 3630 5309 3646
rect 5321 3638 5357 3659
rect 5418 3654 5607 3678
rect 5652 3677 5699 3678
rect 5665 3672 5699 3677
rect 5433 3651 5607 3654
rect 5426 3648 5607 3651
rect 5635 3671 5699 3672
rect 5229 3628 5248 3630
rect 5263 3628 5297 3630
rect 5229 3612 5309 3628
rect 5229 3606 5248 3612
rect 4945 3580 5048 3590
rect 4899 3578 5048 3580
rect 5069 3578 5104 3590
rect 4738 3576 4900 3578
rect 4750 3556 4769 3576
rect 4784 3574 4814 3576
rect 4633 3548 4674 3556
rect 4756 3552 4769 3556
rect 4821 3560 4900 3576
rect 4932 3576 5104 3578
rect 4932 3560 5011 3576
rect 5018 3574 5048 3576
rect 4596 3538 4625 3548
rect 4639 3538 4668 3548
rect 4683 3538 4713 3552
rect 4756 3538 4799 3552
rect 4821 3548 5011 3560
rect 5076 3556 5082 3576
rect 4806 3538 4836 3548
rect 4837 3538 4995 3548
rect 4999 3538 5029 3548
rect 5033 3538 5063 3552
rect 5091 3538 5104 3576
rect 5176 3590 5205 3606
rect 5219 3590 5248 3606
rect 5263 3596 5293 3612
rect 5321 3590 5327 3638
rect 5330 3632 5349 3638
rect 5364 3632 5394 3640
rect 5330 3624 5394 3632
rect 5330 3608 5410 3624
rect 5426 3617 5488 3648
rect 5504 3617 5566 3648
rect 5635 3646 5684 3671
rect 5699 3646 5729 3662
rect 5598 3632 5628 3640
rect 5635 3638 5745 3646
rect 5598 3624 5643 3632
rect 5330 3606 5349 3608
rect 5364 3606 5410 3608
rect 5330 3590 5410 3606
rect 5437 3604 5472 3617
rect 5513 3614 5550 3617
rect 5513 3612 5555 3614
rect 5442 3601 5472 3604
rect 5451 3597 5458 3601
rect 5458 3596 5459 3597
rect 5417 3590 5427 3596
rect 5176 3582 5211 3590
rect 5176 3556 5177 3582
rect 5184 3556 5211 3582
rect 5119 3538 5149 3552
rect 5176 3548 5211 3556
rect 5213 3582 5254 3590
rect 5213 3556 5228 3582
rect 5235 3556 5254 3582
rect 5318 3578 5349 3590
rect 5364 3578 5467 3590
rect 5479 3580 5505 3606
rect 5520 3601 5550 3612
rect 5582 3608 5644 3624
rect 5582 3606 5628 3608
rect 5582 3590 5644 3606
rect 5656 3590 5662 3638
rect 5665 3630 5745 3638
rect 5665 3628 5684 3630
rect 5699 3628 5733 3630
rect 5665 3612 5745 3628
rect 5665 3590 5684 3612
rect 5699 3596 5729 3612
rect 5757 3606 5763 3680
rect 5766 3606 5785 3750
rect 5800 3606 5806 3750
rect 5815 3680 5828 3750
rect 5880 3746 5902 3750
rect 5873 3724 5902 3738
rect 5955 3724 5971 3738
rect 6009 3734 6015 3736
rect 6022 3734 6130 3750
rect 6137 3734 6143 3736
rect 6151 3734 6166 3750
rect 6232 3744 6251 3747
rect 5873 3722 5971 3724
rect 5998 3722 6166 3734
rect 6181 3724 6197 3738
rect 6232 3725 6254 3744
rect 6264 3738 6280 3739
rect 6263 3736 6280 3738
rect 6264 3731 6280 3736
rect 6254 3724 6260 3725
rect 6263 3724 6292 3731
rect 6181 3723 6292 3724
rect 6181 3722 6298 3723
rect 5857 3714 5908 3722
rect 5955 3714 5989 3722
rect 5857 3702 5882 3714
rect 5889 3702 5908 3714
rect 5962 3712 5989 3714
rect 5998 3712 6219 3722
rect 6254 3719 6260 3722
rect 5962 3708 6219 3712
rect 5857 3694 5908 3702
rect 5955 3694 6219 3708
rect 6263 3714 6298 3722
rect 5809 3646 5828 3680
rect 5873 3686 5902 3694
rect 5873 3680 5890 3686
rect 5873 3678 5907 3680
rect 5955 3678 5971 3694
rect 5972 3684 6180 3694
rect 6181 3684 6197 3694
rect 6245 3690 6260 3705
rect 6263 3702 6264 3714
rect 6271 3702 6298 3714
rect 6263 3694 6298 3702
rect 6263 3693 6292 3694
rect 5983 3680 6197 3684
rect 5998 3678 6197 3680
rect 6232 3680 6245 3690
rect 6263 3680 6280 3693
rect 6232 3678 6280 3680
rect 5874 3674 5907 3678
rect 5870 3672 5907 3674
rect 5870 3671 5937 3672
rect 5870 3666 5901 3671
rect 5907 3666 5937 3671
rect 5870 3662 5937 3666
rect 5843 3659 5937 3662
rect 5843 3652 5892 3659
rect 5843 3646 5873 3652
rect 5892 3647 5897 3652
rect 5809 3630 5889 3646
rect 5901 3638 5937 3659
rect 5998 3654 6187 3678
rect 6232 3677 6279 3678
rect 6245 3672 6279 3677
rect 6013 3651 6187 3654
rect 6006 3648 6187 3651
rect 6215 3671 6279 3672
rect 5809 3628 5828 3630
rect 5843 3628 5877 3630
rect 5809 3612 5889 3628
rect 5809 3606 5828 3612
rect 5525 3580 5628 3590
rect 5479 3578 5628 3580
rect 5649 3578 5684 3590
rect 5318 3576 5480 3578
rect 5330 3556 5349 3576
rect 5364 3574 5394 3576
rect 5213 3548 5254 3556
rect 5336 3552 5349 3556
rect 5401 3560 5480 3576
rect 5512 3576 5684 3578
rect 5512 3560 5591 3576
rect 5598 3574 5628 3576
rect 5176 3538 5205 3548
rect 5219 3538 5248 3548
rect 5263 3538 5293 3552
rect 5336 3538 5379 3552
rect 5401 3548 5591 3560
rect 5656 3556 5662 3576
rect 5386 3538 5416 3548
rect 5417 3538 5575 3548
rect 5579 3538 5609 3548
rect 5613 3538 5643 3552
rect 5671 3538 5684 3576
rect 5756 3590 5785 3606
rect 5799 3590 5828 3606
rect 5843 3596 5873 3612
rect 5901 3590 5907 3638
rect 5910 3632 5929 3638
rect 5944 3632 5974 3640
rect 5910 3624 5974 3632
rect 5910 3608 5990 3624
rect 6006 3617 6068 3648
rect 6084 3617 6146 3648
rect 6215 3646 6264 3671
rect 6279 3646 6309 3662
rect 6178 3632 6208 3640
rect 6215 3638 6325 3646
rect 6178 3624 6223 3632
rect 5910 3606 5929 3608
rect 5944 3606 5990 3608
rect 5910 3590 5990 3606
rect 6017 3604 6052 3617
rect 6093 3614 6130 3617
rect 6093 3612 6135 3614
rect 6022 3601 6052 3604
rect 6031 3597 6038 3601
rect 6038 3596 6039 3597
rect 5997 3590 6007 3596
rect 5756 3582 5791 3590
rect 5756 3556 5757 3582
rect 5764 3556 5791 3582
rect 5699 3538 5729 3552
rect 5756 3548 5791 3556
rect 5793 3582 5834 3590
rect 5793 3556 5808 3582
rect 5815 3556 5834 3582
rect 5898 3578 5929 3590
rect 5944 3578 6047 3590
rect 6059 3580 6085 3606
rect 6100 3601 6130 3612
rect 6162 3608 6224 3624
rect 6162 3606 6208 3608
rect 6162 3590 6224 3606
rect 6236 3590 6242 3638
rect 6245 3630 6325 3638
rect 6245 3628 6264 3630
rect 6279 3628 6313 3630
rect 6245 3612 6325 3628
rect 6245 3590 6264 3612
rect 6279 3596 6309 3612
rect 6337 3606 6343 3680
rect 6346 3606 6365 3750
rect 6380 3606 6386 3750
rect 6395 3680 6408 3750
rect 6460 3746 6482 3750
rect 6453 3724 6482 3738
rect 6535 3724 6551 3738
rect 6589 3734 6595 3736
rect 6602 3734 6710 3750
rect 6717 3734 6723 3736
rect 6731 3734 6746 3750
rect 6812 3744 6831 3747
rect 6453 3722 6551 3724
rect 6578 3722 6746 3734
rect 6761 3724 6777 3738
rect 6812 3725 6834 3744
rect 6844 3738 6860 3739
rect 6843 3736 6860 3738
rect 6844 3731 6860 3736
rect 6834 3724 6840 3725
rect 6843 3724 6872 3731
rect 6761 3723 6872 3724
rect 6761 3722 6878 3723
rect 6437 3714 6488 3722
rect 6535 3714 6569 3722
rect 6437 3702 6462 3714
rect 6469 3702 6488 3714
rect 6542 3712 6569 3714
rect 6578 3712 6799 3722
rect 6834 3719 6840 3722
rect 6542 3708 6799 3712
rect 6437 3694 6488 3702
rect 6535 3694 6799 3708
rect 6843 3714 6878 3722
rect 6389 3646 6408 3680
rect 6453 3686 6482 3694
rect 6453 3680 6470 3686
rect 6453 3678 6487 3680
rect 6535 3678 6551 3694
rect 6552 3684 6760 3694
rect 6761 3684 6777 3694
rect 6825 3690 6840 3705
rect 6843 3702 6844 3714
rect 6851 3702 6878 3714
rect 6843 3694 6878 3702
rect 6843 3693 6872 3694
rect 6563 3680 6777 3684
rect 6578 3678 6777 3680
rect 6812 3680 6825 3690
rect 6843 3680 6860 3693
rect 6812 3678 6860 3680
rect 6454 3674 6487 3678
rect 6450 3672 6487 3674
rect 6450 3671 6517 3672
rect 6450 3666 6481 3671
rect 6487 3666 6517 3671
rect 6450 3662 6517 3666
rect 6423 3659 6517 3662
rect 6423 3652 6472 3659
rect 6423 3646 6453 3652
rect 6472 3647 6477 3652
rect 6389 3630 6469 3646
rect 6481 3638 6517 3659
rect 6578 3654 6767 3678
rect 6812 3677 6859 3678
rect 6825 3672 6859 3677
rect 6593 3651 6767 3654
rect 6586 3648 6767 3651
rect 6795 3671 6859 3672
rect 6389 3628 6408 3630
rect 6423 3628 6457 3630
rect 6389 3612 6469 3628
rect 6389 3606 6408 3612
rect 6105 3580 6208 3590
rect 6059 3578 6208 3580
rect 6229 3578 6264 3590
rect 5898 3576 6060 3578
rect 5910 3556 5929 3576
rect 5944 3574 5974 3576
rect 5793 3548 5834 3556
rect 5916 3552 5929 3556
rect 5981 3560 6060 3576
rect 6092 3576 6264 3578
rect 6092 3560 6171 3576
rect 6178 3574 6208 3576
rect 5756 3538 5785 3548
rect 5799 3538 5828 3548
rect 5843 3538 5873 3552
rect 5916 3538 5959 3552
rect 5981 3548 6171 3560
rect 6236 3556 6242 3576
rect 5966 3538 5996 3548
rect 5997 3538 6155 3548
rect 6159 3538 6189 3548
rect 6193 3538 6223 3552
rect 6251 3538 6264 3576
rect 6336 3590 6365 3606
rect 6379 3590 6408 3606
rect 6423 3596 6453 3612
rect 6481 3590 6487 3638
rect 6490 3632 6509 3638
rect 6524 3632 6554 3640
rect 6490 3624 6554 3632
rect 6490 3608 6570 3624
rect 6586 3617 6648 3648
rect 6664 3617 6726 3648
rect 6795 3646 6844 3671
rect 6859 3646 6889 3662
rect 6758 3632 6788 3640
rect 6795 3638 6905 3646
rect 6758 3624 6803 3632
rect 6490 3606 6509 3608
rect 6524 3606 6570 3608
rect 6490 3590 6570 3606
rect 6597 3604 6632 3617
rect 6673 3614 6710 3617
rect 6673 3612 6715 3614
rect 6602 3601 6632 3604
rect 6611 3597 6618 3601
rect 6618 3596 6619 3597
rect 6577 3590 6587 3596
rect 6336 3582 6371 3590
rect 6336 3556 6337 3582
rect 6344 3556 6371 3582
rect 6279 3538 6309 3552
rect 6336 3548 6371 3556
rect 6373 3582 6414 3590
rect 6373 3556 6388 3582
rect 6395 3556 6414 3582
rect 6478 3578 6509 3590
rect 6524 3578 6627 3590
rect 6639 3580 6665 3606
rect 6680 3601 6710 3612
rect 6742 3608 6804 3624
rect 6742 3606 6788 3608
rect 6742 3590 6804 3606
rect 6816 3590 6822 3638
rect 6825 3630 6905 3638
rect 6825 3628 6844 3630
rect 6859 3628 6893 3630
rect 6825 3612 6905 3628
rect 6825 3590 6844 3612
rect 6859 3596 6889 3612
rect 6917 3606 6923 3680
rect 6926 3606 6945 3750
rect 6960 3606 6966 3750
rect 6975 3680 6988 3750
rect 7040 3746 7062 3750
rect 7033 3724 7062 3738
rect 7115 3724 7131 3738
rect 7169 3734 7175 3736
rect 7182 3734 7290 3750
rect 7297 3734 7303 3736
rect 7311 3734 7326 3750
rect 7392 3744 7411 3747
rect 7033 3722 7131 3724
rect 7158 3722 7326 3734
rect 7341 3724 7357 3738
rect 7392 3725 7414 3744
rect 7424 3738 7440 3739
rect 7423 3736 7440 3738
rect 7424 3731 7440 3736
rect 7414 3724 7420 3725
rect 7423 3724 7452 3731
rect 7341 3723 7452 3724
rect 7341 3722 7458 3723
rect 7017 3714 7068 3722
rect 7115 3714 7149 3722
rect 7017 3702 7042 3714
rect 7049 3702 7068 3714
rect 7122 3712 7149 3714
rect 7158 3712 7379 3722
rect 7414 3719 7420 3722
rect 7122 3708 7379 3712
rect 7017 3694 7068 3702
rect 7115 3694 7379 3708
rect 7423 3714 7458 3722
rect 6969 3646 6988 3680
rect 7033 3686 7062 3694
rect 7033 3680 7050 3686
rect 7033 3678 7067 3680
rect 7115 3678 7131 3694
rect 7132 3684 7340 3694
rect 7341 3684 7357 3694
rect 7405 3690 7420 3705
rect 7423 3702 7424 3714
rect 7431 3702 7458 3714
rect 7423 3694 7458 3702
rect 7423 3693 7452 3694
rect 7143 3680 7357 3684
rect 7158 3678 7357 3680
rect 7392 3680 7405 3690
rect 7423 3680 7440 3693
rect 7392 3678 7440 3680
rect 7034 3674 7067 3678
rect 7030 3672 7067 3674
rect 7030 3671 7097 3672
rect 7030 3666 7061 3671
rect 7067 3666 7097 3671
rect 7030 3662 7097 3666
rect 7003 3659 7097 3662
rect 7003 3652 7052 3659
rect 7003 3646 7033 3652
rect 7052 3647 7057 3652
rect 6969 3630 7049 3646
rect 7061 3638 7097 3659
rect 7158 3654 7347 3678
rect 7392 3677 7439 3678
rect 7405 3672 7439 3677
rect 7173 3651 7347 3654
rect 7166 3648 7347 3651
rect 7375 3671 7439 3672
rect 6969 3628 6988 3630
rect 7003 3628 7037 3630
rect 6969 3612 7049 3628
rect 6969 3606 6988 3612
rect 6685 3580 6788 3590
rect 6639 3578 6788 3580
rect 6809 3578 6844 3590
rect 6478 3576 6640 3578
rect 6490 3556 6509 3576
rect 6524 3574 6554 3576
rect 6373 3548 6414 3556
rect 6496 3552 6509 3556
rect 6561 3560 6640 3576
rect 6672 3576 6844 3578
rect 6672 3560 6751 3576
rect 6758 3574 6788 3576
rect 6336 3538 6365 3548
rect 6379 3538 6408 3548
rect 6423 3538 6453 3552
rect 6496 3538 6539 3552
rect 6561 3548 6751 3560
rect 6816 3556 6822 3576
rect 6546 3538 6576 3548
rect 6577 3538 6735 3548
rect 6739 3538 6769 3548
rect 6773 3538 6803 3552
rect 6831 3538 6844 3576
rect 6916 3590 6945 3606
rect 6959 3590 6988 3606
rect 7003 3596 7033 3612
rect 7061 3590 7067 3638
rect 7070 3632 7089 3638
rect 7104 3632 7134 3640
rect 7070 3624 7134 3632
rect 7070 3608 7150 3624
rect 7166 3617 7228 3648
rect 7244 3617 7306 3648
rect 7375 3646 7424 3671
rect 7439 3646 7469 3662
rect 7338 3632 7368 3640
rect 7375 3638 7485 3646
rect 7338 3624 7383 3632
rect 7070 3606 7089 3608
rect 7104 3606 7150 3608
rect 7070 3590 7150 3606
rect 7177 3604 7212 3617
rect 7253 3614 7290 3617
rect 7253 3612 7295 3614
rect 7182 3601 7212 3604
rect 7191 3597 7198 3601
rect 7198 3596 7199 3597
rect 7157 3590 7167 3596
rect 6916 3582 6951 3590
rect 6916 3556 6917 3582
rect 6924 3556 6951 3582
rect 6859 3538 6889 3552
rect 6916 3548 6951 3556
rect 6953 3582 6994 3590
rect 6953 3556 6968 3582
rect 6975 3556 6994 3582
rect 7058 3578 7089 3590
rect 7104 3578 7207 3590
rect 7219 3580 7245 3606
rect 7260 3601 7290 3612
rect 7322 3608 7384 3624
rect 7322 3606 7368 3608
rect 7322 3590 7384 3606
rect 7396 3590 7402 3638
rect 7405 3630 7485 3638
rect 7405 3628 7424 3630
rect 7439 3628 7473 3630
rect 7405 3612 7485 3628
rect 7405 3590 7424 3612
rect 7439 3596 7469 3612
rect 7497 3606 7503 3680
rect 7506 3606 7525 3750
rect 7540 3606 7546 3750
rect 7555 3680 7568 3750
rect 7613 3728 7614 3738
rect 7629 3728 7642 3738
rect 7613 3724 7642 3728
rect 7647 3724 7677 3750
rect 7695 3736 7711 3738
rect 7783 3736 7836 3750
rect 7784 3734 7848 3736
rect 7891 3734 7906 3750
rect 7955 3747 7985 3750
rect 7955 3744 7991 3747
rect 7921 3736 7937 3738
rect 7695 3724 7710 3728
rect 7613 3722 7710 3724
rect 7738 3722 7906 3734
rect 7922 3724 7937 3728
rect 7955 3725 7994 3744
rect 8013 3738 8020 3739
rect 8019 3731 8020 3738
rect 8003 3728 8004 3731
rect 8019 3728 8032 3731
rect 7955 3724 7985 3725
rect 7994 3724 8000 3725
rect 8003 3724 8032 3728
rect 7922 3723 8032 3724
rect 7922 3722 8038 3723
rect 7597 3714 7648 3722
rect 7597 3702 7622 3714
rect 7629 3702 7648 3714
rect 7679 3714 7729 3722
rect 7679 3706 7695 3714
rect 7702 3712 7729 3714
rect 7738 3712 7959 3722
rect 7702 3702 7959 3712
rect 7988 3714 8038 3722
rect 7988 3705 8004 3714
rect 7597 3694 7648 3702
rect 7695 3694 7959 3702
rect 7985 3702 8004 3705
rect 8011 3702 8038 3714
rect 7985 3694 8038 3702
rect 7549 3646 7568 3680
rect 7613 3686 7614 3694
rect 7629 3686 7642 3694
rect 7613 3678 7629 3686
rect 7610 3671 7629 3674
rect 7610 3662 7632 3671
rect 7583 3652 7632 3662
rect 7583 3646 7613 3652
rect 7632 3647 7637 3652
rect 7549 3630 7629 3646
rect 7647 3638 7677 3694
rect 7712 3684 7920 3694
rect 7955 3690 8000 3694
rect 8003 3693 8004 3694
rect 8019 3693 8032 3694
rect 7738 3654 7927 3684
rect 7753 3651 7927 3654
rect 7746 3648 7927 3651
rect 7549 3628 7568 3630
rect 7583 3628 7617 3630
rect 7549 3612 7629 3628
rect 7656 3624 7669 3638
rect 7684 3624 7700 3640
rect 7746 3635 7757 3648
rect 7549 3606 7568 3612
rect 7265 3580 7368 3590
rect 7219 3578 7368 3580
rect 7389 3578 7424 3590
rect 7058 3576 7220 3578
rect 7070 3556 7089 3576
rect 7104 3574 7134 3576
rect 6953 3548 6994 3556
rect 7076 3552 7089 3556
rect 7141 3560 7220 3576
rect 7252 3576 7424 3578
rect 7252 3560 7331 3576
rect 7338 3574 7368 3576
rect 6916 3538 6945 3548
rect 6959 3538 6988 3548
rect 7003 3538 7033 3552
rect 7076 3538 7119 3552
rect 7141 3548 7331 3560
rect 7396 3556 7402 3576
rect 7126 3538 7156 3548
rect 7157 3538 7315 3548
rect 7319 3538 7349 3548
rect 7353 3538 7383 3552
rect 7411 3538 7424 3576
rect 7496 3590 7525 3606
rect 7539 3590 7568 3606
rect 7583 3590 7613 3612
rect 7656 3608 7718 3624
rect 7746 3617 7757 3633
rect 7762 3628 7772 3648
rect 7782 3628 7796 3648
rect 7799 3635 7808 3648
rect 7824 3635 7833 3648
rect 7762 3617 7796 3628
rect 7799 3617 7808 3633
rect 7824 3617 7833 3633
rect 7840 3628 7850 3648
rect 7860 3628 7874 3648
rect 7875 3635 7886 3648
rect 7840 3617 7874 3628
rect 7875 3617 7886 3633
rect 7932 3624 7948 3640
rect 7955 3638 7985 3690
rect 8019 3686 8020 3693
rect 8004 3678 8020 3686
rect 7991 3646 8004 3665
rect 8019 3646 8049 3662
rect 7991 3630 8065 3646
rect 7991 3628 8004 3630
rect 8019 3628 8053 3630
rect 7656 3606 7669 3608
rect 7684 3606 7718 3608
rect 7656 3590 7718 3606
rect 7762 3601 7778 3604
rect 7840 3601 7870 3612
rect 7918 3608 7964 3624
rect 7991 3612 8065 3628
rect 7918 3606 7952 3608
rect 7917 3590 7964 3606
rect 7991 3590 8004 3612
rect 8019 3590 8049 3612
rect 8076 3590 8077 3606
rect 8092 3590 8105 3750
rect 8135 3646 8148 3750
rect 8193 3728 8194 3738
rect 8209 3728 8222 3738
rect 8193 3724 8222 3728
rect 8227 3724 8257 3750
rect 8275 3736 8291 3738
rect 8363 3736 8416 3750
rect 8364 3734 8428 3736
rect 8471 3734 8486 3750
rect 8535 3747 8565 3750
rect 8535 3744 8571 3747
rect 8501 3736 8517 3738
rect 8275 3724 8290 3728
rect 8193 3722 8290 3724
rect 8318 3722 8486 3734
rect 8502 3724 8517 3728
rect 8535 3725 8574 3744
rect 8593 3738 8600 3739
rect 8599 3731 8600 3738
rect 8583 3728 8584 3731
rect 8599 3728 8612 3731
rect 8535 3724 8565 3725
rect 8574 3724 8580 3725
rect 8583 3724 8612 3728
rect 8502 3723 8612 3724
rect 8502 3722 8618 3723
rect 8177 3714 8228 3722
rect 8177 3702 8202 3714
rect 8209 3702 8228 3714
rect 8259 3714 8309 3722
rect 8259 3706 8275 3714
rect 8282 3712 8309 3714
rect 8318 3712 8539 3722
rect 8282 3702 8539 3712
rect 8568 3714 8618 3722
rect 8568 3705 8584 3714
rect 8177 3694 8228 3702
rect 8275 3694 8539 3702
rect 8565 3702 8584 3705
rect 8591 3702 8618 3714
rect 8565 3694 8618 3702
rect 8193 3686 8194 3694
rect 8209 3686 8222 3694
rect 8193 3678 8209 3686
rect 8190 3671 8209 3674
rect 8190 3662 8212 3671
rect 8163 3652 8212 3662
rect 8163 3646 8193 3652
rect 8212 3647 8217 3652
rect 8135 3630 8209 3646
rect 8227 3638 8257 3694
rect 8292 3684 8500 3694
rect 8535 3690 8580 3694
rect 8583 3693 8584 3694
rect 8599 3693 8612 3694
rect 8318 3654 8507 3684
rect 8333 3651 8507 3654
rect 8326 3648 8507 3651
rect 8135 3628 8148 3630
rect 8163 3628 8197 3630
rect 8135 3612 8209 3628
rect 8236 3624 8249 3638
rect 8264 3624 8280 3640
rect 8326 3635 8337 3648
rect 8119 3590 8120 3606
rect 8135 3590 8148 3612
rect 8163 3590 8193 3612
rect 8236 3608 8298 3624
rect 8326 3617 8337 3633
rect 8342 3628 8352 3648
rect 8362 3628 8376 3648
rect 8379 3635 8388 3648
rect 8404 3635 8413 3648
rect 8342 3617 8376 3628
rect 8379 3617 8388 3633
rect 8404 3617 8413 3633
rect 8420 3628 8430 3648
rect 8440 3628 8454 3648
rect 8455 3635 8466 3648
rect 8420 3617 8454 3628
rect 8455 3617 8466 3633
rect 8512 3624 8528 3640
rect 8535 3638 8565 3690
rect 8599 3686 8600 3693
rect 8584 3678 8600 3686
rect 8571 3646 8584 3665
rect 8599 3646 8629 3662
rect 8571 3630 8645 3646
rect 8571 3628 8584 3630
rect 8599 3628 8633 3630
rect 8236 3606 8249 3608
rect 8264 3606 8298 3608
rect 8236 3590 8298 3606
rect 8342 3601 8358 3604
rect 8420 3601 8450 3612
rect 8498 3608 8544 3624
rect 8571 3612 8645 3628
rect 8498 3606 8532 3608
rect 8497 3590 8544 3606
rect 8571 3590 8584 3612
rect 8599 3590 8629 3612
rect 8656 3590 8657 3606
rect 8672 3590 8685 3750
rect 8715 3646 8728 3750
rect 8773 3728 8774 3738
rect 8789 3728 8802 3738
rect 8773 3724 8802 3728
rect 8807 3724 8837 3750
rect 8855 3736 8871 3738
rect 8943 3736 8996 3750
rect 8944 3734 9008 3736
rect 9051 3734 9066 3750
rect 9115 3747 9145 3750
rect 9115 3744 9151 3747
rect 9081 3736 9097 3738
rect 8855 3724 8870 3728
rect 8773 3722 8870 3724
rect 8898 3722 9066 3734
rect 9082 3724 9097 3728
rect 9115 3725 9154 3744
rect 9173 3738 9180 3739
rect 9179 3731 9180 3738
rect 9163 3728 9164 3731
rect 9179 3728 9192 3731
rect 9115 3724 9145 3725
rect 9154 3724 9160 3725
rect 9163 3724 9192 3728
rect 9082 3723 9192 3724
rect 9082 3722 9198 3723
rect 8757 3714 8808 3722
rect 8757 3702 8782 3714
rect 8789 3702 8808 3714
rect 8839 3714 8889 3722
rect 8839 3706 8855 3714
rect 8862 3712 8889 3714
rect 8898 3712 9119 3722
rect 8862 3702 9119 3712
rect 9148 3714 9198 3722
rect 9148 3705 9164 3714
rect 8757 3694 8808 3702
rect 8855 3694 9119 3702
rect 9145 3702 9164 3705
rect 9171 3702 9198 3714
rect 9145 3694 9198 3702
rect 8773 3686 8774 3694
rect 8789 3686 8802 3694
rect 8773 3678 8789 3686
rect 8770 3671 8789 3674
rect 8770 3662 8792 3671
rect 8743 3652 8792 3662
rect 8743 3646 8773 3652
rect 8792 3647 8797 3652
rect 8715 3630 8789 3646
rect 8807 3638 8837 3694
rect 8872 3684 9080 3694
rect 9115 3690 9160 3694
rect 9163 3693 9164 3694
rect 9179 3693 9192 3694
rect 8898 3654 9087 3684
rect 8913 3651 9087 3654
rect 8906 3648 9087 3651
rect 8715 3628 8728 3630
rect 8743 3628 8777 3630
rect 8715 3612 8789 3628
rect 8816 3624 8829 3638
rect 8844 3624 8860 3640
rect 8906 3635 8917 3648
rect 8699 3590 8700 3606
rect 8715 3590 8728 3612
rect 8743 3590 8773 3612
rect 8816 3608 8878 3624
rect 8906 3617 8917 3633
rect 8922 3628 8932 3648
rect 8942 3628 8956 3648
rect 8959 3635 8968 3648
rect 8984 3635 8993 3648
rect 8922 3617 8956 3628
rect 8959 3617 8968 3633
rect 8984 3617 8993 3633
rect 9000 3628 9010 3648
rect 9020 3628 9034 3648
rect 9035 3635 9046 3648
rect 9000 3617 9034 3628
rect 9035 3617 9046 3633
rect 9092 3624 9108 3640
rect 9115 3638 9145 3690
rect 9179 3686 9180 3693
rect 9164 3678 9180 3686
rect 9151 3646 9164 3665
rect 9179 3646 9209 3662
rect 9151 3630 9225 3646
rect 9151 3628 9164 3630
rect 9179 3628 9213 3630
rect 8816 3606 8829 3608
rect 8844 3606 8878 3608
rect 8816 3590 8878 3606
rect 8922 3601 8938 3604
rect 9000 3601 9030 3612
rect 9078 3608 9124 3624
rect 9151 3612 9225 3628
rect 9078 3606 9112 3608
rect 9077 3590 9124 3606
rect 9151 3590 9164 3612
rect 9179 3590 9209 3612
rect 9236 3590 9237 3606
rect 9252 3590 9265 3750
rect 7496 3582 7531 3590
rect 7496 3556 7497 3582
rect 7504 3556 7531 3582
rect 7439 3538 7469 3552
rect 7496 3548 7531 3556
rect 7533 3582 7574 3590
rect 7533 3556 7548 3582
rect 7555 3556 7574 3582
rect 7638 3578 7700 3590
rect 7712 3578 7787 3590
rect 7845 3578 7920 3590
rect 7932 3578 7963 3590
rect 7969 3578 8004 3590
rect 7638 3576 7800 3578
rect 7533 3548 7574 3556
rect 7656 3552 7669 3576
rect 7684 3574 7699 3576
rect 7496 3538 7525 3548
rect 7539 3538 7568 3548
rect 7583 3538 7613 3552
rect 7656 3538 7699 3552
rect 7723 3549 7730 3556
rect 7733 3552 7800 3576
rect 7832 3576 8004 3578
rect 7802 3554 7830 3558
rect 7832 3554 7912 3576
rect 7933 3574 7948 3576
rect 7802 3552 7912 3554
rect 7733 3548 7912 3552
rect 7706 3538 7736 3548
rect 7738 3538 7891 3548
rect 7899 3538 7929 3548
rect 7933 3538 7963 3552
rect 7991 3538 8004 3576
rect 8076 3582 8111 3590
rect 8076 3556 8077 3582
rect 8084 3556 8111 3582
rect 8019 3538 8049 3552
rect 8076 3548 8111 3556
rect 8113 3582 8154 3590
rect 8113 3556 8128 3582
rect 8135 3556 8154 3582
rect 8218 3578 8280 3590
rect 8292 3578 8367 3590
rect 8425 3578 8500 3590
rect 8512 3578 8543 3590
rect 8549 3578 8584 3590
rect 8218 3576 8380 3578
rect 8113 3548 8154 3556
rect 8236 3552 8249 3576
rect 8264 3574 8279 3576
rect 8076 3538 8077 3548
rect 8092 3538 8105 3548
rect 8119 3538 8120 3548
rect 8135 3538 8148 3548
rect 8163 3538 8193 3552
rect 8236 3538 8279 3552
rect 8303 3549 8310 3556
rect 8313 3552 8380 3576
rect 8412 3576 8584 3578
rect 8382 3554 8410 3558
rect 8412 3554 8492 3576
rect 8513 3574 8528 3576
rect 8382 3552 8492 3554
rect 8313 3548 8492 3552
rect 8286 3538 8316 3548
rect 8318 3538 8471 3548
rect 8479 3538 8509 3548
rect 8513 3538 8543 3552
rect 8571 3538 8584 3576
rect 8656 3582 8691 3590
rect 8656 3556 8657 3582
rect 8664 3556 8691 3582
rect 8599 3538 8629 3552
rect 8656 3548 8691 3556
rect 8693 3582 8734 3590
rect 8693 3556 8708 3582
rect 8715 3556 8734 3582
rect 8798 3578 8860 3590
rect 8872 3578 8947 3590
rect 9005 3578 9080 3590
rect 9092 3578 9123 3590
rect 9129 3578 9164 3590
rect 8798 3576 8960 3578
rect 8693 3548 8734 3556
rect 8816 3552 8829 3576
rect 8844 3574 8859 3576
rect 8656 3538 8657 3548
rect 8672 3538 8685 3548
rect 8699 3538 8700 3548
rect 8715 3538 8728 3548
rect 8743 3538 8773 3552
rect 8816 3538 8859 3552
rect 8883 3549 8890 3556
rect 8893 3552 8960 3576
rect 8992 3576 9164 3578
rect 8962 3554 8990 3558
rect 8992 3554 9072 3576
rect 9093 3574 9108 3576
rect 8962 3552 9072 3554
rect 8893 3548 9072 3552
rect 8866 3538 8896 3548
rect 8898 3538 9051 3548
rect 9059 3538 9089 3548
rect 9093 3538 9123 3552
rect 9151 3538 9164 3576
rect 9236 3582 9271 3590
rect 9236 3556 9237 3582
rect 9244 3556 9271 3582
rect 9179 3538 9209 3552
rect 9236 3548 9271 3556
rect 9236 3538 9237 3548
rect 9252 3538 9265 3548
rect -1 3532 9265 3538
rect 0 3524 9265 3532
rect 15 3494 28 3524
rect 43 3510 73 3524
rect 116 3510 159 3524
rect 166 3510 386 3524
rect 393 3510 423 3524
rect 83 3496 98 3508
rect 117 3496 130 3510
rect 198 3506 351 3510
rect 80 3494 102 3496
rect 180 3494 372 3506
rect 451 3494 464 3524
rect 479 3510 509 3524
rect 546 3494 565 3524
rect 580 3494 586 3524
rect 595 3494 608 3524
rect 623 3510 653 3524
rect 696 3510 739 3524
rect 746 3510 966 3524
rect 973 3510 1003 3524
rect 663 3496 678 3508
rect 697 3496 710 3510
rect 778 3506 931 3510
rect 660 3494 682 3496
rect 760 3494 952 3506
rect 1031 3494 1044 3524
rect 1059 3510 1089 3524
rect 1126 3494 1145 3524
rect 1160 3494 1166 3524
rect 1175 3494 1188 3524
rect 1203 3510 1233 3524
rect 1276 3510 1319 3524
rect 1326 3510 1546 3524
rect 1553 3510 1583 3524
rect 1243 3496 1258 3508
rect 1277 3496 1290 3510
rect 1358 3506 1511 3510
rect 1240 3494 1262 3496
rect 1340 3494 1532 3506
rect 1611 3494 1624 3524
rect 1639 3510 1669 3524
rect 1706 3494 1725 3524
rect 1740 3494 1746 3524
rect 1755 3494 1768 3524
rect 1783 3510 1813 3524
rect 1856 3510 1899 3524
rect 1906 3510 2126 3524
rect 2133 3510 2163 3524
rect 1823 3496 1838 3508
rect 1857 3496 1870 3510
rect 1938 3506 2091 3510
rect 1820 3494 1842 3496
rect 1920 3494 2112 3506
rect 2191 3494 2204 3524
rect 2219 3510 2249 3524
rect 2286 3494 2305 3524
rect 2320 3494 2326 3524
rect 2335 3494 2348 3524
rect 2363 3510 2393 3524
rect 2436 3510 2479 3524
rect 2486 3510 2706 3524
rect 2713 3510 2743 3524
rect 2403 3496 2418 3508
rect 2437 3496 2450 3510
rect 2518 3506 2671 3510
rect 2400 3494 2422 3496
rect 2500 3494 2692 3506
rect 2771 3494 2784 3524
rect 2799 3510 2829 3524
rect 2866 3494 2885 3524
rect 2900 3494 2906 3524
rect 2915 3494 2928 3524
rect 2943 3510 2973 3524
rect 3016 3510 3059 3524
rect 3066 3510 3286 3524
rect 3293 3510 3323 3524
rect 2983 3496 2998 3508
rect 3017 3496 3030 3510
rect 3098 3506 3251 3510
rect 2980 3494 3002 3496
rect 3080 3494 3272 3506
rect 3351 3494 3364 3524
rect 3379 3510 3409 3524
rect 3446 3494 3465 3524
rect 3480 3494 3486 3524
rect 3495 3494 3508 3524
rect 3523 3510 3553 3524
rect 3596 3510 3639 3524
rect 3646 3510 3866 3524
rect 3873 3510 3903 3524
rect 3563 3496 3578 3508
rect 3597 3496 3610 3510
rect 3678 3506 3831 3510
rect 3560 3494 3582 3496
rect 3660 3494 3852 3506
rect 3931 3494 3944 3524
rect 3959 3510 3989 3524
rect 4026 3494 4045 3524
rect 4060 3494 4066 3524
rect 4075 3494 4088 3524
rect 4103 3510 4133 3524
rect 4176 3510 4219 3524
rect 4226 3510 4446 3524
rect 4453 3510 4483 3524
rect 4143 3496 4158 3508
rect 4177 3496 4190 3510
rect 4258 3506 4411 3510
rect 4140 3494 4162 3496
rect 4240 3494 4432 3506
rect 4511 3494 4524 3524
rect 4539 3510 4569 3524
rect 4606 3494 4625 3524
rect 4640 3494 4646 3524
rect 4655 3494 4668 3524
rect 4683 3510 4713 3524
rect 4756 3510 4799 3524
rect 4806 3510 5026 3524
rect 5033 3510 5063 3524
rect 4723 3496 4738 3508
rect 4757 3496 4770 3510
rect 4838 3506 4991 3510
rect 4720 3494 4742 3496
rect 4820 3494 5012 3506
rect 5091 3494 5104 3524
rect 5119 3510 5149 3524
rect 5186 3494 5205 3524
rect 5220 3494 5226 3524
rect 5235 3494 5248 3524
rect 5263 3510 5293 3524
rect 5336 3510 5379 3524
rect 5386 3510 5606 3524
rect 5613 3510 5643 3524
rect 5303 3496 5318 3508
rect 5337 3496 5350 3510
rect 5418 3506 5571 3510
rect 5300 3494 5322 3496
rect 5400 3494 5592 3506
rect 5671 3494 5684 3524
rect 5699 3510 5729 3524
rect 5766 3494 5785 3524
rect 5800 3494 5806 3524
rect 5815 3494 5828 3524
rect 5843 3510 5873 3524
rect 5916 3510 5959 3524
rect 5966 3510 6186 3524
rect 6193 3510 6223 3524
rect 5883 3496 5898 3508
rect 5917 3496 5930 3510
rect 5998 3506 6151 3510
rect 5880 3494 5902 3496
rect 5980 3494 6172 3506
rect 6251 3494 6264 3524
rect 6279 3510 6309 3524
rect 6346 3494 6365 3524
rect 6380 3494 6386 3524
rect 6395 3494 6408 3524
rect 6423 3510 6453 3524
rect 6496 3510 6539 3524
rect 6546 3510 6766 3524
rect 6773 3510 6803 3524
rect 6463 3496 6478 3508
rect 6497 3496 6510 3510
rect 6578 3506 6731 3510
rect 6460 3494 6482 3496
rect 6560 3494 6752 3506
rect 6831 3494 6844 3524
rect 6859 3510 6889 3524
rect 6926 3494 6945 3524
rect 6960 3494 6966 3524
rect 6975 3494 6988 3524
rect 7003 3510 7033 3524
rect 7076 3510 7119 3524
rect 7126 3510 7346 3524
rect 7353 3510 7383 3524
rect 7043 3496 7058 3508
rect 7077 3496 7090 3510
rect 7158 3506 7311 3510
rect 7040 3494 7062 3496
rect 7140 3494 7332 3506
rect 7411 3494 7424 3524
rect 7439 3510 7469 3524
rect 7506 3494 7525 3524
rect 7540 3494 7546 3524
rect 7555 3494 7568 3524
rect 7583 3506 7613 3524
rect 7656 3510 7670 3524
rect 7706 3510 7926 3524
rect 7657 3508 7670 3510
rect 7623 3496 7638 3508
rect 7620 3494 7642 3496
rect 7647 3494 7677 3508
rect 7738 3506 7891 3510
rect 7720 3494 7912 3506
rect 7955 3494 7985 3508
rect 7991 3494 8004 3524
rect 8019 3506 8049 3524
rect 8092 3494 8105 3524
rect 8135 3494 8148 3524
rect 8163 3506 8193 3524
rect 8236 3510 8250 3524
rect 8286 3510 8506 3524
rect 8237 3508 8250 3510
rect 8203 3496 8218 3508
rect 8200 3494 8222 3496
rect 8227 3494 8257 3508
rect 8318 3506 8471 3510
rect 8300 3494 8492 3506
rect 8535 3494 8565 3508
rect 8571 3494 8584 3524
rect 8599 3506 8629 3524
rect 8672 3494 8685 3524
rect 8715 3494 8728 3524
rect 8743 3506 8773 3524
rect 8816 3510 8830 3524
rect 8866 3510 9086 3524
rect 8817 3508 8830 3510
rect 8783 3496 8798 3508
rect 8780 3494 8802 3496
rect 8807 3494 8837 3508
rect 8898 3506 9051 3510
rect 8880 3494 9072 3506
rect 9115 3494 9145 3508
rect 9151 3494 9164 3524
rect 9179 3506 9209 3524
rect 9252 3494 9265 3524
rect 0 3480 9265 3494
rect 15 3410 28 3480
rect 80 3476 102 3480
rect 73 3454 102 3468
rect 155 3454 171 3468
rect 209 3464 215 3466
rect 222 3464 330 3480
rect 337 3464 343 3466
rect 351 3464 366 3480
rect 432 3474 451 3477
rect 73 3452 171 3454
rect 198 3452 366 3464
rect 381 3454 397 3468
rect 432 3455 454 3474
rect 464 3468 480 3469
rect 463 3466 480 3468
rect 464 3461 480 3466
rect 454 3454 460 3455
rect 463 3454 492 3461
rect 381 3453 492 3454
rect 381 3452 498 3453
rect 57 3444 108 3452
rect 155 3444 189 3452
rect 57 3432 82 3444
rect 89 3432 108 3444
rect 162 3442 189 3444
rect 198 3442 419 3452
rect 454 3449 460 3452
rect 162 3438 419 3442
rect 57 3424 108 3432
rect 155 3424 419 3438
rect 463 3444 498 3452
rect 9 3376 28 3410
rect 73 3416 102 3424
rect 73 3410 90 3416
rect 73 3408 107 3410
rect 155 3408 171 3424
rect 172 3414 380 3424
rect 381 3414 397 3424
rect 445 3420 460 3435
rect 463 3432 464 3444
rect 471 3432 498 3444
rect 463 3424 498 3432
rect 463 3423 492 3424
rect 183 3410 397 3414
rect 198 3408 397 3410
rect 432 3410 445 3420
rect 463 3410 480 3423
rect 432 3408 480 3410
rect 74 3404 107 3408
rect 70 3402 107 3404
rect 70 3401 137 3402
rect 70 3396 101 3401
rect 107 3396 137 3401
rect 70 3392 137 3396
rect 43 3389 137 3392
rect 43 3382 92 3389
rect 43 3376 73 3382
rect 92 3377 97 3382
rect 9 3360 89 3376
rect 101 3368 137 3389
rect 198 3384 387 3408
rect 432 3407 479 3408
rect 445 3402 479 3407
rect 213 3381 387 3384
rect 206 3378 387 3381
rect 415 3401 479 3402
rect 9 3358 28 3360
rect 43 3358 77 3360
rect 9 3342 89 3358
rect 9 3336 28 3342
rect -1 3320 28 3336
rect 43 3326 73 3342
rect 101 3320 107 3368
rect 110 3362 129 3368
rect 144 3362 174 3370
rect 110 3354 174 3362
rect 110 3338 190 3354
rect 206 3347 268 3378
rect 284 3347 346 3378
rect 415 3376 464 3401
rect 479 3376 509 3392
rect 378 3362 408 3370
rect 415 3368 525 3376
rect 378 3354 423 3362
rect 110 3336 129 3338
rect 144 3336 190 3338
rect 110 3320 190 3336
rect 217 3334 252 3347
rect 293 3344 330 3347
rect 293 3342 335 3344
rect 222 3331 252 3334
rect 231 3327 238 3331
rect 238 3326 239 3327
rect 197 3320 207 3326
rect -7 3312 34 3320
rect -7 3286 8 3312
rect 15 3286 34 3312
rect 98 3308 129 3320
rect 144 3308 247 3320
rect 259 3310 285 3336
rect 300 3331 330 3342
rect 362 3338 424 3354
rect 362 3336 408 3338
rect 362 3320 424 3336
rect 436 3320 442 3368
rect 445 3360 525 3368
rect 445 3358 464 3360
rect 479 3358 513 3360
rect 445 3342 525 3358
rect 445 3320 464 3342
rect 479 3326 509 3342
rect 537 3336 543 3410
rect 546 3336 565 3480
rect 580 3336 586 3480
rect 595 3410 608 3480
rect 660 3476 682 3480
rect 653 3454 682 3468
rect 735 3454 751 3468
rect 789 3464 795 3466
rect 802 3464 910 3480
rect 917 3464 923 3466
rect 931 3464 946 3480
rect 1012 3474 1031 3477
rect 653 3452 751 3454
rect 778 3452 946 3464
rect 961 3454 977 3468
rect 1012 3455 1034 3474
rect 1044 3468 1060 3469
rect 1043 3466 1060 3468
rect 1044 3461 1060 3466
rect 1034 3454 1040 3455
rect 1043 3454 1072 3461
rect 961 3453 1072 3454
rect 961 3452 1078 3453
rect 637 3444 688 3452
rect 735 3444 769 3452
rect 637 3432 662 3444
rect 669 3432 688 3444
rect 742 3442 769 3444
rect 778 3442 999 3452
rect 1034 3449 1040 3452
rect 742 3438 999 3442
rect 637 3424 688 3432
rect 735 3424 999 3438
rect 1043 3444 1078 3452
rect 589 3376 608 3410
rect 653 3416 682 3424
rect 653 3410 670 3416
rect 653 3408 687 3410
rect 735 3408 751 3424
rect 752 3414 960 3424
rect 961 3414 977 3424
rect 1025 3420 1040 3435
rect 1043 3432 1044 3444
rect 1051 3432 1078 3444
rect 1043 3424 1078 3432
rect 1043 3423 1072 3424
rect 763 3410 977 3414
rect 778 3408 977 3410
rect 1012 3410 1025 3420
rect 1043 3410 1060 3423
rect 1012 3408 1060 3410
rect 654 3404 687 3408
rect 650 3402 687 3404
rect 650 3401 717 3402
rect 650 3396 681 3401
rect 687 3396 717 3401
rect 650 3392 717 3396
rect 623 3389 717 3392
rect 623 3382 672 3389
rect 623 3376 653 3382
rect 672 3377 677 3382
rect 589 3360 669 3376
rect 681 3368 717 3389
rect 778 3384 967 3408
rect 1012 3407 1059 3408
rect 1025 3402 1059 3407
rect 793 3381 967 3384
rect 786 3378 967 3381
rect 995 3401 1059 3402
rect 589 3358 608 3360
rect 623 3358 657 3360
rect 589 3342 669 3358
rect 589 3336 608 3342
rect 305 3310 408 3320
rect 259 3308 408 3310
rect 429 3308 464 3320
rect 98 3306 260 3308
rect 110 3286 129 3306
rect 144 3304 174 3306
rect -7 3278 34 3286
rect 116 3282 129 3286
rect 181 3290 260 3306
rect 292 3306 464 3308
rect 292 3290 371 3306
rect 378 3304 408 3306
rect -1 3268 28 3278
rect 43 3268 73 3282
rect 116 3268 159 3282
rect 181 3278 371 3290
rect 436 3286 442 3306
rect 166 3268 196 3278
rect 197 3268 355 3278
rect 359 3268 389 3278
rect 393 3268 423 3282
rect 451 3268 464 3306
rect 536 3320 565 3336
rect 579 3320 608 3336
rect 623 3326 653 3342
rect 681 3320 687 3368
rect 690 3362 709 3368
rect 724 3362 754 3370
rect 690 3354 754 3362
rect 690 3338 770 3354
rect 786 3347 848 3378
rect 864 3347 926 3378
rect 995 3376 1044 3401
rect 1059 3376 1089 3392
rect 958 3362 988 3370
rect 995 3368 1105 3376
rect 958 3354 1003 3362
rect 690 3336 709 3338
rect 724 3336 770 3338
rect 690 3320 770 3336
rect 797 3334 832 3347
rect 873 3344 910 3347
rect 873 3342 915 3344
rect 802 3331 832 3334
rect 811 3327 818 3331
rect 818 3326 819 3327
rect 777 3320 787 3326
rect 536 3312 571 3320
rect 536 3286 537 3312
rect 544 3286 571 3312
rect 479 3268 509 3282
rect 536 3278 571 3286
rect 573 3312 614 3320
rect 573 3286 588 3312
rect 595 3286 614 3312
rect 678 3308 709 3320
rect 724 3308 827 3320
rect 839 3310 865 3336
rect 880 3331 910 3342
rect 942 3338 1004 3354
rect 942 3336 988 3338
rect 942 3320 1004 3336
rect 1016 3320 1022 3368
rect 1025 3360 1105 3368
rect 1025 3358 1044 3360
rect 1059 3358 1093 3360
rect 1025 3342 1105 3358
rect 1025 3320 1044 3342
rect 1059 3326 1089 3342
rect 1117 3336 1123 3410
rect 1126 3336 1145 3480
rect 1160 3336 1166 3480
rect 1175 3410 1188 3480
rect 1240 3476 1262 3480
rect 1233 3454 1262 3468
rect 1315 3454 1331 3468
rect 1369 3464 1375 3466
rect 1382 3464 1490 3480
rect 1497 3464 1503 3466
rect 1511 3464 1526 3480
rect 1592 3474 1611 3477
rect 1233 3452 1331 3454
rect 1358 3452 1526 3464
rect 1541 3454 1557 3468
rect 1592 3455 1614 3474
rect 1624 3468 1640 3469
rect 1623 3466 1640 3468
rect 1624 3461 1640 3466
rect 1614 3454 1620 3455
rect 1623 3454 1652 3461
rect 1541 3453 1652 3454
rect 1541 3452 1658 3453
rect 1217 3444 1268 3452
rect 1315 3444 1349 3452
rect 1217 3432 1242 3444
rect 1249 3432 1268 3444
rect 1322 3442 1349 3444
rect 1358 3442 1579 3452
rect 1614 3449 1620 3452
rect 1322 3438 1579 3442
rect 1217 3424 1268 3432
rect 1315 3424 1579 3438
rect 1623 3444 1658 3452
rect 1169 3376 1188 3410
rect 1233 3416 1262 3424
rect 1233 3410 1250 3416
rect 1233 3408 1267 3410
rect 1315 3408 1331 3424
rect 1332 3414 1540 3424
rect 1541 3414 1557 3424
rect 1605 3420 1620 3435
rect 1623 3432 1624 3444
rect 1631 3432 1658 3444
rect 1623 3424 1658 3432
rect 1623 3423 1652 3424
rect 1343 3410 1557 3414
rect 1358 3408 1557 3410
rect 1592 3410 1605 3420
rect 1623 3410 1640 3423
rect 1592 3408 1640 3410
rect 1234 3404 1267 3408
rect 1230 3402 1267 3404
rect 1230 3401 1297 3402
rect 1230 3396 1261 3401
rect 1267 3396 1297 3401
rect 1230 3392 1297 3396
rect 1203 3389 1297 3392
rect 1203 3382 1252 3389
rect 1203 3376 1233 3382
rect 1252 3377 1257 3382
rect 1169 3360 1249 3376
rect 1261 3368 1297 3389
rect 1358 3384 1547 3408
rect 1592 3407 1639 3408
rect 1605 3402 1639 3407
rect 1373 3381 1547 3384
rect 1366 3378 1547 3381
rect 1575 3401 1639 3402
rect 1169 3358 1188 3360
rect 1203 3358 1237 3360
rect 1169 3342 1249 3358
rect 1169 3336 1188 3342
rect 885 3310 988 3320
rect 839 3308 988 3310
rect 1009 3308 1044 3320
rect 678 3306 840 3308
rect 690 3286 709 3306
rect 724 3304 754 3306
rect 573 3278 614 3286
rect 696 3282 709 3286
rect 761 3290 840 3306
rect 872 3306 1044 3308
rect 872 3290 951 3306
rect 958 3304 988 3306
rect 536 3268 565 3278
rect 579 3268 608 3278
rect 623 3268 653 3282
rect 696 3268 739 3282
rect 761 3278 951 3290
rect 1016 3286 1022 3306
rect 746 3268 776 3278
rect 777 3268 935 3278
rect 939 3268 969 3278
rect 973 3268 1003 3282
rect 1031 3268 1044 3306
rect 1116 3320 1145 3336
rect 1159 3320 1188 3336
rect 1203 3326 1233 3342
rect 1261 3320 1267 3368
rect 1270 3362 1289 3368
rect 1304 3362 1334 3370
rect 1270 3354 1334 3362
rect 1270 3338 1350 3354
rect 1366 3347 1428 3378
rect 1444 3347 1506 3378
rect 1575 3376 1624 3401
rect 1639 3376 1669 3392
rect 1538 3362 1568 3370
rect 1575 3368 1685 3376
rect 1538 3354 1583 3362
rect 1270 3336 1289 3338
rect 1304 3336 1350 3338
rect 1270 3320 1350 3336
rect 1377 3334 1412 3347
rect 1453 3344 1490 3347
rect 1453 3342 1495 3344
rect 1382 3331 1412 3334
rect 1391 3327 1398 3331
rect 1398 3326 1399 3327
rect 1357 3320 1367 3326
rect 1116 3312 1151 3320
rect 1116 3286 1117 3312
rect 1124 3286 1151 3312
rect 1059 3268 1089 3282
rect 1116 3278 1151 3286
rect 1153 3312 1194 3320
rect 1153 3286 1168 3312
rect 1175 3286 1194 3312
rect 1258 3308 1289 3320
rect 1304 3308 1407 3320
rect 1419 3310 1445 3336
rect 1460 3331 1490 3342
rect 1522 3338 1584 3354
rect 1522 3336 1568 3338
rect 1522 3320 1584 3336
rect 1596 3320 1602 3368
rect 1605 3360 1685 3368
rect 1605 3358 1624 3360
rect 1639 3358 1673 3360
rect 1605 3342 1685 3358
rect 1605 3320 1624 3342
rect 1639 3326 1669 3342
rect 1697 3336 1703 3410
rect 1706 3336 1725 3480
rect 1740 3336 1746 3480
rect 1755 3410 1768 3480
rect 1820 3476 1842 3480
rect 1813 3454 1842 3468
rect 1895 3454 1911 3468
rect 1949 3464 1955 3466
rect 1962 3464 2070 3480
rect 2077 3464 2083 3466
rect 2091 3464 2106 3480
rect 2172 3474 2191 3477
rect 1813 3452 1911 3454
rect 1938 3452 2106 3464
rect 2121 3454 2137 3468
rect 2172 3455 2194 3474
rect 2204 3468 2220 3469
rect 2203 3466 2220 3468
rect 2204 3461 2220 3466
rect 2194 3454 2200 3455
rect 2203 3454 2232 3461
rect 2121 3453 2232 3454
rect 2121 3452 2238 3453
rect 1797 3444 1848 3452
rect 1895 3444 1929 3452
rect 1797 3432 1822 3444
rect 1829 3432 1848 3444
rect 1902 3442 1929 3444
rect 1938 3442 2159 3452
rect 2194 3449 2200 3452
rect 1902 3438 2159 3442
rect 1797 3424 1848 3432
rect 1895 3424 2159 3438
rect 2203 3444 2238 3452
rect 1749 3376 1768 3410
rect 1813 3416 1842 3424
rect 1813 3410 1830 3416
rect 1813 3408 1847 3410
rect 1895 3408 1911 3424
rect 1912 3414 2120 3424
rect 2121 3414 2137 3424
rect 2185 3420 2200 3435
rect 2203 3432 2204 3444
rect 2211 3432 2238 3444
rect 2203 3424 2238 3432
rect 2203 3423 2232 3424
rect 1923 3410 2137 3414
rect 1938 3408 2137 3410
rect 2172 3410 2185 3420
rect 2203 3410 2220 3423
rect 2172 3408 2220 3410
rect 1814 3404 1847 3408
rect 1810 3402 1847 3404
rect 1810 3401 1877 3402
rect 1810 3396 1841 3401
rect 1847 3396 1877 3401
rect 1810 3392 1877 3396
rect 1783 3389 1877 3392
rect 1783 3382 1832 3389
rect 1783 3376 1813 3382
rect 1832 3377 1837 3382
rect 1749 3360 1829 3376
rect 1841 3368 1877 3389
rect 1938 3384 2127 3408
rect 2172 3407 2219 3408
rect 2185 3402 2219 3407
rect 1953 3381 2127 3384
rect 1946 3378 2127 3381
rect 2155 3401 2219 3402
rect 1749 3358 1768 3360
rect 1783 3358 1817 3360
rect 1749 3342 1829 3358
rect 1749 3336 1768 3342
rect 1465 3310 1568 3320
rect 1419 3308 1568 3310
rect 1589 3308 1624 3320
rect 1258 3306 1420 3308
rect 1270 3286 1289 3306
rect 1304 3304 1334 3306
rect 1153 3278 1194 3286
rect 1276 3282 1289 3286
rect 1341 3290 1420 3306
rect 1452 3306 1624 3308
rect 1452 3290 1531 3306
rect 1538 3304 1568 3306
rect 1116 3268 1145 3278
rect 1159 3268 1188 3278
rect 1203 3268 1233 3282
rect 1276 3268 1319 3282
rect 1341 3278 1531 3290
rect 1596 3286 1602 3306
rect 1326 3268 1356 3278
rect 1357 3268 1515 3278
rect 1519 3268 1549 3278
rect 1553 3268 1583 3282
rect 1611 3268 1624 3306
rect 1696 3320 1725 3336
rect 1739 3320 1768 3336
rect 1783 3326 1813 3342
rect 1841 3320 1847 3368
rect 1850 3362 1869 3368
rect 1884 3362 1914 3370
rect 1850 3354 1914 3362
rect 1850 3338 1930 3354
rect 1946 3347 2008 3378
rect 2024 3347 2086 3378
rect 2155 3376 2204 3401
rect 2219 3376 2249 3392
rect 2118 3362 2148 3370
rect 2155 3368 2265 3376
rect 2118 3354 2163 3362
rect 1850 3336 1869 3338
rect 1884 3336 1930 3338
rect 1850 3320 1930 3336
rect 1957 3334 1992 3347
rect 2033 3344 2070 3347
rect 2033 3342 2075 3344
rect 1962 3331 1992 3334
rect 1971 3327 1978 3331
rect 1978 3326 1979 3327
rect 1937 3320 1947 3326
rect 1696 3312 1731 3320
rect 1696 3286 1697 3312
rect 1704 3286 1731 3312
rect 1639 3268 1669 3282
rect 1696 3278 1731 3286
rect 1733 3312 1774 3320
rect 1733 3286 1748 3312
rect 1755 3286 1774 3312
rect 1838 3308 1869 3320
rect 1884 3308 1987 3320
rect 1999 3310 2025 3336
rect 2040 3331 2070 3342
rect 2102 3338 2164 3354
rect 2102 3336 2148 3338
rect 2102 3320 2164 3336
rect 2176 3320 2182 3368
rect 2185 3360 2265 3368
rect 2185 3358 2204 3360
rect 2219 3358 2253 3360
rect 2185 3342 2265 3358
rect 2185 3320 2204 3342
rect 2219 3326 2249 3342
rect 2277 3336 2283 3410
rect 2286 3336 2305 3480
rect 2320 3336 2326 3480
rect 2335 3410 2348 3480
rect 2400 3476 2422 3480
rect 2393 3454 2422 3468
rect 2475 3454 2491 3468
rect 2529 3464 2535 3466
rect 2542 3464 2650 3480
rect 2657 3464 2663 3466
rect 2671 3464 2686 3480
rect 2752 3474 2771 3477
rect 2393 3452 2491 3454
rect 2518 3452 2686 3464
rect 2701 3454 2717 3468
rect 2752 3455 2774 3474
rect 2784 3468 2800 3469
rect 2783 3466 2800 3468
rect 2784 3461 2800 3466
rect 2774 3454 2780 3455
rect 2783 3454 2812 3461
rect 2701 3453 2812 3454
rect 2701 3452 2818 3453
rect 2377 3444 2428 3452
rect 2475 3444 2509 3452
rect 2377 3432 2402 3444
rect 2409 3432 2428 3444
rect 2482 3442 2509 3444
rect 2518 3442 2739 3452
rect 2774 3449 2780 3452
rect 2482 3438 2739 3442
rect 2377 3424 2428 3432
rect 2475 3424 2739 3438
rect 2783 3444 2818 3452
rect 2329 3376 2348 3410
rect 2393 3416 2422 3424
rect 2393 3410 2410 3416
rect 2393 3408 2427 3410
rect 2475 3408 2491 3424
rect 2492 3414 2700 3424
rect 2701 3414 2717 3424
rect 2765 3420 2780 3435
rect 2783 3432 2784 3444
rect 2791 3432 2818 3444
rect 2783 3424 2818 3432
rect 2783 3423 2812 3424
rect 2503 3410 2717 3414
rect 2518 3408 2717 3410
rect 2752 3410 2765 3420
rect 2783 3410 2800 3423
rect 2752 3408 2800 3410
rect 2394 3404 2427 3408
rect 2390 3402 2427 3404
rect 2390 3401 2457 3402
rect 2390 3396 2421 3401
rect 2427 3396 2457 3401
rect 2390 3392 2457 3396
rect 2363 3389 2457 3392
rect 2363 3382 2412 3389
rect 2363 3376 2393 3382
rect 2412 3377 2417 3382
rect 2329 3360 2409 3376
rect 2421 3368 2457 3389
rect 2518 3384 2707 3408
rect 2752 3407 2799 3408
rect 2765 3402 2799 3407
rect 2533 3381 2707 3384
rect 2526 3378 2707 3381
rect 2735 3401 2799 3402
rect 2329 3358 2348 3360
rect 2363 3358 2397 3360
rect 2329 3342 2409 3358
rect 2329 3336 2348 3342
rect 2045 3310 2148 3320
rect 1999 3308 2148 3310
rect 2169 3308 2204 3320
rect 1838 3306 2000 3308
rect 1850 3286 1869 3306
rect 1884 3304 1914 3306
rect 1733 3278 1774 3286
rect 1856 3282 1869 3286
rect 1921 3290 2000 3306
rect 2032 3306 2204 3308
rect 2032 3290 2111 3306
rect 2118 3304 2148 3306
rect 1696 3268 1725 3278
rect 1739 3268 1768 3278
rect 1783 3268 1813 3282
rect 1856 3268 1899 3282
rect 1921 3278 2111 3290
rect 2176 3286 2182 3306
rect 1906 3268 1936 3278
rect 1937 3268 2095 3278
rect 2099 3268 2129 3278
rect 2133 3268 2163 3282
rect 2191 3268 2204 3306
rect 2276 3320 2305 3336
rect 2319 3320 2348 3336
rect 2363 3326 2393 3342
rect 2421 3320 2427 3368
rect 2430 3362 2449 3368
rect 2464 3362 2494 3370
rect 2430 3354 2494 3362
rect 2430 3338 2510 3354
rect 2526 3347 2588 3378
rect 2604 3347 2666 3378
rect 2735 3376 2784 3401
rect 2799 3376 2829 3392
rect 2698 3362 2728 3370
rect 2735 3368 2845 3376
rect 2698 3354 2743 3362
rect 2430 3336 2449 3338
rect 2464 3336 2510 3338
rect 2430 3320 2510 3336
rect 2537 3334 2572 3347
rect 2613 3344 2650 3347
rect 2613 3342 2655 3344
rect 2542 3331 2572 3334
rect 2551 3327 2558 3331
rect 2558 3326 2559 3327
rect 2517 3320 2527 3326
rect 2276 3312 2311 3320
rect 2276 3286 2277 3312
rect 2284 3286 2311 3312
rect 2219 3268 2249 3282
rect 2276 3278 2311 3286
rect 2313 3312 2354 3320
rect 2313 3286 2328 3312
rect 2335 3286 2354 3312
rect 2418 3308 2449 3320
rect 2464 3308 2567 3320
rect 2579 3310 2605 3336
rect 2620 3331 2650 3342
rect 2682 3338 2744 3354
rect 2682 3336 2728 3338
rect 2682 3320 2744 3336
rect 2756 3320 2762 3368
rect 2765 3360 2845 3368
rect 2765 3358 2784 3360
rect 2799 3358 2833 3360
rect 2765 3342 2845 3358
rect 2765 3320 2784 3342
rect 2799 3326 2829 3342
rect 2857 3336 2863 3410
rect 2866 3336 2885 3480
rect 2900 3336 2906 3480
rect 2915 3410 2928 3480
rect 2980 3476 3002 3480
rect 2973 3454 3002 3468
rect 3055 3454 3071 3468
rect 3109 3464 3115 3466
rect 3122 3464 3230 3480
rect 3237 3464 3243 3466
rect 3251 3464 3266 3480
rect 3332 3474 3351 3477
rect 2973 3452 3071 3454
rect 3098 3452 3266 3464
rect 3281 3454 3297 3468
rect 3332 3455 3354 3474
rect 3364 3468 3380 3469
rect 3363 3466 3380 3468
rect 3364 3461 3380 3466
rect 3354 3454 3360 3455
rect 3363 3454 3392 3461
rect 3281 3453 3392 3454
rect 3281 3452 3398 3453
rect 2957 3444 3008 3452
rect 3055 3444 3089 3452
rect 2957 3432 2982 3444
rect 2989 3432 3008 3444
rect 3062 3442 3089 3444
rect 3098 3442 3319 3452
rect 3354 3449 3360 3452
rect 3062 3438 3319 3442
rect 2957 3424 3008 3432
rect 3055 3424 3319 3438
rect 3363 3444 3398 3452
rect 2909 3376 2928 3410
rect 2973 3416 3002 3424
rect 2973 3410 2990 3416
rect 2973 3408 3007 3410
rect 3055 3408 3071 3424
rect 3072 3414 3280 3424
rect 3281 3414 3297 3424
rect 3345 3420 3360 3435
rect 3363 3432 3364 3444
rect 3371 3432 3398 3444
rect 3363 3424 3398 3432
rect 3363 3423 3392 3424
rect 3083 3410 3297 3414
rect 3098 3408 3297 3410
rect 3332 3410 3345 3420
rect 3363 3410 3380 3423
rect 3332 3408 3380 3410
rect 2974 3404 3007 3408
rect 2970 3402 3007 3404
rect 2970 3401 3037 3402
rect 2970 3396 3001 3401
rect 3007 3396 3037 3401
rect 2970 3392 3037 3396
rect 2943 3389 3037 3392
rect 2943 3382 2992 3389
rect 2943 3376 2973 3382
rect 2992 3377 2997 3382
rect 2909 3360 2989 3376
rect 3001 3368 3037 3389
rect 3098 3384 3287 3408
rect 3332 3407 3379 3408
rect 3345 3402 3379 3407
rect 3113 3381 3287 3384
rect 3106 3378 3287 3381
rect 3315 3401 3379 3402
rect 2909 3358 2928 3360
rect 2943 3358 2977 3360
rect 2909 3342 2989 3358
rect 2909 3336 2928 3342
rect 2625 3310 2728 3320
rect 2579 3308 2728 3310
rect 2749 3308 2784 3320
rect 2418 3306 2580 3308
rect 2430 3286 2449 3306
rect 2464 3304 2494 3306
rect 2313 3278 2354 3286
rect 2436 3282 2449 3286
rect 2501 3290 2580 3306
rect 2612 3306 2784 3308
rect 2612 3290 2691 3306
rect 2698 3304 2728 3306
rect 2276 3268 2305 3278
rect 2319 3268 2348 3278
rect 2363 3268 2393 3282
rect 2436 3268 2479 3282
rect 2501 3278 2691 3290
rect 2756 3286 2762 3306
rect 2486 3268 2516 3278
rect 2517 3268 2675 3278
rect 2679 3268 2709 3278
rect 2713 3268 2743 3282
rect 2771 3268 2784 3306
rect 2856 3320 2885 3336
rect 2899 3320 2928 3336
rect 2943 3326 2973 3342
rect 3001 3320 3007 3368
rect 3010 3362 3029 3368
rect 3044 3362 3074 3370
rect 3010 3354 3074 3362
rect 3010 3338 3090 3354
rect 3106 3347 3168 3378
rect 3184 3347 3246 3378
rect 3315 3376 3364 3401
rect 3379 3376 3409 3392
rect 3278 3362 3308 3370
rect 3315 3368 3425 3376
rect 3278 3354 3323 3362
rect 3010 3336 3029 3338
rect 3044 3336 3090 3338
rect 3010 3320 3090 3336
rect 3117 3334 3152 3347
rect 3193 3344 3230 3347
rect 3193 3342 3235 3344
rect 3122 3331 3152 3334
rect 3131 3327 3138 3331
rect 3138 3326 3139 3327
rect 3097 3320 3107 3326
rect 2856 3312 2891 3320
rect 2856 3286 2857 3312
rect 2864 3286 2891 3312
rect 2799 3268 2829 3282
rect 2856 3278 2891 3286
rect 2893 3312 2934 3320
rect 2893 3286 2908 3312
rect 2915 3286 2934 3312
rect 2998 3308 3029 3320
rect 3044 3308 3147 3320
rect 3159 3310 3185 3336
rect 3200 3331 3230 3342
rect 3262 3338 3324 3354
rect 3262 3336 3308 3338
rect 3262 3320 3324 3336
rect 3336 3320 3342 3368
rect 3345 3360 3425 3368
rect 3345 3358 3364 3360
rect 3379 3358 3413 3360
rect 3345 3342 3425 3358
rect 3345 3320 3364 3342
rect 3379 3326 3409 3342
rect 3437 3336 3443 3410
rect 3446 3336 3465 3480
rect 3480 3336 3486 3480
rect 3495 3410 3508 3480
rect 3560 3476 3582 3480
rect 3553 3454 3582 3468
rect 3635 3454 3651 3468
rect 3689 3464 3695 3466
rect 3702 3464 3810 3480
rect 3817 3464 3823 3466
rect 3831 3464 3846 3480
rect 3912 3474 3931 3477
rect 3553 3452 3651 3454
rect 3678 3452 3846 3464
rect 3861 3454 3877 3468
rect 3912 3455 3934 3474
rect 3944 3468 3960 3469
rect 3943 3466 3960 3468
rect 3944 3461 3960 3466
rect 3934 3454 3940 3455
rect 3943 3454 3972 3461
rect 3861 3453 3972 3454
rect 3861 3452 3978 3453
rect 3537 3444 3588 3452
rect 3635 3444 3669 3452
rect 3537 3432 3562 3444
rect 3569 3432 3588 3444
rect 3642 3442 3669 3444
rect 3678 3442 3899 3452
rect 3934 3449 3940 3452
rect 3642 3438 3899 3442
rect 3537 3424 3588 3432
rect 3635 3424 3899 3438
rect 3943 3444 3978 3452
rect 3489 3376 3508 3410
rect 3553 3416 3582 3424
rect 3553 3410 3570 3416
rect 3553 3408 3587 3410
rect 3635 3408 3651 3424
rect 3652 3414 3860 3424
rect 3861 3414 3877 3424
rect 3925 3420 3940 3435
rect 3943 3432 3944 3444
rect 3951 3432 3978 3444
rect 3943 3424 3978 3432
rect 3943 3423 3972 3424
rect 3663 3410 3877 3414
rect 3678 3408 3877 3410
rect 3912 3410 3925 3420
rect 3943 3410 3960 3423
rect 3912 3408 3960 3410
rect 3554 3404 3587 3408
rect 3550 3402 3587 3404
rect 3550 3401 3617 3402
rect 3550 3396 3581 3401
rect 3587 3396 3617 3401
rect 3550 3392 3617 3396
rect 3523 3389 3617 3392
rect 3523 3382 3572 3389
rect 3523 3376 3553 3382
rect 3572 3377 3577 3382
rect 3489 3360 3569 3376
rect 3581 3368 3617 3389
rect 3678 3384 3867 3408
rect 3912 3407 3959 3408
rect 3925 3402 3959 3407
rect 3693 3381 3867 3384
rect 3686 3378 3867 3381
rect 3895 3401 3959 3402
rect 3489 3358 3508 3360
rect 3523 3358 3557 3360
rect 3489 3342 3569 3358
rect 3489 3336 3508 3342
rect 3205 3310 3308 3320
rect 3159 3308 3308 3310
rect 3329 3308 3364 3320
rect 2998 3306 3160 3308
rect 3010 3286 3029 3306
rect 3044 3304 3074 3306
rect 2893 3278 2934 3286
rect 3016 3282 3029 3286
rect 3081 3290 3160 3306
rect 3192 3306 3364 3308
rect 3192 3290 3271 3306
rect 3278 3304 3308 3306
rect 2856 3268 2885 3278
rect 2899 3268 2928 3278
rect 2943 3268 2973 3282
rect 3016 3268 3059 3282
rect 3081 3278 3271 3290
rect 3336 3286 3342 3306
rect 3066 3268 3096 3278
rect 3097 3268 3255 3278
rect 3259 3268 3289 3278
rect 3293 3268 3323 3282
rect 3351 3268 3364 3306
rect 3436 3320 3465 3336
rect 3479 3320 3508 3336
rect 3523 3326 3553 3342
rect 3581 3320 3587 3368
rect 3590 3362 3609 3368
rect 3624 3362 3654 3370
rect 3590 3354 3654 3362
rect 3590 3338 3670 3354
rect 3686 3347 3748 3378
rect 3764 3347 3826 3378
rect 3895 3376 3944 3401
rect 3959 3376 3989 3392
rect 3858 3362 3888 3370
rect 3895 3368 4005 3376
rect 3858 3354 3903 3362
rect 3590 3336 3609 3338
rect 3624 3336 3670 3338
rect 3590 3320 3670 3336
rect 3697 3334 3732 3347
rect 3773 3344 3810 3347
rect 3773 3342 3815 3344
rect 3702 3331 3732 3334
rect 3711 3327 3718 3331
rect 3718 3326 3719 3327
rect 3677 3320 3687 3326
rect 3436 3312 3471 3320
rect 3436 3286 3437 3312
rect 3444 3286 3471 3312
rect 3379 3268 3409 3282
rect 3436 3278 3471 3286
rect 3473 3312 3514 3320
rect 3473 3286 3488 3312
rect 3495 3286 3514 3312
rect 3578 3308 3609 3320
rect 3624 3308 3727 3320
rect 3739 3310 3765 3336
rect 3780 3331 3810 3342
rect 3842 3338 3904 3354
rect 3842 3336 3888 3338
rect 3842 3320 3904 3336
rect 3916 3320 3922 3368
rect 3925 3360 4005 3368
rect 3925 3358 3944 3360
rect 3959 3358 3993 3360
rect 3925 3342 4005 3358
rect 3925 3320 3944 3342
rect 3959 3326 3989 3342
rect 4017 3336 4023 3410
rect 4026 3336 4045 3480
rect 4060 3336 4066 3480
rect 4075 3410 4088 3480
rect 4140 3476 4162 3480
rect 4133 3454 4162 3468
rect 4215 3454 4231 3468
rect 4269 3464 4275 3466
rect 4282 3464 4390 3480
rect 4397 3464 4403 3466
rect 4411 3464 4426 3480
rect 4492 3474 4511 3477
rect 4133 3452 4231 3454
rect 4258 3452 4426 3464
rect 4441 3454 4457 3468
rect 4492 3455 4514 3474
rect 4524 3468 4540 3469
rect 4523 3466 4540 3468
rect 4524 3461 4540 3466
rect 4514 3454 4520 3455
rect 4523 3454 4552 3461
rect 4441 3453 4552 3454
rect 4441 3452 4558 3453
rect 4117 3444 4168 3452
rect 4215 3444 4249 3452
rect 4117 3432 4142 3444
rect 4149 3432 4168 3444
rect 4222 3442 4249 3444
rect 4258 3442 4479 3452
rect 4514 3449 4520 3452
rect 4222 3438 4479 3442
rect 4117 3424 4168 3432
rect 4215 3424 4479 3438
rect 4523 3444 4558 3452
rect 4069 3376 4088 3410
rect 4133 3416 4162 3424
rect 4133 3410 4150 3416
rect 4133 3408 4167 3410
rect 4215 3408 4231 3424
rect 4232 3414 4440 3424
rect 4441 3414 4457 3424
rect 4505 3420 4520 3435
rect 4523 3432 4524 3444
rect 4531 3432 4558 3444
rect 4523 3424 4558 3432
rect 4523 3423 4552 3424
rect 4243 3410 4457 3414
rect 4258 3408 4457 3410
rect 4492 3410 4505 3420
rect 4523 3410 4540 3423
rect 4492 3408 4540 3410
rect 4134 3404 4167 3408
rect 4130 3402 4167 3404
rect 4130 3401 4197 3402
rect 4130 3396 4161 3401
rect 4167 3396 4197 3401
rect 4130 3392 4197 3396
rect 4103 3389 4197 3392
rect 4103 3382 4152 3389
rect 4103 3376 4133 3382
rect 4152 3377 4157 3382
rect 4069 3360 4149 3376
rect 4161 3368 4197 3389
rect 4258 3384 4447 3408
rect 4492 3407 4539 3408
rect 4505 3402 4539 3407
rect 4273 3381 4447 3384
rect 4266 3378 4447 3381
rect 4475 3401 4539 3402
rect 4069 3358 4088 3360
rect 4103 3358 4137 3360
rect 4069 3342 4149 3358
rect 4069 3336 4088 3342
rect 3785 3310 3888 3320
rect 3739 3308 3888 3310
rect 3909 3308 3944 3320
rect 3578 3306 3740 3308
rect 3590 3286 3609 3306
rect 3624 3304 3654 3306
rect 3473 3278 3514 3286
rect 3596 3282 3609 3286
rect 3661 3290 3740 3306
rect 3772 3306 3944 3308
rect 3772 3290 3851 3306
rect 3858 3304 3888 3306
rect 3436 3268 3465 3278
rect 3479 3268 3508 3278
rect 3523 3268 3553 3282
rect 3596 3268 3639 3282
rect 3661 3278 3851 3290
rect 3916 3286 3922 3306
rect 3646 3268 3676 3278
rect 3677 3268 3835 3278
rect 3839 3268 3869 3278
rect 3873 3268 3903 3282
rect 3931 3268 3944 3306
rect 4016 3320 4045 3336
rect 4059 3320 4088 3336
rect 4103 3326 4133 3342
rect 4161 3320 4167 3368
rect 4170 3362 4189 3368
rect 4204 3362 4234 3370
rect 4170 3354 4234 3362
rect 4170 3338 4250 3354
rect 4266 3347 4328 3378
rect 4344 3347 4406 3378
rect 4475 3376 4524 3401
rect 4539 3376 4569 3392
rect 4438 3362 4468 3370
rect 4475 3368 4585 3376
rect 4438 3354 4483 3362
rect 4170 3336 4189 3338
rect 4204 3336 4250 3338
rect 4170 3320 4250 3336
rect 4277 3334 4312 3347
rect 4353 3344 4390 3347
rect 4353 3342 4395 3344
rect 4282 3331 4312 3334
rect 4291 3327 4298 3331
rect 4298 3326 4299 3327
rect 4257 3320 4267 3326
rect 4016 3312 4051 3320
rect 4016 3286 4017 3312
rect 4024 3286 4051 3312
rect 3959 3268 3989 3282
rect 4016 3278 4051 3286
rect 4053 3312 4094 3320
rect 4053 3286 4068 3312
rect 4075 3286 4094 3312
rect 4158 3308 4189 3320
rect 4204 3308 4307 3320
rect 4319 3310 4345 3336
rect 4360 3331 4390 3342
rect 4422 3338 4484 3354
rect 4422 3336 4468 3338
rect 4422 3320 4484 3336
rect 4496 3320 4502 3368
rect 4505 3360 4585 3368
rect 4505 3358 4524 3360
rect 4539 3358 4573 3360
rect 4505 3342 4585 3358
rect 4505 3320 4524 3342
rect 4539 3326 4569 3342
rect 4597 3336 4603 3410
rect 4606 3336 4625 3480
rect 4640 3336 4646 3480
rect 4655 3410 4668 3480
rect 4720 3476 4742 3480
rect 4713 3454 4742 3468
rect 4795 3454 4811 3468
rect 4849 3464 4855 3466
rect 4862 3464 4970 3480
rect 4977 3464 4983 3466
rect 4991 3464 5006 3480
rect 5072 3474 5091 3477
rect 4713 3452 4811 3454
rect 4838 3452 5006 3464
rect 5021 3454 5037 3468
rect 5072 3455 5094 3474
rect 5104 3468 5120 3469
rect 5103 3466 5120 3468
rect 5104 3461 5120 3466
rect 5094 3454 5100 3455
rect 5103 3454 5132 3461
rect 5021 3453 5132 3454
rect 5021 3452 5138 3453
rect 4697 3444 4748 3452
rect 4795 3444 4829 3452
rect 4697 3432 4722 3444
rect 4729 3432 4748 3444
rect 4802 3442 4829 3444
rect 4838 3442 5059 3452
rect 5094 3449 5100 3452
rect 4802 3438 5059 3442
rect 4697 3424 4748 3432
rect 4795 3424 5059 3438
rect 5103 3444 5138 3452
rect 4649 3376 4668 3410
rect 4713 3416 4742 3424
rect 4713 3410 4730 3416
rect 4713 3408 4747 3410
rect 4795 3408 4811 3424
rect 4812 3414 5020 3424
rect 5021 3414 5037 3424
rect 5085 3420 5100 3435
rect 5103 3432 5104 3444
rect 5111 3432 5138 3444
rect 5103 3424 5138 3432
rect 5103 3423 5132 3424
rect 4823 3410 5037 3414
rect 4838 3408 5037 3410
rect 5072 3410 5085 3420
rect 5103 3410 5120 3423
rect 5072 3408 5120 3410
rect 4714 3404 4747 3408
rect 4710 3402 4747 3404
rect 4710 3401 4777 3402
rect 4710 3396 4741 3401
rect 4747 3396 4777 3401
rect 4710 3392 4777 3396
rect 4683 3389 4777 3392
rect 4683 3382 4732 3389
rect 4683 3376 4713 3382
rect 4732 3377 4737 3382
rect 4649 3360 4729 3376
rect 4741 3368 4777 3389
rect 4838 3384 5027 3408
rect 5072 3407 5119 3408
rect 5085 3402 5119 3407
rect 4853 3381 5027 3384
rect 4846 3378 5027 3381
rect 5055 3401 5119 3402
rect 4649 3358 4668 3360
rect 4683 3358 4717 3360
rect 4649 3342 4729 3358
rect 4649 3336 4668 3342
rect 4365 3310 4468 3320
rect 4319 3308 4468 3310
rect 4489 3308 4524 3320
rect 4158 3306 4320 3308
rect 4170 3286 4189 3306
rect 4204 3304 4234 3306
rect 4053 3278 4094 3286
rect 4176 3282 4189 3286
rect 4241 3290 4320 3306
rect 4352 3306 4524 3308
rect 4352 3290 4431 3306
rect 4438 3304 4468 3306
rect 4016 3268 4045 3278
rect 4059 3268 4088 3278
rect 4103 3268 4133 3282
rect 4176 3268 4219 3282
rect 4241 3278 4431 3290
rect 4496 3286 4502 3306
rect 4226 3268 4256 3278
rect 4257 3268 4415 3278
rect 4419 3268 4449 3278
rect 4453 3268 4483 3282
rect 4511 3268 4524 3306
rect 4596 3320 4625 3336
rect 4639 3320 4668 3336
rect 4683 3326 4713 3342
rect 4741 3320 4747 3368
rect 4750 3362 4769 3368
rect 4784 3362 4814 3370
rect 4750 3354 4814 3362
rect 4750 3338 4830 3354
rect 4846 3347 4908 3378
rect 4924 3347 4986 3378
rect 5055 3376 5104 3401
rect 5119 3376 5149 3392
rect 5018 3362 5048 3370
rect 5055 3368 5165 3376
rect 5018 3354 5063 3362
rect 4750 3336 4769 3338
rect 4784 3336 4830 3338
rect 4750 3320 4830 3336
rect 4857 3334 4892 3347
rect 4933 3344 4970 3347
rect 4933 3342 4975 3344
rect 4862 3331 4892 3334
rect 4871 3327 4878 3331
rect 4878 3326 4879 3327
rect 4837 3320 4847 3326
rect 4596 3312 4631 3320
rect 4596 3286 4597 3312
rect 4604 3286 4631 3312
rect 4539 3268 4569 3282
rect 4596 3278 4631 3286
rect 4633 3312 4674 3320
rect 4633 3286 4648 3312
rect 4655 3286 4674 3312
rect 4738 3308 4769 3320
rect 4784 3308 4887 3320
rect 4899 3310 4925 3336
rect 4940 3331 4970 3342
rect 5002 3338 5064 3354
rect 5002 3336 5048 3338
rect 5002 3320 5064 3336
rect 5076 3320 5082 3368
rect 5085 3360 5165 3368
rect 5085 3358 5104 3360
rect 5119 3358 5153 3360
rect 5085 3342 5165 3358
rect 5085 3320 5104 3342
rect 5119 3326 5149 3342
rect 5177 3336 5183 3410
rect 5186 3336 5205 3480
rect 5220 3336 5226 3480
rect 5235 3410 5248 3480
rect 5300 3476 5322 3480
rect 5293 3454 5322 3468
rect 5375 3454 5391 3468
rect 5429 3464 5435 3466
rect 5442 3464 5550 3480
rect 5557 3464 5563 3466
rect 5571 3464 5586 3480
rect 5652 3474 5671 3477
rect 5293 3452 5391 3454
rect 5418 3452 5586 3464
rect 5601 3454 5617 3468
rect 5652 3455 5674 3474
rect 5684 3468 5700 3469
rect 5683 3466 5700 3468
rect 5684 3461 5700 3466
rect 5674 3454 5680 3455
rect 5683 3454 5712 3461
rect 5601 3453 5712 3454
rect 5601 3452 5718 3453
rect 5277 3444 5328 3452
rect 5375 3444 5409 3452
rect 5277 3432 5302 3444
rect 5309 3432 5328 3444
rect 5382 3442 5409 3444
rect 5418 3442 5639 3452
rect 5674 3449 5680 3452
rect 5382 3438 5639 3442
rect 5277 3424 5328 3432
rect 5375 3424 5639 3438
rect 5683 3444 5718 3452
rect 5229 3376 5248 3410
rect 5293 3416 5322 3424
rect 5293 3410 5310 3416
rect 5293 3408 5327 3410
rect 5375 3408 5391 3424
rect 5392 3414 5600 3424
rect 5601 3414 5617 3424
rect 5665 3420 5680 3435
rect 5683 3432 5684 3444
rect 5691 3432 5718 3444
rect 5683 3424 5718 3432
rect 5683 3423 5712 3424
rect 5403 3410 5617 3414
rect 5418 3408 5617 3410
rect 5652 3410 5665 3420
rect 5683 3410 5700 3423
rect 5652 3408 5700 3410
rect 5294 3404 5327 3408
rect 5290 3402 5327 3404
rect 5290 3401 5357 3402
rect 5290 3396 5321 3401
rect 5327 3396 5357 3401
rect 5290 3392 5357 3396
rect 5263 3389 5357 3392
rect 5263 3382 5312 3389
rect 5263 3376 5293 3382
rect 5312 3377 5317 3382
rect 5229 3360 5309 3376
rect 5321 3368 5357 3389
rect 5418 3384 5607 3408
rect 5652 3407 5699 3408
rect 5665 3402 5699 3407
rect 5433 3381 5607 3384
rect 5426 3378 5607 3381
rect 5635 3401 5699 3402
rect 5229 3358 5248 3360
rect 5263 3358 5297 3360
rect 5229 3342 5309 3358
rect 5229 3336 5248 3342
rect 4945 3310 5048 3320
rect 4899 3308 5048 3310
rect 5069 3308 5104 3320
rect 4738 3306 4900 3308
rect 4750 3286 4769 3306
rect 4784 3304 4814 3306
rect 4633 3278 4674 3286
rect 4756 3282 4769 3286
rect 4821 3290 4900 3306
rect 4932 3306 5104 3308
rect 4932 3290 5011 3306
rect 5018 3304 5048 3306
rect 4596 3268 4625 3278
rect 4639 3268 4668 3278
rect 4683 3268 4713 3282
rect 4756 3268 4799 3282
rect 4821 3278 5011 3290
rect 5076 3286 5082 3306
rect 4806 3268 4836 3278
rect 4837 3268 4995 3278
rect 4999 3268 5029 3278
rect 5033 3268 5063 3282
rect 5091 3268 5104 3306
rect 5176 3320 5205 3336
rect 5219 3320 5248 3336
rect 5263 3326 5293 3342
rect 5321 3320 5327 3368
rect 5330 3362 5349 3368
rect 5364 3362 5394 3370
rect 5330 3354 5394 3362
rect 5330 3338 5410 3354
rect 5426 3347 5488 3378
rect 5504 3347 5566 3378
rect 5635 3376 5684 3401
rect 5699 3376 5729 3392
rect 5598 3362 5628 3370
rect 5635 3368 5745 3376
rect 5598 3354 5643 3362
rect 5330 3336 5349 3338
rect 5364 3336 5410 3338
rect 5330 3320 5410 3336
rect 5437 3334 5472 3347
rect 5513 3344 5550 3347
rect 5513 3342 5555 3344
rect 5442 3331 5472 3334
rect 5451 3327 5458 3331
rect 5458 3326 5459 3327
rect 5417 3320 5427 3326
rect 5176 3312 5211 3320
rect 5176 3286 5177 3312
rect 5184 3286 5211 3312
rect 5119 3268 5149 3282
rect 5176 3278 5211 3286
rect 5213 3312 5254 3320
rect 5213 3286 5228 3312
rect 5235 3286 5254 3312
rect 5318 3308 5349 3320
rect 5364 3308 5467 3320
rect 5479 3310 5505 3336
rect 5520 3331 5550 3342
rect 5582 3338 5644 3354
rect 5582 3336 5628 3338
rect 5582 3320 5644 3336
rect 5656 3320 5662 3368
rect 5665 3360 5745 3368
rect 5665 3358 5684 3360
rect 5699 3358 5733 3360
rect 5665 3342 5745 3358
rect 5665 3320 5684 3342
rect 5699 3326 5729 3342
rect 5757 3336 5763 3410
rect 5766 3336 5785 3480
rect 5800 3336 5806 3480
rect 5815 3410 5828 3480
rect 5880 3476 5902 3480
rect 5873 3454 5902 3468
rect 5955 3454 5971 3468
rect 6009 3464 6015 3466
rect 6022 3464 6130 3480
rect 6137 3464 6143 3466
rect 6151 3464 6166 3480
rect 6232 3474 6251 3477
rect 5873 3452 5971 3454
rect 5998 3452 6166 3464
rect 6181 3454 6197 3468
rect 6232 3455 6254 3474
rect 6264 3468 6280 3469
rect 6263 3466 6280 3468
rect 6264 3461 6280 3466
rect 6254 3454 6260 3455
rect 6263 3454 6292 3461
rect 6181 3453 6292 3454
rect 6181 3452 6298 3453
rect 5857 3444 5908 3452
rect 5955 3444 5989 3452
rect 5857 3432 5882 3444
rect 5889 3432 5908 3444
rect 5962 3442 5989 3444
rect 5998 3442 6219 3452
rect 6254 3449 6260 3452
rect 5962 3438 6219 3442
rect 5857 3424 5908 3432
rect 5955 3424 6219 3438
rect 6263 3444 6298 3452
rect 5809 3376 5828 3410
rect 5873 3416 5902 3424
rect 5873 3410 5890 3416
rect 5873 3408 5907 3410
rect 5955 3408 5971 3424
rect 5972 3414 6180 3424
rect 6181 3414 6197 3424
rect 6245 3420 6260 3435
rect 6263 3432 6264 3444
rect 6271 3432 6298 3444
rect 6263 3424 6298 3432
rect 6263 3423 6292 3424
rect 5983 3410 6197 3414
rect 5998 3408 6197 3410
rect 6232 3410 6245 3420
rect 6263 3410 6280 3423
rect 6232 3408 6280 3410
rect 5874 3404 5907 3408
rect 5870 3402 5907 3404
rect 5870 3401 5937 3402
rect 5870 3396 5901 3401
rect 5907 3396 5937 3401
rect 5870 3392 5937 3396
rect 5843 3389 5937 3392
rect 5843 3382 5892 3389
rect 5843 3376 5873 3382
rect 5892 3377 5897 3382
rect 5809 3360 5889 3376
rect 5901 3368 5937 3389
rect 5998 3384 6187 3408
rect 6232 3407 6279 3408
rect 6245 3402 6279 3407
rect 6013 3381 6187 3384
rect 6006 3378 6187 3381
rect 6215 3401 6279 3402
rect 5809 3358 5828 3360
rect 5843 3358 5877 3360
rect 5809 3342 5889 3358
rect 5809 3336 5828 3342
rect 5525 3310 5628 3320
rect 5479 3308 5628 3310
rect 5649 3308 5684 3320
rect 5318 3306 5480 3308
rect 5330 3286 5349 3306
rect 5364 3304 5394 3306
rect 5213 3278 5254 3286
rect 5336 3282 5349 3286
rect 5401 3290 5480 3306
rect 5512 3306 5684 3308
rect 5512 3290 5591 3306
rect 5598 3304 5628 3306
rect 5176 3268 5205 3278
rect 5219 3268 5248 3278
rect 5263 3268 5293 3282
rect 5336 3268 5379 3282
rect 5401 3278 5591 3290
rect 5656 3286 5662 3306
rect 5386 3268 5416 3278
rect 5417 3268 5575 3278
rect 5579 3268 5609 3278
rect 5613 3268 5643 3282
rect 5671 3268 5684 3306
rect 5756 3320 5785 3336
rect 5799 3320 5828 3336
rect 5843 3326 5873 3342
rect 5901 3320 5907 3368
rect 5910 3362 5929 3368
rect 5944 3362 5974 3370
rect 5910 3354 5974 3362
rect 5910 3338 5990 3354
rect 6006 3347 6068 3378
rect 6084 3347 6146 3378
rect 6215 3376 6264 3401
rect 6279 3376 6309 3392
rect 6178 3362 6208 3370
rect 6215 3368 6325 3376
rect 6178 3354 6223 3362
rect 5910 3336 5929 3338
rect 5944 3336 5990 3338
rect 5910 3320 5990 3336
rect 6017 3334 6052 3347
rect 6093 3344 6130 3347
rect 6093 3342 6135 3344
rect 6022 3331 6052 3334
rect 6031 3327 6038 3331
rect 6038 3326 6039 3327
rect 5997 3320 6007 3326
rect 5756 3312 5791 3320
rect 5756 3286 5757 3312
rect 5764 3286 5791 3312
rect 5699 3268 5729 3282
rect 5756 3278 5791 3286
rect 5793 3312 5834 3320
rect 5793 3286 5808 3312
rect 5815 3286 5834 3312
rect 5898 3308 5929 3320
rect 5944 3308 6047 3320
rect 6059 3310 6085 3336
rect 6100 3331 6130 3342
rect 6162 3338 6224 3354
rect 6162 3336 6208 3338
rect 6162 3320 6224 3336
rect 6236 3320 6242 3368
rect 6245 3360 6325 3368
rect 6245 3358 6264 3360
rect 6279 3358 6313 3360
rect 6245 3342 6325 3358
rect 6245 3320 6264 3342
rect 6279 3326 6309 3342
rect 6337 3336 6343 3410
rect 6346 3336 6365 3480
rect 6380 3336 6386 3480
rect 6395 3410 6408 3480
rect 6460 3476 6482 3480
rect 6453 3454 6482 3468
rect 6535 3454 6551 3468
rect 6589 3464 6595 3466
rect 6602 3464 6710 3480
rect 6717 3464 6723 3466
rect 6731 3464 6746 3480
rect 6812 3474 6831 3477
rect 6453 3452 6551 3454
rect 6578 3452 6746 3464
rect 6761 3454 6777 3468
rect 6812 3455 6834 3474
rect 6844 3468 6860 3469
rect 6843 3466 6860 3468
rect 6844 3461 6860 3466
rect 6834 3454 6840 3455
rect 6843 3454 6872 3461
rect 6761 3453 6872 3454
rect 6761 3452 6878 3453
rect 6437 3444 6488 3452
rect 6535 3444 6569 3452
rect 6437 3432 6462 3444
rect 6469 3432 6488 3444
rect 6542 3442 6569 3444
rect 6578 3442 6799 3452
rect 6834 3449 6840 3452
rect 6542 3438 6799 3442
rect 6437 3424 6488 3432
rect 6535 3424 6799 3438
rect 6843 3444 6878 3452
rect 6389 3376 6408 3410
rect 6453 3416 6482 3424
rect 6453 3410 6470 3416
rect 6453 3408 6487 3410
rect 6535 3408 6551 3424
rect 6552 3414 6760 3424
rect 6761 3414 6777 3424
rect 6825 3420 6840 3435
rect 6843 3432 6844 3444
rect 6851 3432 6878 3444
rect 6843 3424 6878 3432
rect 6843 3423 6872 3424
rect 6563 3410 6777 3414
rect 6578 3408 6777 3410
rect 6812 3410 6825 3420
rect 6843 3410 6860 3423
rect 6812 3408 6860 3410
rect 6454 3404 6487 3408
rect 6450 3402 6487 3404
rect 6450 3401 6517 3402
rect 6450 3396 6481 3401
rect 6487 3396 6517 3401
rect 6450 3392 6517 3396
rect 6423 3389 6517 3392
rect 6423 3382 6472 3389
rect 6423 3376 6453 3382
rect 6472 3377 6477 3382
rect 6389 3360 6469 3376
rect 6481 3368 6517 3389
rect 6578 3384 6767 3408
rect 6812 3407 6859 3408
rect 6825 3402 6859 3407
rect 6593 3381 6767 3384
rect 6586 3378 6767 3381
rect 6795 3401 6859 3402
rect 6389 3358 6408 3360
rect 6423 3358 6457 3360
rect 6389 3342 6469 3358
rect 6389 3336 6408 3342
rect 6105 3310 6208 3320
rect 6059 3308 6208 3310
rect 6229 3308 6264 3320
rect 5898 3306 6060 3308
rect 5910 3286 5929 3306
rect 5944 3304 5974 3306
rect 5793 3278 5834 3286
rect 5916 3282 5929 3286
rect 5981 3290 6060 3306
rect 6092 3306 6264 3308
rect 6092 3290 6171 3306
rect 6178 3304 6208 3306
rect 5756 3268 5785 3278
rect 5799 3268 5828 3278
rect 5843 3268 5873 3282
rect 5916 3268 5959 3282
rect 5981 3278 6171 3290
rect 6236 3286 6242 3306
rect 5966 3268 5996 3278
rect 5997 3268 6155 3278
rect 6159 3268 6189 3278
rect 6193 3268 6223 3282
rect 6251 3268 6264 3306
rect 6336 3320 6365 3336
rect 6379 3320 6408 3336
rect 6423 3326 6453 3342
rect 6481 3320 6487 3368
rect 6490 3362 6509 3368
rect 6524 3362 6554 3370
rect 6490 3354 6554 3362
rect 6490 3338 6570 3354
rect 6586 3347 6648 3378
rect 6664 3347 6726 3378
rect 6795 3376 6844 3401
rect 6859 3376 6889 3392
rect 6758 3362 6788 3370
rect 6795 3368 6905 3376
rect 6758 3354 6803 3362
rect 6490 3336 6509 3338
rect 6524 3336 6570 3338
rect 6490 3320 6570 3336
rect 6597 3334 6632 3347
rect 6673 3344 6710 3347
rect 6673 3342 6715 3344
rect 6602 3331 6632 3334
rect 6611 3327 6618 3331
rect 6618 3326 6619 3327
rect 6577 3320 6587 3326
rect 6336 3312 6371 3320
rect 6336 3286 6337 3312
rect 6344 3286 6371 3312
rect 6279 3268 6309 3282
rect 6336 3278 6371 3286
rect 6373 3312 6414 3320
rect 6373 3286 6388 3312
rect 6395 3286 6414 3312
rect 6478 3308 6509 3320
rect 6524 3308 6627 3320
rect 6639 3310 6665 3336
rect 6680 3331 6710 3342
rect 6742 3338 6804 3354
rect 6742 3336 6788 3338
rect 6742 3320 6804 3336
rect 6816 3320 6822 3368
rect 6825 3360 6905 3368
rect 6825 3358 6844 3360
rect 6859 3358 6893 3360
rect 6825 3342 6905 3358
rect 6825 3320 6844 3342
rect 6859 3326 6889 3342
rect 6917 3336 6923 3410
rect 6926 3336 6945 3480
rect 6960 3336 6966 3480
rect 6975 3410 6988 3480
rect 7040 3476 7062 3480
rect 7033 3454 7062 3468
rect 7115 3454 7131 3468
rect 7169 3464 7175 3466
rect 7182 3464 7290 3480
rect 7297 3464 7303 3466
rect 7311 3464 7326 3480
rect 7392 3474 7411 3477
rect 7033 3452 7131 3454
rect 7158 3452 7326 3464
rect 7341 3454 7357 3468
rect 7392 3455 7414 3474
rect 7424 3468 7440 3469
rect 7423 3466 7440 3468
rect 7424 3461 7440 3466
rect 7414 3454 7420 3455
rect 7423 3454 7452 3461
rect 7341 3453 7452 3454
rect 7341 3452 7458 3453
rect 7017 3444 7068 3452
rect 7115 3444 7149 3452
rect 7017 3432 7042 3444
rect 7049 3432 7068 3444
rect 7122 3442 7149 3444
rect 7158 3442 7379 3452
rect 7414 3449 7420 3452
rect 7122 3438 7379 3442
rect 7017 3424 7068 3432
rect 7115 3424 7379 3438
rect 7423 3444 7458 3452
rect 6969 3376 6988 3410
rect 7033 3416 7062 3424
rect 7033 3410 7050 3416
rect 7033 3408 7067 3410
rect 7115 3408 7131 3424
rect 7132 3414 7340 3424
rect 7341 3414 7357 3424
rect 7405 3420 7420 3435
rect 7423 3432 7424 3444
rect 7431 3432 7458 3444
rect 7423 3424 7458 3432
rect 7423 3423 7452 3424
rect 7143 3410 7357 3414
rect 7158 3408 7357 3410
rect 7392 3410 7405 3420
rect 7423 3410 7440 3423
rect 7392 3408 7440 3410
rect 7034 3404 7067 3408
rect 7030 3402 7067 3404
rect 7030 3401 7097 3402
rect 7030 3396 7061 3401
rect 7067 3396 7097 3401
rect 7030 3392 7097 3396
rect 7003 3389 7097 3392
rect 7003 3382 7052 3389
rect 7003 3376 7033 3382
rect 7052 3377 7057 3382
rect 6969 3360 7049 3376
rect 7061 3368 7097 3389
rect 7158 3384 7347 3408
rect 7392 3407 7439 3408
rect 7405 3402 7439 3407
rect 7173 3381 7347 3384
rect 7166 3378 7347 3381
rect 7375 3401 7439 3402
rect 6969 3358 6988 3360
rect 7003 3358 7037 3360
rect 6969 3342 7049 3358
rect 6969 3336 6988 3342
rect 6685 3310 6788 3320
rect 6639 3308 6788 3310
rect 6809 3308 6844 3320
rect 6478 3306 6640 3308
rect 6490 3286 6509 3306
rect 6524 3304 6554 3306
rect 6373 3278 6414 3286
rect 6496 3282 6509 3286
rect 6561 3290 6640 3306
rect 6672 3306 6844 3308
rect 6672 3290 6751 3306
rect 6758 3304 6788 3306
rect 6336 3268 6365 3278
rect 6379 3268 6408 3278
rect 6423 3268 6453 3282
rect 6496 3268 6539 3282
rect 6561 3278 6751 3290
rect 6816 3286 6822 3306
rect 6546 3268 6576 3278
rect 6577 3268 6735 3278
rect 6739 3268 6769 3278
rect 6773 3268 6803 3282
rect 6831 3268 6844 3306
rect 6916 3320 6945 3336
rect 6959 3320 6988 3336
rect 7003 3326 7033 3342
rect 7061 3320 7067 3368
rect 7070 3362 7089 3368
rect 7104 3362 7134 3370
rect 7070 3354 7134 3362
rect 7070 3338 7150 3354
rect 7166 3347 7228 3378
rect 7244 3347 7306 3378
rect 7375 3376 7424 3401
rect 7439 3376 7469 3392
rect 7338 3362 7368 3370
rect 7375 3368 7485 3376
rect 7338 3354 7383 3362
rect 7070 3336 7089 3338
rect 7104 3336 7150 3338
rect 7070 3320 7150 3336
rect 7177 3334 7212 3347
rect 7253 3344 7290 3347
rect 7253 3342 7295 3344
rect 7182 3331 7212 3334
rect 7191 3327 7198 3331
rect 7198 3326 7199 3327
rect 7157 3320 7167 3326
rect 6916 3312 6951 3320
rect 6916 3286 6917 3312
rect 6924 3286 6951 3312
rect 6859 3268 6889 3282
rect 6916 3278 6951 3286
rect 6953 3312 6994 3320
rect 6953 3286 6968 3312
rect 6975 3286 6994 3312
rect 7058 3308 7089 3320
rect 7104 3308 7207 3320
rect 7219 3310 7245 3336
rect 7260 3331 7290 3342
rect 7322 3338 7384 3354
rect 7322 3336 7368 3338
rect 7322 3320 7384 3336
rect 7396 3320 7402 3368
rect 7405 3360 7485 3368
rect 7405 3358 7424 3360
rect 7439 3358 7473 3360
rect 7405 3342 7485 3358
rect 7405 3320 7424 3342
rect 7439 3326 7469 3342
rect 7497 3336 7503 3410
rect 7506 3336 7525 3480
rect 7540 3336 7546 3480
rect 7555 3410 7568 3480
rect 7613 3458 7614 3468
rect 7629 3458 7642 3468
rect 7613 3454 7642 3458
rect 7647 3454 7677 3480
rect 7695 3466 7711 3468
rect 7783 3466 7836 3480
rect 7784 3464 7848 3466
rect 7891 3464 7906 3480
rect 7955 3477 7985 3480
rect 7955 3474 7991 3477
rect 7921 3466 7937 3468
rect 7695 3454 7710 3458
rect 7613 3452 7710 3454
rect 7738 3452 7906 3464
rect 7922 3454 7937 3458
rect 7955 3455 7994 3474
rect 8013 3468 8020 3469
rect 8019 3461 8020 3468
rect 8003 3458 8004 3461
rect 8019 3458 8032 3461
rect 7955 3454 7985 3455
rect 7994 3454 8000 3455
rect 8003 3454 8032 3458
rect 7922 3453 8032 3454
rect 7922 3452 8038 3453
rect 7597 3444 7648 3452
rect 7597 3432 7622 3444
rect 7629 3432 7648 3444
rect 7679 3444 7729 3452
rect 7679 3436 7695 3444
rect 7702 3442 7729 3444
rect 7738 3442 7959 3452
rect 7702 3432 7959 3442
rect 7988 3444 8038 3452
rect 7988 3435 8004 3444
rect 7597 3424 7648 3432
rect 7695 3424 7959 3432
rect 7985 3432 8004 3435
rect 8011 3432 8038 3444
rect 7985 3424 8038 3432
rect 7549 3376 7568 3410
rect 7613 3416 7614 3424
rect 7629 3416 7642 3424
rect 7613 3408 7629 3416
rect 7610 3401 7629 3404
rect 7610 3392 7632 3401
rect 7583 3382 7632 3392
rect 7583 3376 7613 3382
rect 7632 3377 7637 3382
rect 7549 3360 7629 3376
rect 7647 3368 7677 3424
rect 7712 3414 7920 3424
rect 7955 3420 8000 3424
rect 8003 3423 8004 3424
rect 8019 3423 8032 3424
rect 7738 3384 7927 3414
rect 7753 3381 7927 3384
rect 7746 3378 7927 3381
rect 7549 3358 7568 3360
rect 7583 3358 7617 3360
rect 7549 3342 7629 3358
rect 7656 3354 7669 3368
rect 7684 3354 7700 3370
rect 7746 3365 7757 3378
rect 7549 3336 7568 3342
rect 7265 3310 7368 3320
rect 7219 3308 7368 3310
rect 7389 3308 7424 3320
rect 7058 3306 7220 3308
rect 7070 3286 7089 3306
rect 7104 3304 7134 3306
rect 6953 3278 6994 3286
rect 7076 3282 7089 3286
rect 7141 3290 7220 3306
rect 7252 3306 7424 3308
rect 7252 3290 7331 3306
rect 7338 3304 7368 3306
rect 6916 3268 6945 3278
rect 6959 3268 6988 3278
rect 7003 3268 7033 3282
rect 7076 3268 7119 3282
rect 7141 3278 7331 3290
rect 7396 3286 7402 3306
rect 7126 3268 7156 3278
rect 7157 3268 7315 3278
rect 7319 3268 7349 3278
rect 7353 3268 7383 3282
rect 7411 3268 7424 3306
rect 7496 3320 7525 3336
rect 7539 3320 7568 3336
rect 7583 3320 7613 3342
rect 7656 3338 7718 3354
rect 7746 3347 7757 3363
rect 7762 3358 7772 3378
rect 7782 3358 7796 3378
rect 7799 3365 7808 3378
rect 7824 3365 7833 3378
rect 7762 3347 7796 3358
rect 7799 3347 7808 3363
rect 7824 3347 7833 3363
rect 7840 3358 7850 3378
rect 7860 3358 7874 3378
rect 7875 3365 7886 3378
rect 7840 3347 7874 3358
rect 7875 3347 7886 3363
rect 7932 3354 7948 3370
rect 7955 3368 7985 3420
rect 8019 3416 8020 3423
rect 8004 3408 8020 3416
rect 7991 3376 8004 3395
rect 8019 3376 8049 3392
rect 7991 3360 8065 3376
rect 7991 3358 8004 3360
rect 8019 3358 8053 3360
rect 7656 3336 7669 3338
rect 7684 3336 7718 3338
rect 7656 3320 7718 3336
rect 7762 3331 7778 3334
rect 7840 3331 7870 3342
rect 7918 3338 7964 3354
rect 7991 3342 8065 3358
rect 7918 3336 7952 3338
rect 7917 3320 7964 3336
rect 7991 3320 8004 3342
rect 8019 3320 8049 3342
rect 8076 3320 8077 3336
rect 8092 3320 8105 3480
rect 8135 3376 8148 3480
rect 8193 3458 8194 3468
rect 8209 3458 8222 3468
rect 8193 3454 8222 3458
rect 8227 3454 8257 3480
rect 8275 3466 8291 3468
rect 8363 3466 8416 3480
rect 8364 3464 8428 3466
rect 8471 3464 8486 3480
rect 8535 3477 8565 3480
rect 8535 3474 8571 3477
rect 8501 3466 8517 3468
rect 8275 3454 8290 3458
rect 8193 3452 8290 3454
rect 8318 3452 8486 3464
rect 8502 3454 8517 3458
rect 8535 3455 8574 3474
rect 8593 3468 8600 3469
rect 8599 3461 8600 3468
rect 8583 3458 8584 3461
rect 8599 3458 8612 3461
rect 8535 3454 8565 3455
rect 8574 3454 8580 3455
rect 8583 3454 8612 3458
rect 8502 3453 8612 3454
rect 8502 3452 8618 3453
rect 8177 3444 8228 3452
rect 8177 3432 8202 3444
rect 8209 3432 8228 3444
rect 8259 3444 8309 3452
rect 8259 3436 8275 3444
rect 8282 3442 8309 3444
rect 8318 3442 8539 3452
rect 8282 3432 8539 3442
rect 8568 3444 8618 3452
rect 8568 3435 8584 3444
rect 8177 3424 8228 3432
rect 8275 3424 8539 3432
rect 8565 3432 8584 3435
rect 8591 3432 8618 3444
rect 8565 3424 8618 3432
rect 8193 3416 8194 3424
rect 8209 3416 8222 3424
rect 8193 3408 8209 3416
rect 8190 3401 8209 3404
rect 8190 3392 8212 3401
rect 8163 3382 8212 3392
rect 8163 3376 8193 3382
rect 8212 3377 8217 3382
rect 8135 3360 8209 3376
rect 8227 3368 8257 3424
rect 8292 3414 8500 3424
rect 8535 3420 8580 3424
rect 8583 3423 8584 3424
rect 8599 3423 8612 3424
rect 8318 3384 8507 3414
rect 8333 3381 8507 3384
rect 8326 3378 8507 3381
rect 8135 3358 8148 3360
rect 8163 3358 8197 3360
rect 8135 3342 8209 3358
rect 8236 3354 8249 3368
rect 8264 3354 8280 3370
rect 8326 3365 8337 3378
rect 8119 3320 8120 3336
rect 8135 3320 8148 3342
rect 8163 3320 8193 3342
rect 8236 3338 8298 3354
rect 8326 3347 8337 3363
rect 8342 3358 8352 3378
rect 8362 3358 8376 3378
rect 8379 3365 8388 3378
rect 8404 3365 8413 3378
rect 8342 3347 8376 3358
rect 8379 3347 8388 3363
rect 8404 3347 8413 3363
rect 8420 3358 8430 3378
rect 8440 3358 8454 3378
rect 8455 3365 8466 3378
rect 8420 3347 8454 3358
rect 8455 3347 8466 3363
rect 8512 3354 8528 3370
rect 8535 3368 8565 3420
rect 8599 3416 8600 3423
rect 8584 3408 8600 3416
rect 8571 3376 8584 3395
rect 8599 3376 8629 3392
rect 8571 3360 8645 3376
rect 8571 3358 8584 3360
rect 8599 3358 8633 3360
rect 8236 3336 8249 3338
rect 8264 3336 8298 3338
rect 8236 3320 8298 3336
rect 8342 3331 8358 3334
rect 8420 3331 8450 3342
rect 8498 3338 8544 3354
rect 8571 3342 8645 3358
rect 8498 3336 8532 3338
rect 8497 3320 8544 3336
rect 8571 3320 8584 3342
rect 8599 3320 8629 3342
rect 8656 3320 8657 3336
rect 8672 3320 8685 3480
rect 8715 3376 8728 3480
rect 8773 3458 8774 3468
rect 8789 3458 8802 3468
rect 8773 3454 8802 3458
rect 8807 3454 8837 3480
rect 8855 3466 8871 3468
rect 8943 3466 8996 3480
rect 8944 3464 9008 3466
rect 9051 3464 9066 3480
rect 9115 3477 9145 3480
rect 9115 3474 9151 3477
rect 9081 3466 9097 3468
rect 8855 3454 8870 3458
rect 8773 3452 8870 3454
rect 8898 3452 9066 3464
rect 9082 3454 9097 3458
rect 9115 3455 9154 3474
rect 9173 3468 9180 3469
rect 9179 3461 9180 3468
rect 9163 3458 9164 3461
rect 9179 3458 9192 3461
rect 9115 3454 9145 3455
rect 9154 3454 9160 3455
rect 9163 3454 9192 3458
rect 9082 3453 9192 3454
rect 9082 3452 9198 3453
rect 8757 3444 8808 3452
rect 8757 3432 8782 3444
rect 8789 3432 8808 3444
rect 8839 3444 8889 3452
rect 8839 3436 8855 3444
rect 8862 3442 8889 3444
rect 8898 3442 9119 3452
rect 8862 3432 9119 3442
rect 9148 3444 9198 3452
rect 9148 3435 9164 3444
rect 8757 3424 8808 3432
rect 8855 3424 9119 3432
rect 9145 3432 9164 3435
rect 9171 3432 9198 3444
rect 9145 3424 9198 3432
rect 8773 3416 8774 3424
rect 8789 3416 8802 3424
rect 8773 3408 8789 3416
rect 8770 3401 8789 3404
rect 8770 3392 8792 3401
rect 8743 3382 8792 3392
rect 8743 3376 8773 3382
rect 8792 3377 8797 3382
rect 8715 3360 8789 3376
rect 8807 3368 8837 3424
rect 8872 3414 9080 3424
rect 9115 3420 9160 3424
rect 9163 3423 9164 3424
rect 9179 3423 9192 3424
rect 8898 3384 9087 3414
rect 8913 3381 9087 3384
rect 8906 3378 9087 3381
rect 8715 3358 8728 3360
rect 8743 3358 8777 3360
rect 8715 3342 8789 3358
rect 8816 3354 8829 3368
rect 8844 3354 8860 3370
rect 8906 3365 8917 3378
rect 8699 3320 8700 3336
rect 8715 3320 8728 3342
rect 8743 3320 8773 3342
rect 8816 3338 8878 3354
rect 8906 3347 8917 3363
rect 8922 3358 8932 3378
rect 8942 3358 8956 3378
rect 8959 3365 8968 3378
rect 8984 3365 8993 3378
rect 8922 3347 8956 3358
rect 8959 3347 8968 3363
rect 8984 3347 8993 3363
rect 9000 3358 9010 3378
rect 9020 3358 9034 3378
rect 9035 3365 9046 3378
rect 9000 3347 9034 3358
rect 9035 3347 9046 3363
rect 9092 3354 9108 3370
rect 9115 3368 9145 3420
rect 9179 3416 9180 3423
rect 9164 3408 9180 3416
rect 9151 3376 9164 3395
rect 9179 3376 9209 3392
rect 9151 3360 9225 3376
rect 9151 3358 9164 3360
rect 9179 3358 9213 3360
rect 8816 3336 8829 3338
rect 8844 3336 8878 3338
rect 8816 3320 8878 3336
rect 8922 3331 8938 3334
rect 9000 3331 9030 3342
rect 9078 3338 9124 3354
rect 9151 3342 9225 3358
rect 9078 3336 9112 3338
rect 9077 3320 9124 3336
rect 9151 3320 9164 3342
rect 9179 3320 9209 3342
rect 9236 3320 9237 3336
rect 9252 3320 9265 3480
rect 7496 3312 7531 3320
rect 7496 3286 7497 3312
rect 7504 3286 7531 3312
rect 7439 3268 7469 3282
rect 7496 3278 7531 3286
rect 7533 3312 7574 3320
rect 7533 3286 7548 3312
rect 7555 3286 7574 3312
rect 7638 3308 7700 3320
rect 7712 3308 7787 3320
rect 7845 3308 7920 3320
rect 7932 3308 7963 3320
rect 7969 3308 8004 3320
rect 7638 3306 7800 3308
rect 7533 3278 7574 3286
rect 7656 3282 7669 3306
rect 7684 3304 7699 3306
rect 7496 3268 7525 3278
rect 7539 3268 7568 3278
rect 7583 3268 7613 3282
rect 7656 3268 7699 3282
rect 7723 3279 7730 3286
rect 7733 3282 7800 3306
rect 7832 3306 8004 3308
rect 7802 3284 7830 3288
rect 7832 3284 7912 3306
rect 7933 3304 7948 3306
rect 7802 3282 7912 3284
rect 7733 3278 7912 3282
rect 7706 3268 7736 3278
rect 7738 3268 7891 3278
rect 7899 3268 7929 3278
rect 7933 3268 7963 3282
rect 7991 3268 8004 3306
rect 8076 3312 8111 3320
rect 8076 3286 8077 3312
rect 8084 3286 8111 3312
rect 8019 3268 8049 3282
rect 8076 3278 8111 3286
rect 8113 3312 8154 3320
rect 8113 3286 8128 3312
rect 8135 3286 8154 3312
rect 8218 3308 8280 3320
rect 8292 3308 8367 3320
rect 8425 3308 8500 3320
rect 8512 3308 8543 3320
rect 8549 3308 8584 3320
rect 8218 3306 8380 3308
rect 8113 3278 8154 3286
rect 8236 3282 8249 3306
rect 8264 3304 8279 3306
rect 8076 3268 8077 3278
rect 8092 3268 8105 3278
rect 8119 3268 8120 3278
rect 8135 3268 8148 3278
rect 8163 3268 8193 3282
rect 8236 3268 8279 3282
rect 8303 3279 8310 3286
rect 8313 3282 8380 3306
rect 8412 3306 8584 3308
rect 8382 3284 8410 3288
rect 8412 3284 8492 3306
rect 8513 3304 8528 3306
rect 8382 3282 8492 3284
rect 8313 3278 8492 3282
rect 8286 3268 8316 3278
rect 8318 3268 8471 3278
rect 8479 3268 8509 3278
rect 8513 3268 8543 3282
rect 8571 3268 8584 3306
rect 8656 3312 8691 3320
rect 8656 3286 8657 3312
rect 8664 3286 8691 3312
rect 8599 3268 8629 3282
rect 8656 3278 8691 3286
rect 8693 3312 8734 3320
rect 8693 3286 8708 3312
rect 8715 3286 8734 3312
rect 8798 3308 8860 3320
rect 8872 3308 8947 3320
rect 9005 3308 9080 3320
rect 9092 3308 9123 3320
rect 9129 3308 9164 3320
rect 8798 3306 8960 3308
rect 8693 3278 8734 3286
rect 8816 3282 8829 3306
rect 8844 3304 8859 3306
rect 8656 3268 8657 3278
rect 8672 3268 8685 3278
rect 8699 3268 8700 3278
rect 8715 3268 8728 3278
rect 8743 3268 8773 3282
rect 8816 3268 8859 3282
rect 8883 3279 8890 3286
rect 8893 3282 8960 3306
rect 8992 3306 9164 3308
rect 8962 3284 8990 3288
rect 8992 3284 9072 3306
rect 9093 3304 9108 3306
rect 8962 3282 9072 3284
rect 8893 3278 9072 3282
rect 8866 3268 8896 3278
rect 8898 3268 9051 3278
rect 9059 3268 9089 3278
rect 9093 3268 9123 3282
rect 9151 3268 9164 3306
rect 9236 3312 9271 3320
rect 9236 3286 9237 3312
rect 9244 3286 9271 3312
rect 9179 3268 9209 3282
rect 9236 3278 9271 3286
rect 9236 3268 9237 3278
rect 9252 3268 9265 3278
rect -1 3262 9265 3268
rect 0 3254 9265 3262
rect 15 3224 28 3254
rect 43 3240 73 3254
rect 116 3240 159 3254
rect 166 3240 386 3254
rect 393 3240 423 3254
rect 83 3226 98 3238
rect 117 3226 130 3240
rect 198 3236 351 3240
rect 80 3224 102 3226
rect 180 3224 372 3236
rect 451 3224 464 3254
rect 479 3240 509 3254
rect 546 3224 565 3254
rect 580 3224 586 3254
rect 595 3224 608 3254
rect 623 3240 653 3254
rect 696 3240 739 3254
rect 746 3240 966 3254
rect 973 3240 1003 3254
rect 663 3226 678 3238
rect 697 3226 710 3240
rect 778 3236 931 3240
rect 660 3224 682 3226
rect 760 3224 952 3236
rect 1031 3224 1044 3254
rect 1059 3240 1089 3254
rect 1126 3224 1145 3254
rect 1160 3224 1166 3254
rect 1175 3224 1188 3254
rect 1203 3240 1233 3254
rect 1276 3240 1319 3254
rect 1326 3240 1546 3254
rect 1553 3240 1583 3254
rect 1243 3226 1258 3238
rect 1277 3226 1290 3240
rect 1358 3236 1511 3240
rect 1240 3224 1262 3226
rect 1340 3224 1532 3236
rect 1611 3224 1624 3254
rect 1639 3240 1669 3254
rect 1706 3224 1725 3254
rect 1740 3224 1746 3254
rect 1755 3224 1768 3254
rect 1783 3240 1813 3254
rect 1856 3240 1899 3254
rect 1906 3240 2126 3254
rect 2133 3240 2163 3254
rect 1823 3226 1838 3238
rect 1857 3226 1870 3240
rect 1938 3236 2091 3240
rect 1820 3224 1842 3226
rect 1920 3224 2112 3236
rect 2191 3224 2204 3254
rect 2219 3240 2249 3254
rect 2286 3224 2305 3254
rect 2320 3224 2326 3254
rect 2335 3224 2348 3254
rect 2363 3240 2393 3254
rect 2436 3240 2479 3254
rect 2486 3240 2706 3254
rect 2713 3240 2743 3254
rect 2403 3226 2418 3238
rect 2437 3226 2450 3240
rect 2518 3236 2671 3240
rect 2400 3224 2422 3226
rect 2500 3224 2692 3236
rect 2771 3224 2784 3254
rect 2799 3240 2829 3254
rect 2866 3224 2885 3254
rect 2900 3224 2906 3254
rect 2915 3224 2928 3254
rect 2943 3240 2973 3254
rect 3016 3240 3059 3254
rect 3066 3240 3286 3254
rect 3293 3240 3323 3254
rect 2983 3226 2998 3238
rect 3017 3226 3030 3240
rect 3098 3236 3251 3240
rect 2980 3224 3002 3226
rect 3080 3224 3272 3236
rect 3351 3224 3364 3254
rect 3379 3240 3409 3254
rect 3446 3224 3465 3254
rect 3480 3224 3486 3254
rect 3495 3224 3508 3254
rect 3523 3240 3553 3254
rect 3596 3240 3639 3254
rect 3646 3240 3866 3254
rect 3873 3240 3903 3254
rect 3563 3226 3578 3238
rect 3597 3226 3610 3240
rect 3678 3236 3831 3240
rect 3560 3224 3582 3226
rect 3660 3224 3852 3236
rect 3931 3224 3944 3254
rect 3959 3240 3989 3254
rect 4026 3224 4045 3254
rect 4060 3224 4066 3254
rect 4075 3224 4088 3254
rect 4103 3240 4133 3254
rect 4176 3240 4219 3254
rect 4226 3240 4446 3254
rect 4453 3240 4483 3254
rect 4143 3226 4158 3238
rect 4177 3226 4190 3240
rect 4258 3236 4411 3240
rect 4140 3224 4162 3226
rect 4240 3224 4432 3236
rect 4511 3224 4524 3254
rect 4539 3240 4569 3254
rect 4606 3224 4625 3254
rect 4640 3224 4646 3254
rect 4655 3224 4668 3254
rect 4683 3240 4713 3254
rect 4756 3240 4799 3254
rect 4806 3240 5026 3254
rect 5033 3240 5063 3254
rect 4723 3226 4738 3238
rect 4757 3226 4770 3240
rect 4838 3236 4991 3240
rect 4720 3224 4742 3226
rect 4820 3224 5012 3236
rect 5091 3224 5104 3254
rect 5119 3240 5149 3254
rect 5186 3224 5205 3254
rect 5220 3224 5226 3254
rect 5235 3224 5248 3254
rect 5263 3240 5293 3254
rect 5336 3240 5379 3254
rect 5386 3240 5606 3254
rect 5613 3240 5643 3254
rect 5303 3226 5318 3238
rect 5337 3226 5350 3240
rect 5418 3236 5571 3240
rect 5300 3224 5322 3226
rect 5400 3224 5592 3236
rect 5671 3224 5684 3254
rect 5699 3240 5729 3254
rect 5766 3224 5785 3254
rect 5800 3224 5806 3254
rect 5815 3224 5828 3254
rect 5843 3240 5873 3254
rect 5916 3240 5959 3254
rect 5966 3240 6186 3254
rect 6193 3240 6223 3254
rect 5883 3226 5898 3238
rect 5917 3226 5930 3240
rect 5998 3236 6151 3240
rect 5880 3224 5902 3226
rect 5980 3224 6172 3236
rect 6251 3224 6264 3254
rect 6279 3240 6309 3254
rect 6346 3224 6365 3254
rect 6380 3224 6386 3254
rect 6395 3224 6408 3254
rect 6423 3240 6453 3254
rect 6496 3240 6539 3254
rect 6546 3240 6766 3254
rect 6773 3240 6803 3254
rect 6463 3226 6478 3238
rect 6497 3226 6510 3240
rect 6578 3236 6731 3240
rect 6460 3224 6482 3226
rect 6560 3224 6752 3236
rect 6831 3224 6844 3254
rect 6859 3240 6889 3254
rect 6926 3224 6945 3254
rect 6960 3224 6966 3254
rect 6975 3224 6988 3254
rect 7003 3240 7033 3254
rect 7076 3240 7119 3254
rect 7126 3240 7346 3254
rect 7353 3240 7383 3254
rect 7043 3226 7058 3238
rect 7077 3226 7090 3240
rect 7158 3236 7311 3240
rect 7040 3224 7062 3226
rect 7140 3224 7332 3236
rect 7411 3224 7424 3254
rect 7439 3240 7469 3254
rect 7506 3224 7525 3254
rect 7540 3224 7546 3254
rect 7555 3224 7568 3254
rect 7583 3236 7613 3254
rect 7656 3240 7670 3254
rect 7706 3240 7926 3254
rect 7657 3238 7670 3240
rect 7623 3226 7638 3238
rect 7620 3224 7642 3226
rect 7647 3224 7677 3238
rect 7738 3236 7891 3240
rect 7720 3224 7912 3236
rect 7955 3224 7985 3238
rect 7991 3224 8004 3254
rect 8019 3236 8049 3254
rect 8092 3224 8105 3254
rect 8135 3224 8148 3254
rect 8163 3236 8193 3254
rect 8236 3240 8250 3254
rect 8286 3240 8506 3254
rect 8237 3238 8250 3240
rect 8203 3226 8218 3238
rect 8200 3224 8222 3226
rect 8227 3224 8257 3238
rect 8318 3236 8471 3240
rect 8300 3224 8492 3236
rect 8535 3224 8565 3238
rect 8571 3224 8584 3254
rect 8599 3236 8629 3254
rect 8672 3224 8685 3254
rect 8715 3224 8728 3254
rect 8743 3236 8773 3254
rect 8816 3240 8830 3254
rect 8866 3240 9086 3254
rect 8817 3238 8830 3240
rect 8783 3226 8798 3238
rect 8780 3224 8802 3226
rect 8807 3224 8837 3238
rect 8898 3236 9051 3240
rect 8880 3224 9072 3236
rect 9115 3224 9145 3238
rect 9151 3224 9164 3254
rect 9179 3236 9209 3254
rect 9252 3224 9265 3254
rect 0 3210 9265 3224
rect 15 3140 28 3210
rect 80 3206 102 3210
rect 73 3184 102 3198
rect 155 3184 171 3198
rect 209 3194 215 3196
rect 222 3194 330 3210
rect 337 3194 343 3196
rect 351 3194 366 3210
rect 432 3204 451 3207
rect 73 3182 171 3184
rect 198 3182 366 3194
rect 381 3184 397 3198
rect 432 3185 454 3204
rect 464 3198 480 3199
rect 463 3196 480 3198
rect 464 3191 480 3196
rect 454 3184 460 3185
rect 463 3184 492 3191
rect 381 3183 492 3184
rect 381 3182 498 3183
rect 57 3174 108 3182
rect 155 3174 189 3182
rect 57 3162 82 3174
rect 89 3162 108 3174
rect 162 3172 189 3174
rect 198 3172 419 3182
rect 454 3179 460 3182
rect 162 3168 419 3172
rect 57 3154 108 3162
rect 155 3154 419 3168
rect 463 3174 498 3182
rect 9 3106 28 3140
rect 73 3146 102 3154
rect 73 3140 90 3146
rect 73 3138 107 3140
rect 155 3138 171 3154
rect 172 3144 380 3154
rect 381 3144 397 3154
rect 445 3150 460 3165
rect 463 3162 464 3174
rect 471 3162 498 3174
rect 463 3154 498 3162
rect 463 3153 492 3154
rect 183 3140 397 3144
rect 198 3138 397 3140
rect 432 3140 445 3150
rect 463 3140 480 3153
rect 432 3138 480 3140
rect 74 3134 107 3138
rect 70 3132 107 3134
rect 70 3131 137 3132
rect 70 3126 101 3131
rect 107 3126 137 3131
rect 70 3122 137 3126
rect 43 3119 137 3122
rect 43 3112 92 3119
rect 43 3106 73 3112
rect 92 3107 97 3112
rect 9 3090 89 3106
rect 101 3098 137 3119
rect 198 3114 387 3138
rect 432 3137 479 3138
rect 445 3132 479 3137
rect 213 3111 387 3114
rect 206 3108 387 3111
rect 415 3131 479 3132
rect 9 3088 28 3090
rect 43 3088 77 3090
rect 9 3072 89 3088
rect 9 3066 28 3072
rect -1 3050 28 3066
rect 43 3056 73 3072
rect 101 3050 107 3098
rect 110 3092 129 3098
rect 144 3092 174 3100
rect 110 3084 174 3092
rect 110 3068 190 3084
rect 206 3077 268 3108
rect 284 3077 346 3108
rect 415 3106 464 3131
rect 479 3106 509 3122
rect 378 3092 408 3100
rect 415 3098 525 3106
rect 378 3084 423 3092
rect 110 3066 129 3068
rect 144 3066 190 3068
rect 110 3050 190 3066
rect 217 3064 252 3077
rect 293 3074 330 3077
rect 293 3072 335 3074
rect 222 3061 252 3064
rect 231 3057 238 3061
rect 238 3056 239 3057
rect 197 3050 207 3056
rect -7 3042 34 3050
rect -7 3016 8 3042
rect 15 3016 34 3042
rect 98 3038 129 3050
rect 144 3038 247 3050
rect 259 3040 285 3066
rect 300 3061 330 3072
rect 362 3068 424 3084
rect 362 3066 408 3068
rect 362 3050 424 3066
rect 436 3050 442 3098
rect 445 3090 525 3098
rect 445 3088 464 3090
rect 479 3088 513 3090
rect 445 3072 525 3088
rect 445 3050 464 3072
rect 479 3056 509 3072
rect 537 3066 543 3140
rect 546 3066 565 3210
rect 580 3066 586 3210
rect 595 3140 608 3210
rect 660 3206 682 3210
rect 653 3184 682 3198
rect 735 3184 751 3198
rect 789 3194 795 3196
rect 802 3194 910 3210
rect 917 3194 923 3196
rect 931 3194 946 3210
rect 1012 3204 1031 3207
rect 653 3182 751 3184
rect 778 3182 946 3194
rect 961 3184 977 3198
rect 1012 3185 1034 3204
rect 1044 3198 1060 3199
rect 1043 3196 1060 3198
rect 1044 3191 1060 3196
rect 1034 3184 1040 3185
rect 1043 3184 1072 3191
rect 961 3183 1072 3184
rect 961 3182 1078 3183
rect 637 3174 688 3182
rect 735 3174 769 3182
rect 637 3162 662 3174
rect 669 3162 688 3174
rect 742 3172 769 3174
rect 778 3172 999 3182
rect 1034 3179 1040 3182
rect 742 3168 999 3172
rect 637 3154 688 3162
rect 735 3154 999 3168
rect 1043 3174 1078 3182
rect 589 3106 608 3140
rect 653 3146 682 3154
rect 653 3140 670 3146
rect 653 3138 687 3140
rect 735 3138 751 3154
rect 752 3144 960 3154
rect 961 3144 977 3154
rect 1025 3150 1040 3165
rect 1043 3162 1044 3174
rect 1051 3162 1078 3174
rect 1043 3154 1078 3162
rect 1043 3153 1072 3154
rect 763 3140 977 3144
rect 778 3138 977 3140
rect 1012 3140 1025 3150
rect 1043 3140 1060 3153
rect 1012 3138 1060 3140
rect 654 3134 687 3138
rect 650 3132 687 3134
rect 650 3131 717 3132
rect 650 3126 681 3131
rect 687 3126 717 3131
rect 650 3122 717 3126
rect 623 3119 717 3122
rect 623 3112 672 3119
rect 623 3106 653 3112
rect 672 3107 677 3112
rect 589 3090 669 3106
rect 681 3098 717 3119
rect 778 3114 967 3138
rect 1012 3137 1059 3138
rect 1025 3132 1059 3137
rect 793 3111 967 3114
rect 786 3108 967 3111
rect 995 3131 1059 3132
rect 589 3088 608 3090
rect 623 3088 657 3090
rect 589 3072 669 3088
rect 589 3066 608 3072
rect 305 3040 408 3050
rect 259 3038 408 3040
rect 429 3038 464 3050
rect 98 3036 260 3038
rect 110 3016 129 3036
rect 144 3034 174 3036
rect -7 3008 34 3016
rect 116 3012 129 3016
rect 181 3020 260 3036
rect 292 3036 464 3038
rect 292 3020 371 3036
rect 378 3034 408 3036
rect -1 2998 28 3008
rect 43 2998 73 3012
rect 116 2998 159 3012
rect 181 3008 371 3020
rect 436 3016 442 3036
rect 166 2998 196 3008
rect 197 2998 355 3008
rect 359 2998 389 3008
rect 393 2998 423 3012
rect 451 2998 464 3036
rect 536 3050 565 3066
rect 579 3050 608 3066
rect 623 3056 653 3072
rect 681 3050 687 3098
rect 690 3092 709 3098
rect 724 3092 754 3100
rect 690 3084 754 3092
rect 690 3068 770 3084
rect 786 3077 848 3108
rect 864 3077 926 3108
rect 995 3106 1044 3131
rect 1059 3106 1089 3122
rect 958 3092 988 3100
rect 995 3098 1105 3106
rect 958 3084 1003 3092
rect 690 3066 709 3068
rect 724 3066 770 3068
rect 690 3050 770 3066
rect 797 3064 832 3077
rect 873 3074 910 3077
rect 873 3072 915 3074
rect 802 3061 832 3064
rect 811 3057 818 3061
rect 818 3056 819 3057
rect 777 3050 787 3056
rect 536 3042 571 3050
rect 536 3016 537 3042
rect 544 3016 571 3042
rect 479 2998 509 3012
rect 536 3008 571 3016
rect 573 3042 614 3050
rect 573 3016 588 3042
rect 595 3016 614 3042
rect 678 3038 709 3050
rect 724 3038 827 3050
rect 839 3040 865 3066
rect 880 3061 910 3072
rect 942 3068 1004 3084
rect 942 3066 988 3068
rect 942 3050 1004 3066
rect 1016 3050 1022 3098
rect 1025 3090 1105 3098
rect 1025 3088 1044 3090
rect 1059 3088 1093 3090
rect 1025 3072 1105 3088
rect 1025 3050 1044 3072
rect 1059 3056 1089 3072
rect 1117 3066 1123 3140
rect 1126 3066 1145 3210
rect 1160 3066 1166 3210
rect 1175 3140 1188 3210
rect 1240 3206 1262 3210
rect 1233 3184 1262 3198
rect 1315 3184 1331 3198
rect 1369 3194 1375 3196
rect 1382 3194 1490 3210
rect 1497 3194 1503 3196
rect 1511 3194 1526 3210
rect 1592 3204 1611 3207
rect 1233 3182 1331 3184
rect 1358 3182 1526 3194
rect 1541 3184 1557 3198
rect 1592 3185 1614 3204
rect 1624 3198 1640 3199
rect 1623 3196 1640 3198
rect 1624 3191 1640 3196
rect 1614 3184 1620 3185
rect 1623 3184 1652 3191
rect 1541 3183 1652 3184
rect 1541 3182 1658 3183
rect 1217 3174 1268 3182
rect 1315 3174 1349 3182
rect 1217 3162 1242 3174
rect 1249 3162 1268 3174
rect 1322 3172 1349 3174
rect 1358 3172 1579 3182
rect 1614 3179 1620 3182
rect 1322 3168 1579 3172
rect 1217 3154 1268 3162
rect 1315 3154 1579 3168
rect 1623 3174 1658 3182
rect 1169 3106 1188 3140
rect 1233 3146 1262 3154
rect 1233 3140 1250 3146
rect 1233 3138 1267 3140
rect 1315 3138 1331 3154
rect 1332 3144 1540 3154
rect 1541 3144 1557 3154
rect 1605 3150 1620 3165
rect 1623 3162 1624 3174
rect 1631 3162 1658 3174
rect 1623 3154 1658 3162
rect 1623 3153 1652 3154
rect 1343 3140 1557 3144
rect 1358 3138 1557 3140
rect 1592 3140 1605 3150
rect 1623 3140 1640 3153
rect 1592 3138 1640 3140
rect 1234 3134 1267 3138
rect 1230 3132 1267 3134
rect 1230 3131 1297 3132
rect 1230 3126 1261 3131
rect 1267 3126 1297 3131
rect 1230 3122 1297 3126
rect 1203 3119 1297 3122
rect 1203 3112 1252 3119
rect 1203 3106 1233 3112
rect 1252 3107 1257 3112
rect 1169 3090 1249 3106
rect 1261 3098 1297 3119
rect 1358 3114 1547 3138
rect 1592 3137 1639 3138
rect 1605 3132 1639 3137
rect 1373 3111 1547 3114
rect 1366 3108 1547 3111
rect 1575 3131 1639 3132
rect 1169 3088 1188 3090
rect 1203 3088 1237 3090
rect 1169 3072 1249 3088
rect 1169 3066 1188 3072
rect 885 3040 988 3050
rect 839 3038 988 3040
rect 1009 3038 1044 3050
rect 678 3036 840 3038
rect 690 3016 709 3036
rect 724 3034 754 3036
rect 573 3008 614 3016
rect 696 3012 709 3016
rect 761 3020 840 3036
rect 872 3036 1044 3038
rect 872 3020 951 3036
rect 958 3034 988 3036
rect 536 2998 565 3008
rect 579 2998 608 3008
rect 623 2998 653 3012
rect 696 2998 739 3012
rect 761 3008 951 3020
rect 1016 3016 1022 3036
rect 746 2998 776 3008
rect 777 2998 935 3008
rect 939 2998 969 3008
rect 973 2998 1003 3012
rect 1031 2998 1044 3036
rect 1116 3050 1145 3066
rect 1159 3050 1188 3066
rect 1203 3056 1233 3072
rect 1261 3050 1267 3098
rect 1270 3092 1289 3098
rect 1304 3092 1334 3100
rect 1270 3084 1334 3092
rect 1270 3068 1350 3084
rect 1366 3077 1428 3108
rect 1444 3077 1506 3108
rect 1575 3106 1624 3131
rect 1639 3106 1669 3122
rect 1538 3092 1568 3100
rect 1575 3098 1685 3106
rect 1538 3084 1583 3092
rect 1270 3066 1289 3068
rect 1304 3066 1350 3068
rect 1270 3050 1350 3066
rect 1377 3064 1412 3077
rect 1453 3074 1490 3077
rect 1453 3072 1495 3074
rect 1382 3061 1412 3064
rect 1391 3057 1398 3061
rect 1398 3056 1399 3057
rect 1357 3050 1367 3056
rect 1116 3042 1151 3050
rect 1116 3016 1117 3042
rect 1124 3016 1151 3042
rect 1059 2998 1089 3012
rect 1116 3008 1151 3016
rect 1153 3042 1194 3050
rect 1153 3016 1168 3042
rect 1175 3016 1194 3042
rect 1258 3038 1289 3050
rect 1304 3038 1407 3050
rect 1419 3040 1445 3066
rect 1460 3061 1490 3072
rect 1522 3068 1584 3084
rect 1522 3066 1568 3068
rect 1522 3050 1584 3066
rect 1596 3050 1602 3098
rect 1605 3090 1685 3098
rect 1605 3088 1624 3090
rect 1639 3088 1673 3090
rect 1605 3072 1685 3088
rect 1605 3050 1624 3072
rect 1639 3056 1669 3072
rect 1697 3066 1703 3140
rect 1706 3066 1725 3210
rect 1740 3066 1746 3210
rect 1755 3140 1768 3210
rect 1820 3206 1842 3210
rect 1813 3184 1842 3198
rect 1895 3184 1911 3198
rect 1949 3194 1955 3196
rect 1962 3194 2070 3210
rect 2077 3194 2083 3196
rect 2091 3194 2106 3210
rect 2172 3204 2191 3207
rect 1813 3182 1911 3184
rect 1938 3182 2106 3194
rect 2121 3184 2137 3198
rect 2172 3185 2194 3204
rect 2204 3198 2220 3199
rect 2203 3196 2220 3198
rect 2204 3191 2220 3196
rect 2194 3184 2200 3185
rect 2203 3184 2232 3191
rect 2121 3183 2232 3184
rect 2121 3182 2238 3183
rect 1797 3174 1848 3182
rect 1895 3174 1929 3182
rect 1797 3162 1822 3174
rect 1829 3162 1848 3174
rect 1902 3172 1929 3174
rect 1938 3172 2159 3182
rect 2194 3179 2200 3182
rect 1902 3168 2159 3172
rect 1797 3154 1848 3162
rect 1895 3154 2159 3168
rect 2203 3174 2238 3182
rect 1749 3106 1768 3140
rect 1813 3146 1842 3154
rect 1813 3140 1830 3146
rect 1813 3138 1847 3140
rect 1895 3138 1911 3154
rect 1912 3144 2120 3154
rect 2121 3144 2137 3154
rect 2185 3150 2200 3165
rect 2203 3162 2204 3174
rect 2211 3162 2238 3174
rect 2203 3154 2238 3162
rect 2203 3153 2232 3154
rect 1923 3140 2137 3144
rect 1938 3138 2137 3140
rect 2172 3140 2185 3150
rect 2203 3140 2220 3153
rect 2172 3138 2220 3140
rect 1814 3134 1847 3138
rect 1810 3132 1847 3134
rect 1810 3131 1877 3132
rect 1810 3126 1841 3131
rect 1847 3126 1877 3131
rect 1810 3122 1877 3126
rect 1783 3119 1877 3122
rect 1783 3112 1832 3119
rect 1783 3106 1813 3112
rect 1832 3107 1837 3112
rect 1749 3090 1829 3106
rect 1841 3098 1877 3119
rect 1938 3114 2127 3138
rect 2172 3137 2219 3138
rect 2185 3132 2219 3137
rect 1953 3111 2127 3114
rect 1946 3108 2127 3111
rect 2155 3131 2219 3132
rect 1749 3088 1768 3090
rect 1783 3088 1817 3090
rect 1749 3072 1829 3088
rect 1749 3066 1768 3072
rect 1465 3040 1568 3050
rect 1419 3038 1568 3040
rect 1589 3038 1624 3050
rect 1258 3036 1420 3038
rect 1270 3016 1289 3036
rect 1304 3034 1334 3036
rect 1153 3008 1194 3016
rect 1276 3012 1289 3016
rect 1341 3020 1420 3036
rect 1452 3036 1624 3038
rect 1452 3020 1531 3036
rect 1538 3034 1568 3036
rect 1116 2998 1145 3008
rect 1159 2998 1188 3008
rect 1203 2998 1233 3012
rect 1276 2998 1319 3012
rect 1341 3008 1531 3020
rect 1596 3016 1602 3036
rect 1326 2998 1356 3008
rect 1357 2998 1515 3008
rect 1519 2998 1549 3008
rect 1553 2998 1583 3012
rect 1611 2998 1624 3036
rect 1696 3050 1725 3066
rect 1739 3050 1768 3066
rect 1783 3056 1813 3072
rect 1841 3050 1847 3098
rect 1850 3092 1869 3098
rect 1884 3092 1914 3100
rect 1850 3084 1914 3092
rect 1850 3068 1930 3084
rect 1946 3077 2008 3108
rect 2024 3077 2086 3108
rect 2155 3106 2204 3131
rect 2219 3106 2249 3122
rect 2118 3092 2148 3100
rect 2155 3098 2265 3106
rect 2118 3084 2163 3092
rect 1850 3066 1869 3068
rect 1884 3066 1930 3068
rect 1850 3050 1930 3066
rect 1957 3064 1992 3077
rect 2033 3074 2070 3077
rect 2033 3072 2075 3074
rect 1962 3061 1992 3064
rect 1971 3057 1978 3061
rect 1978 3056 1979 3057
rect 1937 3050 1947 3056
rect 1696 3042 1731 3050
rect 1696 3016 1697 3042
rect 1704 3016 1731 3042
rect 1639 2998 1669 3012
rect 1696 3008 1731 3016
rect 1733 3042 1774 3050
rect 1733 3016 1748 3042
rect 1755 3016 1774 3042
rect 1838 3038 1869 3050
rect 1884 3038 1987 3050
rect 1999 3040 2025 3066
rect 2040 3061 2070 3072
rect 2102 3068 2164 3084
rect 2102 3066 2148 3068
rect 2102 3050 2164 3066
rect 2176 3050 2182 3098
rect 2185 3090 2265 3098
rect 2185 3088 2204 3090
rect 2219 3088 2253 3090
rect 2185 3072 2265 3088
rect 2185 3050 2204 3072
rect 2219 3056 2249 3072
rect 2277 3066 2283 3140
rect 2286 3066 2305 3210
rect 2320 3066 2326 3210
rect 2335 3140 2348 3210
rect 2400 3206 2422 3210
rect 2393 3184 2422 3198
rect 2475 3184 2491 3198
rect 2529 3194 2535 3196
rect 2542 3194 2650 3210
rect 2657 3194 2663 3196
rect 2671 3194 2686 3210
rect 2752 3204 2771 3207
rect 2393 3182 2491 3184
rect 2518 3182 2686 3194
rect 2701 3184 2717 3198
rect 2752 3185 2774 3204
rect 2784 3198 2800 3199
rect 2783 3196 2800 3198
rect 2784 3191 2800 3196
rect 2774 3184 2780 3185
rect 2783 3184 2812 3191
rect 2701 3183 2812 3184
rect 2701 3182 2818 3183
rect 2377 3174 2428 3182
rect 2475 3174 2509 3182
rect 2377 3162 2402 3174
rect 2409 3162 2428 3174
rect 2482 3172 2509 3174
rect 2518 3172 2739 3182
rect 2774 3179 2780 3182
rect 2482 3168 2739 3172
rect 2377 3154 2428 3162
rect 2475 3154 2739 3168
rect 2783 3174 2818 3182
rect 2329 3106 2348 3140
rect 2393 3146 2422 3154
rect 2393 3140 2410 3146
rect 2393 3138 2427 3140
rect 2475 3138 2491 3154
rect 2492 3144 2700 3154
rect 2701 3144 2717 3154
rect 2765 3150 2780 3165
rect 2783 3162 2784 3174
rect 2791 3162 2818 3174
rect 2783 3154 2818 3162
rect 2783 3153 2812 3154
rect 2503 3140 2717 3144
rect 2518 3138 2717 3140
rect 2752 3140 2765 3150
rect 2783 3140 2800 3153
rect 2752 3138 2800 3140
rect 2394 3134 2427 3138
rect 2390 3132 2427 3134
rect 2390 3131 2457 3132
rect 2390 3126 2421 3131
rect 2427 3126 2457 3131
rect 2390 3122 2457 3126
rect 2363 3119 2457 3122
rect 2363 3112 2412 3119
rect 2363 3106 2393 3112
rect 2412 3107 2417 3112
rect 2329 3090 2409 3106
rect 2421 3098 2457 3119
rect 2518 3114 2707 3138
rect 2752 3137 2799 3138
rect 2765 3132 2799 3137
rect 2533 3111 2707 3114
rect 2526 3108 2707 3111
rect 2735 3131 2799 3132
rect 2329 3088 2348 3090
rect 2363 3088 2397 3090
rect 2329 3072 2409 3088
rect 2329 3066 2348 3072
rect 2045 3040 2148 3050
rect 1999 3038 2148 3040
rect 2169 3038 2204 3050
rect 1838 3036 2000 3038
rect 1850 3016 1869 3036
rect 1884 3034 1914 3036
rect 1733 3008 1774 3016
rect 1856 3012 1869 3016
rect 1921 3020 2000 3036
rect 2032 3036 2204 3038
rect 2032 3020 2111 3036
rect 2118 3034 2148 3036
rect 1696 2998 1725 3008
rect 1739 2998 1768 3008
rect 1783 2998 1813 3012
rect 1856 2998 1899 3012
rect 1921 3008 2111 3020
rect 2176 3016 2182 3036
rect 1906 2998 1936 3008
rect 1937 2998 2095 3008
rect 2099 2998 2129 3008
rect 2133 2998 2163 3012
rect 2191 2998 2204 3036
rect 2276 3050 2305 3066
rect 2319 3050 2348 3066
rect 2363 3056 2393 3072
rect 2421 3050 2427 3098
rect 2430 3092 2449 3098
rect 2464 3092 2494 3100
rect 2430 3084 2494 3092
rect 2430 3068 2510 3084
rect 2526 3077 2588 3108
rect 2604 3077 2666 3108
rect 2735 3106 2784 3131
rect 2799 3106 2829 3122
rect 2698 3092 2728 3100
rect 2735 3098 2845 3106
rect 2698 3084 2743 3092
rect 2430 3066 2449 3068
rect 2464 3066 2510 3068
rect 2430 3050 2510 3066
rect 2537 3064 2572 3077
rect 2613 3074 2650 3077
rect 2613 3072 2655 3074
rect 2542 3061 2572 3064
rect 2551 3057 2558 3061
rect 2558 3056 2559 3057
rect 2517 3050 2527 3056
rect 2276 3042 2311 3050
rect 2276 3016 2277 3042
rect 2284 3016 2311 3042
rect 2219 2998 2249 3012
rect 2276 3008 2311 3016
rect 2313 3042 2354 3050
rect 2313 3016 2328 3042
rect 2335 3016 2354 3042
rect 2418 3038 2449 3050
rect 2464 3038 2567 3050
rect 2579 3040 2605 3066
rect 2620 3061 2650 3072
rect 2682 3068 2744 3084
rect 2682 3066 2728 3068
rect 2682 3050 2744 3066
rect 2756 3050 2762 3098
rect 2765 3090 2845 3098
rect 2765 3088 2784 3090
rect 2799 3088 2833 3090
rect 2765 3072 2845 3088
rect 2765 3050 2784 3072
rect 2799 3056 2829 3072
rect 2857 3066 2863 3140
rect 2866 3066 2885 3210
rect 2900 3066 2906 3210
rect 2915 3140 2928 3210
rect 2980 3206 3002 3210
rect 2973 3184 3002 3198
rect 3055 3184 3071 3198
rect 3109 3194 3115 3196
rect 3122 3194 3230 3210
rect 3237 3194 3243 3196
rect 3251 3194 3266 3210
rect 3332 3204 3351 3207
rect 2973 3182 3071 3184
rect 3098 3182 3266 3194
rect 3281 3184 3297 3198
rect 3332 3185 3354 3204
rect 3364 3198 3380 3199
rect 3363 3196 3380 3198
rect 3364 3191 3380 3196
rect 3354 3184 3360 3185
rect 3363 3184 3392 3191
rect 3281 3183 3392 3184
rect 3281 3182 3398 3183
rect 2957 3174 3008 3182
rect 3055 3174 3089 3182
rect 2957 3162 2982 3174
rect 2989 3162 3008 3174
rect 3062 3172 3089 3174
rect 3098 3172 3319 3182
rect 3354 3179 3360 3182
rect 3062 3168 3319 3172
rect 2957 3154 3008 3162
rect 3055 3154 3319 3168
rect 3363 3174 3398 3182
rect 2909 3106 2928 3140
rect 2973 3146 3002 3154
rect 2973 3140 2990 3146
rect 2973 3138 3007 3140
rect 3055 3138 3071 3154
rect 3072 3144 3280 3154
rect 3281 3144 3297 3154
rect 3345 3150 3360 3165
rect 3363 3162 3364 3174
rect 3371 3162 3398 3174
rect 3363 3154 3398 3162
rect 3363 3153 3392 3154
rect 3083 3140 3297 3144
rect 3098 3138 3297 3140
rect 3332 3140 3345 3150
rect 3363 3140 3380 3153
rect 3332 3138 3380 3140
rect 2974 3134 3007 3138
rect 2970 3132 3007 3134
rect 2970 3131 3037 3132
rect 2970 3126 3001 3131
rect 3007 3126 3037 3131
rect 2970 3122 3037 3126
rect 2943 3119 3037 3122
rect 2943 3112 2992 3119
rect 2943 3106 2973 3112
rect 2992 3107 2997 3112
rect 2909 3090 2989 3106
rect 3001 3098 3037 3119
rect 3098 3114 3287 3138
rect 3332 3137 3379 3138
rect 3345 3132 3379 3137
rect 3113 3111 3287 3114
rect 3106 3108 3287 3111
rect 3315 3131 3379 3132
rect 2909 3088 2928 3090
rect 2943 3088 2977 3090
rect 2909 3072 2989 3088
rect 2909 3066 2928 3072
rect 2625 3040 2728 3050
rect 2579 3038 2728 3040
rect 2749 3038 2784 3050
rect 2418 3036 2580 3038
rect 2430 3016 2449 3036
rect 2464 3034 2494 3036
rect 2313 3008 2354 3016
rect 2436 3012 2449 3016
rect 2501 3020 2580 3036
rect 2612 3036 2784 3038
rect 2612 3020 2691 3036
rect 2698 3034 2728 3036
rect 2276 2998 2305 3008
rect 2319 2998 2348 3008
rect 2363 2998 2393 3012
rect 2436 2998 2479 3012
rect 2501 3008 2691 3020
rect 2756 3016 2762 3036
rect 2486 2998 2516 3008
rect 2517 2998 2675 3008
rect 2679 2998 2709 3008
rect 2713 2998 2743 3012
rect 2771 2998 2784 3036
rect 2856 3050 2885 3066
rect 2899 3050 2928 3066
rect 2943 3056 2973 3072
rect 3001 3050 3007 3098
rect 3010 3092 3029 3098
rect 3044 3092 3074 3100
rect 3010 3084 3074 3092
rect 3010 3068 3090 3084
rect 3106 3077 3168 3108
rect 3184 3077 3246 3108
rect 3315 3106 3364 3131
rect 3379 3106 3409 3122
rect 3278 3092 3308 3100
rect 3315 3098 3425 3106
rect 3278 3084 3323 3092
rect 3010 3066 3029 3068
rect 3044 3066 3090 3068
rect 3010 3050 3090 3066
rect 3117 3064 3152 3077
rect 3193 3074 3230 3077
rect 3193 3072 3235 3074
rect 3122 3061 3152 3064
rect 3131 3057 3138 3061
rect 3138 3056 3139 3057
rect 3097 3050 3107 3056
rect 2856 3042 2891 3050
rect 2856 3016 2857 3042
rect 2864 3016 2891 3042
rect 2799 2998 2829 3012
rect 2856 3008 2891 3016
rect 2893 3042 2934 3050
rect 2893 3016 2908 3042
rect 2915 3016 2934 3042
rect 2998 3038 3029 3050
rect 3044 3038 3147 3050
rect 3159 3040 3185 3066
rect 3200 3061 3230 3072
rect 3262 3068 3324 3084
rect 3262 3066 3308 3068
rect 3262 3050 3324 3066
rect 3336 3050 3342 3098
rect 3345 3090 3425 3098
rect 3345 3088 3364 3090
rect 3379 3088 3413 3090
rect 3345 3072 3425 3088
rect 3345 3050 3364 3072
rect 3379 3056 3409 3072
rect 3437 3066 3443 3140
rect 3446 3066 3465 3210
rect 3480 3066 3486 3210
rect 3495 3140 3508 3210
rect 3560 3206 3582 3210
rect 3553 3184 3582 3198
rect 3635 3184 3651 3198
rect 3689 3194 3695 3196
rect 3702 3194 3810 3210
rect 3817 3194 3823 3196
rect 3831 3194 3846 3210
rect 3912 3204 3931 3207
rect 3553 3182 3651 3184
rect 3678 3182 3846 3194
rect 3861 3184 3877 3198
rect 3912 3185 3934 3204
rect 3944 3198 3960 3199
rect 3943 3196 3960 3198
rect 3944 3191 3960 3196
rect 3934 3184 3940 3185
rect 3943 3184 3972 3191
rect 3861 3183 3972 3184
rect 3861 3182 3978 3183
rect 3537 3174 3588 3182
rect 3635 3174 3669 3182
rect 3537 3162 3562 3174
rect 3569 3162 3588 3174
rect 3642 3172 3669 3174
rect 3678 3172 3899 3182
rect 3934 3179 3940 3182
rect 3642 3168 3899 3172
rect 3537 3154 3588 3162
rect 3635 3154 3899 3168
rect 3943 3174 3978 3182
rect 3489 3106 3508 3140
rect 3553 3146 3582 3154
rect 3553 3140 3570 3146
rect 3553 3138 3587 3140
rect 3635 3138 3651 3154
rect 3652 3144 3860 3154
rect 3861 3144 3877 3154
rect 3925 3150 3940 3165
rect 3943 3162 3944 3174
rect 3951 3162 3978 3174
rect 3943 3154 3978 3162
rect 3943 3153 3972 3154
rect 3663 3140 3877 3144
rect 3678 3138 3877 3140
rect 3912 3140 3925 3150
rect 3943 3140 3960 3153
rect 3912 3138 3960 3140
rect 3554 3134 3587 3138
rect 3550 3132 3587 3134
rect 3550 3131 3617 3132
rect 3550 3126 3581 3131
rect 3587 3126 3617 3131
rect 3550 3122 3617 3126
rect 3523 3119 3617 3122
rect 3523 3112 3572 3119
rect 3523 3106 3553 3112
rect 3572 3107 3577 3112
rect 3489 3090 3569 3106
rect 3581 3098 3617 3119
rect 3678 3114 3867 3138
rect 3912 3137 3959 3138
rect 3925 3132 3959 3137
rect 3693 3111 3867 3114
rect 3686 3108 3867 3111
rect 3895 3131 3959 3132
rect 3489 3088 3508 3090
rect 3523 3088 3557 3090
rect 3489 3072 3569 3088
rect 3489 3066 3508 3072
rect 3205 3040 3308 3050
rect 3159 3038 3308 3040
rect 3329 3038 3364 3050
rect 2998 3036 3160 3038
rect 3010 3016 3029 3036
rect 3044 3034 3074 3036
rect 2893 3008 2934 3016
rect 3016 3012 3029 3016
rect 3081 3020 3160 3036
rect 3192 3036 3364 3038
rect 3192 3020 3271 3036
rect 3278 3034 3308 3036
rect 2856 2998 2885 3008
rect 2899 2998 2928 3008
rect 2943 2998 2973 3012
rect 3016 2998 3059 3012
rect 3081 3008 3271 3020
rect 3336 3016 3342 3036
rect 3066 2998 3096 3008
rect 3097 2998 3255 3008
rect 3259 2998 3289 3008
rect 3293 2998 3323 3012
rect 3351 2998 3364 3036
rect 3436 3050 3465 3066
rect 3479 3050 3508 3066
rect 3523 3056 3553 3072
rect 3581 3050 3587 3098
rect 3590 3092 3609 3098
rect 3624 3092 3654 3100
rect 3590 3084 3654 3092
rect 3590 3068 3670 3084
rect 3686 3077 3748 3108
rect 3764 3077 3826 3108
rect 3895 3106 3944 3131
rect 3959 3106 3989 3122
rect 3858 3092 3888 3100
rect 3895 3098 4005 3106
rect 3858 3084 3903 3092
rect 3590 3066 3609 3068
rect 3624 3066 3670 3068
rect 3590 3050 3670 3066
rect 3697 3064 3732 3077
rect 3773 3074 3810 3077
rect 3773 3072 3815 3074
rect 3702 3061 3732 3064
rect 3711 3057 3718 3061
rect 3718 3056 3719 3057
rect 3677 3050 3687 3056
rect 3436 3042 3471 3050
rect 3436 3016 3437 3042
rect 3444 3016 3471 3042
rect 3379 2998 3409 3012
rect 3436 3008 3471 3016
rect 3473 3042 3514 3050
rect 3473 3016 3488 3042
rect 3495 3016 3514 3042
rect 3578 3038 3609 3050
rect 3624 3038 3727 3050
rect 3739 3040 3765 3066
rect 3780 3061 3810 3072
rect 3842 3068 3904 3084
rect 3842 3066 3888 3068
rect 3842 3050 3904 3066
rect 3916 3050 3922 3098
rect 3925 3090 4005 3098
rect 3925 3088 3944 3090
rect 3959 3088 3993 3090
rect 3925 3072 4005 3088
rect 3925 3050 3944 3072
rect 3959 3056 3989 3072
rect 4017 3066 4023 3140
rect 4026 3066 4045 3210
rect 4060 3066 4066 3210
rect 4075 3140 4088 3210
rect 4140 3206 4162 3210
rect 4133 3184 4162 3198
rect 4215 3184 4231 3198
rect 4269 3194 4275 3196
rect 4282 3194 4390 3210
rect 4397 3194 4403 3196
rect 4411 3194 4426 3210
rect 4492 3204 4511 3207
rect 4133 3182 4231 3184
rect 4258 3182 4426 3194
rect 4441 3184 4457 3198
rect 4492 3185 4514 3204
rect 4524 3198 4540 3199
rect 4523 3196 4540 3198
rect 4524 3191 4540 3196
rect 4514 3184 4520 3185
rect 4523 3184 4552 3191
rect 4441 3183 4552 3184
rect 4441 3182 4558 3183
rect 4117 3174 4168 3182
rect 4215 3174 4249 3182
rect 4117 3162 4142 3174
rect 4149 3162 4168 3174
rect 4222 3172 4249 3174
rect 4258 3172 4479 3182
rect 4514 3179 4520 3182
rect 4222 3168 4479 3172
rect 4117 3154 4168 3162
rect 4215 3154 4479 3168
rect 4523 3174 4558 3182
rect 4069 3106 4088 3140
rect 4133 3146 4162 3154
rect 4133 3140 4150 3146
rect 4133 3138 4167 3140
rect 4215 3138 4231 3154
rect 4232 3144 4440 3154
rect 4441 3144 4457 3154
rect 4505 3150 4520 3165
rect 4523 3162 4524 3174
rect 4531 3162 4558 3174
rect 4523 3154 4558 3162
rect 4523 3153 4552 3154
rect 4243 3140 4457 3144
rect 4258 3138 4457 3140
rect 4492 3140 4505 3150
rect 4523 3140 4540 3153
rect 4492 3138 4540 3140
rect 4134 3134 4167 3138
rect 4130 3132 4167 3134
rect 4130 3131 4197 3132
rect 4130 3126 4161 3131
rect 4167 3126 4197 3131
rect 4130 3122 4197 3126
rect 4103 3119 4197 3122
rect 4103 3112 4152 3119
rect 4103 3106 4133 3112
rect 4152 3107 4157 3112
rect 4069 3090 4149 3106
rect 4161 3098 4197 3119
rect 4258 3114 4447 3138
rect 4492 3137 4539 3138
rect 4505 3132 4539 3137
rect 4273 3111 4447 3114
rect 4266 3108 4447 3111
rect 4475 3131 4539 3132
rect 4069 3088 4088 3090
rect 4103 3088 4137 3090
rect 4069 3072 4149 3088
rect 4069 3066 4088 3072
rect 3785 3040 3888 3050
rect 3739 3038 3888 3040
rect 3909 3038 3944 3050
rect 3578 3036 3740 3038
rect 3590 3016 3609 3036
rect 3624 3034 3654 3036
rect 3473 3008 3514 3016
rect 3596 3012 3609 3016
rect 3661 3020 3740 3036
rect 3772 3036 3944 3038
rect 3772 3020 3851 3036
rect 3858 3034 3888 3036
rect 3436 2998 3465 3008
rect 3479 2998 3508 3008
rect 3523 2998 3553 3012
rect 3596 2998 3639 3012
rect 3661 3008 3851 3020
rect 3916 3016 3922 3036
rect 3646 2998 3676 3008
rect 3677 2998 3835 3008
rect 3839 2998 3869 3008
rect 3873 2998 3903 3012
rect 3931 2998 3944 3036
rect 4016 3050 4045 3066
rect 4059 3050 4088 3066
rect 4103 3056 4133 3072
rect 4161 3050 4167 3098
rect 4170 3092 4189 3098
rect 4204 3092 4234 3100
rect 4170 3084 4234 3092
rect 4170 3068 4250 3084
rect 4266 3077 4328 3108
rect 4344 3077 4406 3108
rect 4475 3106 4524 3131
rect 4539 3106 4569 3122
rect 4438 3092 4468 3100
rect 4475 3098 4585 3106
rect 4438 3084 4483 3092
rect 4170 3066 4189 3068
rect 4204 3066 4250 3068
rect 4170 3050 4250 3066
rect 4277 3064 4312 3077
rect 4353 3074 4390 3077
rect 4353 3072 4395 3074
rect 4282 3061 4312 3064
rect 4291 3057 4298 3061
rect 4298 3056 4299 3057
rect 4257 3050 4267 3056
rect 4016 3042 4051 3050
rect 4016 3016 4017 3042
rect 4024 3016 4051 3042
rect 3959 2998 3989 3012
rect 4016 3008 4051 3016
rect 4053 3042 4094 3050
rect 4053 3016 4068 3042
rect 4075 3016 4094 3042
rect 4158 3038 4189 3050
rect 4204 3038 4307 3050
rect 4319 3040 4345 3066
rect 4360 3061 4390 3072
rect 4422 3068 4484 3084
rect 4422 3066 4468 3068
rect 4422 3050 4484 3066
rect 4496 3050 4502 3098
rect 4505 3090 4585 3098
rect 4505 3088 4524 3090
rect 4539 3088 4573 3090
rect 4505 3072 4585 3088
rect 4505 3050 4524 3072
rect 4539 3056 4569 3072
rect 4597 3066 4603 3140
rect 4606 3066 4625 3210
rect 4640 3066 4646 3210
rect 4655 3140 4668 3210
rect 4720 3206 4742 3210
rect 4713 3184 4742 3198
rect 4795 3184 4811 3198
rect 4849 3194 4855 3196
rect 4862 3194 4970 3210
rect 4977 3194 4983 3196
rect 4991 3194 5006 3210
rect 5072 3204 5091 3207
rect 4713 3182 4811 3184
rect 4838 3182 5006 3194
rect 5021 3184 5037 3198
rect 5072 3185 5094 3204
rect 5104 3198 5120 3199
rect 5103 3196 5120 3198
rect 5104 3191 5120 3196
rect 5094 3184 5100 3185
rect 5103 3184 5132 3191
rect 5021 3183 5132 3184
rect 5021 3182 5138 3183
rect 4697 3174 4748 3182
rect 4795 3174 4829 3182
rect 4697 3162 4722 3174
rect 4729 3162 4748 3174
rect 4802 3172 4829 3174
rect 4838 3172 5059 3182
rect 5094 3179 5100 3182
rect 4802 3168 5059 3172
rect 4697 3154 4748 3162
rect 4795 3154 5059 3168
rect 5103 3174 5138 3182
rect 4649 3106 4668 3140
rect 4713 3146 4742 3154
rect 4713 3140 4730 3146
rect 4713 3138 4747 3140
rect 4795 3138 4811 3154
rect 4812 3144 5020 3154
rect 5021 3144 5037 3154
rect 5085 3150 5100 3165
rect 5103 3162 5104 3174
rect 5111 3162 5138 3174
rect 5103 3154 5138 3162
rect 5103 3153 5132 3154
rect 4823 3140 5037 3144
rect 4838 3138 5037 3140
rect 5072 3140 5085 3150
rect 5103 3140 5120 3153
rect 5072 3138 5120 3140
rect 4714 3134 4747 3138
rect 4710 3132 4747 3134
rect 4710 3131 4777 3132
rect 4710 3126 4741 3131
rect 4747 3126 4777 3131
rect 4710 3122 4777 3126
rect 4683 3119 4777 3122
rect 4683 3112 4732 3119
rect 4683 3106 4713 3112
rect 4732 3107 4737 3112
rect 4649 3090 4729 3106
rect 4741 3098 4777 3119
rect 4838 3114 5027 3138
rect 5072 3137 5119 3138
rect 5085 3132 5119 3137
rect 4853 3111 5027 3114
rect 4846 3108 5027 3111
rect 5055 3131 5119 3132
rect 4649 3088 4668 3090
rect 4683 3088 4717 3090
rect 4649 3072 4729 3088
rect 4649 3066 4668 3072
rect 4365 3040 4468 3050
rect 4319 3038 4468 3040
rect 4489 3038 4524 3050
rect 4158 3036 4320 3038
rect 4170 3016 4189 3036
rect 4204 3034 4234 3036
rect 4053 3008 4094 3016
rect 4176 3012 4189 3016
rect 4241 3020 4320 3036
rect 4352 3036 4524 3038
rect 4352 3020 4431 3036
rect 4438 3034 4468 3036
rect 4016 2998 4045 3008
rect 4059 2998 4088 3008
rect 4103 2998 4133 3012
rect 4176 2998 4219 3012
rect 4241 3008 4431 3020
rect 4496 3016 4502 3036
rect 4226 2998 4256 3008
rect 4257 2998 4415 3008
rect 4419 2998 4449 3008
rect 4453 2998 4483 3012
rect 4511 2998 4524 3036
rect 4596 3050 4625 3066
rect 4639 3050 4668 3066
rect 4683 3056 4713 3072
rect 4741 3050 4747 3098
rect 4750 3092 4769 3098
rect 4784 3092 4814 3100
rect 4750 3084 4814 3092
rect 4750 3068 4830 3084
rect 4846 3077 4908 3108
rect 4924 3077 4986 3108
rect 5055 3106 5104 3131
rect 5119 3106 5149 3122
rect 5018 3092 5048 3100
rect 5055 3098 5165 3106
rect 5018 3084 5063 3092
rect 4750 3066 4769 3068
rect 4784 3066 4830 3068
rect 4750 3050 4830 3066
rect 4857 3064 4892 3077
rect 4933 3074 4970 3077
rect 4933 3072 4975 3074
rect 4862 3061 4892 3064
rect 4871 3057 4878 3061
rect 4878 3056 4879 3057
rect 4837 3050 4847 3056
rect 4596 3042 4631 3050
rect 4596 3016 4597 3042
rect 4604 3016 4631 3042
rect 4539 2998 4569 3012
rect 4596 3008 4631 3016
rect 4633 3042 4674 3050
rect 4633 3016 4648 3042
rect 4655 3016 4674 3042
rect 4738 3038 4769 3050
rect 4784 3038 4887 3050
rect 4899 3040 4925 3066
rect 4940 3061 4970 3072
rect 5002 3068 5064 3084
rect 5002 3066 5048 3068
rect 5002 3050 5064 3066
rect 5076 3050 5082 3098
rect 5085 3090 5165 3098
rect 5085 3088 5104 3090
rect 5119 3088 5153 3090
rect 5085 3072 5165 3088
rect 5085 3050 5104 3072
rect 5119 3056 5149 3072
rect 5177 3066 5183 3140
rect 5186 3066 5205 3210
rect 5220 3066 5226 3210
rect 5235 3140 5248 3210
rect 5300 3206 5322 3210
rect 5293 3184 5322 3198
rect 5375 3184 5391 3198
rect 5429 3194 5435 3196
rect 5442 3194 5550 3210
rect 5557 3194 5563 3196
rect 5571 3194 5586 3210
rect 5652 3204 5671 3207
rect 5293 3182 5391 3184
rect 5418 3182 5586 3194
rect 5601 3184 5617 3198
rect 5652 3185 5674 3204
rect 5684 3198 5700 3199
rect 5683 3196 5700 3198
rect 5684 3191 5700 3196
rect 5674 3184 5680 3185
rect 5683 3184 5712 3191
rect 5601 3183 5712 3184
rect 5601 3182 5718 3183
rect 5277 3174 5328 3182
rect 5375 3174 5409 3182
rect 5277 3162 5302 3174
rect 5309 3162 5328 3174
rect 5382 3172 5409 3174
rect 5418 3172 5639 3182
rect 5674 3179 5680 3182
rect 5382 3168 5639 3172
rect 5277 3154 5328 3162
rect 5375 3154 5639 3168
rect 5683 3174 5718 3182
rect 5229 3106 5248 3140
rect 5293 3146 5322 3154
rect 5293 3140 5310 3146
rect 5293 3138 5327 3140
rect 5375 3138 5391 3154
rect 5392 3144 5600 3154
rect 5601 3144 5617 3154
rect 5665 3150 5680 3165
rect 5683 3162 5684 3174
rect 5691 3162 5718 3174
rect 5683 3154 5718 3162
rect 5683 3153 5712 3154
rect 5403 3140 5617 3144
rect 5418 3138 5617 3140
rect 5652 3140 5665 3150
rect 5683 3140 5700 3153
rect 5652 3138 5700 3140
rect 5294 3134 5327 3138
rect 5290 3132 5327 3134
rect 5290 3131 5357 3132
rect 5290 3126 5321 3131
rect 5327 3126 5357 3131
rect 5290 3122 5357 3126
rect 5263 3119 5357 3122
rect 5263 3112 5312 3119
rect 5263 3106 5293 3112
rect 5312 3107 5317 3112
rect 5229 3090 5309 3106
rect 5321 3098 5357 3119
rect 5418 3114 5607 3138
rect 5652 3137 5699 3138
rect 5665 3132 5699 3137
rect 5433 3111 5607 3114
rect 5426 3108 5607 3111
rect 5635 3131 5699 3132
rect 5229 3088 5248 3090
rect 5263 3088 5297 3090
rect 5229 3072 5309 3088
rect 5229 3066 5248 3072
rect 4945 3040 5048 3050
rect 4899 3038 5048 3040
rect 5069 3038 5104 3050
rect 4738 3036 4900 3038
rect 4750 3016 4769 3036
rect 4784 3034 4814 3036
rect 4633 3008 4674 3016
rect 4756 3012 4769 3016
rect 4821 3020 4900 3036
rect 4932 3036 5104 3038
rect 4932 3020 5011 3036
rect 5018 3034 5048 3036
rect 4596 2998 4625 3008
rect 4639 2998 4668 3008
rect 4683 2998 4713 3012
rect 4756 2998 4799 3012
rect 4821 3008 5011 3020
rect 5076 3016 5082 3036
rect 4806 2998 4836 3008
rect 4837 2998 4995 3008
rect 4999 2998 5029 3008
rect 5033 2998 5063 3012
rect 5091 2998 5104 3036
rect 5176 3050 5205 3066
rect 5219 3050 5248 3066
rect 5263 3056 5293 3072
rect 5321 3050 5327 3098
rect 5330 3092 5349 3098
rect 5364 3092 5394 3100
rect 5330 3084 5394 3092
rect 5330 3068 5410 3084
rect 5426 3077 5488 3108
rect 5504 3077 5566 3108
rect 5635 3106 5684 3131
rect 5699 3106 5729 3122
rect 5598 3092 5628 3100
rect 5635 3098 5745 3106
rect 5598 3084 5643 3092
rect 5330 3066 5349 3068
rect 5364 3066 5410 3068
rect 5330 3050 5410 3066
rect 5437 3064 5472 3077
rect 5513 3074 5550 3077
rect 5513 3072 5555 3074
rect 5442 3061 5472 3064
rect 5451 3057 5458 3061
rect 5458 3056 5459 3057
rect 5417 3050 5427 3056
rect 5176 3042 5211 3050
rect 5176 3016 5177 3042
rect 5184 3016 5211 3042
rect 5119 2998 5149 3012
rect 5176 3008 5211 3016
rect 5213 3042 5254 3050
rect 5213 3016 5228 3042
rect 5235 3016 5254 3042
rect 5318 3038 5349 3050
rect 5364 3038 5467 3050
rect 5479 3040 5505 3066
rect 5520 3061 5550 3072
rect 5582 3068 5644 3084
rect 5582 3066 5628 3068
rect 5582 3050 5644 3066
rect 5656 3050 5662 3098
rect 5665 3090 5745 3098
rect 5665 3088 5684 3090
rect 5699 3088 5733 3090
rect 5665 3072 5745 3088
rect 5665 3050 5684 3072
rect 5699 3056 5729 3072
rect 5757 3066 5763 3140
rect 5766 3066 5785 3210
rect 5800 3066 5806 3210
rect 5815 3140 5828 3210
rect 5880 3206 5902 3210
rect 5873 3184 5902 3198
rect 5955 3184 5971 3198
rect 6009 3194 6015 3196
rect 6022 3194 6130 3210
rect 6137 3194 6143 3196
rect 6151 3194 6166 3210
rect 6232 3204 6251 3207
rect 5873 3182 5971 3184
rect 5998 3182 6166 3194
rect 6181 3184 6197 3198
rect 6232 3185 6254 3204
rect 6264 3198 6280 3199
rect 6263 3196 6280 3198
rect 6264 3191 6280 3196
rect 6254 3184 6260 3185
rect 6263 3184 6292 3191
rect 6181 3183 6292 3184
rect 6181 3182 6298 3183
rect 5857 3174 5908 3182
rect 5955 3174 5989 3182
rect 5857 3162 5882 3174
rect 5889 3162 5908 3174
rect 5962 3172 5989 3174
rect 5998 3172 6219 3182
rect 6254 3179 6260 3182
rect 5962 3168 6219 3172
rect 5857 3154 5908 3162
rect 5955 3154 6219 3168
rect 6263 3174 6298 3182
rect 5809 3106 5828 3140
rect 5873 3146 5902 3154
rect 5873 3140 5890 3146
rect 5873 3138 5907 3140
rect 5955 3138 5971 3154
rect 5972 3144 6180 3154
rect 6181 3144 6197 3154
rect 6245 3150 6260 3165
rect 6263 3162 6264 3174
rect 6271 3162 6298 3174
rect 6263 3154 6298 3162
rect 6263 3153 6292 3154
rect 5983 3140 6197 3144
rect 5998 3138 6197 3140
rect 6232 3140 6245 3150
rect 6263 3140 6280 3153
rect 6232 3138 6280 3140
rect 5874 3134 5907 3138
rect 5870 3132 5907 3134
rect 5870 3131 5937 3132
rect 5870 3126 5901 3131
rect 5907 3126 5937 3131
rect 5870 3122 5937 3126
rect 5843 3119 5937 3122
rect 5843 3112 5892 3119
rect 5843 3106 5873 3112
rect 5892 3107 5897 3112
rect 5809 3090 5889 3106
rect 5901 3098 5937 3119
rect 5998 3114 6187 3138
rect 6232 3137 6279 3138
rect 6245 3132 6279 3137
rect 6013 3111 6187 3114
rect 6006 3108 6187 3111
rect 6215 3131 6279 3132
rect 5809 3088 5828 3090
rect 5843 3088 5877 3090
rect 5809 3072 5889 3088
rect 5809 3066 5828 3072
rect 5525 3040 5628 3050
rect 5479 3038 5628 3040
rect 5649 3038 5684 3050
rect 5318 3036 5480 3038
rect 5330 3016 5349 3036
rect 5364 3034 5394 3036
rect 5213 3008 5254 3016
rect 5336 3012 5349 3016
rect 5401 3020 5480 3036
rect 5512 3036 5684 3038
rect 5512 3020 5591 3036
rect 5598 3034 5628 3036
rect 5176 2998 5205 3008
rect 5219 2998 5248 3008
rect 5263 2998 5293 3012
rect 5336 2998 5379 3012
rect 5401 3008 5591 3020
rect 5656 3016 5662 3036
rect 5386 2998 5416 3008
rect 5417 2998 5575 3008
rect 5579 2998 5609 3008
rect 5613 2998 5643 3012
rect 5671 2998 5684 3036
rect 5756 3050 5785 3066
rect 5799 3050 5828 3066
rect 5843 3056 5873 3072
rect 5901 3050 5907 3098
rect 5910 3092 5929 3098
rect 5944 3092 5974 3100
rect 5910 3084 5974 3092
rect 5910 3068 5990 3084
rect 6006 3077 6068 3108
rect 6084 3077 6146 3108
rect 6215 3106 6264 3131
rect 6279 3106 6309 3122
rect 6178 3092 6208 3100
rect 6215 3098 6325 3106
rect 6178 3084 6223 3092
rect 5910 3066 5929 3068
rect 5944 3066 5990 3068
rect 5910 3050 5990 3066
rect 6017 3064 6052 3077
rect 6093 3074 6130 3077
rect 6093 3072 6135 3074
rect 6022 3061 6052 3064
rect 6031 3057 6038 3061
rect 6038 3056 6039 3057
rect 5997 3050 6007 3056
rect 5756 3042 5791 3050
rect 5756 3016 5757 3042
rect 5764 3016 5791 3042
rect 5699 2998 5729 3012
rect 5756 3008 5791 3016
rect 5793 3042 5834 3050
rect 5793 3016 5808 3042
rect 5815 3016 5834 3042
rect 5898 3038 5929 3050
rect 5944 3038 6047 3050
rect 6059 3040 6085 3066
rect 6100 3061 6130 3072
rect 6162 3068 6224 3084
rect 6162 3066 6208 3068
rect 6162 3050 6224 3066
rect 6236 3050 6242 3098
rect 6245 3090 6325 3098
rect 6245 3088 6264 3090
rect 6279 3088 6313 3090
rect 6245 3072 6325 3088
rect 6245 3050 6264 3072
rect 6279 3056 6309 3072
rect 6337 3066 6343 3140
rect 6346 3066 6365 3210
rect 6380 3066 6386 3210
rect 6395 3140 6408 3210
rect 6460 3206 6482 3210
rect 6453 3184 6482 3198
rect 6535 3184 6551 3198
rect 6589 3194 6595 3196
rect 6602 3194 6710 3210
rect 6717 3194 6723 3196
rect 6731 3194 6746 3210
rect 6812 3204 6831 3207
rect 6453 3182 6551 3184
rect 6578 3182 6746 3194
rect 6761 3184 6777 3198
rect 6812 3185 6834 3204
rect 6844 3198 6860 3199
rect 6843 3196 6860 3198
rect 6844 3191 6860 3196
rect 6834 3184 6840 3185
rect 6843 3184 6872 3191
rect 6761 3183 6872 3184
rect 6761 3182 6878 3183
rect 6437 3174 6488 3182
rect 6535 3174 6569 3182
rect 6437 3162 6462 3174
rect 6469 3162 6488 3174
rect 6542 3172 6569 3174
rect 6578 3172 6799 3182
rect 6834 3179 6840 3182
rect 6542 3168 6799 3172
rect 6437 3154 6488 3162
rect 6535 3154 6799 3168
rect 6843 3174 6878 3182
rect 6389 3106 6408 3140
rect 6453 3146 6482 3154
rect 6453 3140 6470 3146
rect 6453 3138 6487 3140
rect 6535 3138 6551 3154
rect 6552 3144 6760 3154
rect 6761 3144 6777 3154
rect 6825 3150 6840 3165
rect 6843 3162 6844 3174
rect 6851 3162 6878 3174
rect 6843 3154 6878 3162
rect 6843 3153 6872 3154
rect 6563 3140 6777 3144
rect 6578 3138 6777 3140
rect 6812 3140 6825 3150
rect 6843 3140 6860 3153
rect 6812 3138 6860 3140
rect 6454 3134 6487 3138
rect 6450 3132 6487 3134
rect 6450 3131 6517 3132
rect 6450 3126 6481 3131
rect 6487 3126 6517 3131
rect 6450 3122 6517 3126
rect 6423 3119 6517 3122
rect 6423 3112 6472 3119
rect 6423 3106 6453 3112
rect 6472 3107 6477 3112
rect 6389 3090 6469 3106
rect 6481 3098 6517 3119
rect 6578 3114 6767 3138
rect 6812 3137 6859 3138
rect 6825 3132 6859 3137
rect 6593 3111 6767 3114
rect 6586 3108 6767 3111
rect 6795 3131 6859 3132
rect 6389 3088 6408 3090
rect 6423 3088 6457 3090
rect 6389 3072 6469 3088
rect 6389 3066 6408 3072
rect 6105 3040 6208 3050
rect 6059 3038 6208 3040
rect 6229 3038 6264 3050
rect 5898 3036 6060 3038
rect 5910 3016 5929 3036
rect 5944 3034 5974 3036
rect 5793 3008 5834 3016
rect 5916 3012 5929 3016
rect 5981 3020 6060 3036
rect 6092 3036 6264 3038
rect 6092 3020 6171 3036
rect 6178 3034 6208 3036
rect 5756 2998 5785 3008
rect 5799 2998 5828 3008
rect 5843 2998 5873 3012
rect 5916 2998 5959 3012
rect 5981 3008 6171 3020
rect 6236 3016 6242 3036
rect 5966 2998 5996 3008
rect 5997 2998 6155 3008
rect 6159 2998 6189 3008
rect 6193 2998 6223 3012
rect 6251 2998 6264 3036
rect 6336 3050 6365 3066
rect 6379 3050 6408 3066
rect 6423 3056 6453 3072
rect 6481 3050 6487 3098
rect 6490 3092 6509 3098
rect 6524 3092 6554 3100
rect 6490 3084 6554 3092
rect 6490 3068 6570 3084
rect 6586 3077 6648 3108
rect 6664 3077 6726 3108
rect 6795 3106 6844 3131
rect 6859 3106 6889 3122
rect 6758 3092 6788 3100
rect 6795 3098 6905 3106
rect 6758 3084 6803 3092
rect 6490 3066 6509 3068
rect 6524 3066 6570 3068
rect 6490 3050 6570 3066
rect 6597 3064 6632 3077
rect 6673 3074 6710 3077
rect 6673 3072 6715 3074
rect 6602 3061 6632 3064
rect 6611 3057 6618 3061
rect 6618 3056 6619 3057
rect 6577 3050 6587 3056
rect 6336 3042 6371 3050
rect 6336 3016 6337 3042
rect 6344 3016 6371 3042
rect 6279 2998 6309 3012
rect 6336 3008 6371 3016
rect 6373 3042 6414 3050
rect 6373 3016 6388 3042
rect 6395 3016 6414 3042
rect 6478 3038 6509 3050
rect 6524 3038 6627 3050
rect 6639 3040 6665 3066
rect 6680 3061 6710 3072
rect 6742 3068 6804 3084
rect 6742 3066 6788 3068
rect 6742 3050 6804 3066
rect 6816 3050 6822 3098
rect 6825 3090 6905 3098
rect 6825 3088 6844 3090
rect 6859 3088 6893 3090
rect 6825 3072 6905 3088
rect 6825 3050 6844 3072
rect 6859 3056 6889 3072
rect 6917 3066 6923 3140
rect 6926 3066 6945 3210
rect 6960 3066 6966 3210
rect 6975 3140 6988 3210
rect 7040 3206 7062 3210
rect 7033 3184 7062 3198
rect 7115 3184 7131 3198
rect 7169 3194 7175 3196
rect 7182 3194 7290 3210
rect 7297 3194 7303 3196
rect 7311 3194 7326 3210
rect 7392 3204 7411 3207
rect 7033 3182 7131 3184
rect 7158 3182 7326 3194
rect 7341 3184 7357 3198
rect 7392 3185 7414 3204
rect 7424 3198 7440 3199
rect 7423 3196 7440 3198
rect 7424 3191 7440 3196
rect 7414 3184 7420 3185
rect 7423 3184 7452 3191
rect 7341 3183 7452 3184
rect 7341 3182 7458 3183
rect 7017 3174 7068 3182
rect 7115 3174 7149 3182
rect 7017 3162 7042 3174
rect 7049 3162 7068 3174
rect 7122 3172 7149 3174
rect 7158 3172 7379 3182
rect 7414 3179 7420 3182
rect 7122 3168 7379 3172
rect 7017 3154 7068 3162
rect 7115 3154 7379 3168
rect 7423 3174 7458 3182
rect 6969 3106 6988 3140
rect 7033 3146 7062 3154
rect 7033 3140 7050 3146
rect 7033 3138 7067 3140
rect 7115 3138 7131 3154
rect 7132 3144 7340 3154
rect 7341 3144 7357 3154
rect 7405 3150 7420 3165
rect 7423 3162 7424 3174
rect 7431 3162 7458 3174
rect 7423 3154 7458 3162
rect 7423 3153 7452 3154
rect 7143 3140 7357 3144
rect 7158 3138 7357 3140
rect 7392 3140 7405 3150
rect 7423 3140 7440 3153
rect 7392 3138 7440 3140
rect 7034 3134 7067 3138
rect 7030 3132 7067 3134
rect 7030 3131 7097 3132
rect 7030 3126 7061 3131
rect 7067 3126 7097 3131
rect 7030 3122 7097 3126
rect 7003 3119 7097 3122
rect 7003 3112 7052 3119
rect 7003 3106 7033 3112
rect 7052 3107 7057 3112
rect 6969 3090 7049 3106
rect 7061 3098 7097 3119
rect 7158 3114 7347 3138
rect 7392 3137 7439 3138
rect 7405 3132 7439 3137
rect 7173 3111 7347 3114
rect 7166 3108 7347 3111
rect 7375 3131 7439 3132
rect 6969 3088 6988 3090
rect 7003 3088 7037 3090
rect 6969 3072 7049 3088
rect 6969 3066 6988 3072
rect 6685 3040 6788 3050
rect 6639 3038 6788 3040
rect 6809 3038 6844 3050
rect 6478 3036 6640 3038
rect 6490 3016 6509 3036
rect 6524 3034 6554 3036
rect 6373 3008 6414 3016
rect 6496 3012 6509 3016
rect 6561 3020 6640 3036
rect 6672 3036 6844 3038
rect 6672 3020 6751 3036
rect 6758 3034 6788 3036
rect 6336 2998 6365 3008
rect 6379 2998 6408 3008
rect 6423 2998 6453 3012
rect 6496 2998 6539 3012
rect 6561 3008 6751 3020
rect 6816 3016 6822 3036
rect 6546 2998 6576 3008
rect 6577 2998 6735 3008
rect 6739 2998 6769 3008
rect 6773 2998 6803 3012
rect 6831 2998 6844 3036
rect 6916 3050 6945 3066
rect 6959 3050 6988 3066
rect 7003 3056 7033 3072
rect 7061 3050 7067 3098
rect 7070 3092 7089 3098
rect 7104 3092 7134 3100
rect 7070 3084 7134 3092
rect 7070 3068 7150 3084
rect 7166 3077 7228 3108
rect 7244 3077 7306 3108
rect 7375 3106 7424 3131
rect 7439 3106 7469 3122
rect 7338 3092 7368 3100
rect 7375 3098 7485 3106
rect 7338 3084 7383 3092
rect 7070 3066 7089 3068
rect 7104 3066 7150 3068
rect 7070 3050 7150 3066
rect 7177 3064 7212 3077
rect 7253 3074 7290 3077
rect 7253 3072 7295 3074
rect 7182 3061 7212 3064
rect 7191 3057 7198 3061
rect 7198 3056 7199 3057
rect 7157 3050 7167 3056
rect 6916 3042 6951 3050
rect 6916 3016 6917 3042
rect 6924 3016 6951 3042
rect 6859 2998 6889 3012
rect 6916 3008 6951 3016
rect 6953 3042 6994 3050
rect 6953 3016 6968 3042
rect 6975 3016 6994 3042
rect 7058 3038 7089 3050
rect 7104 3038 7207 3050
rect 7219 3040 7245 3066
rect 7260 3061 7290 3072
rect 7322 3068 7384 3084
rect 7322 3066 7368 3068
rect 7322 3050 7384 3066
rect 7396 3050 7402 3098
rect 7405 3090 7485 3098
rect 7405 3088 7424 3090
rect 7439 3088 7473 3090
rect 7405 3072 7485 3088
rect 7405 3050 7424 3072
rect 7439 3056 7469 3072
rect 7497 3066 7503 3140
rect 7506 3066 7525 3210
rect 7540 3066 7546 3210
rect 7555 3140 7568 3210
rect 7613 3188 7614 3198
rect 7629 3188 7642 3198
rect 7613 3184 7642 3188
rect 7647 3184 7677 3210
rect 7695 3196 7711 3198
rect 7783 3196 7836 3210
rect 7784 3194 7848 3196
rect 7891 3194 7906 3210
rect 7955 3207 7985 3210
rect 7955 3204 7991 3207
rect 7921 3196 7937 3198
rect 7695 3184 7710 3188
rect 7613 3182 7710 3184
rect 7738 3182 7906 3194
rect 7922 3184 7937 3188
rect 7955 3185 7994 3204
rect 8013 3198 8020 3199
rect 8019 3191 8020 3198
rect 8003 3188 8004 3191
rect 8019 3188 8032 3191
rect 7955 3184 7985 3185
rect 7994 3184 8000 3185
rect 8003 3184 8032 3188
rect 7922 3183 8032 3184
rect 7922 3182 8038 3183
rect 7597 3174 7648 3182
rect 7597 3162 7622 3174
rect 7629 3162 7648 3174
rect 7679 3174 7729 3182
rect 7679 3166 7695 3174
rect 7702 3172 7729 3174
rect 7738 3172 7959 3182
rect 7702 3162 7959 3172
rect 7988 3174 8038 3182
rect 7988 3165 8004 3174
rect 7597 3154 7648 3162
rect 7695 3154 7959 3162
rect 7985 3162 8004 3165
rect 8011 3162 8038 3174
rect 7985 3154 8038 3162
rect 7549 3106 7568 3140
rect 7613 3146 7614 3154
rect 7629 3146 7642 3154
rect 7613 3138 7629 3146
rect 7610 3131 7629 3134
rect 7610 3122 7632 3131
rect 7583 3112 7632 3122
rect 7583 3106 7613 3112
rect 7632 3107 7637 3112
rect 7549 3090 7629 3106
rect 7647 3103 7677 3154
rect 7712 3144 7920 3154
rect 7955 3150 8000 3154
rect 8003 3153 8004 3154
rect 8019 3153 8032 3154
rect 7738 3114 7927 3144
rect 7753 3111 7927 3114
rect 7641 3098 7677 3103
rect 7746 3108 7927 3111
rect 7746 3103 7757 3108
rect 7762 3103 7772 3108
rect 7782 3103 7796 3108
rect 7799 3103 7808 3108
rect 7549 3088 7568 3090
rect 7583 3088 7617 3090
rect 7549 3072 7629 3088
rect 7549 3066 7568 3072
rect 7265 3040 7368 3050
rect 7219 3038 7368 3040
rect 7389 3038 7424 3050
rect 7058 3036 7220 3038
rect 7070 3016 7089 3036
rect 7104 3034 7134 3036
rect 6953 3008 6994 3016
rect 7076 3012 7089 3016
rect 7141 3020 7220 3036
rect 7252 3036 7424 3038
rect 7252 3020 7331 3036
rect 7338 3034 7368 3036
rect 6916 2998 6945 3008
rect 6959 2998 6988 3008
rect 7003 2998 7033 3012
rect 7076 2998 7119 3012
rect 7141 3008 7331 3020
rect 7396 3016 7402 3036
rect 7126 2998 7156 3008
rect 7157 2998 7315 3008
rect 7319 2998 7349 3008
rect 7353 2998 7383 3012
rect 7411 2998 7424 3036
rect 7496 3050 7525 3066
rect 7539 3050 7568 3066
rect 7583 3056 7613 3072
rect 7641 3050 7647 3098
rect 7650 3092 7669 3098
rect 7684 3092 7714 3100
rect 7650 3084 7714 3092
rect 7650 3068 7730 3084
rect 7746 3077 7808 3103
rect 7824 3103 7833 3108
rect 7840 3103 7850 3108
rect 7860 3103 7874 3108
rect 7875 3103 7886 3108
rect 7824 3077 7886 3103
rect 7955 3103 7985 3150
rect 8019 3146 8020 3153
rect 8004 3138 8020 3146
rect 7991 3106 8004 3125
rect 8019 3106 8049 3122
rect 7991 3103 8065 3106
rect 8092 3103 8105 3210
rect 8135 3106 8148 3210
rect 8193 3188 8194 3198
rect 8209 3188 8222 3198
rect 8193 3184 8222 3188
rect 8227 3184 8257 3210
rect 8275 3196 8291 3198
rect 8363 3196 8416 3210
rect 8364 3194 8428 3196
rect 8471 3194 8486 3210
rect 8535 3207 8565 3210
rect 8535 3204 8571 3207
rect 8501 3196 8517 3198
rect 8275 3184 8290 3188
rect 8193 3182 8290 3184
rect 8318 3182 8486 3194
rect 8502 3184 8517 3188
rect 8535 3185 8574 3204
rect 8593 3198 8600 3199
rect 8599 3191 8600 3198
rect 8583 3188 8584 3191
rect 8599 3188 8612 3191
rect 8535 3184 8565 3185
rect 8574 3184 8580 3185
rect 8583 3184 8612 3188
rect 8502 3183 8612 3184
rect 8502 3182 8618 3183
rect 8177 3174 8228 3182
rect 8177 3162 8202 3174
rect 8209 3162 8228 3174
rect 8259 3174 8309 3182
rect 8259 3166 8275 3174
rect 8282 3172 8309 3174
rect 8318 3172 8539 3182
rect 8282 3162 8539 3172
rect 8568 3174 8618 3182
rect 8568 3165 8584 3174
rect 8177 3154 8228 3162
rect 8275 3154 8539 3162
rect 8565 3162 8584 3165
rect 8591 3162 8618 3174
rect 8565 3154 8618 3162
rect 8193 3146 8194 3154
rect 8209 3146 8222 3154
rect 8193 3138 8209 3146
rect 8190 3131 8209 3134
rect 8190 3122 8212 3131
rect 8163 3112 8212 3122
rect 8163 3106 8193 3112
rect 8212 3107 8217 3112
rect 8135 3103 8209 3106
rect 8227 3103 8257 3154
rect 8292 3144 8500 3154
rect 8535 3150 8580 3154
rect 8583 3153 8584 3154
rect 8599 3153 8612 3154
rect 8318 3114 8507 3144
rect 8333 3111 8507 3114
rect 7918 3092 7948 3100
rect 7955 3098 8065 3103
rect 7918 3084 7963 3092
rect 7650 3066 7669 3068
rect 7684 3066 7730 3068
rect 7650 3050 7730 3066
rect 7757 3064 7792 3077
rect 7833 3074 7870 3077
rect 7833 3072 7875 3074
rect 7762 3061 7792 3064
rect 7771 3057 7778 3061
rect 7778 3056 7779 3057
rect 7737 3050 7747 3056
rect 7496 3042 7531 3050
rect 7496 3016 7497 3042
rect 7504 3016 7531 3042
rect 7439 2998 7469 3012
rect 7496 3008 7531 3016
rect 7533 3042 7574 3050
rect 7533 3016 7548 3042
rect 7555 3016 7574 3042
rect 7638 3038 7669 3050
rect 7684 3038 7787 3050
rect 7799 3040 7825 3066
rect 7840 3061 7870 3072
rect 7902 3068 7964 3084
rect 7902 3066 7948 3068
rect 7902 3050 7964 3066
rect 7976 3050 7982 3098
rect 7985 3090 8065 3098
rect 7985 3088 8004 3090
rect 8019 3088 8053 3090
rect 7985 3072 8065 3088
rect 7985 3050 8004 3072
rect 8019 3056 8049 3072
rect 8077 3066 8083 3103
rect 8086 3066 8105 3103
rect 8120 3066 8126 3103
rect 8129 3090 8209 3103
rect 8221 3098 8257 3103
rect 8326 3108 8507 3111
rect 8326 3103 8337 3108
rect 8342 3103 8352 3108
rect 8362 3103 8376 3108
rect 8379 3103 8388 3108
rect 8129 3088 8148 3090
rect 8163 3088 8197 3090
rect 8129 3072 8209 3088
rect 8129 3066 8148 3072
rect 7845 3040 7948 3050
rect 7799 3038 7948 3040
rect 7969 3038 8004 3050
rect 7638 3036 7800 3038
rect 7650 3016 7669 3036
rect 7684 3034 7714 3036
rect 7533 3008 7574 3016
rect 7656 3012 7669 3016
rect 7721 3020 7800 3036
rect 7832 3036 8004 3038
rect 7832 3020 7911 3036
rect 7918 3034 7948 3036
rect 7496 2998 7525 3008
rect 7539 2998 7568 3008
rect 7583 2998 7613 3012
rect 7656 2998 7699 3012
rect 7721 3008 7911 3020
rect 7976 3016 7982 3036
rect 7706 2998 7736 3008
rect 7737 2998 7895 3008
rect 7899 2998 7929 3008
rect 7933 2998 7963 3012
rect 7991 2998 8004 3036
rect 8076 3050 8105 3066
rect 8119 3050 8148 3066
rect 8163 3056 8193 3072
rect 8221 3050 8227 3098
rect 8230 3092 8249 3098
rect 8264 3092 8294 3100
rect 8230 3084 8294 3092
rect 8230 3068 8310 3084
rect 8326 3077 8388 3103
rect 8404 3103 8413 3108
rect 8420 3103 8430 3108
rect 8440 3103 8454 3108
rect 8455 3103 8466 3108
rect 8404 3077 8466 3103
rect 8535 3103 8565 3150
rect 8599 3146 8600 3153
rect 8584 3138 8600 3146
rect 8571 3106 8584 3125
rect 8599 3106 8629 3122
rect 8571 3103 8645 3106
rect 8672 3103 8685 3210
rect 8715 3106 8728 3210
rect 8773 3188 8774 3198
rect 8789 3188 8802 3198
rect 8773 3184 8802 3188
rect 8807 3184 8837 3210
rect 8855 3196 8871 3198
rect 8943 3196 8996 3210
rect 8944 3194 9008 3196
rect 9051 3194 9066 3210
rect 9115 3207 9145 3210
rect 9115 3204 9151 3207
rect 9081 3196 9097 3198
rect 8855 3184 8870 3188
rect 8773 3182 8870 3184
rect 8898 3182 9066 3194
rect 9082 3184 9097 3188
rect 9115 3185 9154 3204
rect 9173 3198 9180 3199
rect 9179 3191 9180 3198
rect 9163 3188 9164 3191
rect 9179 3188 9192 3191
rect 9115 3184 9145 3185
rect 9154 3184 9160 3185
rect 9163 3184 9192 3188
rect 9082 3183 9192 3184
rect 9082 3182 9198 3183
rect 8757 3174 8808 3182
rect 8757 3162 8782 3174
rect 8789 3162 8808 3174
rect 8839 3174 8889 3182
rect 8839 3166 8855 3174
rect 8862 3172 8889 3174
rect 8898 3172 9119 3182
rect 8862 3162 9119 3172
rect 9148 3174 9198 3182
rect 9148 3165 9164 3174
rect 8757 3154 8808 3162
rect 8855 3154 9119 3162
rect 9145 3162 9164 3165
rect 9171 3162 9198 3174
rect 9145 3154 9198 3162
rect 8773 3146 8774 3154
rect 8789 3146 8802 3154
rect 8773 3138 8789 3146
rect 8770 3131 8789 3134
rect 8770 3122 8792 3131
rect 8743 3112 8792 3122
rect 8743 3106 8773 3112
rect 8792 3107 8797 3112
rect 8715 3103 8789 3106
rect 8807 3103 8837 3154
rect 8872 3144 9080 3154
rect 9115 3150 9160 3154
rect 9163 3153 9164 3154
rect 9179 3153 9192 3154
rect 8898 3114 9087 3144
rect 8913 3111 9087 3114
rect 8498 3092 8528 3100
rect 8535 3098 8645 3103
rect 8498 3084 8543 3092
rect 8230 3066 8249 3068
rect 8264 3066 8310 3068
rect 8230 3050 8310 3066
rect 8337 3064 8372 3077
rect 8413 3074 8450 3077
rect 8413 3072 8455 3074
rect 8342 3061 8372 3064
rect 8351 3057 8358 3061
rect 8358 3056 8359 3057
rect 8317 3050 8327 3056
rect 8076 3042 8111 3050
rect 8076 3016 8077 3042
rect 8084 3016 8111 3042
rect 8019 2998 8049 3012
rect 8076 3008 8111 3016
rect 8113 3042 8154 3050
rect 8113 3016 8128 3042
rect 8135 3016 8154 3042
rect 8218 3038 8249 3050
rect 8264 3038 8367 3050
rect 8379 3040 8405 3066
rect 8420 3061 8450 3072
rect 8482 3068 8544 3084
rect 8482 3066 8528 3068
rect 8482 3050 8544 3066
rect 8556 3050 8562 3098
rect 8565 3090 8645 3098
rect 8565 3088 8584 3090
rect 8599 3088 8633 3090
rect 8565 3072 8645 3088
rect 8565 3050 8584 3072
rect 8599 3056 8629 3072
rect 8657 3066 8663 3103
rect 8666 3066 8685 3103
rect 8700 3066 8706 3103
rect 8709 3090 8789 3103
rect 8801 3098 8837 3103
rect 8906 3108 9087 3111
rect 8906 3103 8917 3108
rect 8922 3103 8932 3108
rect 8942 3103 8956 3108
rect 8959 3103 8968 3108
rect 8709 3088 8728 3090
rect 8743 3088 8777 3090
rect 8709 3072 8789 3088
rect 8709 3066 8728 3072
rect 8425 3040 8528 3050
rect 8379 3038 8528 3040
rect 8549 3038 8584 3050
rect 8218 3036 8380 3038
rect 8230 3016 8249 3036
rect 8264 3034 8294 3036
rect 8113 3008 8154 3016
rect 8236 3012 8249 3016
rect 8301 3020 8380 3036
rect 8412 3036 8584 3038
rect 8412 3020 8491 3036
rect 8498 3034 8528 3036
rect 8076 2998 8105 3008
rect 8119 2998 8148 3008
rect 8163 2998 8193 3012
rect 8236 2998 8279 3012
rect 8301 3008 8491 3020
rect 8556 3016 8562 3036
rect 8286 2998 8316 3008
rect 8317 2998 8475 3008
rect 8479 2998 8509 3008
rect 8513 2998 8543 3012
rect 8571 2998 8584 3036
rect 8656 3050 8685 3066
rect 8699 3050 8728 3066
rect 8743 3056 8773 3072
rect 8801 3050 8807 3098
rect 8810 3092 8829 3098
rect 8844 3092 8874 3100
rect 8810 3084 8874 3092
rect 8810 3068 8890 3084
rect 8906 3077 8968 3103
rect 8984 3103 8993 3108
rect 9000 3103 9010 3108
rect 9020 3103 9034 3108
rect 9035 3103 9046 3108
rect 8984 3077 9046 3103
rect 9115 3103 9145 3150
rect 9179 3146 9180 3153
rect 9164 3138 9180 3146
rect 9151 3106 9164 3125
rect 9179 3106 9209 3122
rect 9151 3103 9225 3106
rect 9078 3092 9108 3100
rect 9115 3098 9225 3103
rect 9078 3084 9123 3092
rect 8810 3066 8829 3068
rect 8844 3066 8890 3068
rect 8810 3050 8890 3066
rect 8917 3064 8952 3077
rect 8993 3074 9030 3077
rect 8993 3072 9035 3074
rect 8922 3061 8952 3064
rect 8931 3057 8938 3061
rect 8938 3056 8939 3057
rect 8897 3050 8907 3056
rect 8656 3042 8691 3050
rect 8656 3016 8657 3042
rect 8664 3016 8691 3042
rect 8599 2998 8629 3012
rect 8656 3008 8691 3016
rect 8693 3042 8734 3050
rect 8693 3016 8708 3042
rect 8715 3016 8734 3042
rect 8798 3038 8829 3050
rect 8844 3038 8947 3050
rect 8959 3040 8985 3066
rect 9000 3061 9030 3072
rect 9062 3068 9124 3084
rect 9062 3066 9108 3068
rect 9062 3050 9124 3066
rect 9136 3050 9142 3098
rect 9145 3090 9225 3098
rect 9145 3088 9164 3090
rect 9179 3088 9213 3090
rect 9145 3072 9225 3088
rect 9145 3050 9164 3072
rect 9179 3056 9209 3072
rect 9237 3066 9243 3103
rect 9252 3066 9265 3210
rect 9005 3040 9108 3050
rect 8959 3038 9108 3040
rect 9129 3038 9164 3050
rect 8798 3036 8960 3038
rect 8810 3016 8829 3036
rect 8844 3034 8874 3036
rect 8693 3008 8734 3016
rect 8816 3012 8829 3016
rect 8881 3020 8960 3036
rect 8992 3036 9164 3038
rect 8992 3020 9071 3036
rect 9078 3034 9108 3036
rect 8656 2998 8685 3008
rect 8699 2998 8728 3008
rect 8743 2998 8773 3012
rect 8816 2998 8859 3012
rect 8881 3008 9071 3020
rect 9136 3016 9142 3036
rect 8866 2998 8896 3008
rect 8897 2998 9055 3008
rect 9059 2998 9089 3008
rect 9093 2998 9123 3012
rect 9151 2998 9164 3036
rect 9236 3050 9265 3066
rect 9236 3042 9271 3050
rect 9236 3016 9237 3042
rect 9244 3016 9271 3042
rect 9179 2998 9209 3012
rect 9236 3008 9271 3016
rect 9236 2998 9265 3008
rect -1 2992 9265 2998
rect 0 2984 9265 2992
rect 15 2954 28 2984
rect 43 2970 73 2984
rect 116 2970 159 2984
rect 166 2970 386 2984
rect 393 2970 423 2984
rect 83 2956 98 2968
rect 117 2956 130 2970
rect 198 2966 351 2970
rect 80 2954 102 2956
rect 180 2954 372 2966
rect 451 2954 464 2984
rect 479 2970 509 2984
rect 546 2954 565 2984
rect 580 2954 586 2984
rect 595 2954 608 2984
rect 623 2970 653 2984
rect 696 2970 739 2984
rect 746 2970 966 2984
rect 973 2970 1003 2984
rect 663 2956 678 2968
rect 697 2956 710 2970
rect 778 2966 931 2970
rect 660 2954 682 2956
rect 760 2954 952 2966
rect 1031 2954 1044 2984
rect 1059 2970 1089 2984
rect 1126 2954 1145 2984
rect 1160 2954 1166 2984
rect 1175 2954 1188 2984
rect 1203 2970 1233 2984
rect 1276 2970 1319 2984
rect 1326 2970 1546 2984
rect 1553 2970 1583 2984
rect 1243 2956 1258 2968
rect 1277 2956 1290 2970
rect 1358 2966 1511 2970
rect 1240 2954 1262 2956
rect 1340 2954 1532 2966
rect 1611 2954 1624 2984
rect 1639 2970 1669 2984
rect 1706 2954 1725 2984
rect 1740 2954 1746 2984
rect 1755 2954 1768 2984
rect 1783 2970 1813 2984
rect 1856 2970 1899 2984
rect 1906 2970 2126 2984
rect 2133 2970 2163 2984
rect 1823 2956 1838 2968
rect 1857 2956 1870 2970
rect 1938 2966 2091 2970
rect 1820 2954 1842 2956
rect 1920 2954 2112 2966
rect 2191 2954 2204 2984
rect 2219 2970 2249 2984
rect 2286 2954 2305 2984
rect 2320 2954 2326 2984
rect 2335 2954 2348 2984
rect 2363 2970 2393 2984
rect 2436 2970 2479 2984
rect 2486 2970 2706 2984
rect 2713 2970 2743 2984
rect 2403 2956 2418 2968
rect 2437 2956 2450 2970
rect 2518 2966 2671 2970
rect 2400 2954 2422 2956
rect 2500 2954 2692 2966
rect 2771 2954 2784 2984
rect 2799 2970 2829 2984
rect 2866 2954 2885 2984
rect 2900 2954 2906 2984
rect 2915 2954 2928 2984
rect 2943 2970 2973 2984
rect 3016 2970 3059 2984
rect 3066 2970 3286 2984
rect 3293 2970 3323 2984
rect 2983 2956 2998 2968
rect 3017 2956 3030 2970
rect 3098 2966 3251 2970
rect 2980 2954 3002 2956
rect 3080 2954 3272 2966
rect 3351 2954 3364 2984
rect 3379 2970 3409 2984
rect 3446 2954 3465 2984
rect 3480 2954 3486 2984
rect 3495 2954 3508 2984
rect 3523 2970 3553 2984
rect 3596 2970 3639 2984
rect 3646 2970 3866 2984
rect 3873 2970 3903 2984
rect 3563 2956 3578 2968
rect 3597 2956 3610 2970
rect 3678 2966 3831 2970
rect 3560 2954 3582 2956
rect 3660 2954 3852 2966
rect 3931 2954 3944 2984
rect 3959 2970 3989 2984
rect 4026 2954 4045 2984
rect 4060 2954 4066 2984
rect 4075 2954 4088 2984
rect 4103 2970 4133 2984
rect 4176 2970 4219 2984
rect 4226 2970 4446 2984
rect 4453 2970 4483 2984
rect 4143 2956 4158 2968
rect 4177 2956 4190 2970
rect 4258 2966 4411 2970
rect 4140 2954 4162 2956
rect 4240 2954 4432 2966
rect 4511 2954 4524 2984
rect 4539 2970 4569 2984
rect 4606 2954 4625 2984
rect 4640 2954 4646 2984
rect 4655 2954 4668 2984
rect 4683 2970 4713 2984
rect 4756 2970 4799 2984
rect 4806 2970 5026 2984
rect 5033 2970 5063 2984
rect 4723 2956 4738 2968
rect 4757 2956 4770 2970
rect 4838 2966 4991 2970
rect 4720 2954 4742 2956
rect 4820 2954 5012 2966
rect 5091 2954 5104 2984
rect 5119 2970 5149 2984
rect 5186 2954 5205 2984
rect 5220 2954 5226 2984
rect 5235 2954 5248 2984
rect 5263 2970 5293 2984
rect 5336 2970 5379 2984
rect 5386 2970 5606 2984
rect 5613 2970 5643 2984
rect 5303 2956 5318 2968
rect 5337 2956 5350 2970
rect 5418 2966 5571 2970
rect 5300 2954 5322 2956
rect 5400 2954 5592 2966
rect 5671 2954 5684 2984
rect 5699 2970 5729 2984
rect 5766 2954 5785 2984
rect 5800 2954 5806 2984
rect 5815 2954 5828 2984
rect 5843 2970 5873 2984
rect 5916 2970 5959 2984
rect 5966 2970 6186 2984
rect 6193 2970 6223 2984
rect 5883 2956 5898 2968
rect 5917 2956 5930 2970
rect 5998 2966 6151 2970
rect 5880 2954 5902 2956
rect 5980 2954 6172 2966
rect 6251 2954 6264 2984
rect 6279 2970 6309 2984
rect 6346 2954 6365 2984
rect 6380 2954 6386 2984
rect 6395 2954 6408 2984
rect 6423 2970 6453 2984
rect 6496 2970 6539 2984
rect 6546 2970 6766 2984
rect 6773 2970 6803 2984
rect 6463 2956 6478 2968
rect 6497 2956 6510 2970
rect 6578 2966 6731 2970
rect 6460 2954 6482 2956
rect 6560 2954 6752 2966
rect 6831 2954 6844 2984
rect 6859 2970 6889 2984
rect 6926 2954 6945 2984
rect 6960 2954 6966 2984
rect 6975 2954 6988 2984
rect 7003 2970 7033 2984
rect 7076 2970 7119 2984
rect 7126 2970 7346 2984
rect 7353 2970 7383 2984
rect 7043 2956 7058 2968
rect 7077 2956 7090 2970
rect 7158 2966 7311 2970
rect 7040 2954 7062 2956
rect 7140 2954 7332 2966
rect 7411 2954 7424 2984
rect 7439 2970 7469 2984
rect 7506 2954 7525 2984
rect 7540 2954 7546 2984
rect 7555 2954 7568 2984
rect 7583 2970 7613 2984
rect 7656 2970 7699 2984
rect 7706 2970 7926 2984
rect 7933 2970 7963 2984
rect 7623 2956 7638 2968
rect 7657 2956 7670 2970
rect 7738 2966 7891 2970
rect 7620 2954 7642 2956
rect 7720 2954 7912 2966
rect 7991 2954 8004 2984
rect 8019 2970 8049 2984
rect 8086 2954 8105 2984
rect 8120 2954 8126 2984
rect 8135 2954 8148 2984
rect 8163 2970 8193 2984
rect 8236 2970 8279 2984
rect 8286 2970 8506 2984
rect 8513 2970 8543 2984
rect 8203 2956 8218 2968
rect 8237 2956 8250 2970
rect 8318 2966 8471 2970
rect 8200 2954 8222 2956
rect 8300 2954 8492 2966
rect 8571 2954 8584 2984
rect 8599 2970 8629 2984
rect 8666 2954 8685 2984
rect 8700 2954 8706 2984
rect 8715 2954 8728 2984
rect 8743 2970 8773 2984
rect 8816 2970 8859 2984
rect 8866 2970 9086 2984
rect 9093 2970 9123 2984
rect 8783 2956 8798 2968
rect 8817 2956 8830 2970
rect 8898 2966 9051 2970
rect 8780 2954 8802 2956
rect 8880 2954 9072 2966
rect 9151 2954 9164 2984
rect 9179 2970 9209 2984
rect 9252 2954 9265 2984
rect 0 2940 9265 2954
rect 15 2870 28 2940
rect 80 2936 102 2940
rect 73 2914 102 2928
rect 155 2914 171 2928
rect 209 2924 215 2926
rect 222 2924 330 2940
rect 337 2924 343 2926
rect 351 2924 366 2940
rect 432 2934 451 2937
rect 73 2912 171 2914
rect 198 2912 366 2924
rect 381 2914 397 2928
rect 432 2915 454 2934
rect 464 2928 480 2929
rect 463 2926 480 2928
rect 464 2921 480 2926
rect 454 2914 460 2915
rect 463 2914 492 2921
rect 381 2913 492 2914
rect 381 2912 498 2913
rect 57 2904 108 2912
rect 155 2904 189 2912
rect 57 2892 82 2904
rect 89 2892 108 2904
rect 162 2902 189 2904
rect 198 2902 419 2912
rect 454 2909 460 2912
rect 162 2898 419 2902
rect 57 2884 108 2892
rect 155 2884 419 2898
rect 463 2904 498 2912
rect 9 2836 28 2870
rect 73 2876 102 2884
rect 73 2870 90 2876
rect 73 2868 107 2870
rect 155 2868 171 2884
rect 172 2874 380 2884
rect 381 2874 397 2884
rect 445 2880 460 2895
rect 463 2892 464 2904
rect 471 2892 498 2904
rect 463 2884 498 2892
rect 463 2883 492 2884
rect 183 2870 397 2874
rect 198 2868 397 2870
rect 432 2870 445 2880
rect 463 2870 480 2883
rect 432 2868 480 2870
rect 74 2864 107 2868
rect 70 2862 107 2864
rect 70 2861 137 2862
rect 70 2856 101 2861
rect 107 2856 137 2861
rect 70 2852 137 2856
rect 43 2849 137 2852
rect 43 2842 92 2849
rect 43 2836 73 2842
rect 92 2837 97 2842
rect 9 2820 89 2836
rect 101 2828 137 2849
rect 198 2844 387 2868
rect 432 2867 479 2868
rect 445 2862 479 2867
rect 213 2841 387 2844
rect 206 2838 387 2841
rect 415 2861 479 2862
rect 9 2818 28 2820
rect 43 2818 77 2820
rect 9 2802 89 2818
rect 9 2796 28 2802
rect -1 2780 28 2796
rect 43 2786 73 2802
rect 101 2780 107 2828
rect 110 2822 129 2828
rect 144 2822 174 2830
rect 110 2814 174 2822
rect 110 2798 190 2814
rect 206 2807 268 2838
rect 284 2807 346 2838
rect 415 2836 464 2861
rect 479 2836 509 2852
rect 378 2822 408 2830
rect 415 2828 525 2836
rect 378 2814 423 2822
rect 110 2796 129 2798
rect 144 2796 190 2798
rect 110 2780 190 2796
rect 217 2794 252 2807
rect 293 2804 330 2807
rect 293 2802 335 2804
rect 222 2791 252 2794
rect 231 2787 238 2791
rect 238 2786 239 2787
rect 197 2780 207 2786
rect -7 2772 34 2780
rect -7 2746 8 2772
rect 15 2746 34 2772
rect 98 2768 129 2780
rect 144 2768 247 2780
rect 259 2770 285 2796
rect 300 2791 330 2802
rect 362 2798 424 2814
rect 362 2796 408 2798
rect 362 2780 424 2796
rect 436 2780 442 2828
rect 445 2820 525 2828
rect 445 2818 464 2820
rect 479 2818 513 2820
rect 445 2802 525 2818
rect 445 2780 464 2802
rect 479 2786 509 2802
rect 537 2796 543 2870
rect 546 2796 565 2940
rect 580 2796 586 2940
rect 595 2870 608 2940
rect 660 2936 682 2940
rect 653 2914 682 2928
rect 735 2914 751 2928
rect 789 2924 795 2926
rect 802 2924 910 2940
rect 917 2924 923 2926
rect 931 2924 946 2940
rect 1012 2934 1031 2937
rect 653 2912 751 2914
rect 778 2912 946 2924
rect 961 2914 977 2928
rect 1012 2915 1034 2934
rect 1044 2928 1060 2929
rect 1043 2926 1060 2928
rect 1044 2921 1060 2926
rect 1034 2914 1040 2915
rect 1043 2914 1072 2921
rect 961 2913 1072 2914
rect 961 2912 1078 2913
rect 637 2904 688 2912
rect 735 2904 769 2912
rect 637 2892 662 2904
rect 669 2892 688 2904
rect 742 2902 769 2904
rect 778 2902 999 2912
rect 1034 2909 1040 2912
rect 742 2898 999 2902
rect 637 2884 688 2892
rect 735 2884 999 2898
rect 1043 2904 1078 2912
rect 589 2836 608 2870
rect 653 2876 682 2884
rect 653 2870 670 2876
rect 653 2868 687 2870
rect 735 2868 751 2884
rect 752 2874 960 2884
rect 961 2874 977 2884
rect 1025 2880 1040 2895
rect 1043 2892 1044 2904
rect 1051 2892 1078 2904
rect 1043 2884 1078 2892
rect 1043 2883 1072 2884
rect 763 2870 977 2874
rect 778 2868 977 2870
rect 1012 2870 1025 2880
rect 1043 2870 1060 2883
rect 1012 2868 1060 2870
rect 654 2864 687 2868
rect 650 2862 687 2864
rect 650 2861 717 2862
rect 650 2856 681 2861
rect 687 2856 717 2861
rect 650 2852 717 2856
rect 623 2849 717 2852
rect 623 2842 672 2849
rect 623 2836 653 2842
rect 672 2837 677 2842
rect 589 2820 669 2836
rect 681 2828 717 2849
rect 778 2844 967 2868
rect 1012 2867 1059 2868
rect 1025 2862 1059 2867
rect 793 2841 967 2844
rect 786 2838 967 2841
rect 995 2861 1059 2862
rect 589 2818 608 2820
rect 623 2818 657 2820
rect 589 2802 669 2818
rect 589 2796 608 2802
rect 305 2770 408 2780
rect 259 2768 408 2770
rect 429 2768 464 2780
rect 98 2766 260 2768
rect 110 2746 129 2766
rect 144 2764 174 2766
rect -7 2738 34 2746
rect 116 2742 129 2746
rect 181 2750 260 2766
rect 292 2766 464 2768
rect 292 2750 371 2766
rect 378 2764 408 2766
rect -1 2728 28 2738
rect 43 2728 73 2742
rect 116 2728 159 2742
rect 181 2738 371 2750
rect 436 2746 442 2766
rect 166 2728 196 2738
rect 197 2728 355 2738
rect 359 2728 389 2738
rect 393 2728 423 2742
rect 451 2728 464 2766
rect 536 2780 565 2796
rect 579 2780 608 2796
rect 623 2786 653 2802
rect 681 2780 687 2828
rect 690 2822 709 2828
rect 724 2822 754 2830
rect 690 2814 754 2822
rect 690 2798 770 2814
rect 786 2807 848 2838
rect 864 2807 926 2838
rect 995 2836 1044 2861
rect 1059 2836 1089 2852
rect 958 2822 988 2830
rect 995 2828 1105 2836
rect 958 2814 1003 2822
rect 690 2796 709 2798
rect 724 2796 770 2798
rect 690 2780 770 2796
rect 797 2794 832 2807
rect 873 2804 910 2807
rect 873 2802 915 2804
rect 802 2791 832 2794
rect 811 2787 818 2791
rect 818 2786 819 2787
rect 777 2780 787 2786
rect 536 2772 571 2780
rect 536 2746 537 2772
rect 544 2746 571 2772
rect 479 2728 509 2742
rect 536 2738 571 2746
rect 573 2772 614 2780
rect 573 2746 588 2772
rect 595 2746 614 2772
rect 678 2768 709 2780
rect 724 2768 827 2780
rect 839 2770 865 2796
rect 880 2791 910 2802
rect 942 2798 1004 2814
rect 942 2796 988 2798
rect 942 2780 1004 2796
rect 1016 2780 1022 2828
rect 1025 2820 1105 2828
rect 1025 2818 1044 2820
rect 1059 2818 1093 2820
rect 1025 2802 1105 2818
rect 1025 2780 1044 2802
rect 1059 2786 1089 2802
rect 1117 2796 1123 2870
rect 1126 2796 1145 2940
rect 1160 2796 1166 2940
rect 1175 2870 1188 2940
rect 1240 2936 1262 2940
rect 1233 2914 1262 2928
rect 1315 2914 1331 2928
rect 1369 2924 1375 2926
rect 1382 2924 1490 2940
rect 1497 2924 1503 2926
rect 1511 2924 1526 2940
rect 1592 2934 1611 2937
rect 1233 2912 1331 2914
rect 1358 2912 1526 2924
rect 1541 2914 1557 2928
rect 1592 2915 1614 2934
rect 1624 2928 1640 2929
rect 1623 2926 1640 2928
rect 1624 2921 1640 2926
rect 1614 2914 1620 2915
rect 1623 2914 1652 2921
rect 1541 2913 1652 2914
rect 1541 2912 1658 2913
rect 1217 2904 1268 2912
rect 1315 2904 1349 2912
rect 1217 2892 1242 2904
rect 1249 2892 1268 2904
rect 1322 2902 1349 2904
rect 1358 2902 1579 2912
rect 1614 2909 1620 2912
rect 1322 2898 1579 2902
rect 1217 2884 1268 2892
rect 1315 2884 1579 2898
rect 1623 2904 1658 2912
rect 1169 2836 1188 2870
rect 1233 2876 1262 2884
rect 1233 2870 1250 2876
rect 1233 2868 1267 2870
rect 1315 2868 1331 2884
rect 1332 2874 1540 2884
rect 1541 2874 1557 2884
rect 1605 2880 1620 2895
rect 1623 2892 1624 2904
rect 1631 2892 1658 2904
rect 1623 2884 1658 2892
rect 1623 2883 1652 2884
rect 1343 2870 1557 2874
rect 1358 2868 1557 2870
rect 1592 2870 1605 2880
rect 1623 2870 1640 2883
rect 1592 2868 1640 2870
rect 1234 2864 1267 2868
rect 1230 2862 1267 2864
rect 1230 2861 1297 2862
rect 1230 2856 1261 2861
rect 1267 2856 1297 2861
rect 1230 2852 1297 2856
rect 1203 2849 1297 2852
rect 1203 2842 1252 2849
rect 1203 2836 1233 2842
rect 1252 2837 1257 2842
rect 1169 2820 1249 2836
rect 1261 2828 1297 2849
rect 1358 2844 1547 2868
rect 1592 2867 1639 2868
rect 1605 2862 1639 2867
rect 1373 2841 1547 2844
rect 1366 2838 1547 2841
rect 1575 2861 1639 2862
rect 1169 2818 1188 2820
rect 1203 2818 1237 2820
rect 1169 2802 1249 2818
rect 1169 2796 1188 2802
rect 885 2770 988 2780
rect 839 2768 988 2770
rect 1009 2768 1044 2780
rect 678 2766 840 2768
rect 690 2746 709 2766
rect 724 2764 754 2766
rect 573 2738 614 2746
rect 696 2742 709 2746
rect 761 2750 840 2766
rect 872 2766 1044 2768
rect 872 2750 951 2766
rect 958 2764 988 2766
rect 536 2728 565 2738
rect 579 2728 608 2738
rect 623 2728 653 2742
rect 696 2728 739 2742
rect 761 2738 951 2750
rect 1016 2746 1022 2766
rect 746 2728 776 2738
rect 777 2728 935 2738
rect 939 2728 969 2738
rect 973 2728 1003 2742
rect 1031 2728 1044 2766
rect 1116 2780 1145 2796
rect 1159 2780 1188 2796
rect 1203 2786 1233 2802
rect 1261 2780 1267 2828
rect 1270 2822 1289 2828
rect 1304 2822 1334 2830
rect 1270 2814 1334 2822
rect 1270 2798 1350 2814
rect 1366 2807 1428 2838
rect 1444 2807 1506 2838
rect 1575 2836 1624 2861
rect 1639 2836 1669 2852
rect 1538 2822 1568 2830
rect 1575 2828 1685 2836
rect 1538 2814 1583 2822
rect 1270 2796 1289 2798
rect 1304 2796 1350 2798
rect 1270 2780 1350 2796
rect 1377 2794 1412 2807
rect 1453 2804 1490 2807
rect 1453 2802 1495 2804
rect 1382 2791 1412 2794
rect 1391 2787 1398 2791
rect 1398 2786 1399 2787
rect 1357 2780 1367 2786
rect 1116 2772 1151 2780
rect 1116 2746 1117 2772
rect 1124 2746 1151 2772
rect 1059 2728 1089 2742
rect 1116 2738 1151 2746
rect 1153 2772 1194 2780
rect 1153 2746 1168 2772
rect 1175 2746 1194 2772
rect 1258 2768 1289 2780
rect 1304 2768 1407 2780
rect 1419 2770 1445 2796
rect 1460 2791 1490 2802
rect 1522 2798 1584 2814
rect 1522 2796 1568 2798
rect 1522 2780 1584 2796
rect 1596 2780 1602 2828
rect 1605 2820 1685 2828
rect 1605 2818 1624 2820
rect 1639 2818 1673 2820
rect 1605 2802 1685 2818
rect 1605 2780 1624 2802
rect 1639 2786 1669 2802
rect 1697 2796 1703 2870
rect 1706 2796 1725 2940
rect 1740 2796 1746 2940
rect 1755 2870 1768 2940
rect 1820 2936 1842 2940
rect 1813 2914 1842 2928
rect 1895 2914 1911 2928
rect 1949 2924 1955 2926
rect 1962 2924 2070 2940
rect 2077 2924 2083 2926
rect 2091 2924 2106 2940
rect 2172 2934 2191 2937
rect 1813 2912 1911 2914
rect 1938 2912 2106 2924
rect 2121 2914 2137 2928
rect 2172 2915 2194 2934
rect 2204 2928 2220 2929
rect 2203 2926 2220 2928
rect 2204 2921 2220 2926
rect 2194 2914 2200 2915
rect 2203 2914 2232 2921
rect 2121 2913 2232 2914
rect 2121 2912 2238 2913
rect 1797 2904 1848 2912
rect 1895 2904 1929 2912
rect 1797 2892 1822 2904
rect 1829 2892 1848 2904
rect 1902 2902 1929 2904
rect 1938 2902 2159 2912
rect 2194 2909 2200 2912
rect 1902 2898 2159 2902
rect 1797 2884 1848 2892
rect 1895 2884 2159 2898
rect 2203 2904 2238 2912
rect 1749 2836 1768 2870
rect 1813 2876 1842 2884
rect 1813 2870 1830 2876
rect 1813 2868 1847 2870
rect 1895 2868 1911 2884
rect 1912 2874 2120 2884
rect 2121 2874 2137 2884
rect 2185 2880 2200 2895
rect 2203 2892 2204 2904
rect 2211 2892 2238 2904
rect 2203 2884 2238 2892
rect 2203 2883 2232 2884
rect 1923 2870 2137 2874
rect 1938 2868 2137 2870
rect 2172 2870 2185 2880
rect 2203 2870 2220 2883
rect 2172 2868 2220 2870
rect 1814 2864 1847 2868
rect 1810 2862 1847 2864
rect 1810 2861 1877 2862
rect 1810 2856 1841 2861
rect 1847 2856 1877 2861
rect 1810 2852 1877 2856
rect 1783 2849 1877 2852
rect 1783 2842 1832 2849
rect 1783 2836 1813 2842
rect 1832 2837 1837 2842
rect 1749 2820 1829 2836
rect 1841 2828 1877 2849
rect 1938 2844 2127 2868
rect 2172 2867 2219 2868
rect 2185 2862 2219 2867
rect 1953 2841 2127 2844
rect 1946 2838 2127 2841
rect 2155 2861 2219 2862
rect 1749 2818 1768 2820
rect 1783 2818 1817 2820
rect 1749 2802 1829 2818
rect 1749 2796 1768 2802
rect 1465 2770 1568 2780
rect 1419 2768 1568 2770
rect 1589 2768 1624 2780
rect 1258 2766 1420 2768
rect 1270 2746 1289 2766
rect 1304 2764 1334 2766
rect 1153 2738 1194 2746
rect 1276 2742 1289 2746
rect 1341 2750 1420 2766
rect 1452 2766 1624 2768
rect 1452 2750 1531 2766
rect 1538 2764 1568 2766
rect 1116 2728 1145 2738
rect 1159 2728 1188 2738
rect 1203 2728 1233 2742
rect 1276 2728 1319 2742
rect 1341 2738 1531 2750
rect 1596 2746 1602 2766
rect 1326 2728 1356 2738
rect 1357 2728 1515 2738
rect 1519 2728 1549 2738
rect 1553 2728 1583 2742
rect 1611 2728 1624 2766
rect 1696 2780 1725 2796
rect 1739 2780 1768 2796
rect 1783 2786 1813 2802
rect 1841 2780 1847 2828
rect 1850 2822 1869 2828
rect 1884 2822 1914 2830
rect 1850 2814 1914 2822
rect 1850 2798 1930 2814
rect 1946 2807 2008 2838
rect 2024 2807 2086 2838
rect 2155 2836 2204 2861
rect 2219 2836 2249 2852
rect 2118 2822 2148 2830
rect 2155 2828 2265 2836
rect 2118 2814 2163 2822
rect 1850 2796 1869 2798
rect 1884 2796 1930 2798
rect 1850 2780 1930 2796
rect 1957 2794 1992 2807
rect 2033 2804 2070 2807
rect 2033 2802 2075 2804
rect 1962 2791 1992 2794
rect 1971 2787 1978 2791
rect 1978 2786 1979 2787
rect 1937 2780 1947 2786
rect 1696 2772 1731 2780
rect 1696 2746 1697 2772
rect 1704 2746 1731 2772
rect 1639 2728 1669 2742
rect 1696 2738 1731 2746
rect 1733 2772 1774 2780
rect 1733 2746 1748 2772
rect 1755 2746 1774 2772
rect 1838 2768 1869 2780
rect 1884 2768 1987 2780
rect 1999 2770 2025 2796
rect 2040 2791 2070 2802
rect 2102 2798 2164 2814
rect 2102 2796 2148 2798
rect 2102 2780 2164 2796
rect 2176 2780 2182 2828
rect 2185 2820 2265 2828
rect 2185 2818 2204 2820
rect 2219 2818 2253 2820
rect 2185 2802 2265 2818
rect 2185 2780 2204 2802
rect 2219 2786 2249 2802
rect 2277 2796 2283 2870
rect 2286 2796 2305 2940
rect 2320 2796 2326 2940
rect 2335 2870 2348 2940
rect 2400 2936 2422 2940
rect 2393 2914 2422 2928
rect 2475 2914 2491 2928
rect 2529 2924 2535 2926
rect 2542 2924 2650 2940
rect 2657 2924 2663 2926
rect 2671 2924 2686 2940
rect 2752 2934 2771 2937
rect 2393 2912 2491 2914
rect 2518 2912 2686 2924
rect 2701 2914 2717 2928
rect 2752 2915 2774 2934
rect 2784 2928 2800 2929
rect 2783 2926 2800 2928
rect 2784 2921 2800 2926
rect 2774 2914 2780 2915
rect 2783 2914 2812 2921
rect 2701 2913 2812 2914
rect 2701 2912 2818 2913
rect 2377 2904 2428 2912
rect 2475 2904 2509 2912
rect 2377 2892 2402 2904
rect 2409 2892 2428 2904
rect 2482 2902 2509 2904
rect 2518 2902 2739 2912
rect 2774 2909 2780 2912
rect 2482 2898 2739 2902
rect 2377 2884 2428 2892
rect 2475 2884 2739 2898
rect 2783 2904 2818 2912
rect 2329 2836 2348 2870
rect 2393 2876 2422 2884
rect 2393 2870 2410 2876
rect 2393 2868 2427 2870
rect 2475 2868 2491 2884
rect 2492 2874 2700 2884
rect 2701 2874 2717 2884
rect 2765 2880 2780 2895
rect 2783 2892 2784 2904
rect 2791 2892 2818 2904
rect 2783 2884 2818 2892
rect 2783 2883 2812 2884
rect 2503 2870 2717 2874
rect 2518 2868 2717 2870
rect 2752 2870 2765 2880
rect 2783 2870 2800 2883
rect 2752 2868 2800 2870
rect 2394 2864 2427 2868
rect 2390 2862 2427 2864
rect 2390 2861 2457 2862
rect 2390 2856 2421 2861
rect 2427 2856 2457 2861
rect 2390 2852 2457 2856
rect 2363 2849 2457 2852
rect 2363 2842 2412 2849
rect 2363 2836 2393 2842
rect 2412 2837 2417 2842
rect 2329 2820 2409 2836
rect 2421 2828 2457 2849
rect 2518 2844 2707 2868
rect 2752 2867 2799 2868
rect 2765 2862 2799 2867
rect 2533 2841 2707 2844
rect 2526 2838 2707 2841
rect 2735 2861 2799 2862
rect 2329 2818 2348 2820
rect 2363 2818 2397 2820
rect 2329 2802 2409 2818
rect 2329 2796 2348 2802
rect 2045 2770 2148 2780
rect 1999 2768 2148 2770
rect 2169 2768 2204 2780
rect 1838 2766 2000 2768
rect 1850 2746 1869 2766
rect 1884 2764 1914 2766
rect 1733 2738 1774 2746
rect 1856 2742 1869 2746
rect 1921 2750 2000 2766
rect 2032 2766 2204 2768
rect 2032 2750 2111 2766
rect 2118 2764 2148 2766
rect 1696 2728 1725 2738
rect 1739 2728 1768 2738
rect 1783 2728 1813 2742
rect 1856 2728 1899 2742
rect 1921 2738 2111 2750
rect 2176 2746 2182 2766
rect 1906 2728 1936 2738
rect 1937 2728 2095 2738
rect 2099 2728 2129 2738
rect 2133 2728 2163 2742
rect 2191 2728 2204 2766
rect 2276 2780 2305 2796
rect 2319 2780 2348 2796
rect 2363 2786 2393 2802
rect 2421 2780 2427 2828
rect 2430 2822 2449 2828
rect 2464 2822 2494 2830
rect 2430 2814 2494 2822
rect 2430 2798 2510 2814
rect 2526 2807 2588 2838
rect 2604 2807 2666 2838
rect 2735 2836 2784 2861
rect 2799 2836 2829 2852
rect 2698 2822 2728 2830
rect 2735 2828 2845 2836
rect 2698 2814 2743 2822
rect 2430 2796 2449 2798
rect 2464 2796 2510 2798
rect 2430 2780 2510 2796
rect 2537 2794 2572 2807
rect 2613 2804 2650 2807
rect 2613 2802 2655 2804
rect 2542 2791 2572 2794
rect 2551 2787 2558 2791
rect 2558 2786 2559 2787
rect 2517 2780 2527 2786
rect 2276 2772 2311 2780
rect 2276 2746 2277 2772
rect 2284 2746 2311 2772
rect 2219 2728 2249 2742
rect 2276 2738 2311 2746
rect 2313 2772 2354 2780
rect 2313 2746 2328 2772
rect 2335 2746 2354 2772
rect 2418 2768 2449 2780
rect 2464 2768 2567 2780
rect 2579 2770 2605 2796
rect 2620 2791 2650 2802
rect 2682 2798 2744 2814
rect 2682 2796 2728 2798
rect 2682 2780 2744 2796
rect 2756 2780 2762 2828
rect 2765 2820 2845 2828
rect 2765 2818 2784 2820
rect 2799 2818 2833 2820
rect 2765 2802 2845 2818
rect 2765 2780 2784 2802
rect 2799 2786 2829 2802
rect 2857 2796 2863 2870
rect 2866 2796 2885 2940
rect 2900 2796 2906 2940
rect 2915 2870 2928 2940
rect 2980 2936 3002 2940
rect 2973 2914 3002 2928
rect 3055 2914 3071 2928
rect 3109 2924 3115 2926
rect 3122 2924 3230 2940
rect 3237 2924 3243 2926
rect 3251 2924 3266 2940
rect 3332 2934 3351 2937
rect 2973 2912 3071 2914
rect 3098 2912 3266 2924
rect 3281 2914 3297 2928
rect 3332 2915 3354 2934
rect 3364 2928 3380 2929
rect 3363 2926 3380 2928
rect 3364 2921 3380 2926
rect 3354 2914 3360 2915
rect 3363 2914 3392 2921
rect 3281 2913 3392 2914
rect 3281 2912 3398 2913
rect 2957 2904 3008 2912
rect 3055 2904 3089 2912
rect 2957 2892 2982 2904
rect 2989 2892 3008 2904
rect 3062 2902 3089 2904
rect 3098 2902 3319 2912
rect 3354 2909 3360 2912
rect 3062 2898 3319 2902
rect 2957 2884 3008 2892
rect 3055 2884 3319 2898
rect 3363 2904 3398 2912
rect 2909 2836 2928 2870
rect 2973 2876 3002 2884
rect 2973 2870 2990 2876
rect 2973 2868 3007 2870
rect 3055 2868 3071 2884
rect 3072 2874 3280 2884
rect 3281 2874 3297 2884
rect 3345 2880 3360 2895
rect 3363 2892 3364 2904
rect 3371 2892 3398 2904
rect 3363 2884 3398 2892
rect 3363 2883 3392 2884
rect 3083 2870 3297 2874
rect 3098 2868 3297 2870
rect 3332 2870 3345 2880
rect 3363 2870 3380 2883
rect 3332 2868 3380 2870
rect 2974 2864 3007 2868
rect 2970 2862 3007 2864
rect 2970 2861 3037 2862
rect 2970 2856 3001 2861
rect 3007 2856 3037 2861
rect 2970 2852 3037 2856
rect 2943 2849 3037 2852
rect 2943 2842 2992 2849
rect 2943 2836 2973 2842
rect 2992 2837 2997 2842
rect 2909 2820 2989 2836
rect 3001 2828 3037 2849
rect 3098 2844 3287 2868
rect 3332 2867 3379 2868
rect 3345 2862 3379 2867
rect 3113 2841 3287 2844
rect 3106 2838 3287 2841
rect 3315 2861 3379 2862
rect 2909 2818 2928 2820
rect 2943 2818 2977 2820
rect 2909 2802 2989 2818
rect 2909 2796 2928 2802
rect 2625 2770 2728 2780
rect 2579 2768 2728 2770
rect 2749 2768 2784 2780
rect 2418 2766 2580 2768
rect 2430 2746 2449 2766
rect 2464 2764 2494 2766
rect 2313 2738 2354 2746
rect 2436 2742 2449 2746
rect 2501 2750 2580 2766
rect 2612 2766 2784 2768
rect 2612 2750 2691 2766
rect 2698 2764 2728 2766
rect 2276 2728 2305 2738
rect 2319 2728 2348 2738
rect 2363 2728 2393 2742
rect 2436 2728 2479 2742
rect 2501 2738 2691 2750
rect 2756 2746 2762 2766
rect 2486 2728 2516 2738
rect 2517 2728 2675 2738
rect 2679 2728 2709 2738
rect 2713 2728 2743 2742
rect 2771 2728 2784 2766
rect 2856 2780 2885 2796
rect 2899 2780 2928 2796
rect 2943 2786 2973 2802
rect 3001 2780 3007 2828
rect 3010 2822 3029 2828
rect 3044 2822 3074 2830
rect 3010 2814 3074 2822
rect 3010 2798 3090 2814
rect 3106 2807 3168 2838
rect 3184 2807 3246 2838
rect 3315 2836 3364 2861
rect 3379 2836 3409 2852
rect 3278 2822 3308 2830
rect 3315 2828 3425 2836
rect 3278 2814 3323 2822
rect 3010 2796 3029 2798
rect 3044 2796 3090 2798
rect 3010 2780 3090 2796
rect 3117 2794 3152 2807
rect 3193 2804 3230 2807
rect 3193 2802 3235 2804
rect 3122 2791 3152 2794
rect 3131 2787 3138 2791
rect 3138 2786 3139 2787
rect 3097 2780 3107 2786
rect 2856 2772 2891 2780
rect 2856 2746 2857 2772
rect 2864 2746 2891 2772
rect 2799 2728 2829 2742
rect 2856 2738 2891 2746
rect 2893 2772 2934 2780
rect 2893 2746 2908 2772
rect 2915 2746 2934 2772
rect 2998 2768 3029 2780
rect 3044 2768 3147 2780
rect 3159 2770 3185 2796
rect 3200 2791 3230 2802
rect 3262 2798 3324 2814
rect 3262 2796 3308 2798
rect 3262 2780 3324 2796
rect 3336 2780 3342 2828
rect 3345 2820 3425 2828
rect 3345 2818 3364 2820
rect 3379 2818 3413 2820
rect 3345 2802 3425 2818
rect 3345 2780 3364 2802
rect 3379 2786 3409 2802
rect 3437 2796 3443 2870
rect 3446 2796 3465 2940
rect 3480 2796 3486 2940
rect 3495 2870 3508 2940
rect 3560 2936 3582 2940
rect 3553 2914 3582 2928
rect 3635 2914 3651 2928
rect 3689 2924 3695 2926
rect 3702 2924 3810 2940
rect 3817 2924 3823 2926
rect 3831 2924 3846 2940
rect 3912 2934 3931 2937
rect 3553 2912 3651 2914
rect 3678 2912 3846 2924
rect 3861 2914 3877 2928
rect 3912 2915 3934 2934
rect 3944 2928 3960 2929
rect 3943 2926 3960 2928
rect 3944 2921 3960 2926
rect 3934 2914 3940 2915
rect 3943 2914 3972 2921
rect 3861 2913 3972 2914
rect 3861 2912 3978 2913
rect 3537 2904 3588 2912
rect 3635 2904 3669 2912
rect 3537 2892 3562 2904
rect 3569 2892 3588 2904
rect 3642 2902 3669 2904
rect 3678 2902 3899 2912
rect 3934 2909 3940 2912
rect 3642 2898 3899 2902
rect 3537 2884 3588 2892
rect 3635 2884 3899 2898
rect 3943 2904 3978 2912
rect 3489 2836 3508 2870
rect 3553 2876 3582 2884
rect 3553 2870 3570 2876
rect 3553 2868 3587 2870
rect 3635 2868 3651 2884
rect 3652 2874 3860 2884
rect 3861 2874 3877 2884
rect 3925 2880 3940 2895
rect 3943 2892 3944 2904
rect 3951 2892 3978 2904
rect 3943 2884 3978 2892
rect 3943 2883 3972 2884
rect 3663 2870 3877 2874
rect 3678 2868 3877 2870
rect 3912 2870 3925 2880
rect 3943 2870 3960 2883
rect 3912 2868 3960 2870
rect 3554 2864 3587 2868
rect 3550 2862 3587 2864
rect 3550 2861 3617 2862
rect 3550 2856 3581 2861
rect 3587 2856 3617 2861
rect 3550 2852 3617 2856
rect 3523 2849 3617 2852
rect 3523 2842 3572 2849
rect 3523 2836 3553 2842
rect 3572 2837 3577 2842
rect 3489 2820 3569 2836
rect 3581 2828 3617 2849
rect 3678 2844 3867 2868
rect 3912 2867 3959 2868
rect 3925 2862 3959 2867
rect 3693 2841 3867 2844
rect 3686 2838 3867 2841
rect 3895 2861 3959 2862
rect 3489 2818 3508 2820
rect 3523 2818 3557 2820
rect 3489 2802 3569 2818
rect 3489 2796 3508 2802
rect 3205 2770 3308 2780
rect 3159 2768 3308 2770
rect 3329 2768 3364 2780
rect 2998 2766 3160 2768
rect 3010 2746 3029 2766
rect 3044 2764 3074 2766
rect 2893 2738 2934 2746
rect 3016 2742 3029 2746
rect 3081 2750 3160 2766
rect 3192 2766 3364 2768
rect 3192 2750 3271 2766
rect 3278 2764 3308 2766
rect 2856 2728 2885 2738
rect 2899 2728 2928 2738
rect 2943 2728 2973 2742
rect 3016 2728 3059 2742
rect 3081 2738 3271 2750
rect 3336 2746 3342 2766
rect 3066 2728 3096 2738
rect 3097 2728 3255 2738
rect 3259 2728 3289 2738
rect 3293 2728 3323 2742
rect 3351 2728 3364 2766
rect 3436 2780 3465 2796
rect 3479 2780 3508 2796
rect 3523 2786 3553 2802
rect 3581 2780 3587 2828
rect 3590 2822 3609 2828
rect 3624 2822 3654 2830
rect 3590 2814 3654 2822
rect 3590 2798 3670 2814
rect 3686 2807 3748 2838
rect 3764 2807 3826 2838
rect 3895 2836 3944 2861
rect 3959 2836 3989 2852
rect 3858 2822 3888 2830
rect 3895 2828 4005 2836
rect 3858 2814 3903 2822
rect 3590 2796 3609 2798
rect 3624 2796 3670 2798
rect 3590 2780 3670 2796
rect 3697 2794 3732 2807
rect 3773 2804 3810 2807
rect 3773 2802 3815 2804
rect 3702 2791 3732 2794
rect 3711 2787 3718 2791
rect 3718 2786 3719 2787
rect 3677 2780 3687 2786
rect 3436 2772 3471 2780
rect 3436 2746 3437 2772
rect 3444 2746 3471 2772
rect 3379 2728 3409 2742
rect 3436 2738 3471 2746
rect 3473 2772 3514 2780
rect 3473 2746 3488 2772
rect 3495 2746 3514 2772
rect 3578 2768 3609 2780
rect 3624 2768 3727 2780
rect 3739 2770 3765 2796
rect 3780 2791 3810 2802
rect 3842 2798 3904 2814
rect 3842 2796 3888 2798
rect 3842 2780 3904 2796
rect 3916 2780 3922 2828
rect 3925 2820 4005 2828
rect 3925 2818 3944 2820
rect 3959 2818 3993 2820
rect 3925 2802 4005 2818
rect 3925 2780 3944 2802
rect 3959 2786 3989 2802
rect 4017 2796 4023 2870
rect 4026 2796 4045 2940
rect 4060 2796 4066 2940
rect 4075 2870 4088 2940
rect 4140 2936 4162 2940
rect 4133 2914 4162 2928
rect 4215 2914 4231 2928
rect 4269 2924 4275 2926
rect 4282 2924 4390 2940
rect 4397 2924 4403 2926
rect 4411 2924 4426 2940
rect 4492 2934 4511 2937
rect 4133 2912 4231 2914
rect 4258 2912 4426 2924
rect 4441 2914 4457 2928
rect 4492 2915 4514 2934
rect 4524 2928 4540 2929
rect 4523 2926 4540 2928
rect 4524 2921 4540 2926
rect 4514 2914 4520 2915
rect 4523 2914 4552 2921
rect 4441 2913 4552 2914
rect 4441 2912 4558 2913
rect 4117 2904 4168 2912
rect 4215 2904 4249 2912
rect 4117 2892 4142 2904
rect 4149 2892 4168 2904
rect 4222 2902 4249 2904
rect 4258 2902 4479 2912
rect 4514 2909 4520 2912
rect 4222 2898 4479 2902
rect 4117 2884 4168 2892
rect 4215 2884 4479 2898
rect 4523 2904 4558 2912
rect 4069 2836 4088 2870
rect 4133 2876 4162 2884
rect 4133 2870 4150 2876
rect 4133 2868 4167 2870
rect 4215 2868 4231 2884
rect 4232 2874 4440 2884
rect 4441 2874 4457 2884
rect 4505 2880 4520 2895
rect 4523 2892 4524 2904
rect 4531 2892 4558 2904
rect 4523 2884 4558 2892
rect 4523 2883 4552 2884
rect 4243 2870 4457 2874
rect 4258 2868 4457 2870
rect 4492 2870 4505 2880
rect 4523 2870 4540 2883
rect 4492 2868 4540 2870
rect 4134 2864 4167 2868
rect 4130 2862 4167 2864
rect 4130 2861 4197 2862
rect 4130 2856 4161 2861
rect 4167 2856 4197 2861
rect 4130 2852 4197 2856
rect 4103 2849 4197 2852
rect 4103 2842 4152 2849
rect 4103 2836 4133 2842
rect 4152 2837 4157 2842
rect 4069 2820 4149 2836
rect 4161 2828 4197 2849
rect 4258 2844 4447 2868
rect 4492 2867 4539 2868
rect 4505 2862 4539 2867
rect 4273 2841 4447 2844
rect 4266 2838 4447 2841
rect 4475 2861 4539 2862
rect 4069 2818 4088 2820
rect 4103 2818 4137 2820
rect 4069 2802 4149 2818
rect 4069 2796 4088 2802
rect 3785 2770 3888 2780
rect 3739 2768 3888 2770
rect 3909 2768 3944 2780
rect 3578 2766 3740 2768
rect 3590 2746 3609 2766
rect 3624 2764 3654 2766
rect 3473 2738 3514 2746
rect 3596 2742 3609 2746
rect 3661 2750 3740 2766
rect 3772 2766 3944 2768
rect 3772 2750 3851 2766
rect 3858 2764 3888 2766
rect 3436 2728 3465 2738
rect 3479 2728 3508 2738
rect 3523 2728 3553 2742
rect 3596 2728 3639 2742
rect 3661 2738 3851 2750
rect 3916 2746 3922 2766
rect 3646 2728 3676 2738
rect 3677 2728 3835 2738
rect 3839 2728 3869 2738
rect 3873 2728 3903 2742
rect 3931 2728 3944 2766
rect 4016 2780 4045 2796
rect 4059 2780 4088 2796
rect 4103 2786 4133 2802
rect 4161 2780 4167 2828
rect 4170 2822 4189 2828
rect 4204 2822 4234 2830
rect 4170 2814 4234 2822
rect 4170 2798 4250 2814
rect 4266 2807 4328 2838
rect 4344 2807 4406 2838
rect 4475 2836 4524 2861
rect 4539 2836 4569 2852
rect 4438 2822 4468 2830
rect 4475 2828 4585 2836
rect 4438 2814 4483 2822
rect 4170 2796 4189 2798
rect 4204 2796 4250 2798
rect 4170 2780 4250 2796
rect 4277 2794 4312 2807
rect 4353 2804 4390 2807
rect 4353 2802 4395 2804
rect 4282 2791 4312 2794
rect 4291 2787 4298 2791
rect 4298 2786 4299 2787
rect 4257 2780 4267 2786
rect 4016 2772 4051 2780
rect 4016 2746 4017 2772
rect 4024 2746 4051 2772
rect 3959 2728 3989 2742
rect 4016 2738 4051 2746
rect 4053 2772 4094 2780
rect 4053 2746 4068 2772
rect 4075 2746 4094 2772
rect 4158 2768 4189 2780
rect 4204 2768 4307 2780
rect 4319 2770 4345 2796
rect 4360 2791 4390 2802
rect 4422 2798 4484 2814
rect 4422 2796 4468 2798
rect 4422 2780 4484 2796
rect 4496 2780 4502 2828
rect 4505 2820 4585 2828
rect 4505 2818 4524 2820
rect 4539 2818 4573 2820
rect 4505 2802 4585 2818
rect 4505 2780 4524 2802
rect 4539 2786 4569 2802
rect 4597 2796 4603 2870
rect 4606 2796 4625 2940
rect 4640 2796 4646 2940
rect 4655 2870 4668 2940
rect 4720 2936 4742 2940
rect 4713 2914 4742 2928
rect 4795 2914 4811 2928
rect 4849 2924 4855 2926
rect 4862 2924 4970 2940
rect 4977 2924 4983 2926
rect 4991 2924 5006 2940
rect 5072 2934 5091 2937
rect 4713 2912 4811 2914
rect 4838 2912 5006 2924
rect 5021 2914 5037 2928
rect 5072 2915 5094 2934
rect 5104 2928 5120 2929
rect 5103 2926 5120 2928
rect 5104 2921 5120 2926
rect 5094 2914 5100 2915
rect 5103 2914 5132 2921
rect 5021 2913 5132 2914
rect 5021 2912 5138 2913
rect 4697 2904 4748 2912
rect 4795 2904 4829 2912
rect 4697 2892 4722 2904
rect 4729 2892 4748 2904
rect 4802 2902 4829 2904
rect 4838 2902 5059 2912
rect 5094 2909 5100 2912
rect 4802 2898 5059 2902
rect 4697 2884 4748 2892
rect 4795 2884 5059 2898
rect 5103 2904 5138 2912
rect 4649 2836 4668 2870
rect 4713 2876 4742 2884
rect 4713 2870 4730 2876
rect 4713 2868 4747 2870
rect 4795 2868 4811 2884
rect 4812 2874 5020 2884
rect 5021 2874 5037 2884
rect 5085 2880 5100 2895
rect 5103 2892 5104 2904
rect 5111 2892 5138 2904
rect 5103 2884 5138 2892
rect 5103 2883 5132 2884
rect 4823 2870 5037 2874
rect 4838 2868 5037 2870
rect 5072 2870 5085 2880
rect 5103 2870 5120 2883
rect 5072 2868 5120 2870
rect 4714 2864 4747 2868
rect 4710 2862 4747 2864
rect 4710 2861 4777 2862
rect 4710 2856 4741 2861
rect 4747 2856 4777 2861
rect 4710 2852 4777 2856
rect 4683 2849 4777 2852
rect 4683 2842 4732 2849
rect 4683 2836 4713 2842
rect 4732 2837 4737 2842
rect 4649 2820 4729 2836
rect 4741 2828 4777 2849
rect 4838 2844 5027 2868
rect 5072 2867 5119 2868
rect 5085 2862 5119 2867
rect 4853 2841 5027 2844
rect 4846 2838 5027 2841
rect 5055 2861 5119 2862
rect 4649 2818 4668 2820
rect 4683 2818 4717 2820
rect 4649 2802 4729 2818
rect 4649 2796 4668 2802
rect 4365 2770 4468 2780
rect 4319 2768 4468 2770
rect 4489 2768 4524 2780
rect 4158 2766 4320 2768
rect 4170 2746 4189 2766
rect 4204 2764 4234 2766
rect 4053 2738 4094 2746
rect 4176 2742 4189 2746
rect 4241 2750 4320 2766
rect 4352 2766 4524 2768
rect 4352 2750 4431 2766
rect 4438 2764 4468 2766
rect 4016 2728 4045 2738
rect 4059 2728 4088 2738
rect 4103 2728 4133 2742
rect 4176 2728 4219 2742
rect 4241 2738 4431 2750
rect 4496 2746 4502 2766
rect 4226 2728 4256 2738
rect 4257 2728 4415 2738
rect 4419 2728 4449 2738
rect 4453 2728 4483 2742
rect 4511 2728 4524 2766
rect 4596 2780 4625 2796
rect 4639 2780 4668 2796
rect 4683 2786 4713 2802
rect 4741 2780 4747 2828
rect 4750 2822 4769 2828
rect 4784 2822 4814 2830
rect 4750 2814 4814 2822
rect 4750 2798 4830 2814
rect 4846 2807 4908 2838
rect 4924 2807 4986 2838
rect 5055 2836 5104 2861
rect 5119 2836 5149 2852
rect 5018 2822 5048 2830
rect 5055 2828 5165 2836
rect 5018 2814 5063 2822
rect 4750 2796 4769 2798
rect 4784 2796 4830 2798
rect 4750 2780 4830 2796
rect 4857 2794 4892 2807
rect 4933 2804 4970 2807
rect 4933 2802 4975 2804
rect 4862 2791 4892 2794
rect 4871 2787 4878 2791
rect 4878 2786 4879 2787
rect 4837 2780 4847 2786
rect 4596 2772 4631 2780
rect 4596 2746 4597 2772
rect 4604 2746 4631 2772
rect 4539 2728 4569 2742
rect 4596 2738 4631 2746
rect 4633 2772 4674 2780
rect 4633 2746 4648 2772
rect 4655 2746 4674 2772
rect 4738 2768 4769 2780
rect 4784 2768 4887 2780
rect 4899 2770 4925 2796
rect 4940 2791 4970 2802
rect 5002 2798 5064 2814
rect 5002 2796 5048 2798
rect 5002 2780 5064 2796
rect 5076 2780 5082 2828
rect 5085 2820 5165 2828
rect 5085 2818 5104 2820
rect 5119 2818 5153 2820
rect 5085 2802 5165 2818
rect 5085 2780 5104 2802
rect 5119 2786 5149 2802
rect 5177 2796 5183 2870
rect 5186 2796 5205 2940
rect 5220 2796 5226 2940
rect 5235 2870 5248 2940
rect 5300 2936 5322 2940
rect 5293 2914 5322 2928
rect 5375 2914 5391 2928
rect 5429 2924 5435 2926
rect 5442 2924 5550 2940
rect 5557 2924 5563 2926
rect 5571 2924 5586 2940
rect 5652 2934 5671 2937
rect 5293 2912 5391 2914
rect 5418 2912 5586 2924
rect 5601 2914 5617 2928
rect 5652 2915 5674 2934
rect 5684 2928 5700 2929
rect 5683 2926 5700 2928
rect 5684 2921 5700 2926
rect 5674 2914 5680 2915
rect 5683 2914 5712 2921
rect 5601 2913 5712 2914
rect 5601 2912 5718 2913
rect 5277 2904 5328 2912
rect 5375 2904 5409 2912
rect 5277 2892 5302 2904
rect 5309 2892 5328 2904
rect 5382 2902 5409 2904
rect 5418 2902 5639 2912
rect 5674 2909 5680 2912
rect 5382 2898 5639 2902
rect 5277 2884 5328 2892
rect 5375 2884 5639 2898
rect 5683 2904 5718 2912
rect 5229 2836 5248 2870
rect 5293 2876 5322 2884
rect 5293 2870 5310 2876
rect 5293 2868 5327 2870
rect 5375 2868 5391 2884
rect 5392 2874 5600 2884
rect 5601 2874 5617 2884
rect 5665 2880 5680 2895
rect 5683 2892 5684 2904
rect 5691 2892 5718 2904
rect 5683 2884 5718 2892
rect 5683 2883 5712 2884
rect 5403 2870 5617 2874
rect 5418 2868 5617 2870
rect 5652 2870 5665 2880
rect 5683 2870 5700 2883
rect 5652 2868 5700 2870
rect 5294 2864 5327 2868
rect 5290 2862 5327 2864
rect 5290 2861 5357 2862
rect 5290 2856 5321 2861
rect 5327 2856 5357 2861
rect 5290 2852 5357 2856
rect 5263 2849 5357 2852
rect 5263 2842 5312 2849
rect 5263 2836 5293 2842
rect 5312 2837 5317 2842
rect 5229 2820 5309 2836
rect 5321 2828 5357 2849
rect 5418 2844 5607 2868
rect 5652 2867 5699 2868
rect 5665 2862 5699 2867
rect 5433 2841 5607 2844
rect 5426 2838 5607 2841
rect 5635 2861 5699 2862
rect 5229 2818 5248 2820
rect 5263 2818 5297 2820
rect 5229 2802 5309 2818
rect 5229 2796 5248 2802
rect 4945 2770 5048 2780
rect 4899 2768 5048 2770
rect 5069 2768 5104 2780
rect 4738 2766 4900 2768
rect 4750 2746 4769 2766
rect 4784 2764 4814 2766
rect 4633 2738 4674 2746
rect 4756 2742 4769 2746
rect 4821 2750 4900 2766
rect 4932 2766 5104 2768
rect 4932 2750 5011 2766
rect 5018 2764 5048 2766
rect 4596 2728 4625 2738
rect 4639 2728 4668 2738
rect 4683 2728 4713 2742
rect 4756 2728 4799 2742
rect 4821 2738 5011 2750
rect 5076 2746 5082 2766
rect 4806 2728 4836 2738
rect 4837 2728 4995 2738
rect 4999 2728 5029 2738
rect 5033 2728 5063 2742
rect 5091 2728 5104 2766
rect 5176 2780 5205 2796
rect 5219 2780 5248 2796
rect 5263 2786 5293 2802
rect 5321 2780 5327 2828
rect 5330 2822 5349 2828
rect 5364 2822 5394 2830
rect 5330 2814 5394 2822
rect 5330 2798 5410 2814
rect 5426 2807 5488 2838
rect 5504 2807 5566 2838
rect 5635 2836 5684 2861
rect 5699 2836 5729 2852
rect 5598 2822 5628 2830
rect 5635 2828 5745 2836
rect 5598 2814 5643 2822
rect 5330 2796 5349 2798
rect 5364 2796 5410 2798
rect 5330 2780 5410 2796
rect 5437 2794 5472 2807
rect 5513 2804 5550 2807
rect 5513 2802 5555 2804
rect 5442 2791 5472 2794
rect 5451 2787 5458 2791
rect 5458 2786 5459 2787
rect 5417 2780 5427 2786
rect 5176 2772 5211 2780
rect 5176 2746 5177 2772
rect 5184 2746 5211 2772
rect 5119 2728 5149 2742
rect 5176 2738 5211 2746
rect 5213 2772 5254 2780
rect 5213 2746 5228 2772
rect 5235 2746 5254 2772
rect 5318 2768 5349 2780
rect 5364 2768 5467 2780
rect 5479 2770 5505 2796
rect 5520 2791 5550 2802
rect 5582 2798 5644 2814
rect 5582 2796 5628 2798
rect 5582 2780 5644 2796
rect 5656 2780 5662 2828
rect 5665 2820 5745 2828
rect 5665 2818 5684 2820
rect 5699 2818 5733 2820
rect 5665 2802 5745 2818
rect 5665 2780 5684 2802
rect 5699 2786 5729 2802
rect 5757 2796 5763 2870
rect 5766 2796 5785 2940
rect 5800 2796 5806 2940
rect 5815 2870 5828 2940
rect 5880 2936 5902 2940
rect 5873 2914 5902 2928
rect 5955 2914 5971 2928
rect 6009 2924 6015 2926
rect 6022 2924 6130 2940
rect 6137 2924 6143 2926
rect 6151 2924 6166 2940
rect 6232 2934 6251 2937
rect 5873 2912 5971 2914
rect 5998 2912 6166 2924
rect 6181 2914 6197 2928
rect 6232 2915 6254 2934
rect 6264 2928 6280 2929
rect 6263 2926 6280 2928
rect 6264 2921 6280 2926
rect 6254 2914 6260 2915
rect 6263 2914 6292 2921
rect 6181 2913 6292 2914
rect 6181 2912 6298 2913
rect 5857 2904 5908 2912
rect 5955 2904 5989 2912
rect 5857 2892 5882 2904
rect 5889 2892 5908 2904
rect 5962 2902 5989 2904
rect 5998 2902 6219 2912
rect 6254 2909 6260 2912
rect 5962 2898 6219 2902
rect 5857 2884 5908 2892
rect 5955 2884 6219 2898
rect 6263 2904 6298 2912
rect 5809 2836 5828 2870
rect 5873 2876 5902 2884
rect 5873 2870 5890 2876
rect 5873 2868 5907 2870
rect 5955 2868 5971 2884
rect 5972 2874 6180 2884
rect 6181 2874 6197 2884
rect 6245 2880 6260 2895
rect 6263 2892 6264 2904
rect 6271 2892 6298 2904
rect 6263 2884 6298 2892
rect 6263 2883 6292 2884
rect 5983 2870 6197 2874
rect 5998 2868 6197 2870
rect 6232 2870 6245 2880
rect 6263 2870 6280 2883
rect 6232 2868 6280 2870
rect 5874 2864 5907 2868
rect 5870 2862 5907 2864
rect 5870 2861 5937 2862
rect 5870 2856 5901 2861
rect 5907 2856 5937 2861
rect 5870 2852 5937 2856
rect 5843 2849 5937 2852
rect 5843 2842 5892 2849
rect 5843 2836 5873 2842
rect 5892 2837 5897 2842
rect 5809 2820 5889 2836
rect 5901 2828 5937 2849
rect 5998 2844 6187 2868
rect 6232 2867 6279 2868
rect 6245 2862 6279 2867
rect 6013 2841 6187 2844
rect 6006 2838 6187 2841
rect 6215 2861 6279 2862
rect 5809 2818 5828 2820
rect 5843 2818 5877 2820
rect 5809 2802 5889 2818
rect 5809 2796 5828 2802
rect 5525 2770 5628 2780
rect 5479 2768 5628 2770
rect 5649 2768 5684 2780
rect 5318 2766 5480 2768
rect 5330 2746 5349 2766
rect 5364 2764 5394 2766
rect 5213 2738 5254 2746
rect 5336 2742 5349 2746
rect 5401 2750 5480 2766
rect 5512 2766 5684 2768
rect 5512 2750 5591 2766
rect 5598 2764 5628 2766
rect 5176 2728 5205 2738
rect 5219 2728 5248 2738
rect 5263 2728 5293 2742
rect 5336 2728 5379 2742
rect 5401 2738 5591 2750
rect 5656 2746 5662 2766
rect 5386 2728 5416 2738
rect 5417 2728 5575 2738
rect 5579 2728 5609 2738
rect 5613 2728 5643 2742
rect 5671 2728 5684 2766
rect 5756 2780 5785 2796
rect 5799 2780 5828 2796
rect 5843 2786 5873 2802
rect 5901 2780 5907 2828
rect 5910 2822 5929 2828
rect 5944 2822 5974 2830
rect 5910 2814 5974 2822
rect 5910 2798 5990 2814
rect 6006 2807 6068 2838
rect 6084 2807 6146 2838
rect 6215 2836 6264 2861
rect 6279 2836 6309 2852
rect 6178 2822 6208 2830
rect 6215 2828 6325 2836
rect 6178 2814 6223 2822
rect 5910 2796 5929 2798
rect 5944 2796 5990 2798
rect 5910 2780 5990 2796
rect 6017 2794 6052 2807
rect 6093 2804 6130 2807
rect 6093 2802 6135 2804
rect 6022 2791 6052 2794
rect 6031 2787 6038 2791
rect 6038 2786 6039 2787
rect 5997 2780 6007 2786
rect 5756 2772 5791 2780
rect 5756 2746 5757 2772
rect 5764 2746 5791 2772
rect 5699 2728 5729 2742
rect 5756 2738 5791 2746
rect 5793 2772 5834 2780
rect 5793 2746 5808 2772
rect 5815 2746 5834 2772
rect 5898 2768 5929 2780
rect 5944 2768 6047 2780
rect 6059 2770 6085 2796
rect 6100 2791 6130 2802
rect 6162 2798 6224 2814
rect 6162 2796 6208 2798
rect 6162 2780 6224 2796
rect 6236 2780 6242 2828
rect 6245 2820 6325 2828
rect 6245 2818 6264 2820
rect 6279 2818 6313 2820
rect 6245 2802 6325 2818
rect 6245 2780 6264 2802
rect 6279 2786 6309 2802
rect 6337 2796 6343 2870
rect 6346 2796 6365 2940
rect 6380 2796 6386 2940
rect 6395 2870 6408 2940
rect 6460 2936 6482 2940
rect 6453 2914 6482 2928
rect 6535 2914 6551 2928
rect 6589 2924 6595 2926
rect 6602 2924 6710 2940
rect 6717 2924 6723 2926
rect 6731 2924 6746 2940
rect 6812 2934 6831 2937
rect 6453 2912 6551 2914
rect 6578 2912 6746 2924
rect 6761 2914 6777 2928
rect 6812 2915 6834 2934
rect 6844 2928 6860 2929
rect 6843 2926 6860 2928
rect 6844 2921 6860 2926
rect 6834 2914 6840 2915
rect 6843 2914 6872 2921
rect 6761 2913 6872 2914
rect 6761 2912 6878 2913
rect 6437 2904 6488 2912
rect 6535 2904 6569 2912
rect 6437 2892 6462 2904
rect 6469 2892 6488 2904
rect 6542 2902 6569 2904
rect 6578 2902 6799 2912
rect 6834 2909 6840 2912
rect 6542 2898 6799 2902
rect 6437 2884 6488 2892
rect 6535 2884 6799 2898
rect 6843 2904 6878 2912
rect 6389 2836 6408 2870
rect 6453 2876 6482 2884
rect 6453 2870 6470 2876
rect 6453 2868 6487 2870
rect 6535 2868 6551 2884
rect 6552 2874 6760 2884
rect 6761 2874 6777 2884
rect 6825 2880 6840 2895
rect 6843 2892 6844 2904
rect 6851 2892 6878 2904
rect 6843 2884 6878 2892
rect 6843 2883 6872 2884
rect 6563 2870 6777 2874
rect 6578 2868 6777 2870
rect 6812 2870 6825 2880
rect 6843 2870 6860 2883
rect 6812 2868 6860 2870
rect 6454 2864 6487 2868
rect 6450 2862 6487 2864
rect 6450 2861 6517 2862
rect 6450 2856 6481 2861
rect 6487 2856 6517 2861
rect 6450 2852 6517 2856
rect 6423 2849 6517 2852
rect 6423 2842 6472 2849
rect 6423 2836 6453 2842
rect 6472 2837 6477 2842
rect 6389 2820 6469 2836
rect 6481 2828 6517 2849
rect 6578 2844 6767 2868
rect 6812 2867 6859 2868
rect 6825 2862 6859 2867
rect 6593 2841 6767 2844
rect 6586 2838 6767 2841
rect 6795 2861 6859 2862
rect 6389 2818 6408 2820
rect 6423 2818 6457 2820
rect 6389 2802 6469 2818
rect 6389 2796 6408 2802
rect 6105 2770 6208 2780
rect 6059 2768 6208 2770
rect 6229 2768 6264 2780
rect 5898 2766 6060 2768
rect 5910 2746 5929 2766
rect 5944 2764 5974 2766
rect 5793 2738 5834 2746
rect 5916 2742 5929 2746
rect 5981 2750 6060 2766
rect 6092 2766 6264 2768
rect 6092 2750 6171 2766
rect 6178 2764 6208 2766
rect 5756 2728 5785 2738
rect 5799 2728 5828 2738
rect 5843 2728 5873 2742
rect 5916 2728 5959 2742
rect 5981 2738 6171 2750
rect 6236 2746 6242 2766
rect 5966 2728 5996 2738
rect 5997 2728 6155 2738
rect 6159 2728 6189 2738
rect 6193 2728 6223 2742
rect 6251 2728 6264 2766
rect 6336 2780 6365 2796
rect 6379 2780 6408 2796
rect 6423 2786 6453 2802
rect 6481 2780 6487 2828
rect 6490 2822 6509 2828
rect 6524 2822 6554 2830
rect 6490 2814 6554 2822
rect 6490 2798 6570 2814
rect 6586 2807 6648 2838
rect 6664 2807 6726 2838
rect 6795 2836 6844 2861
rect 6859 2836 6889 2852
rect 6758 2822 6788 2830
rect 6795 2828 6905 2836
rect 6758 2814 6803 2822
rect 6490 2796 6509 2798
rect 6524 2796 6570 2798
rect 6490 2780 6570 2796
rect 6597 2794 6632 2807
rect 6673 2804 6710 2807
rect 6673 2802 6715 2804
rect 6602 2791 6632 2794
rect 6611 2787 6618 2791
rect 6618 2786 6619 2787
rect 6577 2780 6587 2786
rect 6336 2772 6371 2780
rect 6336 2746 6337 2772
rect 6344 2746 6371 2772
rect 6279 2728 6309 2742
rect 6336 2738 6371 2746
rect 6373 2772 6414 2780
rect 6373 2746 6388 2772
rect 6395 2746 6414 2772
rect 6478 2768 6509 2780
rect 6524 2768 6627 2780
rect 6639 2770 6665 2796
rect 6680 2791 6710 2802
rect 6742 2798 6804 2814
rect 6742 2796 6788 2798
rect 6742 2780 6804 2796
rect 6816 2780 6822 2828
rect 6825 2820 6905 2828
rect 6825 2818 6844 2820
rect 6859 2818 6893 2820
rect 6825 2802 6905 2818
rect 6825 2780 6844 2802
rect 6859 2786 6889 2802
rect 6917 2796 6923 2870
rect 6926 2796 6945 2940
rect 6960 2796 6966 2940
rect 6975 2870 6988 2940
rect 7040 2936 7062 2940
rect 7033 2914 7062 2928
rect 7115 2914 7131 2928
rect 7169 2924 7175 2926
rect 7182 2924 7290 2940
rect 7297 2924 7303 2926
rect 7311 2924 7326 2940
rect 7392 2934 7411 2937
rect 7033 2912 7131 2914
rect 7158 2912 7326 2924
rect 7341 2914 7357 2928
rect 7392 2915 7414 2934
rect 7424 2928 7440 2929
rect 7423 2926 7440 2928
rect 7424 2921 7440 2926
rect 7414 2914 7420 2915
rect 7423 2914 7452 2921
rect 7341 2913 7452 2914
rect 7341 2912 7458 2913
rect 7017 2904 7068 2912
rect 7115 2904 7149 2912
rect 7017 2892 7042 2904
rect 7049 2892 7068 2904
rect 7122 2902 7149 2904
rect 7158 2902 7379 2912
rect 7414 2909 7420 2912
rect 7122 2898 7379 2902
rect 7017 2884 7068 2892
rect 7115 2884 7379 2898
rect 7423 2904 7458 2912
rect 6969 2836 6988 2870
rect 7033 2876 7062 2884
rect 7033 2870 7050 2876
rect 7033 2868 7067 2870
rect 7115 2868 7131 2884
rect 7132 2874 7340 2884
rect 7341 2874 7357 2884
rect 7405 2880 7420 2895
rect 7423 2892 7424 2904
rect 7431 2892 7458 2904
rect 7423 2884 7458 2892
rect 7423 2883 7452 2884
rect 7143 2870 7357 2874
rect 7158 2868 7357 2870
rect 7392 2870 7405 2880
rect 7423 2870 7440 2883
rect 7392 2868 7440 2870
rect 7034 2864 7067 2868
rect 7030 2862 7067 2864
rect 7030 2861 7097 2862
rect 7030 2856 7061 2861
rect 7067 2856 7097 2861
rect 7030 2852 7097 2856
rect 7003 2849 7097 2852
rect 7003 2842 7052 2849
rect 7003 2836 7033 2842
rect 7052 2837 7057 2842
rect 6969 2820 7049 2836
rect 7061 2828 7097 2849
rect 7158 2844 7347 2868
rect 7392 2867 7439 2868
rect 7405 2862 7439 2867
rect 7173 2841 7347 2844
rect 7166 2838 7347 2841
rect 7375 2861 7439 2862
rect 6969 2818 6988 2820
rect 7003 2818 7037 2820
rect 6969 2802 7049 2818
rect 6969 2796 6988 2802
rect 6685 2770 6788 2780
rect 6639 2768 6788 2770
rect 6809 2768 6844 2780
rect 6478 2766 6640 2768
rect 6490 2746 6509 2766
rect 6524 2764 6554 2766
rect 6373 2738 6414 2746
rect 6496 2742 6509 2746
rect 6561 2750 6640 2766
rect 6672 2766 6844 2768
rect 6672 2750 6751 2766
rect 6758 2764 6788 2766
rect 6336 2728 6365 2738
rect 6379 2728 6408 2738
rect 6423 2728 6453 2742
rect 6496 2728 6539 2742
rect 6561 2738 6751 2750
rect 6816 2746 6822 2766
rect 6546 2728 6576 2738
rect 6577 2728 6735 2738
rect 6739 2728 6769 2738
rect 6773 2728 6803 2742
rect 6831 2728 6844 2766
rect 6916 2780 6945 2796
rect 6959 2780 6988 2796
rect 7003 2786 7033 2802
rect 7061 2780 7067 2828
rect 7070 2822 7089 2828
rect 7104 2822 7134 2830
rect 7070 2814 7134 2822
rect 7070 2798 7150 2814
rect 7166 2807 7228 2838
rect 7244 2807 7306 2838
rect 7375 2836 7424 2861
rect 7439 2836 7469 2852
rect 7338 2822 7368 2830
rect 7375 2828 7485 2836
rect 7338 2814 7383 2822
rect 7070 2796 7089 2798
rect 7104 2796 7150 2798
rect 7070 2780 7150 2796
rect 7177 2794 7212 2807
rect 7253 2804 7290 2807
rect 7253 2802 7295 2804
rect 7182 2791 7212 2794
rect 7191 2787 7198 2791
rect 7198 2786 7199 2787
rect 7157 2780 7167 2786
rect 6916 2772 6951 2780
rect 6916 2746 6917 2772
rect 6924 2746 6951 2772
rect 6859 2728 6889 2742
rect 6916 2738 6951 2746
rect 6953 2772 6994 2780
rect 6953 2746 6968 2772
rect 6975 2746 6994 2772
rect 7058 2768 7089 2780
rect 7104 2768 7207 2780
rect 7219 2770 7245 2796
rect 7260 2791 7290 2802
rect 7322 2798 7384 2814
rect 7322 2796 7368 2798
rect 7322 2780 7384 2796
rect 7396 2780 7402 2828
rect 7405 2820 7485 2828
rect 7405 2818 7424 2820
rect 7439 2818 7473 2820
rect 7405 2802 7485 2818
rect 7405 2780 7424 2802
rect 7439 2786 7469 2802
rect 7497 2796 7503 2870
rect 7506 2796 7525 2940
rect 7540 2796 7546 2940
rect 7555 2870 7568 2940
rect 7620 2936 7642 2940
rect 7613 2914 7642 2928
rect 7695 2914 7711 2928
rect 7749 2924 7755 2926
rect 7762 2924 7870 2940
rect 7877 2924 7883 2926
rect 7891 2924 7906 2940
rect 7972 2934 7991 2937
rect 7613 2912 7711 2914
rect 7738 2912 7906 2924
rect 7921 2914 7937 2928
rect 7972 2915 7994 2934
rect 8004 2928 8020 2929
rect 8003 2926 8020 2928
rect 8004 2921 8020 2926
rect 7994 2914 8000 2915
rect 8003 2914 8032 2921
rect 7921 2913 8032 2914
rect 7921 2912 8038 2913
rect 7597 2904 7648 2912
rect 7695 2904 7729 2912
rect 7597 2892 7622 2904
rect 7629 2892 7648 2904
rect 7702 2902 7729 2904
rect 7738 2902 7959 2912
rect 7994 2909 8000 2912
rect 7702 2898 7959 2902
rect 7597 2884 7648 2892
rect 7695 2884 7959 2898
rect 8003 2904 8038 2912
rect 7549 2836 7568 2870
rect 7613 2876 7642 2884
rect 7613 2870 7630 2876
rect 7613 2868 7647 2870
rect 7695 2868 7711 2884
rect 7712 2874 7920 2884
rect 7921 2874 7937 2884
rect 7985 2880 8000 2895
rect 8003 2892 8004 2904
rect 8011 2892 8038 2904
rect 8003 2884 8038 2892
rect 8003 2883 8032 2884
rect 7723 2870 7937 2874
rect 7738 2868 7937 2870
rect 7972 2870 7985 2880
rect 8003 2870 8020 2883
rect 7972 2868 8020 2870
rect 7614 2864 7647 2868
rect 7610 2862 7647 2864
rect 7610 2861 7677 2862
rect 7610 2856 7641 2861
rect 7647 2856 7677 2861
rect 7610 2852 7677 2856
rect 7583 2849 7677 2852
rect 7583 2842 7632 2849
rect 7583 2836 7613 2842
rect 7632 2837 7637 2842
rect 7549 2820 7629 2836
rect 7641 2828 7677 2849
rect 7738 2844 7927 2868
rect 7972 2867 8019 2868
rect 7985 2862 8019 2867
rect 7753 2841 7927 2844
rect 7746 2838 7927 2841
rect 7955 2861 8019 2862
rect 7549 2818 7568 2820
rect 7583 2818 7617 2820
rect 7549 2802 7629 2818
rect 7549 2796 7568 2802
rect 7265 2770 7368 2780
rect 7219 2768 7368 2770
rect 7389 2768 7424 2780
rect 7058 2766 7220 2768
rect 7070 2746 7089 2766
rect 7104 2764 7134 2766
rect 6953 2738 6994 2746
rect 7076 2742 7089 2746
rect 7141 2750 7220 2766
rect 7252 2766 7424 2768
rect 7252 2750 7331 2766
rect 7338 2764 7368 2766
rect 6916 2728 6945 2738
rect 6959 2728 6988 2738
rect 7003 2728 7033 2742
rect 7076 2728 7119 2742
rect 7141 2738 7331 2750
rect 7396 2746 7402 2766
rect 7126 2728 7156 2738
rect 7157 2728 7315 2738
rect 7319 2728 7349 2738
rect 7353 2728 7383 2742
rect 7411 2728 7424 2766
rect 7496 2780 7525 2796
rect 7539 2780 7568 2796
rect 7583 2786 7613 2802
rect 7641 2780 7647 2828
rect 7650 2822 7669 2828
rect 7684 2822 7714 2830
rect 7650 2814 7714 2822
rect 7650 2798 7730 2814
rect 7746 2807 7808 2838
rect 7824 2807 7886 2838
rect 7955 2836 8004 2861
rect 8019 2836 8049 2852
rect 7918 2822 7948 2830
rect 7955 2828 8065 2836
rect 7918 2814 7963 2822
rect 7650 2796 7669 2798
rect 7684 2796 7730 2798
rect 7650 2780 7730 2796
rect 7757 2794 7792 2807
rect 7833 2804 7870 2807
rect 7833 2802 7875 2804
rect 7762 2791 7792 2794
rect 7771 2787 7778 2791
rect 7778 2786 7779 2787
rect 7737 2780 7747 2786
rect 7496 2772 7531 2780
rect 7496 2746 7497 2772
rect 7504 2746 7531 2772
rect 7439 2728 7469 2742
rect 7496 2738 7531 2746
rect 7533 2772 7574 2780
rect 7533 2746 7548 2772
rect 7555 2746 7574 2772
rect 7638 2768 7669 2780
rect 7684 2768 7787 2780
rect 7799 2770 7825 2796
rect 7840 2791 7870 2802
rect 7902 2798 7964 2814
rect 7902 2796 7948 2798
rect 7902 2780 7964 2796
rect 7976 2780 7982 2828
rect 7985 2820 8065 2828
rect 7985 2818 8004 2820
rect 8019 2818 8053 2820
rect 7985 2802 8065 2818
rect 7985 2780 8004 2802
rect 8019 2786 8049 2802
rect 8077 2796 8083 2870
rect 8086 2796 8105 2940
rect 8120 2796 8126 2940
rect 8135 2870 8148 2940
rect 8200 2936 8222 2940
rect 8193 2914 8222 2928
rect 8275 2914 8291 2928
rect 8329 2924 8335 2926
rect 8342 2924 8450 2940
rect 8457 2924 8463 2926
rect 8471 2924 8486 2940
rect 8552 2934 8571 2937
rect 8193 2912 8291 2914
rect 8318 2912 8486 2924
rect 8501 2914 8517 2928
rect 8552 2915 8574 2934
rect 8584 2928 8600 2929
rect 8583 2926 8600 2928
rect 8584 2921 8600 2926
rect 8574 2914 8580 2915
rect 8583 2914 8612 2921
rect 8501 2913 8612 2914
rect 8501 2912 8618 2913
rect 8177 2904 8228 2912
rect 8275 2904 8309 2912
rect 8177 2892 8202 2904
rect 8209 2892 8228 2904
rect 8282 2902 8309 2904
rect 8318 2902 8539 2912
rect 8574 2909 8580 2912
rect 8282 2898 8539 2902
rect 8177 2884 8228 2892
rect 8275 2884 8539 2898
rect 8583 2904 8618 2912
rect 8129 2836 8148 2870
rect 8193 2876 8222 2884
rect 8193 2870 8210 2876
rect 8193 2868 8227 2870
rect 8275 2868 8291 2884
rect 8292 2874 8500 2884
rect 8501 2874 8517 2884
rect 8565 2880 8580 2895
rect 8583 2892 8584 2904
rect 8591 2892 8618 2904
rect 8583 2884 8618 2892
rect 8583 2883 8612 2884
rect 8303 2870 8517 2874
rect 8318 2868 8517 2870
rect 8552 2870 8565 2880
rect 8583 2870 8600 2883
rect 8552 2868 8600 2870
rect 8194 2864 8227 2868
rect 8190 2862 8227 2864
rect 8190 2861 8257 2862
rect 8190 2856 8221 2861
rect 8227 2856 8257 2861
rect 8190 2852 8257 2856
rect 8163 2849 8257 2852
rect 8163 2842 8212 2849
rect 8163 2836 8193 2842
rect 8212 2837 8217 2842
rect 8129 2820 8209 2836
rect 8221 2828 8257 2849
rect 8318 2844 8507 2868
rect 8552 2867 8599 2868
rect 8565 2862 8599 2867
rect 8333 2841 8507 2844
rect 8326 2838 8507 2841
rect 8535 2861 8599 2862
rect 8129 2818 8148 2820
rect 8163 2818 8197 2820
rect 8129 2802 8209 2818
rect 8129 2796 8148 2802
rect 7845 2770 7948 2780
rect 7799 2768 7948 2770
rect 7969 2768 8004 2780
rect 7638 2766 7800 2768
rect 7650 2746 7669 2766
rect 7684 2764 7714 2766
rect 7533 2738 7574 2746
rect 7656 2742 7669 2746
rect 7721 2750 7800 2766
rect 7832 2766 8004 2768
rect 7832 2750 7911 2766
rect 7918 2764 7948 2766
rect 7496 2728 7525 2738
rect 7539 2728 7568 2738
rect 7583 2728 7613 2742
rect 7656 2728 7699 2742
rect 7721 2738 7911 2750
rect 7976 2746 7982 2766
rect 7706 2728 7736 2738
rect 7737 2728 7895 2738
rect 7899 2728 7929 2738
rect 7933 2728 7963 2742
rect 7991 2728 8004 2766
rect 8076 2780 8105 2796
rect 8119 2780 8148 2796
rect 8163 2786 8193 2802
rect 8221 2780 8227 2828
rect 8230 2822 8249 2828
rect 8264 2822 8294 2830
rect 8230 2814 8294 2822
rect 8230 2798 8310 2814
rect 8326 2807 8388 2838
rect 8404 2807 8466 2838
rect 8535 2836 8584 2861
rect 8599 2836 8629 2852
rect 8498 2822 8528 2830
rect 8535 2828 8645 2836
rect 8498 2814 8543 2822
rect 8230 2796 8249 2798
rect 8264 2796 8310 2798
rect 8230 2780 8310 2796
rect 8337 2794 8372 2807
rect 8413 2804 8450 2807
rect 8413 2802 8455 2804
rect 8342 2791 8372 2794
rect 8351 2787 8358 2791
rect 8358 2786 8359 2787
rect 8317 2780 8327 2786
rect 8076 2772 8111 2780
rect 8076 2746 8077 2772
rect 8084 2746 8111 2772
rect 8019 2728 8049 2742
rect 8076 2738 8111 2746
rect 8113 2772 8154 2780
rect 8113 2746 8128 2772
rect 8135 2746 8154 2772
rect 8218 2768 8249 2780
rect 8264 2768 8367 2780
rect 8379 2770 8405 2796
rect 8420 2791 8450 2802
rect 8482 2798 8544 2814
rect 8482 2796 8528 2798
rect 8482 2780 8544 2796
rect 8556 2780 8562 2828
rect 8565 2820 8645 2828
rect 8565 2818 8584 2820
rect 8599 2818 8633 2820
rect 8565 2802 8645 2818
rect 8565 2780 8584 2802
rect 8599 2786 8629 2802
rect 8657 2796 8663 2870
rect 8666 2796 8685 2940
rect 8700 2796 8706 2940
rect 8715 2870 8728 2940
rect 8780 2936 8802 2940
rect 8773 2914 8802 2928
rect 8855 2914 8871 2928
rect 8909 2924 8915 2926
rect 8922 2924 9030 2940
rect 9037 2924 9043 2926
rect 9051 2924 9066 2940
rect 9132 2934 9151 2937
rect 8773 2912 8871 2914
rect 8898 2912 9066 2924
rect 9081 2914 9097 2928
rect 9132 2915 9154 2934
rect 9164 2928 9180 2929
rect 9163 2926 9180 2928
rect 9164 2921 9180 2926
rect 9154 2914 9160 2915
rect 9163 2914 9192 2921
rect 9081 2913 9192 2914
rect 9081 2912 9198 2913
rect 8757 2904 8808 2912
rect 8855 2904 8889 2912
rect 8757 2892 8782 2904
rect 8789 2892 8808 2904
rect 8862 2902 8889 2904
rect 8898 2902 9119 2912
rect 9154 2909 9160 2912
rect 8862 2898 9119 2902
rect 8757 2884 8808 2892
rect 8855 2884 9119 2898
rect 9163 2904 9198 2912
rect 8709 2836 8728 2870
rect 8773 2876 8802 2884
rect 8773 2870 8790 2876
rect 8773 2868 8807 2870
rect 8855 2868 8871 2884
rect 8872 2874 9080 2884
rect 9081 2874 9097 2884
rect 9145 2880 9160 2895
rect 9163 2892 9164 2904
rect 9171 2892 9198 2904
rect 9163 2884 9198 2892
rect 9163 2883 9192 2884
rect 8883 2870 9097 2874
rect 8898 2868 9097 2870
rect 9132 2870 9145 2880
rect 9163 2870 9180 2883
rect 9132 2868 9180 2870
rect 8774 2864 8807 2868
rect 8770 2862 8807 2864
rect 8770 2861 8837 2862
rect 8770 2856 8801 2861
rect 8807 2856 8837 2861
rect 8770 2852 8837 2856
rect 8743 2849 8837 2852
rect 8743 2842 8792 2849
rect 8743 2836 8773 2842
rect 8792 2837 8797 2842
rect 8709 2820 8789 2836
rect 8801 2828 8837 2849
rect 8898 2844 9087 2868
rect 9132 2867 9179 2868
rect 9145 2862 9179 2867
rect 8913 2841 9087 2844
rect 8906 2838 9087 2841
rect 9115 2861 9179 2862
rect 8709 2818 8728 2820
rect 8743 2818 8777 2820
rect 8709 2802 8789 2818
rect 8709 2796 8728 2802
rect 8425 2770 8528 2780
rect 8379 2768 8528 2770
rect 8549 2768 8584 2780
rect 8218 2766 8380 2768
rect 8230 2746 8249 2766
rect 8264 2764 8294 2766
rect 8113 2738 8154 2746
rect 8236 2742 8249 2746
rect 8301 2750 8380 2766
rect 8412 2766 8584 2768
rect 8412 2750 8491 2766
rect 8498 2764 8528 2766
rect 8076 2728 8105 2738
rect 8119 2728 8148 2738
rect 8163 2728 8193 2742
rect 8236 2728 8279 2742
rect 8301 2738 8491 2750
rect 8556 2746 8562 2766
rect 8286 2728 8316 2738
rect 8317 2728 8475 2738
rect 8479 2728 8509 2738
rect 8513 2728 8543 2742
rect 8571 2728 8584 2766
rect 8656 2780 8685 2796
rect 8699 2780 8728 2796
rect 8743 2786 8773 2802
rect 8801 2780 8807 2828
rect 8810 2822 8829 2828
rect 8844 2822 8874 2830
rect 8810 2814 8874 2822
rect 8810 2798 8890 2814
rect 8906 2807 8968 2838
rect 8984 2807 9046 2838
rect 9115 2836 9164 2861
rect 9179 2836 9209 2852
rect 9078 2822 9108 2830
rect 9115 2828 9225 2836
rect 9078 2814 9123 2822
rect 8810 2796 8829 2798
rect 8844 2796 8890 2798
rect 8810 2780 8890 2796
rect 8917 2794 8952 2807
rect 8993 2804 9030 2807
rect 8993 2802 9035 2804
rect 8922 2791 8952 2794
rect 8931 2787 8938 2791
rect 8938 2786 8939 2787
rect 8897 2780 8907 2786
rect 8656 2772 8691 2780
rect 8656 2746 8657 2772
rect 8664 2746 8691 2772
rect 8599 2728 8629 2742
rect 8656 2738 8691 2746
rect 8693 2772 8734 2780
rect 8693 2746 8708 2772
rect 8715 2746 8734 2772
rect 8798 2768 8829 2780
rect 8844 2768 8947 2780
rect 8959 2770 8985 2796
rect 9000 2791 9030 2802
rect 9062 2798 9124 2814
rect 9062 2796 9108 2798
rect 9062 2780 9124 2796
rect 9136 2780 9142 2828
rect 9145 2820 9225 2828
rect 9145 2818 9164 2820
rect 9179 2818 9213 2820
rect 9145 2802 9225 2818
rect 9145 2780 9164 2802
rect 9179 2786 9209 2802
rect 9237 2796 9243 2870
rect 9252 2796 9265 2940
rect 9005 2770 9108 2780
rect 8959 2768 9108 2770
rect 9129 2768 9164 2780
rect 8798 2766 8960 2768
rect 8810 2746 8829 2766
rect 8844 2764 8874 2766
rect 8693 2738 8734 2746
rect 8816 2742 8829 2746
rect 8881 2750 8960 2766
rect 8992 2766 9164 2768
rect 8992 2750 9071 2766
rect 9078 2764 9108 2766
rect 8656 2728 8685 2738
rect 8699 2728 8728 2738
rect 8743 2728 8773 2742
rect 8816 2728 8859 2742
rect 8881 2738 9071 2750
rect 9136 2746 9142 2766
rect 8866 2728 8896 2738
rect 8897 2728 9055 2738
rect 9059 2728 9089 2738
rect 9093 2728 9123 2742
rect 9151 2728 9164 2766
rect 9236 2780 9265 2796
rect 9236 2772 9271 2780
rect 9236 2746 9237 2772
rect 9244 2746 9271 2772
rect 9179 2728 9209 2742
rect 9236 2738 9271 2746
rect 9236 2728 9265 2738
rect -1 2722 9265 2728
rect 0 2714 9265 2722
rect 15 2684 28 2714
rect 43 2700 73 2714
rect 116 2700 159 2714
rect 166 2700 386 2714
rect 393 2700 423 2714
rect 83 2686 98 2698
rect 117 2686 130 2700
rect 198 2696 351 2700
rect 80 2684 102 2686
rect 180 2684 372 2696
rect 451 2684 464 2714
rect 479 2700 509 2714
rect 546 2684 565 2714
rect 580 2684 586 2714
rect 595 2684 608 2714
rect 623 2700 653 2714
rect 696 2700 739 2714
rect 746 2700 966 2714
rect 973 2700 1003 2714
rect 663 2686 678 2698
rect 697 2686 710 2700
rect 778 2696 931 2700
rect 660 2684 682 2686
rect 760 2684 952 2696
rect 1031 2684 1044 2714
rect 1059 2700 1089 2714
rect 1126 2684 1145 2714
rect 1160 2684 1166 2714
rect 1175 2684 1188 2714
rect 1203 2700 1233 2714
rect 1276 2700 1319 2714
rect 1326 2700 1546 2714
rect 1553 2700 1583 2714
rect 1243 2686 1258 2698
rect 1277 2686 1290 2700
rect 1358 2696 1511 2700
rect 1240 2684 1262 2686
rect 1340 2684 1532 2696
rect 1611 2684 1624 2714
rect 1639 2700 1669 2714
rect 1706 2684 1725 2714
rect 1740 2684 1746 2714
rect 1755 2684 1768 2714
rect 1783 2700 1813 2714
rect 1856 2700 1899 2714
rect 1906 2700 2126 2714
rect 2133 2700 2163 2714
rect 1823 2686 1838 2698
rect 1857 2686 1870 2700
rect 1938 2696 2091 2700
rect 1820 2684 1842 2686
rect 1920 2684 2112 2696
rect 2191 2684 2204 2714
rect 2219 2700 2249 2714
rect 2286 2684 2305 2714
rect 2320 2684 2326 2714
rect 2335 2684 2348 2714
rect 2363 2700 2393 2714
rect 2436 2700 2479 2714
rect 2486 2700 2706 2714
rect 2713 2700 2743 2714
rect 2403 2686 2418 2698
rect 2437 2686 2450 2700
rect 2518 2696 2671 2700
rect 2400 2684 2422 2686
rect 2500 2684 2692 2696
rect 2771 2684 2784 2714
rect 2799 2700 2829 2714
rect 2866 2684 2885 2714
rect 2900 2684 2906 2714
rect 2915 2684 2928 2714
rect 2943 2700 2973 2714
rect 3016 2700 3059 2714
rect 3066 2700 3286 2714
rect 3293 2700 3323 2714
rect 2983 2686 2998 2698
rect 3017 2686 3030 2700
rect 3098 2696 3251 2700
rect 2980 2684 3002 2686
rect 3080 2684 3272 2696
rect 3351 2684 3364 2714
rect 3379 2700 3409 2714
rect 3446 2684 3465 2714
rect 3480 2684 3486 2714
rect 3495 2684 3508 2714
rect 3523 2700 3553 2714
rect 3596 2700 3639 2714
rect 3646 2700 3866 2714
rect 3873 2700 3903 2714
rect 3563 2686 3578 2698
rect 3597 2686 3610 2700
rect 3678 2696 3831 2700
rect 3560 2684 3582 2686
rect 3660 2684 3852 2696
rect 3931 2684 3944 2714
rect 3959 2700 3989 2714
rect 4026 2684 4045 2714
rect 4060 2684 4066 2714
rect 4075 2684 4088 2714
rect 4103 2700 4133 2714
rect 4176 2700 4219 2714
rect 4226 2700 4446 2714
rect 4453 2700 4483 2714
rect 4143 2686 4158 2698
rect 4177 2686 4190 2700
rect 4258 2696 4411 2700
rect 4140 2684 4162 2686
rect 4240 2684 4432 2696
rect 4511 2684 4524 2714
rect 4539 2700 4569 2714
rect 4606 2684 4625 2714
rect 4640 2684 4646 2714
rect 4655 2684 4668 2714
rect 4683 2700 4713 2714
rect 4756 2700 4799 2714
rect 4806 2700 5026 2714
rect 5033 2700 5063 2714
rect 4723 2686 4738 2698
rect 4757 2686 4770 2700
rect 4838 2696 4991 2700
rect 4720 2684 4742 2686
rect 4820 2684 5012 2696
rect 5091 2684 5104 2714
rect 5119 2700 5149 2714
rect 5186 2684 5205 2714
rect 5220 2684 5226 2714
rect 5235 2684 5248 2714
rect 5263 2700 5293 2714
rect 5336 2700 5379 2714
rect 5386 2700 5606 2714
rect 5613 2700 5643 2714
rect 5303 2686 5318 2698
rect 5337 2686 5350 2700
rect 5418 2696 5571 2700
rect 5300 2684 5322 2686
rect 5400 2684 5592 2696
rect 5671 2684 5684 2714
rect 5699 2700 5729 2714
rect 5766 2684 5785 2714
rect 5800 2684 5806 2714
rect 5815 2684 5828 2714
rect 5843 2700 5873 2714
rect 5916 2700 5959 2714
rect 5966 2700 6186 2714
rect 6193 2700 6223 2714
rect 5883 2686 5898 2698
rect 5917 2686 5930 2700
rect 5998 2696 6151 2700
rect 5880 2684 5902 2686
rect 5980 2684 6172 2696
rect 6251 2684 6264 2714
rect 6279 2700 6309 2714
rect 6346 2684 6365 2714
rect 6380 2684 6386 2714
rect 6395 2684 6408 2714
rect 6423 2700 6453 2714
rect 6496 2700 6539 2714
rect 6546 2700 6766 2714
rect 6773 2700 6803 2714
rect 6463 2686 6478 2698
rect 6497 2686 6510 2700
rect 6578 2696 6731 2700
rect 6460 2684 6482 2686
rect 6560 2684 6752 2696
rect 6831 2684 6844 2714
rect 6859 2700 6889 2714
rect 6926 2684 6945 2714
rect 6960 2684 6966 2714
rect 6975 2684 6988 2714
rect 7003 2700 7033 2714
rect 7076 2700 7119 2714
rect 7126 2700 7346 2714
rect 7353 2700 7383 2714
rect 7043 2686 7058 2698
rect 7077 2686 7090 2700
rect 7158 2696 7311 2700
rect 7040 2684 7062 2686
rect 7140 2684 7332 2696
rect 7411 2684 7424 2714
rect 7439 2700 7469 2714
rect 7506 2684 7525 2714
rect 7540 2684 7546 2714
rect 7555 2684 7568 2714
rect 7583 2700 7613 2714
rect 7656 2700 7699 2714
rect 7706 2700 7926 2714
rect 7933 2700 7963 2714
rect 7623 2686 7638 2698
rect 7657 2686 7670 2700
rect 7738 2696 7891 2700
rect 7620 2684 7642 2686
rect 7720 2684 7912 2696
rect 7991 2684 8004 2714
rect 8019 2700 8049 2714
rect 8086 2684 8105 2714
rect 8120 2684 8126 2714
rect 8135 2684 8148 2714
rect 8163 2700 8193 2714
rect 8236 2700 8279 2714
rect 8286 2700 8506 2714
rect 8513 2700 8543 2714
rect 8203 2686 8218 2698
rect 8237 2686 8250 2700
rect 8318 2696 8471 2700
rect 8200 2684 8222 2686
rect 8300 2684 8492 2696
rect 8571 2684 8584 2714
rect 8599 2700 8629 2714
rect 8666 2684 8685 2714
rect 8700 2684 8706 2714
rect 8715 2684 8728 2714
rect 8743 2700 8773 2714
rect 8816 2700 8859 2714
rect 8866 2700 9086 2714
rect 9093 2700 9123 2714
rect 8783 2686 8798 2698
rect 8817 2686 8830 2700
rect 8898 2696 9051 2700
rect 8780 2684 8802 2686
rect 8880 2684 9072 2696
rect 9151 2684 9164 2714
rect 9179 2700 9209 2714
rect 9252 2684 9265 2714
rect 0 2670 9265 2684
rect 15 2600 28 2670
rect 80 2666 102 2670
rect 73 2644 102 2658
rect 155 2644 171 2658
rect 209 2654 215 2656
rect 222 2654 330 2670
rect 337 2654 343 2656
rect 351 2654 366 2670
rect 432 2664 451 2667
rect 73 2642 171 2644
rect 198 2642 366 2654
rect 381 2644 397 2658
rect 432 2645 454 2664
rect 464 2658 480 2659
rect 463 2656 480 2658
rect 464 2651 480 2656
rect 454 2644 460 2645
rect 463 2644 492 2651
rect 381 2643 492 2644
rect 381 2642 498 2643
rect 57 2634 108 2642
rect 155 2634 189 2642
rect 57 2622 82 2634
rect 89 2622 108 2634
rect 162 2632 189 2634
rect 198 2632 419 2642
rect 454 2639 460 2642
rect 162 2628 419 2632
rect 57 2614 108 2622
rect 155 2614 419 2628
rect 463 2634 498 2642
rect 9 2566 28 2600
rect 73 2606 102 2614
rect 73 2600 90 2606
rect 73 2598 107 2600
rect 155 2598 171 2614
rect 172 2604 380 2614
rect 381 2604 397 2614
rect 445 2610 460 2625
rect 463 2622 464 2634
rect 471 2622 498 2634
rect 463 2614 498 2622
rect 463 2613 492 2614
rect 183 2600 397 2604
rect 198 2598 397 2600
rect 432 2600 445 2610
rect 463 2600 480 2613
rect 432 2598 480 2600
rect 74 2594 107 2598
rect 70 2592 107 2594
rect 70 2591 137 2592
rect 70 2586 101 2591
rect 107 2586 137 2591
rect 70 2582 137 2586
rect 43 2579 137 2582
rect 43 2572 92 2579
rect 43 2566 73 2572
rect 92 2567 97 2572
rect 9 2550 89 2566
rect 101 2558 137 2579
rect 198 2574 387 2598
rect 432 2597 479 2598
rect 445 2592 479 2597
rect 213 2571 387 2574
rect 206 2568 387 2571
rect 415 2591 479 2592
rect 9 2548 28 2550
rect 43 2548 77 2550
rect 9 2532 89 2548
rect 9 2526 28 2532
rect -1 2510 28 2526
rect 43 2516 73 2532
rect 101 2510 107 2558
rect 110 2552 129 2558
rect 144 2552 174 2560
rect 110 2544 174 2552
rect 110 2528 190 2544
rect 206 2537 268 2568
rect 284 2537 346 2568
rect 415 2566 464 2591
rect 479 2566 509 2582
rect 378 2552 408 2560
rect 415 2558 525 2566
rect 378 2544 423 2552
rect 110 2526 129 2528
rect 144 2526 190 2528
rect 110 2510 190 2526
rect 217 2524 252 2537
rect 293 2534 330 2537
rect 293 2532 335 2534
rect 222 2521 252 2524
rect 231 2517 238 2521
rect 238 2516 239 2517
rect 197 2510 207 2516
rect -7 2502 34 2510
rect -7 2476 8 2502
rect 15 2476 34 2502
rect 98 2498 129 2510
rect 144 2498 247 2510
rect 259 2500 285 2526
rect 300 2521 330 2532
rect 362 2528 424 2544
rect 362 2526 408 2528
rect 362 2510 424 2526
rect 436 2510 442 2558
rect 445 2550 525 2558
rect 445 2548 464 2550
rect 479 2548 513 2550
rect 445 2532 525 2548
rect 445 2510 464 2532
rect 479 2516 509 2532
rect 537 2526 543 2600
rect 546 2526 565 2670
rect 580 2526 586 2670
rect 595 2600 608 2670
rect 660 2666 682 2670
rect 653 2644 682 2658
rect 735 2644 751 2658
rect 789 2654 795 2656
rect 802 2654 910 2670
rect 917 2654 923 2656
rect 931 2654 946 2670
rect 1012 2664 1031 2667
rect 653 2642 751 2644
rect 778 2642 946 2654
rect 961 2644 977 2658
rect 1012 2645 1034 2664
rect 1044 2658 1060 2659
rect 1043 2656 1060 2658
rect 1044 2651 1060 2656
rect 1034 2644 1040 2645
rect 1043 2644 1072 2651
rect 961 2643 1072 2644
rect 961 2642 1078 2643
rect 637 2634 688 2642
rect 735 2634 769 2642
rect 637 2622 662 2634
rect 669 2622 688 2634
rect 742 2632 769 2634
rect 778 2632 999 2642
rect 1034 2639 1040 2642
rect 742 2628 999 2632
rect 637 2614 688 2622
rect 735 2614 999 2628
rect 1043 2634 1078 2642
rect 589 2566 608 2600
rect 653 2606 682 2614
rect 653 2600 670 2606
rect 653 2598 687 2600
rect 735 2598 751 2614
rect 752 2604 960 2614
rect 961 2604 977 2614
rect 1025 2610 1040 2625
rect 1043 2622 1044 2634
rect 1051 2622 1078 2634
rect 1043 2614 1078 2622
rect 1043 2613 1072 2614
rect 763 2600 977 2604
rect 778 2598 977 2600
rect 1012 2600 1025 2610
rect 1043 2600 1060 2613
rect 1012 2598 1060 2600
rect 654 2594 687 2598
rect 650 2592 687 2594
rect 650 2591 717 2592
rect 650 2586 681 2591
rect 687 2586 717 2591
rect 650 2582 717 2586
rect 623 2579 717 2582
rect 623 2572 672 2579
rect 623 2566 653 2572
rect 672 2567 677 2572
rect 589 2550 669 2566
rect 681 2558 717 2579
rect 778 2574 967 2598
rect 1012 2597 1059 2598
rect 1025 2592 1059 2597
rect 793 2571 967 2574
rect 786 2568 967 2571
rect 995 2591 1059 2592
rect 589 2548 608 2550
rect 623 2548 657 2550
rect 589 2532 669 2548
rect 589 2526 608 2532
rect 305 2500 408 2510
rect 259 2498 408 2500
rect 429 2498 464 2510
rect 98 2496 260 2498
rect 110 2476 129 2496
rect 144 2494 174 2496
rect -7 2468 34 2476
rect 116 2472 129 2476
rect 181 2480 260 2496
rect 292 2496 464 2498
rect 292 2480 371 2496
rect 378 2494 408 2496
rect -1 2458 28 2468
rect 43 2458 73 2472
rect 116 2458 159 2472
rect 181 2468 371 2480
rect 436 2476 442 2496
rect 166 2458 196 2468
rect 197 2458 355 2468
rect 359 2458 389 2468
rect 393 2458 423 2472
rect 451 2458 464 2496
rect 536 2510 565 2526
rect 579 2510 608 2526
rect 623 2516 653 2532
rect 681 2510 687 2558
rect 690 2552 709 2558
rect 724 2552 754 2560
rect 690 2544 754 2552
rect 690 2528 770 2544
rect 786 2537 848 2568
rect 864 2537 926 2568
rect 995 2566 1044 2591
rect 1059 2566 1089 2582
rect 958 2552 988 2560
rect 995 2558 1105 2566
rect 958 2544 1003 2552
rect 690 2526 709 2528
rect 724 2526 770 2528
rect 690 2510 770 2526
rect 797 2524 832 2537
rect 873 2534 910 2537
rect 873 2532 915 2534
rect 802 2521 832 2524
rect 811 2517 818 2521
rect 818 2516 819 2517
rect 777 2510 787 2516
rect 536 2502 571 2510
rect 536 2476 537 2502
rect 544 2476 571 2502
rect 479 2458 509 2472
rect 536 2468 571 2476
rect 573 2502 614 2510
rect 573 2476 588 2502
rect 595 2476 614 2502
rect 678 2498 709 2510
rect 724 2498 827 2510
rect 839 2500 865 2526
rect 880 2521 910 2532
rect 942 2528 1004 2544
rect 942 2526 988 2528
rect 942 2510 1004 2526
rect 1016 2510 1022 2558
rect 1025 2550 1105 2558
rect 1025 2548 1044 2550
rect 1059 2548 1093 2550
rect 1025 2532 1105 2548
rect 1025 2510 1044 2532
rect 1059 2516 1089 2532
rect 1117 2526 1123 2600
rect 1126 2526 1145 2670
rect 1160 2526 1166 2670
rect 1175 2600 1188 2670
rect 1240 2666 1262 2670
rect 1233 2644 1262 2658
rect 1315 2644 1331 2658
rect 1369 2654 1375 2656
rect 1382 2654 1490 2670
rect 1497 2654 1503 2656
rect 1511 2654 1526 2670
rect 1592 2664 1611 2667
rect 1233 2642 1331 2644
rect 1358 2642 1526 2654
rect 1541 2644 1557 2658
rect 1592 2645 1614 2664
rect 1624 2658 1640 2659
rect 1623 2656 1640 2658
rect 1624 2651 1640 2656
rect 1614 2644 1620 2645
rect 1623 2644 1652 2651
rect 1541 2643 1652 2644
rect 1541 2642 1658 2643
rect 1217 2634 1268 2642
rect 1315 2634 1349 2642
rect 1217 2622 1242 2634
rect 1249 2622 1268 2634
rect 1322 2632 1349 2634
rect 1358 2632 1579 2642
rect 1614 2639 1620 2642
rect 1322 2628 1579 2632
rect 1217 2614 1268 2622
rect 1315 2614 1579 2628
rect 1623 2634 1658 2642
rect 1169 2566 1188 2600
rect 1233 2606 1262 2614
rect 1233 2600 1250 2606
rect 1233 2598 1267 2600
rect 1315 2598 1331 2614
rect 1332 2604 1540 2614
rect 1541 2604 1557 2614
rect 1605 2610 1620 2625
rect 1623 2622 1624 2634
rect 1631 2622 1658 2634
rect 1623 2614 1658 2622
rect 1623 2613 1652 2614
rect 1343 2600 1557 2604
rect 1358 2598 1557 2600
rect 1592 2600 1605 2610
rect 1623 2600 1640 2613
rect 1592 2598 1640 2600
rect 1234 2594 1267 2598
rect 1230 2592 1267 2594
rect 1230 2591 1297 2592
rect 1230 2586 1261 2591
rect 1267 2586 1297 2591
rect 1230 2582 1297 2586
rect 1203 2579 1297 2582
rect 1203 2572 1252 2579
rect 1203 2566 1233 2572
rect 1252 2567 1257 2572
rect 1169 2550 1249 2566
rect 1261 2558 1297 2579
rect 1358 2574 1547 2598
rect 1592 2597 1639 2598
rect 1605 2592 1639 2597
rect 1373 2571 1547 2574
rect 1366 2568 1547 2571
rect 1575 2591 1639 2592
rect 1169 2548 1188 2550
rect 1203 2548 1237 2550
rect 1169 2532 1249 2548
rect 1169 2526 1188 2532
rect 885 2500 988 2510
rect 839 2498 988 2500
rect 1009 2498 1044 2510
rect 678 2496 840 2498
rect 690 2476 709 2496
rect 724 2494 754 2496
rect 573 2468 614 2476
rect 696 2472 709 2476
rect 761 2480 840 2496
rect 872 2496 1044 2498
rect 872 2480 951 2496
rect 958 2494 988 2496
rect 536 2458 565 2468
rect 579 2458 608 2468
rect 623 2458 653 2472
rect 696 2458 739 2472
rect 761 2468 951 2480
rect 1016 2476 1022 2496
rect 746 2458 776 2468
rect 777 2458 935 2468
rect 939 2458 969 2468
rect 973 2458 1003 2472
rect 1031 2458 1044 2496
rect 1116 2510 1145 2526
rect 1159 2510 1188 2526
rect 1203 2516 1233 2532
rect 1261 2510 1267 2558
rect 1270 2552 1289 2558
rect 1304 2552 1334 2560
rect 1270 2544 1334 2552
rect 1270 2528 1350 2544
rect 1366 2537 1428 2568
rect 1444 2537 1506 2568
rect 1575 2566 1624 2591
rect 1639 2566 1669 2582
rect 1538 2552 1568 2560
rect 1575 2558 1685 2566
rect 1538 2544 1583 2552
rect 1270 2526 1289 2528
rect 1304 2526 1350 2528
rect 1270 2510 1350 2526
rect 1377 2524 1412 2537
rect 1453 2534 1490 2537
rect 1453 2532 1495 2534
rect 1382 2521 1412 2524
rect 1391 2517 1398 2521
rect 1398 2516 1399 2517
rect 1357 2510 1367 2516
rect 1116 2502 1151 2510
rect 1116 2476 1117 2502
rect 1124 2476 1151 2502
rect 1059 2458 1089 2472
rect 1116 2468 1151 2476
rect 1153 2502 1194 2510
rect 1153 2476 1168 2502
rect 1175 2476 1194 2502
rect 1258 2498 1289 2510
rect 1304 2498 1407 2510
rect 1419 2500 1445 2526
rect 1460 2521 1490 2532
rect 1522 2528 1584 2544
rect 1522 2526 1568 2528
rect 1522 2510 1584 2526
rect 1596 2510 1602 2558
rect 1605 2550 1685 2558
rect 1605 2548 1624 2550
rect 1639 2548 1673 2550
rect 1605 2532 1685 2548
rect 1605 2510 1624 2532
rect 1639 2516 1669 2532
rect 1697 2526 1703 2600
rect 1706 2526 1725 2670
rect 1740 2526 1746 2670
rect 1755 2600 1768 2670
rect 1820 2666 1842 2670
rect 1813 2644 1842 2658
rect 1895 2644 1911 2658
rect 1949 2654 1955 2656
rect 1962 2654 2070 2670
rect 2077 2654 2083 2656
rect 2091 2654 2106 2670
rect 2172 2664 2191 2667
rect 1813 2642 1911 2644
rect 1938 2642 2106 2654
rect 2121 2644 2137 2658
rect 2172 2645 2194 2664
rect 2204 2658 2220 2659
rect 2203 2656 2220 2658
rect 2204 2651 2220 2656
rect 2194 2644 2200 2645
rect 2203 2644 2232 2651
rect 2121 2643 2232 2644
rect 2121 2642 2238 2643
rect 1797 2634 1848 2642
rect 1895 2634 1929 2642
rect 1797 2622 1822 2634
rect 1829 2622 1848 2634
rect 1902 2632 1929 2634
rect 1938 2632 2159 2642
rect 2194 2639 2200 2642
rect 1902 2628 2159 2632
rect 1797 2614 1848 2622
rect 1895 2614 2159 2628
rect 2203 2634 2238 2642
rect 1749 2566 1768 2600
rect 1813 2606 1842 2614
rect 1813 2600 1830 2606
rect 1813 2598 1847 2600
rect 1895 2598 1911 2614
rect 1912 2604 2120 2614
rect 2121 2604 2137 2614
rect 2185 2610 2200 2625
rect 2203 2622 2204 2634
rect 2211 2622 2238 2634
rect 2203 2614 2238 2622
rect 2203 2613 2232 2614
rect 1923 2600 2137 2604
rect 1938 2598 2137 2600
rect 2172 2600 2185 2610
rect 2203 2600 2220 2613
rect 2172 2598 2220 2600
rect 1814 2594 1847 2598
rect 1810 2592 1847 2594
rect 1810 2591 1877 2592
rect 1810 2586 1841 2591
rect 1847 2586 1877 2591
rect 1810 2582 1877 2586
rect 1783 2579 1877 2582
rect 1783 2572 1832 2579
rect 1783 2566 1813 2572
rect 1832 2567 1837 2572
rect 1749 2550 1829 2566
rect 1841 2558 1877 2579
rect 1938 2574 2127 2598
rect 2172 2597 2219 2598
rect 2185 2592 2219 2597
rect 1953 2571 2127 2574
rect 1946 2568 2127 2571
rect 2155 2591 2219 2592
rect 1749 2548 1768 2550
rect 1783 2548 1817 2550
rect 1749 2532 1829 2548
rect 1749 2526 1768 2532
rect 1465 2500 1568 2510
rect 1419 2498 1568 2500
rect 1589 2498 1624 2510
rect 1258 2496 1420 2498
rect 1270 2476 1289 2496
rect 1304 2494 1334 2496
rect 1153 2468 1194 2476
rect 1276 2472 1289 2476
rect 1341 2480 1420 2496
rect 1452 2496 1624 2498
rect 1452 2480 1531 2496
rect 1538 2494 1568 2496
rect 1116 2458 1145 2468
rect 1159 2458 1188 2468
rect 1203 2458 1233 2472
rect 1276 2458 1319 2472
rect 1341 2468 1531 2480
rect 1596 2476 1602 2496
rect 1326 2458 1356 2468
rect 1357 2458 1515 2468
rect 1519 2458 1549 2468
rect 1553 2458 1583 2472
rect 1611 2458 1624 2496
rect 1696 2510 1725 2526
rect 1739 2510 1768 2526
rect 1783 2516 1813 2532
rect 1841 2510 1847 2558
rect 1850 2552 1869 2558
rect 1884 2552 1914 2560
rect 1850 2544 1914 2552
rect 1850 2528 1930 2544
rect 1946 2537 2008 2568
rect 2024 2537 2086 2568
rect 2155 2566 2204 2591
rect 2219 2566 2249 2582
rect 2118 2552 2148 2560
rect 2155 2558 2265 2566
rect 2118 2544 2163 2552
rect 1850 2526 1869 2528
rect 1884 2526 1930 2528
rect 1850 2510 1930 2526
rect 1957 2524 1992 2537
rect 2033 2534 2070 2537
rect 2033 2532 2075 2534
rect 1962 2521 1992 2524
rect 1971 2517 1978 2521
rect 1978 2516 1979 2517
rect 1937 2510 1947 2516
rect 1696 2502 1731 2510
rect 1696 2476 1697 2502
rect 1704 2476 1731 2502
rect 1639 2458 1669 2472
rect 1696 2468 1731 2476
rect 1733 2502 1774 2510
rect 1733 2476 1748 2502
rect 1755 2476 1774 2502
rect 1838 2498 1869 2510
rect 1884 2498 1987 2510
rect 1999 2500 2025 2526
rect 2040 2521 2070 2532
rect 2102 2528 2164 2544
rect 2102 2526 2148 2528
rect 2102 2510 2164 2526
rect 2176 2510 2182 2558
rect 2185 2550 2265 2558
rect 2185 2548 2204 2550
rect 2219 2548 2253 2550
rect 2185 2532 2265 2548
rect 2185 2510 2204 2532
rect 2219 2516 2249 2532
rect 2277 2526 2283 2600
rect 2286 2526 2305 2670
rect 2320 2526 2326 2670
rect 2335 2600 2348 2670
rect 2400 2666 2422 2670
rect 2393 2644 2422 2658
rect 2475 2644 2491 2658
rect 2529 2654 2535 2656
rect 2542 2654 2650 2670
rect 2657 2654 2663 2656
rect 2671 2654 2686 2670
rect 2752 2664 2771 2667
rect 2393 2642 2491 2644
rect 2518 2642 2686 2654
rect 2701 2644 2717 2658
rect 2752 2645 2774 2664
rect 2784 2658 2800 2659
rect 2783 2656 2800 2658
rect 2784 2651 2800 2656
rect 2774 2644 2780 2645
rect 2783 2644 2812 2651
rect 2701 2643 2812 2644
rect 2701 2642 2818 2643
rect 2377 2634 2428 2642
rect 2475 2634 2509 2642
rect 2377 2622 2402 2634
rect 2409 2622 2428 2634
rect 2482 2632 2509 2634
rect 2518 2632 2739 2642
rect 2774 2639 2780 2642
rect 2482 2628 2739 2632
rect 2377 2614 2428 2622
rect 2475 2614 2739 2628
rect 2783 2634 2818 2642
rect 2329 2566 2348 2600
rect 2393 2606 2422 2614
rect 2393 2600 2410 2606
rect 2393 2598 2427 2600
rect 2475 2598 2491 2614
rect 2492 2604 2700 2614
rect 2701 2604 2717 2614
rect 2765 2610 2780 2625
rect 2783 2622 2784 2634
rect 2791 2622 2818 2634
rect 2783 2614 2818 2622
rect 2783 2613 2812 2614
rect 2503 2600 2717 2604
rect 2518 2598 2717 2600
rect 2752 2600 2765 2610
rect 2783 2600 2800 2613
rect 2752 2598 2800 2600
rect 2394 2594 2427 2598
rect 2390 2592 2427 2594
rect 2390 2591 2457 2592
rect 2390 2586 2421 2591
rect 2427 2586 2457 2591
rect 2390 2582 2457 2586
rect 2363 2579 2457 2582
rect 2363 2572 2412 2579
rect 2363 2566 2393 2572
rect 2412 2567 2417 2572
rect 2329 2550 2409 2566
rect 2421 2558 2457 2579
rect 2518 2574 2707 2598
rect 2752 2597 2799 2598
rect 2765 2592 2799 2597
rect 2533 2571 2707 2574
rect 2526 2568 2707 2571
rect 2735 2591 2799 2592
rect 2329 2548 2348 2550
rect 2363 2548 2397 2550
rect 2329 2532 2409 2548
rect 2329 2526 2348 2532
rect 2045 2500 2148 2510
rect 1999 2498 2148 2500
rect 2169 2498 2204 2510
rect 1838 2496 2000 2498
rect 1850 2476 1869 2496
rect 1884 2494 1914 2496
rect 1733 2468 1774 2476
rect 1856 2472 1869 2476
rect 1921 2480 2000 2496
rect 2032 2496 2204 2498
rect 2032 2480 2111 2496
rect 2118 2494 2148 2496
rect 1696 2458 1725 2468
rect 1739 2458 1768 2468
rect 1783 2458 1813 2472
rect 1856 2458 1899 2472
rect 1921 2468 2111 2480
rect 2176 2476 2182 2496
rect 1906 2458 1936 2468
rect 1937 2458 2095 2468
rect 2099 2458 2129 2468
rect 2133 2458 2163 2472
rect 2191 2458 2204 2496
rect 2276 2510 2305 2526
rect 2319 2510 2348 2526
rect 2363 2516 2393 2532
rect 2421 2510 2427 2558
rect 2430 2552 2449 2558
rect 2464 2552 2494 2560
rect 2430 2544 2494 2552
rect 2430 2528 2510 2544
rect 2526 2537 2588 2568
rect 2604 2537 2666 2568
rect 2735 2566 2784 2591
rect 2799 2566 2829 2582
rect 2698 2552 2728 2560
rect 2735 2558 2845 2566
rect 2698 2544 2743 2552
rect 2430 2526 2449 2528
rect 2464 2526 2510 2528
rect 2430 2510 2510 2526
rect 2537 2524 2572 2537
rect 2613 2534 2650 2537
rect 2613 2532 2655 2534
rect 2542 2521 2572 2524
rect 2551 2517 2558 2521
rect 2558 2516 2559 2517
rect 2517 2510 2527 2516
rect 2276 2502 2311 2510
rect 2276 2476 2277 2502
rect 2284 2476 2311 2502
rect 2219 2458 2249 2472
rect 2276 2468 2311 2476
rect 2313 2502 2354 2510
rect 2313 2476 2328 2502
rect 2335 2476 2354 2502
rect 2418 2498 2449 2510
rect 2464 2498 2567 2510
rect 2579 2500 2605 2526
rect 2620 2521 2650 2532
rect 2682 2528 2744 2544
rect 2682 2526 2728 2528
rect 2682 2510 2744 2526
rect 2756 2510 2762 2558
rect 2765 2550 2845 2558
rect 2765 2548 2784 2550
rect 2799 2548 2833 2550
rect 2765 2532 2845 2548
rect 2765 2510 2784 2532
rect 2799 2516 2829 2532
rect 2857 2526 2863 2600
rect 2866 2526 2885 2670
rect 2900 2526 2906 2670
rect 2915 2600 2928 2670
rect 2980 2666 3002 2670
rect 2973 2644 3002 2658
rect 3055 2644 3071 2658
rect 3109 2654 3115 2656
rect 3122 2654 3230 2670
rect 3237 2654 3243 2656
rect 3251 2654 3266 2670
rect 3332 2664 3351 2667
rect 2973 2642 3071 2644
rect 3098 2642 3266 2654
rect 3281 2644 3297 2658
rect 3332 2645 3354 2664
rect 3364 2658 3380 2659
rect 3363 2656 3380 2658
rect 3364 2651 3380 2656
rect 3354 2644 3360 2645
rect 3363 2644 3392 2651
rect 3281 2643 3392 2644
rect 3281 2642 3398 2643
rect 2957 2634 3008 2642
rect 3055 2634 3089 2642
rect 2957 2622 2982 2634
rect 2989 2622 3008 2634
rect 3062 2632 3089 2634
rect 3098 2632 3319 2642
rect 3354 2639 3360 2642
rect 3062 2628 3319 2632
rect 2957 2614 3008 2622
rect 3055 2614 3319 2628
rect 3363 2634 3398 2642
rect 2909 2566 2928 2600
rect 2973 2606 3002 2614
rect 2973 2600 2990 2606
rect 2973 2598 3007 2600
rect 3055 2598 3071 2614
rect 3072 2604 3280 2614
rect 3281 2604 3297 2614
rect 3345 2610 3360 2625
rect 3363 2622 3364 2634
rect 3371 2622 3398 2634
rect 3363 2614 3398 2622
rect 3363 2613 3392 2614
rect 3083 2600 3297 2604
rect 3098 2598 3297 2600
rect 3332 2600 3345 2610
rect 3363 2600 3380 2613
rect 3332 2598 3380 2600
rect 2974 2594 3007 2598
rect 2970 2592 3007 2594
rect 2970 2591 3037 2592
rect 2970 2586 3001 2591
rect 3007 2586 3037 2591
rect 2970 2582 3037 2586
rect 2943 2579 3037 2582
rect 2943 2572 2992 2579
rect 2943 2566 2973 2572
rect 2992 2567 2997 2572
rect 2909 2550 2989 2566
rect 3001 2558 3037 2579
rect 3098 2574 3287 2598
rect 3332 2597 3379 2598
rect 3345 2592 3379 2597
rect 3113 2571 3287 2574
rect 3106 2568 3287 2571
rect 3315 2591 3379 2592
rect 2909 2548 2928 2550
rect 2943 2548 2977 2550
rect 2909 2532 2989 2548
rect 2909 2526 2928 2532
rect 2625 2500 2728 2510
rect 2579 2498 2728 2500
rect 2749 2498 2784 2510
rect 2418 2496 2580 2498
rect 2430 2476 2449 2496
rect 2464 2494 2494 2496
rect 2313 2468 2354 2476
rect 2436 2472 2449 2476
rect 2501 2480 2580 2496
rect 2612 2496 2784 2498
rect 2612 2480 2691 2496
rect 2698 2494 2728 2496
rect 2276 2458 2305 2468
rect 2319 2458 2348 2468
rect 2363 2458 2393 2472
rect 2436 2458 2479 2472
rect 2501 2468 2691 2480
rect 2756 2476 2762 2496
rect 2486 2458 2516 2468
rect 2517 2458 2675 2468
rect 2679 2458 2709 2468
rect 2713 2458 2743 2472
rect 2771 2458 2784 2496
rect 2856 2510 2885 2526
rect 2899 2510 2928 2526
rect 2943 2516 2973 2532
rect 3001 2510 3007 2558
rect 3010 2552 3029 2558
rect 3044 2552 3074 2560
rect 3010 2544 3074 2552
rect 3010 2528 3090 2544
rect 3106 2537 3168 2568
rect 3184 2537 3246 2568
rect 3315 2566 3364 2591
rect 3379 2566 3409 2582
rect 3278 2552 3308 2560
rect 3315 2558 3425 2566
rect 3278 2544 3323 2552
rect 3010 2526 3029 2528
rect 3044 2526 3090 2528
rect 3010 2510 3090 2526
rect 3117 2524 3152 2537
rect 3193 2534 3230 2537
rect 3193 2532 3235 2534
rect 3122 2521 3152 2524
rect 3131 2517 3138 2521
rect 3138 2516 3139 2517
rect 3097 2510 3107 2516
rect 2856 2502 2891 2510
rect 2856 2476 2857 2502
rect 2864 2476 2891 2502
rect 2799 2458 2829 2472
rect 2856 2468 2891 2476
rect 2893 2502 2934 2510
rect 2893 2476 2908 2502
rect 2915 2476 2934 2502
rect 2998 2498 3029 2510
rect 3044 2498 3147 2510
rect 3159 2500 3185 2526
rect 3200 2521 3230 2532
rect 3262 2528 3324 2544
rect 3262 2526 3308 2528
rect 3262 2510 3324 2526
rect 3336 2510 3342 2558
rect 3345 2550 3425 2558
rect 3345 2548 3364 2550
rect 3379 2548 3413 2550
rect 3345 2532 3425 2548
rect 3345 2510 3364 2532
rect 3379 2516 3409 2532
rect 3437 2526 3443 2600
rect 3446 2526 3465 2670
rect 3480 2526 3486 2670
rect 3495 2600 3508 2670
rect 3560 2666 3582 2670
rect 3553 2644 3582 2658
rect 3635 2644 3651 2658
rect 3689 2654 3695 2656
rect 3702 2654 3810 2670
rect 3817 2654 3823 2656
rect 3831 2654 3846 2670
rect 3912 2664 3931 2667
rect 3553 2642 3651 2644
rect 3678 2642 3846 2654
rect 3861 2644 3877 2658
rect 3912 2645 3934 2664
rect 3944 2658 3960 2659
rect 3943 2656 3960 2658
rect 3944 2651 3960 2656
rect 3934 2644 3940 2645
rect 3943 2644 3972 2651
rect 3861 2643 3972 2644
rect 3861 2642 3978 2643
rect 3537 2634 3588 2642
rect 3635 2634 3669 2642
rect 3537 2622 3562 2634
rect 3569 2622 3588 2634
rect 3642 2632 3669 2634
rect 3678 2632 3899 2642
rect 3934 2639 3940 2642
rect 3642 2628 3899 2632
rect 3537 2614 3588 2622
rect 3635 2614 3899 2628
rect 3943 2634 3978 2642
rect 3489 2566 3508 2600
rect 3553 2606 3582 2614
rect 3553 2600 3570 2606
rect 3553 2598 3587 2600
rect 3635 2598 3651 2614
rect 3652 2604 3860 2614
rect 3861 2604 3877 2614
rect 3925 2610 3940 2625
rect 3943 2622 3944 2634
rect 3951 2622 3978 2634
rect 3943 2614 3978 2622
rect 3943 2613 3972 2614
rect 3663 2600 3877 2604
rect 3678 2598 3877 2600
rect 3912 2600 3925 2610
rect 3943 2600 3960 2613
rect 3912 2598 3960 2600
rect 3554 2594 3587 2598
rect 3550 2592 3587 2594
rect 3550 2591 3617 2592
rect 3550 2586 3581 2591
rect 3587 2586 3617 2591
rect 3550 2582 3617 2586
rect 3523 2579 3617 2582
rect 3523 2572 3572 2579
rect 3523 2566 3553 2572
rect 3572 2567 3577 2572
rect 3489 2550 3569 2566
rect 3581 2558 3617 2579
rect 3678 2574 3867 2598
rect 3912 2597 3959 2598
rect 3925 2592 3959 2597
rect 3693 2571 3867 2574
rect 3686 2568 3867 2571
rect 3895 2591 3959 2592
rect 3489 2548 3508 2550
rect 3523 2548 3557 2550
rect 3489 2532 3569 2548
rect 3489 2526 3508 2532
rect 3205 2500 3308 2510
rect 3159 2498 3308 2500
rect 3329 2498 3364 2510
rect 2998 2496 3160 2498
rect 3010 2476 3029 2496
rect 3044 2494 3074 2496
rect 2893 2468 2934 2476
rect 3016 2472 3029 2476
rect 3081 2480 3160 2496
rect 3192 2496 3364 2498
rect 3192 2480 3271 2496
rect 3278 2494 3308 2496
rect 2856 2458 2885 2468
rect 2899 2458 2928 2468
rect 2943 2458 2973 2472
rect 3016 2458 3059 2472
rect 3081 2468 3271 2480
rect 3336 2476 3342 2496
rect 3066 2458 3096 2468
rect 3097 2458 3255 2468
rect 3259 2458 3289 2468
rect 3293 2458 3323 2472
rect 3351 2458 3364 2496
rect 3436 2510 3465 2526
rect 3479 2510 3508 2526
rect 3523 2516 3553 2532
rect 3581 2510 3587 2558
rect 3590 2552 3609 2558
rect 3624 2552 3654 2560
rect 3590 2544 3654 2552
rect 3590 2528 3670 2544
rect 3686 2537 3748 2568
rect 3764 2537 3826 2568
rect 3895 2566 3944 2591
rect 3959 2566 3989 2582
rect 3858 2552 3888 2560
rect 3895 2558 4005 2566
rect 3858 2544 3903 2552
rect 3590 2526 3609 2528
rect 3624 2526 3670 2528
rect 3590 2510 3670 2526
rect 3697 2524 3732 2537
rect 3773 2534 3810 2537
rect 3773 2532 3815 2534
rect 3702 2521 3732 2524
rect 3711 2517 3718 2521
rect 3718 2516 3719 2517
rect 3677 2510 3687 2516
rect 3436 2502 3471 2510
rect 3436 2476 3437 2502
rect 3444 2476 3471 2502
rect 3379 2458 3409 2472
rect 3436 2468 3471 2476
rect 3473 2502 3514 2510
rect 3473 2476 3488 2502
rect 3495 2476 3514 2502
rect 3578 2498 3609 2510
rect 3624 2498 3727 2510
rect 3739 2500 3765 2526
rect 3780 2521 3810 2532
rect 3842 2528 3904 2544
rect 3842 2526 3888 2528
rect 3842 2510 3904 2526
rect 3916 2510 3922 2558
rect 3925 2550 4005 2558
rect 3925 2548 3944 2550
rect 3959 2548 3993 2550
rect 3925 2532 4005 2548
rect 3925 2510 3944 2532
rect 3959 2516 3989 2532
rect 4017 2526 4023 2600
rect 4026 2526 4045 2670
rect 4060 2526 4066 2670
rect 4075 2600 4088 2670
rect 4140 2666 4162 2670
rect 4133 2644 4162 2658
rect 4215 2644 4231 2658
rect 4269 2654 4275 2656
rect 4282 2654 4390 2670
rect 4397 2654 4403 2656
rect 4411 2654 4426 2670
rect 4492 2664 4511 2667
rect 4133 2642 4231 2644
rect 4258 2642 4426 2654
rect 4441 2644 4457 2658
rect 4492 2645 4514 2664
rect 4524 2658 4540 2659
rect 4523 2656 4540 2658
rect 4524 2651 4540 2656
rect 4514 2644 4520 2645
rect 4523 2644 4552 2651
rect 4441 2643 4552 2644
rect 4441 2642 4558 2643
rect 4117 2634 4168 2642
rect 4215 2634 4249 2642
rect 4117 2622 4142 2634
rect 4149 2622 4168 2634
rect 4222 2632 4249 2634
rect 4258 2632 4479 2642
rect 4514 2639 4520 2642
rect 4222 2628 4479 2632
rect 4117 2614 4168 2622
rect 4215 2614 4479 2628
rect 4523 2634 4558 2642
rect 4069 2566 4088 2600
rect 4133 2606 4162 2614
rect 4133 2600 4150 2606
rect 4133 2598 4167 2600
rect 4215 2598 4231 2614
rect 4232 2604 4440 2614
rect 4441 2604 4457 2614
rect 4505 2610 4520 2625
rect 4523 2622 4524 2634
rect 4531 2622 4558 2634
rect 4523 2614 4558 2622
rect 4523 2613 4552 2614
rect 4243 2600 4457 2604
rect 4258 2598 4457 2600
rect 4492 2600 4505 2610
rect 4523 2600 4540 2613
rect 4492 2598 4540 2600
rect 4134 2594 4167 2598
rect 4130 2592 4167 2594
rect 4130 2591 4197 2592
rect 4130 2586 4161 2591
rect 4167 2586 4197 2591
rect 4130 2582 4197 2586
rect 4103 2579 4197 2582
rect 4103 2572 4152 2579
rect 4103 2566 4133 2572
rect 4152 2567 4157 2572
rect 4069 2550 4149 2566
rect 4161 2558 4197 2579
rect 4258 2574 4447 2598
rect 4492 2597 4539 2598
rect 4505 2592 4539 2597
rect 4273 2571 4447 2574
rect 4266 2568 4447 2571
rect 4475 2591 4539 2592
rect 4069 2548 4088 2550
rect 4103 2548 4137 2550
rect 4069 2532 4149 2548
rect 4069 2526 4088 2532
rect 3785 2500 3888 2510
rect 3739 2498 3888 2500
rect 3909 2498 3944 2510
rect 3578 2496 3740 2498
rect 3590 2476 3609 2496
rect 3624 2494 3654 2496
rect 3473 2468 3514 2476
rect 3596 2472 3609 2476
rect 3661 2480 3740 2496
rect 3772 2496 3944 2498
rect 3772 2480 3851 2496
rect 3858 2494 3888 2496
rect 3436 2458 3465 2468
rect 3479 2458 3508 2468
rect 3523 2458 3553 2472
rect 3596 2458 3639 2472
rect 3661 2468 3851 2480
rect 3916 2476 3922 2496
rect 3646 2458 3676 2468
rect 3677 2458 3835 2468
rect 3839 2458 3869 2468
rect 3873 2458 3903 2472
rect 3931 2458 3944 2496
rect 4016 2510 4045 2526
rect 4059 2510 4088 2526
rect 4103 2516 4133 2532
rect 4161 2510 4167 2558
rect 4170 2552 4189 2558
rect 4204 2552 4234 2560
rect 4170 2544 4234 2552
rect 4170 2528 4250 2544
rect 4266 2537 4328 2568
rect 4344 2537 4406 2568
rect 4475 2566 4524 2591
rect 4539 2566 4569 2582
rect 4438 2552 4468 2560
rect 4475 2558 4585 2566
rect 4438 2544 4483 2552
rect 4170 2526 4189 2528
rect 4204 2526 4250 2528
rect 4170 2510 4250 2526
rect 4277 2524 4312 2537
rect 4353 2534 4390 2537
rect 4353 2532 4395 2534
rect 4282 2521 4312 2524
rect 4291 2517 4298 2521
rect 4298 2516 4299 2517
rect 4257 2510 4267 2516
rect 4016 2502 4051 2510
rect 4016 2476 4017 2502
rect 4024 2476 4051 2502
rect 3959 2458 3989 2472
rect 4016 2468 4051 2476
rect 4053 2502 4094 2510
rect 4053 2476 4068 2502
rect 4075 2476 4094 2502
rect 4158 2498 4189 2510
rect 4204 2498 4307 2510
rect 4319 2500 4345 2526
rect 4360 2521 4390 2532
rect 4422 2528 4484 2544
rect 4422 2526 4468 2528
rect 4422 2510 4484 2526
rect 4496 2510 4502 2558
rect 4505 2550 4585 2558
rect 4505 2548 4524 2550
rect 4539 2548 4573 2550
rect 4505 2532 4585 2548
rect 4505 2510 4524 2532
rect 4539 2516 4569 2532
rect 4597 2526 4603 2600
rect 4606 2526 4625 2670
rect 4640 2526 4646 2670
rect 4655 2600 4668 2670
rect 4720 2666 4742 2670
rect 4713 2644 4742 2658
rect 4795 2644 4811 2658
rect 4849 2654 4855 2656
rect 4862 2654 4970 2670
rect 4977 2654 4983 2656
rect 4991 2654 5006 2670
rect 5072 2664 5091 2667
rect 4713 2642 4811 2644
rect 4838 2642 5006 2654
rect 5021 2644 5037 2658
rect 5072 2645 5094 2664
rect 5104 2658 5120 2659
rect 5103 2656 5120 2658
rect 5104 2651 5120 2656
rect 5094 2644 5100 2645
rect 5103 2644 5132 2651
rect 5021 2643 5132 2644
rect 5021 2642 5138 2643
rect 4697 2634 4748 2642
rect 4795 2634 4829 2642
rect 4697 2622 4722 2634
rect 4729 2622 4748 2634
rect 4802 2632 4829 2634
rect 4838 2632 5059 2642
rect 5094 2639 5100 2642
rect 4802 2628 5059 2632
rect 4697 2614 4748 2622
rect 4795 2614 5059 2628
rect 5103 2634 5138 2642
rect 4649 2566 4668 2600
rect 4713 2606 4742 2614
rect 4713 2600 4730 2606
rect 4713 2598 4747 2600
rect 4795 2598 4811 2614
rect 4812 2604 5020 2614
rect 5021 2604 5037 2614
rect 5085 2610 5100 2625
rect 5103 2622 5104 2634
rect 5111 2622 5138 2634
rect 5103 2614 5138 2622
rect 5103 2613 5132 2614
rect 4823 2600 5037 2604
rect 4838 2598 5037 2600
rect 5072 2600 5085 2610
rect 5103 2600 5120 2613
rect 5072 2598 5120 2600
rect 4714 2594 4747 2598
rect 4710 2592 4747 2594
rect 4710 2591 4777 2592
rect 4710 2586 4741 2591
rect 4747 2586 4777 2591
rect 4710 2582 4777 2586
rect 4683 2579 4777 2582
rect 4683 2572 4732 2579
rect 4683 2566 4713 2572
rect 4732 2567 4737 2572
rect 4649 2550 4729 2566
rect 4741 2558 4777 2579
rect 4838 2574 5027 2598
rect 5072 2597 5119 2598
rect 5085 2592 5119 2597
rect 4853 2571 5027 2574
rect 4846 2568 5027 2571
rect 5055 2591 5119 2592
rect 4649 2548 4668 2550
rect 4683 2548 4717 2550
rect 4649 2532 4729 2548
rect 4649 2526 4668 2532
rect 4365 2500 4468 2510
rect 4319 2498 4468 2500
rect 4489 2498 4524 2510
rect 4158 2496 4320 2498
rect 4170 2476 4189 2496
rect 4204 2494 4234 2496
rect 4053 2468 4094 2476
rect 4176 2472 4189 2476
rect 4241 2480 4320 2496
rect 4352 2496 4524 2498
rect 4352 2480 4431 2496
rect 4438 2494 4468 2496
rect 4016 2458 4045 2468
rect 4059 2458 4088 2468
rect 4103 2458 4133 2472
rect 4176 2458 4219 2472
rect 4241 2468 4431 2480
rect 4496 2476 4502 2496
rect 4226 2458 4256 2468
rect 4257 2458 4415 2468
rect 4419 2458 4449 2468
rect 4453 2458 4483 2472
rect 4511 2458 4524 2496
rect 4596 2510 4625 2526
rect 4639 2510 4668 2526
rect 4683 2516 4713 2532
rect 4741 2510 4747 2558
rect 4750 2552 4769 2558
rect 4784 2552 4814 2560
rect 4750 2544 4814 2552
rect 4750 2528 4830 2544
rect 4846 2537 4908 2568
rect 4924 2537 4986 2568
rect 5055 2566 5104 2591
rect 5119 2566 5149 2582
rect 5018 2552 5048 2560
rect 5055 2558 5165 2566
rect 5018 2544 5063 2552
rect 4750 2526 4769 2528
rect 4784 2526 4830 2528
rect 4750 2510 4830 2526
rect 4857 2524 4892 2537
rect 4933 2534 4970 2537
rect 4933 2532 4975 2534
rect 4862 2521 4892 2524
rect 4871 2517 4878 2521
rect 4878 2516 4879 2517
rect 4837 2510 4847 2516
rect 4596 2502 4631 2510
rect 4596 2476 4597 2502
rect 4604 2476 4631 2502
rect 4539 2458 4569 2472
rect 4596 2468 4631 2476
rect 4633 2502 4674 2510
rect 4633 2476 4648 2502
rect 4655 2476 4674 2502
rect 4738 2498 4769 2510
rect 4784 2498 4887 2510
rect 4899 2500 4925 2526
rect 4940 2521 4970 2532
rect 5002 2528 5064 2544
rect 5002 2526 5048 2528
rect 5002 2510 5064 2526
rect 5076 2510 5082 2558
rect 5085 2550 5165 2558
rect 5085 2548 5104 2550
rect 5119 2548 5153 2550
rect 5085 2532 5165 2548
rect 5085 2510 5104 2532
rect 5119 2516 5149 2532
rect 5177 2526 5183 2600
rect 5186 2526 5205 2670
rect 5220 2526 5226 2670
rect 5235 2600 5248 2670
rect 5300 2666 5322 2670
rect 5293 2644 5322 2658
rect 5375 2644 5391 2658
rect 5429 2654 5435 2656
rect 5442 2654 5550 2670
rect 5557 2654 5563 2656
rect 5571 2654 5586 2670
rect 5652 2664 5671 2667
rect 5293 2642 5391 2644
rect 5418 2642 5586 2654
rect 5601 2644 5617 2658
rect 5652 2645 5674 2664
rect 5684 2658 5700 2659
rect 5683 2656 5700 2658
rect 5684 2651 5700 2656
rect 5674 2644 5680 2645
rect 5683 2644 5712 2651
rect 5601 2643 5712 2644
rect 5601 2642 5718 2643
rect 5277 2634 5328 2642
rect 5375 2634 5409 2642
rect 5277 2622 5302 2634
rect 5309 2622 5328 2634
rect 5382 2632 5409 2634
rect 5418 2632 5639 2642
rect 5674 2639 5680 2642
rect 5382 2628 5639 2632
rect 5277 2614 5328 2622
rect 5375 2614 5639 2628
rect 5683 2634 5718 2642
rect 5229 2566 5248 2600
rect 5293 2606 5322 2614
rect 5293 2600 5310 2606
rect 5293 2598 5327 2600
rect 5375 2598 5391 2614
rect 5392 2604 5600 2614
rect 5601 2604 5617 2614
rect 5665 2610 5680 2625
rect 5683 2622 5684 2634
rect 5691 2622 5718 2634
rect 5683 2614 5718 2622
rect 5683 2613 5712 2614
rect 5403 2600 5617 2604
rect 5418 2598 5617 2600
rect 5652 2600 5665 2610
rect 5683 2600 5700 2613
rect 5652 2598 5700 2600
rect 5294 2594 5327 2598
rect 5290 2592 5327 2594
rect 5290 2591 5357 2592
rect 5290 2586 5321 2591
rect 5327 2586 5357 2591
rect 5290 2582 5357 2586
rect 5263 2579 5357 2582
rect 5263 2572 5312 2579
rect 5263 2566 5293 2572
rect 5312 2567 5317 2572
rect 5229 2550 5309 2566
rect 5321 2558 5357 2579
rect 5418 2574 5607 2598
rect 5652 2597 5699 2598
rect 5665 2592 5699 2597
rect 5433 2571 5607 2574
rect 5426 2568 5607 2571
rect 5635 2591 5699 2592
rect 5229 2548 5248 2550
rect 5263 2548 5297 2550
rect 5229 2532 5309 2548
rect 5229 2526 5248 2532
rect 4945 2500 5048 2510
rect 4899 2498 5048 2500
rect 5069 2498 5104 2510
rect 4738 2496 4900 2498
rect 4750 2476 4769 2496
rect 4784 2494 4814 2496
rect 4633 2468 4674 2476
rect 4756 2472 4769 2476
rect 4821 2480 4900 2496
rect 4932 2496 5104 2498
rect 4932 2480 5011 2496
rect 5018 2494 5048 2496
rect 4596 2458 4625 2468
rect 4639 2458 4668 2468
rect 4683 2458 4713 2472
rect 4756 2458 4799 2472
rect 4821 2468 5011 2480
rect 5076 2476 5082 2496
rect 4806 2458 4836 2468
rect 4837 2458 4995 2468
rect 4999 2458 5029 2468
rect 5033 2458 5063 2472
rect 5091 2458 5104 2496
rect 5176 2510 5205 2526
rect 5219 2510 5248 2526
rect 5263 2516 5293 2532
rect 5321 2510 5327 2558
rect 5330 2552 5349 2558
rect 5364 2552 5394 2560
rect 5330 2544 5394 2552
rect 5330 2528 5410 2544
rect 5426 2537 5488 2568
rect 5504 2537 5566 2568
rect 5635 2566 5684 2591
rect 5699 2566 5729 2582
rect 5598 2552 5628 2560
rect 5635 2558 5745 2566
rect 5598 2544 5643 2552
rect 5330 2526 5349 2528
rect 5364 2526 5410 2528
rect 5330 2510 5410 2526
rect 5437 2524 5472 2537
rect 5513 2534 5550 2537
rect 5513 2532 5555 2534
rect 5442 2521 5472 2524
rect 5451 2517 5458 2521
rect 5458 2516 5459 2517
rect 5417 2510 5427 2516
rect 5176 2502 5211 2510
rect 5176 2476 5177 2502
rect 5184 2476 5211 2502
rect 5119 2458 5149 2472
rect 5176 2468 5211 2476
rect 5213 2502 5254 2510
rect 5213 2476 5228 2502
rect 5235 2476 5254 2502
rect 5318 2498 5349 2510
rect 5364 2498 5467 2510
rect 5479 2500 5505 2526
rect 5520 2521 5550 2532
rect 5582 2528 5644 2544
rect 5582 2526 5628 2528
rect 5582 2510 5644 2526
rect 5656 2510 5662 2558
rect 5665 2550 5745 2558
rect 5665 2548 5684 2550
rect 5699 2548 5733 2550
rect 5665 2532 5745 2548
rect 5665 2510 5684 2532
rect 5699 2516 5729 2532
rect 5757 2526 5763 2600
rect 5766 2526 5785 2670
rect 5800 2526 5806 2670
rect 5815 2600 5828 2670
rect 5880 2666 5902 2670
rect 5873 2644 5902 2658
rect 5955 2644 5971 2658
rect 6009 2654 6015 2656
rect 6022 2654 6130 2670
rect 6137 2654 6143 2656
rect 6151 2654 6166 2670
rect 6232 2664 6251 2667
rect 5873 2642 5971 2644
rect 5998 2642 6166 2654
rect 6181 2644 6197 2658
rect 6232 2645 6254 2664
rect 6264 2658 6280 2659
rect 6263 2656 6280 2658
rect 6264 2651 6280 2656
rect 6254 2644 6260 2645
rect 6263 2644 6292 2651
rect 6181 2643 6292 2644
rect 6181 2642 6298 2643
rect 5857 2634 5908 2642
rect 5955 2634 5989 2642
rect 5857 2622 5882 2634
rect 5889 2622 5908 2634
rect 5962 2632 5989 2634
rect 5998 2632 6219 2642
rect 6254 2639 6260 2642
rect 5962 2628 6219 2632
rect 5857 2614 5908 2622
rect 5955 2614 6219 2628
rect 6263 2634 6298 2642
rect 5809 2566 5828 2600
rect 5873 2606 5902 2614
rect 5873 2600 5890 2606
rect 5873 2598 5907 2600
rect 5955 2598 5971 2614
rect 5972 2604 6180 2614
rect 6181 2604 6197 2614
rect 6245 2610 6260 2625
rect 6263 2622 6264 2634
rect 6271 2622 6298 2634
rect 6263 2614 6298 2622
rect 6263 2613 6292 2614
rect 5983 2600 6197 2604
rect 5998 2598 6197 2600
rect 6232 2600 6245 2610
rect 6263 2600 6280 2613
rect 6232 2598 6280 2600
rect 5874 2594 5907 2598
rect 5870 2592 5907 2594
rect 5870 2591 5937 2592
rect 5870 2586 5901 2591
rect 5907 2586 5937 2591
rect 5870 2582 5937 2586
rect 5843 2579 5937 2582
rect 5843 2572 5892 2579
rect 5843 2566 5873 2572
rect 5892 2567 5897 2572
rect 5809 2550 5889 2566
rect 5901 2558 5937 2579
rect 5998 2574 6187 2598
rect 6232 2597 6279 2598
rect 6245 2592 6279 2597
rect 6013 2571 6187 2574
rect 6006 2568 6187 2571
rect 6215 2591 6279 2592
rect 5809 2548 5828 2550
rect 5843 2548 5877 2550
rect 5809 2532 5889 2548
rect 5809 2526 5828 2532
rect 5525 2500 5628 2510
rect 5479 2498 5628 2500
rect 5649 2498 5684 2510
rect 5318 2496 5480 2498
rect 5330 2476 5349 2496
rect 5364 2494 5394 2496
rect 5213 2468 5254 2476
rect 5336 2472 5349 2476
rect 5401 2480 5480 2496
rect 5512 2496 5684 2498
rect 5512 2480 5591 2496
rect 5598 2494 5628 2496
rect 5176 2458 5205 2468
rect 5219 2458 5248 2468
rect 5263 2458 5293 2472
rect 5336 2458 5379 2472
rect 5401 2468 5591 2480
rect 5656 2476 5662 2496
rect 5386 2458 5416 2468
rect 5417 2458 5575 2468
rect 5579 2458 5609 2468
rect 5613 2458 5643 2472
rect 5671 2458 5684 2496
rect 5756 2510 5785 2526
rect 5799 2510 5828 2526
rect 5843 2516 5873 2532
rect 5901 2510 5907 2558
rect 5910 2552 5929 2558
rect 5944 2552 5974 2560
rect 5910 2544 5974 2552
rect 5910 2528 5990 2544
rect 6006 2537 6068 2568
rect 6084 2537 6146 2568
rect 6215 2566 6264 2591
rect 6279 2566 6309 2582
rect 6178 2552 6208 2560
rect 6215 2558 6325 2566
rect 6178 2544 6223 2552
rect 5910 2526 5929 2528
rect 5944 2526 5990 2528
rect 5910 2510 5990 2526
rect 6017 2524 6052 2537
rect 6093 2534 6130 2537
rect 6093 2532 6135 2534
rect 6022 2521 6052 2524
rect 6031 2517 6038 2521
rect 6038 2516 6039 2517
rect 5997 2510 6007 2516
rect 5756 2502 5791 2510
rect 5756 2476 5757 2502
rect 5764 2476 5791 2502
rect 5699 2458 5729 2472
rect 5756 2468 5791 2476
rect 5793 2502 5834 2510
rect 5793 2476 5808 2502
rect 5815 2476 5834 2502
rect 5898 2498 5929 2510
rect 5944 2498 6047 2510
rect 6059 2500 6085 2526
rect 6100 2521 6130 2532
rect 6162 2528 6224 2544
rect 6162 2526 6208 2528
rect 6162 2510 6224 2526
rect 6236 2510 6242 2558
rect 6245 2550 6325 2558
rect 6245 2548 6264 2550
rect 6279 2548 6313 2550
rect 6245 2532 6325 2548
rect 6245 2510 6264 2532
rect 6279 2516 6309 2532
rect 6337 2526 6343 2600
rect 6346 2526 6365 2670
rect 6380 2526 6386 2670
rect 6395 2600 6408 2670
rect 6460 2666 6482 2670
rect 6453 2644 6482 2658
rect 6535 2644 6551 2658
rect 6589 2654 6595 2656
rect 6602 2654 6710 2670
rect 6717 2654 6723 2656
rect 6731 2654 6746 2670
rect 6812 2664 6831 2667
rect 6453 2642 6551 2644
rect 6578 2642 6746 2654
rect 6761 2644 6777 2658
rect 6812 2645 6834 2664
rect 6844 2658 6860 2659
rect 6843 2656 6860 2658
rect 6844 2651 6860 2656
rect 6834 2644 6840 2645
rect 6843 2644 6872 2651
rect 6761 2643 6872 2644
rect 6761 2642 6878 2643
rect 6437 2634 6488 2642
rect 6535 2634 6569 2642
rect 6437 2622 6462 2634
rect 6469 2622 6488 2634
rect 6542 2632 6569 2634
rect 6578 2632 6799 2642
rect 6834 2639 6840 2642
rect 6542 2628 6799 2632
rect 6437 2614 6488 2622
rect 6535 2614 6799 2628
rect 6843 2634 6878 2642
rect 6389 2566 6408 2600
rect 6453 2606 6482 2614
rect 6453 2600 6470 2606
rect 6453 2598 6487 2600
rect 6535 2598 6551 2614
rect 6552 2604 6760 2614
rect 6761 2604 6777 2614
rect 6825 2610 6840 2625
rect 6843 2622 6844 2634
rect 6851 2622 6878 2634
rect 6843 2614 6878 2622
rect 6843 2613 6872 2614
rect 6563 2600 6777 2604
rect 6578 2598 6777 2600
rect 6812 2600 6825 2610
rect 6843 2600 6860 2613
rect 6812 2598 6860 2600
rect 6454 2594 6487 2598
rect 6450 2592 6487 2594
rect 6450 2591 6517 2592
rect 6450 2586 6481 2591
rect 6487 2586 6517 2591
rect 6450 2582 6517 2586
rect 6423 2579 6517 2582
rect 6423 2572 6472 2579
rect 6423 2566 6453 2572
rect 6472 2567 6477 2572
rect 6389 2550 6469 2566
rect 6481 2558 6517 2579
rect 6578 2574 6767 2598
rect 6812 2597 6859 2598
rect 6825 2592 6859 2597
rect 6593 2571 6767 2574
rect 6586 2568 6767 2571
rect 6795 2591 6859 2592
rect 6389 2548 6408 2550
rect 6423 2548 6457 2550
rect 6389 2532 6469 2548
rect 6389 2526 6408 2532
rect 6105 2500 6208 2510
rect 6059 2498 6208 2500
rect 6229 2498 6264 2510
rect 5898 2496 6060 2498
rect 5910 2476 5929 2496
rect 5944 2494 5974 2496
rect 5793 2468 5834 2476
rect 5916 2472 5929 2476
rect 5981 2480 6060 2496
rect 6092 2496 6264 2498
rect 6092 2480 6171 2496
rect 6178 2494 6208 2496
rect 5756 2458 5785 2468
rect 5799 2458 5828 2468
rect 5843 2458 5873 2472
rect 5916 2458 5959 2472
rect 5981 2468 6171 2480
rect 6236 2476 6242 2496
rect 5966 2458 5996 2468
rect 5997 2458 6155 2468
rect 6159 2458 6189 2468
rect 6193 2458 6223 2472
rect 6251 2458 6264 2496
rect 6336 2510 6365 2526
rect 6379 2510 6408 2526
rect 6423 2516 6453 2532
rect 6481 2510 6487 2558
rect 6490 2552 6509 2558
rect 6524 2552 6554 2560
rect 6490 2544 6554 2552
rect 6490 2528 6570 2544
rect 6586 2537 6648 2568
rect 6664 2537 6726 2568
rect 6795 2566 6844 2591
rect 6859 2566 6889 2582
rect 6758 2552 6788 2560
rect 6795 2558 6905 2566
rect 6758 2544 6803 2552
rect 6490 2526 6509 2528
rect 6524 2526 6570 2528
rect 6490 2510 6570 2526
rect 6597 2524 6632 2537
rect 6673 2534 6710 2537
rect 6673 2532 6715 2534
rect 6602 2521 6632 2524
rect 6611 2517 6618 2521
rect 6618 2516 6619 2517
rect 6577 2510 6587 2516
rect 6336 2502 6371 2510
rect 6336 2476 6337 2502
rect 6344 2476 6371 2502
rect 6279 2458 6309 2472
rect 6336 2468 6371 2476
rect 6373 2502 6414 2510
rect 6373 2476 6388 2502
rect 6395 2476 6414 2502
rect 6478 2498 6509 2510
rect 6524 2498 6627 2510
rect 6639 2500 6665 2526
rect 6680 2521 6710 2532
rect 6742 2528 6804 2544
rect 6742 2526 6788 2528
rect 6742 2510 6804 2526
rect 6816 2510 6822 2558
rect 6825 2550 6905 2558
rect 6825 2548 6844 2550
rect 6859 2548 6893 2550
rect 6825 2532 6905 2548
rect 6825 2510 6844 2532
rect 6859 2516 6889 2532
rect 6917 2526 6923 2600
rect 6926 2526 6945 2670
rect 6960 2526 6966 2670
rect 6975 2600 6988 2670
rect 7040 2666 7062 2670
rect 7033 2644 7062 2658
rect 7115 2644 7131 2658
rect 7169 2654 7175 2656
rect 7182 2654 7290 2670
rect 7297 2654 7303 2656
rect 7311 2654 7326 2670
rect 7392 2664 7411 2667
rect 7033 2642 7131 2644
rect 7158 2642 7326 2654
rect 7341 2644 7357 2658
rect 7392 2645 7414 2664
rect 7424 2658 7440 2659
rect 7423 2656 7440 2658
rect 7424 2651 7440 2656
rect 7414 2644 7420 2645
rect 7423 2644 7452 2651
rect 7341 2643 7452 2644
rect 7341 2642 7458 2643
rect 7017 2634 7068 2642
rect 7115 2634 7149 2642
rect 7017 2622 7042 2634
rect 7049 2622 7068 2634
rect 7122 2632 7149 2634
rect 7158 2632 7379 2642
rect 7414 2639 7420 2642
rect 7122 2628 7379 2632
rect 7017 2614 7068 2622
rect 7115 2614 7379 2628
rect 7423 2634 7458 2642
rect 6969 2566 6988 2600
rect 7033 2606 7062 2614
rect 7033 2600 7050 2606
rect 7033 2598 7067 2600
rect 7115 2598 7131 2614
rect 7132 2604 7340 2614
rect 7341 2604 7357 2614
rect 7405 2610 7420 2625
rect 7423 2622 7424 2634
rect 7431 2622 7458 2634
rect 7423 2614 7458 2622
rect 7423 2613 7452 2614
rect 7143 2600 7357 2604
rect 7158 2598 7357 2600
rect 7392 2600 7405 2610
rect 7423 2600 7440 2613
rect 7392 2598 7440 2600
rect 7034 2594 7067 2598
rect 7030 2592 7067 2594
rect 7030 2591 7097 2592
rect 7030 2586 7061 2591
rect 7067 2586 7097 2591
rect 7030 2582 7097 2586
rect 7003 2579 7097 2582
rect 7003 2572 7052 2579
rect 7003 2566 7033 2572
rect 7052 2567 7057 2572
rect 6969 2550 7049 2566
rect 7061 2558 7097 2579
rect 7158 2574 7347 2598
rect 7392 2597 7439 2598
rect 7405 2592 7439 2597
rect 7173 2571 7347 2574
rect 7166 2568 7347 2571
rect 7375 2591 7439 2592
rect 6969 2548 6988 2550
rect 7003 2548 7037 2550
rect 6969 2532 7049 2548
rect 6969 2526 6988 2532
rect 6685 2500 6788 2510
rect 6639 2498 6788 2500
rect 6809 2498 6844 2510
rect 6478 2496 6640 2498
rect 6490 2476 6509 2496
rect 6524 2494 6554 2496
rect 6373 2468 6414 2476
rect 6496 2472 6509 2476
rect 6561 2480 6640 2496
rect 6672 2496 6844 2498
rect 6672 2480 6751 2496
rect 6758 2494 6788 2496
rect 6336 2458 6365 2468
rect 6379 2458 6408 2468
rect 6423 2458 6453 2472
rect 6496 2458 6539 2472
rect 6561 2468 6751 2480
rect 6816 2476 6822 2496
rect 6546 2458 6576 2468
rect 6577 2458 6735 2468
rect 6739 2458 6769 2468
rect 6773 2458 6803 2472
rect 6831 2458 6844 2496
rect 6916 2510 6945 2526
rect 6959 2510 6988 2526
rect 7003 2516 7033 2532
rect 7061 2510 7067 2558
rect 7070 2552 7089 2558
rect 7104 2552 7134 2560
rect 7070 2544 7134 2552
rect 7070 2528 7150 2544
rect 7166 2537 7228 2568
rect 7244 2537 7306 2568
rect 7375 2566 7424 2591
rect 7439 2566 7469 2582
rect 7338 2552 7368 2560
rect 7375 2558 7485 2566
rect 7338 2544 7383 2552
rect 7070 2526 7089 2528
rect 7104 2526 7150 2528
rect 7070 2510 7150 2526
rect 7177 2524 7212 2537
rect 7253 2534 7290 2537
rect 7253 2532 7295 2534
rect 7182 2521 7212 2524
rect 7191 2517 7198 2521
rect 7198 2516 7199 2517
rect 7157 2510 7167 2516
rect 6916 2502 6951 2510
rect 6916 2476 6917 2502
rect 6924 2476 6951 2502
rect 6859 2458 6889 2472
rect 6916 2468 6951 2476
rect 6953 2502 6994 2510
rect 6953 2476 6968 2502
rect 6975 2476 6994 2502
rect 7058 2498 7089 2510
rect 7104 2498 7207 2510
rect 7219 2500 7245 2526
rect 7260 2521 7290 2532
rect 7322 2528 7384 2544
rect 7322 2526 7368 2528
rect 7322 2510 7384 2526
rect 7396 2510 7402 2558
rect 7405 2550 7485 2558
rect 7405 2548 7424 2550
rect 7439 2548 7473 2550
rect 7405 2532 7485 2548
rect 7405 2510 7424 2532
rect 7439 2516 7469 2532
rect 7497 2526 7503 2600
rect 7506 2526 7525 2670
rect 7540 2526 7546 2670
rect 7555 2600 7568 2670
rect 7620 2666 7642 2670
rect 7613 2644 7642 2658
rect 7695 2644 7711 2658
rect 7749 2654 7755 2656
rect 7762 2654 7870 2670
rect 7877 2654 7883 2656
rect 7891 2654 7906 2670
rect 7972 2664 7991 2667
rect 7613 2642 7711 2644
rect 7738 2642 7906 2654
rect 7921 2644 7937 2658
rect 7972 2645 7994 2664
rect 8004 2658 8020 2659
rect 8003 2656 8020 2658
rect 8004 2651 8020 2656
rect 7994 2644 8000 2645
rect 8003 2644 8032 2651
rect 7921 2643 8032 2644
rect 7921 2642 8038 2643
rect 7597 2634 7648 2642
rect 7695 2634 7729 2642
rect 7597 2622 7622 2634
rect 7629 2622 7648 2634
rect 7702 2632 7729 2634
rect 7738 2632 7959 2642
rect 7994 2639 8000 2642
rect 7702 2628 7959 2632
rect 7597 2614 7648 2622
rect 7695 2614 7959 2628
rect 8003 2634 8038 2642
rect 7549 2566 7568 2600
rect 7613 2606 7642 2614
rect 7613 2600 7630 2606
rect 7613 2598 7647 2600
rect 7695 2598 7711 2614
rect 7712 2604 7920 2614
rect 7921 2604 7937 2614
rect 7985 2610 8000 2625
rect 8003 2622 8004 2634
rect 8011 2622 8038 2634
rect 8003 2614 8038 2622
rect 8003 2613 8032 2614
rect 7723 2600 7937 2604
rect 7738 2598 7937 2600
rect 7972 2600 7985 2610
rect 8003 2600 8020 2613
rect 7972 2598 8020 2600
rect 7614 2594 7647 2598
rect 7610 2592 7647 2594
rect 7610 2591 7677 2592
rect 7610 2586 7641 2591
rect 7647 2586 7677 2591
rect 7610 2582 7677 2586
rect 7583 2579 7677 2582
rect 7583 2572 7632 2579
rect 7583 2566 7613 2572
rect 7632 2567 7637 2572
rect 7549 2550 7629 2566
rect 7641 2558 7677 2579
rect 7738 2574 7927 2598
rect 7972 2597 8019 2598
rect 7985 2592 8019 2597
rect 7753 2571 7927 2574
rect 7746 2568 7927 2571
rect 7955 2591 8019 2592
rect 7549 2548 7568 2550
rect 7583 2548 7617 2550
rect 7549 2532 7629 2548
rect 7549 2526 7568 2532
rect 7265 2500 7368 2510
rect 7219 2498 7368 2500
rect 7389 2498 7424 2510
rect 7058 2496 7220 2498
rect 7070 2476 7089 2496
rect 7104 2494 7134 2496
rect 6953 2468 6994 2476
rect 7076 2472 7089 2476
rect 7141 2480 7220 2496
rect 7252 2496 7424 2498
rect 7252 2480 7331 2496
rect 7338 2494 7368 2496
rect 6916 2458 6945 2468
rect 6959 2458 6988 2468
rect 7003 2458 7033 2472
rect 7076 2458 7119 2472
rect 7141 2468 7331 2480
rect 7396 2476 7402 2496
rect 7126 2458 7156 2468
rect 7157 2458 7315 2468
rect 7319 2458 7349 2468
rect 7353 2458 7383 2472
rect 7411 2458 7424 2496
rect 7496 2510 7525 2526
rect 7539 2510 7568 2526
rect 7583 2516 7613 2532
rect 7641 2510 7647 2558
rect 7650 2552 7669 2558
rect 7684 2552 7714 2560
rect 7650 2544 7714 2552
rect 7650 2528 7730 2544
rect 7746 2537 7808 2568
rect 7824 2537 7886 2568
rect 7955 2566 8004 2591
rect 8019 2566 8049 2582
rect 7918 2552 7948 2560
rect 7955 2558 8065 2566
rect 7918 2544 7963 2552
rect 7650 2526 7669 2528
rect 7684 2526 7730 2528
rect 7650 2510 7730 2526
rect 7757 2524 7792 2537
rect 7833 2534 7870 2537
rect 7833 2532 7875 2534
rect 7762 2521 7792 2524
rect 7771 2517 7778 2521
rect 7778 2516 7779 2517
rect 7737 2510 7747 2516
rect 7496 2502 7531 2510
rect 7496 2476 7497 2502
rect 7504 2476 7531 2502
rect 7439 2458 7469 2472
rect 7496 2468 7531 2476
rect 7533 2502 7574 2510
rect 7533 2476 7548 2502
rect 7555 2476 7574 2502
rect 7638 2498 7669 2510
rect 7684 2498 7787 2510
rect 7799 2500 7825 2526
rect 7840 2521 7870 2532
rect 7902 2528 7964 2544
rect 7902 2526 7948 2528
rect 7902 2510 7964 2526
rect 7976 2510 7982 2558
rect 7985 2550 8065 2558
rect 7985 2548 8004 2550
rect 8019 2548 8053 2550
rect 7985 2532 8065 2548
rect 7985 2510 8004 2532
rect 8019 2516 8049 2532
rect 8077 2526 8083 2600
rect 8086 2526 8105 2670
rect 8120 2526 8126 2670
rect 8135 2600 8148 2670
rect 8200 2666 8222 2670
rect 8193 2644 8222 2658
rect 8275 2644 8291 2658
rect 8329 2654 8335 2656
rect 8342 2654 8450 2670
rect 8457 2654 8463 2656
rect 8471 2654 8486 2670
rect 8552 2664 8571 2667
rect 8193 2642 8291 2644
rect 8318 2642 8486 2654
rect 8501 2644 8517 2658
rect 8552 2645 8574 2664
rect 8584 2658 8600 2659
rect 8583 2656 8600 2658
rect 8584 2651 8600 2656
rect 8574 2644 8580 2645
rect 8583 2644 8612 2651
rect 8501 2643 8612 2644
rect 8501 2642 8618 2643
rect 8177 2634 8228 2642
rect 8275 2634 8309 2642
rect 8177 2622 8202 2634
rect 8209 2622 8228 2634
rect 8282 2632 8309 2634
rect 8318 2632 8539 2642
rect 8574 2639 8580 2642
rect 8282 2628 8539 2632
rect 8177 2614 8228 2622
rect 8275 2614 8539 2628
rect 8583 2634 8618 2642
rect 8129 2566 8148 2600
rect 8193 2606 8222 2614
rect 8193 2600 8210 2606
rect 8193 2598 8227 2600
rect 8275 2598 8291 2614
rect 8292 2604 8500 2614
rect 8501 2604 8517 2614
rect 8565 2610 8580 2625
rect 8583 2622 8584 2634
rect 8591 2622 8618 2634
rect 8583 2614 8618 2622
rect 8583 2613 8612 2614
rect 8303 2600 8517 2604
rect 8318 2598 8517 2600
rect 8552 2600 8565 2610
rect 8583 2600 8600 2613
rect 8552 2598 8600 2600
rect 8194 2594 8227 2598
rect 8190 2592 8227 2594
rect 8190 2591 8257 2592
rect 8190 2586 8221 2591
rect 8227 2586 8257 2591
rect 8190 2582 8257 2586
rect 8163 2579 8257 2582
rect 8163 2572 8212 2579
rect 8163 2566 8193 2572
rect 8212 2567 8217 2572
rect 8129 2550 8209 2566
rect 8221 2558 8257 2579
rect 8318 2574 8507 2598
rect 8552 2597 8599 2598
rect 8565 2592 8599 2597
rect 8333 2571 8507 2574
rect 8326 2568 8507 2571
rect 8535 2591 8599 2592
rect 8129 2548 8148 2550
rect 8163 2548 8197 2550
rect 8129 2532 8209 2548
rect 8129 2526 8148 2532
rect 7845 2500 7948 2510
rect 7799 2498 7948 2500
rect 7969 2498 8004 2510
rect 7638 2496 7800 2498
rect 7650 2476 7669 2496
rect 7684 2494 7714 2496
rect 7533 2468 7574 2476
rect 7656 2472 7669 2476
rect 7721 2480 7800 2496
rect 7832 2496 8004 2498
rect 7832 2480 7911 2496
rect 7918 2494 7948 2496
rect 7496 2458 7525 2468
rect 7539 2458 7568 2468
rect 7583 2458 7613 2472
rect 7656 2458 7699 2472
rect 7721 2468 7911 2480
rect 7976 2476 7982 2496
rect 7706 2458 7736 2468
rect 7737 2458 7895 2468
rect 7899 2458 7929 2468
rect 7933 2458 7963 2472
rect 7991 2458 8004 2496
rect 8076 2510 8105 2526
rect 8119 2510 8148 2526
rect 8163 2516 8193 2532
rect 8221 2510 8227 2558
rect 8230 2552 8249 2558
rect 8264 2552 8294 2560
rect 8230 2544 8294 2552
rect 8230 2528 8310 2544
rect 8326 2537 8388 2568
rect 8404 2537 8466 2568
rect 8535 2566 8584 2591
rect 8599 2566 8629 2582
rect 8498 2552 8528 2560
rect 8535 2558 8645 2566
rect 8498 2544 8543 2552
rect 8230 2526 8249 2528
rect 8264 2526 8310 2528
rect 8230 2510 8310 2526
rect 8337 2524 8372 2537
rect 8413 2534 8450 2537
rect 8413 2532 8455 2534
rect 8342 2521 8372 2524
rect 8351 2517 8358 2521
rect 8358 2516 8359 2517
rect 8317 2510 8327 2516
rect 8076 2502 8111 2510
rect 8076 2476 8077 2502
rect 8084 2476 8111 2502
rect 8019 2458 8049 2472
rect 8076 2468 8111 2476
rect 8113 2502 8154 2510
rect 8113 2476 8128 2502
rect 8135 2476 8154 2502
rect 8218 2498 8249 2510
rect 8264 2498 8367 2510
rect 8379 2500 8405 2526
rect 8420 2521 8450 2532
rect 8482 2528 8544 2544
rect 8482 2526 8528 2528
rect 8482 2510 8544 2526
rect 8556 2510 8562 2558
rect 8565 2550 8645 2558
rect 8565 2548 8584 2550
rect 8599 2548 8633 2550
rect 8565 2532 8645 2548
rect 8565 2510 8584 2532
rect 8599 2516 8629 2532
rect 8657 2526 8663 2600
rect 8666 2526 8685 2670
rect 8700 2526 8706 2670
rect 8715 2600 8728 2670
rect 8780 2666 8802 2670
rect 8773 2644 8802 2658
rect 8855 2644 8871 2658
rect 8909 2654 8915 2656
rect 8922 2654 9030 2670
rect 9037 2654 9043 2656
rect 9051 2654 9066 2670
rect 9132 2664 9151 2667
rect 8773 2642 8871 2644
rect 8898 2642 9066 2654
rect 9081 2644 9097 2658
rect 9132 2645 9154 2664
rect 9164 2658 9180 2659
rect 9163 2656 9180 2658
rect 9164 2651 9180 2656
rect 9154 2644 9160 2645
rect 9163 2644 9192 2651
rect 9081 2643 9192 2644
rect 9081 2642 9198 2643
rect 8757 2634 8808 2642
rect 8855 2634 8889 2642
rect 8757 2622 8782 2634
rect 8789 2622 8808 2634
rect 8862 2632 8889 2634
rect 8898 2632 9119 2642
rect 9154 2639 9160 2642
rect 8862 2628 9119 2632
rect 8757 2614 8808 2622
rect 8855 2614 9119 2628
rect 9163 2634 9198 2642
rect 8709 2566 8728 2600
rect 8773 2606 8802 2614
rect 8773 2600 8790 2606
rect 8773 2598 8807 2600
rect 8855 2598 8871 2614
rect 8872 2604 9080 2614
rect 9081 2604 9097 2614
rect 9145 2610 9160 2625
rect 9163 2622 9164 2634
rect 9171 2622 9198 2634
rect 9163 2614 9198 2622
rect 9163 2613 9192 2614
rect 8883 2600 9097 2604
rect 8898 2598 9097 2600
rect 9132 2600 9145 2610
rect 9163 2600 9180 2613
rect 9132 2598 9180 2600
rect 8774 2594 8807 2598
rect 8770 2592 8807 2594
rect 8770 2591 8837 2592
rect 8770 2586 8801 2591
rect 8807 2586 8837 2591
rect 8770 2582 8837 2586
rect 8743 2579 8837 2582
rect 8743 2572 8792 2579
rect 8743 2566 8773 2572
rect 8792 2567 8797 2572
rect 8709 2550 8789 2566
rect 8801 2558 8837 2579
rect 8898 2574 9087 2598
rect 9132 2597 9179 2598
rect 9145 2592 9179 2597
rect 8913 2571 9087 2574
rect 8906 2568 9087 2571
rect 9115 2591 9179 2592
rect 8709 2548 8728 2550
rect 8743 2548 8777 2550
rect 8709 2532 8789 2548
rect 8709 2526 8728 2532
rect 8425 2500 8528 2510
rect 8379 2498 8528 2500
rect 8549 2498 8584 2510
rect 8218 2496 8380 2498
rect 8230 2476 8249 2496
rect 8264 2494 8294 2496
rect 8113 2468 8154 2476
rect 8236 2472 8249 2476
rect 8301 2480 8380 2496
rect 8412 2496 8584 2498
rect 8412 2480 8491 2496
rect 8498 2494 8528 2496
rect 8076 2458 8105 2468
rect 8119 2458 8148 2468
rect 8163 2458 8193 2472
rect 8236 2458 8279 2472
rect 8301 2468 8491 2480
rect 8556 2476 8562 2496
rect 8286 2458 8316 2468
rect 8317 2458 8475 2468
rect 8479 2458 8509 2468
rect 8513 2458 8543 2472
rect 8571 2458 8584 2496
rect 8656 2510 8685 2526
rect 8699 2510 8728 2526
rect 8743 2516 8773 2532
rect 8801 2510 8807 2558
rect 8810 2552 8829 2558
rect 8844 2552 8874 2560
rect 8810 2544 8874 2552
rect 8810 2528 8890 2544
rect 8906 2537 8968 2568
rect 8984 2537 9046 2568
rect 9115 2566 9164 2591
rect 9179 2566 9209 2582
rect 9078 2552 9108 2560
rect 9115 2558 9225 2566
rect 9078 2544 9123 2552
rect 8810 2526 8829 2528
rect 8844 2526 8890 2528
rect 8810 2510 8890 2526
rect 8917 2524 8952 2537
rect 8993 2534 9030 2537
rect 8993 2532 9035 2534
rect 8922 2521 8952 2524
rect 8931 2517 8938 2521
rect 8938 2516 8939 2517
rect 8897 2510 8907 2516
rect 8656 2502 8691 2510
rect 8656 2476 8657 2502
rect 8664 2476 8691 2502
rect 8599 2458 8629 2472
rect 8656 2468 8691 2476
rect 8693 2502 8734 2510
rect 8693 2476 8708 2502
rect 8715 2476 8734 2502
rect 8798 2498 8829 2510
rect 8844 2498 8947 2510
rect 8959 2500 8985 2526
rect 9000 2521 9030 2532
rect 9062 2528 9124 2544
rect 9062 2526 9108 2528
rect 9062 2510 9124 2526
rect 9136 2510 9142 2558
rect 9145 2550 9225 2558
rect 9145 2548 9164 2550
rect 9179 2548 9213 2550
rect 9145 2532 9225 2548
rect 9145 2510 9164 2532
rect 9179 2516 9209 2532
rect 9237 2526 9243 2600
rect 9252 2526 9265 2670
rect 9005 2500 9108 2510
rect 8959 2498 9108 2500
rect 9129 2498 9164 2510
rect 8798 2496 8960 2498
rect 8810 2476 8829 2496
rect 8844 2494 8874 2496
rect 8693 2468 8734 2476
rect 8816 2472 8829 2476
rect 8881 2480 8960 2496
rect 8992 2496 9164 2498
rect 8992 2480 9071 2496
rect 9078 2494 9108 2496
rect 8656 2458 8685 2468
rect 8699 2458 8728 2468
rect 8743 2458 8773 2472
rect 8816 2458 8859 2472
rect 8881 2468 9071 2480
rect 9136 2476 9142 2496
rect 8866 2458 8896 2468
rect 8897 2458 9055 2468
rect 9059 2458 9089 2468
rect 9093 2458 9123 2472
rect 9151 2458 9164 2496
rect 9236 2510 9265 2526
rect 9236 2502 9271 2510
rect 9236 2476 9237 2502
rect 9244 2476 9271 2502
rect 9179 2458 9209 2472
rect 9236 2468 9271 2476
rect 9236 2458 9265 2468
rect -1 2452 9265 2458
rect 0 2444 9265 2452
rect 15 2414 28 2444
rect 43 2430 73 2444
rect 116 2430 159 2444
rect 166 2430 386 2444
rect 393 2430 423 2444
rect 83 2416 98 2428
rect 117 2416 130 2430
rect 198 2426 351 2430
rect 80 2414 102 2416
rect 180 2414 372 2426
rect 451 2414 464 2444
rect 479 2430 509 2444
rect 546 2414 565 2444
rect 580 2414 586 2444
rect 595 2414 608 2444
rect 623 2430 653 2444
rect 696 2430 739 2444
rect 746 2430 966 2444
rect 973 2430 1003 2444
rect 663 2416 678 2428
rect 697 2416 710 2430
rect 778 2426 931 2430
rect 660 2414 682 2416
rect 760 2414 952 2426
rect 1031 2414 1044 2444
rect 1059 2430 1089 2444
rect 1126 2414 1145 2444
rect 1160 2414 1166 2444
rect 1175 2414 1188 2444
rect 1203 2430 1233 2444
rect 1276 2430 1319 2444
rect 1326 2430 1546 2444
rect 1553 2430 1583 2444
rect 1243 2416 1258 2428
rect 1277 2416 1290 2430
rect 1358 2426 1511 2430
rect 1240 2414 1262 2416
rect 1340 2414 1532 2426
rect 1611 2414 1624 2444
rect 1639 2430 1669 2444
rect 1706 2414 1725 2444
rect 1740 2414 1746 2444
rect 1755 2414 1768 2444
rect 1783 2430 1813 2444
rect 1856 2430 1899 2444
rect 1906 2430 2126 2444
rect 2133 2430 2163 2444
rect 1823 2416 1838 2428
rect 1857 2416 1870 2430
rect 1938 2426 2091 2430
rect 1820 2414 1842 2416
rect 1920 2414 2112 2426
rect 2191 2414 2204 2444
rect 2219 2430 2249 2444
rect 2286 2414 2305 2444
rect 2320 2414 2326 2444
rect 2335 2414 2348 2444
rect 2363 2430 2393 2444
rect 2436 2430 2479 2444
rect 2486 2430 2706 2444
rect 2713 2430 2743 2444
rect 2403 2416 2418 2428
rect 2437 2416 2450 2430
rect 2518 2426 2671 2430
rect 2400 2414 2422 2416
rect 2500 2414 2692 2426
rect 2771 2414 2784 2444
rect 2799 2430 2829 2444
rect 2866 2414 2885 2444
rect 2900 2414 2906 2444
rect 2915 2414 2928 2444
rect 2943 2430 2973 2444
rect 3016 2430 3059 2444
rect 3066 2430 3286 2444
rect 3293 2430 3323 2444
rect 2983 2416 2998 2428
rect 3017 2416 3030 2430
rect 3098 2426 3251 2430
rect 2980 2414 3002 2416
rect 3080 2414 3272 2426
rect 3351 2414 3364 2444
rect 3379 2430 3409 2444
rect 3446 2414 3465 2444
rect 3480 2414 3486 2444
rect 3495 2414 3508 2444
rect 3523 2430 3553 2444
rect 3596 2430 3639 2444
rect 3646 2430 3866 2444
rect 3873 2430 3903 2444
rect 3563 2416 3578 2428
rect 3597 2416 3610 2430
rect 3678 2426 3831 2430
rect 3560 2414 3582 2416
rect 3660 2414 3852 2426
rect 3931 2414 3944 2444
rect 3959 2430 3989 2444
rect 4026 2414 4045 2444
rect 4060 2414 4066 2444
rect 4075 2414 4088 2444
rect 4103 2430 4133 2444
rect 4176 2430 4219 2444
rect 4226 2430 4446 2444
rect 4453 2430 4483 2444
rect 4143 2416 4158 2428
rect 4177 2416 4190 2430
rect 4258 2426 4411 2430
rect 4140 2414 4162 2416
rect 4240 2414 4432 2426
rect 4511 2414 4524 2444
rect 4539 2430 4569 2444
rect 4606 2414 4625 2444
rect 4640 2414 4646 2444
rect 4655 2414 4668 2444
rect 4683 2430 4713 2444
rect 4756 2430 4799 2444
rect 4806 2430 5026 2444
rect 5033 2430 5063 2444
rect 4723 2416 4738 2428
rect 4757 2416 4770 2430
rect 4838 2426 4991 2430
rect 4720 2414 4742 2416
rect 4820 2414 5012 2426
rect 5091 2414 5104 2444
rect 5119 2430 5149 2444
rect 5186 2414 5205 2444
rect 5220 2414 5226 2444
rect 5235 2414 5248 2444
rect 5263 2430 5293 2444
rect 5336 2430 5379 2444
rect 5386 2430 5606 2444
rect 5613 2430 5643 2444
rect 5303 2416 5318 2428
rect 5337 2416 5350 2430
rect 5418 2426 5571 2430
rect 5300 2414 5322 2416
rect 5400 2414 5592 2426
rect 5671 2414 5684 2444
rect 5699 2430 5729 2444
rect 5766 2414 5785 2444
rect 5800 2414 5806 2444
rect 5815 2414 5828 2444
rect 5843 2430 5873 2444
rect 5916 2430 5959 2444
rect 5966 2430 6186 2444
rect 6193 2430 6223 2444
rect 5883 2416 5898 2428
rect 5917 2416 5930 2430
rect 5998 2426 6151 2430
rect 5880 2414 5902 2416
rect 5980 2414 6172 2426
rect 6251 2414 6264 2444
rect 6279 2430 6309 2444
rect 6346 2414 6365 2444
rect 6380 2414 6386 2444
rect 6395 2414 6408 2444
rect 6423 2430 6453 2444
rect 6496 2430 6539 2444
rect 6546 2430 6766 2444
rect 6773 2430 6803 2444
rect 6463 2416 6478 2428
rect 6497 2416 6510 2430
rect 6578 2426 6731 2430
rect 6460 2414 6482 2416
rect 6560 2414 6752 2426
rect 6831 2414 6844 2444
rect 6859 2430 6889 2444
rect 6926 2414 6945 2444
rect 6960 2414 6966 2444
rect 6975 2414 6988 2444
rect 7003 2430 7033 2444
rect 7076 2430 7119 2444
rect 7126 2430 7346 2444
rect 7353 2430 7383 2444
rect 7043 2416 7058 2428
rect 7077 2416 7090 2430
rect 7158 2426 7311 2430
rect 7040 2414 7062 2416
rect 7140 2414 7332 2426
rect 7411 2414 7424 2444
rect 7439 2430 7469 2444
rect 7506 2414 7525 2444
rect 7540 2414 7546 2444
rect 7555 2414 7568 2444
rect 7583 2430 7613 2444
rect 7656 2430 7699 2444
rect 7706 2430 7926 2444
rect 7933 2430 7963 2444
rect 7623 2416 7638 2428
rect 7657 2416 7670 2430
rect 7738 2426 7891 2430
rect 7620 2414 7642 2416
rect 7720 2414 7912 2426
rect 7991 2414 8004 2444
rect 8019 2430 8049 2444
rect 8086 2414 8105 2444
rect 8120 2414 8126 2444
rect 8135 2414 8148 2444
rect 8163 2430 8193 2444
rect 8236 2430 8279 2444
rect 8286 2430 8506 2444
rect 8513 2430 8543 2444
rect 8203 2416 8218 2428
rect 8237 2416 8250 2430
rect 8318 2426 8471 2430
rect 8200 2414 8222 2416
rect 8300 2414 8492 2426
rect 8571 2414 8584 2444
rect 8599 2430 8629 2444
rect 8666 2414 8685 2444
rect 8700 2414 8706 2444
rect 8715 2414 8728 2444
rect 8743 2430 8773 2444
rect 8816 2430 8859 2444
rect 8866 2430 9086 2444
rect 9093 2430 9123 2444
rect 8783 2416 8798 2428
rect 8817 2416 8830 2430
rect 8898 2426 9051 2430
rect 8780 2414 8802 2416
rect 8880 2414 9072 2426
rect 9151 2414 9164 2444
rect 9179 2430 9209 2444
rect 9252 2414 9265 2444
rect 0 2400 9265 2414
rect 15 2330 28 2400
rect 80 2396 102 2400
rect 73 2374 102 2388
rect 155 2374 171 2388
rect 209 2384 215 2386
rect 222 2384 330 2400
rect 337 2384 343 2386
rect 351 2384 366 2400
rect 432 2394 451 2397
rect 73 2372 171 2374
rect 198 2372 366 2384
rect 381 2374 397 2388
rect 432 2375 454 2394
rect 464 2388 480 2389
rect 463 2386 480 2388
rect 464 2381 480 2386
rect 454 2374 460 2375
rect 463 2374 492 2381
rect 381 2373 492 2374
rect 381 2372 498 2373
rect 57 2364 108 2372
rect 155 2364 189 2372
rect 57 2352 82 2364
rect 89 2352 108 2364
rect 162 2362 189 2364
rect 198 2362 419 2372
rect 454 2369 460 2372
rect 162 2358 419 2362
rect 57 2344 108 2352
rect 155 2344 419 2358
rect 463 2364 498 2372
rect 9 2296 28 2330
rect 73 2336 102 2344
rect 73 2330 90 2336
rect 73 2328 107 2330
rect 155 2328 171 2344
rect 172 2334 380 2344
rect 381 2334 397 2344
rect 445 2340 460 2355
rect 463 2352 464 2364
rect 471 2352 498 2364
rect 463 2344 498 2352
rect 463 2343 492 2344
rect 183 2330 397 2334
rect 198 2328 397 2330
rect 432 2330 445 2340
rect 463 2330 480 2343
rect 432 2328 480 2330
rect 74 2324 107 2328
rect 70 2322 107 2324
rect 70 2321 137 2322
rect 70 2316 101 2321
rect 107 2316 137 2321
rect 70 2312 137 2316
rect 43 2309 137 2312
rect 43 2302 92 2309
rect 43 2296 73 2302
rect 92 2297 97 2302
rect 9 2280 89 2296
rect 101 2288 137 2309
rect 198 2304 387 2328
rect 432 2327 479 2328
rect 445 2322 479 2327
rect 213 2301 387 2304
rect 206 2298 387 2301
rect 415 2321 479 2322
rect 9 2278 28 2280
rect 43 2278 77 2280
rect 9 2262 89 2278
rect 9 2256 28 2262
rect -1 2240 28 2256
rect 43 2246 73 2262
rect 101 2240 107 2288
rect 110 2282 129 2288
rect 144 2282 174 2290
rect 110 2274 174 2282
rect 110 2258 190 2274
rect 206 2267 268 2298
rect 284 2267 346 2298
rect 415 2296 464 2321
rect 479 2296 509 2312
rect 378 2282 408 2290
rect 415 2288 525 2296
rect 378 2274 423 2282
rect 110 2256 129 2258
rect 144 2256 190 2258
rect 110 2240 190 2256
rect 217 2254 252 2267
rect 293 2264 330 2267
rect 293 2262 335 2264
rect 222 2251 252 2254
rect 231 2247 238 2251
rect 238 2246 239 2247
rect 197 2240 207 2246
rect -7 2232 34 2240
rect -7 2206 8 2232
rect 15 2206 34 2232
rect 98 2228 129 2240
rect 144 2228 247 2240
rect 259 2230 285 2256
rect 300 2251 330 2262
rect 362 2258 424 2274
rect 362 2256 408 2258
rect 362 2240 424 2256
rect 436 2240 442 2288
rect 445 2280 525 2288
rect 445 2278 464 2280
rect 479 2278 513 2280
rect 445 2262 525 2278
rect 445 2240 464 2262
rect 479 2246 509 2262
rect 537 2256 543 2330
rect 546 2256 565 2400
rect 580 2256 586 2400
rect 595 2330 608 2400
rect 660 2396 682 2400
rect 653 2374 682 2388
rect 735 2374 751 2388
rect 789 2384 795 2386
rect 802 2384 910 2400
rect 917 2384 923 2386
rect 931 2384 946 2400
rect 1012 2394 1031 2397
rect 653 2372 751 2374
rect 778 2372 946 2384
rect 961 2374 977 2388
rect 1012 2375 1034 2394
rect 1044 2388 1060 2389
rect 1043 2386 1060 2388
rect 1044 2381 1060 2386
rect 1034 2374 1040 2375
rect 1043 2374 1072 2381
rect 961 2373 1072 2374
rect 961 2372 1078 2373
rect 637 2364 688 2372
rect 735 2364 769 2372
rect 637 2352 662 2364
rect 669 2352 688 2364
rect 742 2362 769 2364
rect 778 2362 999 2372
rect 1034 2369 1040 2372
rect 742 2358 999 2362
rect 637 2344 688 2352
rect 735 2344 999 2358
rect 1043 2364 1078 2372
rect 589 2296 608 2330
rect 653 2336 682 2344
rect 653 2330 670 2336
rect 653 2328 687 2330
rect 735 2328 751 2344
rect 752 2334 960 2344
rect 961 2334 977 2344
rect 1025 2340 1040 2355
rect 1043 2352 1044 2364
rect 1051 2352 1078 2364
rect 1043 2344 1078 2352
rect 1043 2343 1072 2344
rect 763 2330 977 2334
rect 778 2328 977 2330
rect 1012 2330 1025 2340
rect 1043 2330 1060 2343
rect 1012 2328 1060 2330
rect 654 2324 687 2328
rect 650 2322 687 2324
rect 650 2321 717 2322
rect 650 2316 681 2321
rect 687 2316 717 2321
rect 650 2312 717 2316
rect 623 2309 717 2312
rect 623 2302 672 2309
rect 623 2296 653 2302
rect 672 2297 677 2302
rect 589 2280 669 2296
rect 681 2288 717 2309
rect 778 2304 967 2328
rect 1012 2327 1059 2328
rect 1025 2322 1059 2327
rect 793 2301 967 2304
rect 786 2298 967 2301
rect 995 2321 1059 2322
rect 589 2278 608 2280
rect 623 2278 657 2280
rect 589 2262 669 2278
rect 589 2256 608 2262
rect 305 2230 408 2240
rect 259 2228 408 2230
rect 429 2228 464 2240
rect 98 2226 260 2228
rect 110 2206 129 2226
rect 144 2224 174 2226
rect -7 2198 34 2206
rect 116 2202 129 2206
rect 181 2210 260 2226
rect 292 2226 464 2228
rect 292 2210 371 2226
rect 378 2224 408 2226
rect -1 2188 28 2198
rect 43 2188 73 2202
rect 116 2188 159 2202
rect 181 2198 371 2210
rect 436 2206 442 2226
rect 166 2188 196 2198
rect 197 2188 355 2198
rect 359 2188 389 2198
rect 393 2188 423 2202
rect 451 2188 464 2226
rect 536 2240 565 2256
rect 579 2240 608 2256
rect 623 2246 653 2262
rect 681 2240 687 2288
rect 690 2282 709 2288
rect 724 2282 754 2290
rect 690 2274 754 2282
rect 690 2258 770 2274
rect 786 2267 848 2298
rect 864 2267 926 2298
rect 995 2296 1044 2321
rect 1059 2296 1089 2312
rect 958 2282 988 2290
rect 995 2288 1105 2296
rect 958 2274 1003 2282
rect 690 2256 709 2258
rect 724 2256 770 2258
rect 690 2240 770 2256
rect 797 2254 832 2267
rect 873 2264 910 2267
rect 873 2262 915 2264
rect 802 2251 832 2254
rect 811 2247 818 2251
rect 818 2246 819 2247
rect 777 2240 787 2246
rect 536 2232 571 2240
rect 536 2206 537 2232
rect 544 2206 571 2232
rect 479 2188 509 2202
rect 536 2198 571 2206
rect 573 2232 614 2240
rect 573 2206 588 2232
rect 595 2206 614 2232
rect 678 2228 709 2240
rect 724 2228 827 2240
rect 839 2230 865 2256
rect 880 2251 910 2262
rect 942 2258 1004 2274
rect 942 2256 988 2258
rect 942 2240 1004 2256
rect 1016 2240 1022 2288
rect 1025 2280 1105 2288
rect 1025 2278 1044 2280
rect 1059 2278 1093 2280
rect 1025 2262 1105 2278
rect 1025 2240 1044 2262
rect 1059 2246 1089 2262
rect 1117 2256 1123 2330
rect 1126 2256 1145 2400
rect 1160 2256 1166 2400
rect 1175 2330 1188 2400
rect 1240 2396 1262 2400
rect 1233 2374 1262 2388
rect 1315 2374 1331 2388
rect 1369 2384 1375 2386
rect 1382 2384 1490 2400
rect 1497 2384 1503 2386
rect 1511 2384 1526 2400
rect 1592 2394 1611 2397
rect 1233 2372 1331 2374
rect 1358 2372 1526 2384
rect 1541 2374 1557 2388
rect 1592 2375 1614 2394
rect 1624 2388 1640 2389
rect 1623 2386 1640 2388
rect 1624 2381 1640 2386
rect 1614 2374 1620 2375
rect 1623 2374 1652 2381
rect 1541 2373 1652 2374
rect 1541 2372 1658 2373
rect 1217 2364 1268 2372
rect 1315 2364 1349 2372
rect 1217 2352 1242 2364
rect 1249 2352 1268 2364
rect 1322 2362 1349 2364
rect 1358 2362 1579 2372
rect 1614 2369 1620 2372
rect 1322 2358 1579 2362
rect 1217 2344 1268 2352
rect 1315 2344 1579 2358
rect 1623 2364 1658 2372
rect 1169 2296 1188 2330
rect 1233 2336 1262 2344
rect 1233 2330 1250 2336
rect 1233 2328 1267 2330
rect 1315 2328 1331 2344
rect 1332 2334 1540 2344
rect 1541 2334 1557 2344
rect 1605 2340 1620 2355
rect 1623 2352 1624 2364
rect 1631 2352 1658 2364
rect 1623 2344 1658 2352
rect 1623 2343 1652 2344
rect 1343 2330 1557 2334
rect 1358 2328 1557 2330
rect 1592 2330 1605 2340
rect 1623 2330 1640 2343
rect 1592 2328 1640 2330
rect 1234 2324 1267 2328
rect 1230 2322 1267 2324
rect 1230 2321 1297 2322
rect 1230 2316 1261 2321
rect 1267 2316 1297 2321
rect 1230 2312 1297 2316
rect 1203 2309 1297 2312
rect 1203 2302 1252 2309
rect 1203 2296 1233 2302
rect 1252 2297 1257 2302
rect 1169 2280 1249 2296
rect 1261 2288 1297 2309
rect 1358 2304 1547 2328
rect 1592 2327 1639 2328
rect 1605 2322 1639 2327
rect 1373 2301 1547 2304
rect 1366 2298 1547 2301
rect 1575 2321 1639 2322
rect 1169 2278 1188 2280
rect 1203 2278 1237 2280
rect 1169 2262 1249 2278
rect 1169 2256 1188 2262
rect 885 2230 988 2240
rect 839 2228 988 2230
rect 1009 2228 1044 2240
rect 678 2226 840 2228
rect 690 2206 709 2226
rect 724 2224 754 2226
rect 573 2198 614 2206
rect 696 2202 709 2206
rect 761 2210 840 2226
rect 872 2226 1044 2228
rect 872 2210 951 2226
rect 958 2224 988 2226
rect 536 2188 565 2198
rect 579 2188 608 2198
rect 623 2188 653 2202
rect 696 2188 739 2202
rect 761 2198 951 2210
rect 1016 2206 1022 2226
rect 746 2188 776 2198
rect 777 2188 935 2198
rect 939 2188 969 2198
rect 973 2188 1003 2202
rect 1031 2188 1044 2226
rect 1116 2240 1145 2256
rect 1159 2240 1188 2256
rect 1203 2246 1233 2262
rect 1261 2240 1267 2288
rect 1270 2282 1289 2288
rect 1304 2282 1334 2290
rect 1270 2274 1334 2282
rect 1270 2258 1350 2274
rect 1366 2267 1428 2298
rect 1444 2267 1506 2298
rect 1575 2296 1624 2321
rect 1639 2296 1669 2312
rect 1538 2282 1568 2290
rect 1575 2288 1685 2296
rect 1538 2274 1583 2282
rect 1270 2256 1289 2258
rect 1304 2256 1350 2258
rect 1270 2240 1350 2256
rect 1377 2254 1412 2267
rect 1453 2264 1490 2267
rect 1453 2262 1495 2264
rect 1382 2251 1412 2254
rect 1391 2247 1398 2251
rect 1398 2246 1399 2247
rect 1357 2240 1367 2246
rect 1116 2232 1151 2240
rect 1116 2206 1117 2232
rect 1124 2206 1151 2232
rect 1059 2188 1089 2202
rect 1116 2198 1151 2206
rect 1153 2232 1194 2240
rect 1153 2206 1168 2232
rect 1175 2206 1194 2232
rect 1258 2228 1289 2240
rect 1304 2228 1407 2240
rect 1419 2230 1445 2256
rect 1460 2251 1490 2262
rect 1522 2258 1584 2274
rect 1522 2256 1568 2258
rect 1522 2240 1584 2256
rect 1596 2240 1602 2288
rect 1605 2280 1685 2288
rect 1605 2278 1624 2280
rect 1639 2278 1673 2280
rect 1605 2262 1685 2278
rect 1605 2240 1624 2262
rect 1639 2246 1669 2262
rect 1697 2256 1703 2330
rect 1706 2256 1725 2400
rect 1740 2256 1746 2400
rect 1755 2330 1768 2400
rect 1820 2396 1842 2400
rect 1813 2374 1842 2388
rect 1895 2374 1911 2388
rect 1949 2384 1955 2386
rect 1962 2384 2070 2400
rect 2077 2384 2083 2386
rect 2091 2384 2106 2400
rect 2172 2394 2191 2397
rect 1813 2372 1911 2374
rect 1938 2372 2106 2384
rect 2121 2374 2137 2388
rect 2172 2375 2194 2394
rect 2204 2388 2220 2389
rect 2203 2386 2220 2388
rect 2204 2381 2220 2386
rect 2194 2374 2200 2375
rect 2203 2374 2232 2381
rect 2121 2373 2232 2374
rect 2121 2372 2238 2373
rect 1797 2364 1848 2372
rect 1895 2364 1929 2372
rect 1797 2352 1822 2364
rect 1829 2352 1848 2364
rect 1902 2362 1929 2364
rect 1938 2362 2159 2372
rect 2194 2369 2200 2372
rect 1902 2358 2159 2362
rect 1797 2344 1848 2352
rect 1895 2344 2159 2358
rect 2203 2364 2238 2372
rect 1749 2296 1768 2330
rect 1813 2336 1842 2344
rect 1813 2330 1830 2336
rect 1813 2328 1847 2330
rect 1895 2328 1911 2344
rect 1912 2334 2120 2344
rect 2121 2334 2137 2344
rect 2185 2340 2200 2355
rect 2203 2352 2204 2364
rect 2211 2352 2238 2364
rect 2203 2344 2238 2352
rect 2203 2343 2232 2344
rect 1923 2330 2137 2334
rect 1938 2328 2137 2330
rect 2172 2330 2185 2340
rect 2203 2330 2220 2343
rect 2172 2328 2220 2330
rect 1814 2324 1847 2328
rect 1810 2322 1847 2324
rect 1810 2321 1877 2322
rect 1810 2316 1841 2321
rect 1847 2316 1877 2321
rect 1810 2312 1877 2316
rect 1783 2309 1877 2312
rect 1783 2302 1832 2309
rect 1783 2296 1813 2302
rect 1832 2297 1837 2302
rect 1749 2280 1829 2296
rect 1841 2288 1877 2309
rect 1938 2304 2127 2328
rect 2172 2327 2219 2328
rect 2185 2322 2219 2327
rect 1953 2301 2127 2304
rect 1946 2298 2127 2301
rect 2155 2321 2219 2322
rect 1749 2278 1768 2280
rect 1783 2278 1817 2280
rect 1749 2262 1829 2278
rect 1749 2256 1768 2262
rect 1465 2230 1568 2240
rect 1419 2228 1568 2230
rect 1589 2228 1624 2240
rect 1258 2226 1420 2228
rect 1270 2206 1289 2226
rect 1304 2224 1334 2226
rect 1153 2198 1194 2206
rect 1276 2202 1289 2206
rect 1341 2210 1420 2226
rect 1452 2226 1624 2228
rect 1452 2210 1531 2226
rect 1538 2224 1568 2226
rect 1116 2188 1145 2198
rect 1159 2188 1188 2198
rect 1203 2188 1233 2202
rect 1276 2188 1319 2202
rect 1341 2198 1531 2210
rect 1596 2206 1602 2226
rect 1326 2188 1356 2198
rect 1357 2188 1515 2198
rect 1519 2188 1549 2198
rect 1553 2188 1583 2202
rect 1611 2188 1624 2226
rect 1696 2240 1725 2256
rect 1739 2240 1768 2256
rect 1783 2246 1813 2262
rect 1841 2240 1847 2288
rect 1850 2282 1869 2288
rect 1884 2282 1914 2290
rect 1850 2274 1914 2282
rect 1850 2258 1930 2274
rect 1946 2267 2008 2298
rect 2024 2267 2086 2298
rect 2155 2296 2204 2321
rect 2219 2296 2249 2312
rect 2118 2282 2148 2290
rect 2155 2288 2265 2296
rect 2118 2274 2163 2282
rect 1850 2256 1869 2258
rect 1884 2256 1930 2258
rect 1850 2240 1930 2256
rect 1957 2254 1992 2267
rect 2033 2264 2070 2267
rect 2033 2262 2075 2264
rect 1962 2251 1992 2254
rect 1971 2247 1978 2251
rect 1978 2246 1979 2247
rect 1937 2240 1947 2246
rect 1696 2232 1731 2240
rect 1696 2206 1697 2232
rect 1704 2206 1731 2232
rect 1639 2188 1669 2202
rect 1696 2198 1731 2206
rect 1733 2232 1774 2240
rect 1733 2206 1748 2232
rect 1755 2206 1774 2232
rect 1838 2228 1869 2240
rect 1884 2228 1987 2240
rect 1999 2230 2025 2256
rect 2040 2251 2070 2262
rect 2102 2258 2164 2274
rect 2102 2256 2148 2258
rect 2102 2240 2164 2256
rect 2176 2240 2182 2288
rect 2185 2280 2265 2288
rect 2185 2278 2204 2280
rect 2219 2278 2253 2280
rect 2185 2262 2265 2278
rect 2185 2240 2204 2262
rect 2219 2246 2249 2262
rect 2277 2256 2283 2330
rect 2286 2256 2305 2400
rect 2320 2256 2326 2400
rect 2335 2330 2348 2400
rect 2400 2396 2422 2400
rect 2393 2374 2422 2388
rect 2475 2374 2491 2388
rect 2529 2384 2535 2386
rect 2542 2384 2650 2400
rect 2657 2384 2663 2386
rect 2671 2384 2686 2400
rect 2752 2394 2771 2397
rect 2393 2372 2491 2374
rect 2518 2372 2686 2384
rect 2701 2374 2717 2388
rect 2752 2375 2774 2394
rect 2784 2388 2800 2389
rect 2783 2386 2800 2388
rect 2784 2381 2800 2386
rect 2774 2374 2780 2375
rect 2783 2374 2812 2381
rect 2701 2373 2812 2374
rect 2701 2372 2818 2373
rect 2377 2364 2428 2372
rect 2475 2364 2509 2372
rect 2377 2352 2402 2364
rect 2409 2352 2428 2364
rect 2482 2362 2509 2364
rect 2518 2362 2739 2372
rect 2774 2369 2780 2372
rect 2482 2358 2739 2362
rect 2377 2344 2428 2352
rect 2475 2344 2739 2358
rect 2783 2364 2818 2372
rect 2329 2296 2348 2330
rect 2393 2336 2422 2344
rect 2393 2330 2410 2336
rect 2393 2328 2427 2330
rect 2475 2328 2491 2344
rect 2492 2334 2700 2344
rect 2701 2334 2717 2344
rect 2765 2340 2780 2355
rect 2783 2352 2784 2364
rect 2791 2352 2818 2364
rect 2783 2344 2818 2352
rect 2783 2343 2812 2344
rect 2503 2330 2717 2334
rect 2518 2328 2717 2330
rect 2752 2330 2765 2340
rect 2783 2330 2800 2343
rect 2752 2328 2800 2330
rect 2394 2324 2427 2328
rect 2390 2322 2427 2324
rect 2390 2321 2457 2322
rect 2390 2316 2421 2321
rect 2427 2316 2457 2321
rect 2390 2312 2457 2316
rect 2363 2309 2457 2312
rect 2363 2302 2412 2309
rect 2363 2296 2393 2302
rect 2412 2297 2417 2302
rect 2329 2280 2409 2296
rect 2421 2288 2457 2309
rect 2518 2304 2707 2328
rect 2752 2327 2799 2328
rect 2765 2322 2799 2327
rect 2533 2301 2707 2304
rect 2526 2298 2707 2301
rect 2735 2321 2799 2322
rect 2329 2278 2348 2280
rect 2363 2278 2397 2280
rect 2329 2262 2409 2278
rect 2329 2256 2348 2262
rect 2045 2230 2148 2240
rect 1999 2228 2148 2230
rect 2169 2228 2204 2240
rect 1838 2226 2000 2228
rect 1850 2206 1869 2226
rect 1884 2224 1914 2226
rect 1733 2198 1774 2206
rect 1856 2202 1869 2206
rect 1921 2210 2000 2226
rect 2032 2226 2204 2228
rect 2032 2210 2111 2226
rect 2118 2224 2148 2226
rect 1696 2188 1725 2198
rect 1739 2188 1768 2198
rect 1783 2188 1813 2202
rect 1856 2188 1899 2202
rect 1921 2198 2111 2210
rect 2176 2206 2182 2226
rect 1906 2188 1936 2198
rect 1937 2188 2095 2198
rect 2099 2188 2129 2198
rect 2133 2188 2163 2202
rect 2191 2188 2204 2226
rect 2276 2240 2305 2256
rect 2319 2240 2348 2256
rect 2363 2246 2393 2262
rect 2421 2240 2427 2288
rect 2430 2282 2449 2288
rect 2464 2282 2494 2290
rect 2430 2274 2494 2282
rect 2430 2258 2510 2274
rect 2526 2267 2588 2298
rect 2604 2267 2666 2298
rect 2735 2296 2784 2321
rect 2799 2296 2829 2312
rect 2698 2282 2728 2290
rect 2735 2288 2845 2296
rect 2698 2274 2743 2282
rect 2430 2256 2449 2258
rect 2464 2256 2510 2258
rect 2430 2240 2510 2256
rect 2537 2254 2572 2267
rect 2613 2264 2650 2267
rect 2613 2262 2655 2264
rect 2542 2251 2572 2254
rect 2551 2247 2558 2251
rect 2558 2246 2559 2247
rect 2517 2240 2527 2246
rect 2276 2232 2311 2240
rect 2276 2206 2277 2232
rect 2284 2206 2311 2232
rect 2219 2188 2249 2202
rect 2276 2198 2311 2206
rect 2313 2232 2354 2240
rect 2313 2206 2328 2232
rect 2335 2206 2354 2232
rect 2418 2228 2449 2240
rect 2464 2228 2567 2240
rect 2579 2230 2605 2256
rect 2620 2251 2650 2262
rect 2682 2258 2744 2274
rect 2682 2256 2728 2258
rect 2682 2240 2744 2256
rect 2756 2240 2762 2288
rect 2765 2280 2845 2288
rect 2765 2278 2784 2280
rect 2799 2278 2833 2280
rect 2765 2262 2845 2278
rect 2765 2240 2784 2262
rect 2799 2246 2829 2262
rect 2857 2256 2863 2330
rect 2866 2256 2885 2400
rect 2900 2256 2906 2400
rect 2915 2330 2928 2400
rect 2980 2396 3002 2400
rect 2973 2374 3002 2388
rect 3055 2374 3071 2388
rect 3109 2384 3115 2386
rect 3122 2384 3230 2400
rect 3237 2384 3243 2386
rect 3251 2384 3266 2400
rect 3332 2394 3351 2397
rect 2973 2372 3071 2374
rect 3098 2372 3266 2384
rect 3281 2374 3297 2388
rect 3332 2375 3354 2394
rect 3364 2388 3380 2389
rect 3363 2386 3380 2388
rect 3364 2381 3380 2386
rect 3354 2374 3360 2375
rect 3363 2374 3392 2381
rect 3281 2373 3392 2374
rect 3281 2372 3398 2373
rect 2957 2364 3008 2372
rect 3055 2364 3089 2372
rect 2957 2352 2982 2364
rect 2989 2352 3008 2364
rect 3062 2362 3089 2364
rect 3098 2362 3319 2372
rect 3354 2369 3360 2372
rect 3062 2358 3319 2362
rect 2957 2344 3008 2352
rect 3055 2344 3319 2358
rect 3363 2364 3398 2372
rect 2909 2296 2928 2330
rect 2973 2336 3002 2344
rect 2973 2330 2990 2336
rect 2973 2328 3007 2330
rect 3055 2328 3071 2344
rect 3072 2334 3280 2344
rect 3281 2334 3297 2344
rect 3345 2340 3360 2355
rect 3363 2352 3364 2364
rect 3371 2352 3398 2364
rect 3363 2344 3398 2352
rect 3363 2343 3392 2344
rect 3083 2330 3297 2334
rect 3098 2328 3297 2330
rect 3332 2330 3345 2340
rect 3363 2330 3380 2343
rect 3332 2328 3380 2330
rect 2974 2324 3007 2328
rect 2970 2322 3007 2324
rect 2970 2321 3037 2322
rect 2970 2316 3001 2321
rect 3007 2316 3037 2321
rect 2970 2312 3037 2316
rect 2943 2309 3037 2312
rect 2943 2302 2992 2309
rect 2943 2296 2973 2302
rect 2992 2297 2997 2302
rect 2909 2280 2989 2296
rect 3001 2288 3037 2309
rect 3098 2304 3287 2328
rect 3332 2327 3379 2328
rect 3345 2322 3379 2327
rect 3113 2301 3287 2304
rect 3106 2298 3287 2301
rect 3315 2321 3379 2322
rect 2909 2278 2928 2280
rect 2943 2278 2977 2280
rect 2909 2262 2989 2278
rect 2909 2256 2928 2262
rect 2625 2230 2728 2240
rect 2579 2228 2728 2230
rect 2749 2228 2784 2240
rect 2418 2226 2580 2228
rect 2430 2206 2449 2226
rect 2464 2224 2494 2226
rect 2313 2198 2354 2206
rect 2436 2202 2449 2206
rect 2501 2210 2580 2226
rect 2612 2226 2784 2228
rect 2612 2210 2691 2226
rect 2698 2224 2728 2226
rect 2276 2188 2305 2198
rect 2319 2188 2348 2198
rect 2363 2188 2393 2202
rect 2436 2188 2479 2202
rect 2501 2198 2691 2210
rect 2756 2206 2762 2226
rect 2486 2188 2516 2198
rect 2517 2188 2675 2198
rect 2679 2188 2709 2198
rect 2713 2188 2743 2202
rect 2771 2188 2784 2226
rect 2856 2240 2885 2256
rect 2899 2240 2928 2256
rect 2943 2246 2973 2262
rect 3001 2240 3007 2288
rect 3010 2282 3029 2288
rect 3044 2282 3074 2290
rect 3010 2274 3074 2282
rect 3010 2258 3090 2274
rect 3106 2267 3168 2298
rect 3184 2267 3246 2298
rect 3315 2296 3364 2321
rect 3379 2296 3409 2312
rect 3278 2282 3308 2290
rect 3315 2288 3425 2296
rect 3278 2274 3323 2282
rect 3010 2256 3029 2258
rect 3044 2256 3090 2258
rect 3010 2240 3090 2256
rect 3117 2254 3152 2267
rect 3193 2264 3230 2267
rect 3193 2262 3235 2264
rect 3122 2251 3152 2254
rect 3131 2247 3138 2251
rect 3138 2246 3139 2247
rect 3097 2240 3107 2246
rect 2856 2232 2891 2240
rect 2856 2206 2857 2232
rect 2864 2206 2891 2232
rect 2799 2188 2829 2202
rect 2856 2198 2891 2206
rect 2893 2232 2934 2240
rect 2893 2206 2908 2232
rect 2915 2206 2934 2232
rect 2998 2228 3029 2240
rect 3044 2228 3147 2240
rect 3159 2230 3185 2256
rect 3200 2251 3230 2262
rect 3262 2258 3324 2274
rect 3262 2256 3308 2258
rect 3262 2240 3324 2256
rect 3336 2240 3342 2288
rect 3345 2280 3425 2288
rect 3345 2278 3364 2280
rect 3379 2278 3413 2280
rect 3345 2262 3425 2278
rect 3345 2240 3364 2262
rect 3379 2246 3409 2262
rect 3437 2256 3443 2330
rect 3446 2256 3465 2400
rect 3480 2256 3486 2400
rect 3495 2330 3508 2400
rect 3560 2396 3582 2400
rect 3553 2374 3582 2388
rect 3635 2374 3651 2388
rect 3689 2384 3695 2386
rect 3702 2384 3810 2400
rect 3817 2384 3823 2386
rect 3831 2384 3846 2400
rect 3912 2394 3931 2397
rect 3553 2372 3651 2374
rect 3678 2372 3846 2384
rect 3861 2374 3877 2388
rect 3912 2375 3934 2394
rect 3944 2388 3960 2389
rect 3943 2386 3960 2388
rect 3944 2381 3960 2386
rect 3934 2374 3940 2375
rect 3943 2374 3972 2381
rect 3861 2373 3972 2374
rect 3861 2372 3978 2373
rect 3537 2364 3588 2372
rect 3635 2364 3669 2372
rect 3537 2352 3562 2364
rect 3569 2352 3588 2364
rect 3642 2362 3669 2364
rect 3678 2362 3899 2372
rect 3934 2369 3940 2372
rect 3642 2358 3899 2362
rect 3537 2344 3588 2352
rect 3635 2344 3899 2358
rect 3943 2364 3978 2372
rect 3489 2296 3508 2330
rect 3553 2336 3582 2344
rect 3553 2330 3570 2336
rect 3553 2328 3587 2330
rect 3635 2328 3651 2344
rect 3652 2334 3860 2344
rect 3861 2334 3877 2344
rect 3925 2340 3940 2355
rect 3943 2352 3944 2364
rect 3951 2352 3978 2364
rect 3943 2344 3978 2352
rect 3943 2343 3972 2344
rect 3663 2330 3877 2334
rect 3678 2328 3877 2330
rect 3912 2330 3925 2340
rect 3943 2330 3960 2343
rect 3912 2328 3960 2330
rect 3554 2324 3587 2328
rect 3550 2322 3587 2324
rect 3550 2321 3617 2322
rect 3550 2316 3581 2321
rect 3587 2316 3617 2321
rect 3550 2312 3617 2316
rect 3523 2309 3617 2312
rect 3523 2302 3572 2309
rect 3523 2296 3553 2302
rect 3572 2297 3577 2302
rect 3489 2280 3569 2296
rect 3581 2288 3617 2309
rect 3678 2304 3867 2328
rect 3912 2327 3959 2328
rect 3925 2322 3959 2327
rect 3693 2301 3867 2304
rect 3686 2298 3867 2301
rect 3895 2321 3959 2322
rect 3489 2278 3508 2280
rect 3523 2278 3557 2280
rect 3489 2262 3569 2278
rect 3489 2256 3508 2262
rect 3205 2230 3308 2240
rect 3159 2228 3308 2230
rect 3329 2228 3364 2240
rect 2998 2226 3160 2228
rect 3010 2206 3029 2226
rect 3044 2224 3074 2226
rect 2893 2198 2934 2206
rect 3016 2202 3029 2206
rect 3081 2210 3160 2226
rect 3192 2226 3364 2228
rect 3192 2210 3271 2226
rect 3278 2224 3308 2226
rect 2856 2188 2885 2198
rect 2899 2188 2928 2198
rect 2943 2188 2973 2202
rect 3016 2188 3059 2202
rect 3081 2198 3271 2210
rect 3336 2206 3342 2226
rect 3066 2188 3096 2198
rect 3097 2188 3255 2198
rect 3259 2188 3289 2198
rect 3293 2188 3323 2202
rect 3351 2188 3364 2226
rect 3436 2240 3465 2256
rect 3479 2240 3508 2256
rect 3523 2246 3553 2262
rect 3581 2240 3587 2288
rect 3590 2282 3609 2288
rect 3624 2282 3654 2290
rect 3590 2274 3654 2282
rect 3590 2258 3670 2274
rect 3686 2267 3748 2298
rect 3764 2267 3826 2298
rect 3895 2296 3944 2321
rect 3959 2296 3989 2312
rect 3858 2282 3888 2290
rect 3895 2288 4005 2296
rect 3858 2274 3903 2282
rect 3590 2256 3609 2258
rect 3624 2256 3670 2258
rect 3590 2240 3670 2256
rect 3697 2254 3732 2267
rect 3773 2264 3810 2267
rect 3773 2262 3815 2264
rect 3702 2251 3732 2254
rect 3711 2247 3718 2251
rect 3718 2246 3719 2247
rect 3677 2240 3687 2246
rect 3436 2232 3471 2240
rect 3436 2206 3437 2232
rect 3444 2206 3471 2232
rect 3379 2188 3409 2202
rect 3436 2198 3471 2206
rect 3473 2232 3514 2240
rect 3473 2206 3488 2232
rect 3495 2206 3514 2232
rect 3578 2228 3609 2240
rect 3624 2228 3727 2240
rect 3739 2230 3765 2256
rect 3780 2251 3810 2262
rect 3842 2258 3904 2274
rect 3842 2256 3888 2258
rect 3842 2240 3904 2256
rect 3916 2240 3922 2288
rect 3925 2280 4005 2288
rect 3925 2278 3944 2280
rect 3959 2278 3993 2280
rect 3925 2262 4005 2278
rect 3925 2240 3944 2262
rect 3959 2246 3989 2262
rect 4017 2256 4023 2330
rect 4026 2256 4045 2400
rect 4060 2256 4066 2400
rect 4075 2330 4088 2400
rect 4140 2396 4162 2400
rect 4133 2374 4162 2388
rect 4215 2374 4231 2388
rect 4269 2384 4275 2386
rect 4282 2384 4390 2400
rect 4397 2384 4403 2386
rect 4411 2384 4426 2400
rect 4492 2394 4511 2397
rect 4133 2372 4231 2374
rect 4258 2372 4426 2384
rect 4441 2374 4457 2388
rect 4492 2375 4514 2394
rect 4524 2388 4540 2389
rect 4523 2386 4540 2388
rect 4524 2381 4540 2386
rect 4514 2374 4520 2375
rect 4523 2374 4552 2381
rect 4441 2373 4552 2374
rect 4441 2372 4558 2373
rect 4117 2364 4168 2372
rect 4215 2364 4249 2372
rect 4117 2352 4142 2364
rect 4149 2352 4168 2364
rect 4222 2362 4249 2364
rect 4258 2362 4479 2372
rect 4514 2369 4520 2372
rect 4222 2358 4479 2362
rect 4117 2344 4168 2352
rect 4215 2344 4479 2358
rect 4523 2364 4558 2372
rect 4069 2296 4088 2330
rect 4133 2336 4162 2344
rect 4133 2330 4150 2336
rect 4133 2328 4167 2330
rect 4215 2328 4231 2344
rect 4232 2334 4440 2344
rect 4441 2334 4457 2344
rect 4505 2340 4520 2355
rect 4523 2352 4524 2364
rect 4531 2352 4558 2364
rect 4523 2344 4558 2352
rect 4523 2343 4552 2344
rect 4243 2330 4457 2334
rect 4258 2328 4457 2330
rect 4492 2330 4505 2340
rect 4523 2330 4540 2343
rect 4492 2328 4540 2330
rect 4134 2324 4167 2328
rect 4130 2322 4167 2324
rect 4130 2321 4197 2322
rect 4130 2316 4161 2321
rect 4167 2316 4197 2321
rect 4130 2312 4197 2316
rect 4103 2309 4197 2312
rect 4103 2302 4152 2309
rect 4103 2296 4133 2302
rect 4152 2297 4157 2302
rect 4069 2280 4149 2296
rect 4161 2288 4197 2309
rect 4258 2304 4447 2328
rect 4492 2327 4539 2328
rect 4505 2322 4539 2327
rect 4273 2301 4447 2304
rect 4266 2298 4447 2301
rect 4475 2321 4539 2322
rect 4069 2278 4088 2280
rect 4103 2278 4137 2280
rect 4069 2262 4149 2278
rect 4069 2256 4088 2262
rect 3785 2230 3888 2240
rect 3739 2228 3888 2230
rect 3909 2228 3944 2240
rect 3578 2226 3740 2228
rect 3590 2206 3609 2226
rect 3624 2224 3654 2226
rect 3473 2198 3514 2206
rect 3596 2202 3609 2206
rect 3661 2210 3740 2226
rect 3772 2226 3944 2228
rect 3772 2210 3851 2226
rect 3858 2224 3888 2226
rect 3436 2188 3465 2198
rect 3479 2188 3508 2198
rect 3523 2188 3553 2202
rect 3596 2188 3639 2202
rect 3661 2198 3851 2210
rect 3916 2206 3922 2226
rect 3646 2188 3676 2198
rect 3677 2188 3835 2198
rect 3839 2188 3869 2198
rect 3873 2188 3903 2202
rect 3931 2188 3944 2226
rect 4016 2240 4045 2256
rect 4059 2240 4088 2256
rect 4103 2246 4133 2262
rect 4161 2240 4167 2288
rect 4170 2282 4189 2288
rect 4204 2282 4234 2290
rect 4170 2274 4234 2282
rect 4170 2258 4250 2274
rect 4266 2267 4328 2298
rect 4344 2267 4406 2298
rect 4475 2296 4524 2321
rect 4539 2296 4569 2312
rect 4438 2282 4468 2290
rect 4475 2288 4585 2296
rect 4438 2274 4483 2282
rect 4170 2256 4189 2258
rect 4204 2256 4250 2258
rect 4170 2240 4250 2256
rect 4277 2254 4312 2267
rect 4353 2264 4390 2267
rect 4353 2262 4395 2264
rect 4282 2251 4312 2254
rect 4291 2247 4298 2251
rect 4298 2246 4299 2247
rect 4257 2240 4267 2246
rect 4016 2232 4051 2240
rect 4016 2206 4017 2232
rect 4024 2206 4051 2232
rect 3959 2188 3989 2202
rect 4016 2198 4051 2206
rect 4053 2232 4094 2240
rect 4053 2206 4068 2232
rect 4075 2206 4094 2232
rect 4158 2228 4189 2240
rect 4204 2228 4307 2240
rect 4319 2230 4345 2256
rect 4360 2251 4390 2262
rect 4422 2258 4484 2274
rect 4422 2256 4468 2258
rect 4422 2240 4484 2256
rect 4496 2240 4502 2288
rect 4505 2280 4585 2288
rect 4505 2278 4524 2280
rect 4539 2278 4573 2280
rect 4505 2262 4585 2278
rect 4505 2240 4524 2262
rect 4539 2246 4569 2262
rect 4597 2256 4603 2330
rect 4606 2256 4625 2400
rect 4640 2256 4646 2400
rect 4655 2330 4668 2400
rect 4720 2396 4742 2400
rect 4713 2374 4742 2388
rect 4795 2374 4811 2388
rect 4849 2384 4855 2386
rect 4862 2384 4970 2400
rect 4977 2384 4983 2386
rect 4991 2384 5006 2400
rect 5072 2394 5091 2397
rect 4713 2372 4811 2374
rect 4838 2372 5006 2384
rect 5021 2374 5037 2388
rect 5072 2375 5094 2394
rect 5104 2388 5120 2389
rect 5103 2386 5120 2388
rect 5104 2381 5120 2386
rect 5094 2374 5100 2375
rect 5103 2374 5132 2381
rect 5021 2373 5132 2374
rect 5021 2372 5138 2373
rect 4697 2364 4748 2372
rect 4795 2364 4829 2372
rect 4697 2352 4722 2364
rect 4729 2352 4748 2364
rect 4802 2362 4829 2364
rect 4838 2362 5059 2372
rect 5094 2369 5100 2372
rect 4802 2358 5059 2362
rect 4697 2344 4748 2352
rect 4795 2344 5059 2358
rect 5103 2364 5138 2372
rect 4649 2296 4668 2330
rect 4713 2336 4742 2344
rect 4713 2330 4730 2336
rect 4713 2328 4747 2330
rect 4795 2328 4811 2344
rect 4812 2334 5020 2344
rect 5021 2334 5037 2344
rect 5085 2340 5100 2355
rect 5103 2352 5104 2364
rect 5111 2352 5138 2364
rect 5103 2344 5138 2352
rect 5103 2343 5132 2344
rect 4823 2330 5037 2334
rect 4838 2328 5037 2330
rect 5072 2330 5085 2340
rect 5103 2330 5120 2343
rect 5072 2328 5120 2330
rect 4714 2324 4747 2328
rect 4710 2322 4747 2324
rect 4710 2321 4777 2322
rect 4710 2316 4741 2321
rect 4747 2316 4777 2321
rect 4710 2312 4777 2316
rect 4683 2309 4777 2312
rect 4683 2302 4732 2309
rect 4683 2296 4713 2302
rect 4732 2297 4737 2302
rect 4649 2280 4729 2296
rect 4741 2288 4777 2309
rect 4838 2304 5027 2328
rect 5072 2327 5119 2328
rect 5085 2322 5119 2327
rect 4853 2301 5027 2304
rect 4846 2298 5027 2301
rect 5055 2321 5119 2322
rect 4649 2278 4668 2280
rect 4683 2278 4717 2280
rect 4649 2262 4729 2278
rect 4649 2256 4668 2262
rect 4365 2230 4468 2240
rect 4319 2228 4468 2230
rect 4489 2228 4524 2240
rect 4158 2226 4320 2228
rect 4170 2206 4189 2226
rect 4204 2224 4234 2226
rect 4053 2198 4094 2206
rect 4176 2202 4189 2206
rect 4241 2210 4320 2226
rect 4352 2226 4524 2228
rect 4352 2210 4431 2226
rect 4438 2224 4468 2226
rect 4016 2188 4045 2198
rect 4059 2188 4088 2198
rect 4103 2188 4133 2202
rect 4176 2188 4219 2202
rect 4241 2198 4431 2210
rect 4496 2206 4502 2226
rect 4226 2188 4256 2198
rect 4257 2188 4415 2198
rect 4419 2188 4449 2198
rect 4453 2188 4483 2202
rect 4511 2188 4524 2226
rect 4596 2240 4625 2256
rect 4639 2240 4668 2256
rect 4683 2246 4713 2262
rect 4741 2240 4747 2288
rect 4750 2282 4769 2288
rect 4784 2282 4814 2290
rect 4750 2274 4814 2282
rect 4750 2258 4830 2274
rect 4846 2267 4908 2298
rect 4924 2267 4986 2298
rect 5055 2296 5104 2321
rect 5119 2296 5149 2312
rect 5018 2282 5048 2290
rect 5055 2288 5165 2296
rect 5018 2274 5063 2282
rect 4750 2256 4769 2258
rect 4784 2256 4830 2258
rect 4750 2240 4830 2256
rect 4857 2254 4892 2267
rect 4933 2264 4970 2267
rect 4933 2262 4975 2264
rect 4862 2251 4892 2254
rect 4871 2247 4878 2251
rect 4878 2246 4879 2247
rect 4837 2240 4847 2246
rect 4596 2232 4631 2240
rect 4596 2206 4597 2232
rect 4604 2206 4631 2232
rect 4539 2188 4569 2202
rect 4596 2198 4631 2206
rect 4633 2232 4674 2240
rect 4633 2206 4648 2232
rect 4655 2206 4674 2232
rect 4738 2228 4769 2240
rect 4784 2228 4887 2240
rect 4899 2230 4925 2256
rect 4940 2251 4970 2262
rect 5002 2258 5064 2274
rect 5002 2256 5048 2258
rect 5002 2240 5064 2256
rect 5076 2240 5082 2288
rect 5085 2280 5165 2288
rect 5085 2278 5104 2280
rect 5119 2278 5153 2280
rect 5085 2262 5165 2278
rect 5085 2240 5104 2262
rect 5119 2246 5149 2262
rect 5177 2256 5183 2330
rect 5186 2256 5205 2400
rect 5220 2256 5226 2400
rect 5235 2330 5248 2400
rect 5300 2396 5322 2400
rect 5293 2374 5322 2388
rect 5375 2374 5391 2388
rect 5429 2384 5435 2386
rect 5442 2384 5550 2400
rect 5557 2384 5563 2386
rect 5571 2384 5586 2400
rect 5652 2394 5671 2397
rect 5293 2372 5391 2374
rect 5418 2372 5586 2384
rect 5601 2374 5617 2388
rect 5652 2375 5674 2394
rect 5684 2388 5700 2389
rect 5683 2386 5700 2388
rect 5684 2381 5700 2386
rect 5674 2374 5680 2375
rect 5683 2374 5712 2381
rect 5601 2373 5712 2374
rect 5601 2372 5718 2373
rect 5277 2364 5328 2372
rect 5375 2364 5409 2372
rect 5277 2352 5302 2364
rect 5309 2352 5328 2364
rect 5382 2362 5409 2364
rect 5418 2362 5639 2372
rect 5674 2369 5680 2372
rect 5382 2358 5639 2362
rect 5277 2344 5328 2352
rect 5375 2344 5639 2358
rect 5683 2364 5718 2372
rect 5229 2296 5248 2330
rect 5293 2336 5322 2344
rect 5293 2330 5310 2336
rect 5293 2328 5327 2330
rect 5375 2328 5391 2344
rect 5392 2334 5600 2344
rect 5601 2334 5617 2344
rect 5665 2340 5680 2355
rect 5683 2352 5684 2364
rect 5691 2352 5718 2364
rect 5683 2344 5718 2352
rect 5683 2343 5712 2344
rect 5403 2330 5617 2334
rect 5418 2328 5617 2330
rect 5652 2330 5665 2340
rect 5683 2330 5700 2343
rect 5652 2328 5700 2330
rect 5294 2324 5327 2328
rect 5290 2322 5327 2324
rect 5290 2321 5357 2322
rect 5290 2316 5321 2321
rect 5327 2316 5357 2321
rect 5290 2312 5357 2316
rect 5263 2309 5357 2312
rect 5263 2302 5312 2309
rect 5263 2296 5293 2302
rect 5312 2297 5317 2302
rect 5229 2280 5309 2296
rect 5321 2288 5357 2309
rect 5418 2304 5607 2328
rect 5652 2327 5699 2328
rect 5665 2322 5699 2327
rect 5433 2301 5607 2304
rect 5426 2298 5607 2301
rect 5635 2321 5699 2322
rect 5229 2278 5248 2280
rect 5263 2278 5297 2280
rect 5229 2262 5309 2278
rect 5229 2256 5248 2262
rect 4945 2230 5048 2240
rect 4899 2228 5048 2230
rect 5069 2228 5104 2240
rect 4738 2226 4900 2228
rect 4750 2206 4769 2226
rect 4784 2224 4814 2226
rect 4633 2198 4674 2206
rect 4756 2202 4769 2206
rect 4821 2210 4900 2226
rect 4932 2226 5104 2228
rect 4932 2210 5011 2226
rect 5018 2224 5048 2226
rect 4596 2188 4625 2198
rect 4639 2188 4668 2198
rect 4683 2188 4713 2202
rect 4756 2188 4799 2202
rect 4821 2198 5011 2210
rect 5076 2206 5082 2226
rect 4806 2188 4836 2198
rect 4837 2188 4995 2198
rect 4999 2188 5029 2198
rect 5033 2188 5063 2202
rect 5091 2188 5104 2226
rect 5176 2240 5205 2256
rect 5219 2240 5248 2256
rect 5263 2246 5293 2262
rect 5321 2240 5327 2288
rect 5330 2282 5349 2288
rect 5364 2282 5394 2290
rect 5330 2274 5394 2282
rect 5330 2258 5410 2274
rect 5426 2267 5488 2298
rect 5504 2267 5566 2298
rect 5635 2296 5684 2321
rect 5699 2296 5729 2312
rect 5598 2282 5628 2290
rect 5635 2288 5745 2296
rect 5598 2274 5643 2282
rect 5330 2256 5349 2258
rect 5364 2256 5410 2258
rect 5330 2240 5410 2256
rect 5437 2254 5472 2267
rect 5513 2264 5550 2267
rect 5513 2262 5555 2264
rect 5442 2251 5472 2254
rect 5451 2247 5458 2251
rect 5458 2246 5459 2247
rect 5417 2240 5427 2246
rect 5176 2232 5211 2240
rect 5176 2206 5177 2232
rect 5184 2206 5211 2232
rect 5119 2188 5149 2202
rect 5176 2198 5211 2206
rect 5213 2232 5254 2240
rect 5213 2206 5228 2232
rect 5235 2206 5254 2232
rect 5318 2228 5349 2240
rect 5364 2228 5467 2240
rect 5479 2230 5505 2256
rect 5520 2251 5550 2262
rect 5582 2258 5644 2274
rect 5582 2256 5628 2258
rect 5582 2240 5644 2256
rect 5656 2240 5662 2288
rect 5665 2280 5745 2288
rect 5665 2278 5684 2280
rect 5699 2278 5733 2280
rect 5665 2262 5745 2278
rect 5665 2240 5684 2262
rect 5699 2246 5729 2262
rect 5757 2256 5763 2330
rect 5766 2256 5785 2400
rect 5800 2256 5806 2400
rect 5815 2330 5828 2400
rect 5880 2396 5902 2400
rect 5873 2374 5902 2388
rect 5955 2374 5971 2388
rect 6009 2384 6015 2386
rect 6022 2384 6130 2400
rect 6137 2384 6143 2386
rect 6151 2384 6166 2400
rect 6232 2394 6251 2397
rect 5873 2372 5971 2374
rect 5998 2372 6166 2384
rect 6181 2374 6197 2388
rect 6232 2375 6254 2394
rect 6264 2388 6280 2389
rect 6263 2386 6280 2388
rect 6264 2381 6280 2386
rect 6254 2374 6260 2375
rect 6263 2374 6292 2381
rect 6181 2373 6292 2374
rect 6181 2372 6298 2373
rect 5857 2364 5908 2372
rect 5955 2364 5989 2372
rect 5857 2352 5882 2364
rect 5889 2352 5908 2364
rect 5962 2362 5989 2364
rect 5998 2362 6219 2372
rect 6254 2369 6260 2372
rect 5962 2358 6219 2362
rect 5857 2344 5908 2352
rect 5955 2344 6219 2358
rect 6263 2364 6298 2372
rect 5809 2296 5828 2330
rect 5873 2336 5902 2344
rect 5873 2330 5890 2336
rect 5873 2328 5907 2330
rect 5955 2328 5971 2344
rect 5972 2334 6180 2344
rect 6181 2334 6197 2344
rect 6245 2340 6260 2355
rect 6263 2352 6264 2364
rect 6271 2352 6298 2364
rect 6263 2344 6298 2352
rect 6263 2343 6292 2344
rect 5983 2330 6197 2334
rect 5998 2328 6197 2330
rect 6232 2330 6245 2340
rect 6263 2330 6280 2343
rect 6232 2328 6280 2330
rect 5874 2324 5907 2328
rect 5870 2322 5907 2324
rect 5870 2321 5937 2322
rect 5870 2316 5901 2321
rect 5907 2316 5937 2321
rect 5870 2312 5937 2316
rect 5843 2309 5937 2312
rect 5843 2302 5892 2309
rect 5843 2296 5873 2302
rect 5892 2297 5897 2302
rect 5809 2280 5889 2296
rect 5901 2288 5937 2309
rect 5998 2304 6187 2328
rect 6232 2327 6279 2328
rect 6245 2322 6279 2327
rect 6013 2301 6187 2304
rect 6006 2298 6187 2301
rect 6215 2321 6279 2322
rect 5809 2278 5828 2280
rect 5843 2278 5877 2280
rect 5809 2262 5889 2278
rect 5809 2256 5828 2262
rect 5525 2230 5628 2240
rect 5479 2228 5628 2230
rect 5649 2228 5684 2240
rect 5318 2226 5480 2228
rect 5330 2206 5349 2226
rect 5364 2224 5394 2226
rect 5213 2198 5254 2206
rect 5336 2202 5349 2206
rect 5401 2210 5480 2226
rect 5512 2226 5684 2228
rect 5512 2210 5591 2226
rect 5598 2224 5628 2226
rect 5176 2188 5205 2198
rect 5219 2188 5248 2198
rect 5263 2188 5293 2202
rect 5336 2188 5379 2202
rect 5401 2198 5591 2210
rect 5656 2206 5662 2226
rect 5386 2188 5416 2198
rect 5417 2188 5575 2198
rect 5579 2188 5609 2198
rect 5613 2188 5643 2202
rect 5671 2188 5684 2226
rect 5756 2240 5785 2256
rect 5799 2240 5828 2256
rect 5843 2246 5873 2262
rect 5901 2240 5907 2288
rect 5910 2282 5929 2288
rect 5944 2282 5974 2290
rect 5910 2274 5974 2282
rect 5910 2258 5990 2274
rect 6006 2267 6068 2298
rect 6084 2267 6146 2298
rect 6215 2296 6264 2321
rect 6279 2296 6309 2312
rect 6178 2282 6208 2290
rect 6215 2288 6325 2296
rect 6178 2274 6223 2282
rect 5910 2256 5929 2258
rect 5944 2256 5990 2258
rect 5910 2240 5990 2256
rect 6017 2254 6052 2267
rect 6093 2264 6130 2267
rect 6093 2262 6135 2264
rect 6022 2251 6052 2254
rect 6031 2247 6038 2251
rect 6038 2246 6039 2247
rect 5997 2240 6007 2246
rect 5756 2232 5791 2240
rect 5756 2206 5757 2232
rect 5764 2206 5791 2232
rect 5699 2188 5729 2202
rect 5756 2198 5791 2206
rect 5793 2232 5834 2240
rect 5793 2206 5808 2232
rect 5815 2206 5834 2232
rect 5898 2228 5929 2240
rect 5944 2228 6047 2240
rect 6059 2230 6085 2256
rect 6100 2251 6130 2262
rect 6162 2258 6224 2274
rect 6162 2256 6208 2258
rect 6162 2240 6224 2256
rect 6236 2240 6242 2288
rect 6245 2280 6325 2288
rect 6245 2278 6264 2280
rect 6279 2278 6313 2280
rect 6245 2262 6325 2278
rect 6245 2240 6264 2262
rect 6279 2246 6309 2262
rect 6337 2256 6343 2330
rect 6346 2256 6365 2400
rect 6380 2256 6386 2400
rect 6395 2330 6408 2400
rect 6460 2396 6482 2400
rect 6453 2374 6482 2388
rect 6535 2374 6551 2388
rect 6589 2384 6595 2386
rect 6602 2384 6710 2400
rect 6717 2384 6723 2386
rect 6731 2384 6746 2400
rect 6812 2394 6831 2397
rect 6453 2372 6551 2374
rect 6578 2372 6746 2384
rect 6761 2374 6777 2388
rect 6812 2375 6834 2394
rect 6844 2388 6860 2389
rect 6843 2386 6860 2388
rect 6844 2381 6860 2386
rect 6834 2374 6840 2375
rect 6843 2374 6872 2381
rect 6761 2373 6872 2374
rect 6761 2372 6878 2373
rect 6437 2364 6488 2372
rect 6535 2364 6569 2372
rect 6437 2352 6462 2364
rect 6469 2352 6488 2364
rect 6542 2362 6569 2364
rect 6578 2362 6799 2372
rect 6834 2369 6840 2372
rect 6542 2358 6799 2362
rect 6437 2344 6488 2352
rect 6535 2344 6799 2358
rect 6843 2364 6878 2372
rect 6389 2296 6408 2330
rect 6453 2336 6482 2344
rect 6453 2330 6470 2336
rect 6453 2328 6487 2330
rect 6535 2328 6551 2344
rect 6552 2334 6760 2344
rect 6761 2334 6777 2344
rect 6825 2340 6840 2355
rect 6843 2352 6844 2364
rect 6851 2352 6878 2364
rect 6843 2344 6878 2352
rect 6843 2343 6872 2344
rect 6563 2330 6777 2334
rect 6578 2328 6777 2330
rect 6812 2330 6825 2340
rect 6843 2330 6860 2343
rect 6812 2328 6860 2330
rect 6454 2324 6487 2328
rect 6450 2322 6487 2324
rect 6450 2321 6517 2322
rect 6450 2316 6481 2321
rect 6487 2316 6517 2321
rect 6450 2312 6517 2316
rect 6423 2309 6517 2312
rect 6423 2302 6472 2309
rect 6423 2296 6453 2302
rect 6472 2297 6477 2302
rect 6389 2280 6469 2296
rect 6481 2288 6517 2309
rect 6578 2304 6767 2328
rect 6812 2327 6859 2328
rect 6825 2322 6859 2327
rect 6593 2301 6767 2304
rect 6586 2298 6767 2301
rect 6795 2321 6859 2322
rect 6389 2278 6408 2280
rect 6423 2278 6457 2280
rect 6389 2262 6469 2278
rect 6389 2256 6408 2262
rect 6105 2230 6208 2240
rect 6059 2228 6208 2230
rect 6229 2228 6264 2240
rect 5898 2226 6060 2228
rect 5910 2206 5929 2226
rect 5944 2224 5974 2226
rect 5793 2198 5834 2206
rect 5916 2202 5929 2206
rect 5981 2210 6060 2226
rect 6092 2226 6264 2228
rect 6092 2210 6171 2226
rect 6178 2224 6208 2226
rect 5756 2188 5785 2198
rect 5799 2188 5828 2198
rect 5843 2188 5873 2202
rect 5916 2188 5959 2202
rect 5981 2198 6171 2210
rect 6236 2206 6242 2226
rect 5966 2188 5996 2198
rect 5997 2188 6155 2198
rect 6159 2188 6189 2198
rect 6193 2188 6223 2202
rect 6251 2188 6264 2226
rect 6336 2240 6365 2256
rect 6379 2240 6408 2256
rect 6423 2246 6453 2262
rect 6481 2240 6487 2288
rect 6490 2282 6509 2288
rect 6524 2282 6554 2290
rect 6490 2274 6554 2282
rect 6490 2258 6570 2274
rect 6586 2267 6648 2298
rect 6664 2267 6726 2298
rect 6795 2296 6844 2321
rect 6859 2296 6889 2312
rect 6758 2282 6788 2290
rect 6795 2288 6905 2296
rect 6758 2274 6803 2282
rect 6490 2256 6509 2258
rect 6524 2256 6570 2258
rect 6490 2240 6570 2256
rect 6597 2254 6632 2267
rect 6673 2264 6710 2267
rect 6673 2262 6715 2264
rect 6602 2251 6632 2254
rect 6611 2247 6618 2251
rect 6618 2246 6619 2247
rect 6577 2240 6587 2246
rect 6336 2232 6371 2240
rect 6336 2206 6337 2232
rect 6344 2206 6371 2232
rect 6279 2188 6309 2202
rect 6336 2198 6371 2206
rect 6373 2232 6414 2240
rect 6373 2206 6388 2232
rect 6395 2206 6414 2232
rect 6478 2228 6509 2240
rect 6524 2228 6627 2240
rect 6639 2230 6665 2256
rect 6680 2251 6710 2262
rect 6742 2258 6804 2274
rect 6742 2256 6788 2258
rect 6742 2240 6804 2256
rect 6816 2240 6822 2288
rect 6825 2280 6905 2288
rect 6825 2278 6844 2280
rect 6859 2278 6893 2280
rect 6825 2262 6905 2278
rect 6825 2240 6844 2262
rect 6859 2246 6889 2262
rect 6917 2256 6923 2330
rect 6926 2256 6945 2400
rect 6960 2256 6966 2400
rect 6975 2330 6988 2400
rect 7040 2396 7062 2400
rect 7033 2374 7062 2388
rect 7115 2374 7131 2388
rect 7169 2384 7175 2386
rect 7182 2384 7290 2400
rect 7297 2384 7303 2386
rect 7311 2384 7326 2400
rect 7392 2394 7411 2397
rect 7033 2372 7131 2374
rect 7158 2372 7326 2384
rect 7341 2374 7357 2388
rect 7392 2375 7414 2394
rect 7424 2388 7440 2389
rect 7423 2386 7440 2388
rect 7424 2381 7440 2386
rect 7414 2374 7420 2375
rect 7423 2374 7452 2381
rect 7341 2373 7452 2374
rect 7341 2372 7458 2373
rect 7017 2364 7068 2372
rect 7115 2364 7149 2372
rect 7017 2352 7042 2364
rect 7049 2352 7068 2364
rect 7122 2362 7149 2364
rect 7158 2362 7379 2372
rect 7414 2369 7420 2372
rect 7122 2358 7379 2362
rect 7017 2344 7068 2352
rect 7115 2344 7379 2358
rect 7423 2364 7458 2372
rect 6969 2296 6988 2330
rect 7033 2336 7062 2344
rect 7033 2330 7050 2336
rect 7033 2328 7067 2330
rect 7115 2328 7131 2344
rect 7132 2334 7340 2344
rect 7341 2334 7357 2344
rect 7405 2340 7420 2355
rect 7423 2352 7424 2364
rect 7431 2352 7458 2364
rect 7423 2344 7458 2352
rect 7423 2343 7452 2344
rect 7143 2330 7357 2334
rect 7158 2328 7357 2330
rect 7392 2330 7405 2340
rect 7423 2330 7440 2343
rect 7392 2328 7440 2330
rect 7034 2324 7067 2328
rect 7030 2322 7067 2324
rect 7030 2321 7097 2322
rect 7030 2316 7061 2321
rect 7067 2316 7097 2321
rect 7030 2312 7097 2316
rect 7003 2309 7097 2312
rect 7003 2302 7052 2309
rect 7003 2296 7033 2302
rect 7052 2297 7057 2302
rect 6969 2280 7049 2296
rect 7061 2288 7097 2309
rect 7158 2304 7347 2328
rect 7392 2327 7439 2328
rect 7405 2322 7439 2327
rect 7173 2301 7347 2304
rect 7166 2298 7347 2301
rect 7375 2321 7439 2322
rect 6969 2278 6988 2280
rect 7003 2278 7037 2280
rect 6969 2262 7049 2278
rect 6969 2256 6988 2262
rect 6685 2230 6788 2240
rect 6639 2228 6788 2230
rect 6809 2228 6844 2240
rect 6478 2226 6640 2228
rect 6490 2206 6509 2226
rect 6524 2224 6554 2226
rect 6373 2198 6414 2206
rect 6496 2202 6509 2206
rect 6561 2210 6640 2226
rect 6672 2226 6844 2228
rect 6672 2210 6751 2226
rect 6758 2224 6788 2226
rect 6336 2188 6365 2198
rect 6379 2188 6408 2198
rect 6423 2188 6453 2202
rect 6496 2188 6539 2202
rect 6561 2198 6751 2210
rect 6816 2206 6822 2226
rect 6546 2188 6576 2198
rect 6577 2188 6735 2198
rect 6739 2188 6769 2198
rect 6773 2188 6803 2202
rect 6831 2188 6844 2226
rect 6916 2240 6945 2256
rect 6959 2240 6988 2256
rect 7003 2246 7033 2262
rect 7061 2240 7067 2288
rect 7070 2282 7089 2288
rect 7104 2282 7134 2290
rect 7070 2274 7134 2282
rect 7070 2258 7150 2274
rect 7166 2267 7228 2298
rect 7244 2267 7306 2298
rect 7375 2296 7424 2321
rect 7439 2296 7469 2312
rect 7338 2282 7368 2290
rect 7375 2288 7485 2296
rect 7338 2274 7383 2282
rect 7070 2256 7089 2258
rect 7104 2256 7150 2258
rect 7070 2240 7150 2256
rect 7177 2254 7212 2267
rect 7253 2264 7290 2267
rect 7253 2262 7295 2264
rect 7182 2251 7212 2254
rect 7191 2247 7198 2251
rect 7198 2246 7199 2247
rect 7157 2240 7167 2246
rect 6916 2232 6951 2240
rect 6916 2206 6917 2232
rect 6924 2206 6951 2232
rect 6859 2188 6889 2202
rect 6916 2198 6951 2206
rect 6953 2232 6994 2240
rect 6953 2206 6968 2232
rect 6975 2206 6994 2232
rect 7058 2228 7089 2240
rect 7104 2228 7207 2240
rect 7219 2230 7245 2256
rect 7260 2251 7290 2262
rect 7322 2258 7384 2274
rect 7322 2256 7368 2258
rect 7322 2240 7384 2256
rect 7396 2240 7402 2288
rect 7405 2280 7485 2288
rect 7405 2278 7424 2280
rect 7439 2278 7473 2280
rect 7405 2262 7485 2278
rect 7405 2240 7424 2262
rect 7439 2246 7469 2262
rect 7497 2256 7503 2330
rect 7506 2256 7525 2400
rect 7540 2256 7546 2400
rect 7555 2330 7568 2400
rect 7620 2396 7642 2400
rect 7613 2374 7642 2388
rect 7695 2374 7711 2388
rect 7749 2384 7755 2386
rect 7762 2384 7870 2400
rect 7877 2384 7883 2386
rect 7891 2384 7906 2400
rect 7972 2394 7991 2397
rect 7613 2372 7711 2374
rect 7738 2372 7906 2384
rect 7921 2374 7937 2388
rect 7972 2375 7994 2394
rect 8004 2388 8020 2389
rect 8003 2386 8020 2388
rect 8004 2381 8020 2386
rect 7994 2374 8000 2375
rect 8003 2374 8032 2381
rect 7921 2373 8032 2374
rect 7921 2372 8038 2373
rect 7597 2364 7648 2372
rect 7695 2364 7729 2372
rect 7597 2352 7622 2364
rect 7629 2352 7648 2364
rect 7702 2362 7729 2364
rect 7738 2362 7959 2372
rect 7994 2369 8000 2372
rect 7702 2358 7959 2362
rect 7597 2344 7648 2352
rect 7695 2344 7959 2358
rect 8003 2364 8038 2372
rect 7549 2296 7568 2330
rect 7613 2336 7642 2344
rect 7613 2330 7630 2336
rect 7613 2328 7647 2330
rect 7695 2328 7711 2344
rect 7712 2334 7920 2344
rect 7921 2334 7937 2344
rect 7985 2340 8000 2355
rect 8003 2352 8004 2364
rect 8011 2352 8038 2364
rect 8003 2344 8038 2352
rect 8003 2343 8032 2344
rect 7723 2330 7937 2334
rect 7738 2328 7937 2330
rect 7972 2330 7985 2340
rect 8003 2330 8020 2343
rect 7972 2328 8020 2330
rect 7614 2324 7647 2328
rect 7610 2322 7647 2324
rect 7610 2321 7677 2322
rect 7610 2316 7641 2321
rect 7647 2316 7677 2321
rect 7610 2312 7677 2316
rect 7583 2309 7677 2312
rect 7583 2302 7632 2309
rect 7583 2296 7613 2302
rect 7632 2297 7637 2302
rect 7549 2280 7629 2296
rect 7641 2288 7677 2309
rect 7738 2304 7927 2328
rect 7972 2327 8019 2328
rect 7985 2322 8019 2327
rect 7753 2301 7927 2304
rect 7746 2298 7927 2301
rect 7955 2321 8019 2322
rect 7549 2278 7568 2280
rect 7583 2278 7617 2280
rect 7549 2262 7629 2278
rect 7549 2256 7568 2262
rect 7265 2230 7368 2240
rect 7219 2228 7368 2230
rect 7389 2228 7424 2240
rect 7058 2226 7220 2228
rect 7070 2206 7089 2226
rect 7104 2224 7134 2226
rect 6953 2198 6994 2206
rect 7076 2202 7089 2206
rect 7141 2210 7220 2226
rect 7252 2226 7424 2228
rect 7252 2210 7331 2226
rect 7338 2224 7368 2226
rect 6916 2188 6945 2198
rect 6959 2188 6988 2198
rect 7003 2188 7033 2202
rect 7076 2188 7119 2202
rect 7141 2198 7331 2210
rect 7396 2206 7402 2226
rect 7126 2188 7156 2198
rect 7157 2188 7315 2198
rect 7319 2188 7349 2198
rect 7353 2188 7383 2202
rect 7411 2188 7424 2226
rect 7496 2240 7525 2256
rect 7539 2240 7568 2256
rect 7583 2246 7613 2262
rect 7641 2240 7647 2288
rect 7650 2282 7669 2288
rect 7684 2282 7714 2290
rect 7650 2274 7714 2282
rect 7650 2258 7730 2274
rect 7746 2267 7808 2298
rect 7824 2267 7886 2298
rect 7955 2296 8004 2321
rect 8019 2296 8049 2312
rect 7918 2282 7948 2290
rect 7955 2288 8065 2296
rect 7918 2274 7963 2282
rect 7650 2256 7669 2258
rect 7684 2256 7730 2258
rect 7650 2240 7730 2256
rect 7757 2254 7792 2267
rect 7833 2264 7870 2267
rect 7833 2262 7875 2264
rect 7762 2251 7792 2254
rect 7771 2247 7778 2251
rect 7778 2246 7779 2247
rect 7737 2240 7747 2246
rect 7496 2232 7531 2240
rect 7496 2206 7497 2232
rect 7504 2206 7531 2232
rect 7439 2188 7469 2202
rect 7496 2198 7531 2206
rect 7533 2232 7574 2240
rect 7533 2206 7548 2232
rect 7555 2206 7574 2232
rect 7638 2228 7669 2240
rect 7684 2228 7787 2240
rect 7799 2230 7825 2256
rect 7840 2251 7870 2262
rect 7902 2258 7964 2274
rect 7902 2256 7948 2258
rect 7902 2240 7964 2256
rect 7976 2240 7982 2288
rect 7985 2280 8065 2288
rect 7985 2278 8004 2280
rect 8019 2278 8053 2280
rect 7985 2262 8065 2278
rect 7985 2240 8004 2262
rect 8019 2246 8049 2262
rect 8077 2256 8083 2330
rect 8086 2256 8105 2400
rect 8120 2256 8126 2400
rect 8135 2330 8148 2400
rect 8200 2396 8222 2400
rect 8193 2374 8222 2388
rect 8275 2374 8291 2388
rect 8329 2384 8335 2386
rect 8342 2384 8450 2400
rect 8457 2384 8463 2386
rect 8471 2384 8486 2400
rect 8552 2394 8571 2397
rect 8193 2372 8291 2374
rect 8318 2372 8486 2384
rect 8501 2374 8517 2388
rect 8552 2375 8574 2394
rect 8584 2388 8600 2389
rect 8583 2386 8600 2388
rect 8584 2381 8600 2386
rect 8574 2374 8580 2375
rect 8583 2374 8612 2381
rect 8501 2373 8612 2374
rect 8501 2372 8618 2373
rect 8177 2364 8228 2372
rect 8275 2364 8309 2372
rect 8177 2352 8202 2364
rect 8209 2352 8228 2364
rect 8282 2362 8309 2364
rect 8318 2362 8539 2372
rect 8574 2369 8580 2372
rect 8282 2358 8539 2362
rect 8177 2344 8228 2352
rect 8275 2344 8539 2358
rect 8583 2364 8618 2372
rect 8129 2296 8148 2330
rect 8193 2336 8222 2344
rect 8193 2330 8210 2336
rect 8193 2328 8227 2330
rect 8275 2328 8291 2344
rect 8292 2334 8500 2344
rect 8501 2334 8517 2344
rect 8565 2340 8580 2355
rect 8583 2352 8584 2364
rect 8591 2352 8618 2364
rect 8583 2344 8618 2352
rect 8583 2343 8612 2344
rect 8303 2330 8517 2334
rect 8318 2328 8517 2330
rect 8552 2330 8565 2340
rect 8583 2330 8600 2343
rect 8552 2328 8600 2330
rect 8194 2324 8227 2328
rect 8190 2322 8227 2324
rect 8190 2321 8257 2322
rect 8190 2316 8221 2321
rect 8227 2316 8257 2321
rect 8190 2312 8257 2316
rect 8163 2309 8257 2312
rect 8163 2302 8212 2309
rect 8163 2296 8193 2302
rect 8212 2297 8217 2302
rect 8129 2280 8209 2296
rect 8221 2288 8257 2309
rect 8318 2304 8507 2328
rect 8552 2327 8599 2328
rect 8565 2322 8599 2327
rect 8333 2301 8507 2304
rect 8326 2298 8507 2301
rect 8535 2321 8599 2322
rect 8129 2278 8148 2280
rect 8163 2278 8197 2280
rect 8129 2262 8209 2278
rect 8129 2256 8148 2262
rect 7845 2230 7948 2240
rect 7799 2228 7948 2230
rect 7969 2228 8004 2240
rect 7638 2226 7800 2228
rect 7650 2206 7669 2226
rect 7684 2224 7714 2226
rect 7533 2198 7574 2206
rect 7656 2202 7669 2206
rect 7721 2210 7800 2226
rect 7832 2226 8004 2228
rect 7832 2210 7911 2226
rect 7918 2224 7948 2226
rect 7496 2188 7525 2198
rect 7539 2188 7568 2198
rect 7583 2188 7613 2202
rect 7656 2188 7699 2202
rect 7721 2198 7911 2210
rect 7976 2206 7982 2226
rect 7706 2188 7736 2198
rect 7737 2188 7895 2198
rect 7899 2188 7929 2198
rect 7933 2188 7963 2202
rect 7991 2188 8004 2226
rect 8076 2240 8105 2256
rect 8119 2240 8148 2256
rect 8163 2246 8193 2262
rect 8221 2240 8227 2288
rect 8230 2282 8249 2288
rect 8264 2282 8294 2290
rect 8230 2274 8294 2282
rect 8230 2258 8310 2274
rect 8326 2267 8388 2298
rect 8404 2267 8466 2298
rect 8535 2296 8584 2321
rect 8599 2296 8629 2312
rect 8498 2282 8528 2290
rect 8535 2288 8645 2296
rect 8498 2274 8543 2282
rect 8230 2256 8249 2258
rect 8264 2256 8310 2258
rect 8230 2240 8310 2256
rect 8337 2254 8372 2267
rect 8413 2264 8450 2267
rect 8413 2262 8455 2264
rect 8342 2251 8372 2254
rect 8351 2247 8358 2251
rect 8358 2246 8359 2247
rect 8317 2240 8327 2246
rect 8076 2232 8111 2240
rect 8076 2206 8077 2232
rect 8084 2206 8111 2232
rect 8019 2188 8049 2202
rect 8076 2198 8111 2206
rect 8113 2232 8154 2240
rect 8113 2206 8128 2232
rect 8135 2206 8154 2232
rect 8218 2228 8249 2240
rect 8264 2228 8367 2240
rect 8379 2230 8405 2256
rect 8420 2251 8450 2262
rect 8482 2258 8544 2274
rect 8482 2256 8528 2258
rect 8482 2240 8544 2256
rect 8556 2240 8562 2288
rect 8565 2280 8645 2288
rect 8565 2278 8584 2280
rect 8599 2278 8633 2280
rect 8565 2262 8645 2278
rect 8565 2240 8584 2262
rect 8599 2246 8629 2262
rect 8657 2256 8663 2330
rect 8666 2256 8685 2400
rect 8700 2256 8706 2400
rect 8715 2330 8728 2400
rect 8780 2396 8802 2400
rect 8773 2374 8802 2388
rect 8855 2374 8871 2388
rect 8909 2384 8915 2386
rect 8922 2384 9030 2400
rect 9037 2384 9043 2386
rect 9051 2384 9066 2400
rect 9132 2394 9151 2397
rect 8773 2372 8871 2374
rect 8898 2372 9066 2384
rect 9081 2374 9097 2388
rect 9132 2375 9154 2394
rect 9164 2388 9180 2389
rect 9163 2386 9180 2388
rect 9164 2381 9180 2386
rect 9154 2374 9160 2375
rect 9163 2374 9192 2381
rect 9081 2373 9192 2374
rect 9081 2372 9198 2373
rect 8757 2364 8808 2372
rect 8855 2364 8889 2372
rect 8757 2352 8782 2364
rect 8789 2352 8808 2364
rect 8862 2362 8889 2364
rect 8898 2362 9119 2372
rect 9154 2369 9160 2372
rect 8862 2358 9119 2362
rect 8757 2344 8808 2352
rect 8855 2344 9119 2358
rect 9163 2364 9198 2372
rect 8709 2296 8728 2330
rect 8773 2336 8802 2344
rect 8773 2330 8790 2336
rect 8773 2328 8807 2330
rect 8855 2328 8871 2344
rect 8872 2334 9080 2344
rect 9081 2334 9097 2344
rect 9145 2340 9160 2355
rect 9163 2352 9164 2364
rect 9171 2352 9198 2364
rect 9163 2344 9198 2352
rect 9163 2343 9192 2344
rect 8883 2330 9097 2334
rect 8898 2328 9097 2330
rect 9132 2330 9145 2340
rect 9163 2330 9180 2343
rect 9132 2328 9180 2330
rect 8774 2324 8807 2328
rect 8770 2322 8807 2324
rect 8770 2321 8837 2322
rect 8770 2316 8801 2321
rect 8807 2316 8837 2321
rect 8770 2312 8837 2316
rect 8743 2309 8837 2312
rect 8743 2302 8792 2309
rect 8743 2296 8773 2302
rect 8792 2297 8797 2302
rect 8709 2280 8789 2296
rect 8801 2288 8837 2309
rect 8898 2304 9087 2328
rect 9132 2327 9179 2328
rect 9145 2322 9179 2327
rect 8913 2301 9087 2304
rect 8906 2298 9087 2301
rect 9115 2321 9179 2322
rect 8709 2278 8728 2280
rect 8743 2278 8777 2280
rect 8709 2262 8789 2278
rect 8709 2256 8728 2262
rect 8425 2230 8528 2240
rect 8379 2228 8528 2230
rect 8549 2228 8584 2240
rect 8218 2226 8380 2228
rect 8230 2206 8249 2226
rect 8264 2224 8294 2226
rect 8113 2198 8154 2206
rect 8236 2202 8249 2206
rect 8301 2210 8380 2226
rect 8412 2226 8584 2228
rect 8412 2210 8491 2226
rect 8498 2224 8528 2226
rect 8076 2188 8105 2198
rect 8119 2188 8148 2198
rect 8163 2188 8193 2202
rect 8236 2188 8279 2202
rect 8301 2198 8491 2210
rect 8556 2206 8562 2226
rect 8286 2188 8316 2198
rect 8317 2188 8475 2198
rect 8479 2188 8509 2198
rect 8513 2188 8543 2202
rect 8571 2188 8584 2226
rect 8656 2240 8685 2256
rect 8699 2240 8728 2256
rect 8743 2246 8773 2262
rect 8801 2240 8807 2288
rect 8810 2282 8829 2288
rect 8844 2282 8874 2290
rect 8810 2274 8874 2282
rect 8810 2258 8890 2274
rect 8906 2267 8968 2298
rect 8984 2267 9046 2298
rect 9115 2296 9164 2321
rect 9179 2296 9209 2312
rect 9078 2282 9108 2290
rect 9115 2288 9225 2296
rect 9078 2274 9123 2282
rect 8810 2256 8829 2258
rect 8844 2256 8890 2258
rect 8810 2240 8890 2256
rect 8917 2254 8952 2267
rect 8993 2264 9030 2267
rect 8993 2262 9035 2264
rect 8922 2251 8952 2254
rect 8931 2247 8938 2251
rect 8938 2246 8939 2247
rect 8897 2240 8907 2246
rect 8656 2232 8691 2240
rect 8656 2206 8657 2232
rect 8664 2206 8691 2232
rect 8599 2188 8629 2202
rect 8656 2198 8691 2206
rect 8693 2232 8734 2240
rect 8693 2206 8708 2232
rect 8715 2206 8734 2232
rect 8798 2228 8829 2240
rect 8844 2228 8947 2240
rect 8959 2230 8985 2256
rect 9000 2251 9030 2262
rect 9062 2258 9124 2274
rect 9062 2256 9108 2258
rect 9062 2240 9124 2256
rect 9136 2240 9142 2288
rect 9145 2280 9225 2288
rect 9145 2278 9164 2280
rect 9179 2278 9213 2280
rect 9145 2262 9225 2278
rect 9145 2240 9164 2262
rect 9179 2246 9209 2262
rect 9237 2256 9243 2330
rect 9252 2256 9265 2400
rect 9005 2230 9108 2240
rect 8959 2228 9108 2230
rect 9129 2228 9164 2240
rect 8798 2226 8960 2228
rect 8810 2206 8829 2226
rect 8844 2224 8874 2226
rect 8693 2198 8734 2206
rect 8816 2202 8829 2206
rect 8881 2210 8960 2226
rect 8992 2226 9164 2228
rect 8992 2210 9071 2226
rect 9078 2224 9108 2226
rect 8656 2188 8685 2198
rect 8699 2188 8728 2198
rect 8743 2188 8773 2202
rect 8816 2188 8859 2202
rect 8881 2198 9071 2210
rect 9136 2206 9142 2226
rect 8866 2188 8896 2198
rect 8897 2188 9055 2198
rect 9059 2188 9089 2198
rect 9093 2188 9123 2202
rect 9151 2188 9164 2226
rect 9236 2240 9265 2256
rect 9236 2232 9271 2240
rect 9236 2206 9237 2232
rect 9244 2206 9271 2232
rect 9179 2188 9209 2202
rect 9236 2198 9271 2206
rect 9236 2188 9265 2198
rect -1 2182 9265 2188
rect 0 2174 9265 2182
rect 15 2144 28 2174
rect 43 2160 73 2174
rect 116 2160 159 2174
rect 166 2160 386 2174
rect 393 2160 423 2174
rect 83 2146 98 2158
rect 117 2146 130 2160
rect 198 2156 351 2160
rect 80 2144 102 2146
rect 180 2144 372 2156
rect 451 2144 464 2174
rect 479 2160 509 2174
rect 546 2144 565 2174
rect 580 2144 586 2174
rect 595 2144 608 2174
rect 623 2160 653 2174
rect 696 2160 739 2174
rect 746 2160 966 2174
rect 973 2160 1003 2174
rect 663 2146 678 2158
rect 697 2146 710 2160
rect 778 2156 931 2160
rect 660 2144 682 2146
rect 760 2144 952 2156
rect 1031 2144 1044 2174
rect 1059 2160 1089 2174
rect 1126 2144 1145 2174
rect 1160 2144 1166 2174
rect 1175 2144 1188 2174
rect 1203 2160 1233 2174
rect 1276 2160 1319 2174
rect 1326 2160 1546 2174
rect 1553 2160 1583 2174
rect 1243 2146 1258 2158
rect 1277 2146 1290 2160
rect 1358 2156 1511 2160
rect 1240 2144 1262 2146
rect 1340 2144 1532 2156
rect 1611 2144 1624 2174
rect 1639 2160 1669 2174
rect 1706 2144 1725 2174
rect 1740 2144 1746 2174
rect 1755 2144 1768 2174
rect 1783 2160 1813 2174
rect 1856 2160 1899 2174
rect 1906 2160 2126 2174
rect 2133 2160 2163 2174
rect 1823 2146 1838 2158
rect 1857 2146 1870 2160
rect 1938 2156 2091 2160
rect 1820 2144 1842 2146
rect 1920 2144 2112 2156
rect 2191 2144 2204 2174
rect 2219 2160 2249 2174
rect 2286 2144 2305 2174
rect 2320 2144 2326 2174
rect 2335 2144 2348 2174
rect 2363 2160 2393 2174
rect 2436 2160 2479 2174
rect 2486 2160 2706 2174
rect 2713 2160 2743 2174
rect 2403 2146 2418 2158
rect 2437 2146 2450 2160
rect 2518 2156 2671 2160
rect 2400 2144 2422 2146
rect 2500 2144 2692 2156
rect 2771 2144 2784 2174
rect 2799 2160 2829 2174
rect 2866 2144 2885 2174
rect 2900 2144 2906 2174
rect 2915 2144 2928 2174
rect 2943 2160 2973 2174
rect 3016 2160 3059 2174
rect 3066 2160 3286 2174
rect 3293 2160 3323 2174
rect 2983 2146 2998 2158
rect 3017 2146 3030 2160
rect 3098 2156 3251 2160
rect 2980 2144 3002 2146
rect 3080 2144 3272 2156
rect 3351 2144 3364 2174
rect 3379 2160 3409 2174
rect 3446 2144 3465 2174
rect 3480 2144 3486 2174
rect 3495 2144 3508 2174
rect 3523 2160 3553 2174
rect 3596 2160 3639 2174
rect 3646 2160 3866 2174
rect 3873 2160 3903 2174
rect 3563 2146 3578 2158
rect 3597 2146 3610 2160
rect 3678 2156 3831 2160
rect 3560 2144 3582 2146
rect 3660 2144 3852 2156
rect 3931 2144 3944 2174
rect 3959 2160 3989 2174
rect 4026 2144 4045 2174
rect 4060 2144 4066 2174
rect 4075 2144 4088 2174
rect 4103 2160 4133 2174
rect 4176 2160 4219 2174
rect 4226 2160 4446 2174
rect 4453 2160 4483 2174
rect 4143 2146 4158 2158
rect 4177 2146 4190 2160
rect 4258 2156 4411 2160
rect 4140 2144 4162 2146
rect 4240 2144 4432 2156
rect 4511 2144 4524 2174
rect 4539 2160 4569 2174
rect 4606 2144 4625 2174
rect 4640 2144 4646 2174
rect 4655 2144 4668 2174
rect 4683 2160 4713 2174
rect 4756 2160 4799 2174
rect 4806 2160 5026 2174
rect 5033 2160 5063 2174
rect 4723 2146 4738 2158
rect 4757 2146 4770 2160
rect 4838 2156 4991 2160
rect 4720 2144 4742 2146
rect 4820 2144 5012 2156
rect 5091 2144 5104 2174
rect 5119 2160 5149 2174
rect 5186 2144 5205 2174
rect 5220 2144 5226 2174
rect 5235 2144 5248 2174
rect 5263 2160 5293 2174
rect 5336 2160 5379 2174
rect 5386 2160 5606 2174
rect 5613 2160 5643 2174
rect 5303 2146 5318 2158
rect 5337 2146 5350 2160
rect 5418 2156 5571 2160
rect 5300 2144 5322 2146
rect 5400 2144 5592 2156
rect 5671 2144 5684 2174
rect 5699 2160 5729 2174
rect 5766 2144 5785 2174
rect 5800 2144 5806 2174
rect 5815 2144 5828 2174
rect 5843 2160 5873 2174
rect 5916 2160 5959 2174
rect 5966 2160 6186 2174
rect 6193 2160 6223 2174
rect 5883 2146 5898 2158
rect 5917 2146 5930 2160
rect 5998 2156 6151 2160
rect 5880 2144 5902 2146
rect 5980 2144 6172 2156
rect 6251 2144 6264 2174
rect 6279 2160 6309 2174
rect 6346 2144 6365 2174
rect 6380 2144 6386 2174
rect 6395 2144 6408 2174
rect 6423 2160 6453 2174
rect 6496 2160 6539 2174
rect 6546 2160 6766 2174
rect 6773 2160 6803 2174
rect 6463 2146 6478 2158
rect 6497 2146 6510 2160
rect 6578 2156 6731 2160
rect 6460 2144 6482 2146
rect 6560 2144 6752 2156
rect 6831 2144 6844 2174
rect 6859 2160 6889 2174
rect 6926 2144 6945 2174
rect 6960 2144 6966 2174
rect 6975 2144 6988 2174
rect 7003 2160 7033 2174
rect 7076 2160 7119 2174
rect 7126 2160 7346 2174
rect 7353 2160 7383 2174
rect 7043 2146 7058 2158
rect 7077 2146 7090 2160
rect 7158 2156 7311 2160
rect 7040 2144 7062 2146
rect 7140 2144 7332 2156
rect 7411 2144 7424 2174
rect 7439 2160 7469 2174
rect 7506 2144 7525 2174
rect 7540 2144 7546 2174
rect 7555 2144 7568 2174
rect 7583 2160 7613 2174
rect 7656 2160 7699 2174
rect 7706 2160 7926 2174
rect 7933 2160 7963 2174
rect 7623 2146 7638 2158
rect 7657 2146 7670 2160
rect 7738 2156 7891 2160
rect 7620 2144 7642 2146
rect 7720 2144 7912 2156
rect 7991 2144 8004 2174
rect 8019 2160 8049 2174
rect 8086 2144 8105 2174
rect 8120 2144 8126 2174
rect 8135 2144 8148 2174
rect 8163 2160 8193 2174
rect 8236 2160 8279 2174
rect 8286 2160 8506 2174
rect 8513 2160 8543 2174
rect 8203 2146 8218 2158
rect 8237 2146 8250 2160
rect 8318 2156 8471 2160
rect 8200 2144 8222 2146
rect 8300 2144 8492 2156
rect 8571 2144 8584 2174
rect 8599 2160 8629 2174
rect 8666 2144 8685 2174
rect 8700 2144 8706 2174
rect 8715 2144 8728 2174
rect 8743 2160 8773 2174
rect 8816 2160 8859 2174
rect 8866 2160 9086 2174
rect 9093 2160 9123 2174
rect 8783 2146 8798 2158
rect 8817 2146 8830 2160
rect 8898 2156 9051 2160
rect 8780 2144 8802 2146
rect 8880 2144 9072 2156
rect 9151 2144 9164 2174
rect 9179 2160 9209 2174
rect 9252 2144 9265 2174
rect 0 2130 9265 2144
rect 15 2060 28 2130
rect 80 2126 102 2130
rect 73 2104 102 2118
rect 155 2104 171 2118
rect 209 2114 215 2116
rect 222 2114 330 2130
rect 337 2114 343 2116
rect 351 2114 366 2130
rect 432 2124 451 2127
rect 73 2102 171 2104
rect 198 2102 366 2114
rect 381 2104 397 2118
rect 432 2105 454 2124
rect 464 2118 480 2119
rect 463 2116 480 2118
rect 464 2111 480 2116
rect 454 2104 460 2105
rect 463 2104 492 2111
rect 381 2103 492 2104
rect 381 2102 498 2103
rect 57 2094 108 2102
rect 155 2094 189 2102
rect 57 2082 82 2094
rect 89 2082 108 2094
rect 162 2092 189 2094
rect 198 2092 419 2102
rect 454 2099 460 2102
rect 162 2088 419 2092
rect 57 2074 108 2082
rect 155 2074 419 2088
rect 463 2094 498 2102
rect 9 2026 28 2060
rect 73 2066 102 2074
rect 73 2060 90 2066
rect 73 2058 107 2060
rect 155 2058 171 2074
rect 172 2064 380 2074
rect 381 2064 397 2074
rect 445 2070 460 2085
rect 463 2082 464 2094
rect 471 2082 498 2094
rect 463 2074 498 2082
rect 463 2073 492 2074
rect 183 2060 397 2064
rect 198 2058 397 2060
rect 432 2060 445 2070
rect 463 2060 480 2073
rect 432 2058 480 2060
rect 74 2054 107 2058
rect 70 2052 107 2054
rect 70 2051 137 2052
rect 70 2046 101 2051
rect 107 2046 137 2051
rect 70 2042 137 2046
rect 43 2039 137 2042
rect 43 2032 92 2039
rect 43 2026 73 2032
rect 92 2027 97 2032
rect 9 2010 89 2026
rect 101 2018 137 2039
rect 198 2034 387 2058
rect 432 2057 479 2058
rect 445 2052 479 2057
rect 213 2031 387 2034
rect 206 2028 387 2031
rect 415 2051 479 2052
rect 9 2008 28 2010
rect 43 2008 77 2010
rect 9 1992 89 2008
rect 9 1986 28 1992
rect -1 1970 28 1986
rect 43 1976 73 1992
rect 101 1970 107 2018
rect 110 2012 129 2018
rect 144 2012 174 2020
rect 110 2004 174 2012
rect 110 1988 190 2004
rect 206 1997 268 2028
rect 284 1997 346 2028
rect 415 2026 464 2051
rect 479 2026 509 2042
rect 378 2012 408 2020
rect 415 2018 525 2026
rect 378 2004 423 2012
rect 110 1986 129 1988
rect 144 1986 190 1988
rect 110 1970 190 1986
rect 217 1984 252 1997
rect 293 1994 330 1997
rect 293 1992 335 1994
rect 222 1981 252 1984
rect 231 1977 238 1981
rect 238 1976 239 1977
rect 197 1970 207 1976
rect -7 1962 34 1970
rect -7 1936 8 1962
rect 15 1936 34 1962
rect 98 1958 129 1970
rect 144 1958 247 1970
rect 259 1960 285 1986
rect 300 1981 330 1992
rect 362 1988 424 2004
rect 362 1986 408 1988
rect 362 1970 424 1986
rect 436 1970 442 2018
rect 445 2010 525 2018
rect 445 2008 464 2010
rect 479 2008 513 2010
rect 445 1992 525 2008
rect 445 1970 464 1992
rect 479 1976 509 1992
rect 537 1986 543 2060
rect 546 1986 565 2130
rect 580 1986 586 2130
rect 595 2060 608 2130
rect 660 2126 682 2130
rect 653 2104 682 2118
rect 735 2104 751 2118
rect 789 2114 795 2116
rect 802 2114 910 2130
rect 917 2114 923 2116
rect 931 2114 946 2130
rect 1012 2124 1031 2127
rect 653 2102 751 2104
rect 778 2102 946 2114
rect 961 2104 977 2118
rect 1012 2105 1034 2124
rect 1044 2118 1060 2119
rect 1043 2116 1060 2118
rect 1044 2111 1060 2116
rect 1034 2104 1040 2105
rect 1043 2104 1072 2111
rect 961 2103 1072 2104
rect 961 2102 1078 2103
rect 637 2094 688 2102
rect 735 2094 769 2102
rect 637 2082 662 2094
rect 669 2082 688 2094
rect 742 2092 769 2094
rect 778 2092 999 2102
rect 1034 2099 1040 2102
rect 742 2088 999 2092
rect 637 2074 688 2082
rect 735 2074 999 2088
rect 1043 2094 1078 2102
rect 589 2026 608 2060
rect 653 2066 682 2074
rect 653 2060 670 2066
rect 653 2058 687 2060
rect 735 2058 751 2074
rect 752 2064 960 2074
rect 961 2064 977 2074
rect 1025 2070 1040 2085
rect 1043 2082 1044 2094
rect 1051 2082 1078 2094
rect 1043 2074 1078 2082
rect 1043 2073 1072 2074
rect 763 2060 977 2064
rect 778 2058 977 2060
rect 1012 2060 1025 2070
rect 1043 2060 1060 2073
rect 1012 2058 1060 2060
rect 654 2054 687 2058
rect 650 2052 687 2054
rect 650 2051 717 2052
rect 650 2046 681 2051
rect 687 2046 717 2051
rect 650 2042 717 2046
rect 623 2039 717 2042
rect 623 2032 672 2039
rect 623 2026 653 2032
rect 672 2027 677 2032
rect 589 2010 669 2026
rect 681 2018 717 2039
rect 778 2034 967 2058
rect 1012 2057 1059 2058
rect 1025 2052 1059 2057
rect 793 2031 967 2034
rect 786 2028 967 2031
rect 995 2051 1059 2052
rect 589 2008 608 2010
rect 623 2008 657 2010
rect 589 1992 669 2008
rect 589 1986 608 1992
rect 305 1960 408 1970
rect 259 1958 408 1960
rect 429 1958 464 1970
rect 98 1956 260 1958
rect 110 1936 129 1956
rect 144 1954 174 1956
rect -7 1928 34 1936
rect 116 1932 129 1936
rect 181 1940 260 1956
rect 292 1956 464 1958
rect 292 1940 371 1956
rect 378 1954 408 1956
rect -1 1918 28 1928
rect 43 1918 73 1932
rect 116 1918 159 1932
rect 181 1928 371 1940
rect 436 1936 442 1956
rect 166 1918 196 1928
rect 197 1918 355 1928
rect 359 1918 389 1928
rect 393 1918 423 1932
rect 451 1918 464 1956
rect 536 1970 565 1986
rect 579 1970 608 1986
rect 623 1976 653 1992
rect 681 1970 687 2018
rect 690 2012 709 2018
rect 724 2012 754 2020
rect 690 2004 754 2012
rect 690 1988 770 2004
rect 786 1997 848 2028
rect 864 1997 926 2028
rect 995 2026 1044 2051
rect 1059 2026 1089 2042
rect 958 2012 988 2020
rect 995 2018 1105 2026
rect 958 2004 1003 2012
rect 690 1986 709 1988
rect 724 1986 770 1988
rect 690 1970 770 1986
rect 797 1984 832 1997
rect 873 1994 910 1997
rect 873 1992 915 1994
rect 802 1981 832 1984
rect 811 1977 818 1981
rect 818 1976 819 1977
rect 777 1970 787 1976
rect 536 1962 571 1970
rect 536 1936 537 1962
rect 544 1936 571 1962
rect 479 1918 509 1932
rect 536 1928 571 1936
rect 573 1962 614 1970
rect 573 1936 588 1962
rect 595 1936 614 1962
rect 678 1958 709 1970
rect 724 1958 827 1970
rect 839 1960 865 1986
rect 880 1981 910 1992
rect 942 1988 1004 2004
rect 942 1986 988 1988
rect 942 1970 1004 1986
rect 1016 1970 1022 2018
rect 1025 2010 1105 2018
rect 1025 2008 1044 2010
rect 1059 2008 1093 2010
rect 1025 1992 1105 2008
rect 1025 1970 1044 1992
rect 1059 1976 1089 1992
rect 1117 1986 1123 2060
rect 1126 1986 1145 2130
rect 1160 1986 1166 2130
rect 1175 2060 1188 2130
rect 1240 2126 1262 2130
rect 1233 2104 1262 2118
rect 1315 2104 1331 2118
rect 1369 2114 1375 2116
rect 1382 2114 1490 2130
rect 1497 2114 1503 2116
rect 1511 2114 1526 2130
rect 1592 2124 1611 2127
rect 1233 2102 1331 2104
rect 1358 2102 1526 2114
rect 1541 2104 1557 2118
rect 1592 2105 1614 2124
rect 1624 2118 1640 2119
rect 1623 2116 1640 2118
rect 1624 2111 1640 2116
rect 1614 2104 1620 2105
rect 1623 2104 1652 2111
rect 1541 2103 1652 2104
rect 1541 2102 1658 2103
rect 1217 2094 1268 2102
rect 1315 2094 1349 2102
rect 1217 2082 1242 2094
rect 1249 2082 1268 2094
rect 1322 2092 1349 2094
rect 1358 2092 1579 2102
rect 1614 2099 1620 2102
rect 1322 2088 1579 2092
rect 1217 2074 1268 2082
rect 1315 2074 1579 2088
rect 1623 2094 1658 2102
rect 1169 2026 1188 2060
rect 1233 2066 1262 2074
rect 1233 2060 1250 2066
rect 1233 2058 1267 2060
rect 1315 2058 1331 2074
rect 1332 2064 1540 2074
rect 1541 2064 1557 2074
rect 1605 2070 1620 2085
rect 1623 2082 1624 2094
rect 1631 2082 1658 2094
rect 1623 2074 1658 2082
rect 1623 2073 1652 2074
rect 1343 2060 1557 2064
rect 1358 2058 1557 2060
rect 1592 2060 1605 2070
rect 1623 2060 1640 2073
rect 1592 2058 1640 2060
rect 1234 2054 1267 2058
rect 1230 2052 1267 2054
rect 1230 2051 1297 2052
rect 1230 2046 1261 2051
rect 1267 2046 1297 2051
rect 1230 2042 1297 2046
rect 1203 2039 1297 2042
rect 1203 2032 1252 2039
rect 1203 2026 1233 2032
rect 1252 2027 1257 2032
rect 1169 2010 1249 2026
rect 1261 2018 1297 2039
rect 1358 2034 1547 2058
rect 1592 2057 1639 2058
rect 1605 2052 1639 2057
rect 1373 2031 1547 2034
rect 1366 2028 1547 2031
rect 1575 2051 1639 2052
rect 1169 2008 1188 2010
rect 1203 2008 1237 2010
rect 1169 1992 1249 2008
rect 1169 1986 1188 1992
rect 885 1960 988 1970
rect 839 1958 988 1960
rect 1009 1958 1044 1970
rect 678 1956 840 1958
rect 690 1936 709 1956
rect 724 1954 754 1956
rect 573 1928 614 1936
rect 696 1932 709 1936
rect 761 1940 840 1956
rect 872 1956 1044 1958
rect 872 1940 951 1956
rect 958 1954 988 1956
rect 536 1918 565 1928
rect 579 1918 608 1928
rect 623 1918 653 1932
rect 696 1918 739 1932
rect 761 1928 951 1940
rect 1016 1936 1022 1956
rect 746 1918 776 1928
rect 777 1918 935 1928
rect 939 1918 969 1928
rect 973 1918 1003 1932
rect 1031 1918 1044 1956
rect 1116 1970 1145 1986
rect 1159 1970 1188 1986
rect 1203 1976 1233 1992
rect 1261 1970 1267 2018
rect 1270 2012 1289 2018
rect 1304 2012 1334 2020
rect 1270 2004 1334 2012
rect 1270 1988 1350 2004
rect 1366 1997 1428 2028
rect 1444 1997 1506 2028
rect 1575 2026 1624 2051
rect 1639 2026 1669 2042
rect 1538 2012 1568 2020
rect 1575 2018 1685 2026
rect 1538 2004 1583 2012
rect 1270 1986 1289 1988
rect 1304 1986 1350 1988
rect 1270 1970 1350 1986
rect 1377 1984 1412 1997
rect 1453 1994 1490 1997
rect 1453 1992 1495 1994
rect 1382 1981 1412 1984
rect 1391 1977 1398 1981
rect 1398 1976 1399 1977
rect 1357 1970 1367 1976
rect 1116 1962 1151 1970
rect 1116 1936 1117 1962
rect 1124 1936 1151 1962
rect 1059 1918 1089 1932
rect 1116 1928 1151 1936
rect 1153 1962 1194 1970
rect 1153 1936 1168 1962
rect 1175 1936 1194 1962
rect 1258 1958 1289 1970
rect 1304 1958 1407 1970
rect 1419 1960 1445 1986
rect 1460 1981 1490 1992
rect 1522 1988 1584 2004
rect 1522 1986 1568 1988
rect 1522 1970 1584 1986
rect 1596 1970 1602 2018
rect 1605 2010 1685 2018
rect 1605 2008 1624 2010
rect 1639 2008 1673 2010
rect 1605 1992 1685 2008
rect 1605 1970 1624 1992
rect 1639 1976 1669 1992
rect 1697 1986 1703 2060
rect 1706 1986 1725 2130
rect 1740 1986 1746 2130
rect 1755 2060 1768 2130
rect 1820 2126 1842 2130
rect 1813 2104 1842 2118
rect 1895 2104 1911 2118
rect 1949 2114 1955 2116
rect 1962 2114 2070 2130
rect 2077 2114 2083 2116
rect 2091 2114 2106 2130
rect 2172 2124 2191 2127
rect 1813 2102 1911 2104
rect 1938 2102 2106 2114
rect 2121 2104 2137 2118
rect 2172 2105 2194 2124
rect 2204 2118 2220 2119
rect 2203 2116 2220 2118
rect 2204 2111 2220 2116
rect 2194 2104 2200 2105
rect 2203 2104 2232 2111
rect 2121 2103 2232 2104
rect 2121 2102 2238 2103
rect 1797 2094 1848 2102
rect 1895 2094 1929 2102
rect 1797 2082 1822 2094
rect 1829 2082 1848 2094
rect 1902 2092 1929 2094
rect 1938 2092 2159 2102
rect 2194 2099 2200 2102
rect 1902 2088 2159 2092
rect 1797 2074 1848 2082
rect 1895 2074 2159 2088
rect 2203 2094 2238 2102
rect 1749 2026 1768 2060
rect 1813 2066 1842 2074
rect 1813 2060 1830 2066
rect 1813 2058 1847 2060
rect 1895 2058 1911 2074
rect 1912 2064 2120 2074
rect 2121 2064 2137 2074
rect 2185 2070 2200 2085
rect 2203 2082 2204 2094
rect 2211 2082 2238 2094
rect 2203 2074 2238 2082
rect 2203 2073 2232 2074
rect 1923 2060 2137 2064
rect 1938 2058 2137 2060
rect 2172 2060 2185 2070
rect 2203 2060 2220 2073
rect 2172 2058 2220 2060
rect 1814 2054 1847 2058
rect 1810 2052 1847 2054
rect 1810 2051 1877 2052
rect 1810 2046 1841 2051
rect 1847 2046 1877 2051
rect 1810 2042 1877 2046
rect 1783 2039 1877 2042
rect 1783 2032 1832 2039
rect 1783 2026 1813 2032
rect 1832 2027 1837 2032
rect 1749 2010 1829 2026
rect 1841 2018 1877 2039
rect 1938 2034 2127 2058
rect 2172 2057 2219 2058
rect 2185 2052 2219 2057
rect 1953 2031 2127 2034
rect 1946 2028 2127 2031
rect 2155 2051 2219 2052
rect 1749 2008 1768 2010
rect 1783 2008 1817 2010
rect 1749 1992 1829 2008
rect 1749 1986 1768 1992
rect 1465 1960 1568 1970
rect 1419 1958 1568 1960
rect 1589 1958 1624 1970
rect 1258 1956 1420 1958
rect 1270 1936 1289 1956
rect 1304 1954 1334 1956
rect 1153 1928 1194 1936
rect 1276 1932 1289 1936
rect 1341 1940 1420 1956
rect 1452 1956 1624 1958
rect 1452 1940 1531 1956
rect 1538 1954 1568 1956
rect 1116 1918 1145 1928
rect 1159 1918 1188 1928
rect 1203 1918 1233 1932
rect 1276 1918 1319 1932
rect 1341 1928 1531 1940
rect 1596 1936 1602 1956
rect 1326 1918 1356 1928
rect 1357 1918 1515 1928
rect 1519 1918 1549 1928
rect 1553 1918 1583 1932
rect 1611 1918 1624 1956
rect 1696 1970 1725 1986
rect 1739 1970 1768 1986
rect 1783 1976 1813 1992
rect 1841 1970 1847 2018
rect 1850 2012 1869 2018
rect 1884 2012 1914 2020
rect 1850 2004 1914 2012
rect 1850 1988 1930 2004
rect 1946 1997 2008 2028
rect 2024 1997 2086 2028
rect 2155 2026 2204 2051
rect 2219 2026 2249 2042
rect 2118 2012 2148 2020
rect 2155 2018 2265 2026
rect 2118 2004 2163 2012
rect 1850 1986 1869 1988
rect 1884 1986 1930 1988
rect 1850 1970 1930 1986
rect 1957 1984 1992 1997
rect 2033 1994 2070 1997
rect 2033 1992 2075 1994
rect 1962 1981 1992 1984
rect 1971 1977 1978 1981
rect 1978 1976 1979 1977
rect 1937 1970 1947 1976
rect 1696 1962 1731 1970
rect 1696 1936 1697 1962
rect 1704 1936 1731 1962
rect 1639 1918 1669 1932
rect 1696 1928 1731 1936
rect 1733 1962 1774 1970
rect 1733 1936 1748 1962
rect 1755 1936 1774 1962
rect 1838 1958 1869 1970
rect 1884 1958 1987 1970
rect 1999 1960 2025 1986
rect 2040 1981 2070 1992
rect 2102 1988 2164 2004
rect 2102 1986 2148 1988
rect 2102 1970 2164 1986
rect 2176 1970 2182 2018
rect 2185 2010 2265 2018
rect 2185 2008 2204 2010
rect 2219 2008 2253 2010
rect 2185 1992 2265 2008
rect 2185 1970 2204 1992
rect 2219 1976 2249 1992
rect 2277 1986 2283 2060
rect 2286 1986 2305 2130
rect 2320 1986 2326 2130
rect 2335 2060 2348 2130
rect 2400 2126 2422 2130
rect 2393 2104 2422 2118
rect 2475 2104 2491 2118
rect 2529 2114 2535 2116
rect 2542 2114 2650 2130
rect 2657 2114 2663 2116
rect 2671 2114 2686 2130
rect 2752 2124 2771 2127
rect 2393 2102 2491 2104
rect 2518 2102 2686 2114
rect 2701 2104 2717 2118
rect 2752 2105 2774 2124
rect 2784 2118 2800 2119
rect 2783 2116 2800 2118
rect 2784 2111 2800 2116
rect 2774 2104 2780 2105
rect 2783 2104 2812 2111
rect 2701 2103 2812 2104
rect 2701 2102 2818 2103
rect 2377 2094 2428 2102
rect 2475 2094 2509 2102
rect 2377 2082 2402 2094
rect 2409 2082 2428 2094
rect 2482 2092 2509 2094
rect 2518 2092 2739 2102
rect 2774 2099 2780 2102
rect 2482 2088 2739 2092
rect 2377 2074 2428 2082
rect 2475 2074 2739 2088
rect 2783 2094 2818 2102
rect 2329 2026 2348 2060
rect 2393 2066 2422 2074
rect 2393 2060 2410 2066
rect 2393 2058 2427 2060
rect 2475 2058 2491 2074
rect 2492 2064 2700 2074
rect 2701 2064 2717 2074
rect 2765 2070 2780 2085
rect 2783 2082 2784 2094
rect 2791 2082 2818 2094
rect 2783 2074 2818 2082
rect 2783 2073 2812 2074
rect 2503 2060 2717 2064
rect 2518 2058 2717 2060
rect 2752 2060 2765 2070
rect 2783 2060 2800 2073
rect 2752 2058 2800 2060
rect 2394 2054 2427 2058
rect 2390 2052 2427 2054
rect 2390 2051 2457 2052
rect 2390 2046 2421 2051
rect 2427 2046 2457 2051
rect 2390 2042 2457 2046
rect 2363 2039 2457 2042
rect 2363 2032 2412 2039
rect 2363 2026 2393 2032
rect 2412 2027 2417 2032
rect 2329 2010 2409 2026
rect 2421 2018 2457 2039
rect 2518 2034 2707 2058
rect 2752 2057 2799 2058
rect 2765 2052 2799 2057
rect 2533 2031 2707 2034
rect 2526 2028 2707 2031
rect 2735 2051 2799 2052
rect 2329 2008 2348 2010
rect 2363 2008 2397 2010
rect 2329 1992 2409 2008
rect 2329 1986 2348 1992
rect 2045 1960 2148 1970
rect 1999 1958 2148 1960
rect 2169 1958 2204 1970
rect 1838 1956 2000 1958
rect 1850 1936 1869 1956
rect 1884 1954 1914 1956
rect 1733 1928 1774 1936
rect 1856 1932 1869 1936
rect 1921 1940 2000 1956
rect 2032 1956 2204 1958
rect 2032 1940 2111 1956
rect 2118 1954 2148 1956
rect 1696 1918 1725 1928
rect 1739 1918 1768 1928
rect 1783 1918 1813 1932
rect 1856 1918 1899 1932
rect 1921 1928 2111 1940
rect 2176 1936 2182 1956
rect 1906 1918 1936 1928
rect 1937 1918 2095 1928
rect 2099 1918 2129 1928
rect 2133 1918 2163 1932
rect 2191 1918 2204 1956
rect 2276 1970 2305 1986
rect 2319 1970 2348 1986
rect 2363 1976 2393 1992
rect 2421 1970 2427 2018
rect 2430 2012 2449 2018
rect 2464 2012 2494 2020
rect 2430 2004 2494 2012
rect 2430 1988 2510 2004
rect 2526 1997 2588 2028
rect 2604 1997 2666 2028
rect 2735 2026 2784 2051
rect 2799 2026 2829 2042
rect 2698 2012 2728 2020
rect 2735 2018 2845 2026
rect 2698 2004 2743 2012
rect 2430 1986 2449 1988
rect 2464 1986 2510 1988
rect 2430 1970 2510 1986
rect 2537 1984 2572 1997
rect 2613 1994 2650 1997
rect 2613 1992 2655 1994
rect 2542 1981 2572 1984
rect 2551 1977 2558 1981
rect 2558 1976 2559 1977
rect 2517 1970 2527 1976
rect 2276 1962 2311 1970
rect 2276 1936 2277 1962
rect 2284 1936 2311 1962
rect 2219 1918 2249 1932
rect 2276 1928 2311 1936
rect 2313 1962 2354 1970
rect 2313 1936 2328 1962
rect 2335 1936 2354 1962
rect 2418 1958 2449 1970
rect 2464 1958 2567 1970
rect 2579 1960 2605 1986
rect 2620 1981 2650 1992
rect 2682 1988 2744 2004
rect 2682 1986 2728 1988
rect 2682 1970 2744 1986
rect 2756 1970 2762 2018
rect 2765 2010 2845 2018
rect 2765 2008 2784 2010
rect 2799 2008 2833 2010
rect 2765 1992 2845 2008
rect 2765 1970 2784 1992
rect 2799 1976 2829 1992
rect 2857 1986 2863 2060
rect 2866 1986 2885 2130
rect 2900 1986 2906 2130
rect 2915 2060 2928 2130
rect 2980 2126 3002 2130
rect 2973 2104 3002 2118
rect 3055 2104 3071 2118
rect 3109 2114 3115 2116
rect 3122 2114 3230 2130
rect 3237 2114 3243 2116
rect 3251 2114 3266 2130
rect 3332 2124 3351 2127
rect 2973 2102 3071 2104
rect 3098 2102 3266 2114
rect 3281 2104 3297 2118
rect 3332 2105 3354 2124
rect 3364 2118 3380 2119
rect 3363 2116 3380 2118
rect 3364 2111 3380 2116
rect 3354 2104 3360 2105
rect 3363 2104 3392 2111
rect 3281 2103 3392 2104
rect 3281 2102 3398 2103
rect 2957 2094 3008 2102
rect 3055 2094 3089 2102
rect 2957 2082 2982 2094
rect 2989 2082 3008 2094
rect 3062 2092 3089 2094
rect 3098 2092 3319 2102
rect 3354 2099 3360 2102
rect 3062 2088 3319 2092
rect 2957 2074 3008 2082
rect 3055 2074 3319 2088
rect 3363 2094 3398 2102
rect 2909 2026 2928 2060
rect 2973 2066 3002 2074
rect 2973 2060 2990 2066
rect 2973 2058 3007 2060
rect 3055 2058 3071 2074
rect 3072 2064 3280 2074
rect 3281 2064 3297 2074
rect 3345 2070 3360 2085
rect 3363 2082 3364 2094
rect 3371 2082 3398 2094
rect 3363 2074 3398 2082
rect 3363 2073 3392 2074
rect 3083 2060 3297 2064
rect 3098 2058 3297 2060
rect 3332 2060 3345 2070
rect 3363 2060 3380 2073
rect 3332 2058 3380 2060
rect 2974 2054 3007 2058
rect 2970 2052 3007 2054
rect 2970 2051 3037 2052
rect 2970 2046 3001 2051
rect 3007 2046 3037 2051
rect 2970 2042 3037 2046
rect 2943 2039 3037 2042
rect 2943 2032 2992 2039
rect 2943 2026 2973 2032
rect 2992 2027 2997 2032
rect 2909 2010 2989 2026
rect 3001 2018 3037 2039
rect 3098 2034 3287 2058
rect 3332 2057 3379 2058
rect 3345 2052 3379 2057
rect 3113 2031 3287 2034
rect 3106 2028 3287 2031
rect 3315 2051 3379 2052
rect 2909 2008 2928 2010
rect 2943 2008 2977 2010
rect 2909 1992 2989 2008
rect 2909 1986 2928 1992
rect 2625 1960 2728 1970
rect 2579 1958 2728 1960
rect 2749 1958 2784 1970
rect 2418 1956 2580 1958
rect 2430 1936 2449 1956
rect 2464 1954 2494 1956
rect 2313 1928 2354 1936
rect 2436 1932 2449 1936
rect 2501 1940 2580 1956
rect 2612 1956 2784 1958
rect 2612 1940 2691 1956
rect 2698 1954 2728 1956
rect 2276 1918 2305 1928
rect 2319 1918 2348 1928
rect 2363 1918 2393 1932
rect 2436 1918 2479 1932
rect 2501 1928 2691 1940
rect 2756 1936 2762 1956
rect 2486 1918 2516 1928
rect 2517 1918 2675 1928
rect 2679 1918 2709 1928
rect 2713 1918 2743 1932
rect 2771 1918 2784 1956
rect 2856 1970 2885 1986
rect 2899 1970 2928 1986
rect 2943 1976 2973 1992
rect 3001 1970 3007 2018
rect 3010 2012 3029 2018
rect 3044 2012 3074 2020
rect 3010 2004 3074 2012
rect 3010 1988 3090 2004
rect 3106 1997 3168 2028
rect 3184 1997 3246 2028
rect 3315 2026 3364 2051
rect 3379 2026 3409 2042
rect 3278 2012 3308 2020
rect 3315 2018 3425 2026
rect 3278 2004 3323 2012
rect 3010 1986 3029 1988
rect 3044 1986 3090 1988
rect 3010 1970 3090 1986
rect 3117 1984 3152 1997
rect 3193 1994 3230 1997
rect 3193 1992 3235 1994
rect 3122 1981 3152 1984
rect 3131 1977 3138 1981
rect 3138 1976 3139 1977
rect 3097 1970 3107 1976
rect 2856 1962 2891 1970
rect 2856 1936 2857 1962
rect 2864 1936 2891 1962
rect 2799 1918 2829 1932
rect 2856 1928 2891 1936
rect 2893 1962 2934 1970
rect 2893 1936 2908 1962
rect 2915 1936 2934 1962
rect 2998 1958 3029 1970
rect 3044 1958 3147 1970
rect 3159 1960 3185 1986
rect 3200 1981 3230 1992
rect 3262 1988 3324 2004
rect 3262 1986 3308 1988
rect 3262 1970 3324 1986
rect 3336 1970 3342 2018
rect 3345 2010 3425 2018
rect 3345 2008 3364 2010
rect 3379 2008 3413 2010
rect 3345 1992 3425 2008
rect 3345 1970 3364 1992
rect 3379 1976 3409 1992
rect 3437 1986 3443 2060
rect 3446 1986 3465 2130
rect 3480 1986 3486 2130
rect 3495 2060 3508 2130
rect 3560 2126 3582 2130
rect 3553 2104 3582 2118
rect 3635 2104 3651 2118
rect 3689 2114 3695 2116
rect 3702 2114 3810 2130
rect 3817 2114 3823 2116
rect 3831 2114 3846 2130
rect 3912 2124 3931 2127
rect 3553 2102 3651 2104
rect 3678 2102 3846 2114
rect 3861 2104 3877 2118
rect 3912 2105 3934 2124
rect 3944 2118 3960 2119
rect 3943 2116 3960 2118
rect 3944 2111 3960 2116
rect 3934 2104 3940 2105
rect 3943 2104 3972 2111
rect 3861 2103 3972 2104
rect 3861 2102 3978 2103
rect 3537 2094 3588 2102
rect 3635 2094 3669 2102
rect 3537 2082 3562 2094
rect 3569 2082 3588 2094
rect 3642 2092 3669 2094
rect 3678 2092 3899 2102
rect 3934 2099 3940 2102
rect 3642 2088 3899 2092
rect 3537 2074 3588 2082
rect 3635 2074 3899 2088
rect 3943 2094 3978 2102
rect 3489 2026 3508 2060
rect 3553 2066 3582 2074
rect 3553 2060 3570 2066
rect 3553 2058 3587 2060
rect 3635 2058 3651 2074
rect 3652 2064 3860 2074
rect 3861 2064 3877 2074
rect 3925 2070 3940 2085
rect 3943 2082 3944 2094
rect 3951 2082 3978 2094
rect 3943 2074 3978 2082
rect 3943 2073 3972 2074
rect 3663 2060 3877 2064
rect 3678 2058 3877 2060
rect 3912 2060 3925 2070
rect 3943 2060 3960 2073
rect 3912 2058 3960 2060
rect 3554 2054 3587 2058
rect 3550 2052 3587 2054
rect 3550 2051 3617 2052
rect 3550 2046 3581 2051
rect 3587 2046 3617 2051
rect 3550 2042 3617 2046
rect 3523 2039 3617 2042
rect 3523 2032 3572 2039
rect 3523 2026 3553 2032
rect 3572 2027 3577 2032
rect 3489 2010 3569 2026
rect 3581 2018 3617 2039
rect 3678 2034 3867 2058
rect 3912 2057 3959 2058
rect 3925 2052 3959 2057
rect 3693 2031 3867 2034
rect 3686 2028 3867 2031
rect 3895 2051 3959 2052
rect 3489 2008 3508 2010
rect 3523 2008 3557 2010
rect 3489 1992 3569 2008
rect 3489 1986 3508 1992
rect 3205 1960 3308 1970
rect 3159 1958 3308 1960
rect 3329 1958 3364 1970
rect 2998 1956 3160 1958
rect 3010 1936 3029 1956
rect 3044 1954 3074 1956
rect 2893 1928 2934 1936
rect 3016 1932 3029 1936
rect 3081 1940 3160 1956
rect 3192 1956 3364 1958
rect 3192 1940 3271 1956
rect 3278 1954 3308 1956
rect 2856 1918 2885 1928
rect 2899 1918 2928 1928
rect 2943 1918 2973 1932
rect 3016 1918 3059 1932
rect 3081 1928 3271 1940
rect 3336 1936 3342 1956
rect 3066 1918 3096 1928
rect 3097 1918 3255 1928
rect 3259 1918 3289 1928
rect 3293 1918 3323 1932
rect 3351 1918 3364 1956
rect 3436 1970 3465 1986
rect 3479 1970 3508 1986
rect 3523 1976 3553 1992
rect 3581 1970 3587 2018
rect 3590 2012 3609 2018
rect 3624 2012 3654 2020
rect 3590 2004 3654 2012
rect 3590 1988 3670 2004
rect 3686 1997 3748 2028
rect 3764 1997 3826 2028
rect 3895 2026 3944 2051
rect 3959 2026 3989 2042
rect 3858 2012 3888 2020
rect 3895 2018 4005 2026
rect 3858 2004 3903 2012
rect 3590 1986 3609 1988
rect 3624 1986 3670 1988
rect 3590 1970 3670 1986
rect 3697 1984 3732 1997
rect 3773 1994 3810 1997
rect 3773 1992 3815 1994
rect 3702 1981 3732 1984
rect 3711 1977 3718 1981
rect 3718 1976 3719 1977
rect 3677 1970 3687 1976
rect 3436 1962 3471 1970
rect 3436 1936 3437 1962
rect 3444 1936 3471 1962
rect 3379 1918 3409 1932
rect 3436 1928 3471 1936
rect 3473 1962 3514 1970
rect 3473 1936 3488 1962
rect 3495 1936 3514 1962
rect 3578 1958 3609 1970
rect 3624 1958 3727 1970
rect 3739 1960 3765 1986
rect 3780 1981 3810 1992
rect 3842 1988 3904 2004
rect 3842 1986 3888 1988
rect 3842 1970 3904 1986
rect 3916 1970 3922 2018
rect 3925 2010 4005 2018
rect 3925 2008 3944 2010
rect 3959 2008 3993 2010
rect 3925 1992 4005 2008
rect 3925 1970 3944 1992
rect 3959 1976 3989 1992
rect 4017 1986 4023 2060
rect 4026 1986 4045 2130
rect 4060 1986 4066 2130
rect 4075 2060 4088 2130
rect 4140 2126 4162 2130
rect 4133 2104 4162 2118
rect 4215 2104 4231 2118
rect 4269 2114 4275 2116
rect 4282 2114 4390 2130
rect 4397 2114 4403 2116
rect 4411 2114 4426 2130
rect 4492 2124 4511 2127
rect 4133 2102 4231 2104
rect 4258 2102 4426 2114
rect 4441 2104 4457 2118
rect 4492 2105 4514 2124
rect 4524 2118 4540 2119
rect 4523 2116 4540 2118
rect 4524 2111 4540 2116
rect 4514 2104 4520 2105
rect 4523 2104 4552 2111
rect 4441 2103 4552 2104
rect 4441 2102 4558 2103
rect 4117 2094 4168 2102
rect 4215 2094 4249 2102
rect 4117 2082 4142 2094
rect 4149 2082 4168 2094
rect 4222 2092 4249 2094
rect 4258 2092 4479 2102
rect 4514 2099 4520 2102
rect 4222 2088 4479 2092
rect 4117 2074 4168 2082
rect 4215 2074 4479 2088
rect 4523 2094 4558 2102
rect 4069 2026 4088 2060
rect 4133 2066 4162 2074
rect 4133 2060 4150 2066
rect 4133 2058 4167 2060
rect 4215 2058 4231 2074
rect 4232 2064 4440 2074
rect 4441 2064 4457 2074
rect 4505 2070 4520 2085
rect 4523 2082 4524 2094
rect 4531 2082 4558 2094
rect 4523 2074 4558 2082
rect 4523 2073 4552 2074
rect 4243 2060 4457 2064
rect 4258 2058 4457 2060
rect 4492 2060 4505 2070
rect 4523 2060 4540 2073
rect 4492 2058 4540 2060
rect 4134 2054 4167 2058
rect 4130 2052 4167 2054
rect 4130 2051 4197 2052
rect 4130 2046 4161 2051
rect 4167 2046 4197 2051
rect 4130 2042 4197 2046
rect 4103 2039 4197 2042
rect 4103 2032 4152 2039
rect 4103 2026 4133 2032
rect 4152 2027 4157 2032
rect 4069 2010 4149 2026
rect 4161 2018 4197 2039
rect 4258 2034 4447 2058
rect 4492 2057 4539 2058
rect 4505 2052 4539 2057
rect 4273 2031 4447 2034
rect 4266 2028 4447 2031
rect 4475 2051 4539 2052
rect 4069 2008 4088 2010
rect 4103 2008 4137 2010
rect 4069 1992 4149 2008
rect 4069 1986 4088 1992
rect 3785 1960 3888 1970
rect 3739 1958 3888 1960
rect 3909 1958 3944 1970
rect 3578 1956 3740 1958
rect 3590 1936 3609 1956
rect 3624 1954 3654 1956
rect 3473 1928 3514 1936
rect 3596 1932 3609 1936
rect 3661 1940 3740 1956
rect 3772 1956 3944 1958
rect 3772 1940 3851 1956
rect 3858 1954 3888 1956
rect 3436 1918 3465 1928
rect 3479 1918 3508 1928
rect 3523 1918 3553 1932
rect 3596 1918 3639 1932
rect 3661 1928 3851 1940
rect 3916 1936 3922 1956
rect 3646 1918 3676 1928
rect 3677 1918 3835 1928
rect 3839 1918 3869 1928
rect 3873 1918 3903 1932
rect 3931 1918 3944 1956
rect 4016 1970 4045 1986
rect 4059 1970 4088 1986
rect 4103 1976 4133 1992
rect 4161 1970 4167 2018
rect 4170 2012 4189 2018
rect 4204 2012 4234 2020
rect 4170 2004 4234 2012
rect 4170 1988 4250 2004
rect 4266 1997 4328 2028
rect 4344 1997 4406 2028
rect 4475 2026 4524 2051
rect 4539 2026 4569 2042
rect 4438 2012 4468 2020
rect 4475 2018 4585 2026
rect 4438 2004 4483 2012
rect 4170 1986 4189 1988
rect 4204 1986 4250 1988
rect 4170 1970 4250 1986
rect 4277 1984 4312 1997
rect 4353 1994 4390 1997
rect 4353 1992 4395 1994
rect 4282 1981 4312 1984
rect 4291 1977 4298 1981
rect 4298 1976 4299 1977
rect 4257 1970 4267 1976
rect 4016 1962 4051 1970
rect 4016 1936 4017 1962
rect 4024 1936 4051 1962
rect 3959 1918 3989 1932
rect 4016 1928 4051 1936
rect 4053 1962 4094 1970
rect 4053 1936 4068 1962
rect 4075 1936 4094 1962
rect 4158 1958 4189 1970
rect 4204 1958 4307 1970
rect 4319 1960 4345 1986
rect 4360 1981 4390 1992
rect 4422 1988 4484 2004
rect 4422 1986 4468 1988
rect 4422 1970 4484 1986
rect 4496 1970 4502 2018
rect 4505 2010 4585 2018
rect 4505 2008 4524 2010
rect 4539 2008 4573 2010
rect 4505 1992 4585 2008
rect 4505 1970 4524 1992
rect 4539 1976 4569 1992
rect 4597 1986 4603 2060
rect 4606 1986 4625 2130
rect 4640 1986 4646 2130
rect 4655 2060 4668 2130
rect 4720 2126 4742 2130
rect 4713 2104 4742 2118
rect 4795 2104 4811 2118
rect 4849 2114 4855 2116
rect 4862 2114 4970 2130
rect 4977 2114 4983 2116
rect 4991 2114 5006 2130
rect 5072 2124 5091 2127
rect 4713 2102 4811 2104
rect 4838 2102 5006 2114
rect 5021 2104 5037 2118
rect 5072 2105 5094 2124
rect 5104 2118 5120 2119
rect 5103 2116 5120 2118
rect 5104 2111 5120 2116
rect 5094 2104 5100 2105
rect 5103 2104 5132 2111
rect 5021 2103 5132 2104
rect 5021 2102 5138 2103
rect 4697 2094 4748 2102
rect 4795 2094 4829 2102
rect 4697 2082 4722 2094
rect 4729 2082 4748 2094
rect 4802 2092 4829 2094
rect 4838 2092 5059 2102
rect 5094 2099 5100 2102
rect 4802 2088 5059 2092
rect 4697 2074 4748 2082
rect 4795 2074 5059 2088
rect 5103 2094 5138 2102
rect 4649 2026 4668 2060
rect 4713 2066 4742 2074
rect 4713 2060 4730 2066
rect 4713 2058 4747 2060
rect 4795 2058 4811 2074
rect 4812 2064 5020 2074
rect 5021 2064 5037 2074
rect 5085 2070 5100 2085
rect 5103 2082 5104 2094
rect 5111 2082 5138 2094
rect 5103 2074 5138 2082
rect 5103 2073 5132 2074
rect 4823 2060 5037 2064
rect 4838 2058 5037 2060
rect 5072 2060 5085 2070
rect 5103 2060 5120 2073
rect 5072 2058 5120 2060
rect 4714 2054 4747 2058
rect 4710 2052 4747 2054
rect 4710 2051 4777 2052
rect 4710 2046 4741 2051
rect 4747 2046 4777 2051
rect 4710 2042 4777 2046
rect 4683 2039 4777 2042
rect 4683 2032 4732 2039
rect 4683 2026 4713 2032
rect 4732 2027 4737 2032
rect 4649 2010 4729 2026
rect 4741 2018 4777 2039
rect 4838 2034 5027 2058
rect 5072 2057 5119 2058
rect 5085 2052 5119 2057
rect 4853 2031 5027 2034
rect 4846 2028 5027 2031
rect 5055 2051 5119 2052
rect 4649 2008 4668 2010
rect 4683 2008 4717 2010
rect 4649 1992 4729 2008
rect 4649 1986 4668 1992
rect 4365 1960 4468 1970
rect 4319 1958 4468 1960
rect 4489 1958 4524 1970
rect 4158 1956 4320 1958
rect 4170 1936 4189 1956
rect 4204 1954 4234 1956
rect 4053 1928 4094 1936
rect 4176 1932 4189 1936
rect 4241 1940 4320 1956
rect 4352 1956 4524 1958
rect 4352 1940 4431 1956
rect 4438 1954 4468 1956
rect 4016 1918 4045 1928
rect 4059 1918 4088 1928
rect 4103 1918 4133 1932
rect 4176 1918 4219 1932
rect 4241 1928 4431 1940
rect 4496 1936 4502 1956
rect 4226 1918 4256 1928
rect 4257 1918 4415 1928
rect 4419 1918 4449 1928
rect 4453 1918 4483 1932
rect 4511 1918 4524 1956
rect 4596 1970 4625 1986
rect 4639 1970 4668 1986
rect 4683 1976 4713 1992
rect 4741 1970 4747 2018
rect 4750 2012 4769 2018
rect 4784 2012 4814 2020
rect 4750 2004 4814 2012
rect 4750 1988 4830 2004
rect 4846 1997 4908 2028
rect 4924 1997 4986 2028
rect 5055 2026 5104 2051
rect 5119 2026 5149 2042
rect 5018 2012 5048 2020
rect 5055 2018 5165 2026
rect 5018 2004 5063 2012
rect 4750 1986 4769 1988
rect 4784 1986 4830 1988
rect 4750 1970 4830 1986
rect 4857 1984 4892 1997
rect 4933 1994 4970 1997
rect 4933 1992 4975 1994
rect 4862 1981 4892 1984
rect 4871 1977 4878 1981
rect 4878 1976 4879 1977
rect 4837 1970 4847 1976
rect 4596 1962 4631 1970
rect 4596 1936 4597 1962
rect 4604 1936 4631 1962
rect 4539 1918 4569 1932
rect 4596 1928 4631 1936
rect 4633 1962 4674 1970
rect 4633 1936 4648 1962
rect 4655 1936 4674 1962
rect 4738 1958 4769 1970
rect 4784 1958 4887 1970
rect 4899 1960 4925 1986
rect 4940 1981 4970 1992
rect 5002 1988 5064 2004
rect 5002 1986 5048 1988
rect 5002 1970 5064 1986
rect 5076 1970 5082 2018
rect 5085 2010 5165 2018
rect 5085 2008 5104 2010
rect 5119 2008 5153 2010
rect 5085 1992 5165 2008
rect 5085 1970 5104 1992
rect 5119 1976 5149 1992
rect 5177 1986 5183 2060
rect 5186 1986 5205 2130
rect 5220 1986 5226 2130
rect 5235 2060 5248 2130
rect 5300 2126 5322 2130
rect 5293 2104 5322 2118
rect 5375 2104 5391 2118
rect 5429 2114 5435 2116
rect 5442 2114 5550 2130
rect 5557 2114 5563 2116
rect 5571 2114 5586 2130
rect 5652 2124 5671 2127
rect 5293 2102 5391 2104
rect 5418 2102 5586 2114
rect 5601 2104 5617 2118
rect 5652 2105 5674 2124
rect 5684 2118 5700 2119
rect 5683 2116 5700 2118
rect 5684 2111 5700 2116
rect 5674 2104 5680 2105
rect 5683 2104 5712 2111
rect 5601 2103 5712 2104
rect 5601 2102 5718 2103
rect 5277 2094 5328 2102
rect 5375 2094 5409 2102
rect 5277 2082 5302 2094
rect 5309 2082 5328 2094
rect 5382 2092 5409 2094
rect 5418 2092 5639 2102
rect 5674 2099 5680 2102
rect 5382 2088 5639 2092
rect 5277 2074 5328 2082
rect 5375 2074 5639 2088
rect 5683 2094 5718 2102
rect 5229 2026 5248 2060
rect 5293 2066 5322 2074
rect 5293 2060 5310 2066
rect 5293 2058 5327 2060
rect 5375 2058 5391 2074
rect 5392 2064 5600 2074
rect 5601 2064 5617 2074
rect 5665 2070 5680 2085
rect 5683 2082 5684 2094
rect 5691 2082 5718 2094
rect 5683 2074 5718 2082
rect 5683 2073 5712 2074
rect 5403 2060 5617 2064
rect 5418 2058 5617 2060
rect 5652 2060 5665 2070
rect 5683 2060 5700 2073
rect 5652 2058 5700 2060
rect 5294 2054 5327 2058
rect 5290 2052 5327 2054
rect 5290 2051 5357 2052
rect 5290 2046 5321 2051
rect 5327 2046 5357 2051
rect 5290 2042 5357 2046
rect 5263 2039 5357 2042
rect 5263 2032 5312 2039
rect 5263 2026 5293 2032
rect 5312 2027 5317 2032
rect 5229 2010 5309 2026
rect 5321 2018 5357 2039
rect 5418 2034 5607 2058
rect 5652 2057 5699 2058
rect 5665 2052 5699 2057
rect 5433 2031 5607 2034
rect 5426 2028 5607 2031
rect 5635 2051 5699 2052
rect 5229 2008 5248 2010
rect 5263 2008 5297 2010
rect 5229 1992 5309 2008
rect 5229 1986 5248 1992
rect 4945 1960 5048 1970
rect 4899 1958 5048 1960
rect 5069 1958 5104 1970
rect 4738 1956 4900 1958
rect 4750 1936 4769 1956
rect 4784 1954 4814 1956
rect 4633 1928 4674 1936
rect 4756 1932 4769 1936
rect 4821 1940 4900 1956
rect 4932 1956 5104 1958
rect 4932 1940 5011 1956
rect 5018 1954 5048 1956
rect 4596 1918 4625 1928
rect 4639 1918 4668 1928
rect 4683 1918 4713 1932
rect 4756 1918 4799 1932
rect 4821 1928 5011 1940
rect 5076 1936 5082 1956
rect 4806 1918 4836 1928
rect 4837 1918 4995 1928
rect 4999 1918 5029 1928
rect 5033 1918 5063 1932
rect 5091 1918 5104 1956
rect 5176 1970 5205 1986
rect 5219 1970 5248 1986
rect 5263 1976 5293 1992
rect 5321 1970 5327 2018
rect 5330 2012 5349 2018
rect 5364 2012 5394 2020
rect 5330 2004 5394 2012
rect 5330 1988 5410 2004
rect 5426 1997 5488 2028
rect 5504 1997 5566 2028
rect 5635 2026 5684 2051
rect 5699 2026 5729 2042
rect 5598 2012 5628 2020
rect 5635 2018 5745 2026
rect 5598 2004 5643 2012
rect 5330 1986 5349 1988
rect 5364 1986 5410 1988
rect 5330 1970 5410 1986
rect 5437 1984 5472 1997
rect 5513 1994 5550 1997
rect 5513 1992 5555 1994
rect 5442 1981 5472 1984
rect 5451 1977 5458 1981
rect 5458 1976 5459 1977
rect 5417 1970 5427 1976
rect 5176 1962 5211 1970
rect 5176 1936 5177 1962
rect 5184 1936 5211 1962
rect 5119 1918 5149 1932
rect 5176 1928 5211 1936
rect 5213 1962 5254 1970
rect 5213 1936 5228 1962
rect 5235 1936 5254 1962
rect 5318 1958 5349 1970
rect 5364 1958 5467 1970
rect 5479 1960 5505 1986
rect 5520 1981 5550 1992
rect 5582 1988 5644 2004
rect 5582 1986 5628 1988
rect 5582 1970 5644 1986
rect 5656 1970 5662 2018
rect 5665 2010 5745 2018
rect 5665 2008 5684 2010
rect 5699 2008 5733 2010
rect 5665 1992 5745 2008
rect 5665 1970 5684 1992
rect 5699 1976 5729 1992
rect 5757 1986 5763 2060
rect 5766 1986 5785 2130
rect 5800 1986 5806 2130
rect 5815 2060 5828 2130
rect 5880 2126 5902 2130
rect 5873 2104 5902 2118
rect 5955 2104 5971 2118
rect 6009 2114 6015 2116
rect 6022 2114 6130 2130
rect 6137 2114 6143 2116
rect 6151 2114 6166 2130
rect 6232 2124 6251 2127
rect 5873 2102 5971 2104
rect 5998 2102 6166 2114
rect 6181 2104 6197 2118
rect 6232 2105 6254 2124
rect 6264 2118 6280 2119
rect 6263 2116 6280 2118
rect 6264 2111 6280 2116
rect 6254 2104 6260 2105
rect 6263 2104 6292 2111
rect 6181 2103 6292 2104
rect 6181 2102 6298 2103
rect 5857 2094 5908 2102
rect 5955 2094 5989 2102
rect 5857 2082 5882 2094
rect 5889 2082 5908 2094
rect 5962 2092 5989 2094
rect 5998 2092 6219 2102
rect 6254 2099 6260 2102
rect 5962 2088 6219 2092
rect 5857 2074 5908 2082
rect 5955 2074 6219 2088
rect 6263 2094 6298 2102
rect 5809 2026 5828 2060
rect 5873 2066 5902 2074
rect 5873 2060 5890 2066
rect 5873 2058 5907 2060
rect 5955 2058 5971 2074
rect 5972 2064 6180 2074
rect 6181 2064 6197 2074
rect 6245 2070 6260 2085
rect 6263 2082 6264 2094
rect 6271 2082 6298 2094
rect 6263 2074 6298 2082
rect 6263 2073 6292 2074
rect 5983 2060 6197 2064
rect 5998 2058 6197 2060
rect 6232 2060 6245 2070
rect 6263 2060 6280 2073
rect 6232 2058 6280 2060
rect 5874 2054 5907 2058
rect 5870 2052 5907 2054
rect 5870 2051 5937 2052
rect 5870 2046 5901 2051
rect 5907 2046 5937 2051
rect 5870 2042 5937 2046
rect 5843 2039 5937 2042
rect 5843 2032 5892 2039
rect 5843 2026 5873 2032
rect 5892 2027 5897 2032
rect 5809 2010 5889 2026
rect 5901 2018 5937 2039
rect 5998 2034 6187 2058
rect 6232 2057 6279 2058
rect 6245 2052 6279 2057
rect 6013 2031 6187 2034
rect 6006 2028 6187 2031
rect 6215 2051 6279 2052
rect 5809 2008 5828 2010
rect 5843 2008 5877 2010
rect 5809 1992 5889 2008
rect 5809 1986 5828 1992
rect 5525 1960 5628 1970
rect 5479 1958 5628 1960
rect 5649 1958 5684 1970
rect 5318 1956 5480 1958
rect 5330 1936 5349 1956
rect 5364 1954 5394 1956
rect 5213 1928 5254 1936
rect 5336 1932 5349 1936
rect 5401 1940 5480 1956
rect 5512 1956 5684 1958
rect 5512 1940 5591 1956
rect 5598 1954 5628 1956
rect 5176 1918 5205 1928
rect 5219 1918 5248 1928
rect 5263 1918 5293 1932
rect 5336 1918 5379 1932
rect 5401 1928 5591 1940
rect 5656 1936 5662 1956
rect 5386 1918 5416 1928
rect 5417 1918 5575 1928
rect 5579 1918 5609 1928
rect 5613 1918 5643 1932
rect 5671 1918 5684 1956
rect 5756 1970 5785 1986
rect 5799 1970 5828 1986
rect 5843 1976 5873 1992
rect 5901 1970 5907 2018
rect 5910 2012 5929 2018
rect 5944 2012 5974 2020
rect 5910 2004 5974 2012
rect 5910 1988 5990 2004
rect 6006 1997 6068 2028
rect 6084 1997 6146 2028
rect 6215 2026 6264 2051
rect 6279 2026 6309 2042
rect 6178 2012 6208 2020
rect 6215 2018 6325 2026
rect 6178 2004 6223 2012
rect 5910 1986 5929 1988
rect 5944 1986 5990 1988
rect 5910 1970 5990 1986
rect 6017 1984 6052 1997
rect 6093 1994 6130 1997
rect 6093 1992 6135 1994
rect 6022 1981 6052 1984
rect 6031 1977 6038 1981
rect 6038 1976 6039 1977
rect 5997 1970 6007 1976
rect 5756 1962 5791 1970
rect 5756 1936 5757 1962
rect 5764 1936 5791 1962
rect 5699 1918 5729 1932
rect 5756 1928 5791 1936
rect 5793 1962 5834 1970
rect 5793 1936 5808 1962
rect 5815 1936 5834 1962
rect 5898 1958 5929 1970
rect 5944 1958 6047 1970
rect 6059 1960 6085 1986
rect 6100 1981 6130 1992
rect 6162 1988 6224 2004
rect 6162 1986 6208 1988
rect 6162 1970 6224 1986
rect 6236 1970 6242 2018
rect 6245 2010 6325 2018
rect 6245 2008 6264 2010
rect 6279 2008 6313 2010
rect 6245 1992 6325 2008
rect 6245 1970 6264 1992
rect 6279 1976 6309 1992
rect 6337 1986 6343 2060
rect 6346 1986 6365 2130
rect 6380 1986 6386 2130
rect 6395 2060 6408 2130
rect 6460 2126 6482 2130
rect 6453 2104 6482 2118
rect 6535 2104 6551 2118
rect 6589 2114 6595 2116
rect 6602 2114 6710 2130
rect 6717 2114 6723 2116
rect 6731 2114 6746 2130
rect 6812 2124 6831 2127
rect 6453 2102 6551 2104
rect 6578 2102 6746 2114
rect 6761 2104 6777 2118
rect 6812 2105 6834 2124
rect 6844 2118 6860 2119
rect 6843 2116 6860 2118
rect 6844 2111 6860 2116
rect 6834 2104 6840 2105
rect 6843 2104 6872 2111
rect 6761 2103 6872 2104
rect 6761 2102 6878 2103
rect 6437 2094 6488 2102
rect 6535 2094 6569 2102
rect 6437 2082 6462 2094
rect 6469 2082 6488 2094
rect 6542 2092 6569 2094
rect 6578 2092 6799 2102
rect 6834 2099 6840 2102
rect 6542 2088 6799 2092
rect 6437 2074 6488 2082
rect 6535 2074 6799 2088
rect 6843 2094 6878 2102
rect 6389 2026 6408 2060
rect 6453 2066 6482 2074
rect 6453 2060 6470 2066
rect 6453 2058 6487 2060
rect 6535 2058 6551 2074
rect 6552 2064 6760 2074
rect 6761 2064 6777 2074
rect 6825 2070 6840 2085
rect 6843 2082 6844 2094
rect 6851 2082 6878 2094
rect 6843 2074 6878 2082
rect 6843 2073 6872 2074
rect 6563 2060 6777 2064
rect 6578 2058 6777 2060
rect 6812 2060 6825 2070
rect 6843 2060 6860 2073
rect 6812 2058 6860 2060
rect 6454 2054 6487 2058
rect 6450 2052 6487 2054
rect 6450 2051 6517 2052
rect 6450 2046 6481 2051
rect 6487 2046 6517 2051
rect 6450 2042 6517 2046
rect 6423 2039 6517 2042
rect 6423 2032 6472 2039
rect 6423 2026 6453 2032
rect 6472 2027 6477 2032
rect 6389 2010 6469 2026
rect 6481 2018 6517 2039
rect 6578 2034 6767 2058
rect 6812 2057 6859 2058
rect 6825 2052 6859 2057
rect 6593 2031 6767 2034
rect 6586 2028 6767 2031
rect 6795 2051 6859 2052
rect 6389 2008 6408 2010
rect 6423 2008 6457 2010
rect 6389 1992 6469 2008
rect 6389 1986 6408 1992
rect 6105 1960 6208 1970
rect 6059 1958 6208 1960
rect 6229 1958 6264 1970
rect 5898 1956 6060 1958
rect 5910 1936 5929 1956
rect 5944 1954 5974 1956
rect 5793 1928 5834 1936
rect 5916 1932 5929 1936
rect 5981 1940 6060 1956
rect 6092 1956 6264 1958
rect 6092 1940 6171 1956
rect 6178 1954 6208 1956
rect 5756 1918 5785 1928
rect 5799 1918 5828 1928
rect 5843 1918 5873 1932
rect 5916 1918 5959 1932
rect 5981 1928 6171 1940
rect 6236 1936 6242 1956
rect 5966 1918 5996 1928
rect 5997 1918 6155 1928
rect 6159 1918 6189 1928
rect 6193 1918 6223 1932
rect 6251 1918 6264 1956
rect 6336 1970 6365 1986
rect 6379 1970 6408 1986
rect 6423 1976 6453 1992
rect 6481 1970 6487 2018
rect 6490 2012 6509 2018
rect 6524 2012 6554 2020
rect 6490 2004 6554 2012
rect 6490 1988 6570 2004
rect 6586 1997 6648 2028
rect 6664 1997 6726 2028
rect 6795 2026 6844 2051
rect 6859 2026 6889 2042
rect 6758 2012 6788 2020
rect 6795 2018 6905 2026
rect 6758 2004 6803 2012
rect 6490 1986 6509 1988
rect 6524 1986 6570 1988
rect 6490 1970 6570 1986
rect 6597 1984 6632 1997
rect 6673 1994 6710 1997
rect 6673 1992 6715 1994
rect 6602 1981 6632 1984
rect 6611 1977 6618 1981
rect 6618 1976 6619 1977
rect 6577 1970 6587 1976
rect 6336 1962 6371 1970
rect 6336 1936 6337 1962
rect 6344 1936 6371 1962
rect 6279 1918 6309 1932
rect 6336 1928 6371 1936
rect 6373 1962 6414 1970
rect 6373 1936 6388 1962
rect 6395 1936 6414 1962
rect 6478 1958 6509 1970
rect 6524 1958 6627 1970
rect 6639 1960 6665 1986
rect 6680 1981 6710 1992
rect 6742 1988 6804 2004
rect 6742 1986 6788 1988
rect 6742 1970 6804 1986
rect 6816 1970 6822 2018
rect 6825 2010 6905 2018
rect 6825 2008 6844 2010
rect 6859 2008 6893 2010
rect 6825 1992 6905 2008
rect 6825 1970 6844 1992
rect 6859 1976 6889 1992
rect 6917 1986 6923 2060
rect 6926 1986 6945 2130
rect 6960 1986 6966 2130
rect 6975 2060 6988 2130
rect 7040 2126 7062 2130
rect 7033 2104 7062 2118
rect 7115 2104 7131 2118
rect 7169 2114 7175 2116
rect 7182 2114 7290 2130
rect 7297 2114 7303 2116
rect 7311 2114 7326 2130
rect 7392 2124 7411 2127
rect 7033 2102 7131 2104
rect 7158 2102 7326 2114
rect 7341 2104 7357 2118
rect 7392 2105 7414 2124
rect 7424 2118 7440 2119
rect 7423 2116 7440 2118
rect 7424 2111 7440 2116
rect 7414 2104 7420 2105
rect 7423 2104 7452 2111
rect 7341 2103 7452 2104
rect 7341 2102 7458 2103
rect 7017 2094 7068 2102
rect 7115 2094 7149 2102
rect 7017 2082 7042 2094
rect 7049 2082 7068 2094
rect 7122 2092 7149 2094
rect 7158 2092 7379 2102
rect 7414 2099 7420 2102
rect 7122 2088 7379 2092
rect 7017 2074 7068 2082
rect 7115 2074 7379 2088
rect 7423 2094 7458 2102
rect 6969 2026 6988 2060
rect 7033 2066 7062 2074
rect 7033 2060 7050 2066
rect 7033 2058 7067 2060
rect 7115 2058 7131 2074
rect 7132 2064 7340 2074
rect 7341 2064 7357 2074
rect 7405 2070 7420 2085
rect 7423 2082 7424 2094
rect 7431 2082 7458 2094
rect 7423 2074 7458 2082
rect 7423 2073 7452 2074
rect 7143 2060 7357 2064
rect 7158 2058 7357 2060
rect 7392 2060 7405 2070
rect 7423 2060 7440 2073
rect 7392 2058 7440 2060
rect 7034 2054 7067 2058
rect 7030 2052 7067 2054
rect 7030 2051 7097 2052
rect 7030 2046 7061 2051
rect 7067 2046 7097 2051
rect 7030 2042 7097 2046
rect 7003 2039 7097 2042
rect 7003 2032 7052 2039
rect 7003 2026 7033 2032
rect 7052 2027 7057 2032
rect 6969 2010 7049 2026
rect 7061 2018 7097 2039
rect 7158 2034 7347 2058
rect 7392 2057 7439 2058
rect 7405 2052 7439 2057
rect 7173 2031 7347 2034
rect 7166 2028 7347 2031
rect 7375 2051 7439 2052
rect 6969 2008 6988 2010
rect 7003 2008 7037 2010
rect 6969 1992 7049 2008
rect 6969 1986 6988 1992
rect 6685 1960 6788 1970
rect 6639 1958 6788 1960
rect 6809 1958 6844 1970
rect 6478 1956 6640 1958
rect 6490 1936 6509 1956
rect 6524 1954 6554 1956
rect 6373 1928 6414 1936
rect 6496 1932 6509 1936
rect 6561 1940 6640 1956
rect 6672 1956 6844 1958
rect 6672 1940 6751 1956
rect 6758 1954 6788 1956
rect 6336 1918 6365 1928
rect 6379 1918 6408 1928
rect 6423 1918 6453 1932
rect 6496 1918 6539 1932
rect 6561 1928 6751 1940
rect 6816 1936 6822 1956
rect 6546 1918 6576 1928
rect 6577 1918 6735 1928
rect 6739 1918 6769 1928
rect 6773 1918 6803 1932
rect 6831 1918 6844 1956
rect 6916 1970 6945 1986
rect 6959 1970 6988 1986
rect 7003 1976 7033 1992
rect 7061 1970 7067 2018
rect 7070 2012 7089 2018
rect 7104 2012 7134 2020
rect 7070 2004 7134 2012
rect 7070 1988 7150 2004
rect 7166 1997 7228 2028
rect 7244 1997 7306 2028
rect 7375 2026 7424 2051
rect 7439 2026 7469 2042
rect 7338 2012 7368 2020
rect 7375 2018 7485 2026
rect 7338 2004 7383 2012
rect 7070 1986 7089 1988
rect 7104 1986 7150 1988
rect 7070 1970 7150 1986
rect 7177 1984 7212 1997
rect 7253 1994 7290 1997
rect 7253 1992 7295 1994
rect 7182 1981 7212 1984
rect 7191 1977 7198 1981
rect 7198 1976 7199 1977
rect 7157 1970 7167 1976
rect 6916 1962 6951 1970
rect 6916 1936 6917 1962
rect 6924 1936 6951 1962
rect 6859 1918 6889 1932
rect 6916 1928 6951 1936
rect 6953 1962 6994 1970
rect 6953 1936 6968 1962
rect 6975 1936 6994 1962
rect 7058 1958 7089 1970
rect 7104 1958 7207 1970
rect 7219 1960 7245 1986
rect 7260 1981 7290 1992
rect 7322 1988 7384 2004
rect 7322 1986 7368 1988
rect 7322 1970 7384 1986
rect 7396 1970 7402 2018
rect 7405 2010 7485 2018
rect 7405 2008 7424 2010
rect 7439 2008 7473 2010
rect 7405 1992 7485 2008
rect 7405 1970 7424 1992
rect 7439 1976 7469 1992
rect 7497 1986 7503 2060
rect 7506 1986 7525 2130
rect 7540 1986 7546 2130
rect 7555 2060 7568 2130
rect 7620 2126 7642 2130
rect 7613 2104 7642 2118
rect 7695 2104 7711 2118
rect 7749 2114 7755 2116
rect 7762 2114 7870 2130
rect 7877 2114 7883 2116
rect 7891 2114 7906 2130
rect 7972 2124 7991 2127
rect 7613 2102 7711 2104
rect 7738 2102 7906 2114
rect 7921 2104 7937 2118
rect 7972 2105 7994 2124
rect 8004 2118 8020 2119
rect 8003 2116 8020 2118
rect 8004 2111 8020 2116
rect 7994 2104 8000 2105
rect 8003 2104 8032 2111
rect 7921 2103 8032 2104
rect 7921 2102 8038 2103
rect 7597 2094 7648 2102
rect 7695 2094 7729 2102
rect 7597 2082 7622 2094
rect 7629 2082 7648 2094
rect 7702 2092 7729 2094
rect 7738 2092 7959 2102
rect 7994 2099 8000 2102
rect 7702 2088 7959 2092
rect 7597 2074 7648 2082
rect 7695 2074 7959 2088
rect 8003 2094 8038 2102
rect 7549 2026 7568 2060
rect 7613 2066 7642 2074
rect 7613 2060 7630 2066
rect 7613 2058 7647 2060
rect 7695 2058 7711 2074
rect 7712 2064 7920 2074
rect 7921 2064 7937 2074
rect 7985 2070 8000 2085
rect 8003 2082 8004 2094
rect 8011 2082 8038 2094
rect 8003 2074 8038 2082
rect 8003 2073 8032 2074
rect 7723 2060 7937 2064
rect 7738 2058 7937 2060
rect 7972 2060 7985 2070
rect 8003 2060 8020 2073
rect 7972 2058 8020 2060
rect 7614 2054 7647 2058
rect 7610 2052 7647 2054
rect 7610 2051 7677 2052
rect 7610 2046 7641 2051
rect 7647 2046 7677 2051
rect 7610 2042 7677 2046
rect 7583 2039 7677 2042
rect 7583 2032 7632 2039
rect 7583 2026 7613 2032
rect 7632 2027 7637 2032
rect 7549 2010 7629 2026
rect 7641 2018 7677 2039
rect 7738 2034 7927 2058
rect 7972 2057 8019 2058
rect 7985 2052 8019 2057
rect 7753 2031 7927 2034
rect 7746 2028 7927 2031
rect 7955 2051 8019 2052
rect 7549 2008 7568 2010
rect 7583 2008 7617 2010
rect 7549 1992 7629 2008
rect 7549 1986 7568 1992
rect 7265 1960 7368 1970
rect 7219 1958 7368 1960
rect 7389 1958 7424 1970
rect 7058 1956 7220 1958
rect 7070 1936 7089 1956
rect 7104 1954 7134 1956
rect 6953 1928 6994 1936
rect 7076 1932 7089 1936
rect 7141 1940 7220 1956
rect 7252 1956 7424 1958
rect 7252 1940 7331 1956
rect 7338 1954 7368 1956
rect 6916 1918 6945 1928
rect 6959 1918 6988 1928
rect 7003 1918 7033 1932
rect 7076 1918 7119 1932
rect 7141 1928 7331 1940
rect 7396 1936 7402 1956
rect 7126 1918 7156 1928
rect 7157 1918 7315 1928
rect 7319 1918 7349 1928
rect 7353 1918 7383 1932
rect 7411 1918 7424 1956
rect 7496 1970 7525 1986
rect 7539 1970 7568 1986
rect 7583 1976 7613 1992
rect 7641 1970 7647 2018
rect 7650 2012 7669 2018
rect 7684 2012 7714 2020
rect 7650 2004 7714 2012
rect 7650 1988 7730 2004
rect 7746 1997 7808 2028
rect 7824 1997 7886 2028
rect 7955 2026 8004 2051
rect 8019 2026 8049 2042
rect 7918 2012 7948 2020
rect 7955 2018 8065 2026
rect 7918 2004 7963 2012
rect 7650 1986 7669 1988
rect 7684 1986 7730 1988
rect 7650 1970 7730 1986
rect 7757 1984 7792 1997
rect 7833 1994 7870 1997
rect 7833 1992 7875 1994
rect 7762 1981 7792 1984
rect 7771 1977 7778 1981
rect 7778 1976 7779 1977
rect 7737 1970 7747 1976
rect 7496 1962 7531 1970
rect 7496 1936 7497 1962
rect 7504 1936 7531 1962
rect 7439 1918 7469 1932
rect 7496 1928 7531 1936
rect 7533 1962 7574 1970
rect 7533 1936 7548 1962
rect 7555 1936 7574 1962
rect 7638 1958 7669 1970
rect 7684 1958 7787 1970
rect 7799 1960 7825 1986
rect 7840 1981 7870 1992
rect 7902 1988 7964 2004
rect 7902 1986 7948 1988
rect 7902 1970 7964 1986
rect 7976 1970 7982 2018
rect 7985 2010 8065 2018
rect 7985 2008 8004 2010
rect 8019 2008 8053 2010
rect 7985 1992 8065 2008
rect 7985 1970 8004 1992
rect 8019 1976 8049 1992
rect 8077 1986 8083 2060
rect 8086 1986 8105 2130
rect 8120 1986 8126 2130
rect 8135 2060 8148 2130
rect 8200 2126 8222 2130
rect 8193 2104 8222 2118
rect 8275 2104 8291 2118
rect 8329 2114 8335 2116
rect 8342 2114 8450 2130
rect 8457 2114 8463 2116
rect 8471 2114 8486 2130
rect 8552 2124 8571 2127
rect 8193 2102 8291 2104
rect 8318 2102 8486 2114
rect 8501 2104 8517 2118
rect 8552 2105 8574 2124
rect 8584 2118 8600 2119
rect 8583 2116 8600 2118
rect 8584 2111 8600 2116
rect 8574 2104 8580 2105
rect 8583 2104 8612 2111
rect 8501 2103 8612 2104
rect 8501 2102 8618 2103
rect 8177 2094 8228 2102
rect 8275 2094 8309 2102
rect 8177 2082 8202 2094
rect 8209 2082 8228 2094
rect 8282 2092 8309 2094
rect 8318 2092 8539 2102
rect 8574 2099 8580 2102
rect 8282 2088 8539 2092
rect 8177 2074 8228 2082
rect 8275 2074 8539 2088
rect 8583 2094 8618 2102
rect 8129 2026 8148 2060
rect 8193 2066 8222 2074
rect 8193 2060 8210 2066
rect 8193 2058 8227 2060
rect 8275 2058 8291 2074
rect 8292 2064 8500 2074
rect 8501 2064 8517 2074
rect 8565 2070 8580 2085
rect 8583 2082 8584 2094
rect 8591 2082 8618 2094
rect 8583 2074 8618 2082
rect 8583 2073 8612 2074
rect 8303 2060 8517 2064
rect 8318 2058 8517 2060
rect 8552 2060 8565 2070
rect 8583 2060 8600 2073
rect 8552 2058 8600 2060
rect 8194 2054 8227 2058
rect 8190 2052 8227 2054
rect 8190 2051 8257 2052
rect 8190 2046 8221 2051
rect 8227 2046 8257 2051
rect 8190 2042 8257 2046
rect 8163 2039 8257 2042
rect 8163 2032 8212 2039
rect 8163 2026 8193 2032
rect 8212 2027 8217 2032
rect 8129 2010 8209 2026
rect 8221 2018 8257 2039
rect 8318 2034 8507 2058
rect 8552 2057 8599 2058
rect 8565 2052 8599 2057
rect 8333 2031 8507 2034
rect 8326 2028 8507 2031
rect 8535 2051 8599 2052
rect 8129 2008 8148 2010
rect 8163 2008 8197 2010
rect 8129 1992 8209 2008
rect 8129 1986 8148 1992
rect 7845 1960 7948 1970
rect 7799 1958 7948 1960
rect 7969 1958 8004 1970
rect 7638 1956 7800 1958
rect 7650 1936 7669 1956
rect 7684 1954 7714 1956
rect 7533 1928 7574 1936
rect 7656 1932 7669 1936
rect 7721 1940 7800 1956
rect 7832 1956 8004 1958
rect 7832 1940 7911 1956
rect 7918 1954 7948 1956
rect 7496 1918 7525 1928
rect 7539 1918 7568 1928
rect 7583 1918 7613 1932
rect 7656 1918 7699 1932
rect 7721 1928 7911 1940
rect 7976 1936 7982 1956
rect 7706 1918 7736 1928
rect 7737 1918 7895 1928
rect 7899 1918 7929 1928
rect 7933 1918 7963 1932
rect 7991 1918 8004 1956
rect 8076 1970 8105 1986
rect 8119 1970 8148 1986
rect 8163 1976 8193 1992
rect 8221 1970 8227 2018
rect 8230 2012 8249 2018
rect 8264 2012 8294 2020
rect 8230 2004 8294 2012
rect 8230 1988 8310 2004
rect 8326 1997 8388 2028
rect 8404 1997 8466 2028
rect 8535 2026 8584 2051
rect 8599 2026 8629 2042
rect 8498 2012 8528 2020
rect 8535 2018 8645 2026
rect 8498 2004 8543 2012
rect 8230 1986 8249 1988
rect 8264 1986 8310 1988
rect 8230 1970 8310 1986
rect 8337 1984 8372 1997
rect 8413 1994 8450 1997
rect 8413 1992 8455 1994
rect 8342 1981 8372 1984
rect 8351 1977 8358 1981
rect 8358 1976 8359 1977
rect 8317 1970 8327 1976
rect 8076 1962 8111 1970
rect 8076 1936 8077 1962
rect 8084 1936 8111 1962
rect 8019 1918 8049 1932
rect 8076 1928 8111 1936
rect 8113 1962 8154 1970
rect 8113 1936 8128 1962
rect 8135 1936 8154 1962
rect 8218 1958 8249 1970
rect 8264 1958 8367 1970
rect 8379 1960 8405 1986
rect 8420 1981 8450 1992
rect 8482 1988 8544 2004
rect 8482 1986 8528 1988
rect 8482 1970 8544 1986
rect 8556 1970 8562 2018
rect 8565 2010 8645 2018
rect 8565 2008 8584 2010
rect 8599 2008 8633 2010
rect 8565 1992 8645 2008
rect 8565 1970 8584 1992
rect 8599 1976 8629 1992
rect 8657 1986 8663 2060
rect 8666 1986 8685 2130
rect 8700 1986 8706 2130
rect 8715 2060 8728 2130
rect 8780 2126 8802 2130
rect 8773 2104 8802 2118
rect 8855 2104 8871 2118
rect 8909 2114 8915 2116
rect 8922 2114 9030 2130
rect 9037 2114 9043 2116
rect 9051 2114 9066 2130
rect 9132 2124 9151 2127
rect 8773 2102 8871 2104
rect 8898 2102 9066 2114
rect 9081 2104 9097 2118
rect 9132 2105 9154 2124
rect 9164 2118 9180 2119
rect 9163 2116 9180 2118
rect 9164 2111 9180 2116
rect 9154 2104 9160 2105
rect 9163 2104 9192 2111
rect 9081 2103 9192 2104
rect 9081 2102 9198 2103
rect 8757 2094 8808 2102
rect 8855 2094 8889 2102
rect 8757 2082 8782 2094
rect 8789 2082 8808 2094
rect 8862 2092 8889 2094
rect 8898 2092 9119 2102
rect 9154 2099 9160 2102
rect 8862 2088 9119 2092
rect 8757 2074 8808 2082
rect 8855 2074 9119 2088
rect 9163 2094 9198 2102
rect 8709 2026 8728 2060
rect 8773 2066 8802 2074
rect 8773 2060 8790 2066
rect 8773 2058 8807 2060
rect 8855 2058 8871 2074
rect 8872 2064 9080 2074
rect 9081 2064 9097 2074
rect 9145 2070 9160 2085
rect 9163 2082 9164 2094
rect 9171 2082 9198 2094
rect 9163 2074 9198 2082
rect 9163 2073 9192 2074
rect 8883 2060 9097 2064
rect 8898 2058 9097 2060
rect 9132 2060 9145 2070
rect 9163 2060 9180 2073
rect 9132 2058 9180 2060
rect 8774 2054 8807 2058
rect 8770 2052 8807 2054
rect 8770 2051 8837 2052
rect 8770 2046 8801 2051
rect 8807 2046 8837 2051
rect 8770 2042 8837 2046
rect 8743 2039 8837 2042
rect 8743 2032 8792 2039
rect 8743 2026 8773 2032
rect 8792 2027 8797 2032
rect 8709 2010 8789 2026
rect 8801 2018 8837 2039
rect 8898 2034 9087 2058
rect 9132 2057 9179 2058
rect 9145 2052 9179 2057
rect 8913 2031 9087 2034
rect 8906 2028 9087 2031
rect 9115 2051 9179 2052
rect 8709 2008 8728 2010
rect 8743 2008 8777 2010
rect 8709 1992 8789 2008
rect 8709 1986 8728 1992
rect 8425 1960 8528 1970
rect 8379 1958 8528 1960
rect 8549 1958 8584 1970
rect 8218 1956 8380 1958
rect 8230 1936 8249 1956
rect 8264 1954 8294 1956
rect 8113 1928 8154 1936
rect 8236 1932 8249 1936
rect 8301 1940 8380 1956
rect 8412 1956 8584 1958
rect 8412 1940 8491 1956
rect 8498 1954 8528 1956
rect 8076 1918 8105 1928
rect 8119 1918 8148 1928
rect 8163 1918 8193 1932
rect 8236 1918 8279 1932
rect 8301 1928 8491 1940
rect 8556 1936 8562 1956
rect 8286 1918 8316 1928
rect 8317 1918 8475 1928
rect 8479 1918 8509 1928
rect 8513 1918 8543 1932
rect 8571 1918 8584 1956
rect 8656 1970 8685 1986
rect 8699 1970 8728 1986
rect 8743 1976 8773 1992
rect 8801 1970 8807 2018
rect 8810 2012 8829 2018
rect 8844 2012 8874 2020
rect 8810 2004 8874 2012
rect 8810 1988 8890 2004
rect 8906 1997 8968 2028
rect 8984 1997 9046 2028
rect 9115 2026 9164 2051
rect 9179 2026 9209 2042
rect 9078 2012 9108 2020
rect 9115 2018 9225 2026
rect 9078 2004 9123 2012
rect 8810 1986 8829 1988
rect 8844 1986 8890 1988
rect 8810 1970 8890 1986
rect 8917 1984 8952 1997
rect 8993 1994 9030 1997
rect 8993 1992 9035 1994
rect 8922 1981 8952 1984
rect 8931 1977 8938 1981
rect 8938 1976 8939 1977
rect 8897 1970 8907 1976
rect 8656 1962 8691 1970
rect 8656 1936 8657 1962
rect 8664 1936 8691 1962
rect 8599 1918 8629 1932
rect 8656 1928 8691 1936
rect 8693 1962 8734 1970
rect 8693 1936 8708 1962
rect 8715 1936 8734 1962
rect 8798 1958 8829 1970
rect 8844 1958 8947 1970
rect 8959 1960 8985 1986
rect 9000 1981 9030 1992
rect 9062 1988 9124 2004
rect 9062 1986 9108 1988
rect 9062 1970 9124 1986
rect 9136 1970 9142 2018
rect 9145 2010 9225 2018
rect 9145 2008 9164 2010
rect 9179 2008 9213 2010
rect 9145 1992 9225 2008
rect 9145 1970 9164 1992
rect 9179 1976 9209 1992
rect 9237 1986 9243 2060
rect 9252 1986 9265 2130
rect 9005 1960 9108 1970
rect 8959 1958 9108 1960
rect 9129 1958 9164 1970
rect 8798 1956 8960 1958
rect 8810 1936 8829 1956
rect 8844 1954 8874 1956
rect 8693 1928 8734 1936
rect 8816 1932 8829 1936
rect 8881 1940 8960 1956
rect 8992 1956 9164 1958
rect 8992 1940 9071 1956
rect 9078 1954 9108 1956
rect 8656 1918 8685 1928
rect 8699 1918 8728 1928
rect 8743 1918 8773 1932
rect 8816 1918 8859 1932
rect 8881 1928 9071 1940
rect 9136 1936 9142 1956
rect 8866 1918 8896 1928
rect 8897 1918 9055 1928
rect 9059 1918 9089 1928
rect 9093 1918 9123 1932
rect 9151 1918 9164 1956
rect 9236 1970 9265 1986
rect 9236 1962 9271 1970
rect 9236 1936 9237 1962
rect 9244 1936 9271 1962
rect 9179 1918 9209 1932
rect 9236 1928 9271 1936
rect 9236 1918 9265 1928
rect -1 1912 9265 1918
rect 0 1904 9265 1912
rect 15 1874 28 1904
rect 43 1890 73 1904
rect 116 1890 159 1904
rect 166 1890 386 1904
rect 393 1890 423 1904
rect 83 1876 98 1888
rect 117 1876 130 1890
rect 198 1886 351 1890
rect 80 1874 102 1876
rect 180 1874 372 1886
rect 451 1874 464 1904
rect 479 1890 509 1904
rect 546 1874 565 1904
rect 580 1874 586 1904
rect 595 1874 608 1904
rect 623 1890 653 1904
rect 696 1890 739 1904
rect 746 1890 966 1904
rect 973 1890 1003 1904
rect 663 1876 678 1888
rect 697 1876 710 1890
rect 778 1886 931 1890
rect 660 1874 682 1876
rect 760 1874 952 1886
rect 1031 1874 1044 1904
rect 1059 1890 1089 1904
rect 1126 1874 1145 1904
rect 1160 1874 1166 1904
rect 1175 1874 1188 1904
rect 1203 1890 1233 1904
rect 1276 1890 1319 1904
rect 1326 1890 1546 1904
rect 1553 1890 1583 1904
rect 1243 1876 1258 1888
rect 1277 1876 1290 1890
rect 1358 1886 1511 1890
rect 1240 1874 1262 1876
rect 1340 1874 1532 1886
rect 1611 1874 1624 1904
rect 1639 1890 1669 1904
rect 1706 1874 1725 1904
rect 1740 1874 1746 1904
rect 1755 1874 1768 1904
rect 1783 1890 1813 1904
rect 1856 1890 1899 1904
rect 1906 1890 2126 1904
rect 2133 1890 2163 1904
rect 1823 1876 1838 1888
rect 1857 1876 1870 1890
rect 1938 1886 2091 1890
rect 1820 1874 1842 1876
rect 1920 1874 2112 1886
rect 2191 1874 2204 1904
rect 2219 1890 2249 1904
rect 2286 1874 2305 1904
rect 2320 1874 2326 1904
rect 2335 1874 2348 1904
rect 2363 1890 2393 1904
rect 2436 1890 2479 1904
rect 2486 1890 2706 1904
rect 2713 1890 2743 1904
rect 2403 1876 2418 1888
rect 2437 1876 2450 1890
rect 2518 1886 2671 1890
rect 2400 1874 2422 1876
rect 2500 1874 2692 1886
rect 2771 1874 2784 1904
rect 2799 1890 2829 1904
rect 2866 1874 2885 1904
rect 2900 1874 2906 1904
rect 2915 1874 2928 1904
rect 2943 1890 2973 1904
rect 3016 1890 3059 1904
rect 3066 1890 3286 1904
rect 3293 1890 3323 1904
rect 2983 1876 2998 1888
rect 3017 1876 3030 1890
rect 3098 1886 3251 1890
rect 2980 1874 3002 1876
rect 3080 1874 3272 1886
rect 3351 1874 3364 1904
rect 3379 1890 3409 1904
rect 3446 1874 3465 1904
rect 3480 1874 3486 1904
rect 3495 1874 3508 1904
rect 3523 1890 3553 1904
rect 3596 1890 3639 1904
rect 3646 1890 3866 1904
rect 3873 1890 3903 1904
rect 3563 1876 3578 1888
rect 3597 1876 3610 1890
rect 3678 1886 3831 1890
rect 3560 1874 3582 1876
rect 3660 1874 3852 1886
rect 3931 1874 3944 1904
rect 3959 1890 3989 1904
rect 4026 1874 4045 1904
rect 4060 1874 4066 1904
rect 4075 1874 4088 1904
rect 4103 1890 4133 1904
rect 4176 1890 4219 1904
rect 4226 1890 4446 1904
rect 4453 1890 4483 1904
rect 4143 1876 4158 1888
rect 4177 1876 4190 1890
rect 4258 1886 4411 1890
rect 4140 1874 4162 1876
rect 4240 1874 4432 1886
rect 4511 1874 4524 1904
rect 4539 1890 4569 1904
rect 4606 1874 4625 1904
rect 4640 1874 4646 1904
rect 4655 1874 4668 1904
rect 4683 1890 4713 1904
rect 4756 1890 4799 1904
rect 4806 1890 5026 1904
rect 5033 1890 5063 1904
rect 4723 1876 4738 1888
rect 4757 1876 4770 1890
rect 4838 1886 4991 1890
rect 4720 1874 4742 1876
rect 4820 1874 5012 1886
rect 5091 1874 5104 1904
rect 5119 1890 5149 1904
rect 5186 1874 5205 1904
rect 5220 1874 5226 1904
rect 5235 1874 5248 1904
rect 5263 1890 5293 1904
rect 5336 1890 5379 1904
rect 5386 1890 5606 1904
rect 5613 1890 5643 1904
rect 5303 1876 5318 1888
rect 5337 1876 5350 1890
rect 5418 1886 5571 1890
rect 5300 1874 5322 1876
rect 5400 1874 5592 1886
rect 5671 1874 5684 1904
rect 5699 1890 5729 1904
rect 5766 1874 5785 1904
rect 5800 1874 5806 1904
rect 5815 1874 5828 1904
rect 5843 1890 5873 1904
rect 5916 1890 5959 1904
rect 5966 1890 6186 1904
rect 6193 1890 6223 1904
rect 5883 1876 5898 1888
rect 5917 1876 5930 1890
rect 5998 1886 6151 1890
rect 5880 1874 5902 1876
rect 5980 1874 6172 1886
rect 6251 1874 6264 1904
rect 6279 1890 6309 1904
rect 6346 1874 6365 1904
rect 6380 1874 6386 1904
rect 6395 1874 6408 1904
rect 6423 1890 6453 1904
rect 6496 1890 6539 1904
rect 6546 1890 6766 1904
rect 6773 1890 6803 1904
rect 6463 1876 6478 1888
rect 6497 1876 6510 1890
rect 6578 1886 6731 1890
rect 6460 1874 6482 1876
rect 6560 1874 6752 1886
rect 6831 1874 6844 1904
rect 6859 1890 6889 1904
rect 6926 1874 6945 1904
rect 6960 1874 6966 1904
rect 6975 1874 6988 1904
rect 7003 1890 7033 1904
rect 7076 1890 7119 1904
rect 7126 1890 7346 1904
rect 7353 1890 7383 1904
rect 7043 1876 7058 1888
rect 7077 1876 7090 1890
rect 7158 1886 7311 1890
rect 7040 1874 7062 1876
rect 7140 1874 7332 1886
rect 7411 1874 7424 1904
rect 7439 1890 7469 1904
rect 7506 1874 7525 1904
rect 7540 1874 7546 1904
rect 7555 1874 7568 1904
rect 7583 1890 7613 1904
rect 7656 1890 7699 1904
rect 7706 1890 7926 1904
rect 7933 1890 7963 1904
rect 7623 1876 7638 1888
rect 7657 1876 7670 1890
rect 7738 1886 7891 1890
rect 7620 1874 7642 1876
rect 7720 1874 7912 1886
rect 7991 1874 8004 1904
rect 8019 1890 8049 1904
rect 8086 1874 8105 1904
rect 8120 1874 8126 1904
rect 8135 1874 8148 1904
rect 8163 1890 8193 1904
rect 8236 1890 8279 1904
rect 8286 1890 8506 1904
rect 8513 1890 8543 1904
rect 8203 1876 8218 1888
rect 8237 1876 8250 1890
rect 8318 1886 8471 1890
rect 8200 1874 8222 1876
rect 8300 1874 8492 1886
rect 8571 1874 8584 1904
rect 8599 1890 8629 1904
rect 8666 1874 8685 1904
rect 8700 1874 8706 1904
rect 8715 1874 8728 1904
rect 8743 1890 8773 1904
rect 8816 1890 8859 1904
rect 8866 1890 9086 1904
rect 9093 1890 9123 1904
rect 8783 1876 8798 1888
rect 8817 1876 8830 1890
rect 8898 1886 9051 1890
rect 8780 1874 8802 1876
rect 8880 1874 9072 1886
rect 9151 1874 9164 1904
rect 9179 1890 9209 1904
rect 9252 1874 9265 1904
rect 0 1860 9265 1874
rect 15 1790 28 1860
rect 80 1856 102 1860
rect 73 1834 102 1848
rect 155 1834 171 1848
rect 209 1844 215 1846
rect 222 1844 330 1860
rect 337 1844 343 1846
rect 351 1844 366 1860
rect 432 1854 451 1857
rect 73 1832 171 1834
rect 198 1832 366 1844
rect 381 1834 397 1848
rect 432 1835 454 1854
rect 464 1848 480 1849
rect 463 1846 480 1848
rect 464 1841 480 1846
rect 454 1834 460 1835
rect 463 1834 492 1841
rect 381 1833 492 1834
rect 381 1832 498 1833
rect 57 1824 108 1832
rect 155 1824 189 1832
rect 57 1812 82 1824
rect 89 1812 108 1824
rect 162 1822 189 1824
rect 198 1822 419 1832
rect 454 1829 460 1832
rect 162 1818 419 1822
rect 57 1804 108 1812
rect 155 1804 419 1818
rect 463 1824 498 1832
rect 9 1756 28 1790
rect 73 1796 102 1804
rect 73 1790 90 1796
rect 73 1788 107 1790
rect 155 1788 171 1804
rect 172 1794 380 1804
rect 381 1794 397 1804
rect 445 1800 460 1815
rect 463 1812 464 1824
rect 471 1812 498 1824
rect 463 1804 498 1812
rect 463 1803 492 1804
rect 183 1790 397 1794
rect 198 1788 397 1790
rect 432 1790 445 1800
rect 463 1790 480 1803
rect 432 1788 480 1790
rect 74 1784 107 1788
rect 70 1782 107 1784
rect 70 1781 137 1782
rect 70 1776 101 1781
rect 107 1776 137 1781
rect 70 1772 137 1776
rect 43 1769 137 1772
rect 43 1762 92 1769
rect 43 1756 73 1762
rect 92 1757 97 1762
rect 9 1740 89 1756
rect 101 1748 137 1769
rect 198 1764 387 1788
rect 432 1787 479 1788
rect 445 1782 479 1787
rect 213 1761 387 1764
rect 206 1758 387 1761
rect 415 1781 479 1782
rect 9 1738 28 1740
rect 43 1738 77 1740
rect 9 1722 89 1738
rect 9 1716 28 1722
rect -1 1700 28 1716
rect 43 1706 73 1722
rect 101 1700 107 1748
rect 110 1742 129 1748
rect 144 1742 174 1750
rect 110 1734 174 1742
rect 110 1718 190 1734
rect 206 1727 268 1758
rect 284 1727 346 1758
rect 415 1756 464 1781
rect 479 1756 509 1772
rect 378 1742 408 1750
rect 415 1748 525 1756
rect 378 1734 423 1742
rect 110 1716 129 1718
rect 144 1716 190 1718
rect 110 1700 190 1716
rect 217 1714 252 1727
rect 293 1724 330 1727
rect 293 1722 335 1724
rect 222 1711 252 1714
rect 231 1707 238 1711
rect 238 1706 239 1707
rect 197 1700 207 1706
rect -7 1692 34 1700
rect -7 1666 8 1692
rect 15 1666 34 1692
rect 98 1688 129 1700
rect 144 1688 247 1700
rect 259 1690 285 1716
rect 300 1711 330 1722
rect 362 1718 424 1734
rect 362 1716 408 1718
rect 362 1700 424 1716
rect 436 1700 442 1748
rect 445 1740 525 1748
rect 445 1738 464 1740
rect 479 1738 513 1740
rect 445 1722 525 1738
rect 445 1700 464 1722
rect 479 1706 509 1722
rect 537 1716 543 1790
rect 546 1716 565 1860
rect 580 1716 586 1860
rect 595 1790 608 1860
rect 660 1856 682 1860
rect 653 1834 682 1848
rect 735 1834 751 1848
rect 789 1844 795 1846
rect 802 1844 910 1860
rect 917 1844 923 1846
rect 931 1844 946 1860
rect 1012 1854 1031 1857
rect 653 1832 751 1834
rect 778 1832 946 1844
rect 961 1834 977 1848
rect 1012 1835 1034 1854
rect 1044 1848 1060 1849
rect 1043 1846 1060 1848
rect 1044 1841 1060 1846
rect 1034 1834 1040 1835
rect 1043 1834 1072 1841
rect 961 1833 1072 1834
rect 961 1832 1078 1833
rect 637 1824 688 1832
rect 735 1824 769 1832
rect 637 1812 662 1824
rect 669 1812 688 1824
rect 742 1822 769 1824
rect 778 1822 999 1832
rect 1034 1829 1040 1832
rect 742 1818 999 1822
rect 637 1804 688 1812
rect 735 1804 999 1818
rect 1043 1824 1078 1832
rect 589 1756 608 1790
rect 653 1796 682 1804
rect 653 1790 670 1796
rect 653 1788 687 1790
rect 735 1788 751 1804
rect 752 1794 960 1804
rect 961 1794 977 1804
rect 1025 1800 1040 1815
rect 1043 1812 1044 1824
rect 1051 1812 1078 1824
rect 1043 1804 1078 1812
rect 1043 1803 1072 1804
rect 763 1790 977 1794
rect 778 1788 977 1790
rect 1012 1790 1025 1800
rect 1043 1790 1060 1803
rect 1012 1788 1060 1790
rect 654 1784 687 1788
rect 650 1782 687 1784
rect 650 1781 717 1782
rect 650 1776 681 1781
rect 687 1776 717 1781
rect 650 1772 717 1776
rect 623 1769 717 1772
rect 623 1762 672 1769
rect 623 1756 653 1762
rect 672 1757 677 1762
rect 589 1740 669 1756
rect 681 1748 717 1769
rect 778 1764 967 1788
rect 1012 1787 1059 1788
rect 1025 1782 1059 1787
rect 793 1761 967 1764
rect 786 1758 967 1761
rect 995 1781 1059 1782
rect 589 1738 608 1740
rect 623 1738 657 1740
rect 589 1722 669 1738
rect 589 1716 608 1722
rect 305 1690 408 1700
rect 259 1688 408 1690
rect 429 1688 464 1700
rect 98 1686 260 1688
rect 110 1666 129 1686
rect 144 1684 174 1686
rect -7 1658 34 1666
rect 116 1662 129 1666
rect 181 1670 260 1686
rect 292 1686 464 1688
rect 292 1670 371 1686
rect 378 1684 408 1686
rect -1 1648 28 1658
rect 43 1648 73 1662
rect 116 1648 159 1662
rect 181 1658 371 1670
rect 436 1666 442 1686
rect 166 1648 196 1658
rect 197 1648 355 1658
rect 359 1648 389 1658
rect 393 1648 423 1662
rect 451 1648 464 1686
rect 536 1700 565 1716
rect 579 1700 608 1716
rect 623 1706 653 1722
rect 681 1700 687 1748
rect 690 1742 709 1748
rect 724 1742 754 1750
rect 690 1734 754 1742
rect 690 1718 770 1734
rect 786 1727 848 1758
rect 864 1727 926 1758
rect 995 1756 1044 1781
rect 1059 1756 1089 1772
rect 958 1742 988 1750
rect 995 1748 1105 1756
rect 958 1734 1003 1742
rect 690 1716 709 1718
rect 724 1716 770 1718
rect 690 1700 770 1716
rect 797 1714 832 1727
rect 873 1724 910 1727
rect 873 1722 915 1724
rect 802 1711 832 1714
rect 811 1707 818 1711
rect 818 1706 819 1707
rect 777 1700 787 1706
rect 536 1692 571 1700
rect 536 1666 537 1692
rect 544 1666 571 1692
rect 479 1648 509 1662
rect 536 1658 571 1666
rect 573 1692 614 1700
rect 573 1666 588 1692
rect 595 1666 614 1692
rect 678 1688 709 1700
rect 724 1688 827 1700
rect 839 1690 865 1716
rect 880 1711 910 1722
rect 942 1718 1004 1734
rect 942 1716 988 1718
rect 942 1700 1004 1716
rect 1016 1700 1022 1748
rect 1025 1740 1105 1748
rect 1025 1738 1044 1740
rect 1059 1738 1093 1740
rect 1025 1722 1105 1738
rect 1025 1700 1044 1722
rect 1059 1706 1089 1722
rect 1117 1716 1123 1790
rect 1126 1716 1145 1860
rect 1160 1716 1166 1860
rect 1175 1790 1188 1860
rect 1240 1856 1262 1860
rect 1233 1834 1262 1848
rect 1315 1834 1331 1848
rect 1369 1844 1375 1846
rect 1382 1844 1490 1860
rect 1497 1844 1503 1846
rect 1511 1844 1526 1860
rect 1592 1854 1611 1857
rect 1233 1832 1331 1834
rect 1358 1832 1526 1844
rect 1541 1834 1557 1848
rect 1592 1835 1614 1854
rect 1624 1848 1640 1849
rect 1623 1846 1640 1848
rect 1624 1841 1640 1846
rect 1614 1834 1620 1835
rect 1623 1834 1652 1841
rect 1541 1833 1652 1834
rect 1541 1832 1658 1833
rect 1217 1824 1268 1832
rect 1315 1824 1349 1832
rect 1217 1812 1242 1824
rect 1249 1812 1268 1824
rect 1322 1822 1349 1824
rect 1358 1822 1579 1832
rect 1614 1829 1620 1832
rect 1322 1818 1579 1822
rect 1217 1804 1268 1812
rect 1315 1804 1579 1818
rect 1623 1824 1658 1832
rect 1169 1756 1188 1790
rect 1233 1796 1262 1804
rect 1233 1790 1250 1796
rect 1233 1788 1267 1790
rect 1315 1788 1331 1804
rect 1332 1794 1540 1804
rect 1541 1794 1557 1804
rect 1605 1800 1620 1815
rect 1623 1812 1624 1824
rect 1631 1812 1658 1824
rect 1623 1804 1658 1812
rect 1623 1803 1652 1804
rect 1343 1790 1557 1794
rect 1358 1788 1557 1790
rect 1592 1790 1605 1800
rect 1623 1790 1640 1803
rect 1592 1788 1640 1790
rect 1234 1784 1267 1788
rect 1230 1782 1267 1784
rect 1230 1781 1297 1782
rect 1230 1776 1261 1781
rect 1267 1776 1297 1781
rect 1230 1772 1297 1776
rect 1203 1769 1297 1772
rect 1203 1762 1252 1769
rect 1203 1756 1233 1762
rect 1252 1757 1257 1762
rect 1169 1740 1249 1756
rect 1261 1748 1297 1769
rect 1358 1764 1547 1788
rect 1592 1787 1639 1788
rect 1605 1782 1639 1787
rect 1373 1761 1547 1764
rect 1366 1758 1547 1761
rect 1575 1781 1639 1782
rect 1169 1738 1188 1740
rect 1203 1738 1237 1740
rect 1169 1722 1249 1738
rect 1169 1716 1188 1722
rect 885 1690 988 1700
rect 839 1688 988 1690
rect 1009 1688 1044 1700
rect 678 1686 840 1688
rect 690 1666 709 1686
rect 724 1684 754 1686
rect 573 1658 614 1666
rect 696 1662 709 1666
rect 761 1670 840 1686
rect 872 1686 1044 1688
rect 872 1670 951 1686
rect 958 1684 988 1686
rect 536 1648 565 1658
rect 579 1648 608 1658
rect 623 1648 653 1662
rect 696 1648 739 1662
rect 761 1658 951 1670
rect 1016 1666 1022 1686
rect 746 1648 776 1658
rect 777 1648 935 1658
rect 939 1648 969 1658
rect 973 1648 1003 1662
rect 1031 1648 1044 1686
rect 1116 1700 1145 1716
rect 1159 1700 1188 1716
rect 1203 1706 1233 1722
rect 1261 1700 1267 1748
rect 1270 1742 1289 1748
rect 1304 1742 1334 1750
rect 1270 1734 1334 1742
rect 1270 1718 1350 1734
rect 1366 1727 1428 1758
rect 1444 1727 1506 1758
rect 1575 1756 1624 1781
rect 1639 1756 1669 1772
rect 1538 1742 1568 1750
rect 1575 1748 1685 1756
rect 1538 1734 1583 1742
rect 1270 1716 1289 1718
rect 1304 1716 1350 1718
rect 1270 1700 1350 1716
rect 1377 1714 1412 1727
rect 1453 1724 1490 1727
rect 1453 1722 1495 1724
rect 1382 1711 1412 1714
rect 1391 1707 1398 1711
rect 1398 1706 1399 1707
rect 1357 1700 1367 1706
rect 1116 1692 1151 1700
rect 1116 1666 1117 1692
rect 1124 1666 1151 1692
rect 1059 1648 1089 1662
rect 1116 1658 1151 1666
rect 1153 1692 1194 1700
rect 1153 1666 1168 1692
rect 1175 1666 1194 1692
rect 1258 1688 1289 1700
rect 1304 1688 1407 1700
rect 1419 1690 1445 1716
rect 1460 1711 1490 1722
rect 1522 1718 1584 1734
rect 1522 1716 1568 1718
rect 1522 1700 1584 1716
rect 1596 1700 1602 1748
rect 1605 1740 1685 1748
rect 1605 1738 1624 1740
rect 1639 1738 1673 1740
rect 1605 1722 1685 1738
rect 1605 1700 1624 1722
rect 1639 1706 1669 1722
rect 1697 1716 1703 1790
rect 1706 1716 1725 1860
rect 1740 1716 1746 1860
rect 1755 1790 1768 1860
rect 1820 1856 1842 1860
rect 1813 1834 1842 1848
rect 1895 1834 1911 1848
rect 1949 1844 1955 1846
rect 1962 1844 2070 1860
rect 2077 1844 2083 1846
rect 2091 1844 2106 1860
rect 2172 1854 2191 1857
rect 1813 1832 1911 1834
rect 1938 1832 2106 1844
rect 2121 1834 2137 1848
rect 2172 1835 2194 1854
rect 2204 1848 2220 1849
rect 2203 1846 2220 1848
rect 2204 1841 2220 1846
rect 2194 1834 2200 1835
rect 2203 1834 2232 1841
rect 2121 1833 2232 1834
rect 2121 1832 2238 1833
rect 1797 1824 1848 1832
rect 1895 1824 1929 1832
rect 1797 1812 1822 1824
rect 1829 1812 1848 1824
rect 1902 1822 1929 1824
rect 1938 1822 2159 1832
rect 2194 1829 2200 1832
rect 1902 1818 2159 1822
rect 1797 1804 1848 1812
rect 1895 1804 2159 1818
rect 2203 1824 2238 1832
rect 1749 1756 1768 1790
rect 1813 1796 1842 1804
rect 1813 1790 1830 1796
rect 1813 1788 1847 1790
rect 1895 1788 1911 1804
rect 1912 1794 2120 1804
rect 2121 1794 2137 1804
rect 2185 1800 2200 1815
rect 2203 1812 2204 1824
rect 2211 1812 2238 1824
rect 2203 1804 2238 1812
rect 2203 1803 2232 1804
rect 1923 1790 2137 1794
rect 1938 1788 2137 1790
rect 2172 1790 2185 1800
rect 2203 1790 2220 1803
rect 2172 1788 2220 1790
rect 1814 1784 1847 1788
rect 1810 1782 1847 1784
rect 1810 1781 1877 1782
rect 1810 1776 1841 1781
rect 1847 1776 1877 1781
rect 1810 1772 1877 1776
rect 1783 1769 1877 1772
rect 1783 1762 1832 1769
rect 1783 1756 1813 1762
rect 1832 1757 1837 1762
rect 1749 1740 1829 1756
rect 1841 1748 1877 1769
rect 1938 1764 2127 1788
rect 2172 1787 2219 1788
rect 2185 1782 2219 1787
rect 1953 1761 2127 1764
rect 1946 1758 2127 1761
rect 2155 1781 2219 1782
rect 1749 1738 1768 1740
rect 1783 1738 1817 1740
rect 1749 1722 1829 1738
rect 1749 1716 1768 1722
rect 1465 1690 1568 1700
rect 1419 1688 1568 1690
rect 1589 1688 1624 1700
rect 1258 1686 1420 1688
rect 1270 1666 1289 1686
rect 1304 1684 1334 1686
rect 1153 1658 1194 1666
rect 1276 1662 1289 1666
rect 1341 1670 1420 1686
rect 1452 1686 1624 1688
rect 1452 1670 1531 1686
rect 1538 1684 1568 1686
rect 1116 1648 1145 1658
rect 1159 1648 1188 1658
rect 1203 1648 1233 1662
rect 1276 1648 1319 1662
rect 1341 1658 1531 1670
rect 1596 1666 1602 1686
rect 1326 1648 1356 1658
rect 1357 1648 1515 1658
rect 1519 1648 1549 1658
rect 1553 1648 1583 1662
rect 1611 1648 1624 1686
rect 1696 1700 1725 1716
rect 1739 1700 1768 1716
rect 1783 1706 1813 1722
rect 1841 1700 1847 1748
rect 1850 1742 1869 1748
rect 1884 1742 1914 1750
rect 1850 1734 1914 1742
rect 1850 1718 1930 1734
rect 1946 1727 2008 1758
rect 2024 1727 2086 1758
rect 2155 1756 2204 1781
rect 2219 1756 2249 1772
rect 2118 1742 2148 1750
rect 2155 1748 2265 1756
rect 2118 1734 2163 1742
rect 1850 1716 1869 1718
rect 1884 1716 1930 1718
rect 1850 1700 1930 1716
rect 1957 1714 1992 1727
rect 2033 1724 2070 1727
rect 2033 1722 2075 1724
rect 1962 1711 1992 1714
rect 1971 1707 1978 1711
rect 1978 1706 1979 1707
rect 1937 1700 1947 1706
rect 1696 1692 1731 1700
rect 1696 1666 1697 1692
rect 1704 1666 1731 1692
rect 1639 1648 1669 1662
rect 1696 1658 1731 1666
rect 1733 1692 1774 1700
rect 1733 1666 1748 1692
rect 1755 1666 1774 1692
rect 1838 1688 1869 1700
rect 1884 1688 1987 1700
rect 1999 1690 2025 1716
rect 2040 1711 2070 1722
rect 2102 1718 2164 1734
rect 2102 1716 2148 1718
rect 2102 1700 2164 1716
rect 2176 1700 2182 1748
rect 2185 1740 2265 1748
rect 2185 1738 2204 1740
rect 2219 1738 2253 1740
rect 2185 1722 2265 1738
rect 2185 1700 2204 1722
rect 2219 1706 2249 1722
rect 2277 1716 2283 1790
rect 2286 1716 2305 1860
rect 2320 1716 2326 1860
rect 2335 1790 2348 1860
rect 2400 1856 2422 1860
rect 2393 1834 2422 1848
rect 2475 1834 2491 1848
rect 2529 1844 2535 1846
rect 2542 1844 2650 1860
rect 2657 1844 2663 1846
rect 2671 1844 2686 1860
rect 2752 1854 2771 1857
rect 2393 1832 2491 1834
rect 2518 1832 2686 1844
rect 2701 1834 2717 1848
rect 2752 1835 2774 1854
rect 2784 1848 2800 1849
rect 2783 1846 2800 1848
rect 2784 1841 2800 1846
rect 2774 1834 2780 1835
rect 2783 1834 2812 1841
rect 2701 1833 2812 1834
rect 2701 1832 2818 1833
rect 2377 1824 2428 1832
rect 2475 1824 2509 1832
rect 2377 1812 2402 1824
rect 2409 1812 2428 1824
rect 2482 1822 2509 1824
rect 2518 1822 2739 1832
rect 2774 1829 2780 1832
rect 2482 1818 2739 1822
rect 2377 1804 2428 1812
rect 2475 1804 2739 1818
rect 2783 1824 2818 1832
rect 2329 1756 2348 1790
rect 2393 1796 2422 1804
rect 2393 1790 2410 1796
rect 2393 1788 2427 1790
rect 2475 1788 2491 1804
rect 2492 1794 2700 1804
rect 2701 1794 2717 1804
rect 2765 1800 2780 1815
rect 2783 1812 2784 1824
rect 2791 1812 2818 1824
rect 2783 1804 2818 1812
rect 2783 1803 2812 1804
rect 2503 1790 2717 1794
rect 2518 1788 2717 1790
rect 2752 1790 2765 1800
rect 2783 1790 2800 1803
rect 2752 1788 2800 1790
rect 2394 1784 2427 1788
rect 2390 1782 2427 1784
rect 2390 1781 2457 1782
rect 2390 1776 2421 1781
rect 2427 1776 2457 1781
rect 2390 1772 2457 1776
rect 2363 1769 2457 1772
rect 2363 1762 2412 1769
rect 2363 1756 2393 1762
rect 2412 1757 2417 1762
rect 2329 1740 2409 1756
rect 2421 1748 2457 1769
rect 2518 1764 2707 1788
rect 2752 1787 2799 1788
rect 2765 1782 2799 1787
rect 2533 1761 2707 1764
rect 2526 1758 2707 1761
rect 2735 1781 2799 1782
rect 2329 1738 2348 1740
rect 2363 1738 2397 1740
rect 2329 1722 2409 1738
rect 2329 1716 2348 1722
rect 2045 1690 2148 1700
rect 1999 1688 2148 1690
rect 2169 1688 2204 1700
rect 1838 1686 2000 1688
rect 1850 1666 1869 1686
rect 1884 1684 1914 1686
rect 1733 1658 1774 1666
rect 1856 1662 1869 1666
rect 1921 1670 2000 1686
rect 2032 1686 2204 1688
rect 2032 1670 2111 1686
rect 2118 1684 2148 1686
rect 1696 1648 1725 1658
rect 1739 1648 1768 1658
rect 1783 1648 1813 1662
rect 1856 1648 1899 1662
rect 1921 1658 2111 1670
rect 2176 1666 2182 1686
rect 1906 1648 1936 1658
rect 1937 1648 2095 1658
rect 2099 1648 2129 1658
rect 2133 1648 2163 1662
rect 2191 1648 2204 1686
rect 2276 1700 2305 1716
rect 2319 1700 2348 1716
rect 2363 1706 2393 1722
rect 2421 1700 2427 1748
rect 2430 1742 2449 1748
rect 2464 1742 2494 1750
rect 2430 1734 2494 1742
rect 2430 1718 2510 1734
rect 2526 1727 2588 1758
rect 2604 1727 2666 1758
rect 2735 1756 2784 1781
rect 2799 1756 2829 1772
rect 2698 1742 2728 1750
rect 2735 1748 2845 1756
rect 2698 1734 2743 1742
rect 2430 1716 2449 1718
rect 2464 1716 2510 1718
rect 2430 1700 2510 1716
rect 2537 1714 2572 1727
rect 2613 1724 2650 1727
rect 2613 1722 2655 1724
rect 2542 1711 2572 1714
rect 2551 1707 2558 1711
rect 2558 1706 2559 1707
rect 2517 1700 2527 1706
rect 2276 1692 2311 1700
rect 2276 1666 2277 1692
rect 2284 1666 2311 1692
rect 2219 1648 2249 1662
rect 2276 1658 2311 1666
rect 2313 1692 2354 1700
rect 2313 1666 2328 1692
rect 2335 1666 2354 1692
rect 2418 1688 2449 1700
rect 2464 1688 2567 1700
rect 2579 1690 2605 1716
rect 2620 1711 2650 1722
rect 2682 1718 2744 1734
rect 2682 1716 2728 1718
rect 2682 1700 2744 1716
rect 2756 1700 2762 1748
rect 2765 1740 2845 1748
rect 2765 1738 2784 1740
rect 2799 1738 2833 1740
rect 2765 1722 2845 1738
rect 2765 1700 2784 1722
rect 2799 1706 2829 1722
rect 2857 1716 2863 1790
rect 2866 1716 2885 1860
rect 2900 1716 2906 1860
rect 2915 1790 2928 1860
rect 2980 1856 3002 1860
rect 2973 1834 3002 1848
rect 3055 1834 3071 1848
rect 3109 1844 3115 1846
rect 3122 1844 3230 1860
rect 3237 1844 3243 1846
rect 3251 1844 3266 1860
rect 3332 1854 3351 1857
rect 2973 1832 3071 1834
rect 3098 1832 3266 1844
rect 3281 1834 3297 1848
rect 3332 1835 3354 1854
rect 3364 1848 3380 1849
rect 3363 1846 3380 1848
rect 3364 1841 3380 1846
rect 3354 1834 3360 1835
rect 3363 1834 3392 1841
rect 3281 1833 3392 1834
rect 3281 1832 3398 1833
rect 2957 1824 3008 1832
rect 3055 1824 3089 1832
rect 2957 1812 2982 1824
rect 2989 1812 3008 1824
rect 3062 1822 3089 1824
rect 3098 1822 3319 1832
rect 3354 1829 3360 1832
rect 3062 1818 3319 1822
rect 2957 1804 3008 1812
rect 3055 1804 3319 1818
rect 3363 1824 3398 1832
rect 2909 1756 2928 1790
rect 2973 1796 3002 1804
rect 2973 1790 2990 1796
rect 2973 1788 3007 1790
rect 3055 1788 3071 1804
rect 3072 1794 3280 1804
rect 3281 1794 3297 1804
rect 3345 1800 3360 1815
rect 3363 1812 3364 1824
rect 3371 1812 3398 1824
rect 3363 1804 3398 1812
rect 3363 1803 3392 1804
rect 3083 1790 3297 1794
rect 3098 1788 3297 1790
rect 3332 1790 3345 1800
rect 3363 1790 3380 1803
rect 3332 1788 3380 1790
rect 2974 1784 3007 1788
rect 2970 1782 3007 1784
rect 2970 1781 3037 1782
rect 2970 1776 3001 1781
rect 3007 1776 3037 1781
rect 2970 1772 3037 1776
rect 2943 1769 3037 1772
rect 2943 1762 2992 1769
rect 2943 1756 2973 1762
rect 2992 1757 2997 1762
rect 2909 1740 2989 1756
rect 3001 1748 3037 1769
rect 3098 1764 3287 1788
rect 3332 1787 3379 1788
rect 3345 1782 3379 1787
rect 3113 1761 3287 1764
rect 3106 1758 3287 1761
rect 3315 1781 3379 1782
rect 2909 1738 2928 1740
rect 2943 1738 2977 1740
rect 2909 1722 2989 1738
rect 2909 1716 2928 1722
rect 2625 1690 2728 1700
rect 2579 1688 2728 1690
rect 2749 1688 2784 1700
rect 2418 1686 2580 1688
rect 2430 1666 2449 1686
rect 2464 1684 2494 1686
rect 2313 1658 2354 1666
rect 2436 1662 2449 1666
rect 2501 1670 2580 1686
rect 2612 1686 2784 1688
rect 2612 1670 2691 1686
rect 2698 1684 2728 1686
rect 2276 1648 2305 1658
rect 2319 1648 2348 1658
rect 2363 1648 2393 1662
rect 2436 1648 2479 1662
rect 2501 1658 2691 1670
rect 2756 1666 2762 1686
rect 2486 1648 2516 1658
rect 2517 1648 2675 1658
rect 2679 1648 2709 1658
rect 2713 1648 2743 1662
rect 2771 1648 2784 1686
rect 2856 1700 2885 1716
rect 2899 1700 2928 1716
rect 2943 1706 2973 1722
rect 3001 1700 3007 1748
rect 3010 1742 3029 1748
rect 3044 1742 3074 1750
rect 3010 1734 3074 1742
rect 3010 1718 3090 1734
rect 3106 1727 3168 1758
rect 3184 1727 3246 1758
rect 3315 1756 3364 1781
rect 3379 1756 3409 1772
rect 3278 1742 3308 1750
rect 3315 1748 3425 1756
rect 3278 1734 3323 1742
rect 3010 1716 3029 1718
rect 3044 1716 3090 1718
rect 3010 1700 3090 1716
rect 3117 1714 3152 1727
rect 3193 1724 3230 1727
rect 3193 1722 3235 1724
rect 3122 1711 3152 1714
rect 3131 1707 3138 1711
rect 3138 1706 3139 1707
rect 3097 1700 3107 1706
rect 2856 1692 2891 1700
rect 2856 1666 2857 1692
rect 2864 1666 2891 1692
rect 2799 1648 2829 1662
rect 2856 1658 2891 1666
rect 2893 1692 2934 1700
rect 2893 1666 2908 1692
rect 2915 1666 2934 1692
rect 2998 1688 3029 1700
rect 3044 1688 3147 1700
rect 3159 1690 3185 1716
rect 3200 1711 3230 1722
rect 3262 1718 3324 1734
rect 3262 1716 3308 1718
rect 3262 1700 3324 1716
rect 3336 1700 3342 1748
rect 3345 1740 3425 1748
rect 3345 1738 3364 1740
rect 3379 1738 3413 1740
rect 3345 1722 3425 1738
rect 3345 1700 3364 1722
rect 3379 1706 3409 1722
rect 3437 1716 3443 1790
rect 3446 1716 3465 1860
rect 3480 1716 3486 1860
rect 3495 1790 3508 1860
rect 3560 1856 3582 1860
rect 3553 1834 3582 1848
rect 3635 1834 3651 1848
rect 3689 1844 3695 1846
rect 3702 1844 3810 1860
rect 3817 1844 3823 1846
rect 3831 1844 3846 1860
rect 3912 1854 3931 1857
rect 3553 1832 3651 1834
rect 3678 1832 3846 1844
rect 3861 1834 3877 1848
rect 3912 1835 3934 1854
rect 3944 1848 3960 1849
rect 3943 1846 3960 1848
rect 3944 1841 3960 1846
rect 3934 1834 3940 1835
rect 3943 1834 3972 1841
rect 3861 1833 3972 1834
rect 3861 1832 3978 1833
rect 3537 1824 3588 1832
rect 3635 1824 3669 1832
rect 3537 1812 3562 1824
rect 3569 1812 3588 1824
rect 3642 1822 3669 1824
rect 3678 1822 3899 1832
rect 3934 1829 3940 1832
rect 3642 1818 3899 1822
rect 3537 1804 3588 1812
rect 3635 1804 3899 1818
rect 3943 1824 3978 1832
rect 3489 1756 3508 1790
rect 3553 1796 3582 1804
rect 3553 1790 3570 1796
rect 3553 1788 3587 1790
rect 3635 1788 3651 1804
rect 3652 1794 3860 1804
rect 3861 1794 3877 1804
rect 3925 1800 3940 1815
rect 3943 1812 3944 1824
rect 3951 1812 3978 1824
rect 3943 1804 3978 1812
rect 3943 1803 3972 1804
rect 3663 1790 3877 1794
rect 3678 1788 3877 1790
rect 3912 1790 3925 1800
rect 3943 1790 3960 1803
rect 3912 1788 3960 1790
rect 3554 1784 3587 1788
rect 3550 1782 3587 1784
rect 3550 1781 3617 1782
rect 3550 1776 3581 1781
rect 3587 1776 3617 1781
rect 3550 1772 3617 1776
rect 3523 1769 3617 1772
rect 3523 1762 3572 1769
rect 3523 1756 3553 1762
rect 3572 1757 3577 1762
rect 3489 1740 3569 1756
rect 3581 1748 3617 1769
rect 3678 1764 3867 1788
rect 3912 1787 3959 1788
rect 3925 1782 3959 1787
rect 3693 1761 3867 1764
rect 3686 1758 3867 1761
rect 3895 1781 3959 1782
rect 3489 1738 3508 1740
rect 3523 1738 3557 1740
rect 3489 1722 3569 1738
rect 3489 1716 3508 1722
rect 3205 1690 3308 1700
rect 3159 1688 3308 1690
rect 3329 1688 3364 1700
rect 2998 1686 3160 1688
rect 3010 1666 3029 1686
rect 3044 1684 3074 1686
rect 2893 1658 2934 1666
rect 3016 1662 3029 1666
rect 3081 1670 3160 1686
rect 3192 1686 3364 1688
rect 3192 1670 3271 1686
rect 3278 1684 3308 1686
rect 2856 1648 2885 1658
rect 2899 1648 2928 1658
rect 2943 1648 2973 1662
rect 3016 1648 3059 1662
rect 3081 1658 3271 1670
rect 3336 1666 3342 1686
rect 3066 1648 3096 1658
rect 3097 1648 3255 1658
rect 3259 1648 3289 1658
rect 3293 1648 3323 1662
rect 3351 1648 3364 1686
rect 3436 1700 3465 1716
rect 3479 1700 3508 1716
rect 3523 1706 3553 1722
rect 3581 1700 3587 1748
rect 3590 1742 3609 1748
rect 3624 1742 3654 1750
rect 3590 1734 3654 1742
rect 3590 1718 3670 1734
rect 3686 1727 3748 1758
rect 3764 1727 3826 1758
rect 3895 1756 3944 1781
rect 3959 1756 3989 1772
rect 3858 1742 3888 1750
rect 3895 1748 4005 1756
rect 3858 1734 3903 1742
rect 3590 1716 3609 1718
rect 3624 1716 3670 1718
rect 3590 1700 3670 1716
rect 3697 1714 3732 1727
rect 3773 1724 3810 1727
rect 3773 1722 3815 1724
rect 3702 1711 3732 1714
rect 3711 1707 3718 1711
rect 3718 1706 3719 1707
rect 3677 1700 3687 1706
rect 3436 1692 3471 1700
rect 3436 1666 3437 1692
rect 3444 1666 3471 1692
rect 3379 1648 3409 1662
rect 3436 1658 3471 1666
rect 3473 1692 3514 1700
rect 3473 1666 3488 1692
rect 3495 1666 3514 1692
rect 3578 1688 3609 1700
rect 3624 1688 3727 1700
rect 3739 1690 3765 1716
rect 3780 1711 3810 1722
rect 3842 1718 3904 1734
rect 3842 1716 3888 1718
rect 3842 1700 3904 1716
rect 3916 1700 3922 1748
rect 3925 1740 4005 1748
rect 3925 1738 3944 1740
rect 3959 1738 3993 1740
rect 3925 1722 4005 1738
rect 3925 1700 3944 1722
rect 3959 1706 3989 1722
rect 4017 1716 4023 1790
rect 4026 1716 4045 1860
rect 4060 1716 4066 1860
rect 4075 1790 4088 1860
rect 4140 1856 4162 1860
rect 4133 1834 4162 1848
rect 4215 1834 4231 1848
rect 4269 1844 4275 1846
rect 4282 1844 4390 1860
rect 4397 1844 4403 1846
rect 4411 1844 4426 1860
rect 4492 1854 4511 1857
rect 4133 1832 4231 1834
rect 4258 1832 4426 1844
rect 4441 1834 4457 1848
rect 4492 1835 4514 1854
rect 4524 1848 4540 1849
rect 4523 1846 4540 1848
rect 4524 1841 4540 1846
rect 4514 1834 4520 1835
rect 4523 1834 4552 1841
rect 4441 1833 4552 1834
rect 4441 1832 4558 1833
rect 4117 1824 4168 1832
rect 4215 1824 4249 1832
rect 4117 1812 4142 1824
rect 4149 1812 4168 1824
rect 4222 1822 4249 1824
rect 4258 1822 4479 1832
rect 4514 1829 4520 1832
rect 4222 1818 4479 1822
rect 4117 1804 4168 1812
rect 4215 1804 4479 1818
rect 4523 1824 4558 1832
rect 4069 1756 4088 1790
rect 4133 1796 4162 1804
rect 4133 1790 4150 1796
rect 4133 1788 4167 1790
rect 4215 1788 4231 1804
rect 4232 1794 4440 1804
rect 4441 1794 4457 1804
rect 4505 1800 4520 1815
rect 4523 1812 4524 1824
rect 4531 1812 4558 1824
rect 4523 1804 4558 1812
rect 4523 1803 4552 1804
rect 4243 1790 4457 1794
rect 4258 1788 4457 1790
rect 4492 1790 4505 1800
rect 4523 1790 4540 1803
rect 4492 1788 4540 1790
rect 4134 1784 4167 1788
rect 4130 1782 4167 1784
rect 4130 1781 4197 1782
rect 4130 1776 4161 1781
rect 4167 1776 4197 1781
rect 4130 1772 4197 1776
rect 4103 1769 4197 1772
rect 4103 1762 4152 1769
rect 4103 1756 4133 1762
rect 4152 1757 4157 1762
rect 4069 1740 4149 1756
rect 4161 1748 4197 1769
rect 4258 1764 4447 1788
rect 4492 1787 4539 1788
rect 4505 1782 4539 1787
rect 4273 1761 4447 1764
rect 4266 1758 4447 1761
rect 4475 1781 4539 1782
rect 4069 1738 4088 1740
rect 4103 1738 4137 1740
rect 4069 1722 4149 1738
rect 4069 1716 4088 1722
rect 3785 1690 3888 1700
rect 3739 1688 3888 1690
rect 3909 1688 3944 1700
rect 3578 1686 3740 1688
rect 3590 1666 3609 1686
rect 3624 1684 3654 1686
rect 3473 1658 3514 1666
rect 3596 1662 3609 1666
rect 3661 1670 3740 1686
rect 3772 1686 3944 1688
rect 3772 1670 3851 1686
rect 3858 1684 3888 1686
rect 3436 1648 3465 1658
rect 3479 1648 3508 1658
rect 3523 1648 3553 1662
rect 3596 1648 3639 1662
rect 3661 1658 3851 1670
rect 3916 1666 3922 1686
rect 3646 1648 3676 1658
rect 3677 1648 3835 1658
rect 3839 1648 3869 1658
rect 3873 1648 3903 1662
rect 3931 1648 3944 1686
rect 4016 1700 4045 1716
rect 4059 1700 4088 1716
rect 4103 1706 4133 1722
rect 4161 1700 4167 1748
rect 4170 1742 4189 1748
rect 4204 1742 4234 1750
rect 4170 1734 4234 1742
rect 4170 1718 4250 1734
rect 4266 1727 4328 1758
rect 4344 1727 4406 1758
rect 4475 1756 4524 1781
rect 4539 1756 4569 1772
rect 4438 1742 4468 1750
rect 4475 1748 4585 1756
rect 4438 1734 4483 1742
rect 4170 1716 4189 1718
rect 4204 1716 4250 1718
rect 4170 1700 4250 1716
rect 4277 1714 4312 1727
rect 4353 1724 4390 1727
rect 4353 1722 4395 1724
rect 4282 1711 4312 1714
rect 4291 1707 4298 1711
rect 4298 1706 4299 1707
rect 4257 1700 4267 1706
rect 4016 1692 4051 1700
rect 4016 1666 4017 1692
rect 4024 1666 4051 1692
rect 3959 1648 3989 1662
rect 4016 1658 4051 1666
rect 4053 1692 4094 1700
rect 4053 1666 4068 1692
rect 4075 1666 4094 1692
rect 4158 1688 4189 1700
rect 4204 1688 4307 1700
rect 4319 1690 4345 1716
rect 4360 1711 4390 1722
rect 4422 1718 4484 1734
rect 4422 1716 4468 1718
rect 4422 1700 4484 1716
rect 4496 1700 4502 1748
rect 4505 1740 4585 1748
rect 4505 1738 4524 1740
rect 4539 1738 4573 1740
rect 4505 1722 4585 1738
rect 4505 1700 4524 1722
rect 4539 1706 4569 1722
rect 4597 1716 4603 1790
rect 4606 1716 4625 1860
rect 4640 1716 4646 1860
rect 4655 1790 4668 1860
rect 4720 1856 4742 1860
rect 4713 1834 4742 1848
rect 4795 1834 4811 1848
rect 4849 1844 4855 1846
rect 4862 1844 4970 1860
rect 4977 1844 4983 1846
rect 4991 1844 5006 1860
rect 5072 1854 5091 1857
rect 4713 1832 4811 1834
rect 4838 1832 5006 1844
rect 5021 1834 5037 1848
rect 5072 1835 5094 1854
rect 5104 1848 5120 1849
rect 5103 1846 5120 1848
rect 5104 1841 5120 1846
rect 5094 1834 5100 1835
rect 5103 1834 5132 1841
rect 5021 1833 5132 1834
rect 5021 1832 5138 1833
rect 4697 1824 4748 1832
rect 4795 1824 4829 1832
rect 4697 1812 4722 1824
rect 4729 1812 4748 1824
rect 4802 1822 4829 1824
rect 4838 1822 5059 1832
rect 5094 1829 5100 1832
rect 4802 1818 5059 1822
rect 4697 1804 4748 1812
rect 4795 1804 5059 1818
rect 5103 1824 5138 1832
rect 4649 1756 4668 1790
rect 4713 1796 4742 1804
rect 4713 1790 4730 1796
rect 4713 1788 4747 1790
rect 4795 1788 4811 1804
rect 4812 1794 5020 1804
rect 5021 1794 5037 1804
rect 5085 1800 5100 1815
rect 5103 1812 5104 1824
rect 5111 1812 5138 1824
rect 5103 1804 5138 1812
rect 5103 1803 5132 1804
rect 4823 1790 5037 1794
rect 4838 1788 5037 1790
rect 5072 1790 5085 1800
rect 5103 1790 5120 1803
rect 5072 1788 5120 1790
rect 4714 1784 4747 1788
rect 4710 1782 4747 1784
rect 4710 1781 4777 1782
rect 4710 1776 4741 1781
rect 4747 1776 4777 1781
rect 4710 1772 4777 1776
rect 4683 1769 4777 1772
rect 4683 1762 4732 1769
rect 4683 1756 4713 1762
rect 4732 1757 4737 1762
rect 4649 1740 4729 1756
rect 4741 1748 4777 1769
rect 4838 1764 5027 1788
rect 5072 1787 5119 1788
rect 5085 1782 5119 1787
rect 4853 1761 5027 1764
rect 4846 1758 5027 1761
rect 5055 1781 5119 1782
rect 4649 1738 4668 1740
rect 4683 1738 4717 1740
rect 4649 1722 4729 1738
rect 4649 1716 4668 1722
rect 4365 1690 4468 1700
rect 4319 1688 4468 1690
rect 4489 1688 4524 1700
rect 4158 1686 4320 1688
rect 4170 1666 4189 1686
rect 4204 1684 4234 1686
rect 4053 1658 4094 1666
rect 4176 1662 4189 1666
rect 4241 1670 4320 1686
rect 4352 1686 4524 1688
rect 4352 1670 4431 1686
rect 4438 1684 4468 1686
rect 4016 1648 4045 1658
rect 4059 1648 4088 1658
rect 4103 1648 4133 1662
rect 4176 1648 4219 1662
rect 4241 1658 4431 1670
rect 4496 1666 4502 1686
rect 4226 1648 4256 1658
rect 4257 1648 4415 1658
rect 4419 1648 4449 1658
rect 4453 1648 4483 1662
rect 4511 1648 4524 1686
rect 4596 1700 4625 1716
rect 4639 1700 4668 1716
rect 4683 1706 4713 1722
rect 4741 1700 4747 1748
rect 4750 1742 4769 1748
rect 4784 1742 4814 1750
rect 4750 1734 4814 1742
rect 4750 1718 4830 1734
rect 4846 1727 4908 1758
rect 4924 1727 4986 1758
rect 5055 1756 5104 1781
rect 5119 1756 5149 1772
rect 5018 1742 5048 1750
rect 5055 1748 5165 1756
rect 5018 1734 5063 1742
rect 4750 1716 4769 1718
rect 4784 1716 4830 1718
rect 4750 1700 4830 1716
rect 4857 1714 4892 1727
rect 4933 1724 4970 1727
rect 4933 1722 4975 1724
rect 4862 1711 4892 1714
rect 4871 1707 4878 1711
rect 4878 1706 4879 1707
rect 4837 1700 4847 1706
rect 4596 1692 4631 1700
rect 4596 1666 4597 1692
rect 4604 1666 4631 1692
rect 4539 1648 4569 1662
rect 4596 1658 4631 1666
rect 4633 1692 4674 1700
rect 4633 1666 4648 1692
rect 4655 1666 4674 1692
rect 4738 1688 4769 1700
rect 4784 1688 4887 1700
rect 4899 1690 4925 1716
rect 4940 1711 4970 1722
rect 5002 1718 5064 1734
rect 5002 1716 5048 1718
rect 5002 1700 5064 1716
rect 5076 1700 5082 1748
rect 5085 1740 5165 1748
rect 5085 1738 5104 1740
rect 5119 1738 5153 1740
rect 5085 1722 5165 1738
rect 5085 1700 5104 1722
rect 5119 1706 5149 1722
rect 5177 1716 5183 1790
rect 5186 1716 5205 1860
rect 5220 1716 5226 1860
rect 5235 1790 5248 1860
rect 5300 1856 5322 1860
rect 5293 1834 5322 1848
rect 5375 1834 5391 1848
rect 5429 1844 5435 1846
rect 5442 1844 5550 1860
rect 5557 1844 5563 1846
rect 5571 1844 5586 1860
rect 5652 1854 5671 1857
rect 5293 1832 5391 1834
rect 5418 1832 5586 1844
rect 5601 1834 5617 1848
rect 5652 1835 5674 1854
rect 5684 1848 5700 1849
rect 5683 1846 5700 1848
rect 5684 1841 5700 1846
rect 5674 1834 5680 1835
rect 5683 1834 5712 1841
rect 5601 1833 5712 1834
rect 5601 1832 5718 1833
rect 5277 1824 5328 1832
rect 5375 1824 5409 1832
rect 5277 1812 5302 1824
rect 5309 1812 5328 1824
rect 5382 1822 5409 1824
rect 5418 1822 5639 1832
rect 5674 1829 5680 1832
rect 5382 1818 5639 1822
rect 5277 1804 5328 1812
rect 5375 1804 5639 1818
rect 5683 1824 5718 1832
rect 5229 1756 5248 1790
rect 5293 1796 5322 1804
rect 5293 1790 5310 1796
rect 5293 1788 5327 1790
rect 5375 1788 5391 1804
rect 5392 1794 5600 1804
rect 5601 1794 5617 1804
rect 5665 1800 5680 1815
rect 5683 1812 5684 1824
rect 5691 1812 5718 1824
rect 5683 1804 5718 1812
rect 5683 1803 5712 1804
rect 5403 1790 5617 1794
rect 5418 1788 5617 1790
rect 5652 1790 5665 1800
rect 5683 1790 5700 1803
rect 5652 1788 5700 1790
rect 5294 1784 5327 1788
rect 5290 1782 5327 1784
rect 5290 1781 5357 1782
rect 5290 1776 5321 1781
rect 5327 1776 5357 1781
rect 5290 1772 5357 1776
rect 5263 1769 5357 1772
rect 5263 1762 5312 1769
rect 5263 1756 5293 1762
rect 5312 1757 5317 1762
rect 5229 1740 5309 1756
rect 5321 1748 5357 1769
rect 5418 1764 5607 1788
rect 5652 1787 5699 1788
rect 5665 1782 5699 1787
rect 5433 1761 5607 1764
rect 5426 1758 5607 1761
rect 5635 1781 5699 1782
rect 5229 1738 5248 1740
rect 5263 1738 5297 1740
rect 5229 1722 5309 1738
rect 5229 1716 5248 1722
rect 4945 1690 5048 1700
rect 4899 1688 5048 1690
rect 5069 1688 5104 1700
rect 4738 1686 4900 1688
rect 4750 1666 4769 1686
rect 4784 1684 4814 1686
rect 4633 1658 4674 1666
rect 4756 1662 4769 1666
rect 4821 1670 4900 1686
rect 4932 1686 5104 1688
rect 4932 1670 5011 1686
rect 5018 1684 5048 1686
rect 4596 1648 4625 1658
rect 4639 1648 4668 1658
rect 4683 1648 4713 1662
rect 4756 1648 4799 1662
rect 4821 1658 5011 1670
rect 5076 1666 5082 1686
rect 4806 1648 4836 1658
rect 4837 1648 4995 1658
rect 4999 1648 5029 1658
rect 5033 1648 5063 1662
rect 5091 1648 5104 1686
rect 5176 1700 5205 1716
rect 5219 1700 5248 1716
rect 5263 1706 5293 1722
rect 5321 1700 5327 1748
rect 5330 1742 5349 1748
rect 5364 1742 5394 1750
rect 5330 1734 5394 1742
rect 5330 1718 5410 1734
rect 5426 1727 5488 1758
rect 5504 1727 5566 1758
rect 5635 1756 5684 1781
rect 5699 1756 5729 1772
rect 5598 1742 5628 1750
rect 5635 1748 5745 1756
rect 5598 1734 5643 1742
rect 5330 1716 5349 1718
rect 5364 1716 5410 1718
rect 5330 1700 5410 1716
rect 5437 1714 5472 1727
rect 5513 1724 5550 1727
rect 5513 1722 5555 1724
rect 5442 1711 5472 1714
rect 5451 1707 5458 1711
rect 5458 1706 5459 1707
rect 5417 1700 5427 1706
rect 5176 1692 5211 1700
rect 5176 1666 5177 1692
rect 5184 1666 5211 1692
rect 5119 1648 5149 1662
rect 5176 1658 5211 1666
rect 5213 1692 5254 1700
rect 5213 1666 5228 1692
rect 5235 1666 5254 1692
rect 5318 1688 5349 1700
rect 5364 1688 5467 1700
rect 5479 1690 5505 1716
rect 5520 1711 5550 1722
rect 5582 1718 5644 1734
rect 5582 1716 5628 1718
rect 5582 1700 5644 1716
rect 5656 1700 5662 1748
rect 5665 1740 5745 1748
rect 5665 1738 5684 1740
rect 5699 1738 5733 1740
rect 5665 1722 5745 1738
rect 5665 1700 5684 1722
rect 5699 1706 5729 1722
rect 5757 1716 5763 1790
rect 5766 1716 5785 1860
rect 5800 1716 5806 1860
rect 5815 1790 5828 1860
rect 5880 1856 5902 1860
rect 5873 1834 5902 1848
rect 5955 1834 5971 1848
rect 6009 1844 6015 1846
rect 6022 1844 6130 1860
rect 6137 1844 6143 1846
rect 6151 1844 6166 1860
rect 6232 1854 6251 1857
rect 5873 1832 5971 1834
rect 5998 1832 6166 1844
rect 6181 1834 6197 1848
rect 6232 1835 6254 1854
rect 6264 1848 6280 1849
rect 6263 1846 6280 1848
rect 6264 1841 6280 1846
rect 6254 1834 6260 1835
rect 6263 1834 6292 1841
rect 6181 1833 6292 1834
rect 6181 1832 6298 1833
rect 5857 1824 5908 1832
rect 5955 1824 5989 1832
rect 5857 1812 5882 1824
rect 5889 1812 5908 1824
rect 5962 1822 5989 1824
rect 5998 1822 6219 1832
rect 6254 1829 6260 1832
rect 5962 1818 6219 1822
rect 5857 1804 5908 1812
rect 5955 1804 6219 1818
rect 6263 1824 6298 1832
rect 5809 1756 5828 1790
rect 5873 1796 5902 1804
rect 5873 1790 5890 1796
rect 5873 1788 5907 1790
rect 5955 1788 5971 1804
rect 5972 1794 6180 1804
rect 6181 1794 6197 1804
rect 6245 1800 6260 1815
rect 6263 1812 6264 1824
rect 6271 1812 6298 1824
rect 6263 1804 6298 1812
rect 6263 1803 6292 1804
rect 5983 1790 6197 1794
rect 5998 1788 6197 1790
rect 6232 1790 6245 1800
rect 6263 1790 6280 1803
rect 6232 1788 6280 1790
rect 5874 1784 5907 1788
rect 5870 1782 5907 1784
rect 5870 1781 5937 1782
rect 5870 1776 5901 1781
rect 5907 1776 5937 1781
rect 5870 1772 5937 1776
rect 5843 1769 5937 1772
rect 5843 1762 5892 1769
rect 5843 1756 5873 1762
rect 5892 1757 5897 1762
rect 5809 1740 5889 1756
rect 5901 1748 5937 1769
rect 5998 1764 6187 1788
rect 6232 1787 6279 1788
rect 6245 1782 6279 1787
rect 6013 1761 6187 1764
rect 6006 1758 6187 1761
rect 6215 1781 6279 1782
rect 5809 1738 5828 1740
rect 5843 1738 5877 1740
rect 5809 1722 5889 1738
rect 5809 1716 5828 1722
rect 5525 1690 5628 1700
rect 5479 1688 5628 1690
rect 5649 1688 5684 1700
rect 5318 1686 5480 1688
rect 5330 1666 5349 1686
rect 5364 1684 5394 1686
rect 5213 1658 5254 1666
rect 5336 1662 5349 1666
rect 5401 1670 5480 1686
rect 5512 1686 5684 1688
rect 5512 1670 5591 1686
rect 5598 1684 5628 1686
rect 5176 1648 5205 1658
rect 5219 1648 5248 1658
rect 5263 1648 5293 1662
rect 5336 1648 5379 1662
rect 5401 1658 5591 1670
rect 5656 1666 5662 1686
rect 5386 1648 5416 1658
rect 5417 1648 5575 1658
rect 5579 1648 5609 1658
rect 5613 1648 5643 1662
rect 5671 1648 5684 1686
rect 5756 1700 5785 1716
rect 5799 1700 5828 1716
rect 5843 1706 5873 1722
rect 5901 1700 5907 1748
rect 5910 1742 5929 1748
rect 5944 1742 5974 1750
rect 5910 1734 5974 1742
rect 5910 1718 5990 1734
rect 6006 1727 6068 1758
rect 6084 1727 6146 1758
rect 6215 1756 6264 1781
rect 6279 1756 6309 1772
rect 6178 1742 6208 1750
rect 6215 1748 6325 1756
rect 6178 1734 6223 1742
rect 5910 1716 5929 1718
rect 5944 1716 5990 1718
rect 5910 1700 5990 1716
rect 6017 1714 6052 1727
rect 6093 1724 6130 1727
rect 6093 1722 6135 1724
rect 6022 1711 6052 1714
rect 6031 1707 6038 1711
rect 6038 1706 6039 1707
rect 5997 1700 6007 1706
rect 5756 1692 5791 1700
rect 5756 1666 5757 1692
rect 5764 1666 5791 1692
rect 5699 1648 5729 1662
rect 5756 1658 5791 1666
rect 5793 1692 5834 1700
rect 5793 1666 5808 1692
rect 5815 1666 5834 1692
rect 5898 1688 5929 1700
rect 5944 1688 6047 1700
rect 6059 1690 6085 1716
rect 6100 1711 6130 1722
rect 6162 1718 6224 1734
rect 6162 1716 6208 1718
rect 6162 1700 6224 1716
rect 6236 1700 6242 1748
rect 6245 1740 6325 1748
rect 6245 1738 6264 1740
rect 6279 1738 6313 1740
rect 6245 1722 6325 1738
rect 6245 1700 6264 1722
rect 6279 1706 6309 1722
rect 6337 1716 6343 1790
rect 6346 1716 6365 1860
rect 6380 1716 6386 1860
rect 6395 1790 6408 1860
rect 6460 1856 6482 1860
rect 6453 1834 6482 1848
rect 6535 1834 6551 1848
rect 6589 1844 6595 1846
rect 6602 1844 6710 1860
rect 6717 1844 6723 1846
rect 6731 1844 6746 1860
rect 6812 1854 6831 1857
rect 6453 1832 6551 1834
rect 6578 1832 6746 1844
rect 6761 1834 6777 1848
rect 6812 1835 6834 1854
rect 6844 1848 6860 1849
rect 6843 1846 6860 1848
rect 6844 1841 6860 1846
rect 6834 1834 6840 1835
rect 6843 1834 6872 1841
rect 6761 1833 6872 1834
rect 6761 1832 6878 1833
rect 6437 1824 6488 1832
rect 6535 1824 6569 1832
rect 6437 1812 6462 1824
rect 6469 1812 6488 1824
rect 6542 1822 6569 1824
rect 6578 1822 6799 1832
rect 6834 1829 6840 1832
rect 6542 1818 6799 1822
rect 6437 1804 6488 1812
rect 6535 1804 6799 1818
rect 6843 1824 6878 1832
rect 6389 1756 6408 1790
rect 6453 1796 6482 1804
rect 6453 1790 6470 1796
rect 6453 1788 6487 1790
rect 6535 1788 6551 1804
rect 6552 1794 6760 1804
rect 6761 1794 6777 1804
rect 6825 1800 6840 1815
rect 6843 1812 6844 1824
rect 6851 1812 6878 1824
rect 6843 1804 6878 1812
rect 6843 1803 6872 1804
rect 6563 1790 6777 1794
rect 6578 1788 6777 1790
rect 6812 1790 6825 1800
rect 6843 1790 6860 1803
rect 6812 1788 6860 1790
rect 6454 1784 6487 1788
rect 6450 1782 6487 1784
rect 6450 1781 6517 1782
rect 6450 1776 6481 1781
rect 6487 1776 6517 1781
rect 6450 1772 6517 1776
rect 6423 1769 6517 1772
rect 6423 1762 6472 1769
rect 6423 1756 6453 1762
rect 6472 1757 6477 1762
rect 6389 1740 6469 1756
rect 6481 1748 6517 1769
rect 6578 1764 6767 1788
rect 6812 1787 6859 1788
rect 6825 1782 6859 1787
rect 6593 1761 6767 1764
rect 6586 1758 6767 1761
rect 6795 1781 6859 1782
rect 6389 1738 6408 1740
rect 6423 1738 6457 1740
rect 6389 1722 6469 1738
rect 6389 1716 6408 1722
rect 6105 1690 6208 1700
rect 6059 1688 6208 1690
rect 6229 1688 6264 1700
rect 5898 1686 6060 1688
rect 5910 1666 5929 1686
rect 5944 1684 5974 1686
rect 5793 1658 5834 1666
rect 5916 1662 5929 1666
rect 5981 1670 6060 1686
rect 6092 1686 6264 1688
rect 6092 1670 6171 1686
rect 6178 1684 6208 1686
rect 5756 1648 5785 1658
rect 5799 1648 5828 1658
rect 5843 1648 5873 1662
rect 5916 1648 5959 1662
rect 5981 1658 6171 1670
rect 6236 1666 6242 1686
rect 5966 1648 5996 1658
rect 5997 1648 6155 1658
rect 6159 1648 6189 1658
rect 6193 1648 6223 1662
rect 6251 1648 6264 1686
rect 6336 1700 6365 1716
rect 6379 1700 6408 1716
rect 6423 1706 6453 1722
rect 6481 1700 6487 1748
rect 6490 1742 6509 1748
rect 6524 1742 6554 1750
rect 6490 1734 6554 1742
rect 6490 1718 6570 1734
rect 6586 1727 6648 1758
rect 6664 1727 6726 1758
rect 6795 1756 6844 1781
rect 6859 1756 6889 1772
rect 6758 1742 6788 1750
rect 6795 1748 6905 1756
rect 6758 1734 6803 1742
rect 6490 1716 6509 1718
rect 6524 1716 6570 1718
rect 6490 1700 6570 1716
rect 6597 1714 6632 1727
rect 6673 1724 6710 1727
rect 6673 1722 6715 1724
rect 6602 1711 6632 1714
rect 6611 1707 6618 1711
rect 6618 1706 6619 1707
rect 6577 1700 6587 1706
rect 6336 1692 6371 1700
rect 6336 1666 6337 1692
rect 6344 1666 6371 1692
rect 6279 1648 6309 1662
rect 6336 1658 6371 1666
rect 6373 1692 6414 1700
rect 6373 1666 6388 1692
rect 6395 1666 6414 1692
rect 6478 1688 6509 1700
rect 6524 1688 6627 1700
rect 6639 1690 6665 1716
rect 6680 1711 6710 1722
rect 6742 1718 6804 1734
rect 6742 1716 6788 1718
rect 6742 1700 6804 1716
rect 6816 1700 6822 1748
rect 6825 1740 6905 1748
rect 6825 1738 6844 1740
rect 6859 1738 6893 1740
rect 6825 1722 6905 1738
rect 6825 1700 6844 1722
rect 6859 1706 6889 1722
rect 6917 1716 6923 1790
rect 6926 1716 6945 1860
rect 6960 1716 6966 1860
rect 6975 1790 6988 1860
rect 7040 1856 7062 1860
rect 7033 1834 7062 1848
rect 7115 1834 7131 1848
rect 7169 1844 7175 1846
rect 7182 1844 7290 1860
rect 7297 1844 7303 1846
rect 7311 1844 7326 1860
rect 7392 1854 7411 1857
rect 7033 1832 7131 1834
rect 7158 1832 7326 1844
rect 7341 1834 7357 1848
rect 7392 1835 7414 1854
rect 7424 1848 7440 1849
rect 7423 1846 7440 1848
rect 7424 1841 7440 1846
rect 7414 1834 7420 1835
rect 7423 1834 7452 1841
rect 7341 1833 7452 1834
rect 7341 1832 7458 1833
rect 7017 1824 7068 1832
rect 7115 1824 7149 1832
rect 7017 1812 7042 1824
rect 7049 1812 7068 1824
rect 7122 1822 7149 1824
rect 7158 1822 7379 1832
rect 7414 1829 7420 1832
rect 7122 1818 7379 1822
rect 7017 1804 7068 1812
rect 7115 1804 7379 1818
rect 7423 1824 7458 1832
rect 6969 1756 6988 1790
rect 7033 1796 7062 1804
rect 7033 1790 7050 1796
rect 7033 1788 7067 1790
rect 7115 1788 7131 1804
rect 7132 1794 7340 1804
rect 7341 1794 7357 1804
rect 7405 1800 7420 1815
rect 7423 1812 7424 1824
rect 7431 1812 7458 1824
rect 7423 1804 7458 1812
rect 7423 1803 7452 1804
rect 7143 1790 7357 1794
rect 7158 1788 7357 1790
rect 7392 1790 7405 1800
rect 7423 1790 7440 1803
rect 7392 1788 7440 1790
rect 7034 1784 7067 1788
rect 7030 1782 7067 1784
rect 7030 1781 7097 1782
rect 7030 1776 7061 1781
rect 7067 1776 7097 1781
rect 7030 1772 7097 1776
rect 7003 1769 7097 1772
rect 7003 1762 7052 1769
rect 7003 1756 7033 1762
rect 7052 1757 7057 1762
rect 6969 1740 7049 1756
rect 7061 1748 7097 1769
rect 7158 1764 7347 1788
rect 7392 1787 7439 1788
rect 7405 1782 7439 1787
rect 7173 1761 7347 1764
rect 7166 1758 7347 1761
rect 7375 1781 7439 1782
rect 6969 1738 6988 1740
rect 7003 1738 7037 1740
rect 6969 1722 7049 1738
rect 6969 1716 6988 1722
rect 6685 1690 6788 1700
rect 6639 1688 6788 1690
rect 6809 1688 6844 1700
rect 6478 1686 6640 1688
rect 6490 1666 6509 1686
rect 6524 1684 6554 1686
rect 6373 1658 6414 1666
rect 6496 1662 6509 1666
rect 6561 1670 6640 1686
rect 6672 1686 6844 1688
rect 6672 1670 6751 1686
rect 6758 1684 6788 1686
rect 6336 1648 6365 1658
rect 6379 1648 6408 1658
rect 6423 1648 6453 1662
rect 6496 1648 6539 1662
rect 6561 1658 6751 1670
rect 6816 1666 6822 1686
rect 6546 1648 6576 1658
rect 6577 1648 6735 1658
rect 6739 1648 6769 1658
rect 6773 1648 6803 1662
rect 6831 1648 6844 1686
rect 6916 1700 6945 1716
rect 6959 1700 6988 1716
rect 7003 1706 7033 1722
rect 7061 1700 7067 1748
rect 7070 1742 7089 1748
rect 7104 1742 7134 1750
rect 7070 1734 7134 1742
rect 7070 1718 7150 1734
rect 7166 1727 7228 1758
rect 7244 1727 7306 1758
rect 7375 1756 7424 1781
rect 7439 1756 7469 1772
rect 7338 1742 7368 1750
rect 7375 1748 7485 1756
rect 7338 1734 7383 1742
rect 7070 1716 7089 1718
rect 7104 1716 7150 1718
rect 7070 1700 7150 1716
rect 7177 1714 7212 1727
rect 7253 1724 7290 1727
rect 7253 1722 7295 1724
rect 7182 1711 7212 1714
rect 7191 1707 7198 1711
rect 7198 1706 7199 1707
rect 7157 1700 7167 1706
rect 6916 1692 6951 1700
rect 6916 1666 6917 1692
rect 6924 1666 6951 1692
rect 6859 1648 6889 1662
rect 6916 1658 6951 1666
rect 6953 1692 6994 1700
rect 6953 1666 6968 1692
rect 6975 1666 6994 1692
rect 7058 1688 7089 1700
rect 7104 1688 7207 1700
rect 7219 1690 7245 1716
rect 7260 1711 7290 1722
rect 7322 1718 7384 1734
rect 7322 1716 7368 1718
rect 7322 1700 7384 1716
rect 7396 1700 7402 1748
rect 7405 1740 7485 1748
rect 7405 1738 7424 1740
rect 7439 1738 7473 1740
rect 7405 1722 7485 1738
rect 7405 1700 7424 1722
rect 7439 1706 7469 1722
rect 7497 1716 7503 1790
rect 7506 1716 7525 1860
rect 7540 1716 7546 1860
rect 7555 1790 7568 1860
rect 7620 1856 7642 1860
rect 7613 1834 7642 1848
rect 7695 1834 7711 1848
rect 7749 1844 7755 1846
rect 7762 1844 7870 1860
rect 7877 1844 7883 1846
rect 7891 1844 7906 1860
rect 7972 1854 7991 1857
rect 7613 1832 7711 1834
rect 7738 1832 7906 1844
rect 7921 1834 7937 1848
rect 7972 1835 7994 1854
rect 8004 1848 8020 1849
rect 8003 1846 8020 1848
rect 8004 1841 8020 1846
rect 7994 1834 8000 1835
rect 8003 1834 8032 1841
rect 7921 1833 8032 1834
rect 7921 1832 8038 1833
rect 7597 1824 7648 1832
rect 7695 1824 7729 1832
rect 7597 1812 7622 1824
rect 7629 1812 7648 1824
rect 7702 1822 7729 1824
rect 7738 1822 7959 1832
rect 7994 1829 8000 1832
rect 7702 1818 7959 1822
rect 7597 1804 7648 1812
rect 7695 1804 7959 1818
rect 8003 1824 8038 1832
rect 7549 1756 7568 1790
rect 7613 1796 7642 1804
rect 7613 1790 7630 1796
rect 7613 1788 7647 1790
rect 7695 1788 7711 1804
rect 7712 1794 7920 1804
rect 7921 1794 7937 1804
rect 7985 1800 8000 1815
rect 8003 1812 8004 1824
rect 8011 1812 8038 1824
rect 8003 1804 8038 1812
rect 8003 1803 8032 1804
rect 7723 1790 7937 1794
rect 7738 1788 7937 1790
rect 7972 1790 7985 1800
rect 8003 1790 8020 1803
rect 7972 1788 8020 1790
rect 7614 1784 7647 1788
rect 7610 1782 7647 1784
rect 7610 1781 7677 1782
rect 7610 1776 7641 1781
rect 7647 1776 7677 1781
rect 7610 1772 7677 1776
rect 7583 1769 7677 1772
rect 7583 1762 7632 1769
rect 7583 1756 7613 1762
rect 7632 1757 7637 1762
rect 7549 1740 7629 1756
rect 7641 1748 7677 1769
rect 7738 1764 7927 1788
rect 7972 1787 8019 1788
rect 7985 1782 8019 1787
rect 7753 1761 7927 1764
rect 7746 1758 7927 1761
rect 7955 1781 8019 1782
rect 7549 1738 7568 1740
rect 7583 1738 7617 1740
rect 7549 1722 7629 1738
rect 7549 1716 7568 1722
rect 7265 1690 7368 1700
rect 7219 1688 7368 1690
rect 7389 1688 7424 1700
rect 7058 1686 7220 1688
rect 7070 1666 7089 1686
rect 7104 1684 7134 1686
rect 6953 1658 6994 1666
rect 7076 1662 7089 1666
rect 7141 1670 7220 1686
rect 7252 1686 7424 1688
rect 7252 1670 7331 1686
rect 7338 1684 7368 1686
rect 6916 1648 6945 1658
rect 6959 1648 6988 1658
rect 7003 1648 7033 1662
rect 7076 1648 7119 1662
rect 7141 1658 7331 1670
rect 7396 1666 7402 1686
rect 7126 1648 7156 1658
rect 7157 1648 7315 1658
rect 7319 1648 7349 1658
rect 7353 1648 7383 1662
rect 7411 1648 7424 1686
rect 7496 1700 7525 1716
rect 7539 1700 7568 1716
rect 7583 1706 7613 1722
rect 7641 1700 7647 1748
rect 7650 1742 7669 1748
rect 7684 1742 7714 1750
rect 7650 1734 7714 1742
rect 7650 1718 7730 1734
rect 7746 1727 7808 1758
rect 7824 1727 7886 1758
rect 7955 1756 8004 1781
rect 8019 1756 8049 1772
rect 7918 1742 7948 1750
rect 7955 1748 8065 1756
rect 7918 1734 7963 1742
rect 7650 1716 7669 1718
rect 7684 1716 7730 1718
rect 7650 1700 7730 1716
rect 7757 1714 7792 1727
rect 7833 1724 7870 1727
rect 7833 1722 7875 1724
rect 7762 1711 7792 1714
rect 7771 1707 7778 1711
rect 7778 1706 7779 1707
rect 7737 1700 7747 1706
rect 7496 1692 7531 1700
rect 7496 1666 7497 1692
rect 7504 1666 7531 1692
rect 7439 1648 7469 1662
rect 7496 1658 7531 1666
rect 7533 1692 7574 1700
rect 7533 1666 7548 1692
rect 7555 1666 7574 1692
rect 7638 1688 7669 1700
rect 7684 1688 7787 1700
rect 7799 1690 7825 1716
rect 7840 1711 7870 1722
rect 7902 1718 7964 1734
rect 7902 1716 7948 1718
rect 7902 1700 7964 1716
rect 7976 1700 7982 1748
rect 7985 1740 8065 1748
rect 7985 1738 8004 1740
rect 8019 1738 8053 1740
rect 7985 1722 8065 1738
rect 7985 1700 8004 1722
rect 8019 1706 8049 1722
rect 8077 1716 8083 1790
rect 8086 1716 8105 1860
rect 8120 1716 8126 1860
rect 8135 1790 8148 1860
rect 8200 1856 8222 1860
rect 8193 1834 8222 1848
rect 8275 1834 8291 1848
rect 8329 1844 8335 1846
rect 8342 1844 8450 1860
rect 8457 1844 8463 1846
rect 8471 1844 8486 1860
rect 8552 1854 8571 1857
rect 8193 1832 8291 1834
rect 8318 1832 8486 1844
rect 8501 1834 8517 1848
rect 8552 1835 8574 1854
rect 8584 1848 8600 1849
rect 8583 1846 8600 1848
rect 8584 1841 8600 1846
rect 8574 1834 8580 1835
rect 8583 1834 8612 1841
rect 8501 1833 8612 1834
rect 8501 1832 8618 1833
rect 8177 1824 8228 1832
rect 8275 1824 8309 1832
rect 8177 1812 8202 1824
rect 8209 1812 8228 1824
rect 8282 1822 8309 1824
rect 8318 1822 8539 1832
rect 8574 1829 8580 1832
rect 8282 1818 8539 1822
rect 8177 1804 8228 1812
rect 8275 1804 8539 1818
rect 8583 1824 8618 1832
rect 8129 1756 8148 1790
rect 8193 1796 8222 1804
rect 8193 1790 8210 1796
rect 8193 1788 8227 1790
rect 8275 1788 8291 1804
rect 8292 1794 8500 1804
rect 8501 1794 8517 1804
rect 8565 1800 8580 1815
rect 8583 1812 8584 1824
rect 8591 1812 8618 1824
rect 8583 1804 8618 1812
rect 8583 1803 8612 1804
rect 8303 1790 8517 1794
rect 8318 1788 8517 1790
rect 8552 1790 8565 1800
rect 8583 1790 8600 1803
rect 8552 1788 8600 1790
rect 8194 1784 8227 1788
rect 8190 1782 8227 1784
rect 8190 1781 8257 1782
rect 8190 1776 8221 1781
rect 8227 1776 8257 1781
rect 8190 1772 8257 1776
rect 8163 1769 8257 1772
rect 8163 1762 8212 1769
rect 8163 1756 8193 1762
rect 8212 1757 8217 1762
rect 8129 1740 8209 1756
rect 8221 1748 8257 1769
rect 8318 1764 8507 1788
rect 8552 1787 8599 1788
rect 8565 1782 8599 1787
rect 8333 1761 8507 1764
rect 8326 1758 8507 1761
rect 8535 1781 8599 1782
rect 8129 1738 8148 1740
rect 8163 1738 8197 1740
rect 8129 1722 8209 1738
rect 8129 1716 8148 1722
rect 7845 1690 7948 1700
rect 7799 1688 7948 1690
rect 7969 1688 8004 1700
rect 7638 1686 7800 1688
rect 7650 1666 7669 1686
rect 7684 1684 7714 1686
rect 7533 1658 7574 1666
rect 7656 1662 7669 1666
rect 7721 1670 7800 1686
rect 7832 1686 8004 1688
rect 7832 1670 7911 1686
rect 7918 1684 7948 1686
rect 7496 1648 7525 1658
rect 7539 1648 7568 1658
rect 7583 1648 7613 1662
rect 7656 1648 7699 1662
rect 7721 1658 7911 1670
rect 7976 1666 7982 1686
rect 7706 1648 7736 1658
rect 7737 1648 7895 1658
rect 7899 1648 7929 1658
rect 7933 1648 7963 1662
rect 7991 1648 8004 1686
rect 8076 1700 8105 1716
rect 8119 1700 8148 1716
rect 8163 1706 8193 1722
rect 8221 1700 8227 1748
rect 8230 1742 8249 1748
rect 8264 1742 8294 1750
rect 8230 1734 8294 1742
rect 8230 1718 8310 1734
rect 8326 1727 8388 1758
rect 8404 1727 8466 1758
rect 8535 1756 8584 1781
rect 8599 1756 8629 1772
rect 8498 1742 8528 1750
rect 8535 1748 8645 1756
rect 8498 1734 8543 1742
rect 8230 1716 8249 1718
rect 8264 1716 8310 1718
rect 8230 1700 8310 1716
rect 8337 1714 8372 1727
rect 8413 1724 8450 1727
rect 8413 1722 8455 1724
rect 8342 1711 8372 1714
rect 8351 1707 8358 1711
rect 8358 1706 8359 1707
rect 8317 1700 8327 1706
rect 8076 1692 8111 1700
rect 8076 1666 8077 1692
rect 8084 1666 8111 1692
rect 8019 1648 8049 1662
rect 8076 1658 8111 1666
rect 8113 1692 8154 1700
rect 8113 1666 8128 1692
rect 8135 1666 8154 1692
rect 8218 1688 8249 1700
rect 8264 1688 8367 1700
rect 8379 1690 8405 1716
rect 8420 1711 8450 1722
rect 8482 1718 8544 1734
rect 8482 1716 8528 1718
rect 8482 1700 8544 1716
rect 8556 1700 8562 1748
rect 8565 1740 8645 1748
rect 8565 1738 8584 1740
rect 8599 1738 8633 1740
rect 8565 1722 8645 1738
rect 8565 1700 8584 1722
rect 8599 1706 8629 1722
rect 8657 1716 8663 1790
rect 8666 1716 8685 1860
rect 8700 1716 8706 1860
rect 8715 1790 8728 1860
rect 8780 1856 8802 1860
rect 8773 1834 8802 1848
rect 8855 1834 8871 1848
rect 8909 1844 8915 1846
rect 8922 1844 9030 1860
rect 9037 1844 9043 1846
rect 9051 1844 9066 1860
rect 9132 1854 9151 1857
rect 8773 1832 8871 1834
rect 8898 1832 9066 1844
rect 9081 1834 9097 1848
rect 9132 1835 9154 1854
rect 9164 1848 9180 1849
rect 9163 1846 9180 1848
rect 9164 1841 9180 1846
rect 9154 1834 9160 1835
rect 9163 1834 9192 1841
rect 9081 1833 9192 1834
rect 9081 1832 9198 1833
rect 8757 1824 8808 1832
rect 8855 1824 8889 1832
rect 8757 1812 8782 1824
rect 8789 1812 8808 1824
rect 8862 1822 8889 1824
rect 8898 1822 9119 1832
rect 9154 1829 9160 1832
rect 8862 1818 9119 1822
rect 8757 1804 8808 1812
rect 8855 1804 9119 1818
rect 9163 1824 9198 1832
rect 8709 1756 8728 1790
rect 8773 1796 8802 1804
rect 8773 1790 8790 1796
rect 8773 1788 8807 1790
rect 8855 1788 8871 1804
rect 8872 1794 9080 1804
rect 9081 1794 9097 1804
rect 9145 1800 9160 1815
rect 9163 1812 9164 1824
rect 9171 1812 9198 1824
rect 9163 1804 9198 1812
rect 9163 1803 9192 1804
rect 8883 1790 9097 1794
rect 8898 1788 9097 1790
rect 9132 1790 9145 1800
rect 9163 1790 9180 1803
rect 9132 1788 9180 1790
rect 8774 1784 8807 1788
rect 8770 1782 8807 1784
rect 8770 1781 8837 1782
rect 8770 1776 8801 1781
rect 8807 1776 8837 1781
rect 8770 1772 8837 1776
rect 8743 1769 8837 1772
rect 8743 1762 8792 1769
rect 8743 1756 8773 1762
rect 8792 1757 8797 1762
rect 8709 1740 8789 1756
rect 8801 1748 8837 1769
rect 8898 1764 9087 1788
rect 9132 1787 9179 1788
rect 9145 1782 9179 1787
rect 8913 1761 9087 1764
rect 8906 1758 9087 1761
rect 9115 1781 9179 1782
rect 8709 1738 8728 1740
rect 8743 1738 8777 1740
rect 8709 1722 8789 1738
rect 8709 1716 8728 1722
rect 8425 1690 8528 1700
rect 8379 1688 8528 1690
rect 8549 1688 8584 1700
rect 8218 1686 8380 1688
rect 8230 1666 8249 1686
rect 8264 1684 8294 1686
rect 8113 1658 8154 1666
rect 8236 1662 8249 1666
rect 8301 1670 8380 1686
rect 8412 1686 8584 1688
rect 8412 1670 8491 1686
rect 8498 1684 8528 1686
rect 8076 1648 8105 1658
rect 8119 1648 8148 1658
rect 8163 1648 8193 1662
rect 8236 1648 8279 1662
rect 8301 1658 8491 1670
rect 8556 1666 8562 1686
rect 8286 1648 8316 1658
rect 8317 1648 8475 1658
rect 8479 1648 8509 1658
rect 8513 1648 8543 1662
rect 8571 1648 8584 1686
rect 8656 1700 8685 1716
rect 8699 1700 8728 1716
rect 8743 1706 8773 1722
rect 8801 1700 8807 1748
rect 8810 1742 8829 1748
rect 8844 1742 8874 1750
rect 8810 1734 8874 1742
rect 8810 1718 8890 1734
rect 8906 1727 8968 1758
rect 8984 1727 9046 1758
rect 9115 1756 9164 1781
rect 9179 1756 9209 1772
rect 9078 1742 9108 1750
rect 9115 1748 9225 1756
rect 9078 1734 9123 1742
rect 8810 1716 8829 1718
rect 8844 1716 8890 1718
rect 8810 1700 8890 1716
rect 8917 1714 8952 1727
rect 8993 1724 9030 1727
rect 8993 1722 9035 1724
rect 8922 1711 8952 1714
rect 8931 1707 8938 1711
rect 8938 1706 8939 1707
rect 8897 1700 8907 1706
rect 8656 1692 8691 1700
rect 8656 1666 8657 1692
rect 8664 1666 8691 1692
rect 8599 1648 8629 1662
rect 8656 1658 8691 1666
rect 8693 1692 8734 1700
rect 8693 1666 8708 1692
rect 8715 1666 8734 1692
rect 8798 1688 8829 1700
rect 8844 1688 8947 1700
rect 8959 1690 8985 1716
rect 9000 1711 9030 1722
rect 9062 1718 9124 1734
rect 9062 1716 9108 1718
rect 9062 1700 9124 1716
rect 9136 1700 9142 1748
rect 9145 1740 9225 1748
rect 9145 1738 9164 1740
rect 9179 1738 9213 1740
rect 9145 1722 9225 1738
rect 9145 1700 9164 1722
rect 9179 1706 9209 1722
rect 9237 1716 9243 1790
rect 9252 1716 9265 1860
rect 9005 1690 9108 1700
rect 8959 1688 9108 1690
rect 9129 1688 9164 1700
rect 8798 1686 8960 1688
rect 8810 1666 8829 1686
rect 8844 1684 8874 1686
rect 8693 1658 8734 1666
rect 8816 1662 8829 1666
rect 8881 1670 8960 1686
rect 8992 1686 9164 1688
rect 8992 1670 9071 1686
rect 9078 1684 9108 1686
rect 8656 1648 8685 1658
rect 8699 1648 8728 1658
rect 8743 1648 8773 1662
rect 8816 1648 8859 1662
rect 8881 1658 9071 1670
rect 9136 1666 9142 1686
rect 8866 1648 8896 1658
rect 8897 1648 9055 1658
rect 9059 1648 9089 1658
rect 9093 1648 9123 1662
rect 9151 1648 9164 1686
rect 9236 1700 9265 1716
rect 9236 1692 9271 1700
rect 9236 1666 9237 1692
rect 9244 1666 9271 1692
rect 9179 1648 9209 1662
rect 9236 1658 9271 1666
rect 9236 1648 9265 1658
rect -1 1642 9265 1648
rect 0 1634 9265 1642
rect 15 1604 28 1634
rect 43 1620 73 1634
rect 116 1620 159 1634
rect 166 1620 386 1634
rect 393 1620 423 1634
rect 83 1606 98 1618
rect 117 1606 130 1620
rect 198 1616 351 1620
rect 80 1604 102 1606
rect 180 1604 372 1616
rect 451 1604 464 1634
rect 479 1620 509 1634
rect 546 1604 565 1634
rect 580 1604 586 1634
rect 595 1604 608 1634
rect 623 1620 653 1634
rect 696 1620 739 1634
rect 746 1620 966 1634
rect 973 1620 1003 1634
rect 663 1606 678 1618
rect 697 1606 710 1620
rect 778 1616 931 1620
rect 660 1604 682 1606
rect 760 1604 952 1616
rect 1031 1604 1044 1634
rect 1059 1620 1089 1634
rect 1126 1604 1145 1634
rect 1160 1604 1166 1634
rect 1175 1604 1188 1634
rect 1203 1620 1233 1634
rect 1276 1620 1319 1634
rect 1326 1620 1546 1634
rect 1553 1620 1583 1634
rect 1243 1606 1258 1618
rect 1277 1606 1290 1620
rect 1358 1616 1511 1620
rect 1240 1604 1262 1606
rect 1340 1604 1532 1616
rect 1611 1604 1624 1634
rect 1639 1620 1669 1634
rect 1706 1604 1725 1634
rect 1740 1604 1746 1634
rect 1755 1604 1768 1634
rect 1783 1620 1813 1634
rect 1856 1620 1899 1634
rect 1906 1620 2126 1634
rect 2133 1620 2163 1634
rect 1823 1606 1838 1618
rect 1857 1606 1870 1620
rect 1938 1616 2091 1620
rect 1820 1604 1842 1606
rect 1920 1604 2112 1616
rect 2191 1604 2204 1634
rect 2219 1620 2249 1634
rect 2286 1604 2305 1634
rect 2320 1604 2326 1634
rect 2335 1604 2348 1634
rect 2363 1620 2393 1634
rect 2436 1620 2479 1634
rect 2486 1620 2706 1634
rect 2713 1620 2743 1634
rect 2403 1606 2418 1618
rect 2437 1606 2450 1620
rect 2518 1616 2671 1620
rect 2400 1604 2422 1606
rect 2500 1604 2692 1616
rect 2771 1604 2784 1634
rect 2799 1620 2829 1634
rect 2866 1604 2885 1634
rect 2900 1604 2906 1634
rect 2915 1604 2928 1634
rect 2943 1620 2973 1634
rect 3016 1620 3059 1634
rect 3066 1620 3286 1634
rect 3293 1620 3323 1634
rect 2983 1606 2998 1618
rect 3017 1606 3030 1620
rect 3098 1616 3251 1620
rect 2980 1604 3002 1606
rect 3080 1604 3272 1616
rect 3351 1604 3364 1634
rect 3379 1620 3409 1634
rect 3446 1604 3465 1634
rect 3480 1604 3486 1634
rect 3495 1604 3508 1634
rect 3523 1620 3553 1634
rect 3596 1620 3639 1634
rect 3646 1620 3866 1634
rect 3873 1620 3903 1634
rect 3563 1606 3578 1618
rect 3597 1606 3610 1620
rect 3678 1616 3831 1620
rect 3560 1604 3582 1606
rect 3660 1604 3852 1616
rect 3931 1604 3944 1634
rect 3959 1620 3989 1634
rect 4026 1604 4045 1634
rect 4060 1604 4066 1634
rect 4075 1604 4088 1634
rect 4103 1620 4133 1634
rect 4176 1620 4219 1634
rect 4226 1620 4446 1634
rect 4453 1620 4483 1634
rect 4143 1606 4158 1618
rect 4177 1606 4190 1620
rect 4258 1616 4411 1620
rect 4140 1604 4162 1606
rect 4240 1604 4432 1616
rect 4511 1604 4524 1634
rect 4539 1620 4569 1634
rect 4606 1604 4625 1634
rect 4640 1604 4646 1634
rect 4655 1604 4668 1634
rect 4683 1620 4713 1634
rect 4756 1620 4799 1634
rect 4806 1620 5026 1634
rect 5033 1620 5063 1634
rect 4723 1606 4738 1618
rect 4757 1606 4770 1620
rect 4838 1616 4991 1620
rect 4720 1604 4742 1606
rect 4820 1604 5012 1616
rect 5091 1604 5104 1634
rect 5119 1620 5149 1634
rect 5186 1604 5205 1634
rect 5220 1604 5226 1634
rect 5235 1604 5248 1634
rect 5263 1620 5293 1634
rect 5336 1620 5379 1634
rect 5386 1620 5606 1634
rect 5613 1620 5643 1634
rect 5303 1606 5318 1618
rect 5337 1606 5350 1620
rect 5418 1616 5571 1620
rect 5300 1604 5322 1606
rect 5400 1604 5592 1616
rect 5671 1604 5684 1634
rect 5699 1620 5729 1634
rect 5766 1604 5785 1634
rect 5800 1604 5806 1634
rect 5815 1604 5828 1634
rect 5843 1620 5873 1634
rect 5916 1620 5959 1634
rect 5966 1620 6186 1634
rect 6193 1620 6223 1634
rect 5883 1606 5898 1618
rect 5917 1606 5930 1620
rect 5998 1616 6151 1620
rect 5880 1604 5902 1606
rect 5980 1604 6172 1616
rect 6251 1604 6264 1634
rect 6279 1620 6309 1634
rect 6346 1604 6365 1634
rect 6380 1604 6386 1634
rect 6395 1604 6408 1634
rect 6423 1620 6453 1634
rect 6496 1620 6539 1634
rect 6546 1620 6766 1634
rect 6773 1620 6803 1634
rect 6463 1606 6478 1618
rect 6497 1606 6510 1620
rect 6578 1616 6731 1620
rect 6460 1604 6482 1606
rect 6560 1604 6752 1616
rect 6831 1604 6844 1634
rect 6859 1620 6889 1634
rect 6926 1604 6945 1634
rect 6960 1604 6966 1634
rect 6975 1604 6988 1634
rect 7003 1620 7033 1634
rect 7076 1620 7119 1634
rect 7126 1620 7346 1634
rect 7353 1620 7383 1634
rect 7043 1606 7058 1618
rect 7077 1606 7090 1620
rect 7158 1616 7311 1620
rect 7040 1604 7062 1606
rect 7140 1604 7332 1616
rect 7411 1604 7424 1634
rect 7439 1620 7469 1634
rect 7506 1604 7525 1634
rect 7540 1604 7546 1634
rect 7555 1604 7568 1634
rect 7583 1620 7613 1634
rect 7656 1620 7699 1634
rect 7706 1620 7926 1634
rect 7933 1620 7963 1634
rect 7623 1606 7638 1618
rect 7657 1606 7670 1620
rect 7738 1616 7891 1620
rect 7620 1604 7642 1606
rect 7720 1604 7912 1616
rect 7991 1604 8004 1634
rect 8019 1620 8049 1634
rect 8086 1604 8105 1634
rect 8120 1604 8126 1634
rect 8135 1604 8148 1634
rect 8163 1620 8193 1634
rect 8236 1620 8279 1634
rect 8286 1620 8506 1634
rect 8513 1620 8543 1634
rect 8203 1606 8218 1618
rect 8237 1606 8250 1620
rect 8318 1616 8471 1620
rect 8200 1604 8222 1606
rect 8300 1604 8492 1616
rect 8571 1604 8584 1634
rect 8599 1620 8629 1634
rect 8666 1604 8685 1634
rect 8700 1604 8706 1634
rect 8715 1604 8728 1634
rect 8743 1620 8773 1634
rect 8816 1620 8859 1634
rect 8866 1620 9086 1634
rect 9093 1620 9123 1634
rect 8783 1606 8798 1618
rect 8817 1606 8830 1620
rect 8898 1616 9051 1620
rect 8780 1604 8802 1606
rect 8880 1604 9072 1616
rect 9151 1604 9164 1634
rect 9179 1620 9209 1634
rect 9252 1604 9265 1634
rect 0 1590 9265 1604
rect 15 1520 28 1590
rect 80 1586 102 1590
rect 73 1564 102 1578
rect 155 1564 171 1578
rect 209 1574 215 1576
rect 222 1574 330 1590
rect 337 1574 343 1576
rect 351 1574 366 1590
rect 432 1584 451 1587
rect 73 1562 171 1564
rect 198 1562 366 1574
rect 381 1564 397 1578
rect 432 1565 454 1584
rect 464 1578 480 1579
rect 463 1576 480 1578
rect 464 1571 480 1576
rect 454 1564 460 1565
rect 463 1564 492 1571
rect 381 1563 492 1564
rect 381 1562 498 1563
rect 57 1554 108 1562
rect 155 1554 189 1562
rect 57 1542 82 1554
rect 89 1542 108 1554
rect 162 1552 189 1554
rect 198 1552 419 1562
rect 454 1559 460 1562
rect 162 1548 419 1552
rect 57 1534 108 1542
rect 155 1534 419 1548
rect 463 1554 498 1562
rect 9 1486 28 1520
rect 73 1526 102 1534
rect 73 1520 90 1526
rect 73 1518 107 1520
rect 155 1518 171 1534
rect 172 1524 380 1534
rect 381 1524 397 1534
rect 445 1530 460 1545
rect 463 1542 464 1554
rect 471 1542 498 1554
rect 463 1534 498 1542
rect 463 1533 492 1534
rect 183 1520 397 1524
rect 198 1518 397 1520
rect 432 1520 445 1530
rect 463 1520 480 1533
rect 432 1518 480 1520
rect 74 1514 107 1518
rect 70 1512 107 1514
rect 70 1511 137 1512
rect 70 1506 101 1511
rect 107 1506 137 1511
rect 70 1502 137 1506
rect 43 1499 137 1502
rect 43 1492 92 1499
rect 43 1486 73 1492
rect 92 1487 97 1492
rect 9 1470 89 1486
rect 101 1478 137 1499
rect 198 1494 387 1518
rect 432 1517 479 1518
rect 445 1512 479 1517
rect 213 1491 387 1494
rect 206 1488 387 1491
rect 415 1511 479 1512
rect 9 1468 28 1470
rect 43 1468 77 1470
rect 9 1452 89 1468
rect 9 1446 28 1452
rect -1 1430 28 1446
rect 43 1436 73 1452
rect 101 1430 107 1478
rect 110 1472 129 1478
rect 144 1472 174 1480
rect 110 1464 174 1472
rect 110 1448 190 1464
rect 206 1457 268 1488
rect 284 1457 346 1488
rect 415 1486 464 1511
rect 479 1486 509 1502
rect 378 1472 408 1480
rect 415 1478 525 1486
rect 378 1464 423 1472
rect 110 1446 129 1448
rect 144 1446 190 1448
rect 110 1430 190 1446
rect 217 1444 252 1457
rect 293 1454 330 1457
rect 293 1452 335 1454
rect 222 1441 252 1444
rect 231 1437 238 1441
rect 238 1436 239 1437
rect 197 1430 207 1436
rect -7 1422 34 1430
rect -7 1396 8 1422
rect 15 1396 34 1422
rect 98 1418 129 1430
rect 144 1418 247 1430
rect 259 1420 285 1446
rect 300 1441 330 1452
rect 362 1448 424 1464
rect 362 1446 408 1448
rect 362 1430 424 1446
rect 436 1430 442 1478
rect 445 1470 525 1478
rect 445 1468 464 1470
rect 479 1468 513 1470
rect 445 1452 525 1468
rect 445 1430 464 1452
rect 479 1436 509 1452
rect 537 1446 543 1520
rect 546 1446 565 1590
rect 580 1446 586 1590
rect 595 1520 608 1590
rect 660 1586 682 1590
rect 653 1564 682 1578
rect 735 1564 751 1578
rect 789 1574 795 1576
rect 802 1574 910 1590
rect 917 1574 923 1576
rect 931 1574 946 1590
rect 1012 1584 1031 1587
rect 653 1562 751 1564
rect 778 1562 946 1574
rect 961 1564 977 1578
rect 1012 1565 1034 1584
rect 1044 1578 1060 1579
rect 1043 1576 1060 1578
rect 1044 1571 1060 1576
rect 1034 1564 1040 1565
rect 1043 1564 1072 1571
rect 961 1563 1072 1564
rect 961 1562 1078 1563
rect 637 1554 688 1562
rect 735 1554 769 1562
rect 637 1542 662 1554
rect 669 1542 688 1554
rect 742 1552 769 1554
rect 778 1552 999 1562
rect 1034 1559 1040 1562
rect 742 1548 999 1552
rect 637 1534 688 1542
rect 735 1534 999 1548
rect 1043 1554 1078 1562
rect 589 1486 608 1520
rect 653 1526 682 1534
rect 653 1520 670 1526
rect 653 1518 687 1520
rect 735 1518 751 1534
rect 752 1524 960 1534
rect 961 1524 977 1534
rect 1025 1530 1040 1545
rect 1043 1542 1044 1554
rect 1051 1542 1078 1554
rect 1043 1534 1078 1542
rect 1043 1533 1072 1534
rect 763 1520 977 1524
rect 778 1518 977 1520
rect 1012 1520 1025 1530
rect 1043 1520 1060 1533
rect 1012 1518 1060 1520
rect 654 1514 687 1518
rect 650 1512 687 1514
rect 650 1511 717 1512
rect 650 1506 681 1511
rect 687 1506 717 1511
rect 650 1502 717 1506
rect 623 1499 717 1502
rect 623 1492 672 1499
rect 623 1486 653 1492
rect 672 1487 677 1492
rect 589 1470 669 1486
rect 681 1478 717 1499
rect 778 1494 967 1518
rect 1012 1517 1059 1518
rect 1025 1512 1059 1517
rect 793 1491 967 1494
rect 786 1488 967 1491
rect 995 1511 1059 1512
rect 589 1468 608 1470
rect 623 1468 657 1470
rect 589 1452 669 1468
rect 589 1446 608 1452
rect 305 1420 408 1430
rect 259 1418 408 1420
rect 429 1418 464 1430
rect 98 1416 260 1418
rect 110 1396 129 1416
rect 144 1414 174 1416
rect -7 1388 34 1396
rect 116 1392 129 1396
rect 181 1400 260 1416
rect 292 1416 464 1418
rect 292 1400 371 1416
rect 378 1414 408 1416
rect -1 1378 28 1388
rect 43 1378 73 1392
rect 116 1378 159 1392
rect 181 1388 371 1400
rect 436 1396 442 1416
rect 166 1378 196 1388
rect 197 1378 355 1388
rect 359 1378 389 1388
rect 393 1378 423 1392
rect 451 1378 464 1416
rect 536 1430 565 1446
rect 579 1430 608 1446
rect 623 1436 653 1452
rect 681 1430 687 1478
rect 690 1472 709 1478
rect 724 1472 754 1480
rect 690 1464 754 1472
rect 690 1448 770 1464
rect 786 1457 848 1488
rect 864 1457 926 1488
rect 995 1486 1044 1511
rect 1059 1486 1089 1502
rect 958 1472 988 1480
rect 995 1478 1105 1486
rect 958 1464 1003 1472
rect 690 1446 709 1448
rect 724 1446 770 1448
rect 690 1430 770 1446
rect 797 1444 832 1457
rect 873 1454 910 1457
rect 873 1452 915 1454
rect 802 1441 832 1444
rect 811 1437 818 1441
rect 818 1436 819 1437
rect 777 1430 787 1436
rect 536 1422 571 1430
rect 536 1396 537 1422
rect 544 1396 571 1422
rect 479 1378 509 1392
rect 536 1388 571 1396
rect 573 1422 614 1430
rect 573 1396 588 1422
rect 595 1396 614 1422
rect 678 1418 709 1430
rect 724 1418 827 1430
rect 839 1420 865 1446
rect 880 1441 910 1452
rect 942 1448 1004 1464
rect 942 1446 988 1448
rect 942 1430 1004 1446
rect 1016 1430 1022 1478
rect 1025 1470 1105 1478
rect 1025 1468 1044 1470
rect 1059 1468 1093 1470
rect 1025 1452 1105 1468
rect 1025 1430 1044 1452
rect 1059 1436 1089 1452
rect 1117 1446 1123 1520
rect 1126 1446 1145 1590
rect 1160 1446 1166 1590
rect 1175 1520 1188 1590
rect 1240 1586 1262 1590
rect 1233 1564 1262 1578
rect 1315 1564 1331 1578
rect 1369 1574 1375 1576
rect 1382 1574 1490 1590
rect 1497 1574 1503 1576
rect 1511 1574 1526 1590
rect 1592 1584 1611 1587
rect 1233 1562 1331 1564
rect 1358 1562 1526 1574
rect 1541 1564 1557 1578
rect 1592 1565 1614 1584
rect 1624 1578 1640 1579
rect 1623 1576 1640 1578
rect 1624 1571 1640 1576
rect 1614 1564 1620 1565
rect 1623 1564 1652 1571
rect 1541 1563 1652 1564
rect 1541 1562 1658 1563
rect 1217 1554 1268 1562
rect 1315 1554 1349 1562
rect 1217 1542 1242 1554
rect 1249 1542 1268 1554
rect 1322 1552 1349 1554
rect 1358 1552 1579 1562
rect 1614 1559 1620 1562
rect 1322 1548 1579 1552
rect 1217 1534 1268 1542
rect 1315 1534 1579 1548
rect 1623 1554 1658 1562
rect 1169 1486 1188 1520
rect 1233 1526 1262 1534
rect 1233 1520 1250 1526
rect 1233 1518 1267 1520
rect 1315 1518 1331 1534
rect 1332 1524 1540 1534
rect 1541 1524 1557 1534
rect 1605 1530 1620 1545
rect 1623 1542 1624 1554
rect 1631 1542 1658 1554
rect 1623 1534 1658 1542
rect 1623 1533 1652 1534
rect 1343 1520 1557 1524
rect 1358 1518 1557 1520
rect 1592 1520 1605 1530
rect 1623 1520 1640 1533
rect 1592 1518 1640 1520
rect 1234 1514 1267 1518
rect 1230 1512 1267 1514
rect 1230 1511 1297 1512
rect 1230 1506 1261 1511
rect 1267 1506 1297 1511
rect 1230 1502 1297 1506
rect 1203 1499 1297 1502
rect 1203 1492 1252 1499
rect 1203 1486 1233 1492
rect 1252 1487 1257 1492
rect 1169 1470 1249 1486
rect 1261 1478 1297 1499
rect 1358 1494 1547 1518
rect 1592 1517 1639 1518
rect 1605 1512 1639 1517
rect 1373 1491 1547 1494
rect 1366 1488 1547 1491
rect 1575 1511 1639 1512
rect 1169 1468 1188 1470
rect 1203 1468 1237 1470
rect 1169 1452 1249 1468
rect 1169 1446 1188 1452
rect 885 1420 988 1430
rect 839 1418 988 1420
rect 1009 1418 1044 1430
rect 678 1416 840 1418
rect 690 1396 709 1416
rect 724 1414 754 1416
rect 573 1388 614 1396
rect 696 1392 709 1396
rect 761 1400 840 1416
rect 872 1416 1044 1418
rect 872 1400 951 1416
rect 958 1414 988 1416
rect 536 1378 565 1388
rect 579 1378 608 1388
rect 623 1378 653 1392
rect 696 1378 739 1392
rect 761 1388 951 1400
rect 1016 1396 1022 1416
rect 746 1378 776 1388
rect 777 1378 935 1388
rect 939 1378 969 1388
rect 973 1378 1003 1392
rect 1031 1378 1044 1416
rect 1116 1430 1145 1446
rect 1159 1430 1188 1446
rect 1203 1436 1233 1452
rect 1261 1430 1267 1478
rect 1270 1472 1289 1478
rect 1304 1472 1334 1480
rect 1270 1464 1334 1472
rect 1270 1448 1350 1464
rect 1366 1457 1428 1488
rect 1444 1457 1506 1488
rect 1575 1486 1624 1511
rect 1639 1486 1669 1502
rect 1538 1472 1568 1480
rect 1575 1478 1685 1486
rect 1538 1464 1583 1472
rect 1270 1446 1289 1448
rect 1304 1446 1350 1448
rect 1270 1430 1350 1446
rect 1377 1444 1412 1457
rect 1453 1454 1490 1457
rect 1453 1452 1495 1454
rect 1382 1441 1412 1444
rect 1391 1437 1398 1441
rect 1398 1436 1399 1437
rect 1357 1430 1367 1436
rect 1116 1422 1151 1430
rect 1116 1396 1117 1422
rect 1124 1396 1151 1422
rect 1059 1378 1089 1392
rect 1116 1388 1151 1396
rect 1153 1422 1194 1430
rect 1153 1396 1168 1422
rect 1175 1396 1194 1422
rect 1258 1418 1289 1430
rect 1304 1418 1407 1430
rect 1419 1420 1445 1446
rect 1460 1441 1490 1452
rect 1522 1448 1584 1464
rect 1522 1446 1568 1448
rect 1522 1430 1584 1446
rect 1596 1430 1602 1478
rect 1605 1470 1685 1478
rect 1605 1468 1624 1470
rect 1639 1468 1673 1470
rect 1605 1452 1685 1468
rect 1605 1430 1624 1452
rect 1639 1436 1669 1452
rect 1697 1446 1703 1520
rect 1706 1446 1725 1590
rect 1740 1446 1746 1590
rect 1755 1520 1768 1590
rect 1820 1586 1842 1590
rect 1813 1564 1842 1578
rect 1895 1564 1911 1578
rect 1949 1574 1955 1576
rect 1962 1574 2070 1590
rect 2077 1574 2083 1576
rect 2091 1574 2106 1590
rect 2172 1584 2191 1587
rect 1813 1562 1911 1564
rect 1938 1562 2106 1574
rect 2121 1564 2137 1578
rect 2172 1565 2194 1584
rect 2204 1578 2220 1579
rect 2203 1576 2220 1578
rect 2204 1571 2220 1576
rect 2194 1564 2200 1565
rect 2203 1564 2232 1571
rect 2121 1563 2232 1564
rect 2121 1562 2238 1563
rect 1797 1554 1848 1562
rect 1895 1554 1929 1562
rect 1797 1542 1822 1554
rect 1829 1542 1848 1554
rect 1902 1552 1929 1554
rect 1938 1552 2159 1562
rect 2194 1559 2200 1562
rect 1902 1548 2159 1552
rect 1797 1534 1848 1542
rect 1895 1534 2159 1548
rect 2203 1554 2238 1562
rect 1749 1486 1768 1520
rect 1813 1526 1842 1534
rect 1813 1520 1830 1526
rect 1813 1518 1847 1520
rect 1895 1518 1911 1534
rect 1912 1524 2120 1534
rect 2121 1524 2137 1534
rect 2185 1530 2200 1545
rect 2203 1542 2204 1554
rect 2211 1542 2238 1554
rect 2203 1534 2238 1542
rect 2203 1533 2232 1534
rect 1923 1520 2137 1524
rect 1938 1518 2137 1520
rect 2172 1520 2185 1530
rect 2203 1520 2220 1533
rect 2172 1518 2220 1520
rect 1814 1514 1847 1518
rect 1810 1512 1847 1514
rect 1810 1511 1877 1512
rect 1810 1506 1841 1511
rect 1847 1506 1877 1511
rect 1810 1502 1877 1506
rect 1783 1499 1877 1502
rect 1783 1492 1832 1499
rect 1783 1486 1813 1492
rect 1832 1487 1837 1492
rect 1749 1470 1829 1486
rect 1841 1478 1877 1499
rect 1938 1494 2127 1518
rect 2172 1517 2219 1518
rect 2185 1512 2219 1517
rect 1953 1491 2127 1494
rect 1946 1488 2127 1491
rect 2155 1511 2219 1512
rect 1749 1468 1768 1470
rect 1783 1468 1817 1470
rect 1749 1452 1829 1468
rect 1749 1446 1768 1452
rect 1465 1420 1568 1430
rect 1419 1418 1568 1420
rect 1589 1418 1624 1430
rect 1258 1416 1420 1418
rect 1270 1396 1289 1416
rect 1304 1414 1334 1416
rect 1153 1388 1194 1396
rect 1276 1392 1289 1396
rect 1341 1400 1420 1416
rect 1452 1416 1624 1418
rect 1452 1400 1531 1416
rect 1538 1414 1568 1416
rect 1116 1378 1145 1388
rect 1159 1378 1188 1388
rect 1203 1378 1233 1392
rect 1276 1378 1319 1392
rect 1341 1388 1531 1400
rect 1596 1396 1602 1416
rect 1326 1378 1356 1388
rect 1357 1378 1515 1388
rect 1519 1378 1549 1388
rect 1553 1378 1583 1392
rect 1611 1378 1624 1416
rect 1696 1430 1725 1446
rect 1739 1430 1768 1446
rect 1783 1436 1813 1452
rect 1841 1430 1847 1478
rect 1850 1472 1869 1478
rect 1884 1472 1914 1480
rect 1850 1464 1914 1472
rect 1850 1448 1930 1464
rect 1946 1457 2008 1488
rect 2024 1457 2086 1488
rect 2155 1486 2204 1511
rect 2219 1486 2249 1502
rect 2118 1472 2148 1480
rect 2155 1478 2265 1486
rect 2118 1464 2163 1472
rect 1850 1446 1869 1448
rect 1884 1446 1930 1448
rect 1850 1430 1930 1446
rect 1957 1444 1992 1457
rect 2033 1454 2070 1457
rect 2033 1452 2075 1454
rect 1962 1441 1992 1444
rect 1971 1437 1978 1441
rect 1978 1436 1979 1437
rect 1937 1430 1947 1436
rect 1696 1422 1731 1430
rect 1696 1396 1697 1422
rect 1704 1396 1731 1422
rect 1639 1378 1669 1392
rect 1696 1388 1731 1396
rect 1733 1422 1774 1430
rect 1733 1396 1748 1422
rect 1755 1396 1774 1422
rect 1838 1418 1869 1430
rect 1884 1418 1987 1430
rect 1999 1420 2025 1446
rect 2040 1441 2070 1452
rect 2102 1448 2164 1464
rect 2102 1446 2148 1448
rect 2102 1430 2164 1446
rect 2176 1430 2182 1478
rect 2185 1470 2265 1478
rect 2185 1468 2204 1470
rect 2219 1468 2253 1470
rect 2185 1452 2265 1468
rect 2185 1430 2204 1452
rect 2219 1436 2249 1452
rect 2277 1446 2283 1520
rect 2286 1446 2305 1590
rect 2320 1446 2326 1590
rect 2335 1520 2348 1590
rect 2400 1586 2422 1590
rect 2393 1564 2422 1578
rect 2475 1564 2491 1578
rect 2529 1574 2535 1576
rect 2542 1574 2650 1590
rect 2657 1574 2663 1576
rect 2671 1574 2686 1590
rect 2752 1584 2771 1587
rect 2393 1562 2491 1564
rect 2518 1562 2686 1574
rect 2701 1564 2717 1578
rect 2752 1565 2774 1584
rect 2784 1578 2800 1579
rect 2783 1576 2800 1578
rect 2784 1571 2800 1576
rect 2774 1564 2780 1565
rect 2783 1564 2812 1571
rect 2701 1563 2812 1564
rect 2701 1562 2818 1563
rect 2377 1554 2428 1562
rect 2475 1554 2509 1562
rect 2377 1542 2402 1554
rect 2409 1542 2428 1554
rect 2482 1552 2509 1554
rect 2518 1552 2739 1562
rect 2774 1559 2780 1562
rect 2482 1548 2739 1552
rect 2377 1534 2428 1542
rect 2475 1534 2739 1548
rect 2783 1554 2818 1562
rect 2329 1486 2348 1520
rect 2393 1526 2422 1534
rect 2393 1520 2410 1526
rect 2393 1518 2427 1520
rect 2475 1518 2491 1534
rect 2492 1524 2700 1534
rect 2701 1524 2717 1534
rect 2765 1530 2780 1545
rect 2783 1542 2784 1554
rect 2791 1542 2818 1554
rect 2783 1534 2818 1542
rect 2783 1533 2812 1534
rect 2503 1520 2717 1524
rect 2518 1518 2717 1520
rect 2752 1520 2765 1530
rect 2783 1520 2800 1533
rect 2752 1518 2800 1520
rect 2394 1514 2427 1518
rect 2390 1512 2427 1514
rect 2390 1511 2457 1512
rect 2390 1506 2421 1511
rect 2427 1506 2457 1511
rect 2390 1502 2457 1506
rect 2363 1499 2457 1502
rect 2363 1492 2412 1499
rect 2363 1486 2393 1492
rect 2412 1487 2417 1492
rect 2329 1470 2409 1486
rect 2421 1478 2457 1499
rect 2518 1494 2707 1518
rect 2752 1517 2799 1518
rect 2765 1512 2799 1517
rect 2533 1491 2707 1494
rect 2526 1488 2707 1491
rect 2735 1511 2799 1512
rect 2329 1468 2348 1470
rect 2363 1468 2397 1470
rect 2329 1452 2409 1468
rect 2329 1446 2348 1452
rect 2045 1420 2148 1430
rect 1999 1418 2148 1420
rect 2169 1418 2204 1430
rect 1838 1416 2000 1418
rect 1850 1396 1869 1416
rect 1884 1414 1914 1416
rect 1733 1388 1774 1396
rect 1856 1392 1869 1396
rect 1921 1400 2000 1416
rect 2032 1416 2204 1418
rect 2032 1400 2111 1416
rect 2118 1414 2148 1416
rect 1696 1378 1725 1388
rect 1739 1378 1768 1388
rect 1783 1378 1813 1392
rect 1856 1378 1899 1392
rect 1921 1388 2111 1400
rect 2176 1396 2182 1416
rect 1906 1378 1936 1388
rect 1937 1378 2095 1388
rect 2099 1378 2129 1388
rect 2133 1378 2163 1392
rect 2191 1378 2204 1416
rect 2276 1430 2305 1446
rect 2319 1430 2348 1446
rect 2363 1436 2393 1452
rect 2421 1430 2427 1478
rect 2430 1472 2449 1478
rect 2464 1472 2494 1480
rect 2430 1464 2494 1472
rect 2430 1448 2510 1464
rect 2526 1457 2588 1488
rect 2604 1457 2666 1488
rect 2735 1486 2784 1511
rect 2799 1486 2829 1502
rect 2698 1472 2728 1480
rect 2735 1478 2845 1486
rect 2698 1464 2743 1472
rect 2430 1446 2449 1448
rect 2464 1446 2510 1448
rect 2430 1430 2510 1446
rect 2537 1444 2572 1457
rect 2613 1454 2650 1457
rect 2613 1452 2655 1454
rect 2542 1441 2572 1444
rect 2551 1437 2558 1441
rect 2558 1436 2559 1437
rect 2517 1430 2527 1436
rect 2276 1422 2311 1430
rect 2276 1396 2277 1422
rect 2284 1396 2311 1422
rect 2219 1378 2249 1392
rect 2276 1388 2311 1396
rect 2313 1422 2354 1430
rect 2313 1396 2328 1422
rect 2335 1396 2354 1422
rect 2418 1418 2449 1430
rect 2464 1418 2567 1430
rect 2579 1420 2605 1446
rect 2620 1441 2650 1452
rect 2682 1448 2744 1464
rect 2682 1446 2728 1448
rect 2682 1430 2744 1446
rect 2756 1430 2762 1478
rect 2765 1470 2845 1478
rect 2765 1468 2784 1470
rect 2799 1468 2833 1470
rect 2765 1452 2845 1468
rect 2765 1430 2784 1452
rect 2799 1436 2829 1452
rect 2857 1446 2863 1520
rect 2866 1446 2885 1590
rect 2900 1446 2906 1590
rect 2915 1520 2928 1590
rect 2980 1586 3002 1590
rect 2973 1564 3002 1578
rect 3055 1564 3071 1578
rect 3109 1574 3115 1576
rect 3122 1574 3230 1590
rect 3237 1574 3243 1576
rect 3251 1574 3266 1590
rect 3332 1584 3351 1587
rect 2973 1562 3071 1564
rect 3098 1562 3266 1574
rect 3281 1564 3297 1578
rect 3332 1565 3354 1584
rect 3364 1578 3380 1579
rect 3363 1576 3380 1578
rect 3364 1571 3380 1576
rect 3354 1564 3360 1565
rect 3363 1564 3392 1571
rect 3281 1563 3392 1564
rect 3281 1562 3398 1563
rect 2957 1554 3008 1562
rect 3055 1554 3089 1562
rect 2957 1542 2982 1554
rect 2989 1542 3008 1554
rect 3062 1552 3089 1554
rect 3098 1552 3319 1562
rect 3354 1559 3360 1562
rect 3062 1548 3319 1552
rect 2957 1534 3008 1542
rect 3055 1534 3319 1548
rect 3363 1554 3398 1562
rect 2909 1486 2928 1520
rect 2973 1526 3002 1534
rect 2973 1520 2990 1526
rect 2973 1518 3007 1520
rect 3055 1518 3071 1534
rect 3072 1524 3280 1534
rect 3281 1524 3297 1534
rect 3345 1530 3360 1545
rect 3363 1542 3364 1554
rect 3371 1542 3398 1554
rect 3363 1534 3398 1542
rect 3363 1533 3392 1534
rect 3083 1520 3297 1524
rect 3098 1518 3297 1520
rect 3332 1520 3345 1530
rect 3363 1520 3380 1533
rect 3332 1518 3380 1520
rect 2974 1514 3007 1518
rect 2970 1512 3007 1514
rect 2970 1511 3037 1512
rect 2970 1506 3001 1511
rect 3007 1506 3037 1511
rect 2970 1502 3037 1506
rect 2943 1499 3037 1502
rect 2943 1492 2992 1499
rect 2943 1486 2973 1492
rect 2992 1487 2997 1492
rect 2909 1470 2989 1486
rect 3001 1478 3037 1499
rect 3098 1494 3287 1518
rect 3332 1517 3379 1518
rect 3345 1512 3379 1517
rect 3113 1491 3287 1494
rect 3106 1488 3287 1491
rect 3315 1511 3379 1512
rect 2909 1468 2928 1470
rect 2943 1468 2977 1470
rect 2909 1452 2989 1468
rect 2909 1446 2928 1452
rect 2625 1420 2728 1430
rect 2579 1418 2728 1420
rect 2749 1418 2784 1430
rect 2418 1416 2580 1418
rect 2430 1396 2449 1416
rect 2464 1414 2494 1416
rect 2313 1388 2354 1396
rect 2436 1392 2449 1396
rect 2501 1400 2580 1416
rect 2612 1416 2784 1418
rect 2612 1400 2691 1416
rect 2698 1414 2728 1416
rect 2276 1378 2305 1388
rect 2319 1378 2348 1388
rect 2363 1378 2393 1392
rect 2436 1378 2479 1392
rect 2501 1388 2691 1400
rect 2756 1396 2762 1416
rect 2486 1378 2516 1388
rect 2517 1378 2675 1388
rect 2679 1378 2709 1388
rect 2713 1378 2743 1392
rect 2771 1378 2784 1416
rect 2856 1430 2885 1446
rect 2899 1430 2928 1446
rect 2943 1436 2973 1452
rect 3001 1430 3007 1478
rect 3010 1472 3029 1478
rect 3044 1472 3074 1480
rect 3010 1464 3074 1472
rect 3010 1448 3090 1464
rect 3106 1457 3168 1488
rect 3184 1457 3246 1488
rect 3315 1486 3364 1511
rect 3379 1486 3409 1502
rect 3278 1472 3308 1480
rect 3315 1478 3425 1486
rect 3278 1464 3323 1472
rect 3010 1446 3029 1448
rect 3044 1446 3090 1448
rect 3010 1430 3090 1446
rect 3117 1444 3152 1457
rect 3193 1454 3230 1457
rect 3193 1452 3235 1454
rect 3122 1441 3152 1444
rect 3131 1437 3138 1441
rect 3138 1436 3139 1437
rect 3097 1430 3107 1436
rect 2856 1422 2891 1430
rect 2856 1396 2857 1422
rect 2864 1396 2891 1422
rect 2799 1378 2829 1392
rect 2856 1388 2891 1396
rect 2893 1422 2934 1430
rect 2893 1396 2908 1422
rect 2915 1396 2934 1422
rect 2998 1418 3029 1430
rect 3044 1418 3147 1430
rect 3159 1420 3185 1446
rect 3200 1441 3230 1452
rect 3262 1448 3324 1464
rect 3262 1446 3308 1448
rect 3262 1430 3324 1446
rect 3336 1430 3342 1478
rect 3345 1470 3425 1478
rect 3345 1468 3364 1470
rect 3379 1468 3413 1470
rect 3345 1452 3425 1468
rect 3345 1430 3364 1452
rect 3379 1436 3409 1452
rect 3437 1446 3443 1520
rect 3446 1446 3465 1590
rect 3480 1446 3486 1590
rect 3495 1520 3508 1590
rect 3560 1586 3582 1590
rect 3553 1564 3582 1578
rect 3635 1564 3651 1578
rect 3689 1574 3695 1576
rect 3702 1574 3810 1590
rect 3817 1574 3823 1576
rect 3831 1574 3846 1590
rect 3912 1584 3931 1587
rect 3553 1562 3651 1564
rect 3678 1562 3846 1574
rect 3861 1564 3877 1578
rect 3912 1565 3934 1584
rect 3944 1578 3960 1579
rect 3943 1576 3960 1578
rect 3944 1571 3960 1576
rect 3934 1564 3940 1565
rect 3943 1564 3972 1571
rect 3861 1563 3972 1564
rect 3861 1562 3978 1563
rect 3537 1554 3588 1562
rect 3635 1554 3669 1562
rect 3537 1542 3562 1554
rect 3569 1542 3588 1554
rect 3642 1552 3669 1554
rect 3678 1552 3899 1562
rect 3934 1559 3940 1562
rect 3642 1548 3899 1552
rect 3537 1534 3588 1542
rect 3635 1534 3899 1548
rect 3943 1554 3978 1562
rect 3489 1486 3508 1520
rect 3553 1526 3582 1534
rect 3553 1520 3570 1526
rect 3553 1518 3587 1520
rect 3635 1518 3651 1534
rect 3652 1524 3860 1534
rect 3861 1524 3877 1534
rect 3925 1530 3940 1545
rect 3943 1542 3944 1554
rect 3951 1542 3978 1554
rect 3943 1534 3978 1542
rect 3943 1533 3972 1534
rect 3663 1520 3877 1524
rect 3678 1518 3877 1520
rect 3912 1520 3925 1530
rect 3943 1520 3960 1533
rect 3912 1518 3960 1520
rect 3554 1514 3587 1518
rect 3550 1512 3587 1514
rect 3550 1511 3617 1512
rect 3550 1506 3581 1511
rect 3587 1506 3617 1511
rect 3550 1502 3617 1506
rect 3523 1499 3617 1502
rect 3523 1492 3572 1499
rect 3523 1486 3553 1492
rect 3572 1487 3577 1492
rect 3489 1470 3569 1486
rect 3581 1478 3617 1499
rect 3678 1494 3867 1518
rect 3912 1517 3959 1518
rect 3925 1512 3959 1517
rect 3693 1491 3867 1494
rect 3686 1488 3867 1491
rect 3895 1511 3959 1512
rect 3489 1468 3508 1470
rect 3523 1468 3557 1470
rect 3489 1452 3569 1468
rect 3489 1446 3508 1452
rect 3205 1420 3308 1430
rect 3159 1418 3308 1420
rect 3329 1418 3364 1430
rect 2998 1416 3160 1418
rect 3010 1396 3029 1416
rect 3044 1414 3074 1416
rect 2893 1388 2934 1396
rect 3016 1392 3029 1396
rect 3081 1400 3160 1416
rect 3192 1416 3364 1418
rect 3192 1400 3271 1416
rect 3278 1414 3308 1416
rect 2856 1378 2885 1388
rect 2899 1378 2928 1388
rect 2943 1378 2973 1392
rect 3016 1378 3059 1392
rect 3081 1388 3271 1400
rect 3336 1396 3342 1416
rect 3066 1378 3096 1388
rect 3097 1378 3255 1388
rect 3259 1378 3289 1388
rect 3293 1378 3323 1392
rect 3351 1378 3364 1416
rect 3436 1430 3465 1446
rect 3479 1430 3508 1446
rect 3523 1436 3553 1452
rect 3581 1430 3587 1478
rect 3590 1472 3609 1478
rect 3624 1472 3654 1480
rect 3590 1464 3654 1472
rect 3590 1448 3670 1464
rect 3686 1457 3748 1488
rect 3764 1457 3826 1488
rect 3895 1486 3944 1511
rect 3959 1486 3989 1502
rect 3858 1472 3888 1480
rect 3895 1478 4005 1486
rect 3858 1464 3903 1472
rect 3590 1446 3609 1448
rect 3624 1446 3670 1448
rect 3590 1430 3670 1446
rect 3697 1444 3732 1457
rect 3773 1454 3810 1457
rect 3773 1452 3815 1454
rect 3702 1441 3732 1444
rect 3711 1437 3718 1441
rect 3718 1436 3719 1437
rect 3677 1430 3687 1436
rect 3436 1422 3471 1430
rect 3436 1396 3437 1422
rect 3444 1396 3471 1422
rect 3379 1378 3409 1392
rect 3436 1388 3471 1396
rect 3473 1422 3514 1430
rect 3473 1396 3488 1422
rect 3495 1396 3514 1422
rect 3578 1418 3609 1430
rect 3624 1418 3727 1430
rect 3739 1420 3765 1446
rect 3780 1441 3810 1452
rect 3842 1448 3904 1464
rect 3842 1446 3888 1448
rect 3842 1430 3904 1446
rect 3916 1430 3922 1478
rect 3925 1470 4005 1478
rect 3925 1468 3944 1470
rect 3959 1468 3993 1470
rect 3925 1452 4005 1468
rect 3925 1430 3944 1452
rect 3959 1436 3989 1452
rect 4017 1446 4023 1520
rect 4026 1446 4045 1590
rect 4060 1446 4066 1590
rect 4075 1520 4088 1590
rect 4140 1586 4162 1590
rect 4133 1564 4162 1578
rect 4215 1564 4231 1578
rect 4269 1574 4275 1576
rect 4282 1574 4390 1590
rect 4397 1574 4403 1576
rect 4411 1574 4426 1590
rect 4492 1584 4511 1587
rect 4133 1562 4231 1564
rect 4258 1562 4426 1574
rect 4441 1564 4457 1578
rect 4492 1565 4514 1584
rect 4524 1578 4540 1579
rect 4523 1576 4540 1578
rect 4524 1571 4540 1576
rect 4514 1564 4520 1565
rect 4523 1564 4552 1571
rect 4441 1563 4552 1564
rect 4441 1562 4558 1563
rect 4117 1554 4168 1562
rect 4215 1554 4249 1562
rect 4117 1542 4142 1554
rect 4149 1542 4168 1554
rect 4222 1552 4249 1554
rect 4258 1552 4479 1562
rect 4514 1559 4520 1562
rect 4222 1548 4479 1552
rect 4117 1534 4168 1542
rect 4215 1534 4479 1548
rect 4523 1554 4558 1562
rect 4069 1486 4088 1520
rect 4133 1526 4162 1534
rect 4133 1520 4150 1526
rect 4133 1518 4167 1520
rect 4215 1518 4231 1534
rect 4232 1524 4440 1534
rect 4441 1524 4457 1534
rect 4505 1530 4520 1545
rect 4523 1542 4524 1554
rect 4531 1542 4558 1554
rect 4523 1534 4558 1542
rect 4523 1533 4552 1534
rect 4243 1520 4457 1524
rect 4258 1518 4457 1520
rect 4492 1520 4505 1530
rect 4523 1520 4540 1533
rect 4492 1518 4540 1520
rect 4134 1514 4167 1518
rect 4130 1512 4167 1514
rect 4130 1511 4197 1512
rect 4130 1506 4161 1511
rect 4167 1506 4197 1511
rect 4130 1502 4197 1506
rect 4103 1499 4197 1502
rect 4103 1492 4152 1499
rect 4103 1486 4133 1492
rect 4152 1487 4157 1492
rect 4069 1470 4149 1486
rect 4161 1478 4197 1499
rect 4258 1494 4447 1518
rect 4492 1517 4539 1518
rect 4505 1512 4539 1517
rect 4273 1491 4447 1494
rect 4266 1488 4447 1491
rect 4475 1511 4539 1512
rect 4069 1468 4088 1470
rect 4103 1468 4137 1470
rect 4069 1452 4149 1468
rect 4069 1446 4088 1452
rect 3785 1420 3888 1430
rect 3739 1418 3888 1420
rect 3909 1418 3944 1430
rect 3578 1416 3740 1418
rect 3590 1396 3609 1416
rect 3624 1414 3654 1416
rect 3473 1388 3514 1396
rect 3596 1392 3609 1396
rect 3661 1400 3740 1416
rect 3772 1416 3944 1418
rect 3772 1400 3851 1416
rect 3858 1414 3888 1416
rect 3436 1378 3465 1388
rect 3479 1378 3508 1388
rect 3523 1378 3553 1392
rect 3596 1378 3639 1392
rect 3661 1388 3851 1400
rect 3916 1396 3922 1416
rect 3646 1378 3676 1388
rect 3677 1378 3835 1388
rect 3839 1378 3869 1388
rect 3873 1378 3903 1392
rect 3931 1378 3944 1416
rect 4016 1430 4045 1446
rect 4059 1430 4088 1446
rect 4103 1436 4133 1452
rect 4161 1430 4167 1478
rect 4170 1472 4189 1478
rect 4204 1472 4234 1480
rect 4170 1464 4234 1472
rect 4170 1448 4250 1464
rect 4266 1457 4328 1488
rect 4344 1457 4406 1488
rect 4475 1486 4524 1511
rect 4539 1486 4569 1502
rect 4438 1472 4468 1480
rect 4475 1478 4585 1486
rect 4438 1464 4483 1472
rect 4170 1446 4189 1448
rect 4204 1446 4250 1448
rect 4170 1430 4250 1446
rect 4277 1444 4312 1457
rect 4353 1454 4390 1457
rect 4353 1452 4395 1454
rect 4282 1441 4312 1444
rect 4291 1437 4298 1441
rect 4298 1436 4299 1437
rect 4257 1430 4267 1436
rect 4016 1422 4051 1430
rect 4016 1396 4017 1422
rect 4024 1396 4051 1422
rect 3959 1378 3989 1392
rect 4016 1388 4051 1396
rect 4053 1422 4094 1430
rect 4053 1396 4068 1422
rect 4075 1396 4094 1422
rect 4158 1418 4189 1430
rect 4204 1418 4307 1430
rect 4319 1420 4345 1446
rect 4360 1441 4390 1452
rect 4422 1448 4484 1464
rect 4422 1446 4468 1448
rect 4422 1430 4484 1446
rect 4496 1430 4502 1478
rect 4505 1470 4585 1478
rect 4505 1468 4524 1470
rect 4539 1468 4573 1470
rect 4505 1452 4585 1468
rect 4505 1430 4524 1452
rect 4539 1436 4569 1452
rect 4597 1446 4603 1520
rect 4606 1446 4625 1590
rect 4640 1446 4646 1590
rect 4655 1520 4668 1590
rect 4720 1586 4742 1590
rect 4713 1564 4742 1578
rect 4795 1564 4811 1578
rect 4849 1574 4855 1576
rect 4862 1574 4970 1590
rect 4977 1574 4983 1576
rect 4991 1574 5006 1590
rect 5072 1584 5091 1587
rect 4713 1562 4811 1564
rect 4838 1562 5006 1574
rect 5021 1564 5037 1578
rect 5072 1565 5094 1584
rect 5104 1578 5120 1579
rect 5103 1576 5120 1578
rect 5104 1571 5120 1576
rect 5094 1564 5100 1565
rect 5103 1564 5132 1571
rect 5021 1563 5132 1564
rect 5021 1562 5138 1563
rect 4697 1554 4748 1562
rect 4795 1554 4829 1562
rect 4697 1542 4722 1554
rect 4729 1542 4748 1554
rect 4802 1552 4829 1554
rect 4838 1552 5059 1562
rect 5094 1559 5100 1562
rect 4802 1548 5059 1552
rect 4697 1534 4748 1542
rect 4795 1534 5059 1548
rect 5103 1554 5138 1562
rect 4649 1486 4668 1520
rect 4713 1526 4742 1534
rect 4713 1520 4730 1526
rect 4713 1518 4747 1520
rect 4795 1518 4811 1534
rect 4812 1524 5020 1534
rect 5021 1524 5037 1534
rect 5085 1530 5100 1545
rect 5103 1542 5104 1554
rect 5111 1542 5138 1554
rect 5103 1534 5138 1542
rect 5103 1533 5132 1534
rect 4823 1520 5037 1524
rect 4838 1518 5037 1520
rect 5072 1520 5085 1530
rect 5103 1520 5120 1533
rect 5072 1518 5120 1520
rect 4714 1514 4747 1518
rect 4710 1512 4747 1514
rect 4710 1511 4777 1512
rect 4710 1506 4741 1511
rect 4747 1506 4777 1511
rect 4710 1502 4777 1506
rect 4683 1499 4777 1502
rect 4683 1492 4732 1499
rect 4683 1486 4713 1492
rect 4732 1487 4737 1492
rect 4649 1470 4729 1486
rect 4741 1478 4777 1499
rect 4838 1494 5027 1518
rect 5072 1517 5119 1518
rect 5085 1512 5119 1517
rect 4853 1491 5027 1494
rect 4846 1488 5027 1491
rect 5055 1511 5119 1512
rect 4649 1468 4668 1470
rect 4683 1468 4717 1470
rect 4649 1452 4729 1468
rect 4649 1446 4668 1452
rect 4365 1420 4468 1430
rect 4319 1418 4468 1420
rect 4489 1418 4524 1430
rect 4158 1416 4320 1418
rect 4170 1396 4189 1416
rect 4204 1414 4234 1416
rect 4053 1388 4094 1396
rect 4176 1392 4189 1396
rect 4241 1400 4320 1416
rect 4352 1416 4524 1418
rect 4352 1400 4431 1416
rect 4438 1414 4468 1416
rect 4016 1378 4045 1388
rect 4059 1378 4088 1388
rect 4103 1378 4133 1392
rect 4176 1378 4219 1392
rect 4241 1388 4431 1400
rect 4496 1396 4502 1416
rect 4226 1378 4256 1388
rect 4257 1378 4415 1388
rect 4419 1378 4449 1388
rect 4453 1378 4483 1392
rect 4511 1378 4524 1416
rect 4596 1430 4625 1446
rect 4639 1430 4668 1446
rect 4683 1436 4713 1452
rect 4741 1430 4747 1478
rect 4750 1472 4769 1478
rect 4784 1472 4814 1480
rect 4750 1464 4814 1472
rect 4750 1448 4830 1464
rect 4846 1457 4908 1488
rect 4924 1457 4986 1488
rect 5055 1486 5104 1511
rect 5119 1486 5149 1502
rect 5018 1472 5048 1480
rect 5055 1478 5165 1486
rect 5018 1464 5063 1472
rect 4750 1446 4769 1448
rect 4784 1446 4830 1448
rect 4750 1430 4830 1446
rect 4857 1444 4892 1457
rect 4933 1454 4970 1457
rect 4933 1452 4975 1454
rect 4862 1441 4892 1444
rect 4871 1437 4878 1441
rect 4878 1436 4879 1437
rect 4837 1430 4847 1436
rect 4596 1422 4631 1430
rect 4596 1396 4597 1422
rect 4604 1396 4631 1422
rect 4539 1378 4569 1392
rect 4596 1388 4631 1396
rect 4633 1422 4674 1430
rect 4633 1396 4648 1422
rect 4655 1396 4674 1422
rect 4738 1418 4769 1430
rect 4784 1418 4887 1430
rect 4899 1420 4925 1446
rect 4940 1441 4970 1452
rect 5002 1448 5064 1464
rect 5002 1446 5048 1448
rect 5002 1430 5064 1446
rect 5076 1430 5082 1478
rect 5085 1470 5165 1478
rect 5085 1468 5104 1470
rect 5119 1468 5153 1470
rect 5085 1452 5165 1468
rect 5085 1430 5104 1452
rect 5119 1436 5149 1452
rect 5177 1446 5183 1520
rect 5186 1446 5205 1590
rect 5220 1446 5226 1590
rect 5235 1520 5248 1590
rect 5300 1586 5322 1590
rect 5293 1564 5322 1578
rect 5375 1564 5391 1578
rect 5429 1574 5435 1576
rect 5442 1574 5550 1590
rect 5557 1574 5563 1576
rect 5571 1574 5586 1590
rect 5652 1584 5671 1587
rect 5293 1562 5391 1564
rect 5418 1562 5586 1574
rect 5601 1564 5617 1578
rect 5652 1565 5674 1584
rect 5684 1578 5700 1579
rect 5683 1576 5700 1578
rect 5684 1571 5700 1576
rect 5674 1564 5680 1565
rect 5683 1564 5712 1571
rect 5601 1563 5712 1564
rect 5601 1562 5718 1563
rect 5277 1554 5328 1562
rect 5375 1554 5409 1562
rect 5277 1542 5302 1554
rect 5309 1542 5328 1554
rect 5382 1552 5409 1554
rect 5418 1552 5639 1562
rect 5674 1559 5680 1562
rect 5382 1548 5639 1552
rect 5277 1534 5328 1542
rect 5375 1534 5639 1548
rect 5683 1554 5718 1562
rect 5229 1486 5248 1520
rect 5293 1526 5322 1534
rect 5293 1520 5310 1526
rect 5293 1518 5327 1520
rect 5375 1518 5391 1534
rect 5392 1524 5600 1534
rect 5601 1524 5617 1534
rect 5665 1530 5680 1545
rect 5683 1542 5684 1554
rect 5691 1542 5718 1554
rect 5683 1534 5718 1542
rect 5683 1533 5712 1534
rect 5403 1520 5617 1524
rect 5418 1518 5617 1520
rect 5652 1520 5665 1530
rect 5683 1520 5700 1533
rect 5652 1518 5700 1520
rect 5294 1514 5327 1518
rect 5290 1512 5327 1514
rect 5290 1511 5357 1512
rect 5290 1506 5321 1511
rect 5327 1506 5357 1511
rect 5290 1502 5357 1506
rect 5263 1499 5357 1502
rect 5263 1492 5312 1499
rect 5263 1486 5293 1492
rect 5312 1487 5317 1492
rect 5229 1470 5309 1486
rect 5321 1478 5357 1499
rect 5418 1494 5607 1518
rect 5652 1517 5699 1518
rect 5665 1512 5699 1517
rect 5433 1491 5607 1494
rect 5426 1488 5607 1491
rect 5635 1511 5699 1512
rect 5229 1468 5248 1470
rect 5263 1468 5297 1470
rect 5229 1452 5309 1468
rect 5229 1446 5248 1452
rect 4945 1420 5048 1430
rect 4899 1418 5048 1420
rect 5069 1418 5104 1430
rect 4738 1416 4900 1418
rect 4750 1396 4769 1416
rect 4784 1414 4814 1416
rect 4633 1388 4674 1396
rect 4756 1392 4769 1396
rect 4821 1400 4900 1416
rect 4932 1416 5104 1418
rect 4932 1400 5011 1416
rect 5018 1414 5048 1416
rect 4596 1378 4625 1388
rect 4639 1378 4668 1388
rect 4683 1378 4713 1392
rect 4756 1378 4799 1392
rect 4821 1388 5011 1400
rect 5076 1396 5082 1416
rect 4806 1378 4836 1388
rect 4837 1378 4995 1388
rect 4999 1378 5029 1388
rect 5033 1378 5063 1392
rect 5091 1378 5104 1416
rect 5176 1430 5205 1446
rect 5219 1430 5248 1446
rect 5263 1436 5293 1452
rect 5321 1430 5327 1478
rect 5330 1472 5349 1478
rect 5364 1472 5394 1480
rect 5330 1464 5394 1472
rect 5330 1448 5410 1464
rect 5426 1457 5488 1488
rect 5504 1457 5566 1488
rect 5635 1486 5684 1511
rect 5699 1486 5729 1502
rect 5598 1472 5628 1480
rect 5635 1478 5745 1486
rect 5598 1464 5643 1472
rect 5330 1446 5349 1448
rect 5364 1446 5410 1448
rect 5330 1430 5410 1446
rect 5437 1444 5472 1457
rect 5513 1454 5550 1457
rect 5513 1452 5555 1454
rect 5442 1441 5472 1444
rect 5451 1437 5458 1441
rect 5458 1436 5459 1437
rect 5417 1430 5427 1436
rect 5176 1422 5211 1430
rect 5176 1396 5177 1422
rect 5184 1396 5211 1422
rect 5119 1378 5149 1392
rect 5176 1388 5211 1396
rect 5213 1422 5254 1430
rect 5213 1396 5228 1422
rect 5235 1396 5254 1422
rect 5318 1418 5349 1430
rect 5364 1418 5467 1430
rect 5479 1420 5505 1446
rect 5520 1441 5550 1452
rect 5582 1448 5644 1464
rect 5582 1446 5628 1448
rect 5582 1430 5644 1446
rect 5656 1430 5662 1478
rect 5665 1470 5745 1478
rect 5665 1468 5684 1470
rect 5699 1468 5733 1470
rect 5665 1452 5745 1468
rect 5665 1430 5684 1452
rect 5699 1436 5729 1452
rect 5757 1446 5763 1520
rect 5766 1446 5785 1590
rect 5800 1446 5806 1590
rect 5815 1520 5828 1590
rect 5880 1586 5902 1590
rect 5873 1564 5902 1578
rect 5955 1564 5971 1578
rect 6009 1574 6015 1576
rect 6022 1574 6130 1590
rect 6137 1574 6143 1576
rect 6151 1574 6166 1590
rect 6232 1584 6251 1587
rect 5873 1562 5971 1564
rect 5998 1562 6166 1574
rect 6181 1564 6197 1578
rect 6232 1565 6254 1584
rect 6264 1578 6280 1579
rect 6263 1576 6280 1578
rect 6264 1571 6280 1576
rect 6254 1564 6260 1565
rect 6263 1564 6292 1571
rect 6181 1563 6292 1564
rect 6181 1562 6298 1563
rect 5857 1554 5908 1562
rect 5955 1554 5989 1562
rect 5857 1542 5882 1554
rect 5889 1542 5908 1554
rect 5962 1552 5989 1554
rect 5998 1552 6219 1562
rect 6254 1559 6260 1562
rect 5962 1548 6219 1552
rect 5857 1534 5908 1542
rect 5955 1534 6219 1548
rect 6263 1554 6298 1562
rect 5809 1486 5828 1520
rect 5873 1526 5902 1534
rect 5873 1520 5890 1526
rect 5873 1518 5907 1520
rect 5955 1518 5971 1534
rect 5972 1524 6180 1534
rect 6181 1524 6197 1534
rect 6245 1530 6260 1545
rect 6263 1542 6264 1554
rect 6271 1542 6298 1554
rect 6263 1534 6298 1542
rect 6263 1533 6292 1534
rect 5983 1520 6197 1524
rect 5998 1518 6197 1520
rect 6232 1520 6245 1530
rect 6263 1520 6280 1533
rect 6232 1518 6280 1520
rect 5874 1514 5907 1518
rect 5870 1512 5907 1514
rect 5870 1511 5937 1512
rect 5870 1506 5901 1511
rect 5907 1506 5937 1511
rect 5870 1502 5937 1506
rect 5843 1499 5937 1502
rect 5843 1492 5892 1499
rect 5843 1486 5873 1492
rect 5892 1487 5897 1492
rect 5809 1470 5889 1486
rect 5901 1478 5937 1499
rect 5998 1494 6187 1518
rect 6232 1517 6279 1518
rect 6245 1512 6279 1517
rect 6013 1491 6187 1494
rect 6006 1488 6187 1491
rect 6215 1511 6279 1512
rect 5809 1468 5828 1470
rect 5843 1468 5877 1470
rect 5809 1452 5889 1468
rect 5809 1446 5828 1452
rect 5525 1420 5628 1430
rect 5479 1418 5628 1420
rect 5649 1418 5684 1430
rect 5318 1416 5480 1418
rect 5330 1396 5349 1416
rect 5364 1414 5394 1416
rect 5213 1388 5254 1396
rect 5336 1392 5349 1396
rect 5401 1400 5480 1416
rect 5512 1416 5684 1418
rect 5512 1400 5591 1416
rect 5598 1414 5628 1416
rect 5176 1378 5205 1388
rect 5219 1378 5248 1388
rect 5263 1378 5293 1392
rect 5336 1378 5379 1392
rect 5401 1388 5591 1400
rect 5656 1396 5662 1416
rect 5386 1378 5416 1388
rect 5417 1378 5575 1388
rect 5579 1378 5609 1388
rect 5613 1378 5643 1392
rect 5671 1378 5684 1416
rect 5756 1430 5785 1446
rect 5799 1430 5828 1446
rect 5843 1436 5873 1452
rect 5901 1430 5907 1478
rect 5910 1472 5929 1478
rect 5944 1472 5974 1480
rect 5910 1464 5974 1472
rect 5910 1448 5990 1464
rect 6006 1457 6068 1488
rect 6084 1457 6146 1488
rect 6215 1486 6264 1511
rect 6279 1486 6309 1502
rect 6178 1472 6208 1480
rect 6215 1478 6325 1486
rect 6178 1464 6223 1472
rect 5910 1446 5929 1448
rect 5944 1446 5990 1448
rect 5910 1430 5990 1446
rect 6017 1444 6052 1457
rect 6093 1454 6130 1457
rect 6093 1452 6135 1454
rect 6022 1441 6052 1444
rect 6031 1437 6038 1441
rect 6038 1436 6039 1437
rect 5997 1430 6007 1436
rect 5756 1422 5791 1430
rect 5756 1396 5757 1422
rect 5764 1396 5791 1422
rect 5699 1378 5729 1392
rect 5756 1388 5791 1396
rect 5793 1422 5834 1430
rect 5793 1396 5808 1422
rect 5815 1396 5834 1422
rect 5898 1418 5929 1430
rect 5944 1418 6047 1430
rect 6059 1420 6085 1446
rect 6100 1441 6130 1452
rect 6162 1448 6224 1464
rect 6162 1446 6208 1448
rect 6162 1430 6224 1446
rect 6236 1430 6242 1478
rect 6245 1470 6325 1478
rect 6245 1468 6264 1470
rect 6279 1468 6313 1470
rect 6245 1452 6325 1468
rect 6245 1430 6264 1452
rect 6279 1436 6309 1452
rect 6337 1446 6343 1520
rect 6346 1446 6365 1590
rect 6380 1446 6386 1590
rect 6395 1520 6408 1590
rect 6460 1586 6482 1590
rect 6453 1564 6482 1578
rect 6535 1564 6551 1578
rect 6589 1574 6595 1576
rect 6602 1574 6710 1590
rect 6717 1574 6723 1576
rect 6731 1574 6746 1590
rect 6812 1584 6831 1587
rect 6453 1562 6551 1564
rect 6578 1562 6746 1574
rect 6761 1564 6777 1578
rect 6812 1565 6834 1584
rect 6844 1578 6860 1579
rect 6843 1576 6860 1578
rect 6844 1571 6860 1576
rect 6834 1564 6840 1565
rect 6843 1564 6872 1571
rect 6761 1563 6872 1564
rect 6761 1562 6878 1563
rect 6437 1554 6488 1562
rect 6535 1554 6569 1562
rect 6437 1542 6462 1554
rect 6469 1542 6488 1554
rect 6542 1552 6569 1554
rect 6578 1552 6799 1562
rect 6834 1559 6840 1562
rect 6542 1548 6799 1552
rect 6437 1534 6488 1542
rect 6535 1534 6799 1548
rect 6843 1554 6878 1562
rect 6389 1486 6408 1520
rect 6453 1526 6482 1534
rect 6453 1520 6470 1526
rect 6453 1518 6487 1520
rect 6535 1518 6551 1534
rect 6552 1524 6760 1534
rect 6761 1524 6777 1534
rect 6825 1530 6840 1545
rect 6843 1542 6844 1554
rect 6851 1542 6878 1554
rect 6843 1534 6878 1542
rect 6843 1533 6872 1534
rect 6563 1520 6777 1524
rect 6578 1518 6777 1520
rect 6812 1520 6825 1530
rect 6843 1520 6860 1533
rect 6812 1518 6860 1520
rect 6454 1514 6487 1518
rect 6450 1512 6487 1514
rect 6450 1511 6517 1512
rect 6450 1506 6481 1511
rect 6487 1506 6517 1511
rect 6450 1502 6517 1506
rect 6423 1499 6517 1502
rect 6423 1492 6472 1499
rect 6423 1486 6453 1492
rect 6472 1487 6477 1492
rect 6389 1470 6469 1486
rect 6481 1478 6517 1499
rect 6578 1494 6767 1518
rect 6812 1517 6859 1518
rect 6825 1512 6859 1517
rect 6593 1491 6767 1494
rect 6586 1488 6767 1491
rect 6795 1511 6859 1512
rect 6389 1468 6408 1470
rect 6423 1468 6457 1470
rect 6389 1452 6469 1468
rect 6389 1446 6408 1452
rect 6105 1420 6208 1430
rect 6059 1418 6208 1420
rect 6229 1418 6264 1430
rect 5898 1416 6060 1418
rect 5910 1396 5929 1416
rect 5944 1414 5974 1416
rect 5793 1388 5834 1396
rect 5916 1392 5929 1396
rect 5981 1400 6060 1416
rect 6092 1416 6264 1418
rect 6092 1400 6171 1416
rect 6178 1414 6208 1416
rect 5756 1378 5785 1388
rect 5799 1378 5828 1388
rect 5843 1378 5873 1392
rect 5916 1378 5959 1392
rect 5981 1388 6171 1400
rect 6236 1396 6242 1416
rect 5966 1378 5996 1388
rect 5997 1378 6155 1388
rect 6159 1378 6189 1388
rect 6193 1378 6223 1392
rect 6251 1378 6264 1416
rect 6336 1430 6365 1446
rect 6379 1430 6408 1446
rect 6423 1436 6453 1452
rect 6481 1430 6487 1478
rect 6490 1472 6509 1478
rect 6524 1472 6554 1480
rect 6490 1464 6554 1472
rect 6490 1448 6570 1464
rect 6586 1457 6648 1488
rect 6664 1457 6726 1488
rect 6795 1486 6844 1511
rect 6859 1486 6889 1502
rect 6758 1472 6788 1480
rect 6795 1478 6905 1486
rect 6758 1464 6803 1472
rect 6490 1446 6509 1448
rect 6524 1446 6570 1448
rect 6490 1430 6570 1446
rect 6597 1444 6632 1457
rect 6673 1454 6710 1457
rect 6673 1452 6715 1454
rect 6602 1441 6632 1444
rect 6611 1437 6618 1441
rect 6618 1436 6619 1437
rect 6577 1430 6587 1436
rect 6336 1422 6371 1430
rect 6336 1396 6337 1422
rect 6344 1396 6371 1422
rect 6279 1378 6309 1392
rect 6336 1388 6371 1396
rect 6373 1422 6414 1430
rect 6373 1396 6388 1422
rect 6395 1396 6414 1422
rect 6478 1418 6509 1430
rect 6524 1418 6627 1430
rect 6639 1420 6665 1446
rect 6680 1441 6710 1452
rect 6742 1448 6804 1464
rect 6742 1446 6788 1448
rect 6742 1430 6804 1446
rect 6816 1430 6822 1478
rect 6825 1470 6905 1478
rect 6825 1468 6844 1470
rect 6859 1468 6893 1470
rect 6825 1452 6905 1468
rect 6825 1430 6844 1452
rect 6859 1436 6889 1452
rect 6917 1446 6923 1520
rect 6926 1446 6945 1590
rect 6960 1446 6966 1590
rect 6975 1520 6988 1590
rect 7040 1586 7062 1590
rect 7033 1564 7062 1578
rect 7115 1564 7131 1578
rect 7169 1574 7175 1576
rect 7182 1574 7290 1590
rect 7297 1574 7303 1576
rect 7311 1574 7326 1590
rect 7392 1584 7411 1587
rect 7033 1562 7131 1564
rect 7158 1562 7326 1574
rect 7341 1564 7357 1578
rect 7392 1565 7414 1584
rect 7424 1578 7440 1579
rect 7423 1576 7440 1578
rect 7424 1571 7440 1576
rect 7414 1564 7420 1565
rect 7423 1564 7452 1571
rect 7341 1563 7452 1564
rect 7341 1562 7458 1563
rect 7017 1554 7068 1562
rect 7115 1554 7149 1562
rect 7017 1542 7042 1554
rect 7049 1542 7068 1554
rect 7122 1552 7149 1554
rect 7158 1552 7379 1562
rect 7414 1559 7420 1562
rect 7122 1548 7379 1552
rect 7017 1534 7068 1542
rect 7115 1534 7379 1548
rect 7423 1554 7458 1562
rect 6969 1486 6988 1520
rect 7033 1526 7062 1534
rect 7033 1520 7050 1526
rect 7033 1518 7067 1520
rect 7115 1518 7131 1534
rect 7132 1524 7340 1534
rect 7341 1524 7357 1534
rect 7405 1530 7420 1545
rect 7423 1542 7424 1554
rect 7431 1542 7458 1554
rect 7423 1534 7458 1542
rect 7423 1533 7452 1534
rect 7143 1520 7357 1524
rect 7158 1518 7357 1520
rect 7392 1520 7405 1530
rect 7423 1520 7440 1533
rect 7392 1518 7440 1520
rect 7034 1514 7067 1518
rect 7030 1512 7067 1514
rect 7030 1511 7097 1512
rect 7030 1506 7061 1511
rect 7067 1506 7097 1511
rect 7030 1502 7097 1506
rect 7003 1499 7097 1502
rect 7003 1492 7052 1499
rect 7003 1486 7033 1492
rect 7052 1487 7057 1492
rect 6969 1470 7049 1486
rect 7061 1478 7097 1499
rect 7158 1494 7347 1518
rect 7392 1517 7439 1518
rect 7405 1512 7439 1517
rect 7173 1491 7347 1494
rect 7166 1488 7347 1491
rect 7375 1511 7439 1512
rect 6969 1468 6988 1470
rect 7003 1468 7037 1470
rect 6969 1452 7049 1468
rect 6969 1446 6988 1452
rect 6685 1420 6788 1430
rect 6639 1418 6788 1420
rect 6809 1418 6844 1430
rect 6478 1416 6640 1418
rect 6490 1396 6509 1416
rect 6524 1414 6554 1416
rect 6373 1388 6414 1396
rect 6496 1392 6509 1396
rect 6561 1400 6640 1416
rect 6672 1416 6844 1418
rect 6672 1400 6751 1416
rect 6758 1414 6788 1416
rect 6336 1378 6365 1388
rect 6379 1378 6408 1388
rect 6423 1378 6453 1392
rect 6496 1378 6539 1392
rect 6561 1388 6751 1400
rect 6816 1396 6822 1416
rect 6546 1378 6576 1388
rect 6577 1378 6735 1388
rect 6739 1378 6769 1388
rect 6773 1378 6803 1392
rect 6831 1378 6844 1416
rect 6916 1430 6945 1446
rect 6959 1430 6988 1446
rect 7003 1436 7033 1452
rect 7061 1430 7067 1478
rect 7070 1472 7089 1478
rect 7104 1472 7134 1480
rect 7070 1464 7134 1472
rect 7070 1448 7150 1464
rect 7166 1457 7228 1488
rect 7244 1457 7306 1488
rect 7375 1486 7424 1511
rect 7439 1486 7469 1502
rect 7338 1472 7368 1480
rect 7375 1478 7485 1486
rect 7338 1464 7383 1472
rect 7070 1446 7089 1448
rect 7104 1446 7150 1448
rect 7070 1430 7150 1446
rect 7177 1444 7212 1457
rect 7253 1454 7290 1457
rect 7253 1452 7295 1454
rect 7182 1441 7212 1444
rect 7191 1437 7198 1441
rect 7198 1436 7199 1437
rect 7157 1430 7167 1436
rect 6916 1422 6951 1430
rect 6916 1396 6917 1422
rect 6924 1396 6951 1422
rect 6859 1378 6889 1392
rect 6916 1388 6951 1396
rect 6953 1422 6994 1430
rect 6953 1396 6968 1422
rect 6975 1396 6994 1422
rect 7058 1418 7089 1430
rect 7104 1418 7207 1430
rect 7219 1420 7245 1446
rect 7260 1441 7290 1452
rect 7322 1448 7384 1464
rect 7322 1446 7368 1448
rect 7322 1430 7384 1446
rect 7396 1430 7402 1478
rect 7405 1470 7485 1478
rect 7405 1468 7424 1470
rect 7439 1468 7473 1470
rect 7405 1452 7485 1468
rect 7405 1430 7424 1452
rect 7439 1436 7469 1452
rect 7497 1446 7503 1520
rect 7506 1446 7525 1590
rect 7540 1446 7546 1590
rect 7555 1520 7568 1590
rect 7620 1586 7642 1590
rect 7613 1564 7642 1578
rect 7695 1564 7711 1578
rect 7749 1574 7755 1576
rect 7762 1574 7870 1590
rect 7877 1574 7883 1576
rect 7891 1574 7906 1590
rect 7972 1584 7991 1587
rect 7613 1562 7711 1564
rect 7738 1562 7906 1574
rect 7921 1564 7937 1578
rect 7972 1565 7994 1584
rect 8004 1578 8020 1579
rect 8003 1576 8020 1578
rect 8004 1571 8020 1576
rect 7994 1564 8000 1565
rect 8003 1564 8032 1571
rect 7921 1563 8032 1564
rect 7921 1562 8038 1563
rect 7597 1554 7648 1562
rect 7695 1554 7729 1562
rect 7597 1542 7622 1554
rect 7629 1542 7648 1554
rect 7702 1552 7729 1554
rect 7738 1552 7959 1562
rect 7994 1559 8000 1562
rect 7702 1548 7959 1552
rect 7597 1534 7648 1542
rect 7695 1534 7959 1548
rect 8003 1554 8038 1562
rect 7549 1486 7568 1520
rect 7613 1526 7642 1534
rect 7613 1520 7630 1526
rect 7613 1518 7647 1520
rect 7695 1518 7711 1534
rect 7712 1524 7920 1534
rect 7921 1524 7937 1534
rect 7985 1530 8000 1545
rect 8003 1542 8004 1554
rect 8011 1542 8038 1554
rect 8003 1534 8038 1542
rect 8003 1533 8032 1534
rect 7723 1520 7937 1524
rect 7738 1518 7937 1520
rect 7972 1520 7985 1530
rect 8003 1520 8020 1533
rect 7972 1518 8020 1520
rect 7614 1514 7647 1518
rect 7610 1512 7647 1514
rect 7610 1511 7677 1512
rect 7610 1506 7641 1511
rect 7647 1506 7677 1511
rect 7610 1502 7677 1506
rect 7583 1499 7677 1502
rect 7583 1492 7632 1499
rect 7583 1486 7613 1492
rect 7632 1487 7637 1492
rect 7549 1470 7629 1486
rect 7641 1478 7677 1499
rect 7738 1494 7927 1518
rect 7972 1517 8019 1518
rect 7985 1512 8019 1517
rect 7753 1491 7927 1494
rect 7746 1488 7927 1491
rect 7955 1511 8019 1512
rect 7549 1468 7568 1470
rect 7583 1468 7617 1470
rect 7549 1452 7629 1468
rect 7549 1446 7568 1452
rect 7265 1420 7368 1430
rect 7219 1418 7368 1420
rect 7389 1418 7424 1430
rect 7058 1416 7220 1418
rect 7070 1396 7089 1416
rect 7104 1414 7134 1416
rect 6953 1388 6994 1396
rect 7076 1392 7089 1396
rect 7141 1400 7220 1416
rect 7252 1416 7424 1418
rect 7252 1400 7331 1416
rect 7338 1414 7368 1416
rect 6916 1378 6945 1388
rect 6959 1378 6988 1388
rect 7003 1378 7033 1392
rect 7076 1378 7119 1392
rect 7141 1388 7331 1400
rect 7396 1396 7402 1416
rect 7126 1378 7156 1388
rect 7157 1378 7315 1388
rect 7319 1378 7349 1388
rect 7353 1378 7383 1392
rect 7411 1378 7424 1416
rect 7496 1430 7525 1446
rect 7539 1430 7568 1446
rect 7583 1436 7613 1452
rect 7641 1430 7647 1478
rect 7650 1472 7669 1478
rect 7684 1472 7714 1480
rect 7650 1464 7714 1472
rect 7650 1448 7730 1464
rect 7746 1457 7808 1488
rect 7824 1457 7886 1488
rect 7955 1486 8004 1511
rect 8019 1486 8049 1502
rect 7918 1472 7948 1480
rect 7955 1478 8065 1486
rect 7918 1464 7963 1472
rect 7650 1446 7669 1448
rect 7684 1446 7730 1448
rect 7650 1430 7730 1446
rect 7757 1444 7792 1457
rect 7833 1454 7870 1457
rect 7833 1452 7875 1454
rect 7762 1441 7792 1444
rect 7771 1437 7778 1441
rect 7778 1436 7779 1437
rect 7737 1430 7747 1436
rect 7496 1422 7531 1430
rect 7496 1396 7497 1422
rect 7504 1396 7531 1422
rect 7439 1378 7469 1392
rect 7496 1388 7531 1396
rect 7533 1422 7574 1430
rect 7533 1396 7548 1422
rect 7555 1396 7574 1422
rect 7638 1418 7669 1430
rect 7684 1418 7787 1430
rect 7799 1420 7825 1446
rect 7840 1441 7870 1452
rect 7902 1448 7964 1464
rect 7902 1446 7948 1448
rect 7902 1430 7964 1446
rect 7976 1430 7982 1478
rect 7985 1470 8065 1478
rect 7985 1468 8004 1470
rect 8019 1468 8053 1470
rect 7985 1452 8065 1468
rect 7985 1430 8004 1452
rect 8019 1436 8049 1452
rect 8077 1446 8083 1520
rect 8086 1446 8105 1590
rect 8120 1446 8126 1590
rect 8135 1520 8148 1590
rect 8200 1586 8222 1590
rect 8193 1564 8222 1578
rect 8275 1564 8291 1578
rect 8329 1574 8335 1576
rect 8342 1574 8450 1590
rect 8457 1574 8463 1576
rect 8471 1574 8486 1590
rect 8552 1584 8571 1587
rect 8193 1562 8291 1564
rect 8318 1562 8486 1574
rect 8501 1564 8517 1578
rect 8552 1565 8574 1584
rect 8584 1578 8600 1579
rect 8583 1576 8600 1578
rect 8584 1571 8600 1576
rect 8574 1564 8580 1565
rect 8583 1564 8612 1571
rect 8501 1563 8612 1564
rect 8501 1562 8618 1563
rect 8177 1554 8228 1562
rect 8275 1554 8309 1562
rect 8177 1542 8202 1554
rect 8209 1542 8228 1554
rect 8282 1552 8309 1554
rect 8318 1552 8539 1562
rect 8574 1559 8580 1562
rect 8282 1548 8539 1552
rect 8177 1534 8228 1542
rect 8275 1534 8539 1548
rect 8583 1554 8618 1562
rect 8129 1486 8148 1520
rect 8193 1526 8222 1534
rect 8193 1520 8210 1526
rect 8193 1518 8227 1520
rect 8275 1518 8291 1534
rect 8292 1524 8500 1534
rect 8501 1524 8517 1534
rect 8565 1530 8580 1545
rect 8583 1542 8584 1554
rect 8591 1542 8618 1554
rect 8583 1534 8618 1542
rect 8583 1533 8612 1534
rect 8303 1520 8517 1524
rect 8318 1518 8517 1520
rect 8552 1520 8565 1530
rect 8583 1520 8600 1533
rect 8552 1518 8600 1520
rect 8194 1514 8227 1518
rect 8190 1512 8227 1514
rect 8190 1511 8257 1512
rect 8190 1506 8221 1511
rect 8227 1506 8257 1511
rect 8190 1502 8257 1506
rect 8163 1499 8257 1502
rect 8163 1492 8212 1499
rect 8163 1486 8193 1492
rect 8212 1487 8217 1492
rect 8129 1470 8209 1486
rect 8221 1478 8257 1499
rect 8318 1494 8507 1518
rect 8552 1517 8599 1518
rect 8565 1512 8599 1517
rect 8333 1491 8507 1494
rect 8326 1488 8507 1491
rect 8535 1511 8599 1512
rect 8129 1468 8148 1470
rect 8163 1468 8197 1470
rect 8129 1452 8209 1468
rect 8129 1446 8148 1452
rect 7845 1420 7948 1430
rect 7799 1418 7948 1420
rect 7969 1418 8004 1430
rect 7638 1416 7800 1418
rect 7650 1396 7669 1416
rect 7684 1414 7714 1416
rect 7533 1388 7574 1396
rect 7656 1392 7669 1396
rect 7721 1400 7800 1416
rect 7832 1416 8004 1418
rect 7832 1400 7911 1416
rect 7918 1414 7948 1416
rect 7496 1378 7525 1388
rect 7539 1378 7568 1388
rect 7583 1378 7613 1392
rect 7656 1378 7699 1392
rect 7721 1388 7911 1400
rect 7976 1396 7982 1416
rect 7706 1378 7736 1388
rect 7737 1378 7895 1388
rect 7899 1378 7929 1388
rect 7933 1378 7963 1392
rect 7991 1378 8004 1416
rect 8076 1430 8105 1446
rect 8119 1430 8148 1446
rect 8163 1436 8193 1452
rect 8221 1430 8227 1478
rect 8230 1472 8249 1478
rect 8264 1472 8294 1480
rect 8230 1464 8294 1472
rect 8230 1448 8310 1464
rect 8326 1457 8388 1488
rect 8404 1457 8466 1488
rect 8535 1486 8584 1511
rect 8599 1486 8629 1502
rect 8498 1472 8528 1480
rect 8535 1478 8645 1486
rect 8498 1464 8543 1472
rect 8230 1446 8249 1448
rect 8264 1446 8310 1448
rect 8230 1430 8310 1446
rect 8337 1444 8372 1457
rect 8413 1454 8450 1457
rect 8413 1452 8455 1454
rect 8342 1441 8372 1444
rect 8351 1437 8358 1441
rect 8358 1436 8359 1437
rect 8317 1430 8327 1436
rect 8076 1422 8111 1430
rect 8076 1396 8077 1422
rect 8084 1396 8111 1422
rect 8019 1378 8049 1392
rect 8076 1388 8111 1396
rect 8113 1422 8154 1430
rect 8113 1396 8128 1422
rect 8135 1396 8154 1422
rect 8218 1418 8249 1430
rect 8264 1418 8367 1430
rect 8379 1420 8405 1446
rect 8420 1441 8450 1452
rect 8482 1448 8544 1464
rect 8482 1446 8528 1448
rect 8482 1430 8544 1446
rect 8556 1430 8562 1478
rect 8565 1470 8645 1478
rect 8565 1468 8584 1470
rect 8599 1468 8633 1470
rect 8565 1452 8645 1468
rect 8565 1430 8584 1452
rect 8599 1436 8629 1452
rect 8657 1446 8663 1520
rect 8666 1446 8685 1590
rect 8700 1446 8706 1590
rect 8715 1520 8728 1590
rect 8780 1586 8802 1590
rect 8773 1564 8802 1578
rect 8855 1564 8871 1578
rect 8909 1574 8915 1576
rect 8922 1574 9030 1590
rect 9037 1574 9043 1576
rect 9051 1574 9066 1590
rect 9132 1584 9151 1587
rect 8773 1562 8871 1564
rect 8898 1562 9066 1574
rect 9081 1564 9097 1578
rect 9132 1565 9154 1584
rect 9164 1578 9180 1579
rect 9163 1576 9180 1578
rect 9164 1571 9180 1576
rect 9154 1564 9160 1565
rect 9163 1564 9192 1571
rect 9081 1563 9192 1564
rect 9081 1562 9198 1563
rect 8757 1554 8808 1562
rect 8855 1554 8889 1562
rect 8757 1542 8782 1554
rect 8789 1542 8808 1554
rect 8862 1552 8889 1554
rect 8898 1552 9119 1562
rect 9154 1559 9160 1562
rect 8862 1548 9119 1552
rect 8757 1534 8808 1542
rect 8855 1534 9119 1548
rect 9163 1554 9198 1562
rect 8709 1486 8728 1520
rect 8773 1526 8802 1534
rect 8773 1520 8790 1526
rect 8773 1518 8807 1520
rect 8855 1518 8871 1534
rect 8872 1524 9080 1534
rect 9081 1524 9097 1534
rect 9145 1530 9160 1545
rect 9163 1542 9164 1554
rect 9171 1542 9198 1554
rect 9163 1534 9198 1542
rect 9163 1533 9192 1534
rect 8883 1520 9097 1524
rect 8898 1518 9097 1520
rect 9132 1520 9145 1530
rect 9163 1520 9180 1533
rect 9132 1518 9180 1520
rect 8774 1514 8807 1518
rect 8770 1512 8807 1514
rect 8770 1511 8837 1512
rect 8770 1506 8801 1511
rect 8807 1506 8837 1511
rect 8770 1502 8837 1506
rect 8743 1499 8837 1502
rect 8743 1492 8792 1499
rect 8743 1486 8773 1492
rect 8792 1487 8797 1492
rect 8709 1470 8789 1486
rect 8801 1478 8837 1499
rect 8898 1494 9087 1518
rect 9132 1517 9179 1518
rect 9145 1512 9179 1517
rect 8913 1491 9087 1494
rect 8906 1488 9087 1491
rect 9115 1511 9179 1512
rect 8709 1468 8728 1470
rect 8743 1468 8777 1470
rect 8709 1452 8789 1468
rect 8709 1446 8728 1452
rect 8425 1420 8528 1430
rect 8379 1418 8528 1420
rect 8549 1418 8584 1430
rect 8218 1416 8380 1418
rect 8230 1396 8249 1416
rect 8264 1414 8294 1416
rect 8113 1388 8154 1396
rect 8236 1392 8249 1396
rect 8301 1400 8380 1416
rect 8412 1416 8584 1418
rect 8412 1400 8491 1416
rect 8498 1414 8528 1416
rect 8076 1378 8105 1388
rect 8119 1378 8148 1388
rect 8163 1378 8193 1392
rect 8236 1378 8279 1392
rect 8301 1388 8491 1400
rect 8556 1396 8562 1416
rect 8286 1378 8316 1388
rect 8317 1378 8475 1388
rect 8479 1378 8509 1388
rect 8513 1378 8543 1392
rect 8571 1378 8584 1416
rect 8656 1430 8685 1446
rect 8699 1430 8728 1446
rect 8743 1436 8773 1452
rect 8801 1430 8807 1478
rect 8810 1472 8829 1478
rect 8844 1472 8874 1480
rect 8810 1464 8874 1472
rect 8810 1448 8890 1464
rect 8906 1457 8968 1488
rect 8984 1457 9046 1488
rect 9115 1486 9164 1511
rect 9179 1486 9209 1502
rect 9078 1472 9108 1480
rect 9115 1478 9225 1486
rect 9078 1464 9123 1472
rect 8810 1446 8829 1448
rect 8844 1446 8890 1448
rect 8810 1430 8890 1446
rect 8917 1444 8952 1457
rect 8993 1454 9030 1457
rect 8993 1452 9035 1454
rect 8922 1441 8952 1444
rect 8931 1437 8938 1441
rect 8938 1436 8939 1437
rect 8897 1430 8907 1436
rect 8656 1422 8691 1430
rect 8656 1396 8657 1422
rect 8664 1396 8691 1422
rect 8599 1378 8629 1392
rect 8656 1388 8691 1396
rect 8693 1422 8734 1430
rect 8693 1396 8708 1422
rect 8715 1396 8734 1422
rect 8798 1418 8829 1430
rect 8844 1418 8947 1430
rect 8959 1420 8985 1446
rect 9000 1441 9030 1452
rect 9062 1448 9124 1464
rect 9062 1446 9108 1448
rect 9062 1430 9124 1446
rect 9136 1430 9142 1478
rect 9145 1470 9225 1478
rect 9145 1468 9164 1470
rect 9179 1468 9213 1470
rect 9145 1452 9225 1468
rect 9145 1430 9164 1452
rect 9179 1436 9209 1452
rect 9237 1446 9243 1520
rect 9252 1446 9265 1590
rect 9005 1420 9108 1430
rect 8959 1418 9108 1420
rect 9129 1418 9164 1430
rect 8798 1416 8960 1418
rect 8810 1396 8829 1416
rect 8844 1414 8874 1416
rect 8693 1388 8734 1396
rect 8816 1392 8829 1396
rect 8881 1400 8960 1416
rect 8992 1416 9164 1418
rect 8992 1400 9071 1416
rect 9078 1414 9108 1416
rect 8656 1378 8685 1388
rect 8699 1378 8728 1388
rect 8743 1378 8773 1392
rect 8816 1378 8859 1392
rect 8881 1388 9071 1400
rect 9136 1396 9142 1416
rect 8866 1378 8896 1388
rect 8897 1378 9055 1388
rect 9059 1378 9089 1388
rect 9093 1378 9123 1392
rect 9151 1378 9164 1416
rect 9236 1430 9265 1446
rect 9236 1422 9271 1430
rect 9236 1396 9237 1422
rect 9244 1396 9271 1422
rect 9179 1378 9209 1392
rect 9236 1388 9271 1396
rect 9236 1378 9265 1388
rect -1 1372 9265 1378
rect 0 1364 9265 1372
rect 15 1334 28 1364
rect 43 1350 73 1364
rect 116 1350 159 1364
rect 166 1350 386 1364
rect 393 1350 423 1364
rect 83 1336 98 1348
rect 117 1336 130 1350
rect 198 1346 351 1350
rect 80 1334 102 1336
rect 180 1334 372 1346
rect 451 1334 464 1364
rect 479 1350 509 1364
rect 546 1334 565 1364
rect 580 1334 586 1364
rect 595 1334 608 1364
rect 623 1350 653 1364
rect 696 1350 739 1364
rect 746 1350 966 1364
rect 973 1350 1003 1364
rect 663 1336 678 1348
rect 697 1336 710 1350
rect 778 1346 931 1350
rect 660 1334 682 1336
rect 760 1334 952 1346
rect 1031 1334 1044 1364
rect 1059 1350 1089 1364
rect 1126 1334 1145 1364
rect 1160 1334 1166 1364
rect 1175 1334 1188 1364
rect 1203 1350 1233 1364
rect 1276 1350 1319 1364
rect 1326 1350 1546 1364
rect 1553 1350 1583 1364
rect 1243 1336 1258 1348
rect 1277 1336 1290 1350
rect 1358 1346 1511 1350
rect 1240 1334 1262 1336
rect 1340 1334 1532 1346
rect 1611 1334 1624 1364
rect 1639 1350 1669 1364
rect 1706 1334 1725 1364
rect 1740 1334 1746 1364
rect 1755 1334 1768 1364
rect 1783 1350 1813 1364
rect 1856 1350 1899 1364
rect 1906 1350 2126 1364
rect 2133 1350 2163 1364
rect 1823 1336 1838 1348
rect 1857 1336 1870 1350
rect 1938 1346 2091 1350
rect 1820 1334 1842 1336
rect 1920 1334 2112 1346
rect 2191 1334 2204 1364
rect 2219 1350 2249 1364
rect 2286 1334 2305 1364
rect 2320 1334 2326 1364
rect 2335 1334 2348 1364
rect 2363 1350 2393 1364
rect 2436 1350 2479 1364
rect 2486 1350 2706 1364
rect 2713 1350 2743 1364
rect 2403 1336 2418 1348
rect 2437 1336 2450 1350
rect 2518 1346 2671 1350
rect 2400 1334 2422 1336
rect 2500 1334 2692 1346
rect 2771 1334 2784 1364
rect 2799 1350 2829 1364
rect 2866 1334 2885 1364
rect 2900 1334 2906 1364
rect 2915 1334 2928 1364
rect 2943 1350 2973 1364
rect 3016 1350 3059 1364
rect 3066 1350 3286 1364
rect 3293 1350 3323 1364
rect 2983 1336 2998 1348
rect 3017 1336 3030 1350
rect 3098 1346 3251 1350
rect 2980 1334 3002 1336
rect 3080 1334 3272 1346
rect 3351 1334 3364 1364
rect 3379 1350 3409 1364
rect 3446 1334 3465 1364
rect 3480 1334 3486 1364
rect 3495 1334 3508 1364
rect 3523 1350 3553 1364
rect 3596 1350 3639 1364
rect 3646 1350 3866 1364
rect 3873 1350 3903 1364
rect 3563 1336 3578 1348
rect 3597 1336 3610 1350
rect 3678 1346 3831 1350
rect 3560 1334 3582 1336
rect 3660 1334 3852 1346
rect 3931 1334 3944 1364
rect 3959 1350 3989 1364
rect 4026 1334 4045 1364
rect 4060 1334 4066 1364
rect 4075 1334 4088 1364
rect 4103 1350 4133 1364
rect 4176 1350 4219 1364
rect 4226 1350 4446 1364
rect 4453 1350 4483 1364
rect 4143 1336 4158 1348
rect 4177 1336 4190 1350
rect 4258 1346 4411 1350
rect 4140 1334 4162 1336
rect 4240 1334 4432 1346
rect 4511 1334 4524 1364
rect 4539 1350 4569 1364
rect 4606 1334 4625 1364
rect 4640 1334 4646 1364
rect 4655 1334 4668 1364
rect 4683 1350 4713 1364
rect 4756 1350 4799 1364
rect 4806 1350 5026 1364
rect 5033 1350 5063 1364
rect 4723 1336 4738 1348
rect 4757 1336 4770 1350
rect 4838 1346 4991 1350
rect 4720 1334 4742 1336
rect 4820 1334 5012 1346
rect 5091 1334 5104 1364
rect 5119 1350 5149 1364
rect 5186 1334 5205 1364
rect 5220 1334 5226 1364
rect 5235 1334 5248 1364
rect 5263 1350 5293 1364
rect 5336 1350 5379 1364
rect 5386 1350 5606 1364
rect 5613 1350 5643 1364
rect 5303 1336 5318 1348
rect 5337 1336 5350 1350
rect 5418 1346 5571 1350
rect 5300 1334 5322 1336
rect 5400 1334 5592 1346
rect 5671 1334 5684 1364
rect 5699 1350 5729 1364
rect 5766 1334 5785 1364
rect 5800 1334 5806 1364
rect 5815 1334 5828 1364
rect 5843 1350 5873 1364
rect 5916 1350 5959 1364
rect 5966 1350 6186 1364
rect 6193 1350 6223 1364
rect 5883 1336 5898 1348
rect 5917 1336 5930 1350
rect 5998 1346 6151 1350
rect 5880 1334 5902 1336
rect 5980 1334 6172 1346
rect 6251 1334 6264 1364
rect 6279 1350 6309 1364
rect 6346 1334 6365 1364
rect 6380 1334 6386 1364
rect 6395 1334 6408 1364
rect 6423 1350 6453 1364
rect 6496 1350 6539 1364
rect 6546 1350 6766 1364
rect 6773 1350 6803 1364
rect 6463 1336 6478 1348
rect 6497 1336 6510 1350
rect 6578 1346 6731 1350
rect 6460 1334 6482 1336
rect 6560 1334 6752 1346
rect 6831 1334 6844 1364
rect 6859 1350 6889 1364
rect 6926 1334 6945 1364
rect 6960 1334 6966 1364
rect 6975 1334 6988 1364
rect 7003 1350 7033 1364
rect 7076 1350 7119 1364
rect 7126 1350 7346 1364
rect 7353 1350 7383 1364
rect 7043 1336 7058 1348
rect 7077 1336 7090 1350
rect 7158 1346 7311 1350
rect 7040 1334 7062 1336
rect 7140 1334 7332 1346
rect 7411 1334 7424 1364
rect 7439 1350 7469 1364
rect 7506 1334 7525 1364
rect 7540 1334 7546 1364
rect 7555 1334 7568 1364
rect 7583 1350 7613 1364
rect 7656 1350 7699 1364
rect 7706 1350 7926 1364
rect 7933 1350 7963 1364
rect 7623 1336 7638 1348
rect 7657 1336 7670 1350
rect 7738 1346 7891 1350
rect 7620 1334 7642 1336
rect 7720 1334 7912 1346
rect 7991 1334 8004 1364
rect 8019 1350 8049 1364
rect 8086 1334 8105 1364
rect 8120 1334 8126 1364
rect 8135 1334 8148 1364
rect 8163 1350 8193 1364
rect 8236 1350 8279 1364
rect 8286 1350 8506 1364
rect 8513 1350 8543 1364
rect 8203 1336 8218 1348
rect 8237 1336 8250 1350
rect 8318 1346 8471 1350
rect 8200 1334 8222 1336
rect 8300 1334 8492 1346
rect 8571 1334 8584 1364
rect 8599 1350 8629 1364
rect 8666 1334 8685 1364
rect 8700 1334 8706 1364
rect 8715 1334 8728 1364
rect 8743 1350 8773 1364
rect 8816 1350 8859 1364
rect 8866 1350 9086 1364
rect 9093 1350 9123 1364
rect 8783 1336 8798 1348
rect 8817 1336 8830 1350
rect 8898 1346 9051 1350
rect 8780 1334 8802 1336
rect 8880 1334 9072 1346
rect 9151 1334 9164 1364
rect 9179 1350 9209 1364
rect 9252 1334 9265 1364
rect 0 1320 9265 1334
rect 15 1250 28 1320
rect 80 1316 102 1320
rect 73 1294 102 1308
rect 155 1294 171 1308
rect 209 1304 215 1306
rect 222 1304 330 1320
rect 337 1304 343 1306
rect 351 1304 366 1320
rect 432 1314 451 1317
rect 73 1292 171 1294
rect 198 1292 366 1304
rect 381 1294 397 1308
rect 432 1295 454 1314
rect 464 1308 480 1309
rect 463 1306 480 1308
rect 464 1301 480 1306
rect 454 1294 460 1295
rect 463 1294 492 1301
rect 381 1293 492 1294
rect 381 1292 498 1293
rect 57 1284 108 1292
rect 155 1284 189 1292
rect 57 1272 82 1284
rect 89 1272 108 1284
rect 162 1282 189 1284
rect 198 1282 419 1292
rect 454 1289 460 1292
rect 162 1278 419 1282
rect 57 1264 108 1272
rect 155 1264 419 1278
rect 463 1284 498 1292
rect 9 1216 28 1250
rect 73 1256 102 1264
rect 73 1250 90 1256
rect 73 1248 107 1250
rect 155 1248 171 1264
rect 172 1254 380 1264
rect 381 1254 397 1264
rect 445 1260 460 1275
rect 463 1272 464 1284
rect 471 1272 498 1284
rect 463 1264 498 1272
rect 463 1263 492 1264
rect 183 1250 397 1254
rect 198 1248 397 1250
rect 432 1250 445 1260
rect 463 1250 480 1263
rect 432 1248 480 1250
rect 74 1244 107 1248
rect 70 1242 107 1244
rect 70 1241 137 1242
rect 70 1236 101 1241
rect 107 1236 137 1241
rect 70 1232 137 1236
rect 43 1229 137 1232
rect 43 1222 92 1229
rect 43 1216 73 1222
rect 92 1217 97 1222
rect 9 1200 89 1216
rect 101 1208 137 1229
rect 198 1224 387 1248
rect 432 1247 479 1248
rect 445 1242 479 1247
rect 213 1221 387 1224
rect 206 1218 387 1221
rect 415 1241 479 1242
rect 9 1198 28 1200
rect 43 1198 77 1200
rect 9 1182 89 1198
rect 9 1176 28 1182
rect -1 1160 28 1176
rect 43 1166 73 1182
rect 101 1160 107 1208
rect 110 1202 129 1208
rect 144 1202 174 1210
rect 110 1194 174 1202
rect 110 1178 190 1194
rect 206 1187 268 1218
rect 284 1187 346 1218
rect 415 1216 464 1241
rect 479 1216 509 1232
rect 378 1202 408 1210
rect 415 1208 525 1216
rect 378 1194 423 1202
rect 110 1176 129 1178
rect 144 1176 190 1178
rect 110 1160 190 1176
rect 217 1174 252 1187
rect 293 1184 330 1187
rect 293 1182 335 1184
rect 222 1171 252 1174
rect 231 1167 238 1171
rect 238 1166 239 1167
rect 197 1160 207 1166
rect -7 1152 34 1160
rect -7 1126 8 1152
rect 15 1126 34 1152
rect 98 1148 129 1160
rect 144 1148 247 1160
rect 259 1150 285 1176
rect 300 1171 330 1182
rect 362 1178 424 1194
rect 362 1176 408 1178
rect 362 1160 424 1176
rect 436 1160 442 1208
rect 445 1200 525 1208
rect 445 1198 464 1200
rect 479 1198 513 1200
rect 445 1182 525 1198
rect 445 1160 464 1182
rect 479 1166 509 1182
rect 537 1176 543 1250
rect 546 1176 565 1320
rect 580 1176 586 1320
rect 595 1250 608 1320
rect 660 1316 682 1320
rect 653 1294 682 1308
rect 735 1294 751 1308
rect 789 1304 795 1306
rect 802 1304 910 1320
rect 917 1304 923 1306
rect 931 1304 946 1320
rect 1012 1314 1031 1317
rect 653 1292 751 1294
rect 778 1292 946 1304
rect 961 1294 977 1308
rect 1012 1295 1034 1314
rect 1044 1308 1060 1309
rect 1043 1306 1060 1308
rect 1044 1301 1060 1306
rect 1034 1294 1040 1295
rect 1043 1294 1072 1301
rect 961 1293 1072 1294
rect 961 1292 1078 1293
rect 637 1284 688 1292
rect 735 1284 769 1292
rect 637 1272 662 1284
rect 669 1272 688 1284
rect 742 1282 769 1284
rect 778 1282 999 1292
rect 1034 1289 1040 1292
rect 742 1278 999 1282
rect 637 1264 688 1272
rect 735 1264 999 1278
rect 1043 1284 1078 1292
rect 589 1216 608 1250
rect 653 1256 682 1264
rect 653 1250 670 1256
rect 653 1248 687 1250
rect 735 1248 751 1264
rect 752 1254 960 1264
rect 961 1254 977 1264
rect 1025 1260 1040 1275
rect 1043 1272 1044 1284
rect 1051 1272 1078 1284
rect 1043 1264 1078 1272
rect 1043 1263 1072 1264
rect 763 1250 977 1254
rect 778 1248 977 1250
rect 1012 1250 1025 1260
rect 1043 1250 1060 1263
rect 1012 1248 1060 1250
rect 654 1244 687 1248
rect 650 1242 687 1244
rect 650 1241 717 1242
rect 650 1236 681 1241
rect 687 1236 717 1241
rect 650 1232 717 1236
rect 623 1229 717 1232
rect 623 1222 672 1229
rect 623 1216 653 1222
rect 672 1217 677 1222
rect 589 1200 669 1216
rect 681 1208 717 1229
rect 778 1224 967 1248
rect 1012 1247 1059 1248
rect 1025 1242 1059 1247
rect 793 1221 967 1224
rect 786 1218 967 1221
rect 995 1241 1059 1242
rect 589 1198 608 1200
rect 623 1198 657 1200
rect 589 1182 669 1198
rect 589 1176 608 1182
rect 305 1150 408 1160
rect 259 1148 408 1150
rect 429 1148 464 1160
rect 98 1146 260 1148
rect 110 1126 129 1146
rect 144 1144 174 1146
rect -7 1118 34 1126
rect 116 1122 129 1126
rect 181 1130 260 1146
rect 292 1146 464 1148
rect 292 1130 371 1146
rect 378 1144 408 1146
rect -1 1108 28 1118
rect 43 1108 73 1122
rect 116 1108 159 1122
rect 181 1118 371 1130
rect 436 1126 442 1146
rect 166 1108 196 1118
rect 197 1108 355 1118
rect 359 1108 389 1118
rect 393 1108 423 1122
rect 451 1108 464 1146
rect 536 1160 565 1176
rect 579 1160 608 1176
rect 623 1166 653 1182
rect 681 1160 687 1208
rect 690 1202 709 1208
rect 724 1202 754 1210
rect 690 1194 754 1202
rect 690 1178 770 1194
rect 786 1187 848 1218
rect 864 1187 926 1218
rect 995 1216 1044 1241
rect 1059 1216 1089 1232
rect 958 1202 988 1210
rect 995 1208 1105 1216
rect 958 1194 1003 1202
rect 690 1176 709 1178
rect 724 1176 770 1178
rect 690 1160 770 1176
rect 797 1174 832 1187
rect 873 1184 910 1187
rect 873 1182 915 1184
rect 802 1171 832 1174
rect 811 1167 818 1171
rect 818 1166 819 1167
rect 777 1160 787 1166
rect 536 1152 571 1160
rect 536 1126 537 1152
rect 544 1126 571 1152
rect 479 1108 509 1122
rect 536 1118 571 1126
rect 573 1152 614 1160
rect 573 1126 588 1152
rect 595 1126 614 1152
rect 678 1148 709 1160
rect 724 1148 827 1160
rect 839 1150 865 1176
rect 880 1171 910 1182
rect 942 1178 1004 1194
rect 942 1176 988 1178
rect 942 1160 1004 1176
rect 1016 1160 1022 1208
rect 1025 1200 1105 1208
rect 1025 1198 1044 1200
rect 1059 1198 1093 1200
rect 1025 1182 1105 1198
rect 1025 1160 1044 1182
rect 1059 1166 1089 1182
rect 1117 1176 1123 1250
rect 1126 1176 1145 1320
rect 1160 1176 1166 1320
rect 1175 1250 1188 1320
rect 1240 1316 1262 1320
rect 1233 1294 1262 1308
rect 1315 1294 1331 1308
rect 1369 1304 1375 1306
rect 1382 1304 1490 1320
rect 1497 1304 1503 1306
rect 1511 1304 1526 1320
rect 1592 1314 1611 1317
rect 1233 1292 1331 1294
rect 1358 1292 1526 1304
rect 1541 1294 1557 1308
rect 1592 1295 1614 1314
rect 1624 1308 1640 1309
rect 1623 1306 1640 1308
rect 1624 1301 1640 1306
rect 1614 1294 1620 1295
rect 1623 1294 1652 1301
rect 1541 1293 1652 1294
rect 1541 1292 1658 1293
rect 1217 1284 1268 1292
rect 1315 1284 1349 1292
rect 1217 1272 1242 1284
rect 1249 1272 1268 1284
rect 1322 1282 1349 1284
rect 1358 1282 1579 1292
rect 1614 1289 1620 1292
rect 1322 1278 1579 1282
rect 1217 1264 1268 1272
rect 1315 1264 1579 1278
rect 1623 1284 1658 1292
rect 1169 1216 1188 1250
rect 1233 1256 1262 1264
rect 1233 1250 1250 1256
rect 1233 1248 1267 1250
rect 1315 1248 1331 1264
rect 1332 1254 1540 1264
rect 1541 1254 1557 1264
rect 1605 1260 1620 1275
rect 1623 1272 1624 1284
rect 1631 1272 1658 1284
rect 1623 1264 1658 1272
rect 1623 1263 1652 1264
rect 1343 1250 1557 1254
rect 1358 1248 1557 1250
rect 1592 1250 1605 1260
rect 1623 1250 1640 1263
rect 1592 1248 1640 1250
rect 1234 1244 1267 1248
rect 1230 1242 1267 1244
rect 1230 1241 1297 1242
rect 1230 1236 1261 1241
rect 1267 1236 1297 1241
rect 1230 1232 1297 1236
rect 1203 1229 1297 1232
rect 1203 1222 1252 1229
rect 1203 1216 1233 1222
rect 1252 1217 1257 1222
rect 1169 1200 1249 1216
rect 1261 1208 1297 1229
rect 1358 1224 1547 1248
rect 1592 1247 1639 1248
rect 1605 1242 1639 1247
rect 1373 1221 1547 1224
rect 1366 1218 1547 1221
rect 1575 1241 1639 1242
rect 1169 1198 1188 1200
rect 1203 1198 1237 1200
rect 1169 1182 1249 1198
rect 1169 1176 1188 1182
rect 885 1150 988 1160
rect 839 1148 988 1150
rect 1009 1148 1044 1160
rect 678 1146 840 1148
rect 690 1126 709 1146
rect 724 1144 754 1146
rect 573 1118 614 1126
rect 696 1122 709 1126
rect 761 1130 840 1146
rect 872 1146 1044 1148
rect 872 1130 951 1146
rect 958 1144 988 1146
rect 536 1108 565 1118
rect 579 1108 608 1118
rect 623 1108 653 1122
rect 696 1108 739 1122
rect 761 1118 951 1130
rect 1016 1126 1022 1146
rect 746 1108 776 1118
rect 777 1108 935 1118
rect 939 1108 969 1118
rect 973 1108 1003 1122
rect 1031 1108 1044 1146
rect 1116 1160 1145 1176
rect 1159 1160 1188 1176
rect 1203 1166 1233 1182
rect 1261 1160 1267 1208
rect 1270 1202 1289 1208
rect 1304 1202 1334 1210
rect 1270 1194 1334 1202
rect 1270 1178 1350 1194
rect 1366 1187 1428 1218
rect 1444 1187 1506 1218
rect 1575 1216 1624 1241
rect 1639 1216 1669 1232
rect 1538 1202 1568 1210
rect 1575 1208 1685 1216
rect 1538 1194 1583 1202
rect 1270 1176 1289 1178
rect 1304 1176 1350 1178
rect 1270 1160 1350 1176
rect 1377 1174 1412 1187
rect 1453 1184 1490 1187
rect 1453 1182 1495 1184
rect 1382 1171 1412 1174
rect 1391 1167 1398 1171
rect 1398 1166 1399 1167
rect 1357 1160 1367 1166
rect 1116 1152 1151 1160
rect 1116 1126 1117 1152
rect 1124 1126 1151 1152
rect 1059 1108 1089 1122
rect 1116 1118 1151 1126
rect 1153 1152 1194 1160
rect 1153 1126 1168 1152
rect 1175 1126 1194 1152
rect 1258 1148 1289 1160
rect 1304 1148 1407 1160
rect 1419 1150 1445 1176
rect 1460 1171 1490 1182
rect 1522 1178 1584 1194
rect 1522 1176 1568 1178
rect 1522 1160 1584 1176
rect 1596 1160 1602 1208
rect 1605 1200 1685 1208
rect 1605 1198 1624 1200
rect 1639 1198 1673 1200
rect 1605 1182 1685 1198
rect 1605 1160 1624 1182
rect 1639 1166 1669 1182
rect 1697 1176 1703 1250
rect 1706 1176 1725 1320
rect 1740 1176 1746 1320
rect 1755 1250 1768 1320
rect 1820 1316 1842 1320
rect 1813 1294 1842 1308
rect 1895 1294 1911 1308
rect 1949 1304 1955 1306
rect 1962 1304 2070 1320
rect 2077 1304 2083 1306
rect 2091 1304 2106 1320
rect 2172 1314 2191 1317
rect 1813 1292 1911 1294
rect 1938 1292 2106 1304
rect 2121 1294 2137 1308
rect 2172 1295 2194 1314
rect 2204 1308 2220 1309
rect 2203 1306 2220 1308
rect 2204 1301 2220 1306
rect 2194 1294 2200 1295
rect 2203 1294 2232 1301
rect 2121 1293 2232 1294
rect 2121 1292 2238 1293
rect 1797 1284 1848 1292
rect 1895 1284 1929 1292
rect 1797 1272 1822 1284
rect 1829 1272 1848 1284
rect 1902 1282 1929 1284
rect 1938 1282 2159 1292
rect 2194 1289 2200 1292
rect 1902 1278 2159 1282
rect 1797 1264 1848 1272
rect 1895 1264 2159 1278
rect 2203 1284 2238 1292
rect 1749 1216 1768 1250
rect 1813 1256 1842 1264
rect 1813 1250 1830 1256
rect 1813 1248 1847 1250
rect 1895 1248 1911 1264
rect 1912 1254 2120 1264
rect 2121 1254 2137 1264
rect 2185 1260 2200 1275
rect 2203 1272 2204 1284
rect 2211 1272 2238 1284
rect 2203 1264 2238 1272
rect 2203 1263 2232 1264
rect 1923 1250 2137 1254
rect 1938 1248 2137 1250
rect 2172 1250 2185 1260
rect 2203 1250 2220 1263
rect 2172 1248 2220 1250
rect 1814 1244 1847 1248
rect 1810 1242 1847 1244
rect 1810 1241 1877 1242
rect 1810 1236 1841 1241
rect 1847 1236 1877 1241
rect 1810 1232 1877 1236
rect 1783 1229 1877 1232
rect 1783 1222 1832 1229
rect 1783 1216 1813 1222
rect 1832 1217 1837 1222
rect 1749 1200 1829 1216
rect 1841 1208 1877 1229
rect 1938 1224 2127 1248
rect 2172 1247 2219 1248
rect 2185 1242 2219 1247
rect 1953 1221 2127 1224
rect 1946 1218 2127 1221
rect 2155 1241 2219 1242
rect 1749 1198 1768 1200
rect 1783 1198 1817 1200
rect 1749 1182 1829 1198
rect 1749 1176 1768 1182
rect 1465 1150 1568 1160
rect 1419 1148 1568 1150
rect 1589 1148 1624 1160
rect 1258 1146 1420 1148
rect 1270 1126 1289 1146
rect 1304 1144 1334 1146
rect 1153 1118 1194 1126
rect 1276 1122 1289 1126
rect 1341 1130 1420 1146
rect 1452 1146 1624 1148
rect 1452 1130 1531 1146
rect 1538 1144 1568 1146
rect 1116 1108 1145 1118
rect 1159 1108 1188 1118
rect 1203 1108 1233 1122
rect 1276 1108 1319 1122
rect 1341 1118 1531 1130
rect 1596 1126 1602 1146
rect 1326 1108 1356 1118
rect 1357 1108 1515 1118
rect 1519 1108 1549 1118
rect 1553 1108 1583 1122
rect 1611 1108 1624 1146
rect 1696 1160 1725 1176
rect 1739 1160 1768 1176
rect 1783 1166 1813 1182
rect 1841 1160 1847 1208
rect 1850 1202 1869 1208
rect 1884 1202 1914 1210
rect 1850 1194 1914 1202
rect 1850 1178 1930 1194
rect 1946 1187 2008 1218
rect 2024 1187 2086 1218
rect 2155 1216 2204 1241
rect 2219 1216 2249 1232
rect 2118 1202 2148 1210
rect 2155 1208 2265 1216
rect 2118 1194 2163 1202
rect 1850 1176 1869 1178
rect 1884 1176 1930 1178
rect 1850 1160 1930 1176
rect 1957 1174 1992 1187
rect 2033 1184 2070 1187
rect 2033 1182 2075 1184
rect 1962 1171 1992 1174
rect 1971 1167 1978 1171
rect 1978 1166 1979 1167
rect 1937 1160 1947 1166
rect 1696 1152 1731 1160
rect 1696 1126 1697 1152
rect 1704 1126 1731 1152
rect 1639 1108 1669 1122
rect 1696 1118 1731 1126
rect 1733 1152 1774 1160
rect 1733 1126 1748 1152
rect 1755 1126 1774 1152
rect 1838 1148 1869 1160
rect 1884 1148 1987 1160
rect 1999 1150 2025 1176
rect 2040 1171 2070 1182
rect 2102 1178 2164 1194
rect 2102 1176 2148 1178
rect 2102 1160 2164 1176
rect 2176 1160 2182 1208
rect 2185 1200 2265 1208
rect 2185 1198 2204 1200
rect 2219 1198 2253 1200
rect 2185 1182 2265 1198
rect 2185 1160 2204 1182
rect 2219 1166 2249 1182
rect 2277 1176 2283 1250
rect 2286 1176 2305 1320
rect 2320 1176 2326 1320
rect 2335 1250 2348 1320
rect 2400 1316 2422 1320
rect 2393 1294 2422 1308
rect 2475 1294 2491 1308
rect 2529 1304 2535 1306
rect 2542 1304 2650 1320
rect 2657 1304 2663 1306
rect 2671 1304 2686 1320
rect 2752 1314 2771 1317
rect 2393 1292 2491 1294
rect 2518 1292 2686 1304
rect 2701 1294 2717 1308
rect 2752 1295 2774 1314
rect 2784 1308 2800 1309
rect 2783 1306 2800 1308
rect 2784 1301 2800 1306
rect 2774 1294 2780 1295
rect 2783 1294 2812 1301
rect 2701 1293 2812 1294
rect 2701 1292 2818 1293
rect 2377 1284 2428 1292
rect 2475 1284 2509 1292
rect 2377 1272 2402 1284
rect 2409 1272 2428 1284
rect 2482 1282 2509 1284
rect 2518 1282 2739 1292
rect 2774 1289 2780 1292
rect 2482 1278 2739 1282
rect 2377 1264 2428 1272
rect 2475 1264 2739 1278
rect 2783 1284 2818 1292
rect 2329 1216 2348 1250
rect 2393 1256 2422 1264
rect 2393 1250 2410 1256
rect 2393 1248 2427 1250
rect 2475 1248 2491 1264
rect 2492 1254 2700 1264
rect 2701 1254 2717 1264
rect 2765 1260 2780 1275
rect 2783 1272 2784 1284
rect 2791 1272 2818 1284
rect 2783 1264 2818 1272
rect 2783 1263 2812 1264
rect 2503 1250 2717 1254
rect 2518 1248 2717 1250
rect 2752 1250 2765 1260
rect 2783 1250 2800 1263
rect 2752 1248 2800 1250
rect 2394 1244 2427 1248
rect 2390 1242 2427 1244
rect 2390 1241 2457 1242
rect 2390 1236 2421 1241
rect 2427 1236 2457 1241
rect 2390 1232 2457 1236
rect 2363 1229 2457 1232
rect 2363 1222 2412 1229
rect 2363 1216 2393 1222
rect 2412 1217 2417 1222
rect 2329 1200 2409 1216
rect 2421 1208 2457 1229
rect 2518 1224 2707 1248
rect 2752 1247 2799 1248
rect 2765 1242 2799 1247
rect 2533 1221 2707 1224
rect 2526 1218 2707 1221
rect 2735 1241 2799 1242
rect 2329 1198 2348 1200
rect 2363 1198 2397 1200
rect 2329 1182 2409 1198
rect 2329 1176 2348 1182
rect 2045 1150 2148 1160
rect 1999 1148 2148 1150
rect 2169 1148 2204 1160
rect 1838 1146 2000 1148
rect 1850 1126 1869 1146
rect 1884 1144 1914 1146
rect 1733 1118 1774 1126
rect 1856 1122 1869 1126
rect 1921 1130 2000 1146
rect 2032 1146 2204 1148
rect 2032 1130 2111 1146
rect 2118 1144 2148 1146
rect 1696 1108 1725 1118
rect 1739 1108 1768 1118
rect 1783 1108 1813 1122
rect 1856 1108 1899 1122
rect 1921 1118 2111 1130
rect 2176 1126 2182 1146
rect 1906 1108 1936 1118
rect 1937 1108 2095 1118
rect 2099 1108 2129 1118
rect 2133 1108 2163 1122
rect 2191 1108 2204 1146
rect 2276 1160 2305 1176
rect 2319 1160 2348 1176
rect 2363 1166 2393 1182
rect 2421 1160 2427 1208
rect 2430 1202 2449 1208
rect 2464 1202 2494 1210
rect 2430 1194 2494 1202
rect 2430 1178 2510 1194
rect 2526 1187 2588 1218
rect 2604 1187 2666 1218
rect 2735 1216 2784 1241
rect 2799 1216 2829 1232
rect 2698 1202 2728 1210
rect 2735 1208 2845 1216
rect 2698 1194 2743 1202
rect 2430 1176 2449 1178
rect 2464 1176 2510 1178
rect 2430 1160 2510 1176
rect 2537 1174 2572 1187
rect 2613 1184 2650 1187
rect 2613 1182 2655 1184
rect 2542 1171 2572 1174
rect 2551 1167 2558 1171
rect 2558 1166 2559 1167
rect 2517 1160 2527 1166
rect 2276 1152 2311 1160
rect 2276 1126 2277 1152
rect 2284 1126 2311 1152
rect 2219 1108 2249 1122
rect 2276 1118 2311 1126
rect 2313 1152 2354 1160
rect 2313 1126 2328 1152
rect 2335 1126 2354 1152
rect 2418 1148 2449 1160
rect 2464 1148 2567 1160
rect 2579 1150 2605 1176
rect 2620 1171 2650 1182
rect 2682 1178 2744 1194
rect 2682 1176 2728 1178
rect 2682 1160 2744 1176
rect 2756 1160 2762 1208
rect 2765 1200 2845 1208
rect 2765 1198 2784 1200
rect 2799 1198 2833 1200
rect 2765 1182 2845 1198
rect 2765 1160 2784 1182
rect 2799 1166 2829 1182
rect 2857 1176 2863 1250
rect 2866 1176 2885 1320
rect 2900 1176 2906 1320
rect 2915 1250 2928 1320
rect 2980 1316 3002 1320
rect 2973 1294 3002 1308
rect 3055 1294 3071 1308
rect 3109 1304 3115 1306
rect 3122 1304 3230 1320
rect 3237 1304 3243 1306
rect 3251 1304 3266 1320
rect 3332 1314 3351 1317
rect 2973 1292 3071 1294
rect 3098 1292 3266 1304
rect 3281 1294 3297 1308
rect 3332 1295 3354 1314
rect 3364 1308 3380 1309
rect 3363 1306 3380 1308
rect 3364 1301 3380 1306
rect 3354 1294 3360 1295
rect 3363 1294 3392 1301
rect 3281 1293 3392 1294
rect 3281 1292 3398 1293
rect 2957 1284 3008 1292
rect 3055 1284 3089 1292
rect 2957 1272 2982 1284
rect 2989 1272 3008 1284
rect 3062 1282 3089 1284
rect 3098 1282 3319 1292
rect 3354 1289 3360 1292
rect 3062 1278 3319 1282
rect 2957 1264 3008 1272
rect 3055 1264 3319 1278
rect 3363 1284 3398 1292
rect 2909 1216 2928 1250
rect 2973 1256 3002 1264
rect 2973 1250 2990 1256
rect 2973 1248 3007 1250
rect 3055 1248 3071 1264
rect 3072 1254 3280 1264
rect 3281 1254 3297 1264
rect 3345 1260 3360 1275
rect 3363 1272 3364 1284
rect 3371 1272 3398 1284
rect 3363 1264 3398 1272
rect 3363 1263 3392 1264
rect 3083 1250 3297 1254
rect 3098 1248 3297 1250
rect 3332 1250 3345 1260
rect 3363 1250 3380 1263
rect 3332 1248 3380 1250
rect 2974 1244 3007 1248
rect 2970 1242 3007 1244
rect 2970 1241 3037 1242
rect 2970 1236 3001 1241
rect 3007 1236 3037 1241
rect 2970 1232 3037 1236
rect 2943 1229 3037 1232
rect 2943 1222 2992 1229
rect 2943 1216 2973 1222
rect 2992 1217 2997 1222
rect 2909 1200 2989 1216
rect 3001 1208 3037 1229
rect 3098 1224 3287 1248
rect 3332 1247 3379 1248
rect 3345 1242 3379 1247
rect 3113 1221 3287 1224
rect 3106 1218 3287 1221
rect 3315 1241 3379 1242
rect 2909 1198 2928 1200
rect 2943 1198 2977 1200
rect 2909 1182 2989 1198
rect 2909 1176 2928 1182
rect 2625 1150 2728 1160
rect 2579 1148 2728 1150
rect 2749 1148 2784 1160
rect 2418 1146 2580 1148
rect 2430 1126 2449 1146
rect 2464 1144 2494 1146
rect 2313 1118 2354 1126
rect 2436 1122 2449 1126
rect 2501 1130 2580 1146
rect 2612 1146 2784 1148
rect 2612 1130 2691 1146
rect 2698 1144 2728 1146
rect 2276 1108 2305 1118
rect 2319 1108 2348 1118
rect 2363 1108 2393 1122
rect 2436 1108 2479 1122
rect 2501 1118 2691 1130
rect 2756 1126 2762 1146
rect 2486 1108 2516 1118
rect 2517 1108 2675 1118
rect 2679 1108 2709 1118
rect 2713 1108 2743 1122
rect 2771 1108 2784 1146
rect 2856 1160 2885 1176
rect 2899 1160 2928 1176
rect 2943 1166 2973 1182
rect 3001 1160 3007 1208
rect 3010 1202 3029 1208
rect 3044 1202 3074 1210
rect 3010 1194 3074 1202
rect 3010 1178 3090 1194
rect 3106 1187 3168 1218
rect 3184 1187 3246 1218
rect 3315 1216 3364 1241
rect 3379 1216 3409 1232
rect 3278 1202 3308 1210
rect 3315 1208 3425 1216
rect 3278 1194 3323 1202
rect 3010 1176 3029 1178
rect 3044 1176 3090 1178
rect 3010 1160 3090 1176
rect 3117 1174 3152 1187
rect 3193 1184 3230 1187
rect 3193 1182 3235 1184
rect 3122 1171 3152 1174
rect 3131 1167 3138 1171
rect 3138 1166 3139 1167
rect 3097 1160 3107 1166
rect 2856 1152 2891 1160
rect 2856 1126 2857 1152
rect 2864 1126 2891 1152
rect 2799 1108 2829 1122
rect 2856 1118 2891 1126
rect 2893 1152 2934 1160
rect 2893 1126 2908 1152
rect 2915 1126 2934 1152
rect 2998 1148 3029 1160
rect 3044 1148 3147 1160
rect 3159 1150 3185 1176
rect 3200 1171 3230 1182
rect 3262 1178 3324 1194
rect 3262 1176 3308 1178
rect 3262 1160 3324 1176
rect 3336 1160 3342 1208
rect 3345 1200 3425 1208
rect 3345 1198 3364 1200
rect 3379 1198 3413 1200
rect 3345 1182 3425 1198
rect 3345 1160 3364 1182
rect 3379 1166 3409 1182
rect 3437 1176 3443 1250
rect 3446 1176 3465 1320
rect 3480 1176 3486 1320
rect 3495 1250 3508 1320
rect 3560 1316 3582 1320
rect 3553 1294 3582 1308
rect 3635 1294 3651 1308
rect 3689 1304 3695 1306
rect 3702 1304 3810 1320
rect 3817 1304 3823 1306
rect 3831 1304 3846 1320
rect 3912 1314 3931 1317
rect 3553 1292 3651 1294
rect 3678 1292 3846 1304
rect 3861 1294 3877 1308
rect 3912 1295 3934 1314
rect 3944 1308 3960 1309
rect 3943 1306 3960 1308
rect 3944 1301 3960 1306
rect 3934 1294 3940 1295
rect 3943 1294 3972 1301
rect 3861 1293 3972 1294
rect 3861 1292 3978 1293
rect 3537 1284 3588 1292
rect 3635 1284 3669 1292
rect 3537 1272 3562 1284
rect 3569 1272 3588 1284
rect 3642 1282 3669 1284
rect 3678 1282 3899 1292
rect 3934 1289 3940 1292
rect 3642 1278 3899 1282
rect 3537 1264 3588 1272
rect 3635 1264 3899 1278
rect 3943 1284 3978 1292
rect 3489 1216 3508 1250
rect 3553 1256 3582 1264
rect 3553 1250 3570 1256
rect 3553 1248 3587 1250
rect 3635 1248 3651 1264
rect 3652 1254 3860 1264
rect 3861 1254 3877 1264
rect 3925 1260 3940 1275
rect 3943 1272 3944 1284
rect 3951 1272 3978 1284
rect 3943 1264 3978 1272
rect 3943 1263 3972 1264
rect 3663 1250 3877 1254
rect 3678 1248 3877 1250
rect 3912 1250 3925 1260
rect 3943 1250 3960 1263
rect 3912 1248 3960 1250
rect 3554 1244 3587 1248
rect 3550 1242 3587 1244
rect 3550 1241 3617 1242
rect 3550 1236 3581 1241
rect 3587 1236 3617 1241
rect 3550 1232 3617 1236
rect 3523 1229 3617 1232
rect 3523 1222 3572 1229
rect 3523 1216 3553 1222
rect 3572 1217 3577 1222
rect 3489 1200 3569 1216
rect 3581 1208 3617 1229
rect 3678 1224 3867 1248
rect 3912 1247 3959 1248
rect 3925 1242 3959 1247
rect 3693 1221 3867 1224
rect 3686 1218 3867 1221
rect 3895 1241 3959 1242
rect 3489 1198 3508 1200
rect 3523 1198 3557 1200
rect 3489 1182 3569 1198
rect 3489 1176 3508 1182
rect 3205 1150 3308 1160
rect 3159 1148 3308 1150
rect 3329 1148 3364 1160
rect 2998 1146 3160 1148
rect 3010 1126 3029 1146
rect 3044 1144 3074 1146
rect 2893 1118 2934 1126
rect 3016 1122 3029 1126
rect 3081 1130 3160 1146
rect 3192 1146 3364 1148
rect 3192 1130 3271 1146
rect 3278 1144 3308 1146
rect 2856 1108 2885 1118
rect 2899 1108 2928 1118
rect 2943 1108 2973 1122
rect 3016 1108 3059 1122
rect 3081 1118 3271 1130
rect 3336 1126 3342 1146
rect 3066 1108 3096 1118
rect 3097 1108 3255 1118
rect 3259 1108 3289 1118
rect 3293 1108 3323 1122
rect 3351 1108 3364 1146
rect 3436 1160 3465 1176
rect 3479 1160 3508 1176
rect 3523 1166 3553 1182
rect 3581 1160 3587 1208
rect 3590 1202 3609 1208
rect 3624 1202 3654 1210
rect 3590 1194 3654 1202
rect 3590 1178 3670 1194
rect 3686 1187 3748 1218
rect 3764 1187 3826 1218
rect 3895 1216 3944 1241
rect 3959 1216 3989 1232
rect 3858 1202 3888 1210
rect 3895 1208 4005 1216
rect 3858 1194 3903 1202
rect 3590 1176 3609 1178
rect 3624 1176 3670 1178
rect 3590 1160 3670 1176
rect 3697 1174 3732 1187
rect 3773 1184 3810 1187
rect 3773 1182 3815 1184
rect 3702 1171 3732 1174
rect 3711 1167 3718 1171
rect 3718 1166 3719 1167
rect 3677 1160 3687 1166
rect 3436 1152 3471 1160
rect 3436 1126 3437 1152
rect 3444 1126 3471 1152
rect 3379 1108 3409 1122
rect 3436 1118 3471 1126
rect 3473 1152 3514 1160
rect 3473 1126 3488 1152
rect 3495 1126 3514 1152
rect 3578 1148 3609 1160
rect 3624 1148 3727 1160
rect 3739 1150 3765 1176
rect 3780 1171 3810 1182
rect 3842 1178 3904 1194
rect 3842 1176 3888 1178
rect 3842 1160 3904 1176
rect 3916 1160 3922 1208
rect 3925 1200 4005 1208
rect 3925 1198 3944 1200
rect 3959 1198 3993 1200
rect 3925 1182 4005 1198
rect 3925 1160 3944 1182
rect 3959 1166 3989 1182
rect 4017 1176 4023 1250
rect 4026 1176 4045 1320
rect 4060 1176 4066 1320
rect 4075 1250 4088 1320
rect 4140 1316 4162 1320
rect 4133 1294 4162 1308
rect 4215 1294 4231 1308
rect 4269 1304 4275 1306
rect 4282 1304 4390 1320
rect 4397 1304 4403 1306
rect 4411 1304 4426 1320
rect 4492 1314 4511 1317
rect 4133 1292 4231 1294
rect 4258 1292 4426 1304
rect 4441 1294 4457 1308
rect 4492 1295 4514 1314
rect 4524 1308 4540 1309
rect 4523 1306 4540 1308
rect 4524 1301 4540 1306
rect 4514 1294 4520 1295
rect 4523 1294 4552 1301
rect 4441 1293 4552 1294
rect 4441 1292 4558 1293
rect 4117 1284 4168 1292
rect 4215 1284 4249 1292
rect 4117 1272 4142 1284
rect 4149 1272 4168 1284
rect 4222 1282 4249 1284
rect 4258 1282 4479 1292
rect 4514 1289 4520 1292
rect 4222 1278 4479 1282
rect 4117 1264 4168 1272
rect 4215 1264 4479 1278
rect 4523 1284 4558 1292
rect 4069 1216 4088 1250
rect 4133 1256 4162 1264
rect 4133 1250 4150 1256
rect 4133 1248 4167 1250
rect 4215 1248 4231 1264
rect 4232 1254 4440 1264
rect 4441 1254 4457 1264
rect 4505 1260 4520 1275
rect 4523 1272 4524 1284
rect 4531 1272 4558 1284
rect 4523 1264 4558 1272
rect 4523 1263 4552 1264
rect 4243 1250 4457 1254
rect 4258 1248 4457 1250
rect 4492 1250 4505 1260
rect 4523 1250 4540 1263
rect 4492 1248 4540 1250
rect 4134 1244 4167 1248
rect 4130 1242 4167 1244
rect 4130 1241 4197 1242
rect 4130 1236 4161 1241
rect 4167 1236 4197 1241
rect 4130 1232 4197 1236
rect 4103 1229 4197 1232
rect 4103 1222 4152 1229
rect 4103 1216 4133 1222
rect 4152 1217 4157 1222
rect 4069 1200 4149 1216
rect 4161 1208 4197 1229
rect 4258 1224 4447 1248
rect 4492 1247 4539 1248
rect 4505 1242 4539 1247
rect 4273 1221 4447 1224
rect 4266 1218 4447 1221
rect 4475 1241 4539 1242
rect 4069 1198 4088 1200
rect 4103 1198 4137 1200
rect 4069 1182 4149 1198
rect 4069 1176 4088 1182
rect 3785 1150 3888 1160
rect 3739 1148 3888 1150
rect 3909 1148 3944 1160
rect 3578 1146 3740 1148
rect 3590 1126 3609 1146
rect 3624 1144 3654 1146
rect 3473 1118 3514 1126
rect 3596 1122 3609 1126
rect 3661 1130 3740 1146
rect 3772 1146 3944 1148
rect 3772 1130 3851 1146
rect 3858 1144 3888 1146
rect 3436 1108 3465 1118
rect 3479 1108 3508 1118
rect 3523 1108 3553 1122
rect 3596 1108 3639 1122
rect 3661 1118 3851 1130
rect 3916 1126 3922 1146
rect 3646 1108 3676 1118
rect 3677 1108 3835 1118
rect 3839 1108 3869 1118
rect 3873 1108 3903 1122
rect 3931 1108 3944 1146
rect 4016 1160 4045 1176
rect 4059 1160 4088 1176
rect 4103 1166 4133 1182
rect 4161 1160 4167 1208
rect 4170 1202 4189 1208
rect 4204 1202 4234 1210
rect 4170 1194 4234 1202
rect 4170 1178 4250 1194
rect 4266 1187 4328 1218
rect 4344 1187 4406 1218
rect 4475 1216 4524 1241
rect 4539 1216 4569 1232
rect 4438 1202 4468 1210
rect 4475 1208 4585 1216
rect 4438 1194 4483 1202
rect 4170 1176 4189 1178
rect 4204 1176 4250 1178
rect 4170 1160 4250 1176
rect 4277 1174 4312 1187
rect 4353 1184 4390 1187
rect 4353 1182 4395 1184
rect 4282 1171 4312 1174
rect 4291 1167 4298 1171
rect 4298 1166 4299 1167
rect 4257 1160 4267 1166
rect 4016 1152 4051 1160
rect 4016 1126 4017 1152
rect 4024 1126 4051 1152
rect 3959 1108 3989 1122
rect 4016 1118 4051 1126
rect 4053 1152 4094 1160
rect 4053 1126 4068 1152
rect 4075 1126 4094 1152
rect 4158 1148 4189 1160
rect 4204 1148 4307 1160
rect 4319 1150 4345 1176
rect 4360 1171 4390 1182
rect 4422 1178 4484 1194
rect 4422 1176 4468 1178
rect 4422 1160 4484 1176
rect 4496 1160 4502 1208
rect 4505 1200 4585 1208
rect 4505 1198 4524 1200
rect 4539 1198 4573 1200
rect 4505 1182 4585 1198
rect 4505 1160 4524 1182
rect 4539 1166 4569 1182
rect 4597 1176 4603 1250
rect 4606 1176 4625 1320
rect 4640 1176 4646 1320
rect 4655 1250 4668 1320
rect 4720 1316 4742 1320
rect 4713 1294 4742 1308
rect 4795 1294 4811 1308
rect 4849 1304 4855 1306
rect 4862 1304 4970 1320
rect 4977 1304 4983 1306
rect 4991 1304 5006 1320
rect 5072 1314 5091 1317
rect 4713 1292 4811 1294
rect 4838 1292 5006 1304
rect 5021 1294 5037 1308
rect 5072 1295 5094 1314
rect 5104 1308 5120 1309
rect 5103 1306 5120 1308
rect 5104 1301 5120 1306
rect 5094 1294 5100 1295
rect 5103 1294 5132 1301
rect 5021 1293 5132 1294
rect 5021 1292 5138 1293
rect 4697 1284 4748 1292
rect 4795 1284 4829 1292
rect 4697 1272 4722 1284
rect 4729 1272 4748 1284
rect 4802 1282 4829 1284
rect 4838 1282 5059 1292
rect 5094 1289 5100 1292
rect 4802 1278 5059 1282
rect 4697 1264 4748 1272
rect 4795 1264 5059 1278
rect 5103 1284 5138 1292
rect 4649 1216 4668 1250
rect 4713 1256 4742 1264
rect 4713 1250 4730 1256
rect 4713 1248 4747 1250
rect 4795 1248 4811 1264
rect 4812 1254 5020 1264
rect 5021 1254 5037 1264
rect 5085 1260 5100 1275
rect 5103 1272 5104 1284
rect 5111 1272 5138 1284
rect 5103 1264 5138 1272
rect 5103 1263 5132 1264
rect 4823 1250 5037 1254
rect 4838 1248 5037 1250
rect 5072 1250 5085 1260
rect 5103 1250 5120 1263
rect 5072 1248 5120 1250
rect 4714 1244 4747 1248
rect 4710 1242 4747 1244
rect 4710 1241 4777 1242
rect 4710 1236 4741 1241
rect 4747 1236 4777 1241
rect 4710 1232 4777 1236
rect 4683 1229 4777 1232
rect 4683 1222 4732 1229
rect 4683 1216 4713 1222
rect 4732 1217 4737 1222
rect 4649 1200 4729 1216
rect 4741 1208 4777 1229
rect 4838 1224 5027 1248
rect 5072 1247 5119 1248
rect 5085 1242 5119 1247
rect 4853 1221 5027 1224
rect 4846 1218 5027 1221
rect 5055 1241 5119 1242
rect 4649 1198 4668 1200
rect 4683 1198 4717 1200
rect 4649 1182 4729 1198
rect 4649 1176 4668 1182
rect 4365 1150 4468 1160
rect 4319 1148 4468 1150
rect 4489 1148 4524 1160
rect 4158 1146 4320 1148
rect 4170 1126 4189 1146
rect 4204 1144 4234 1146
rect 4053 1118 4094 1126
rect 4176 1122 4189 1126
rect 4241 1130 4320 1146
rect 4352 1146 4524 1148
rect 4352 1130 4431 1146
rect 4438 1144 4468 1146
rect 4016 1108 4045 1118
rect 4059 1108 4088 1118
rect 4103 1108 4133 1122
rect 4176 1108 4219 1122
rect 4241 1118 4431 1130
rect 4496 1126 4502 1146
rect 4226 1108 4256 1118
rect 4257 1108 4415 1118
rect 4419 1108 4449 1118
rect 4453 1108 4483 1122
rect 4511 1108 4524 1146
rect 4596 1160 4625 1176
rect 4639 1160 4668 1176
rect 4683 1166 4713 1182
rect 4741 1160 4747 1208
rect 4750 1202 4769 1208
rect 4784 1202 4814 1210
rect 4750 1194 4814 1202
rect 4750 1178 4830 1194
rect 4846 1187 4908 1218
rect 4924 1187 4986 1218
rect 5055 1216 5104 1241
rect 5119 1216 5149 1232
rect 5018 1202 5048 1210
rect 5055 1208 5165 1216
rect 5018 1194 5063 1202
rect 4750 1176 4769 1178
rect 4784 1176 4830 1178
rect 4750 1160 4830 1176
rect 4857 1174 4892 1187
rect 4933 1184 4970 1187
rect 4933 1182 4975 1184
rect 4862 1171 4892 1174
rect 4871 1167 4878 1171
rect 4878 1166 4879 1167
rect 4837 1160 4847 1166
rect 4596 1152 4631 1160
rect 4596 1126 4597 1152
rect 4604 1126 4631 1152
rect 4539 1108 4569 1122
rect 4596 1118 4631 1126
rect 4633 1152 4674 1160
rect 4633 1126 4648 1152
rect 4655 1126 4674 1152
rect 4738 1148 4769 1160
rect 4784 1148 4887 1160
rect 4899 1150 4925 1176
rect 4940 1171 4970 1182
rect 5002 1178 5064 1194
rect 5002 1176 5048 1178
rect 5002 1160 5064 1176
rect 5076 1160 5082 1208
rect 5085 1200 5165 1208
rect 5085 1198 5104 1200
rect 5119 1198 5153 1200
rect 5085 1182 5165 1198
rect 5085 1160 5104 1182
rect 5119 1166 5149 1182
rect 5177 1176 5183 1250
rect 5186 1176 5205 1320
rect 5220 1176 5226 1320
rect 5235 1250 5248 1320
rect 5300 1316 5322 1320
rect 5293 1294 5322 1308
rect 5375 1294 5391 1308
rect 5429 1304 5435 1306
rect 5442 1304 5550 1320
rect 5557 1304 5563 1306
rect 5571 1304 5586 1320
rect 5652 1314 5671 1317
rect 5293 1292 5391 1294
rect 5418 1292 5586 1304
rect 5601 1294 5617 1308
rect 5652 1295 5674 1314
rect 5684 1308 5700 1309
rect 5683 1306 5700 1308
rect 5684 1301 5700 1306
rect 5674 1294 5680 1295
rect 5683 1294 5712 1301
rect 5601 1293 5712 1294
rect 5601 1292 5718 1293
rect 5277 1284 5328 1292
rect 5375 1284 5409 1292
rect 5277 1272 5302 1284
rect 5309 1272 5328 1284
rect 5382 1282 5409 1284
rect 5418 1282 5639 1292
rect 5674 1289 5680 1292
rect 5382 1278 5639 1282
rect 5277 1264 5328 1272
rect 5375 1264 5639 1278
rect 5683 1284 5718 1292
rect 5229 1216 5248 1250
rect 5293 1256 5322 1264
rect 5293 1250 5310 1256
rect 5293 1248 5327 1250
rect 5375 1248 5391 1264
rect 5392 1254 5600 1264
rect 5601 1254 5617 1264
rect 5665 1260 5680 1275
rect 5683 1272 5684 1284
rect 5691 1272 5718 1284
rect 5683 1264 5718 1272
rect 5683 1263 5712 1264
rect 5403 1250 5617 1254
rect 5418 1248 5617 1250
rect 5652 1250 5665 1260
rect 5683 1250 5700 1263
rect 5652 1248 5700 1250
rect 5294 1244 5327 1248
rect 5290 1242 5327 1244
rect 5290 1241 5357 1242
rect 5290 1236 5321 1241
rect 5327 1236 5357 1241
rect 5290 1232 5357 1236
rect 5263 1229 5357 1232
rect 5263 1222 5312 1229
rect 5263 1216 5293 1222
rect 5312 1217 5317 1222
rect 5229 1200 5309 1216
rect 5321 1208 5357 1229
rect 5418 1224 5607 1248
rect 5652 1247 5699 1248
rect 5665 1242 5699 1247
rect 5433 1221 5607 1224
rect 5426 1218 5607 1221
rect 5635 1241 5699 1242
rect 5229 1198 5248 1200
rect 5263 1198 5297 1200
rect 5229 1182 5309 1198
rect 5229 1176 5248 1182
rect 4945 1150 5048 1160
rect 4899 1148 5048 1150
rect 5069 1148 5104 1160
rect 4738 1146 4900 1148
rect 4750 1126 4769 1146
rect 4784 1144 4814 1146
rect 4633 1118 4674 1126
rect 4756 1122 4769 1126
rect 4821 1130 4900 1146
rect 4932 1146 5104 1148
rect 4932 1130 5011 1146
rect 5018 1144 5048 1146
rect 4596 1108 4625 1118
rect 4639 1108 4668 1118
rect 4683 1108 4713 1122
rect 4756 1108 4799 1122
rect 4821 1118 5011 1130
rect 5076 1126 5082 1146
rect 4806 1108 4836 1118
rect 4837 1108 4995 1118
rect 4999 1108 5029 1118
rect 5033 1108 5063 1122
rect 5091 1108 5104 1146
rect 5176 1160 5205 1176
rect 5219 1160 5248 1176
rect 5263 1166 5293 1182
rect 5321 1160 5327 1208
rect 5330 1202 5349 1208
rect 5364 1202 5394 1210
rect 5330 1194 5394 1202
rect 5330 1178 5410 1194
rect 5426 1187 5488 1218
rect 5504 1187 5566 1218
rect 5635 1216 5684 1241
rect 5699 1216 5729 1232
rect 5598 1202 5628 1210
rect 5635 1208 5745 1216
rect 5598 1194 5643 1202
rect 5330 1176 5349 1178
rect 5364 1176 5410 1178
rect 5330 1160 5410 1176
rect 5437 1174 5472 1187
rect 5513 1184 5550 1187
rect 5513 1182 5555 1184
rect 5442 1171 5472 1174
rect 5451 1167 5458 1171
rect 5458 1166 5459 1167
rect 5417 1160 5427 1166
rect 5176 1152 5211 1160
rect 5176 1126 5177 1152
rect 5184 1126 5211 1152
rect 5119 1108 5149 1122
rect 5176 1118 5211 1126
rect 5213 1152 5254 1160
rect 5213 1126 5228 1152
rect 5235 1126 5254 1152
rect 5318 1148 5349 1160
rect 5364 1148 5467 1160
rect 5479 1150 5505 1176
rect 5520 1171 5550 1182
rect 5582 1178 5644 1194
rect 5582 1176 5628 1178
rect 5582 1160 5644 1176
rect 5656 1160 5662 1208
rect 5665 1200 5745 1208
rect 5665 1198 5684 1200
rect 5699 1198 5733 1200
rect 5665 1182 5745 1198
rect 5665 1160 5684 1182
rect 5699 1166 5729 1182
rect 5757 1176 5763 1250
rect 5766 1176 5785 1320
rect 5800 1176 5806 1320
rect 5815 1250 5828 1320
rect 5880 1316 5902 1320
rect 5873 1294 5902 1308
rect 5955 1294 5971 1308
rect 6009 1304 6015 1306
rect 6022 1304 6130 1320
rect 6137 1304 6143 1306
rect 6151 1304 6166 1320
rect 6232 1314 6251 1317
rect 5873 1292 5971 1294
rect 5998 1292 6166 1304
rect 6181 1294 6197 1308
rect 6232 1295 6254 1314
rect 6264 1308 6280 1309
rect 6263 1306 6280 1308
rect 6264 1301 6280 1306
rect 6254 1294 6260 1295
rect 6263 1294 6292 1301
rect 6181 1293 6292 1294
rect 6181 1292 6298 1293
rect 5857 1284 5908 1292
rect 5955 1284 5989 1292
rect 5857 1272 5882 1284
rect 5889 1272 5908 1284
rect 5962 1282 5989 1284
rect 5998 1282 6219 1292
rect 6254 1289 6260 1292
rect 5962 1278 6219 1282
rect 5857 1264 5908 1272
rect 5955 1264 6219 1278
rect 6263 1284 6298 1292
rect 5809 1216 5828 1250
rect 5873 1256 5902 1264
rect 5873 1250 5890 1256
rect 5873 1248 5907 1250
rect 5955 1248 5971 1264
rect 5972 1254 6180 1264
rect 6181 1254 6197 1264
rect 6245 1260 6260 1275
rect 6263 1272 6264 1284
rect 6271 1272 6298 1284
rect 6263 1264 6298 1272
rect 6263 1263 6292 1264
rect 5983 1250 6197 1254
rect 5998 1248 6197 1250
rect 6232 1250 6245 1260
rect 6263 1250 6280 1263
rect 6232 1248 6280 1250
rect 5874 1244 5907 1248
rect 5870 1242 5907 1244
rect 5870 1241 5937 1242
rect 5870 1236 5901 1241
rect 5907 1236 5937 1241
rect 5870 1232 5937 1236
rect 5843 1229 5937 1232
rect 5843 1222 5892 1229
rect 5843 1216 5873 1222
rect 5892 1217 5897 1222
rect 5809 1200 5889 1216
rect 5901 1208 5937 1229
rect 5998 1224 6187 1248
rect 6232 1247 6279 1248
rect 6245 1242 6279 1247
rect 6013 1221 6187 1224
rect 6006 1218 6187 1221
rect 6215 1241 6279 1242
rect 5809 1198 5828 1200
rect 5843 1198 5877 1200
rect 5809 1182 5889 1198
rect 5809 1176 5828 1182
rect 5525 1150 5628 1160
rect 5479 1148 5628 1150
rect 5649 1148 5684 1160
rect 5318 1146 5480 1148
rect 5330 1126 5349 1146
rect 5364 1144 5394 1146
rect 5213 1118 5254 1126
rect 5336 1122 5349 1126
rect 5401 1130 5480 1146
rect 5512 1146 5684 1148
rect 5512 1130 5591 1146
rect 5598 1144 5628 1146
rect 5176 1108 5205 1118
rect 5219 1108 5248 1118
rect 5263 1108 5293 1122
rect 5336 1108 5379 1122
rect 5401 1118 5591 1130
rect 5656 1126 5662 1146
rect 5386 1108 5416 1118
rect 5417 1108 5575 1118
rect 5579 1108 5609 1118
rect 5613 1108 5643 1122
rect 5671 1108 5684 1146
rect 5756 1160 5785 1176
rect 5799 1160 5828 1176
rect 5843 1166 5873 1182
rect 5901 1160 5907 1208
rect 5910 1202 5929 1208
rect 5944 1202 5974 1210
rect 5910 1194 5974 1202
rect 5910 1178 5990 1194
rect 6006 1187 6068 1218
rect 6084 1187 6146 1218
rect 6215 1216 6264 1241
rect 6279 1216 6309 1232
rect 6178 1202 6208 1210
rect 6215 1208 6325 1216
rect 6178 1194 6223 1202
rect 5910 1176 5929 1178
rect 5944 1176 5990 1178
rect 5910 1160 5990 1176
rect 6017 1174 6052 1187
rect 6093 1184 6130 1187
rect 6093 1182 6135 1184
rect 6022 1171 6052 1174
rect 6031 1167 6038 1171
rect 6038 1166 6039 1167
rect 5997 1160 6007 1166
rect 5756 1152 5791 1160
rect 5756 1126 5757 1152
rect 5764 1126 5791 1152
rect 5699 1108 5729 1122
rect 5756 1118 5791 1126
rect 5793 1152 5834 1160
rect 5793 1126 5808 1152
rect 5815 1126 5834 1152
rect 5898 1148 5929 1160
rect 5944 1148 6047 1160
rect 6059 1150 6085 1176
rect 6100 1171 6130 1182
rect 6162 1178 6224 1194
rect 6162 1176 6208 1178
rect 6162 1160 6224 1176
rect 6236 1160 6242 1208
rect 6245 1200 6325 1208
rect 6245 1198 6264 1200
rect 6279 1198 6313 1200
rect 6245 1182 6325 1198
rect 6245 1160 6264 1182
rect 6279 1166 6309 1182
rect 6337 1176 6343 1250
rect 6346 1176 6365 1320
rect 6380 1176 6386 1320
rect 6395 1250 6408 1320
rect 6460 1316 6482 1320
rect 6453 1294 6482 1308
rect 6535 1294 6551 1308
rect 6589 1304 6595 1306
rect 6602 1304 6710 1320
rect 6717 1304 6723 1306
rect 6731 1304 6746 1320
rect 6812 1314 6831 1317
rect 6453 1292 6551 1294
rect 6578 1292 6746 1304
rect 6761 1294 6777 1308
rect 6812 1295 6834 1314
rect 6844 1308 6860 1309
rect 6843 1306 6860 1308
rect 6844 1301 6860 1306
rect 6834 1294 6840 1295
rect 6843 1294 6872 1301
rect 6761 1293 6872 1294
rect 6761 1292 6878 1293
rect 6437 1284 6488 1292
rect 6535 1284 6569 1292
rect 6437 1272 6462 1284
rect 6469 1272 6488 1284
rect 6542 1282 6569 1284
rect 6578 1282 6799 1292
rect 6834 1289 6840 1292
rect 6542 1278 6799 1282
rect 6437 1264 6488 1272
rect 6535 1264 6799 1278
rect 6843 1284 6878 1292
rect 6389 1216 6408 1250
rect 6453 1256 6482 1264
rect 6453 1250 6470 1256
rect 6453 1248 6487 1250
rect 6535 1248 6551 1264
rect 6552 1254 6760 1264
rect 6761 1254 6777 1264
rect 6825 1260 6840 1275
rect 6843 1272 6844 1284
rect 6851 1272 6878 1284
rect 6843 1264 6878 1272
rect 6843 1263 6872 1264
rect 6563 1250 6777 1254
rect 6578 1248 6777 1250
rect 6812 1250 6825 1260
rect 6843 1250 6860 1263
rect 6812 1248 6860 1250
rect 6454 1244 6487 1248
rect 6450 1242 6487 1244
rect 6450 1241 6517 1242
rect 6450 1236 6481 1241
rect 6487 1236 6517 1241
rect 6450 1232 6517 1236
rect 6423 1229 6517 1232
rect 6423 1222 6472 1229
rect 6423 1216 6453 1222
rect 6472 1217 6477 1222
rect 6389 1200 6469 1216
rect 6481 1208 6517 1229
rect 6578 1224 6767 1248
rect 6812 1247 6859 1248
rect 6825 1242 6859 1247
rect 6593 1221 6767 1224
rect 6586 1218 6767 1221
rect 6795 1241 6859 1242
rect 6389 1198 6408 1200
rect 6423 1198 6457 1200
rect 6389 1182 6469 1198
rect 6389 1176 6408 1182
rect 6105 1150 6208 1160
rect 6059 1148 6208 1150
rect 6229 1148 6264 1160
rect 5898 1146 6060 1148
rect 5910 1126 5929 1146
rect 5944 1144 5974 1146
rect 5793 1118 5834 1126
rect 5916 1122 5929 1126
rect 5981 1130 6060 1146
rect 6092 1146 6264 1148
rect 6092 1130 6171 1146
rect 6178 1144 6208 1146
rect 5756 1108 5785 1118
rect 5799 1108 5828 1118
rect 5843 1108 5873 1122
rect 5916 1108 5959 1122
rect 5981 1118 6171 1130
rect 6236 1126 6242 1146
rect 5966 1108 5996 1118
rect 5997 1108 6155 1118
rect 6159 1108 6189 1118
rect 6193 1108 6223 1122
rect 6251 1108 6264 1146
rect 6336 1160 6365 1176
rect 6379 1160 6408 1176
rect 6423 1166 6453 1182
rect 6481 1160 6487 1208
rect 6490 1202 6509 1208
rect 6524 1202 6554 1210
rect 6490 1194 6554 1202
rect 6490 1178 6570 1194
rect 6586 1187 6648 1218
rect 6664 1187 6726 1218
rect 6795 1216 6844 1241
rect 6859 1216 6889 1232
rect 6758 1202 6788 1210
rect 6795 1208 6905 1216
rect 6758 1194 6803 1202
rect 6490 1176 6509 1178
rect 6524 1176 6570 1178
rect 6490 1160 6570 1176
rect 6597 1174 6632 1187
rect 6673 1184 6710 1187
rect 6673 1182 6715 1184
rect 6602 1171 6632 1174
rect 6611 1167 6618 1171
rect 6618 1166 6619 1167
rect 6577 1160 6587 1166
rect 6336 1152 6371 1160
rect 6336 1126 6337 1152
rect 6344 1126 6371 1152
rect 6279 1108 6309 1122
rect 6336 1118 6371 1126
rect 6373 1152 6414 1160
rect 6373 1126 6388 1152
rect 6395 1126 6414 1152
rect 6478 1148 6509 1160
rect 6524 1148 6627 1160
rect 6639 1150 6665 1176
rect 6680 1171 6710 1182
rect 6742 1178 6804 1194
rect 6742 1176 6788 1178
rect 6742 1160 6804 1176
rect 6816 1160 6822 1208
rect 6825 1200 6905 1208
rect 6825 1198 6844 1200
rect 6859 1198 6893 1200
rect 6825 1182 6905 1198
rect 6825 1160 6844 1182
rect 6859 1166 6889 1182
rect 6917 1176 6923 1250
rect 6926 1176 6945 1320
rect 6960 1176 6966 1320
rect 6975 1250 6988 1320
rect 7040 1316 7062 1320
rect 7033 1294 7062 1308
rect 7115 1294 7131 1308
rect 7169 1304 7175 1306
rect 7182 1304 7290 1320
rect 7297 1304 7303 1306
rect 7311 1304 7326 1320
rect 7392 1314 7411 1317
rect 7033 1292 7131 1294
rect 7158 1292 7326 1304
rect 7341 1294 7357 1308
rect 7392 1295 7414 1314
rect 7424 1308 7440 1309
rect 7423 1306 7440 1308
rect 7424 1301 7440 1306
rect 7414 1294 7420 1295
rect 7423 1294 7452 1301
rect 7341 1293 7452 1294
rect 7341 1292 7458 1293
rect 7017 1284 7068 1292
rect 7115 1284 7149 1292
rect 7017 1272 7042 1284
rect 7049 1272 7068 1284
rect 7122 1282 7149 1284
rect 7158 1282 7379 1292
rect 7414 1289 7420 1292
rect 7122 1278 7379 1282
rect 7017 1264 7068 1272
rect 7115 1264 7379 1278
rect 7423 1284 7458 1292
rect 6969 1216 6988 1250
rect 7033 1256 7062 1264
rect 7033 1250 7050 1256
rect 7033 1248 7067 1250
rect 7115 1248 7131 1264
rect 7132 1254 7340 1264
rect 7341 1254 7357 1264
rect 7405 1260 7420 1275
rect 7423 1272 7424 1284
rect 7431 1272 7458 1284
rect 7423 1264 7458 1272
rect 7423 1263 7452 1264
rect 7143 1250 7357 1254
rect 7158 1248 7357 1250
rect 7392 1250 7405 1260
rect 7423 1250 7440 1263
rect 7392 1248 7440 1250
rect 7034 1244 7067 1248
rect 7030 1242 7067 1244
rect 7030 1241 7097 1242
rect 7030 1236 7061 1241
rect 7067 1236 7097 1241
rect 7030 1232 7097 1236
rect 7003 1229 7097 1232
rect 7003 1222 7052 1229
rect 7003 1216 7033 1222
rect 7052 1217 7057 1222
rect 6969 1200 7049 1216
rect 7061 1208 7097 1229
rect 7158 1224 7347 1248
rect 7392 1247 7439 1248
rect 7405 1242 7439 1247
rect 7173 1221 7347 1224
rect 7166 1218 7347 1221
rect 7375 1241 7439 1242
rect 6969 1198 6988 1200
rect 7003 1198 7037 1200
rect 6969 1182 7049 1198
rect 6969 1176 6988 1182
rect 6685 1150 6788 1160
rect 6639 1148 6788 1150
rect 6809 1148 6844 1160
rect 6478 1146 6640 1148
rect 6490 1126 6509 1146
rect 6524 1144 6554 1146
rect 6373 1118 6414 1126
rect 6496 1122 6509 1126
rect 6561 1130 6640 1146
rect 6672 1146 6844 1148
rect 6672 1130 6751 1146
rect 6758 1144 6788 1146
rect 6336 1108 6365 1118
rect 6379 1108 6408 1118
rect 6423 1108 6453 1122
rect 6496 1108 6539 1122
rect 6561 1118 6751 1130
rect 6816 1126 6822 1146
rect 6546 1108 6576 1118
rect 6577 1108 6735 1118
rect 6739 1108 6769 1118
rect 6773 1108 6803 1122
rect 6831 1108 6844 1146
rect 6916 1160 6945 1176
rect 6959 1160 6988 1176
rect 7003 1166 7033 1182
rect 7061 1160 7067 1208
rect 7070 1202 7089 1208
rect 7104 1202 7134 1210
rect 7070 1194 7134 1202
rect 7070 1178 7150 1194
rect 7166 1187 7228 1218
rect 7244 1187 7306 1218
rect 7375 1216 7424 1241
rect 7439 1216 7469 1232
rect 7338 1202 7368 1210
rect 7375 1208 7485 1216
rect 7338 1194 7383 1202
rect 7070 1176 7089 1178
rect 7104 1176 7150 1178
rect 7070 1160 7150 1176
rect 7177 1174 7212 1187
rect 7253 1184 7290 1187
rect 7253 1182 7295 1184
rect 7182 1171 7212 1174
rect 7191 1167 7198 1171
rect 7198 1166 7199 1167
rect 7157 1160 7167 1166
rect 6916 1152 6951 1160
rect 6916 1126 6917 1152
rect 6924 1126 6951 1152
rect 6859 1108 6889 1122
rect 6916 1118 6951 1126
rect 6953 1152 6994 1160
rect 6953 1126 6968 1152
rect 6975 1126 6994 1152
rect 7058 1148 7089 1160
rect 7104 1148 7207 1160
rect 7219 1150 7245 1176
rect 7260 1171 7290 1182
rect 7322 1178 7384 1194
rect 7322 1176 7368 1178
rect 7322 1160 7384 1176
rect 7396 1160 7402 1208
rect 7405 1200 7485 1208
rect 7405 1198 7424 1200
rect 7439 1198 7473 1200
rect 7405 1182 7485 1198
rect 7405 1160 7424 1182
rect 7439 1166 7469 1182
rect 7497 1176 7503 1250
rect 7506 1176 7525 1320
rect 7540 1176 7546 1320
rect 7555 1250 7568 1320
rect 7620 1316 7642 1320
rect 7613 1294 7642 1308
rect 7695 1294 7711 1308
rect 7749 1304 7755 1306
rect 7762 1304 7870 1320
rect 7877 1304 7883 1306
rect 7891 1304 7906 1320
rect 7972 1314 7991 1317
rect 7613 1292 7711 1294
rect 7738 1292 7906 1304
rect 7921 1294 7937 1308
rect 7972 1295 7994 1314
rect 8004 1308 8020 1309
rect 8003 1306 8020 1308
rect 8004 1301 8020 1306
rect 7994 1294 8000 1295
rect 8003 1294 8032 1301
rect 7921 1293 8032 1294
rect 7921 1292 8038 1293
rect 7597 1284 7648 1292
rect 7695 1284 7729 1292
rect 7597 1272 7622 1284
rect 7629 1272 7648 1284
rect 7702 1282 7729 1284
rect 7738 1282 7959 1292
rect 7994 1289 8000 1292
rect 7702 1278 7959 1282
rect 7597 1264 7648 1272
rect 7695 1264 7959 1278
rect 8003 1284 8038 1292
rect 7549 1216 7568 1250
rect 7613 1256 7642 1264
rect 7613 1250 7630 1256
rect 7613 1248 7647 1250
rect 7695 1248 7711 1264
rect 7712 1254 7920 1264
rect 7921 1254 7937 1264
rect 7985 1260 8000 1275
rect 8003 1272 8004 1284
rect 8011 1272 8038 1284
rect 8003 1264 8038 1272
rect 8003 1263 8032 1264
rect 7723 1250 7937 1254
rect 7738 1248 7937 1250
rect 7972 1250 7985 1260
rect 8003 1250 8020 1263
rect 7972 1248 8020 1250
rect 7614 1244 7647 1248
rect 7610 1242 7647 1244
rect 7610 1241 7677 1242
rect 7610 1236 7641 1241
rect 7647 1236 7677 1241
rect 7610 1232 7677 1236
rect 7583 1229 7677 1232
rect 7583 1222 7632 1229
rect 7583 1216 7613 1222
rect 7632 1217 7637 1222
rect 7549 1200 7629 1216
rect 7641 1208 7677 1229
rect 7738 1224 7927 1248
rect 7972 1247 8019 1248
rect 7985 1242 8019 1247
rect 7753 1221 7927 1224
rect 7746 1218 7927 1221
rect 7955 1241 8019 1242
rect 7549 1198 7568 1200
rect 7583 1198 7617 1200
rect 7549 1182 7629 1198
rect 7549 1176 7568 1182
rect 7265 1150 7368 1160
rect 7219 1148 7368 1150
rect 7389 1148 7424 1160
rect 7058 1146 7220 1148
rect 7070 1126 7089 1146
rect 7104 1144 7134 1146
rect 6953 1118 6994 1126
rect 7076 1122 7089 1126
rect 7141 1130 7220 1146
rect 7252 1146 7424 1148
rect 7252 1130 7331 1146
rect 7338 1144 7368 1146
rect 6916 1108 6945 1118
rect 6959 1108 6988 1118
rect 7003 1108 7033 1122
rect 7076 1108 7119 1122
rect 7141 1118 7331 1130
rect 7396 1126 7402 1146
rect 7126 1108 7156 1118
rect 7157 1108 7315 1118
rect 7319 1108 7349 1118
rect 7353 1108 7383 1122
rect 7411 1108 7424 1146
rect 7496 1160 7525 1176
rect 7539 1160 7568 1176
rect 7583 1166 7613 1182
rect 7641 1160 7647 1208
rect 7650 1202 7669 1208
rect 7684 1202 7714 1210
rect 7650 1194 7714 1202
rect 7650 1178 7730 1194
rect 7746 1187 7808 1218
rect 7824 1187 7886 1218
rect 7955 1216 8004 1241
rect 8019 1216 8049 1232
rect 7918 1202 7948 1210
rect 7955 1208 8065 1216
rect 7918 1194 7963 1202
rect 7650 1176 7669 1178
rect 7684 1176 7730 1178
rect 7650 1160 7730 1176
rect 7757 1174 7792 1187
rect 7833 1184 7870 1187
rect 7833 1182 7875 1184
rect 7762 1171 7792 1174
rect 7771 1167 7778 1171
rect 7778 1166 7779 1167
rect 7737 1160 7747 1166
rect 7496 1152 7531 1160
rect 7496 1126 7497 1152
rect 7504 1126 7531 1152
rect 7439 1108 7469 1122
rect 7496 1118 7531 1126
rect 7533 1152 7574 1160
rect 7533 1126 7548 1152
rect 7555 1126 7574 1152
rect 7638 1148 7669 1160
rect 7684 1148 7787 1160
rect 7799 1150 7825 1176
rect 7840 1171 7870 1182
rect 7902 1178 7964 1194
rect 7902 1176 7948 1178
rect 7902 1160 7964 1176
rect 7976 1160 7982 1208
rect 7985 1200 8065 1208
rect 7985 1198 8004 1200
rect 8019 1198 8053 1200
rect 7985 1182 8065 1198
rect 7985 1160 8004 1182
rect 8019 1166 8049 1182
rect 8077 1176 8083 1250
rect 8086 1176 8105 1320
rect 8120 1176 8126 1320
rect 8135 1250 8148 1320
rect 8200 1316 8222 1320
rect 8193 1294 8222 1308
rect 8275 1294 8291 1308
rect 8329 1304 8335 1306
rect 8342 1304 8450 1320
rect 8457 1304 8463 1306
rect 8471 1304 8486 1320
rect 8552 1314 8571 1317
rect 8193 1292 8291 1294
rect 8318 1292 8486 1304
rect 8501 1294 8517 1308
rect 8552 1295 8574 1314
rect 8584 1308 8600 1309
rect 8583 1306 8600 1308
rect 8584 1301 8600 1306
rect 8574 1294 8580 1295
rect 8583 1294 8612 1301
rect 8501 1293 8612 1294
rect 8501 1292 8618 1293
rect 8177 1284 8228 1292
rect 8275 1284 8309 1292
rect 8177 1272 8202 1284
rect 8209 1272 8228 1284
rect 8282 1282 8309 1284
rect 8318 1282 8539 1292
rect 8574 1289 8580 1292
rect 8282 1278 8539 1282
rect 8177 1264 8228 1272
rect 8275 1264 8539 1278
rect 8583 1284 8618 1292
rect 8129 1216 8148 1250
rect 8193 1256 8222 1264
rect 8193 1250 8210 1256
rect 8193 1248 8227 1250
rect 8275 1248 8291 1264
rect 8292 1254 8500 1264
rect 8501 1254 8517 1264
rect 8565 1260 8580 1275
rect 8583 1272 8584 1284
rect 8591 1272 8618 1284
rect 8583 1264 8618 1272
rect 8583 1263 8612 1264
rect 8303 1250 8517 1254
rect 8318 1248 8517 1250
rect 8552 1250 8565 1260
rect 8583 1250 8600 1263
rect 8552 1248 8600 1250
rect 8194 1244 8227 1248
rect 8190 1242 8227 1244
rect 8190 1241 8257 1242
rect 8190 1236 8221 1241
rect 8227 1236 8257 1241
rect 8190 1232 8257 1236
rect 8163 1229 8257 1232
rect 8163 1222 8212 1229
rect 8163 1216 8193 1222
rect 8212 1217 8217 1222
rect 8129 1200 8209 1216
rect 8221 1208 8257 1229
rect 8318 1224 8507 1248
rect 8552 1247 8599 1248
rect 8565 1242 8599 1247
rect 8333 1221 8507 1224
rect 8326 1218 8507 1221
rect 8535 1241 8599 1242
rect 8129 1198 8148 1200
rect 8163 1198 8197 1200
rect 8129 1182 8209 1198
rect 8129 1176 8148 1182
rect 7845 1150 7948 1160
rect 7799 1148 7948 1150
rect 7969 1148 8004 1160
rect 7638 1146 7800 1148
rect 7650 1126 7669 1146
rect 7684 1144 7714 1146
rect 7533 1118 7574 1126
rect 7656 1122 7669 1126
rect 7721 1130 7800 1146
rect 7832 1146 8004 1148
rect 7832 1130 7911 1146
rect 7918 1144 7948 1146
rect 7496 1108 7525 1118
rect 7539 1108 7568 1118
rect 7583 1108 7613 1122
rect 7656 1108 7699 1122
rect 7721 1118 7911 1130
rect 7976 1126 7982 1146
rect 7706 1108 7736 1118
rect 7737 1108 7895 1118
rect 7899 1108 7929 1118
rect 7933 1108 7963 1122
rect 7991 1108 8004 1146
rect 8076 1160 8105 1176
rect 8119 1160 8148 1176
rect 8163 1166 8193 1182
rect 8221 1160 8227 1208
rect 8230 1202 8249 1208
rect 8264 1202 8294 1210
rect 8230 1194 8294 1202
rect 8230 1178 8310 1194
rect 8326 1187 8388 1218
rect 8404 1187 8466 1218
rect 8535 1216 8584 1241
rect 8599 1216 8629 1232
rect 8498 1202 8528 1210
rect 8535 1208 8645 1216
rect 8498 1194 8543 1202
rect 8230 1176 8249 1178
rect 8264 1176 8310 1178
rect 8230 1160 8310 1176
rect 8337 1174 8372 1187
rect 8413 1184 8450 1187
rect 8413 1182 8455 1184
rect 8342 1171 8372 1174
rect 8351 1167 8358 1171
rect 8358 1166 8359 1167
rect 8317 1160 8327 1166
rect 8076 1152 8111 1160
rect 8076 1126 8077 1152
rect 8084 1126 8111 1152
rect 8019 1108 8049 1122
rect 8076 1118 8111 1126
rect 8113 1152 8154 1160
rect 8113 1126 8128 1152
rect 8135 1126 8154 1152
rect 8218 1148 8249 1160
rect 8264 1148 8367 1160
rect 8379 1150 8405 1176
rect 8420 1171 8450 1182
rect 8482 1178 8544 1194
rect 8482 1176 8528 1178
rect 8482 1160 8544 1176
rect 8556 1160 8562 1208
rect 8565 1200 8645 1208
rect 8565 1198 8584 1200
rect 8599 1198 8633 1200
rect 8565 1182 8645 1198
rect 8565 1160 8584 1182
rect 8599 1166 8629 1182
rect 8657 1176 8663 1250
rect 8666 1176 8685 1320
rect 8700 1176 8706 1320
rect 8715 1250 8728 1320
rect 8780 1316 8802 1320
rect 8773 1294 8802 1308
rect 8855 1294 8871 1308
rect 8909 1304 8915 1306
rect 8922 1304 9030 1320
rect 9037 1304 9043 1306
rect 9051 1304 9066 1320
rect 9132 1314 9151 1317
rect 8773 1292 8871 1294
rect 8898 1292 9066 1304
rect 9081 1294 9097 1308
rect 9132 1295 9154 1314
rect 9164 1308 9180 1309
rect 9163 1306 9180 1308
rect 9164 1301 9180 1306
rect 9154 1294 9160 1295
rect 9163 1294 9192 1301
rect 9081 1293 9192 1294
rect 9081 1292 9198 1293
rect 8757 1284 8808 1292
rect 8855 1284 8889 1292
rect 8757 1272 8782 1284
rect 8789 1272 8808 1284
rect 8862 1282 8889 1284
rect 8898 1282 9119 1292
rect 9154 1289 9160 1292
rect 8862 1278 9119 1282
rect 8757 1264 8808 1272
rect 8855 1264 9119 1278
rect 9163 1284 9198 1292
rect 8709 1216 8728 1250
rect 8773 1256 8802 1264
rect 8773 1250 8790 1256
rect 8773 1248 8807 1250
rect 8855 1248 8871 1264
rect 8872 1254 9080 1264
rect 9081 1254 9097 1264
rect 9145 1260 9160 1275
rect 9163 1272 9164 1284
rect 9171 1272 9198 1284
rect 9163 1264 9198 1272
rect 9163 1263 9192 1264
rect 8883 1250 9097 1254
rect 8898 1248 9097 1250
rect 9132 1250 9145 1260
rect 9163 1250 9180 1263
rect 9132 1248 9180 1250
rect 8774 1244 8807 1248
rect 8770 1242 8807 1244
rect 8770 1241 8837 1242
rect 8770 1236 8801 1241
rect 8807 1236 8837 1241
rect 8770 1232 8837 1236
rect 8743 1229 8837 1232
rect 8743 1222 8792 1229
rect 8743 1216 8773 1222
rect 8792 1217 8797 1222
rect 8709 1200 8789 1216
rect 8801 1208 8837 1229
rect 8898 1224 9087 1248
rect 9132 1247 9179 1248
rect 9145 1242 9179 1247
rect 8913 1221 9087 1224
rect 8906 1218 9087 1221
rect 9115 1241 9179 1242
rect 8709 1198 8728 1200
rect 8743 1198 8777 1200
rect 8709 1182 8789 1198
rect 8709 1176 8728 1182
rect 8425 1150 8528 1160
rect 8379 1148 8528 1150
rect 8549 1148 8584 1160
rect 8218 1146 8380 1148
rect 8230 1126 8249 1146
rect 8264 1144 8294 1146
rect 8113 1118 8154 1126
rect 8236 1122 8249 1126
rect 8301 1130 8380 1146
rect 8412 1146 8584 1148
rect 8412 1130 8491 1146
rect 8498 1144 8528 1146
rect 8076 1108 8105 1118
rect 8119 1108 8148 1118
rect 8163 1108 8193 1122
rect 8236 1108 8279 1122
rect 8301 1118 8491 1130
rect 8556 1126 8562 1146
rect 8286 1108 8316 1118
rect 8317 1108 8475 1118
rect 8479 1108 8509 1118
rect 8513 1108 8543 1122
rect 8571 1108 8584 1146
rect 8656 1160 8685 1176
rect 8699 1160 8728 1176
rect 8743 1166 8773 1182
rect 8801 1160 8807 1208
rect 8810 1202 8829 1208
rect 8844 1202 8874 1210
rect 8810 1194 8874 1202
rect 8810 1178 8890 1194
rect 8906 1187 8968 1218
rect 8984 1187 9046 1218
rect 9115 1216 9164 1241
rect 9179 1216 9209 1232
rect 9078 1202 9108 1210
rect 9115 1208 9225 1216
rect 9078 1194 9123 1202
rect 8810 1176 8829 1178
rect 8844 1176 8890 1178
rect 8810 1160 8890 1176
rect 8917 1174 8952 1187
rect 8993 1184 9030 1187
rect 8993 1182 9035 1184
rect 8922 1171 8952 1174
rect 8931 1167 8938 1171
rect 8938 1166 8939 1167
rect 8897 1160 8907 1166
rect 8656 1152 8691 1160
rect 8656 1126 8657 1152
rect 8664 1126 8691 1152
rect 8599 1108 8629 1122
rect 8656 1118 8691 1126
rect 8693 1152 8734 1160
rect 8693 1126 8708 1152
rect 8715 1126 8734 1152
rect 8798 1148 8829 1160
rect 8844 1148 8947 1160
rect 8959 1150 8985 1176
rect 9000 1171 9030 1182
rect 9062 1178 9124 1194
rect 9062 1176 9108 1178
rect 9062 1160 9124 1176
rect 9136 1160 9142 1208
rect 9145 1200 9225 1208
rect 9145 1198 9164 1200
rect 9179 1198 9213 1200
rect 9145 1182 9225 1198
rect 9145 1160 9164 1182
rect 9179 1166 9209 1182
rect 9237 1176 9243 1250
rect 9252 1176 9265 1320
rect 9005 1150 9108 1160
rect 8959 1148 9108 1150
rect 9129 1148 9164 1160
rect 8798 1146 8960 1148
rect 8810 1126 8829 1146
rect 8844 1144 8874 1146
rect 8693 1118 8734 1126
rect 8816 1122 8829 1126
rect 8881 1130 8960 1146
rect 8992 1146 9164 1148
rect 8992 1130 9071 1146
rect 9078 1144 9108 1146
rect 8656 1108 8685 1118
rect 8699 1108 8728 1118
rect 8743 1108 8773 1122
rect 8816 1108 8859 1122
rect 8881 1118 9071 1130
rect 9136 1126 9142 1146
rect 8866 1108 8896 1118
rect 8897 1108 9055 1118
rect 9059 1108 9089 1118
rect 9093 1108 9123 1122
rect 9151 1108 9164 1146
rect 9236 1160 9265 1176
rect 9236 1152 9271 1160
rect 9236 1126 9237 1152
rect 9244 1126 9271 1152
rect 9179 1108 9209 1122
rect 9236 1118 9271 1126
rect 9236 1108 9265 1118
rect -1 1102 9265 1108
rect 0 1094 9265 1102
rect 15 1064 28 1094
rect 43 1080 73 1094
rect 116 1080 159 1094
rect 166 1080 386 1094
rect 393 1080 423 1094
rect 83 1066 98 1078
rect 117 1066 130 1080
rect 198 1076 351 1080
rect 80 1064 102 1066
rect 180 1064 372 1076
rect 451 1064 464 1094
rect 479 1080 509 1094
rect 546 1064 565 1094
rect 580 1064 586 1094
rect 595 1064 608 1094
rect 623 1080 653 1094
rect 696 1080 739 1094
rect 746 1080 966 1094
rect 973 1080 1003 1094
rect 663 1066 678 1078
rect 697 1066 710 1080
rect 778 1076 931 1080
rect 660 1064 682 1066
rect 760 1064 952 1076
rect 1031 1064 1044 1094
rect 1059 1080 1089 1094
rect 1126 1064 1145 1094
rect 1160 1064 1166 1094
rect 1175 1064 1188 1094
rect 1203 1080 1233 1094
rect 1276 1080 1319 1094
rect 1326 1080 1546 1094
rect 1553 1080 1583 1094
rect 1243 1066 1258 1078
rect 1277 1066 1290 1080
rect 1358 1076 1511 1080
rect 1240 1064 1262 1066
rect 1340 1064 1532 1076
rect 1611 1064 1624 1094
rect 1639 1080 1669 1094
rect 1706 1064 1725 1094
rect 1740 1064 1746 1094
rect 1755 1064 1768 1094
rect 1783 1080 1813 1094
rect 1856 1080 1899 1094
rect 1906 1080 2126 1094
rect 2133 1080 2163 1094
rect 1823 1066 1838 1078
rect 1857 1066 1870 1080
rect 1938 1076 2091 1080
rect 1820 1064 1842 1066
rect 1920 1064 2112 1076
rect 2191 1064 2204 1094
rect 2219 1080 2249 1094
rect 2286 1064 2305 1094
rect 2320 1064 2326 1094
rect 2335 1064 2348 1094
rect 2363 1080 2393 1094
rect 2436 1080 2479 1094
rect 2486 1080 2706 1094
rect 2713 1080 2743 1094
rect 2403 1066 2418 1078
rect 2437 1066 2450 1080
rect 2518 1076 2671 1080
rect 2400 1064 2422 1066
rect 2500 1064 2692 1076
rect 2771 1064 2784 1094
rect 2799 1080 2829 1094
rect 2866 1064 2885 1094
rect 2900 1064 2906 1094
rect 2915 1064 2928 1094
rect 2943 1080 2973 1094
rect 3016 1080 3059 1094
rect 3066 1080 3286 1094
rect 3293 1080 3323 1094
rect 2983 1066 2998 1078
rect 3017 1066 3030 1080
rect 3098 1076 3251 1080
rect 2980 1064 3002 1066
rect 3080 1064 3272 1076
rect 3351 1064 3364 1094
rect 3379 1080 3409 1094
rect 3446 1064 3465 1094
rect 3480 1064 3486 1094
rect 3495 1064 3508 1094
rect 3523 1080 3553 1094
rect 3596 1080 3639 1094
rect 3646 1080 3866 1094
rect 3873 1080 3903 1094
rect 3563 1066 3578 1078
rect 3597 1066 3610 1080
rect 3678 1076 3831 1080
rect 3560 1064 3582 1066
rect 3660 1064 3852 1076
rect 3931 1064 3944 1094
rect 3959 1080 3989 1094
rect 4026 1064 4045 1094
rect 4060 1064 4066 1094
rect 4075 1064 4088 1094
rect 4103 1080 4133 1094
rect 4176 1080 4219 1094
rect 4226 1080 4446 1094
rect 4453 1080 4483 1094
rect 4143 1066 4158 1078
rect 4177 1066 4190 1080
rect 4258 1076 4411 1080
rect 4140 1064 4162 1066
rect 4240 1064 4432 1076
rect 4511 1064 4524 1094
rect 4539 1080 4569 1094
rect 4606 1064 4625 1094
rect 4640 1064 4646 1094
rect 4655 1064 4668 1094
rect 4683 1080 4713 1094
rect 4756 1080 4799 1094
rect 4806 1080 5026 1094
rect 5033 1080 5063 1094
rect 4723 1066 4738 1078
rect 4757 1066 4770 1080
rect 4838 1076 4991 1080
rect 4720 1064 4742 1066
rect 4820 1064 5012 1076
rect 5091 1064 5104 1094
rect 5119 1080 5149 1094
rect 5186 1064 5205 1094
rect 5220 1064 5226 1094
rect 5235 1064 5248 1094
rect 5263 1080 5293 1094
rect 5336 1080 5379 1094
rect 5386 1080 5606 1094
rect 5613 1080 5643 1094
rect 5303 1066 5318 1078
rect 5337 1066 5350 1080
rect 5418 1076 5571 1080
rect 5300 1064 5322 1066
rect 5400 1064 5592 1076
rect 5671 1064 5684 1094
rect 5699 1080 5729 1094
rect 5766 1064 5785 1094
rect 5800 1064 5806 1094
rect 5815 1064 5828 1094
rect 5843 1080 5873 1094
rect 5916 1080 5959 1094
rect 5966 1080 6186 1094
rect 6193 1080 6223 1094
rect 5883 1066 5898 1078
rect 5917 1066 5930 1080
rect 5998 1076 6151 1080
rect 5880 1064 5902 1066
rect 5980 1064 6172 1076
rect 6251 1064 6264 1094
rect 6279 1080 6309 1094
rect 6346 1064 6365 1094
rect 6380 1064 6386 1094
rect 6395 1064 6408 1094
rect 6423 1080 6453 1094
rect 6496 1080 6539 1094
rect 6546 1080 6766 1094
rect 6773 1080 6803 1094
rect 6463 1066 6478 1078
rect 6497 1066 6510 1080
rect 6578 1076 6731 1080
rect 6460 1064 6482 1066
rect 6560 1064 6752 1076
rect 6831 1064 6844 1094
rect 6859 1080 6889 1094
rect 6926 1064 6945 1094
rect 6960 1064 6966 1094
rect 6975 1064 6988 1094
rect 7003 1080 7033 1094
rect 7076 1080 7119 1094
rect 7126 1080 7346 1094
rect 7353 1080 7383 1094
rect 7043 1066 7058 1078
rect 7077 1066 7090 1080
rect 7158 1076 7311 1080
rect 7040 1064 7062 1066
rect 7140 1064 7332 1076
rect 7411 1064 7424 1094
rect 7439 1080 7469 1094
rect 7506 1064 7525 1094
rect 7540 1064 7546 1094
rect 7555 1064 7568 1094
rect 7583 1080 7613 1094
rect 7656 1080 7699 1094
rect 7706 1080 7926 1094
rect 7933 1080 7963 1094
rect 7623 1066 7638 1078
rect 7657 1066 7670 1080
rect 7738 1076 7891 1080
rect 7620 1064 7642 1066
rect 7720 1064 7912 1076
rect 7991 1064 8004 1094
rect 8019 1080 8049 1094
rect 8086 1064 8105 1094
rect 8120 1064 8126 1094
rect 8135 1064 8148 1094
rect 8163 1080 8193 1094
rect 8236 1080 8279 1094
rect 8286 1080 8506 1094
rect 8513 1080 8543 1094
rect 8203 1066 8218 1078
rect 8237 1066 8250 1080
rect 8318 1076 8471 1080
rect 8200 1064 8222 1066
rect 8300 1064 8492 1076
rect 8571 1064 8584 1094
rect 8599 1080 8629 1094
rect 8666 1064 8685 1094
rect 8700 1064 8706 1094
rect 8715 1064 8728 1094
rect 8743 1080 8773 1094
rect 8816 1080 8859 1094
rect 8866 1080 9086 1094
rect 9093 1080 9123 1094
rect 8783 1066 8798 1078
rect 8817 1066 8830 1080
rect 8898 1076 9051 1080
rect 8780 1064 8802 1066
rect 8880 1064 9072 1076
rect 9151 1064 9164 1094
rect 9179 1080 9209 1094
rect 9252 1064 9265 1094
rect 0 1050 9265 1064
rect 15 980 28 1050
rect 80 1046 102 1050
rect 73 1024 102 1038
rect 155 1024 171 1038
rect 209 1034 215 1036
rect 222 1034 330 1050
rect 337 1034 343 1036
rect 351 1034 366 1050
rect 432 1044 451 1047
rect 73 1022 171 1024
rect 198 1022 366 1034
rect 381 1024 397 1038
rect 432 1025 454 1044
rect 464 1038 480 1039
rect 463 1036 480 1038
rect 464 1031 480 1036
rect 454 1024 460 1025
rect 463 1024 492 1031
rect 381 1023 492 1024
rect 381 1022 498 1023
rect 57 1014 108 1022
rect 155 1014 189 1022
rect 57 1002 82 1014
rect 89 1002 108 1014
rect 162 1012 189 1014
rect 198 1012 419 1022
rect 454 1019 460 1022
rect 162 1008 419 1012
rect 57 994 108 1002
rect 155 994 419 1008
rect 463 1014 498 1022
rect 9 946 28 980
rect 73 986 102 994
rect 73 980 90 986
rect 73 978 107 980
rect 155 978 171 994
rect 172 984 380 994
rect 381 984 397 994
rect 445 990 460 1005
rect 463 1002 464 1014
rect 471 1002 498 1014
rect 463 994 498 1002
rect 463 993 492 994
rect 183 980 397 984
rect 198 978 397 980
rect 432 980 445 990
rect 463 980 480 993
rect 432 978 480 980
rect 74 974 107 978
rect 70 972 107 974
rect 70 971 137 972
rect 70 966 101 971
rect 107 966 137 971
rect 70 962 137 966
rect 43 959 137 962
rect 43 952 92 959
rect 43 946 73 952
rect 92 947 97 952
rect 9 930 89 946
rect 101 938 137 959
rect 198 954 387 978
rect 432 977 479 978
rect 445 972 479 977
rect 213 951 387 954
rect 206 948 387 951
rect 415 971 479 972
rect 9 928 28 930
rect 43 928 77 930
rect 9 912 89 928
rect 9 906 28 912
rect -1 890 28 906
rect 43 896 73 912
rect 101 890 107 938
rect 110 932 129 938
rect 144 932 174 940
rect 110 924 174 932
rect 110 908 190 924
rect 206 917 268 948
rect 284 917 346 948
rect 415 946 464 971
rect 479 946 509 962
rect 378 932 408 940
rect 415 938 525 946
rect 378 924 423 932
rect 110 906 129 908
rect 144 906 190 908
rect 110 890 190 906
rect 217 904 252 917
rect 293 914 330 917
rect 293 912 335 914
rect 222 901 252 904
rect 231 897 238 901
rect 238 896 239 897
rect 197 890 207 896
rect -7 882 34 890
rect -7 856 8 882
rect 15 856 34 882
rect 98 878 129 890
rect 144 878 247 890
rect 259 880 285 906
rect 300 901 330 912
rect 362 908 424 924
rect 362 906 408 908
rect 362 890 424 906
rect 436 890 442 938
rect 445 930 525 938
rect 445 928 464 930
rect 479 928 513 930
rect 445 912 525 928
rect 445 890 464 912
rect 479 896 509 912
rect 537 906 543 980
rect 546 906 565 1050
rect 580 906 586 1050
rect 595 980 608 1050
rect 660 1046 682 1050
rect 653 1024 682 1038
rect 735 1024 751 1038
rect 789 1034 795 1036
rect 802 1034 910 1050
rect 917 1034 923 1036
rect 931 1034 946 1050
rect 1012 1044 1031 1047
rect 653 1022 751 1024
rect 778 1022 946 1034
rect 961 1024 977 1038
rect 1012 1025 1034 1044
rect 1044 1038 1060 1039
rect 1043 1036 1060 1038
rect 1044 1031 1060 1036
rect 1034 1024 1040 1025
rect 1043 1024 1072 1031
rect 961 1023 1072 1024
rect 961 1022 1078 1023
rect 637 1014 688 1022
rect 735 1014 769 1022
rect 637 1002 662 1014
rect 669 1002 688 1014
rect 742 1012 769 1014
rect 778 1012 999 1022
rect 1034 1019 1040 1022
rect 742 1008 999 1012
rect 637 994 688 1002
rect 735 994 999 1008
rect 1043 1014 1078 1022
rect 589 946 608 980
rect 653 986 682 994
rect 653 980 670 986
rect 653 978 687 980
rect 735 978 751 994
rect 752 984 960 994
rect 961 984 977 994
rect 1025 990 1040 1005
rect 1043 1002 1044 1014
rect 1051 1002 1078 1014
rect 1043 994 1078 1002
rect 1043 993 1072 994
rect 763 980 977 984
rect 778 978 977 980
rect 1012 980 1025 990
rect 1043 980 1060 993
rect 1012 978 1060 980
rect 654 974 687 978
rect 650 972 687 974
rect 650 971 717 972
rect 650 966 681 971
rect 687 966 717 971
rect 650 962 717 966
rect 623 959 717 962
rect 623 952 672 959
rect 623 946 653 952
rect 672 947 677 952
rect 589 930 669 946
rect 681 938 717 959
rect 778 954 967 978
rect 1012 977 1059 978
rect 1025 972 1059 977
rect 793 951 967 954
rect 786 948 967 951
rect 995 971 1059 972
rect 589 928 608 930
rect 623 928 657 930
rect 589 912 669 928
rect 589 906 608 912
rect 305 880 408 890
rect 259 878 408 880
rect 429 878 464 890
rect 98 876 260 878
rect 110 856 129 876
rect 144 874 174 876
rect -7 848 34 856
rect 116 852 129 856
rect 181 860 260 876
rect 292 876 464 878
rect 292 860 371 876
rect 378 874 408 876
rect -1 838 28 848
rect 43 838 73 852
rect 116 838 159 852
rect 181 848 371 860
rect 436 856 442 876
rect 166 838 196 848
rect 197 838 355 848
rect 359 838 389 848
rect 393 838 423 852
rect 451 838 464 876
rect 536 890 565 906
rect 579 890 608 906
rect 623 896 653 912
rect 681 890 687 938
rect 690 932 709 938
rect 724 932 754 940
rect 690 924 754 932
rect 690 908 770 924
rect 786 917 848 948
rect 864 917 926 948
rect 995 946 1044 971
rect 1059 946 1089 962
rect 958 932 988 940
rect 995 938 1105 946
rect 958 924 1003 932
rect 690 906 709 908
rect 724 906 770 908
rect 690 890 770 906
rect 797 904 832 917
rect 873 914 910 917
rect 873 912 915 914
rect 802 901 832 904
rect 811 897 818 901
rect 818 896 819 897
rect 777 890 787 896
rect 536 882 571 890
rect 536 856 537 882
rect 544 856 571 882
rect 479 838 509 852
rect 536 848 571 856
rect 573 882 614 890
rect 573 856 588 882
rect 595 856 614 882
rect 678 878 709 890
rect 724 878 827 890
rect 839 880 865 906
rect 880 901 910 912
rect 942 908 1004 924
rect 942 906 988 908
rect 942 890 1004 906
rect 1016 890 1022 938
rect 1025 930 1105 938
rect 1025 928 1044 930
rect 1059 928 1093 930
rect 1025 912 1105 928
rect 1025 890 1044 912
rect 1059 896 1089 912
rect 1117 906 1123 980
rect 1126 906 1145 1050
rect 1160 906 1166 1050
rect 1175 980 1188 1050
rect 1240 1046 1262 1050
rect 1233 1024 1262 1038
rect 1315 1024 1331 1038
rect 1369 1034 1375 1036
rect 1382 1034 1490 1050
rect 1497 1034 1503 1036
rect 1511 1034 1526 1050
rect 1592 1044 1611 1047
rect 1233 1022 1331 1024
rect 1358 1022 1526 1034
rect 1541 1024 1557 1038
rect 1592 1025 1614 1044
rect 1624 1038 1640 1039
rect 1623 1036 1640 1038
rect 1624 1031 1640 1036
rect 1614 1024 1620 1025
rect 1623 1024 1652 1031
rect 1541 1023 1652 1024
rect 1541 1022 1658 1023
rect 1217 1014 1268 1022
rect 1315 1014 1349 1022
rect 1217 1002 1242 1014
rect 1249 1002 1268 1014
rect 1322 1012 1349 1014
rect 1358 1012 1579 1022
rect 1614 1019 1620 1022
rect 1322 1008 1579 1012
rect 1217 994 1268 1002
rect 1315 994 1579 1008
rect 1623 1014 1658 1022
rect 1169 946 1188 980
rect 1233 986 1262 994
rect 1233 980 1250 986
rect 1233 978 1267 980
rect 1315 978 1331 994
rect 1332 984 1540 994
rect 1541 984 1557 994
rect 1605 990 1620 1005
rect 1623 1002 1624 1014
rect 1631 1002 1658 1014
rect 1623 994 1658 1002
rect 1623 993 1652 994
rect 1343 980 1557 984
rect 1358 978 1557 980
rect 1592 980 1605 990
rect 1623 980 1640 993
rect 1592 978 1640 980
rect 1234 974 1267 978
rect 1230 972 1267 974
rect 1230 971 1297 972
rect 1230 966 1261 971
rect 1267 966 1297 971
rect 1230 962 1297 966
rect 1203 959 1297 962
rect 1203 952 1252 959
rect 1203 946 1233 952
rect 1252 947 1257 952
rect 1169 930 1249 946
rect 1261 938 1297 959
rect 1358 954 1547 978
rect 1592 977 1639 978
rect 1605 972 1639 977
rect 1373 951 1547 954
rect 1366 948 1547 951
rect 1575 971 1639 972
rect 1169 928 1188 930
rect 1203 928 1237 930
rect 1169 912 1249 928
rect 1169 906 1188 912
rect 885 880 988 890
rect 839 878 988 880
rect 1009 878 1044 890
rect 678 876 840 878
rect 690 856 709 876
rect 724 874 754 876
rect 573 848 614 856
rect 696 852 709 856
rect 761 860 840 876
rect 872 876 1044 878
rect 872 860 951 876
rect 958 874 988 876
rect 536 838 565 848
rect 579 838 608 848
rect 623 838 653 852
rect 696 838 739 852
rect 761 848 951 860
rect 1016 856 1022 876
rect 746 838 776 848
rect 777 838 935 848
rect 939 838 969 848
rect 973 838 1003 852
rect 1031 838 1044 876
rect 1116 890 1145 906
rect 1159 890 1188 906
rect 1203 896 1233 912
rect 1261 890 1267 938
rect 1270 932 1289 938
rect 1304 932 1334 940
rect 1270 924 1334 932
rect 1270 908 1350 924
rect 1366 917 1428 948
rect 1444 917 1506 948
rect 1575 946 1624 971
rect 1639 946 1669 962
rect 1538 932 1568 940
rect 1575 938 1685 946
rect 1538 924 1583 932
rect 1270 906 1289 908
rect 1304 906 1350 908
rect 1270 890 1350 906
rect 1377 904 1412 917
rect 1453 914 1490 917
rect 1453 912 1495 914
rect 1382 901 1412 904
rect 1391 897 1398 901
rect 1398 896 1399 897
rect 1357 890 1367 896
rect 1116 882 1151 890
rect 1116 856 1117 882
rect 1124 856 1151 882
rect 1059 838 1089 852
rect 1116 848 1151 856
rect 1153 882 1194 890
rect 1153 856 1168 882
rect 1175 856 1194 882
rect 1258 878 1289 890
rect 1304 878 1407 890
rect 1419 880 1445 906
rect 1460 901 1490 912
rect 1522 908 1584 924
rect 1522 906 1568 908
rect 1522 890 1584 906
rect 1596 890 1602 938
rect 1605 930 1685 938
rect 1605 928 1624 930
rect 1639 928 1673 930
rect 1605 912 1685 928
rect 1605 890 1624 912
rect 1639 896 1669 912
rect 1697 906 1703 980
rect 1706 906 1725 1050
rect 1740 906 1746 1050
rect 1755 980 1768 1050
rect 1820 1046 1842 1050
rect 1813 1024 1842 1038
rect 1895 1024 1911 1038
rect 1949 1034 1955 1036
rect 1962 1034 2070 1050
rect 2077 1034 2083 1036
rect 2091 1034 2106 1050
rect 2172 1044 2191 1047
rect 1813 1022 1911 1024
rect 1938 1022 2106 1034
rect 2121 1024 2137 1038
rect 2172 1025 2194 1044
rect 2204 1038 2220 1039
rect 2203 1036 2220 1038
rect 2204 1031 2220 1036
rect 2194 1024 2200 1025
rect 2203 1024 2232 1031
rect 2121 1023 2232 1024
rect 2121 1022 2238 1023
rect 1797 1014 1848 1022
rect 1895 1014 1929 1022
rect 1797 1002 1822 1014
rect 1829 1002 1848 1014
rect 1902 1012 1929 1014
rect 1938 1012 2159 1022
rect 2194 1019 2200 1022
rect 1902 1008 2159 1012
rect 1797 994 1848 1002
rect 1895 994 2159 1008
rect 2203 1014 2238 1022
rect 1749 946 1768 980
rect 1813 986 1842 994
rect 1813 980 1830 986
rect 1813 978 1847 980
rect 1895 978 1911 994
rect 1912 984 2120 994
rect 2121 984 2137 994
rect 2185 990 2200 1005
rect 2203 1002 2204 1014
rect 2211 1002 2238 1014
rect 2203 994 2238 1002
rect 2203 993 2232 994
rect 1923 980 2137 984
rect 1938 978 2137 980
rect 2172 980 2185 990
rect 2203 980 2220 993
rect 2172 978 2220 980
rect 1814 974 1847 978
rect 1810 972 1847 974
rect 1810 971 1877 972
rect 1810 966 1841 971
rect 1847 966 1877 971
rect 1810 962 1877 966
rect 1783 959 1877 962
rect 1783 952 1832 959
rect 1783 946 1813 952
rect 1832 947 1837 952
rect 1749 930 1829 946
rect 1841 938 1877 959
rect 1938 954 2127 978
rect 2172 977 2219 978
rect 2185 972 2219 977
rect 1953 951 2127 954
rect 1946 948 2127 951
rect 2155 971 2219 972
rect 1749 928 1768 930
rect 1783 928 1817 930
rect 1749 912 1829 928
rect 1749 906 1768 912
rect 1465 880 1568 890
rect 1419 878 1568 880
rect 1589 878 1624 890
rect 1258 876 1420 878
rect 1270 856 1289 876
rect 1304 874 1334 876
rect 1153 848 1194 856
rect 1276 852 1289 856
rect 1341 860 1420 876
rect 1452 876 1624 878
rect 1452 860 1531 876
rect 1538 874 1568 876
rect 1116 838 1145 848
rect 1159 838 1188 848
rect 1203 838 1233 852
rect 1276 838 1319 852
rect 1341 848 1531 860
rect 1596 856 1602 876
rect 1326 838 1356 848
rect 1357 838 1515 848
rect 1519 838 1549 848
rect 1553 838 1583 852
rect 1611 838 1624 876
rect 1696 890 1725 906
rect 1739 890 1768 906
rect 1783 896 1813 912
rect 1841 890 1847 938
rect 1850 932 1869 938
rect 1884 932 1914 940
rect 1850 924 1914 932
rect 1850 908 1930 924
rect 1946 917 2008 948
rect 2024 917 2086 948
rect 2155 946 2204 971
rect 2219 946 2249 962
rect 2118 932 2148 940
rect 2155 938 2265 946
rect 2118 924 2163 932
rect 1850 906 1869 908
rect 1884 906 1930 908
rect 1850 890 1930 906
rect 1957 904 1992 917
rect 2033 914 2070 917
rect 2033 912 2075 914
rect 1962 901 1992 904
rect 1971 897 1978 901
rect 1978 896 1979 897
rect 1937 890 1947 896
rect 1696 882 1731 890
rect 1696 856 1697 882
rect 1704 856 1731 882
rect 1639 838 1669 852
rect 1696 848 1731 856
rect 1733 882 1774 890
rect 1733 856 1748 882
rect 1755 856 1774 882
rect 1838 878 1869 890
rect 1884 878 1987 890
rect 1999 880 2025 906
rect 2040 901 2070 912
rect 2102 908 2164 924
rect 2102 906 2148 908
rect 2102 890 2164 906
rect 2176 890 2182 938
rect 2185 930 2265 938
rect 2185 928 2204 930
rect 2219 928 2253 930
rect 2185 912 2265 928
rect 2185 890 2204 912
rect 2219 896 2249 912
rect 2277 906 2283 980
rect 2286 906 2305 1050
rect 2320 906 2326 1050
rect 2335 980 2348 1050
rect 2400 1046 2422 1050
rect 2393 1024 2422 1038
rect 2475 1024 2491 1038
rect 2529 1034 2535 1036
rect 2542 1034 2650 1050
rect 2657 1034 2663 1036
rect 2671 1034 2686 1050
rect 2752 1044 2771 1047
rect 2393 1022 2491 1024
rect 2518 1022 2686 1034
rect 2701 1024 2717 1038
rect 2752 1025 2774 1044
rect 2784 1038 2800 1039
rect 2783 1036 2800 1038
rect 2784 1031 2800 1036
rect 2774 1024 2780 1025
rect 2783 1024 2812 1031
rect 2701 1023 2812 1024
rect 2701 1022 2818 1023
rect 2377 1014 2428 1022
rect 2475 1014 2509 1022
rect 2377 1002 2402 1014
rect 2409 1002 2428 1014
rect 2482 1012 2509 1014
rect 2518 1012 2739 1022
rect 2774 1019 2780 1022
rect 2482 1008 2739 1012
rect 2377 994 2428 1002
rect 2475 994 2739 1008
rect 2783 1014 2818 1022
rect 2329 946 2348 980
rect 2393 986 2422 994
rect 2393 980 2410 986
rect 2393 978 2427 980
rect 2475 978 2491 994
rect 2492 984 2700 994
rect 2701 984 2717 994
rect 2765 990 2780 1005
rect 2783 1002 2784 1014
rect 2791 1002 2818 1014
rect 2783 994 2818 1002
rect 2783 993 2812 994
rect 2503 980 2717 984
rect 2518 978 2717 980
rect 2752 980 2765 990
rect 2783 980 2800 993
rect 2752 978 2800 980
rect 2394 974 2427 978
rect 2390 972 2427 974
rect 2390 971 2457 972
rect 2390 966 2421 971
rect 2427 966 2457 971
rect 2390 962 2457 966
rect 2363 959 2457 962
rect 2363 952 2412 959
rect 2363 946 2393 952
rect 2412 947 2417 952
rect 2329 930 2409 946
rect 2421 938 2457 959
rect 2518 954 2707 978
rect 2752 977 2799 978
rect 2765 972 2799 977
rect 2533 951 2707 954
rect 2526 948 2707 951
rect 2735 971 2799 972
rect 2329 928 2348 930
rect 2363 928 2397 930
rect 2329 912 2409 928
rect 2329 906 2348 912
rect 2045 880 2148 890
rect 1999 878 2148 880
rect 2169 878 2204 890
rect 1838 876 2000 878
rect 1850 856 1869 876
rect 1884 874 1914 876
rect 1733 848 1774 856
rect 1856 852 1869 856
rect 1921 860 2000 876
rect 2032 876 2204 878
rect 2032 860 2111 876
rect 2118 874 2148 876
rect 1696 838 1725 848
rect 1739 838 1768 848
rect 1783 838 1813 852
rect 1856 838 1899 852
rect 1921 848 2111 860
rect 2176 856 2182 876
rect 1906 838 1936 848
rect 1937 838 2095 848
rect 2099 838 2129 848
rect 2133 838 2163 852
rect 2191 838 2204 876
rect 2276 890 2305 906
rect 2319 890 2348 906
rect 2363 896 2393 912
rect 2421 890 2427 938
rect 2430 932 2449 938
rect 2464 932 2494 940
rect 2430 924 2494 932
rect 2430 908 2510 924
rect 2526 917 2588 948
rect 2604 917 2666 948
rect 2735 946 2784 971
rect 2799 946 2829 962
rect 2698 932 2728 940
rect 2735 938 2845 946
rect 2698 924 2743 932
rect 2430 906 2449 908
rect 2464 906 2510 908
rect 2430 890 2510 906
rect 2537 904 2572 917
rect 2613 914 2650 917
rect 2613 912 2655 914
rect 2542 901 2572 904
rect 2551 897 2558 901
rect 2558 896 2559 897
rect 2517 890 2527 896
rect 2276 882 2311 890
rect 2276 856 2277 882
rect 2284 856 2311 882
rect 2219 838 2249 852
rect 2276 848 2311 856
rect 2313 882 2354 890
rect 2313 856 2328 882
rect 2335 856 2354 882
rect 2418 878 2449 890
rect 2464 878 2567 890
rect 2579 880 2605 906
rect 2620 901 2650 912
rect 2682 908 2744 924
rect 2682 906 2728 908
rect 2682 890 2744 906
rect 2756 890 2762 938
rect 2765 930 2845 938
rect 2765 928 2784 930
rect 2799 928 2833 930
rect 2765 912 2845 928
rect 2765 890 2784 912
rect 2799 896 2829 912
rect 2857 906 2863 980
rect 2866 906 2885 1050
rect 2900 906 2906 1050
rect 2915 980 2928 1050
rect 2980 1046 3002 1050
rect 2973 1024 3002 1038
rect 3055 1024 3071 1038
rect 3109 1034 3115 1036
rect 3122 1034 3230 1050
rect 3237 1034 3243 1036
rect 3251 1034 3266 1050
rect 3332 1044 3351 1047
rect 2973 1022 3071 1024
rect 3098 1022 3266 1034
rect 3281 1024 3297 1038
rect 3332 1025 3354 1044
rect 3364 1038 3380 1039
rect 3363 1036 3380 1038
rect 3364 1031 3380 1036
rect 3354 1024 3360 1025
rect 3363 1024 3392 1031
rect 3281 1023 3392 1024
rect 3281 1022 3398 1023
rect 2957 1014 3008 1022
rect 3055 1014 3089 1022
rect 2957 1002 2982 1014
rect 2989 1002 3008 1014
rect 3062 1012 3089 1014
rect 3098 1012 3319 1022
rect 3354 1019 3360 1022
rect 3062 1008 3319 1012
rect 2957 994 3008 1002
rect 3055 994 3319 1008
rect 3363 1014 3398 1022
rect 2909 946 2928 980
rect 2973 986 3002 994
rect 2973 980 2990 986
rect 2973 978 3007 980
rect 3055 978 3071 994
rect 3072 984 3280 994
rect 3281 984 3297 994
rect 3345 990 3360 1005
rect 3363 1002 3364 1014
rect 3371 1002 3398 1014
rect 3363 994 3398 1002
rect 3363 993 3392 994
rect 3083 980 3297 984
rect 3098 978 3297 980
rect 3332 980 3345 990
rect 3363 980 3380 993
rect 3332 978 3380 980
rect 2974 974 3007 978
rect 2970 972 3007 974
rect 2970 971 3037 972
rect 2970 966 3001 971
rect 3007 966 3037 971
rect 2970 962 3037 966
rect 2943 959 3037 962
rect 2943 952 2992 959
rect 2943 946 2973 952
rect 2992 947 2997 952
rect 2909 930 2989 946
rect 3001 938 3037 959
rect 3098 954 3287 978
rect 3332 977 3379 978
rect 3345 972 3379 977
rect 3113 951 3287 954
rect 3106 948 3287 951
rect 3315 971 3379 972
rect 2909 928 2928 930
rect 2943 928 2977 930
rect 2909 912 2989 928
rect 2909 906 2928 912
rect 2625 880 2728 890
rect 2579 878 2728 880
rect 2749 878 2784 890
rect 2418 876 2580 878
rect 2430 856 2449 876
rect 2464 874 2494 876
rect 2313 848 2354 856
rect 2436 852 2449 856
rect 2501 860 2580 876
rect 2612 876 2784 878
rect 2612 860 2691 876
rect 2698 874 2728 876
rect 2276 838 2305 848
rect 2319 838 2348 848
rect 2363 838 2393 852
rect 2436 838 2479 852
rect 2501 848 2691 860
rect 2756 856 2762 876
rect 2486 838 2516 848
rect 2517 838 2675 848
rect 2679 838 2709 848
rect 2713 838 2743 852
rect 2771 838 2784 876
rect 2856 890 2885 906
rect 2899 890 2928 906
rect 2943 896 2973 912
rect 3001 890 3007 938
rect 3010 932 3029 938
rect 3044 932 3074 940
rect 3010 924 3074 932
rect 3010 908 3090 924
rect 3106 917 3168 948
rect 3184 917 3246 948
rect 3315 946 3364 971
rect 3379 946 3409 962
rect 3278 932 3308 940
rect 3315 938 3425 946
rect 3278 924 3323 932
rect 3010 906 3029 908
rect 3044 906 3090 908
rect 3010 890 3090 906
rect 3117 904 3152 917
rect 3193 914 3230 917
rect 3193 912 3235 914
rect 3122 901 3152 904
rect 3131 897 3138 901
rect 3138 896 3139 897
rect 3097 890 3107 896
rect 2856 882 2891 890
rect 2856 856 2857 882
rect 2864 856 2891 882
rect 2799 838 2829 852
rect 2856 848 2891 856
rect 2893 882 2934 890
rect 2893 856 2908 882
rect 2915 856 2934 882
rect 2998 878 3029 890
rect 3044 878 3147 890
rect 3159 880 3185 906
rect 3200 901 3230 912
rect 3262 908 3324 924
rect 3262 906 3308 908
rect 3262 890 3324 906
rect 3336 890 3342 938
rect 3345 930 3425 938
rect 3345 928 3364 930
rect 3379 928 3413 930
rect 3345 912 3425 928
rect 3345 890 3364 912
rect 3379 896 3409 912
rect 3437 906 3443 980
rect 3446 906 3465 1050
rect 3480 906 3486 1050
rect 3495 980 3508 1050
rect 3560 1046 3582 1050
rect 3553 1024 3582 1038
rect 3635 1024 3651 1038
rect 3689 1034 3695 1036
rect 3702 1034 3810 1050
rect 3817 1034 3823 1036
rect 3831 1034 3846 1050
rect 3912 1044 3931 1047
rect 3553 1022 3651 1024
rect 3678 1022 3846 1034
rect 3861 1024 3877 1038
rect 3912 1025 3934 1044
rect 3944 1038 3960 1039
rect 3943 1036 3960 1038
rect 3944 1031 3960 1036
rect 3934 1024 3940 1025
rect 3943 1024 3972 1031
rect 3861 1023 3972 1024
rect 3861 1022 3978 1023
rect 3537 1014 3588 1022
rect 3635 1014 3669 1022
rect 3537 1002 3562 1014
rect 3569 1002 3588 1014
rect 3642 1012 3669 1014
rect 3678 1012 3899 1022
rect 3934 1019 3940 1022
rect 3642 1008 3899 1012
rect 3537 994 3588 1002
rect 3635 994 3899 1008
rect 3943 1014 3978 1022
rect 3489 946 3508 980
rect 3553 986 3582 994
rect 3553 980 3570 986
rect 3553 978 3587 980
rect 3635 978 3651 994
rect 3652 984 3860 994
rect 3861 984 3877 994
rect 3925 990 3940 1005
rect 3943 1002 3944 1014
rect 3951 1002 3978 1014
rect 3943 994 3978 1002
rect 3943 993 3972 994
rect 3663 980 3877 984
rect 3678 978 3877 980
rect 3912 980 3925 990
rect 3943 980 3960 993
rect 3912 978 3960 980
rect 3554 974 3587 978
rect 3550 972 3587 974
rect 3550 971 3617 972
rect 3550 966 3581 971
rect 3587 966 3617 971
rect 3550 962 3617 966
rect 3523 959 3617 962
rect 3523 952 3572 959
rect 3523 946 3553 952
rect 3572 947 3577 952
rect 3489 930 3569 946
rect 3581 938 3617 959
rect 3678 954 3867 978
rect 3912 977 3959 978
rect 3925 972 3959 977
rect 3693 951 3867 954
rect 3686 948 3867 951
rect 3895 971 3959 972
rect 3489 928 3508 930
rect 3523 928 3557 930
rect 3489 912 3569 928
rect 3489 906 3508 912
rect 3205 880 3308 890
rect 3159 878 3308 880
rect 3329 878 3364 890
rect 2998 876 3160 878
rect 3010 856 3029 876
rect 3044 874 3074 876
rect 2893 848 2934 856
rect 3016 852 3029 856
rect 3081 860 3160 876
rect 3192 876 3364 878
rect 3192 860 3271 876
rect 3278 874 3308 876
rect 2856 838 2885 848
rect 2899 838 2928 848
rect 2943 838 2973 852
rect 3016 838 3059 852
rect 3081 848 3271 860
rect 3336 856 3342 876
rect 3066 838 3096 848
rect 3097 838 3255 848
rect 3259 838 3289 848
rect 3293 838 3323 852
rect 3351 838 3364 876
rect 3436 890 3465 906
rect 3479 890 3508 906
rect 3523 896 3553 912
rect 3581 890 3587 938
rect 3590 932 3609 938
rect 3624 932 3654 940
rect 3590 924 3654 932
rect 3590 908 3670 924
rect 3686 917 3748 948
rect 3764 917 3826 948
rect 3895 946 3944 971
rect 3959 946 3989 962
rect 3858 932 3888 940
rect 3895 938 4005 946
rect 3858 924 3903 932
rect 3590 906 3609 908
rect 3624 906 3670 908
rect 3590 890 3670 906
rect 3697 904 3732 917
rect 3773 914 3810 917
rect 3773 912 3815 914
rect 3702 901 3732 904
rect 3711 897 3718 901
rect 3718 896 3719 897
rect 3677 890 3687 896
rect 3436 882 3471 890
rect 3436 856 3437 882
rect 3444 856 3471 882
rect 3379 838 3409 852
rect 3436 848 3471 856
rect 3473 882 3514 890
rect 3473 856 3488 882
rect 3495 856 3514 882
rect 3578 878 3609 890
rect 3624 878 3727 890
rect 3739 880 3765 906
rect 3780 901 3810 912
rect 3842 908 3904 924
rect 3842 906 3888 908
rect 3842 890 3904 906
rect 3916 890 3922 938
rect 3925 930 4005 938
rect 3925 928 3944 930
rect 3959 928 3993 930
rect 3925 912 4005 928
rect 3925 890 3944 912
rect 3959 896 3989 912
rect 4017 906 4023 980
rect 4026 906 4045 1050
rect 4060 906 4066 1050
rect 4075 980 4088 1050
rect 4140 1046 4162 1050
rect 4133 1024 4162 1038
rect 4215 1024 4231 1038
rect 4269 1034 4275 1036
rect 4282 1034 4390 1050
rect 4397 1034 4403 1036
rect 4411 1034 4426 1050
rect 4492 1044 4511 1047
rect 4133 1022 4231 1024
rect 4258 1022 4426 1034
rect 4441 1024 4457 1038
rect 4492 1025 4514 1044
rect 4524 1038 4540 1039
rect 4523 1036 4540 1038
rect 4524 1031 4540 1036
rect 4514 1024 4520 1025
rect 4523 1024 4552 1031
rect 4441 1023 4552 1024
rect 4441 1022 4558 1023
rect 4117 1014 4168 1022
rect 4215 1014 4249 1022
rect 4117 1002 4142 1014
rect 4149 1002 4168 1014
rect 4222 1012 4249 1014
rect 4258 1012 4479 1022
rect 4514 1019 4520 1022
rect 4222 1008 4479 1012
rect 4117 994 4168 1002
rect 4215 994 4479 1008
rect 4523 1014 4558 1022
rect 4069 946 4088 980
rect 4133 986 4162 994
rect 4133 980 4150 986
rect 4133 978 4167 980
rect 4215 978 4231 994
rect 4232 984 4440 994
rect 4441 984 4457 994
rect 4505 990 4520 1005
rect 4523 1002 4524 1014
rect 4531 1002 4558 1014
rect 4523 994 4558 1002
rect 4523 993 4552 994
rect 4243 980 4457 984
rect 4258 978 4457 980
rect 4492 980 4505 990
rect 4523 980 4540 993
rect 4492 978 4540 980
rect 4134 974 4167 978
rect 4130 972 4167 974
rect 4130 971 4197 972
rect 4130 966 4161 971
rect 4167 966 4197 971
rect 4130 962 4197 966
rect 4103 959 4197 962
rect 4103 952 4152 959
rect 4103 946 4133 952
rect 4152 947 4157 952
rect 4069 930 4149 946
rect 4161 938 4197 959
rect 4258 954 4447 978
rect 4492 977 4539 978
rect 4505 972 4539 977
rect 4273 951 4447 954
rect 4266 948 4447 951
rect 4475 971 4539 972
rect 4069 928 4088 930
rect 4103 928 4137 930
rect 4069 912 4149 928
rect 4069 906 4088 912
rect 3785 880 3888 890
rect 3739 878 3888 880
rect 3909 878 3944 890
rect 3578 876 3740 878
rect 3590 856 3609 876
rect 3624 874 3654 876
rect 3473 848 3514 856
rect 3596 852 3609 856
rect 3661 860 3740 876
rect 3772 876 3944 878
rect 3772 860 3851 876
rect 3858 874 3888 876
rect 3436 838 3465 848
rect 3479 838 3508 848
rect 3523 838 3553 852
rect 3596 838 3639 852
rect 3661 848 3851 860
rect 3916 856 3922 876
rect 3646 838 3676 848
rect 3677 838 3835 848
rect 3839 838 3869 848
rect 3873 838 3903 852
rect 3931 838 3944 876
rect 4016 890 4045 906
rect 4059 890 4088 906
rect 4103 896 4133 912
rect 4161 890 4167 938
rect 4170 932 4189 938
rect 4204 932 4234 940
rect 4170 924 4234 932
rect 4170 908 4250 924
rect 4266 917 4328 948
rect 4344 917 4406 948
rect 4475 946 4524 971
rect 4539 946 4569 962
rect 4438 932 4468 940
rect 4475 938 4585 946
rect 4438 924 4483 932
rect 4170 906 4189 908
rect 4204 906 4250 908
rect 4170 890 4250 906
rect 4277 904 4312 917
rect 4353 914 4390 917
rect 4353 912 4395 914
rect 4282 901 4312 904
rect 4291 897 4298 901
rect 4298 896 4299 897
rect 4257 890 4267 896
rect 4016 882 4051 890
rect 4016 856 4017 882
rect 4024 856 4051 882
rect 3959 838 3989 852
rect 4016 848 4051 856
rect 4053 882 4094 890
rect 4053 856 4068 882
rect 4075 856 4094 882
rect 4158 878 4189 890
rect 4204 878 4307 890
rect 4319 880 4345 906
rect 4360 901 4390 912
rect 4422 908 4484 924
rect 4422 906 4468 908
rect 4422 890 4484 906
rect 4496 890 4502 938
rect 4505 930 4585 938
rect 4505 928 4524 930
rect 4539 928 4573 930
rect 4505 912 4585 928
rect 4505 890 4524 912
rect 4539 896 4569 912
rect 4597 906 4603 980
rect 4606 906 4625 1050
rect 4640 906 4646 1050
rect 4655 980 4668 1050
rect 4720 1046 4742 1050
rect 4713 1024 4742 1038
rect 4795 1024 4811 1038
rect 4849 1034 4855 1036
rect 4862 1034 4970 1050
rect 4977 1034 4983 1036
rect 4991 1034 5006 1050
rect 5072 1044 5091 1047
rect 4713 1022 4811 1024
rect 4838 1022 5006 1034
rect 5021 1024 5037 1038
rect 5072 1025 5094 1044
rect 5104 1038 5120 1039
rect 5103 1036 5120 1038
rect 5104 1031 5120 1036
rect 5094 1024 5100 1025
rect 5103 1024 5132 1031
rect 5021 1023 5132 1024
rect 5021 1022 5138 1023
rect 4697 1014 4748 1022
rect 4795 1014 4829 1022
rect 4697 1002 4722 1014
rect 4729 1002 4748 1014
rect 4802 1012 4829 1014
rect 4838 1012 5059 1022
rect 5094 1019 5100 1022
rect 4802 1008 5059 1012
rect 4697 994 4748 1002
rect 4795 994 5059 1008
rect 5103 1014 5138 1022
rect 4649 946 4668 980
rect 4713 986 4742 994
rect 4713 980 4730 986
rect 4713 978 4747 980
rect 4795 978 4811 994
rect 4812 984 5020 994
rect 5021 984 5037 994
rect 5085 990 5100 1005
rect 5103 1002 5104 1014
rect 5111 1002 5138 1014
rect 5103 994 5138 1002
rect 5103 993 5132 994
rect 4823 980 5037 984
rect 4838 978 5037 980
rect 5072 980 5085 990
rect 5103 980 5120 993
rect 5072 978 5120 980
rect 4714 974 4747 978
rect 4710 972 4747 974
rect 4710 971 4777 972
rect 4710 966 4741 971
rect 4747 966 4777 971
rect 4710 962 4777 966
rect 4683 959 4777 962
rect 4683 952 4732 959
rect 4683 946 4713 952
rect 4732 947 4737 952
rect 4649 930 4729 946
rect 4741 938 4777 959
rect 4838 954 5027 978
rect 5072 977 5119 978
rect 5085 972 5119 977
rect 4853 951 5027 954
rect 4846 948 5027 951
rect 5055 971 5119 972
rect 4649 928 4668 930
rect 4683 928 4717 930
rect 4649 912 4729 928
rect 4649 906 4668 912
rect 4365 880 4468 890
rect 4319 878 4468 880
rect 4489 878 4524 890
rect 4158 876 4320 878
rect 4170 856 4189 876
rect 4204 874 4234 876
rect 4053 848 4094 856
rect 4176 852 4189 856
rect 4241 860 4320 876
rect 4352 876 4524 878
rect 4352 860 4431 876
rect 4438 874 4468 876
rect 4016 838 4045 848
rect 4059 838 4088 848
rect 4103 838 4133 852
rect 4176 838 4219 852
rect 4241 848 4431 860
rect 4496 856 4502 876
rect 4226 838 4256 848
rect 4257 838 4415 848
rect 4419 838 4449 848
rect 4453 838 4483 852
rect 4511 838 4524 876
rect 4596 890 4625 906
rect 4639 890 4668 906
rect 4683 896 4713 912
rect 4741 890 4747 938
rect 4750 932 4769 938
rect 4784 932 4814 940
rect 4750 924 4814 932
rect 4750 908 4830 924
rect 4846 917 4908 948
rect 4924 917 4986 948
rect 5055 946 5104 971
rect 5119 946 5149 962
rect 5018 932 5048 940
rect 5055 938 5165 946
rect 5018 924 5063 932
rect 4750 906 4769 908
rect 4784 906 4830 908
rect 4750 890 4830 906
rect 4857 904 4892 917
rect 4933 914 4970 917
rect 4933 912 4975 914
rect 4862 901 4892 904
rect 4871 897 4878 901
rect 4878 896 4879 897
rect 4837 890 4847 896
rect 4596 882 4631 890
rect 4596 856 4597 882
rect 4604 856 4631 882
rect 4539 838 4569 852
rect 4596 848 4631 856
rect 4633 882 4674 890
rect 4633 856 4648 882
rect 4655 856 4674 882
rect 4738 878 4769 890
rect 4784 878 4887 890
rect 4899 880 4925 906
rect 4940 901 4970 912
rect 5002 908 5064 924
rect 5002 906 5048 908
rect 5002 890 5064 906
rect 5076 890 5082 938
rect 5085 930 5165 938
rect 5085 928 5104 930
rect 5119 928 5153 930
rect 5085 912 5165 928
rect 5085 890 5104 912
rect 5119 896 5149 912
rect 5177 906 5183 980
rect 5186 906 5205 1050
rect 5220 906 5226 1050
rect 5235 980 5248 1050
rect 5300 1046 5322 1050
rect 5293 1024 5322 1038
rect 5375 1024 5391 1038
rect 5429 1034 5435 1036
rect 5442 1034 5550 1050
rect 5557 1034 5563 1036
rect 5571 1034 5586 1050
rect 5652 1044 5671 1047
rect 5293 1022 5391 1024
rect 5418 1022 5586 1034
rect 5601 1024 5617 1038
rect 5652 1025 5674 1044
rect 5684 1038 5700 1039
rect 5683 1036 5700 1038
rect 5684 1031 5700 1036
rect 5674 1024 5680 1025
rect 5683 1024 5712 1031
rect 5601 1023 5712 1024
rect 5601 1022 5718 1023
rect 5277 1014 5328 1022
rect 5375 1014 5409 1022
rect 5277 1002 5302 1014
rect 5309 1002 5328 1014
rect 5382 1012 5409 1014
rect 5418 1012 5639 1022
rect 5674 1019 5680 1022
rect 5382 1008 5639 1012
rect 5277 994 5328 1002
rect 5375 994 5639 1008
rect 5683 1014 5718 1022
rect 5229 946 5248 980
rect 5293 986 5322 994
rect 5293 980 5310 986
rect 5293 978 5327 980
rect 5375 978 5391 994
rect 5392 984 5600 994
rect 5601 984 5617 994
rect 5665 990 5680 1005
rect 5683 1002 5684 1014
rect 5691 1002 5718 1014
rect 5683 994 5718 1002
rect 5683 993 5712 994
rect 5403 980 5617 984
rect 5418 978 5617 980
rect 5652 980 5665 990
rect 5683 980 5700 993
rect 5652 978 5700 980
rect 5294 974 5327 978
rect 5290 972 5327 974
rect 5290 971 5357 972
rect 5290 966 5321 971
rect 5327 966 5357 971
rect 5290 962 5357 966
rect 5263 959 5357 962
rect 5263 952 5312 959
rect 5263 946 5293 952
rect 5312 947 5317 952
rect 5229 930 5309 946
rect 5321 938 5357 959
rect 5418 954 5607 978
rect 5652 977 5699 978
rect 5665 972 5699 977
rect 5433 951 5607 954
rect 5426 948 5607 951
rect 5635 971 5699 972
rect 5229 928 5248 930
rect 5263 928 5297 930
rect 5229 912 5309 928
rect 5229 906 5248 912
rect 4945 880 5048 890
rect 4899 878 5048 880
rect 5069 878 5104 890
rect 4738 876 4900 878
rect 4750 856 4769 876
rect 4784 874 4814 876
rect 4633 848 4674 856
rect 4756 852 4769 856
rect 4821 860 4900 876
rect 4932 876 5104 878
rect 4932 860 5011 876
rect 5018 874 5048 876
rect 4596 838 4625 848
rect 4639 838 4668 848
rect 4683 838 4713 852
rect 4756 838 4799 852
rect 4821 848 5011 860
rect 5076 856 5082 876
rect 4806 838 4836 848
rect 4837 838 4995 848
rect 4999 838 5029 848
rect 5033 838 5063 852
rect 5091 838 5104 876
rect 5176 890 5205 906
rect 5219 890 5248 906
rect 5263 896 5293 912
rect 5321 890 5327 938
rect 5330 932 5349 938
rect 5364 932 5394 940
rect 5330 924 5394 932
rect 5330 908 5410 924
rect 5426 917 5488 948
rect 5504 917 5566 948
rect 5635 946 5684 971
rect 5699 946 5729 962
rect 5598 932 5628 940
rect 5635 938 5745 946
rect 5598 924 5643 932
rect 5330 906 5349 908
rect 5364 906 5410 908
rect 5330 890 5410 906
rect 5437 904 5472 917
rect 5513 914 5550 917
rect 5513 912 5555 914
rect 5442 901 5472 904
rect 5451 897 5458 901
rect 5458 896 5459 897
rect 5417 890 5427 896
rect 5176 882 5211 890
rect 5176 856 5177 882
rect 5184 856 5211 882
rect 5119 838 5149 852
rect 5176 848 5211 856
rect 5213 882 5254 890
rect 5213 856 5228 882
rect 5235 856 5254 882
rect 5318 878 5349 890
rect 5364 878 5467 890
rect 5479 880 5505 906
rect 5520 901 5550 912
rect 5582 908 5644 924
rect 5582 906 5628 908
rect 5582 890 5644 906
rect 5656 890 5662 938
rect 5665 930 5745 938
rect 5665 928 5684 930
rect 5699 928 5733 930
rect 5665 912 5745 928
rect 5665 890 5684 912
rect 5699 896 5729 912
rect 5757 906 5763 980
rect 5766 906 5785 1050
rect 5800 906 5806 1050
rect 5815 980 5828 1050
rect 5880 1046 5902 1050
rect 5873 1024 5902 1038
rect 5955 1024 5971 1038
rect 6009 1034 6015 1036
rect 6022 1034 6130 1050
rect 6137 1034 6143 1036
rect 6151 1034 6166 1050
rect 6232 1044 6251 1047
rect 5873 1022 5971 1024
rect 5998 1022 6166 1034
rect 6181 1024 6197 1038
rect 6232 1025 6254 1044
rect 6264 1038 6280 1039
rect 6263 1036 6280 1038
rect 6264 1031 6280 1036
rect 6254 1024 6260 1025
rect 6263 1024 6292 1031
rect 6181 1023 6292 1024
rect 6181 1022 6298 1023
rect 5857 1014 5908 1022
rect 5955 1014 5989 1022
rect 5857 1002 5882 1014
rect 5889 1002 5908 1014
rect 5962 1012 5989 1014
rect 5998 1012 6219 1022
rect 6254 1019 6260 1022
rect 5962 1008 6219 1012
rect 5857 994 5908 1002
rect 5955 994 6219 1008
rect 6263 1014 6298 1022
rect 5809 946 5828 980
rect 5873 986 5902 994
rect 5873 980 5890 986
rect 5873 978 5907 980
rect 5955 978 5971 994
rect 5972 984 6180 994
rect 6181 984 6197 994
rect 6245 990 6260 1005
rect 6263 1002 6264 1014
rect 6271 1002 6298 1014
rect 6263 994 6298 1002
rect 6263 993 6292 994
rect 5983 980 6197 984
rect 5998 978 6197 980
rect 6232 980 6245 990
rect 6263 980 6280 993
rect 6232 978 6280 980
rect 5874 974 5907 978
rect 5870 972 5907 974
rect 5870 971 5937 972
rect 5870 966 5901 971
rect 5907 966 5937 971
rect 5870 962 5937 966
rect 5843 959 5937 962
rect 5843 952 5892 959
rect 5843 946 5873 952
rect 5892 947 5897 952
rect 5809 930 5889 946
rect 5901 938 5937 959
rect 5998 954 6187 978
rect 6232 977 6279 978
rect 6245 972 6279 977
rect 6013 951 6187 954
rect 6006 948 6187 951
rect 6215 971 6279 972
rect 5809 928 5828 930
rect 5843 928 5877 930
rect 5809 912 5889 928
rect 5809 906 5828 912
rect 5525 880 5628 890
rect 5479 878 5628 880
rect 5649 878 5684 890
rect 5318 876 5480 878
rect 5330 856 5349 876
rect 5364 874 5394 876
rect 5213 848 5254 856
rect 5336 852 5349 856
rect 5401 860 5480 876
rect 5512 876 5684 878
rect 5512 860 5591 876
rect 5598 874 5628 876
rect 5176 838 5205 848
rect 5219 838 5248 848
rect 5263 838 5293 852
rect 5336 838 5379 852
rect 5401 848 5591 860
rect 5656 856 5662 876
rect 5386 838 5416 848
rect 5417 838 5575 848
rect 5579 838 5609 848
rect 5613 838 5643 852
rect 5671 838 5684 876
rect 5756 890 5785 906
rect 5799 890 5828 906
rect 5843 896 5873 912
rect 5901 890 5907 938
rect 5910 932 5929 938
rect 5944 932 5974 940
rect 5910 924 5974 932
rect 5910 908 5990 924
rect 6006 917 6068 948
rect 6084 917 6146 948
rect 6215 946 6264 971
rect 6279 946 6309 962
rect 6178 932 6208 940
rect 6215 938 6325 946
rect 6178 924 6223 932
rect 5910 906 5929 908
rect 5944 906 5990 908
rect 5910 890 5990 906
rect 6017 904 6052 917
rect 6093 914 6130 917
rect 6093 912 6135 914
rect 6022 901 6052 904
rect 6031 897 6038 901
rect 6038 896 6039 897
rect 5997 890 6007 896
rect 5756 882 5791 890
rect 5756 856 5757 882
rect 5764 856 5791 882
rect 5699 838 5729 852
rect 5756 848 5791 856
rect 5793 882 5834 890
rect 5793 856 5808 882
rect 5815 856 5834 882
rect 5898 878 5929 890
rect 5944 878 6047 890
rect 6059 880 6085 906
rect 6100 901 6130 912
rect 6162 908 6224 924
rect 6162 906 6208 908
rect 6162 890 6224 906
rect 6236 890 6242 938
rect 6245 930 6325 938
rect 6245 928 6264 930
rect 6279 928 6313 930
rect 6245 912 6325 928
rect 6245 890 6264 912
rect 6279 896 6309 912
rect 6337 906 6343 980
rect 6346 906 6365 1050
rect 6380 906 6386 1050
rect 6395 980 6408 1050
rect 6460 1046 6482 1050
rect 6453 1024 6482 1038
rect 6535 1024 6551 1038
rect 6589 1034 6595 1036
rect 6602 1034 6710 1050
rect 6717 1034 6723 1036
rect 6731 1034 6746 1050
rect 6812 1044 6831 1047
rect 6453 1022 6551 1024
rect 6578 1022 6746 1034
rect 6761 1024 6777 1038
rect 6812 1025 6834 1044
rect 6844 1038 6860 1039
rect 6843 1036 6860 1038
rect 6844 1031 6860 1036
rect 6834 1024 6840 1025
rect 6843 1024 6872 1031
rect 6761 1023 6872 1024
rect 6761 1022 6878 1023
rect 6437 1014 6488 1022
rect 6535 1014 6569 1022
rect 6437 1002 6462 1014
rect 6469 1002 6488 1014
rect 6542 1012 6569 1014
rect 6578 1012 6799 1022
rect 6834 1019 6840 1022
rect 6542 1008 6799 1012
rect 6437 994 6488 1002
rect 6535 994 6799 1008
rect 6843 1014 6878 1022
rect 6389 946 6408 980
rect 6453 986 6482 994
rect 6453 980 6470 986
rect 6453 978 6487 980
rect 6535 978 6551 994
rect 6552 984 6760 994
rect 6761 984 6777 994
rect 6825 990 6840 1005
rect 6843 1002 6844 1014
rect 6851 1002 6878 1014
rect 6843 994 6878 1002
rect 6843 993 6872 994
rect 6563 980 6777 984
rect 6578 978 6777 980
rect 6812 980 6825 990
rect 6843 980 6860 993
rect 6812 978 6860 980
rect 6454 974 6487 978
rect 6450 972 6487 974
rect 6450 971 6517 972
rect 6450 966 6481 971
rect 6487 966 6517 971
rect 6450 962 6517 966
rect 6423 959 6517 962
rect 6423 952 6472 959
rect 6423 946 6453 952
rect 6472 947 6477 952
rect 6389 930 6469 946
rect 6481 938 6517 959
rect 6578 954 6767 978
rect 6812 977 6859 978
rect 6825 972 6859 977
rect 6593 951 6767 954
rect 6586 948 6767 951
rect 6795 971 6859 972
rect 6389 928 6408 930
rect 6423 928 6457 930
rect 6389 912 6469 928
rect 6389 906 6408 912
rect 6105 880 6208 890
rect 6059 878 6208 880
rect 6229 878 6264 890
rect 5898 876 6060 878
rect 5910 856 5929 876
rect 5944 874 5974 876
rect 5793 848 5834 856
rect 5916 852 5929 856
rect 5981 860 6060 876
rect 6092 876 6264 878
rect 6092 860 6171 876
rect 6178 874 6208 876
rect 5756 838 5785 848
rect 5799 838 5828 848
rect 5843 838 5873 852
rect 5916 838 5959 852
rect 5981 848 6171 860
rect 6236 856 6242 876
rect 5966 838 5996 848
rect 5997 838 6155 848
rect 6159 838 6189 848
rect 6193 838 6223 852
rect 6251 838 6264 876
rect 6336 890 6365 906
rect 6379 890 6408 906
rect 6423 896 6453 912
rect 6481 890 6487 938
rect 6490 932 6509 938
rect 6524 932 6554 940
rect 6490 924 6554 932
rect 6490 908 6570 924
rect 6586 917 6648 948
rect 6664 917 6726 948
rect 6795 946 6844 971
rect 6859 946 6889 962
rect 6758 932 6788 940
rect 6795 938 6905 946
rect 6758 924 6803 932
rect 6490 906 6509 908
rect 6524 906 6570 908
rect 6490 890 6570 906
rect 6597 904 6632 917
rect 6673 914 6710 917
rect 6673 912 6715 914
rect 6602 901 6632 904
rect 6611 897 6618 901
rect 6618 896 6619 897
rect 6577 890 6587 896
rect 6336 882 6371 890
rect 6336 856 6337 882
rect 6344 856 6371 882
rect 6279 838 6309 852
rect 6336 848 6371 856
rect 6373 882 6414 890
rect 6373 856 6388 882
rect 6395 856 6414 882
rect 6478 878 6509 890
rect 6524 878 6627 890
rect 6639 880 6665 906
rect 6680 901 6710 912
rect 6742 908 6804 924
rect 6742 906 6788 908
rect 6742 890 6804 906
rect 6816 890 6822 938
rect 6825 930 6905 938
rect 6825 928 6844 930
rect 6859 928 6893 930
rect 6825 912 6905 928
rect 6825 890 6844 912
rect 6859 896 6889 912
rect 6917 906 6923 980
rect 6926 906 6945 1050
rect 6960 906 6966 1050
rect 6975 980 6988 1050
rect 7040 1046 7062 1050
rect 7033 1024 7062 1038
rect 7115 1024 7131 1038
rect 7169 1034 7175 1036
rect 7182 1034 7290 1050
rect 7297 1034 7303 1036
rect 7311 1034 7326 1050
rect 7392 1044 7411 1047
rect 7033 1022 7131 1024
rect 7158 1022 7326 1034
rect 7341 1024 7357 1038
rect 7392 1025 7414 1044
rect 7424 1038 7440 1039
rect 7423 1036 7440 1038
rect 7424 1031 7440 1036
rect 7414 1024 7420 1025
rect 7423 1024 7452 1031
rect 7341 1023 7452 1024
rect 7341 1022 7458 1023
rect 7017 1014 7068 1022
rect 7115 1014 7149 1022
rect 7017 1002 7042 1014
rect 7049 1002 7068 1014
rect 7122 1012 7149 1014
rect 7158 1012 7379 1022
rect 7414 1019 7420 1022
rect 7122 1008 7379 1012
rect 7017 994 7068 1002
rect 7115 994 7379 1008
rect 7423 1014 7458 1022
rect 6969 946 6988 980
rect 7033 986 7062 994
rect 7033 980 7050 986
rect 7033 978 7067 980
rect 7115 978 7131 994
rect 7132 984 7340 994
rect 7341 984 7357 994
rect 7405 990 7420 1005
rect 7423 1002 7424 1014
rect 7431 1002 7458 1014
rect 7423 994 7458 1002
rect 7423 993 7452 994
rect 7143 980 7357 984
rect 7158 978 7357 980
rect 7392 980 7405 990
rect 7423 980 7440 993
rect 7392 978 7440 980
rect 7034 974 7067 978
rect 7030 972 7067 974
rect 7030 971 7097 972
rect 7030 966 7061 971
rect 7067 966 7097 971
rect 7030 962 7097 966
rect 7003 959 7097 962
rect 7003 952 7052 959
rect 7003 946 7033 952
rect 7052 947 7057 952
rect 6969 930 7049 946
rect 7061 938 7097 959
rect 7158 954 7347 978
rect 7392 977 7439 978
rect 7405 972 7439 977
rect 7173 951 7347 954
rect 7166 948 7347 951
rect 7375 971 7439 972
rect 6969 928 6988 930
rect 7003 928 7037 930
rect 6969 912 7049 928
rect 6969 906 6988 912
rect 6685 880 6788 890
rect 6639 878 6788 880
rect 6809 878 6844 890
rect 6478 876 6640 878
rect 6490 856 6509 876
rect 6524 874 6554 876
rect 6373 848 6414 856
rect 6496 852 6509 856
rect 6561 860 6640 876
rect 6672 876 6844 878
rect 6672 860 6751 876
rect 6758 874 6788 876
rect 6336 838 6365 848
rect 6379 838 6408 848
rect 6423 838 6453 852
rect 6496 838 6539 852
rect 6561 848 6751 860
rect 6816 856 6822 876
rect 6546 838 6576 848
rect 6577 838 6735 848
rect 6739 838 6769 848
rect 6773 838 6803 852
rect 6831 838 6844 876
rect 6916 890 6945 906
rect 6959 890 6988 906
rect 7003 896 7033 912
rect 7061 890 7067 938
rect 7070 932 7089 938
rect 7104 932 7134 940
rect 7070 924 7134 932
rect 7070 908 7150 924
rect 7166 917 7228 948
rect 7244 917 7306 948
rect 7375 946 7424 971
rect 7439 946 7469 962
rect 7338 932 7368 940
rect 7375 938 7485 946
rect 7338 924 7383 932
rect 7070 906 7089 908
rect 7104 906 7150 908
rect 7070 890 7150 906
rect 7177 904 7212 917
rect 7253 914 7290 917
rect 7253 912 7295 914
rect 7182 901 7212 904
rect 7191 897 7198 901
rect 7198 896 7199 897
rect 7157 890 7167 896
rect 6916 882 6951 890
rect 6916 856 6917 882
rect 6924 856 6951 882
rect 6859 838 6889 852
rect 6916 848 6951 856
rect 6953 882 6994 890
rect 6953 856 6968 882
rect 6975 856 6994 882
rect 7058 878 7089 890
rect 7104 878 7207 890
rect 7219 880 7245 906
rect 7260 901 7290 912
rect 7322 908 7384 924
rect 7322 906 7368 908
rect 7322 890 7384 906
rect 7396 890 7402 938
rect 7405 930 7485 938
rect 7405 928 7424 930
rect 7439 928 7473 930
rect 7405 912 7485 928
rect 7405 890 7424 912
rect 7439 896 7469 912
rect 7497 906 7503 980
rect 7506 906 7525 1050
rect 7540 906 7546 1050
rect 7555 980 7568 1050
rect 7620 1046 7642 1050
rect 7613 1024 7642 1038
rect 7695 1024 7711 1038
rect 7749 1034 7755 1036
rect 7762 1034 7870 1050
rect 7877 1034 7883 1036
rect 7891 1034 7906 1050
rect 7972 1044 7991 1047
rect 7613 1022 7711 1024
rect 7738 1022 7906 1034
rect 7921 1024 7937 1038
rect 7972 1025 7994 1044
rect 8004 1038 8020 1039
rect 8003 1036 8020 1038
rect 8004 1031 8020 1036
rect 7994 1024 8000 1025
rect 8003 1024 8032 1031
rect 7921 1023 8032 1024
rect 7921 1022 8038 1023
rect 7597 1014 7648 1022
rect 7695 1014 7729 1022
rect 7597 1002 7622 1014
rect 7629 1002 7648 1014
rect 7702 1012 7729 1014
rect 7738 1012 7959 1022
rect 7994 1019 8000 1022
rect 7702 1008 7959 1012
rect 7597 994 7648 1002
rect 7695 994 7959 1008
rect 8003 1014 8038 1022
rect 7549 946 7568 980
rect 7613 986 7642 994
rect 7613 980 7630 986
rect 7613 978 7647 980
rect 7695 978 7711 994
rect 7712 984 7920 994
rect 7921 984 7937 994
rect 7985 990 8000 1005
rect 8003 1002 8004 1014
rect 8011 1002 8038 1014
rect 8003 994 8038 1002
rect 8003 993 8032 994
rect 7723 980 7937 984
rect 7738 978 7937 980
rect 7972 980 7985 990
rect 8003 980 8020 993
rect 7972 978 8020 980
rect 7614 974 7647 978
rect 7610 972 7647 974
rect 7610 971 7677 972
rect 7610 966 7641 971
rect 7647 966 7677 971
rect 7610 962 7677 966
rect 7583 959 7677 962
rect 7583 952 7632 959
rect 7583 946 7613 952
rect 7632 947 7637 952
rect 7549 930 7629 946
rect 7641 938 7677 959
rect 7738 954 7927 978
rect 7972 977 8019 978
rect 7985 972 8019 977
rect 7753 951 7927 954
rect 7746 948 7927 951
rect 7955 971 8019 972
rect 7549 928 7568 930
rect 7583 928 7617 930
rect 7549 912 7629 928
rect 7549 906 7568 912
rect 7265 880 7368 890
rect 7219 878 7368 880
rect 7389 878 7424 890
rect 7058 876 7220 878
rect 7070 856 7089 876
rect 7104 874 7134 876
rect 6953 848 6994 856
rect 7076 852 7089 856
rect 7141 860 7220 876
rect 7252 876 7424 878
rect 7252 860 7331 876
rect 7338 874 7368 876
rect 6916 838 6945 848
rect 6959 838 6988 848
rect 7003 838 7033 852
rect 7076 838 7119 852
rect 7141 848 7331 860
rect 7396 856 7402 876
rect 7126 838 7156 848
rect 7157 838 7315 848
rect 7319 838 7349 848
rect 7353 838 7383 852
rect 7411 838 7424 876
rect 7496 890 7525 906
rect 7539 890 7568 906
rect 7583 896 7613 912
rect 7641 890 7647 938
rect 7650 932 7669 938
rect 7684 932 7714 940
rect 7650 924 7714 932
rect 7650 908 7730 924
rect 7746 917 7808 948
rect 7824 917 7886 948
rect 7955 946 8004 971
rect 8019 946 8049 962
rect 7918 932 7948 940
rect 7955 938 8065 946
rect 7918 924 7963 932
rect 7650 906 7669 908
rect 7684 906 7730 908
rect 7650 890 7730 906
rect 7757 904 7792 917
rect 7833 914 7870 917
rect 7833 912 7875 914
rect 7762 901 7792 904
rect 7771 897 7778 901
rect 7778 896 7779 897
rect 7737 890 7747 896
rect 7496 882 7531 890
rect 7496 856 7497 882
rect 7504 856 7531 882
rect 7439 838 7469 852
rect 7496 848 7531 856
rect 7533 882 7574 890
rect 7533 856 7548 882
rect 7555 856 7574 882
rect 7638 878 7669 890
rect 7684 878 7787 890
rect 7799 880 7825 906
rect 7840 901 7870 912
rect 7902 908 7964 924
rect 7902 906 7948 908
rect 7902 890 7964 906
rect 7976 890 7982 938
rect 7985 930 8065 938
rect 7985 928 8004 930
rect 8019 928 8053 930
rect 7985 912 8065 928
rect 7985 890 8004 912
rect 8019 896 8049 912
rect 8077 906 8083 980
rect 8086 906 8105 1050
rect 8120 906 8126 1050
rect 8135 980 8148 1050
rect 8200 1046 8222 1050
rect 8193 1024 8222 1038
rect 8275 1024 8291 1038
rect 8329 1034 8335 1036
rect 8342 1034 8450 1050
rect 8457 1034 8463 1036
rect 8471 1034 8486 1050
rect 8552 1044 8571 1047
rect 8193 1022 8291 1024
rect 8318 1022 8486 1034
rect 8501 1024 8517 1038
rect 8552 1025 8574 1044
rect 8584 1038 8600 1039
rect 8583 1036 8600 1038
rect 8584 1031 8600 1036
rect 8574 1024 8580 1025
rect 8583 1024 8612 1031
rect 8501 1023 8612 1024
rect 8501 1022 8618 1023
rect 8177 1014 8228 1022
rect 8275 1014 8309 1022
rect 8177 1002 8202 1014
rect 8209 1002 8228 1014
rect 8282 1012 8309 1014
rect 8318 1012 8539 1022
rect 8574 1019 8580 1022
rect 8282 1008 8539 1012
rect 8177 994 8228 1002
rect 8275 994 8539 1008
rect 8583 1014 8618 1022
rect 8129 946 8148 980
rect 8193 986 8222 994
rect 8193 980 8210 986
rect 8193 978 8227 980
rect 8275 978 8291 994
rect 8292 984 8500 994
rect 8501 984 8517 994
rect 8565 990 8580 1005
rect 8583 1002 8584 1014
rect 8591 1002 8618 1014
rect 8583 994 8618 1002
rect 8583 993 8612 994
rect 8303 980 8517 984
rect 8318 978 8517 980
rect 8552 980 8565 990
rect 8583 980 8600 993
rect 8552 978 8600 980
rect 8194 974 8227 978
rect 8190 972 8227 974
rect 8190 971 8257 972
rect 8190 966 8221 971
rect 8227 966 8257 971
rect 8190 962 8257 966
rect 8163 959 8257 962
rect 8163 952 8212 959
rect 8163 946 8193 952
rect 8212 947 8217 952
rect 8129 930 8209 946
rect 8221 938 8257 959
rect 8318 954 8507 978
rect 8552 977 8599 978
rect 8565 972 8599 977
rect 8333 951 8507 954
rect 8326 948 8507 951
rect 8535 971 8599 972
rect 8129 928 8148 930
rect 8163 928 8197 930
rect 8129 912 8209 928
rect 8129 906 8148 912
rect 7845 880 7948 890
rect 7799 878 7948 880
rect 7969 878 8004 890
rect 7638 876 7800 878
rect 7650 856 7669 876
rect 7684 874 7714 876
rect 7533 848 7574 856
rect 7656 852 7669 856
rect 7721 860 7800 876
rect 7832 876 8004 878
rect 7832 860 7911 876
rect 7918 874 7948 876
rect 7496 838 7525 848
rect 7539 838 7568 848
rect 7583 838 7613 852
rect 7656 838 7699 852
rect 7721 848 7911 860
rect 7976 856 7982 876
rect 7706 838 7736 848
rect 7737 838 7895 848
rect 7899 838 7929 848
rect 7933 838 7963 852
rect 7991 838 8004 876
rect 8076 890 8105 906
rect 8119 890 8148 906
rect 8163 896 8193 912
rect 8221 890 8227 938
rect 8230 932 8249 938
rect 8264 932 8294 940
rect 8230 924 8294 932
rect 8230 908 8310 924
rect 8326 917 8388 948
rect 8404 917 8466 948
rect 8535 946 8584 971
rect 8599 946 8629 962
rect 8498 932 8528 940
rect 8535 938 8645 946
rect 8498 924 8543 932
rect 8230 906 8249 908
rect 8264 906 8310 908
rect 8230 890 8310 906
rect 8337 904 8372 917
rect 8413 914 8450 917
rect 8413 912 8455 914
rect 8342 901 8372 904
rect 8351 897 8358 901
rect 8358 896 8359 897
rect 8317 890 8327 896
rect 8076 882 8111 890
rect 8076 856 8077 882
rect 8084 856 8111 882
rect 8019 838 8049 852
rect 8076 848 8111 856
rect 8113 882 8154 890
rect 8113 856 8128 882
rect 8135 856 8154 882
rect 8218 878 8249 890
rect 8264 878 8367 890
rect 8379 880 8405 906
rect 8420 901 8450 912
rect 8482 908 8544 924
rect 8482 906 8528 908
rect 8482 890 8544 906
rect 8556 890 8562 938
rect 8565 930 8645 938
rect 8565 928 8584 930
rect 8599 928 8633 930
rect 8565 912 8645 928
rect 8565 890 8584 912
rect 8599 896 8629 912
rect 8657 906 8663 980
rect 8666 906 8685 1050
rect 8700 906 8706 1050
rect 8715 980 8728 1050
rect 8780 1046 8802 1050
rect 8773 1024 8802 1038
rect 8855 1024 8871 1038
rect 8909 1034 8915 1036
rect 8922 1034 9030 1050
rect 9037 1034 9043 1036
rect 9051 1034 9066 1050
rect 9132 1044 9151 1047
rect 8773 1022 8871 1024
rect 8898 1022 9066 1034
rect 9081 1024 9097 1038
rect 9132 1025 9154 1044
rect 9164 1038 9180 1039
rect 9163 1036 9180 1038
rect 9164 1031 9180 1036
rect 9154 1024 9160 1025
rect 9163 1024 9192 1031
rect 9081 1023 9192 1024
rect 9081 1022 9198 1023
rect 8757 1014 8808 1022
rect 8855 1014 8889 1022
rect 8757 1002 8782 1014
rect 8789 1002 8808 1014
rect 8862 1012 8889 1014
rect 8898 1012 9119 1022
rect 9154 1019 9160 1022
rect 8862 1008 9119 1012
rect 8757 994 8808 1002
rect 8855 994 9119 1008
rect 9163 1014 9198 1022
rect 8709 946 8728 980
rect 8773 986 8802 994
rect 8773 980 8790 986
rect 8773 978 8807 980
rect 8855 978 8871 994
rect 8872 984 9080 994
rect 9081 984 9097 994
rect 9145 990 9160 1005
rect 9163 1002 9164 1014
rect 9171 1002 9198 1014
rect 9163 994 9198 1002
rect 9163 993 9192 994
rect 8883 980 9097 984
rect 8898 978 9097 980
rect 9132 980 9145 990
rect 9163 980 9180 993
rect 9132 978 9180 980
rect 8774 974 8807 978
rect 8770 972 8807 974
rect 8770 971 8837 972
rect 8770 966 8801 971
rect 8807 966 8837 971
rect 8770 962 8837 966
rect 8743 959 8837 962
rect 8743 952 8792 959
rect 8743 946 8773 952
rect 8792 947 8797 952
rect 8709 930 8789 946
rect 8801 938 8837 959
rect 8898 954 9087 978
rect 9132 977 9179 978
rect 9145 972 9179 977
rect 8913 951 9087 954
rect 8906 948 9087 951
rect 9115 971 9179 972
rect 8709 928 8728 930
rect 8743 928 8777 930
rect 8709 912 8789 928
rect 8709 906 8728 912
rect 8425 880 8528 890
rect 8379 878 8528 880
rect 8549 878 8584 890
rect 8218 876 8380 878
rect 8230 856 8249 876
rect 8264 874 8294 876
rect 8113 848 8154 856
rect 8236 852 8249 856
rect 8301 860 8380 876
rect 8412 876 8584 878
rect 8412 860 8491 876
rect 8498 874 8528 876
rect 8076 838 8105 848
rect 8119 838 8148 848
rect 8163 838 8193 852
rect 8236 838 8279 852
rect 8301 848 8491 860
rect 8556 856 8562 876
rect 8286 838 8316 848
rect 8317 838 8475 848
rect 8479 838 8509 848
rect 8513 838 8543 852
rect 8571 838 8584 876
rect 8656 890 8685 906
rect 8699 890 8728 906
rect 8743 896 8773 912
rect 8801 890 8807 938
rect 8810 932 8829 938
rect 8844 932 8874 940
rect 8810 924 8874 932
rect 8810 908 8890 924
rect 8906 917 8968 948
rect 8984 917 9046 948
rect 9115 946 9164 971
rect 9179 946 9209 962
rect 9078 932 9108 940
rect 9115 938 9225 946
rect 9078 924 9123 932
rect 8810 906 8829 908
rect 8844 906 8890 908
rect 8810 890 8890 906
rect 8917 904 8952 917
rect 8993 914 9030 917
rect 8993 912 9035 914
rect 8922 901 8952 904
rect 8931 897 8938 901
rect 8938 896 8939 897
rect 8897 890 8907 896
rect 8656 882 8691 890
rect 8656 856 8657 882
rect 8664 856 8691 882
rect 8599 838 8629 852
rect 8656 848 8691 856
rect 8693 882 8734 890
rect 8693 856 8708 882
rect 8715 856 8734 882
rect 8798 878 8829 890
rect 8844 878 8947 890
rect 8959 880 8985 906
rect 9000 901 9030 912
rect 9062 908 9124 924
rect 9062 906 9108 908
rect 9062 890 9124 906
rect 9136 890 9142 938
rect 9145 930 9225 938
rect 9145 928 9164 930
rect 9179 928 9213 930
rect 9145 912 9225 928
rect 9145 890 9164 912
rect 9179 896 9209 912
rect 9237 906 9243 980
rect 9252 906 9265 1050
rect 9005 880 9108 890
rect 8959 878 9108 880
rect 9129 878 9164 890
rect 8798 876 8960 878
rect 8810 856 8829 876
rect 8844 874 8874 876
rect 8693 848 8734 856
rect 8816 852 8829 856
rect 8881 860 8960 876
rect 8992 876 9164 878
rect 8992 860 9071 876
rect 9078 874 9108 876
rect 8656 838 8685 848
rect 8699 838 8728 848
rect 8743 838 8773 852
rect 8816 838 8859 852
rect 8881 848 9071 860
rect 9136 856 9142 876
rect 8866 838 8896 848
rect 8897 838 9055 848
rect 9059 838 9089 848
rect 9093 838 9123 852
rect 9151 838 9164 876
rect 9236 890 9265 906
rect 9236 882 9271 890
rect 9236 856 9237 882
rect 9244 856 9271 882
rect 9179 838 9209 852
rect 9236 848 9271 856
rect 9236 838 9265 848
rect -1 832 9265 838
rect 0 824 9265 832
rect 15 794 28 824
rect 43 810 73 824
rect 116 810 159 824
rect 166 810 386 824
rect 393 810 423 824
rect 83 796 98 808
rect 117 796 130 810
rect 198 806 351 810
rect 80 794 102 796
rect 180 794 372 806
rect 451 794 464 824
rect 479 810 509 824
rect 546 794 565 824
rect 580 794 586 824
rect 595 794 608 824
rect 623 810 653 824
rect 696 810 739 824
rect 746 810 966 824
rect 973 810 1003 824
rect 663 796 678 808
rect 697 796 710 810
rect 778 806 931 810
rect 660 794 682 796
rect 760 794 952 806
rect 1031 794 1044 824
rect 1059 810 1089 824
rect 1126 794 1145 824
rect 1160 794 1166 824
rect 1175 794 1188 824
rect 1203 810 1233 824
rect 1276 810 1319 824
rect 1326 810 1546 824
rect 1553 810 1583 824
rect 1243 796 1258 808
rect 1277 796 1290 810
rect 1358 806 1511 810
rect 1240 794 1262 796
rect 1340 794 1532 806
rect 1611 794 1624 824
rect 1639 810 1669 824
rect 1706 794 1725 824
rect 1740 794 1746 824
rect 1755 794 1768 824
rect 1783 810 1813 824
rect 1856 810 1899 824
rect 1906 810 2126 824
rect 2133 810 2163 824
rect 1823 796 1838 808
rect 1857 796 1870 810
rect 1938 806 2091 810
rect 1820 794 1842 796
rect 1920 794 2112 806
rect 2191 794 2204 824
rect 2219 810 2249 824
rect 2286 794 2305 824
rect 2320 794 2326 824
rect 2335 794 2348 824
rect 2363 810 2393 824
rect 2436 810 2479 824
rect 2486 810 2706 824
rect 2713 810 2743 824
rect 2403 796 2418 808
rect 2437 796 2450 810
rect 2518 806 2671 810
rect 2400 794 2422 796
rect 2500 794 2692 806
rect 2771 794 2784 824
rect 2799 810 2829 824
rect 2866 794 2885 824
rect 2900 794 2906 824
rect 2915 794 2928 824
rect 2943 810 2973 824
rect 3016 810 3059 824
rect 3066 810 3286 824
rect 3293 810 3323 824
rect 2983 796 2998 808
rect 3017 796 3030 810
rect 3098 806 3251 810
rect 2980 794 3002 796
rect 3080 794 3272 806
rect 3351 794 3364 824
rect 3379 810 3409 824
rect 3446 794 3465 824
rect 3480 794 3486 824
rect 3495 794 3508 824
rect 3523 810 3553 824
rect 3596 810 3639 824
rect 3646 810 3866 824
rect 3873 810 3903 824
rect 3563 796 3578 808
rect 3597 796 3610 810
rect 3678 806 3831 810
rect 3560 794 3582 796
rect 3660 794 3852 806
rect 3931 794 3944 824
rect 3959 810 3989 824
rect 4026 794 4045 824
rect 4060 794 4066 824
rect 4075 794 4088 824
rect 4103 810 4133 824
rect 4176 810 4219 824
rect 4226 810 4446 824
rect 4453 810 4483 824
rect 4143 796 4158 808
rect 4177 796 4190 810
rect 4258 806 4411 810
rect 4140 794 4162 796
rect 4240 794 4432 806
rect 4511 794 4524 824
rect 4539 810 4569 824
rect 4606 794 4625 824
rect 4640 794 4646 824
rect 4655 794 4668 824
rect 4683 810 4713 824
rect 4756 810 4799 824
rect 4806 810 5026 824
rect 5033 810 5063 824
rect 4723 796 4738 808
rect 4757 796 4770 810
rect 4838 806 4991 810
rect 4720 794 4742 796
rect 4820 794 5012 806
rect 5091 794 5104 824
rect 5119 810 5149 824
rect 5186 794 5205 824
rect 5220 794 5226 824
rect 5235 794 5248 824
rect 5263 810 5293 824
rect 5336 810 5379 824
rect 5386 810 5606 824
rect 5613 810 5643 824
rect 5303 796 5318 808
rect 5337 796 5350 810
rect 5418 806 5571 810
rect 5300 794 5322 796
rect 5400 794 5592 806
rect 5671 794 5684 824
rect 5699 810 5729 824
rect 5766 794 5785 824
rect 5800 794 5806 824
rect 5815 794 5828 824
rect 5843 810 5873 824
rect 5916 810 5959 824
rect 5966 810 6186 824
rect 6193 810 6223 824
rect 5883 796 5898 808
rect 5917 796 5930 810
rect 5998 806 6151 810
rect 5880 794 5902 796
rect 5980 794 6172 806
rect 6251 794 6264 824
rect 6279 810 6309 824
rect 6346 794 6365 824
rect 6380 794 6386 824
rect 6395 794 6408 824
rect 6423 810 6453 824
rect 6496 810 6539 824
rect 6546 810 6766 824
rect 6773 810 6803 824
rect 6463 796 6478 808
rect 6497 796 6510 810
rect 6578 806 6731 810
rect 6460 794 6482 796
rect 6560 794 6752 806
rect 6831 794 6844 824
rect 6859 810 6889 824
rect 6926 794 6945 824
rect 6960 794 6966 824
rect 6975 794 6988 824
rect 7003 810 7033 824
rect 7076 810 7119 824
rect 7126 810 7346 824
rect 7353 810 7383 824
rect 7043 796 7058 808
rect 7077 796 7090 810
rect 7158 806 7311 810
rect 7040 794 7062 796
rect 7140 794 7332 806
rect 7411 794 7424 824
rect 7439 810 7469 824
rect 7506 794 7525 824
rect 7540 794 7546 824
rect 7555 794 7568 824
rect 7583 810 7613 824
rect 7656 810 7699 824
rect 7706 810 7926 824
rect 7933 810 7963 824
rect 7623 796 7638 808
rect 7657 796 7670 810
rect 7738 806 7891 810
rect 7620 794 7642 796
rect 7720 794 7912 806
rect 7991 794 8004 824
rect 8019 810 8049 824
rect 8086 794 8105 824
rect 8120 794 8126 824
rect 8135 794 8148 824
rect 8163 810 8193 824
rect 8236 810 8279 824
rect 8286 810 8506 824
rect 8513 810 8543 824
rect 8203 796 8218 808
rect 8237 796 8250 810
rect 8318 806 8471 810
rect 8200 794 8222 796
rect 8300 794 8492 806
rect 8571 794 8584 824
rect 8599 810 8629 824
rect 8666 794 8685 824
rect 8700 794 8706 824
rect 8715 794 8728 824
rect 8743 810 8773 824
rect 8816 810 8859 824
rect 8866 810 9086 824
rect 9093 810 9123 824
rect 8783 796 8798 808
rect 8817 796 8830 810
rect 8898 806 9051 810
rect 8780 794 8802 796
rect 8880 794 9072 806
rect 9151 794 9164 824
rect 9179 810 9209 824
rect 9252 794 9265 824
rect 0 780 9265 794
rect 15 710 28 780
rect 80 776 102 780
rect 73 754 102 768
rect 155 754 171 768
rect 209 765 215 766
rect 222 765 330 780
rect 337 765 343 766
rect 351 765 366 780
rect 432 774 451 777
rect 73 752 171 754
rect 198 752 366 765
rect 381 754 397 768
rect 432 755 454 774
rect 464 768 480 769
rect 463 766 480 768
rect 464 761 480 766
rect 454 754 460 755
rect 463 754 492 761
rect 381 753 492 754
rect 381 752 498 753
rect 57 744 108 752
rect 155 744 189 752
rect 57 732 82 744
rect 89 732 108 744
rect 162 742 189 744
rect 198 742 419 752
rect 454 749 460 752
rect 162 738 419 742
rect 57 724 108 732
rect 155 724 419 738
rect 463 744 498 752
rect 9 676 28 710
rect 73 716 102 724
rect 73 710 90 716
rect 73 708 107 710
rect 155 708 171 724
rect 172 714 380 724
rect 381 714 397 724
rect 445 720 460 735
rect 463 732 464 744
rect 471 732 498 744
rect 463 724 498 732
rect 463 723 492 724
rect 183 710 397 714
rect 198 708 397 710
rect 432 710 445 720
rect 463 710 480 723
rect 432 708 480 710
rect 74 704 107 708
rect 70 702 107 704
rect 70 701 137 702
rect 70 696 101 701
rect 107 696 137 701
rect 70 692 137 696
rect 43 689 137 692
rect 43 682 92 689
rect 43 676 73 682
rect 92 677 97 682
rect 9 660 89 676
rect 101 668 137 689
rect 198 684 387 708
rect 432 707 479 708
rect 445 702 479 707
rect 213 681 387 684
rect 206 678 387 681
rect 415 701 479 702
rect 9 658 28 660
rect 43 658 77 660
rect 9 642 89 658
rect 9 636 28 642
rect -1 620 28 636
rect 43 626 73 642
rect 101 620 107 668
rect 110 662 129 668
rect 144 662 174 670
rect 110 654 174 662
rect 110 638 190 654
rect 206 647 268 678
rect 284 647 346 678
rect 415 676 464 701
rect 479 676 509 692
rect 378 662 408 670
rect 415 668 525 676
rect 378 654 423 662
rect 110 636 129 638
rect 144 636 190 638
rect 110 620 190 636
rect 217 634 252 647
rect 293 644 330 647
rect 293 642 335 644
rect 222 631 252 634
rect 231 627 238 631
rect 238 626 239 627
rect 197 620 207 626
rect -7 612 34 620
rect -7 586 8 612
rect 15 586 34 612
rect 98 608 129 620
rect 144 608 247 620
rect 259 610 285 636
rect 300 631 330 642
rect 362 638 424 654
rect 362 636 408 638
rect 362 620 424 636
rect 436 620 442 668
rect 445 660 525 668
rect 445 658 464 660
rect 479 658 513 660
rect 445 642 525 658
rect 445 620 464 642
rect 479 626 509 642
rect 537 636 543 710
rect 546 636 565 780
rect 580 636 586 780
rect 595 710 608 780
rect 660 776 682 780
rect 653 754 682 768
rect 735 754 751 768
rect 789 765 795 766
rect 802 765 910 780
rect 917 765 923 766
rect 931 765 946 780
rect 1012 774 1031 777
rect 653 752 751 754
rect 778 752 946 765
rect 961 754 977 768
rect 1012 755 1034 774
rect 1044 768 1060 769
rect 1043 766 1060 768
rect 1044 761 1060 766
rect 1034 754 1040 755
rect 1043 754 1072 761
rect 961 753 1072 754
rect 961 752 1078 753
rect 637 744 688 752
rect 735 744 769 752
rect 637 732 662 744
rect 669 732 688 744
rect 742 742 769 744
rect 778 742 999 752
rect 1034 749 1040 752
rect 742 738 999 742
rect 637 724 688 732
rect 735 724 999 738
rect 1043 744 1078 752
rect 589 676 608 710
rect 653 716 682 724
rect 653 710 670 716
rect 653 708 687 710
rect 735 708 751 724
rect 752 714 960 724
rect 961 714 977 724
rect 1025 720 1040 735
rect 1043 732 1044 744
rect 1051 732 1078 744
rect 1043 724 1078 732
rect 1043 723 1072 724
rect 763 710 977 714
rect 778 708 977 710
rect 1012 710 1025 720
rect 1043 710 1060 723
rect 1012 708 1060 710
rect 654 704 687 708
rect 650 702 687 704
rect 650 701 717 702
rect 650 696 681 701
rect 687 696 717 701
rect 650 692 717 696
rect 623 689 717 692
rect 623 682 672 689
rect 623 676 653 682
rect 672 677 677 682
rect 589 660 669 676
rect 681 668 717 689
rect 778 684 967 708
rect 1012 707 1059 708
rect 1025 702 1059 707
rect 793 681 967 684
rect 786 678 967 681
rect 995 701 1059 702
rect 589 658 608 660
rect 623 658 657 660
rect 589 642 669 658
rect 589 636 608 642
rect 305 610 408 620
rect 259 608 408 610
rect 429 608 464 620
rect 98 606 260 608
rect 110 586 129 606
rect 144 604 174 606
rect -7 578 34 586
rect 116 583 129 586
rect 181 590 260 606
rect 292 606 464 608
rect 292 590 371 606
rect 378 604 408 606
rect -1 568 28 578
rect 43 568 73 583
rect 116 579 159 583
rect 181 579 371 590
rect 436 586 442 606
rect 393 579 423 583
rect 116 578 423 579
rect 116 568 159 578
rect 166 568 196 578
rect 197 568 355 578
rect 359 568 389 578
rect 393 568 423 578
rect 451 568 464 606
rect 536 620 565 636
rect 579 620 608 636
rect 623 626 653 642
rect 681 620 687 668
rect 690 662 709 668
rect 724 662 754 670
rect 690 654 754 662
rect 690 638 770 654
rect 786 647 848 678
rect 864 647 926 678
rect 995 676 1044 701
rect 1059 676 1089 692
rect 958 662 988 670
rect 995 668 1105 676
rect 958 654 1003 662
rect 690 636 709 638
rect 724 636 770 638
rect 690 620 770 636
rect 797 634 832 647
rect 873 644 910 647
rect 873 642 915 644
rect 802 631 832 634
rect 811 627 818 631
rect 818 626 819 627
rect 777 620 787 626
rect 536 612 571 620
rect 536 586 537 612
rect 544 586 571 612
rect 479 568 509 583
rect 536 578 571 586
rect 573 612 614 620
rect 573 586 588 612
rect 595 586 614 612
rect 678 608 709 620
rect 724 608 827 620
rect 839 610 865 636
rect 880 631 910 642
rect 942 638 1004 654
rect 942 636 988 638
rect 942 620 1004 636
rect 1016 620 1022 668
rect 1025 660 1105 668
rect 1025 658 1044 660
rect 1059 658 1093 660
rect 1025 642 1105 658
rect 1025 620 1044 642
rect 1059 626 1089 642
rect 1117 636 1123 710
rect 1126 636 1145 780
rect 1160 636 1166 780
rect 1175 710 1188 780
rect 1240 776 1262 780
rect 1233 754 1262 768
rect 1315 754 1331 768
rect 1369 765 1375 766
rect 1382 765 1490 780
rect 1497 765 1503 766
rect 1511 765 1526 780
rect 1592 774 1611 777
rect 1233 752 1331 754
rect 1358 752 1526 765
rect 1541 754 1557 768
rect 1592 755 1614 774
rect 1624 768 1640 769
rect 1623 766 1640 768
rect 1624 761 1640 766
rect 1614 754 1620 755
rect 1623 754 1652 761
rect 1541 753 1652 754
rect 1541 752 1658 753
rect 1217 744 1268 752
rect 1315 744 1349 752
rect 1217 732 1242 744
rect 1249 732 1268 744
rect 1322 742 1349 744
rect 1358 742 1579 752
rect 1614 749 1620 752
rect 1322 738 1579 742
rect 1217 724 1268 732
rect 1315 724 1579 738
rect 1623 744 1658 752
rect 1169 676 1188 710
rect 1233 716 1262 724
rect 1233 710 1250 716
rect 1233 708 1267 710
rect 1315 708 1331 724
rect 1332 714 1540 724
rect 1541 714 1557 724
rect 1605 720 1620 735
rect 1623 732 1624 744
rect 1631 732 1658 744
rect 1623 724 1658 732
rect 1623 723 1652 724
rect 1343 710 1557 714
rect 1358 708 1557 710
rect 1592 710 1605 720
rect 1623 710 1640 723
rect 1592 708 1640 710
rect 1234 704 1267 708
rect 1230 702 1267 704
rect 1230 701 1297 702
rect 1230 696 1261 701
rect 1267 696 1297 701
rect 1230 692 1297 696
rect 1203 689 1297 692
rect 1203 682 1252 689
rect 1203 676 1233 682
rect 1252 677 1257 682
rect 1169 660 1249 676
rect 1261 668 1297 689
rect 1358 684 1547 708
rect 1592 707 1639 708
rect 1605 702 1639 707
rect 1373 681 1547 684
rect 1366 678 1547 681
rect 1575 701 1639 702
rect 1169 658 1188 660
rect 1203 658 1237 660
rect 1169 642 1249 658
rect 1169 636 1188 642
rect 885 610 988 620
rect 839 608 988 610
rect 1009 608 1044 620
rect 678 606 840 608
rect 690 586 709 606
rect 724 604 754 606
rect 573 578 614 586
rect 696 583 709 586
rect 761 590 840 606
rect 872 606 1044 608
rect 872 590 951 606
rect 958 604 988 606
rect 536 568 565 578
rect 579 568 608 578
rect 623 568 653 583
rect 696 579 739 583
rect 761 579 951 590
rect 1016 586 1022 606
rect 973 579 1003 583
rect 696 578 1003 579
rect 696 568 739 578
rect 746 568 776 578
rect 777 568 935 578
rect 939 568 969 578
rect 973 568 1003 578
rect 1031 568 1044 606
rect 1116 620 1145 636
rect 1159 620 1188 636
rect 1203 626 1233 642
rect 1261 620 1267 668
rect 1270 662 1289 668
rect 1304 662 1334 670
rect 1270 654 1334 662
rect 1270 638 1350 654
rect 1366 647 1428 678
rect 1444 647 1506 678
rect 1575 676 1624 701
rect 1639 676 1669 692
rect 1538 662 1568 670
rect 1575 668 1685 676
rect 1538 654 1583 662
rect 1270 636 1289 638
rect 1304 636 1350 638
rect 1270 620 1350 636
rect 1377 634 1412 647
rect 1453 644 1490 647
rect 1453 642 1495 644
rect 1382 631 1412 634
rect 1391 627 1398 631
rect 1398 626 1399 627
rect 1357 620 1367 626
rect 1116 612 1151 620
rect 1116 586 1117 612
rect 1124 586 1151 612
rect 1059 568 1089 583
rect 1116 578 1151 586
rect 1153 612 1194 620
rect 1153 586 1168 612
rect 1175 586 1194 612
rect 1258 608 1289 620
rect 1304 608 1407 620
rect 1419 610 1445 636
rect 1460 631 1490 642
rect 1522 638 1584 654
rect 1522 636 1568 638
rect 1522 620 1584 636
rect 1596 620 1602 668
rect 1605 660 1685 668
rect 1605 658 1624 660
rect 1639 658 1673 660
rect 1605 642 1685 658
rect 1605 620 1624 642
rect 1639 626 1669 642
rect 1697 636 1703 710
rect 1706 636 1725 780
rect 1740 636 1746 780
rect 1755 710 1768 780
rect 1820 776 1842 780
rect 1813 754 1842 768
rect 1895 754 1911 768
rect 1949 765 1955 766
rect 1962 765 2070 780
rect 2077 765 2083 766
rect 2091 765 2106 780
rect 2172 774 2191 777
rect 1813 752 1911 754
rect 1938 752 2106 765
rect 2121 754 2137 768
rect 2172 755 2194 774
rect 2204 768 2220 769
rect 2203 766 2220 768
rect 2204 761 2220 766
rect 2194 754 2200 755
rect 2203 754 2232 761
rect 2121 753 2232 754
rect 2121 752 2238 753
rect 1797 744 1848 752
rect 1895 744 1929 752
rect 1797 732 1822 744
rect 1829 732 1848 744
rect 1902 742 1929 744
rect 1938 742 2159 752
rect 2194 749 2200 752
rect 1902 738 2159 742
rect 1797 724 1848 732
rect 1895 724 2159 738
rect 2203 744 2238 752
rect 1749 676 1768 710
rect 1813 716 1842 724
rect 1813 710 1830 716
rect 1813 708 1847 710
rect 1895 708 1911 724
rect 1912 714 2120 724
rect 2121 714 2137 724
rect 2185 720 2200 735
rect 2203 732 2204 744
rect 2211 732 2238 744
rect 2203 724 2238 732
rect 2203 723 2232 724
rect 1923 710 2137 714
rect 1938 708 2137 710
rect 2172 710 2185 720
rect 2203 710 2220 723
rect 2172 708 2220 710
rect 1814 704 1847 708
rect 1810 702 1847 704
rect 1810 701 1877 702
rect 1810 696 1841 701
rect 1847 696 1877 701
rect 1810 692 1877 696
rect 1783 689 1877 692
rect 1783 682 1832 689
rect 1783 676 1813 682
rect 1832 677 1837 682
rect 1749 660 1829 676
rect 1841 668 1877 689
rect 1938 684 2127 708
rect 2172 707 2219 708
rect 2185 702 2219 707
rect 1953 681 2127 684
rect 1946 678 2127 681
rect 2155 701 2219 702
rect 1749 658 1768 660
rect 1783 658 1817 660
rect 1749 642 1829 658
rect 1749 636 1768 642
rect 1465 610 1568 620
rect 1419 608 1568 610
rect 1589 608 1624 620
rect 1258 606 1420 608
rect 1270 586 1289 606
rect 1304 604 1334 606
rect 1153 578 1194 586
rect 1276 583 1289 586
rect 1341 590 1420 606
rect 1452 606 1624 608
rect 1452 590 1531 606
rect 1538 604 1568 606
rect 1116 568 1145 578
rect 1159 568 1188 578
rect 1203 568 1233 583
rect 1276 579 1319 583
rect 1341 579 1531 590
rect 1596 586 1602 606
rect 1553 579 1583 583
rect 1276 578 1583 579
rect 1276 568 1319 578
rect 1326 568 1356 578
rect 1357 568 1515 578
rect 1519 568 1549 578
rect 1553 568 1583 578
rect 1611 568 1624 606
rect 1696 620 1725 636
rect 1739 620 1768 636
rect 1783 626 1813 642
rect 1841 620 1847 668
rect 1850 662 1869 668
rect 1884 662 1914 670
rect 1850 654 1914 662
rect 1850 638 1930 654
rect 1946 647 2008 678
rect 2024 647 2086 678
rect 2155 676 2204 701
rect 2219 676 2249 692
rect 2118 662 2148 670
rect 2155 668 2265 676
rect 2118 654 2163 662
rect 1850 636 1869 638
rect 1884 636 1930 638
rect 1850 620 1930 636
rect 1957 634 1992 647
rect 2033 644 2070 647
rect 2033 642 2075 644
rect 1962 631 1992 634
rect 1971 627 1978 631
rect 1978 626 1979 627
rect 1937 620 1947 626
rect 1696 612 1731 620
rect 1696 586 1697 612
rect 1704 586 1731 612
rect 1639 568 1669 583
rect 1696 578 1731 586
rect 1733 612 1774 620
rect 1733 586 1748 612
rect 1755 586 1774 612
rect 1838 608 1869 620
rect 1884 608 1987 620
rect 1999 610 2025 636
rect 2040 631 2070 642
rect 2102 638 2164 654
rect 2102 636 2148 638
rect 2102 620 2164 636
rect 2176 620 2182 668
rect 2185 660 2265 668
rect 2185 658 2204 660
rect 2219 658 2253 660
rect 2185 642 2265 658
rect 2185 620 2204 642
rect 2219 626 2249 642
rect 2277 636 2283 710
rect 2286 636 2305 780
rect 2320 636 2326 780
rect 2335 710 2348 780
rect 2400 776 2422 780
rect 2393 754 2422 768
rect 2475 754 2491 768
rect 2529 765 2535 766
rect 2542 765 2650 780
rect 2657 765 2663 766
rect 2671 765 2686 780
rect 2752 774 2771 777
rect 2393 752 2491 754
rect 2518 752 2686 765
rect 2701 754 2717 768
rect 2752 755 2774 774
rect 2784 768 2800 769
rect 2783 766 2800 768
rect 2784 761 2800 766
rect 2774 754 2780 755
rect 2783 754 2812 761
rect 2701 753 2812 754
rect 2701 752 2818 753
rect 2377 744 2428 752
rect 2475 744 2509 752
rect 2377 732 2402 744
rect 2409 732 2428 744
rect 2482 742 2509 744
rect 2518 742 2739 752
rect 2774 749 2780 752
rect 2482 738 2739 742
rect 2377 724 2428 732
rect 2475 724 2739 738
rect 2783 744 2818 752
rect 2329 676 2348 710
rect 2393 716 2422 724
rect 2393 710 2410 716
rect 2393 708 2427 710
rect 2475 708 2491 724
rect 2492 714 2700 724
rect 2701 714 2717 724
rect 2765 720 2780 735
rect 2783 732 2784 744
rect 2791 732 2818 744
rect 2783 724 2818 732
rect 2783 723 2812 724
rect 2503 710 2717 714
rect 2518 708 2717 710
rect 2752 710 2765 720
rect 2783 710 2800 723
rect 2752 708 2800 710
rect 2394 704 2427 708
rect 2390 702 2427 704
rect 2390 701 2457 702
rect 2390 696 2421 701
rect 2427 696 2457 701
rect 2390 692 2457 696
rect 2363 689 2457 692
rect 2363 682 2412 689
rect 2363 676 2393 682
rect 2412 677 2417 682
rect 2329 660 2409 676
rect 2421 668 2457 689
rect 2518 684 2707 708
rect 2752 707 2799 708
rect 2765 702 2799 707
rect 2533 681 2707 684
rect 2526 678 2707 681
rect 2735 701 2799 702
rect 2329 658 2348 660
rect 2363 658 2397 660
rect 2329 642 2409 658
rect 2329 636 2348 642
rect 2045 610 2148 620
rect 1999 608 2148 610
rect 2169 608 2204 620
rect 1838 606 2000 608
rect 1850 586 1869 606
rect 1884 604 1914 606
rect 1733 578 1774 586
rect 1856 583 1869 586
rect 1921 590 2000 606
rect 2032 606 2204 608
rect 2032 590 2111 606
rect 2118 604 2148 606
rect 1696 568 1725 578
rect 1739 568 1768 578
rect 1783 568 1813 583
rect 1856 579 1899 583
rect 1921 579 2111 590
rect 2176 586 2182 606
rect 2133 579 2163 583
rect 1856 578 2163 579
rect 1856 568 1899 578
rect 1906 568 1936 578
rect 1937 568 2095 578
rect 2099 568 2129 578
rect 2133 568 2163 578
rect 2191 568 2204 606
rect 2276 620 2305 636
rect 2319 620 2348 636
rect 2363 626 2393 642
rect 2421 620 2427 668
rect 2430 662 2449 668
rect 2464 662 2494 670
rect 2430 654 2494 662
rect 2430 638 2510 654
rect 2526 647 2588 678
rect 2604 647 2666 678
rect 2735 676 2784 701
rect 2799 676 2829 692
rect 2698 662 2728 670
rect 2735 668 2845 676
rect 2698 654 2743 662
rect 2430 636 2449 638
rect 2464 636 2510 638
rect 2430 620 2510 636
rect 2537 634 2572 647
rect 2613 644 2650 647
rect 2613 642 2655 644
rect 2542 631 2572 634
rect 2551 627 2558 631
rect 2558 626 2559 627
rect 2517 620 2527 626
rect 2276 612 2311 620
rect 2276 586 2277 612
rect 2284 586 2311 612
rect 2219 568 2249 583
rect 2276 578 2311 586
rect 2313 612 2354 620
rect 2313 586 2328 612
rect 2335 586 2354 612
rect 2418 608 2449 620
rect 2464 608 2567 620
rect 2579 610 2605 636
rect 2620 631 2650 642
rect 2682 638 2744 654
rect 2682 636 2728 638
rect 2682 620 2744 636
rect 2756 620 2762 668
rect 2765 660 2845 668
rect 2765 658 2784 660
rect 2799 658 2833 660
rect 2765 642 2845 658
rect 2765 620 2784 642
rect 2799 626 2829 642
rect 2857 636 2863 710
rect 2866 636 2885 780
rect 2900 636 2906 780
rect 2915 710 2928 780
rect 2980 776 3002 780
rect 2973 754 3002 768
rect 3055 754 3071 768
rect 3109 765 3115 766
rect 3122 765 3230 780
rect 3237 765 3243 766
rect 3251 765 3266 780
rect 3332 774 3351 777
rect 2973 752 3071 754
rect 3098 752 3266 765
rect 3281 754 3297 768
rect 3332 755 3354 774
rect 3364 768 3380 769
rect 3363 766 3380 768
rect 3364 761 3380 766
rect 3354 754 3360 755
rect 3363 754 3392 761
rect 3281 753 3392 754
rect 3281 752 3398 753
rect 2957 744 3008 752
rect 3055 744 3089 752
rect 2957 732 2982 744
rect 2989 732 3008 744
rect 3062 742 3089 744
rect 3098 742 3319 752
rect 3354 749 3360 752
rect 3062 738 3319 742
rect 2957 724 3008 732
rect 3055 724 3319 738
rect 3363 744 3398 752
rect 2909 676 2928 710
rect 2973 716 3002 724
rect 2973 710 2990 716
rect 2973 708 3007 710
rect 3055 708 3071 724
rect 3072 714 3280 724
rect 3281 714 3297 724
rect 3345 720 3360 735
rect 3363 732 3364 744
rect 3371 732 3398 744
rect 3363 724 3398 732
rect 3363 723 3392 724
rect 3083 710 3297 714
rect 3098 708 3297 710
rect 3332 710 3345 720
rect 3363 710 3380 723
rect 3332 708 3380 710
rect 2974 704 3007 708
rect 2970 702 3007 704
rect 2970 701 3037 702
rect 2970 696 3001 701
rect 3007 696 3037 701
rect 2970 692 3037 696
rect 2943 689 3037 692
rect 2943 682 2992 689
rect 2943 676 2973 682
rect 2992 677 2997 682
rect 2909 660 2989 676
rect 3001 668 3037 689
rect 3098 684 3287 708
rect 3332 707 3379 708
rect 3345 702 3379 707
rect 3113 681 3287 684
rect 3106 678 3287 681
rect 3315 701 3379 702
rect 2909 658 2928 660
rect 2943 658 2977 660
rect 2909 642 2989 658
rect 2909 636 2928 642
rect 2625 610 2728 620
rect 2579 608 2728 610
rect 2749 608 2784 620
rect 2418 606 2580 608
rect 2430 586 2449 606
rect 2464 604 2494 606
rect 2313 578 2354 586
rect 2436 583 2449 586
rect 2501 590 2580 606
rect 2612 606 2784 608
rect 2612 590 2691 606
rect 2698 604 2728 606
rect 2276 568 2305 578
rect 2319 568 2348 578
rect 2363 568 2393 583
rect 2436 579 2479 583
rect 2501 579 2691 590
rect 2756 586 2762 606
rect 2713 579 2743 583
rect 2436 578 2743 579
rect 2436 568 2479 578
rect 2486 568 2516 578
rect 2517 568 2675 578
rect 2679 568 2709 578
rect 2713 568 2743 578
rect 2771 568 2784 606
rect 2856 620 2885 636
rect 2899 620 2928 636
rect 2943 626 2973 642
rect 3001 620 3007 668
rect 3010 662 3029 668
rect 3044 662 3074 670
rect 3010 654 3074 662
rect 3010 638 3090 654
rect 3106 647 3168 678
rect 3184 647 3246 678
rect 3315 676 3364 701
rect 3379 676 3409 692
rect 3278 662 3308 670
rect 3315 668 3425 676
rect 3278 654 3323 662
rect 3010 636 3029 638
rect 3044 636 3090 638
rect 3010 620 3090 636
rect 3117 634 3152 647
rect 3193 644 3230 647
rect 3193 642 3235 644
rect 3122 631 3152 634
rect 3131 627 3138 631
rect 3138 626 3139 627
rect 3097 620 3107 626
rect 2856 612 2891 620
rect 2856 586 2857 612
rect 2864 586 2891 612
rect 2799 568 2829 583
rect 2856 578 2891 586
rect 2893 612 2934 620
rect 2893 586 2908 612
rect 2915 586 2934 612
rect 2998 608 3029 620
rect 3044 608 3147 620
rect 3159 610 3185 636
rect 3200 631 3230 642
rect 3262 638 3324 654
rect 3262 636 3308 638
rect 3262 620 3324 636
rect 3336 620 3342 668
rect 3345 660 3425 668
rect 3345 658 3364 660
rect 3379 658 3413 660
rect 3345 642 3425 658
rect 3345 620 3364 642
rect 3379 626 3409 642
rect 3437 636 3443 710
rect 3446 636 3465 780
rect 3480 636 3486 780
rect 3495 710 3508 780
rect 3560 776 3582 780
rect 3553 754 3582 768
rect 3635 754 3651 768
rect 3689 765 3695 766
rect 3702 765 3810 780
rect 3817 765 3823 766
rect 3831 765 3846 780
rect 3912 774 3931 777
rect 3553 752 3651 754
rect 3678 752 3846 765
rect 3861 754 3877 768
rect 3912 755 3934 774
rect 3944 768 3960 769
rect 3943 766 3960 768
rect 3944 761 3960 766
rect 3934 754 3940 755
rect 3943 754 3972 761
rect 3861 753 3972 754
rect 3861 752 3978 753
rect 3537 744 3588 752
rect 3635 744 3669 752
rect 3537 732 3562 744
rect 3569 732 3588 744
rect 3642 742 3669 744
rect 3678 742 3899 752
rect 3934 749 3940 752
rect 3642 738 3899 742
rect 3537 724 3588 732
rect 3635 724 3899 738
rect 3943 744 3978 752
rect 3489 676 3508 710
rect 3553 716 3582 724
rect 3553 710 3570 716
rect 3553 708 3587 710
rect 3635 708 3651 724
rect 3652 714 3860 724
rect 3861 714 3877 724
rect 3925 720 3940 735
rect 3943 732 3944 744
rect 3951 732 3978 744
rect 3943 724 3978 732
rect 3943 723 3972 724
rect 3663 710 3877 714
rect 3678 708 3877 710
rect 3912 710 3925 720
rect 3943 710 3960 723
rect 3912 708 3960 710
rect 3554 704 3587 708
rect 3550 702 3587 704
rect 3550 701 3617 702
rect 3550 696 3581 701
rect 3587 696 3617 701
rect 3550 692 3617 696
rect 3523 689 3617 692
rect 3523 682 3572 689
rect 3523 676 3553 682
rect 3572 677 3577 682
rect 3489 660 3569 676
rect 3581 668 3617 689
rect 3678 684 3867 708
rect 3912 707 3959 708
rect 3925 702 3959 707
rect 3693 681 3867 684
rect 3686 678 3867 681
rect 3895 701 3959 702
rect 3489 658 3508 660
rect 3523 658 3557 660
rect 3489 642 3569 658
rect 3489 636 3508 642
rect 3205 610 3308 620
rect 3159 608 3308 610
rect 3329 608 3364 620
rect 2998 606 3160 608
rect 3010 586 3029 606
rect 3044 604 3074 606
rect 2893 578 2934 586
rect 3016 583 3029 586
rect 3081 590 3160 606
rect 3192 606 3364 608
rect 3192 590 3271 606
rect 3278 604 3308 606
rect 2856 568 2885 578
rect 2899 568 2928 578
rect 2943 568 2973 583
rect 3016 579 3059 583
rect 3081 579 3271 590
rect 3336 586 3342 606
rect 3293 579 3323 583
rect 3016 578 3323 579
rect 3016 568 3059 578
rect 3066 568 3096 578
rect 3097 568 3255 578
rect 3259 568 3289 578
rect 3293 568 3323 578
rect 3351 568 3364 606
rect 3436 620 3465 636
rect 3479 620 3508 636
rect 3523 626 3553 642
rect 3581 620 3587 668
rect 3590 662 3609 668
rect 3624 662 3654 670
rect 3590 654 3654 662
rect 3590 638 3670 654
rect 3686 647 3748 678
rect 3764 647 3826 678
rect 3895 676 3944 701
rect 3959 676 3989 692
rect 3858 662 3888 670
rect 3895 668 4005 676
rect 3858 654 3903 662
rect 3590 636 3609 638
rect 3624 636 3670 638
rect 3590 620 3670 636
rect 3697 634 3732 647
rect 3773 644 3810 647
rect 3773 642 3815 644
rect 3702 631 3732 634
rect 3711 627 3718 631
rect 3718 626 3719 627
rect 3677 620 3687 626
rect 3436 612 3471 620
rect 3436 586 3437 612
rect 3444 586 3471 612
rect 3379 568 3409 583
rect 3436 578 3471 586
rect 3473 612 3514 620
rect 3473 586 3488 612
rect 3495 586 3514 612
rect 3578 608 3609 620
rect 3624 608 3727 620
rect 3739 610 3765 636
rect 3780 631 3810 642
rect 3842 638 3904 654
rect 3842 636 3888 638
rect 3842 620 3904 636
rect 3916 620 3922 668
rect 3925 660 4005 668
rect 3925 658 3944 660
rect 3959 658 3993 660
rect 3925 642 4005 658
rect 3925 620 3944 642
rect 3959 626 3989 642
rect 4017 636 4023 710
rect 4026 636 4045 780
rect 4060 636 4066 780
rect 4075 710 4088 780
rect 4140 776 4162 780
rect 4133 754 4162 768
rect 4215 754 4231 768
rect 4269 765 4275 766
rect 4282 765 4390 780
rect 4397 765 4403 766
rect 4411 765 4426 780
rect 4492 774 4511 777
rect 4133 752 4231 754
rect 4258 752 4426 765
rect 4441 754 4457 768
rect 4492 755 4514 774
rect 4524 768 4540 769
rect 4523 766 4540 768
rect 4524 761 4540 766
rect 4514 754 4520 755
rect 4523 754 4552 761
rect 4441 753 4552 754
rect 4441 752 4558 753
rect 4117 744 4168 752
rect 4215 744 4249 752
rect 4117 732 4142 744
rect 4149 732 4168 744
rect 4222 742 4249 744
rect 4258 742 4479 752
rect 4514 749 4520 752
rect 4222 738 4479 742
rect 4117 724 4168 732
rect 4215 724 4479 738
rect 4523 744 4558 752
rect 4069 676 4088 710
rect 4133 716 4162 724
rect 4133 710 4150 716
rect 4133 708 4167 710
rect 4215 708 4231 724
rect 4232 714 4440 724
rect 4441 714 4457 724
rect 4505 720 4520 735
rect 4523 732 4524 744
rect 4531 732 4558 744
rect 4523 724 4558 732
rect 4523 723 4552 724
rect 4243 710 4457 714
rect 4258 708 4457 710
rect 4492 710 4505 720
rect 4523 710 4540 723
rect 4492 708 4540 710
rect 4134 704 4167 708
rect 4130 702 4167 704
rect 4130 701 4197 702
rect 4130 696 4161 701
rect 4167 696 4197 701
rect 4130 692 4197 696
rect 4103 689 4197 692
rect 4103 682 4152 689
rect 4103 676 4133 682
rect 4152 677 4157 682
rect 4069 660 4149 676
rect 4161 668 4197 689
rect 4258 684 4447 708
rect 4492 707 4539 708
rect 4505 702 4539 707
rect 4273 681 4447 684
rect 4266 678 4447 681
rect 4475 701 4539 702
rect 4069 658 4088 660
rect 4103 658 4137 660
rect 4069 642 4149 658
rect 4069 636 4088 642
rect 3785 610 3888 620
rect 3739 608 3888 610
rect 3909 608 3944 620
rect 3578 606 3740 608
rect 3590 586 3609 606
rect 3624 604 3654 606
rect 3473 578 3514 586
rect 3596 583 3609 586
rect 3661 590 3740 606
rect 3772 606 3944 608
rect 3772 590 3851 606
rect 3858 604 3888 606
rect 3436 568 3465 578
rect 3479 568 3508 578
rect 3523 568 3553 583
rect 3596 579 3639 583
rect 3661 579 3851 590
rect 3916 586 3922 606
rect 3873 579 3903 583
rect 3596 578 3903 579
rect 3596 568 3639 578
rect 3646 568 3676 578
rect 3677 568 3835 578
rect 3839 568 3869 578
rect 3873 568 3903 578
rect 3931 568 3944 606
rect 4016 620 4045 636
rect 4059 620 4088 636
rect 4103 626 4133 642
rect 4161 620 4167 668
rect 4170 662 4189 668
rect 4204 662 4234 670
rect 4170 654 4234 662
rect 4170 638 4250 654
rect 4266 647 4328 678
rect 4344 647 4406 678
rect 4475 676 4524 701
rect 4539 676 4569 692
rect 4438 662 4468 670
rect 4475 668 4585 676
rect 4438 654 4483 662
rect 4170 636 4189 638
rect 4204 636 4250 638
rect 4170 620 4250 636
rect 4277 634 4312 647
rect 4353 644 4390 647
rect 4353 642 4395 644
rect 4282 631 4312 634
rect 4291 627 4298 631
rect 4298 626 4299 627
rect 4257 620 4267 626
rect 4016 612 4051 620
rect 4016 586 4017 612
rect 4024 586 4051 612
rect 3959 568 3989 583
rect 4016 578 4051 586
rect 4053 612 4094 620
rect 4053 586 4068 612
rect 4075 586 4094 612
rect 4158 608 4189 620
rect 4204 608 4307 620
rect 4319 610 4345 636
rect 4360 631 4390 642
rect 4422 638 4484 654
rect 4422 636 4468 638
rect 4422 620 4484 636
rect 4496 620 4502 668
rect 4505 660 4585 668
rect 4505 658 4524 660
rect 4539 658 4573 660
rect 4505 642 4585 658
rect 4505 620 4524 642
rect 4539 626 4569 642
rect 4597 636 4603 710
rect 4606 636 4625 780
rect 4640 636 4646 780
rect 4655 710 4668 780
rect 4720 776 4742 780
rect 4713 754 4742 768
rect 4795 754 4811 768
rect 4849 765 4855 766
rect 4862 765 4970 780
rect 4977 765 4983 766
rect 4991 765 5006 780
rect 5072 774 5091 777
rect 4713 752 4811 754
rect 4838 752 5006 765
rect 5021 754 5037 768
rect 5072 755 5094 774
rect 5104 768 5120 769
rect 5103 766 5120 768
rect 5104 761 5120 766
rect 5094 754 5100 755
rect 5103 754 5132 761
rect 5021 753 5132 754
rect 5021 752 5138 753
rect 4697 744 4748 752
rect 4795 744 4829 752
rect 4697 732 4722 744
rect 4729 732 4748 744
rect 4802 742 4829 744
rect 4838 742 5059 752
rect 5094 749 5100 752
rect 4802 738 5059 742
rect 4697 724 4748 732
rect 4795 724 5059 738
rect 5103 744 5138 752
rect 4649 676 4668 710
rect 4713 716 4742 724
rect 4713 710 4730 716
rect 4713 708 4747 710
rect 4795 708 4811 724
rect 4812 714 5020 724
rect 5021 714 5037 724
rect 5085 720 5100 735
rect 5103 732 5104 744
rect 5111 732 5138 744
rect 5103 724 5138 732
rect 5103 723 5132 724
rect 4823 710 5037 714
rect 4838 708 5037 710
rect 5072 710 5085 720
rect 5103 710 5120 723
rect 5072 708 5120 710
rect 4714 704 4747 708
rect 4710 702 4747 704
rect 4710 701 4777 702
rect 4710 696 4741 701
rect 4747 696 4777 701
rect 4710 692 4777 696
rect 4683 689 4777 692
rect 4683 682 4732 689
rect 4683 676 4713 682
rect 4732 677 4737 682
rect 4649 660 4729 676
rect 4741 668 4777 689
rect 4838 684 5027 708
rect 5072 707 5119 708
rect 5085 702 5119 707
rect 4853 681 5027 684
rect 4846 678 5027 681
rect 5055 701 5119 702
rect 4649 658 4668 660
rect 4683 658 4717 660
rect 4649 642 4729 658
rect 4649 636 4668 642
rect 4365 610 4468 620
rect 4319 608 4468 610
rect 4489 608 4524 620
rect 4158 606 4320 608
rect 4170 586 4189 606
rect 4204 604 4234 606
rect 4053 578 4094 586
rect 4176 583 4189 586
rect 4241 590 4320 606
rect 4352 606 4524 608
rect 4352 590 4431 606
rect 4438 604 4468 606
rect 4016 568 4045 578
rect 4059 568 4088 578
rect 4103 568 4133 583
rect 4176 579 4219 583
rect 4241 579 4431 590
rect 4496 586 4502 606
rect 4453 579 4483 583
rect 4176 578 4483 579
rect 4176 568 4219 578
rect 4226 568 4256 578
rect 4257 568 4415 578
rect 4419 568 4449 578
rect 4453 568 4483 578
rect 4511 568 4524 606
rect 4596 620 4625 636
rect 4639 620 4668 636
rect 4683 626 4713 642
rect 4741 620 4747 668
rect 4750 662 4769 668
rect 4784 662 4814 670
rect 4750 654 4814 662
rect 4750 638 4830 654
rect 4846 647 4908 678
rect 4924 647 4986 678
rect 5055 676 5104 701
rect 5119 676 5149 692
rect 5018 662 5048 670
rect 5055 668 5165 676
rect 5018 654 5063 662
rect 4750 636 4769 638
rect 4784 636 4830 638
rect 4750 620 4830 636
rect 4857 634 4892 647
rect 4933 644 4970 647
rect 4933 642 4975 644
rect 4862 631 4892 634
rect 4871 627 4878 631
rect 4878 626 4879 627
rect 4837 620 4847 626
rect 4596 612 4631 620
rect 4596 586 4597 612
rect 4604 586 4631 612
rect 4539 568 4569 583
rect 4596 578 4631 586
rect 4633 612 4674 620
rect 4633 586 4648 612
rect 4655 586 4674 612
rect 4738 608 4769 620
rect 4784 608 4887 620
rect 4899 610 4925 636
rect 4940 631 4970 642
rect 5002 638 5064 654
rect 5002 636 5048 638
rect 5002 620 5064 636
rect 5076 620 5082 668
rect 5085 660 5165 668
rect 5085 658 5104 660
rect 5119 658 5153 660
rect 5085 642 5165 658
rect 5085 620 5104 642
rect 5119 626 5149 642
rect 5177 636 5183 710
rect 5186 636 5205 780
rect 5220 636 5226 780
rect 5235 710 5248 780
rect 5300 776 5322 780
rect 5293 754 5322 768
rect 5375 754 5391 768
rect 5429 765 5435 766
rect 5442 765 5550 780
rect 5557 765 5563 766
rect 5571 765 5586 780
rect 5652 774 5671 777
rect 5293 752 5391 754
rect 5418 752 5586 765
rect 5601 754 5617 768
rect 5652 755 5674 774
rect 5684 768 5700 769
rect 5683 766 5700 768
rect 5684 761 5700 766
rect 5674 754 5680 755
rect 5683 754 5712 761
rect 5601 753 5712 754
rect 5601 752 5718 753
rect 5277 744 5328 752
rect 5375 744 5409 752
rect 5277 732 5302 744
rect 5309 732 5328 744
rect 5382 742 5409 744
rect 5418 742 5639 752
rect 5674 749 5680 752
rect 5382 738 5639 742
rect 5277 724 5328 732
rect 5375 724 5639 738
rect 5683 744 5718 752
rect 5229 676 5248 710
rect 5293 716 5322 724
rect 5293 710 5310 716
rect 5293 708 5327 710
rect 5375 708 5391 724
rect 5392 714 5600 724
rect 5601 714 5617 724
rect 5665 720 5680 735
rect 5683 732 5684 744
rect 5691 732 5718 744
rect 5683 724 5718 732
rect 5683 723 5712 724
rect 5403 710 5617 714
rect 5418 708 5617 710
rect 5652 710 5665 720
rect 5683 710 5700 723
rect 5652 708 5700 710
rect 5294 704 5327 708
rect 5290 702 5327 704
rect 5290 701 5357 702
rect 5290 696 5321 701
rect 5327 696 5357 701
rect 5290 692 5357 696
rect 5263 689 5357 692
rect 5263 682 5312 689
rect 5263 676 5293 682
rect 5312 677 5317 682
rect 5229 660 5309 676
rect 5321 668 5357 689
rect 5418 684 5607 708
rect 5652 707 5699 708
rect 5665 702 5699 707
rect 5433 681 5607 684
rect 5426 678 5607 681
rect 5635 701 5699 702
rect 5229 658 5248 660
rect 5263 658 5297 660
rect 5229 642 5309 658
rect 5229 636 5248 642
rect 4945 610 5048 620
rect 4899 608 5048 610
rect 5069 608 5104 620
rect 4738 606 4900 608
rect 4750 586 4769 606
rect 4784 604 4814 606
rect 4633 578 4674 586
rect 4756 583 4769 586
rect 4821 590 4900 606
rect 4932 606 5104 608
rect 4932 590 5011 606
rect 5018 604 5048 606
rect 4596 568 4625 578
rect 4639 568 4668 578
rect 4683 568 4713 583
rect 4756 579 4799 583
rect 4821 579 5011 590
rect 5076 586 5082 606
rect 5033 579 5063 583
rect 4756 578 5063 579
rect 4756 568 4799 578
rect 4806 568 4836 578
rect 4837 568 4995 578
rect 4999 568 5029 578
rect 5033 568 5063 578
rect 5091 568 5104 606
rect 5176 620 5205 636
rect 5219 620 5248 636
rect 5263 626 5293 642
rect 5321 620 5327 668
rect 5330 662 5349 668
rect 5364 662 5394 670
rect 5330 654 5394 662
rect 5330 638 5410 654
rect 5426 647 5488 678
rect 5504 647 5566 678
rect 5635 676 5684 701
rect 5699 676 5729 692
rect 5598 662 5628 670
rect 5635 668 5745 676
rect 5598 654 5643 662
rect 5330 636 5349 638
rect 5364 636 5410 638
rect 5330 620 5410 636
rect 5437 634 5472 647
rect 5513 644 5550 647
rect 5513 642 5555 644
rect 5442 631 5472 634
rect 5451 627 5458 631
rect 5458 626 5459 627
rect 5417 620 5427 626
rect 5176 612 5211 620
rect 5176 586 5177 612
rect 5184 586 5211 612
rect 5119 568 5149 583
rect 5176 578 5211 586
rect 5213 612 5254 620
rect 5213 586 5228 612
rect 5235 586 5254 612
rect 5318 608 5349 620
rect 5364 608 5467 620
rect 5479 610 5505 636
rect 5520 631 5550 642
rect 5582 638 5644 654
rect 5582 636 5628 638
rect 5582 620 5644 636
rect 5656 620 5662 668
rect 5665 660 5745 668
rect 5665 658 5684 660
rect 5699 658 5733 660
rect 5665 642 5745 658
rect 5665 620 5684 642
rect 5699 626 5729 642
rect 5757 636 5763 710
rect 5766 636 5785 780
rect 5800 636 5806 780
rect 5815 710 5828 780
rect 5880 776 5902 780
rect 5873 754 5902 768
rect 5955 754 5971 768
rect 6009 765 6015 766
rect 6022 765 6130 780
rect 6137 765 6143 766
rect 6151 765 6166 780
rect 6232 774 6251 777
rect 5873 752 5971 754
rect 5998 752 6166 765
rect 6181 754 6197 768
rect 6232 755 6254 774
rect 6264 768 6280 769
rect 6263 766 6280 768
rect 6264 761 6280 766
rect 6254 754 6260 755
rect 6263 754 6292 761
rect 6181 753 6292 754
rect 6181 752 6298 753
rect 5857 744 5908 752
rect 5955 744 5989 752
rect 5857 732 5882 744
rect 5889 732 5908 744
rect 5962 742 5989 744
rect 5998 742 6219 752
rect 6254 749 6260 752
rect 5962 738 6219 742
rect 5857 724 5908 732
rect 5955 724 6219 738
rect 6263 744 6298 752
rect 5809 676 5828 710
rect 5873 716 5902 724
rect 5873 710 5890 716
rect 5873 708 5907 710
rect 5955 708 5971 724
rect 5972 714 6180 724
rect 6181 714 6197 724
rect 6245 720 6260 735
rect 6263 732 6264 744
rect 6271 732 6298 744
rect 6263 724 6298 732
rect 6263 723 6292 724
rect 5983 710 6197 714
rect 5998 708 6197 710
rect 6232 710 6245 720
rect 6263 710 6280 723
rect 6232 708 6280 710
rect 5874 704 5907 708
rect 5870 702 5907 704
rect 5870 701 5937 702
rect 5870 696 5901 701
rect 5907 696 5937 701
rect 5870 692 5937 696
rect 5843 689 5937 692
rect 5843 682 5892 689
rect 5843 676 5873 682
rect 5892 677 5897 682
rect 5809 660 5889 676
rect 5901 668 5937 689
rect 5998 684 6187 708
rect 6232 707 6279 708
rect 6245 702 6279 707
rect 6013 681 6187 684
rect 6006 678 6187 681
rect 6215 701 6279 702
rect 5809 658 5828 660
rect 5843 658 5877 660
rect 5809 642 5889 658
rect 5809 636 5828 642
rect 5525 610 5628 620
rect 5479 608 5628 610
rect 5649 608 5684 620
rect 5318 606 5480 608
rect 5330 586 5349 606
rect 5364 604 5394 606
rect 5213 578 5254 586
rect 5336 583 5349 586
rect 5401 590 5480 606
rect 5512 606 5684 608
rect 5512 590 5591 606
rect 5598 604 5628 606
rect 5176 568 5205 578
rect 5219 568 5248 578
rect 5263 568 5293 583
rect 5336 579 5379 583
rect 5401 579 5591 590
rect 5656 586 5662 606
rect 5613 579 5643 583
rect 5336 578 5643 579
rect 5336 568 5379 578
rect 5386 568 5416 578
rect 5417 568 5575 578
rect 5579 568 5609 578
rect 5613 568 5643 578
rect 5671 568 5684 606
rect 5756 620 5785 636
rect 5799 620 5828 636
rect 5843 626 5873 642
rect 5901 620 5907 668
rect 5910 662 5929 668
rect 5944 662 5974 670
rect 5910 654 5974 662
rect 5910 638 5990 654
rect 6006 647 6068 678
rect 6084 647 6146 678
rect 6215 676 6264 701
rect 6279 676 6309 692
rect 6178 662 6208 670
rect 6215 668 6325 676
rect 6178 654 6223 662
rect 5910 636 5929 638
rect 5944 636 5990 638
rect 5910 620 5990 636
rect 6017 634 6052 647
rect 6093 644 6130 647
rect 6093 642 6135 644
rect 6022 631 6052 634
rect 6031 627 6038 631
rect 6038 626 6039 627
rect 5997 620 6007 626
rect 5756 612 5791 620
rect 5756 586 5757 612
rect 5764 586 5791 612
rect 5699 568 5729 583
rect 5756 578 5791 586
rect 5793 612 5834 620
rect 5793 586 5808 612
rect 5815 586 5834 612
rect 5898 608 5929 620
rect 5944 608 6047 620
rect 6059 610 6085 636
rect 6100 631 6130 642
rect 6162 638 6224 654
rect 6162 636 6208 638
rect 6162 620 6224 636
rect 6236 620 6242 668
rect 6245 660 6325 668
rect 6245 658 6264 660
rect 6279 658 6313 660
rect 6245 642 6325 658
rect 6245 620 6264 642
rect 6279 626 6309 642
rect 6337 636 6343 710
rect 6346 636 6365 780
rect 6380 636 6386 780
rect 6395 710 6408 780
rect 6460 776 6482 780
rect 6453 754 6482 768
rect 6535 754 6551 768
rect 6589 765 6595 766
rect 6602 765 6710 780
rect 6717 765 6723 766
rect 6731 765 6746 780
rect 6812 774 6831 777
rect 6453 752 6551 754
rect 6578 752 6746 765
rect 6761 754 6777 768
rect 6812 755 6834 774
rect 6844 768 6860 769
rect 6843 766 6860 768
rect 6844 761 6860 766
rect 6834 754 6840 755
rect 6843 754 6872 761
rect 6761 753 6872 754
rect 6761 752 6878 753
rect 6437 744 6488 752
rect 6535 744 6569 752
rect 6437 732 6462 744
rect 6469 732 6488 744
rect 6542 742 6569 744
rect 6578 742 6799 752
rect 6834 749 6840 752
rect 6542 738 6799 742
rect 6437 724 6488 732
rect 6535 724 6799 738
rect 6843 744 6878 752
rect 6389 676 6408 710
rect 6453 716 6482 724
rect 6453 710 6470 716
rect 6453 708 6487 710
rect 6535 708 6551 724
rect 6552 714 6760 724
rect 6761 714 6777 724
rect 6825 720 6840 735
rect 6843 732 6844 744
rect 6851 732 6878 744
rect 6843 724 6878 732
rect 6843 723 6872 724
rect 6563 710 6777 714
rect 6578 708 6777 710
rect 6812 710 6825 720
rect 6843 710 6860 723
rect 6812 708 6860 710
rect 6454 704 6487 708
rect 6450 702 6487 704
rect 6450 701 6517 702
rect 6450 696 6481 701
rect 6487 696 6517 701
rect 6450 692 6517 696
rect 6423 689 6517 692
rect 6423 682 6472 689
rect 6423 676 6453 682
rect 6472 677 6477 682
rect 6389 660 6469 676
rect 6481 668 6517 689
rect 6578 684 6767 708
rect 6812 707 6859 708
rect 6825 702 6859 707
rect 6593 681 6767 684
rect 6586 678 6767 681
rect 6795 701 6859 702
rect 6389 658 6408 660
rect 6423 658 6457 660
rect 6389 642 6469 658
rect 6389 636 6408 642
rect 6105 610 6208 620
rect 6059 608 6208 610
rect 6229 608 6264 620
rect 5898 606 6060 608
rect 5910 586 5929 606
rect 5944 604 5974 606
rect 5793 578 5834 586
rect 5916 583 5929 586
rect 5981 590 6060 606
rect 6092 606 6264 608
rect 6092 590 6171 606
rect 6178 604 6208 606
rect 5756 568 5785 578
rect 5799 568 5828 578
rect 5843 568 5873 583
rect 5916 579 5959 583
rect 5981 579 6171 590
rect 6236 586 6242 606
rect 6193 579 6223 583
rect 5916 578 6223 579
rect 5916 568 5959 578
rect 5966 568 5996 578
rect 5997 568 6155 578
rect 6159 568 6189 578
rect 6193 568 6223 578
rect 6251 568 6264 606
rect 6336 620 6365 636
rect 6379 620 6408 636
rect 6423 626 6453 642
rect 6481 620 6487 668
rect 6490 662 6509 668
rect 6524 662 6554 670
rect 6490 654 6554 662
rect 6490 638 6570 654
rect 6586 647 6648 678
rect 6664 647 6726 678
rect 6795 676 6844 701
rect 6859 676 6889 692
rect 6758 662 6788 670
rect 6795 668 6905 676
rect 6758 654 6803 662
rect 6490 636 6509 638
rect 6524 636 6570 638
rect 6490 620 6570 636
rect 6597 634 6632 647
rect 6673 644 6710 647
rect 6673 642 6715 644
rect 6602 631 6632 634
rect 6611 627 6618 631
rect 6618 626 6619 627
rect 6577 620 6587 626
rect 6336 612 6371 620
rect 6336 586 6337 612
rect 6344 586 6371 612
rect 6279 568 6309 583
rect 6336 578 6371 586
rect 6373 612 6414 620
rect 6373 586 6388 612
rect 6395 586 6414 612
rect 6478 608 6509 620
rect 6524 608 6627 620
rect 6639 610 6665 636
rect 6680 631 6710 642
rect 6742 638 6804 654
rect 6742 636 6788 638
rect 6742 620 6804 636
rect 6816 620 6822 668
rect 6825 660 6905 668
rect 6825 658 6844 660
rect 6859 658 6893 660
rect 6825 642 6905 658
rect 6825 620 6844 642
rect 6859 626 6889 642
rect 6917 636 6923 710
rect 6926 636 6945 780
rect 6960 636 6966 780
rect 6975 710 6988 780
rect 7040 776 7062 780
rect 7033 754 7062 768
rect 7115 754 7131 768
rect 7169 765 7175 766
rect 7182 765 7290 780
rect 7297 765 7303 766
rect 7311 765 7326 780
rect 7392 774 7411 777
rect 7033 752 7131 754
rect 7158 752 7326 765
rect 7341 754 7357 768
rect 7392 755 7414 774
rect 7424 768 7440 769
rect 7423 766 7440 768
rect 7424 761 7440 766
rect 7414 754 7420 755
rect 7423 754 7452 761
rect 7341 753 7452 754
rect 7341 752 7458 753
rect 7017 744 7068 752
rect 7115 744 7149 752
rect 7017 732 7042 744
rect 7049 732 7068 744
rect 7122 742 7149 744
rect 7158 742 7379 752
rect 7414 749 7420 752
rect 7122 738 7379 742
rect 7017 724 7068 732
rect 7115 724 7379 738
rect 7423 744 7458 752
rect 6969 676 6988 710
rect 7033 716 7062 724
rect 7033 710 7050 716
rect 7033 708 7067 710
rect 7115 708 7131 724
rect 7132 714 7340 724
rect 7341 714 7357 724
rect 7405 720 7420 735
rect 7423 732 7424 744
rect 7431 732 7458 744
rect 7423 724 7458 732
rect 7423 723 7452 724
rect 7143 710 7357 714
rect 7158 708 7357 710
rect 7392 710 7405 720
rect 7423 710 7440 723
rect 7392 708 7440 710
rect 7034 704 7067 708
rect 7030 702 7067 704
rect 7030 701 7097 702
rect 7030 696 7061 701
rect 7067 696 7097 701
rect 7030 692 7097 696
rect 7003 689 7097 692
rect 7003 682 7052 689
rect 7003 676 7033 682
rect 7052 677 7057 682
rect 6969 660 7049 676
rect 7061 668 7097 689
rect 7158 684 7347 708
rect 7392 707 7439 708
rect 7405 702 7439 707
rect 7173 681 7347 684
rect 7166 678 7347 681
rect 7375 701 7439 702
rect 6969 658 6988 660
rect 7003 658 7037 660
rect 6969 642 7049 658
rect 6969 636 6988 642
rect 6685 610 6788 620
rect 6639 608 6788 610
rect 6809 608 6844 620
rect 6478 606 6640 608
rect 6490 586 6509 606
rect 6524 604 6554 606
rect 6373 578 6414 586
rect 6496 583 6509 586
rect 6561 590 6640 606
rect 6672 606 6844 608
rect 6672 590 6751 606
rect 6758 604 6788 606
rect 6336 568 6365 578
rect 6379 568 6408 578
rect 6423 568 6453 583
rect 6496 579 6539 583
rect 6561 579 6751 590
rect 6816 586 6822 606
rect 6773 579 6803 583
rect 6496 578 6803 579
rect 6496 568 6539 578
rect 6546 568 6576 578
rect 6577 568 6735 578
rect 6739 568 6769 578
rect 6773 568 6803 578
rect 6831 568 6844 606
rect 6916 620 6945 636
rect 6959 620 6988 636
rect 7003 626 7033 642
rect 7061 620 7067 668
rect 7070 662 7089 668
rect 7104 662 7134 670
rect 7070 654 7134 662
rect 7070 638 7150 654
rect 7166 647 7228 678
rect 7244 647 7306 678
rect 7375 676 7424 701
rect 7439 676 7469 692
rect 7338 662 7368 670
rect 7375 668 7485 676
rect 7338 654 7383 662
rect 7070 636 7089 638
rect 7104 636 7150 638
rect 7070 620 7150 636
rect 7177 634 7212 647
rect 7253 644 7290 647
rect 7253 642 7295 644
rect 7182 631 7212 634
rect 7191 627 7198 631
rect 7198 626 7199 627
rect 7157 620 7167 626
rect 6916 612 6951 620
rect 6916 586 6917 612
rect 6924 586 6951 612
rect 6859 568 6889 583
rect 6916 578 6951 586
rect 6953 612 6994 620
rect 6953 586 6968 612
rect 6975 586 6994 612
rect 7058 608 7089 620
rect 7104 608 7207 620
rect 7219 610 7245 636
rect 7260 631 7290 642
rect 7322 638 7384 654
rect 7322 636 7368 638
rect 7322 620 7384 636
rect 7396 620 7402 668
rect 7405 660 7485 668
rect 7405 658 7424 660
rect 7439 658 7473 660
rect 7405 642 7485 658
rect 7405 620 7424 642
rect 7439 626 7469 642
rect 7497 636 7503 710
rect 7506 636 7525 780
rect 7540 636 7546 780
rect 7555 710 7568 780
rect 7620 776 7642 780
rect 7613 754 7642 768
rect 7695 754 7711 768
rect 7749 765 7755 766
rect 7762 765 7870 780
rect 7877 765 7883 766
rect 7891 765 7906 780
rect 7972 774 7991 777
rect 7613 752 7711 754
rect 7738 752 7906 765
rect 7921 754 7937 768
rect 7972 755 7994 774
rect 8004 768 8020 769
rect 8003 766 8020 768
rect 8004 761 8020 766
rect 7994 754 8000 755
rect 8003 754 8032 761
rect 7921 753 8032 754
rect 7921 752 8038 753
rect 7597 744 7648 752
rect 7695 744 7729 752
rect 7597 732 7622 744
rect 7629 732 7648 744
rect 7702 742 7729 744
rect 7738 742 7959 752
rect 7994 749 8000 752
rect 7702 738 7959 742
rect 7597 724 7648 732
rect 7695 724 7959 738
rect 8003 744 8038 752
rect 7549 676 7568 710
rect 7613 716 7642 724
rect 7613 710 7630 716
rect 7613 708 7647 710
rect 7695 708 7711 724
rect 7712 714 7920 724
rect 7921 714 7937 724
rect 7985 720 8000 735
rect 8003 732 8004 744
rect 8011 732 8038 744
rect 8003 724 8038 732
rect 8003 723 8032 724
rect 7723 710 7937 714
rect 7738 708 7937 710
rect 7972 710 7985 720
rect 8003 710 8020 723
rect 7972 708 8020 710
rect 7614 704 7647 708
rect 7610 702 7647 704
rect 7610 701 7677 702
rect 7610 696 7641 701
rect 7647 696 7677 701
rect 7610 692 7677 696
rect 7583 689 7677 692
rect 7583 682 7632 689
rect 7583 676 7613 682
rect 7632 677 7637 682
rect 7549 660 7629 676
rect 7641 668 7677 689
rect 7738 684 7927 708
rect 7972 707 8019 708
rect 7985 702 8019 707
rect 7753 681 7927 684
rect 7746 678 7927 681
rect 7955 701 8019 702
rect 7549 658 7568 660
rect 7583 658 7617 660
rect 7549 642 7629 658
rect 7549 636 7568 642
rect 7265 610 7368 620
rect 7219 608 7368 610
rect 7389 608 7424 620
rect 7058 606 7220 608
rect 7070 586 7089 606
rect 7104 604 7134 606
rect 6953 578 6994 586
rect 7076 583 7089 586
rect 7141 590 7220 606
rect 7252 606 7424 608
rect 7252 590 7331 606
rect 7338 604 7368 606
rect 6916 568 6945 578
rect 6959 568 6988 578
rect 7003 568 7033 583
rect 7076 579 7119 583
rect 7141 579 7331 590
rect 7396 586 7402 606
rect 7353 579 7383 583
rect 7076 578 7383 579
rect 7076 568 7119 578
rect 7126 568 7156 578
rect 7157 568 7315 578
rect 7319 568 7349 578
rect 7353 568 7383 578
rect 7411 568 7424 606
rect 7496 620 7525 636
rect 7539 620 7568 636
rect 7583 626 7613 642
rect 7641 620 7647 668
rect 7650 662 7669 668
rect 7684 662 7714 670
rect 7650 654 7714 662
rect 7650 638 7730 654
rect 7746 647 7808 678
rect 7824 647 7886 678
rect 7955 676 8004 701
rect 8019 676 8049 692
rect 7918 662 7948 670
rect 7955 668 8065 676
rect 7918 654 7963 662
rect 7650 636 7669 638
rect 7684 636 7730 638
rect 7650 620 7730 636
rect 7757 634 7792 647
rect 7833 644 7870 647
rect 7833 642 7875 644
rect 7762 631 7792 634
rect 7771 627 7778 631
rect 7778 626 7779 627
rect 7737 620 7747 626
rect 7496 612 7531 620
rect 7496 586 7497 612
rect 7504 586 7531 612
rect 7439 568 7469 583
rect 7496 578 7531 586
rect 7533 612 7574 620
rect 7533 586 7548 612
rect 7555 586 7574 612
rect 7638 608 7669 620
rect 7684 608 7787 620
rect 7799 610 7825 636
rect 7840 631 7870 642
rect 7902 638 7964 654
rect 7902 636 7948 638
rect 7902 620 7964 636
rect 7976 620 7982 668
rect 7985 660 8065 668
rect 7985 658 8004 660
rect 8019 658 8053 660
rect 7985 642 8065 658
rect 7985 620 8004 642
rect 8019 626 8049 642
rect 8077 636 8083 710
rect 8086 636 8105 780
rect 8120 636 8126 780
rect 8135 710 8148 780
rect 8200 776 8222 780
rect 8193 754 8222 768
rect 8275 754 8291 768
rect 8329 765 8335 766
rect 8342 765 8450 780
rect 8457 765 8463 766
rect 8471 765 8486 780
rect 8552 774 8571 777
rect 8193 752 8291 754
rect 8318 752 8486 765
rect 8501 754 8517 768
rect 8552 755 8574 774
rect 8584 768 8600 769
rect 8583 766 8600 768
rect 8584 761 8600 766
rect 8574 754 8580 755
rect 8583 754 8612 761
rect 8501 753 8612 754
rect 8501 752 8618 753
rect 8177 744 8228 752
rect 8275 744 8309 752
rect 8177 732 8202 744
rect 8209 732 8228 744
rect 8282 742 8309 744
rect 8318 742 8539 752
rect 8574 749 8580 752
rect 8282 738 8539 742
rect 8177 724 8228 732
rect 8275 724 8539 738
rect 8583 744 8618 752
rect 8129 676 8148 710
rect 8193 716 8222 724
rect 8193 710 8210 716
rect 8193 708 8227 710
rect 8275 708 8291 724
rect 8292 714 8500 724
rect 8501 714 8517 724
rect 8565 720 8580 735
rect 8583 732 8584 744
rect 8591 732 8618 744
rect 8583 724 8618 732
rect 8583 723 8612 724
rect 8303 710 8517 714
rect 8318 708 8517 710
rect 8552 710 8565 720
rect 8583 710 8600 723
rect 8552 708 8600 710
rect 8194 704 8227 708
rect 8190 702 8227 704
rect 8190 701 8257 702
rect 8190 696 8221 701
rect 8227 696 8257 701
rect 8190 692 8257 696
rect 8163 689 8257 692
rect 8163 682 8212 689
rect 8163 676 8193 682
rect 8212 677 8217 682
rect 8129 660 8209 676
rect 8221 668 8257 689
rect 8318 684 8507 708
rect 8552 707 8599 708
rect 8565 702 8599 707
rect 8333 681 8507 684
rect 8326 678 8507 681
rect 8535 701 8599 702
rect 8129 658 8148 660
rect 8163 658 8197 660
rect 8129 642 8209 658
rect 8129 636 8148 642
rect 7845 610 7948 620
rect 7799 608 7948 610
rect 7969 608 8004 620
rect 7638 606 7800 608
rect 7650 586 7669 606
rect 7684 604 7714 606
rect 7533 578 7574 586
rect 7656 583 7669 586
rect 7721 590 7800 606
rect 7832 606 8004 608
rect 7832 590 7911 606
rect 7918 604 7948 606
rect 7496 568 7525 578
rect 7539 568 7568 578
rect 7583 568 7613 583
rect 7656 579 7699 583
rect 7721 579 7911 590
rect 7976 586 7982 606
rect 7933 579 7963 583
rect 7656 578 7963 579
rect 7656 568 7699 578
rect 7706 568 7736 578
rect 7737 568 7895 578
rect 7899 568 7929 578
rect 7933 568 7963 578
rect 7991 568 8004 606
rect 8076 620 8105 636
rect 8119 620 8148 636
rect 8163 626 8193 642
rect 8221 620 8227 668
rect 8230 662 8249 668
rect 8264 662 8294 670
rect 8230 654 8294 662
rect 8230 638 8310 654
rect 8326 647 8388 678
rect 8404 647 8466 678
rect 8535 676 8584 701
rect 8599 676 8629 692
rect 8498 662 8528 670
rect 8535 668 8645 676
rect 8498 654 8543 662
rect 8230 636 8249 638
rect 8264 636 8310 638
rect 8230 620 8310 636
rect 8337 634 8372 647
rect 8413 644 8450 647
rect 8413 642 8455 644
rect 8342 631 8372 634
rect 8351 627 8358 631
rect 8358 626 8359 627
rect 8317 620 8327 626
rect 8076 612 8111 620
rect 8076 586 8077 612
rect 8084 586 8111 612
rect 8019 568 8049 583
rect 8076 578 8111 586
rect 8113 612 8154 620
rect 8113 586 8128 612
rect 8135 586 8154 612
rect 8218 608 8249 620
rect 8264 608 8367 620
rect 8379 610 8405 636
rect 8420 631 8450 642
rect 8482 638 8544 654
rect 8482 636 8528 638
rect 8482 620 8544 636
rect 8556 620 8562 668
rect 8565 660 8645 668
rect 8565 658 8584 660
rect 8599 658 8633 660
rect 8565 642 8645 658
rect 8565 620 8584 642
rect 8599 626 8629 642
rect 8657 636 8663 710
rect 8666 636 8685 780
rect 8700 636 8706 780
rect 8715 710 8728 780
rect 8780 776 8802 780
rect 8773 754 8802 768
rect 8855 754 8871 768
rect 8909 765 8915 766
rect 8922 765 9030 780
rect 9037 765 9043 766
rect 9051 765 9066 780
rect 9132 774 9151 777
rect 8773 752 8871 754
rect 8898 752 9066 765
rect 9081 754 9097 768
rect 9132 755 9154 774
rect 9164 768 9180 769
rect 9163 766 9180 768
rect 9164 761 9180 766
rect 9154 754 9160 755
rect 9163 754 9192 761
rect 9081 753 9192 754
rect 9081 752 9198 753
rect 8757 744 8808 752
rect 8855 744 8889 752
rect 8757 732 8782 744
rect 8789 732 8808 744
rect 8862 742 8889 744
rect 8898 742 9119 752
rect 9154 749 9160 752
rect 8862 738 9119 742
rect 8757 724 8808 732
rect 8855 724 9119 738
rect 9163 744 9198 752
rect 8709 676 8728 710
rect 8773 716 8802 724
rect 8773 710 8790 716
rect 8773 708 8807 710
rect 8855 708 8871 724
rect 8872 714 9080 724
rect 9081 714 9097 724
rect 9145 720 9160 735
rect 9163 732 9164 744
rect 9171 732 9198 744
rect 9163 724 9198 732
rect 9163 723 9192 724
rect 8883 710 9097 714
rect 8898 708 9097 710
rect 9132 710 9145 720
rect 9163 710 9180 723
rect 9132 708 9180 710
rect 8774 704 8807 708
rect 8770 702 8807 704
rect 8770 701 8837 702
rect 8770 696 8801 701
rect 8807 696 8837 701
rect 8770 692 8837 696
rect 8743 689 8837 692
rect 8743 682 8792 689
rect 8743 676 8773 682
rect 8792 677 8797 682
rect 8709 660 8789 676
rect 8801 668 8837 689
rect 8898 684 9087 708
rect 9132 707 9179 708
rect 9145 702 9179 707
rect 8913 681 9087 684
rect 8906 678 9087 681
rect 9115 701 9179 702
rect 8709 658 8728 660
rect 8743 658 8777 660
rect 8709 642 8789 658
rect 8709 636 8728 642
rect 8425 610 8528 620
rect 8379 608 8528 610
rect 8549 608 8584 620
rect 8218 606 8380 608
rect 8230 586 8249 606
rect 8264 604 8294 606
rect 8113 578 8154 586
rect 8236 583 8249 586
rect 8301 590 8380 606
rect 8412 606 8584 608
rect 8412 590 8491 606
rect 8498 604 8528 606
rect 8076 568 8105 578
rect 8119 568 8148 578
rect 8163 568 8193 583
rect 8236 579 8279 583
rect 8301 579 8491 590
rect 8556 586 8562 606
rect 8513 579 8543 583
rect 8236 578 8543 579
rect 8236 568 8279 578
rect 8286 568 8316 578
rect 8317 568 8475 578
rect 8479 568 8509 578
rect 8513 568 8543 578
rect 8571 568 8584 606
rect 8656 620 8685 636
rect 8699 620 8728 636
rect 8743 626 8773 642
rect 8801 620 8807 668
rect 8810 662 8829 668
rect 8844 662 8874 670
rect 8810 654 8874 662
rect 8810 638 8890 654
rect 8906 647 8968 678
rect 8984 647 9046 678
rect 9115 676 9164 701
rect 9179 676 9209 692
rect 9078 662 9108 670
rect 9115 668 9225 676
rect 9078 654 9123 662
rect 8810 636 8829 638
rect 8844 636 8890 638
rect 8810 620 8890 636
rect 8917 634 8952 647
rect 8993 644 9030 647
rect 8993 642 9035 644
rect 8922 631 8952 634
rect 8931 627 8938 631
rect 8938 626 8939 627
rect 8897 620 8907 626
rect 8656 612 8691 620
rect 8656 586 8657 612
rect 8664 586 8691 612
rect 8599 568 8629 583
rect 8656 578 8691 586
rect 8693 612 8734 620
rect 8693 586 8708 612
rect 8715 586 8734 612
rect 8798 608 8829 620
rect 8844 608 8947 620
rect 8959 610 8985 636
rect 9000 631 9030 642
rect 9062 638 9124 654
rect 9062 636 9108 638
rect 9062 620 9124 636
rect 9136 620 9142 668
rect 9145 660 9225 668
rect 9145 658 9164 660
rect 9179 658 9213 660
rect 9145 642 9225 658
rect 9145 620 9164 642
rect 9179 626 9209 642
rect 9237 636 9243 710
rect 9252 636 9265 780
rect 9005 610 9108 620
rect 8959 608 9108 610
rect 9129 608 9164 620
rect 8798 606 8960 608
rect 8810 586 8829 606
rect 8844 604 8874 606
rect 8693 578 8734 586
rect 8816 583 8829 586
rect 8881 590 8960 606
rect 8992 606 9164 608
rect 8992 590 9071 606
rect 9078 604 9108 606
rect 8656 568 8685 578
rect 8699 568 8728 578
rect 8743 568 8773 583
rect 8816 579 8859 583
rect 8881 579 9071 590
rect 9136 586 9142 606
rect 9093 579 9123 583
rect 8816 578 9123 579
rect 8816 568 8859 578
rect 8866 568 8896 578
rect 8897 568 9055 578
rect 9059 568 9089 578
rect 9093 568 9123 578
rect 9151 568 9164 606
rect 9236 620 9265 636
rect 9236 612 9271 620
rect 9236 586 9237 612
rect 9244 586 9271 612
rect 9179 568 9209 583
rect 9236 578 9271 586
rect 9236 568 9265 578
rect -1 562 9265 568
rect 0 554 9265 562
rect 15 525 28 554
rect 43 541 73 554
rect 116 541 159 554
rect 83 527 98 539
rect 117 527 130 541
rect 166 540 386 554
rect 393 541 423 554
rect 198 537 351 540
rect 80 525 102 527
rect 180 525 372 537
rect 451 525 464 554
rect 479 541 509 554
rect 546 525 565 554
rect 580 525 586 554
rect 595 525 608 554
rect 623 541 653 554
rect 696 541 739 554
rect 663 527 678 539
rect 697 527 710 541
rect 746 540 966 554
rect 973 541 1003 554
rect 778 537 931 540
rect 660 525 682 527
rect 760 525 952 537
rect 1031 525 1044 554
rect 1059 541 1089 554
rect 1126 525 1145 554
rect 1160 525 1166 554
rect 1175 525 1188 554
rect 1203 541 1233 554
rect 1276 541 1319 554
rect 1243 527 1258 539
rect 1277 527 1290 541
rect 1326 540 1546 554
rect 1553 541 1583 554
rect 1358 537 1511 540
rect 1240 525 1262 527
rect 1340 525 1532 537
rect 1611 525 1624 554
rect 1639 541 1669 554
rect 1706 525 1725 554
rect 1740 525 1746 554
rect 1755 525 1768 554
rect 1783 541 1813 554
rect 1856 541 1899 554
rect 1823 527 1838 539
rect 1857 527 1870 541
rect 1906 540 2126 554
rect 2133 541 2163 554
rect 1938 537 2091 540
rect 1820 525 1842 527
rect 1920 525 2112 537
rect 2191 525 2204 554
rect 2219 541 2249 554
rect 2286 525 2305 554
rect 2320 525 2326 554
rect 2335 525 2348 554
rect 2363 541 2393 554
rect 2436 541 2479 554
rect 2403 527 2418 539
rect 2437 527 2450 541
rect 2486 540 2706 554
rect 2713 541 2743 554
rect 2518 537 2671 540
rect 2400 525 2422 527
rect 2500 525 2692 537
rect 2771 525 2784 554
rect 2799 541 2829 554
rect 2866 525 2885 554
rect 2900 525 2906 554
rect 2915 525 2928 554
rect 2943 541 2973 554
rect 3016 541 3059 554
rect 2983 527 2998 539
rect 3017 527 3030 541
rect 3066 540 3286 554
rect 3293 541 3323 554
rect 3098 537 3251 540
rect 2980 525 3002 527
rect 3080 525 3272 537
rect 3351 525 3364 554
rect 3379 541 3409 554
rect 3446 525 3465 554
rect 3480 525 3486 554
rect 3495 525 3508 554
rect 3523 541 3553 554
rect 3596 541 3639 554
rect 3563 527 3578 539
rect 3597 527 3610 541
rect 3646 540 3866 554
rect 3873 541 3903 554
rect 3678 537 3831 540
rect 3560 525 3582 527
rect 3660 525 3852 537
rect 3931 525 3944 554
rect 3959 541 3989 554
rect 4026 525 4045 554
rect 4060 525 4066 554
rect 4075 525 4088 554
rect 4103 541 4133 554
rect 4176 541 4219 554
rect 4143 527 4158 539
rect 4177 527 4190 541
rect 4226 540 4446 554
rect 4453 541 4483 554
rect 4258 537 4411 540
rect 4140 525 4162 527
rect 4240 525 4432 537
rect 4511 525 4524 554
rect 4539 541 4569 554
rect 4606 525 4625 554
rect 4640 541 4646 554
rect 4640 540 4654 541
rect 4640 525 4646 540
rect 4655 525 4668 554
rect 4683 541 4713 554
rect 4756 541 4799 554
rect 4723 527 4738 539
rect 4757 527 4770 541
rect 4806 540 5026 554
rect 5033 541 5063 554
rect 4838 537 4991 540
rect 4720 525 4742 527
rect 4820 525 5012 537
rect 5091 525 5104 554
rect 5119 541 5149 554
rect 5186 525 5205 554
rect 5220 525 5226 554
rect 5235 525 5248 554
rect 5263 541 5293 554
rect 5336 541 5379 554
rect 5303 527 5318 539
rect 5337 527 5350 541
rect 5386 540 5606 554
rect 5613 541 5643 554
rect 5418 537 5571 540
rect 5300 525 5322 527
rect 5400 525 5592 537
rect 5671 525 5684 554
rect 5699 541 5729 554
rect 5766 525 5785 554
rect 5800 525 5806 554
rect 5815 525 5828 554
rect 5843 541 5873 554
rect 5916 541 5959 554
rect 5883 527 5898 539
rect 5917 527 5930 541
rect 5966 540 6186 554
rect 6193 541 6223 554
rect 5998 537 6151 540
rect 5880 525 5902 527
rect 5980 525 6172 537
rect 6251 525 6264 554
rect 6279 541 6309 554
rect 6346 525 6365 554
rect 6380 525 6386 554
rect 6395 525 6408 554
rect 6423 541 6453 554
rect 6496 541 6539 554
rect 6463 527 6478 539
rect 6497 527 6510 541
rect 6546 540 6766 554
rect 6773 541 6803 554
rect 6578 537 6731 540
rect 6460 525 6482 527
rect 6560 525 6752 537
rect 6831 525 6844 554
rect 6859 541 6889 554
rect 6926 525 6945 554
rect 6960 525 6966 554
rect 6975 525 6988 554
rect 7003 541 7033 554
rect 7076 541 7119 554
rect 7043 527 7058 539
rect 7077 527 7090 541
rect 7126 540 7346 554
rect 7353 541 7383 554
rect 7158 537 7311 540
rect 7040 525 7062 527
rect 7140 525 7332 537
rect 7411 525 7424 554
rect 7439 541 7469 554
rect 7506 525 7525 554
rect 7540 525 7546 554
rect 7555 525 7568 554
rect 7583 541 7613 554
rect 7656 541 7699 554
rect 7623 527 7638 539
rect 7657 527 7670 541
rect 7706 540 7926 554
rect 7933 541 7963 554
rect 7738 537 7891 540
rect 7620 525 7642 527
rect 7720 525 7912 537
rect 7991 525 8004 554
rect 8019 541 8049 554
rect 8086 525 8105 554
rect 8120 525 8126 554
rect 8135 525 8148 554
rect 8163 541 8193 554
rect 8236 541 8279 554
rect 8203 527 8218 539
rect 8237 527 8250 541
rect 8286 540 8506 554
rect 8513 541 8543 554
rect 8318 537 8471 540
rect 8200 525 8222 527
rect 8300 525 8492 537
rect 8571 525 8584 554
rect 8599 541 8629 554
rect 8666 525 8685 554
rect 8700 525 8706 554
rect 8715 525 8728 554
rect 8743 541 8773 554
rect 8816 541 8859 554
rect 8783 527 8798 539
rect 8817 527 8830 541
rect 8866 540 9086 554
rect 9093 541 9123 554
rect 8898 537 9051 540
rect 8780 525 8802 527
rect 8880 525 9072 537
rect 9151 525 9164 554
rect 9179 541 9209 554
rect 9252 525 9265 554
rect -13 511 9265 525
rect -13 497 0 511
rect 15 441 28 511
rect 80 506 102 511
rect 73 485 102 499
rect 155 485 171 499
rect 209 495 215 497
rect 222 495 330 511
rect 337 495 343 497
rect 351 495 366 511
rect 432 505 451 508
rect 73 483 171 485
rect 198 483 366 495
rect 381 485 397 499
rect 432 486 454 505
rect 464 499 480 500
rect 463 497 480 499
rect 464 492 480 497
rect 454 485 460 486
rect 463 485 492 492
rect 381 484 492 485
rect 381 483 498 484
rect 57 475 108 483
rect 155 475 189 483
rect 57 463 82 475
rect 89 463 108 475
rect 162 473 189 475
rect 198 473 419 483
rect 454 480 460 483
rect 162 469 419 473
rect 57 455 108 463
rect 155 455 419 469
rect 463 475 498 483
rect 9 407 28 441
rect 73 447 102 455
rect 73 441 90 447
rect 73 439 107 441
rect 155 439 171 455
rect 172 445 380 455
rect 381 445 397 455
rect 445 451 460 466
rect 463 463 464 475
rect 471 463 498 475
rect 463 455 498 463
rect 463 454 492 455
rect 183 441 397 445
rect 198 439 397 441
rect 432 441 445 451
rect 463 441 480 454
rect 432 439 480 441
rect 74 435 107 439
rect 70 433 107 435
rect 70 432 137 433
rect 70 427 101 432
rect 107 427 137 432
rect 70 423 137 427
rect 43 420 137 423
rect 43 413 92 420
rect 43 407 73 413
rect 92 408 97 413
rect -13 373 0 401
rect 9 391 89 407
rect 101 399 137 420
rect 198 415 387 439
rect 432 438 479 439
rect 445 433 479 438
rect 213 412 387 415
rect 206 409 387 412
rect 415 432 479 433
rect 9 389 28 391
rect 43 389 77 391
rect 9 373 89 389
rect 9 367 28 373
rect -1 351 28 367
rect 43 357 73 373
rect 101 351 107 399
rect 110 393 129 399
rect 144 393 174 401
rect 110 385 174 393
rect 110 369 190 385
rect 206 378 268 409
rect 284 378 346 409
rect 415 407 464 432
rect 479 407 509 423
rect 378 393 408 401
rect 415 399 525 407
rect 378 385 423 393
rect 110 367 129 369
rect 144 367 190 369
rect 110 351 190 367
rect 217 365 252 378
rect 293 375 330 378
rect 293 373 335 375
rect 222 362 252 365
rect 231 358 238 362
rect 238 357 239 358
rect 197 351 207 357
rect -7 343 34 351
rect -7 317 8 343
rect 15 317 34 343
rect 98 339 129 351
rect 144 339 247 351
rect 259 341 285 367
rect 300 362 330 373
rect 362 369 424 385
rect 362 367 408 369
rect 362 351 424 367
rect 436 351 442 399
rect 445 391 525 399
rect 445 389 464 391
rect 479 389 513 391
rect 445 373 525 389
rect 445 351 464 373
rect 479 357 509 373
rect 537 367 543 441
rect 546 367 565 511
rect 580 367 586 511
rect 595 441 608 511
rect 660 506 682 511
rect 653 485 682 499
rect 735 485 751 499
rect 789 495 795 497
rect 802 495 910 511
rect 917 495 923 497
rect 931 495 946 511
rect 1012 505 1031 508
rect 653 483 751 485
rect 778 483 946 495
rect 961 485 977 499
rect 1012 486 1034 505
rect 1044 499 1060 500
rect 1043 497 1060 499
rect 1044 492 1060 497
rect 1034 485 1040 486
rect 1043 485 1072 492
rect 961 484 1072 485
rect 961 483 1078 484
rect 637 475 688 483
rect 735 475 769 483
rect 637 463 662 475
rect 669 463 688 475
rect 742 473 769 475
rect 778 473 999 483
rect 1034 480 1040 483
rect 742 469 999 473
rect 637 455 688 463
rect 735 455 999 469
rect 1043 475 1078 483
rect 589 407 608 441
rect 653 447 682 455
rect 653 441 670 447
rect 653 439 687 441
rect 735 439 751 455
rect 752 445 960 455
rect 961 445 977 455
rect 1025 451 1040 466
rect 1043 463 1044 475
rect 1051 463 1078 475
rect 1043 455 1078 463
rect 1043 454 1072 455
rect 763 441 977 445
rect 778 439 977 441
rect 1012 441 1025 451
rect 1043 441 1060 454
rect 1012 439 1060 441
rect 654 435 687 439
rect 650 433 687 435
rect 650 432 717 433
rect 650 427 681 432
rect 687 427 717 432
rect 650 423 717 427
rect 623 420 717 423
rect 623 413 672 420
rect 623 407 653 413
rect 672 408 677 413
rect 589 391 669 407
rect 681 399 717 420
rect 778 415 967 439
rect 1012 438 1059 439
rect 1025 433 1059 438
rect 793 412 967 415
rect 786 409 967 412
rect 995 432 1059 433
rect 589 389 608 391
rect 623 389 657 391
rect 589 373 669 389
rect 589 367 608 373
rect 305 341 408 351
rect 259 339 408 341
rect 429 339 464 351
rect 98 337 260 339
rect 110 317 129 337
rect 144 335 174 337
rect -7 309 34 317
rect 116 313 129 317
rect 181 321 260 337
rect 292 337 464 339
rect 292 321 371 337
rect 378 335 408 337
rect -1 299 28 309
rect 43 299 73 313
rect 116 299 159 313
rect 181 309 371 321
rect 436 317 442 337
rect 166 299 196 309
rect 197 299 355 309
rect 359 299 389 309
rect 393 299 423 313
rect 451 299 464 337
rect 536 351 565 367
rect 579 351 608 367
rect 623 357 653 373
rect 681 351 687 399
rect 690 393 709 399
rect 724 393 754 401
rect 690 385 754 393
rect 690 369 770 385
rect 786 378 848 409
rect 864 378 926 409
rect 995 407 1044 432
rect 1059 407 1089 423
rect 958 393 988 401
rect 995 399 1105 407
rect 958 385 1003 393
rect 690 367 709 369
rect 724 367 770 369
rect 690 351 770 367
rect 797 365 832 378
rect 873 375 910 378
rect 873 373 915 375
rect 802 362 832 365
rect 811 358 818 362
rect 818 357 819 358
rect 777 351 787 357
rect 536 343 571 351
rect 536 317 537 343
rect 544 317 571 343
rect 479 299 509 313
rect 536 309 571 317
rect 573 343 614 351
rect 573 317 588 343
rect 595 317 614 343
rect 678 339 709 351
rect 724 339 827 351
rect 839 341 865 367
rect 880 362 910 373
rect 942 369 1004 385
rect 942 367 988 369
rect 942 351 1004 367
rect 1016 351 1022 399
rect 1025 391 1105 399
rect 1025 389 1044 391
rect 1059 389 1093 391
rect 1025 373 1105 389
rect 1025 351 1044 373
rect 1059 357 1089 373
rect 1117 367 1123 441
rect 1126 367 1145 511
rect 1160 367 1166 511
rect 1175 441 1188 511
rect 1240 506 1262 511
rect 1233 485 1262 499
rect 1315 485 1331 499
rect 1369 495 1375 497
rect 1382 495 1490 511
rect 1497 495 1503 497
rect 1511 495 1526 511
rect 1592 505 1611 508
rect 1233 483 1331 485
rect 1358 483 1526 495
rect 1541 485 1557 499
rect 1592 486 1614 505
rect 1624 499 1640 500
rect 1623 497 1640 499
rect 1624 492 1640 497
rect 1614 485 1620 486
rect 1623 485 1652 492
rect 1541 484 1652 485
rect 1541 483 1658 484
rect 1217 475 1268 483
rect 1315 475 1349 483
rect 1217 463 1242 475
rect 1249 463 1268 475
rect 1322 473 1349 475
rect 1358 473 1579 483
rect 1614 480 1620 483
rect 1322 469 1579 473
rect 1217 455 1268 463
rect 1315 455 1579 469
rect 1623 475 1658 483
rect 1169 407 1188 441
rect 1233 447 1262 455
rect 1233 441 1250 447
rect 1233 439 1267 441
rect 1315 439 1331 455
rect 1332 445 1540 455
rect 1541 445 1557 455
rect 1605 451 1620 466
rect 1623 463 1624 475
rect 1631 463 1658 475
rect 1623 455 1658 463
rect 1623 454 1652 455
rect 1343 441 1557 445
rect 1358 439 1557 441
rect 1592 441 1605 451
rect 1623 441 1640 454
rect 1592 439 1640 441
rect 1234 435 1267 439
rect 1230 433 1267 435
rect 1230 432 1297 433
rect 1230 427 1261 432
rect 1267 427 1297 432
rect 1230 423 1297 427
rect 1203 420 1297 423
rect 1203 413 1252 420
rect 1203 407 1233 413
rect 1252 408 1257 413
rect 1169 391 1249 407
rect 1261 399 1297 420
rect 1358 415 1547 439
rect 1592 438 1639 439
rect 1605 433 1639 438
rect 1373 412 1547 415
rect 1366 409 1547 412
rect 1575 432 1639 433
rect 1169 389 1188 391
rect 1203 389 1237 391
rect 1169 373 1249 389
rect 1169 367 1188 373
rect 885 341 988 351
rect 839 339 988 341
rect 1009 339 1044 351
rect 678 337 840 339
rect 690 317 709 337
rect 724 335 754 337
rect 573 309 614 317
rect 696 313 709 317
rect 761 321 840 337
rect 872 337 1044 339
rect 872 321 951 337
rect 958 335 988 337
rect 536 299 565 309
rect 579 299 608 309
rect 623 299 653 313
rect 696 299 739 313
rect 761 309 951 321
rect 1016 317 1022 337
rect 746 299 776 309
rect 777 299 935 309
rect 939 299 969 309
rect 973 299 1003 313
rect 1031 299 1044 337
rect 1116 351 1145 367
rect 1159 351 1188 367
rect 1203 357 1233 373
rect 1261 351 1267 399
rect 1270 393 1289 399
rect 1304 393 1334 401
rect 1270 385 1334 393
rect 1270 369 1350 385
rect 1366 378 1428 409
rect 1444 378 1506 409
rect 1575 407 1624 432
rect 1639 407 1669 423
rect 1538 393 1568 401
rect 1575 399 1685 407
rect 1538 385 1583 393
rect 1270 367 1289 369
rect 1304 367 1350 369
rect 1270 351 1350 367
rect 1377 365 1412 378
rect 1453 375 1490 378
rect 1453 373 1495 375
rect 1382 362 1412 365
rect 1391 358 1398 362
rect 1398 357 1399 358
rect 1357 351 1367 357
rect 1116 343 1151 351
rect 1116 317 1117 343
rect 1124 317 1151 343
rect 1059 299 1089 313
rect 1116 309 1151 317
rect 1153 343 1194 351
rect 1153 317 1168 343
rect 1175 317 1194 343
rect 1258 339 1289 351
rect 1304 339 1407 351
rect 1419 341 1445 367
rect 1460 362 1490 373
rect 1522 369 1584 385
rect 1522 367 1568 369
rect 1522 351 1584 367
rect 1596 351 1602 399
rect 1605 391 1685 399
rect 1605 389 1624 391
rect 1639 389 1673 391
rect 1605 373 1685 389
rect 1605 351 1624 373
rect 1639 357 1669 373
rect 1697 367 1703 441
rect 1706 367 1725 511
rect 1740 367 1746 511
rect 1755 441 1768 511
rect 1820 506 1842 511
rect 1813 485 1842 499
rect 1895 485 1911 499
rect 1949 495 1955 497
rect 1962 495 2070 511
rect 2077 495 2083 497
rect 2091 495 2106 511
rect 2172 505 2191 508
rect 1813 483 1911 485
rect 1938 483 2106 495
rect 2121 485 2137 499
rect 2172 486 2194 505
rect 2204 499 2220 500
rect 2203 497 2220 499
rect 2204 492 2220 497
rect 2194 485 2200 486
rect 2203 485 2232 492
rect 2121 484 2232 485
rect 2121 483 2238 484
rect 1797 475 1848 483
rect 1895 475 1929 483
rect 1797 463 1822 475
rect 1829 463 1848 475
rect 1902 473 1929 475
rect 1938 473 2159 483
rect 2194 480 2200 483
rect 1902 469 2159 473
rect 1797 455 1848 463
rect 1895 455 2159 469
rect 2203 475 2238 483
rect 1749 407 1768 441
rect 1813 447 1842 455
rect 1813 441 1830 447
rect 1813 439 1847 441
rect 1895 439 1911 455
rect 1912 445 2120 455
rect 2121 445 2137 455
rect 2185 451 2200 466
rect 2203 463 2204 475
rect 2211 463 2238 475
rect 2203 455 2238 463
rect 2203 454 2232 455
rect 1923 441 2137 445
rect 1938 439 2137 441
rect 2172 441 2185 451
rect 2203 441 2220 454
rect 2172 439 2220 441
rect 1814 435 1847 439
rect 1810 433 1847 435
rect 1810 432 1877 433
rect 1810 427 1841 432
rect 1847 427 1877 432
rect 1810 423 1877 427
rect 1783 420 1877 423
rect 1783 413 1832 420
rect 1783 407 1813 413
rect 1832 408 1837 413
rect 1749 391 1829 407
rect 1841 399 1877 420
rect 1938 415 2127 439
rect 2172 438 2219 439
rect 2185 433 2219 438
rect 1953 412 2127 415
rect 1946 409 2127 412
rect 2155 432 2219 433
rect 1749 389 1768 391
rect 1783 389 1817 391
rect 1749 373 1829 389
rect 1749 367 1768 373
rect 1465 341 1568 351
rect 1419 339 1568 341
rect 1589 339 1624 351
rect 1258 337 1420 339
rect 1270 317 1289 337
rect 1304 335 1334 337
rect 1153 309 1194 317
rect 1276 313 1289 317
rect 1341 321 1420 337
rect 1452 337 1624 339
rect 1452 321 1531 337
rect 1538 335 1568 337
rect 1116 299 1145 309
rect 1159 299 1188 309
rect 1203 299 1233 313
rect 1276 299 1319 313
rect 1341 309 1531 321
rect 1596 317 1602 337
rect 1326 299 1356 309
rect 1357 299 1515 309
rect 1519 299 1549 309
rect 1553 299 1583 313
rect 1611 299 1624 337
rect 1696 351 1725 367
rect 1739 351 1768 367
rect 1783 357 1813 373
rect 1841 351 1847 399
rect 1850 393 1869 399
rect 1884 393 1914 401
rect 1850 385 1914 393
rect 1850 369 1930 385
rect 1946 378 2008 409
rect 2024 378 2086 409
rect 2155 407 2204 432
rect 2219 407 2249 423
rect 2118 393 2148 401
rect 2155 399 2265 407
rect 2118 385 2163 393
rect 1850 367 1869 369
rect 1884 367 1930 369
rect 1850 351 1930 367
rect 1957 365 1992 378
rect 2033 375 2070 378
rect 2033 373 2075 375
rect 1962 362 1992 365
rect 1971 358 1978 362
rect 1978 357 1979 358
rect 1937 351 1947 357
rect 1696 343 1731 351
rect 1696 317 1697 343
rect 1704 317 1731 343
rect 1639 299 1669 313
rect 1696 309 1731 317
rect 1733 343 1774 351
rect 1733 317 1748 343
rect 1755 317 1774 343
rect 1838 339 1869 351
rect 1884 339 1987 351
rect 1999 341 2025 367
rect 2040 362 2070 373
rect 2102 369 2164 385
rect 2102 367 2148 369
rect 2102 351 2164 367
rect 2176 351 2182 399
rect 2185 391 2265 399
rect 2185 389 2204 391
rect 2219 389 2253 391
rect 2185 373 2265 389
rect 2185 351 2204 373
rect 2219 357 2249 373
rect 2277 367 2283 441
rect 2286 367 2305 511
rect 2320 367 2326 511
rect 2335 441 2348 511
rect 2400 506 2422 511
rect 2393 485 2422 499
rect 2475 485 2491 499
rect 2529 495 2535 497
rect 2542 495 2650 511
rect 2657 495 2663 497
rect 2671 495 2686 511
rect 2752 505 2771 508
rect 2393 483 2491 485
rect 2518 483 2686 495
rect 2701 485 2717 499
rect 2752 486 2774 505
rect 2784 499 2800 500
rect 2783 497 2800 499
rect 2784 492 2800 497
rect 2774 485 2780 486
rect 2783 485 2812 492
rect 2701 484 2812 485
rect 2701 483 2818 484
rect 2377 475 2428 483
rect 2475 475 2509 483
rect 2377 463 2402 475
rect 2409 463 2428 475
rect 2482 473 2509 475
rect 2518 473 2739 483
rect 2774 480 2780 483
rect 2482 469 2739 473
rect 2377 455 2428 463
rect 2475 455 2739 469
rect 2783 475 2818 483
rect 2329 407 2348 441
rect 2393 447 2422 455
rect 2393 441 2410 447
rect 2393 439 2427 441
rect 2475 439 2491 455
rect 2492 445 2700 455
rect 2701 445 2717 455
rect 2765 451 2780 466
rect 2783 463 2784 475
rect 2791 463 2818 475
rect 2783 455 2818 463
rect 2783 454 2812 455
rect 2503 441 2717 445
rect 2518 439 2717 441
rect 2752 441 2765 451
rect 2783 441 2800 454
rect 2752 439 2800 441
rect 2394 435 2427 439
rect 2390 433 2427 435
rect 2390 432 2457 433
rect 2390 427 2421 432
rect 2427 427 2457 432
rect 2390 423 2457 427
rect 2363 420 2457 423
rect 2363 413 2412 420
rect 2363 407 2393 413
rect 2412 408 2417 413
rect 2329 391 2409 407
rect 2421 399 2457 420
rect 2518 415 2707 439
rect 2752 438 2799 439
rect 2765 433 2799 438
rect 2533 412 2707 415
rect 2526 409 2707 412
rect 2735 432 2799 433
rect 2329 389 2348 391
rect 2363 389 2397 391
rect 2329 373 2409 389
rect 2329 367 2348 373
rect 2045 341 2148 351
rect 1999 339 2148 341
rect 2169 339 2204 351
rect 1838 337 2000 339
rect 1850 317 1869 337
rect 1884 335 1914 337
rect 1733 309 1774 317
rect 1856 313 1869 317
rect 1921 321 2000 337
rect 2032 337 2204 339
rect 2032 321 2111 337
rect 2118 335 2148 337
rect 1696 299 1725 309
rect 1739 299 1768 309
rect 1783 299 1813 313
rect 1856 299 1899 313
rect 1921 309 2111 321
rect 2176 317 2182 337
rect 1906 299 1936 309
rect 1937 299 2095 309
rect 2099 299 2129 309
rect 2133 299 2163 313
rect 2191 299 2204 337
rect 2276 351 2305 367
rect 2319 351 2348 367
rect 2363 357 2393 373
rect 2421 351 2427 399
rect 2430 393 2449 399
rect 2464 393 2494 401
rect 2430 385 2494 393
rect 2430 369 2510 385
rect 2526 378 2588 409
rect 2604 378 2666 409
rect 2735 407 2784 432
rect 2799 407 2829 423
rect 2698 393 2728 401
rect 2735 399 2845 407
rect 2698 385 2743 393
rect 2430 367 2449 369
rect 2464 367 2510 369
rect 2430 351 2510 367
rect 2537 365 2572 378
rect 2613 375 2650 378
rect 2613 373 2655 375
rect 2542 362 2572 365
rect 2551 358 2558 362
rect 2558 357 2559 358
rect 2517 351 2527 357
rect 2276 343 2311 351
rect 2276 317 2277 343
rect 2284 317 2311 343
rect 2219 299 2249 313
rect 2276 309 2311 317
rect 2313 343 2354 351
rect 2313 317 2328 343
rect 2335 317 2354 343
rect 2418 339 2449 351
rect 2464 339 2567 351
rect 2579 341 2605 367
rect 2620 362 2650 373
rect 2682 369 2744 385
rect 2682 367 2728 369
rect 2682 351 2744 367
rect 2756 351 2762 399
rect 2765 391 2845 399
rect 2765 389 2784 391
rect 2799 389 2833 391
rect 2765 373 2845 389
rect 2765 351 2784 373
rect 2799 357 2829 373
rect 2857 367 2863 441
rect 2866 367 2885 511
rect 2900 367 2906 511
rect 2915 441 2928 511
rect 2980 506 3002 511
rect 2973 485 3002 499
rect 3055 485 3071 499
rect 3109 495 3115 497
rect 3122 495 3230 511
rect 3237 495 3243 497
rect 3251 495 3266 511
rect 3332 505 3351 508
rect 2973 483 3071 485
rect 3098 483 3266 495
rect 3281 485 3297 499
rect 3332 486 3354 505
rect 3364 499 3380 500
rect 3363 497 3380 499
rect 3364 492 3380 497
rect 3354 485 3360 486
rect 3363 485 3392 492
rect 3281 484 3392 485
rect 3281 483 3398 484
rect 2957 475 3008 483
rect 3055 475 3089 483
rect 2957 463 2982 475
rect 2989 463 3008 475
rect 3062 473 3089 475
rect 3098 473 3319 483
rect 3354 480 3360 483
rect 3062 469 3319 473
rect 2957 455 3008 463
rect 3055 455 3319 469
rect 3363 475 3398 483
rect 2909 407 2928 441
rect 2973 447 3002 455
rect 2973 441 2990 447
rect 2973 439 3007 441
rect 3055 439 3071 455
rect 3072 445 3280 455
rect 3281 445 3297 455
rect 3345 451 3360 466
rect 3363 463 3364 475
rect 3371 463 3398 475
rect 3363 455 3398 463
rect 3363 454 3392 455
rect 3083 441 3297 445
rect 3098 439 3297 441
rect 3332 441 3345 451
rect 3363 441 3380 454
rect 3332 439 3380 441
rect 2974 435 3007 439
rect 2970 433 3007 435
rect 2970 432 3037 433
rect 2970 427 3001 432
rect 3007 427 3037 432
rect 2970 423 3037 427
rect 2943 420 3037 423
rect 2943 413 2992 420
rect 2943 407 2973 413
rect 2992 408 2997 413
rect 2909 391 2989 407
rect 3001 399 3037 420
rect 3098 415 3287 439
rect 3332 438 3379 439
rect 3345 433 3379 438
rect 3113 412 3287 415
rect 3106 409 3287 412
rect 3315 432 3379 433
rect 2909 389 2928 391
rect 2943 389 2977 391
rect 2909 373 2989 389
rect 2909 367 2928 373
rect 2625 341 2728 351
rect 2579 339 2728 341
rect 2749 339 2784 351
rect 2418 337 2580 339
rect 2430 317 2449 337
rect 2464 335 2494 337
rect 2313 309 2354 317
rect 2436 313 2449 317
rect 2501 321 2580 337
rect 2612 337 2784 339
rect 2612 321 2691 337
rect 2698 335 2728 337
rect 2276 299 2305 309
rect 2319 299 2348 309
rect 2363 299 2393 313
rect 2436 299 2479 313
rect 2501 309 2691 321
rect 2756 317 2762 337
rect 2486 299 2516 309
rect 2517 299 2675 309
rect 2679 299 2709 309
rect 2713 299 2743 313
rect 2771 299 2784 337
rect 2856 351 2885 367
rect 2899 351 2928 367
rect 2943 357 2973 373
rect 3001 351 3007 399
rect 3010 393 3029 399
rect 3044 393 3074 401
rect 3010 385 3074 393
rect 3010 369 3090 385
rect 3106 378 3168 409
rect 3184 378 3246 409
rect 3315 407 3364 432
rect 3379 407 3409 423
rect 3278 393 3308 401
rect 3315 399 3425 407
rect 3278 385 3323 393
rect 3010 367 3029 369
rect 3044 367 3090 369
rect 3010 351 3090 367
rect 3117 365 3152 378
rect 3193 375 3230 378
rect 3193 373 3235 375
rect 3122 362 3152 365
rect 3131 358 3138 362
rect 3138 357 3139 358
rect 3097 351 3107 357
rect 2856 343 2891 351
rect 2856 317 2857 343
rect 2864 317 2891 343
rect 2799 299 2829 313
rect 2856 309 2891 317
rect 2893 343 2934 351
rect 2893 317 2908 343
rect 2915 317 2934 343
rect 2998 339 3029 351
rect 3044 339 3147 351
rect 3159 341 3185 367
rect 3200 362 3230 373
rect 3262 369 3324 385
rect 3262 367 3308 369
rect 3262 351 3324 367
rect 3336 351 3342 399
rect 3345 391 3425 399
rect 3345 389 3364 391
rect 3379 389 3413 391
rect 3345 373 3425 389
rect 3345 351 3364 373
rect 3379 357 3409 373
rect 3437 367 3443 441
rect 3446 367 3465 511
rect 3480 367 3486 511
rect 3495 441 3508 511
rect 3560 506 3582 511
rect 3553 485 3582 499
rect 3635 485 3651 499
rect 3689 495 3695 497
rect 3702 495 3810 511
rect 3817 495 3823 497
rect 3831 495 3846 511
rect 3912 505 3931 508
rect 3553 483 3651 485
rect 3678 483 3846 495
rect 3861 485 3877 499
rect 3912 486 3934 505
rect 3944 499 3960 500
rect 3943 497 3960 499
rect 3944 492 3960 497
rect 3934 485 3940 486
rect 3943 485 3972 492
rect 3861 484 3972 485
rect 3861 483 3978 484
rect 3537 475 3588 483
rect 3635 475 3669 483
rect 3537 463 3562 475
rect 3569 463 3588 475
rect 3642 473 3669 475
rect 3678 473 3899 483
rect 3934 480 3940 483
rect 3642 469 3899 473
rect 3537 455 3588 463
rect 3635 455 3899 469
rect 3943 475 3978 483
rect 3489 407 3508 441
rect 3553 447 3582 455
rect 3553 441 3570 447
rect 3553 439 3587 441
rect 3635 439 3651 455
rect 3652 445 3860 455
rect 3861 445 3877 455
rect 3925 451 3940 466
rect 3943 463 3944 475
rect 3951 463 3978 475
rect 3943 455 3978 463
rect 3943 454 3972 455
rect 3663 441 3877 445
rect 3678 439 3877 441
rect 3912 441 3925 451
rect 3943 441 3960 454
rect 3912 439 3960 441
rect 3554 435 3587 439
rect 3550 433 3587 435
rect 3550 432 3617 433
rect 3550 427 3581 432
rect 3587 427 3617 432
rect 3550 423 3617 427
rect 3523 420 3617 423
rect 3523 413 3572 420
rect 3523 407 3553 413
rect 3572 408 3577 413
rect 3489 391 3569 407
rect 3581 399 3617 420
rect 3678 415 3867 439
rect 3912 438 3959 439
rect 3925 433 3959 438
rect 3693 412 3867 415
rect 3686 409 3867 412
rect 3895 432 3959 433
rect 3489 389 3508 391
rect 3523 389 3557 391
rect 3489 373 3569 389
rect 3489 367 3508 373
rect 3205 341 3308 351
rect 3159 339 3308 341
rect 3329 339 3364 351
rect 2998 337 3160 339
rect 3010 317 3029 337
rect 3044 335 3074 337
rect 2893 309 2934 317
rect 3016 313 3029 317
rect 3081 321 3160 337
rect 3192 337 3364 339
rect 3192 321 3271 337
rect 3278 335 3308 337
rect 2856 299 2885 309
rect 2899 299 2928 309
rect 2943 299 2973 313
rect 3016 299 3059 313
rect 3081 309 3271 321
rect 3336 317 3342 337
rect 3066 299 3096 309
rect 3097 299 3255 309
rect 3259 299 3289 309
rect 3293 299 3323 313
rect 3351 299 3364 337
rect 3436 351 3465 367
rect 3479 351 3508 367
rect 3523 357 3553 373
rect 3581 351 3587 399
rect 3590 393 3609 399
rect 3624 393 3654 401
rect 3590 385 3654 393
rect 3590 369 3670 385
rect 3686 378 3748 409
rect 3764 378 3826 409
rect 3895 407 3944 432
rect 3959 407 3989 423
rect 3858 393 3888 401
rect 3895 399 4005 407
rect 3858 385 3903 393
rect 3590 367 3609 369
rect 3624 367 3670 369
rect 3590 351 3670 367
rect 3697 365 3732 378
rect 3773 375 3810 378
rect 3773 373 3815 375
rect 3702 362 3732 365
rect 3711 358 3718 362
rect 3718 357 3719 358
rect 3677 351 3687 357
rect 3436 343 3471 351
rect 3436 317 3437 343
rect 3444 317 3471 343
rect 3379 299 3409 313
rect 3436 309 3471 317
rect 3473 343 3514 351
rect 3473 317 3488 343
rect 3495 317 3514 343
rect 3578 339 3609 351
rect 3624 339 3727 351
rect 3739 341 3765 367
rect 3780 362 3810 373
rect 3842 369 3904 385
rect 3842 367 3888 369
rect 3842 351 3904 367
rect 3916 351 3922 399
rect 3925 391 4005 399
rect 3925 389 3944 391
rect 3959 389 3993 391
rect 3925 373 4005 389
rect 3925 351 3944 373
rect 3959 357 3989 373
rect 4017 367 4023 441
rect 4026 367 4045 511
rect 4060 367 4066 511
rect 4075 441 4088 511
rect 4140 506 4162 511
rect 4133 485 4162 499
rect 4215 485 4231 499
rect 4269 495 4275 497
rect 4282 495 4390 511
rect 4397 495 4403 497
rect 4411 495 4426 511
rect 4606 510 4646 511
rect 4492 505 4511 508
rect 4133 483 4231 485
rect 4258 483 4426 495
rect 4441 485 4457 499
rect 4492 486 4514 505
rect 4524 499 4540 500
rect 4523 497 4540 499
rect 4524 492 4540 497
rect 4514 485 4520 486
rect 4523 485 4552 492
rect 4441 484 4552 485
rect 4441 483 4558 484
rect 4117 475 4168 483
rect 4215 475 4249 483
rect 4117 463 4142 475
rect 4149 463 4168 475
rect 4222 473 4249 475
rect 4258 473 4479 483
rect 4514 480 4520 483
rect 4222 469 4479 473
rect 4117 455 4168 463
rect 4215 455 4479 469
rect 4523 475 4558 483
rect 4069 407 4088 441
rect 4133 447 4162 455
rect 4133 441 4150 447
rect 4133 439 4167 441
rect 4215 439 4231 455
rect 4232 445 4440 455
rect 4441 445 4457 455
rect 4505 451 4520 466
rect 4523 463 4524 475
rect 4531 463 4558 475
rect 4523 455 4558 463
rect 4523 454 4552 455
rect 4243 441 4457 445
rect 4258 439 4457 441
rect 4492 441 4505 451
rect 4523 441 4540 454
rect 4492 439 4540 441
rect 4134 435 4167 439
rect 4130 433 4167 435
rect 4130 432 4197 433
rect 4130 427 4161 432
rect 4167 427 4197 432
rect 4130 423 4197 427
rect 4103 420 4197 423
rect 4103 413 4152 420
rect 4103 407 4133 413
rect 4152 408 4157 413
rect 4069 391 4149 407
rect 4161 399 4197 420
rect 4258 415 4447 439
rect 4492 438 4539 439
rect 4505 433 4539 438
rect 4273 412 4447 415
rect 4266 409 4447 412
rect 4475 432 4539 433
rect 4069 389 4088 391
rect 4103 389 4137 391
rect 4069 373 4149 389
rect 4069 367 4088 373
rect 3785 341 3888 351
rect 3739 339 3888 341
rect 3909 339 3944 351
rect 3578 337 3740 339
rect 3590 317 3609 337
rect 3624 335 3654 337
rect 3473 309 3514 317
rect 3596 313 3609 317
rect 3661 321 3740 337
rect 3772 337 3944 339
rect 3772 321 3851 337
rect 3858 335 3888 337
rect 3436 299 3465 309
rect 3479 299 3508 309
rect 3523 299 3553 313
rect 3596 299 3639 313
rect 3661 309 3851 321
rect 3916 317 3922 337
rect 3646 299 3676 309
rect 3677 299 3835 309
rect 3839 299 3869 309
rect 3873 299 3903 313
rect 3931 299 3944 337
rect 4016 351 4045 367
rect 4059 351 4088 367
rect 4103 357 4133 373
rect 4161 351 4167 399
rect 4170 393 4189 399
rect 4204 393 4234 401
rect 4170 385 4234 393
rect 4170 369 4250 385
rect 4266 378 4328 409
rect 4344 378 4406 409
rect 4475 407 4524 432
rect 4539 407 4569 423
rect 4438 393 4468 401
rect 4475 399 4585 407
rect 4438 385 4483 393
rect 4170 367 4189 369
rect 4204 367 4250 369
rect 4170 351 4250 367
rect 4277 365 4312 378
rect 4353 375 4390 378
rect 4353 373 4395 375
rect 4282 362 4312 365
rect 4291 358 4298 362
rect 4298 357 4299 358
rect 4257 351 4267 357
rect 4016 343 4051 351
rect 4016 317 4017 343
rect 4024 317 4051 343
rect 3959 299 3989 313
rect 4016 309 4051 317
rect 4053 343 4094 351
rect 4053 317 4068 343
rect 4075 317 4094 343
rect 4158 339 4189 351
rect 4204 339 4307 351
rect 4319 341 4345 367
rect 4360 362 4390 373
rect 4422 369 4484 385
rect 4422 367 4468 369
rect 4422 351 4484 367
rect 4496 351 4502 399
rect 4505 391 4585 399
rect 4505 389 4524 391
rect 4539 389 4573 391
rect 4505 373 4585 389
rect 4505 351 4524 373
rect 4539 357 4569 373
rect 4597 367 4603 441
rect 4606 367 4625 510
rect 4640 367 4646 510
rect 4655 441 4668 511
rect 4720 506 4742 511
rect 4713 485 4742 499
rect 4795 485 4811 499
rect 4849 495 4855 497
rect 4862 495 4970 511
rect 4977 495 4983 497
rect 4991 495 5006 511
rect 5072 505 5091 508
rect 4713 483 4811 485
rect 4838 483 5006 495
rect 5021 485 5037 499
rect 5072 486 5094 505
rect 5104 499 5120 500
rect 5103 497 5120 499
rect 5104 492 5120 497
rect 5094 485 5100 486
rect 5103 485 5132 492
rect 5021 484 5132 485
rect 5021 483 5138 484
rect 4697 475 4748 483
rect 4795 475 4829 483
rect 4697 463 4722 475
rect 4729 463 4748 475
rect 4802 473 4829 475
rect 4838 473 5059 483
rect 5094 480 5100 483
rect 4802 469 5059 473
rect 4697 455 4748 463
rect 4795 455 5059 469
rect 5103 475 5138 483
rect 4649 407 4668 441
rect 4713 447 4742 455
rect 4713 441 4730 447
rect 4713 439 4747 441
rect 4795 439 4811 455
rect 4812 445 5020 455
rect 5021 445 5037 455
rect 5085 451 5100 466
rect 5103 463 5104 475
rect 5111 463 5138 475
rect 5103 455 5138 463
rect 5103 454 5132 455
rect 4823 441 5037 445
rect 4838 439 5037 441
rect 5072 441 5085 451
rect 5103 441 5120 454
rect 5072 439 5120 441
rect 4714 435 4747 439
rect 4710 433 4747 435
rect 4710 432 4777 433
rect 4710 427 4741 432
rect 4747 427 4777 432
rect 4710 423 4777 427
rect 4683 420 4777 423
rect 4683 413 4732 420
rect 4683 407 4713 413
rect 4732 408 4737 413
rect 4649 391 4729 407
rect 4741 399 4777 420
rect 4838 415 5027 439
rect 5072 438 5119 439
rect 5085 433 5119 438
rect 4853 412 5027 415
rect 4846 409 5027 412
rect 5055 432 5119 433
rect 4649 389 4668 391
rect 4683 389 4717 391
rect 4649 373 4729 389
rect 4649 367 4668 373
rect 4365 341 4468 351
rect 4319 339 4468 341
rect 4489 339 4524 351
rect 4158 337 4320 339
rect 4170 317 4189 337
rect 4204 335 4234 337
rect 4053 309 4094 317
rect 4176 313 4189 317
rect 4241 321 4320 337
rect 4352 337 4524 339
rect 4352 321 4431 337
rect 4438 335 4468 337
rect 4016 299 4045 309
rect 4059 299 4088 309
rect 4103 299 4133 313
rect 4176 299 4219 313
rect 4241 309 4431 321
rect 4496 317 4502 337
rect 4226 299 4256 309
rect 4257 299 4415 309
rect 4419 299 4449 309
rect 4453 299 4483 313
rect 4511 299 4524 337
rect 4596 351 4625 367
rect 4639 351 4668 367
rect 4683 357 4713 373
rect 4741 351 4747 399
rect 4750 393 4769 399
rect 4784 393 4814 401
rect 4750 385 4814 393
rect 4750 369 4830 385
rect 4846 378 4908 409
rect 4924 378 4986 409
rect 5055 407 5104 432
rect 5119 407 5149 423
rect 5018 393 5048 401
rect 5055 399 5165 407
rect 5018 385 5063 393
rect 4750 367 4769 369
rect 4784 367 4830 369
rect 4750 351 4830 367
rect 4857 365 4892 378
rect 4933 375 4970 378
rect 4933 373 4975 375
rect 4862 362 4892 365
rect 4871 358 4878 362
rect 4878 357 4879 358
rect 4837 351 4847 357
rect 4596 343 4631 351
rect 4596 317 4597 343
rect 4604 317 4631 343
rect 4539 299 4569 313
rect 4596 309 4631 317
rect 4633 343 4674 351
rect 4633 317 4648 343
rect 4655 317 4674 343
rect 4738 339 4769 351
rect 4784 339 4887 351
rect 4899 341 4925 367
rect 4940 362 4970 373
rect 5002 369 5064 385
rect 5002 367 5048 369
rect 5002 351 5064 367
rect 5076 351 5082 399
rect 5085 391 5165 399
rect 5085 389 5104 391
rect 5119 389 5153 391
rect 5085 373 5165 389
rect 5085 351 5104 373
rect 5119 357 5149 373
rect 5177 367 5183 441
rect 5186 367 5205 511
rect 5220 367 5226 511
rect 5235 441 5248 511
rect 5300 506 5322 511
rect 5293 485 5322 499
rect 5375 485 5391 499
rect 5429 495 5435 497
rect 5442 495 5550 511
rect 5557 495 5563 497
rect 5571 495 5586 511
rect 5652 505 5671 508
rect 5293 483 5391 485
rect 5418 483 5586 495
rect 5601 485 5617 499
rect 5652 486 5674 505
rect 5684 499 5700 500
rect 5683 497 5700 499
rect 5684 492 5700 497
rect 5674 485 5680 486
rect 5683 485 5712 492
rect 5601 484 5712 485
rect 5601 483 5718 484
rect 5277 475 5328 483
rect 5375 475 5409 483
rect 5277 463 5302 475
rect 5309 463 5328 475
rect 5382 473 5409 475
rect 5418 473 5639 483
rect 5674 480 5680 483
rect 5382 469 5639 473
rect 5277 455 5328 463
rect 5375 455 5639 469
rect 5683 475 5718 483
rect 5229 407 5248 441
rect 5293 447 5322 455
rect 5293 441 5310 447
rect 5293 439 5327 441
rect 5375 439 5391 455
rect 5392 445 5600 455
rect 5601 445 5617 455
rect 5665 451 5680 466
rect 5683 463 5684 475
rect 5691 463 5718 475
rect 5683 455 5718 463
rect 5683 454 5712 455
rect 5403 441 5617 445
rect 5418 439 5617 441
rect 5652 441 5665 451
rect 5683 441 5700 454
rect 5652 439 5700 441
rect 5294 435 5327 439
rect 5290 433 5327 435
rect 5290 432 5357 433
rect 5290 427 5321 432
rect 5327 427 5357 432
rect 5290 423 5357 427
rect 5263 420 5357 423
rect 5263 413 5312 420
rect 5263 407 5293 413
rect 5312 408 5317 413
rect 5229 391 5309 407
rect 5321 399 5357 420
rect 5418 415 5607 439
rect 5652 438 5699 439
rect 5665 433 5699 438
rect 5433 412 5607 415
rect 5426 409 5607 412
rect 5635 432 5699 433
rect 5229 389 5248 391
rect 5263 389 5297 391
rect 5229 373 5309 389
rect 5229 367 5248 373
rect 4945 341 5048 351
rect 4899 339 5048 341
rect 5069 339 5104 351
rect 4738 337 4900 339
rect 4750 317 4769 337
rect 4784 335 4814 337
rect 4633 309 4674 317
rect 4756 313 4769 317
rect 4821 321 4900 337
rect 4932 337 5104 339
rect 4932 321 5011 337
rect 5018 335 5048 337
rect 4596 299 4625 309
rect 4639 299 4668 309
rect 4683 299 4713 313
rect 4756 299 4799 313
rect 4821 309 5011 321
rect 5076 317 5082 337
rect 4806 299 4836 309
rect 4837 299 4995 309
rect 4999 299 5029 309
rect 5033 299 5063 313
rect 5091 299 5104 337
rect 5176 351 5205 367
rect 5219 351 5248 367
rect 5263 357 5293 373
rect 5321 351 5327 399
rect 5330 393 5349 399
rect 5364 393 5394 401
rect 5330 385 5394 393
rect 5330 369 5410 385
rect 5426 378 5488 409
rect 5504 378 5566 409
rect 5635 407 5684 432
rect 5699 407 5729 423
rect 5598 393 5628 401
rect 5635 399 5745 407
rect 5598 385 5643 393
rect 5330 367 5349 369
rect 5364 367 5410 369
rect 5330 351 5410 367
rect 5437 365 5472 378
rect 5513 375 5550 378
rect 5513 373 5555 375
rect 5442 362 5472 365
rect 5451 358 5458 362
rect 5458 357 5459 358
rect 5417 351 5427 357
rect 5176 343 5211 351
rect 5176 317 5177 343
rect 5184 317 5211 343
rect 5119 299 5149 313
rect 5176 309 5211 317
rect 5213 343 5254 351
rect 5213 317 5228 343
rect 5235 317 5254 343
rect 5318 339 5349 351
rect 5364 339 5467 351
rect 5479 341 5505 367
rect 5520 362 5550 373
rect 5582 369 5644 385
rect 5582 367 5628 369
rect 5582 351 5644 367
rect 5656 351 5662 399
rect 5665 391 5745 399
rect 5665 389 5684 391
rect 5699 389 5733 391
rect 5665 373 5745 389
rect 5665 351 5684 373
rect 5699 357 5729 373
rect 5757 367 5763 441
rect 5766 367 5785 511
rect 5800 367 5806 511
rect 5815 441 5828 511
rect 5880 506 5902 511
rect 5873 485 5902 499
rect 5955 485 5971 499
rect 6009 495 6015 497
rect 6022 495 6130 511
rect 6137 495 6143 497
rect 6151 495 6166 511
rect 6232 505 6251 508
rect 5873 483 5971 485
rect 5998 483 6166 495
rect 6181 485 6197 499
rect 6232 486 6254 505
rect 6264 499 6280 500
rect 6263 497 6280 499
rect 6264 492 6280 497
rect 6254 485 6260 486
rect 6263 485 6292 492
rect 6181 484 6292 485
rect 6181 483 6298 484
rect 5857 475 5908 483
rect 5955 475 5989 483
rect 5857 463 5882 475
rect 5889 463 5908 475
rect 5962 473 5989 475
rect 5998 473 6219 483
rect 6254 480 6260 483
rect 5962 469 6219 473
rect 5857 455 5908 463
rect 5955 455 6219 469
rect 6263 475 6298 483
rect 5809 407 5828 441
rect 5873 447 5902 455
rect 5873 441 5890 447
rect 5873 439 5907 441
rect 5955 439 5971 455
rect 5972 445 6180 455
rect 6181 445 6197 455
rect 6245 451 6260 466
rect 6263 463 6264 475
rect 6271 463 6298 475
rect 6263 455 6298 463
rect 6263 454 6292 455
rect 5983 441 6197 445
rect 5998 439 6197 441
rect 6232 441 6245 451
rect 6263 441 6280 454
rect 6232 439 6280 441
rect 5874 435 5907 439
rect 5870 433 5907 435
rect 5870 432 5937 433
rect 5870 427 5901 432
rect 5907 427 5937 432
rect 5870 423 5937 427
rect 5843 420 5937 423
rect 5843 413 5892 420
rect 5843 407 5873 413
rect 5892 408 5897 413
rect 5809 391 5889 407
rect 5901 399 5937 420
rect 5998 415 6187 439
rect 6232 438 6279 439
rect 6245 433 6279 438
rect 6013 412 6187 415
rect 6006 409 6187 412
rect 6215 432 6279 433
rect 5809 389 5828 391
rect 5843 389 5877 391
rect 5809 373 5889 389
rect 5809 367 5828 373
rect 5525 341 5628 351
rect 5479 339 5628 341
rect 5649 339 5684 351
rect 5318 337 5480 339
rect 5330 317 5349 337
rect 5364 335 5394 337
rect 5213 309 5254 317
rect 5336 313 5349 317
rect 5401 321 5480 337
rect 5512 337 5684 339
rect 5512 321 5591 337
rect 5598 335 5628 337
rect 5176 299 5205 309
rect 5219 299 5248 309
rect 5263 299 5293 313
rect 5336 299 5379 313
rect 5401 309 5591 321
rect 5656 317 5662 337
rect 5386 299 5416 309
rect 5417 299 5575 309
rect 5579 299 5609 309
rect 5613 299 5643 313
rect 5671 299 5684 337
rect 5756 351 5785 367
rect 5799 351 5828 367
rect 5843 357 5873 373
rect 5901 351 5907 399
rect 5910 393 5929 399
rect 5944 393 5974 401
rect 5910 385 5974 393
rect 5910 369 5990 385
rect 6006 378 6068 409
rect 6084 378 6146 409
rect 6215 407 6264 432
rect 6279 407 6309 423
rect 6178 393 6208 401
rect 6215 399 6325 407
rect 6178 385 6223 393
rect 5910 367 5929 369
rect 5944 367 5990 369
rect 5910 351 5990 367
rect 6017 365 6052 378
rect 6093 375 6130 378
rect 6093 373 6135 375
rect 6022 362 6052 365
rect 6031 358 6038 362
rect 6038 357 6039 358
rect 5997 351 6007 357
rect 5756 343 5791 351
rect 5756 317 5757 343
rect 5764 317 5791 343
rect 5699 299 5729 313
rect 5756 309 5791 317
rect 5793 343 5834 351
rect 5793 317 5808 343
rect 5815 317 5834 343
rect 5898 339 5929 351
rect 5944 339 6047 351
rect 6059 341 6085 367
rect 6100 362 6130 373
rect 6162 369 6224 385
rect 6162 367 6208 369
rect 6162 351 6224 367
rect 6236 351 6242 399
rect 6245 391 6325 399
rect 6245 389 6264 391
rect 6279 389 6313 391
rect 6245 373 6325 389
rect 6245 351 6264 373
rect 6279 357 6309 373
rect 6337 367 6343 441
rect 6346 367 6365 511
rect 6380 367 6386 511
rect 6395 441 6408 511
rect 6460 506 6482 511
rect 6453 485 6482 499
rect 6535 485 6551 499
rect 6589 495 6595 497
rect 6602 495 6710 511
rect 6717 495 6723 497
rect 6731 495 6746 511
rect 6812 505 6831 508
rect 6453 483 6551 485
rect 6578 483 6746 495
rect 6761 485 6777 499
rect 6812 486 6834 505
rect 6844 499 6860 500
rect 6843 497 6860 499
rect 6844 492 6860 497
rect 6834 485 6840 486
rect 6843 485 6872 492
rect 6761 484 6872 485
rect 6761 483 6878 484
rect 6437 475 6488 483
rect 6535 475 6569 483
rect 6437 463 6462 475
rect 6469 463 6488 475
rect 6542 473 6569 475
rect 6578 473 6799 483
rect 6834 480 6840 483
rect 6542 469 6799 473
rect 6437 455 6488 463
rect 6535 455 6799 469
rect 6843 475 6878 483
rect 6389 407 6408 441
rect 6453 447 6482 455
rect 6453 441 6470 447
rect 6453 439 6487 441
rect 6535 439 6551 455
rect 6552 445 6760 455
rect 6761 445 6777 455
rect 6825 451 6840 466
rect 6843 463 6844 475
rect 6851 463 6878 475
rect 6843 455 6878 463
rect 6843 454 6872 455
rect 6563 441 6777 445
rect 6578 439 6777 441
rect 6812 441 6825 451
rect 6843 441 6860 454
rect 6812 439 6860 441
rect 6454 435 6487 439
rect 6450 433 6487 435
rect 6450 432 6517 433
rect 6450 427 6481 432
rect 6487 427 6517 432
rect 6450 423 6517 427
rect 6423 420 6517 423
rect 6423 413 6472 420
rect 6423 407 6453 413
rect 6472 408 6477 413
rect 6389 391 6469 407
rect 6481 399 6517 420
rect 6578 415 6767 439
rect 6812 438 6859 439
rect 6825 433 6859 438
rect 6593 412 6767 415
rect 6586 409 6767 412
rect 6795 432 6859 433
rect 6389 389 6408 391
rect 6423 389 6457 391
rect 6389 373 6469 389
rect 6389 367 6408 373
rect 6105 341 6208 351
rect 6059 339 6208 341
rect 6229 339 6264 351
rect 5898 337 6060 339
rect 5910 317 5929 337
rect 5944 335 5974 337
rect 5793 309 5834 317
rect 5916 313 5929 317
rect 5981 321 6060 337
rect 6092 337 6264 339
rect 6092 321 6171 337
rect 6178 335 6208 337
rect 5756 299 5785 309
rect 5799 299 5828 309
rect 5843 299 5873 313
rect 5916 299 5959 313
rect 5981 309 6171 321
rect 6236 317 6242 337
rect 5966 299 5996 309
rect 5997 299 6155 309
rect 6159 299 6189 309
rect 6193 299 6223 313
rect 6251 299 6264 337
rect 6336 351 6365 367
rect 6379 351 6408 367
rect 6423 357 6453 373
rect 6481 351 6487 399
rect 6490 393 6509 399
rect 6524 393 6554 401
rect 6490 385 6554 393
rect 6490 369 6570 385
rect 6586 378 6648 409
rect 6664 378 6726 409
rect 6795 407 6844 432
rect 6859 407 6889 423
rect 6758 393 6788 401
rect 6795 399 6905 407
rect 6758 385 6803 393
rect 6490 367 6509 369
rect 6524 367 6570 369
rect 6490 351 6570 367
rect 6597 365 6632 378
rect 6673 375 6710 378
rect 6673 373 6715 375
rect 6602 362 6632 365
rect 6611 358 6618 362
rect 6618 357 6619 358
rect 6577 351 6587 357
rect 6336 343 6371 351
rect 6336 317 6337 343
rect 6344 317 6371 343
rect 6279 299 6309 313
rect 6336 309 6371 317
rect 6373 343 6414 351
rect 6373 317 6388 343
rect 6395 317 6414 343
rect 6478 339 6509 351
rect 6524 339 6627 351
rect 6639 341 6665 367
rect 6680 362 6710 373
rect 6742 369 6804 385
rect 6742 367 6788 369
rect 6742 351 6804 367
rect 6816 351 6822 399
rect 6825 391 6905 399
rect 6825 389 6844 391
rect 6859 389 6893 391
rect 6825 373 6905 389
rect 6825 351 6844 373
rect 6859 357 6889 373
rect 6917 367 6923 441
rect 6926 367 6945 511
rect 6960 367 6966 511
rect 6975 441 6988 511
rect 7040 506 7062 511
rect 7033 485 7062 499
rect 7115 485 7131 499
rect 7169 495 7175 497
rect 7182 495 7290 511
rect 7297 495 7303 497
rect 7311 495 7326 511
rect 7392 505 7411 508
rect 7033 483 7131 485
rect 7158 483 7326 495
rect 7341 485 7357 499
rect 7392 486 7414 505
rect 7424 499 7440 500
rect 7423 497 7440 499
rect 7424 492 7440 497
rect 7414 485 7420 486
rect 7423 485 7452 492
rect 7341 484 7452 485
rect 7341 483 7458 484
rect 7017 475 7068 483
rect 7115 475 7149 483
rect 7017 463 7042 475
rect 7049 463 7068 475
rect 7122 473 7149 475
rect 7158 473 7379 483
rect 7414 480 7420 483
rect 7122 469 7379 473
rect 7017 455 7068 463
rect 7115 455 7379 469
rect 7423 475 7458 483
rect 6969 407 6988 441
rect 7033 447 7062 455
rect 7033 441 7050 447
rect 7033 439 7067 441
rect 7115 439 7131 455
rect 7132 445 7340 455
rect 7341 445 7357 455
rect 7405 451 7420 466
rect 7423 463 7424 475
rect 7431 463 7458 475
rect 7423 455 7458 463
rect 7423 454 7452 455
rect 7143 441 7357 445
rect 7158 439 7357 441
rect 7392 441 7405 451
rect 7423 441 7440 454
rect 7392 439 7440 441
rect 7034 435 7067 439
rect 7030 433 7067 435
rect 7030 432 7097 433
rect 7030 427 7061 432
rect 7067 427 7097 432
rect 7030 423 7097 427
rect 7003 420 7097 423
rect 7003 413 7052 420
rect 7003 407 7033 413
rect 7052 408 7057 413
rect 6969 391 7049 407
rect 7061 399 7097 420
rect 7158 415 7347 439
rect 7392 438 7439 439
rect 7405 433 7439 438
rect 7173 412 7347 415
rect 7166 409 7347 412
rect 7375 432 7439 433
rect 6969 389 6988 391
rect 7003 389 7037 391
rect 6969 373 7049 389
rect 6969 367 6988 373
rect 6685 341 6788 351
rect 6639 339 6788 341
rect 6809 339 6844 351
rect 6478 337 6640 339
rect 6490 317 6509 337
rect 6524 335 6554 337
rect 6373 309 6414 317
rect 6496 313 6509 317
rect 6561 321 6640 337
rect 6672 337 6844 339
rect 6672 321 6751 337
rect 6758 335 6788 337
rect 6336 299 6365 309
rect 6379 299 6408 309
rect 6423 299 6453 313
rect 6496 299 6539 313
rect 6561 309 6751 321
rect 6816 317 6822 337
rect 6546 299 6576 309
rect 6577 299 6735 309
rect 6739 299 6769 309
rect 6773 299 6803 313
rect 6831 299 6844 337
rect 6916 351 6945 367
rect 6959 351 6988 367
rect 7003 357 7033 373
rect 7061 351 7067 399
rect 7070 393 7089 399
rect 7104 393 7134 401
rect 7070 385 7134 393
rect 7070 369 7150 385
rect 7166 378 7228 409
rect 7244 378 7306 409
rect 7375 407 7424 432
rect 7439 407 7469 423
rect 7338 393 7368 401
rect 7375 399 7485 407
rect 7338 385 7383 393
rect 7070 367 7089 369
rect 7104 367 7150 369
rect 7070 351 7150 367
rect 7177 365 7212 378
rect 7253 375 7290 378
rect 7253 373 7295 375
rect 7182 362 7212 365
rect 7191 358 7198 362
rect 7198 357 7199 358
rect 7157 351 7167 357
rect 6916 343 6951 351
rect 6916 317 6917 343
rect 6924 317 6951 343
rect 6859 299 6889 313
rect 6916 309 6951 317
rect 6953 343 6994 351
rect 6953 317 6968 343
rect 6975 317 6994 343
rect 7058 339 7089 351
rect 7104 339 7207 351
rect 7219 341 7245 367
rect 7260 362 7290 373
rect 7322 369 7384 385
rect 7322 367 7368 369
rect 7322 351 7384 367
rect 7396 351 7402 399
rect 7405 391 7485 399
rect 7405 389 7424 391
rect 7439 389 7473 391
rect 7405 373 7485 389
rect 7405 351 7424 373
rect 7439 357 7469 373
rect 7497 367 7503 441
rect 7506 367 7525 511
rect 7540 367 7546 511
rect 7555 441 7568 511
rect 7620 506 7642 511
rect 7613 485 7642 499
rect 7695 485 7711 499
rect 7749 495 7755 497
rect 7762 495 7870 511
rect 7877 495 7883 497
rect 7891 495 7906 511
rect 7972 505 7991 508
rect 7613 483 7711 485
rect 7738 483 7906 495
rect 7921 485 7937 499
rect 7972 486 7994 505
rect 8004 499 8020 500
rect 8003 497 8020 499
rect 8004 492 8020 497
rect 7994 485 8000 486
rect 8003 485 8032 492
rect 7921 484 8032 485
rect 7921 483 8038 484
rect 7597 475 7648 483
rect 7695 475 7729 483
rect 7597 463 7622 475
rect 7629 463 7648 475
rect 7702 473 7729 475
rect 7738 473 7959 483
rect 7994 480 8000 483
rect 7702 469 7959 473
rect 7597 455 7648 463
rect 7695 455 7959 469
rect 8003 475 8038 483
rect 7549 407 7568 441
rect 7613 447 7642 455
rect 7613 441 7630 447
rect 7613 439 7647 441
rect 7695 439 7711 455
rect 7712 445 7920 455
rect 7921 445 7937 455
rect 7985 451 8000 466
rect 8003 463 8004 475
rect 8011 463 8038 475
rect 8003 455 8038 463
rect 8003 454 8032 455
rect 7723 441 7937 445
rect 7738 439 7937 441
rect 7972 441 7985 451
rect 8003 441 8020 454
rect 7972 439 8020 441
rect 7614 435 7647 439
rect 7610 433 7647 435
rect 7610 432 7677 433
rect 7610 427 7641 432
rect 7647 427 7677 432
rect 7610 423 7677 427
rect 7583 420 7677 423
rect 7583 413 7632 420
rect 7583 407 7613 413
rect 7632 408 7637 413
rect 7549 391 7629 407
rect 7641 399 7677 420
rect 7738 415 7927 439
rect 7972 438 8019 439
rect 7985 433 8019 438
rect 7753 412 7927 415
rect 7746 409 7927 412
rect 7955 432 8019 433
rect 7549 389 7568 391
rect 7583 389 7617 391
rect 7549 373 7629 389
rect 7549 367 7568 373
rect 7265 341 7368 351
rect 7219 339 7368 341
rect 7389 339 7424 351
rect 7058 337 7220 339
rect 7070 317 7089 337
rect 7104 335 7134 337
rect 6953 309 6994 317
rect 7076 313 7089 317
rect 7141 321 7220 337
rect 7252 337 7424 339
rect 7252 321 7331 337
rect 7338 335 7368 337
rect 6916 299 6945 309
rect 6959 299 6988 309
rect 7003 299 7033 313
rect 7076 299 7119 313
rect 7141 309 7331 321
rect 7396 317 7402 337
rect 7126 299 7156 309
rect 7157 299 7315 309
rect 7319 299 7349 309
rect 7353 299 7383 313
rect 7411 299 7424 337
rect 7496 351 7525 367
rect 7539 351 7568 367
rect 7583 357 7613 373
rect 7641 351 7647 399
rect 7650 393 7669 399
rect 7684 393 7714 401
rect 7650 385 7714 393
rect 7650 369 7730 385
rect 7746 378 7808 409
rect 7824 378 7886 409
rect 7955 407 8004 432
rect 8019 407 8049 423
rect 7918 393 7948 401
rect 7955 399 8065 407
rect 7918 385 7963 393
rect 7650 367 7669 369
rect 7684 367 7730 369
rect 7650 351 7730 367
rect 7757 365 7792 378
rect 7833 375 7870 378
rect 7833 373 7875 375
rect 7762 362 7792 365
rect 7771 358 7778 362
rect 7778 357 7779 358
rect 7737 351 7747 357
rect 7496 343 7531 351
rect 7496 317 7497 343
rect 7504 317 7531 343
rect 7439 299 7469 313
rect 7496 309 7531 317
rect 7533 343 7574 351
rect 7533 317 7548 343
rect 7555 317 7574 343
rect 7638 339 7669 351
rect 7684 339 7787 351
rect 7799 341 7825 367
rect 7840 362 7870 373
rect 7902 369 7964 385
rect 7902 367 7948 369
rect 7902 351 7964 367
rect 7976 351 7982 399
rect 7985 391 8065 399
rect 7985 389 8004 391
rect 8019 389 8053 391
rect 7985 373 8065 389
rect 7985 351 8004 373
rect 8019 357 8049 373
rect 8077 367 8083 441
rect 8086 367 8105 511
rect 8120 367 8126 511
rect 8135 441 8148 511
rect 8200 506 8222 511
rect 8193 485 8222 499
rect 8275 485 8291 499
rect 8329 495 8335 497
rect 8342 495 8450 511
rect 8457 495 8463 497
rect 8471 495 8486 511
rect 8552 505 8571 508
rect 8193 483 8291 485
rect 8318 483 8486 495
rect 8501 485 8517 499
rect 8552 486 8574 505
rect 8584 499 8600 500
rect 8583 497 8600 499
rect 8584 492 8600 497
rect 8574 485 8580 486
rect 8583 485 8612 492
rect 8501 484 8612 485
rect 8501 483 8618 484
rect 8177 475 8228 483
rect 8275 475 8309 483
rect 8177 463 8202 475
rect 8209 463 8228 475
rect 8282 473 8309 475
rect 8318 473 8539 483
rect 8574 480 8580 483
rect 8282 469 8539 473
rect 8177 455 8228 463
rect 8275 455 8539 469
rect 8583 475 8618 483
rect 8129 407 8148 441
rect 8193 447 8222 455
rect 8193 441 8210 447
rect 8193 439 8227 441
rect 8275 439 8291 455
rect 8292 445 8500 455
rect 8501 445 8517 455
rect 8565 451 8580 466
rect 8583 463 8584 475
rect 8591 463 8618 475
rect 8583 455 8618 463
rect 8583 454 8612 455
rect 8303 441 8517 445
rect 8318 439 8517 441
rect 8552 441 8565 451
rect 8583 441 8600 454
rect 8552 439 8600 441
rect 8194 435 8227 439
rect 8190 433 8227 435
rect 8190 432 8257 433
rect 8190 427 8221 432
rect 8227 427 8257 432
rect 8190 423 8257 427
rect 8163 420 8257 423
rect 8163 413 8212 420
rect 8163 407 8193 413
rect 8212 408 8217 413
rect 8129 391 8209 407
rect 8221 399 8257 420
rect 8318 415 8507 439
rect 8552 438 8599 439
rect 8565 433 8599 438
rect 8333 412 8507 415
rect 8326 409 8507 412
rect 8535 432 8599 433
rect 8129 389 8148 391
rect 8163 389 8197 391
rect 8129 373 8209 389
rect 8129 367 8148 373
rect 7845 341 7948 351
rect 7799 339 7948 341
rect 7969 339 8004 351
rect 7638 337 7800 339
rect 7650 317 7669 337
rect 7684 335 7714 337
rect 7533 309 7574 317
rect 7656 313 7669 317
rect 7721 321 7800 337
rect 7832 337 8004 339
rect 7832 321 7911 337
rect 7918 335 7948 337
rect 7496 299 7525 309
rect 7539 299 7568 309
rect 7583 299 7613 313
rect 7656 299 7699 313
rect 7721 309 7911 321
rect 7976 317 7982 337
rect 7706 299 7736 309
rect 7737 299 7895 309
rect 7899 299 7929 309
rect 7933 299 7963 313
rect 7991 299 8004 337
rect 8076 351 8105 367
rect 8119 351 8148 367
rect 8163 357 8193 373
rect 8221 351 8227 399
rect 8230 393 8249 399
rect 8264 393 8294 401
rect 8230 385 8294 393
rect 8230 369 8310 385
rect 8326 378 8388 409
rect 8404 378 8466 409
rect 8535 407 8584 432
rect 8599 407 8629 423
rect 8498 393 8528 401
rect 8535 399 8645 407
rect 8498 385 8543 393
rect 8230 367 8249 369
rect 8264 367 8310 369
rect 8230 351 8310 367
rect 8337 365 8372 378
rect 8413 375 8450 378
rect 8413 373 8455 375
rect 8342 362 8372 365
rect 8351 358 8358 362
rect 8358 357 8359 358
rect 8317 351 8327 357
rect 8076 343 8111 351
rect 8076 317 8077 343
rect 8084 317 8111 343
rect 8019 299 8049 313
rect 8076 309 8111 317
rect 8113 343 8154 351
rect 8113 317 8128 343
rect 8135 317 8154 343
rect 8218 339 8249 351
rect 8264 339 8367 351
rect 8379 341 8405 367
rect 8420 362 8450 373
rect 8482 369 8544 385
rect 8482 367 8528 369
rect 8482 351 8544 367
rect 8556 351 8562 399
rect 8565 391 8645 399
rect 8565 389 8584 391
rect 8599 389 8633 391
rect 8565 373 8645 389
rect 8565 351 8584 373
rect 8599 357 8629 373
rect 8657 367 8663 441
rect 8666 367 8685 511
rect 8700 367 8706 511
rect 8715 441 8728 511
rect 8780 506 8802 511
rect 8773 485 8802 499
rect 8855 485 8871 499
rect 8909 495 8915 497
rect 8922 495 9030 511
rect 9037 495 9043 497
rect 9051 495 9066 511
rect 9132 505 9151 508
rect 8773 483 8871 485
rect 8898 483 9066 495
rect 9081 485 9097 499
rect 9132 486 9154 505
rect 9164 499 9180 500
rect 9163 497 9180 499
rect 9164 492 9180 497
rect 9154 485 9160 486
rect 9163 485 9192 492
rect 9081 484 9192 485
rect 9081 483 9198 484
rect 8757 475 8808 483
rect 8855 475 8889 483
rect 8757 463 8782 475
rect 8789 463 8808 475
rect 8862 473 8889 475
rect 8898 473 9119 483
rect 9154 480 9160 483
rect 8862 469 9119 473
rect 8757 455 8808 463
rect 8855 455 9119 469
rect 9163 475 9198 483
rect 8709 407 8728 441
rect 8773 447 8802 455
rect 8773 441 8790 447
rect 8773 439 8807 441
rect 8855 439 8871 455
rect 8872 445 9080 455
rect 9081 445 9097 455
rect 9145 451 9160 466
rect 9163 463 9164 475
rect 9171 463 9198 475
rect 9163 455 9198 463
rect 9163 454 9192 455
rect 8883 441 9097 445
rect 8898 439 9097 441
rect 9132 441 9145 451
rect 9163 441 9180 454
rect 9132 439 9180 441
rect 8774 435 8807 439
rect 8770 433 8807 435
rect 8770 432 8837 433
rect 8770 427 8801 432
rect 8807 427 8837 432
rect 8770 423 8837 427
rect 8743 420 8837 423
rect 8743 413 8792 420
rect 8743 407 8773 413
rect 8792 408 8797 413
rect 8709 391 8789 407
rect 8801 399 8837 420
rect 8898 415 9087 439
rect 9132 438 9179 439
rect 9145 433 9179 438
rect 8913 412 9087 415
rect 8906 409 9087 412
rect 9115 432 9179 433
rect 8709 389 8728 391
rect 8743 389 8777 391
rect 8709 373 8789 389
rect 8709 367 8728 373
rect 8425 341 8528 351
rect 8379 339 8528 341
rect 8549 339 8584 351
rect 8218 337 8380 339
rect 8230 317 8249 337
rect 8264 335 8294 337
rect 8113 309 8154 317
rect 8236 313 8249 317
rect 8301 321 8380 337
rect 8412 337 8584 339
rect 8412 321 8491 337
rect 8498 335 8528 337
rect 8076 299 8105 309
rect 8119 299 8148 309
rect 8163 299 8193 313
rect 8236 299 8279 313
rect 8301 309 8491 321
rect 8556 317 8562 337
rect 8286 299 8316 309
rect 8317 299 8475 309
rect 8479 299 8509 309
rect 8513 299 8543 313
rect 8571 299 8584 337
rect 8656 351 8685 367
rect 8699 351 8728 367
rect 8743 357 8773 373
rect 8801 351 8807 399
rect 8810 393 8829 399
rect 8844 393 8874 401
rect 8810 385 8874 393
rect 8810 369 8890 385
rect 8906 378 8968 409
rect 8984 378 9046 409
rect 9115 407 9164 432
rect 9179 407 9209 423
rect 9078 393 9108 401
rect 9115 399 9225 407
rect 9078 385 9123 393
rect 8810 367 8829 369
rect 8844 367 8890 369
rect 8810 351 8890 367
rect 8917 365 8952 378
rect 8993 375 9030 378
rect 8993 373 9035 375
rect 8922 362 8952 365
rect 8931 358 8938 362
rect 8938 357 8939 358
rect 8897 351 8907 357
rect 8656 343 8691 351
rect 8656 317 8657 343
rect 8664 317 8691 343
rect 8599 299 8629 313
rect 8656 309 8691 317
rect 8693 343 8734 351
rect 8693 317 8708 343
rect 8715 317 8734 343
rect 8798 339 8829 351
rect 8844 339 8947 351
rect 8959 341 8985 367
rect 9000 362 9030 373
rect 9062 369 9124 385
rect 9062 367 9108 369
rect 9062 351 9124 367
rect 9136 351 9142 399
rect 9145 391 9225 399
rect 9145 389 9164 391
rect 9179 389 9213 391
rect 9145 373 9225 389
rect 9145 351 9164 373
rect 9179 357 9209 373
rect 9237 367 9243 441
rect 9252 367 9265 511
rect 9005 341 9108 351
rect 8959 339 9108 341
rect 9129 339 9164 351
rect 8798 337 8960 339
rect 8810 317 8829 337
rect 8844 335 8874 337
rect 8693 309 8734 317
rect 8816 313 8829 317
rect 8881 321 8960 337
rect 8992 337 9164 339
rect 8992 321 9071 337
rect 9078 335 9108 337
rect 8656 299 8685 309
rect 8699 299 8728 309
rect 8743 299 8773 313
rect 8816 299 8859 313
rect 8881 309 9071 321
rect 9136 317 9142 337
rect 8866 299 8896 309
rect 8897 299 9055 309
rect 9059 299 9089 309
rect 9093 299 9123 313
rect 9151 299 9164 337
rect 9236 351 9265 367
rect 9236 343 9271 351
rect 9236 317 9237 343
rect 9244 317 9271 343
rect 9179 299 9209 313
rect 9236 309 9271 317
rect 9236 299 9265 309
rect -1 293 9265 299
rect 0 285 9265 293
rect 15 255 28 285
rect 43 271 73 285
rect 116 271 159 285
rect 166 271 386 285
rect 393 271 423 285
rect 83 257 98 269
rect 117 257 130 271
rect 198 267 351 271
rect 80 255 102 257
rect 180 255 372 267
rect 451 255 464 285
rect 479 271 509 285
rect 546 255 565 285
rect 580 255 586 285
rect 595 255 608 285
rect 623 271 653 285
rect 696 271 739 285
rect 746 271 966 285
rect 973 271 1003 285
rect 663 257 678 269
rect 697 257 710 271
rect 778 267 931 271
rect 660 255 682 257
rect 760 255 952 267
rect 1031 255 1044 285
rect 1059 271 1089 285
rect 1126 255 1145 285
rect 1160 255 1166 285
rect 1175 255 1188 285
rect 1203 271 1233 285
rect 1276 271 1319 285
rect 1326 271 1546 285
rect 1553 271 1583 285
rect 1243 257 1258 269
rect 1277 257 1290 271
rect 1358 267 1511 271
rect 1240 255 1262 257
rect 1340 255 1532 267
rect 1611 255 1624 285
rect 1639 271 1669 285
rect 1706 255 1725 285
rect 1740 255 1746 285
rect 1755 255 1768 285
rect 1783 271 1813 285
rect 1856 271 1899 285
rect 1906 271 2126 285
rect 2133 271 2163 285
rect 1823 257 1838 269
rect 1857 257 1870 271
rect 1938 267 2091 271
rect 1820 255 1842 257
rect 1920 255 2112 267
rect 2191 255 2204 285
rect 2219 271 2249 285
rect 2286 255 2305 285
rect 2320 255 2326 285
rect 2335 255 2348 285
rect 2363 271 2393 285
rect 2436 271 2479 285
rect 2486 271 2706 285
rect 2713 271 2743 285
rect 2403 257 2418 269
rect 2437 257 2450 271
rect 2518 267 2671 271
rect 2400 255 2422 257
rect 2500 255 2692 267
rect 2771 255 2784 285
rect 2799 271 2829 285
rect 2866 255 2885 285
rect 2900 255 2906 285
rect 2915 255 2928 285
rect 2943 271 2973 285
rect 3016 271 3059 285
rect 3066 271 3286 285
rect 3293 271 3323 285
rect 2983 257 2998 269
rect 3017 257 3030 271
rect 3098 267 3251 271
rect 2980 255 3002 257
rect 3080 255 3272 267
rect 3351 255 3364 285
rect 3379 271 3409 285
rect 3446 255 3465 285
rect 3480 255 3486 285
rect 3495 255 3508 285
rect 3523 271 3553 285
rect 3596 271 3639 285
rect 3646 271 3866 285
rect 3873 271 3903 285
rect 3563 257 3578 269
rect 3597 257 3610 271
rect 3678 267 3831 271
rect 3560 255 3582 257
rect 3660 255 3852 267
rect 3931 255 3944 285
rect 3959 271 3989 285
rect 4026 255 4045 285
rect 4060 255 4066 285
rect 4075 255 4088 285
rect 4103 271 4133 285
rect 4176 271 4219 285
rect 4226 271 4446 285
rect 4453 271 4483 285
rect 4143 257 4158 269
rect 4177 257 4190 271
rect 4258 267 4411 271
rect 4140 255 4162 257
rect 4240 255 4432 267
rect 4511 255 4524 285
rect 4539 271 4569 285
rect 4606 284 4646 285
rect 4606 255 4625 284
rect 4640 255 4646 284
rect 4655 255 4668 285
rect 4683 271 4713 285
rect 4756 271 4799 285
rect 4806 271 5026 285
rect 5033 271 5063 285
rect 4723 257 4738 269
rect 4757 257 4770 271
rect 4838 267 4991 271
rect 4720 255 4742 257
rect 4820 255 5012 267
rect 5091 255 5104 285
rect 5119 271 5149 285
rect 5186 255 5205 285
rect 5220 255 5226 285
rect 5235 255 5248 285
rect 5263 271 5293 285
rect 5336 271 5379 285
rect 5386 271 5606 285
rect 5613 271 5643 285
rect 5303 257 5318 269
rect 5337 257 5350 271
rect 5418 267 5571 271
rect 5300 255 5322 257
rect 5400 255 5592 267
rect 5671 255 5684 285
rect 5699 271 5729 285
rect 5766 255 5785 285
rect 5800 255 5806 285
rect 5815 255 5828 285
rect 5843 271 5873 285
rect 5916 271 5959 285
rect 5966 271 6186 285
rect 6193 271 6223 285
rect 5883 257 5898 269
rect 5917 257 5930 271
rect 5998 267 6151 271
rect 5880 255 5902 257
rect 5980 255 6172 267
rect 6251 255 6264 285
rect 6279 271 6309 285
rect 6346 255 6365 285
rect 6380 255 6386 285
rect 6395 255 6408 285
rect 6423 271 6453 285
rect 6496 271 6539 285
rect 6546 271 6766 285
rect 6773 271 6803 285
rect 6463 257 6478 269
rect 6497 257 6510 271
rect 6578 267 6731 271
rect 6460 255 6482 257
rect 6560 255 6752 267
rect 6831 255 6844 285
rect 6859 271 6889 285
rect 6926 255 6945 285
rect 6960 255 6966 285
rect 6975 255 6988 285
rect 7003 271 7033 285
rect 7076 271 7119 285
rect 7126 271 7346 285
rect 7353 271 7383 285
rect 7043 257 7058 269
rect 7077 257 7090 271
rect 7158 267 7311 271
rect 7040 255 7062 257
rect 7140 255 7332 267
rect 7411 255 7424 285
rect 7439 271 7469 285
rect 7506 255 7525 285
rect 7540 255 7546 285
rect 7555 255 7568 285
rect 7583 271 7613 285
rect 7656 271 7699 285
rect 7706 271 7926 285
rect 7933 271 7963 285
rect 7623 257 7638 269
rect 7657 257 7670 271
rect 7738 267 7891 271
rect 7620 255 7642 257
rect 7720 255 7912 267
rect 7991 255 8004 285
rect 8019 271 8049 285
rect 8086 255 8105 285
rect 8120 255 8126 285
rect 8135 255 8148 285
rect 8163 271 8193 285
rect 8236 271 8279 285
rect 8286 271 8506 285
rect 8513 271 8543 285
rect 8203 257 8218 269
rect 8237 257 8250 271
rect 8318 267 8471 271
rect 8200 255 8222 257
rect 8300 255 8492 267
rect 8571 255 8584 285
rect 8599 271 8629 285
rect 8666 255 8685 285
rect 8700 255 8706 285
rect 8715 255 8728 285
rect 8743 271 8773 285
rect 8816 271 8859 285
rect 8866 271 9086 285
rect 9093 271 9123 285
rect 8783 257 8798 269
rect 8817 257 8830 271
rect 8898 267 9051 271
rect 8780 255 8802 257
rect 8880 255 9072 267
rect 9151 255 9164 285
rect 9179 271 9209 285
rect 9252 255 9265 285
rect 0 241 9265 255
rect 15 171 28 241
rect 80 237 102 241
rect 73 215 102 229
rect 155 215 171 229
rect 209 219 215 227
rect 222 225 330 241
rect 73 213 171 215
rect 57 205 108 213
rect 155 205 189 213
rect 57 193 82 205
rect 89 193 108 205
rect 162 203 189 205
rect 198 205 215 219
rect 260 205 292 225
rect 337 219 343 227
rect 351 219 366 241
rect 432 235 451 238
rect 337 213 366 219
rect 381 215 397 229
rect 432 216 454 235
rect 464 229 480 230
rect 463 227 480 229
rect 464 222 480 227
rect 454 215 460 216
rect 463 215 492 222
rect 381 214 492 215
rect 381 213 498 214
rect 337 205 419 213
rect 454 210 460 213
rect 198 203 419 205
rect 162 199 234 203
rect 262 201 290 203
rect 57 185 108 193
rect 155 191 287 199
rect 290 191 301 199
rect 155 189 234 191
rect 315 189 419 203
rect 463 205 498 213
rect 155 185 252 189
rect 9 137 28 171
rect 73 177 102 185
rect 73 171 90 177
rect 73 169 107 171
rect 155 169 171 185
rect 172 181 252 185
rect 300 185 419 189
rect 300 181 380 185
rect 172 175 380 181
rect 381 175 397 185
rect 445 181 460 196
rect 463 193 464 205
rect 471 193 498 205
rect 463 185 498 193
rect 463 184 492 185
rect 183 171 293 175
rect 74 165 107 169
rect 70 163 107 165
rect 70 162 137 163
rect 70 157 101 162
rect 107 157 137 162
rect 198 159 213 171
rect 70 153 137 157
rect 43 150 137 153
rect 43 143 92 150
rect 43 137 73 143
rect 92 138 97 143
rect 9 121 89 137
rect 101 129 137 150
rect 222 149 252 158
rect 275 153 293 171
rect 351 169 397 175
rect 432 171 445 181
rect 463 171 480 184
rect 432 169 480 171
rect 313 163 315 165
rect 315 161 317 163
rect 317 158 327 161
rect 300 151 330 158
rect 300 149 331 151
rect 351 149 387 169
rect 432 168 479 169
rect 445 163 479 168
rect 198 145 387 149
rect 213 142 387 145
rect 206 139 387 142
rect 415 162 479 163
rect 9 119 28 121
rect 43 119 77 121
rect 9 103 89 119
rect 9 97 28 103
rect -1 81 28 97
rect 43 87 73 103
rect 101 81 107 129
rect 110 123 129 129
rect 144 123 174 131
rect 110 115 174 123
rect 110 99 190 115
rect 206 108 268 139
rect 284 108 346 139
rect 415 137 464 162
rect 479 137 509 153
rect 378 123 408 131
rect 415 129 525 137
rect 378 115 423 123
rect 217 105 221 108
rect 222 105 252 108
rect 110 97 129 99
rect 144 97 190 99
rect 110 81 190 97
rect 221 95 252 105
rect 293 105 299 108
rect 300 105 330 108
rect 293 103 335 105
rect 222 92 252 95
rect 231 88 238 92
rect 238 87 239 88
rect 197 81 207 87
rect 259 81 275 97
rect 300 92 330 103
rect 362 99 424 115
rect 362 97 408 99
rect 362 81 424 97
rect 436 81 442 129
rect 445 121 525 129
rect 445 119 464 121
rect 479 119 513 121
rect 445 103 525 119
rect 445 81 464 103
rect 479 87 509 103
rect 537 97 543 171
rect 546 97 565 241
rect 580 97 586 241
rect 595 171 608 241
rect 660 237 682 241
rect 653 215 682 229
rect 735 215 751 229
rect 789 219 795 227
rect 802 225 910 241
rect 653 213 751 215
rect 637 205 688 213
rect 735 205 769 213
rect 637 193 662 205
rect 669 193 688 205
rect 742 203 769 205
rect 778 205 795 219
rect 840 205 872 225
rect 917 219 923 227
rect 931 219 946 241
rect 1012 235 1031 238
rect 917 213 946 219
rect 961 215 977 229
rect 1012 216 1034 235
rect 1044 229 1060 230
rect 1043 227 1060 229
rect 1044 222 1060 227
rect 1034 215 1040 216
rect 1043 215 1072 222
rect 961 214 1072 215
rect 961 213 1078 214
rect 917 205 999 213
rect 1034 210 1040 213
rect 778 203 999 205
rect 742 199 814 203
rect 842 201 870 203
rect 637 185 688 193
rect 735 191 867 199
rect 870 191 881 199
rect 735 189 814 191
rect 895 189 999 203
rect 1043 205 1078 213
rect 735 185 832 189
rect 589 137 608 171
rect 653 177 682 185
rect 653 171 670 177
rect 653 169 687 171
rect 735 169 751 185
rect 752 181 832 185
rect 880 185 999 189
rect 880 181 960 185
rect 752 175 960 181
rect 961 175 977 185
rect 1025 181 1040 196
rect 1043 193 1044 205
rect 1051 193 1078 205
rect 1043 185 1078 193
rect 1043 184 1072 185
rect 763 171 873 175
rect 654 165 687 169
rect 650 163 687 165
rect 650 162 717 163
rect 650 157 681 162
rect 687 157 717 162
rect 778 159 793 171
rect 650 153 717 157
rect 623 150 717 153
rect 623 143 672 150
rect 623 137 653 143
rect 672 138 677 143
rect 589 121 669 137
rect 681 129 717 150
rect 802 149 832 158
rect 855 153 873 171
rect 931 169 977 175
rect 1012 171 1025 181
rect 1043 171 1060 184
rect 1012 169 1060 171
rect 893 163 895 165
rect 895 161 897 163
rect 897 158 907 161
rect 880 151 910 158
rect 880 149 911 151
rect 931 149 967 169
rect 1012 168 1059 169
rect 1025 163 1059 168
rect 778 145 967 149
rect 793 142 967 145
rect 786 139 967 142
rect 995 162 1059 163
rect 589 119 608 121
rect 623 119 657 121
rect 589 103 669 119
rect 589 97 608 103
rect -7 73 34 81
rect -7 47 8 73
rect 15 47 34 73
rect 98 69 129 81
rect 144 69 247 81
rect 259 71 285 81
rect 305 71 408 81
rect 259 69 408 71
rect 429 69 464 81
rect 98 67 260 69
rect 110 47 129 67
rect 144 65 174 67
rect -7 39 34 47
rect -1 29 28 39
rect 116 29 129 47
rect 181 51 260 67
rect 292 67 464 69
rect 292 51 371 67
rect 378 65 408 67
rect 181 43 371 51
rect 436 47 442 67
rect 181 39 260 43
rect 262 39 290 43
rect 292 39 371 43
rect 166 29 174 39
rect 193 31 196 39
rect 197 31 215 39
rect 260 31 292 39
rect 337 31 355 39
rect 193 29 359 31
rect 378 29 389 39
rect 451 29 464 67
rect 536 81 565 97
rect 579 81 608 97
rect 623 87 653 103
rect 681 81 687 129
rect 690 123 709 129
rect 724 123 754 131
rect 690 115 754 123
rect 690 99 770 115
rect 786 108 848 139
rect 864 108 926 139
rect 995 137 1044 162
rect 1059 137 1089 153
rect 958 123 988 131
rect 995 129 1105 137
rect 958 115 1003 123
rect 797 105 801 108
rect 802 105 832 108
rect 690 97 709 99
rect 724 97 770 99
rect 690 81 770 97
rect 801 95 832 105
rect 873 105 879 108
rect 880 105 910 108
rect 873 103 915 105
rect 802 92 832 95
rect 811 88 818 92
rect 818 87 819 88
rect 777 81 787 87
rect 839 81 855 97
rect 880 92 910 103
rect 942 99 1004 115
rect 942 97 988 99
rect 942 81 1004 97
rect 1016 81 1022 129
rect 1025 121 1105 129
rect 1025 119 1044 121
rect 1059 119 1093 121
rect 1025 103 1105 119
rect 1025 81 1044 103
rect 1059 87 1089 103
rect 1117 97 1123 171
rect 1126 97 1145 241
rect 1160 97 1166 241
rect 1175 171 1188 241
rect 1240 237 1262 241
rect 1233 215 1262 229
rect 1315 215 1331 229
rect 1369 219 1375 227
rect 1382 225 1490 241
rect 1233 213 1331 215
rect 1217 205 1268 213
rect 1315 205 1349 213
rect 1217 193 1242 205
rect 1249 193 1268 205
rect 1322 203 1349 205
rect 1358 205 1375 219
rect 1420 205 1452 225
rect 1497 219 1503 227
rect 1511 219 1526 241
rect 1592 235 1611 238
rect 1497 213 1526 219
rect 1541 215 1557 229
rect 1592 216 1614 235
rect 1624 229 1640 230
rect 1623 227 1640 229
rect 1624 222 1640 227
rect 1614 215 1620 216
rect 1623 215 1652 222
rect 1541 214 1652 215
rect 1541 213 1658 214
rect 1497 205 1579 213
rect 1614 210 1620 213
rect 1358 203 1579 205
rect 1322 199 1394 203
rect 1422 201 1450 203
rect 1217 185 1268 193
rect 1315 191 1447 199
rect 1450 191 1461 199
rect 1315 189 1394 191
rect 1475 189 1579 203
rect 1623 205 1658 213
rect 1315 185 1412 189
rect 1169 137 1188 171
rect 1233 177 1262 185
rect 1233 171 1250 177
rect 1233 169 1267 171
rect 1315 169 1331 185
rect 1332 181 1412 185
rect 1460 185 1579 189
rect 1460 181 1540 185
rect 1332 175 1540 181
rect 1541 175 1557 185
rect 1605 181 1620 196
rect 1623 193 1624 205
rect 1631 193 1658 205
rect 1623 185 1658 193
rect 1623 184 1652 185
rect 1343 171 1453 175
rect 1234 165 1267 169
rect 1230 163 1267 165
rect 1230 162 1297 163
rect 1230 157 1261 162
rect 1267 157 1297 162
rect 1358 159 1373 171
rect 1230 153 1297 157
rect 1203 150 1297 153
rect 1203 143 1252 150
rect 1203 137 1233 143
rect 1252 138 1257 143
rect 1169 121 1249 137
rect 1261 129 1297 150
rect 1382 149 1412 158
rect 1435 153 1453 171
rect 1511 169 1557 175
rect 1592 171 1605 181
rect 1623 171 1640 184
rect 1592 169 1640 171
rect 1473 163 1475 165
rect 1475 161 1477 163
rect 1477 158 1487 161
rect 1460 151 1490 158
rect 1460 149 1491 151
rect 1511 149 1547 169
rect 1592 168 1639 169
rect 1605 163 1639 168
rect 1358 145 1547 149
rect 1373 142 1547 145
rect 1366 139 1547 142
rect 1575 162 1639 163
rect 1169 119 1188 121
rect 1203 119 1237 121
rect 1169 103 1249 119
rect 1169 97 1188 103
rect 536 73 571 81
rect 536 47 537 73
rect 544 47 571 73
rect 536 39 571 47
rect 573 73 614 81
rect 573 47 588 73
rect 595 47 614 73
rect 678 69 709 81
rect 724 69 827 81
rect 839 71 865 81
rect 885 71 988 81
rect 839 69 988 71
rect 1009 69 1044 81
rect 678 67 840 69
rect 690 47 709 67
rect 724 65 754 67
rect 573 39 614 47
rect 536 29 565 39
rect 579 29 608 39
rect 696 29 709 47
rect 761 51 840 67
rect 872 67 1044 69
rect 872 51 951 67
rect 958 65 988 67
rect 761 43 951 51
rect 1016 47 1022 67
rect 761 39 840 43
rect 842 39 870 43
rect 872 39 951 43
rect 746 29 754 39
rect 773 31 776 39
rect 777 31 795 39
rect 840 31 872 39
rect 917 31 935 39
rect 773 29 939 31
rect 958 29 969 39
rect 1031 29 1044 67
rect 1116 81 1145 97
rect 1159 81 1188 97
rect 1203 87 1233 103
rect 1261 81 1267 129
rect 1270 123 1289 129
rect 1304 123 1334 131
rect 1270 115 1334 123
rect 1270 99 1350 115
rect 1366 108 1428 139
rect 1444 108 1506 139
rect 1575 137 1624 162
rect 1639 137 1669 153
rect 1538 123 1568 131
rect 1575 129 1685 137
rect 1538 115 1583 123
rect 1377 105 1381 108
rect 1382 105 1412 108
rect 1270 97 1289 99
rect 1304 97 1350 99
rect 1270 81 1350 97
rect 1381 95 1412 105
rect 1453 105 1459 108
rect 1460 105 1490 108
rect 1453 103 1495 105
rect 1382 92 1412 95
rect 1391 88 1398 92
rect 1398 87 1399 88
rect 1357 81 1367 87
rect 1419 81 1435 97
rect 1460 92 1490 103
rect 1522 99 1584 115
rect 1522 97 1568 99
rect 1522 81 1584 97
rect 1596 81 1602 129
rect 1605 121 1685 129
rect 1605 119 1624 121
rect 1639 119 1673 121
rect 1605 103 1685 119
rect 1605 81 1624 103
rect 1639 87 1669 103
rect 1697 97 1703 171
rect 1706 97 1725 241
rect 1740 97 1746 241
rect 1755 171 1768 241
rect 1820 237 1842 241
rect 1813 215 1842 229
rect 1895 215 1911 229
rect 1949 219 1955 227
rect 1962 225 2070 241
rect 1813 213 1911 215
rect 1797 205 1848 213
rect 1895 205 1929 213
rect 1797 193 1822 205
rect 1829 193 1848 205
rect 1902 203 1929 205
rect 1938 205 1955 219
rect 2000 205 2032 225
rect 2077 219 2083 227
rect 2091 219 2106 241
rect 2172 235 2191 238
rect 2077 213 2106 219
rect 2121 215 2137 229
rect 2172 216 2194 235
rect 2204 229 2220 230
rect 2203 227 2220 229
rect 2204 222 2220 227
rect 2194 215 2200 216
rect 2203 215 2232 222
rect 2121 214 2232 215
rect 2121 213 2238 214
rect 2077 205 2159 213
rect 2194 210 2200 213
rect 1938 203 2159 205
rect 1902 199 1974 203
rect 2002 201 2030 203
rect 1797 185 1848 193
rect 1895 191 2027 199
rect 2030 191 2041 199
rect 1895 189 1974 191
rect 2055 189 2159 203
rect 2203 205 2238 213
rect 1895 185 1992 189
rect 1749 137 1768 171
rect 1813 177 1842 185
rect 1813 171 1830 177
rect 1813 169 1847 171
rect 1895 169 1911 185
rect 1912 181 1992 185
rect 2040 185 2159 189
rect 2040 181 2120 185
rect 1912 175 2120 181
rect 2121 175 2137 185
rect 2185 181 2200 196
rect 2203 193 2204 205
rect 2211 193 2238 205
rect 2203 185 2238 193
rect 2203 184 2232 185
rect 1923 171 2033 175
rect 1814 165 1847 169
rect 1810 163 1847 165
rect 1810 162 1877 163
rect 1810 157 1841 162
rect 1847 157 1877 162
rect 1938 159 1953 171
rect 1810 153 1877 157
rect 1783 150 1877 153
rect 1783 143 1832 150
rect 1783 137 1813 143
rect 1832 138 1837 143
rect 1749 121 1829 137
rect 1841 129 1877 150
rect 1962 149 1992 158
rect 2015 153 2033 171
rect 2091 169 2137 175
rect 2172 171 2185 181
rect 2203 171 2220 184
rect 2172 169 2220 171
rect 2053 163 2055 165
rect 2055 161 2057 163
rect 2057 158 2067 161
rect 2040 151 2070 158
rect 2040 149 2071 151
rect 2091 149 2127 169
rect 2172 168 2219 169
rect 2185 163 2219 168
rect 1938 145 2127 149
rect 1953 142 2127 145
rect 1946 139 2127 142
rect 2155 162 2219 163
rect 1749 119 1768 121
rect 1783 119 1817 121
rect 1749 103 1829 119
rect 1749 97 1768 103
rect 1116 73 1151 81
rect 1116 47 1117 73
rect 1124 47 1151 73
rect 1116 39 1151 47
rect 1153 73 1194 81
rect 1153 47 1168 73
rect 1175 47 1194 73
rect 1258 69 1289 81
rect 1304 69 1407 81
rect 1419 71 1445 81
rect 1465 71 1568 81
rect 1419 69 1568 71
rect 1589 69 1624 81
rect 1258 67 1420 69
rect 1270 47 1289 67
rect 1304 65 1334 67
rect 1153 39 1194 47
rect 1116 29 1145 39
rect 1159 29 1188 39
rect 1276 29 1289 47
rect 1341 51 1420 67
rect 1452 67 1624 69
rect 1452 51 1531 67
rect 1538 65 1568 67
rect 1341 43 1531 51
rect 1596 47 1602 67
rect 1341 39 1420 43
rect 1422 39 1450 43
rect 1452 39 1531 43
rect 1326 29 1334 39
rect 1353 31 1356 39
rect 1357 31 1375 39
rect 1420 31 1452 39
rect 1497 31 1515 39
rect 1353 29 1519 31
rect 1538 29 1549 39
rect 1611 29 1624 67
rect 1696 81 1725 97
rect 1739 81 1768 97
rect 1783 87 1813 103
rect 1841 81 1847 129
rect 1850 123 1869 129
rect 1884 123 1914 131
rect 1850 115 1914 123
rect 1850 99 1930 115
rect 1946 108 2008 139
rect 2024 108 2086 139
rect 2155 137 2204 162
rect 2219 137 2249 153
rect 2118 123 2148 131
rect 2155 129 2265 137
rect 2118 115 2163 123
rect 1957 105 1961 108
rect 1962 105 1992 108
rect 1850 97 1869 99
rect 1884 97 1930 99
rect 1850 81 1930 97
rect 1961 95 1992 105
rect 2033 105 2039 108
rect 2040 105 2070 108
rect 2033 103 2075 105
rect 1962 92 1992 95
rect 1971 88 1978 92
rect 1978 87 1979 88
rect 1937 81 1947 87
rect 1999 81 2015 97
rect 2040 92 2070 103
rect 2102 99 2164 115
rect 2102 97 2148 99
rect 2102 81 2164 97
rect 2176 81 2182 129
rect 2185 121 2265 129
rect 2185 119 2204 121
rect 2219 119 2253 121
rect 2185 103 2265 119
rect 2185 81 2204 103
rect 2219 87 2249 103
rect 2277 97 2283 171
rect 2286 97 2305 241
rect 2320 97 2326 241
rect 2335 171 2348 241
rect 2400 237 2422 241
rect 2393 215 2422 229
rect 2475 215 2491 229
rect 2529 219 2535 227
rect 2542 225 2650 241
rect 2393 213 2491 215
rect 2377 205 2428 213
rect 2475 205 2509 213
rect 2377 193 2402 205
rect 2409 193 2428 205
rect 2482 203 2509 205
rect 2518 205 2535 219
rect 2580 205 2612 225
rect 2657 219 2663 227
rect 2671 219 2686 241
rect 2752 235 2771 238
rect 2657 213 2686 219
rect 2701 215 2717 229
rect 2752 216 2774 235
rect 2784 229 2800 230
rect 2783 227 2800 229
rect 2784 222 2800 227
rect 2774 215 2780 216
rect 2783 215 2812 222
rect 2701 214 2812 215
rect 2701 213 2818 214
rect 2657 205 2739 213
rect 2774 210 2780 213
rect 2518 203 2739 205
rect 2482 199 2554 203
rect 2582 201 2610 203
rect 2377 185 2428 193
rect 2475 191 2607 199
rect 2610 191 2621 199
rect 2475 189 2554 191
rect 2635 189 2739 203
rect 2783 205 2818 213
rect 2475 185 2572 189
rect 2329 137 2348 171
rect 2393 177 2422 185
rect 2393 171 2410 177
rect 2393 169 2427 171
rect 2475 169 2491 185
rect 2492 181 2572 185
rect 2620 185 2739 189
rect 2620 181 2700 185
rect 2492 175 2700 181
rect 2701 175 2717 185
rect 2765 181 2780 196
rect 2783 193 2784 205
rect 2791 193 2818 205
rect 2783 185 2818 193
rect 2783 184 2812 185
rect 2503 171 2613 175
rect 2394 165 2427 169
rect 2390 163 2427 165
rect 2390 162 2457 163
rect 2390 157 2421 162
rect 2427 157 2457 162
rect 2518 159 2533 171
rect 2390 153 2457 157
rect 2363 150 2457 153
rect 2363 143 2412 150
rect 2363 137 2393 143
rect 2412 138 2417 143
rect 2329 121 2409 137
rect 2421 129 2457 150
rect 2542 149 2572 158
rect 2595 153 2613 171
rect 2671 169 2717 175
rect 2752 171 2765 181
rect 2783 171 2800 184
rect 2752 169 2800 171
rect 2633 163 2635 165
rect 2635 161 2637 163
rect 2637 158 2647 161
rect 2620 151 2650 158
rect 2620 149 2651 151
rect 2671 149 2707 169
rect 2752 168 2799 169
rect 2765 163 2799 168
rect 2518 145 2707 149
rect 2533 142 2707 145
rect 2526 139 2707 142
rect 2735 162 2799 163
rect 2329 119 2348 121
rect 2363 119 2397 121
rect 2329 103 2409 119
rect 2329 97 2348 103
rect 1696 73 1731 81
rect 1696 47 1697 73
rect 1704 47 1731 73
rect 1696 39 1731 47
rect 1733 73 1774 81
rect 1733 47 1748 73
rect 1755 47 1774 73
rect 1838 69 1869 81
rect 1884 69 1987 81
rect 1999 71 2025 81
rect 2045 71 2148 81
rect 1999 69 2148 71
rect 2169 69 2204 81
rect 1838 67 2000 69
rect 1850 47 1869 67
rect 1884 65 1914 67
rect 1733 39 1774 47
rect 1696 29 1725 39
rect 1739 29 1768 39
rect 1856 29 1869 47
rect 1921 51 2000 67
rect 2032 67 2204 69
rect 2032 51 2111 67
rect 2118 65 2148 67
rect 1921 43 2111 51
rect 2176 47 2182 67
rect 1921 39 2000 43
rect 2002 39 2030 43
rect 2032 39 2111 43
rect 1906 29 1914 39
rect 1933 31 1936 39
rect 1937 31 1955 39
rect 2000 31 2032 39
rect 2077 31 2095 39
rect 1933 29 2099 31
rect 2118 29 2129 39
rect 2191 29 2204 67
rect 2276 81 2305 97
rect 2319 81 2348 97
rect 2363 87 2393 103
rect 2421 81 2427 129
rect 2430 123 2449 129
rect 2464 123 2494 131
rect 2430 115 2494 123
rect 2430 99 2510 115
rect 2526 108 2588 139
rect 2604 108 2666 139
rect 2735 137 2784 162
rect 2799 137 2829 153
rect 2698 123 2728 131
rect 2735 129 2845 137
rect 2698 115 2743 123
rect 2537 105 2541 108
rect 2542 105 2572 108
rect 2430 97 2449 99
rect 2464 97 2510 99
rect 2430 81 2510 97
rect 2541 95 2572 105
rect 2613 105 2619 108
rect 2620 105 2650 108
rect 2613 103 2655 105
rect 2542 92 2572 95
rect 2551 88 2558 92
rect 2558 87 2559 88
rect 2517 81 2527 87
rect 2579 81 2595 97
rect 2620 92 2650 103
rect 2682 99 2744 115
rect 2682 97 2728 99
rect 2682 81 2744 97
rect 2756 81 2762 129
rect 2765 121 2845 129
rect 2765 119 2784 121
rect 2799 119 2833 121
rect 2765 103 2845 119
rect 2765 81 2784 103
rect 2799 87 2829 103
rect 2857 97 2863 171
rect 2866 97 2885 241
rect 2900 97 2906 241
rect 2915 171 2928 241
rect 2980 237 3002 241
rect 2973 215 3002 229
rect 3055 215 3071 229
rect 3109 219 3115 227
rect 3122 225 3230 241
rect 2973 213 3071 215
rect 2957 205 3008 213
rect 3055 205 3089 213
rect 2957 193 2982 205
rect 2989 193 3008 205
rect 3062 203 3089 205
rect 3098 205 3115 219
rect 3160 205 3192 225
rect 3237 219 3243 227
rect 3251 219 3266 241
rect 3332 235 3351 238
rect 3237 213 3266 219
rect 3281 215 3297 229
rect 3332 216 3354 235
rect 3364 229 3380 230
rect 3363 227 3380 229
rect 3364 222 3380 227
rect 3354 215 3360 216
rect 3363 215 3392 222
rect 3281 214 3392 215
rect 3281 213 3398 214
rect 3237 205 3319 213
rect 3354 210 3360 213
rect 3098 203 3319 205
rect 3062 199 3134 203
rect 3162 201 3190 203
rect 2957 185 3008 193
rect 3055 191 3187 199
rect 3190 191 3201 199
rect 3055 189 3134 191
rect 3215 189 3319 203
rect 3363 205 3398 213
rect 3055 185 3152 189
rect 2909 137 2928 171
rect 2973 177 3002 185
rect 2973 171 2990 177
rect 2973 169 3007 171
rect 3055 169 3071 185
rect 3072 181 3152 185
rect 3200 185 3319 189
rect 3200 181 3280 185
rect 3072 175 3280 181
rect 3281 175 3297 185
rect 3345 181 3360 196
rect 3363 193 3364 205
rect 3371 193 3398 205
rect 3363 185 3398 193
rect 3363 184 3392 185
rect 3083 171 3193 175
rect 2974 165 3007 169
rect 2970 163 3007 165
rect 2970 162 3037 163
rect 2970 157 3001 162
rect 3007 157 3037 162
rect 3098 159 3113 171
rect 2970 153 3037 157
rect 2943 150 3037 153
rect 2943 143 2992 150
rect 2943 137 2973 143
rect 2992 138 2997 143
rect 2909 121 2989 137
rect 3001 129 3037 150
rect 3122 149 3152 158
rect 3175 153 3193 171
rect 3251 169 3297 175
rect 3332 171 3345 181
rect 3363 171 3380 184
rect 3332 169 3380 171
rect 3213 163 3215 165
rect 3215 161 3217 163
rect 3217 158 3227 161
rect 3200 151 3230 158
rect 3200 149 3231 151
rect 3251 149 3287 169
rect 3332 168 3379 169
rect 3345 163 3379 168
rect 3098 145 3287 149
rect 3113 142 3287 145
rect 3106 139 3287 142
rect 3315 162 3379 163
rect 2909 119 2928 121
rect 2943 119 2977 121
rect 2909 103 2989 119
rect 2909 97 2928 103
rect 2276 73 2311 81
rect 2276 47 2277 73
rect 2284 47 2311 73
rect 2276 39 2311 47
rect 2313 73 2354 81
rect 2313 47 2328 73
rect 2335 47 2354 73
rect 2418 69 2449 81
rect 2464 69 2567 81
rect 2579 71 2605 81
rect 2625 71 2728 81
rect 2579 69 2728 71
rect 2749 69 2784 81
rect 2418 67 2580 69
rect 2430 47 2449 67
rect 2464 65 2494 67
rect 2313 39 2354 47
rect 2276 29 2305 39
rect 2319 29 2348 39
rect 2436 29 2449 47
rect 2501 51 2580 67
rect 2612 67 2784 69
rect 2612 51 2691 67
rect 2698 65 2728 67
rect 2501 43 2691 51
rect 2756 47 2762 67
rect 2501 39 2580 43
rect 2582 39 2610 43
rect 2612 39 2691 43
rect 2486 29 2494 39
rect 2513 31 2516 39
rect 2517 31 2535 39
rect 2580 31 2612 39
rect 2657 31 2675 39
rect 2513 29 2679 31
rect 2698 29 2709 39
rect 2771 29 2784 67
rect 2856 81 2885 97
rect 2899 81 2928 97
rect 2943 87 2973 103
rect 3001 81 3007 129
rect 3010 123 3029 129
rect 3044 123 3074 131
rect 3010 115 3074 123
rect 3010 99 3090 115
rect 3106 108 3168 139
rect 3184 108 3246 139
rect 3315 137 3364 162
rect 3379 137 3409 153
rect 3278 123 3308 131
rect 3315 129 3425 137
rect 3278 115 3323 123
rect 3117 105 3121 108
rect 3122 105 3152 108
rect 3010 97 3029 99
rect 3044 97 3090 99
rect 3010 81 3090 97
rect 3121 95 3152 105
rect 3193 105 3199 108
rect 3200 105 3230 108
rect 3193 103 3235 105
rect 3122 92 3152 95
rect 3131 88 3138 92
rect 3138 87 3139 88
rect 3097 81 3107 87
rect 3159 81 3175 97
rect 3200 92 3230 103
rect 3262 99 3324 115
rect 3262 97 3308 99
rect 3262 81 3324 97
rect 3336 81 3342 129
rect 3345 121 3425 129
rect 3345 119 3364 121
rect 3379 119 3413 121
rect 3345 103 3425 119
rect 3345 81 3364 103
rect 3379 87 3409 103
rect 3437 97 3443 171
rect 3446 97 3465 241
rect 3480 97 3486 241
rect 3495 171 3508 241
rect 3560 237 3582 241
rect 3553 215 3582 229
rect 3635 215 3651 229
rect 3689 219 3695 227
rect 3702 225 3810 241
rect 3553 213 3651 215
rect 3537 205 3588 213
rect 3635 205 3669 213
rect 3537 193 3562 205
rect 3569 193 3588 205
rect 3642 203 3669 205
rect 3678 205 3695 219
rect 3740 205 3772 225
rect 3817 219 3823 227
rect 3831 219 3846 241
rect 3912 235 3931 238
rect 3817 213 3846 219
rect 3861 215 3877 229
rect 3912 216 3934 235
rect 3944 229 3960 230
rect 3943 227 3960 229
rect 3944 222 3960 227
rect 3934 215 3940 216
rect 3943 215 3972 222
rect 3861 214 3972 215
rect 3861 213 3978 214
rect 3817 205 3899 213
rect 3934 210 3940 213
rect 3678 203 3899 205
rect 3642 199 3714 203
rect 3742 201 3770 203
rect 3537 185 3588 193
rect 3635 191 3767 199
rect 3770 191 3781 199
rect 3635 189 3714 191
rect 3795 189 3899 203
rect 3943 205 3978 213
rect 3635 185 3732 189
rect 3489 137 3508 171
rect 3553 177 3582 185
rect 3553 171 3570 177
rect 3553 169 3587 171
rect 3635 169 3651 185
rect 3652 181 3732 185
rect 3780 185 3899 189
rect 3780 181 3860 185
rect 3652 175 3860 181
rect 3861 175 3877 185
rect 3925 181 3940 196
rect 3943 193 3944 205
rect 3951 193 3978 205
rect 3943 185 3978 193
rect 3943 184 3972 185
rect 3663 171 3773 175
rect 3554 165 3587 169
rect 3550 163 3587 165
rect 3550 162 3617 163
rect 3550 157 3581 162
rect 3587 157 3617 162
rect 3678 159 3693 171
rect 3550 153 3617 157
rect 3523 150 3617 153
rect 3523 143 3572 150
rect 3523 137 3553 143
rect 3572 138 3577 143
rect 3489 121 3569 137
rect 3581 129 3617 150
rect 3702 149 3732 158
rect 3755 153 3773 171
rect 3831 169 3877 175
rect 3912 171 3925 181
rect 3943 171 3960 184
rect 3912 169 3960 171
rect 3793 163 3795 165
rect 3795 161 3797 163
rect 3797 160 3798 161
rect 3798 158 3807 160
rect 3780 151 3810 158
rect 3780 149 3811 151
rect 3831 149 3867 169
rect 3912 168 3959 169
rect 3925 163 3959 168
rect 3678 145 3867 149
rect 3693 142 3867 145
rect 3686 139 3867 142
rect 3895 162 3959 163
rect 3489 119 3508 121
rect 3523 119 3557 121
rect 3489 103 3569 119
rect 3489 97 3508 103
rect 2856 73 2891 81
rect 2856 47 2857 73
rect 2864 47 2891 73
rect 2856 39 2891 47
rect 2893 73 2934 81
rect 2893 47 2908 73
rect 2915 47 2934 73
rect 2998 69 3029 81
rect 3044 69 3147 81
rect 3159 71 3185 81
rect 3205 71 3308 81
rect 3159 69 3308 71
rect 3329 69 3364 81
rect 2998 67 3160 69
rect 3010 47 3029 67
rect 3044 65 3074 67
rect 2893 39 2934 47
rect 2856 29 2885 39
rect 2899 29 2928 39
rect 3016 29 3029 47
rect 3081 51 3160 67
rect 3192 67 3364 69
rect 3192 51 3271 67
rect 3278 65 3308 67
rect 3081 43 3271 51
rect 3336 47 3342 67
rect 3081 39 3160 43
rect 3162 39 3190 43
rect 3192 39 3271 43
rect 3066 29 3074 39
rect 3093 31 3096 39
rect 3097 31 3115 39
rect 3160 31 3192 39
rect 3237 31 3255 39
rect 3093 29 3259 31
rect 3278 29 3289 39
rect 3351 29 3364 67
rect 3436 81 3465 97
rect 3479 81 3508 97
rect 3523 87 3553 103
rect 3581 81 3587 129
rect 3590 123 3609 129
rect 3624 123 3654 131
rect 3590 115 3654 123
rect 3590 99 3670 115
rect 3686 108 3748 139
rect 3764 108 3826 139
rect 3895 137 3944 162
rect 3959 137 3989 153
rect 3858 123 3888 131
rect 3895 129 4005 137
rect 3858 115 3903 123
rect 3697 105 3701 108
rect 3702 105 3732 108
rect 3590 97 3609 99
rect 3624 97 3670 99
rect 3590 81 3670 97
rect 3701 95 3732 105
rect 3773 105 3779 108
rect 3780 105 3810 108
rect 3773 103 3815 105
rect 3702 92 3732 95
rect 3711 88 3718 92
rect 3718 87 3719 88
rect 3677 81 3687 87
rect 3739 81 3755 97
rect 3780 92 3810 103
rect 3842 99 3904 115
rect 3842 97 3888 99
rect 3842 81 3904 97
rect 3916 81 3922 129
rect 3925 121 4005 129
rect 3925 119 3944 121
rect 3959 119 3993 121
rect 3925 103 4005 119
rect 3925 81 3944 103
rect 3959 87 3989 103
rect 4017 97 4023 171
rect 4026 97 4045 241
rect 4060 97 4066 241
rect 4075 171 4088 241
rect 4140 237 4162 241
rect 4133 215 4162 229
rect 4215 215 4231 229
rect 4269 219 4275 227
rect 4282 225 4390 241
rect 4133 213 4231 215
rect 4117 205 4168 213
rect 4215 205 4249 213
rect 4117 193 4142 205
rect 4149 193 4168 205
rect 4222 203 4249 205
rect 4258 205 4275 219
rect 4320 205 4352 225
rect 4397 219 4403 227
rect 4411 219 4426 241
rect 4492 235 4511 238
rect 4397 213 4426 219
rect 4441 215 4457 229
rect 4492 216 4514 235
rect 4524 229 4540 230
rect 4523 227 4540 229
rect 4524 222 4540 227
rect 4514 215 4520 216
rect 4523 215 4552 222
rect 4441 214 4552 215
rect 4441 213 4558 214
rect 4397 205 4479 213
rect 4514 210 4520 213
rect 4258 203 4479 205
rect 4222 199 4294 203
rect 4322 201 4350 203
rect 4117 185 4168 193
rect 4215 191 4347 199
rect 4350 191 4361 199
rect 4215 189 4294 191
rect 4375 189 4479 203
rect 4523 205 4558 213
rect 4215 185 4312 189
rect 4069 137 4088 171
rect 4133 177 4162 185
rect 4133 171 4150 177
rect 4133 169 4167 171
rect 4215 169 4231 185
rect 4232 181 4312 185
rect 4360 185 4479 189
rect 4360 181 4440 185
rect 4232 175 4440 181
rect 4441 175 4457 185
rect 4505 181 4520 196
rect 4523 193 4524 205
rect 4531 193 4558 205
rect 4523 185 4558 193
rect 4523 184 4552 185
rect 4243 171 4353 175
rect 4134 165 4167 169
rect 4130 163 4167 165
rect 4130 162 4197 163
rect 4130 157 4161 162
rect 4167 157 4197 162
rect 4258 159 4273 171
rect 4130 153 4197 157
rect 4103 150 4197 153
rect 4103 143 4152 150
rect 4103 137 4133 143
rect 4152 138 4157 143
rect 4069 121 4149 137
rect 4161 129 4197 150
rect 4282 149 4312 158
rect 4335 153 4353 171
rect 4411 169 4457 175
rect 4492 171 4505 181
rect 4523 171 4540 184
rect 4492 169 4540 171
rect 4373 163 4375 165
rect 4375 161 4377 163
rect 4377 160 4378 161
rect 4378 158 4387 160
rect 4360 151 4390 158
rect 4360 149 4391 151
rect 4411 149 4447 169
rect 4492 168 4539 169
rect 4505 163 4539 168
rect 4258 145 4447 149
rect 4273 142 4447 145
rect 4266 139 4447 142
rect 4475 162 4539 163
rect 4069 119 4088 121
rect 4103 119 4137 121
rect 4069 103 4149 119
rect 4069 97 4088 103
rect 3436 73 3471 81
rect 3436 47 3437 73
rect 3444 47 3471 73
rect 3436 39 3471 47
rect 3473 73 3514 81
rect 3473 47 3488 73
rect 3495 47 3514 73
rect 3578 69 3609 81
rect 3624 69 3727 81
rect 3739 71 3765 81
rect 3785 71 3888 81
rect 3739 69 3888 71
rect 3909 69 3944 81
rect 3578 67 3740 69
rect 3590 47 3609 67
rect 3624 65 3654 67
rect 3473 39 3514 47
rect 3436 29 3465 39
rect 3479 29 3508 39
rect 3596 29 3609 47
rect 3661 51 3740 67
rect 3772 67 3944 69
rect 3772 51 3851 67
rect 3858 65 3888 67
rect 3661 43 3851 51
rect 3916 47 3922 67
rect 3661 39 3740 43
rect 3742 39 3770 43
rect 3772 39 3851 43
rect 3646 29 3654 39
rect 3673 31 3676 39
rect 3677 31 3695 39
rect 3740 31 3772 39
rect 3817 31 3835 39
rect 3673 29 3839 31
rect 3858 29 3869 39
rect 3931 29 3944 67
rect 4016 81 4045 97
rect 4059 81 4088 97
rect 4103 87 4133 103
rect 4161 81 4167 129
rect 4170 123 4189 129
rect 4204 123 4234 131
rect 4170 115 4234 123
rect 4170 99 4250 115
rect 4266 108 4328 139
rect 4344 108 4406 139
rect 4475 137 4524 162
rect 4539 137 4569 153
rect 4438 123 4468 131
rect 4475 129 4585 137
rect 4438 115 4483 123
rect 4277 105 4281 108
rect 4282 105 4312 108
rect 4170 97 4189 99
rect 4204 97 4250 99
rect 4170 81 4250 97
rect 4281 95 4312 105
rect 4353 105 4359 108
rect 4360 105 4390 108
rect 4353 103 4395 105
rect 4282 92 4312 95
rect 4291 88 4298 92
rect 4298 87 4299 88
rect 4257 81 4267 87
rect 4319 81 4335 97
rect 4360 92 4390 103
rect 4422 99 4484 115
rect 4422 97 4468 99
rect 4422 81 4484 97
rect 4496 81 4502 129
rect 4505 121 4585 129
rect 4505 119 4524 121
rect 4539 119 4573 121
rect 4505 103 4585 119
rect 4505 81 4524 103
rect 4539 87 4569 103
rect 4597 97 4603 171
rect 4606 97 4625 241
rect 4640 97 4646 241
rect 4655 171 4668 241
rect 4720 237 4742 241
rect 4713 215 4742 229
rect 4795 215 4811 229
rect 4849 219 4855 227
rect 4862 225 4970 241
rect 4713 213 4811 215
rect 4697 205 4748 213
rect 4795 205 4829 213
rect 4697 193 4722 205
rect 4729 193 4748 205
rect 4802 203 4829 205
rect 4838 205 4855 219
rect 4900 205 4932 225
rect 4977 219 4983 227
rect 4991 219 5006 241
rect 5072 235 5091 238
rect 4977 213 5006 219
rect 5021 215 5037 229
rect 5072 216 5094 235
rect 5104 229 5120 230
rect 5103 227 5120 229
rect 5104 222 5120 227
rect 5094 215 5100 216
rect 5103 215 5132 222
rect 5021 214 5132 215
rect 5021 213 5138 214
rect 4977 205 5059 213
rect 5094 210 5100 213
rect 4838 203 5059 205
rect 4802 199 4874 203
rect 4902 201 4930 203
rect 4697 185 4748 193
rect 4795 191 4927 199
rect 4930 191 4942 199
rect 4795 189 4874 191
rect 4955 189 5059 203
rect 4795 185 4892 189
rect 4649 137 4668 171
rect 4713 177 4742 185
rect 4713 171 4730 177
rect 4713 169 4747 171
rect 4795 169 4811 185
rect 4812 181 4892 185
rect 4940 185 5059 189
rect 4940 181 5020 185
rect 4812 175 5020 181
rect 5021 175 5037 185
rect 5085 181 5100 196
rect 5103 184 5138 213
rect 4823 171 4933 175
rect 4714 165 4747 169
rect 4710 163 4747 165
rect 4710 162 4777 163
rect 4710 157 4741 162
rect 4747 157 4777 162
rect 4838 159 4853 171
rect 4710 153 4777 157
rect 4683 150 4777 153
rect 4683 143 4732 150
rect 4683 137 4713 143
rect 4732 138 4737 143
rect 4649 121 4729 137
rect 4741 129 4777 150
rect 4862 149 4892 158
rect 4915 153 4933 171
rect 4991 169 5037 175
rect 5072 171 5085 181
rect 5103 171 5120 184
rect 4953 163 4955 165
rect 4955 160 4958 163
rect 4958 158 4967 160
rect 4940 151 4970 158
rect 4940 149 4971 151
rect 4991 149 5027 169
rect 5072 168 5120 171
rect 5085 163 5119 168
rect 4838 145 5027 149
rect 4853 142 5027 145
rect 4846 139 5027 142
rect 5055 162 5119 163
rect 4649 119 4668 121
rect 4683 119 4717 121
rect 4649 103 4729 119
rect 4649 97 4668 103
rect 4016 73 4051 81
rect 4016 47 4017 73
rect 4024 47 4051 73
rect 4016 39 4051 47
rect 4053 73 4094 81
rect 4053 47 4068 73
rect 4075 47 4094 73
rect 4158 69 4189 81
rect 4204 69 4307 81
rect 4319 71 4345 81
rect 4365 71 4468 81
rect 4319 69 4468 71
rect 4489 69 4524 81
rect 4158 67 4320 69
rect 4170 47 4189 67
rect 4204 65 4234 67
rect 4053 39 4094 47
rect 4016 29 4045 39
rect 4059 29 4088 39
rect 4176 29 4189 47
rect 4241 51 4320 67
rect 4352 67 4524 69
rect 4352 51 4431 67
rect 4438 65 4468 67
rect 4241 43 4431 51
rect 4496 47 4502 67
rect 4241 39 4320 43
rect 4322 39 4350 43
rect 4352 39 4431 43
rect 4226 29 4234 39
rect 4253 31 4256 39
rect 4257 31 4275 39
rect 4320 31 4352 39
rect 4397 31 4415 39
rect 4253 29 4419 31
rect 4438 29 4449 39
rect 4511 29 4524 67
rect 4596 81 4625 97
rect 4639 81 4668 97
rect 4683 87 4713 103
rect 4741 81 4747 129
rect 4750 123 4769 129
rect 4784 123 4814 131
rect 4750 115 4814 123
rect 4750 99 4830 115
rect 4846 108 4908 139
rect 4924 108 4986 139
rect 5055 137 5104 162
rect 5119 137 5149 153
rect 5018 123 5048 131
rect 5055 129 5165 137
rect 5018 115 5063 123
rect 4857 104 4892 108
rect 4750 97 4769 99
rect 4784 97 4830 99
rect 4750 81 4830 97
rect 4862 92 4892 104
rect 4933 105 4970 108
rect 4933 103 4975 105
rect 4871 88 4878 92
rect 4878 87 4879 88
rect 4837 81 4847 87
rect 4596 73 4631 81
rect 4596 47 4597 73
rect 4604 47 4631 73
rect 4596 39 4631 47
rect 4633 73 4674 81
rect 4633 47 4648 73
rect 4655 47 4674 73
rect 4738 69 4769 81
rect 4784 69 4887 81
rect 4899 80 4916 97
rect 4940 92 4970 103
rect 5002 99 5064 115
rect 5002 97 5048 99
rect 5002 81 5064 97
rect 5076 81 5082 129
rect 5085 121 5165 129
rect 5085 119 5104 121
rect 5119 119 5153 121
rect 5085 103 5165 119
rect 5085 81 5104 103
rect 5119 87 5149 103
rect 5177 97 5183 171
rect 5186 97 5205 241
rect 5220 97 5226 241
rect 5235 171 5248 241
rect 5300 237 5322 241
rect 5293 215 5322 229
rect 5375 215 5391 229
rect 5429 219 5435 227
rect 5442 225 5550 241
rect 5279 213 5391 215
rect 5277 185 5328 213
rect 5375 205 5409 213
rect 5382 203 5409 205
rect 5418 205 5435 219
rect 5480 205 5512 225
rect 5557 219 5563 227
rect 5571 219 5586 241
rect 5652 235 5671 238
rect 5557 213 5586 219
rect 5601 215 5617 229
rect 5652 216 5674 235
rect 5684 229 5700 230
rect 5683 227 5700 229
rect 5684 222 5700 227
rect 5674 215 5680 216
rect 5683 215 5712 222
rect 5601 214 5712 215
rect 5601 213 5718 214
rect 5557 205 5639 213
rect 5674 210 5680 213
rect 5418 203 5639 205
rect 5382 199 5454 203
rect 5482 201 5510 203
rect 5229 137 5248 171
rect 5293 184 5328 185
rect 5375 191 5507 199
rect 5510 191 5522 199
rect 5375 189 5454 191
rect 5535 189 5639 203
rect 5375 185 5472 189
rect 5293 177 5322 184
rect 5293 171 5310 177
rect 5293 168 5327 171
rect 5375 169 5391 185
rect 5392 181 5472 185
rect 5520 185 5639 189
rect 5520 181 5600 185
rect 5392 175 5600 181
rect 5601 175 5617 185
rect 5665 181 5680 196
rect 5683 184 5718 213
rect 5403 171 5513 175
rect 5294 165 5327 168
rect 5290 163 5327 165
rect 5290 162 5357 163
rect 5290 157 5321 162
rect 5327 157 5357 162
rect 5418 159 5433 171
rect 5290 153 5357 157
rect 5263 150 5357 153
rect 5263 143 5312 150
rect 5263 137 5293 143
rect 5312 138 5317 143
rect 5229 121 5309 137
rect 5321 129 5357 150
rect 5442 149 5472 158
rect 5495 153 5513 171
rect 5571 169 5617 175
rect 5652 171 5665 181
rect 5683 171 5700 184
rect 5533 163 5535 165
rect 5535 160 5538 163
rect 5538 158 5547 160
rect 5520 151 5550 158
rect 5520 149 5551 151
rect 5571 149 5607 169
rect 5652 168 5700 171
rect 5665 163 5699 168
rect 5418 145 5607 149
rect 5433 142 5607 145
rect 5426 139 5607 142
rect 5635 162 5699 163
rect 5229 119 5248 121
rect 5263 119 5297 121
rect 5229 103 5309 119
rect 5229 97 5248 103
rect 4899 71 4925 80
rect 4945 71 5048 81
rect 4899 69 5048 71
rect 5069 69 5104 81
rect 4738 67 4900 69
rect 4750 47 4769 67
rect 4784 65 4814 67
rect 4633 39 4674 47
rect 4596 29 4625 39
rect 4639 29 4668 39
rect 4756 29 4769 47
rect 4821 51 4900 67
rect 4932 67 5104 69
rect 4932 51 5011 67
rect 5018 65 5048 67
rect 4821 43 5011 51
rect 5076 47 5082 67
rect 4821 39 4900 43
rect 4902 39 4930 43
rect 4932 39 5011 43
rect 4806 29 4814 39
rect 4833 31 4836 39
rect 4837 31 4855 39
rect 4900 31 4932 39
rect 4977 31 4995 39
rect 4833 29 4999 31
rect 5018 29 5029 39
rect 5091 29 5104 67
rect 5176 81 5205 97
rect 5219 81 5248 97
rect 5263 87 5293 103
rect 5321 81 5327 129
rect 5330 123 5349 129
rect 5364 123 5394 131
rect 5330 115 5394 123
rect 5330 99 5410 115
rect 5426 108 5488 139
rect 5504 108 5566 139
rect 5635 137 5684 162
rect 5699 137 5729 153
rect 5598 123 5628 131
rect 5635 129 5745 137
rect 5598 115 5643 123
rect 5437 104 5472 108
rect 5330 97 5349 99
rect 5364 97 5410 99
rect 5330 81 5410 97
rect 5442 92 5472 104
rect 5513 105 5550 108
rect 5513 103 5555 105
rect 5451 88 5458 92
rect 5458 87 5459 88
rect 5417 81 5427 87
rect 5176 69 5211 81
rect 5213 69 5254 81
rect 5176 39 5254 69
rect 5318 69 5349 81
rect 5364 69 5467 81
rect 5479 80 5496 97
rect 5520 92 5550 103
rect 5582 99 5644 115
rect 5582 97 5628 99
rect 5582 81 5644 97
rect 5656 81 5662 129
rect 5665 121 5745 129
rect 5665 119 5684 121
rect 5699 119 5733 121
rect 5665 103 5745 119
rect 5665 81 5684 103
rect 5699 87 5729 103
rect 5757 97 5763 171
rect 5766 97 5785 241
rect 5800 97 5806 241
rect 5815 171 5828 241
rect 5880 237 5902 241
rect 5873 215 5902 229
rect 5955 215 5971 229
rect 6009 219 6015 227
rect 6022 225 6130 241
rect 5859 213 5971 215
rect 5857 185 5908 213
rect 5955 205 5989 213
rect 5962 203 5989 205
rect 5998 205 6015 219
rect 6060 205 6092 225
rect 6137 219 6143 227
rect 6151 219 6166 241
rect 6232 235 6251 238
rect 6137 213 6166 219
rect 6181 215 6197 229
rect 6232 216 6254 235
rect 6264 229 6280 230
rect 6263 227 6280 229
rect 6264 222 6280 227
rect 6254 215 6260 216
rect 6263 215 6292 222
rect 6181 214 6292 215
rect 6181 213 6298 214
rect 6137 205 6219 213
rect 6254 210 6260 213
rect 5998 203 6219 205
rect 5962 199 6034 203
rect 6062 201 6090 203
rect 5809 137 5828 171
rect 5873 184 5908 185
rect 5955 191 6087 199
rect 6090 191 6102 199
rect 5955 189 6034 191
rect 6115 189 6219 203
rect 5955 185 6052 189
rect 5873 177 5902 184
rect 5873 171 5890 177
rect 5873 168 5907 171
rect 5955 169 5971 185
rect 5972 181 6052 185
rect 6100 185 6219 189
rect 6100 181 6180 185
rect 5972 175 6180 181
rect 6181 175 6197 185
rect 6245 181 6260 196
rect 6263 184 6298 213
rect 5983 171 6093 175
rect 5874 165 5907 168
rect 5870 163 5907 165
rect 5870 162 5937 163
rect 5870 157 5901 162
rect 5907 157 5937 162
rect 5998 159 6013 171
rect 5870 153 5937 157
rect 5843 150 5937 153
rect 5843 143 5892 150
rect 5843 137 5873 143
rect 5892 138 5897 143
rect 5809 121 5889 137
rect 5901 129 5937 150
rect 6022 149 6052 158
rect 6075 153 6093 171
rect 6151 169 6197 175
rect 6232 171 6245 181
rect 6263 171 6280 184
rect 6113 163 6115 165
rect 6115 160 6118 163
rect 6118 158 6127 160
rect 6100 151 6130 158
rect 6100 149 6131 151
rect 6151 149 6187 169
rect 6232 168 6280 171
rect 6245 163 6279 168
rect 5998 145 6187 149
rect 6013 142 6187 145
rect 6006 139 6187 142
rect 6215 162 6279 163
rect 5809 119 5828 121
rect 5843 119 5877 121
rect 5809 103 5889 119
rect 5809 97 5828 103
rect 5479 71 5505 80
rect 5525 71 5628 81
rect 5479 69 5628 71
rect 5649 69 5684 81
rect 5318 67 5480 69
rect 5330 47 5349 67
rect 5364 65 5394 67
rect 5176 38 5211 39
rect 5219 38 5254 39
rect 5176 29 5205 38
rect 5219 29 5248 38
rect 5336 29 5349 47
rect 5401 51 5480 67
rect 5512 67 5684 69
rect 5512 51 5591 67
rect 5598 65 5628 67
rect 5401 43 5591 51
rect 5656 47 5662 67
rect 5401 39 5480 43
rect 5482 39 5510 43
rect 5512 39 5591 43
rect 5386 29 5394 39
rect 5413 31 5416 39
rect 5417 31 5435 39
rect 5480 31 5512 39
rect 5557 31 5575 39
rect 5413 29 5579 31
rect 5598 29 5609 39
rect 5671 29 5684 67
rect 5756 81 5785 97
rect 5799 81 5828 97
rect 5843 87 5873 103
rect 5901 81 5907 129
rect 5910 123 5929 129
rect 5944 123 5974 131
rect 5910 115 5974 123
rect 5910 99 5990 115
rect 6006 108 6068 139
rect 6084 108 6146 139
rect 6215 137 6264 162
rect 6279 137 6309 153
rect 6178 123 6208 131
rect 6215 129 6325 137
rect 6178 115 6223 123
rect 6017 104 6052 108
rect 5910 97 5929 99
rect 5944 97 5990 99
rect 5910 81 5990 97
rect 6022 92 6052 104
rect 6093 105 6130 108
rect 6093 103 6135 105
rect 6031 88 6038 92
rect 6038 87 6039 88
rect 5997 81 6007 87
rect 5756 69 5791 81
rect 5793 69 5834 81
rect 5756 39 5834 69
rect 5898 69 5929 81
rect 5944 69 6047 81
rect 6059 80 6076 97
rect 6100 92 6130 103
rect 6162 99 6224 115
rect 6162 97 6208 99
rect 6162 81 6224 97
rect 6236 81 6242 129
rect 6245 121 6325 129
rect 6245 119 6264 121
rect 6279 119 6313 121
rect 6245 103 6325 119
rect 6245 81 6264 103
rect 6279 87 6309 103
rect 6337 97 6343 171
rect 6346 97 6365 241
rect 6380 97 6386 241
rect 6395 171 6408 241
rect 6460 237 6482 241
rect 6453 215 6482 229
rect 6535 215 6551 229
rect 6589 219 6595 227
rect 6602 225 6710 241
rect 6439 213 6551 215
rect 6437 185 6488 213
rect 6535 205 6569 213
rect 6542 203 6569 205
rect 6578 205 6595 219
rect 6640 205 6672 225
rect 6717 219 6723 227
rect 6731 219 6746 241
rect 6812 235 6831 238
rect 6717 213 6746 219
rect 6761 215 6777 229
rect 6812 216 6834 235
rect 6844 229 6860 230
rect 6843 227 6860 229
rect 6844 222 6860 227
rect 6834 215 6840 216
rect 6843 215 6872 222
rect 6761 214 6872 215
rect 6761 213 6878 214
rect 6717 205 6799 213
rect 6834 210 6840 213
rect 6578 203 6799 205
rect 6542 199 6614 203
rect 6642 201 6670 203
rect 6389 137 6408 171
rect 6453 184 6488 185
rect 6535 191 6667 199
rect 6670 191 6682 199
rect 6535 189 6614 191
rect 6695 189 6799 203
rect 6535 185 6632 189
rect 6453 177 6482 184
rect 6453 171 6470 177
rect 6453 168 6487 171
rect 6535 169 6551 185
rect 6552 181 6632 185
rect 6680 185 6799 189
rect 6680 181 6760 185
rect 6552 175 6760 181
rect 6761 175 6777 185
rect 6825 181 6840 196
rect 6843 184 6878 213
rect 6563 171 6673 175
rect 6454 165 6487 168
rect 6450 163 6487 165
rect 6450 162 6517 163
rect 6450 157 6481 162
rect 6487 157 6517 162
rect 6578 159 6593 171
rect 6450 153 6517 157
rect 6423 150 6517 153
rect 6423 143 6472 150
rect 6423 137 6453 143
rect 6472 138 6477 143
rect 6389 121 6469 137
rect 6481 129 6517 150
rect 6602 149 6632 158
rect 6655 153 6673 171
rect 6731 169 6777 175
rect 6812 171 6825 181
rect 6843 171 6860 184
rect 6693 163 6695 165
rect 6695 160 6698 163
rect 6698 158 6707 160
rect 6680 151 6710 158
rect 6680 149 6711 151
rect 6731 149 6767 169
rect 6812 168 6860 171
rect 6825 163 6859 168
rect 6578 145 6767 149
rect 6593 142 6767 145
rect 6586 139 6767 142
rect 6795 162 6859 163
rect 6389 119 6408 121
rect 6423 119 6457 121
rect 6389 103 6469 119
rect 6389 97 6408 103
rect 6059 71 6085 80
rect 6105 71 6208 81
rect 6059 69 6208 71
rect 6229 69 6264 81
rect 5898 67 6060 69
rect 5910 47 5929 67
rect 5944 65 5974 67
rect 5756 38 5791 39
rect 5799 38 5834 39
rect 5756 29 5785 38
rect 5799 29 5828 38
rect 5916 29 5929 47
rect 5981 51 6060 67
rect 6092 67 6264 69
rect 6092 51 6171 67
rect 6178 65 6208 67
rect 5981 43 6171 51
rect 6236 47 6242 67
rect 5981 39 6060 43
rect 6062 39 6090 43
rect 6092 39 6171 43
rect 5966 29 5974 39
rect 5993 31 5996 39
rect 5997 31 6015 39
rect 6060 31 6092 39
rect 6137 31 6155 39
rect 5993 29 6159 31
rect 6178 29 6189 39
rect 6251 29 6264 67
rect 6336 81 6365 97
rect 6379 81 6408 97
rect 6423 87 6453 103
rect 6481 81 6487 129
rect 6490 123 6509 129
rect 6524 123 6554 131
rect 6490 115 6554 123
rect 6490 99 6570 115
rect 6586 108 6648 139
rect 6664 108 6726 139
rect 6795 137 6844 162
rect 6859 137 6889 153
rect 6758 123 6788 131
rect 6795 129 6905 137
rect 6758 115 6803 123
rect 6597 104 6632 108
rect 6490 97 6509 99
rect 6524 97 6570 99
rect 6490 81 6570 97
rect 6602 92 6632 104
rect 6673 105 6710 108
rect 6673 103 6715 105
rect 6611 88 6618 92
rect 6618 87 6619 88
rect 6577 81 6587 87
rect 6336 69 6371 81
rect 6373 69 6414 81
rect 6336 39 6414 69
rect 6478 69 6509 81
rect 6524 69 6627 81
rect 6639 80 6656 97
rect 6680 92 6710 103
rect 6742 99 6804 115
rect 6742 97 6788 99
rect 6742 81 6804 97
rect 6816 81 6822 129
rect 6825 121 6905 129
rect 6825 119 6844 121
rect 6859 119 6893 121
rect 6825 103 6905 119
rect 6825 81 6844 103
rect 6859 87 6889 103
rect 6917 97 6923 171
rect 6926 97 6945 241
rect 6960 97 6966 241
rect 6975 171 6988 241
rect 7040 237 7062 241
rect 7033 215 7062 229
rect 7115 215 7131 229
rect 7169 219 7175 227
rect 7182 225 7290 241
rect 7019 213 7131 215
rect 7017 185 7068 213
rect 7115 205 7149 213
rect 7122 203 7149 205
rect 7158 205 7175 219
rect 7220 205 7252 225
rect 7297 219 7303 227
rect 7311 219 7326 241
rect 7392 235 7411 238
rect 7297 213 7326 219
rect 7341 215 7357 229
rect 7392 216 7414 235
rect 7424 229 7440 230
rect 7423 227 7440 229
rect 7424 222 7440 227
rect 7414 215 7420 216
rect 7423 215 7452 222
rect 7341 214 7452 215
rect 7341 213 7458 214
rect 7297 205 7379 213
rect 7414 210 7420 213
rect 7158 203 7379 205
rect 7122 199 7194 203
rect 7222 201 7250 203
rect 6969 137 6988 171
rect 7033 184 7068 185
rect 7115 191 7247 199
rect 7250 191 7262 199
rect 7115 189 7194 191
rect 7275 189 7379 203
rect 7115 185 7212 189
rect 7033 177 7062 184
rect 7033 171 7050 177
rect 7033 168 7067 171
rect 7115 169 7131 185
rect 7132 181 7212 185
rect 7260 185 7379 189
rect 7260 181 7340 185
rect 7132 175 7340 181
rect 7341 175 7357 185
rect 7405 181 7420 196
rect 7423 184 7458 213
rect 7143 171 7253 175
rect 7034 165 7067 168
rect 7030 163 7067 165
rect 7030 162 7097 163
rect 7030 157 7061 162
rect 7067 157 7097 162
rect 7158 159 7173 171
rect 7030 153 7097 157
rect 7003 150 7097 153
rect 7003 143 7052 150
rect 7003 137 7033 143
rect 7052 138 7057 143
rect 6969 121 7049 137
rect 7061 129 7097 150
rect 7182 149 7212 158
rect 7235 153 7253 171
rect 7311 169 7357 175
rect 7392 171 7405 181
rect 7423 171 7440 184
rect 7273 163 7275 165
rect 7275 160 7278 163
rect 7278 158 7287 160
rect 7260 151 7290 158
rect 7260 149 7291 151
rect 7311 149 7347 169
rect 7392 168 7440 171
rect 7405 163 7439 168
rect 7158 145 7347 149
rect 7173 142 7347 145
rect 7166 139 7347 142
rect 7375 162 7439 163
rect 6969 119 6988 121
rect 7003 119 7037 121
rect 6969 103 7049 119
rect 6969 97 6988 103
rect 6639 71 6665 80
rect 6685 71 6788 81
rect 6639 69 6788 71
rect 6809 69 6844 81
rect 6478 67 6640 69
rect 6490 47 6509 67
rect 6524 65 6554 67
rect 6336 38 6371 39
rect 6379 38 6414 39
rect 6336 29 6365 38
rect 6379 29 6408 38
rect 6496 29 6509 47
rect 6561 51 6640 67
rect 6672 67 6844 69
rect 6672 51 6751 67
rect 6758 65 6788 67
rect 6561 43 6751 51
rect 6816 47 6822 67
rect 6561 39 6640 43
rect 6642 39 6670 43
rect 6672 39 6751 43
rect 6546 29 6554 39
rect 6573 31 6576 39
rect 6577 31 6595 39
rect 6640 31 6672 39
rect 6717 31 6735 39
rect 6573 29 6739 31
rect 6758 29 6769 39
rect 6831 29 6844 67
rect 6916 81 6945 97
rect 6959 81 6988 97
rect 7003 87 7033 103
rect 7061 81 7067 129
rect 7070 123 7089 129
rect 7104 123 7134 131
rect 7070 115 7134 123
rect 7070 99 7150 115
rect 7166 108 7228 139
rect 7244 108 7306 139
rect 7375 137 7424 162
rect 7439 137 7469 153
rect 7338 123 7368 131
rect 7375 129 7485 137
rect 7338 115 7383 123
rect 7177 104 7212 108
rect 7070 97 7089 99
rect 7104 97 7150 99
rect 7070 81 7150 97
rect 7182 92 7212 104
rect 7253 105 7290 108
rect 7253 103 7295 105
rect 7191 88 7198 92
rect 7198 87 7199 88
rect 7157 81 7167 87
rect 6916 69 6951 81
rect 6953 69 6994 81
rect 6916 39 6994 69
rect 7058 69 7089 81
rect 7104 69 7207 81
rect 7219 80 7236 97
rect 7260 92 7290 103
rect 7322 99 7384 115
rect 7322 97 7368 99
rect 7322 81 7384 97
rect 7396 81 7402 129
rect 7405 121 7485 129
rect 7405 119 7424 121
rect 7439 119 7473 121
rect 7405 103 7485 119
rect 7405 81 7424 103
rect 7439 87 7469 103
rect 7497 97 7503 171
rect 7506 97 7525 241
rect 7540 97 7546 241
rect 7555 171 7568 241
rect 7620 237 7642 241
rect 7613 215 7642 229
rect 7695 215 7711 229
rect 7749 219 7755 227
rect 7762 225 7870 241
rect 7599 213 7711 215
rect 7597 185 7648 213
rect 7695 205 7729 213
rect 7702 203 7729 205
rect 7738 205 7755 219
rect 7800 205 7832 225
rect 7877 219 7883 227
rect 7891 219 7906 241
rect 7972 235 7991 238
rect 7877 213 7906 219
rect 7921 215 7937 229
rect 7972 216 7994 235
rect 8004 229 8020 230
rect 8003 227 8020 229
rect 8004 222 8020 227
rect 7994 215 8000 216
rect 8003 215 8032 222
rect 7921 214 8032 215
rect 7921 213 8038 214
rect 7877 205 7959 213
rect 7994 210 8000 213
rect 7738 203 7959 205
rect 7702 199 7774 203
rect 7802 201 7830 203
rect 7549 137 7568 171
rect 7613 184 7648 185
rect 7695 191 7827 199
rect 7830 191 7842 199
rect 7695 189 7774 191
rect 7855 189 7959 203
rect 7695 185 7792 189
rect 7613 177 7642 184
rect 7613 171 7630 177
rect 7613 168 7647 171
rect 7695 169 7711 185
rect 7712 181 7792 185
rect 7840 185 7959 189
rect 7840 181 7920 185
rect 7712 175 7920 181
rect 7921 175 7937 185
rect 7985 181 8000 196
rect 8003 184 8038 213
rect 7723 171 7833 175
rect 7614 165 7647 168
rect 7610 163 7647 165
rect 7610 162 7677 163
rect 7610 157 7641 162
rect 7647 157 7677 162
rect 7738 159 7753 171
rect 7610 153 7677 157
rect 7583 150 7677 153
rect 7583 143 7632 150
rect 7583 137 7613 143
rect 7632 138 7637 143
rect 7549 121 7629 137
rect 7641 129 7677 150
rect 7762 149 7792 158
rect 7815 153 7833 171
rect 7891 169 7937 175
rect 7972 171 7985 181
rect 8003 171 8020 184
rect 7853 163 7855 165
rect 7855 160 7858 163
rect 7858 158 7867 160
rect 7840 151 7870 158
rect 7840 149 7871 151
rect 7891 149 7927 169
rect 7972 168 8020 171
rect 7985 163 8019 168
rect 7738 145 7927 149
rect 7753 142 7927 145
rect 7746 139 7927 142
rect 7955 162 8019 163
rect 7549 119 7568 121
rect 7583 119 7617 121
rect 7549 103 7629 119
rect 7549 97 7568 103
rect 7219 71 7245 80
rect 7265 71 7368 81
rect 7219 69 7368 71
rect 7389 69 7424 81
rect 7058 67 7220 69
rect 7070 47 7089 67
rect 7104 65 7134 67
rect 6916 38 6951 39
rect 6959 38 6994 39
rect 6916 29 6945 38
rect 6959 29 6988 38
rect 7076 29 7089 47
rect 7141 51 7220 67
rect 7252 67 7424 69
rect 7252 51 7331 67
rect 7338 65 7368 67
rect 7141 43 7331 51
rect 7396 47 7402 67
rect 7141 39 7220 43
rect 7222 39 7250 43
rect 7252 39 7331 43
rect 7126 29 7134 39
rect 7153 31 7156 39
rect 7157 31 7175 39
rect 7220 31 7252 39
rect 7297 31 7315 39
rect 7153 29 7319 31
rect 7338 29 7349 39
rect 7411 29 7424 67
rect 7496 81 7525 97
rect 7539 81 7568 97
rect 7583 87 7613 103
rect 7641 81 7647 129
rect 7650 123 7669 129
rect 7684 123 7714 131
rect 7650 115 7714 123
rect 7650 99 7730 115
rect 7746 108 7808 139
rect 7824 108 7886 139
rect 7955 137 8004 162
rect 8019 137 8049 153
rect 7918 123 7948 131
rect 7955 129 8065 137
rect 7918 115 7963 123
rect 7757 104 7792 108
rect 7650 97 7669 99
rect 7684 97 7730 99
rect 7650 81 7730 97
rect 7762 92 7792 104
rect 7833 105 7870 108
rect 7833 103 7875 105
rect 7771 88 7778 92
rect 7778 87 7779 88
rect 7737 81 7747 87
rect 7496 69 7531 81
rect 7533 69 7574 81
rect 7496 39 7574 69
rect 7638 69 7669 81
rect 7684 69 7787 81
rect 7799 80 7816 97
rect 7840 92 7870 103
rect 7902 99 7964 115
rect 7902 97 7948 99
rect 7902 81 7964 97
rect 7976 81 7982 129
rect 7985 121 8065 129
rect 7985 119 8004 121
rect 8019 119 8053 121
rect 7985 103 8065 119
rect 7985 81 8004 103
rect 8019 87 8049 103
rect 8077 97 8083 171
rect 8086 97 8105 241
rect 8120 97 8126 241
rect 8135 171 8148 241
rect 8200 237 8222 241
rect 8193 215 8222 229
rect 8275 215 8291 229
rect 8329 219 8335 227
rect 8342 225 8450 241
rect 8179 213 8291 215
rect 8177 185 8228 213
rect 8275 205 8309 213
rect 8282 203 8309 205
rect 8318 205 8335 219
rect 8380 205 8412 225
rect 8457 219 8463 227
rect 8471 219 8486 241
rect 8552 235 8571 238
rect 8457 213 8486 219
rect 8501 215 8517 229
rect 8552 216 8574 235
rect 8584 229 8600 230
rect 8583 227 8600 229
rect 8584 222 8600 227
rect 8574 215 8580 216
rect 8583 215 8612 222
rect 8501 214 8612 215
rect 8501 213 8618 214
rect 8457 205 8539 213
rect 8574 210 8580 213
rect 8318 203 8539 205
rect 8282 199 8354 203
rect 8382 201 8410 203
rect 8129 137 8148 171
rect 8193 184 8228 185
rect 8275 191 8407 199
rect 8410 191 8422 199
rect 8275 189 8354 191
rect 8435 189 8539 203
rect 8275 185 8372 189
rect 8193 177 8222 184
rect 8193 171 8210 177
rect 8193 168 8227 171
rect 8275 169 8291 185
rect 8292 181 8372 185
rect 8420 185 8539 189
rect 8420 181 8500 185
rect 8292 175 8500 181
rect 8501 175 8517 185
rect 8565 181 8580 196
rect 8583 184 8618 213
rect 8303 171 8413 175
rect 8194 165 8227 168
rect 8190 163 8227 165
rect 8190 162 8257 163
rect 8190 157 8221 162
rect 8227 157 8257 162
rect 8318 159 8333 171
rect 8190 153 8257 157
rect 8163 150 8257 153
rect 8163 143 8212 150
rect 8163 137 8193 143
rect 8212 138 8217 143
rect 8129 121 8209 137
rect 8221 129 8257 150
rect 8342 149 8372 158
rect 8395 153 8413 171
rect 8471 169 8517 175
rect 8552 171 8565 181
rect 8583 171 8600 184
rect 8433 163 8435 165
rect 8435 160 8438 163
rect 8438 158 8447 160
rect 8420 151 8450 158
rect 8420 149 8451 151
rect 8471 149 8507 169
rect 8552 168 8600 171
rect 8565 163 8599 168
rect 8318 145 8507 149
rect 8333 142 8507 145
rect 8326 139 8507 142
rect 8535 162 8599 163
rect 8129 119 8148 121
rect 8163 119 8197 121
rect 8129 103 8209 119
rect 8129 97 8148 103
rect 7799 71 7825 80
rect 7845 71 7948 81
rect 7799 69 7948 71
rect 7969 69 8004 81
rect 7638 67 7800 69
rect 7650 47 7669 67
rect 7684 65 7714 67
rect 7496 38 7531 39
rect 7539 38 7574 39
rect 7496 29 7525 38
rect 7539 29 7568 38
rect 7656 29 7669 47
rect 7721 51 7800 67
rect 7832 67 8004 69
rect 7832 51 7911 67
rect 7918 65 7948 67
rect 7721 43 7911 51
rect 7976 47 7982 67
rect 7721 39 7800 43
rect 7802 39 7830 43
rect 7832 39 7911 43
rect 7706 29 7714 39
rect 7733 31 7736 39
rect 7737 31 7755 39
rect 7800 31 7832 39
rect 7877 31 7895 39
rect 7733 29 7899 31
rect 7918 29 7929 39
rect 7991 29 8004 67
rect 8076 81 8105 97
rect 8119 81 8148 97
rect 8163 87 8193 103
rect 8221 81 8227 129
rect 8230 123 8249 129
rect 8264 123 8294 131
rect 8230 115 8294 123
rect 8230 99 8310 115
rect 8326 108 8388 139
rect 8404 108 8466 139
rect 8535 137 8584 162
rect 8599 137 8629 153
rect 8498 123 8528 131
rect 8535 129 8645 137
rect 8498 115 8543 123
rect 8337 104 8372 108
rect 8230 97 8249 99
rect 8264 97 8310 99
rect 8230 81 8310 97
rect 8342 92 8372 104
rect 8413 105 8450 108
rect 8413 103 8455 105
rect 8351 88 8358 92
rect 8358 87 8359 88
rect 8317 81 8327 87
rect 8076 69 8111 81
rect 8113 69 8154 81
rect 8076 39 8154 69
rect 8218 69 8249 81
rect 8264 69 8367 81
rect 8379 80 8396 97
rect 8420 92 8450 103
rect 8482 99 8544 115
rect 8482 97 8528 99
rect 8482 81 8544 97
rect 8556 81 8562 129
rect 8565 121 8645 129
rect 8565 119 8584 121
rect 8599 119 8633 121
rect 8565 103 8645 119
rect 8565 81 8584 103
rect 8599 87 8629 103
rect 8657 97 8663 171
rect 8666 97 8685 241
rect 8700 97 8706 241
rect 8715 171 8728 241
rect 8780 237 8802 241
rect 8773 215 8802 229
rect 8855 215 8871 229
rect 8909 219 8915 227
rect 8922 225 9030 241
rect 8759 213 8871 215
rect 8757 185 8808 213
rect 8855 205 8889 213
rect 8862 203 8889 205
rect 8898 205 8915 219
rect 8960 205 8992 225
rect 9037 219 9043 227
rect 9051 219 9066 241
rect 9132 235 9151 238
rect 9037 213 9066 219
rect 9081 215 9097 229
rect 9132 216 9154 235
rect 9164 229 9180 230
rect 9163 227 9180 229
rect 9164 222 9180 227
rect 9154 215 9160 216
rect 9163 215 9192 222
rect 9081 214 9192 215
rect 9081 213 9198 214
rect 9037 205 9119 213
rect 9154 210 9160 213
rect 8898 203 9119 205
rect 8862 199 8934 203
rect 8962 201 8990 203
rect 8709 137 8728 171
rect 8773 184 8808 185
rect 8855 191 8987 199
rect 8990 191 9002 199
rect 8855 189 8934 191
rect 9015 189 9119 203
rect 8855 185 8952 189
rect 8773 177 8802 184
rect 8773 171 8790 177
rect 8773 168 8807 171
rect 8855 169 8871 185
rect 8872 181 8952 185
rect 9000 185 9119 189
rect 9000 181 9080 185
rect 8872 175 9080 181
rect 9081 175 9097 185
rect 9145 181 9160 196
rect 9163 184 9198 213
rect 8883 171 8993 175
rect 8774 165 8807 168
rect 8770 163 8807 165
rect 8770 162 8837 163
rect 8770 157 8801 162
rect 8807 157 8837 162
rect 8898 159 8913 171
rect 8770 153 8837 157
rect 8743 150 8837 153
rect 8743 143 8792 150
rect 8743 137 8773 143
rect 8792 138 8797 143
rect 8709 121 8789 137
rect 8801 129 8837 150
rect 8922 149 8952 158
rect 8975 153 8993 171
rect 9051 169 9097 175
rect 9132 171 9145 181
rect 9163 171 9180 184
rect 9013 163 9015 165
rect 9015 160 9018 163
rect 9018 158 9027 160
rect 9000 151 9030 158
rect 9000 149 9031 151
rect 9051 149 9087 169
rect 9132 168 9180 171
rect 9145 163 9179 168
rect 8898 145 9087 149
rect 8913 142 9087 145
rect 8906 139 9087 142
rect 9115 162 9179 163
rect 8709 119 8728 121
rect 8743 119 8777 121
rect 8709 103 8789 119
rect 8709 97 8728 103
rect 8379 71 8405 80
rect 8425 71 8528 81
rect 8379 69 8528 71
rect 8549 69 8584 81
rect 8218 67 8380 69
rect 8230 47 8249 67
rect 8264 65 8294 67
rect 8076 38 8111 39
rect 8119 38 8154 39
rect 8076 29 8105 38
rect 8119 29 8148 38
rect 8236 29 8249 47
rect 8301 51 8380 67
rect 8412 67 8584 69
rect 8412 51 8491 67
rect 8498 65 8528 67
rect 8301 43 8491 51
rect 8556 47 8562 67
rect 8301 39 8380 43
rect 8382 39 8410 43
rect 8412 39 8491 43
rect 8286 29 8294 39
rect 8313 31 8316 39
rect 8317 31 8335 39
rect 8380 31 8412 39
rect 8457 31 8475 39
rect 8313 29 8479 31
rect 8498 29 8509 39
rect 8571 29 8584 67
rect 8656 81 8685 97
rect 8699 81 8728 97
rect 8743 87 8773 103
rect 8801 81 8807 129
rect 8810 123 8829 129
rect 8844 123 8874 131
rect 8810 115 8874 123
rect 8810 99 8890 115
rect 8906 108 8968 139
rect 8984 108 9046 139
rect 9115 137 9164 162
rect 9179 137 9209 153
rect 9078 123 9108 131
rect 9115 129 9225 137
rect 9078 115 9123 123
rect 8917 104 8952 108
rect 8810 97 8829 99
rect 8844 97 8890 99
rect 8810 81 8890 97
rect 8922 92 8952 104
rect 8993 105 9030 108
rect 8993 103 9035 105
rect 8931 88 8938 92
rect 8938 87 8939 88
rect 8897 81 8907 87
rect 8656 69 8691 81
rect 8693 69 8734 81
rect 8656 39 8734 69
rect 8798 69 8829 81
rect 8844 69 8947 81
rect 8959 80 8976 97
rect 9000 92 9030 103
rect 9062 99 9124 115
rect 9062 97 9108 99
rect 9062 81 9124 97
rect 9136 81 9142 129
rect 9145 121 9225 129
rect 9145 119 9164 121
rect 9179 119 9213 121
rect 9145 103 9225 119
rect 9145 81 9164 103
rect 9179 87 9209 103
rect 9237 97 9243 171
rect 9252 97 9265 241
rect 8959 71 8985 80
rect 9005 71 9108 81
rect 8959 69 9108 71
rect 9129 69 9164 81
rect 8798 67 8960 69
rect 8810 47 8829 67
rect 8844 65 8874 67
rect 8656 38 8691 39
rect 8699 38 8734 39
rect 8656 29 8685 38
rect 8699 29 8728 38
rect 8816 29 8829 47
rect 8881 51 8960 67
rect 8992 67 9164 69
rect 8992 51 9071 67
rect 9078 65 9108 67
rect 8881 43 9071 51
rect 9136 47 9142 67
rect 8881 39 8960 43
rect 8962 39 8990 43
rect 8992 39 9071 43
rect 8866 29 8874 39
rect 8893 31 8896 39
rect 8897 31 8915 39
rect 8960 31 8992 39
rect 9037 31 9055 39
rect 8893 29 9059 31
rect 9078 29 9089 39
rect 9151 29 9164 67
rect 9236 81 9265 97
rect 9236 38 9271 81
rect 9236 29 9265 38
rect -1 23 9265 29
rect 0 15 9265 23
rect 15 1 28 15
rect 43 -3 73 15
rect 116 1 159 15
rect 166 2 174 15
rect 207 2 345 15
rect 378 2 386 15
rect 129 -17 159 1
rect 222 -1 330 2
rect 222 -3 252 -1
rect 300 -3 330 -1
rect 393 -17 423 15
rect 451 1 464 15
rect 479 -3 509 15
rect 546 1 565 15
rect 580 1 586 15
rect 595 1 608 15
rect 623 -3 653 15
rect 696 1 739 15
rect 746 2 754 15
rect 787 2 925 15
rect 958 2 966 15
rect 709 -17 739 1
rect 802 -1 910 2
rect 802 -3 832 -1
rect 880 -3 910 -1
rect 973 -17 1003 15
rect 1031 1 1044 15
rect 1059 -3 1089 15
rect 1126 1 1145 15
rect 1160 1 1166 15
rect 1175 1 1188 15
rect 1203 -3 1233 15
rect 1276 1 1319 15
rect 1326 2 1334 15
rect 1367 2 1505 15
rect 1538 2 1546 15
rect 1289 -17 1319 1
rect 1382 -1 1490 2
rect 1382 -3 1412 -1
rect 1460 -3 1490 -1
rect 1553 -17 1583 15
rect 1611 1 1624 15
rect 1639 -3 1669 15
rect 1706 1 1725 15
rect 1740 1 1746 15
rect 1755 1 1768 15
rect 1783 -3 1813 15
rect 1856 1 1899 15
rect 1906 2 1914 15
rect 1947 2 2085 15
rect 2118 2 2126 15
rect 1869 -17 1899 1
rect 1962 -1 2070 2
rect 1962 -3 1992 -1
rect 2040 -3 2070 -1
rect 2133 -17 2163 15
rect 2191 1 2204 15
rect 2219 -3 2249 15
rect 2286 1 2305 15
rect 2320 1 2326 15
rect 2335 1 2348 15
rect 2363 -3 2393 15
rect 2436 1 2479 15
rect 2486 2 2494 15
rect 2527 2 2665 15
rect 2698 2 2706 15
rect 2449 -17 2479 1
rect 2542 -1 2650 2
rect 2542 -3 2572 -1
rect 2620 -3 2650 -1
rect 2713 -17 2743 15
rect 2771 1 2784 15
rect 2799 -3 2829 15
rect 2866 1 2885 15
rect 2900 1 2906 15
rect 2915 1 2928 15
rect 2943 -3 2973 15
rect 3016 1 3059 15
rect 3066 2 3074 15
rect 3107 2 3245 15
rect 3278 2 3286 15
rect 3029 -17 3059 1
rect 3122 -1 3230 2
rect 3122 -3 3152 -1
rect 3200 -3 3230 -1
rect 3293 -17 3323 15
rect 3351 1 3364 15
rect 3379 -3 3409 15
rect 3446 1 3465 15
rect 3480 1 3486 15
rect 3495 1 3508 15
rect 3523 -3 3553 15
rect 3596 1 3639 15
rect 3646 2 3654 15
rect 3687 2 3825 15
rect 3858 2 3866 15
rect 3609 -17 3639 1
rect 3702 -1 3810 2
rect 3702 -3 3732 -1
rect 3780 -3 3810 -1
rect 3873 -17 3903 15
rect 3931 1 3944 15
rect 3959 -3 3989 15
rect 4026 1 4045 15
rect 4060 1 4066 15
rect 4075 1 4088 15
rect 4103 -3 4133 15
rect 4176 1 4219 15
rect 4226 2 4234 15
rect 4267 2 4405 15
rect 4438 2 4446 15
rect 4189 -17 4219 1
rect 4282 -1 4390 2
rect 4282 -3 4312 -1
rect 4360 -3 4390 -1
rect 4453 -17 4483 15
rect 4511 1 4524 15
rect 4539 -3 4569 15
rect 4606 1 4625 15
rect 4640 1 4646 15
rect 4655 1 4668 15
rect 4683 -3 4713 15
rect 4756 1 4799 15
rect 4806 2 4814 15
rect 4847 2 4985 15
rect 5018 2 5026 15
rect 4769 -17 4799 1
rect 4862 -1 4970 2
rect 4862 -3 4892 -1
rect 4940 -3 4970 -1
rect 5033 -17 5063 15
rect 5091 1 5104 15
rect 5119 -3 5149 15
rect 5186 1 5205 15
rect 5220 1 5226 15
rect 5235 1 5248 15
rect 5263 -3 5293 15
rect 5336 1 5379 15
rect 5386 2 5394 15
rect 5427 2 5565 15
rect 5598 2 5606 15
rect 5349 -17 5379 1
rect 5442 -1 5550 2
rect 5442 -3 5472 -1
rect 5520 -3 5550 -1
rect 5613 -17 5643 15
rect 5671 1 5684 15
rect 5699 -3 5729 15
rect 5766 1 5785 15
rect 5800 1 5806 15
rect 5815 1 5828 15
rect 5843 -3 5873 15
rect 5916 1 5959 15
rect 5966 2 5974 15
rect 6007 2 6145 15
rect 6178 2 6186 15
rect 5929 -17 5959 1
rect 6022 -1 6130 2
rect 6022 -3 6052 -1
rect 6100 -3 6130 -1
rect 6193 -17 6223 15
rect 6251 1 6264 15
rect 6279 -3 6309 15
rect 6346 1 6365 15
rect 6380 1 6386 15
rect 6395 1 6408 15
rect 6423 -3 6453 15
rect 6496 1 6539 15
rect 6546 2 6554 15
rect 6587 2 6725 15
rect 6758 2 6766 15
rect 6509 -17 6539 1
rect 6602 -1 6710 2
rect 6602 -3 6632 -1
rect 6680 -3 6710 -1
rect 6773 -17 6803 15
rect 6831 1 6844 15
rect 6859 -3 6889 15
rect 6926 1 6945 15
rect 6960 1 6966 15
rect 6975 1 6988 15
rect 7003 -3 7033 15
rect 7076 1 7119 15
rect 7126 2 7134 15
rect 7167 2 7305 15
rect 7338 2 7346 15
rect 7089 -17 7119 1
rect 7182 -1 7290 2
rect 7182 -3 7212 -1
rect 7260 -3 7290 -1
rect 7353 -17 7383 15
rect 7411 1 7424 15
rect 7439 -3 7469 15
rect 7506 1 7525 15
rect 7540 1 7546 15
rect 7555 1 7568 15
rect 7583 -3 7613 15
rect 7656 1 7699 15
rect 7706 2 7714 15
rect 7747 2 7885 15
rect 7918 2 7926 15
rect 7669 -17 7699 1
rect 7762 -1 7870 2
rect 7762 -3 7792 -1
rect 7840 -3 7870 -1
rect 7933 -17 7963 15
rect 7991 1 8004 15
rect 8019 -3 8049 15
rect 8086 1 8105 15
rect 8120 1 8126 15
rect 8135 1 8148 15
rect 8163 -3 8193 15
rect 8236 1 8279 15
rect 8286 2 8294 15
rect 8327 2 8465 15
rect 8498 2 8506 15
rect 8249 -17 8279 1
rect 8342 -1 8450 2
rect 8342 -3 8372 -1
rect 8420 -3 8450 -1
rect 8513 -17 8543 15
rect 8571 1 8584 15
rect 8599 -3 8629 15
rect 8666 1 8685 15
rect 8700 1 8706 15
rect 8715 1 8728 15
rect 8743 -3 8773 15
rect 8816 1 8859 15
rect 8866 2 8874 15
rect 8907 2 9045 15
rect 9078 2 9086 15
rect 8829 -17 8859 1
rect 8922 -1 9030 2
rect 8922 -3 8952 -1
rect 9000 -3 9030 -1
rect 9093 -17 9123 15
rect 9151 1 9164 15
rect 9179 -3 9209 15
rect 9252 1 9265 15
<< pwell >>
rect 4612 7560 4640 7574
rect 4612 7516 4640 7530
rect 4612 7290 4640 7304
rect 4612 7246 4640 7260
rect 4612 7020 4640 7034
rect 4612 6976 4640 6990
rect 4612 6750 4640 6764
rect 4612 6706 4640 6720
rect 4612 6480 4640 6494
rect 4612 6436 4640 6450
rect 4612 6210 4640 6224
rect 4612 6166 4640 6180
rect 4612 5940 4640 5954
rect 4612 5896 4640 5910
rect 4612 5670 4640 5684
rect 4612 5626 4640 5640
rect 4612 5400 4640 5414
rect 4612 5356 4640 5370
rect 4612 5130 4640 5144
rect 4612 5086 4640 5100
rect 4612 4860 4640 4874
rect 4612 4816 4640 4830
rect 4612 4590 4640 4604
rect 4612 4546 4640 4560
rect 4612 4320 4640 4334
rect 4612 4276 4640 4290
rect 4612 4050 4640 4064
rect 4612 4006 4640 4020
rect 4612 3780 4640 3794
rect 4612 3736 4640 3750
rect 4612 3510 4640 3524
rect 4612 3466 4640 3480
rect 4612 3240 4640 3254
rect 4612 3196 4640 3210
rect 4612 2970 4640 2984
rect 4612 2926 4640 2940
rect 4612 2700 4640 2714
rect 4612 2656 4640 2670
rect 4612 2430 4640 2444
rect 4612 2386 4640 2400
rect 4612 2160 4640 2174
rect 4612 2116 4640 2130
rect 4612 1890 4640 1904
rect 4612 1846 4640 1860
rect 4612 1620 4640 1634
rect 4612 1576 4640 1590
rect 4612 1350 4640 1364
rect 4612 1306 4640 1320
rect 4612 1080 4640 1094
rect 4612 1036 4640 1050
rect 4612 810 4640 824
rect 4612 766 4640 780
rect 4612 540 4640 554
rect 4612 496 4640 510
rect 4612 270 4640 284
rect 4612 226 4640 240
rect 74 184 89 212
rect 464 184 479 213
rect 4714 184 4729 212
rect 5104 184 5119 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 4640 38 4655 80
rect 5177 38 5192 80
rect 5220 38 5235 80
rect 4612 0 4640 14
<< ndiffc >>
rect 74 185 89 213
rect 464 185 479 214
rect 654 185 669 213
rect 1044 185 1059 214
rect 1234 185 1249 213
rect 1624 185 1639 214
rect 1814 185 1829 213
rect 2204 185 2219 214
rect 2394 185 2409 213
rect 2784 185 2799 214
rect 2974 185 2989 213
rect 3364 185 3379 214
rect 3554 185 3569 213
rect 3944 185 3959 214
rect 4134 185 4149 213
rect 4524 185 4539 214
rect 4714 185 4729 213
rect 5104 184 5119 213
rect 5294 184 5309 212
rect 5684 184 5699 213
rect 5874 184 5889 212
rect 6264 184 6279 213
rect 6454 184 6469 212
rect 6844 184 6859 213
rect 7034 184 7049 212
rect 7424 184 7439 213
rect 7614 184 7629 212
rect 8004 184 8019 213
rect 8194 184 8209 212
rect 8584 184 8599 213
rect 8774 184 8789 212
rect 9164 184 9179 213
rect 0 39 15 81
rect 537 39 552 81
rect 580 39 595 81
rect 1117 39 1132 81
rect 1160 39 1175 81
rect 1697 39 1712 81
rect 1740 39 1755 81
rect 2277 39 2292 81
rect 2320 39 2335 81
rect 2857 39 2872 81
rect 2900 39 2915 81
rect 3437 39 3452 81
rect 3480 39 3495 81
rect 4017 39 4032 81
rect 4060 39 4075 81
rect 4597 39 4612 81
rect 4640 39 4655 81
rect 5177 38 5192 80
rect 5220 38 5235 80
rect 5757 38 5772 80
rect 5800 38 5815 80
rect 6337 38 6352 80
rect 6380 38 6395 80
rect 6917 38 6932 80
rect 6960 38 6975 80
rect 7497 38 7512 80
rect 7540 38 7555 80
rect 8077 38 8092 80
rect 8120 38 8135 80
rect 8657 38 8672 80
rect 8700 38 8715 80
rect 9237 38 9252 80
<< poly >>
rect 0 8610 30 8640
rect 4561 8610 4708 8640
rect 0 8340 30 8370
rect 4567 8340 4701 8370
rect 0 8070 30 8100
rect 4571 8070 4694 8100
rect 0 7800 30 7830
rect 4574 7800 4724 7830
rect 0 7530 30 7560
rect 4558 7530 4711 7560
rect 0 7260 30 7290
rect 4556 7260 4739 7290
rect 0 6990 30 7020
rect 4554 6990 4707 7020
rect 0 6720 30 6750
rect 4563 6720 4759 6750
rect 0 6450 30 6480
rect 4572 6450 4700 6480
rect 0 6180 30 6210
rect 4575 6180 4747 6210
rect 0 5910 30 5940
rect 4563 5910 4729 5940
rect 0 5640 30 5670
rect 4560 5640 4732 5670
rect 0 5370 30 5400
rect 4563 5370 4700 5400
rect 0 5100 30 5130
rect 4572 5100 4706 5130
rect 0 4830 30 4860
rect 4544 4830 4694 4860
rect 0 4560 30 4590
rect 4561 4560 4714 4590
rect 0 4290 30 4320
rect 4568 4290 4703 4320
rect 0 4020 30 4050
rect 4566 4020 4736 4050
rect 0 3750 30 3780
rect 4563 3750 4719 3780
rect 0 3480 30 3510
rect 4561 3480 4713 3510
rect 0 3210 30 3240
rect 4563 3210 4714 3240
rect 0 2940 30 2970
rect 4565 2940 4704 2970
rect 0 2670 30 2700
rect 4553 2670 4697 2700
rect 0 2400 30 2430
rect 4553 2400 4701 2430
rect 0 2130 30 2160
rect 4562 2130 4697 2160
rect 0 1860 30 1890
rect 4564 1860 4695 1890
rect 0 1590 30 1620
rect 4566 1590 4721 1620
rect 0 1320 30 1350
rect 4569 1320 4706 1350
rect 0 1050 30 1080
rect 4549 1050 4695 1080
rect 0 780 30 810
rect 4564 780 4713 810
rect 0 510 30 540
rect 4577 510 4701 540
rect 0 241 30 271
rect 4570 241 4698 271
<< metal1 >>
rect 0 8596 15 8610
rect 4576 8596 4671 8610
rect 0 8472 15 8506
rect 4505 8472 4691 8506
rect 0 8370 15 8384
rect 4573 8370 4670 8384
rect 0 8326 15 8340
rect 4578 8326 4678 8340
rect 0 8202 15 8236
rect 4502 8202 4701 8236
rect 0 8100 15 8114
rect 4578 8100 4688 8114
rect 0 8056 15 8070
rect 4581 8056 4663 8070
rect 0 7932 15 7966
rect 4505 7932 4727 7966
rect 0 7830 15 7844
rect 4582 7830 4666 7844
rect 0 7786 15 7800
rect 4575 7786 4685 7800
rect 0 7662 15 7696
rect 4640 7662 4655 7696
rect 0 7560 15 7574
rect 4612 7560 4655 7574
rect 0 7516 15 7530
rect 4612 7516 4655 7530
rect 0 7392 15 7426
rect 4504 7392 4727 7426
rect 0 7290 15 7304
rect 4612 7290 4655 7304
rect 0 7246 15 7260
rect 4612 7246 4655 7260
rect 0 7122 15 7156
rect 4496 7122 4683 7156
rect 0 7020 15 7034
rect 4612 7020 4655 7034
rect 0 6976 15 6990
rect 4612 6976 4655 6990
rect 0 6852 15 6886
rect 4505 6852 4734 6886
rect 0 6750 15 6764
rect 4612 6750 4655 6764
rect 0 6706 15 6720
rect 4612 6706 4655 6720
rect 0 6582 15 6616
rect 4502 6582 4705 6616
rect 0 6480 15 6494
rect 4612 6480 4655 6494
rect 0 6436 15 6450
rect 4612 6436 4655 6450
rect 0 6312 15 6346
rect 4505 6312 4722 6346
rect 0 6210 15 6224
rect 4612 6210 4655 6224
rect 0 6166 15 6180
rect 4612 6166 4655 6180
rect 0 6042 15 6076
rect 4499 6042 4731 6076
rect 0 5940 15 5954
rect 4612 5940 4655 5954
rect 0 5896 15 5910
rect 4612 5896 4655 5910
rect 0 5772 15 5806
rect 4505 5772 4740 5806
rect 0 5670 15 5684
rect 4612 5670 4655 5684
rect 0 5626 15 5640
rect 4612 5626 4655 5640
rect 0 5502 15 5536
rect 4505 5502 4728 5536
rect 0 5400 15 5414
rect 4612 5400 4655 5414
rect 0 5356 15 5370
rect 4612 5356 4655 5370
rect 0 5232 15 5266
rect 4496 5232 4728 5266
rect 0 5130 15 5144
rect 4612 5130 4655 5144
rect 0 5086 15 5100
rect 4612 5086 4655 5100
rect 0 4962 15 4996
rect 4502 4962 4746 4996
rect 0 4860 15 4874
rect 4612 4860 4655 4874
rect 0 4816 15 4830
rect 4612 4816 4655 4830
rect 0 4692 15 4726
rect 4505 4692 4716 4726
rect 0 4590 15 4604
rect 4612 4590 4655 4604
rect 0 4546 15 4560
rect 4612 4546 4655 4560
rect 0 4422 15 4456
rect 4503 4422 4753 4456
rect 0 4320 15 4334
rect 4612 4320 4655 4334
rect 0 4276 15 4290
rect 4612 4276 4655 4290
rect 0 4152 15 4186
rect 4505 4152 4724 4186
rect 0 4050 15 4064
rect 4612 4050 4655 4064
rect 0 4006 15 4020
rect 4612 4006 4655 4020
rect 0 3882 15 3916
rect 4503 3882 4731 3916
rect 0 3780 15 3794
rect 4612 3780 4655 3794
rect 0 3736 15 3750
rect 4612 3736 4655 3750
rect 0 3612 15 3646
rect 4505 3612 4736 3646
rect 0 3510 15 3524
rect 4612 3510 4655 3524
rect 0 3466 15 3480
rect 4612 3466 4655 3480
rect 0 3342 15 3376
rect 4496 3342 4727 3376
rect 0 3240 15 3254
rect 4612 3240 4655 3254
rect 0 3196 15 3210
rect 4612 3196 4655 3210
rect 0 3072 15 3106
rect 4502 3072 4741 3106
rect 0 2970 15 2984
rect 4612 2970 4655 2984
rect 0 2926 15 2940
rect 4612 2926 4655 2940
rect 0 2802 15 2836
rect 4502 2802 4734 2836
rect 0 2700 15 2714
rect 4612 2700 4655 2714
rect 0 2656 15 2670
rect 4612 2656 4655 2670
rect 0 2532 15 2566
rect 4505 2532 4736 2566
rect 0 2430 15 2444
rect 4612 2430 4655 2444
rect 0 2386 15 2400
rect 4612 2386 4655 2400
rect 0 2262 15 2296
rect 4497 2262 4740 2296
rect 0 2160 15 2174
rect 4612 2160 4655 2174
rect 0 2116 15 2130
rect 4612 2116 4655 2130
rect 0 1992 15 2026
rect 4505 1992 4710 2026
rect 0 1890 15 1904
rect 4612 1890 4655 1904
rect 0 1846 15 1860
rect 4612 1846 4655 1860
rect 0 1722 15 1756
rect 4505 1722 4688 1756
rect 0 1620 15 1634
rect 4612 1620 4655 1634
rect 0 1576 15 1590
rect 4612 1576 4655 1590
rect 0 1452 15 1486
rect 4501 1452 4708 1486
rect 0 1350 15 1364
rect 4612 1350 4655 1364
rect 0 1306 15 1320
rect 4612 1306 4655 1320
rect 0 1182 15 1216
rect 4505 1182 4701 1216
rect 0 1080 15 1094
rect 4612 1080 4655 1094
rect 0 1036 15 1050
rect 4612 1036 4655 1050
rect 0 912 15 946
rect 4505 912 4725 946
rect 0 810 15 824
rect 4612 810 4655 824
rect 0 766 15 780
rect 4612 766 4655 780
rect 0 642 15 676
rect 4505 642 4741 676
rect 0 540 15 554
rect 4612 540 4655 554
rect 0 496 15 510
rect 4612 496 4655 510
rect 0 372 15 406
rect 4505 372 4683 406
rect 0 271 15 284
rect 4612 271 4655 284
rect 0 227 15 241
rect 4612 227 4655 241
rect 0 103 15 137
rect 4505 103 4705 137
rect 0 1 15 15
rect 4612 1 4655 15
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1656019537
transform 1 0 0 0 1 7830
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1656019537
transform 1 0 0 0 1 7560
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1656019537
transform 1 0 0 0 1 8370
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1656019537
transform 1 0 0 0 1 8100
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1656019537
transform 1 0 0 0 1 6480
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1656019537
transform 1 0 0 0 1 6750
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1656019537
transform 1 0 0 0 1 7290
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1656019537
transform 1 0 0 0 1 7020
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_8
timestamp 1656019537
transform 1 0 0 0 1 4590
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_9
timestamp 1656019537
transform 1 0 0 0 1 4320
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_10
timestamp 1656019537
transform 1 0 0 0 1 4860
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_11
timestamp 1656019537
transform 1 0 0 0 1 5130
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_12
timestamp 1656019537
transform 1 0 0 0 1 5400
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_13
timestamp 1656019537
transform 1 0 0 0 1 5670
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_14
timestamp 1656019537
transform 1 0 0 0 1 6210
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_15
timestamp 1656019537
transform 1 0 0 0 1 5940
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_16
timestamp 1656019537
transform 1 0 0 0 1 1
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_17
timestamp 1656019537
transform 1 0 0 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_18
timestamp 1656019537
transform 1 0 0 0 1 271
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_19
timestamp 1656019537
transform 1 0 0 0 1 1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_20
timestamp 1656019537
transform 1 0 0 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_21
timestamp 1656019537
transform 1 0 0 0 1 1620
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_22
timestamp 1656019537
transform 1 0 0 0 1 1350
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_23
timestamp 1656019537
transform 1 0 0 0 1 2160
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_24
timestamp 1656019537
transform 1 0 0 0 1 1890
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_25
timestamp 1656019537
transform 1 0 0 0 1 2700
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_26
timestamp 1656019537
transform 1 0 0 0 1 2430
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_27
timestamp 1656019537
transform 1 0 0 0 1 3240
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_28
timestamp 1656019537
transform 1 0 0 0 1 2970
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_29
timestamp 1656019537
transform 1 0 0 0 1 3780
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_30
timestamp 1656019537
transform 1 0 0 0 1 3510
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_31
timestamp 1656019537
transform 1 0 0 0 1 4050
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_32
timestamp 1656019537
transform 1 0 4640 0 1 271
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_33
timestamp 1656019537
transform 1 0 4640 0 1 1
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_34
timestamp 1656019537
transform 1 0 4640 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_35
timestamp 1656019537
transform 1 0 4640 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_36
timestamp 1656019537
transform 1 0 4640 0 1 1350
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_37
timestamp 1656019537
transform 1 0 4640 0 1 1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_38
timestamp 1656019537
transform 1 0 4640 0 1 1890
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_39
timestamp 1656019537
transform 1 0 4640 0 1 2160
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_40
timestamp 1656019537
transform 1 0 4640 0 1 1620
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_41
timestamp 1656019537
transform 1 0 4640 0 1 2430
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_42
timestamp 1656019537
transform 1 0 4640 0 1 2700
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_43
timestamp 1656019537
transform 1 0 4640 0 1 2970
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_44
timestamp 1656019537
transform 1 0 4640 0 1 3240
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_45
timestamp 1656019537
transform 1 0 4640 0 1 3780
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_46
timestamp 1656019537
transform 1 0 4640 0 1 3510
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_47
timestamp 1656019537
transform 1 0 4640 0 1 4050
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_48
timestamp 1656019537
transform 1 0 4640 0 1 4320
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_49
timestamp 1656019537
transform 1 0 4640 0 1 4590
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_50
timestamp 1656019537
transform 1 0 4640 0 1 4860
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_51
timestamp 1656019537
transform 1 0 4640 0 1 5130
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_52
timestamp 1656019537
transform 1 0 4640 0 1 5400
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_53
timestamp 1656019537
transform 1 0 4640 0 1 5670
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_54
timestamp 1656019537
transform 1 0 4640 0 1 5940
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_55
timestamp 1656019537
transform 1 0 4640 0 1 6210
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_56
timestamp 1656019537
transform 1 0 4640 0 1 6480
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_57
timestamp 1656019537
transform 1 0 4640 0 1 6750
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_58
timestamp 1656019537
transform 1 0 4640 0 1 7020
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_59
timestamp 1656019537
transform 1 0 4640 0 1 7290
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_60
timestamp 1656019537
transform 1 0 4640 0 1 7560
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_61
timestamp 1656019537
transform 1 0 4640 0 1 7830
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_62
timestamp 1656019537
transform 1 0 4640 0 1 8100
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_63
timestamp 1656019537
transform 1 0 4640 0 1 8370
box -7 -4 4631 312
<< labels >>
rlabel locali 0 39 15 81 1 RBL1_0
port 1 ns signal output
rlabel locali 537 39 552 81 1 RBL0_0
port 2 ns signal output
rlabel locali 580 39 595 81 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 39 1132 81 1 RBL0_1
port 4 ns signal output
rlabel locali 1160 39 1175 81 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 39 1712 81 1 RBL0_2
port 6 ns signal output
rlabel locali 1740 39 1755 81 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 39 2292 81 1 RBL0_3
port 8 ns signal output
rlabel locali 2320 39 2335 81 1 RBL1_4
port 9 ns signal output
rlabel locali 2857 39 2872 81 1 RBL0_4
port 10 ns signal output
rlabel locali 2900 39 2915 81 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 39 3452 81 1 RBL0_5
port 12 ns signal output
rlabel locali 3480 39 3495 81 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 39 4032 81 1 RBL0_6
port 14 ns signal output
rlabel locali 4060 39 4075 81 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 39 4612 81 1 RBL0_7
port 16 ns signal output
rlabel locali 4640 39 4655 81 1 RBL1_8
port 17 ns signal output
rlabel locali 5177 38 5192 80 1 RBL0_8
port 18 ns signal output
rlabel locali 5220 38 5235 80 1 RBL1_9
port 19 ns signal output
rlabel locali 5757 38 5772 80 1 RBL0_9
port 20 ns signal output
rlabel locali 5800 38 5815 80 1 RBL1_10
port 21 ns signal output
rlabel locali 6337 38 6352 80 1 RBL0_10
port 22 ns signal output
rlabel locali 6380 38 6395 80 1 RBL1_11
port 23 ns signal output
rlabel locali 6917 38 6932 80 1 RBL0_11
port 24 ns signal output
rlabel locali 6960 38 6975 80 1 RBL1_12
port 25 ns signal output
rlabel locali 7497 38 7512 80 1 RBL0_12
port 26 ns signal output
rlabel locali 7540 38 7555 80 1 RBL1_13
port 27 ns signal output
rlabel locali 8077 38 8092 80 1 RBL0_13
port 28 ns signal output
rlabel locali 8120 38 8135 80 1 RBL1_14
port 29 ns signal output
rlabel locali 8657 38 8672 80 1 RBL0_14
port 30 ns signal output
rlabel locali 8700 38 8715 80 1 RBL1_15
port 31 ns signal output
rlabel locali 9237 38 9252 80 1 RBL0_15
port 32 ns signal output
rlabel poly 0 8610 30 8640 1 WWL_0
port 33 ew signal input
rlabel metal1 0 8472 15 8506 1 RWL_0
port 34 ew signal input
rlabel poly 0 8340 30 8370 1 WWL_1
port 35 ew signal input
rlabel metal1 0 8202 15 8236 1 RWL_1
port 36 ew signal input
rlabel poly 0 8070 30 8100 1 WWL_2
port 37 ew signal input
rlabel metal1 0 7932 15 7966 1 RWL_2
port 38 ew signal input
rlabel poly 0 7800 30 7830 1 WWL_3
port 39 ew signal input
rlabel metal1 0 7662 15 7696 1 RWL_3
port 40 ew signal input
rlabel poly 0 7530 30 7560 1 WWL_4
port 41 ew signal input
rlabel metal1 0 7392 15 7426 1 RWL_4
port 42 ew signal input
rlabel poly 0 7260 30 7290 1 WWL_5
port 43 ew signal input
rlabel metal1 0 7122 15 7156 1 RWL_5
port 44 ew signal input
rlabel poly 0 6990 30 7020 1 WWL_6
port 45 ew signal input
rlabel metal1 0 6852 15 6886 1 RWL_6
port 46 ew signal input
rlabel poly 0 6720 30 6750 1 WWL_7
port 47 ew signal input
rlabel metal1 0 6582 15 6616 1 RWL_7
port 48 ew signal input
rlabel poly 0 6450 30 6480 1 WWL_8
port 49 ew signal input
rlabel metal1 0 6312 15 6346 1 RWL_8
port 50 ew signal input
rlabel poly 0 6180 30 6210 1 WWL_9
port 51 ew signal input
rlabel metal1 0 6042 15 6076 1 RWL_9
port 52 ew signal input
rlabel poly 0 5910 30 5940 1 WWL_10
port 53 ew signal input
rlabel metal1 0 5772 15 5806 1 RWL_10
port 54 ew signal input
rlabel poly 0 5640 30 5670 1 WWL_11
port 55 ew signal input
rlabel metal1 0 5502 15 5536 1 RWL_11
port 56 ew signal input
rlabel poly 0 5370 30 5400 1 WWL_12
port 57 ew signal input
rlabel metal1 0 5232 15 5266 1 RWL_12
port 58 ew signal input
rlabel poly 0 5100 30 5130 1 WWL_13
port 59 ew signal input
rlabel metal1 0 4962 15 4996 1 RWL_13
port 60 ew signal input
rlabel poly 0 4830 30 4860 1 WWL_14
port 61 ew signal input
rlabel metal1 0 4692 15 4726 1 RWL_14
port 62 ew signal input
rlabel poly 0 4560 30 4590 1 WWL_15
port 63 ew signal input
rlabel metal1 0 4422 15 4456 1 RWL_15
port 64 ew signal input
rlabel poly 0 4290 30 4320 1 WWL_16
port 65 ew signal input
rlabel metal1 0 4152 15 4186 1 RWL_16
port 66 ew signal input
rlabel poly 0 4020 30 4050 1 WWL_17
port 67 ew signal input
rlabel metal1 0 3882 15 3916 1 RWL_17
port 68 ew signal input
rlabel poly 0 3750 30 3780 1 WWL_18
port 69 ew signal input
rlabel metal1 0 3612 15 3646 1 RWL_18
port 70 ew signal input
rlabel poly 0 3480 30 3510 1 WWL_19
port 71 ew signal input
rlabel metal1 0 3342 15 3376 1 RWL_19
port 72 ew signal input
rlabel poly 0 3210 30 3240 1 WWL_20
port 73 ew signal input
rlabel metal1 0 3072 15 3106 1 RWL_20
port 74 ew signal input
rlabel poly 0 2940 30 2970 1 WWL_21
port 75 ew signal input
rlabel metal1 0 2802 15 2836 1 RWL_21
port 76 ew signal input
rlabel poly 0 2670 30 2700 1 WWL_22
port 77 ew signal input
rlabel metal1 0 2532 15 2566 1 RWL_22
port 78 ew signal input
rlabel poly 0 2400 30 2430 1 WWL_23
port 79 ew signal input
rlabel metal1 0 2262 15 2296 1 RWL_23
port 80 ew signal input
rlabel poly 0 2130 30 2160 1 WWL_24
port 81 ew signal input
rlabel metal1 0 1992 15 2026 1 RWL_24
port 82 ew signal input
rlabel poly 0 1860 30 1890 1 WWL_25
port 83 ew signal input
rlabel metal1 0 1722 15 1756 1 RWL_25
port 84 ew signal input
rlabel poly 0 1590 30 1620 1 WWL_26
port 85 ew signal input
rlabel metal1 0 1452 15 1486 1 RWL_26
port 86 ew signal input
rlabel poly 0 1320 30 1350 1 WWL_27
port 87 ew signal input
rlabel metal1 0 1182 15 1216 1 RWL_27
port 88 ew signal input
rlabel poly 0 1050 30 1080 1 WWL_28
port 89 ew signal input
rlabel metal1 0 912 15 946 1 RWL_28
port 90 ew signal input
rlabel poly 0 780 30 810 1 WWL_29
port 91 ew signal input
rlabel metal1 0 642 15 676 1 RWL_29
port 92 ew signal input
rlabel poly 0 510 30 540 1 WWL_30
port 93 ew signal input
rlabel metal1 0 372 15 406 1 RWL_30
port 94 ew signal input
rlabel poly 0 241 30 271 1 WWL_31
port 95 ew signal input
rlabel metal1 0 103 15 137 1 RWL_31
port 96 ew signal input
rlabel locali 464 185 479 214 1 WBL_0
port 97 ns signal input
rlabel locali 74 185 89 213 1 WBLb_0
port 98 ns signal input
rlabel locali 1044 185 1059 214 1 WBL_1
port 99 ns signal input
rlabel locali 654 185 669 213 1 WBLb_1
port 100 ns signal input
rlabel locali 1624 185 1639 214 1 WBL_2
port 101 ns signal input
rlabel locali 1234 185 1249 213 1 WBLb_2
port 102 ns signal input
rlabel locali 2204 185 2219 214 1 WBL_3
port 103 ns signal input
rlabel locali 1814 185 1829 213 1 WBLb_3
port 104 ns signal input
rlabel locali 2784 185 2799 214 1 WBL_4
port 105 ns signal input
rlabel locali 2394 185 2409 213 1 WBLb_4
port 106 ns signal input
rlabel locali 3364 185 3379 214 1 WBL_5
port 107 ns signal input
rlabel locali 2974 185 2989 213 1 WBLb_5
port 108 ns signal input
rlabel locali 3944 185 3959 214 1 WBL_6
port 109 ns signal input
rlabel locali 3554 185 3569 213 1 WBLb_6
port 110 ns signal input
rlabel locali 4524 185 4539 214 1 WBL_7
port 111 ns signal input
rlabel locali 4134 185 4149 213 1 WBLb_7
port 112 ns signal input
rlabel locali 5104 184 5119 213 1 WBL_8
port 113 ns signal input
rlabel locali 4714 185 4729 213 1 WBLb_8
port 114 ns signal input
rlabel locali 5684 184 5699 213 1 WBL_9
port 115 ns signal input
rlabel locali 5294 184 5309 212 1 WBLb_9
port 116 ns signal input
rlabel locali 6264 184 6279 213 1 WBL_10
port 117 ns signal input
rlabel locali 5874 184 5889 212 1 WBLb_10
port 118 ns signal input
rlabel locali 6844 184 6859 213 1 WBL_11
port 119 ns signal input
rlabel locali 6454 184 6469 212 1 WBLb_11
port 120 ns signal input
rlabel locali 7424 184 7439 213 1 WBL_12
port 121 ns signal input
rlabel locali 7034 184 7049 212 1 WBLb_12
port 122 ns signal input
rlabel locali 8004 184 8019 213 1 WBL_13
port 123 ns signal input
rlabel locali 7614 184 7629 212 1 WBLb_13
port 124 ns signal input
rlabel locali 8584 184 8599 213 1 WBL_14
port 125 ns signal input
rlabel locali 8194 184 8209 212 1 WBLb_14
port 126 ns signal input
rlabel locali 9164 184 9179 213 1 WBL_15
port 127 ns signal input
rlabel locali 8774 184 8789 212 1 WBLb_15
port 128 ns signal input
rlabel metal1 0 227 15 241 1 VDD
port 129 ew power bidirectional abutment
rlabel metal1 0 1 15 15 1 GND
port 130 ew ground bidirectional abutment
rlabel metal1 0 8596 15 8610 1 VDD
rlabel metal1 0 8370 15 8384 1 GND
rlabel metal1 0 8326 15 8340 1 VDD
rlabel metal1 0 8100 15 8114 1 GND
rlabel metal1 0 8056 15 8070 1 VDD
rlabel metal1 0 7830 15 7844 1 GND
rlabel metal1 0 7786 15 7800 1 VDD
rlabel metal1 0 7560 15 7574 1 GND
rlabel metal1 0 7516 15 7530 1 VDD
rlabel metal1 0 7290 15 7304 1 GND
rlabel metal1 0 7246 15 7260 1 VDD
rlabel metal1 0 7020 15 7034 1 GND
rlabel metal1 0 6976 15 6990 1 VDD
rlabel metal1 0 6750 15 6764 1 GND
rlabel metal1 0 6706 15 6720 1 VDD
rlabel metal1 0 6480 15 6494 1 GND
rlabel metal1 0 6436 15 6450 1 VDD
rlabel metal1 0 6210 15 6224 1 GND
rlabel metal1 0 6166 15 6180 1 VDD
rlabel metal1 0 5940 15 5954 1 GND
rlabel metal1 0 5896 15 5910 1 VDD
rlabel metal1 0 5670 15 5684 1 GND
rlabel metal1 0 5626 15 5640 1 VDD
rlabel metal1 0 5400 15 5414 1 GND
rlabel metal1 0 5356 15 5370 1 VDD
rlabel metal1 0 5130 15 5144 1 GND
rlabel metal1 0 5086 15 5100 1 VDD
rlabel metal1 0 4860 15 4874 1 GND
rlabel metal1 0 4816 15 4830 1 VDD
rlabel metal1 0 4590 15 4604 1 GND
rlabel metal1 0 4546 15 4560 1 VDD
rlabel metal1 0 4320 15 4334 1 GND
rlabel metal1 0 4276 15 4290 1 VDD
rlabel metal1 0 4050 15 4064 1 GND
rlabel metal1 0 4006 15 4020 1 VDD
rlabel metal1 0 3780 15 3794 1 GND
rlabel metal1 0 3736 15 3750 1 VDD
rlabel metal1 0 3510 15 3524 1 GND
rlabel metal1 0 3466 15 3480 1 VDD
rlabel metal1 0 3240 15 3254 1 GND
rlabel metal1 0 3196 15 3210 1 VDD
rlabel metal1 0 2926 15 2940 1 VDD
rlabel metal1 0 2970 15 2984 1 GND
rlabel metal1 0 2700 15 2714 1 GND
rlabel metal1 0 2656 15 2670 1 VDD
rlabel metal1 0 2430 15 2444 1 GND
rlabel metal1 0 2386 15 2400 1 VDD
rlabel metal1 0 2160 15 2174 1 GND
rlabel metal1 0 2116 15 2130 1 VDD
rlabel metal1 0 1890 15 1904 1 GND
rlabel metal1 0 1846 15 1860 1 VDD
rlabel metal1 0 1620 15 1634 1 GND
rlabel metal1 0 1576 15 1590 1 VDD
rlabel metal1 0 1350 15 1364 1 GND
rlabel metal1 0 1306 15 1320 1 VDD
rlabel metal1 0 1080 15 1094 1 GND
rlabel metal1 0 1036 15 1050 1 VDD
rlabel metal1 0 810 15 824 1 GND
rlabel metal1 0 766 15 780 1 VDD
rlabel metal1 0 540 15 554 1 GND
rlabel metal1 0 496 15 510 1 VDD
rlabel metal1 0 270 15 284 1 GND
<< end >>
