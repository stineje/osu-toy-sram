magic
tech sky130
magscale 1 2
timestamp 1653352002
<< error_p >>
rect -778 991 -776 1004
rect -806 957 -798 991
rect -786 957 -772 991
rect -778 946 -776 957
rect -862 916 -806 946
rect -778 916 -722 946
rect -778 858 -776 916
rect -435 866 -339 931
rect -806 816 -790 832
rect -407 816 -405 826
rect -822 800 -811 816
rect -822 782 -811 798
rect -806 782 -798 816
rect -772 782 -764 816
rect -447 804 -427 816
rect -618 782 -516 799
rect -435 782 -427 804
rect -415 804 -395 816
rect -415 782 -401 804
rect -806 771 -790 782
rect -848 766 -790 771
rect -848 741 -806 766
rect -764 747 -722 771
rect -584 765 -568 781
rect -566 765 -550 781
rect -407 771 -405 782
rect -369 771 -316 863
rect -600 749 -534 765
rect -584 748 -550 749
rect -764 746 -597 747
rect -780 741 -597 746
rect -780 730 -764 741
rect -600 731 -593 741
rect -584 735 -583 748
rect -491 741 -435 771
rect -407 741 -316 771
rect -584 731 -550 735
rect -537 731 -534 741
rect -407 730 -405 741
rect -806 696 -798 730
rect -772 696 -764 730
rect -759 714 -748 730
rect -593 725 -537 727
rect -584 715 -568 725
rect -566 715 -550 725
rect -759 696 -748 712
rect -685 705 -669 713
rect -667 705 -651 713
rect -780 685 -764 696
rect -701 685 -697 697
rect -685 695 -651 697
rect -639 685 -635 697
rect -435 696 -427 730
rect -415 696 -401 730
rect -407 685 -405 696
rect -369 685 -316 741
rect -848 655 -806 685
rect -780 680 -722 685
rect -764 655 -722 680
rect -701 678 -685 679
rect -651 678 -635 679
rect -701 663 -635 678
rect -685 647 -669 663
rect -667 647 -651 663
rect -491 655 -435 685
rect -407 655 -316 685
rect -407 644 -405 655
rect -806 610 -798 644
rect -772 610 -764 644
rect -719 629 -617 644
rect -435 622 -427 644
rect -447 610 -427 622
rect -415 622 -401 644
rect -415 610 -395 622
rect -407 604 -405 610
rect -369 604 -316 655
rect -484 559 -316 604
rect -817 521 -797 533
rect -805 499 -797 521
rect -771 521 -751 533
rect -771 499 -763 521
rect -448 515 -428 527
rect -436 493 -428 515
rect -402 515 -382 527
rect -402 493 -394 515
rect -847 474 -805 482
rect -763 474 -721 482
rect -847 452 -721 474
rect -478 473 -436 482
rect -394 473 -352 482
rect -551 452 -348 473
rect -309 452 -306 524
rect -807 439 -805 452
rect -777 432 -763 447
rect -861 402 -805 432
rect -777 402 -721 432
rect -436 431 -422 446
rect -478 402 -422 431
rect -394 431 -392 452
rect -394 402 -338 431
rect -777 391 -775 402
rect -478 401 -338 402
rect -394 391 -392 401
rect -805 356 -797 391
rect -785 356 -771 391
rect -422 356 -414 391
rect -402 356 -388 391
rect -777 333 -775 356
rect -394 333 -392 356
<< nwell >>
rect -484 559 -369 863
<< nmos >>
rect -806 916 -778 946
rect -435 916 -339 946
rect -806 741 -764 771
rect -806 655 -764 685
rect -805 452 -763 482
rect -436 452 -394 482
rect -805 402 -777 432
rect -422 401 -394 431
<< pmos >>
rect -435 741 -407 771
rect -435 655 -407 685
<< ndiff >>
rect -806 991 -778 1004
rect -806 946 -778 957
rect -435 991 -339 1013
rect -435 957 -417 991
rect -383 957 -339 991
rect -435 946 -339 957
rect -806 858 -778 916
rect -435 907 -339 916
rect -435 873 -417 907
rect -383 873 -339 907
rect -435 866 -339 873
rect -806 816 -764 858
rect -806 771 -764 782
rect -806 730 -764 741
rect -806 685 -764 696
rect -806 644 -764 655
rect -806 595 -764 610
rect -805 533 -763 541
rect -805 482 -763 499
rect -436 527 -394 536
rect -436 482 -394 493
rect -805 439 -763 452
rect -805 432 -777 439
rect -436 437 -394 452
rect -422 431 -394 437
rect -805 391 -777 402
rect -805 333 -777 356
rect -422 391 -394 401
rect -422 333 -394 356
<< pdiff >>
rect -435 816 -407 826
rect -435 771 -407 782
rect -435 730 -407 741
rect -435 685 -407 696
rect -435 644 -407 655
rect -435 599 -407 610
<< ndiffc >>
rect -806 957 -778 991
rect -417 957 -383 991
rect -417 873 -383 907
rect -806 782 -764 816
rect -806 696 -764 730
rect -806 610 -764 644
rect -805 499 -763 533
rect -436 493 -394 527
rect -805 356 -777 391
rect -422 356 -394 391
<< pdiffc >>
rect -435 782 -407 816
rect -435 696 -407 730
rect -435 610 -407 644
<< poly >>
rect -887 916 -806 946
rect -778 916 -435 946
rect -339 916 -278 946
rect -887 741 -806 771
rect -764 765 -435 771
rect -764 741 -584 765
rect -593 731 -584 741
rect -550 741 -435 765
rect -407 741 -279 771
rect -550 731 -537 741
rect -593 725 -537 731
rect -697 697 -639 705
rect -697 685 -685 697
rect -933 655 -806 685
rect -764 663 -685 685
rect -651 685 -639 697
rect -651 663 -435 685
rect -764 655 -435 663
rect -407 655 -368 685
rect -933 432 -903 655
rect -839 452 -805 482
rect -763 452 -727 482
rect -551 452 -436 482
rect -394 452 -348 482
rect -933 402 -805 432
rect -777 402 -727 432
rect -309 431 -279 741
rect -551 401 -422 431
rect -394 401 -279 431
<< polycont >>
rect -584 731 -550 765
rect -685 663 -651 697
<< locali >>
rect -858 957 -806 991
rect -778 957 -727 991
rect -470 957 -417 991
rect -383 957 -278 991
rect -600 873 -584 907
rect -550 873 -417 907
rect -383 873 -278 907
rect -811 782 -806 816
rect -764 782 -435 816
rect -407 782 -364 816
rect -950 696 -934 730
rect -900 696 -806 730
rect -764 696 -759 730
rect -685 697 -651 782
rect -934 391 -899 696
rect -584 644 -550 731
rect -510 696 -435 730
rect -407 696 -279 730
rect -245 696 -229 730
rect -852 610 -806 644
rect -764 610 -584 644
rect -550 610 -435 644
rect -407 610 -367 644
rect -844 499 -805 533
rect -763 499 -716 533
rect -532 493 -436 527
rect -394 493 -350 527
rect -934 356 -805 391
rect -777 356 -422 391
rect -394 356 -355 391
<< viali >>
rect -584 873 -550 907
rect -934 696 -900 730
rect -279 696 -245 730
rect -584 610 -550 644
<< metal1 >>
rect -584 913 -550 919
rect -590 907 -544 913
rect -590 873 -584 907
rect -550 873 -544 907
rect -590 867 -544 873
rect -934 736 -900 742
rect -940 730 -894 736
rect -940 696 -934 730
rect -900 696 -894 730
rect -940 690 -894 696
rect -934 660 -900 690
rect -584 650 -550 867
rect -279 736 -245 766
rect -285 730 -239 736
rect -285 696 -279 730
rect -245 696 -239 730
rect -285 690 -239 696
rect -279 684 -245 690
rect -590 644 -544 650
rect -590 610 -584 644
rect -550 610 -544 644
rect -590 604 -544 610
rect -584 598 -550 604
<< labels >>
rlabel viali -584 610 -550 644 1 VDD
rlabel viali -584 873 -550 907 5 VDD
rlabel space -784 916 -435 946 1 WWL
rlabel ndiffc -417 957 -383 991 1 WBL
rlabel locali -532 493 -429 527 1 RBL1
rlabel poly -551 452 -490 482 1 RWL1
rlabel viali -279 696 -245 730 1 VDD
rlabel viali -934 696 -900 730 1 GND
rlabel locali -794 957 -760 991 1 WBL_b
rlabel locali -844 499 -797 533 1 RBL0
rlabel poly -763 452 -727 482 1 RWL0
<< end >>
