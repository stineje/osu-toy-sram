magic
tech sky130A
magscale 1 2
timestamp 1666997038
<< error_p >>
rect 13 2146 26 2162
rect 115 2160 128 2162
rect 81 2146 96 2160
rect 105 2146 135 2160
rect 196 2158 349 2204
rect 178 2146 370 2158
rect 413 2146 443 2160
rect 449 2146 462 2162
rect 550 2146 563 2162
rect 593 2146 606 2162
rect 695 2160 708 2162
rect 661 2146 676 2160
rect 685 2146 715 2160
rect 776 2158 929 2204
rect 758 2146 950 2158
rect 993 2146 1023 2160
rect 1029 2146 1042 2162
rect 1130 2146 1143 2162
rect 1173 2146 1186 2162
rect 1275 2160 1288 2162
rect 1241 2146 1256 2160
rect 1265 2146 1295 2160
rect 1356 2158 1509 2204
rect 1338 2146 1530 2158
rect 1573 2146 1603 2160
rect 1609 2146 1622 2162
rect 1710 2146 1723 2162
rect 1753 2146 1766 2162
rect 1855 2160 1868 2162
rect 1821 2146 1836 2160
rect 1845 2146 1875 2160
rect 1936 2158 2089 2204
rect 1918 2146 2110 2158
rect 2153 2146 2183 2160
rect 2189 2146 2202 2162
rect 2290 2146 2303 2162
rect 2333 2146 2346 2162
rect 2435 2160 2448 2162
rect 2401 2146 2416 2160
rect 2425 2146 2455 2160
rect 2516 2158 2669 2204
rect 2498 2146 2690 2158
rect 2733 2146 2763 2160
rect 2769 2146 2782 2162
rect 2870 2146 2883 2162
rect 2913 2146 2926 2162
rect 3015 2160 3028 2162
rect 2981 2146 2996 2160
rect 3005 2146 3035 2160
rect 3096 2158 3249 2204
rect 3078 2146 3270 2158
rect 3313 2146 3343 2160
rect 3349 2146 3362 2162
rect 3450 2146 3463 2162
rect 5911 2146 5924 2162
rect 6013 2160 6026 2162
rect 5979 2146 5994 2160
rect 6003 2146 6033 2160
rect 6094 2158 6247 2204
rect 6076 2146 6268 2158
rect 6311 2146 6341 2160
rect 6347 2146 6360 2162
rect 6448 2146 6461 2162
rect 6491 2146 6504 2162
rect 6593 2160 6606 2162
rect 6559 2146 6574 2160
rect 6583 2146 6613 2160
rect 6674 2158 6827 2204
rect 6656 2146 6848 2158
rect 6891 2146 6921 2160
rect 6927 2146 6940 2162
rect 7028 2146 7041 2162
rect 7071 2146 7084 2162
rect 7173 2160 7186 2162
rect 7139 2146 7154 2160
rect 7163 2146 7193 2160
rect 7254 2158 7407 2204
rect 7236 2146 7428 2158
rect 7471 2146 7501 2160
rect 7507 2146 7520 2162
rect 7608 2146 7621 2162
rect 7651 2146 7664 2162
rect 7753 2160 7766 2162
rect 7719 2146 7734 2160
rect 7743 2146 7773 2160
rect 7834 2158 7987 2204
rect 7816 2146 8008 2158
rect 8051 2146 8081 2160
rect 8087 2146 8100 2162
rect 8188 2146 8201 2162
rect 8231 2146 8244 2162
rect 8333 2160 8346 2162
rect 8299 2146 8314 2160
rect 8323 2146 8353 2160
rect 8414 2158 8567 2204
rect 8396 2146 8588 2158
rect 8631 2146 8661 2160
rect 8667 2146 8680 2162
rect 8768 2146 8781 2162
rect 8811 2146 8824 2162
rect 8913 2160 8926 2162
rect 8879 2146 8894 2160
rect 8903 2146 8933 2160
rect 8994 2158 9147 2204
rect 8976 2146 9168 2158
rect 9211 2146 9241 2160
rect 9247 2146 9260 2162
rect 9348 2146 9361 2162
rect -2 2132 3469 2146
rect 5889 2132 9361 2146
rect 13 2028 26 2132
rect 71 2110 72 2120
rect 87 2110 100 2120
rect 71 2106 100 2110
rect 105 2106 135 2132
rect 153 2118 169 2120
rect 241 2118 294 2132
rect 242 2116 306 2118
rect 349 2116 364 2132
rect 413 2129 443 2132
rect 413 2126 449 2129
rect 379 2118 395 2120
rect 153 2106 168 2110
rect 71 2104 168 2106
rect 196 2104 364 2116
rect 380 2106 395 2110
rect 413 2107 452 2126
rect 471 2120 478 2121
rect 477 2113 478 2120
rect 461 2110 462 2113
rect 477 2110 490 2113
rect 413 2106 443 2107
rect 452 2106 458 2107
rect 461 2106 490 2110
rect 380 2105 490 2106
rect 380 2104 496 2105
rect 55 2096 106 2104
rect 55 2084 80 2096
rect 87 2084 106 2096
rect 137 2096 187 2104
rect 137 2088 153 2096
rect 160 2094 187 2096
rect 196 2094 417 2104
rect 160 2084 417 2094
rect 446 2096 496 2104
rect 446 2087 462 2096
rect 55 2076 106 2084
rect 153 2076 417 2084
rect 443 2084 462 2087
rect 469 2084 496 2096
rect 443 2076 496 2084
rect 71 2068 72 2076
rect 87 2068 100 2076
rect 71 2060 87 2068
rect 68 2053 87 2056
rect 68 2044 90 2053
rect 41 2034 90 2044
rect 41 2028 71 2034
rect 90 2029 95 2034
rect 13 2012 87 2028
rect 105 2020 135 2076
rect 170 2066 378 2076
rect 413 2072 458 2076
rect 461 2075 462 2076
rect 477 2075 490 2076
rect 196 2036 385 2066
rect 211 2033 385 2036
rect 204 2030 385 2033
rect 13 2010 26 2012
rect 41 2010 75 2012
rect 13 1994 87 2010
rect 114 2006 127 2020
rect 142 2006 158 2022
rect 204 2017 215 2030
rect -3 1972 -2 1988
rect 13 1972 26 1994
rect 41 1972 71 1994
rect 114 1990 176 2006
rect 204 1999 215 2015
rect 220 2010 230 2030
rect 240 2010 254 2030
rect 257 2017 266 2030
rect 282 2017 291 2030
rect 220 1999 254 2010
rect 257 1999 266 2015
rect 282 1999 291 2015
rect 298 2010 308 2030
rect 318 2010 332 2030
rect 333 2017 344 2030
rect 298 1999 332 2010
rect 333 1999 344 2015
rect 390 2006 406 2022
rect 413 2020 443 2072
rect 477 2068 478 2075
rect 462 2060 478 2068
rect 449 2028 462 2047
rect 477 2028 507 2044
rect 449 2012 523 2028
rect 449 2010 462 2012
rect 477 2010 511 2012
rect 114 1988 127 1990
rect 142 1988 176 1990
rect 114 1972 176 1988
rect 220 1983 236 1986
rect 298 1983 328 1994
rect 376 1990 422 2006
rect 449 1994 523 2010
rect 376 1988 410 1990
rect 375 1972 422 1988
rect 449 1972 462 1994
rect 477 1972 507 1994
rect 534 1972 535 1988
rect 550 1972 563 2132
rect 593 2028 606 2132
rect 651 2110 652 2120
rect 667 2110 680 2120
rect 651 2106 680 2110
rect 685 2106 715 2132
rect 733 2118 749 2120
rect 821 2118 874 2132
rect 822 2116 886 2118
rect 929 2116 944 2132
rect 993 2129 1023 2132
rect 993 2126 1029 2129
rect 959 2118 975 2120
rect 733 2106 748 2110
rect 651 2104 748 2106
rect 776 2104 944 2116
rect 960 2106 975 2110
rect 993 2107 1032 2126
rect 1051 2120 1058 2121
rect 1057 2113 1058 2120
rect 1041 2110 1042 2113
rect 1057 2110 1070 2113
rect 993 2106 1023 2107
rect 1032 2106 1038 2107
rect 1041 2106 1070 2110
rect 960 2105 1070 2106
rect 960 2104 1076 2105
rect 635 2096 686 2104
rect 635 2084 660 2096
rect 667 2084 686 2096
rect 717 2096 767 2104
rect 717 2088 733 2096
rect 740 2094 767 2096
rect 776 2094 997 2104
rect 740 2084 997 2094
rect 1026 2096 1076 2104
rect 1026 2087 1042 2096
rect 635 2076 686 2084
rect 733 2076 997 2084
rect 1023 2084 1042 2087
rect 1049 2084 1076 2096
rect 1023 2076 1076 2084
rect 651 2068 652 2076
rect 667 2068 680 2076
rect 651 2060 667 2068
rect 648 2053 667 2056
rect 648 2044 670 2053
rect 621 2034 670 2044
rect 621 2028 651 2034
rect 670 2029 675 2034
rect 593 2012 667 2028
rect 685 2020 715 2076
rect 750 2066 958 2076
rect 993 2072 1038 2076
rect 1041 2075 1042 2076
rect 1057 2075 1070 2076
rect 776 2036 965 2066
rect 791 2033 965 2036
rect 784 2030 965 2033
rect 593 2010 606 2012
rect 621 2010 655 2012
rect 593 1994 667 2010
rect 694 2006 707 2020
rect 722 2006 738 2022
rect 784 2017 795 2030
rect 577 1972 578 1988
rect 593 1972 606 1994
rect 621 1972 651 1994
rect 694 1990 756 2006
rect 784 1999 795 2015
rect 800 2010 810 2030
rect 820 2010 834 2030
rect 837 2017 846 2030
rect 862 2017 871 2030
rect 800 1999 834 2010
rect 837 1999 846 2015
rect 862 1999 871 2015
rect 878 2010 888 2030
rect 898 2010 912 2030
rect 913 2017 924 2030
rect 878 1999 912 2010
rect 913 1999 924 2015
rect 970 2006 986 2022
rect 993 2020 1023 2072
rect 1057 2068 1058 2075
rect 1042 2060 1058 2068
rect 1029 2028 1042 2047
rect 1057 2028 1087 2044
rect 1029 2012 1103 2028
rect 1029 2010 1042 2012
rect 1057 2010 1091 2012
rect 694 1988 707 1990
rect 722 1988 756 1990
rect 694 1972 756 1988
rect 800 1983 816 1986
rect 878 1983 908 1994
rect 956 1990 1002 2006
rect 1029 1994 1103 2010
rect 956 1988 990 1990
rect 955 1972 1002 1988
rect 1029 1972 1042 1994
rect 1057 1972 1087 1994
rect 1114 1972 1115 1988
rect 1130 1972 1143 2132
rect 1173 2028 1186 2132
rect 1231 2110 1232 2120
rect 1247 2110 1260 2120
rect 1231 2106 1260 2110
rect 1265 2106 1295 2132
rect 1313 2118 1329 2120
rect 1401 2118 1454 2132
rect 1402 2116 1466 2118
rect 1509 2116 1524 2132
rect 1573 2129 1603 2132
rect 1573 2126 1609 2129
rect 1539 2118 1555 2120
rect 1313 2106 1328 2110
rect 1231 2104 1328 2106
rect 1356 2104 1524 2116
rect 1540 2106 1555 2110
rect 1573 2107 1612 2126
rect 1631 2120 1638 2121
rect 1637 2113 1638 2120
rect 1621 2110 1622 2113
rect 1637 2110 1650 2113
rect 1573 2106 1603 2107
rect 1612 2106 1618 2107
rect 1621 2106 1650 2110
rect 1540 2105 1650 2106
rect 1540 2104 1656 2105
rect 1215 2096 1266 2104
rect 1215 2084 1240 2096
rect 1247 2084 1266 2096
rect 1297 2096 1347 2104
rect 1297 2088 1313 2096
rect 1320 2094 1347 2096
rect 1356 2094 1577 2104
rect 1320 2084 1577 2094
rect 1606 2096 1656 2104
rect 1606 2087 1622 2096
rect 1215 2076 1266 2084
rect 1313 2076 1577 2084
rect 1603 2084 1622 2087
rect 1629 2084 1656 2096
rect 1603 2076 1656 2084
rect 1231 2068 1232 2076
rect 1247 2068 1260 2076
rect 1231 2060 1247 2068
rect 1228 2053 1247 2056
rect 1228 2044 1250 2053
rect 1201 2034 1250 2044
rect 1201 2028 1231 2034
rect 1250 2029 1255 2034
rect 1173 2012 1247 2028
rect 1265 2020 1295 2076
rect 1330 2066 1538 2076
rect 1573 2072 1618 2076
rect 1621 2075 1622 2076
rect 1637 2075 1650 2076
rect 1356 2036 1545 2066
rect 1371 2033 1545 2036
rect 1364 2030 1545 2033
rect 1173 2010 1186 2012
rect 1201 2010 1235 2012
rect 1173 1994 1247 2010
rect 1274 2006 1287 2020
rect 1302 2006 1318 2022
rect 1364 2017 1375 2030
rect 1157 1972 1158 1988
rect 1173 1972 1186 1994
rect 1201 1972 1231 1994
rect 1274 1990 1336 2006
rect 1364 1999 1375 2015
rect 1380 2010 1390 2030
rect 1400 2010 1414 2030
rect 1417 2017 1426 2030
rect 1442 2017 1451 2030
rect 1380 1999 1414 2010
rect 1417 1999 1426 2015
rect 1442 1999 1451 2015
rect 1458 2010 1468 2030
rect 1478 2010 1492 2030
rect 1493 2017 1504 2030
rect 1458 1999 1492 2010
rect 1493 1999 1504 2015
rect 1550 2006 1566 2022
rect 1573 2020 1603 2072
rect 1637 2068 1638 2075
rect 1622 2060 1638 2068
rect 1609 2028 1622 2047
rect 1637 2028 1667 2044
rect 1609 2012 1683 2028
rect 1609 2010 1622 2012
rect 1637 2010 1671 2012
rect 1274 1988 1287 1990
rect 1302 1988 1336 1990
rect 1274 1972 1336 1988
rect 1380 1983 1396 1986
rect 1458 1983 1488 1994
rect 1536 1990 1582 2006
rect 1609 1994 1683 2010
rect 1536 1988 1570 1990
rect 1535 1972 1582 1988
rect 1609 1972 1622 1994
rect 1637 1972 1667 1994
rect 1694 1972 1695 1988
rect 1710 1972 1723 2132
rect 1753 2028 1766 2132
rect 1811 2110 1812 2120
rect 1827 2110 1840 2120
rect 1811 2106 1840 2110
rect 1845 2106 1875 2132
rect 1893 2118 1909 2120
rect 1981 2118 2034 2132
rect 1982 2116 2046 2118
rect 2089 2116 2104 2132
rect 2153 2129 2183 2132
rect 2153 2126 2189 2129
rect 2119 2118 2135 2120
rect 1893 2106 1908 2110
rect 1811 2104 1908 2106
rect 1936 2104 2104 2116
rect 2120 2106 2135 2110
rect 2153 2107 2192 2126
rect 2211 2120 2218 2121
rect 2217 2113 2218 2120
rect 2201 2110 2202 2113
rect 2217 2110 2230 2113
rect 2153 2106 2183 2107
rect 2192 2106 2198 2107
rect 2201 2106 2230 2110
rect 2120 2105 2230 2106
rect 2120 2104 2236 2105
rect 1795 2096 1846 2104
rect 1795 2084 1820 2096
rect 1827 2084 1846 2096
rect 1877 2096 1927 2104
rect 1877 2088 1893 2096
rect 1900 2094 1927 2096
rect 1936 2094 2157 2104
rect 1900 2084 2157 2094
rect 2186 2096 2236 2104
rect 2186 2087 2202 2096
rect 1795 2076 1846 2084
rect 1893 2076 2157 2084
rect 2183 2084 2202 2087
rect 2209 2084 2236 2096
rect 2183 2076 2236 2084
rect 1811 2068 1812 2076
rect 1827 2068 1840 2076
rect 1811 2060 1827 2068
rect 1808 2053 1827 2056
rect 1808 2044 1830 2053
rect 1781 2034 1830 2044
rect 1781 2028 1811 2034
rect 1830 2029 1835 2034
rect 1753 2012 1827 2028
rect 1845 2020 1875 2076
rect 1910 2066 2118 2076
rect 2153 2072 2198 2076
rect 2201 2075 2202 2076
rect 2217 2075 2230 2076
rect 1936 2036 2125 2066
rect 1951 2033 2125 2036
rect 1944 2030 2125 2033
rect 1753 2010 1766 2012
rect 1781 2010 1815 2012
rect 1753 1994 1827 2010
rect 1854 2006 1867 2020
rect 1882 2006 1898 2022
rect 1944 2017 1955 2030
rect 1737 1972 1738 1988
rect 1753 1972 1766 1994
rect 1781 1972 1811 1994
rect 1854 1990 1916 2006
rect 1944 1999 1955 2015
rect 1960 2010 1970 2030
rect 1980 2010 1994 2030
rect 1997 2017 2006 2030
rect 2022 2017 2031 2030
rect 1960 1999 1994 2010
rect 1997 1999 2006 2015
rect 2022 1999 2031 2015
rect 2038 2010 2048 2030
rect 2058 2010 2072 2030
rect 2073 2017 2084 2030
rect 2038 1999 2072 2010
rect 2073 1999 2084 2015
rect 2130 2006 2146 2022
rect 2153 2020 2183 2072
rect 2217 2068 2218 2075
rect 2202 2060 2218 2068
rect 2189 2028 2202 2047
rect 2217 2028 2247 2044
rect 2189 2012 2263 2028
rect 2189 2010 2202 2012
rect 2217 2010 2251 2012
rect 1854 1988 1867 1990
rect 1882 1988 1916 1990
rect 1854 1972 1916 1988
rect 1960 1983 1976 1986
rect 2038 1983 2068 1994
rect 2116 1990 2162 2006
rect 2189 1994 2263 2010
rect 2116 1988 2150 1990
rect 2115 1972 2162 1988
rect 2189 1972 2202 1994
rect 2217 1972 2247 1994
rect 2274 1972 2275 1988
rect 2290 1972 2303 2132
rect 2333 2028 2346 2132
rect 2391 2110 2392 2120
rect 2407 2110 2420 2120
rect 2391 2106 2420 2110
rect 2425 2106 2455 2132
rect 2473 2118 2489 2120
rect 2561 2118 2614 2132
rect 2562 2116 2626 2118
rect 2669 2116 2684 2132
rect 2733 2129 2763 2132
rect 2733 2126 2769 2129
rect 2699 2118 2715 2120
rect 2473 2106 2488 2110
rect 2391 2104 2488 2106
rect 2516 2104 2684 2116
rect 2700 2106 2715 2110
rect 2733 2107 2772 2126
rect 2791 2120 2798 2121
rect 2797 2113 2798 2120
rect 2781 2110 2782 2113
rect 2797 2110 2810 2113
rect 2733 2106 2763 2107
rect 2772 2106 2778 2107
rect 2781 2106 2810 2110
rect 2700 2105 2810 2106
rect 2700 2104 2816 2105
rect 2375 2096 2426 2104
rect 2375 2084 2400 2096
rect 2407 2084 2426 2096
rect 2457 2096 2507 2104
rect 2457 2088 2473 2096
rect 2480 2094 2507 2096
rect 2516 2094 2737 2104
rect 2480 2084 2737 2094
rect 2766 2096 2816 2104
rect 2766 2087 2782 2096
rect 2375 2076 2426 2084
rect 2473 2076 2737 2084
rect 2763 2084 2782 2087
rect 2789 2084 2816 2096
rect 2763 2076 2816 2084
rect 2391 2068 2392 2076
rect 2407 2068 2420 2076
rect 2391 2060 2407 2068
rect 2388 2053 2407 2056
rect 2388 2044 2410 2053
rect 2361 2034 2410 2044
rect 2361 2028 2391 2034
rect 2410 2029 2415 2034
rect 2333 2012 2407 2028
rect 2425 2020 2455 2076
rect 2490 2066 2698 2076
rect 2733 2072 2778 2076
rect 2781 2075 2782 2076
rect 2797 2075 2810 2076
rect 2516 2036 2705 2066
rect 2531 2033 2705 2036
rect 2524 2030 2705 2033
rect 2333 2010 2346 2012
rect 2361 2010 2395 2012
rect 2333 1994 2407 2010
rect 2434 2006 2447 2020
rect 2462 2006 2478 2022
rect 2524 2017 2535 2030
rect 2317 1972 2318 1988
rect 2333 1972 2346 1994
rect 2361 1972 2391 1994
rect 2434 1990 2496 2006
rect 2524 1999 2535 2015
rect 2540 2010 2550 2030
rect 2560 2010 2574 2030
rect 2577 2017 2586 2030
rect 2602 2017 2611 2030
rect 2540 1999 2574 2010
rect 2577 1999 2586 2015
rect 2602 1999 2611 2015
rect 2618 2010 2628 2030
rect 2638 2010 2652 2030
rect 2653 2017 2664 2030
rect 2618 1999 2652 2010
rect 2653 1999 2664 2015
rect 2710 2006 2726 2022
rect 2733 2020 2763 2072
rect 2797 2068 2798 2075
rect 2782 2060 2798 2068
rect 2769 2028 2782 2047
rect 2797 2028 2827 2044
rect 2769 2012 2843 2028
rect 2769 2010 2782 2012
rect 2797 2010 2831 2012
rect 2434 1988 2447 1990
rect 2462 1988 2496 1990
rect 2434 1972 2496 1988
rect 2540 1983 2556 1986
rect 2618 1983 2648 1994
rect 2696 1990 2742 2006
rect 2769 1994 2843 2010
rect 2696 1988 2730 1990
rect 2695 1972 2742 1988
rect 2769 1972 2782 1994
rect 2797 1972 2827 1994
rect 2854 1972 2855 1988
rect 2870 1972 2883 2132
rect 2913 2028 2926 2132
rect 2971 2110 2972 2120
rect 2987 2110 3000 2120
rect 2971 2106 3000 2110
rect 3005 2106 3035 2132
rect 3053 2118 3069 2120
rect 3141 2118 3194 2132
rect 3142 2116 3206 2118
rect 3249 2116 3264 2132
rect 3313 2129 3343 2132
rect 3313 2126 3349 2129
rect 3279 2118 3295 2120
rect 3053 2106 3068 2110
rect 2971 2104 3068 2106
rect 3096 2104 3264 2116
rect 3280 2106 3295 2110
rect 3313 2107 3352 2126
rect 3371 2120 3378 2121
rect 3377 2113 3378 2120
rect 3361 2110 3362 2113
rect 3377 2110 3390 2113
rect 3313 2106 3343 2107
rect 3352 2106 3358 2107
rect 3361 2106 3390 2110
rect 3280 2105 3390 2106
rect 3280 2104 3396 2105
rect 2955 2096 3006 2104
rect 2955 2084 2980 2096
rect 2987 2084 3006 2096
rect 3037 2096 3087 2104
rect 3037 2088 3053 2096
rect 3060 2094 3087 2096
rect 3096 2094 3317 2104
rect 3060 2084 3317 2094
rect 3346 2096 3396 2104
rect 3346 2087 3362 2096
rect 2955 2076 3006 2084
rect 3053 2076 3317 2084
rect 3343 2084 3362 2087
rect 3369 2084 3396 2096
rect 3343 2076 3396 2084
rect 2971 2068 2972 2076
rect 2987 2068 3000 2076
rect 2971 2060 2987 2068
rect 2968 2053 2987 2056
rect 2968 2044 2990 2053
rect 2941 2034 2990 2044
rect 2941 2028 2971 2034
rect 2990 2029 2995 2034
rect 2913 2012 2987 2028
rect 3005 2020 3035 2076
rect 3070 2066 3278 2076
rect 3313 2072 3358 2076
rect 3361 2075 3362 2076
rect 3377 2075 3390 2076
rect 3096 2036 3285 2066
rect 3111 2033 3285 2036
rect 3104 2030 3285 2033
rect 2913 2010 2926 2012
rect 2941 2010 2975 2012
rect 2913 1994 2987 2010
rect 3014 2006 3027 2020
rect 3042 2006 3058 2022
rect 3104 2017 3115 2030
rect 2897 1972 2898 1988
rect 2913 1972 2926 1994
rect 2941 1972 2971 1994
rect 3014 1990 3076 2006
rect 3104 1999 3115 2015
rect 3120 2010 3130 2030
rect 3140 2010 3154 2030
rect 3157 2017 3166 2030
rect 3182 2017 3191 2030
rect 3120 1999 3154 2010
rect 3157 1999 3166 2015
rect 3182 1999 3191 2015
rect 3198 2010 3208 2030
rect 3218 2010 3232 2030
rect 3233 2017 3244 2030
rect 3198 1999 3232 2010
rect 3233 1999 3244 2015
rect 3290 2006 3306 2022
rect 3313 2020 3343 2072
rect 3377 2068 3378 2075
rect 3362 2060 3378 2068
rect 3349 2028 3362 2047
rect 3377 2028 3407 2044
rect 3349 2012 3423 2028
rect 3349 2010 3362 2012
rect 3377 2010 3411 2012
rect 3014 1988 3027 1990
rect 3042 1988 3076 1990
rect 3014 1972 3076 1988
rect 3120 1983 3136 1986
rect 3198 1983 3228 1994
rect 3276 1990 3322 2006
rect 3349 1994 3423 2010
rect 3276 1988 3310 1990
rect 3275 1972 3322 1988
rect 3349 1972 3362 1994
rect 3377 1972 3407 1994
rect 3434 1972 3435 1988
rect 3450 1972 3463 2132
rect 5911 2028 5924 2132
rect 5969 2110 5970 2120
rect 5985 2110 5998 2120
rect 5969 2106 5998 2110
rect 6003 2106 6033 2132
rect 6051 2118 6067 2120
rect 6139 2118 6192 2132
rect 6140 2116 6204 2118
rect 6247 2116 6262 2132
rect 6311 2129 6341 2132
rect 6311 2126 6347 2129
rect 6277 2118 6293 2120
rect 6051 2106 6066 2110
rect 5969 2104 6066 2106
rect 6094 2104 6262 2116
rect 6278 2106 6293 2110
rect 6311 2107 6350 2126
rect 6369 2120 6376 2121
rect 6375 2113 6376 2120
rect 6359 2110 6360 2113
rect 6375 2110 6388 2113
rect 6311 2106 6341 2107
rect 6350 2106 6356 2107
rect 6359 2106 6388 2110
rect 6278 2105 6388 2106
rect 6278 2104 6394 2105
rect 5953 2096 6004 2104
rect 5953 2084 5978 2096
rect 5985 2084 6004 2096
rect 6035 2096 6085 2104
rect 6035 2088 6051 2096
rect 6058 2094 6085 2096
rect 6094 2094 6315 2104
rect 6058 2084 6315 2094
rect 6344 2096 6394 2104
rect 6344 2087 6360 2096
rect 5953 2076 6004 2084
rect 6051 2076 6315 2084
rect 6341 2084 6360 2087
rect 6367 2084 6394 2096
rect 6341 2076 6394 2084
rect 5969 2068 5970 2076
rect 5985 2068 5998 2076
rect 5969 2060 5985 2068
rect 5966 2053 5985 2056
rect 5966 2044 5988 2053
rect 5939 2034 5988 2044
rect 5939 2028 5969 2034
rect 5988 2029 5993 2034
rect 5911 2012 5985 2028
rect 6003 2020 6033 2076
rect 6068 2066 6276 2076
rect 6311 2072 6356 2076
rect 6359 2075 6360 2076
rect 6375 2075 6388 2076
rect 6094 2036 6283 2066
rect 6109 2033 6283 2036
rect 6102 2030 6283 2033
rect 5911 2010 5924 2012
rect 5939 2010 5973 2012
rect 5911 1994 5985 2010
rect 6012 2006 6025 2020
rect 6040 2006 6056 2022
rect 6102 2017 6113 2030
rect 5895 1972 5896 1988
rect 5911 1972 5924 1994
rect 5939 1972 5969 1994
rect 6012 1990 6074 2006
rect 6102 1999 6113 2015
rect 6118 2010 6128 2030
rect 6138 2010 6152 2030
rect 6155 2017 6164 2030
rect 6180 2017 6189 2030
rect 6118 1999 6152 2010
rect 6155 1999 6164 2015
rect 6180 1999 6189 2015
rect 6196 2010 6206 2030
rect 6216 2010 6230 2030
rect 6231 2017 6242 2030
rect 6196 1999 6230 2010
rect 6231 1999 6242 2015
rect 6288 2006 6304 2022
rect 6311 2020 6341 2072
rect 6375 2068 6376 2075
rect 6360 2060 6376 2068
rect 6347 2028 6360 2047
rect 6375 2028 6405 2044
rect 6347 2012 6421 2028
rect 6347 2010 6360 2012
rect 6375 2010 6409 2012
rect 6012 1988 6025 1990
rect 6040 1988 6074 1990
rect 6012 1972 6074 1988
rect 6118 1983 6134 1986
rect 6196 1983 6226 1994
rect 6274 1990 6320 2006
rect 6347 1994 6421 2010
rect 6274 1988 6308 1990
rect 6273 1972 6320 1988
rect 6347 1972 6360 1994
rect 6375 1972 6405 1994
rect 6432 1972 6433 1988
rect 6448 1972 6461 2132
rect 6491 2028 6504 2132
rect 6549 2110 6550 2120
rect 6565 2110 6578 2120
rect 6549 2106 6578 2110
rect 6583 2106 6613 2132
rect 6631 2118 6647 2120
rect 6719 2118 6772 2132
rect 6720 2116 6784 2118
rect 6827 2116 6842 2132
rect 6891 2129 6921 2132
rect 6891 2126 6927 2129
rect 6857 2118 6873 2120
rect 6631 2106 6646 2110
rect 6549 2104 6646 2106
rect 6674 2104 6842 2116
rect 6858 2106 6873 2110
rect 6891 2107 6930 2126
rect 6949 2120 6956 2121
rect 6955 2113 6956 2120
rect 6939 2110 6940 2113
rect 6955 2110 6968 2113
rect 6891 2106 6921 2107
rect 6930 2106 6936 2107
rect 6939 2106 6968 2110
rect 6858 2105 6968 2106
rect 6858 2104 6974 2105
rect 6533 2096 6584 2104
rect 6533 2084 6558 2096
rect 6565 2084 6584 2096
rect 6615 2096 6665 2104
rect 6615 2088 6631 2096
rect 6638 2094 6665 2096
rect 6674 2094 6895 2104
rect 6638 2084 6895 2094
rect 6924 2096 6974 2104
rect 6924 2087 6940 2096
rect 6533 2076 6584 2084
rect 6631 2076 6895 2084
rect 6921 2084 6940 2087
rect 6947 2084 6974 2096
rect 6921 2076 6974 2084
rect 6549 2068 6550 2076
rect 6565 2068 6578 2076
rect 6549 2060 6565 2068
rect 6546 2053 6565 2056
rect 6546 2044 6568 2053
rect 6519 2034 6568 2044
rect 6519 2028 6549 2034
rect 6568 2029 6573 2034
rect 6491 2012 6565 2028
rect 6583 2020 6613 2076
rect 6648 2066 6856 2076
rect 6891 2072 6936 2076
rect 6939 2075 6940 2076
rect 6955 2075 6968 2076
rect 6674 2036 6863 2066
rect 6689 2033 6863 2036
rect 6682 2030 6863 2033
rect 6491 2010 6504 2012
rect 6519 2010 6553 2012
rect 6491 1994 6565 2010
rect 6592 2006 6605 2020
rect 6620 2006 6636 2022
rect 6682 2017 6693 2030
rect 6475 1972 6476 1988
rect 6491 1972 6504 1994
rect 6519 1972 6549 1994
rect 6592 1990 6654 2006
rect 6682 1999 6693 2015
rect 6698 2010 6708 2030
rect 6718 2010 6732 2030
rect 6735 2017 6744 2030
rect 6760 2017 6769 2030
rect 6698 1999 6732 2010
rect 6735 1999 6744 2015
rect 6760 1999 6769 2015
rect 6776 2010 6786 2030
rect 6796 2010 6810 2030
rect 6811 2017 6822 2030
rect 6776 1999 6810 2010
rect 6811 1999 6822 2015
rect 6868 2006 6884 2022
rect 6891 2020 6921 2072
rect 6955 2068 6956 2075
rect 6940 2060 6956 2068
rect 6927 2028 6940 2047
rect 6955 2028 6985 2044
rect 6927 2012 7001 2028
rect 6927 2010 6940 2012
rect 6955 2010 6989 2012
rect 6592 1988 6605 1990
rect 6620 1988 6654 1990
rect 6592 1972 6654 1988
rect 6698 1983 6714 1986
rect 6776 1983 6806 1994
rect 6854 1990 6900 2006
rect 6927 1994 7001 2010
rect 6854 1988 6888 1990
rect 6853 1972 6900 1988
rect 6927 1972 6940 1994
rect 6955 1972 6985 1994
rect 7012 1972 7013 1988
rect 7028 1972 7041 2132
rect 7071 2028 7084 2132
rect 7129 2110 7130 2120
rect 7145 2110 7158 2120
rect 7129 2106 7158 2110
rect 7163 2106 7193 2132
rect 7211 2118 7227 2120
rect 7299 2118 7352 2132
rect 7300 2116 7364 2118
rect 7407 2116 7422 2132
rect 7471 2129 7501 2132
rect 7471 2126 7507 2129
rect 7437 2118 7453 2120
rect 7211 2106 7226 2110
rect 7129 2104 7226 2106
rect 7254 2104 7422 2116
rect 7438 2106 7453 2110
rect 7471 2107 7510 2126
rect 7529 2120 7536 2121
rect 7535 2113 7536 2120
rect 7519 2110 7520 2113
rect 7535 2110 7548 2113
rect 7471 2106 7501 2107
rect 7510 2106 7516 2107
rect 7519 2106 7548 2110
rect 7438 2105 7548 2106
rect 7438 2104 7554 2105
rect 7113 2096 7164 2104
rect 7113 2084 7138 2096
rect 7145 2084 7164 2096
rect 7195 2096 7245 2104
rect 7195 2088 7211 2096
rect 7218 2094 7245 2096
rect 7254 2094 7475 2104
rect 7218 2084 7475 2094
rect 7504 2096 7554 2104
rect 7504 2087 7520 2096
rect 7113 2076 7164 2084
rect 7211 2076 7475 2084
rect 7501 2084 7520 2087
rect 7527 2084 7554 2096
rect 7501 2076 7554 2084
rect 7129 2068 7130 2076
rect 7145 2068 7158 2076
rect 7129 2060 7145 2068
rect 7126 2053 7145 2056
rect 7126 2044 7148 2053
rect 7099 2034 7148 2044
rect 7099 2028 7129 2034
rect 7148 2029 7153 2034
rect 7071 2012 7145 2028
rect 7163 2020 7193 2076
rect 7228 2066 7436 2076
rect 7471 2072 7516 2076
rect 7519 2075 7520 2076
rect 7535 2075 7548 2076
rect 7254 2036 7443 2066
rect 7269 2033 7443 2036
rect 7262 2030 7443 2033
rect 7071 2010 7084 2012
rect 7099 2010 7133 2012
rect 7071 1994 7145 2010
rect 7172 2006 7185 2020
rect 7200 2006 7216 2022
rect 7262 2017 7273 2030
rect 7055 1972 7056 1988
rect 7071 1972 7084 1994
rect 7099 1972 7129 1994
rect 7172 1990 7234 2006
rect 7262 1999 7273 2015
rect 7278 2010 7288 2030
rect 7298 2010 7312 2030
rect 7315 2017 7324 2030
rect 7340 2017 7349 2030
rect 7278 1999 7312 2010
rect 7315 1999 7324 2015
rect 7340 1999 7349 2015
rect 7356 2010 7366 2030
rect 7376 2010 7390 2030
rect 7391 2017 7402 2030
rect 7356 1999 7390 2010
rect 7391 1999 7402 2015
rect 7448 2006 7464 2022
rect 7471 2020 7501 2072
rect 7535 2068 7536 2075
rect 7520 2060 7536 2068
rect 7507 2028 7520 2047
rect 7535 2028 7565 2044
rect 7507 2012 7581 2028
rect 7507 2010 7520 2012
rect 7535 2010 7569 2012
rect 7172 1988 7185 1990
rect 7200 1988 7234 1990
rect 7172 1972 7234 1988
rect 7278 1983 7294 1986
rect 7356 1983 7386 1994
rect 7434 1990 7480 2006
rect 7507 1994 7581 2010
rect 7434 1988 7468 1990
rect 7433 1972 7480 1988
rect 7507 1972 7520 1994
rect 7535 1972 7565 1994
rect 7592 1972 7593 1988
rect 7608 1972 7621 2132
rect 7651 2028 7664 2132
rect 7709 2110 7710 2120
rect 7725 2110 7738 2120
rect 7709 2106 7738 2110
rect 7743 2106 7773 2132
rect 7791 2118 7807 2120
rect 7879 2118 7932 2132
rect 7880 2116 7944 2118
rect 7987 2116 8002 2132
rect 8051 2129 8081 2132
rect 8051 2126 8087 2129
rect 8017 2118 8033 2120
rect 7791 2106 7806 2110
rect 7709 2104 7806 2106
rect 7834 2104 8002 2116
rect 8018 2106 8033 2110
rect 8051 2107 8090 2126
rect 8109 2120 8116 2121
rect 8115 2113 8116 2120
rect 8099 2110 8100 2113
rect 8115 2110 8128 2113
rect 8051 2106 8081 2107
rect 8090 2106 8096 2107
rect 8099 2106 8128 2110
rect 8018 2105 8128 2106
rect 8018 2104 8134 2105
rect 7693 2096 7744 2104
rect 7693 2084 7718 2096
rect 7725 2084 7744 2096
rect 7775 2096 7825 2104
rect 7775 2088 7791 2096
rect 7798 2094 7825 2096
rect 7834 2094 8055 2104
rect 7798 2084 8055 2094
rect 8084 2096 8134 2104
rect 8084 2087 8100 2096
rect 7693 2076 7744 2084
rect 7791 2076 8055 2084
rect 8081 2084 8100 2087
rect 8107 2084 8134 2096
rect 8081 2076 8134 2084
rect 7709 2068 7710 2076
rect 7725 2068 7738 2076
rect 7709 2060 7725 2068
rect 7706 2053 7725 2056
rect 7706 2044 7728 2053
rect 7679 2034 7728 2044
rect 7679 2028 7709 2034
rect 7728 2029 7733 2034
rect 7651 2012 7725 2028
rect 7743 2020 7773 2076
rect 7808 2066 8016 2076
rect 8051 2072 8096 2076
rect 8099 2075 8100 2076
rect 8115 2075 8128 2076
rect 7834 2036 8023 2066
rect 7849 2033 8023 2036
rect 7842 2030 8023 2033
rect 7651 2010 7664 2012
rect 7679 2010 7713 2012
rect 7651 1994 7725 2010
rect 7752 2006 7765 2020
rect 7780 2006 7796 2022
rect 7842 2017 7853 2030
rect 7635 1972 7636 1988
rect 7651 1972 7664 1994
rect 7679 1972 7709 1994
rect 7752 1990 7814 2006
rect 7842 1999 7853 2015
rect 7858 2010 7868 2030
rect 7878 2010 7892 2030
rect 7895 2017 7904 2030
rect 7920 2017 7929 2030
rect 7858 1999 7892 2010
rect 7895 1999 7904 2015
rect 7920 1999 7929 2015
rect 7936 2010 7946 2030
rect 7956 2010 7970 2030
rect 7971 2017 7982 2030
rect 7936 1999 7970 2010
rect 7971 1999 7982 2015
rect 8028 2006 8044 2022
rect 8051 2020 8081 2072
rect 8115 2068 8116 2075
rect 8100 2060 8116 2068
rect 8087 2028 8100 2047
rect 8115 2028 8145 2044
rect 8087 2012 8161 2028
rect 8087 2010 8100 2012
rect 8115 2010 8149 2012
rect 7752 1988 7765 1990
rect 7780 1988 7814 1990
rect 7752 1972 7814 1988
rect 7858 1983 7874 1986
rect 7936 1983 7966 1994
rect 8014 1990 8060 2006
rect 8087 1994 8161 2010
rect 8014 1988 8048 1990
rect 8013 1972 8060 1988
rect 8087 1972 8100 1994
rect 8115 1972 8145 1994
rect 8172 1972 8173 1988
rect 8188 1972 8201 2132
rect 8231 2028 8244 2132
rect 8289 2110 8290 2120
rect 8305 2110 8318 2120
rect 8289 2106 8318 2110
rect 8323 2106 8353 2132
rect 8371 2118 8387 2120
rect 8459 2118 8512 2132
rect 8460 2116 8524 2118
rect 8567 2116 8582 2132
rect 8631 2129 8661 2132
rect 8631 2126 8667 2129
rect 8597 2118 8613 2120
rect 8371 2106 8386 2110
rect 8289 2104 8386 2106
rect 8414 2104 8582 2116
rect 8598 2106 8613 2110
rect 8631 2107 8670 2126
rect 8689 2120 8696 2121
rect 8695 2113 8696 2120
rect 8679 2110 8680 2113
rect 8695 2110 8708 2113
rect 8631 2106 8661 2107
rect 8670 2106 8676 2107
rect 8679 2106 8708 2110
rect 8598 2105 8708 2106
rect 8598 2104 8714 2105
rect 8273 2096 8324 2104
rect 8273 2084 8298 2096
rect 8305 2084 8324 2096
rect 8355 2096 8405 2104
rect 8355 2088 8371 2096
rect 8378 2094 8405 2096
rect 8414 2094 8635 2104
rect 8378 2084 8635 2094
rect 8664 2096 8714 2104
rect 8664 2087 8680 2096
rect 8273 2076 8324 2084
rect 8371 2076 8635 2084
rect 8661 2084 8680 2087
rect 8687 2084 8714 2096
rect 8661 2076 8714 2084
rect 8289 2068 8290 2076
rect 8305 2068 8318 2076
rect 8289 2060 8305 2068
rect 8286 2053 8305 2056
rect 8286 2044 8308 2053
rect 8259 2034 8308 2044
rect 8259 2028 8289 2034
rect 8308 2029 8313 2034
rect 8231 2012 8305 2028
rect 8323 2020 8353 2076
rect 8388 2066 8596 2076
rect 8631 2072 8676 2076
rect 8679 2075 8680 2076
rect 8695 2075 8708 2076
rect 8414 2036 8603 2066
rect 8429 2033 8603 2036
rect 8422 2030 8603 2033
rect 8231 2010 8244 2012
rect 8259 2010 8293 2012
rect 8231 1994 8305 2010
rect 8332 2006 8345 2020
rect 8360 2006 8376 2022
rect 8422 2017 8433 2030
rect 8215 1972 8216 1988
rect 8231 1972 8244 1994
rect 8259 1972 8289 1994
rect 8332 1990 8394 2006
rect 8422 1999 8433 2015
rect 8438 2010 8448 2030
rect 8458 2010 8472 2030
rect 8475 2017 8484 2030
rect 8500 2017 8509 2030
rect 8438 1999 8472 2010
rect 8475 1999 8484 2015
rect 8500 1999 8509 2015
rect 8516 2010 8526 2030
rect 8536 2010 8550 2030
rect 8551 2017 8562 2030
rect 8516 1999 8550 2010
rect 8551 1999 8562 2015
rect 8608 2006 8624 2022
rect 8631 2020 8661 2072
rect 8695 2068 8696 2075
rect 8680 2060 8696 2068
rect 8667 2028 8680 2047
rect 8695 2028 8725 2044
rect 8667 2012 8741 2028
rect 8667 2010 8680 2012
rect 8695 2010 8729 2012
rect 8332 1988 8345 1990
rect 8360 1988 8394 1990
rect 8332 1972 8394 1988
rect 8438 1983 8454 1986
rect 8516 1983 8546 1994
rect 8594 1990 8640 2006
rect 8667 1994 8741 2010
rect 8594 1988 8628 1990
rect 8593 1972 8640 1988
rect 8667 1972 8680 1994
rect 8695 1972 8725 1994
rect 8752 1972 8753 1988
rect 8768 1972 8781 2132
rect 8811 2028 8824 2132
rect 8869 2110 8870 2120
rect 8885 2110 8898 2120
rect 8869 2106 8898 2110
rect 8903 2106 8933 2132
rect 8951 2118 8967 2120
rect 9039 2118 9092 2132
rect 9040 2116 9104 2118
rect 9147 2116 9162 2132
rect 9211 2129 9241 2132
rect 9211 2126 9247 2129
rect 9177 2118 9193 2120
rect 8951 2106 8966 2110
rect 8869 2104 8966 2106
rect 8994 2104 9162 2116
rect 9178 2106 9193 2110
rect 9211 2107 9250 2126
rect 9269 2120 9276 2121
rect 9275 2113 9276 2120
rect 9259 2110 9260 2113
rect 9275 2110 9288 2113
rect 9211 2106 9241 2107
rect 9250 2106 9256 2107
rect 9259 2106 9288 2110
rect 9178 2105 9288 2106
rect 9178 2104 9294 2105
rect 8853 2096 8904 2104
rect 8853 2084 8878 2096
rect 8885 2084 8904 2096
rect 8935 2096 8985 2104
rect 8935 2088 8951 2096
rect 8958 2094 8985 2096
rect 8994 2094 9215 2104
rect 8958 2084 9215 2094
rect 9244 2096 9294 2104
rect 9244 2087 9260 2096
rect 8853 2076 8904 2084
rect 8951 2076 9215 2084
rect 9241 2084 9260 2087
rect 9267 2084 9294 2096
rect 9241 2076 9294 2084
rect 8869 2068 8870 2076
rect 8885 2068 8898 2076
rect 8869 2060 8885 2068
rect 8866 2053 8885 2056
rect 8866 2044 8888 2053
rect 8839 2034 8888 2044
rect 8839 2028 8869 2034
rect 8888 2029 8893 2034
rect 8811 2012 8885 2028
rect 8903 2020 8933 2076
rect 8968 2066 9176 2076
rect 9211 2072 9256 2076
rect 9259 2075 9260 2076
rect 9275 2075 9288 2076
rect 8994 2036 9183 2066
rect 9009 2033 9183 2036
rect 9002 2030 9183 2033
rect 8811 2010 8824 2012
rect 8839 2010 8873 2012
rect 8811 1994 8885 2010
rect 8912 2006 8925 2020
rect 8940 2006 8956 2022
rect 9002 2017 9013 2030
rect 8795 1972 8796 1988
rect 8811 1972 8824 1994
rect 8839 1972 8869 1994
rect 8912 1990 8974 2006
rect 9002 1999 9013 2015
rect 9018 2010 9028 2030
rect 9038 2010 9052 2030
rect 9055 2017 9064 2030
rect 9080 2017 9089 2030
rect 9018 1999 9052 2010
rect 9055 1999 9064 2015
rect 9080 1999 9089 2015
rect 9096 2010 9106 2030
rect 9116 2010 9130 2030
rect 9131 2017 9142 2030
rect 9096 1999 9130 2010
rect 9131 1999 9142 2015
rect 9188 2006 9204 2022
rect 9211 2020 9241 2072
rect 9275 2068 9276 2075
rect 9260 2060 9276 2068
rect 9247 2028 9260 2047
rect 9275 2028 9305 2044
rect 9247 2012 9321 2028
rect 9247 2010 9260 2012
rect 9275 2010 9309 2012
rect 8912 1988 8925 1990
rect 8940 1988 8974 1990
rect 8912 1972 8974 1988
rect 9018 1983 9034 1986
rect 9096 1983 9126 1994
rect 9174 1990 9220 2006
rect 9247 1994 9321 2010
rect 9174 1988 9208 1990
rect 9173 1972 9220 1988
rect 9247 1972 9260 1994
rect 9275 1972 9305 1994
rect 9332 1972 9333 1988
rect 9348 1972 9361 2132
rect -9 1964 32 1972
rect -9 1938 6 1964
rect 13 1938 32 1964
rect 96 1960 158 1972
rect 170 1960 245 1972
rect 303 1960 378 1972
rect 390 1960 421 1972
rect 427 1960 462 1972
rect 96 1958 258 1960
rect -9 1930 32 1938
rect 114 1934 127 1958
rect 142 1956 157 1958
rect -3 1920 -2 1930
rect 13 1920 26 1930
rect 41 1920 71 1934
rect 114 1920 157 1934
rect 181 1931 188 1938
rect 191 1934 258 1958
rect 290 1958 462 1960
rect 260 1936 288 1940
rect 290 1936 370 1958
rect 391 1956 406 1958
rect 260 1934 370 1936
rect 191 1930 370 1934
rect 164 1920 194 1930
rect 196 1920 349 1930
rect 357 1920 387 1930
rect 391 1920 421 1934
rect 449 1920 462 1958
rect 534 1964 569 1972
rect 534 1938 535 1964
rect 542 1938 569 1964
rect 477 1920 507 1934
rect 534 1930 569 1938
rect 571 1964 612 1972
rect 571 1938 586 1964
rect 593 1938 612 1964
rect 676 1960 738 1972
rect 750 1960 825 1972
rect 883 1960 958 1972
rect 970 1960 1001 1972
rect 1007 1960 1042 1972
rect 676 1958 838 1960
rect 571 1930 612 1938
rect 694 1934 707 1958
rect 722 1956 737 1958
rect 534 1920 535 1930
rect 550 1920 563 1930
rect 577 1920 578 1930
rect 593 1920 606 1930
rect 621 1920 651 1934
rect 694 1920 737 1934
rect 761 1931 768 1938
rect 771 1934 838 1958
rect 870 1958 1042 1960
rect 840 1936 868 1940
rect 870 1936 950 1958
rect 971 1956 986 1958
rect 840 1934 950 1936
rect 771 1930 950 1934
rect 744 1920 774 1930
rect 776 1920 929 1930
rect 937 1920 967 1930
rect 971 1920 1001 1934
rect 1029 1920 1042 1958
rect 1114 1964 1149 1972
rect 1114 1938 1115 1964
rect 1122 1938 1149 1964
rect 1057 1920 1087 1934
rect 1114 1930 1149 1938
rect 1151 1964 1192 1972
rect 1151 1938 1166 1964
rect 1173 1938 1192 1964
rect 1256 1960 1318 1972
rect 1330 1960 1405 1972
rect 1463 1960 1538 1972
rect 1550 1960 1581 1972
rect 1587 1960 1622 1972
rect 1256 1958 1418 1960
rect 1151 1930 1192 1938
rect 1274 1934 1287 1958
rect 1302 1956 1317 1958
rect 1114 1920 1115 1930
rect 1130 1920 1143 1930
rect 1157 1920 1158 1930
rect 1173 1920 1186 1930
rect 1201 1920 1231 1934
rect 1274 1920 1317 1934
rect 1341 1931 1348 1938
rect 1351 1934 1418 1958
rect 1450 1958 1622 1960
rect 1420 1936 1448 1940
rect 1450 1936 1530 1958
rect 1551 1956 1566 1958
rect 1420 1934 1530 1936
rect 1351 1930 1530 1934
rect 1324 1920 1354 1930
rect 1356 1920 1509 1930
rect 1517 1920 1547 1930
rect 1551 1920 1581 1934
rect 1609 1920 1622 1958
rect 1694 1964 1729 1972
rect 1694 1938 1695 1964
rect 1702 1938 1729 1964
rect 1637 1920 1667 1934
rect 1694 1930 1729 1938
rect 1731 1964 1772 1972
rect 1731 1938 1746 1964
rect 1753 1938 1772 1964
rect 1836 1960 1898 1972
rect 1910 1960 1985 1972
rect 2043 1960 2118 1972
rect 2130 1960 2161 1972
rect 2167 1960 2202 1972
rect 1836 1958 1998 1960
rect 1731 1930 1772 1938
rect 1854 1934 1867 1958
rect 1882 1956 1897 1958
rect 1694 1920 1695 1930
rect 1710 1920 1723 1930
rect 1737 1920 1738 1930
rect 1753 1920 1766 1930
rect 1781 1920 1811 1934
rect 1854 1920 1897 1934
rect 1921 1931 1928 1938
rect 1931 1934 1998 1958
rect 2030 1958 2202 1960
rect 2000 1936 2028 1940
rect 2030 1936 2110 1958
rect 2131 1956 2146 1958
rect 2000 1934 2110 1936
rect 1931 1930 2110 1934
rect 1904 1920 1934 1930
rect 1936 1920 2089 1930
rect 2097 1920 2127 1930
rect 2131 1920 2161 1934
rect 2189 1920 2202 1958
rect 2274 1964 2309 1972
rect 2274 1938 2275 1964
rect 2282 1938 2309 1964
rect 2217 1920 2247 1934
rect 2274 1930 2309 1938
rect 2311 1964 2352 1972
rect 2311 1938 2326 1964
rect 2333 1938 2352 1964
rect 2416 1960 2478 1972
rect 2490 1960 2565 1972
rect 2623 1960 2698 1972
rect 2710 1960 2741 1972
rect 2747 1960 2782 1972
rect 2416 1958 2578 1960
rect 2311 1930 2352 1938
rect 2434 1934 2447 1958
rect 2462 1956 2477 1958
rect 2274 1920 2275 1930
rect 2290 1920 2303 1930
rect 2317 1920 2318 1930
rect 2333 1920 2346 1930
rect 2361 1920 2391 1934
rect 2434 1920 2477 1934
rect 2501 1931 2508 1938
rect 2511 1934 2578 1958
rect 2610 1958 2782 1960
rect 2580 1936 2608 1940
rect 2610 1936 2690 1958
rect 2711 1956 2726 1958
rect 2580 1934 2690 1936
rect 2511 1930 2690 1934
rect 2484 1920 2514 1930
rect 2516 1920 2669 1930
rect 2677 1920 2707 1930
rect 2711 1920 2741 1934
rect 2769 1920 2782 1958
rect 2854 1964 2889 1972
rect 2854 1938 2855 1964
rect 2862 1938 2889 1964
rect 2797 1920 2827 1934
rect 2854 1930 2889 1938
rect 2891 1964 2932 1972
rect 2891 1938 2906 1964
rect 2913 1938 2932 1964
rect 2996 1960 3058 1972
rect 3070 1960 3145 1972
rect 3203 1960 3278 1972
rect 3290 1960 3321 1972
rect 3327 1960 3362 1972
rect 2996 1958 3158 1960
rect 2891 1930 2932 1938
rect 3014 1934 3027 1958
rect 3042 1956 3057 1958
rect 2854 1920 2855 1930
rect 2870 1920 2883 1930
rect 2897 1920 2898 1930
rect 2913 1920 2926 1930
rect 2941 1920 2971 1934
rect 3014 1920 3057 1934
rect 3081 1931 3088 1938
rect 3091 1934 3158 1958
rect 3190 1958 3362 1960
rect 3160 1936 3188 1940
rect 3190 1936 3270 1958
rect 3291 1956 3306 1958
rect 3160 1934 3270 1936
rect 3091 1930 3270 1934
rect 3064 1920 3094 1930
rect 3096 1920 3249 1930
rect 3257 1920 3287 1930
rect 3291 1920 3321 1934
rect 3349 1920 3362 1958
rect 3434 1964 3469 1972
rect 3434 1938 3435 1964
rect 3442 1938 3469 1964
rect 3377 1920 3407 1934
rect 3434 1930 3469 1938
rect 3434 1920 3435 1930
rect 3450 1920 3463 1930
rect -3 1914 3469 1920
rect -2 1906 3469 1914
rect 5889 1964 5930 1972
rect 5889 1938 5904 1964
rect 5911 1938 5930 1964
rect 5994 1960 6056 1972
rect 6068 1960 6143 1972
rect 6201 1960 6276 1972
rect 6288 1960 6319 1972
rect 6325 1960 6360 1972
rect 5994 1958 6156 1960
rect 5889 1930 5930 1938
rect 6012 1934 6025 1958
rect 6040 1956 6055 1958
rect 5895 1920 5896 1930
rect 5911 1920 5924 1930
rect 5939 1920 5969 1934
rect 6012 1920 6055 1934
rect 6079 1931 6086 1938
rect 6089 1934 6156 1958
rect 6188 1958 6360 1960
rect 6158 1936 6186 1940
rect 6188 1936 6268 1958
rect 6289 1956 6304 1958
rect 6158 1934 6268 1936
rect 6089 1930 6268 1934
rect 6062 1920 6092 1930
rect 6094 1920 6247 1930
rect 6255 1920 6285 1930
rect 6289 1920 6319 1934
rect 6347 1920 6360 1958
rect 6432 1964 6467 1972
rect 6432 1938 6433 1964
rect 6440 1938 6467 1964
rect 6375 1920 6405 1934
rect 6432 1930 6467 1938
rect 6469 1964 6510 1972
rect 6469 1938 6484 1964
rect 6491 1938 6510 1964
rect 6574 1960 6636 1972
rect 6648 1960 6723 1972
rect 6781 1960 6856 1972
rect 6868 1960 6899 1972
rect 6905 1960 6940 1972
rect 6574 1958 6736 1960
rect 6469 1930 6510 1938
rect 6592 1934 6605 1958
rect 6620 1956 6635 1958
rect 6432 1920 6433 1930
rect 6448 1920 6461 1930
rect 6475 1920 6476 1930
rect 6491 1920 6504 1930
rect 6519 1920 6549 1934
rect 6592 1920 6635 1934
rect 6659 1931 6666 1938
rect 6669 1934 6736 1958
rect 6768 1958 6940 1960
rect 6738 1936 6766 1940
rect 6768 1936 6848 1958
rect 6869 1956 6884 1958
rect 6738 1934 6848 1936
rect 6669 1930 6848 1934
rect 6642 1920 6672 1930
rect 6674 1920 6827 1930
rect 6835 1920 6865 1930
rect 6869 1920 6899 1934
rect 6927 1920 6940 1958
rect 7012 1964 7047 1972
rect 7012 1938 7013 1964
rect 7020 1938 7047 1964
rect 6955 1920 6985 1934
rect 7012 1930 7047 1938
rect 7049 1964 7090 1972
rect 7049 1938 7064 1964
rect 7071 1938 7090 1964
rect 7154 1960 7216 1972
rect 7228 1960 7303 1972
rect 7361 1960 7436 1972
rect 7448 1960 7479 1972
rect 7485 1960 7520 1972
rect 7154 1958 7316 1960
rect 7049 1930 7090 1938
rect 7172 1934 7185 1958
rect 7200 1956 7215 1958
rect 7012 1920 7013 1930
rect 7028 1920 7041 1930
rect 7055 1920 7056 1930
rect 7071 1920 7084 1930
rect 7099 1920 7129 1934
rect 7172 1920 7215 1934
rect 7239 1931 7246 1938
rect 7249 1934 7316 1958
rect 7348 1958 7520 1960
rect 7318 1936 7346 1940
rect 7348 1936 7428 1958
rect 7449 1956 7464 1958
rect 7318 1934 7428 1936
rect 7249 1930 7428 1934
rect 7222 1920 7252 1930
rect 7254 1920 7407 1930
rect 7415 1920 7445 1930
rect 7449 1920 7479 1934
rect 7507 1920 7520 1958
rect 7592 1964 7627 1972
rect 7592 1938 7593 1964
rect 7600 1938 7627 1964
rect 7535 1920 7565 1934
rect 7592 1930 7627 1938
rect 7629 1964 7670 1972
rect 7629 1938 7644 1964
rect 7651 1938 7670 1964
rect 7734 1960 7796 1972
rect 7808 1960 7883 1972
rect 7941 1960 8016 1972
rect 8028 1960 8059 1972
rect 8065 1960 8100 1972
rect 7734 1958 7896 1960
rect 7629 1930 7670 1938
rect 7752 1934 7765 1958
rect 7780 1956 7795 1958
rect 7592 1920 7593 1930
rect 7608 1920 7621 1930
rect 7635 1920 7636 1930
rect 7651 1920 7664 1930
rect 7679 1920 7709 1934
rect 7752 1920 7795 1934
rect 7819 1931 7826 1938
rect 7829 1934 7896 1958
rect 7928 1958 8100 1960
rect 7898 1936 7926 1940
rect 7928 1936 8008 1958
rect 8029 1956 8044 1958
rect 7898 1934 8008 1936
rect 7829 1930 8008 1934
rect 7802 1920 7832 1930
rect 7834 1920 7987 1930
rect 7995 1920 8025 1930
rect 8029 1920 8059 1934
rect 8087 1920 8100 1958
rect 8172 1964 8207 1972
rect 8172 1938 8173 1964
rect 8180 1938 8207 1964
rect 8115 1920 8145 1934
rect 8172 1930 8207 1938
rect 8209 1964 8250 1972
rect 8209 1938 8224 1964
rect 8231 1938 8250 1964
rect 8314 1960 8376 1972
rect 8388 1960 8463 1972
rect 8521 1960 8596 1972
rect 8608 1960 8639 1972
rect 8645 1960 8680 1972
rect 8314 1958 8476 1960
rect 8209 1930 8250 1938
rect 8332 1934 8345 1958
rect 8360 1956 8375 1958
rect 8172 1920 8173 1930
rect 8188 1920 8201 1930
rect 8215 1920 8216 1930
rect 8231 1920 8244 1930
rect 8259 1920 8289 1934
rect 8332 1920 8375 1934
rect 8399 1931 8406 1938
rect 8409 1934 8476 1958
rect 8508 1958 8680 1960
rect 8478 1936 8506 1940
rect 8508 1936 8588 1958
rect 8609 1956 8624 1958
rect 8478 1934 8588 1936
rect 8409 1930 8588 1934
rect 8382 1920 8412 1930
rect 8414 1920 8567 1930
rect 8575 1920 8605 1930
rect 8609 1920 8639 1934
rect 8667 1920 8680 1958
rect 8752 1964 8787 1972
rect 8752 1938 8753 1964
rect 8760 1938 8787 1964
rect 8695 1920 8725 1934
rect 8752 1930 8787 1938
rect 8789 1964 8830 1972
rect 8789 1938 8804 1964
rect 8811 1938 8830 1964
rect 8894 1960 8956 1972
rect 8968 1960 9043 1972
rect 9101 1960 9176 1972
rect 9188 1960 9219 1972
rect 9225 1960 9260 1972
rect 8894 1958 9056 1960
rect 8789 1930 8830 1938
rect 8912 1934 8925 1958
rect 8940 1956 8955 1958
rect 8752 1920 8753 1930
rect 8768 1920 8781 1930
rect 8795 1920 8796 1930
rect 8811 1920 8824 1930
rect 8839 1920 8869 1934
rect 8912 1920 8955 1934
rect 8979 1931 8986 1938
rect 8989 1934 9056 1958
rect 9088 1958 9260 1960
rect 9058 1936 9086 1940
rect 9088 1936 9168 1958
rect 9189 1956 9204 1958
rect 9058 1934 9168 1936
rect 8989 1930 9168 1934
rect 8962 1920 8992 1930
rect 8994 1920 9147 1930
rect 9155 1920 9185 1930
rect 9189 1920 9219 1934
rect 9247 1920 9260 1958
rect 9332 1964 9367 1972
rect 9332 1938 9333 1964
rect 9340 1938 9367 1964
rect 9275 1920 9305 1934
rect 9332 1930 9367 1938
rect 9332 1920 9333 1930
rect 9348 1920 9361 1930
rect 5889 1906 9361 1920
rect 13 1876 26 1906
rect 41 1888 71 1906
rect 114 1892 128 1906
rect 164 1892 384 1906
rect 115 1890 128 1892
rect 81 1878 96 1890
rect 78 1876 100 1878
rect 105 1876 135 1890
rect 196 1888 349 1892
rect 178 1876 370 1888
rect 413 1876 443 1890
rect 449 1876 462 1906
rect 477 1888 507 1906
rect 550 1876 563 1906
rect 593 1876 606 1906
rect 621 1888 651 1906
rect 694 1892 708 1906
rect 744 1892 964 1906
rect 695 1890 708 1892
rect 661 1878 676 1890
rect 658 1876 680 1878
rect 685 1876 715 1890
rect 776 1888 929 1892
rect 758 1876 950 1888
rect 993 1876 1023 1890
rect 1029 1876 1042 1906
rect 1057 1888 1087 1906
rect 1130 1876 1143 1906
rect 1173 1876 1186 1906
rect 1201 1888 1231 1906
rect 1274 1892 1288 1906
rect 1324 1892 1544 1906
rect 1275 1890 1288 1892
rect 1241 1878 1256 1890
rect 1238 1876 1260 1878
rect 1265 1876 1295 1890
rect 1356 1888 1509 1892
rect 1338 1876 1530 1888
rect 1573 1876 1603 1890
rect 1609 1876 1622 1906
rect 1637 1888 1667 1906
rect 1710 1876 1723 1906
rect 1753 1876 1766 1906
rect 1781 1888 1811 1906
rect 1854 1892 1868 1906
rect 1904 1892 2124 1906
rect 1855 1890 1868 1892
rect 1821 1878 1836 1890
rect 1818 1876 1840 1878
rect 1845 1876 1875 1890
rect 1936 1888 2089 1892
rect 1918 1876 2110 1888
rect 2153 1876 2183 1890
rect 2189 1876 2202 1906
rect 2217 1888 2247 1906
rect 2290 1876 2303 1906
rect 2333 1876 2346 1906
rect 2361 1888 2391 1906
rect 2434 1892 2448 1906
rect 2484 1892 2704 1906
rect 2435 1890 2448 1892
rect 2401 1878 2416 1890
rect 2398 1876 2420 1878
rect 2425 1876 2455 1890
rect 2516 1888 2669 1892
rect 2498 1876 2690 1888
rect 2733 1876 2763 1890
rect 2769 1876 2782 1906
rect 2797 1888 2827 1906
rect 2870 1876 2883 1906
rect 2913 1876 2926 1906
rect 2941 1888 2971 1906
rect 3014 1892 3028 1906
rect 3064 1892 3284 1906
rect 3015 1890 3028 1892
rect 2981 1878 2996 1890
rect 2978 1876 3000 1878
rect 3005 1876 3035 1890
rect 3096 1888 3249 1892
rect 3078 1876 3270 1888
rect 3313 1876 3343 1890
rect 3349 1876 3362 1906
rect 3377 1888 3407 1906
rect 3450 1876 3463 1906
rect 5911 1876 5924 1906
rect 5939 1888 5969 1906
rect 6012 1892 6026 1906
rect 6062 1892 6282 1906
rect 6013 1890 6026 1892
rect 5979 1878 5994 1890
rect 5976 1876 5998 1878
rect 6003 1876 6033 1890
rect 6094 1888 6247 1892
rect 6076 1876 6268 1888
rect 6311 1876 6341 1890
rect 6347 1876 6360 1906
rect 6375 1888 6405 1906
rect 6448 1876 6461 1906
rect 6491 1876 6504 1906
rect 6519 1888 6549 1906
rect 6592 1892 6606 1906
rect 6642 1892 6862 1906
rect 6593 1890 6606 1892
rect 6559 1878 6574 1890
rect 6556 1876 6578 1878
rect 6583 1876 6613 1890
rect 6674 1888 6827 1892
rect 6656 1876 6848 1888
rect 6891 1876 6921 1890
rect 6927 1876 6940 1906
rect 6955 1888 6985 1906
rect 7028 1876 7041 1906
rect 7071 1876 7084 1906
rect 7099 1888 7129 1906
rect 7172 1892 7186 1906
rect 7222 1892 7442 1906
rect 7173 1890 7186 1892
rect 7139 1878 7154 1890
rect 7136 1876 7158 1878
rect 7163 1876 7193 1890
rect 7254 1888 7407 1892
rect 7236 1876 7428 1888
rect 7471 1876 7501 1890
rect 7507 1876 7520 1906
rect 7535 1888 7565 1906
rect 7608 1876 7621 1906
rect 7651 1876 7664 1906
rect 7679 1888 7709 1906
rect 7752 1892 7766 1906
rect 7802 1892 8022 1906
rect 7753 1890 7766 1892
rect 7719 1878 7734 1890
rect 7716 1876 7738 1878
rect 7743 1876 7773 1890
rect 7834 1888 7987 1892
rect 7816 1876 8008 1888
rect 8051 1876 8081 1890
rect 8087 1876 8100 1906
rect 8115 1888 8145 1906
rect 8188 1876 8201 1906
rect 8231 1876 8244 1906
rect 8259 1888 8289 1906
rect 8332 1892 8346 1906
rect 8382 1892 8602 1906
rect 8333 1890 8346 1892
rect 8299 1878 8314 1890
rect 8296 1876 8318 1878
rect 8323 1876 8353 1890
rect 8414 1888 8567 1892
rect 8396 1876 8588 1888
rect 8631 1876 8661 1890
rect 8667 1876 8680 1906
rect 8695 1888 8725 1906
rect 8768 1876 8781 1906
rect 8811 1876 8824 1906
rect 8839 1888 8869 1906
rect 8912 1892 8926 1906
rect 8962 1892 9182 1906
rect 8913 1890 8926 1892
rect 8879 1878 8894 1890
rect 8876 1876 8898 1878
rect 8903 1876 8933 1890
rect 8994 1888 9147 1892
rect 8976 1876 9168 1888
rect 9211 1876 9241 1890
rect 9247 1876 9260 1906
rect 9275 1888 9305 1906
rect 9348 1876 9361 1906
rect -2 1862 3469 1876
rect 5889 1862 9361 1876
rect 13 1758 26 1862
rect 71 1840 72 1850
rect 87 1840 100 1850
rect 71 1836 100 1840
rect 105 1836 135 1862
rect 153 1848 169 1850
rect 241 1848 294 1862
rect 242 1846 306 1848
rect 349 1846 364 1862
rect 413 1859 443 1862
rect 413 1856 449 1859
rect 379 1848 395 1850
rect 153 1836 168 1840
rect 71 1834 168 1836
rect 196 1834 364 1846
rect 380 1836 395 1840
rect 413 1837 452 1856
rect 471 1850 478 1851
rect 477 1843 478 1850
rect 461 1840 462 1843
rect 477 1840 490 1843
rect 413 1836 443 1837
rect 452 1836 458 1837
rect 461 1836 490 1840
rect 380 1835 490 1836
rect 380 1834 496 1835
rect 55 1826 106 1834
rect 55 1814 80 1826
rect 87 1814 106 1826
rect 137 1826 187 1834
rect 137 1818 153 1826
rect 160 1824 187 1826
rect 196 1824 417 1834
rect 160 1814 417 1824
rect 446 1826 496 1834
rect 446 1817 462 1826
rect 55 1806 106 1814
rect 153 1806 417 1814
rect 443 1814 462 1817
rect 469 1814 496 1826
rect 443 1806 496 1814
rect 71 1798 72 1806
rect 87 1798 100 1806
rect 71 1790 87 1798
rect 68 1783 87 1786
rect 68 1774 90 1783
rect 41 1764 90 1774
rect 41 1758 71 1764
rect 90 1759 95 1764
rect 13 1742 87 1758
rect 105 1750 135 1806
rect 170 1796 378 1806
rect 413 1802 458 1806
rect 461 1805 462 1806
rect 477 1805 490 1806
rect 196 1766 385 1796
rect 211 1763 385 1766
rect 204 1760 385 1763
rect 13 1740 26 1742
rect 41 1740 75 1742
rect 13 1724 87 1740
rect 114 1736 127 1750
rect 142 1736 158 1752
rect 204 1747 215 1760
rect -3 1702 -2 1718
rect 13 1702 26 1724
rect 41 1702 71 1724
rect 114 1720 176 1736
rect 204 1729 215 1745
rect 220 1740 230 1760
rect 240 1740 254 1760
rect 257 1747 266 1760
rect 282 1747 291 1760
rect 220 1729 254 1740
rect 257 1729 266 1745
rect 282 1729 291 1745
rect 298 1740 308 1760
rect 318 1740 332 1760
rect 333 1747 344 1760
rect 298 1729 332 1740
rect 333 1729 344 1745
rect 390 1736 406 1752
rect 413 1750 443 1802
rect 477 1798 478 1805
rect 462 1790 478 1798
rect 449 1758 462 1777
rect 477 1758 507 1774
rect 449 1742 523 1758
rect 449 1740 462 1742
rect 477 1740 511 1742
rect 114 1718 127 1720
rect 142 1718 176 1720
rect 114 1702 176 1718
rect 220 1713 236 1716
rect 298 1713 328 1724
rect 376 1720 422 1736
rect 449 1724 523 1740
rect 376 1718 410 1720
rect 375 1702 422 1718
rect 449 1702 462 1724
rect 477 1702 507 1724
rect 534 1702 535 1718
rect 550 1702 563 1862
rect 593 1758 606 1862
rect 651 1840 652 1850
rect 667 1840 680 1850
rect 651 1836 680 1840
rect 685 1836 715 1862
rect 733 1848 749 1850
rect 821 1848 874 1862
rect 822 1846 886 1848
rect 929 1846 944 1862
rect 993 1859 1023 1862
rect 993 1856 1029 1859
rect 959 1848 975 1850
rect 733 1836 748 1840
rect 651 1834 748 1836
rect 776 1834 944 1846
rect 960 1836 975 1840
rect 993 1837 1032 1856
rect 1051 1850 1058 1851
rect 1057 1843 1058 1850
rect 1041 1840 1042 1843
rect 1057 1840 1070 1843
rect 993 1836 1023 1837
rect 1032 1836 1038 1837
rect 1041 1836 1070 1840
rect 960 1835 1070 1836
rect 960 1834 1076 1835
rect 635 1826 686 1834
rect 635 1814 660 1826
rect 667 1814 686 1826
rect 717 1826 767 1834
rect 717 1818 733 1826
rect 740 1824 767 1826
rect 776 1824 997 1834
rect 740 1814 997 1824
rect 1026 1826 1076 1834
rect 1026 1817 1042 1826
rect 635 1806 686 1814
rect 733 1806 997 1814
rect 1023 1814 1042 1817
rect 1049 1814 1076 1826
rect 1023 1806 1076 1814
rect 651 1798 652 1806
rect 667 1798 680 1806
rect 651 1790 667 1798
rect 648 1783 667 1786
rect 648 1774 670 1783
rect 621 1764 670 1774
rect 621 1758 651 1764
rect 670 1759 675 1764
rect 593 1742 667 1758
rect 685 1750 715 1806
rect 750 1796 958 1806
rect 993 1802 1038 1806
rect 1041 1805 1042 1806
rect 1057 1805 1070 1806
rect 776 1766 965 1796
rect 791 1763 965 1766
rect 784 1760 965 1763
rect 593 1740 606 1742
rect 621 1740 655 1742
rect 593 1724 667 1740
rect 694 1736 707 1750
rect 722 1736 738 1752
rect 784 1747 795 1760
rect 577 1702 578 1718
rect 593 1702 606 1724
rect 621 1702 651 1724
rect 694 1720 756 1736
rect 784 1729 795 1745
rect 800 1740 810 1760
rect 820 1740 834 1760
rect 837 1747 846 1760
rect 862 1747 871 1760
rect 800 1729 834 1740
rect 837 1729 846 1745
rect 862 1729 871 1745
rect 878 1740 888 1760
rect 898 1740 912 1760
rect 913 1747 924 1760
rect 878 1729 912 1740
rect 913 1729 924 1745
rect 970 1736 986 1752
rect 993 1750 1023 1802
rect 1057 1798 1058 1805
rect 1042 1790 1058 1798
rect 1029 1758 1042 1777
rect 1057 1758 1087 1774
rect 1029 1742 1103 1758
rect 1029 1740 1042 1742
rect 1057 1740 1091 1742
rect 694 1718 707 1720
rect 722 1718 756 1720
rect 694 1702 756 1718
rect 800 1713 816 1716
rect 878 1713 908 1724
rect 956 1720 1002 1736
rect 1029 1724 1103 1740
rect 956 1718 990 1720
rect 955 1702 1002 1718
rect 1029 1702 1042 1724
rect 1057 1702 1087 1724
rect 1114 1702 1115 1718
rect 1130 1702 1143 1862
rect 1173 1758 1186 1862
rect 1231 1840 1232 1850
rect 1247 1840 1260 1850
rect 1231 1836 1260 1840
rect 1265 1836 1295 1862
rect 1313 1848 1329 1850
rect 1401 1848 1454 1862
rect 1402 1846 1466 1848
rect 1509 1846 1524 1862
rect 1573 1859 1603 1862
rect 1573 1856 1609 1859
rect 1539 1848 1555 1850
rect 1313 1836 1328 1840
rect 1231 1834 1328 1836
rect 1356 1834 1524 1846
rect 1540 1836 1555 1840
rect 1573 1837 1612 1856
rect 1631 1850 1638 1851
rect 1637 1843 1638 1850
rect 1621 1840 1622 1843
rect 1637 1840 1650 1843
rect 1573 1836 1603 1837
rect 1612 1836 1618 1837
rect 1621 1836 1650 1840
rect 1540 1835 1650 1836
rect 1540 1834 1656 1835
rect 1215 1826 1266 1834
rect 1215 1814 1240 1826
rect 1247 1814 1266 1826
rect 1297 1826 1347 1834
rect 1297 1818 1313 1826
rect 1320 1824 1347 1826
rect 1356 1824 1577 1834
rect 1320 1814 1577 1824
rect 1606 1826 1656 1834
rect 1606 1817 1622 1826
rect 1215 1806 1266 1814
rect 1313 1806 1577 1814
rect 1603 1814 1622 1817
rect 1629 1814 1656 1826
rect 1603 1806 1656 1814
rect 1231 1798 1232 1806
rect 1247 1798 1260 1806
rect 1231 1790 1247 1798
rect 1228 1783 1247 1786
rect 1228 1774 1250 1783
rect 1201 1764 1250 1774
rect 1201 1758 1231 1764
rect 1250 1759 1255 1764
rect 1173 1742 1247 1758
rect 1265 1750 1295 1806
rect 1330 1796 1538 1806
rect 1573 1802 1618 1806
rect 1621 1805 1622 1806
rect 1637 1805 1650 1806
rect 1356 1766 1545 1796
rect 1371 1763 1545 1766
rect 1364 1760 1545 1763
rect 1173 1740 1186 1742
rect 1201 1740 1235 1742
rect 1173 1724 1247 1740
rect 1274 1736 1287 1750
rect 1302 1736 1318 1752
rect 1364 1747 1375 1760
rect 1157 1702 1158 1718
rect 1173 1702 1186 1724
rect 1201 1702 1231 1724
rect 1274 1720 1336 1736
rect 1364 1729 1375 1745
rect 1380 1740 1390 1760
rect 1400 1740 1414 1760
rect 1417 1747 1426 1760
rect 1442 1747 1451 1760
rect 1380 1729 1414 1740
rect 1417 1729 1426 1745
rect 1442 1729 1451 1745
rect 1458 1740 1468 1760
rect 1478 1740 1492 1760
rect 1493 1747 1504 1760
rect 1458 1729 1492 1740
rect 1493 1729 1504 1745
rect 1550 1736 1566 1752
rect 1573 1750 1603 1802
rect 1637 1798 1638 1805
rect 1622 1790 1638 1798
rect 1609 1758 1622 1777
rect 1637 1758 1667 1774
rect 1609 1742 1683 1758
rect 1609 1740 1622 1742
rect 1637 1740 1671 1742
rect 1274 1718 1287 1720
rect 1302 1718 1336 1720
rect 1274 1702 1336 1718
rect 1380 1713 1396 1716
rect 1458 1713 1488 1724
rect 1536 1720 1582 1736
rect 1609 1724 1683 1740
rect 1536 1718 1570 1720
rect 1535 1702 1582 1718
rect 1609 1702 1622 1724
rect 1637 1702 1667 1724
rect 1694 1702 1695 1718
rect 1710 1702 1723 1862
rect 1753 1758 1766 1862
rect 1811 1840 1812 1850
rect 1827 1840 1840 1850
rect 1811 1836 1840 1840
rect 1845 1836 1875 1862
rect 1893 1848 1909 1850
rect 1981 1848 2034 1862
rect 1982 1846 2046 1848
rect 2089 1846 2104 1862
rect 2153 1859 2183 1862
rect 2153 1856 2189 1859
rect 2119 1848 2135 1850
rect 1893 1836 1908 1840
rect 1811 1834 1908 1836
rect 1936 1834 2104 1846
rect 2120 1836 2135 1840
rect 2153 1837 2192 1856
rect 2211 1850 2218 1851
rect 2217 1843 2218 1850
rect 2201 1840 2202 1843
rect 2217 1840 2230 1843
rect 2153 1836 2183 1837
rect 2192 1836 2198 1837
rect 2201 1836 2230 1840
rect 2120 1835 2230 1836
rect 2120 1834 2236 1835
rect 1795 1826 1846 1834
rect 1795 1814 1820 1826
rect 1827 1814 1846 1826
rect 1877 1826 1927 1834
rect 1877 1818 1893 1826
rect 1900 1824 1927 1826
rect 1936 1824 2157 1834
rect 1900 1814 2157 1824
rect 2186 1826 2236 1834
rect 2186 1817 2202 1826
rect 1795 1806 1846 1814
rect 1893 1806 2157 1814
rect 2183 1814 2202 1817
rect 2209 1814 2236 1826
rect 2183 1806 2236 1814
rect 1811 1798 1812 1806
rect 1827 1798 1840 1806
rect 1811 1790 1827 1798
rect 1808 1783 1827 1786
rect 1808 1774 1830 1783
rect 1781 1764 1830 1774
rect 1781 1758 1811 1764
rect 1830 1759 1835 1764
rect 1753 1742 1827 1758
rect 1845 1750 1875 1806
rect 1910 1796 2118 1806
rect 2153 1802 2198 1806
rect 2201 1805 2202 1806
rect 2217 1805 2230 1806
rect 1936 1766 2125 1796
rect 1951 1763 2125 1766
rect 1944 1760 2125 1763
rect 1753 1740 1766 1742
rect 1781 1740 1815 1742
rect 1753 1724 1827 1740
rect 1854 1736 1867 1750
rect 1882 1736 1898 1752
rect 1944 1747 1955 1760
rect 1737 1702 1738 1718
rect 1753 1702 1766 1724
rect 1781 1702 1811 1724
rect 1854 1720 1916 1736
rect 1944 1729 1955 1745
rect 1960 1740 1970 1760
rect 1980 1740 1994 1760
rect 1997 1747 2006 1760
rect 2022 1747 2031 1760
rect 1960 1729 1994 1740
rect 1997 1729 2006 1745
rect 2022 1729 2031 1745
rect 2038 1740 2048 1760
rect 2058 1740 2072 1760
rect 2073 1747 2084 1760
rect 2038 1729 2072 1740
rect 2073 1729 2084 1745
rect 2130 1736 2146 1752
rect 2153 1750 2183 1802
rect 2217 1798 2218 1805
rect 2202 1790 2218 1798
rect 2189 1758 2202 1777
rect 2217 1758 2247 1774
rect 2189 1742 2263 1758
rect 2189 1740 2202 1742
rect 2217 1740 2251 1742
rect 1854 1718 1867 1720
rect 1882 1718 1916 1720
rect 1854 1702 1916 1718
rect 1960 1713 1976 1716
rect 2038 1713 2068 1724
rect 2116 1720 2162 1736
rect 2189 1724 2263 1740
rect 2116 1718 2150 1720
rect 2115 1702 2162 1718
rect 2189 1702 2202 1724
rect 2217 1702 2247 1724
rect 2274 1702 2275 1718
rect 2290 1702 2303 1862
rect 2333 1758 2346 1862
rect 2391 1840 2392 1850
rect 2407 1840 2420 1850
rect 2391 1836 2420 1840
rect 2425 1836 2455 1862
rect 2473 1848 2489 1850
rect 2561 1848 2614 1862
rect 2562 1846 2626 1848
rect 2669 1846 2684 1862
rect 2733 1859 2763 1862
rect 2733 1856 2769 1859
rect 2699 1848 2715 1850
rect 2473 1836 2488 1840
rect 2391 1834 2488 1836
rect 2516 1834 2684 1846
rect 2700 1836 2715 1840
rect 2733 1837 2772 1856
rect 2791 1850 2798 1851
rect 2797 1843 2798 1850
rect 2781 1840 2782 1843
rect 2797 1840 2810 1843
rect 2733 1836 2763 1837
rect 2772 1836 2778 1837
rect 2781 1836 2810 1840
rect 2700 1835 2810 1836
rect 2700 1834 2816 1835
rect 2375 1826 2426 1834
rect 2375 1814 2400 1826
rect 2407 1814 2426 1826
rect 2457 1826 2507 1834
rect 2457 1818 2473 1826
rect 2480 1824 2507 1826
rect 2516 1824 2737 1834
rect 2480 1814 2737 1824
rect 2766 1826 2816 1834
rect 2766 1817 2782 1826
rect 2375 1806 2426 1814
rect 2473 1806 2737 1814
rect 2763 1814 2782 1817
rect 2789 1814 2816 1826
rect 2763 1806 2816 1814
rect 2391 1798 2392 1806
rect 2407 1798 2420 1806
rect 2391 1790 2407 1798
rect 2388 1783 2407 1786
rect 2388 1774 2410 1783
rect 2361 1764 2410 1774
rect 2361 1758 2391 1764
rect 2410 1759 2415 1764
rect 2333 1742 2407 1758
rect 2425 1750 2455 1806
rect 2490 1796 2698 1806
rect 2733 1802 2778 1806
rect 2781 1805 2782 1806
rect 2797 1805 2810 1806
rect 2516 1766 2705 1796
rect 2531 1763 2705 1766
rect 2524 1760 2705 1763
rect 2333 1740 2346 1742
rect 2361 1740 2395 1742
rect 2333 1724 2407 1740
rect 2434 1736 2447 1750
rect 2462 1736 2478 1752
rect 2524 1747 2535 1760
rect 2317 1702 2318 1718
rect 2333 1702 2346 1724
rect 2361 1702 2391 1724
rect 2434 1720 2496 1736
rect 2524 1729 2535 1745
rect 2540 1740 2550 1760
rect 2560 1740 2574 1760
rect 2577 1747 2586 1760
rect 2602 1747 2611 1760
rect 2540 1729 2574 1740
rect 2577 1729 2586 1745
rect 2602 1729 2611 1745
rect 2618 1740 2628 1760
rect 2638 1740 2652 1760
rect 2653 1747 2664 1760
rect 2618 1729 2652 1740
rect 2653 1729 2664 1745
rect 2710 1736 2726 1752
rect 2733 1750 2763 1802
rect 2797 1798 2798 1805
rect 2782 1790 2798 1798
rect 2769 1758 2782 1777
rect 2797 1758 2827 1774
rect 2769 1742 2843 1758
rect 2769 1740 2782 1742
rect 2797 1740 2831 1742
rect 2434 1718 2447 1720
rect 2462 1718 2496 1720
rect 2434 1702 2496 1718
rect 2540 1713 2556 1716
rect 2618 1713 2648 1724
rect 2696 1720 2742 1736
rect 2769 1724 2843 1740
rect 2696 1718 2730 1720
rect 2695 1702 2742 1718
rect 2769 1702 2782 1724
rect 2797 1702 2827 1724
rect 2854 1702 2855 1718
rect 2870 1702 2883 1862
rect 2913 1758 2926 1862
rect 2971 1840 2972 1850
rect 2987 1840 3000 1850
rect 2971 1836 3000 1840
rect 3005 1836 3035 1862
rect 3053 1848 3069 1850
rect 3141 1848 3194 1862
rect 3142 1846 3206 1848
rect 3249 1846 3264 1862
rect 3313 1859 3343 1862
rect 3313 1856 3349 1859
rect 3279 1848 3295 1850
rect 3053 1836 3068 1840
rect 2971 1834 3068 1836
rect 3096 1834 3264 1846
rect 3280 1836 3295 1840
rect 3313 1837 3352 1856
rect 3371 1850 3378 1851
rect 3377 1843 3378 1850
rect 3361 1840 3362 1843
rect 3377 1840 3390 1843
rect 3313 1836 3343 1837
rect 3352 1836 3358 1837
rect 3361 1836 3390 1840
rect 3280 1835 3390 1836
rect 3280 1834 3396 1835
rect 2955 1826 3006 1834
rect 2955 1814 2980 1826
rect 2987 1814 3006 1826
rect 3037 1826 3087 1834
rect 3037 1818 3053 1826
rect 3060 1824 3087 1826
rect 3096 1824 3317 1834
rect 3060 1814 3317 1824
rect 3346 1826 3396 1834
rect 3346 1817 3362 1826
rect 2955 1806 3006 1814
rect 3053 1806 3317 1814
rect 3343 1814 3362 1817
rect 3369 1814 3396 1826
rect 3343 1806 3396 1814
rect 2971 1798 2972 1806
rect 2987 1798 3000 1806
rect 2971 1790 2987 1798
rect 2968 1783 2987 1786
rect 2968 1774 2990 1783
rect 2941 1764 2990 1774
rect 2941 1758 2971 1764
rect 2990 1759 2995 1764
rect 2913 1742 2987 1758
rect 3005 1750 3035 1806
rect 3070 1796 3278 1806
rect 3313 1802 3358 1806
rect 3361 1805 3362 1806
rect 3377 1805 3390 1806
rect 3096 1766 3285 1796
rect 3111 1763 3285 1766
rect 3104 1760 3285 1763
rect 2913 1740 2926 1742
rect 2941 1740 2975 1742
rect 2913 1724 2987 1740
rect 3014 1736 3027 1750
rect 3042 1736 3058 1752
rect 3104 1747 3115 1760
rect 2897 1702 2898 1718
rect 2913 1702 2926 1724
rect 2941 1702 2971 1724
rect 3014 1720 3076 1736
rect 3104 1729 3115 1745
rect 3120 1740 3130 1760
rect 3140 1740 3154 1760
rect 3157 1747 3166 1760
rect 3182 1747 3191 1760
rect 3120 1729 3154 1740
rect 3157 1729 3166 1745
rect 3182 1729 3191 1745
rect 3198 1740 3208 1760
rect 3218 1740 3232 1760
rect 3233 1747 3244 1760
rect 3198 1729 3232 1740
rect 3233 1729 3244 1745
rect 3290 1736 3306 1752
rect 3313 1750 3343 1802
rect 3377 1798 3378 1805
rect 3362 1790 3378 1798
rect 3349 1758 3362 1777
rect 3377 1758 3407 1774
rect 3349 1742 3423 1758
rect 3349 1740 3362 1742
rect 3377 1740 3411 1742
rect 3014 1718 3027 1720
rect 3042 1718 3076 1720
rect 3014 1702 3076 1718
rect 3120 1713 3136 1716
rect 3198 1713 3228 1724
rect 3276 1720 3322 1736
rect 3349 1724 3423 1740
rect 3276 1718 3310 1720
rect 3275 1702 3322 1718
rect 3349 1702 3362 1724
rect 3377 1702 3407 1724
rect 3434 1702 3435 1718
rect 3450 1702 3463 1862
rect 5911 1758 5924 1862
rect 5969 1840 5970 1850
rect 5985 1840 5998 1850
rect 5969 1836 5998 1840
rect 6003 1836 6033 1862
rect 6051 1848 6067 1850
rect 6139 1848 6192 1862
rect 6140 1846 6204 1848
rect 6247 1846 6262 1862
rect 6311 1859 6341 1862
rect 6311 1856 6347 1859
rect 6277 1848 6293 1850
rect 6051 1836 6066 1840
rect 5969 1834 6066 1836
rect 6094 1834 6262 1846
rect 6278 1836 6293 1840
rect 6311 1837 6350 1856
rect 6369 1850 6376 1851
rect 6375 1843 6376 1850
rect 6359 1840 6360 1843
rect 6375 1840 6388 1843
rect 6311 1836 6341 1837
rect 6350 1836 6356 1837
rect 6359 1836 6388 1840
rect 6278 1835 6388 1836
rect 6278 1834 6394 1835
rect 5953 1826 6004 1834
rect 5953 1814 5978 1826
rect 5985 1814 6004 1826
rect 6035 1826 6085 1834
rect 6035 1818 6051 1826
rect 6058 1824 6085 1826
rect 6094 1824 6315 1834
rect 6058 1814 6315 1824
rect 6344 1826 6394 1834
rect 6344 1817 6360 1826
rect 5953 1806 6004 1814
rect 6051 1806 6315 1814
rect 6341 1814 6360 1817
rect 6367 1814 6394 1826
rect 6341 1806 6394 1814
rect 5969 1798 5970 1806
rect 5985 1798 5998 1806
rect 5969 1790 5985 1798
rect 5966 1783 5985 1786
rect 5966 1774 5988 1783
rect 5939 1764 5988 1774
rect 5939 1758 5969 1764
rect 5988 1759 5993 1764
rect 5911 1742 5985 1758
rect 6003 1750 6033 1806
rect 6068 1796 6276 1806
rect 6311 1802 6356 1806
rect 6359 1805 6360 1806
rect 6375 1805 6388 1806
rect 6094 1766 6283 1796
rect 6109 1763 6283 1766
rect 6102 1760 6283 1763
rect 5911 1740 5924 1742
rect 5939 1740 5973 1742
rect 5911 1724 5985 1740
rect 6012 1736 6025 1750
rect 6040 1736 6056 1752
rect 6102 1747 6113 1760
rect 5895 1702 5896 1718
rect 5911 1702 5924 1724
rect 5939 1702 5969 1724
rect 6012 1720 6074 1736
rect 6102 1729 6113 1745
rect 6118 1740 6128 1760
rect 6138 1740 6152 1760
rect 6155 1747 6164 1760
rect 6180 1747 6189 1760
rect 6118 1729 6152 1740
rect 6155 1729 6164 1745
rect 6180 1729 6189 1745
rect 6196 1740 6206 1760
rect 6216 1740 6230 1760
rect 6231 1747 6242 1760
rect 6196 1729 6230 1740
rect 6231 1729 6242 1745
rect 6288 1736 6304 1752
rect 6311 1750 6341 1802
rect 6375 1798 6376 1805
rect 6360 1790 6376 1798
rect 6347 1758 6360 1777
rect 6375 1758 6405 1774
rect 6347 1742 6421 1758
rect 6347 1740 6360 1742
rect 6375 1740 6409 1742
rect 6012 1718 6025 1720
rect 6040 1718 6074 1720
rect 6012 1702 6074 1718
rect 6118 1713 6134 1716
rect 6196 1713 6226 1724
rect 6274 1720 6320 1736
rect 6347 1724 6421 1740
rect 6274 1718 6308 1720
rect 6273 1702 6320 1718
rect 6347 1702 6360 1724
rect 6375 1702 6405 1724
rect 6432 1702 6433 1718
rect 6448 1702 6461 1862
rect 6491 1758 6504 1862
rect 6549 1840 6550 1850
rect 6565 1840 6578 1850
rect 6549 1836 6578 1840
rect 6583 1836 6613 1862
rect 6631 1848 6647 1850
rect 6719 1848 6772 1862
rect 6720 1846 6784 1848
rect 6827 1846 6842 1862
rect 6891 1859 6921 1862
rect 6891 1856 6927 1859
rect 6857 1848 6873 1850
rect 6631 1836 6646 1840
rect 6549 1834 6646 1836
rect 6674 1834 6842 1846
rect 6858 1836 6873 1840
rect 6891 1837 6930 1856
rect 6949 1850 6956 1851
rect 6955 1843 6956 1850
rect 6939 1840 6940 1843
rect 6955 1840 6968 1843
rect 6891 1836 6921 1837
rect 6930 1836 6936 1837
rect 6939 1836 6968 1840
rect 6858 1835 6968 1836
rect 6858 1834 6974 1835
rect 6533 1826 6584 1834
rect 6533 1814 6558 1826
rect 6565 1814 6584 1826
rect 6615 1826 6665 1834
rect 6615 1818 6631 1826
rect 6638 1824 6665 1826
rect 6674 1824 6895 1834
rect 6638 1814 6895 1824
rect 6924 1826 6974 1834
rect 6924 1817 6940 1826
rect 6533 1806 6584 1814
rect 6631 1806 6895 1814
rect 6921 1814 6940 1817
rect 6947 1814 6974 1826
rect 6921 1806 6974 1814
rect 6549 1798 6550 1806
rect 6565 1798 6578 1806
rect 6549 1790 6565 1798
rect 6546 1783 6565 1786
rect 6546 1774 6568 1783
rect 6519 1764 6568 1774
rect 6519 1758 6549 1764
rect 6568 1759 6573 1764
rect 6491 1742 6565 1758
rect 6583 1750 6613 1806
rect 6648 1796 6856 1806
rect 6891 1802 6936 1806
rect 6939 1805 6940 1806
rect 6955 1805 6968 1806
rect 6674 1766 6863 1796
rect 6689 1763 6863 1766
rect 6682 1760 6863 1763
rect 6491 1740 6504 1742
rect 6519 1740 6553 1742
rect 6491 1724 6565 1740
rect 6592 1736 6605 1750
rect 6620 1736 6636 1752
rect 6682 1747 6693 1760
rect 6475 1702 6476 1718
rect 6491 1702 6504 1724
rect 6519 1702 6549 1724
rect 6592 1720 6654 1736
rect 6682 1729 6693 1745
rect 6698 1740 6708 1760
rect 6718 1740 6732 1760
rect 6735 1747 6744 1760
rect 6760 1747 6769 1760
rect 6698 1729 6732 1740
rect 6735 1729 6744 1745
rect 6760 1729 6769 1745
rect 6776 1740 6786 1760
rect 6796 1740 6810 1760
rect 6811 1747 6822 1760
rect 6776 1729 6810 1740
rect 6811 1729 6822 1745
rect 6868 1736 6884 1752
rect 6891 1750 6921 1802
rect 6955 1798 6956 1805
rect 6940 1790 6956 1798
rect 6927 1758 6940 1777
rect 6955 1758 6985 1774
rect 6927 1742 7001 1758
rect 6927 1740 6940 1742
rect 6955 1740 6989 1742
rect 6592 1718 6605 1720
rect 6620 1718 6654 1720
rect 6592 1702 6654 1718
rect 6698 1713 6714 1716
rect 6776 1713 6806 1724
rect 6854 1720 6900 1736
rect 6927 1724 7001 1740
rect 6854 1718 6888 1720
rect 6853 1702 6900 1718
rect 6927 1702 6940 1724
rect 6955 1702 6985 1724
rect 7012 1702 7013 1718
rect 7028 1702 7041 1862
rect 7071 1758 7084 1862
rect 7129 1840 7130 1850
rect 7145 1840 7158 1850
rect 7129 1836 7158 1840
rect 7163 1836 7193 1862
rect 7211 1848 7227 1850
rect 7299 1848 7352 1862
rect 7300 1846 7364 1848
rect 7407 1846 7422 1862
rect 7471 1859 7501 1862
rect 7471 1856 7507 1859
rect 7437 1848 7453 1850
rect 7211 1836 7226 1840
rect 7129 1834 7226 1836
rect 7254 1834 7422 1846
rect 7438 1836 7453 1840
rect 7471 1837 7510 1856
rect 7529 1850 7536 1851
rect 7535 1843 7536 1850
rect 7519 1840 7520 1843
rect 7535 1840 7548 1843
rect 7471 1836 7501 1837
rect 7510 1836 7516 1837
rect 7519 1836 7548 1840
rect 7438 1835 7548 1836
rect 7438 1834 7554 1835
rect 7113 1826 7164 1834
rect 7113 1814 7138 1826
rect 7145 1814 7164 1826
rect 7195 1826 7245 1834
rect 7195 1818 7211 1826
rect 7218 1824 7245 1826
rect 7254 1824 7475 1834
rect 7218 1814 7475 1824
rect 7504 1826 7554 1834
rect 7504 1817 7520 1826
rect 7113 1806 7164 1814
rect 7211 1806 7475 1814
rect 7501 1814 7520 1817
rect 7527 1814 7554 1826
rect 7501 1806 7554 1814
rect 7129 1798 7130 1806
rect 7145 1798 7158 1806
rect 7129 1790 7145 1798
rect 7126 1783 7145 1786
rect 7126 1774 7148 1783
rect 7099 1764 7148 1774
rect 7099 1758 7129 1764
rect 7148 1759 7153 1764
rect 7071 1742 7145 1758
rect 7163 1750 7193 1806
rect 7228 1796 7436 1806
rect 7471 1802 7516 1806
rect 7519 1805 7520 1806
rect 7535 1805 7548 1806
rect 7254 1766 7443 1796
rect 7269 1763 7443 1766
rect 7262 1760 7443 1763
rect 7071 1740 7084 1742
rect 7099 1740 7133 1742
rect 7071 1724 7145 1740
rect 7172 1736 7185 1750
rect 7200 1736 7216 1752
rect 7262 1747 7273 1760
rect 7055 1702 7056 1718
rect 7071 1702 7084 1724
rect 7099 1702 7129 1724
rect 7172 1720 7234 1736
rect 7262 1729 7273 1745
rect 7278 1740 7288 1760
rect 7298 1740 7312 1760
rect 7315 1747 7324 1760
rect 7340 1747 7349 1760
rect 7278 1729 7312 1740
rect 7315 1729 7324 1745
rect 7340 1729 7349 1745
rect 7356 1740 7366 1760
rect 7376 1740 7390 1760
rect 7391 1747 7402 1760
rect 7356 1729 7390 1740
rect 7391 1729 7402 1745
rect 7448 1736 7464 1752
rect 7471 1750 7501 1802
rect 7535 1798 7536 1805
rect 7520 1790 7536 1798
rect 7507 1758 7520 1777
rect 7535 1758 7565 1774
rect 7507 1742 7581 1758
rect 7507 1740 7520 1742
rect 7535 1740 7569 1742
rect 7172 1718 7185 1720
rect 7200 1718 7234 1720
rect 7172 1702 7234 1718
rect 7278 1713 7294 1716
rect 7356 1713 7386 1724
rect 7434 1720 7480 1736
rect 7507 1724 7581 1740
rect 7434 1718 7468 1720
rect 7433 1702 7480 1718
rect 7507 1702 7520 1724
rect 7535 1702 7565 1724
rect 7592 1702 7593 1718
rect 7608 1702 7621 1862
rect 7651 1758 7664 1862
rect 7709 1840 7710 1850
rect 7725 1840 7738 1850
rect 7709 1836 7738 1840
rect 7743 1836 7773 1862
rect 7791 1848 7807 1850
rect 7879 1848 7932 1862
rect 7880 1846 7944 1848
rect 7987 1846 8002 1862
rect 8051 1859 8081 1862
rect 8051 1856 8087 1859
rect 8017 1848 8033 1850
rect 7791 1836 7806 1840
rect 7709 1834 7806 1836
rect 7834 1834 8002 1846
rect 8018 1836 8033 1840
rect 8051 1837 8090 1856
rect 8109 1850 8116 1851
rect 8115 1843 8116 1850
rect 8099 1840 8100 1843
rect 8115 1840 8128 1843
rect 8051 1836 8081 1837
rect 8090 1836 8096 1837
rect 8099 1836 8128 1840
rect 8018 1835 8128 1836
rect 8018 1834 8134 1835
rect 7693 1826 7744 1834
rect 7693 1814 7718 1826
rect 7725 1814 7744 1826
rect 7775 1826 7825 1834
rect 7775 1818 7791 1826
rect 7798 1824 7825 1826
rect 7834 1824 8055 1834
rect 7798 1814 8055 1824
rect 8084 1826 8134 1834
rect 8084 1817 8100 1826
rect 7693 1806 7744 1814
rect 7791 1806 8055 1814
rect 8081 1814 8100 1817
rect 8107 1814 8134 1826
rect 8081 1806 8134 1814
rect 7709 1798 7710 1806
rect 7725 1798 7738 1806
rect 7709 1790 7725 1798
rect 7706 1783 7725 1786
rect 7706 1774 7728 1783
rect 7679 1764 7728 1774
rect 7679 1758 7709 1764
rect 7728 1759 7733 1764
rect 7651 1742 7725 1758
rect 7743 1750 7773 1806
rect 7808 1796 8016 1806
rect 8051 1802 8096 1806
rect 8099 1805 8100 1806
rect 8115 1805 8128 1806
rect 7834 1766 8023 1796
rect 7849 1763 8023 1766
rect 7842 1760 8023 1763
rect 7651 1740 7664 1742
rect 7679 1740 7713 1742
rect 7651 1724 7725 1740
rect 7752 1736 7765 1750
rect 7780 1736 7796 1752
rect 7842 1747 7853 1760
rect 7635 1702 7636 1718
rect 7651 1702 7664 1724
rect 7679 1702 7709 1724
rect 7752 1720 7814 1736
rect 7842 1729 7853 1745
rect 7858 1740 7868 1760
rect 7878 1740 7892 1760
rect 7895 1747 7904 1760
rect 7920 1747 7929 1760
rect 7858 1729 7892 1740
rect 7895 1729 7904 1745
rect 7920 1729 7929 1745
rect 7936 1740 7946 1760
rect 7956 1740 7970 1760
rect 7971 1747 7982 1760
rect 7936 1729 7970 1740
rect 7971 1729 7982 1745
rect 8028 1736 8044 1752
rect 8051 1750 8081 1802
rect 8115 1798 8116 1805
rect 8100 1790 8116 1798
rect 8087 1758 8100 1777
rect 8115 1758 8145 1774
rect 8087 1742 8161 1758
rect 8087 1740 8100 1742
rect 8115 1740 8149 1742
rect 7752 1718 7765 1720
rect 7780 1718 7814 1720
rect 7752 1702 7814 1718
rect 7858 1713 7874 1716
rect 7936 1713 7966 1724
rect 8014 1720 8060 1736
rect 8087 1724 8161 1740
rect 8014 1718 8048 1720
rect 8013 1702 8060 1718
rect 8087 1702 8100 1724
rect 8115 1702 8145 1724
rect 8172 1702 8173 1718
rect 8188 1702 8201 1862
rect 8231 1758 8244 1862
rect 8289 1840 8290 1850
rect 8305 1840 8318 1850
rect 8289 1836 8318 1840
rect 8323 1836 8353 1862
rect 8371 1848 8387 1850
rect 8459 1848 8512 1862
rect 8460 1846 8524 1848
rect 8567 1846 8582 1862
rect 8631 1859 8661 1862
rect 8631 1856 8667 1859
rect 8597 1848 8613 1850
rect 8371 1836 8386 1840
rect 8289 1834 8386 1836
rect 8414 1834 8582 1846
rect 8598 1836 8613 1840
rect 8631 1837 8670 1856
rect 8689 1850 8696 1851
rect 8695 1843 8696 1850
rect 8679 1840 8680 1843
rect 8695 1840 8708 1843
rect 8631 1836 8661 1837
rect 8670 1836 8676 1837
rect 8679 1836 8708 1840
rect 8598 1835 8708 1836
rect 8598 1834 8714 1835
rect 8273 1826 8324 1834
rect 8273 1814 8298 1826
rect 8305 1814 8324 1826
rect 8355 1826 8405 1834
rect 8355 1818 8371 1826
rect 8378 1824 8405 1826
rect 8414 1824 8635 1834
rect 8378 1814 8635 1824
rect 8664 1826 8714 1834
rect 8664 1817 8680 1826
rect 8273 1806 8324 1814
rect 8371 1806 8635 1814
rect 8661 1814 8680 1817
rect 8687 1814 8714 1826
rect 8661 1806 8714 1814
rect 8289 1798 8290 1806
rect 8305 1798 8318 1806
rect 8289 1790 8305 1798
rect 8286 1783 8305 1786
rect 8286 1774 8308 1783
rect 8259 1764 8308 1774
rect 8259 1758 8289 1764
rect 8308 1759 8313 1764
rect 8231 1742 8305 1758
rect 8323 1750 8353 1806
rect 8388 1796 8596 1806
rect 8631 1802 8676 1806
rect 8679 1805 8680 1806
rect 8695 1805 8708 1806
rect 8414 1766 8603 1796
rect 8429 1763 8603 1766
rect 8422 1760 8603 1763
rect 8231 1740 8244 1742
rect 8259 1740 8293 1742
rect 8231 1724 8305 1740
rect 8332 1736 8345 1750
rect 8360 1736 8376 1752
rect 8422 1747 8433 1760
rect 8215 1702 8216 1718
rect 8231 1702 8244 1724
rect 8259 1702 8289 1724
rect 8332 1720 8394 1736
rect 8422 1729 8433 1745
rect 8438 1740 8448 1760
rect 8458 1740 8472 1760
rect 8475 1747 8484 1760
rect 8500 1747 8509 1760
rect 8438 1729 8472 1740
rect 8475 1729 8484 1745
rect 8500 1729 8509 1745
rect 8516 1740 8526 1760
rect 8536 1740 8550 1760
rect 8551 1747 8562 1760
rect 8516 1729 8550 1740
rect 8551 1729 8562 1745
rect 8608 1736 8624 1752
rect 8631 1750 8661 1802
rect 8695 1798 8696 1805
rect 8680 1790 8696 1798
rect 8667 1758 8680 1777
rect 8695 1758 8725 1774
rect 8667 1742 8741 1758
rect 8667 1740 8680 1742
rect 8695 1740 8729 1742
rect 8332 1718 8345 1720
rect 8360 1718 8394 1720
rect 8332 1702 8394 1718
rect 8438 1713 8454 1716
rect 8516 1713 8546 1724
rect 8594 1720 8640 1736
rect 8667 1724 8741 1740
rect 8594 1718 8628 1720
rect 8593 1702 8640 1718
rect 8667 1702 8680 1724
rect 8695 1702 8725 1724
rect 8752 1702 8753 1718
rect 8768 1702 8781 1862
rect 8811 1758 8824 1862
rect 8869 1840 8870 1850
rect 8885 1840 8898 1850
rect 8869 1836 8898 1840
rect 8903 1836 8933 1862
rect 8951 1848 8967 1850
rect 9039 1848 9092 1862
rect 9040 1846 9104 1848
rect 9147 1846 9162 1862
rect 9211 1859 9241 1862
rect 9211 1856 9247 1859
rect 9177 1848 9193 1850
rect 8951 1836 8966 1840
rect 8869 1834 8966 1836
rect 8994 1834 9162 1846
rect 9178 1836 9193 1840
rect 9211 1837 9250 1856
rect 9269 1850 9276 1851
rect 9275 1843 9276 1850
rect 9259 1840 9260 1843
rect 9275 1840 9288 1843
rect 9211 1836 9241 1837
rect 9250 1836 9256 1837
rect 9259 1836 9288 1840
rect 9178 1835 9288 1836
rect 9178 1834 9294 1835
rect 8853 1826 8904 1834
rect 8853 1814 8878 1826
rect 8885 1814 8904 1826
rect 8935 1826 8985 1834
rect 8935 1818 8951 1826
rect 8958 1824 8985 1826
rect 8994 1824 9215 1834
rect 8958 1814 9215 1824
rect 9244 1826 9294 1834
rect 9244 1817 9260 1826
rect 8853 1806 8904 1814
rect 8951 1806 9215 1814
rect 9241 1814 9260 1817
rect 9267 1814 9294 1826
rect 9241 1806 9294 1814
rect 8869 1798 8870 1806
rect 8885 1798 8898 1806
rect 8869 1790 8885 1798
rect 8866 1783 8885 1786
rect 8866 1774 8888 1783
rect 8839 1764 8888 1774
rect 8839 1758 8869 1764
rect 8888 1759 8893 1764
rect 8811 1742 8885 1758
rect 8903 1750 8933 1806
rect 8968 1796 9176 1806
rect 9211 1802 9256 1806
rect 9259 1805 9260 1806
rect 9275 1805 9288 1806
rect 8994 1766 9183 1796
rect 9009 1763 9183 1766
rect 9002 1760 9183 1763
rect 8811 1740 8824 1742
rect 8839 1740 8873 1742
rect 8811 1724 8885 1740
rect 8912 1736 8925 1750
rect 8940 1736 8956 1752
rect 9002 1747 9013 1760
rect 8795 1702 8796 1718
rect 8811 1702 8824 1724
rect 8839 1702 8869 1724
rect 8912 1720 8974 1736
rect 9002 1729 9013 1745
rect 9018 1740 9028 1760
rect 9038 1740 9052 1760
rect 9055 1747 9064 1760
rect 9080 1747 9089 1760
rect 9018 1729 9052 1740
rect 9055 1729 9064 1745
rect 9080 1729 9089 1745
rect 9096 1740 9106 1760
rect 9116 1740 9130 1760
rect 9131 1747 9142 1760
rect 9096 1729 9130 1740
rect 9131 1729 9142 1745
rect 9188 1736 9204 1752
rect 9211 1750 9241 1802
rect 9275 1798 9276 1805
rect 9260 1790 9276 1798
rect 9247 1758 9260 1777
rect 9275 1758 9305 1774
rect 9247 1742 9321 1758
rect 9247 1740 9260 1742
rect 9275 1740 9309 1742
rect 8912 1718 8925 1720
rect 8940 1718 8974 1720
rect 8912 1702 8974 1718
rect 9018 1713 9034 1716
rect 9096 1713 9126 1724
rect 9174 1720 9220 1736
rect 9247 1724 9321 1740
rect 9174 1718 9208 1720
rect 9173 1702 9220 1718
rect 9247 1702 9260 1724
rect 9275 1702 9305 1724
rect 9332 1702 9333 1718
rect 9348 1702 9361 1862
rect -9 1694 32 1702
rect -9 1668 6 1694
rect 13 1668 32 1694
rect 96 1690 158 1702
rect 170 1690 245 1702
rect 303 1690 378 1702
rect 390 1690 421 1702
rect 427 1690 462 1702
rect 96 1688 258 1690
rect -9 1660 32 1668
rect 114 1664 127 1688
rect 142 1686 157 1688
rect -3 1650 -2 1660
rect 13 1650 26 1660
rect 41 1650 71 1664
rect 114 1650 157 1664
rect 181 1661 188 1668
rect 191 1664 258 1688
rect 290 1688 462 1690
rect 260 1666 288 1670
rect 290 1666 370 1688
rect 391 1686 406 1688
rect 260 1664 370 1666
rect 191 1660 370 1664
rect 164 1650 194 1660
rect 196 1650 349 1660
rect 357 1650 387 1660
rect 391 1650 421 1664
rect 449 1650 462 1688
rect 534 1694 569 1702
rect 534 1668 535 1694
rect 542 1668 569 1694
rect 477 1650 507 1664
rect 534 1660 569 1668
rect 571 1694 612 1702
rect 571 1668 586 1694
rect 593 1668 612 1694
rect 676 1690 738 1702
rect 750 1690 825 1702
rect 883 1690 958 1702
rect 970 1690 1001 1702
rect 1007 1690 1042 1702
rect 676 1688 838 1690
rect 571 1660 612 1668
rect 694 1664 707 1688
rect 722 1686 737 1688
rect 534 1650 535 1660
rect 550 1650 563 1660
rect 577 1650 578 1660
rect 593 1650 606 1660
rect 621 1650 651 1664
rect 694 1650 737 1664
rect 761 1661 768 1668
rect 771 1664 838 1688
rect 870 1688 1042 1690
rect 840 1666 868 1670
rect 870 1666 950 1688
rect 971 1686 986 1688
rect 840 1664 950 1666
rect 771 1660 950 1664
rect 744 1650 774 1660
rect 776 1650 929 1660
rect 937 1650 967 1660
rect 971 1650 1001 1664
rect 1029 1650 1042 1688
rect 1114 1694 1149 1702
rect 1114 1668 1115 1694
rect 1122 1668 1149 1694
rect 1057 1650 1087 1664
rect 1114 1660 1149 1668
rect 1151 1694 1192 1702
rect 1151 1668 1166 1694
rect 1173 1668 1192 1694
rect 1256 1690 1318 1702
rect 1330 1690 1405 1702
rect 1463 1690 1538 1702
rect 1550 1690 1581 1702
rect 1587 1690 1622 1702
rect 1256 1688 1418 1690
rect 1151 1660 1192 1668
rect 1274 1664 1287 1688
rect 1302 1686 1317 1688
rect 1114 1650 1115 1660
rect 1130 1650 1143 1660
rect 1157 1650 1158 1660
rect 1173 1650 1186 1660
rect 1201 1650 1231 1664
rect 1274 1650 1317 1664
rect 1341 1661 1348 1668
rect 1351 1664 1418 1688
rect 1450 1688 1622 1690
rect 1420 1666 1448 1670
rect 1450 1666 1530 1688
rect 1551 1686 1566 1688
rect 1420 1664 1530 1666
rect 1351 1660 1530 1664
rect 1324 1650 1354 1660
rect 1356 1650 1509 1660
rect 1517 1650 1547 1660
rect 1551 1650 1581 1664
rect 1609 1650 1622 1688
rect 1694 1694 1729 1702
rect 1694 1668 1695 1694
rect 1702 1668 1729 1694
rect 1637 1650 1667 1664
rect 1694 1660 1729 1668
rect 1731 1694 1772 1702
rect 1731 1668 1746 1694
rect 1753 1668 1772 1694
rect 1836 1690 1898 1702
rect 1910 1690 1985 1702
rect 2043 1690 2118 1702
rect 2130 1690 2161 1702
rect 2167 1690 2202 1702
rect 1836 1688 1998 1690
rect 1731 1660 1772 1668
rect 1854 1664 1867 1688
rect 1882 1686 1897 1688
rect 1694 1650 1695 1660
rect 1710 1650 1723 1660
rect 1737 1650 1738 1660
rect 1753 1650 1766 1660
rect 1781 1650 1811 1664
rect 1854 1650 1897 1664
rect 1921 1661 1928 1668
rect 1931 1664 1998 1688
rect 2030 1688 2202 1690
rect 2000 1666 2028 1670
rect 2030 1666 2110 1688
rect 2131 1686 2146 1688
rect 2000 1664 2110 1666
rect 1931 1660 2110 1664
rect 1904 1650 1934 1660
rect 1936 1650 2089 1660
rect 2097 1650 2127 1660
rect 2131 1650 2161 1664
rect 2189 1650 2202 1688
rect 2274 1694 2309 1702
rect 2274 1668 2275 1694
rect 2282 1668 2309 1694
rect 2217 1650 2247 1664
rect 2274 1660 2309 1668
rect 2311 1694 2352 1702
rect 2311 1668 2326 1694
rect 2333 1668 2352 1694
rect 2416 1690 2478 1702
rect 2490 1690 2565 1702
rect 2623 1690 2698 1702
rect 2710 1690 2741 1702
rect 2747 1690 2782 1702
rect 2416 1688 2578 1690
rect 2311 1660 2352 1668
rect 2434 1664 2447 1688
rect 2462 1686 2477 1688
rect 2274 1650 2275 1660
rect 2290 1650 2303 1660
rect 2317 1650 2318 1660
rect 2333 1650 2346 1660
rect 2361 1650 2391 1664
rect 2434 1650 2477 1664
rect 2501 1661 2508 1668
rect 2511 1664 2578 1688
rect 2610 1688 2782 1690
rect 2580 1666 2608 1670
rect 2610 1666 2690 1688
rect 2711 1686 2726 1688
rect 2580 1664 2690 1666
rect 2511 1660 2690 1664
rect 2484 1650 2514 1660
rect 2516 1650 2669 1660
rect 2677 1650 2707 1660
rect 2711 1650 2741 1664
rect 2769 1650 2782 1688
rect 2854 1694 2889 1702
rect 2854 1668 2855 1694
rect 2862 1668 2889 1694
rect 2797 1650 2827 1664
rect 2854 1660 2889 1668
rect 2891 1694 2932 1702
rect 2891 1668 2906 1694
rect 2913 1668 2932 1694
rect 2996 1690 3058 1702
rect 3070 1690 3145 1702
rect 3203 1690 3278 1702
rect 3290 1690 3321 1702
rect 3327 1690 3362 1702
rect 2996 1688 3158 1690
rect 2891 1660 2932 1668
rect 3014 1664 3027 1688
rect 3042 1686 3057 1688
rect 2854 1650 2855 1660
rect 2870 1650 2883 1660
rect 2897 1650 2898 1660
rect 2913 1650 2926 1660
rect 2941 1650 2971 1664
rect 3014 1650 3057 1664
rect 3081 1661 3088 1668
rect 3091 1664 3158 1688
rect 3190 1688 3362 1690
rect 3160 1666 3188 1670
rect 3190 1666 3270 1688
rect 3291 1686 3306 1688
rect 3160 1664 3270 1666
rect 3091 1660 3270 1664
rect 3064 1650 3094 1660
rect 3096 1650 3249 1660
rect 3257 1650 3287 1660
rect 3291 1650 3321 1664
rect 3349 1650 3362 1688
rect 3434 1694 3469 1702
rect 3434 1668 3435 1694
rect 3442 1668 3469 1694
rect 3377 1650 3407 1664
rect 3434 1660 3469 1668
rect 3434 1650 3435 1660
rect 3450 1650 3463 1660
rect -3 1644 3469 1650
rect -2 1636 3469 1644
rect 5889 1694 5930 1702
rect 5889 1668 5904 1694
rect 5911 1668 5930 1694
rect 5994 1690 6056 1702
rect 6068 1690 6143 1702
rect 6201 1690 6276 1702
rect 6288 1690 6319 1702
rect 6325 1690 6360 1702
rect 5994 1688 6156 1690
rect 5889 1660 5930 1668
rect 6012 1664 6025 1688
rect 6040 1686 6055 1688
rect 5895 1650 5896 1660
rect 5911 1650 5924 1660
rect 5939 1650 5969 1664
rect 6012 1650 6055 1664
rect 6079 1661 6086 1668
rect 6089 1664 6156 1688
rect 6188 1688 6360 1690
rect 6158 1666 6186 1670
rect 6188 1666 6268 1688
rect 6289 1686 6304 1688
rect 6158 1664 6268 1666
rect 6089 1660 6268 1664
rect 6062 1650 6092 1660
rect 6094 1650 6247 1660
rect 6255 1650 6285 1660
rect 6289 1650 6319 1664
rect 6347 1650 6360 1688
rect 6432 1694 6467 1702
rect 6432 1668 6433 1694
rect 6440 1668 6467 1694
rect 6375 1650 6405 1664
rect 6432 1660 6467 1668
rect 6469 1694 6510 1702
rect 6469 1668 6484 1694
rect 6491 1668 6510 1694
rect 6574 1690 6636 1702
rect 6648 1690 6723 1702
rect 6781 1690 6856 1702
rect 6868 1690 6899 1702
rect 6905 1690 6940 1702
rect 6574 1688 6736 1690
rect 6469 1660 6510 1668
rect 6592 1664 6605 1688
rect 6620 1686 6635 1688
rect 6432 1650 6433 1660
rect 6448 1650 6461 1660
rect 6475 1650 6476 1660
rect 6491 1650 6504 1660
rect 6519 1650 6549 1664
rect 6592 1650 6635 1664
rect 6659 1661 6666 1668
rect 6669 1664 6736 1688
rect 6768 1688 6940 1690
rect 6738 1666 6766 1670
rect 6768 1666 6848 1688
rect 6869 1686 6884 1688
rect 6738 1664 6848 1666
rect 6669 1660 6848 1664
rect 6642 1650 6672 1660
rect 6674 1650 6827 1660
rect 6835 1650 6865 1660
rect 6869 1650 6899 1664
rect 6927 1650 6940 1688
rect 7012 1694 7047 1702
rect 7012 1668 7013 1694
rect 7020 1668 7047 1694
rect 6955 1650 6985 1664
rect 7012 1660 7047 1668
rect 7049 1694 7090 1702
rect 7049 1668 7064 1694
rect 7071 1668 7090 1694
rect 7154 1690 7216 1702
rect 7228 1690 7303 1702
rect 7361 1690 7436 1702
rect 7448 1690 7479 1702
rect 7485 1690 7520 1702
rect 7154 1688 7316 1690
rect 7049 1660 7090 1668
rect 7172 1664 7185 1688
rect 7200 1686 7215 1688
rect 7012 1650 7013 1660
rect 7028 1650 7041 1660
rect 7055 1650 7056 1660
rect 7071 1650 7084 1660
rect 7099 1650 7129 1664
rect 7172 1650 7215 1664
rect 7239 1661 7246 1668
rect 7249 1664 7316 1688
rect 7348 1688 7520 1690
rect 7318 1666 7346 1670
rect 7348 1666 7428 1688
rect 7449 1686 7464 1688
rect 7318 1664 7428 1666
rect 7249 1660 7428 1664
rect 7222 1650 7252 1660
rect 7254 1650 7407 1660
rect 7415 1650 7445 1660
rect 7449 1650 7479 1664
rect 7507 1650 7520 1688
rect 7592 1694 7627 1702
rect 7592 1668 7593 1694
rect 7600 1668 7627 1694
rect 7535 1650 7565 1664
rect 7592 1660 7627 1668
rect 7629 1694 7670 1702
rect 7629 1668 7644 1694
rect 7651 1668 7670 1694
rect 7734 1690 7796 1702
rect 7808 1690 7883 1702
rect 7941 1690 8016 1702
rect 8028 1690 8059 1702
rect 8065 1690 8100 1702
rect 7734 1688 7896 1690
rect 7629 1660 7670 1668
rect 7752 1664 7765 1688
rect 7780 1686 7795 1688
rect 7592 1650 7593 1660
rect 7608 1650 7621 1660
rect 7635 1650 7636 1660
rect 7651 1650 7664 1660
rect 7679 1650 7709 1664
rect 7752 1650 7795 1664
rect 7819 1661 7826 1668
rect 7829 1664 7896 1688
rect 7928 1688 8100 1690
rect 7898 1666 7926 1670
rect 7928 1666 8008 1688
rect 8029 1686 8044 1688
rect 7898 1664 8008 1666
rect 7829 1660 8008 1664
rect 7802 1650 7832 1660
rect 7834 1650 7987 1660
rect 7995 1650 8025 1660
rect 8029 1650 8059 1664
rect 8087 1650 8100 1688
rect 8172 1694 8207 1702
rect 8172 1668 8173 1694
rect 8180 1668 8207 1694
rect 8115 1650 8145 1664
rect 8172 1660 8207 1668
rect 8209 1694 8250 1702
rect 8209 1668 8224 1694
rect 8231 1668 8250 1694
rect 8314 1690 8376 1702
rect 8388 1690 8463 1702
rect 8521 1690 8596 1702
rect 8608 1690 8639 1702
rect 8645 1690 8680 1702
rect 8314 1688 8476 1690
rect 8209 1660 8250 1668
rect 8332 1664 8345 1688
rect 8360 1686 8375 1688
rect 8172 1650 8173 1660
rect 8188 1650 8201 1660
rect 8215 1650 8216 1660
rect 8231 1650 8244 1660
rect 8259 1650 8289 1664
rect 8332 1650 8375 1664
rect 8399 1661 8406 1668
rect 8409 1664 8476 1688
rect 8508 1688 8680 1690
rect 8478 1666 8506 1670
rect 8508 1666 8588 1688
rect 8609 1686 8624 1688
rect 8478 1664 8588 1666
rect 8409 1660 8588 1664
rect 8382 1650 8412 1660
rect 8414 1650 8567 1660
rect 8575 1650 8605 1660
rect 8609 1650 8639 1664
rect 8667 1650 8680 1688
rect 8752 1694 8787 1702
rect 8752 1668 8753 1694
rect 8760 1668 8787 1694
rect 8695 1650 8725 1664
rect 8752 1660 8787 1668
rect 8789 1694 8830 1702
rect 8789 1668 8804 1694
rect 8811 1668 8830 1694
rect 8894 1690 8956 1702
rect 8968 1690 9043 1702
rect 9101 1690 9176 1702
rect 9188 1690 9219 1702
rect 9225 1690 9260 1702
rect 8894 1688 9056 1690
rect 8789 1660 8830 1668
rect 8912 1664 8925 1688
rect 8940 1686 8955 1688
rect 8752 1650 8753 1660
rect 8768 1650 8781 1660
rect 8795 1650 8796 1660
rect 8811 1650 8824 1660
rect 8839 1650 8869 1664
rect 8912 1650 8955 1664
rect 8979 1661 8986 1668
rect 8989 1664 9056 1688
rect 9088 1688 9260 1690
rect 9058 1666 9086 1670
rect 9088 1666 9168 1688
rect 9189 1686 9204 1688
rect 9058 1664 9168 1666
rect 8989 1660 9168 1664
rect 8962 1650 8992 1660
rect 8994 1650 9147 1660
rect 9155 1650 9185 1660
rect 9189 1650 9219 1664
rect 9247 1650 9260 1688
rect 9332 1694 9367 1702
rect 9332 1668 9333 1694
rect 9340 1668 9367 1694
rect 9275 1650 9305 1664
rect 9332 1660 9367 1668
rect 9332 1650 9333 1660
rect 9348 1650 9361 1660
rect 5889 1636 9361 1650
rect 13 1606 26 1636
rect 41 1618 71 1636
rect 114 1622 128 1636
rect 164 1622 384 1636
rect 115 1620 128 1622
rect 81 1608 96 1620
rect 78 1606 100 1608
rect 105 1606 135 1620
rect 196 1618 349 1622
rect 178 1606 370 1618
rect 413 1606 443 1620
rect 449 1606 462 1636
rect 477 1618 507 1636
rect 550 1606 563 1636
rect 593 1606 606 1636
rect 621 1618 651 1636
rect 694 1622 708 1636
rect 744 1622 964 1636
rect 695 1620 708 1622
rect 661 1608 676 1620
rect 658 1606 680 1608
rect 685 1606 715 1620
rect 776 1618 929 1622
rect 758 1606 950 1618
rect 993 1606 1023 1620
rect 1029 1606 1042 1636
rect 1057 1618 1087 1636
rect 1130 1606 1143 1636
rect 1173 1606 1186 1636
rect 1201 1618 1231 1636
rect 1274 1622 1288 1636
rect 1324 1622 1544 1636
rect 1275 1620 1288 1622
rect 1241 1608 1256 1620
rect 1238 1606 1260 1608
rect 1265 1606 1295 1620
rect 1356 1618 1509 1622
rect 1338 1606 1530 1618
rect 1573 1606 1603 1620
rect 1609 1606 1622 1636
rect 1637 1618 1667 1636
rect 1710 1606 1723 1636
rect 1753 1606 1766 1636
rect 1781 1618 1811 1636
rect 1854 1622 1868 1636
rect 1904 1622 2124 1636
rect 1855 1620 1868 1622
rect 1821 1608 1836 1620
rect 1818 1606 1840 1608
rect 1845 1606 1875 1620
rect 1936 1618 2089 1622
rect 1918 1606 2110 1618
rect 2153 1606 2183 1620
rect 2189 1606 2202 1636
rect 2217 1618 2247 1636
rect 2290 1606 2303 1636
rect 2333 1606 2346 1636
rect 2361 1618 2391 1636
rect 2434 1622 2448 1636
rect 2484 1622 2704 1636
rect 2435 1620 2448 1622
rect 2401 1608 2416 1620
rect 2398 1606 2420 1608
rect 2425 1606 2455 1620
rect 2516 1618 2669 1622
rect 2498 1606 2690 1618
rect 2733 1606 2763 1620
rect 2769 1606 2782 1636
rect 2797 1618 2827 1636
rect 2870 1606 2883 1636
rect 2913 1606 2926 1636
rect 2941 1618 2971 1636
rect 3014 1622 3028 1636
rect 3064 1622 3284 1636
rect 3015 1620 3028 1622
rect 2981 1608 2996 1620
rect 2978 1606 3000 1608
rect 3005 1606 3035 1620
rect 3096 1618 3249 1622
rect 3078 1606 3270 1618
rect 3313 1606 3343 1620
rect 3349 1606 3362 1636
rect 3377 1618 3407 1636
rect 3450 1606 3463 1636
rect 5911 1606 5924 1636
rect 5939 1618 5969 1636
rect 6012 1622 6026 1636
rect 6062 1622 6282 1636
rect 6013 1620 6026 1622
rect 5979 1608 5994 1620
rect 5976 1606 5998 1608
rect 6003 1606 6033 1620
rect 6094 1618 6247 1622
rect 6076 1606 6268 1618
rect 6311 1606 6341 1620
rect 6347 1606 6360 1636
rect 6375 1618 6405 1636
rect 6448 1606 6461 1636
rect 6491 1606 6504 1636
rect 6519 1618 6549 1636
rect 6592 1622 6606 1636
rect 6642 1622 6862 1636
rect 6593 1620 6606 1622
rect 6559 1608 6574 1620
rect 6556 1606 6578 1608
rect 6583 1606 6613 1620
rect 6674 1618 6827 1622
rect 6656 1606 6848 1618
rect 6891 1606 6921 1620
rect 6927 1606 6940 1636
rect 6955 1618 6985 1636
rect 7028 1606 7041 1636
rect 7071 1606 7084 1636
rect 7099 1618 7129 1636
rect 7172 1622 7186 1636
rect 7222 1622 7442 1636
rect 7173 1620 7186 1622
rect 7139 1608 7154 1620
rect 7136 1606 7158 1608
rect 7163 1606 7193 1620
rect 7254 1618 7407 1622
rect 7236 1606 7428 1618
rect 7471 1606 7501 1620
rect 7507 1606 7520 1636
rect 7535 1618 7565 1636
rect 7608 1606 7621 1636
rect 7651 1606 7664 1636
rect 7679 1618 7709 1636
rect 7752 1622 7766 1636
rect 7802 1622 8022 1636
rect 7753 1620 7766 1622
rect 7719 1608 7734 1620
rect 7716 1606 7738 1608
rect 7743 1606 7773 1620
rect 7834 1618 7987 1622
rect 7816 1606 8008 1618
rect 8051 1606 8081 1620
rect 8087 1606 8100 1636
rect 8115 1618 8145 1636
rect 8188 1606 8201 1636
rect 8231 1606 8244 1636
rect 8259 1618 8289 1636
rect 8332 1622 8346 1636
rect 8382 1622 8602 1636
rect 8333 1620 8346 1622
rect 8299 1608 8314 1620
rect 8296 1606 8318 1608
rect 8323 1606 8353 1620
rect 8414 1618 8567 1622
rect 8396 1606 8588 1618
rect 8631 1606 8661 1620
rect 8667 1606 8680 1636
rect 8695 1618 8725 1636
rect 8768 1606 8781 1636
rect 8811 1606 8824 1636
rect 8839 1618 8869 1636
rect 8912 1622 8926 1636
rect 8962 1622 9182 1636
rect 8913 1620 8926 1622
rect 8879 1608 8894 1620
rect 8876 1606 8898 1608
rect 8903 1606 8933 1620
rect 8994 1618 9147 1622
rect 8976 1606 9168 1618
rect 9211 1606 9241 1620
rect 9247 1606 9260 1636
rect 9275 1618 9305 1636
rect 9348 1606 9361 1636
rect -2 1592 3469 1606
rect 5889 1592 9361 1606
rect 13 1488 26 1592
rect 71 1570 72 1580
rect 87 1570 100 1580
rect 71 1566 100 1570
rect 105 1566 135 1592
rect 153 1578 169 1580
rect 241 1578 294 1592
rect 242 1576 306 1578
rect 349 1576 364 1592
rect 413 1589 443 1592
rect 413 1586 449 1589
rect 379 1578 395 1580
rect 153 1566 168 1570
rect 71 1564 168 1566
rect 196 1564 364 1576
rect 380 1566 395 1570
rect 413 1567 452 1586
rect 471 1580 478 1581
rect 477 1573 478 1580
rect 461 1570 462 1573
rect 477 1570 490 1573
rect 413 1566 443 1567
rect 452 1566 458 1567
rect 461 1566 490 1570
rect 380 1565 490 1566
rect 380 1564 496 1565
rect 55 1556 106 1564
rect 55 1544 80 1556
rect 87 1544 106 1556
rect 137 1556 187 1564
rect 137 1548 153 1556
rect 160 1554 187 1556
rect 196 1554 417 1564
rect 160 1544 417 1554
rect 446 1556 496 1564
rect 446 1547 462 1556
rect 55 1536 106 1544
rect 153 1536 417 1544
rect 443 1544 462 1547
rect 469 1544 496 1556
rect 443 1536 496 1544
rect 71 1528 72 1536
rect 87 1528 100 1536
rect 71 1520 87 1528
rect 68 1513 87 1516
rect 68 1504 90 1513
rect 41 1494 90 1504
rect 41 1488 71 1494
rect 90 1489 95 1494
rect 13 1472 87 1488
rect 105 1480 135 1536
rect 170 1526 378 1536
rect 413 1532 458 1536
rect 461 1535 462 1536
rect 477 1535 490 1536
rect 196 1496 385 1526
rect 211 1493 385 1496
rect 204 1490 385 1493
rect 13 1470 26 1472
rect 41 1470 75 1472
rect 13 1454 87 1470
rect 114 1466 127 1480
rect 142 1466 158 1482
rect 204 1477 215 1490
rect -3 1432 -2 1448
rect 13 1432 26 1454
rect 41 1432 71 1454
rect 114 1450 176 1466
rect 204 1459 215 1475
rect 220 1470 230 1490
rect 240 1470 254 1490
rect 257 1477 266 1490
rect 282 1477 291 1490
rect 220 1459 254 1470
rect 257 1459 266 1475
rect 282 1459 291 1475
rect 298 1470 308 1490
rect 318 1470 332 1490
rect 333 1477 344 1490
rect 298 1459 332 1470
rect 333 1459 344 1475
rect 390 1466 406 1482
rect 413 1480 443 1532
rect 477 1528 478 1535
rect 462 1520 478 1528
rect 449 1488 462 1507
rect 477 1488 507 1504
rect 449 1472 523 1488
rect 449 1470 462 1472
rect 477 1470 511 1472
rect 114 1448 127 1450
rect 142 1448 176 1450
rect 114 1432 176 1448
rect 220 1443 236 1446
rect 298 1443 328 1454
rect 376 1450 422 1466
rect 449 1454 523 1470
rect 376 1448 410 1450
rect 375 1432 422 1448
rect 449 1432 462 1454
rect 477 1432 507 1454
rect 534 1432 535 1448
rect 550 1432 563 1592
rect 593 1488 606 1592
rect 651 1570 652 1580
rect 667 1570 680 1580
rect 651 1566 680 1570
rect 685 1566 715 1592
rect 733 1578 749 1580
rect 821 1578 874 1592
rect 822 1576 886 1578
rect 929 1576 944 1592
rect 993 1589 1023 1592
rect 993 1586 1029 1589
rect 959 1578 975 1580
rect 733 1566 748 1570
rect 651 1564 748 1566
rect 776 1564 944 1576
rect 960 1566 975 1570
rect 993 1567 1032 1586
rect 1051 1580 1058 1581
rect 1057 1573 1058 1580
rect 1041 1570 1042 1573
rect 1057 1570 1070 1573
rect 993 1566 1023 1567
rect 1032 1566 1038 1567
rect 1041 1566 1070 1570
rect 960 1565 1070 1566
rect 960 1564 1076 1565
rect 635 1556 686 1564
rect 635 1544 660 1556
rect 667 1544 686 1556
rect 717 1556 767 1564
rect 717 1548 733 1556
rect 740 1554 767 1556
rect 776 1554 997 1564
rect 740 1544 997 1554
rect 1026 1556 1076 1564
rect 1026 1547 1042 1556
rect 635 1536 686 1544
rect 733 1536 997 1544
rect 1023 1544 1042 1547
rect 1049 1544 1076 1556
rect 1023 1536 1076 1544
rect 651 1528 652 1536
rect 667 1528 680 1536
rect 651 1520 667 1528
rect 648 1513 667 1516
rect 648 1504 670 1513
rect 621 1494 670 1504
rect 621 1488 651 1494
rect 670 1489 675 1494
rect 593 1472 667 1488
rect 685 1480 715 1536
rect 750 1526 958 1536
rect 993 1532 1038 1536
rect 1041 1535 1042 1536
rect 1057 1535 1070 1536
rect 776 1496 965 1526
rect 791 1493 965 1496
rect 784 1490 965 1493
rect 593 1470 606 1472
rect 621 1470 655 1472
rect 593 1454 667 1470
rect 694 1466 707 1480
rect 722 1466 738 1482
rect 784 1477 795 1490
rect 577 1432 578 1448
rect 593 1432 606 1454
rect 621 1432 651 1454
rect 694 1450 756 1466
rect 784 1459 795 1475
rect 800 1470 810 1490
rect 820 1470 834 1490
rect 837 1477 846 1490
rect 862 1477 871 1490
rect 800 1459 834 1470
rect 837 1459 846 1475
rect 862 1459 871 1475
rect 878 1470 888 1490
rect 898 1470 912 1490
rect 913 1477 924 1490
rect 878 1459 912 1470
rect 913 1459 924 1475
rect 970 1466 986 1482
rect 993 1480 1023 1532
rect 1057 1528 1058 1535
rect 1042 1520 1058 1528
rect 1029 1488 1042 1507
rect 1057 1488 1087 1504
rect 1029 1472 1103 1488
rect 1029 1470 1042 1472
rect 1057 1470 1091 1472
rect 694 1448 707 1450
rect 722 1448 756 1450
rect 694 1432 756 1448
rect 800 1443 816 1446
rect 878 1443 908 1454
rect 956 1450 1002 1466
rect 1029 1454 1103 1470
rect 956 1448 990 1450
rect 955 1432 1002 1448
rect 1029 1432 1042 1454
rect 1057 1432 1087 1454
rect 1114 1432 1115 1448
rect 1130 1432 1143 1592
rect 1173 1488 1186 1592
rect 1231 1570 1232 1580
rect 1247 1570 1260 1580
rect 1231 1566 1260 1570
rect 1265 1566 1295 1592
rect 1313 1578 1329 1580
rect 1401 1578 1454 1592
rect 1402 1576 1466 1578
rect 1509 1576 1524 1592
rect 1573 1589 1603 1592
rect 1573 1586 1609 1589
rect 1539 1578 1555 1580
rect 1313 1566 1328 1570
rect 1231 1564 1328 1566
rect 1356 1564 1524 1576
rect 1540 1566 1555 1570
rect 1573 1567 1612 1586
rect 1631 1580 1638 1581
rect 1637 1573 1638 1580
rect 1621 1570 1622 1573
rect 1637 1570 1650 1573
rect 1573 1566 1603 1567
rect 1612 1566 1618 1567
rect 1621 1566 1650 1570
rect 1540 1565 1650 1566
rect 1540 1564 1656 1565
rect 1215 1556 1266 1564
rect 1215 1544 1240 1556
rect 1247 1544 1266 1556
rect 1297 1556 1347 1564
rect 1297 1548 1313 1556
rect 1320 1554 1347 1556
rect 1356 1554 1577 1564
rect 1320 1544 1577 1554
rect 1606 1556 1656 1564
rect 1606 1547 1622 1556
rect 1215 1536 1266 1544
rect 1313 1536 1577 1544
rect 1603 1544 1622 1547
rect 1629 1544 1656 1556
rect 1603 1536 1656 1544
rect 1231 1528 1232 1536
rect 1247 1528 1260 1536
rect 1231 1520 1247 1528
rect 1228 1513 1247 1516
rect 1228 1504 1250 1513
rect 1201 1494 1250 1504
rect 1201 1488 1231 1494
rect 1250 1489 1255 1494
rect 1173 1472 1247 1488
rect 1265 1480 1295 1536
rect 1330 1526 1538 1536
rect 1573 1532 1618 1536
rect 1621 1535 1622 1536
rect 1637 1535 1650 1536
rect 1356 1496 1545 1526
rect 1371 1493 1545 1496
rect 1364 1490 1545 1493
rect 1173 1470 1186 1472
rect 1201 1470 1235 1472
rect 1173 1454 1247 1470
rect 1274 1466 1287 1480
rect 1302 1466 1318 1482
rect 1364 1477 1375 1490
rect 1157 1432 1158 1448
rect 1173 1432 1186 1454
rect 1201 1432 1231 1454
rect 1274 1450 1336 1466
rect 1364 1459 1375 1475
rect 1380 1470 1390 1490
rect 1400 1470 1414 1490
rect 1417 1477 1426 1490
rect 1442 1477 1451 1490
rect 1380 1459 1414 1470
rect 1417 1459 1426 1475
rect 1442 1459 1451 1475
rect 1458 1470 1468 1490
rect 1478 1470 1492 1490
rect 1493 1477 1504 1490
rect 1458 1459 1492 1470
rect 1493 1459 1504 1475
rect 1550 1466 1566 1482
rect 1573 1480 1603 1532
rect 1637 1528 1638 1535
rect 1622 1520 1638 1528
rect 1609 1488 1622 1507
rect 1637 1488 1667 1504
rect 1609 1472 1683 1488
rect 1609 1470 1622 1472
rect 1637 1470 1671 1472
rect 1274 1448 1287 1450
rect 1302 1448 1336 1450
rect 1274 1432 1336 1448
rect 1380 1443 1396 1446
rect 1458 1443 1488 1454
rect 1536 1450 1582 1466
rect 1609 1454 1683 1470
rect 1536 1448 1570 1450
rect 1535 1432 1582 1448
rect 1609 1432 1622 1454
rect 1637 1432 1667 1454
rect 1694 1432 1695 1448
rect 1710 1432 1723 1592
rect 1753 1488 1766 1592
rect 1811 1570 1812 1580
rect 1827 1570 1840 1580
rect 1811 1566 1840 1570
rect 1845 1566 1875 1592
rect 1893 1578 1909 1580
rect 1981 1578 2034 1592
rect 1982 1576 2046 1578
rect 2089 1576 2104 1592
rect 2153 1589 2183 1592
rect 2153 1586 2189 1589
rect 2119 1578 2135 1580
rect 1893 1566 1908 1570
rect 1811 1564 1908 1566
rect 1936 1564 2104 1576
rect 2120 1566 2135 1570
rect 2153 1567 2192 1586
rect 2211 1580 2218 1581
rect 2217 1573 2218 1580
rect 2201 1570 2202 1573
rect 2217 1570 2230 1573
rect 2153 1566 2183 1567
rect 2192 1566 2198 1567
rect 2201 1566 2230 1570
rect 2120 1565 2230 1566
rect 2120 1564 2236 1565
rect 1795 1556 1846 1564
rect 1795 1544 1820 1556
rect 1827 1544 1846 1556
rect 1877 1556 1927 1564
rect 1877 1548 1893 1556
rect 1900 1554 1927 1556
rect 1936 1554 2157 1564
rect 1900 1544 2157 1554
rect 2186 1556 2236 1564
rect 2186 1547 2202 1556
rect 1795 1536 1846 1544
rect 1893 1536 2157 1544
rect 2183 1544 2202 1547
rect 2209 1544 2236 1556
rect 2183 1536 2236 1544
rect 1811 1528 1812 1536
rect 1827 1528 1840 1536
rect 1811 1520 1827 1528
rect 1808 1513 1827 1516
rect 1808 1504 1830 1513
rect 1781 1494 1830 1504
rect 1781 1488 1811 1494
rect 1830 1489 1835 1494
rect 1753 1472 1827 1488
rect 1845 1480 1875 1536
rect 1910 1526 2118 1536
rect 2153 1532 2198 1536
rect 2201 1535 2202 1536
rect 2217 1535 2230 1536
rect 1936 1496 2125 1526
rect 1951 1493 2125 1496
rect 1944 1490 2125 1493
rect 1753 1470 1766 1472
rect 1781 1470 1815 1472
rect 1753 1454 1827 1470
rect 1854 1466 1867 1480
rect 1882 1466 1898 1482
rect 1944 1477 1955 1490
rect 1737 1432 1738 1448
rect 1753 1432 1766 1454
rect 1781 1432 1811 1454
rect 1854 1450 1916 1466
rect 1944 1459 1955 1475
rect 1960 1470 1970 1490
rect 1980 1470 1994 1490
rect 1997 1477 2006 1490
rect 2022 1477 2031 1490
rect 1960 1459 1994 1470
rect 1997 1459 2006 1475
rect 2022 1459 2031 1475
rect 2038 1470 2048 1490
rect 2058 1470 2072 1490
rect 2073 1477 2084 1490
rect 2038 1459 2072 1470
rect 2073 1459 2084 1475
rect 2130 1466 2146 1482
rect 2153 1480 2183 1532
rect 2217 1528 2218 1535
rect 2202 1520 2218 1528
rect 2189 1488 2202 1507
rect 2217 1488 2247 1504
rect 2189 1472 2263 1488
rect 2189 1470 2202 1472
rect 2217 1470 2251 1472
rect 1854 1448 1867 1450
rect 1882 1448 1916 1450
rect 1854 1432 1916 1448
rect 1960 1443 1976 1446
rect 2038 1443 2068 1454
rect 2116 1450 2162 1466
rect 2189 1454 2263 1470
rect 2116 1448 2150 1450
rect 2115 1432 2162 1448
rect 2189 1432 2202 1454
rect 2217 1432 2247 1454
rect 2274 1432 2275 1448
rect 2290 1432 2303 1592
rect 2333 1488 2346 1592
rect 2391 1570 2392 1580
rect 2407 1570 2420 1580
rect 2391 1566 2420 1570
rect 2425 1566 2455 1592
rect 2473 1578 2489 1580
rect 2561 1578 2614 1592
rect 2562 1576 2626 1578
rect 2669 1576 2684 1592
rect 2733 1589 2763 1592
rect 2733 1586 2769 1589
rect 2699 1578 2715 1580
rect 2473 1566 2488 1570
rect 2391 1564 2488 1566
rect 2516 1564 2684 1576
rect 2700 1566 2715 1570
rect 2733 1567 2772 1586
rect 2791 1580 2798 1581
rect 2797 1573 2798 1580
rect 2781 1570 2782 1573
rect 2797 1570 2810 1573
rect 2733 1566 2763 1567
rect 2772 1566 2778 1567
rect 2781 1566 2810 1570
rect 2700 1565 2810 1566
rect 2700 1564 2816 1565
rect 2375 1556 2426 1564
rect 2375 1544 2400 1556
rect 2407 1544 2426 1556
rect 2457 1556 2507 1564
rect 2457 1548 2473 1556
rect 2480 1554 2507 1556
rect 2516 1554 2737 1564
rect 2480 1544 2737 1554
rect 2766 1556 2816 1564
rect 2766 1547 2782 1556
rect 2375 1536 2426 1544
rect 2473 1536 2737 1544
rect 2763 1544 2782 1547
rect 2789 1544 2816 1556
rect 2763 1536 2816 1544
rect 2391 1528 2392 1536
rect 2407 1528 2420 1536
rect 2391 1520 2407 1528
rect 2388 1513 2407 1516
rect 2388 1504 2410 1513
rect 2361 1494 2410 1504
rect 2361 1488 2391 1494
rect 2410 1489 2415 1494
rect 2333 1472 2407 1488
rect 2425 1480 2455 1536
rect 2490 1526 2698 1536
rect 2733 1532 2778 1536
rect 2781 1535 2782 1536
rect 2797 1535 2810 1536
rect 2516 1496 2705 1526
rect 2531 1493 2705 1496
rect 2524 1490 2705 1493
rect 2333 1470 2346 1472
rect 2361 1470 2395 1472
rect 2333 1454 2407 1470
rect 2434 1466 2447 1480
rect 2462 1466 2478 1482
rect 2524 1477 2535 1490
rect 2317 1432 2318 1448
rect 2333 1432 2346 1454
rect 2361 1432 2391 1454
rect 2434 1450 2496 1466
rect 2524 1459 2535 1475
rect 2540 1470 2550 1490
rect 2560 1470 2574 1490
rect 2577 1477 2586 1490
rect 2602 1477 2611 1490
rect 2540 1459 2574 1470
rect 2577 1459 2586 1475
rect 2602 1459 2611 1475
rect 2618 1470 2628 1490
rect 2638 1470 2652 1490
rect 2653 1477 2664 1490
rect 2618 1459 2652 1470
rect 2653 1459 2664 1475
rect 2710 1466 2726 1482
rect 2733 1480 2763 1532
rect 2797 1528 2798 1535
rect 2782 1520 2798 1528
rect 2769 1488 2782 1507
rect 2797 1488 2827 1504
rect 2769 1472 2843 1488
rect 2769 1470 2782 1472
rect 2797 1470 2831 1472
rect 2434 1448 2447 1450
rect 2462 1448 2496 1450
rect 2434 1432 2496 1448
rect 2540 1443 2556 1446
rect 2618 1443 2648 1454
rect 2696 1450 2742 1466
rect 2769 1454 2843 1470
rect 2696 1448 2730 1450
rect 2695 1432 2742 1448
rect 2769 1432 2782 1454
rect 2797 1432 2827 1454
rect 2854 1432 2855 1448
rect 2870 1432 2883 1592
rect 2913 1488 2926 1592
rect 2971 1570 2972 1580
rect 2987 1570 3000 1580
rect 2971 1566 3000 1570
rect 3005 1566 3035 1592
rect 3053 1578 3069 1580
rect 3141 1578 3194 1592
rect 3142 1576 3206 1578
rect 3249 1576 3264 1592
rect 3313 1589 3343 1592
rect 3313 1586 3349 1589
rect 3279 1578 3295 1580
rect 3053 1566 3068 1570
rect 2971 1564 3068 1566
rect 3096 1564 3264 1576
rect 3280 1566 3295 1570
rect 3313 1567 3352 1586
rect 3371 1580 3378 1581
rect 3377 1573 3378 1580
rect 3361 1570 3362 1573
rect 3377 1570 3390 1573
rect 3313 1566 3343 1567
rect 3352 1566 3358 1567
rect 3361 1566 3390 1570
rect 3280 1565 3390 1566
rect 3280 1564 3396 1565
rect 2955 1556 3006 1564
rect 2955 1544 2980 1556
rect 2987 1544 3006 1556
rect 3037 1556 3087 1564
rect 3037 1548 3053 1556
rect 3060 1554 3087 1556
rect 3096 1554 3317 1564
rect 3060 1544 3317 1554
rect 3346 1556 3396 1564
rect 3346 1547 3362 1556
rect 2955 1536 3006 1544
rect 3053 1536 3317 1544
rect 3343 1544 3362 1547
rect 3369 1544 3396 1556
rect 3343 1536 3396 1544
rect 2971 1528 2972 1536
rect 2987 1528 3000 1536
rect 2971 1520 2987 1528
rect 2968 1513 2987 1516
rect 2968 1504 2990 1513
rect 2941 1494 2990 1504
rect 2941 1488 2971 1494
rect 2990 1489 2995 1494
rect 2913 1472 2987 1488
rect 3005 1480 3035 1536
rect 3070 1526 3278 1536
rect 3313 1532 3358 1536
rect 3361 1535 3362 1536
rect 3377 1535 3390 1536
rect 3096 1496 3285 1526
rect 3111 1493 3285 1496
rect 3104 1490 3285 1493
rect 2913 1470 2926 1472
rect 2941 1470 2975 1472
rect 2913 1454 2987 1470
rect 3014 1466 3027 1480
rect 3042 1466 3058 1482
rect 3104 1477 3115 1490
rect 2897 1432 2898 1448
rect 2913 1432 2926 1454
rect 2941 1432 2971 1454
rect 3014 1450 3076 1466
rect 3104 1459 3115 1475
rect 3120 1470 3130 1490
rect 3140 1470 3154 1490
rect 3157 1477 3166 1490
rect 3182 1477 3191 1490
rect 3120 1459 3154 1470
rect 3157 1459 3166 1475
rect 3182 1459 3191 1475
rect 3198 1470 3208 1490
rect 3218 1470 3232 1490
rect 3233 1477 3244 1490
rect 3198 1459 3232 1470
rect 3233 1459 3244 1475
rect 3290 1466 3306 1482
rect 3313 1480 3343 1532
rect 3377 1528 3378 1535
rect 3362 1520 3378 1528
rect 3349 1488 3362 1507
rect 3377 1488 3407 1504
rect 3349 1472 3423 1488
rect 3349 1470 3362 1472
rect 3377 1470 3411 1472
rect 3014 1448 3027 1450
rect 3042 1448 3076 1450
rect 3014 1432 3076 1448
rect 3120 1443 3136 1446
rect 3198 1443 3228 1454
rect 3276 1450 3322 1466
rect 3349 1454 3423 1470
rect 3276 1448 3310 1450
rect 3275 1432 3322 1448
rect 3349 1432 3362 1454
rect 3377 1432 3407 1454
rect 3434 1432 3435 1448
rect 3450 1432 3463 1592
rect 5911 1488 5924 1592
rect 5969 1570 5970 1580
rect 5985 1570 5998 1580
rect 5969 1566 5998 1570
rect 6003 1566 6033 1592
rect 6051 1578 6067 1580
rect 6139 1578 6192 1592
rect 6140 1576 6204 1578
rect 6247 1576 6262 1592
rect 6311 1589 6341 1592
rect 6311 1586 6347 1589
rect 6277 1578 6293 1580
rect 6051 1566 6066 1570
rect 5969 1564 6066 1566
rect 6094 1564 6262 1576
rect 6278 1566 6293 1570
rect 6311 1567 6350 1586
rect 6369 1580 6376 1581
rect 6375 1573 6376 1580
rect 6359 1570 6360 1573
rect 6375 1570 6388 1573
rect 6311 1566 6341 1567
rect 6350 1566 6356 1567
rect 6359 1566 6388 1570
rect 6278 1565 6388 1566
rect 6278 1564 6394 1565
rect 5953 1556 6004 1564
rect 5953 1544 5978 1556
rect 5985 1544 6004 1556
rect 6035 1556 6085 1564
rect 6035 1548 6051 1556
rect 6058 1554 6085 1556
rect 6094 1554 6315 1564
rect 6058 1544 6315 1554
rect 6344 1556 6394 1564
rect 6344 1547 6360 1556
rect 5953 1536 6004 1544
rect 6051 1536 6315 1544
rect 6341 1544 6360 1547
rect 6367 1544 6394 1556
rect 6341 1536 6394 1544
rect 5969 1528 5970 1536
rect 5985 1528 5998 1536
rect 5969 1520 5985 1528
rect 5966 1513 5985 1516
rect 5966 1504 5988 1513
rect 5939 1494 5988 1504
rect 5939 1488 5969 1494
rect 5988 1489 5993 1494
rect 5911 1472 5985 1488
rect 6003 1480 6033 1536
rect 6068 1526 6276 1536
rect 6311 1532 6356 1536
rect 6359 1535 6360 1536
rect 6375 1535 6388 1536
rect 6094 1496 6283 1526
rect 6109 1493 6283 1496
rect 6102 1490 6283 1493
rect 5911 1470 5924 1472
rect 5939 1470 5973 1472
rect 5911 1454 5985 1470
rect 6012 1466 6025 1480
rect 6040 1466 6056 1482
rect 6102 1477 6113 1490
rect 5895 1432 5896 1448
rect 5911 1432 5924 1454
rect 5939 1432 5969 1454
rect 6012 1450 6074 1466
rect 6102 1459 6113 1475
rect 6118 1470 6128 1490
rect 6138 1470 6152 1490
rect 6155 1477 6164 1490
rect 6180 1477 6189 1490
rect 6118 1459 6152 1470
rect 6155 1459 6164 1475
rect 6180 1459 6189 1475
rect 6196 1470 6206 1490
rect 6216 1470 6230 1490
rect 6231 1477 6242 1490
rect 6196 1459 6230 1470
rect 6231 1459 6242 1475
rect 6288 1466 6304 1482
rect 6311 1480 6341 1532
rect 6375 1528 6376 1535
rect 6360 1520 6376 1528
rect 6347 1488 6360 1507
rect 6375 1488 6405 1504
rect 6347 1472 6421 1488
rect 6347 1470 6360 1472
rect 6375 1470 6409 1472
rect 6012 1448 6025 1450
rect 6040 1448 6074 1450
rect 6012 1432 6074 1448
rect 6118 1443 6134 1446
rect 6196 1443 6226 1454
rect 6274 1450 6320 1466
rect 6347 1454 6421 1470
rect 6274 1448 6308 1450
rect 6273 1432 6320 1448
rect 6347 1432 6360 1454
rect 6375 1432 6405 1454
rect 6432 1432 6433 1448
rect 6448 1432 6461 1592
rect 6491 1488 6504 1592
rect 6549 1570 6550 1580
rect 6565 1570 6578 1580
rect 6549 1566 6578 1570
rect 6583 1566 6613 1592
rect 6631 1578 6647 1580
rect 6719 1578 6772 1592
rect 6720 1576 6784 1578
rect 6827 1576 6842 1592
rect 6891 1589 6921 1592
rect 6891 1586 6927 1589
rect 6857 1578 6873 1580
rect 6631 1566 6646 1570
rect 6549 1564 6646 1566
rect 6674 1564 6842 1576
rect 6858 1566 6873 1570
rect 6891 1567 6930 1586
rect 6949 1580 6956 1581
rect 6955 1573 6956 1580
rect 6939 1570 6940 1573
rect 6955 1570 6968 1573
rect 6891 1566 6921 1567
rect 6930 1566 6936 1567
rect 6939 1566 6968 1570
rect 6858 1565 6968 1566
rect 6858 1564 6974 1565
rect 6533 1556 6584 1564
rect 6533 1544 6558 1556
rect 6565 1544 6584 1556
rect 6615 1556 6665 1564
rect 6615 1548 6631 1556
rect 6638 1554 6665 1556
rect 6674 1554 6895 1564
rect 6638 1544 6895 1554
rect 6924 1556 6974 1564
rect 6924 1547 6940 1556
rect 6533 1536 6584 1544
rect 6631 1536 6895 1544
rect 6921 1544 6940 1547
rect 6947 1544 6974 1556
rect 6921 1536 6974 1544
rect 6549 1528 6550 1536
rect 6565 1528 6578 1536
rect 6549 1520 6565 1528
rect 6546 1513 6565 1516
rect 6546 1504 6568 1513
rect 6519 1494 6568 1504
rect 6519 1488 6549 1494
rect 6568 1489 6573 1494
rect 6491 1472 6565 1488
rect 6583 1480 6613 1536
rect 6648 1526 6856 1536
rect 6891 1532 6936 1536
rect 6939 1535 6940 1536
rect 6955 1535 6968 1536
rect 6674 1496 6863 1526
rect 6689 1493 6863 1496
rect 6682 1490 6863 1493
rect 6491 1470 6504 1472
rect 6519 1470 6553 1472
rect 6491 1454 6565 1470
rect 6592 1466 6605 1480
rect 6620 1466 6636 1482
rect 6682 1477 6693 1490
rect 6475 1432 6476 1448
rect 6491 1432 6504 1454
rect 6519 1432 6549 1454
rect 6592 1450 6654 1466
rect 6682 1459 6693 1475
rect 6698 1470 6708 1490
rect 6718 1470 6732 1490
rect 6735 1477 6744 1490
rect 6760 1477 6769 1490
rect 6698 1459 6732 1470
rect 6735 1459 6744 1475
rect 6760 1459 6769 1475
rect 6776 1470 6786 1490
rect 6796 1470 6810 1490
rect 6811 1477 6822 1490
rect 6776 1459 6810 1470
rect 6811 1459 6822 1475
rect 6868 1466 6884 1482
rect 6891 1480 6921 1532
rect 6955 1528 6956 1535
rect 6940 1520 6956 1528
rect 6927 1488 6940 1507
rect 6955 1488 6985 1504
rect 6927 1472 7001 1488
rect 6927 1470 6940 1472
rect 6955 1470 6989 1472
rect 6592 1448 6605 1450
rect 6620 1448 6654 1450
rect 6592 1432 6654 1448
rect 6698 1443 6714 1446
rect 6776 1443 6806 1454
rect 6854 1450 6900 1466
rect 6927 1454 7001 1470
rect 6854 1448 6888 1450
rect 6853 1432 6900 1448
rect 6927 1432 6940 1454
rect 6955 1432 6985 1454
rect 7012 1432 7013 1448
rect 7028 1432 7041 1592
rect 7071 1488 7084 1592
rect 7129 1570 7130 1580
rect 7145 1570 7158 1580
rect 7129 1566 7158 1570
rect 7163 1566 7193 1592
rect 7211 1578 7227 1580
rect 7299 1578 7352 1592
rect 7300 1576 7364 1578
rect 7407 1576 7422 1592
rect 7471 1589 7501 1592
rect 7471 1586 7507 1589
rect 7437 1578 7453 1580
rect 7211 1566 7226 1570
rect 7129 1564 7226 1566
rect 7254 1564 7422 1576
rect 7438 1566 7453 1570
rect 7471 1567 7510 1586
rect 7529 1580 7536 1581
rect 7535 1573 7536 1580
rect 7519 1570 7520 1573
rect 7535 1570 7548 1573
rect 7471 1566 7501 1567
rect 7510 1566 7516 1567
rect 7519 1566 7548 1570
rect 7438 1565 7548 1566
rect 7438 1564 7554 1565
rect 7113 1556 7164 1564
rect 7113 1544 7138 1556
rect 7145 1544 7164 1556
rect 7195 1556 7245 1564
rect 7195 1548 7211 1556
rect 7218 1554 7245 1556
rect 7254 1554 7475 1564
rect 7218 1544 7475 1554
rect 7504 1556 7554 1564
rect 7504 1547 7520 1556
rect 7113 1536 7164 1544
rect 7211 1536 7475 1544
rect 7501 1544 7520 1547
rect 7527 1544 7554 1556
rect 7501 1536 7554 1544
rect 7129 1528 7130 1536
rect 7145 1528 7158 1536
rect 7129 1520 7145 1528
rect 7126 1513 7145 1516
rect 7126 1504 7148 1513
rect 7099 1494 7148 1504
rect 7099 1488 7129 1494
rect 7148 1489 7153 1494
rect 7071 1472 7145 1488
rect 7163 1480 7193 1536
rect 7228 1526 7436 1536
rect 7471 1532 7516 1536
rect 7519 1535 7520 1536
rect 7535 1535 7548 1536
rect 7254 1496 7443 1526
rect 7269 1493 7443 1496
rect 7262 1490 7443 1493
rect 7071 1470 7084 1472
rect 7099 1470 7133 1472
rect 7071 1454 7145 1470
rect 7172 1466 7185 1480
rect 7200 1466 7216 1482
rect 7262 1477 7273 1490
rect 7055 1432 7056 1448
rect 7071 1432 7084 1454
rect 7099 1432 7129 1454
rect 7172 1450 7234 1466
rect 7262 1459 7273 1475
rect 7278 1470 7288 1490
rect 7298 1470 7312 1490
rect 7315 1477 7324 1490
rect 7340 1477 7349 1490
rect 7278 1459 7312 1470
rect 7315 1459 7324 1475
rect 7340 1459 7349 1475
rect 7356 1470 7366 1490
rect 7376 1470 7390 1490
rect 7391 1477 7402 1490
rect 7356 1459 7390 1470
rect 7391 1459 7402 1475
rect 7448 1466 7464 1482
rect 7471 1480 7501 1532
rect 7535 1528 7536 1535
rect 7520 1520 7536 1528
rect 7507 1488 7520 1507
rect 7535 1488 7565 1504
rect 7507 1472 7581 1488
rect 7507 1470 7520 1472
rect 7535 1470 7569 1472
rect 7172 1448 7185 1450
rect 7200 1448 7234 1450
rect 7172 1432 7234 1448
rect 7278 1443 7294 1446
rect 7356 1443 7386 1454
rect 7434 1450 7480 1466
rect 7507 1454 7581 1470
rect 7434 1448 7468 1450
rect 7433 1432 7480 1448
rect 7507 1432 7520 1454
rect 7535 1432 7565 1454
rect 7592 1432 7593 1448
rect 7608 1432 7621 1592
rect 7651 1488 7664 1592
rect 7709 1570 7710 1580
rect 7725 1570 7738 1580
rect 7709 1566 7738 1570
rect 7743 1566 7773 1592
rect 7791 1578 7807 1580
rect 7879 1578 7932 1592
rect 7880 1576 7944 1578
rect 7987 1576 8002 1592
rect 8051 1589 8081 1592
rect 8051 1586 8087 1589
rect 8017 1578 8033 1580
rect 7791 1566 7806 1570
rect 7709 1564 7806 1566
rect 7834 1564 8002 1576
rect 8018 1566 8033 1570
rect 8051 1567 8090 1586
rect 8109 1580 8116 1581
rect 8115 1573 8116 1580
rect 8099 1570 8100 1573
rect 8115 1570 8128 1573
rect 8051 1566 8081 1567
rect 8090 1566 8096 1567
rect 8099 1566 8128 1570
rect 8018 1565 8128 1566
rect 8018 1564 8134 1565
rect 7693 1556 7744 1564
rect 7693 1544 7718 1556
rect 7725 1544 7744 1556
rect 7775 1556 7825 1564
rect 7775 1548 7791 1556
rect 7798 1554 7825 1556
rect 7834 1554 8055 1564
rect 7798 1544 8055 1554
rect 8084 1556 8134 1564
rect 8084 1547 8100 1556
rect 7693 1536 7744 1544
rect 7791 1536 8055 1544
rect 8081 1544 8100 1547
rect 8107 1544 8134 1556
rect 8081 1536 8134 1544
rect 7709 1528 7710 1536
rect 7725 1528 7738 1536
rect 7709 1520 7725 1528
rect 7706 1513 7725 1516
rect 7706 1504 7728 1513
rect 7679 1494 7728 1504
rect 7679 1488 7709 1494
rect 7728 1489 7733 1494
rect 7651 1472 7725 1488
rect 7743 1480 7773 1536
rect 7808 1526 8016 1536
rect 8051 1532 8096 1536
rect 8099 1535 8100 1536
rect 8115 1535 8128 1536
rect 7834 1496 8023 1526
rect 7849 1493 8023 1496
rect 7842 1490 8023 1493
rect 7651 1470 7664 1472
rect 7679 1470 7713 1472
rect 7651 1454 7725 1470
rect 7752 1466 7765 1480
rect 7780 1466 7796 1482
rect 7842 1477 7853 1490
rect 7635 1432 7636 1448
rect 7651 1432 7664 1454
rect 7679 1432 7709 1454
rect 7752 1450 7814 1466
rect 7842 1459 7853 1475
rect 7858 1470 7868 1490
rect 7878 1470 7892 1490
rect 7895 1477 7904 1490
rect 7920 1477 7929 1490
rect 7858 1459 7892 1470
rect 7895 1459 7904 1475
rect 7920 1459 7929 1475
rect 7936 1470 7946 1490
rect 7956 1470 7970 1490
rect 7971 1477 7982 1490
rect 7936 1459 7970 1470
rect 7971 1459 7982 1475
rect 8028 1466 8044 1482
rect 8051 1480 8081 1532
rect 8115 1528 8116 1535
rect 8100 1520 8116 1528
rect 8087 1488 8100 1507
rect 8115 1488 8145 1504
rect 8087 1472 8161 1488
rect 8087 1470 8100 1472
rect 8115 1470 8149 1472
rect 7752 1448 7765 1450
rect 7780 1448 7814 1450
rect 7752 1432 7814 1448
rect 7858 1443 7874 1446
rect 7936 1443 7966 1454
rect 8014 1450 8060 1466
rect 8087 1454 8161 1470
rect 8014 1448 8048 1450
rect 8013 1432 8060 1448
rect 8087 1432 8100 1454
rect 8115 1432 8145 1454
rect 8172 1432 8173 1448
rect 8188 1432 8201 1592
rect 8231 1488 8244 1592
rect 8289 1570 8290 1580
rect 8305 1570 8318 1580
rect 8289 1566 8318 1570
rect 8323 1566 8353 1592
rect 8371 1578 8387 1580
rect 8459 1578 8512 1592
rect 8460 1576 8524 1578
rect 8567 1576 8582 1592
rect 8631 1589 8661 1592
rect 8631 1586 8667 1589
rect 8597 1578 8613 1580
rect 8371 1566 8386 1570
rect 8289 1564 8386 1566
rect 8414 1564 8582 1576
rect 8598 1566 8613 1570
rect 8631 1567 8670 1586
rect 8689 1580 8696 1581
rect 8695 1573 8696 1580
rect 8679 1570 8680 1573
rect 8695 1570 8708 1573
rect 8631 1566 8661 1567
rect 8670 1566 8676 1567
rect 8679 1566 8708 1570
rect 8598 1565 8708 1566
rect 8598 1564 8714 1565
rect 8273 1556 8324 1564
rect 8273 1544 8298 1556
rect 8305 1544 8324 1556
rect 8355 1556 8405 1564
rect 8355 1548 8371 1556
rect 8378 1554 8405 1556
rect 8414 1554 8635 1564
rect 8378 1544 8635 1554
rect 8664 1556 8714 1564
rect 8664 1547 8680 1556
rect 8273 1536 8324 1544
rect 8371 1536 8635 1544
rect 8661 1544 8680 1547
rect 8687 1544 8714 1556
rect 8661 1536 8714 1544
rect 8289 1528 8290 1536
rect 8305 1528 8318 1536
rect 8289 1520 8305 1528
rect 8286 1513 8305 1516
rect 8286 1504 8308 1513
rect 8259 1494 8308 1504
rect 8259 1488 8289 1494
rect 8308 1489 8313 1494
rect 8231 1472 8305 1488
rect 8323 1480 8353 1536
rect 8388 1526 8596 1536
rect 8631 1532 8676 1536
rect 8679 1535 8680 1536
rect 8695 1535 8708 1536
rect 8414 1496 8603 1526
rect 8429 1493 8603 1496
rect 8422 1490 8603 1493
rect 8231 1470 8244 1472
rect 8259 1470 8293 1472
rect 8231 1454 8305 1470
rect 8332 1466 8345 1480
rect 8360 1466 8376 1482
rect 8422 1477 8433 1490
rect 8215 1432 8216 1448
rect 8231 1432 8244 1454
rect 8259 1432 8289 1454
rect 8332 1450 8394 1466
rect 8422 1459 8433 1475
rect 8438 1470 8448 1490
rect 8458 1470 8472 1490
rect 8475 1477 8484 1490
rect 8500 1477 8509 1490
rect 8438 1459 8472 1470
rect 8475 1459 8484 1475
rect 8500 1459 8509 1475
rect 8516 1470 8526 1490
rect 8536 1470 8550 1490
rect 8551 1477 8562 1490
rect 8516 1459 8550 1470
rect 8551 1459 8562 1475
rect 8608 1466 8624 1482
rect 8631 1480 8661 1532
rect 8695 1528 8696 1535
rect 8680 1520 8696 1528
rect 8667 1488 8680 1507
rect 8695 1488 8725 1504
rect 8667 1472 8741 1488
rect 8667 1470 8680 1472
rect 8695 1470 8729 1472
rect 8332 1448 8345 1450
rect 8360 1448 8394 1450
rect 8332 1432 8394 1448
rect 8438 1443 8454 1446
rect 8516 1443 8546 1454
rect 8594 1450 8640 1466
rect 8667 1454 8741 1470
rect 8594 1448 8628 1450
rect 8593 1432 8640 1448
rect 8667 1432 8680 1454
rect 8695 1432 8725 1454
rect 8752 1432 8753 1448
rect 8768 1432 8781 1592
rect 8811 1488 8824 1592
rect 8869 1570 8870 1580
rect 8885 1570 8898 1580
rect 8869 1566 8898 1570
rect 8903 1566 8933 1592
rect 8951 1578 8967 1580
rect 9039 1578 9092 1592
rect 9040 1576 9104 1578
rect 9147 1576 9162 1592
rect 9211 1589 9241 1592
rect 9211 1586 9247 1589
rect 9177 1578 9193 1580
rect 8951 1566 8966 1570
rect 8869 1564 8966 1566
rect 8994 1564 9162 1576
rect 9178 1566 9193 1570
rect 9211 1567 9250 1586
rect 9269 1580 9276 1581
rect 9275 1573 9276 1580
rect 9259 1570 9260 1573
rect 9275 1570 9288 1573
rect 9211 1566 9241 1567
rect 9250 1566 9256 1567
rect 9259 1566 9288 1570
rect 9178 1565 9288 1566
rect 9178 1564 9294 1565
rect 8853 1556 8904 1564
rect 8853 1544 8878 1556
rect 8885 1544 8904 1556
rect 8935 1556 8985 1564
rect 8935 1548 8951 1556
rect 8958 1554 8985 1556
rect 8994 1554 9215 1564
rect 8958 1544 9215 1554
rect 9244 1556 9294 1564
rect 9244 1547 9260 1556
rect 8853 1536 8904 1544
rect 8951 1536 9215 1544
rect 9241 1544 9260 1547
rect 9267 1544 9294 1556
rect 9241 1536 9294 1544
rect 8869 1528 8870 1536
rect 8885 1528 8898 1536
rect 8869 1520 8885 1528
rect 8866 1513 8885 1516
rect 8866 1504 8888 1513
rect 8839 1494 8888 1504
rect 8839 1488 8869 1494
rect 8888 1489 8893 1494
rect 8811 1472 8885 1488
rect 8903 1480 8933 1536
rect 8968 1526 9176 1536
rect 9211 1532 9256 1536
rect 9259 1535 9260 1536
rect 9275 1535 9288 1536
rect 8994 1496 9183 1526
rect 9009 1493 9183 1496
rect 9002 1490 9183 1493
rect 8811 1470 8824 1472
rect 8839 1470 8873 1472
rect 8811 1454 8885 1470
rect 8912 1466 8925 1480
rect 8940 1466 8956 1482
rect 9002 1477 9013 1490
rect 8795 1432 8796 1448
rect 8811 1432 8824 1454
rect 8839 1432 8869 1454
rect 8912 1450 8974 1466
rect 9002 1459 9013 1475
rect 9018 1470 9028 1490
rect 9038 1470 9052 1490
rect 9055 1477 9064 1490
rect 9080 1477 9089 1490
rect 9018 1459 9052 1470
rect 9055 1459 9064 1475
rect 9080 1459 9089 1475
rect 9096 1470 9106 1490
rect 9116 1470 9130 1490
rect 9131 1477 9142 1490
rect 9096 1459 9130 1470
rect 9131 1459 9142 1475
rect 9188 1466 9204 1482
rect 9211 1480 9241 1532
rect 9275 1528 9276 1535
rect 9260 1520 9276 1528
rect 9247 1488 9260 1507
rect 9275 1488 9305 1504
rect 9247 1472 9321 1488
rect 9247 1470 9260 1472
rect 9275 1470 9309 1472
rect 8912 1448 8925 1450
rect 8940 1448 8974 1450
rect 8912 1432 8974 1448
rect 9018 1443 9034 1446
rect 9096 1443 9126 1454
rect 9174 1450 9220 1466
rect 9247 1454 9321 1470
rect 9174 1448 9208 1450
rect 9173 1432 9220 1448
rect 9247 1432 9260 1454
rect 9275 1432 9305 1454
rect 9332 1432 9333 1448
rect 9348 1432 9361 1592
rect -9 1424 32 1432
rect -9 1398 6 1424
rect 13 1398 32 1424
rect 96 1420 158 1432
rect 170 1420 245 1432
rect 303 1420 378 1432
rect 390 1420 421 1432
rect 427 1420 462 1432
rect 96 1418 258 1420
rect -9 1390 32 1398
rect 114 1394 127 1418
rect 142 1416 157 1418
rect -3 1380 -2 1390
rect 13 1380 26 1390
rect 41 1380 71 1394
rect 114 1380 157 1394
rect 181 1391 188 1398
rect 191 1394 258 1418
rect 290 1418 462 1420
rect 260 1396 288 1400
rect 290 1396 370 1418
rect 391 1416 406 1418
rect 260 1394 370 1396
rect 191 1390 370 1394
rect 164 1380 194 1390
rect 196 1380 349 1390
rect 357 1380 387 1390
rect 391 1380 421 1394
rect 449 1380 462 1418
rect 534 1424 569 1432
rect 534 1398 535 1424
rect 542 1398 569 1424
rect 477 1380 507 1394
rect 534 1390 569 1398
rect 571 1424 612 1432
rect 571 1398 586 1424
rect 593 1398 612 1424
rect 676 1420 738 1432
rect 750 1420 825 1432
rect 883 1420 958 1432
rect 970 1420 1001 1432
rect 1007 1420 1042 1432
rect 676 1418 838 1420
rect 571 1390 612 1398
rect 694 1394 707 1418
rect 722 1416 737 1418
rect 534 1380 535 1390
rect 550 1380 563 1390
rect 577 1380 578 1390
rect 593 1380 606 1390
rect 621 1380 651 1394
rect 694 1380 737 1394
rect 761 1391 768 1398
rect 771 1394 838 1418
rect 870 1418 1042 1420
rect 840 1396 868 1400
rect 870 1396 950 1418
rect 971 1416 986 1418
rect 840 1394 950 1396
rect 771 1390 950 1394
rect 744 1380 774 1390
rect 776 1380 929 1390
rect 937 1380 967 1390
rect 971 1380 1001 1394
rect 1029 1380 1042 1418
rect 1114 1424 1149 1432
rect 1114 1398 1115 1424
rect 1122 1398 1149 1424
rect 1057 1380 1087 1394
rect 1114 1390 1149 1398
rect 1151 1424 1192 1432
rect 1151 1398 1166 1424
rect 1173 1398 1192 1424
rect 1256 1420 1318 1432
rect 1330 1420 1405 1432
rect 1463 1420 1538 1432
rect 1550 1420 1581 1432
rect 1587 1420 1622 1432
rect 1256 1418 1418 1420
rect 1151 1390 1192 1398
rect 1274 1394 1287 1418
rect 1302 1416 1317 1418
rect 1114 1380 1115 1390
rect 1130 1380 1143 1390
rect 1157 1380 1158 1390
rect 1173 1380 1186 1390
rect 1201 1380 1231 1394
rect 1274 1380 1317 1394
rect 1341 1391 1348 1398
rect 1351 1394 1418 1418
rect 1450 1418 1622 1420
rect 1420 1396 1448 1400
rect 1450 1396 1530 1418
rect 1551 1416 1566 1418
rect 1420 1394 1530 1396
rect 1351 1390 1530 1394
rect 1324 1380 1354 1390
rect 1356 1380 1509 1390
rect 1517 1380 1547 1390
rect 1551 1380 1581 1394
rect 1609 1380 1622 1418
rect 1694 1424 1729 1432
rect 1694 1398 1695 1424
rect 1702 1398 1729 1424
rect 1637 1380 1667 1394
rect 1694 1390 1729 1398
rect 1731 1424 1772 1432
rect 1731 1398 1746 1424
rect 1753 1398 1772 1424
rect 1836 1420 1898 1432
rect 1910 1420 1985 1432
rect 2043 1420 2118 1432
rect 2130 1420 2161 1432
rect 2167 1420 2202 1432
rect 1836 1418 1998 1420
rect 1731 1390 1772 1398
rect 1854 1394 1867 1418
rect 1882 1416 1897 1418
rect 1694 1380 1695 1390
rect 1710 1380 1723 1390
rect 1737 1380 1738 1390
rect 1753 1380 1766 1390
rect 1781 1380 1811 1394
rect 1854 1380 1897 1394
rect 1921 1391 1928 1398
rect 1931 1394 1998 1418
rect 2030 1418 2202 1420
rect 2000 1396 2028 1400
rect 2030 1396 2110 1418
rect 2131 1416 2146 1418
rect 2000 1394 2110 1396
rect 1931 1390 2110 1394
rect 1904 1380 1934 1390
rect 1936 1380 2089 1390
rect 2097 1380 2127 1390
rect 2131 1380 2161 1394
rect 2189 1380 2202 1418
rect 2274 1424 2309 1432
rect 2274 1398 2275 1424
rect 2282 1398 2309 1424
rect 2217 1380 2247 1394
rect 2274 1390 2309 1398
rect 2311 1424 2352 1432
rect 2311 1398 2326 1424
rect 2333 1398 2352 1424
rect 2416 1420 2478 1432
rect 2490 1420 2565 1432
rect 2623 1420 2698 1432
rect 2710 1420 2741 1432
rect 2747 1420 2782 1432
rect 2416 1418 2578 1420
rect 2311 1390 2352 1398
rect 2434 1394 2447 1418
rect 2462 1416 2477 1418
rect 2274 1380 2275 1390
rect 2290 1380 2303 1390
rect 2317 1380 2318 1390
rect 2333 1380 2346 1390
rect 2361 1380 2391 1394
rect 2434 1380 2477 1394
rect 2501 1391 2508 1398
rect 2511 1394 2578 1418
rect 2610 1418 2782 1420
rect 2580 1396 2608 1400
rect 2610 1396 2690 1418
rect 2711 1416 2726 1418
rect 2580 1394 2690 1396
rect 2511 1390 2690 1394
rect 2484 1380 2514 1390
rect 2516 1380 2669 1390
rect 2677 1380 2707 1390
rect 2711 1380 2741 1394
rect 2769 1380 2782 1418
rect 2854 1424 2889 1432
rect 2854 1398 2855 1424
rect 2862 1398 2889 1424
rect 2797 1380 2827 1394
rect 2854 1390 2889 1398
rect 2891 1424 2932 1432
rect 2891 1398 2906 1424
rect 2913 1398 2932 1424
rect 2996 1420 3058 1432
rect 3070 1420 3145 1432
rect 3203 1420 3278 1432
rect 3290 1420 3321 1432
rect 3327 1420 3362 1432
rect 2996 1418 3158 1420
rect 2891 1390 2932 1398
rect 3014 1394 3027 1418
rect 3042 1416 3057 1418
rect 2854 1380 2855 1390
rect 2870 1380 2883 1390
rect 2897 1380 2898 1390
rect 2913 1380 2926 1390
rect 2941 1380 2971 1394
rect 3014 1380 3057 1394
rect 3081 1391 3088 1398
rect 3091 1394 3158 1418
rect 3190 1418 3362 1420
rect 3160 1396 3188 1400
rect 3190 1396 3270 1418
rect 3291 1416 3306 1418
rect 3160 1394 3270 1396
rect 3091 1390 3270 1394
rect 3064 1380 3094 1390
rect 3096 1380 3249 1390
rect 3257 1380 3287 1390
rect 3291 1380 3321 1394
rect 3349 1380 3362 1418
rect 3434 1424 3469 1432
rect 3434 1398 3435 1424
rect 3442 1398 3469 1424
rect 3377 1380 3407 1394
rect 3434 1390 3469 1398
rect 3434 1380 3435 1390
rect 3450 1380 3463 1390
rect -3 1374 3469 1380
rect -2 1366 3469 1374
rect 5889 1424 5930 1432
rect 5889 1398 5904 1424
rect 5911 1398 5930 1424
rect 5994 1420 6056 1432
rect 6068 1420 6143 1432
rect 6201 1420 6276 1432
rect 6288 1420 6319 1432
rect 6325 1420 6360 1432
rect 5994 1418 6156 1420
rect 5889 1390 5930 1398
rect 6012 1394 6025 1418
rect 6040 1416 6055 1418
rect 5895 1380 5896 1390
rect 5911 1380 5924 1390
rect 5939 1380 5969 1394
rect 6012 1380 6055 1394
rect 6079 1391 6086 1398
rect 6089 1394 6156 1418
rect 6188 1418 6360 1420
rect 6158 1396 6186 1400
rect 6188 1396 6268 1418
rect 6289 1416 6304 1418
rect 6158 1394 6268 1396
rect 6089 1390 6268 1394
rect 6062 1380 6092 1390
rect 6094 1380 6247 1390
rect 6255 1380 6285 1390
rect 6289 1380 6319 1394
rect 6347 1380 6360 1418
rect 6432 1424 6467 1432
rect 6432 1398 6433 1424
rect 6440 1398 6467 1424
rect 6375 1380 6405 1394
rect 6432 1390 6467 1398
rect 6469 1424 6510 1432
rect 6469 1398 6484 1424
rect 6491 1398 6510 1424
rect 6574 1420 6636 1432
rect 6648 1420 6723 1432
rect 6781 1420 6856 1432
rect 6868 1420 6899 1432
rect 6905 1420 6940 1432
rect 6574 1418 6736 1420
rect 6469 1390 6510 1398
rect 6592 1394 6605 1418
rect 6620 1416 6635 1418
rect 6432 1380 6433 1390
rect 6448 1380 6461 1390
rect 6475 1380 6476 1390
rect 6491 1380 6504 1390
rect 6519 1380 6549 1394
rect 6592 1380 6635 1394
rect 6659 1391 6666 1398
rect 6669 1394 6736 1418
rect 6768 1418 6940 1420
rect 6738 1396 6766 1400
rect 6768 1396 6848 1418
rect 6869 1416 6884 1418
rect 6738 1394 6848 1396
rect 6669 1390 6848 1394
rect 6642 1380 6672 1390
rect 6674 1380 6827 1390
rect 6835 1380 6865 1390
rect 6869 1380 6899 1394
rect 6927 1380 6940 1418
rect 7012 1424 7047 1432
rect 7012 1398 7013 1424
rect 7020 1398 7047 1424
rect 6955 1380 6985 1394
rect 7012 1390 7047 1398
rect 7049 1424 7090 1432
rect 7049 1398 7064 1424
rect 7071 1398 7090 1424
rect 7154 1420 7216 1432
rect 7228 1420 7303 1432
rect 7361 1420 7436 1432
rect 7448 1420 7479 1432
rect 7485 1420 7520 1432
rect 7154 1418 7316 1420
rect 7049 1390 7090 1398
rect 7172 1394 7185 1418
rect 7200 1416 7215 1418
rect 7012 1380 7013 1390
rect 7028 1380 7041 1390
rect 7055 1380 7056 1390
rect 7071 1380 7084 1390
rect 7099 1380 7129 1394
rect 7172 1380 7215 1394
rect 7239 1391 7246 1398
rect 7249 1394 7316 1418
rect 7348 1418 7520 1420
rect 7318 1396 7346 1400
rect 7348 1396 7428 1418
rect 7449 1416 7464 1418
rect 7318 1394 7428 1396
rect 7249 1390 7428 1394
rect 7222 1380 7252 1390
rect 7254 1380 7407 1390
rect 7415 1380 7445 1390
rect 7449 1380 7479 1394
rect 7507 1380 7520 1418
rect 7592 1424 7627 1432
rect 7592 1398 7593 1424
rect 7600 1398 7627 1424
rect 7535 1380 7565 1394
rect 7592 1390 7627 1398
rect 7629 1424 7670 1432
rect 7629 1398 7644 1424
rect 7651 1398 7670 1424
rect 7734 1420 7796 1432
rect 7808 1420 7883 1432
rect 7941 1420 8016 1432
rect 8028 1420 8059 1432
rect 8065 1420 8100 1432
rect 7734 1418 7896 1420
rect 7629 1390 7670 1398
rect 7752 1394 7765 1418
rect 7780 1416 7795 1418
rect 7592 1380 7593 1390
rect 7608 1380 7621 1390
rect 7635 1380 7636 1390
rect 7651 1380 7664 1390
rect 7679 1380 7709 1394
rect 7752 1380 7795 1394
rect 7819 1391 7826 1398
rect 7829 1394 7896 1418
rect 7928 1418 8100 1420
rect 7898 1396 7926 1400
rect 7928 1396 8008 1418
rect 8029 1416 8044 1418
rect 7898 1394 8008 1396
rect 7829 1390 8008 1394
rect 7802 1380 7832 1390
rect 7834 1380 7987 1390
rect 7995 1380 8025 1390
rect 8029 1380 8059 1394
rect 8087 1380 8100 1418
rect 8172 1424 8207 1432
rect 8172 1398 8173 1424
rect 8180 1398 8207 1424
rect 8115 1380 8145 1394
rect 8172 1390 8207 1398
rect 8209 1424 8250 1432
rect 8209 1398 8224 1424
rect 8231 1398 8250 1424
rect 8314 1420 8376 1432
rect 8388 1420 8463 1432
rect 8521 1420 8596 1432
rect 8608 1420 8639 1432
rect 8645 1420 8680 1432
rect 8314 1418 8476 1420
rect 8209 1390 8250 1398
rect 8332 1394 8345 1418
rect 8360 1416 8375 1418
rect 8172 1380 8173 1390
rect 8188 1380 8201 1390
rect 8215 1380 8216 1390
rect 8231 1380 8244 1390
rect 8259 1380 8289 1394
rect 8332 1380 8375 1394
rect 8399 1391 8406 1398
rect 8409 1394 8476 1418
rect 8508 1418 8680 1420
rect 8478 1396 8506 1400
rect 8508 1396 8588 1418
rect 8609 1416 8624 1418
rect 8478 1394 8588 1396
rect 8409 1390 8588 1394
rect 8382 1380 8412 1390
rect 8414 1380 8567 1390
rect 8575 1380 8605 1390
rect 8609 1380 8639 1394
rect 8667 1380 8680 1418
rect 8752 1424 8787 1432
rect 8752 1398 8753 1424
rect 8760 1398 8787 1424
rect 8695 1380 8725 1394
rect 8752 1390 8787 1398
rect 8789 1424 8830 1432
rect 8789 1398 8804 1424
rect 8811 1398 8830 1424
rect 8894 1420 8956 1432
rect 8968 1420 9043 1432
rect 9101 1420 9176 1432
rect 9188 1420 9219 1432
rect 9225 1420 9260 1432
rect 8894 1418 9056 1420
rect 8789 1390 8830 1398
rect 8912 1394 8925 1418
rect 8940 1416 8955 1418
rect 8752 1380 8753 1390
rect 8768 1380 8781 1390
rect 8795 1380 8796 1390
rect 8811 1380 8824 1390
rect 8839 1380 8869 1394
rect 8912 1380 8955 1394
rect 8979 1391 8986 1398
rect 8989 1394 9056 1418
rect 9088 1418 9260 1420
rect 9058 1396 9086 1400
rect 9088 1396 9168 1418
rect 9189 1416 9204 1418
rect 9058 1394 9168 1396
rect 8989 1390 9168 1394
rect 8962 1380 8992 1390
rect 8994 1380 9147 1390
rect 9155 1380 9185 1390
rect 9189 1380 9219 1394
rect 9247 1380 9260 1418
rect 9332 1424 9367 1432
rect 9332 1398 9333 1424
rect 9340 1398 9367 1424
rect 9275 1380 9305 1394
rect 9332 1390 9367 1398
rect 9332 1380 9333 1390
rect 9348 1380 9361 1390
rect 5889 1366 9361 1380
rect 13 1336 26 1366
rect 41 1348 71 1366
rect 114 1352 128 1366
rect 164 1352 384 1366
rect 115 1350 128 1352
rect 81 1338 96 1350
rect 78 1336 100 1338
rect 105 1336 135 1350
rect 196 1348 349 1352
rect 178 1336 370 1348
rect 413 1336 443 1350
rect 449 1336 462 1366
rect 477 1348 507 1366
rect 550 1336 563 1366
rect 593 1336 606 1366
rect 621 1348 651 1366
rect 694 1352 708 1366
rect 744 1352 964 1366
rect 695 1350 708 1352
rect 661 1338 676 1350
rect 658 1336 680 1338
rect 685 1336 715 1350
rect 776 1348 929 1352
rect 758 1336 950 1348
rect 993 1336 1023 1350
rect 1029 1336 1042 1366
rect 1057 1348 1087 1366
rect 1130 1336 1143 1366
rect 1173 1336 1186 1366
rect 1201 1348 1231 1366
rect 1274 1352 1288 1366
rect 1324 1352 1544 1366
rect 1275 1350 1288 1352
rect 1241 1338 1256 1350
rect 1238 1336 1260 1338
rect 1265 1336 1295 1350
rect 1356 1348 1509 1352
rect 1338 1336 1530 1348
rect 1573 1336 1603 1350
rect 1609 1336 1622 1366
rect 1637 1348 1667 1366
rect 1710 1336 1723 1366
rect 1753 1336 1766 1366
rect 1781 1348 1811 1366
rect 1854 1352 1868 1366
rect 1904 1352 2124 1366
rect 1855 1350 1868 1352
rect 1821 1338 1836 1350
rect 1818 1336 1840 1338
rect 1845 1336 1875 1350
rect 1936 1348 2089 1352
rect 1918 1336 2110 1348
rect 2153 1336 2183 1350
rect 2189 1336 2202 1366
rect 2217 1348 2247 1366
rect 2290 1336 2303 1366
rect 2333 1336 2346 1366
rect 2361 1348 2391 1366
rect 2434 1352 2448 1366
rect 2484 1352 2704 1366
rect 2435 1350 2448 1352
rect 2401 1338 2416 1350
rect 2398 1336 2420 1338
rect 2425 1336 2455 1350
rect 2516 1348 2669 1352
rect 2498 1336 2690 1348
rect 2733 1336 2763 1350
rect 2769 1336 2782 1366
rect 2797 1348 2827 1366
rect 2870 1336 2883 1366
rect 2913 1336 2926 1366
rect 2941 1348 2971 1366
rect 3014 1352 3028 1366
rect 3064 1352 3284 1366
rect 3015 1350 3028 1352
rect 2981 1338 2996 1350
rect 2978 1336 3000 1338
rect 3005 1336 3035 1350
rect 3096 1348 3249 1352
rect 3078 1336 3270 1348
rect 3313 1336 3343 1350
rect 3349 1336 3362 1366
rect 3377 1348 3407 1366
rect 3450 1336 3463 1366
rect 5911 1336 5924 1366
rect 5939 1348 5969 1366
rect 6012 1352 6026 1366
rect 6062 1352 6282 1366
rect 6013 1350 6026 1352
rect 5979 1338 5994 1350
rect 5976 1336 5998 1338
rect 6003 1336 6033 1350
rect 6094 1348 6247 1352
rect 6076 1336 6268 1348
rect 6311 1336 6341 1350
rect 6347 1336 6360 1366
rect 6375 1348 6405 1366
rect 6448 1336 6461 1366
rect 6491 1336 6504 1366
rect 6519 1348 6549 1366
rect 6592 1352 6606 1366
rect 6642 1352 6862 1366
rect 6593 1350 6606 1352
rect 6559 1338 6574 1350
rect 6556 1336 6578 1338
rect 6583 1336 6613 1350
rect 6674 1348 6827 1352
rect 6656 1336 6848 1348
rect 6891 1336 6921 1350
rect 6927 1336 6940 1366
rect 6955 1348 6985 1366
rect 7028 1336 7041 1366
rect 7071 1336 7084 1366
rect 7099 1348 7129 1366
rect 7172 1352 7186 1366
rect 7222 1352 7442 1366
rect 7173 1350 7186 1352
rect 7139 1338 7154 1350
rect 7136 1336 7158 1338
rect 7163 1336 7193 1350
rect 7254 1348 7407 1352
rect 7236 1336 7428 1348
rect 7471 1336 7501 1350
rect 7507 1336 7520 1366
rect 7535 1348 7565 1366
rect 7608 1336 7621 1366
rect 7651 1336 7664 1366
rect 7679 1348 7709 1366
rect 7752 1352 7766 1366
rect 7802 1352 8022 1366
rect 7753 1350 7766 1352
rect 7719 1338 7734 1350
rect 7716 1336 7738 1338
rect 7743 1336 7773 1350
rect 7834 1348 7987 1352
rect 7816 1336 8008 1348
rect 8051 1336 8081 1350
rect 8087 1336 8100 1366
rect 8115 1348 8145 1366
rect 8188 1336 8201 1366
rect 8231 1336 8244 1366
rect 8259 1348 8289 1366
rect 8332 1352 8346 1366
rect 8382 1352 8602 1366
rect 8333 1350 8346 1352
rect 8299 1338 8314 1350
rect 8296 1336 8318 1338
rect 8323 1336 8353 1350
rect 8414 1348 8567 1352
rect 8396 1336 8588 1348
rect 8631 1336 8661 1350
rect 8667 1336 8680 1366
rect 8695 1348 8725 1366
rect 8768 1336 8781 1366
rect 8811 1336 8824 1366
rect 8839 1348 8869 1366
rect 8912 1352 8926 1366
rect 8962 1352 9182 1366
rect 8913 1350 8926 1352
rect 8879 1338 8894 1350
rect 8876 1336 8898 1338
rect 8903 1336 8933 1350
rect 8994 1348 9147 1352
rect 8976 1336 9168 1348
rect 9211 1336 9241 1350
rect 9247 1336 9260 1366
rect 9275 1348 9305 1366
rect 9348 1336 9361 1366
rect -2 1322 3469 1336
rect 5889 1322 9361 1336
rect 13 1218 26 1322
rect 71 1300 72 1310
rect 87 1300 100 1310
rect 71 1296 100 1300
rect 105 1296 135 1322
rect 153 1308 169 1310
rect 241 1308 294 1322
rect 242 1306 306 1308
rect 349 1306 364 1322
rect 413 1319 443 1322
rect 413 1316 449 1319
rect 379 1308 395 1310
rect 153 1296 168 1300
rect 71 1294 168 1296
rect 196 1294 364 1306
rect 380 1296 395 1300
rect 413 1297 452 1316
rect 471 1310 478 1311
rect 477 1303 478 1310
rect 461 1300 462 1303
rect 477 1300 490 1303
rect 413 1296 443 1297
rect 452 1296 458 1297
rect 461 1296 490 1300
rect 380 1295 490 1296
rect 380 1294 496 1295
rect 55 1286 106 1294
rect 55 1274 80 1286
rect 87 1274 106 1286
rect 137 1286 187 1294
rect 137 1278 153 1286
rect 160 1284 187 1286
rect 196 1284 417 1294
rect 160 1274 417 1284
rect 446 1286 496 1294
rect 446 1277 462 1286
rect 55 1266 106 1274
rect 153 1266 417 1274
rect 443 1274 462 1277
rect 469 1274 496 1286
rect 443 1266 496 1274
rect 71 1258 72 1266
rect 87 1258 100 1266
rect 71 1250 87 1258
rect 68 1243 87 1246
rect 68 1234 90 1243
rect 41 1224 90 1234
rect 41 1218 71 1224
rect 90 1219 95 1224
rect 13 1202 87 1218
rect 105 1210 135 1266
rect 170 1256 378 1266
rect 413 1262 458 1266
rect 461 1265 462 1266
rect 477 1265 490 1266
rect 196 1226 385 1256
rect 211 1223 385 1226
rect 204 1220 385 1223
rect 13 1200 26 1202
rect 41 1200 75 1202
rect 13 1184 87 1200
rect 114 1196 127 1210
rect 142 1196 158 1212
rect 204 1207 215 1220
rect -3 1162 -2 1178
rect 13 1162 26 1184
rect 41 1162 71 1184
rect 114 1180 176 1196
rect 204 1189 215 1205
rect 220 1200 230 1220
rect 240 1200 254 1220
rect 257 1207 266 1220
rect 282 1207 291 1220
rect 220 1189 254 1200
rect 257 1189 266 1205
rect 282 1189 291 1205
rect 298 1200 308 1220
rect 318 1200 332 1220
rect 333 1207 344 1220
rect 298 1189 332 1200
rect 333 1189 344 1205
rect 390 1196 406 1212
rect 413 1210 443 1262
rect 477 1258 478 1265
rect 462 1250 478 1258
rect 449 1218 462 1237
rect 477 1218 507 1234
rect 449 1202 523 1218
rect 449 1200 462 1202
rect 477 1200 511 1202
rect 114 1178 127 1180
rect 142 1178 176 1180
rect 114 1162 176 1178
rect 220 1173 236 1176
rect 298 1173 328 1184
rect 376 1180 422 1196
rect 449 1184 523 1200
rect 376 1178 410 1180
rect 375 1162 422 1178
rect 449 1162 462 1184
rect 477 1162 507 1184
rect 534 1162 535 1178
rect 550 1162 563 1322
rect 593 1218 606 1322
rect 651 1300 652 1310
rect 667 1300 680 1310
rect 651 1296 680 1300
rect 685 1296 715 1322
rect 733 1308 749 1310
rect 821 1308 874 1322
rect 822 1306 886 1308
rect 929 1306 944 1322
rect 993 1319 1023 1322
rect 993 1316 1029 1319
rect 959 1308 975 1310
rect 733 1296 748 1300
rect 651 1294 748 1296
rect 776 1294 944 1306
rect 960 1296 975 1300
rect 993 1297 1032 1316
rect 1051 1310 1058 1311
rect 1057 1303 1058 1310
rect 1041 1300 1042 1303
rect 1057 1300 1070 1303
rect 993 1296 1023 1297
rect 1032 1296 1038 1297
rect 1041 1296 1070 1300
rect 960 1295 1070 1296
rect 960 1294 1076 1295
rect 635 1286 686 1294
rect 635 1274 660 1286
rect 667 1274 686 1286
rect 717 1286 767 1294
rect 717 1278 733 1286
rect 740 1284 767 1286
rect 776 1284 997 1294
rect 740 1274 997 1284
rect 1026 1286 1076 1294
rect 1026 1277 1042 1286
rect 635 1266 686 1274
rect 733 1266 997 1274
rect 1023 1274 1042 1277
rect 1049 1274 1076 1286
rect 1023 1266 1076 1274
rect 651 1258 652 1266
rect 667 1258 680 1266
rect 651 1250 667 1258
rect 648 1243 667 1246
rect 648 1234 670 1243
rect 621 1224 670 1234
rect 621 1218 651 1224
rect 670 1219 675 1224
rect 593 1202 667 1218
rect 685 1210 715 1266
rect 750 1256 958 1266
rect 993 1262 1038 1266
rect 1041 1265 1042 1266
rect 1057 1265 1070 1266
rect 776 1226 965 1256
rect 791 1223 965 1226
rect 784 1220 965 1223
rect 593 1200 606 1202
rect 621 1200 655 1202
rect 593 1184 667 1200
rect 694 1196 707 1210
rect 722 1196 738 1212
rect 784 1207 795 1220
rect 577 1162 578 1178
rect 593 1162 606 1184
rect 621 1162 651 1184
rect 694 1180 756 1196
rect 784 1189 795 1205
rect 800 1200 810 1220
rect 820 1200 834 1220
rect 837 1207 846 1220
rect 862 1207 871 1220
rect 800 1189 834 1200
rect 837 1189 846 1205
rect 862 1189 871 1205
rect 878 1200 888 1220
rect 898 1200 912 1220
rect 913 1207 924 1220
rect 878 1189 912 1200
rect 913 1189 924 1205
rect 970 1196 986 1212
rect 993 1210 1023 1262
rect 1057 1258 1058 1265
rect 1042 1250 1058 1258
rect 1029 1218 1042 1237
rect 1057 1218 1087 1234
rect 1029 1202 1103 1218
rect 1029 1200 1042 1202
rect 1057 1200 1091 1202
rect 694 1178 707 1180
rect 722 1178 756 1180
rect 694 1162 756 1178
rect 800 1173 816 1176
rect 878 1173 908 1184
rect 956 1180 1002 1196
rect 1029 1184 1103 1200
rect 956 1178 990 1180
rect 955 1162 1002 1178
rect 1029 1162 1042 1184
rect 1057 1162 1087 1184
rect 1114 1162 1115 1178
rect 1130 1162 1143 1322
rect 1173 1218 1186 1322
rect 1231 1300 1232 1310
rect 1247 1300 1260 1310
rect 1231 1296 1260 1300
rect 1265 1296 1295 1322
rect 1313 1308 1329 1310
rect 1401 1308 1454 1322
rect 1402 1306 1466 1308
rect 1509 1306 1524 1322
rect 1573 1319 1603 1322
rect 1573 1316 1609 1319
rect 1539 1308 1555 1310
rect 1313 1296 1328 1300
rect 1231 1294 1328 1296
rect 1356 1294 1524 1306
rect 1540 1296 1555 1300
rect 1573 1297 1612 1316
rect 1631 1310 1638 1311
rect 1637 1303 1638 1310
rect 1621 1300 1622 1303
rect 1637 1300 1650 1303
rect 1573 1296 1603 1297
rect 1612 1296 1618 1297
rect 1621 1296 1650 1300
rect 1540 1295 1650 1296
rect 1540 1294 1656 1295
rect 1215 1286 1266 1294
rect 1215 1274 1240 1286
rect 1247 1274 1266 1286
rect 1297 1286 1347 1294
rect 1297 1278 1313 1286
rect 1320 1284 1347 1286
rect 1356 1284 1577 1294
rect 1320 1274 1577 1284
rect 1606 1286 1656 1294
rect 1606 1277 1622 1286
rect 1215 1266 1266 1274
rect 1313 1266 1577 1274
rect 1603 1274 1622 1277
rect 1629 1274 1656 1286
rect 1603 1266 1656 1274
rect 1231 1258 1232 1266
rect 1247 1258 1260 1266
rect 1231 1250 1247 1258
rect 1228 1243 1247 1246
rect 1228 1234 1250 1243
rect 1201 1224 1250 1234
rect 1201 1218 1231 1224
rect 1250 1219 1255 1224
rect 1173 1202 1247 1218
rect 1265 1210 1295 1266
rect 1330 1256 1538 1266
rect 1573 1262 1618 1266
rect 1621 1265 1622 1266
rect 1637 1265 1650 1266
rect 1356 1226 1545 1256
rect 1371 1223 1545 1226
rect 1364 1220 1545 1223
rect 1173 1200 1186 1202
rect 1201 1200 1235 1202
rect 1173 1184 1247 1200
rect 1274 1196 1287 1210
rect 1302 1196 1318 1212
rect 1364 1207 1375 1220
rect 1157 1162 1158 1178
rect 1173 1162 1186 1184
rect 1201 1162 1231 1184
rect 1274 1180 1336 1196
rect 1364 1189 1375 1205
rect 1380 1200 1390 1220
rect 1400 1200 1414 1220
rect 1417 1207 1426 1220
rect 1442 1207 1451 1220
rect 1380 1189 1414 1200
rect 1417 1189 1426 1205
rect 1442 1189 1451 1205
rect 1458 1200 1468 1220
rect 1478 1200 1492 1220
rect 1493 1207 1504 1220
rect 1458 1189 1492 1200
rect 1493 1189 1504 1205
rect 1550 1196 1566 1212
rect 1573 1210 1603 1262
rect 1637 1258 1638 1265
rect 1622 1250 1638 1258
rect 1609 1218 1622 1237
rect 1637 1218 1667 1234
rect 1609 1202 1683 1218
rect 1609 1200 1622 1202
rect 1637 1200 1671 1202
rect 1274 1178 1287 1180
rect 1302 1178 1336 1180
rect 1274 1162 1336 1178
rect 1380 1173 1396 1176
rect 1458 1173 1488 1184
rect 1536 1180 1582 1196
rect 1609 1184 1683 1200
rect 1536 1178 1570 1180
rect 1535 1162 1582 1178
rect 1609 1162 1622 1184
rect 1637 1162 1667 1184
rect 1694 1162 1695 1178
rect 1710 1162 1723 1322
rect 1753 1218 1766 1322
rect 1811 1300 1812 1310
rect 1827 1300 1840 1310
rect 1811 1296 1840 1300
rect 1845 1296 1875 1322
rect 1893 1308 1909 1310
rect 1981 1308 2034 1322
rect 1982 1306 2046 1308
rect 2089 1306 2104 1322
rect 2153 1319 2183 1322
rect 2153 1316 2189 1319
rect 2119 1308 2135 1310
rect 1893 1296 1908 1300
rect 1811 1294 1908 1296
rect 1936 1294 2104 1306
rect 2120 1296 2135 1300
rect 2153 1297 2192 1316
rect 2211 1310 2218 1311
rect 2217 1303 2218 1310
rect 2201 1300 2202 1303
rect 2217 1300 2230 1303
rect 2153 1296 2183 1297
rect 2192 1296 2198 1297
rect 2201 1296 2230 1300
rect 2120 1295 2230 1296
rect 2120 1294 2236 1295
rect 1795 1286 1846 1294
rect 1795 1274 1820 1286
rect 1827 1274 1846 1286
rect 1877 1286 1927 1294
rect 1877 1278 1893 1286
rect 1900 1284 1927 1286
rect 1936 1284 2157 1294
rect 1900 1274 2157 1284
rect 2186 1286 2236 1294
rect 2186 1277 2202 1286
rect 1795 1266 1846 1274
rect 1893 1266 2157 1274
rect 2183 1274 2202 1277
rect 2209 1274 2236 1286
rect 2183 1266 2236 1274
rect 1811 1258 1812 1266
rect 1827 1258 1840 1266
rect 1811 1250 1827 1258
rect 1808 1243 1827 1246
rect 1808 1234 1830 1243
rect 1781 1224 1830 1234
rect 1781 1218 1811 1224
rect 1830 1219 1835 1224
rect 1753 1202 1827 1218
rect 1845 1210 1875 1266
rect 1910 1256 2118 1266
rect 2153 1262 2198 1266
rect 2201 1265 2202 1266
rect 2217 1265 2230 1266
rect 1936 1226 2125 1256
rect 1951 1223 2125 1226
rect 1944 1220 2125 1223
rect 1753 1200 1766 1202
rect 1781 1200 1815 1202
rect 1753 1184 1827 1200
rect 1854 1196 1867 1210
rect 1882 1196 1898 1212
rect 1944 1207 1955 1220
rect 1737 1162 1738 1178
rect 1753 1162 1766 1184
rect 1781 1162 1811 1184
rect 1854 1180 1916 1196
rect 1944 1189 1955 1205
rect 1960 1200 1970 1220
rect 1980 1200 1994 1220
rect 1997 1207 2006 1220
rect 2022 1207 2031 1220
rect 1960 1189 1994 1200
rect 1997 1189 2006 1205
rect 2022 1189 2031 1205
rect 2038 1200 2048 1220
rect 2058 1200 2072 1220
rect 2073 1207 2084 1220
rect 2038 1189 2072 1200
rect 2073 1189 2084 1205
rect 2130 1196 2146 1212
rect 2153 1210 2183 1262
rect 2217 1258 2218 1265
rect 2202 1250 2218 1258
rect 2189 1218 2202 1237
rect 2217 1218 2247 1234
rect 2189 1202 2263 1218
rect 2189 1200 2202 1202
rect 2217 1200 2251 1202
rect 1854 1178 1867 1180
rect 1882 1178 1916 1180
rect 1854 1162 1916 1178
rect 1960 1173 1976 1176
rect 2038 1173 2068 1184
rect 2116 1180 2162 1196
rect 2189 1184 2263 1200
rect 2116 1178 2150 1180
rect 2115 1162 2162 1178
rect 2189 1162 2202 1184
rect 2217 1162 2247 1184
rect 2274 1162 2275 1178
rect 2290 1162 2303 1322
rect 2333 1218 2346 1322
rect 2391 1300 2392 1310
rect 2407 1300 2420 1310
rect 2391 1296 2420 1300
rect 2425 1296 2455 1322
rect 2473 1308 2489 1310
rect 2561 1308 2614 1322
rect 2562 1306 2626 1308
rect 2669 1306 2684 1322
rect 2733 1319 2763 1322
rect 2733 1316 2769 1319
rect 2699 1308 2715 1310
rect 2473 1296 2488 1300
rect 2391 1294 2488 1296
rect 2516 1294 2684 1306
rect 2700 1296 2715 1300
rect 2733 1297 2772 1316
rect 2791 1310 2798 1311
rect 2797 1303 2798 1310
rect 2781 1300 2782 1303
rect 2797 1300 2810 1303
rect 2733 1296 2763 1297
rect 2772 1296 2778 1297
rect 2781 1296 2810 1300
rect 2700 1295 2810 1296
rect 2700 1294 2816 1295
rect 2375 1286 2426 1294
rect 2375 1274 2400 1286
rect 2407 1274 2426 1286
rect 2457 1286 2507 1294
rect 2457 1278 2473 1286
rect 2480 1284 2507 1286
rect 2516 1284 2737 1294
rect 2480 1274 2737 1284
rect 2766 1286 2816 1294
rect 2766 1277 2782 1286
rect 2375 1266 2426 1274
rect 2473 1266 2737 1274
rect 2763 1274 2782 1277
rect 2789 1274 2816 1286
rect 2763 1266 2816 1274
rect 2391 1258 2392 1266
rect 2407 1258 2420 1266
rect 2391 1250 2407 1258
rect 2388 1243 2407 1246
rect 2388 1234 2410 1243
rect 2361 1224 2410 1234
rect 2361 1218 2391 1224
rect 2410 1219 2415 1224
rect 2333 1202 2407 1218
rect 2425 1210 2455 1266
rect 2490 1256 2698 1266
rect 2733 1262 2778 1266
rect 2781 1265 2782 1266
rect 2797 1265 2810 1266
rect 2516 1226 2705 1256
rect 2531 1223 2705 1226
rect 2524 1220 2705 1223
rect 2333 1200 2346 1202
rect 2361 1200 2395 1202
rect 2333 1184 2407 1200
rect 2434 1196 2447 1210
rect 2462 1196 2478 1212
rect 2524 1207 2535 1220
rect 2317 1162 2318 1178
rect 2333 1162 2346 1184
rect 2361 1162 2391 1184
rect 2434 1180 2496 1196
rect 2524 1189 2535 1205
rect 2540 1200 2550 1220
rect 2560 1200 2574 1220
rect 2577 1207 2586 1220
rect 2602 1207 2611 1220
rect 2540 1189 2574 1200
rect 2577 1189 2586 1205
rect 2602 1189 2611 1205
rect 2618 1200 2628 1220
rect 2638 1200 2652 1220
rect 2653 1207 2664 1220
rect 2618 1189 2652 1200
rect 2653 1189 2664 1205
rect 2710 1196 2726 1212
rect 2733 1210 2763 1262
rect 2797 1258 2798 1265
rect 2782 1250 2798 1258
rect 2769 1218 2782 1237
rect 2797 1218 2827 1234
rect 2769 1202 2843 1218
rect 2769 1200 2782 1202
rect 2797 1200 2831 1202
rect 2434 1178 2447 1180
rect 2462 1178 2496 1180
rect 2434 1162 2496 1178
rect 2540 1173 2556 1176
rect 2618 1173 2648 1184
rect 2696 1180 2742 1196
rect 2769 1184 2843 1200
rect 2696 1178 2730 1180
rect 2695 1162 2742 1178
rect 2769 1162 2782 1184
rect 2797 1162 2827 1184
rect 2854 1162 2855 1178
rect 2870 1162 2883 1322
rect 2913 1218 2926 1322
rect 2971 1300 2972 1310
rect 2987 1300 3000 1310
rect 2971 1296 3000 1300
rect 3005 1296 3035 1322
rect 3053 1308 3069 1310
rect 3141 1308 3194 1322
rect 3142 1306 3206 1308
rect 3249 1306 3264 1322
rect 3313 1319 3343 1322
rect 3313 1316 3349 1319
rect 3279 1308 3295 1310
rect 3053 1296 3068 1300
rect 2971 1294 3068 1296
rect 3096 1294 3264 1306
rect 3280 1296 3295 1300
rect 3313 1297 3352 1316
rect 3371 1310 3378 1311
rect 3377 1303 3378 1310
rect 3361 1300 3362 1303
rect 3377 1300 3390 1303
rect 3313 1296 3343 1297
rect 3352 1296 3358 1297
rect 3361 1296 3390 1300
rect 3280 1295 3390 1296
rect 3280 1294 3396 1295
rect 2955 1286 3006 1294
rect 2955 1274 2980 1286
rect 2987 1274 3006 1286
rect 3037 1286 3087 1294
rect 3037 1278 3053 1286
rect 3060 1284 3087 1286
rect 3096 1284 3317 1294
rect 3060 1274 3317 1284
rect 3346 1286 3396 1294
rect 3346 1277 3362 1286
rect 2955 1266 3006 1274
rect 3053 1266 3317 1274
rect 3343 1274 3362 1277
rect 3369 1274 3396 1286
rect 3343 1266 3396 1274
rect 2971 1258 2972 1266
rect 2987 1258 3000 1266
rect 2971 1250 2987 1258
rect 2968 1243 2987 1246
rect 2968 1234 2990 1243
rect 2941 1224 2990 1234
rect 2941 1218 2971 1224
rect 2990 1219 2995 1224
rect 2913 1202 2987 1218
rect 3005 1210 3035 1266
rect 3070 1256 3278 1266
rect 3313 1262 3358 1266
rect 3361 1265 3362 1266
rect 3377 1265 3390 1266
rect 3096 1226 3285 1256
rect 3111 1223 3285 1226
rect 3104 1220 3285 1223
rect 2913 1200 2926 1202
rect 2941 1200 2975 1202
rect 2913 1184 2987 1200
rect 3014 1196 3027 1210
rect 3042 1196 3058 1212
rect 3104 1207 3115 1220
rect 2897 1162 2898 1178
rect 2913 1162 2926 1184
rect 2941 1162 2971 1184
rect 3014 1180 3076 1196
rect 3104 1189 3115 1205
rect 3120 1200 3130 1220
rect 3140 1200 3154 1220
rect 3157 1207 3166 1220
rect 3182 1207 3191 1220
rect 3120 1189 3154 1200
rect 3157 1189 3166 1205
rect 3182 1189 3191 1205
rect 3198 1200 3208 1220
rect 3218 1200 3232 1220
rect 3233 1207 3244 1220
rect 3198 1189 3232 1200
rect 3233 1189 3244 1205
rect 3290 1196 3306 1212
rect 3313 1210 3343 1262
rect 3377 1258 3378 1265
rect 3362 1250 3378 1258
rect 3349 1218 3362 1237
rect 3377 1218 3407 1234
rect 3349 1202 3423 1218
rect 3349 1200 3362 1202
rect 3377 1200 3411 1202
rect 3014 1178 3027 1180
rect 3042 1178 3076 1180
rect 3014 1162 3076 1178
rect 3120 1173 3136 1176
rect 3198 1173 3228 1184
rect 3276 1180 3322 1196
rect 3349 1184 3423 1200
rect 3276 1178 3310 1180
rect 3275 1162 3322 1178
rect 3349 1162 3362 1184
rect 3377 1162 3407 1184
rect 3434 1162 3435 1178
rect 3450 1162 3463 1322
rect 5911 1218 5924 1322
rect 5969 1300 5970 1310
rect 5985 1300 5998 1310
rect 5969 1296 5998 1300
rect 6003 1296 6033 1322
rect 6051 1308 6067 1310
rect 6139 1308 6192 1322
rect 6140 1306 6204 1308
rect 6247 1306 6262 1322
rect 6311 1319 6341 1322
rect 6311 1316 6347 1319
rect 6277 1308 6293 1310
rect 6051 1296 6066 1300
rect 5969 1294 6066 1296
rect 6094 1294 6262 1306
rect 6278 1296 6293 1300
rect 6311 1297 6350 1316
rect 6369 1310 6376 1311
rect 6375 1303 6376 1310
rect 6359 1300 6360 1303
rect 6375 1300 6388 1303
rect 6311 1296 6341 1297
rect 6350 1296 6356 1297
rect 6359 1296 6388 1300
rect 6278 1295 6388 1296
rect 6278 1294 6394 1295
rect 5953 1286 6004 1294
rect 5953 1274 5978 1286
rect 5985 1274 6004 1286
rect 6035 1286 6085 1294
rect 6035 1278 6051 1286
rect 6058 1284 6085 1286
rect 6094 1284 6315 1294
rect 6058 1274 6315 1284
rect 6344 1286 6394 1294
rect 6344 1277 6360 1286
rect 5953 1266 6004 1274
rect 6051 1266 6315 1274
rect 6341 1274 6360 1277
rect 6367 1274 6394 1286
rect 6341 1266 6394 1274
rect 5969 1258 5970 1266
rect 5985 1258 5998 1266
rect 5969 1250 5985 1258
rect 5966 1243 5985 1246
rect 5966 1234 5988 1243
rect 5939 1224 5988 1234
rect 5939 1218 5969 1224
rect 5988 1219 5993 1224
rect 5911 1202 5985 1218
rect 6003 1210 6033 1266
rect 6068 1256 6276 1266
rect 6311 1262 6356 1266
rect 6359 1265 6360 1266
rect 6375 1265 6388 1266
rect 6094 1226 6283 1256
rect 6109 1223 6283 1226
rect 6102 1220 6283 1223
rect 5911 1200 5924 1202
rect 5939 1200 5973 1202
rect 5911 1184 5985 1200
rect 6012 1196 6025 1210
rect 6040 1196 6056 1212
rect 6102 1207 6113 1220
rect 5895 1162 5896 1178
rect 5911 1162 5924 1184
rect 5939 1162 5969 1184
rect 6012 1180 6074 1196
rect 6102 1189 6113 1205
rect 6118 1200 6128 1220
rect 6138 1200 6152 1220
rect 6155 1207 6164 1220
rect 6180 1207 6189 1220
rect 6118 1189 6152 1200
rect 6155 1189 6164 1205
rect 6180 1189 6189 1205
rect 6196 1200 6206 1220
rect 6216 1200 6230 1220
rect 6231 1207 6242 1220
rect 6196 1189 6230 1200
rect 6231 1189 6242 1205
rect 6288 1196 6304 1212
rect 6311 1210 6341 1262
rect 6375 1258 6376 1265
rect 6360 1250 6376 1258
rect 6347 1218 6360 1237
rect 6375 1218 6405 1234
rect 6347 1202 6421 1218
rect 6347 1200 6360 1202
rect 6375 1200 6409 1202
rect 6012 1178 6025 1180
rect 6040 1178 6074 1180
rect 6012 1162 6074 1178
rect 6118 1173 6134 1176
rect 6196 1173 6226 1184
rect 6274 1180 6320 1196
rect 6347 1184 6421 1200
rect 6274 1178 6308 1180
rect 6273 1162 6320 1178
rect 6347 1162 6360 1184
rect 6375 1162 6405 1184
rect 6432 1162 6433 1178
rect 6448 1162 6461 1322
rect 6491 1218 6504 1322
rect 6549 1300 6550 1310
rect 6565 1300 6578 1310
rect 6549 1296 6578 1300
rect 6583 1296 6613 1322
rect 6631 1308 6647 1310
rect 6719 1308 6772 1322
rect 6720 1306 6784 1308
rect 6827 1306 6842 1322
rect 6891 1319 6921 1322
rect 6891 1316 6927 1319
rect 6857 1308 6873 1310
rect 6631 1296 6646 1300
rect 6549 1294 6646 1296
rect 6674 1294 6842 1306
rect 6858 1296 6873 1300
rect 6891 1297 6930 1316
rect 6949 1310 6956 1311
rect 6955 1303 6956 1310
rect 6939 1300 6940 1303
rect 6955 1300 6968 1303
rect 6891 1296 6921 1297
rect 6930 1296 6936 1297
rect 6939 1296 6968 1300
rect 6858 1295 6968 1296
rect 6858 1294 6974 1295
rect 6533 1286 6584 1294
rect 6533 1274 6558 1286
rect 6565 1274 6584 1286
rect 6615 1286 6665 1294
rect 6615 1278 6631 1286
rect 6638 1284 6665 1286
rect 6674 1284 6895 1294
rect 6638 1274 6895 1284
rect 6924 1286 6974 1294
rect 6924 1277 6940 1286
rect 6533 1266 6584 1274
rect 6631 1266 6895 1274
rect 6921 1274 6940 1277
rect 6947 1274 6974 1286
rect 6921 1266 6974 1274
rect 6549 1258 6550 1266
rect 6565 1258 6578 1266
rect 6549 1250 6565 1258
rect 6546 1243 6565 1246
rect 6546 1234 6568 1243
rect 6519 1224 6568 1234
rect 6519 1218 6549 1224
rect 6568 1219 6573 1224
rect 6491 1202 6565 1218
rect 6583 1210 6613 1266
rect 6648 1256 6856 1266
rect 6891 1262 6936 1266
rect 6939 1265 6940 1266
rect 6955 1265 6968 1266
rect 6674 1226 6863 1256
rect 6689 1223 6863 1226
rect 6682 1220 6863 1223
rect 6491 1200 6504 1202
rect 6519 1200 6553 1202
rect 6491 1184 6565 1200
rect 6592 1196 6605 1210
rect 6620 1196 6636 1212
rect 6682 1207 6693 1220
rect 6475 1162 6476 1178
rect 6491 1162 6504 1184
rect 6519 1162 6549 1184
rect 6592 1180 6654 1196
rect 6682 1189 6693 1205
rect 6698 1200 6708 1220
rect 6718 1200 6732 1220
rect 6735 1207 6744 1220
rect 6760 1207 6769 1220
rect 6698 1189 6732 1200
rect 6735 1189 6744 1205
rect 6760 1189 6769 1205
rect 6776 1200 6786 1220
rect 6796 1200 6810 1220
rect 6811 1207 6822 1220
rect 6776 1189 6810 1200
rect 6811 1189 6822 1205
rect 6868 1196 6884 1212
rect 6891 1210 6921 1262
rect 6955 1258 6956 1265
rect 6940 1250 6956 1258
rect 6927 1218 6940 1237
rect 6955 1218 6985 1234
rect 6927 1202 7001 1218
rect 6927 1200 6940 1202
rect 6955 1200 6989 1202
rect 6592 1178 6605 1180
rect 6620 1178 6654 1180
rect 6592 1162 6654 1178
rect 6698 1173 6714 1176
rect 6776 1173 6806 1184
rect 6854 1180 6900 1196
rect 6927 1184 7001 1200
rect 6854 1178 6888 1180
rect 6853 1162 6900 1178
rect 6927 1162 6940 1184
rect 6955 1162 6985 1184
rect 7012 1162 7013 1178
rect 7028 1162 7041 1322
rect 7071 1218 7084 1322
rect 7129 1300 7130 1310
rect 7145 1300 7158 1310
rect 7129 1296 7158 1300
rect 7163 1296 7193 1322
rect 7211 1308 7227 1310
rect 7299 1308 7352 1322
rect 7300 1306 7364 1308
rect 7407 1306 7422 1322
rect 7471 1319 7501 1322
rect 7471 1316 7507 1319
rect 7437 1308 7453 1310
rect 7211 1296 7226 1300
rect 7129 1294 7226 1296
rect 7254 1294 7422 1306
rect 7438 1296 7453 1300
rect 7471 1297 7510 1316
rect 7529 1310 7536 1311
rect 7535 1303 7536 1310
rect 7519 1300 7520 1303
rect 7535 1300 7548 1303
rect 7471 1296 7501 1297
rect 7510 1296 7516 1297
rect 7519 1296 7548 1300
rect 7438 1295 7548 1296
rect 7438 1294 7554 1295
rect 7113 1286 7164 1294
rect 7113 1274 7138 1286
rect 7145 1274 7164 1286
rect 7195 1286 7245 1294
rect 7195 1278 7211 1286
rect 7218 1284 7245 1286
rect 7254 1284 7475 1294
rect 7218 1274 7475 1284
rect 7504 1286 7554 1294
rect 7504 1277 7520 1286
rect 7113 1266 7164 1274
rect 7211 1266 7475 1274
rect 7501 1274 7520 1277
rect 7527 1274 7554 1286
rect 7501 1266 7554 1274
rect 7129 1258 7130 1266
rect 7145 1258 7158 1266
rect 7129 1250 7145 1258
rect 7126 1243 7145 1246
rect 7126 1234 7148 1243
rect 7099 1224 7148 1234
rect 7099 1218 7129 1224
rect 7148 1219 7153 1224
rect 7071 1202 7145 1218
rect 7163 1210 7193 1266
rect 7228 1256 7436 1266
rect 7471 1262 7516 1266
rect 7519 1265 7520 1266
rect 7535 1265 7548 1266
rect 7254 1226 7443 1256
rect 7269 1223 7443 1226
rect 7262 1220 7443 1223
rect 7071 1200 7084 1202
rect 7099 1200 7133 1202
rect 7071 1184 7145 1200
rect 7172 1196 7185 1210
rect 7200 1196 7216 1212
rect 7262 1207 7273 1220
rect 7055 1162 7056 1178
rect 7071 1162 7084 1184
rect 7099 1162 7129 1184
rect 7172 1180 7234 1196
rect 7262 1189 7273 1205
rect 7278 1200 7288 1220
rect 7298 1200 7312 1220
rect 7315 1207 7324 1220
rect 7340 1207 7349 1220
rect 7278 1189 7312 1200
rect 7315 1189 7324 1205
rect 7340 1189 7349 1205
rect 7356 1200 7366 1220
rect 7376 1200 7390 1220
rect 7391 1207 7402 1220
rect 7356 1189 7390 1200
rect 7391 1189 7402 1205
rect 7448 1196 7464 1212
rect 7471 1210 7501 1262
rect 7535 1258 7536 1265
rect 7520 1250 7536 1258
rect 7507 1218 7520 1237
rect 7535 1218 7565 1234
rect 7507 1202 7581 1218
rect 7507 1200 7520 1202
rect 7535 1200 7569 1202
rect 7172 1178 7185 1180
rect 7200 1178 7234 1180
rect 7172 1162 7234 1178
rect 7278 1173 7294 1176
rect 7356 1173 7386 1184
rect 7434 1180 7480 1196
rect 7507 1184 7581 1200
rect 7434 1178 7468 1180
rect 7433 1162 7480 1178
rect 7507 1162 7520 1184
rect 7535 1162 7565 1184
rect 7592 1162 7593 1178
rect 7608 1162 7621 1322
rect 7651 1218 7664 1322
rect 7709 1300 7710 1310
rect 7725 1300 7738 1310
rect 7709 1296 7738 1300
rect 7743 1296 7773 1322
rect 7791 1308 7807 1310
rect 7879 1308 7932 1322
rect 7880 1306 7944 1308
rect 7987 1306 8002 1322
rect 8051 1319 8081 1322
rect 8051 1316 8087 1319
rect 8017 1308 8033 1310
rect 7791 1296 7806 1300
rect 7709 1294 7806 1296
rect 7834 1294 8002 1306
rect 8018 1296 8033 1300
rect 8051 1297 8090 1316
rect 8109 1310 8116 1311
rect 8115 1303 8116 1310
rect 8099 1300 8100 1303
rect 8115 1300 8128 1303
rect 8051 1296 8081 1297
rect 8090 1296 8096 1297
rect 8099 1296 8128 1300
rect 8018 1295 8128 1296
rect 8018 1294 8134 1295
rect 7693 1286 7744 1294
rect 7693 1274 7718 1286
rect 7725 1274 7744 1286
rect 7775 1286 7825 1294
rect 7775 1278 7791 1286
rect 7798 1284 7825 1286
rect 7834 1284 8055 1294
rect 7798 1274 8055 1284
rect 8084 1286 8134 1294
rect 8084 1277 8100 1286
rect 7693 1266 7744 1274
rect 7791 1266 8055 1274
rect 8081 1274 8100 1277
rect 8107 1274 8134 1286
rect 8081 1266 8134 1274
rect 7709 1258 7710 1266
rect 7725 1258 7738 1266
rect 7709 1250 7725 1258
rect 7706 1243 7725 1246
rect 7706 1234 7728 1243
rect 7679 1224 7728 1234
rect 7679 1218 7709 1224
rect 7728 1219 7733 1224
rect 7651 1202 7725 1218
rect 7743 1210 7773 1266
rect 7808 1256 8016 1266
rect 8051 1262 8096 1266
rect 8099 1265 8100 1266
rect 8115 1265 8128 1266
rect 7834 1226 8023 1256
rect 7849 1223 8023 1226
rect 7842 1220 8023 1223
rect 7651 1200 7664 1202
rect 7679 1200 7713 1202
rect 7651 1184 7725 1200
rect 7752 1196 7765 1210
rect 7780 1196 7796 1212
rect 7842 1207 7853 1220
rect 7635 1162 7636 1178
rect 7651 1162 7664 1184
rect 7679 1162 7709 1184
rect 7752 1180 7814 1196
rect 7842 1189 7853 1205
rect 7858 1200 7868 1220
rect 7878 1200 7892 1220
rect 7895 1207 7904 1220
rect 7920 1207 7929 1220
rect 7858 1189 7892 1200
rect 7895 1189 7904 1205
rect 7920 1189 7929 1205
rect 7936 1200 7946 1220
rect 7956 1200 7970 1220
rect 7971 1207 7982 1220
rect 7936 1189 7970 1200
rect 7971 1189 7982 1205
rect 8028 1196 8044 1212
rect 8051 1210 8081 1262
rect 8115 1258 8116 1265
rect 8100 1250 8116 1258
rect 8087 1218 8100 1237
rect 8115 1218 8145 1234
rect 8087 1202 8161 1218
rect 8087 1200 8100 1202
rect 8115 1200 8149 1202
rect 7752 1178 7765 1180
rect 7780 1178 7814 1180
rect 7752 1162 7814 1178
rect 7858 1173 7874 1176
rect 7936 1173 7966 1184
rect 8014 1180 8060 1196
rect 8087 1184 8161 1200
rect 8014 1178 8048 1180
rect 8013 1162 8060 1178
rect 8087 1162 8100 1184
rect 8115 1162 8145 1184
rect 8172 1162 8173 1178
rect 8188 1162 8201 1322
rect 8231 1218 8244 1322
rect 8289 1300 8290 1310
rect 8305 1300 8318 1310
rect 8289 1296 8318 1300
rect 8323 1296 8353 1322
rect 8371 1308 8387 1310
rect 8459 1308 8512 1322
rect 8460 1306 8524 1308
rect 8567 1306 8582 1322
rect 8631 1319 8661 1322
rect 8631 1316 8667 1319
rect 8597 1308 8613 1310
rect 8371 1296 8386 1300
rect 8289 1294 8386 1296
rect 8414 1294 8582 1306
rect 8598 1296 8613 1300
rect 8631 1297 8670 1316
rect 8689 1310 8696 1311
rect 8695 1303 8696 1310
rect 8679 1300 8680 1303
rect 8695 1300 8708 1303
rect 8631 1296 8661 1297
rect 8670 1296 8676 1297
rect 8679 1296 8708 1300
rect 8598 1295 8708 1296
rect 8598 1294 8714 1295
rect 8273 1286 8324 1294
rect 8273 1274 8298 1286
rect 8305 1274 8324 1286
rect 8355 1286 8405 1294
rect 8355 1278 8371 1286
rect 8378 1284 8405 1286
rect 8414 1284 8635 1294
rect 8378 1274 8635 1284
rect 8664 1286 8714 1294
rect 8664 1277 8680 1286
rect 8273 1266 8324 1274
rect 8371 1266 8635 1274
rect 8661 1274 8680 1277
rect 8687 1274 8714 1286
rect 8661 1266 8714 1274
rect 8289 1258 8290 1266
rect 8305 1258 8318 1266
rect 8289 1250 8305 1258
rect 8286 1243 8305 1246
rect 8286 1234 8308 1243
rect 8259 1224 8308 1234
rect 8259 1218 8289 1224
rect 8308 1219 8313 1224
rect 8231 1202 8305 1218
rect 8323 1210 8353 1266
rect 8388 1256 8596 1266
rect 8631 1262 8676 1266
rect 8679 1265 8680 1266
rect 8695 1265 8708 1266
rect 8414 1226 8603 1256
rect 8429 1223 8603 1226
rect 8422 1220 8603 1223
rect 8231 1200 8244 1202
rect 8259 1200 8293 1202
rect 8231 1184 8305 1200
rect 8332 1196 8345 1210
rect 8360 1196 8376 1212
rect 8422 1207 8433 1220
rect 8215 1162 8216 1178
rect 8231 1162 8244 1184
rect 8259 1162 8289 1184
rect 8332 1180 8394 1196
rect 8422 1189 8433 1205
rect 8438 1200 8448 1220
rect 8458 1200 8472 1220
rect 8475 1207 8484 1220
rect 8500 1207 8509 1220
rect 8438 1189 8472 1200
rect 8475 1189 8484 1205
rect 8500 1189 8509 1205
rect 8516 1200 8526 1220
rect 8536 1200 8550 1220
rect 8551 1207 8562 1220
rect 8516 1189 8550 1200
rect 8551 1189 8562 1205
rect 8608 1196 8624 1212
rect 8631 1210 8661 1262
rect 8695 1258 8696 1265
rect 8680 1250 8696 1258
rect 8667 1218 8680 1237
rect 8695 1218 8725 1234
rect 8667 1202 8741 1218
rect 8667 1200 8680 1202
rect 8695 1200 8729 1202
rect 8332 1178 8345 1180
rect 8360 1178 8394 1180
rect 8332 1162 8394 1178
rect 8438 1173 8454 1176
rect 8516 1173 8546 1184
rect 8594 1180 8640 1196
rect 8667 1184 8741 1200
rect 8594 1178 8628 1180
rect 8593 1162 8640 1178
rect 8667 1162 8680 1184
rect 8695 1162 8725 1184
rect 8752 1162 8753 1178
rect 8768 1162 8781 1322
rect 8811 1218 8824 1322
rect 8869 1300 8870 1310
rect 8885 1300 8898 1310
rect 8869 1296 8898 1300
rect 8903 1296 8933 1322
rect 8951 1308 8967 1310
rect 9039 1308 9092 1322
rect 9040 1306 9104 1308
rect 9147 1306 9162 1322
rect 9211 1319 9241 1322
rect 9211 1316 9247 1319
rect 9177 1308 9193 1310
rect 8951 1296 8966 1300
rect 8869 1294 8966 1296
rect 8994 1294 9162 1306
rect 9178 1296 9193 1300
rect 9211 1297 9250 1316
rect 9269 1310 9276 1311
rect 9275 1303 9276 1310
rect 9259 1300 9260 1303
rect 9275 1300 9288 1303
rect 9211 1296 9241 1297
rect 9250 1296 9256 1297
rect 9259 1296 9288 1300
rect 9178 1295 9288 1296
rect 9178 1294 9294 1295
rect 8853 1286 8904 1294
rect 8853 1274 8878 1286
rect 8885 1274 8904 1286
rect 8935 1286 8985 1294
rect 8935 1278 8951 1286
rect 8958 1284 8985 1286
rect 8994 1284 9215 1294
rect 8958 1274 9215 1284
rect 9244 1286 9294 1294
rect 9244 1277 9260 1286
rect 8853 1266 8904 1274
rect 8951 1266 9215 1274
rect 9241 1274 9260 1277
rect 9267 1274 9294 1286
rect 9241 1266 9294 1274
rect 8869 1258 8870 1266
rect 8885 1258 8898 1266
rect 8869 1250 8885 1258
rect 8866 1243 8885 1246
rect 8866 1234 8888 1243
rect 8839 1224 8888 1234
rect 8839 1218 8869 1224
rect 8888 1219 8893 1224
rect 8811 1202 8885 1218
rect 8903 1210 8933 1266
rect 8968 1256 9176 1266
rect 9211 1262 9256 1266
rect 9259 1265 9260 1266
rect 9275 1265 9288 1266
rect 8994 1226 9183 1256
rect 9009 1223 9183 1226
rect 9002 1220 9183 1223
rect 8811 1200 8824 1202
rect 8839 1200 8873 1202
rect 8811 1184 8885 1200
rect 8912 1196 8925 1210
rect 8940 1196 8956 1212
rect 9002 1207 9013 1220
rect 8795 1162 8796 1178
rect 8811 1162 8824 1184
rect 8839 1162 8869 1184
rect 8912 1180 8974 1196
rect 9002 1189 9013 1205
rect 9018 1200 9028 1220
rect 9038 1200 9052 1220
rect 9055 1207 9064 1220
rect 9080 1207 9089 1220
rect 9018 1189 9052 1200
rect 9055 1189 9064 1205
rect 9080 1189 9089 1205
rect 9096 1200 9106 1220
rect 9116 1200 9130 1220
rect 9131 1207 9142 1220
rect 9096 1189 9130 1200
rect 9131 1189 9142 1205
rect 9188 1196 9204 1212
rect 9211 1210 9241 1262
rect 9275 1258 9276 1265
rect 9260 1250 9276 1258
rect 9247 1218 9260 1237
rect 9275 1218 9305 1234
rect 9247 1202 9321 1218
rect 9247 1200 9260 1202
rect 9275 1200 9309 1202
rect 8912 1178 8925 1180
rect 8940 1178 8974 1180
rect 8912 1162 8974 1178
rect 9018 1173 9034 1176
rect 9096 1173 9126 1184
rect 9174 1180 9220 1196
rect 9247 1184 9321 1200
rect 9174 1178 9208 1180
rect 9173 1162 9220 1178
rect 9247 1162 9260 1184
rect 9275 1162 9305 1184
rect 9332 1162 9333 1178
rect 9348 1162 9361 1322
rect -9 1154 32 1162
rect -9 1128 6 1154
rect 13 1128 32 1154
rect 96 1150 158 1162
rect 170 1150 245 1162
rect 303 1150 378 1162
rect 390 1150 421 1162
rect 427 1150 462 1162
rect 96 1148 258 1150
rect -9 1120 32 1128
rect 114 1124 127 1148
rect 142 1146 157 1148
rect -3 1110 -2 1120
rect 13 1110 26 1120
rect 41 1110 71 1124
rect 114 1110 157 1124
rect 181 1121 188 1128
rect 191 1124 258 1148
rect 290 1148 462 1150
rect 260 1126 288 1130
rect 290 1126 370 1148
rect 391 1146 406 1148
rect 260 1124 370 1126
rect 191 1120 370 1124
rect 164 1110 194 1120
rect 196 1110 349 1120
rect 357 1110 387 1120
rect 391 1110 421 1124
rect 449 1110 462 1148
rect 534 1154 569 1162
rect 534 1128 535 1154
rect 542 1128 569 1154
rect 477 1110 507 1124
rect 534 1120 569 1128
rect 571 1154 612 1162
rect 571 1128 586 1154
rect 593 1128 612 1154
rect 676 1150 738 1162
rect 750 1150 825 1162
rect 883 1150 958 1162
rect 970 1150 1001 1162
rect 1007 1150 1042 1162
rect 676 1148 838 1150
rect 571 1120 612 1128
rect 694 1124 707 1148
rect 722 1146 737 1148
rect 534 1110 535 1120
rect 550 1110 563 1120
rect 577 1110 578 1120
rect 593 1110 606 1120
rect 621 1110 651 1124
rect 694 1110 737 1124
rect 761 1121 768 1128
rect 771 1124 838 1148
rect 870 1148 1042 1150
rect 840 1126 868 1130
rect 870 1126 950 1148
rect 971 1146 986 1148
rect 840 1124 950 1126
rect 771 1120 950 1124
rect 744 1110 774 1120
rect 776 1110 929 1120
rect 937 1110 967 1120
rect 971 1110 1001 1124
rect 1029 1110 1042 1148
rect 1114 1154 1149 1162
rect 1114 1128 1115 1154
rect 1122 1128 1149 1154
rect 1057 1110 1087 1124
rect 1114 1120 1149 1128
rect 1151 1154 1192 1162
rect 1151 1128 1166 1154
rect 1173 1128 1192 1154
rect 1256 1150 1318 1162
rect 1330 1150 1405 1162
rect 1463 1150 1538 1162
rect 1550 1150 1581 1162
rect 1587 1150 1622 1162
rect 1256 1148 1418 1150
rect 1151 1120 1192 1128
rect 1274 1124 1287 1148
rect 1302 1146 1317 1148
rect 1114 1110 1115 1120
rect 1130 1110 1143 1120
rect 1157 1110 1158 1120
rect 1173 1110 1186 1120
rect 1201 1110 1231 1124
rect 1274 1110 1317 1124
rect 1341 1121 1348 1128
rect 1351 1124 1418 1148
rect 1450 1148 1622 1150
rect 1420 1126 1448 1130
rect 1450 1126 1530 1148
rect 1551 1146 1566 1148
rect 1420 1124 1530 1126
rect 1351 1120 1530 1124
rect 1324 1110 1354 1120
rect 1356 1110 1509 1120
rect 1517 1110 1547 1120
rect 1551 1110 1581 1124
rect 1609 1110 1622 1148
rect 1694 1154 1729 1162
rect 1694 1128 1695 1154
rect 1702 1128 1729 1154
rect 1637 1110 1667 1124
rect 1694 1120 1729 1128
rect 1731 1154 1772 1162
rect 1731 1128 1746 1154
rect 1753 1128 1772 1154
rect 1836 1150 1898 1162
rect 1910 1150 1985 1162
rect 2043 1150 2118 1162
rect 2130 1150 2161 1162
rect 2167 1150 2202 1162
rect 1836 1148 1998 1150
rect 1731 1120 1772 1128
rect 1854 1124 1867 1148
rect 1882 1146 1897 1148
rect 1694 1110 1695 1120
rect 1710 1110 1723 1120
rect 1737 1110 1738 1120
rect 1753 1110 1766 1120
rect 1781 1110 1811 1124
rect 1854 1110 1897 1124
rect 1921 1121 1928 1128
rect 1931 1124 1998 1148
rect 2030 1148 2202 1150
rect 2000 1126 2028 1130
rect 2030 1126 2110 1148
rect 2131 1146 2146 1148
rect 2000 1124 2110 1126
rect 1931 1120 2110 1124
rect 1904 1110 1934 1120
rect 1936 1110 2089 1120
rect 2097 1110 2127 1120
rect 2131 1110 2161 1124
rect 2189 1110 2202 1148
rect 2274 1154 2309 1162
rect 2274 1128 2275 1154
rect 2282 1128 2309 1154
rect 2217 1110 2247 1124
rect 2274 1120 2309 1128
rect 2311 1154 2352 1162
rect 2311 1128 2326 1154
rect 2333 1128 2352 1154
rect 2416 1150 2478 1162
rect 2490 1150 2565 1162
rect 2623 1150 2698 1162
rect 2710 1150 2741 1162
rect 2747 1150 2782 1162
rect 2416 1148 2578 1150
rect 2311 1120 2352 1128
rect 2434 1124 2447 1148
rect 2462 1146 2477 1148
rect 2274 1110 2275 1120
rect 2290 1110 2303 1120
rect 2317 1110 2318 1120
rect 2333 1110 2346 1120
rect 2361 1110 2391 1124
rect 2434 1110 2477 1124
rect 2501 1121 2508 1128
rect 2511 1124 2578 1148
rect 2610 1148 2782 1150
rect 2580 1126 2608 1130
rect 2610 1126 2690 1148
rect 2711 1146 2726 1148
rect 2580 1124 2690 1126
rect 2511 1120 2690 1124
rect 2484 1110 2514 1120
rect 2516 1110 2669 1120
rect 2677 1110 2707 1120
rect 2711 1110 2741 1124
rect 2769 1110 2782 1148
rect 2854 1154 2889 1162
rect 2854 1128 2855 1154
rect 2862 1128 2889 1154
rect 2797 1110 2827 1124
rect 2854 1120 2889 1128
rect 2891 1154 2932 1162
rect 2891 1128 2906 1154
rect 2913 1128 2932 1154
rect 2996 1150 3058 1162
rect 3070 1150 3145 1162
rect 3203 1150 3278 1162
rect 3290 1150 3321 1162
rect 3327 1150 3362 1162
rect 2996 1148 3158 1150
rect 2891 1120 2932 1128
rect 3014 1124 3027 1148
rect 3042 1146 3057 1148
rect 2854 1110 2855 1120
rect 2870 1110 2883 1120
rect 2897 1110 2898 1120
rect 2913 1110 2926 1120
rect 2941 1110 2971 1124
rect 3014 1110 3057 1124
rect 3081 1121 3088 1128
rect 3091 1124 3158 1148
rect 3190 1148 3362 1150
rect 3160 1126 3188 1130
rect 3190 1126 3270 1148
rect 3291 1146 3306 1148
rect 3160 1124 3270 1126
rect 3091 1120 3270 1124
rect 3064 1110 3094 1120
rect 3096 1110 3249 1120
rect 3257 1110 3287 1120
rect 3291 1110 3321 1124
rect 3349 1110 3362 1148
rect 3434 1154 3469 1162
rect 3434 1128 3435 1154
rect 3442 1128 3469 1154
rect 3377 1110 3407 1124
rect 3434 1120 3469 1128
rect 3434 1110 3435 1120
rect 3450 1110 3463 1120
rect -3 1104 3469 1110
rect -2 1096 3469 1104
rect 5889 1154 5930 1162
rect 5889 1128 5904 1154
rect 5911 1128 5930 1154
rect 5994 1150 6056 1162
rect 6068 1150 6143 1162
rect 6201 1150 6276 1162
rect 6288 1150 6319 1162
rect 6325 1150 6360 1162
rect 5994 1148 6156 1150
rect 5889 1120 5930 1128
rect 6012 1124 6025 1148
rect 6040 1146 6055 1148
rect 5895 1110 5896 1120
rect 5911 1110 5924 1120
rect 5939 1110 5969 1124
rect 6012 1110 6055 1124
rect 6079 1121 6086 1128
rect 6089 1124 6156 1148
rect 6188 1148 6360 1150
rect 6158 1126 6186 1130
rect 6188 1126 6268 1148
rect 6289 1146 6304 1148
rect 6158 1124 6268 1126
rect 6089 1120 6268 1124
rect 6062 1110 6092 1120
rect 6094 1110 6247 1120
rect 6255 1110 6285 1120
rect 6289 1110 6319 1124
rect 6347 1110 6360 1148
rect 6432 1154 6467 1162
rect 6432 1128 6433 1154
rect 6440 1128 6467 1154
rect 6375 1110 6405 1124
rect 6432 1120 6467 1128
rect 6469 1154 6510 1162
rect 6469 1128 6484 1154
rect 6491 1128 6510 1154
rect 6574 1150 6636 1162
rect 6648 1150 6723 1162
rect 6781 1150 6856 1162
rect 6868 1150 6899 1162
rect 6905 1150 6940 1162
rect 6574 1148 6736 1150
rect 6469 1120 6510 1128
rect 6592 1124 6605 1148
rect 6620 1146 6635 1148
rect 6432 1110 6433 1120
rect 6448 1110 6461 1120
rect 6475 1110 6476 1120
rect 6491 1110 6504 1120
rect 6519 1110 6549 1124
rect 6592 1110 6635 1124
rect 6659 1121 6666 1128
rect 6669 1124 6736 1148
rect 6768 1148 6940 1150
rect 6738 1126 6766 1130
rect 6768 1126 6848 1148
rect 6869 1146 6884 1148
rect 6738 1124 6848 1126
rect 6669 1120 6848 1124
rect 6642 1110 6672 1120
rect 6674 1110 6827 1120
rect 6835 1110 6865 1120
rect 6869 1110 6899 1124
rect 6927 1110 6940 1148
rect 7012 1154 7047 1162
rect 7012 1128 7013 1154
rect 7020 1128 7047 1154
rect 6955 1110 6985 1124
rect 7012 1120 7047 1128
rect 7049 1154 7090 1162
rect 7049 1128 7064 1154
rect 7071 1128 7090 1154
rect 7154 1150 7216 1162
rect 7228 1150 7303 1162
rect 7361 1150 7436 1162
rect 7448 1150 7479 1162
rect 7485 1150 7520 1162
rect 7154 1148 7316 1150
rect 7049 1120 7090 1128
rect 7172 1124 7185 1148
rect 7200 1146 7215 1148
rect 7012 1110 7013 1120
rect 7028 1110 7041 1120
rect 7055 1110 7056 1120
rect 7071 1110 7084 1120
rect 7099 1110 7129 1124
rect 7172 1110 7215 1124
rect 7239 1121 7246 1128
rect 7249 1124 7316 1148
rect 7348 1148 7520 1150
rect 7318 1126 7346 1130
rect 7348 1126 7428 1148
rect 7449 1146 7464 1148
rect 7318 1124 7428 1126
rect 7249 1120 7428 1124
rect 7222 1110 7252 1120
rect 7254 1110 7407 1120
rect 7415 1110 7445 1120
rect 7449 1110 7479 1124
rect 7507 1110 7520 1148
rect 7592 1154 7627 1162
rect 7592 1128 7593 1154
rect 7600 1128 7627 1154
rect 7535 1110 7565 1124
rect 7592 1120 7627 1128
rect 7629 1154 7670 1162
rect 7629 1128 7644 1154
rect 7651 1128 7670 1154
rect 7734 1150 7796 1162
rect 7808 1150 7883 1162
rect 7941 1150 8016 1162
rect 8028 1150 8059 1162
rect 8065 1150 8100 1162
rect 7734 1148 7896 1150
rect 7629 1120 7670 1128
rect 7752 1124 7765 1148
rect 7780 1146 7795 1148
rect 7592 1110 7593 1120
rect 7608 1110 7621 1120
rect 7635 1110 7636 1120
rect 7651 1110 7664 1120
rect 7679 1110 7709 1124
rect 7752 1110 7795 1124
rect 7819 1121 7826 1128
rect 7829 1124 7896 1148
rect 7928 1148 8100 1150
rect 7898 1126 7926 1130
rect 7928 1126 8008 1148
rect 8029 1146 8044 1148
rect 7898 1124 8008 1126
rect 7829 1120 8008 1124
rect 7802 1110 7832 1120
rect 7834 1110 7987 1120
rect 7995 1110 8025 1120
rect 8029 1110 8059 1124
rect 8087 1110 8100 1148
rect 8172 1154 8207 1162
rect 8172 1128 8173 1154
rect 8180 1128 8207 1154
rect 8115 1110 8145 1124
rect 8172 1120 8207 1128
rect 8209 1154 8250 1162
rect 8209 1128 8224 1154
rect 8231 1128 8250 1154
rect 8314 1150 8376 1162
rect 8388 1150 8463 1162
rect 8521 1150 8596 1162
rect 8608 1150 8639 1162
rect 8645 1150 8680 1162
rect 8314 1148 8476 1150
rect 8209 1120 8250 1128
rect 8332 1124 8345 1148
rect 8360 1146 8375 1148
rect 8172 1110 8173 1120
rect 8188 1110 8201 1120
rect 8215 1110 8216 1120
rect 8231 1110 8244 1120
rect 8259 1110 8289 1124
rect 8332 1110 8375 1124
rect 8399 1121 8406 1128
rect 8409 1124 8476 1148
rect 8508 1148 8680 1150
rect 8478 1126 8506 1130
rect 8508 1126 8588 1148
rect 8609 1146 8624 1148
rect 8478 1124 8588 1126
rect 8409 1120 8588 1124
rect 8382 1110 8412 1120
rect 8414 1110 8567 1120
rect 8575 1110 8605 1120
rect 8609 1110 8639 1124
rect 8667 1110 8680 1148
rect 8752 1154 8787 1162
rect 8752 1128 8753 1154
rect 8760 1128 8787 1154
rect 8695 1110 8725 1124
rect 8752 1120 8787 1128
rect 8789 1154 8830 1162
rect 8789 1128 8804 1154
rect 8811 1128 8830 1154
rect 8894 1150 8956 1162
rect 8968 1150 9043 1162
rect 9101 1150 9176 1162
rect 9188 1150 9219 1162
rect 9225 1150 9260 1162
rect 8894 1148 9056 1150
rect 8789 1120 8830 1128
rect 8912 1124 8925 1148
rect 8940 1146 8955 1148
rect 8752 1110 8753 1120
rect 8768 1110 8781 1120
rect 8795 1110 8796 1120
rect 8811 1110 8824 1120
rect 8839 1110 8869 1124
rect 8912 1110 8955 1124
rect 8979 1121 8986 1128
rect 8989 1124 9056 1148
rect 9088 1148 9260 1150
rect 9058 1126 9086 1130
rect 9088 1126 9168 1148
rect 9189 1146 9204 1148
rect 9058 1124 9168 1126
rect 8989 1120 9168 1124
rect 8962 1110 8992 1120
rect 8994 1110 9147 1120
rect 9155 1110 9185 1120
rect 9189 1110 9219 1124
rect 9247 1110 9260 1148
rect 9332 1154 9367 1162
rect 9332 1128 9333 1154
rect 9340 1128 9367 1154
rect 9275 1110 9305 1124
rect 9332 1120 9367 1128
rect 9332 1110 9333 1120
rect 9348 1110 9361 1120
rect 5889 1096 9361 1110
rect 13 1066 26 1096
rect 41 1078 71 1096
rect 114 1082 128 1096
rect 164 1082 384 1096
rect 115 1080 128 1082
rect 81 1068 96 1080
rect 78 1066 100 1068
rect 105 1066 135 1080
rect 196 1078 349 1082
rect 178 1066 370 1078
rect 413 1066 443 1080
rect 449 1066 462 1096
rect 477 1078 507 1096
rect 550 1066 563 1096
rect 593 1066 606 1096
rect 621 1078 651 1096
rect 694 1082 708 1096
rect 744 1082 964 1096
rect 695 1080 708 1082
rect 661 1068 676 1080
rect 658 1066 680 1068
rect 685 1066 715 1080
rect 776 1078 929 1082
rect 758 1066 950 1078
rect 993 1066 1023 1080
rect 1029 1066 1042 1096
rect 1057 1078 1087 1096
rect 1130 1066 1143 1096
rect 1173 1066 1186 1096
rect 1201 1078 1231 1096
rect 1274 1082 1288 1096
rect 1324 1082 1544 1096
rect 1275 1080 1288 1082
rect 1241 1068 1256 1080
rect 1238 1066 1260 1068
rect 1265 1066 1295 1080
rect 1356 1078 1509 1082
rect 1338 1066 1530 1078
rect 1573 1066 1603 1080
rect 1609 1066 1622 1096
rect 1637 1078 1667 1096
rect 1710 1066 1723 1096
rect 1753 1066 1766 1096
rect 1781 1078 1811 1096
rect 1854 1082 1868 1096
rect 1904 1082 2124 1096
rect 1855 1080 1868 1082
rect 1821 1068 1836 1080
rect 1818 1066 1840 1068
rect 1845 1066 1875 1080
rect 1936 1078 2089 1082
rect 1918 1066 2110 1078
rect 2153 1066 2183 1080
rect 2189 1066 2202 1096
rect 2217 1078 2247 1096
rect 2290 1066 2303 1096
rect 2333 1066 2346 1096
rect 2361 1078 2391 1096
rect 2434 1082 2448 1096
rect 2484 1082 2704 1096
rect 2435 1080 2448 1082
rect 2401 1068 2416 1080
rect 2398 1066 2420 1068
rect 2425 1066 2455 1080
rect 2516 1078 2669 1082
rect 2498 1066 2690 1078
rect 2733 1066 2763 1080
rect 2769 1066 2782 1096
rect 2797 1078 2827 1096
rect 2870 1066 2883 1096
rect 2913 1066 2926 1096
rect 2941 1078 2971 1096
rect 3014 1082 3028 1096
rect 3064 1082 3284 1096
rect 3015 1080 3028 1082
rect 2981 1068 2996 1080
rect 2978 1066 3000 1068
rect 3005 1066 3035 1080
rect 3096 1078 3249 1082
rect 3078 1066 3270 1078
rect 3313 1066 3343 1080
rect 3349 1066 3362 1096
rect 3377 1078 3407 1096
rect 3450 1066 3463 1096
rect 5911 1066 5924 1096
rect 5939 1078 5969 1096
rect 6012 1082 6026 1096
rect 6062 1082 6282 1096
rect 6013 1080 6026 1082
rect 5979 1068 5994 1080
rect 5976 1066 5998 1068
rect 6003 1066 6033 1080
rect 6094 1078 6247 1082
rect 6076 1066 6268 1078
rect 6311 1066 6341 1080
rect 6347 1066 6360 1096
rect 6375 1078 6405 1096
rect 6448 1066 6461 1096
rect 6491 1066 6504 1096
rect 6519 1078 6549 1096
rect 6592 1082 6606 1096
rect 6642 1082 6862 1096
rect 6593 1080 6606 1082
rect 6559 1068 6574 1080
rect 6556 1066 6578 1068
rect 6583 1066 6613 1080
rect 6674 1078 6827 1082
rect 6656 1066 6848 1078
rect 6891 1066 6921 1080
rect 6927 1066 6940 1096
rect 6955 1078 6985 1096
rect 7028 1066 7041 1096
rect 7071 1066 7084 1096
rect 7099 1078 7129 1096
rect 7172 1082 7186 1096
rect 7222 1082 7442 1096
rect 7173 1080 7186 1082
rect 7139 1068 7154 1080
rect 7136 1066 7158 1068
rect 7163 1066 7193 1080
rect 7254 1078 7407 1082
rect 7236 1066 7428 1078
rect 7471 1066 7501 1080
rect 7507 1066 7520 1096
rect 7535 1078 7565 1096
rect 7608 1066 7621 1096
rect 7651 1066 7664 1096
rect 7679 1078 7709 1096
rect 7752 1082 7766 1096
rect 7802 1082 8022 1096
rect 7753 1080 7766 1082
rect 7719 1068 7734 1080
rect 7716 1066 7738 1068
rect 7743 1066 7773 1080
rect 7834 1078 7987 1082
rect 7816 1066 8008 1078
rect 8051 1066 8081 1080
rect 8087 1066 8100 1096
rect 8115 1078 8145 1096
rect 8188 1066 8201 1096
rect 8231 1066 8244 1096
rect 8259 1078 8289 1096
rect 8332 1082 8346 1096
rect 8382 1082 8602 1096
rect 8333 1080 8346 1082
rect 8299 1068 8314 1080
rect 8296 1066 8318 1068
rect 8323 1066 8353 1080
rect 8414 1078 8567 1082
rect 8396 1066 8588 1078
rect 8631 1066 8661 1080
rect 8667 1066 8680 1096
rect 8695 1078 8725 1096
rect 8768 1066 8781 1096
rect 8811 1066 8824 1096
rect 8839 1078 8869 1096
rect 8912 1082 8926 1096
rect 8962 1082 9182 1096
rect 8913 1080 8926 1082
rect 8879 1068 8894 1080
rect 8876 1066 8898 1068
rect 8903 1066 8933 1080
rect 8994 1078 9147 1082
rect 8976 1066 9168 1078
rect 9211 1066 9241 1080
rect 9247 1066 9260 1096
rect 9275 1078 9305 1096
rect 9348 1066 9361 1096
rect -2 1052 3469 1066
rect 5889 1052 9361 1066
rect 13 948 26 1052
rect 71 1030 72 1040
rect 87 1030 100 1040
rect 71 1026 100 1030
rect 105 1026 135 1052
rect 153 1038 169 1040
rect 241 1038 294 1052
rect 242 1036 306 1038
rect 349 1036 364 1052
rect 413 1049 443 1052
rect 413 1046 449 1049
rect 379 1038 395 1040
rect 153 1026 168 1030
rect 71 1024 168 1026
rect 196 1024 364 1036
rect 380 1026 395 1030
rect 413 1027 452 1046
rect 471 1040 478 1041
rect 477 1033 478 1040
rect 461 1030 462 1033
rect 477 1030 490 1033
rect 413 1026 443 1027
rect 452 1026 458 1027
rect 461 1026 490 1030
rect 380 1025 490 1026
rect 380 1024 496 1025
rect 55 1016 106 1024
rect 55 1004 80 1016
rect 87 1004 106 1016
rect 137 1016 187 1024
rect 137 1008 153 1016
rect 160 1014 187 1016
rect 196 1014 417 1024
rect 160 1004 417 1014
rect 446 1016 496 1024
rect 446 1007 462 1016
rect 55 996 106 1004
rect 153 996 417 1004
rect 443 1004 462 1007
rect 469 1004 496 1016
rect 443 996 496 1004
rect 71 988 72 996
rect 87 988 100 996
rect 71 980 87 988
rect 68 973 87 976
rect 68 964 90 973
rect 41 954 90 964
rect 41 948 71 954
rect 90 949 95 954
rect 13 932 87 948
rect 105 940 135 996
rect 170 986 378 996
rect 413 992 458 996
rect 461 995 462 996
rect 477 995 490 996
rect 196 956 385 986
rect 211 953 385 956
rect 204 950 385 953
rect 13 930 26 932
rect 41 930 75 932
rect 13 914 87 930
rect 114 926 127 940
rect 142 926 158 942
rect 204 937 215 950
rect -3 892 -2 908
rect 13 892 26 914
rect 41 892 71 914
rect 114 910 176 926
rect 204 919 215 935
rect 220 930 230 950
rect 240 930 254 950
rect 257 937 266 950
rect 282 937 291 950
rect 220 919 254 930
rect 257 919 266 935
rect 282 919 291 935
rect 298 930 308 950
rect 318 930 332 950
rect 333 937 344 950
rect 298 919 332 930
rect 333 919 344 935
rect 390 926 406 942
rect 413 940 443 992
rect 477 988 478 995
rect 462 980 478 988
rect 449 948 462 967
rect 477 948 507 964
rect 449 932 523 948
rect 449 930 462 932
rect 477 930 511 932
rect 114 908 127 910
rect 142 908 176 910
rect 114 892 176 908
rect 220 903 236 906
rect 298 903 328 914
rect 376 910 422 926
rect 449 914 523 930
rect 376 908 410 910
rect 375 892 422 908
rect 449 892 462 914
rect 477 892 507 914
rect 534 892 535 908
rect 550 892 563 1052
rect 593 948 606 1052
rect 651 1030 652 1040
rect 667 1030 680 1040
rect 651 1026 680 1030
rect 685 1026 715 1052
rect 733 1038 749 1040
rect 821 1038 874 1052
rect 822 1036 886 1038
rect 929 1036 944 1052
rect 993 1049 1023 1052
rect 993 1046 1029 1049
rect 959 1038 975 1040
rect 733 1026 748 1030
rect 651 1024 748 1026
rect 776 1024 944 1036
rect 960 1026 975 1030
rect 993 1027 1032 1046
rect 1051 1040 1058 1041
rect 1057 1033 1058 1040
rect 1041 1030 1042 1033
rect 1057 1030 1070 1033
rect 993 1026 1023 1027
rect 1032 1026 1038 1027
rect 1041 1026 1070 1030
rect 960 1025 1070 1026
rect 960 1024 1076 1025
rect 635 1016 686 1024
rect 635 1004 660 1016
rect 667 1004 686 1016
rect 717 1016 767 1024
rect 717 1008 733 1016
rect 740 1014 767 1016
rect 776 1014 997 1024
rect 740 1004 997 1014
rect 1026 1016 1076 1024
rect 1026 1007 1042 1016
rect 635 996 686 1004
rect 733 996 997 1004
rect 1023 1004 1042 1007
rect 1049 1004 1076 1016
rect 1023 996 1076 1004
rect 651 988 652 996
rect 667 988 680 996
rect 651 980 667 988
rect 648 973 667 976
rect 648 964 670 973
rect 621 954 670 964
rect 621 948 651 954
rect 670 949 675 954
rect 593 932 667 948
rect 685 940 715 996
rect 750 986 958 996
rect 993 992 1038 996
rect 1041 995 1042 996
rect 1057 995 1070 996
rect 776 956 965 986
rect 791 953 965 956
rect 784 950 965 953
rect 593 930 606 932
rect 621 930 655 932
rect 593 914 667 930
rect 694 926 707 940
rect 722 926 738 942
rect 784 937 795 950
rect 577 892 578 908
rect 593 892 606 914
rect 621 892 651 914
rect 694 910 756 926
rect 784 919 795 935
rect 800 930 810 950
rect 820 930 834 950
rect 837 937 846 950
rect 862 937 871 950
rect 800 919 834 930
rect 837 919 846 935
rect 862 919 871 935
rect 878 930 888 950
rect 898 930 912 950
rect 913 937 924 950
rect 878 919 912 930
rect 913 919 924 935
rect 970 926 986 942
rect 993 940 1023 992
rect 1057 988 1058 995
rect 1042 980 1058 988
rect 1029 948 1042 967
rect 1057 948 1087 964
rect 1029 932 1103 948
rect 1029 930 1042 932
rect 1057 930 1091 932
rect 694 908 707 910
rect 722 908 756 910
rect 694 892 756 908
rect 800 903 816 906
rect 878 903 908 914
rect 956 910 1002 926
rect 1029 914 1103 930
rect 956 908 990 910
rect 955 892 1002 908
rect 1029 892 1042 914
rect 1057 892 1087 914
rect 1114 892 1115 908
rect 1130 892 1143 1052
rect 1173 948 1186 1052
rect 1231 1030 1232 1040
rect 1247 1030 1260 1040
rect 1231 1026 1260 1030
rect 1265 1026 1295 1052
rect 1313 1038 1329 1040
rect 1401 1038 1454 1052
rect 1402 1036 1466 1038
rect 1509 1036 1524 1052
rect 1573 1049 1603 1052
rect 1573 1046 1609 1049
rect 1539 1038 1555 1040
rect 1313 1026 1328 1030
rect 1231 1024 1328 1026
rect 1356 1024 1524 1036
rect 1540 1026 1555 1030
rect 1573 1027 1612 1046
rect 1631 1040 1638 1041
rect 1637 1033 1638 1040
rect 1621 1030 1622 1033
rect 1637 1030 1650 1033
rect 1573 1026 1603 1027
rect 1612 1026 1618 1027
rect 1621 1026 1650 1030
rect 1540 1025 1650 1026
rect 1540 1024 1656 1025
rect 1215 1016 1266 1024
rect 1215 1004 1240 1016
rect 1247 1004 1266 1016
rect 1297 1016 1347 1024
rect 1297 1008 1313 1016
rect 1320 1014 1347 1016
rect 1356 1014 1577 1024
rect 1320 1004 1577 1014
rect 1606 1016 1656 1024
rect 1606 1007 1622 1016
rect 1215 996 1266 1004
rect 1313 996 1577 1004
rect 1603 1004 1622 1007
rect 1629 1004 1656 1016
rect 1603 996 1656 1004
rect 1231 988 1232 996
rect 1247 988 1260 996
rect 1231 980 1247 988
rect 1228 973 1247 976
rect 1228 964 1250 973
rect 1201 954 1250 964
rect 1201 948 1231 954
rect 1250 949 1255 954
rect 1173 932 1247 948
rect 1265 940 1295 996
rect 1330 986 1538 996
rect 1573 992 1618 996
rect 1621 995 1622 996
rect 1637 995 1650 996
rect 1356 956 1545 986
rect 1371 953 1545 956
rect 1364 950 1545 953
rect 1173 930 1186 932
rect 1201 930 1235 932
rect 1173 914 1247 930
rect 1274 926 1287 940
rect 1302 926 1318 942
rect 1364 937 1375 950
rect 1157 892 1158 908
rect 1173 892 1186 914
rect 1201 892 1231 914
rect 1274 910 1336 926
rect 1364 919 1375 935
rect 1380 930 1390 950
rect 1400 930 1414 950
rect 1417 937 1426 950
rect 1442 937 1451 950
rect 1380 919 1414 930
rect 1417 919 1426 935
rect 1442 919 1451 935
rect 1458 930 1468 950
rect 1478 930 1492 950
rect 1493 937 1504 950
rect 1458 919 1492 930
rect 1493 919 1504 935
rect 1550 926 1566 942
rect 1573 940 1603 992
rect 1637 988 1638 995
rect 1622 980 1638 988
rect 1609 948 1622 967
rect 1637 948 1667 964
rect 1609 932 1683 948
rect 1609 930 1622 932
rect 1637 930 1671 932
rect 1274 908 1287 910
rect 1302 908 1336 910
rect 1274 892 1336 908
rect 1380 903 1396 906
rect 1458 903 1488 914
rect 1536 910 1582 926
rect 1609 914 1683 930
rect 1536 908 1570 910
rect 1535 892 1582 908
rect 1609 892 1622 914
rect 1637 892 1667 914
rect 1694 892 1695 908
rect 1710 892 1723 1052
rect 1753 948 1766 1052
rect 1811 1030 1812 1040
rect 1827 1030 1840 1040
rect 1811 1026 1840 1030
rect 1845 1026 1875 1052
rect 1893 1038 1909 1040
rect 1981 1038 2034 1052
rect 1982 1036 2046 1038
rect 2089 1036 2104 1052
rect 2153 1049 2183 1052
rect 2153 1046 2189 1049
rect 2119 1038 2135 1040
rect 1893 1026 1908 1030
rect 1811 1024 1908 1026
rect 1936 1024 2104 1036
rect 2120 1026 2135 1030
rect 2153 1027 2192 1046
rect 2211 1040 2218 1041
rect 2217 1033 2218 1040
rect 2201 1030 2202 1033
rect 2217 1030 2230 1033
rect 2153 1026 2183 1027
rect 2192 1026 2198 1027
rect 2201 1026 2230 1030
rect 2120 1025 2230 1026
rect 2120 1024 2236 1025
rect 1795 1016 1846 1024
rect 1795 1004 1820 1016
rect 1827 1004 1846 1016
rect 1877 1016 1927 1024
rect 1877 1008 1893 1016
rect 1900 1014 1927 1016
rect 1936 1014 2157 1024
rect 1900 1004 2157 1014
rect 2186 1016 2236 1024
rect 2186 1007 2202 1016
rect 1795 996 1846 1004
rect 1893 996 2157 1004
rect 2183 1004 2202 1007
rect 2209 1004 2236 1016
rect 2183 996 2236 1004
rect 1811 988 1812 996
rect 1827 988 1840 996
rect 1811 980 1827 988
rect 1808 973 1827 976
rect 1808 964 1830 973
rect 1781 954 1830 964
rect 1781 948 1811 954
rect 1830 949 1835 954
rect 1753 932 1827 948
rect 1845 940 1875 996
rect 1910 986 2118 996
rect 2153 992 2198 996
rect 2201 995 2202 996
rect 2217 995 2230 996
rect 1936 956 2125 986
rect 1951 953 2125 956
rect 1944 950 2125 953
rect 1753 930 1766 932
rect 1781 930 1815 932
rect 1753 914 1827 930
rect 1854 926 1867 940
rect 1882 926 1898 942
rect 1944 937 1955 950
rect 1737 892 1738 908
rect 1753 892 1766 914
rect 1781 892 1811 914
rect 1854 910 1916 926
rect 1944 919 1955 935
rect 1960 930 1970 950
rect 1980 930 1994 950
rect 1997 937 2006 950
rect 2022 937 2031 950
rect 1960 919 1994 930
rect 1997 919 2006 935
rect 2022 919 2031 935
rect 2038 930 2048 950
rect 2058 930 2072 950
rect 2073 937 2084 950
rect 2038 919 2072 930
rect 2073 919 2084 935
rect 2130 926 2146 942
rect 2153 940 2183 992
rect 2217 988 2218 995
rect 2202 980 2218 988
rect 2189 948 2202 967
rect 2217 948 2247 964
rect 2189 932 2263 948
rect 2189 930 2202 932
rect 2217 930 2251 932
rect 1854 908 1867 910
rect 1882 908 1916 910
rect 1854 892 1916 908
rect 1960 903 1976 906
rect 2038 903 2068 914
rect 2116 910 2162 926
rect 2189 914 2263 930
rect 2116 908 2150 910
rect 2115 892 2162 908
rect 2189 892 2202 914
rect 2217 892 2247 914
rect 2274 892 2275 908
rect 2290 892 2303 1052
rect 2333 948 2346 1052
rect 2391 1030 2392 1040
rect 2407 1030 2420 1040
rect 2391 1026 2420 1030
rect 2425 1026 2455 1052
rect 2473 1038 2489 1040
rect 2561 1038 2614 1052
rect 2562 1036 2626 1038
rect 2669 1036 2684 1052
rect 2733 1049 2763 1052
rect 2733 1046 2769 1049
rect 2699 1038 2715 1040
rect 2473 1026 2488 1030
rect 2391 1024 2488 1026
rect 2516 1024 2684 1036
rect 2700 1026 2715 1030
rect 2733 1027 2772 1046
rect 2791 1040 2798 1041
rect 2797 1033 2798 1040
rect 2781 1030 2782 1033
rect 2797 1030 2810 1033
rect 2733 1026 2763 1027
rect 2772 1026 2778 1027
rect 2781 1026 2810 1030
rect 2700 1025 2810 1026
rect 2700 1024 2816 1025
rect 2375 1016 2426 1024
rect 2375 1004 2400 1016
rect 2407 1004 2426 1016
rect 2457 1016 2507 1024
rect 2457 1008 2473 1016
rect 2480 1014 2507 1016
rect 2516 1014 2737 1024
rect 2480 1004 2737 1014
rect 2766 1016 2816 1024
rect 2766 1007 2782 1016
rect 2375 996 2426 1004
rect 2473 996 2737 1004
rect 2763 1004 2782 1007
rect 2789 1004 2816 1016
rect 2763 996 2816 1004
rect 2391 988 2392 996
rect 2407 988 2420 996
rect 2391 980 2407 988
rect 2388 973 2407 976
rect 2388 964 2410 973
rect 2361 954 2410 964
rect 2361 948 2391 954
rect 2410 949 2415 954
rect 2333 932 2407 948
rect 2425 940 2455 996
rect 2490 986 2698 996
rect 2733 992 2778 996
rect 2781 995 2782 996
rect 2797 995 2810 996
rect 2516 956 2705 986
rect 2531 953 2705 956
rect 2524 950 2705 953
rect 2333 930 2346 932
rect 2361 930 2395 932
rect 2333 914 2407 930
rect 2434 926 2447 940
rect 2462 926 2478 942
rect 2524 937 2535 950
rect 2317 892 2318 908
rect 2333 892 2346 914
rect 2361 892 2391 914
rect 2434 910 2496 926
rect 2524 919 2535 935
rect 2540 930 2550 950
rect 2560 930 2574 950
rect 2577 937 2586 950
rect 2602 937 2611 950
rect 2540 919 2574 930
rect 2577 919 2586 935
rect 2602 919 2611 935
rect 2618 930 2628 950
rect 2638 930 2652 950
rect 2653 937 2664 950
rect 2618 919 2652 930
rect 2653 919 2664 935
rect 2710 926 2726 942
rect 2733 940 2763 992
rect 2797 988 2798 995
rect 2782 980 2798 988
rect 2769 948 2782 967
rect 2797 948 2827 964
rect 2769 932 2843 948
rect 2769 930 2782 932
rect 2797 930 2831 932
rect 2434 908 2447 910
rect 2462 908 2496 910
rect 2434 892 2496 908
rect 2540 903 2556 906
rect 2618 903 2648 914
rect 2696 910 2742 926
rect 2769 914 2843 930
rect 2696 908 2730 910
rect 2695 892 2742 908
rect 2769 892 2782 914
rect 2797 892 2827 914
rect 2854 892 2855 908
rect 2870 892 2883 1052
rect 2913 948 2926 1052
rect 2971 1030 2972 1040
rect 2987 1030 3000 1040
rect 2971 1026 3000 1030
rect 3005 1026 3035 1052
rect 3053 1038 3069 1040
rect 3141 1038 3194 1052
rect 3142 1036 3206 1038
rect 3249 1036 3264 1052
rect 3313 1049 3343 1052
rect 3313 1046 3349 1049
rect 3279 1038 3295 1040
rect 3053 1026 3068 1030
rect 2971 1024 3068 1026
rect 3096 1024 3264 1036
rect 3280 1026 3295 1030
rect 3313 1027 3352 1046
rect 3371 1040 3378 1041
rect 3377 1033 3378 1040
rect 3361 1030 3362 1033
rect 3377 1030 3390 1033
rect 3313 1026 3343 1027
rect 3352 1026 3358 1027
rect 3361 1026 3390 1030
rect 3280 1025 3390 1026
rect 3280 1024 3396 1025
rect 2955 1016 3006 1024
rect 2955 1004 2980 1016
rect 2987 1004 3006 1016
rect 3037 1016 3087 1024
rect 3037 1008 3053 1016
rect 3060 1014 3087 1016
rect 3096 1014 3317 1024
rect 3060 1004 3317 1014
rect 3346 1016 3396 1024
rect 3346 1007 3362 1016
rect 2955 996 3006 1004
rect 3053 996 3317 1004
rect 3343 1004 3362 1007
rect 3369 1004 3396 1016
rect 3343 996 3396 1004
rect 2971 988 2972 996
rect 2987 988 3000 996
rect 2971 980 2987 988
rect 2968 973 2987 976
rect 2968 964 2990 973
rect 2941 954 2990 964
rect 2941 948 2971 954
rect 2990 949 2995 954
rect 2913 932 2987 948
rect 3005 940 3035 996
rect 3070 986 3278 996
rect 3313 992 3358 996
rect 3361 995 3362 996
rect 3377 995 3390 996
rect 3096 956 3285 986
rect 3111 953 3285 956
rect 3104 950 3285 953
rect 2913 930 2926 932
rect 2941 930 2975 932
rect 2913 914 2987 930
rect 3014 926 3027 940
rect 3042 926 3058 942
rect 3104 937 3115 950
rect 2897 892 2898 908
rect 2913 892 2926 914
rect 2941 892 2971 914
rect 3014 910 3076 926
rect 3104 919 3115 935
rect 3120 930 3130 950
rect 3140 930 3154 950
rect 3157 937 3166 950
rect 3182 937 3191 950
rect 3120 919 3154 930
rect 3157 919 3166 935
rect 3182 919 3191 935
rect 3198 930 3208 950
rect 3218 930 3232 950
rect 3233 937 3244 950
rect 3198 919 3232 930
rect 3233 919 3244 935
rect 3290 926 3306 942
rect 3313 940 3343 992
rect 3377 988 3378 995
rect 3362 980 3378 988
rect 3349 948 3362 967
rect 3377 948 3407 964
rect 3349 932 3423 948
rect 3349 930 3362 932
rect 3377 930 3411 932
rect 3014 908 3027 910
rect 3042 908 3076 910
rect 3014 892 3076 908
rect 3120 903 3136 906
rect 3198 903 3228 914
rect 3276 910 3322 926
rect 3349 914 3423 930
rect 3276 908 3310 910
rect 3275 892 3322 908
rect 3349 892 3362 914
rect 3377 892 3407 914
rect 3434 892 3435 908
rect 3450 892 3463 1052
rect 5911 948 5924 1052
rect 5969 1030 5970 1040
rect 5985 1030 5998 1040
rect 5969 1026 5998 1030
rect 6003 1026 6033 1052
rect 6051 1038 6067 1040
rect 6139 1038 6192 1052
rect 6140 1036 6204 1038
rect 6247 1036 6262 1052
rect 6311 1049 6341 1052
rect 6311 1046 6347 1049
rect 6277 1038 6293 1040
rect 6051 1026 6066 1030
rect 5969 1024 6066 1026
rect 6094 1024 6262 1036
rect 6278 1026 6293 1030
rect 6311 1027 6350 1046
rect 6369 1040 6376 1041
rect 6375 1033 6376 1040
rect 6359 1030 6360 1033
rect 6375 1030 6388 1033
rect 6311 1026 6341 1027
rect 6350 1026 6356 1027
rect 6359 1026 6388 1030
rect 6278 1025 6388 1026
rect 6278 1024 6394 1025
rect 5953 1016 6004 1024
rect 5953 1004 5978 1016
rect 5985 1004 6004 1016
rect 6035 1016 6085 1024
rect 6035 1008 6051 1016
rect 6058 1014 6085 1016
rect 6094 1014 6315 1024
rect 6058 1004 6315 1014
rect 6344 1016 6394 1024
rect 6344 1007 6360 1016
rect 5953 996 6004 1004
rect 6051 996 6315 1004
rect 6341 1004 6360 1007
rect 6367 1004 6394 1016
rect 6341 996 6394 1004
rect 5969 988 5970 996
rect 5985 988 5998 996
rect 5969 980 5985 988
rect 5966 973 5985 976
rect 5966 964 5988 973
rect 5939 954 5988 964
rect 5939 948 5969 954
rect 5988 949 5993 954
rect 5911 932 5985 948
rect 6003 940 6033 996
rect 6068 986 6276 996
rect 6311 992 6356 996
rect 6359 995 6360 996
rect 6375 995 6388 996
rect 6094 956 6283 986
rect 6109 953 6283 956
rect 6102 950 6283 953
rect 5911 930 5924 932
rect 5939 930 5973 932
rect 5911 914 5985 930
rect 6012 926 6025 940
rect 6040 926 6056 942
rect 6102 937 6113 950
rect 5895 892 5896 908
rect 5911 892 5924 914
rect 5939 892 5969 914
rect 6012 910 6074 926
rect 6102 919 6113 935
rect 6118 930 6128 950
rect 6138 930 6152 950
rect 6155 937 6164 950
rect 6180 937 6189 950
rect 6118 919 6152 930
rect 6155 919 6164 935
rect 6180 919 6189 935
rect 6196 930 6206 950
rect 6216 930 6230 950
rect 6231 937 6242 950
rect 6196 919 6230 930
rect 6231 919 6242 935
rect 6288 926 6304 942
rect 6311 940 6341 992
rect 6375 988 6376 995
rect 6360 980 6376 988
rect 6347 948 6360 967
rect 6375 948 6405 964
rect 6347 932 6421 948
rect 6347 930 6360 932
rect 6375 930 6409 932
rect 6012 908 6025 910
rect 6040 908 6074 910
rect 6012 892 6074 908
rect 6118 903 6134 906
rect 6196 903 6226 914
rect 6274 910 6320 926
rect 6347 914 6421 930
rect 6274 908 6308 910
rect 6273 892 6320 908
rect 6347 892 6360 914
rect 6375 892 6405 914
rect 6432 892 6433 908
rect 6448 892 6461 1052
rect 6491 948 6504 1052
rect 6549 1030 6550 1040
rect 6565 1030 6578 1040
rect 6549 1026 6578 1030
rect 6583 1026 6613 1052
rect 6631 1038 6647 1040
rect 6719 1038 6772 1052
rect 6720 1036 6784 1038
rect 6827 1036 6842 1052
rect 6891 1049 6921 1052
rect 6891 1046 6927 1049
rect 6857 1038 6873 1040
rect 6631 1026 6646 1030
rect 6549 1024 6646 1026
rect 6674 1024 6842 1036
rect 6858 1026 6873 1030
rect 6891 1027 6930 1046
rect 6949 1040 6956 1041
rect 6955 1033 6956 1040
rect 6939 1030 6940 1033
rect 6955 1030 6968 1033
rect 6891 1026 6921 1027
rect 6930 1026 6936 1027
rect 6939 1026 6968 1030
rect 6858 1025 6968 1026
rect 6858 1024 6974 1025
rect 6533 1016 6584 1024
rect 6533 1004 6558 1016
rect 6565 1004 6584 1016
rect 6615 1016 6665 1024
rect 6615 1008 6631 1016
rect 6638 1014 6665 1016
rect 6674 1014 6895 1024
rect 6638 1004 6895 1014
rect 6924 1016 6974 1024
rect 6924 1007 6940 1016
rect 6533 996 6584 1004
rect 6631 996 6895 1004
rect 6921 1004 6940 1007
rect 6947 1004 6974 1016
rect 6921 996 6974 1004
rect 6549 988 6550 996
rect 6565 988 6578 996
rect 6549 980 6565 988
rect 6546 973 6565 976
rect 6546 964 6568 973
rect 6519 954 6568 964
rect 6519 948 6549 954
rect 6568 949 6573 954
rect 6491 932 6565 948
rect 6583 940 6613 996
rect 6648 986 6856 996
rect 6891 992 6936 996
rect 6939 995 6940 996
rect 6955 995 6968 996
rect 6674 956 6863 986
rect 6689 953 6863 956
rect 6682 950 6863 953
rect 6491 930 6504 932
rect 6519 930 6553 932
rect 6491 914 6565 930
rect 6592 926 6605 940
rect 6620 926 6636 942
rect 6682 937 6693 950
rect 6475 892 6476 908
rect 6491 892 6504 914
rect 6519 892 6549 914
rect 6592 910 6654 926
rect 6682 919 6693 935
rect 6698 930 6708 950
rect 6718 930 6732 950
rect 6735 937 6744 950
rect 6760 937 6769 950
rect 6698 919 6732 930
rect 6735 919 6744 935
rect 6760 919 6769 935
rect 6776 930 6786 950
rect 6796 930 6810 950
rect 6811 937 6822 950
rect 6776 919 6810 930
rect 6811 919 6822 935
rect 6868 926 6884 942
rect 6891 940 6921 992
rect 6955 988 6956 995
rect 6940 980 6956 988
rect 6927 948 6940 967
rect 6955 948 6985 964
rect 6927 932 7001 948
rect 6927 930 6940 932
rect 6955 930 6989 932
rect 6592 908 6605 910
rect 6620 908 6654 910
rect 6592 892 6654 908
rect 6698 903 6714 906
rect 6776 903 6806 914
rect 6854 910 6900 926
rect 6927 914 7001 930
rect 6854 908 6888 910
rect 6853 892 6900 908
rect 6927 892 6940 914
rect 6955 892 6985 914
rect 7012 892 7013 908
rect 7028 892 7041 1052
rect 7071 948 7084 1052
rect 7129 1030 7130 1040
rect 7145 1030 7158 1040
rect 7129 1026 7158 1030
rect 7163 1026 7193 1052
rect 7211 1038 7227 1040
rect 7299 1038 7352 1052
rect 7300 1036 7364 1038
rect 7407 1036 7422 1052
rect 7471 1049 7501 1052
rect 7471 1046 7507 1049
rect 7437 1038 7453 1040
rect 7211 1026 7226 1030
rect 7129 1024 7226 1026
rect 7254 1024 7422 1036
rect 7438 1026 7453 1030
rect 7471 1027 7510 1046
rect 7529 1040 7536 1041
rect 7535 1033 7536 1040
rect 7519 1030 7520 1033
rect 7535 1030 7548 1033
rect 7471 1026 7501 1027
rect 7510 1026 7516 1027
rect 7519 1026 7548 1030
rect 7438 1025 7548 1026
rect 7438 1024 7554 1025
rect 7113 1016 7164 1024
rect 7113 1004 7138 1016
rect 7145 1004 7164 1016
rect 7195 1016 7245 1024
rect 7195 1008 7211 1016
rect 7218 1014 7245 1016
rect 7254 1014 7475 1024
rect 7218 1004 7475 1014
rect 7504 1016 7554 1024
rect 7504 1007 7520 1016
rect 7113 996 7164 1004
rect 7211 996 7475 1004
rect 7501 1004 7520 1007
rect 7527 1004 7554 1016
rect 7501 996 7554 1004
rect 7129 988 7130 996
rect 7145 988 7158 996
rect 7129 980 7145 988
rect 7126 973 7145 976
rect 7126 964 7148 973
rect 7099 954 7148 964
rect 7099 948 7129 954
rect 7148 949 7153 954
rect 7071 932 7145 948
rect 7163 940 7193 996
rect 7228 986 7436 996
rect 7471 992 7516 996
rect 7519 995 7520 996
rect 7535 995 7548 996
rect 7254 956 7443 986
rect 7269 953 7443 956
rect 7262 950 7443 953
rect 7071 930 7084 932
rect 7099 930 7133 932
rect 7071 914 7145 930
rect 7172 926 7185 940
rect 7200 926 7216 942
rect 7262 937 7273 950
rect 7055 892 7056 908
rect 7071 892 7084 914
rect 7099 892 7129 914
rect 7172 910 7234 926
rect 7262 919 7273 935
rect 7278 930 7288 950
rect 7298 930 7312 950
rect 7315 937 7324 950
rect 7340 937 7349 950
rect 7278 919 7312 930
rect 7315 919 7324 935
rect 7340 919 7349 935
rect 7356 930 7366 950
rect 7376 930 7390 950
rect 7391 937 7402 950
rect 7356 919 7390 930
rect 7391 919 7402 935
rect 7448 926 7464 942
rect 7471 940 7501 992
rect 7535 988 7536 995
rect 7520 980 7536 988
rect 7507 948 7520 967
rect 7535 948 7565 964
rect 7507 932 7581 948
rect 7507 930 7520 932
rect 7535 930 7569 932
rect 7172 908 7185 910
rect 7200 908 7234 910
rect 7172 892 7234 908
rect 7278 903 7294 906
rect 7356 903 7386 914
rect 7434 910 7480 926
rect 7507 914 7581 930
rect 7434 908 7468 910
rect 7433 892 7480 908
rect 7507 892 7520 914
rect 7535 892 7565 914
rect 7592 892 7593 908
rect 7608 892 7621 1052
rect 7651 948 7664 1052
rect 7709 1030 7710 1040
rect 7725 1030 7738 1040
rect 7709 1026 7738 1030
rect 7743 1026 7773 1052
rect 7791 1038 7807 1040
rect 7879 1038 7932 1052
rect 7880 1036 7944 1038
rect 7987 1036 8002 1052
rect 8051 1049 8081 1052
rect 8051 1046 8087 1049
rect 8017 1038 8033 1040
rect 7791 1026 7806 1030
rect 7709 1024 7806 1026
rect 7834 1024 8002 1036
rect 8018 1026 8033 1030
rect 8051 1027 8090 1046
rect 8109 1040 8116 1041
rect 8115 1033 8116 1040
rect 8099 1030 8100 1033
rect 8115 1030 8128 1033
rect 8051 1026 8081 1027
rect 8090 1026 8096 1027
rect 8099 1026 8128 1030
rect 8018 1025 8128 1026
rect 8018 1024 8134 1025
rect 7693 1016 7744 1024
rect 7693 1004 7718 1016
rect 7725 1004 7744 1016
rect 7775 1016 7825 1024
rect 7775 1008 7791 1016
rect 7798 1014 7825 1016
rect 7834 1014 8055 1024
rect 7798 1004 8055 1014
rect 8084 1016 8134 1024
rect 8084 1007 8100 1016
rect 7693 996 7744 1004
rect 7791 996 8055 1004
rect 8081 1004 8100 1007
rect 8107 1004 8134 1016
rect 8081 996 8134 1004
rect 7709 988 7710 996
rect 7725 988 7738 996
rect 7709 980 7725 988
rect 7706 973 7725 976
rect 7706 964 7728 973
rect 7679 954 7728 964
rect 7679 948 7709 954
rect 7728 949 7733 954
rect 7651 932 7725 948
rect 7743 940 7773 996
rect 7808 986 8016 996
rect 8051 992 8096 996
rect 8099 995 8100 996
rect 8115 995 8128 996
rect 7834 956 8023 986
rect 7849 953 8023 956
rect 7842 950 8023 953
rect 7651 930 7664 932
rect 7679 930 7713 932
rect 7651 914 7725 930
rect 7752 926 7765 940
rect 7780 926 7796 942
rect 7842 937 7853 950
rect 7635 892 7636 908
rect 7651 892 7664 914
rect 7679 892 7709 914
rect 7752 910 7814 926
rect 7842 919 7853 935
rect 7858 930 7868 950
rect 7878 930 7892 950
rect 7895 937 7904 950
rect 7920 937 7929 950
rect 7858 919 7892 930
rect 7895 919 7904 935
rect 7920 919 7929 935
rect 7936 930 7946 950
rect 7956 930 7970 950
rect 7971 937 7982 950
rect 7936 919 7970 930
rect 7971 919 7982 935
rect 8028 926 8044 942
rect 8051 940 8081 992
rect 8115 988 8116 995
rect 8100 980 8116 988
rect 8087 948 8100 967
rect 8115 948 8145 964
rect 8087 932 8161 948
rect 8087 930 8100 932
rect 8115 930 8149 932
rect 7752 908 7765 910
rect 7780 908 7814 910
rect 7752 892 7814 908
rect 7858 903 7874 906
rect 7936 903 7966 914
rect 8014 910 8060 926
rect 8087 914 8161 930
rect 8014 908 8048 910
rect 8013 892 8060 908
rect 8087 892 8100 914
rect 8115 892 8145 914
rect 8172 892 8173 908
rect 8188 892 8201 1052
rect 8231 948 8244 1052
rect 8289 1030 8290 1040
rect 8305 1030 8318 1040
rect 8289 1026 8318 1030
rect 8323 1026 8353 1052
rect 8371 1038 8387 1040
rect 8459 1038 8512 1052
rect 8460 1036 8524 1038
rect 8567 1036 8582 1052
rect 8631 1049 8661 1052
rect 8631 1046 8667 1049
rect 8597 1038 8613 1040
rect 8371 1026 8386 1030
rect 8289 1024 8386 1026
rect 8414 1024 8582 1036
rect 8598 1026 8613 1030
rect 8631 1027 8670 1046
rect 8689 1040 8696 1041
rect 8695 1033 8696 1040
rect 8679 1030 8680 1033
rect 8695 1030 8708 1033
rect 8631 1026 8661 1027
rect 8670 1026 8676 1027
rect 8679 1026 8708 1030
rect 8598 1025 8708 1026
rect 8598 1024 8714 1025
rect 8273 1016 8324 1024
rect 8273 1004 8298 1016
rect 8305 1004 8324 1016
rect 8355 1016 8405 1024
rect 8355 1008 8371 1016
rect 8378 1014 8405 1016
rect 8414 1014 8635 1024
rect 8378 1004 8635 1014
rect 8664 1016 8714 1024
rect 8664 1007 8680 1016
rect 8273 996 8324 1004
rect 8371 996 8635 1004
rect 8661 1004 8680 1007
rect 8687 1004 8714 1016
rect 8661 996 8714 1004
rect 8289 988 8290 996
rect 8305 988 8318 996
rect 8289 980 8305 988
rect 8286 973 8305 976
rect 8286 964 8308 973
rect 8259 954 8308 964
rect 8259 948 8289 954
rect 8308 949 8313 954
rect 8231 932 8305 948
rect 8323 940 8353 996
rect 8388 986 8596 996
rect 8631 992 8676 996
rect 8679 995 8680 996
rect 8695 995 8708 996
rect 8414 956 8603 986
rect 8429 953 8603 956
rect 8422 950 8603 953
rect 8231 930 8244 932
rect 8259 930 8293 932
rect 8231 914 8305 930
rect 8332 926 8345 940
rect 8360 926 8376 942
rect 8422 937 8433 950
rect 8215 892 8216 908
rect 8231 892 8244 914
rect 8259 892 8289 914
rect 8332 910 8394 926
rect 8422 919 8433 935
rect 8438 930 8448 950
rect 8458 930 8472 950
rect 8475 937 8484 950
rect 8500 937 8509 950
rect 8438 919 8472 930
rect 8475 919 8484 935
rect 8500 919 8509 935
rect 8516 930 8526 950
rect 8536 930 8550 950
rect 8551 937 8562 950
rect 8516 919 8550 930
rect 8551 919 8562 935
rect 8608 926 8624 942
rect 8631 940 8661 992
rect 8695 988 8696 995
rect 8680 980 8696 988
rect 8667 948 8680 967
rect 8695 948 8725 964
rect 8667 932 8741 948
rect 8667 930 8680 932
rect 8695 930 8729 932
rect 8332 908 8345 910
rect 8360 908 8394 910
rect 8332 892 8394 908
rect 8438 903 8454 906
rect 8516 903 8546 914
rect 8594 910 8640 926
rect 8667 914 8741 930
rect 8594 908 8628 910
rect 8593 892 8640 908
rect 8667 892 8680 914
rect 8695 892 8725 914
rect 8752 892 8753 908
rect 8768 892 8781 1052
rect 8811 948 8824 1052
rect 8869 1030 8870 1040
rect 8885 1030 8898 1040
rect 8869 1026 8898 1030
rect 8903 1026 8933 1052
rect 8951 1038 8967 1040
rect 9039 1038 9092 1052
rect 9040 1036 9104 1038
rect 9147 1036 9162 1052
rect 9211 1049 9241 1052
rect 9211 1046 9247 1049
rect 9177 1038 9193 1040
rect 8951 1026 8966 1030
rect 8869 1024 8966 1026
rect 8994 1024 9162 1036
rect 9178 1026 9193 1030
rect 9211 1027 9250 1046
rect 9269 1040 9276 1041
rect 9275 1033 9276 1040
rect 9259 1030 9260 1033
rect 9275 1030 9288 1033
rect 9211 1026 9241 1027
rect 9250 1026 9256 1027
rect 9259 1026 9288 1030
rect 9178 1025 9288 1026
rect 9178 1024 9294 1025
rect 8853 1016 8904 1024
rect 8853 1004 8878 1016
rect 8885 1004 8904 1016
rect 8935 1016 8985 1024
rect 8935 1008 8951 1016
rect 8958 1014 8985 1016
rect 8994 1014 9215 1024
rect 8958 1004 9215 1014
rect 9244 1016 9294 1024
rect 9244 1007 9260 1016
rect 8853 996 8904 1004
rect 8951 996 9215 1004
rect 9241 1004 9260 1007
rect 9267 1004 9294 1016
rect 9241 996 9294 1004
rect 8869 988 8870 996
rect 8885 988 8898 996
rect 8869 980 8885 988
rect 8866 973 8885 976
rect 8866 964 8888 973
rect 8839 954 8888 964
rect 8839 948 8869 954
rect 8888 949 8893 954
rect 8811 932 8885 948
rect 8903 940 8933 996
rect 8968 986 9176 996
rect 9211 992 9256 996
rect 9259 995 9260 996
rect 9275 995 9288 996
rect 8994 956 9183 986
rect 9009 953 9183 956
rect 9002 950 9183 953
rect 8811 930 8824 932
rect 8839 930 8873 932
rect 8811 914 8885 930
rect 8912 926 8925 940
rect 8940 926 8956 942
rect 9002 937 9013 950
rect 8795 892 8796 908
rect 8811 892 8824 914
rect 8839 892 8869 914
rect 8912 910 8974 926
rect 9002 919 9013 935
rect 9018 930 9028 950
rect 9038 930 9052 950
rect 9055 937 9064 950
rect 9080 937 9089 950
rect 9018 919 9052 930
rect 9055 919 9064 935
rect 9080 919 9089 935
rect 9096 930 9106 950
rect 9116 930 9130 950
rect 9131 937 9142 950
rect 9096 919 9130 930
rect 9131 919 9142 935
rect 9188 926 9204 942
rect 9211 940 9241 992
rect 9275 988 9276 995
rect 9260 980 9276 988
rect 9247 948 9260 967
rect 9275 948 9305 964
rect 9247 932 9321 948
rect 9247 930 9260 932
rect 9275 930 9309 932
rect 8912 908 8925 910
rect 8940 908 8974 910
rect 8912 892 8974 908
rect 9018 903 9034 906
rect 9096 903 9126 914
rect 9174 910 9220 926
rect 9247 914 9321 930
rect 9174 908 9208 910
rect 9173 892 9220 908
rect 9247 892 9260 914
rect 9275 892 9305 914
rect 9332 892 9333 908
rect 9348 892 9361 1052
rect -9 884 32 892
rect -9 858 6 884
rect 13 858 32 884
rect 96 880 158 892
rect 170 880 245 892
rect 303 880 378 892
rect 390 880 421 892
rect 427 880 462 892
rect 96 878 258 880
rect -9 850 32 858
rect 114 854 127 878
rect 142 876 157 878
rect -3 840 -2 850
rect 13 840 26 850
rect 41 840 71 854
rect 114 840 157 854
rect 181 851 188 858
rect 191 854 258 878
rect 290 878 462 880
rect 260 856 288 860
rect 290 856 370 878
rect 391 876 406 878
rect 260 854 370 856
rect 191 850 370 854
rect 164 840 194 850
rect 196 840 349 850
rect 357 840 387 850
rect 391 840 421 854
rect 449 840 462 878
rect 534 884 569 892
rect 534 858 535 884
rect 542 858 569 884
rect 477 840 507 854
rect 534 850 569 858
rect 571 884 612 892
rect 571 858 586 884
rect 593 858 612 884
rect 676 880 738 892
rect 750 880 825 892
rect 883 880 958 892
rect 970 880 1001 892
rect 1007 880 1042 892
rect 676 878 838 880
rect 571 850 612 858
rect 694 854 707 878
rect 722 876 737 878
rect 534 840 535 850
rect 550 840 563 850
rect 577 840 578 850
rect 593 840 606 850
rect 621 840 651 854
rect 694 840 737 854
rect 761 851 768 858
rect 771 854 838 878
rect 870 878 1042 880
rect 840 856 868 860
rect 870 856 950 878
rect 971 876 986 878
rect 840 854 950 856
rect 771 850 950 854
rect 744 840 774 850
rect 776 840 929 850
rect 937 840 967 850
rect 971 840 1001 854
rect 1029 840 1042 878
rect 1114 884 1149 892
rect 1114 858 1115 884
rect 1122 858 1149 884
rect 1057 840 1087 854
rect 1114 850 1149 858
rect 1151 884 1192 892
rect 1151 858 1166 884
rect 1173 858 1192 884
rect 1256 880 1318 892
rect 1330 880 1405 892
rect 1463 880 1538 892
rect 1550 880 1581 892
rect 1587 880 1622 892
rect 1256 878 1418 880
rect 1151 850 1192 858
rect 1274 854 1287 878
rect 1302 876 1317 878
rect 1114 840 1115 850
rect 1130 840 1143 850
rect 1157 840 1158 850
rect 1173 840 1186 850
rect 1201 840 1231 854
rect 1274 840 1317 854
rect 1341 851 1348 858
rect 1351 854 1418 878
rect 1450 878 1622 880
rect 1420 856 1448 860
rect 1450 856 1530 878
rect 1551 876 1566 878
rect 1420 854 1530 856
rect 1351 850 1530 854
rect 1324 840 1354 850
rect 1356 840 1509 850
rect 1517 840 1547 850
rect 1551 840 1581 854
rect 1609 840 1622 878
rect 1694 884 1729 892
rect 1694 858 1695 884
rect 1702 858 1729 884
rect 1637 840 1667 854
rect 1694 850 1729 858
rect 1731 884 1772 892
rect 1731 858 1746 884
rect 1753 858 1772 884
rect 1836 880 1898 892
rect 1910 880 1985 892
rect 2043 880 2118 892
rect 2130 880 2161 892
rect 2167 880 2202 892
rect 1836 878 1998 880
rect 1731 850 1772 858
rect 1854 854 1867 878
rect 1882 876 1897 878
rect 1694 840 1695 850
rect 1710 840 1723 850
rect 1737 840 1738 850
rect 1753 840 1766 850
rect 1781 840 1811 854
rect 1854 840 1897 854
rect 1921 851 1928 858
rect 1931 854 1998 878
rect 2030 878 2202 880
rect 2000 856 2028 860
rect 2030 856 2110 878
rect 2131 876 2146 878
rect 2000 854 2110 856
rect 1931 850 2110 854
rect 1904 840 1934 850
rect 1936 840 2089 850
rect 2097 840 2127 850
rect 2131 840 2161 854
rect 2189 840 2202 878
rect 2274 884 2309 892
rect 2274 858 2275 884
rect 2282 858 2309 884
rect 2217 840 2247 854
rect 2274 850 2309 858
rect 2311 884 2352 892
rect 2311 858 2326 884
rect 2333 858 2352 884
rect 2416 880 2478 892
rect 2490 880 2565 892
rect 2623 880 2698 892
rect 2710 880 2741 892
rect 2747 880 2782 892
rect 2416 878 2578 880
rect 2311 850 2352 858
rect 2434 854 2447 878
rect 2462 876 2477 878
rect 2274 840 2275 850
rect 2290 840 2303 850
rect 2317 840 2318 850
rect 2333 840 2346 850
rect 2361 840 2391 854
rect 2434 840 2477 854
rect 2501 851 2508 858
rect 2511 854 2578 878
rect 2610 878 2782 880
rect 2580 856 2608 860
rect 2610 856 2690 878
rect 2711 876 2726 878
rect 2580 854 2690 856
rect 2511 850 2690 854
rect 2484 840 2514 850
rect 2516 840 2669 850
rect 2677 840 2707 850
rect 2711 840 2741 854
rect 2769 840 2782 878
rect 2854 884 2889 892
rect 2854 858 2855 884
rect 2862 858 2889 884
rect 2797 840 2827 854
rect 2854 850 2889 858
rect 2891 884 2932 892
rect 2891 858 2906 884
rect 2913 858 2932 884
rect 2996 880 3058 892
rect 3070 880 3145 892
rect 3203 880 3278 892
rect 3290 880 3321 892
rect 3327 880 3362 892
rect 2996 878 3158 880
rect 2891 850 2932 858
rect 3014 854 3027 878
rect 3042 876 3057 878
rect 2854 840 2855 850
rect 2870 840 2883 850
rect 2897 840 2898 850
rect 2913 840 2926 850
rect 2941 840 2971 854
rect 3014 840 3057 854
rect 3081 851 3088 858
rect 3091 854 3158 878
rect 3190 878 3362 880
rect 3160 856 3188 860
rect 3190 856 3270 878
rect 3291 876 3306 878
rect 3160 854 3270 856
rect 3091 850 3270 854
rect 3064 840 3094 850
rect 3096 840 3249 850
rect 3257 840 3287 850
rect 3291 840 3321 854
rect 3349 840 3362 878
rect 3434 884 3469 892
rect 3434 858 3435 884
rect 3442 858 3469 884
rect 3377 840 3407 854
rect 3434 850 3469 858
rect 3434 840 3435 850
rect 3450 840 3463 850
rect -3 834 3469 840
rect -2 826 3469 834
rect 5889 884 5930 892
rect 5889 858 5904 884
rect 5911 858 5930 884
rect 5994 880 6056 892
rect 6068 880 6143 892
rect 6201 880 6276 892
rect 6288 880 6319 892
rect 6325 880 6360 892
rect 5994 878 6156 880
rect 5889 850 5930 858
rect 6012 854 6025 878
rect 6040 876 6055 878
rect 5895 840 5896 850
rect 5911 840 5924 850
rect 5939 840 5969 854
rect 6012 840 6055 854
rect 6079 851 6086 858
rect 6089 854 6156 878
rect 6188 878 6360 880
rect 6158 856 6186 860
rect 6188 856 6268 878
rect 6289 876 6304 878
rect 6158 854 6268 856
rect 6089 850 6268 854
rect 6062 840 6092 850
rect 6094 840 6247 850
rect 6255 840 6285 850
rect 6289 840 6319 854
rect 6347 840 6360 878
rect 6432 884 6467 892
rect 6432 858 6433 884
rect 6440 858 6467 884
rect 6375 840 6405 854
rect 6432 850 6467 858
rect 6469 884 6510 892
rect 6469 858 6484 884
rect 6491 858 6510 884
rect 6574 880 6636 892
rect 6648 880 6723 892
rect 6781 880 6856 892
rect 6868 880 6899 892
rect 6905 880 6940 892
rect 6574 878 6736 880
rect 6469 850 6510 858
rect 6592 854 6605 878
rect 6620 876 6635 878
rect 6432 840 6433 850
rect 6448 840 6461 850
rect 6475 840 6476 850
rect 6491 840 6504 850
rect 6519 840 6549 854
rect 6592 840 6635 854
rect 6659 851 6666 858
rect 6669 854 6736 878
rect 6768 878 6940 880
rect 6738 856 6766 860
rect 6768 856 6848 878
rect 6869 876 6884 878
rect 6738 854 6848 856
rect 6669 850 6848 854
rect 6642 840 6672 850
rect 6674 840 6827 850
rect 6835 840 6865 850
rect 6869 840 6899 854
rect 6927 840 6940 878
rect 7012 884 7047 892
rect 7012 858 7013 884
rect 7020 858 7047 884
rect 6955 840 6985 854
rect 7012 850 7047 858
rect 7049 884 7090 892
rect 7049 858 7064 884
rect 7071 858 7090 884
rect 7154 880 7216 892
rect 7228 880 7303 892
rect 7361 880 7436 892
rect 7448 880 7479 892
rect 7485 880 7520 892
rect 7154 878 7316 880
rect 7049 850 7090 858
rect 7172 854 7185 878
rect 7200 876 7215 878
rect 7012 840 7013 850
rect 7028 840 7041 850
rect 7055 840 7056 850
rect 7071 840 7084 850
rect 7099 840 7129 854
rect 7172 840 7215 854
rect 7239 851 7246 858
rect 7249 854 7316 878
rect 7348 878 7520 880
rect 7318 856 7346 860
rect 7348 856 7428 878
rect 7449 876 7464 878
rect 7318 854 7428 856
rect 7249 850 7428 854
rect 7222 840 7252 850
rect 7254 840 7407 850
rect 7415 840 7445 850
rect 7449 840 7479 854
rect 7507 840 7520 878
rect 7592 884 7627 892
rect 7592 858 7593 884
rect 7600 858 7627 884
rect 7535 840 7565 854
rect 7592 850 7627 858
rect 7629 884 7670 892
rect 7629 858 7644 884
rect 7651 858 7670 884
rect 7734 880 7796 892
rect 7808 880 7883 892
rect 7941 880 8016 892
rect 8028 880 8059 892
rect 8065 880 8100 892
rect 7734 878 7896 880
rect 7629 850 7670 858
rect 7752 854 7765 878
rect 7780 876 7795 878
rect 7592 840 7593 850
rect 7608 840 7621 850
rect 7635 840 7636 850
rect 7651 840 7664 850
rect 7679 840 7709 854
rect 7752 840 7795 854
rect 7819 851 7826 858
rect 7829 854 7896 878
rect 7928 878 8100 880
rect 7898 856 7926 860
rect 7928 856 8008 878
rect 8029 876 8044 878
rect 7898 854 8008 856
rect 7829 850 8008 854
rect 7802 840 7832 850
rect 7834 840 7987 850
rect 7995 840 8025 850
rect 8029 840 8059 854
rect 8087 840 8100 878
rect 8172 884 8207 892
rect 8172 858 8173 884
rect 8180 858 8207 884
rect 8115 840 8145 854
rect 8172 850 8207 858
rect 8209 884 8250 892
rect 8209 858 8224 884
rect 8231 858 8250 884
rect 8314 880 8376 892
rect 8388 880 8463 892
rect 8521 880 8596 892
rect 8608 880 8639 892
rect 8645 880 8680 892
rect 8314 878 8476 880
rect 8209 850 8250 858
rect 8332 854 8345 878
rect 8360 876 8375 878
rect 8172 840 8173 850
rect 8188 840 8201 850
rect 8215 840 8216 850
rect 8231 840 8244 850
rect 8259 840 8289 854
rect 8332 840 8375 854
rect 8399 851 8406 858
rect 8409 854 8476 878
rect 8508 878 8680 880
rect 8478 856 8506 860
rect 8508 856 8588 878
rect 8609 876 8624 878
rect 8478 854 8588 856
rect 8409 850 8588 854
rect 8382 840 8412 850
rect 8414 840 8567 850
rect 8575 840 8605 850
rect 8609 840 8639 854
rect 8667 840 8680 878
rect 8752 884 8787 892
rect 8752 858 8753 884
rect 8760 858 8787 884
rect 8695 840 8725 854
rect 8752 850 8787 858
rect 8789 884 8830 892
rect 8789 858 8804 884
rect 8811 858 8830 884
rect 8894 880 8956 892
rect 8968 880 9043 892
rect 9101 880 9176 892
rect 9188 880 9219 892
rect 9225 880 9260 892
rect 8894 878 9056 880
rect 8789 850 8830 858
rect 8912 854 8925 878
rect 8940 876 8955 878
rect 8752 840 8753 850
rect 8768 840 8781 850
rect 8795 840 8796 850
rect 8811 840 8824 850
rect 8839 840 8869 854
rect 8912 840 8955 854
rect 8979 851 8986 858
rect 8989 854 9056 878
rect 9088 878 9260 880
rect 9058 856 9086 860
rect 9088 856 9168 878
rect 9189 876 9204 878
rect 9058 854 9168 856
rect 8989 850 9168 854
rect 8962 840 8992 850
rect 8994 840 9147 850
rect 9155 840 9185 850
rect 9189 840 9219 854
rect 9247 840 9260 878
rect 9332 884 9367 892
rect 9332 858 9333 884
rect 9340 858 9367 884
rect 9275 840 9305 854
rect 9332 850 9367 858
rect 9332 840 9333 850
rect 9348 840 9361 850
rect 5889 826 9361 840
rect 13 796 26 826
rect 41 808 71 826
rect 114 812 128 826
rect 164 812 384 826
rect 115 810 128 812
rect 81 798 96 810
rect 78 796 100 798
rect 105 796 135 810
rect 196 808 349 812
rect 178 796 370 808
rect 413 796 443 810
rect 449 796 462 826
rect 477 808 507 826
rect 550 796 563 826
rect 593 796 606 826
rect 621 808 651 826
rect 694 812 708 826
rect 744 812 964 826
rect 695 810 708 812
rect 661 798 676 810
rect 658 796 680 798
rect 685 796 715 810
rect 776 808 929 812
rect 758 796 950 808
rect 993 796 1023 810
rect 1029 796 1042 826
rect 1057 808 1087 826
rect 1130 796 1143 826
rect 1173 796 1186 826
rect 1201 808 1231 826
rect 1274 812 1288 826
rect 1324 812 1544 826
rect 1275 810 1288 812
rect 1241 798 1256 810
rect 1238 796 1260 798
rect 1265 796 1295 810
rect 1356 808 1509 812
rect 1338 796 1530 808
rect 1573 796 1603 810
rect 1609 796 1622 826
rect 1637 808 1667 826
rect 1710 796 1723 826
rect 1753 796 1766 826
rect 1781 808 1811 826
rect 1854 812 1868 826
rect 1904 812 2124 826
rect 1855 810 1868 812
rect 1821 798 1836 810
rect 1818 796 1840 798
rect 1845 796 1875 810
rect 1936 808 2089 812
rect 1918 796 2110 808
rect 2153 796 2183 810
rect 2189 796 2202 826
rect 2217 808 2247 826
rect 2290 796 2303 826
rect 2333 796 2346 826
rect 2361 808 2391 826
rect 2434 812 2448 826
rect 2484 812 2704 826
rect 2435 810 2448 812
rect 2401 798 2416 810
rect 2398 796 2420 798
rect 2425 796 2455 810
rect 2516 808 2669 812
rect 2498 796 2690 808
rect 2733 796 2763 810
rect 2769 796 2782 826
rect 2797 808 2827 826
rect 2870 796 2883 826
rect 2913 796 2926 826
rect 2941 808 2971 826
rect 3014 812 3028 826
rect 3064 812 3284 826
rect 3015 810 3028 812
rect 2981 798 2996 810
rect 2978 796 3000 798
rect 3005 796 3035 810
rect 3096 808 3249 812
rect 3078 796 3270 808
rect 3313 796 3343 810
rect 3349 796 3362 826
rect 3377 808 3407 826
rect 3450 796 3463 826
rect 5911 796 5924 826
rect 5939 808 5969 826
rect 6012 812 6026 826
rect 6062 812 6282 826
rect 6013 810 6026 812
rect 5979 798 5994 810
rect 5976 796 5998 798
rect 6003 796 6033 810
rect 6094 808 6247 812
rect 6076 796 6268 808
rect 6311 796 6341 810
rect 6347 796 6360 826
rect 6375 808 6405 826
rect 6448 796 6461 826
rect 6491 796 6504 826
rect 6519 808 6549 826
rect 6592 812 6606 826
rect 6642 812 6862 826
rect 6593 810 6606 812
rect 6559 798 6574 810
rect 6556 796 6578 798
rect 6583 796 6613 810
rect 6674 808 6827 812
rect 6656 796 6848 808
rect 6891 796 6921 810
rect 6927 796 6940 826
rect 6955 808 6985 826
rect 7028 796 7041 826
rect 7071 796 7084 826
rect 7099 808 7129 826
rect 7172 812 7186 826
rect 7222 812 7442 826
rect 7173 810 7186 812
rect 7139 798 7154 810
rect 7136 796 7158 798
rect 7163 796 7193 810
rect 7254 808 7407 812
rect 7236 796 7428 808
rect 7471 796 7501 810
rect 7507 796 7520 826
rect 7535 808 7565 826
rect 7608 796 7621 826
rect 7651 796 7664 826
rect 7679 808 7709 826
rect 7752 812 7766 826
rect 7802 812 8022 826
rect 7753 810 7766 812
rect 7719 798 7734 810
rect 7716 796 7738 798
rect 7743 796 7773 810
rect 7834 808 7987 812
rect 7816 796 8008 808
rect 8051 796 8081 810
rect 8087 796 8100 826
rect 8115 808 8145 826
rect 8188 796 8201 826
rect 8231 796 8244 826
rect 8259 808 8289 826
rect 8332 812 8346 826
rect 8382 812 8602 826
rect 8333 810 8346 812
rect 8299 798 8314 810
rect 8296 796 8318 798
rect 8323 796 8353 810
rect 8414 808 8567 812
rect 8396 796 8588 808
rect 8631 796 8661 810
rect 8667 796 8680 826
rect 8695 808 8725 826
rect 8768 796 8781 826
rect 8811 796 8824 826
rect 8839 808 8869 826
rect 8912 812 8926 826
rect 8962 812 9182 826
rect 8913 810 8926 812
rect 8879 798 8894 810
rect 8876 796 8898 798
rect 8903 796 8933 810
rect 8994 808 9147 812
rect 8976 796 9168 808
rect 9211 796 9241 810
rect 9247 796 9260 826
rect 9275 808 9305 826
rect 9348 796 9361 826
rect -2 782 3469 796
rect 5889 782 9361 796
rect 13 678 26 782
rect 71 760 72 770
rect 87 760 100 770
rect 71 756 100 760
rect 105 756 135 782
rect 153 768 169 770
rect 241 768 294 782
rect 242 766 306 768
rect 349 766 364 782
rect 413 779 443 782
rect 413 776 449 779
rect 379 768 395 770
rect 153 756 168 760
rect 71 754 168 756
rect 196 754 364 766
rect 380 756 395 760
rect 413 757 452 776
rect 471 770 478 771
rect 477 763 478 770
rect 461 760 462 763
rect 477 760 490 763
rect 413 756 443 757
rect 452 756 458 757
rect 461 756 490 760
rect 380 755 490 756
rect 380 754 496 755
rect 55 746 106 754
rect 55 734 80 746
rect 87 734 106 746
rect 137 746 187 754
rect 137 738 153 746
rect 160 744 187 746
rect 196 744 417 754
rect 160 734 417 744
rect 446 746 496 754
rect 446 737 462 746
rect 55 726 106 734
rect 153 726 417 734
rect 443 734 462 737
rect 469 734 496 746
rect 443 726 496 734
rect 71 718 72 726
rect 87 718 100 726
rect 71 710 87 718
rect 68 703 87 706
rect 68 694 90 703
rect 41 684 90 694
rect 41 678 71 684
rect 90 679 95 684
rect 13 662 87 678
rect 105 670 135 726
rect 170 716 378 726
rect 413 722 458 726
rect 461 725 462 726
rect 477 725 490 726
rect 196 686 385 716
rect 211 683 385 686
rect 204 680 385 683
rect 13 660 26 662
rect 41 660 75 662
rect 13 644 87 660
rect 114 656 127 670
rect 142 656 158 672
rect 204 667 215 680
rect -3 622 -2 638
rect 13 622 26 644
rect 41 622 71 644
rect 114 640 176 656
rect 204 649 215 665
rect 220 660 230 680
rect 240 660 254 680
rect 257 667 266 680
rect 282 667 291 680
rect 220 649 254 660
rect 257 649 266 665
rect 282 649 291 665
rect 298 660 308 680
rect 318 660 332 680
rect 333 667 344 680
rect 298 649 332 660
rect 333 649 344 665
rect 390 656 406 672
rect 413 670 443 722
rect 477 718 478 725
rect 462 710 478 718
rect 449 678 462 697
rect 477 678 507 694
rect 449 662 523 678
rect 449 660 462 662
rect 477 660 511 662
rect 114 638 127 640
rect 142 638 176 640
rect 114 622 176 638
rect 220 633 236 636
rect 298 633 328 644
rect 376 640 422 656
rect 449 644 523 660
rect 376 638 410 640
rect 375 622 422 638
rect 449 622 462 644
rect 477 622 507 644
rect 534 622 535 638
rect 550 622 563 782
rect 593 678 606 782
rect 651 760 652 770
rect 667 760 680 770
rect 651 756 680 760
rect 685 756 715 782
rect 733 768 749 770
rect 821 768 874 782
rect 822 766 886 768
rect 929 766 944 782
rect 993 779 1023 782
rect 993 776 1029 779
rect 959 768 975 770
rect 733 756 748 760
rect 651 754 748 756
rect 776 754 944 766
rect 960 756 975 760
rect 993 757 1032 776
rect 1051 770 1058 771
rect 1057 763 1058 770
rect 1041 760 1042 763
rect 1057 760 1070 763
rect 993 756 1023 757
rect 1032 756 1038 757
rect 1041 756 1070 760
rect 960 755 1070 756
rect 960 754 1076 755
rect 635 746 686 754
rect 635 734 660 746
rect 667 734 686 746
rect 717 746 767 754
rect 717 738 733 746
rect 740 744 767 746
rect 776 744 997 754
rect 740 734 997 744
rect 1026 746 1076 754
rect 1026 737 1042 746
rect 635 726 686 734
rect 733 726 997 734
rect 1023 734 1042 737
rect 1049 734 1076 746
rect 1023 726 1076 734
rect 651 718 652 726
rect 667 718 680 726
rect 651 710 667 718
rect 648 703 667 706
rect 648 694 670 703
rect 621 684 670 694
rect 621 678 651 684
rect 670 679 675 684
rect 593 662 667 678
rect 685 670 715 726
rect 750 716 958 726
rect 993 722 1038 726
rect 1041 725 1042 726
rect 1057 725 1070 726
rect 776 686 965 716
rect 791 683 965 686
rect 784 680 965 683
rect 593 660 606 662
rect 621 660 655 662
rect 593 644 667 660
rect 694 656 707 670
rect 722 656 738 672
rect 784 667 795 680
rect 577 622 578 638
rect 593 622 606 644
rect 621 622 651 644
rect 694 640 756 656
rect 784 649 795 665
rect 800 660 810 680
rect 820 660 834 680
rect 837 667 846 680
rect 862 667 871 680
rect 800 649 834 660
rect 837 649 846 665
rect 862 649 871 665
rect 878 660 888 680
rect 898 660 912 680
rect 913 667 924 680
rect 878 649 912 660
rect 913 649 924 665
rect 970 656 986 672
rect 993 670 1023 722
rect 1057 718 1058 725
rect 1042 710 1058 718
rect 1029 678 1042 697
rect 1057 678 1087 694
rect 1029 662 1103 678
rect 1029 660 1042 662
rect 1057 660 1091 662
rect 694 638 707 640
rect 722 638 756 640
rect 694 622 756 638
rect 800 633 816 636
rect 878 633 908 644
rect 956 640 1002 656
rect 1029 644 1103 660
rect 956 638 990 640
rect 955 622 1002 638
rect 1029 622 1042 644
rect 1057 622 1087 644
rect 1114 622 1115 638
rect 1130 622 1143 782
rect 1173 678 1186 782
rect 1231 760 1232 770
rect 1247 760 1260 770
rect 1231 756 1260 760
rect 1265 756 1295 782
rect 1313 768 1329 770
rect 1401 768 1454 782
rect 1402 766 1466 768
rect 1509 766 1524 782
rect 1573 779 1603 782
rect 1573 776 1609 779
rect 1539 768 1555 770
rect 1313 756 1328 760
rect 1231 754 1328 756
rect 1356 754 1524 766
rect 1540 756 1555 760
rect 1573 757 1612 776
rect 1631 770 1638 771
rect 1637 763 1638 770
rect 1621 760 1622 763
rect 1637 760 1650 763
rect 1573 756 1603 757
rect 1612 756 1618 757
rect 1621 756 1650 760
rect 1540 755 1650 756
rect 1540 754 1656 755
rect 1215 746 1266 754
rect 1215 734 1240 746
rect 1247 734 1266 746
rect 1297 746 1347 754
rect 1297 738 1313 746
rect 1320 744 1347 746
rect 1356 744 1577 754
rect 1320 734 1577 744
rect 1606 746 1656 754
rect 1606 737 1622 746
rect 1215 726 1266 734
rect 1313 726 1577 734
rect 1603 734 1622 737
rect 1629 734 1656 746
rect 1603 726 1656 734
rect 1231 718 1232 726
rect 1247 718 1260 726
rect 1231 710 1247 718
rect 1228 703 1247 706
rect 1228 694 1250 703
rect 1201 684 1250 694
rect 1201 678 1231 684
rect 1250 679 1255 684
rect 1173 662 1247 678
rect 1265 670 1295 726
rect 1330 716 1538 726
rect 1573 722 1618 726
rect 1621 725 1622 726
rect 1637 725 1650 726
rect 1356 686 1545 716
rect 1371 683 1545 686
rect 1364 680 1545 683
rect 1173 660 1186 662
rect 1201 660 1235 662
rect 1173 644 1247 660
rect 1274 656 1287 670
rect 1302 656 1318 672
rect 1364 667 1375 680
rect 1157 622 1158 638
rect 1173 622 1186 644
rect 1201 622 1231 644
rect 1274 640 1336 656
rect 1364 649 1375 665
rect 1380 660 1390 680
rect 1400 660 1414 680
rect 1417 667 1426 680
rect 1442 667 1451 680
rect 1380 649 1414 660
rect 1417 649 1426 665
rect 1442 649 1451 665
rect 1458 660 1468 680
rect 1478 660 1492 680
rect 1493 667 1504 680
rect 1458 649 1492 660
rect 1493 649 1504 665
rect 1550 656 1566 672
rect 1573 670 1603 722
rect 1637 718 1638 725
rect 1622 710 1638 718
rect 1609 678 1622 697
rect 1637 678 1667 694
rect 1609 662 1683 678
rect 1609 660 1622 662
rect 1637 660 1671 662
rect 1274 638 1287 640
rect 1302 638 1336 640
rect 1274 622 1336 638
rect 1380 633 1396 636
rect 1458 633 1488 644
rect 1536 640 1582 656
rect 1609 644 1683 660
rect 1536 638 1570 640
rect 1535 622 1582 638
rect 1609 622 1622 644
rect 1637 622 1667 644
rect 1694 622 1695 638
rect 1710 622 1723 782
rect 1753 678 1766 782
rect 1811 760 1812 770
rect 1827 760 1840 770
rect 1811 756 1840 760
rect 1845 756 1875 782
rect 1893 768 1909 770
rect 1981 768 2034 782
rect 1982 766 2046 768
rect 2089 766 2104 782
rect 2153 779 2183 782
rect 2153 776 2189 779
rect 2119 768 2135 770
rect 1893 756 1908 760
rect 1811 754 1908 756
rect 1936 754 2104 766
rect 2120 756 2135 760
rect 2153 757 2192 776
rect 2211 770 2218 771
rect 2217 763 2218 770
rect 2201 760 2202 763
rect 2217 760 2230 763
rect 2153 756 2183 757
rect 2192 756 2198 757
rect 2201 756 2230 760
rect 2120 755 2230 756
rect 2120 754 2236 755
rect 1795 746 1846 754
rect 1795 734 1820 746
rect 1827 734 1846 746
rect 1877 746 1927 754
rect 1877 738 1893 746
rect 1900 744 1927 746
rect 1936 744 2157 754
rect 1900 734 2157 744
rect 2186 746 2236 754
rect 2186 737 2202 746
rect 1795 726 1846 734
rect 1893 726 2157 734
rect 2183 734 2202 737
rect 2209 734 2236 746
rect 2183 726 2236 734
rect 1811 718 1812 726
rect 1827 718 1840 726
rect 1811 710 1827 718
rect 1808 703 1827 706
rect 1808 694 1830 703
rect 1781 684 1830 694
rect 1781 678 1811 684
rect 1830 679 1835 684
rect 1753 662 1827 678
rect 1845 670 1875 726
rect 1910 716 2118 726
rect 2153 722 2198 726
rect 2201 725 2202 726
rect 2217 725 2230 726
rect 1936 686 2125 716
rect 1951 683 2125 686
rect 1944 680 2125 683
rect 1753 660 1766 662
rect 1781 660 1815 662
rect 1753 644 1827 660
rect 1854 656 1867 670
rect 1882 656 1898 672
rect 1944 667 1955 680
rect 1737 622 1738 638
rect 1753 622 1766 644
rect 1781 622 1811 644
rect 1854 640 1916 656
rect 1944 649 1955 665
rect 1960 660 1970 680
rect 1980 660 1994 680
rect 1997 667 2006 680
rect 2022 667 2031 680
rect 1960 649 1994 660
rect 1997 649 2006 665
rect 2022 649 2031 665
rect 2038 660 2048 680
rect 2058 660 2072 680
rect 2073 667 2084 680
rect 2038 649 2072 660
rect 2073 649 2084 665
rect 2130 656 2146 672
rect 2153 670 2183 722
rect 2217 718 2218 725
rect 2202 710 2218 718
rect 2189 678 2202 697
rect 2217 678 2247 694
rect 2189 662 2263 678
rect 2189 660 2202 662
rect 2217 660 2251 662
rect 1854 638 1867 640
rect 1882 638 1916 640
rect 1854 622 1916 638
rect 1960 633 1976 636
rect 2038 633 2068 644
rect 2116 640 2162 656
rect 2189 644 2263 660
rect 2116 638 2150 640
rect 2115 622 2162 638
rect 2189 622 2202 644
rect 2217 622 2247 644
rect 2274 622 2275 638
rect 2290 622 2303 782
rect 2333 678 2346 782
rect 2391 760 2392 770
rect 2407 760 2420 770
rect 2391 756 2420 760
rect 2425 756 2455 782
rect 2473 768 2489 770
rect 2561 768 2614 782
rect 2562 766 2626 768
rect 2669 766 2684 782
rect 2733 779 2763 782
rect 2733 776 2769 779
rect 2699 768 2715 770
rect 2473 756 2488 760
rect 2391 754 2488 756
rect 2516 754 2684 766
rect 2700 756 2715 760
rect 2733 757 2772 776
rect 2791 770 2798 771
rect 2797 763 2798 770
rect 2781 760 2782 763
rect 2797 760 2810 763
rect 2733 756 2763 757
rect 2772 756 2778 757
rect 2781 756 2810 760
rect 2700 755 2810 756
rect 2700 754 2816 755
rect 2375 746 2426 754
rect 2375 734 2400 746
rect 2407 734 2426 746
rect 2457 746 2507 754
rect 2457 738 2473 746
rect 2480 744 2507 746
rect 2516 744 2737 754
rect 2480 734 2737 744
rect 2766 746 2816 754
rect 2766 737 2782 746
rect 2375 726 2426 734
rect 2473 726 2737 734
rect 2763 734 2782 737
rect 2789 734 2816 746
rect 2763 726 2816 734
rect 2391 718 2392 726
rect 2407 718 2420 726
rect 2391 710 2407 718
rect 2388 703 2407 706
rect 2388 694 2410 703
rect 2361 684 2410 694
rect 2361 678 2391 684
rect 2410 679 2415 684
rect 2333 662 2407 678
rect 2425 670 2455 726
rect 2490 716 2698 726
rect 2733 722 2778 726
rect 2781 725 2782 726
rect 2797 725 2810 726
rect 2516 686 2705 716
rect 2531 683 2705 686
rect 2524 680 2705 683
rect 2333 660 2346 662
rect 2361 660 2395 662
rect 2333 644 2407 660
rect 2434 656 2447 670
rect 2462 656 2478 672
rect 2524 667 2535 680
rect 2317 622 2318 638
rect 2333 622 2346 644
rect 2361 622 2391 644
rect 2434 640 2496 656
rect 2524 649 2535 665
rect 2540 660 2550 680
rect 2560 660 2574 680
rect 2577 667 2586 680
rect 2602 667 2611 680
rect 2540 649 2574 660
rect 2577 649 2586 665
rect 2602 649 2611 665
rect 2618 660 2628 680
rect 2638 660 2652 680
rect 2653 667 2664 680
rect 2618 649 2652 660
rect 2653 649 2664 665
rect 2710 656 2726 672
rect 2733 670 2763 722
rect 2797 718 2798 725
rect 2782 710 2798 718
rect 2769 678 2782 697
rect 2797 678 2827 694
rect 2769 662 2843 678
rect 2769 660 2782 662
rect 2797 660 2831 662
rect 2434 638 2447 640
rect 2462 638 2496 640
rect 2434 622 2496 638
rect 2540 633 2556 636
rect 2618 633 2648 644
rect 2696 640 2742 656
rect 2769 644 2843 660
rect 2696 638 2730 640
rect 2695 622 2742 638
rect 2769 622 2782 644
rect 2797 622 2827 644
rect 2854 622 2855 638
rect 2870 622 2883 782
rect 2913 678 2926 782
rect 2971 760 2972 770
rect 2987 760 3000 770
rect 2971 756 3000 760
rect 3005 756 3035 782
rect 3053 768 3069 770
rect 3141 768 3194 782
rect 3142 766 3206 768
rect 3249 766 3264 782
rect 3313 779 3343 782
rect 3313 776 3349 779
rect 3279 768 3295 770
rect 3053 756 3068 760
rect 2971 754 3068 756
rect 3096 754 3264 766
rect 3280 756 3295 760
rect 3313 757 3352 776
rect 3371 770 3378 771
rect 3377 763 3378 770
rect 3361 760 3362 763
rect 3377 760 3390 763
rect 3313 756 3343 757
rect 3352 756 3358 757
rect 3361 756 3390 760
rect 3280 755 3390 756
rect 3280 754 3396 755
rect 2955 746 3006 754
rect 2955 734 2980 746
rect 2987 734 3006 746
rect 3037 746 3087 754
rect 3037 738 3053 746
rect 3060 744 3087 746
rect 3096 744 3317 754
rect 3060 734 3317 744
rect 3346 746 3396 754
rect 3346 737 3362 746
rect 2955 726 3006 734
rect 3053 726 3317 734
rect 3343 734 3362 737
rect 3369 734 3396 746
rect 3343 726 3396 734
rect 2971 718 2972 726
rect 2987 718 3000 726
rect 2971 710 2987 718
rect 2968 703 2987 706
rect 2968 694 2990 703
rect 2941 684 2990 694
rect 2941 678 2971 684
rect 2990 679 2995 684
rect 2913 662 2987 678
rect 3005 670 3035 726
rect 3070 716 3278 726
rect 3313 722 3358 726
rect 3361 725 3362 726
rect 3377 725 3390 726
rect 3096 686 3285 716
rect 3111 683 3285 686
rect 3104 680 3285 683
rect 2913 660 2926 662
rect 2941 660 2975 662
rect 2913 644 2987 660
rect 3014 656 3027 670
rect 3042 656 3058 672
rect 3104 667 3115 680
rect 2897 622 2898 638
rect 2913 622 2926 644
rect 2941 622 2971 644
rect 3014 640 3076 656
rect 3104 649 3115 665
rect 3120 660 3130 680
rect 3140 660 3154 680
rect 3157 667 3166 680
rect 3182 667 3191 680
rect 3120 649 3154 660
rect 3157 649 3166 665
rect 3182 649 3191 665
rect 3198 660 3208 680
rect 3218 660 3232 680
rect 3233 667 3244 680
rect 3198 649 3232 660
rect 3233 649 3244 665
rect 3290 656 3306 672
rect 3313 670 3343 722
rect 3377 718 3378 725
rect 3362 710 3378 718
rect 3349 678 3362 697
rect 3377 678 3407 694
rect 3349 662 3423 678
rect 3349 660 3362 662
rect 3377 660 3411 662
rect 3014 638 3027 640
rect 3042 638 3076 640
rect 3014 622 3076 638
rect 3120 633 3136 636
rect 3198 633 3228 644
rect 3276 640 3322 656
rect 3349 644 3423 660
rect 3276 638 3310 640
rect 3275 622 3322 638
rect 3349 622 3362 644
rect 3377 622 3407 644
rect 3434 622 3435 638
rect 3450 622 3463 782
rect 5911 678 5924 782
rect 5969 760 5970 770
rect 5985 760 5998 770
rect 5969 756 5998 760
rect 6003 756 6033 782
rect 6051 768 6067 770
rect 6139 768 6192 782
rect 6140 766 6204 768
rect 6247 766 6262 782
rect 6311 779 6341 782
rect 6311 776 6347 779
rect 6277 768 6293 770
rect 6051 756 6066 760
rect 5969 754 6066 756
rect 6094 754 6262 766
rect 6278 756 6293 760
rect 6311 757 6350 776
rect 6369 770 6376 771
rect 6375 763 6376 770
rect 6359 760 6360 763
rect 6375 760 6388 763
rect 6311 756 6341 757
rect 6350 756 6356 757
rect 6359 756 6388 760
rect 6278 755 6388 756
rect 6278 754 6394 755
rect 5953 746 6004 754
rect 5953 734 5978 746
rect 5985 734 6004 746
rect 6035 746 6085 754
rect 6035 738 6051 746
rect 6058 744 6085 746
rect 6094 744 6315 754
rect 6058 734 6315 744
rect 6344 746 6394 754
rect 6344 737 6360 746
rect 5953 726 6004 734
rect 6051 726 6315 734
rect 6341 734 6360 737
rect 6367 734 6394 746
rect 6341 726 6394 734
rect 5969 718 5970 726
rect 5985 718 5998 726
rect 5969 710 5985 718
rect 5966 703 5985 706
rect 5966 694 5988 703
rect 5939 684 5988 694
rect 5939 678 5969 684
rect 5988 679 5993 684
rect 5911 662 5985 678
rect 6003 670 6033 726
rect 6068 716 6276 726
rect 6311 722 6356 726
rect 6359 725 6360 726
rect 6375 725 6388 726
rect 6094 686 6283 716
rect 6109 683 6283 686
rect 6102 680 6283 683
rect 5911 660 5924 662
rect 5939 660 5973 662
rect 5911 644 5985 660
rect 6012 656 6025 670
rect 6040 656 6056 672
rect 6102 667 6113 680
rect 5895 622 5896 638
rect 5911 622 5924 644
rect 5939 622 5969 644
rect 6012 640 6074 656
rect 6102 649 6113 665
rect 6118 660 6128 680
rect 6138 660 6152 680
rect 6155 667 6164 680
rect 6180 667 6189 680
rect 6118 649 6152 660
rect 6155 649 6164 665
rect 6180 649 6189 665
rect 6196 660 6206 680
rect 6216 660 6230 680
rect 6231 667 6242 680
rect 6196 649 6230 660
rect 6231 649 6242 665
rect 6288 656 6304 672
rect 6311 670 6341 722
rect 6375 718 6376 725
rect 6360 710 6376 718
rect 6347 678 6360 697
rect 6375 678 6405 694
rect 6347 662 6421 678
rect 6347 660 6360 662
rect 6375 660 6409 662
rect 6012 638 6025 640
rect 6040 638 6074 640
rect 6012 622 6074 638
rect 6118 633 6134 636
rect 6196 633 6226 644
rect 6274 640 6320 656
rect 6347 644 6421 660
rect 6274 638 6308 640
rect 6273 622 6320 638
rect 6347 622 6360 644
rect 6375 622 6405 644
rect 6432 622 6433 638
rect 6448 622 6461 782
rect 6491 678 6504 782
rect 6549 760 6550 770
rect 6565 760 6578 770
rect 6549 756 6578 760
rect 6583 756 6613 782
rect 6631 768 6647 770
rect 6719 768 6772 782
rect 6720 766 6784 768
rect 6827 766 6842 782
rect 6891 779 6921 782
rect 6891 776 6927 779
rect 6857 768 6873 770
rect 6631 756 6646 760
rect 6549 754 6646 756
rect 6674 754 6842 766
rect 6858 756 6873 760
rect 6891 757 6930 776
rect 6949 770 6956 771
rect 6955 763 6956 770
rect 6939 760 6940 763
rect 6955 760 6968 763
rect 6891 756 6921 757
rect 6930 756 6936 757
rect 6939 756 6968 760
rect 6858 755 6968 756
rect 6858 754 6974 755
rect 6533 746 6584 754
rect 6533 734 6558 746
rect 6565 734 6584 746
rect 6615 746 6665 754
rect 6615 738 6631 746
rect 6638 744 6665 746
rect 6674 744 6895 754
rect 6638 734 6895 744
rect 6924 746 6974 754
rect 6924 737 6940 746
rect 6533 726 6584 734
rect 6631 726 6895 734
rect 6921 734 6940 737
rect 6947 734 6974 746
rect 6921 726 6974 734
rect 6549 718 6550 726
rect 6565 718 6578 726
rect 6549 710 6565 718
rect 6546 703 6565 706
rect 6546 694 6568 703
rect 6519 684 6568 694
rect 6519 678 6549 684
rect 6568 679 6573 684
rect 6491 662 6565 678
rect 6583 670 6613 726
rect 6648 716 6856 726
rect 6891 722 6936 726
rect 6939 725 6940 726
rect 6955 725 6968 726
rect 6674 686 6863 716
rect 6689 683 6863 686
rect 6682 680 6863 683
rect 6491 660 6504 662
rect 6519 660 6553 662
rect 6491 644 6565 660
rect 6592 656 6605 670
rect 6620 656 6636 672
rect 6682 667 6693 680
rect 6475 622 6476 638
rect 6491 622 6504 644
rect 6519 622 6549 644
rect 6592 640 6654 656
rect 6682 649 6693 665
rect 6698 660 6708 680
rect 6718 660 6732 680
rect 6735 667 6744 680
rect 6760 667 6769 680
rect 6698 649 6732 660
rect 6735 649 6744 665
rect 6760 649 6769 665
rect 6776 660 6786 680
rect 6796 660 6810 680
rect 6811 667 6822 680
rect 6776 649 6810 660
rect 6811 649 6822 665
rect 6868 656 6884 672
rect 6891 670 6921 722
rect 6955 718 6956 725
rect 6940 710 6956 718
rect 6927 678 6940 697
rect 6955 678 6985 694
rect 6927 662 7001 678
rect 6927 660 6940 662
rect 6955 660 6989 662
rect 6592 638 6605 640
rect 6620 638 6654 640
rect 6592 622 6654 638
rect 6698 633 6714 636
rect 6776 633 6806 644
rect 6854 640 6900 656
rect 6927 644 7001 660
rect 6854 638 6888 640
rect 6853 622 6900 638
rect 6927 622 6940 644
rect 6955 622 6985 644
rect 7012 622 7013 638
rect 7028 622 7041 782
rect 7071 678 7084 782
rect 7129 760 7130 770
rect 7145 760 7158 770
rect 7129 756 7158 760
rect 7163 756 7193 782
rect 7211 768 7227 770
rect 7299 768 7352 782
rect 7300 766 7364 768
rect 7407 766 7422 782
rect 7471 779 7501 782
rect 7471 776 7507 779
rect 7437 768 7453 770
rect 7211 756 7226 760
rect 7129 754 7226 756
rect 7254 754 7422 766
rect 7438 756 7453 760
rect 7471 757 7510 776
rect 7529 770 7536 771
rect 7535 763 7536 770
rect 7519 760 7520 763
rect 7535 760 7548 763
rect 7471 756 7501 757
rect 7510 756 7516 757
rect 7519 756 7548 760
rect 7438 755 7548 756
rect 7438 754 7554 755
rect 7113 746 7164 754
rect 7113 734 7138 746
rect 7145 734 7164 746
rect 7195 746 7245 754
rect 7195 738 7211 746
rect 7218 744 7245 746
rect 7254 744 7475 754
rect 7218 734 7475 744
rect 7504 746 7554 754
rect 7504 737 7520 746
rect 7113 726 7164 734
rect 7211 726 7475 734
rect 7501 734 7520 737
rect 7527 734 7554 746
rect 7501 726 7554 734
rect 7129 718 7130 726
rect 7145 718 7158 726
rect 7129 710 7145 718
rect 7126 703 7145 706
rect 7126 694 7148 703
rect 7099 684 7148 694
rect 7099 678 7129 684
rect 7148 679 7153 684
rect 7071 662 7145 678
rect 7163 670 7193 726
rect 7228 716 7436 726
rect 7471 722 7516 726
rect 7519 725 7520 726
rect 7535 725 7548 726
rect 7254 686 7443 716
rect 7269 683 7443 686
rect 7262 680 7443 683
rect 7071 660 7084 662
rect 7099 660 7133 662
rect 7071 644 7145 660
rect 7172 656 7185 670
rect 7200 656 7216 672
rect 7262 667 7273 680
rect 7055 622 7056 638
rect 7071 622 7084 644
rect 7099 622 7129 644
rect 7172 640 7234 656
rect 7262 649 7273 665
rect 7278 660 7288 680
rect 7298 660 7312 680
rect 7315 667 7324 680
rect 7340 667 7349 680
rect 7278 649 7312 660
rect 7315 649 7324 665
rect 7340 649 7349 665
rect 7356 660 7366 680
rect 7376 660 7390 680
rect 7391 667 7402 680
rect 7356 649 7390 660
rect 7391 649 7402 665
rect 7448 656 7464 672
rect 7471 670 7501 722
rect 7535 718 7536 725
rect 7520 710 7536 718
rect 7507 678 7520 697
rect 7535 678 7565 694
rect 7507 662 7581 678
rect 7507 660 7520 662
rect 7535 660 7569 662
rect 7172 638 7185 640
rect 7200 638 7234 640
rect 7172 622 7234 638
rect 7278 633 7294 636
rect 7356 633 7386 644
rect 7434 640 7480 656
rect 7507 644 7581 660
rect 7434 638 7468 640
rect 7433 622 7480 638
rect 7507 622 7520 644
rect 7535 622 7565 644
rect 7592 622 7593 638
rect 7608 622 7621 782
rect 7651 678 7664 782
rect 7709 760 7710 770
rect 7725 760 7738 770
rect 7709 756 7738 760
rect 7743 756 7773 782
rect 7791 768 7807 770
rect 7879 768 7932 782
rect 7880 766 7944 768
rect 7987 766 8002 782
rect 8051 779 8081 782
rect 8051 776 8087 779
rect 8017 768 8033 770
rect 7791 756 7806 760
rect 7709 754 7806 756
rect 7834 754 8002 766
rect 8018 756 8033 760
rect 8051 757 8090 776
rect 8109 770 8116 771
rect 8115 763 8116 770
rect 8099 760 8100 763
rect 8115 760 8128 763
rect 8051 756 8081 757
rect 8090 756 8096 757
rect 8099 756 8128 760
rect 8018 755 8128 756
rect 8018 754 8134 755
rect 7693 746 7744 754
rect 7693 734 7718 746
rect 7725 734 7744 746
rect 7775 746 7825 754
rect 7775 738 7791 746
rect 7798 744 7825 746
rect 7834 744 8055 754
rect 7798 734 8055 744
rect 8084 746 8134 754
rect 8084 737 8100 746
rect 7693 726 7744 734
rect 7791 726 8055 734
rect 8081 734 8100 737
rect 8107 734 8134 746
rect 8081 726 8134 734
rect 7709 718 7710 726
rect 7725 718 7738 726
rect 7709 710 7725 718
rect 7706 703 7725 706
rect 7706 694 7728 703
rect 7679 684 7728 694
rect 7679 678 7709 684
rect 7728 679 7733 684
rect 7651 662 7725 678
rect 7743 670 7773 726
rect 7808 716 8016 726
rect 8051 722 8096 726
rect 8099 725 8100 726
rect 8115 725 8128 726
rect 7834 686 8023 716
rect 7849 683 8023 686
rect 7842 680 8023 683
rect 7651 660 7664 662
rect 7679 660 7713 662
rect 7651 644 7725 660
rect 7752 656 7765 670
rect 7780 656 7796 672
rect 7842 667 7853 680
rect 7635 622 7636 638
rect 7651 622 7664 644
rect 7679 622 7709 644
rect 7752 640 7814 656
rect 7842 649 7853 665
rect 7858 660 7868 680
rect 7878 660 7892 680
rect 7895 667 7904 680
rect 7920 667 7929 680
rect 7858 649 7892 660
rect 7895 649 7904 665
rect 7920 649 7929 665
rect 7936 660 7946 680
rect 7956 660 7970 680
rect 7971 667 7982 680
rect 7936 649 7970 660
rect 7971 649 7982 665
rect 8028 656 8044 672
rect 8051 670 8081 722
rect 8115 718 8116 725
rect 8100 710 8116 718
rect 8087 678 8100 697
rect 8115 678 8145 694
rect 8087 662 8161 678
rect 8087 660 8100 662
rect 8115 660 8149 662
rect 7752 638 7765 640
rect 7780 638 7814 640
rect 7752 622 7814 638
rect 7858 633 7874 636
rect 7936 633 7966 644
rect 8014 640 8060 656
rect 8087 644 8161 660
rect 8014 638 8048 640
rect 8013 622 8060 638
rect 8087 622 8100 644
rect 8115 622 8145 644
rect 8172 622 8173 638
rect 8188 622 8201 782
rect 8231 678 8244 782
rect 8289 760 8290 770
rect 8305 760 8318 770
rect 8289 756 8318 760
rect 8323 756 8353 782
rect 8371 768 8387 770
rect 8459 768 8512 782
rect 8460 766 8524 768
rect 8567 766 8582 782
rect 8631 779 8661 782
rect 8631 776 8667 779
rect 8597 768 8613 770
rect 8371 756 8386 760
rect 8289 754 8386 756
rect 8414 754 8582 766
rect 8598 756 8613 760
rect 8631 757 8670 776
rect 8689 770 8696 771
rect 8695 763 8696 770
rect 8679 760 8680 763
rect 8695 760 8708 763
rect 8631 756 8661 757
rect 8670 756 8676 757
rect 8679 756 8708 760
rect 8598 755 8708 756
rect 8598 754 8714 755
rect 8273 746 8324 754
rect 8273 734 8298 746
rect 8305 734 8324 746
rect 8355 746 8405 754
rect 8355 738 8371 746
rect 8378 744 8405 746
rect 8414 744 8635 754
rect 8378 734 8635 744
rect 8664 746 8714 754
rect 8664 737 8680 746
rect 8273 726 8324 734
rect 8371 726 8635 734
rect 8661 734 8680 737
rect 8687 734 8714 746
rect 8661 726 8714 734
rect 8289 718 8290 726
rect 8305 718 8318 726
rect 8289 710 8305 718
rect 8286 703 8305 706
rect 8286 694 8308 703
rect 8259 684 8308 694
rect 8259 678 8289 684
rect 8308 679 8313 684
rect 8231 662 8305 678
rect 8323 670 8353 726
rect 8388 716 8596 726
rect 8631 722 8676 726
rect 8679 725 8680 726
rect 8695 725 8708 726
rect 8414 686 8603 716
rect 8429 683 8603 686
rect 8422 680 8603 683
rect 8231 660 8244 662
rect 8259 660 8293 662
rect 8231 644 8305 660
rect 8332 656 8345 670
rect 8360 656 8376 672
rect 8422 667 8433 680
rect 8215 622 8216 638
rect 8231 622 8244 644
rect 8259 622 8289 644
rect 8332 640 8394 656
rect 8422 649 8433 665
rect 8438 660 8448 680
rect 8458 660 8472 680
rect 8475 667 8484 680
rect 8500 667 8509 680
rect 8438 649 8472 660
rect 8475 649 8484 665
rect 8500 649 8509 665
rect 8516 660 8526 680
rect 8536 660 8550 680
rect 8551 667 8562 680
rect 8516 649 8550 660
rect 8551 649 8562 665
rect 8608 656 8624 672
rect 8631 670 8661 722
rect 8695 718 8696 725
rect 8680 710 8696 718
rect 8667 678 8680 697
rect 8695 678 8725 694
rect 8667 662 8741 678
rect 8667 660 8680 662
rect 8695 660 8729 662
rect 8332 638 8345 640
rect 8360 638 8394 640
rect 8332 622 8394 638
rect 8438 633 8454 636
rect 8516 633 8546 644
rect 8594 640 8640 656
rect 8667 644 8741 660
rect 8594 638 8628 640
rect 8593 622 8640 638
rect 8667 622 8680 644
rect 8695 622 8725 644
rect 8752 622 8753 638
rect 8768 622 8781 782
rect 8811 678 8824 782
rect 8869 760 8870 770
rect 8885 760 8898 770
rect 8869 756 8898 760
rect 8903 756 8933 782
rect 8951 768 8967 770
rect 9039 768 9092 782
rect 9040 766 9104 768
rect 9147 766 9162 782
rect 9211 779 9241 782
rect 9211 776 9247 779
rect 9177 768 9193 770
rect 8951 756 8966 760
rect 8869 754 8966 756
rect 8994 754 9162 766
rect 9178 756 9193 760
rect 9211 757 9250 776
rect 9269 770 9276 771
rect 9275 763 9276 770
rect 9259 760 9260 763
rect 9275 760 9288 763
rect 9211 756 9241 757
rect 9250 756 9256 757
rect 9259 756 9288 760
rect 9178 755 9288 756
rect 9178 754 9294 755
rect 8853 746 8904 754
rect 8853 734 8878 746
rect 8885 734 8904 746
rect 8935 746 8985 754
rect 8935 738 8951 746
rect 8958 744 8985 746
rect 8994 744 9215 754
rect 8958 734 9215 744
rect 9244 746 9294 754
rect 9244 737 9260 746
rect 8853 726 8904 734
rect 8951 726 9215 734
rect 9241 734 9260 737
rect 9267 734 9294 746
rect 9241 726 9294 734
rect 8869 718 8870 726
rect 8885 718 8898 726
rect 8869 710 8885 718
rect 8866 703 8885 706
rect 8866 694 8888 703
rect 8839 684 8888 694
rect 8839 678 8869 684
rect 8888 679 8893 684
rect 8811 662 8885 678
rect 8903 670 8933 726
rect 8968 716 9176 726
rect 9211 722 9256 726
rect 9259 725 9260 726
rect 9275 725 9288 726
rect 8994 686 9183 716
rect 9009 683 9183 686
rect 9002 680 9183 683
rect 8811 660 8824 662
rect 8839 660 8873 662
rect 8811 644 8885 660
rect 8912 656 8925 670
rect 8940 656 8956 672
rect 9002 667 9013 680
rect 8795 622 8796 638
rect 8811 622 8824 644
rect 8839 622 8869 644
rect 8912 640 8974 656
rect 9002 649 9013 665
rect 9018 660 9028 680
rect 9038 660 9052 680
rect 9055 667 9064 680
rect 9080 667 9089 680
rect 9018 649 9052 660
rect 9055 649 9064 665
rect 9080 649 9089 665
rect 9096 660 9106 680
rect 9116 660 9130 680
rect 9131 667 9142 680
rect 9096 649 9130 660
rect 9131 649 9142 665
rect 9188 656 9204 672
rect 9211 670 9241 722
rect 9275 718 9276 725
rect 9260 710 9276 718
rect 9247 678 9260 697
rect 9275 678 9305 694
rect 9247 662 9321 678
rect 9247 660 9260 662
rect 9275 660 9309 662
rect 8912 638 8925 640
rect 8940 638 8974 640
rect 8912 622 8974 638
rect 9018 633 9034 636
rect 9096 633 9126 644
rect 9174 640 9220 656
rect 9247 644 9321 660
rect 9174 638 9208 640
rect 9173 622 9220 638
rect 9247 622 9260 644
rect 9275 622 9305 644
rect 9332 622 9333 638
rect 9348 622 9361 782
rect -9 614 32 622
rect -9 588 6 614
rect 13 588 32 614
rect 96 610 158 622
rect 170 610 245 622
rect 303 610 378 622
rect 390 610 421 622
rect 427 610 462 622
rect 96 608 258 610
rect -9 580 32 588
rect 114 584 127 608
rect 142 606 157 608
rect -3 570 -2 580
rect 13 570 26 580
rect 41 570 71 584
rect 114 570 157 584
rect 181 581 188 588
rect 191 584 258 608
rect 290 608 462 610
rect 260 586 288 590
rect 290 586 370 608
rect 391 606 406 608
rect 260 584 370 586
rect 191 580 370 584
rect 164 570 194 580
rect 196 570 349 580
rect 357 570 387 580
rect 391 570 421 584
rect 449 570 462 608
rect 534 614 569 622
rect 534 588 535 614
rect 542 588 569 614
rect 477 570 507 584
rect 534 580 569 588
rect 571 614 612 622
rect 571 588 586 614
rect 593 588 612 614
rect 676 610 738 622
rect 750 610 825 622
rect 883 610 958 622
rect 970 610 1001 622
rect 1007 610 1042 622
rect 676 608 838 610
rect 571 580 612 588
rect 694 584 707 608
rect 722 606 737 608
rect 534 570 535 580
rect 550 570 563 580
rect 577 570 578 580
rect 593 570 606 580
rect 621 570 651 584
rect 694 570 737 584
rect 761 581 768 588
rect 771 584 838 608
rect 870 608 1042 610
rect 840 586 868 590
rect 870 586 950 608
rect 971 606 986 608
rect 840 584 950 586
rect 771 580 950 584
rect 744 570 774 580
rect 776 570 929 580
rect 937 570 967 580
rect 971 570 1001 584
rect 1029 570 1042 608
rect 1114 614 1149 622
rect 1114 588 1115 614
rect 1122 588 1149 614
rect 1057 570 1087 584
rect 1114 580 1149 588
rect 1151 614 1192 622
rect 1151 588 1166 614
rect 1173 588 1192 614
rect 1256 610 1318 622
rect 1330 610 1405 622
rect 1463 610 1538 622
rect 1550 610 1581 622
rect 1587 610 1622 622
rect 1256 608 1418 610
rect 1151 580 1192 588
rect 1274 584 1287 608
rect 1302 606 1317 608
rect 1114 570 1115 580
rect 1130 570 1143 580
rect 1157 570 1158 580
rect 1173 570 1186 580
rect 1201 570 1231 584
rect 1274 570 1317 584
rect 1341 581 1348 588
rect 1351 584 1418 608
rect 1450 608 1622 610
rect 1420 586 1448 590
rect 1450 586 1530 608
rect 1551 606 1566 608
rect 1420 584 1530 586
rect 1351 580 1530 584
rect 1324 570 1354 580
rect 1356 570 1509 580
rect 1517 570 1547 580
rect 1551 570 1581 584
rect 1609 570 1622 608
rect 1694 614 1729 622
rect 1694 588 1695 614
rect 1702 588 1729 614
rect 1637 570 1667 584
rect 1694 580 1729 588
rect 1731 614 1772 622
rect 1731 588 1746 614
rect 1753 588 1772 614
rect 1836 610 1898 622
rect 1910 610 1985 622
rect 2043 610 2118 622
rect 2130 610 2161 622
rect 2167 610 2202 622
rect 1836 608 1998 610
rect 1731 580 1772 588
rect 1854 584 1867 608
rect 1882 606 1897 608
rect 1694 570 1695 580
rect 1710 570 1723 580
rect 1737 570 1738 580
rect 1753 570 1766 580
rect 1781 570 1811 584
rect 1854 570 1897 584
rect 1921 581 1928 588
rect 1931 584 1998 608
rect 2030 608 2202 610
rect 2000 586 2028 590
rect 2030 586 2110 608
rect 2131 606 2146 608
rect 2000 584 2110 586
rect 1931 580 2110 584
rect 1904 570 1934 580
rect 1936 570 2089 580
rect 2097 570 2127 580
rect 2131 570 2161 584
rect 2189 570 2202 608
rect 2274 614 2309 622
rect 2274 588 2275 614
rect 2282 588 2309 614
rect 2217 570 2247 584
rect 2274 580 2309 588
rect 2311 614 2352 622
rect 2311 588 2326 614
rect 2333 588 2352 614
rect 2416 610 2478 622
rect 2490 610 2565 622
rect 2623 610 2698 622
rect 2710 610 2741 622
rect 2747 610 2782 622
rect 2416 608 2578 610
rect 2311 580 2352 588
rect 2434 584 2447 608
rect 2462 606 2477 608
rect 2274 570 2275 580
rect 2290 570 2303 580
rect 2317 570 2318 580
rect 2333 570 2346 580
rect 2361 570 2391 584
rect 2434 570 2477 584
rect 2501 581 2508 588
rect 2511 584 2578 608
rect 2610 608 2782 610
rect 2580 586 2608 590
rect 2610 586 2690 608
rect 2711 606 2726 608
rect 2580 584 2690 586
rect 2511 580 2690 584
rect 2484 570 2514 580
rect 2516 570 2669 580
rect 2677 570 2707 580
rect 2711 570 2741 584
rect 2769 570 2782 608
rect 2854 614 2889 622
rect 2854 588 2855 614
rect 2862 588 2889 614
rect 2797 570 2827 584
rect 2854 580 2889 588
rect 2891 614 2932 622
rect 2891 588 2906 614
rect 2913 588 2932 614
rect 2996 610 3058 622
rect 3070 610 3145 622
rect 3203 610 3278 622
rect 3290 610 3321 622
rect 3327 610 3362 622
rect 2996 608 3158 610
rect 2891 580 2932 588
rect 3014 584 3027 608
rect 3042 606 3057 608
rect 2854 570 2855 580
rect 2870 570 2883 580
rect 2897 570 2898 580
rect 2913 570 2926 580
rect 2941 570 2971 584
rect 3014 570 3057 584
rect 3081 581 3088 588
rect 3091 584 3158 608
rect 3190 608 3362 610
rect 3160 586 3188 590
rect 3190 586 3270 608
rect 3291 606 3306 608
rect 3160 584 3270 586
rect 3091 580 3270 584
rect 3064 570 3094 580
rect 3096 570 3249 580
rect 3257 570 3287 580
rect 3291 570 3321 584
rect 3349 570 3362 608
rect 3434 614 3469 622
rect 3434 588 3435 614
rect 3442 588 3469 614
rect 3377 570 3407 584
rect 3434 580 3469 588
rect 3434 570 3435 580
rect 3450 570 3463 580
rect -3 564 3469 570
rect -2 556 3469 564
rect 5889 614 5930 622
rect 5889 588 5904 614
rect 5911 588 5930 614
rect 5994 610 6056 622
rect 6068 610 6143 622
rect 6201 610 6276 622
rect 6288 610 6319 622
rect 6325 610 6360 622
rect 5994 608 6156 610
rect 5889 580 5930 588
rect 6012 584 6025 608
rect 6040 606 6055 608
rect 5895 570 5896 580
rect 5911 570 5924 580
rect 5939 570 5969 584
rect 6012 570 6055 584
rect 6079 581 6086 588
rect 6089 584 6156 608
rect 6188 608 6360 610
rect 6158 586 6186 590
rect 6188 586 6268 608
rect 6289 606 6304 608
rect 6158 584 6268 586
rect 6089 580 6268 584
rect 6062 570 6092 580
rect 6094 570 6247 580
rect 6255 570 6285 580
rect 6289 570 6319 584
rect 6347 570 6360 608
rect 6432 614 6467 622
rect 6432 588 6433 614
rect 6440 588 6467 614
rect 6375 570 6405 584
rect 6432 580 6467 588
rect 6469 614 6510 622
rect 6469 588 6484 614
rect 6491 588 6510 614
rect 6574 610 6636 622
rect 6648 610 6723 622
rect 6781 610 6856 622
rect 6868 610 6899 622
rect 6905 610 6940 622
rect 6574 608 6736 610
rect 6469 580 6510 588
rect 6592 584 6605 608
rect 6620 606 6635 608
rect 6432 570 6433 580
rect 6448 570 6461 580
rect 6475 570 6476 580
rect 6491 570 6504 580
rect 6519 570 6549 584
rect 6592 570 6635 584
rect 6659 581 6666 588
rect 6669 584 6736 608
rect 6768 608 6940 610
rect 6738 586 6766 590
rect 6768 586 6848 608
rect 6869 606 6884 608
rect 6738 584 6848 586
rect 6669 580 6848 584
rect 6642 570 6672 580
rect 6674 570 6827 580
rect 6835 570 6865 580
rect 6869 570 6899 584
rect 6927 570 6940 608
rect 7012 614 7047 622
rect 7012 588 7013 614
rect 7020 588 7047 614
rect 6955 570 6985 584
rect 7012 580 7047 588
rect 7049 614 7090 622
rect 7049 588 7064 614
rect 7071 588 7090 614
rect 7154 610 7216 622
rect 7228 610 7303 622
rect 7361 610 7436 622
rect 7448 610 7479 622
rect 7485 610 7520 622
rect 7154 608 7316 610
rect 7049 580 7090 588
rect 7172 584 7185 608
rect 7200 606 7215 608
rect 7012 570 7013 580
rect 7028 570 7041 580
rect 7055 570 7056 580
rect 7071 570 7084 580
rect 7099 570 7129 584
rect 7172 570 7215 584
rect 7239 581 7246 588
rect 7249 584 7316 608
rect 7348 608 7520 610
rect 7318 586 7346 590
rect 7348 586 7428 608
rect 7449 606 7464 608
rect 7318 584 7428 586
rect 7249 580 7428 584
rect 7222 570 7252 580
rect 7254 570 7407 580
rect 7415 570 7445 580
rect 7449 570 7479 584
rect 7507 570 7520 608
rect 7592 614 7627 622
rect 7592 588 7593 614
rect 7600 588 7627 614
rect 7535 570 7565 584
rect 7592 580 7627 588
rect 7629 614 7670 622
rect 7629 588 7644 614
rect 7651 588 7670 614
rect 7734 610 7796 622
rect 7808 610 7883 622
rect 7941 610 8016 622
rect 8028 610 8059 622
rect 8065 610 8100 622
rect 7734 608 7896 610
rect 7629 580 7670 588
rect 7752 584 7765 608
rect 7780 606 7795 608
rect 7592 570 7593 580
rect 7608 570 7621 580
rect 7635 570 7636 580
rect 7651 570 7664 580
rect 7679 570 7709 584
rect 7752 570 7795 584
rect 7819 581 7826 588
rect 7829 584 7896 608
rect 7928 608 8100 610
rect 7898 586 7926 590
rect 7928 586 8008 608
rect 8029 606 8044 608
rect 7898 584 8008 586
rect 7829 580 8008 584
rect 7802 570 7832 580
rect 7834 570 7987 580
rect 7995 570 8025 580
rect 8029 570 8059 584
rect 8087 570 8100 608
rect 8172 614 8207 622
rect 8172 588 8173 614
rect 8180 588 8207 614
rect 8115 570 8145 584
rect 8172 580 8207 588
rect 8209 614 8250 622
rect 8209 588 8224 614
rect 8231 588 8250 614
rect 8314 610 8376 622
rect 8388 610 8463 622
rect 8521 610 8596 622
rect 8608 610 8639 622
rect 8645 610 8680 622
rect 8314 608 8476 610
rect 8209 580 8250 588
rect 8332 584 8345 608
rect 8360 606 8375 608
rect 8172 570 8173 580
rect 8188 570 8201 580
rect 8215 570 8216 580
rect 8231 570 8244 580
rect 8259 570 8289 584
rect 8332 570 8375 584
rect 8399 581 8406 588
rect 8409 584 8476 608
rect 8508 608 8680 610
rect 8478 586 8506 590
rect 8508 586 8588 608
rect 8609 606 8624 608
rect 8478 584 8588 586
rect 8409 580 8588 584
rect 8382 570 8412 580
rect 8414 570 8567 580
rect 8575 570 8605 580
rect 8609 570 8639 584
rect 8667 570 8680 608
rect 8752 614 8787 622
rect 8752 588 8753 614
rect 8760 588 8787 614
rect 8695 570 8725 584
rect 8752 580 8787 588
rect 8789 614 8830 622
rect 8789 588 8804 614
rect 8811 588 8830 614
rect 8894 610 8956 622
rect 8968 610 9043 622
rect 9101 610 9176 622
rect 9188 610 9219 622
rect 9225 610 9260 622
rect 8894 608 9056 610
rect 8789 580 8830 588
rect 8912 584 8925 608
rect 8940 606 8955 608
rect 8752 570 8753 580
rect 8768 570 8781 580
rect 8795 570 8796 580
rect 8811 570 8824 580
rect 8839 570 8869 584
rect 8912 570 8955 584
rect 8979 581 8986 588
rect 8989 584 9056 608
rect 9088 608 9260 610
rect 9058 586 9086 590
rect 9088 586 9168 608
rect 9189 606 9204 608
rect 9058 584 9168 586
rect 8989 580 9168 584
rect 8962 570 8992 580
rect 8994 570 9147 580
rect 9155 570 9185 580
rect 9189 570 9219 584
rect 9247 570 9260 608
rect 9332 614 9367 622
rect 9332 588 9333 614
rect 9340 588 9367 614
rect 9275 570 9305 584
rect 9332 580 9367 588
rect 9332 570 9333 580
rect 9348 570 9361 580
rect 5889 556 9361 570
rect 13 526 26 556
rect 41 538 71 556
rect 114 542 128 556
rect 164 542 384 556
rect 115 540 128 542
rect 81 528 96 540
rect 78 526 100 528
rect 105 526 135 540
rect 196 538 349 542
rect 178 526 370 538
rect 413 526 443 540
rect 449 526 462 556
rect 477 538 507 556
rect 550 526 563 556
rect 593 526 606 556
rect 621 538 651 556
rect 694 542 708 556
rect 744 542 964 556
rect 695 540 708 542
rect 661 528 676 540
rect 658 526 680 528
rect 685 526 715 540
rect 776 538 929 542
rect 758 526 950 538
rect 993 526 1023 540
rect 1029 526 1042 556
rect 1057 538 1087 556
rect 1130 526 1143 556
rect 1173 526 1186 556
rect 1201 538 1231 556
rect 1274 542 1288 556
rect 1324 542 1544 556
rect 1275 540 1288 542
rect 1241 528 1256 540
rect 1238 526 1260 528
rect 1265 526 1295 540
rect 1356 538 1509 542
rect 1338 526 1530 538
rect 1573 526 1603 540
rect 1609 526 1622 556
rect 1637 538 1667 556
rect 1710 526 1723 556
rect 1753 526 1766 556
rect 1781 538 1811 556
rect 1854 542 1868 556
rect 1904 542 2124 556
rect 1855 540 1868 542
rect 1821 528 1836 540
rect 1818 526 1840 528
rect 1845 526 1875 540
rect 1936 538 2089 542
rect 1918 526 2110 538
rect 2153 526 2183 540
rect 2189 526 2202 556
rect 2217 538 2247 556
rect 2290 526 2303 556
rect 2333 526 2346 556
rect 2361 538 2391 556
rect 2434 542 2448 556
rect 2484 542 2704 556
rect 2435 540 2448 542
rect 2401 528 2416 540
rect 2398 526 2420 528
rect 2425 526 2455 540
rect 2516 538 2669 542
rect 2498 526 2690 538
rect 2733 526 2763 540
rect 2769 526 2782 556
rect 2797 538 2827 556
rect 2870 526 2883 556
rect 2913 526 2926 556
rect 2941 538 2971 556
rect 3014 542 3028 556
rect 3064 542 3284 556
rect 3015 540 3028 542
rect 2981 528 2996 540
rect 2978 526 3000 528
rect 3005 526 3035 540
rect 3096 538 3249 542
rect 3078 526 3270 538
rect 3313 526 3343 540
rect 3349 526 3362 556
rect 3377 538 3407 556
rect 3450 526 3463 556
rect 5911 526 5924 556
rect 5939 538 5969 556
rect 6012 542 6026 556
rect 6062 542 6282 556
rect 6013 540 6026 542
rect 5979 528 5994 540
rect 5976 526 5998 528
rect 6003 526 6033 540
rect 6094 538 6247 542
rect 6076 526 6268 538
rect 6311 526 6341 540
rect 6347 526 6360 556
rect 6375 538 6405 556
rect 6448 526 6461 556
rect 6491 526 6504 556
rect 6519 538 6549 556
rect 6592 542 6606 556
rect 6642 542 6862 556
rect 6593 540 6606 542
rect 6559 528 6574 540
rect 6556 526 6578 528
rect 6583 526 6613 540
rect 6674 538 6827 542
rect 6656 526 6848 538
rect 6891 526 6921 540
rect 6927 526 6940 556
rect 6955 538 6985 556
rect 7028 526 7041 556
rect 7071 526 7084 556
rect 7099 538 7129 556
rect 7172 542 7186 556
rect 7222 542 7442 556
rect 7173 540 7186 542
rect 7139 528 7154 540
rect 7136 526 7158 528
rect 7163 526 7193 540
rect 7254 538 7407 542
rect 7236 526 7428 538
rect 7471 526 7501 540
rect 7507 526 7520 556
rect 7535 538 7565 556
rect 7608 526 7621 556
rect 7651 526 7664 556
rect 7679 538 7709 556
rect 7752 542 7766 556
rect 7802 542 8022 556
rect 7753 540 7766 542
rect 7719 528 7734 540
rect 7716 526 7738 528
rect 7743 526 7773 540
rect 7834 538 7987 542
rect 7816 526 8008 538
rect 8051 526 8081 540
rect 8087 526 8100 556
rect 8115 538 8145 556
rect 8188 526 8201 556
rect 8231 526 8244 556
rect 8259 538 8289 556
rect 8332 542 8346 556
rect 8382 542 8602 556
rect 8333 540 8346 542
rect 8299 528 8314 540
rect 8296 526 8318 528
rect 8323 526 8353 540
rect 8414 538 8567 542
rect 8396 526 8588 538
rect 8631 526 8661 540
rect 8667 526 8680 556
rect 8695 538 8725 556
rect 8768 526 8781 556
rect 8811 526 8824 556
rect 8839 538 8869 556
rect 8912 542 8926 556
rect 8962 542 9182 556
rect 8913 540 8926 542
rect 8879 528 8894 540
rect 8876 526 8898 528
rect 8903 526 8933 540
rect 8994 538 9147 542
rect 8976 526 9168 538
rect 9211 526 9241 540
rect 9247 526 9260 556
rect 9275 538 9305 556
rect 9348 526 9361 556
rect -2 512 3469 526
rect 5889 512 9361 526
rect 13 408 26 512
rect 71 490 72 500
rect 87 490 100 500
rect 71 486 100 490
rect 105 486 135 512
rect 153 498 169 500
rect 241 498 294 512
rect 242 496 306 498
rect 349 496 364 512
rect 413 509 443 512
rect 413 506 449 509
rect 379 498 395 500
rect 153 486 168 490
rect 71 484 168 486
rect 196 484 364 496
rect 380 486 395 490
rect 413 487 452 506
rect 471 500 478 501
rect 477 493 478 500
rect 461 490 462 493
rect 477 490 490 493
rect 413 486 443 487
rect 452 486 458 487
rect 461 486 490 490
rect 380 485 490 486
rect 380 484 496 485
rect 55 476 106 484
rect 55 464 80 476
rect 87 464 106 476
rect 137 476 187 484
rect 137 468 153 476
rect 160 474 187 476
rect 196 474 417 484
rect 160 464 417 474
rect 446 476 496 484
rect 446 467 462 476
rect 55 456 106 464
rect 153 456 417 464
rect 443 464 462 467
rect 469 464 496 476
rect 443 456 496 464
rect 71 448 72 456
rect 87 448 100 456
rect 71 440 87 448
rect 68 433 87 436
rect 68 424 90 433
rect 41 414 90 424
rect 41 408 71 414
rect 90 409 95 414
rect 13 392 87 408
rect 105 400 135 456
rect 170 446 378 456
rect 413 452 458 456
rect 461 455 462 456
rect 477 455 490 456
rect 196 416 385 446
rect 211 413 385 416
rect 204 410 385 413
rect 13 390 26 392
rect 41 390 75 392
rect 13 374 87 390
rect 114 386 127 400
rect 142 386 158 402
rect 204 397 215 410
rect -3 352 -2 368
rect 13 352 26 374
rect 41 352 71 374
rect 114 370 176 386
rect 204 379 215 395
rect 220 390 230 410
rect 240 390 254 410
rect 257 397 266 410
rect 282 397 291 410
rect 220 379 254 390
rect 257 379 266 395
rect 282 379 291 395
rect 298 390 308 410
rect 318 390 332 410
rect 333 397 344 410
rect 298 379 332 390
rect 333 379 344 395
rect 390 386 406 402
rect 413 400 443 452
rect 477 448 478 455
rect 462 440 478 448
rect 449 408 462 427
rect 477 408 507 424
rect 449 392 523 408
rect 449 390 462 392
rect 477 390 511 392
rect 114 368 127 370
rect 142 368 176 370
rect 114 352 176 368
rect 220 363 236 366
rect 298 363 328 374
rect 376 370 422 386
rect 449 374 523 390
rect 376 368 410 370
rect 375 352 422 368
rect 449 352 462 374
rect 477 352 507 374
rect 534 352 535 368
rect 550 352 563 512
rect 593 408 606 512
rect 651 490 652 500
rect 667 490 680 500
rect 651 486 680 490
rect 685 486 715 512
rect 733 498 749 500
rect 821 498 874 512
rect 822 496 886 498
rect 929 496 944 512
rect 993 509 1023 512
rect 993 506 1029 509
rect 959 498 975 500
rect 733 486 748 490
rect 651 484 748 486
rect 776 484 944 496
rect 960 486 975 490
rect 993 487 1032 506
rect 1051 500 1058 501
rect 1057 493 1058 500
rect 1041 490 1042 493
rect 1057 490 1070 493
rect 993 486 1023 487
rect 1032 486 1038 487
rect 1041 486 1070 490
rect 960 485 1070 486
rect 960 484 1076 485
rect 635 476 686 484
rect 635 464 660 476
rect 667 464 686 476
rect 717 476 767 484
rect 717 468 733 476
rect 740 474 767 476
rect 776 474 997 484
rect 740 464 997 474
rect 1026 476 1076 484
rect 1026 467 1042 476
rect 635 456 686 464
rect 733 456 997 464
rect 1023 464 1042 467
rect 1049 464 1076 476
rect 1023 456 1076 464
rect 651 448 652 456
rect 667 448 680 456
rect 651 440 667 448
rect 648 433 667 436
rect 648 424 670 433
rect 621 414 670 424
rect 621 408 651 414
rect 670 409 675 414
rect 593 392 667 408
rect 685 400 715 456
rect 750 446 958 456
rect 993 452 1038 456
rect 1041 455 1042 456
rect 1057 455 1070 456
rect 776 416 965 446
rect 791 413 965 416
rect 784 410 965 413
rect 593 390 606 392
rect 621 390 655 392
rect 593 374 667 390
rect 694 386 707 400
rect 722 386 738 402
rect 784 397 795 410
rect 577 352 578 368
rect 593 352 606 374
rect 621 352 651 374
rect 694 370 756 386
rect 784 379 795 395
rect 800 390 810 410
rect 820 390 834 410
rect 837 397 846 410
rect 862 397 871 410
rect 800 379 834 390
rect 837 379 846 395
rect 862 379 871 395
rect 878 390 888 410
rect 898 390 912 410
rect 913 397 924 410
rect 878 379 912 390
rect 913 379 924 395
rect 970 386 986 402
rect 993 400 1023 452
rect 1057 448 1058 455
rect 1042 440 1058 448
rect 1029 408 1042 427
rect 1057 408 1087 424
rect 1029 392 1103 408
rect 1029 390 1042 392
rect 1057 390 1091 392
rect 694 368 707 370
rect 722 368 756 370
rect 694 352 756 368
rect 800 363 816 366
rect 878 363 908 374
rect 956 370 1002 386
rect 1029 374 1103 390
rect 956 368 990 370
rect 955 352 1002 368
rect 1029 352 1042 374
rect 1057 352 1087 374
rect 1114 352 1115 368
rect 1130 352 1143 512
rect 1173 408 1186 512
rect 1231 490 1232 500
rect 1247 490 1260 500
rect 1231 486 1260 490
rect 1265 486 1295 512
rect 1313 498 1329 500
rect 1401 498 1454 512
rect 1402 496 1466 498
rect 1509 496 1524 512
rect 1573 509 1603 512
rect 1573 506 1609 509
rect 1539 498 1555 500
rect 1313 486 1328 490
rect 1231 484 1328 486
rect 1356 484 1524 496
rect 1540 486 1555 490
rect 1573 487 1612 506
rect 1631 500 1638 501
rect 1637 493 1638 500
rect 1621 490 1622 493
rect 1637 490 1650 493
rect 1573 486 1603 487
rect 1612 486 1618 487
rect 1621 486 1650 490
rect 1540 485 1650 486
rect 1540 484 1656 485
rect 1215 476 1266 484
rect 1215 464 1240 476
rect 1247 464 1266 476
rect 1297 476 1347 484
rect 1297 468 1313 476
rect 1320 474 1347 476
rect 1356 474 1577 484
rect 1320 464 1577 474
rect 1606 476 1656 484
rect 1606 467 1622 476
rect 1215 456 1266 464
rect 1313 456 1577 464
rect 1603 464 1622 467
rect 1629 464 1656 476
rect 1603 456 1656 464
rect 1231 448 1232 456
rect 1247 448 1260 456
rect 1231 440 1247 448
rect 1228 433 1247 436
rect 1228 424 1250 433
rect 1201 414 1250 424
rect 1201 408 1231 414
rect 1250 409 1255 414
rect 1173 392 1247 408
rect 1265 400 1295 456
rect 1330 446 1538 456
rect 1573 452 1618 456
rect 1621 455 1622 456
rect 1637 455 1650 456
rect 1356 416 1545 446
rect 1371 413 1545 416
rect 1364 410 1545 413
rect 1173 390 1186 392
rect 1201 390 1235 392
rect 1173 374 1247 390
rect 1274 386 1287 400
rect 1302 386 1318 402
rect 1364 397 1375 410
rect 1157 352 1158 368
rect 1173 352 1186 374
rect 1201 352 1231 374
rect 1274 370 1336 386
rect 1364 379 1375 395
rect 1380 390 1390 410
rect 1400 390 1414 410
rect 1417 397 1426 410
rect 1442 397 1451 410
rect 1380 379 1414 390
rect 1417 379 1426 395
rect 1442 379 1451 395
rect 1458 390 1468 410
rect 1478 390 1492 410
rect 1493 397 1504 410
rect 1458 379 1492 390
rect 1493 379 1504 395
rect 1550 386 1566 402
rect 1573 400 1603 452
rect 1637 448 1638 455
rect 1622 440 1638 448
rect 1609 408 1622 427
rect 1637 408 1667 424
rect 1609 392 1683 408
rect 1609 390 1622 392
rect 1637 390 1671 392
rect 1274 368 1287 370
rect 1302 368 1336 370
rect 1274 352 1336 368
rect 1380 363 1396 366
rect 1458 363 1488 374
rect 1536 370 1582 386
rect 1609 374 1683 390
rect 1536 368 1570 370
rect 1535 352 1582 368
rect 1609 352 1622 374
rect 1637 352 1667 374
rect 1694 352 1695 368
rect 1710 352 1723 512
rect 1753 408 1766 512
rect 1811 490 1812 500
rect 1827 490 1840 500
rect 1811 486 1840 490
rect 1845 486 1875 512
rect 1893 498 1909 500
rect 1981 498 2034 512
rect 1982 496 2046 498
rect 2089 496 2104 512
rect 2153 509 2183 512
rect 2153 506 2189 509
rect 2119 498 2135 500
rect 1893 486 1908 490
rect 1811 484 1908 486
rect 1936 484 2104 496
rect 2120 486 2135 490
rect 2153 487 2192 506
rect 2211 500 2218 501
rect 2217 493 2218 500
rect 2201 490 2202 493
rect 2217 490 2230 493
rect 2153 486 2183 487
rect 2192 486 2198 487
rect 2201 486 2230 490
rect 2120 485 2230 486
rect 2120 484 2236 485
rect 1795 476 1846 484
rect 1795 464 1820 476
rect 1827 464 1846 476
rect 1877 476 1927 484
rect 1877 468 1893 476
rect 1900 474 1927 476
rect 1936 474 2157 484
rect 1900 464 2157 474
rect 2186 476 2236 484
rect 2186 467 2202 476
rect 1795 456 1846 464
rect 1893 456 2157 464
rect 2183 464 2202 467
rect 2209 464 2236 476
rect 2183 456 2236 464
rect 1811 448 1812 456
rect 1827 448 1840 456
rect 1811 440 1827 448
rect 1808 433 1827 436
rect 1808 424 1830 433
rect 1781 414 1830 424
rect 1781 408 1811 414
rect 1830 409 1835 414
rect 1753 392 1827 408
rect 1845 400 1875 456
rect 1910 446 2118 456
rect 2153 452 2198 456
rect 2201 455 2202 456
rect 2217 455 2230 456
rect 1936 416 2125 446
rect 1951 413 2125 416
rect 1944 410 2125 413
rect 1753 390 1766 392
rect 1781 390 1815 392
rect 1753 374 1827 390
rect 1854 386 1867 400
rect 1882 386 1898 402
rect 1944 397 1955 410
rect 1737 352 1738 368
rect 1753 352 1766 374
rect 1781 352 1811 374
rect 1854 370 1916 386
rect 1944 379 1955 395
rect 1960 390 1970 410
rect 1980 390 1994 410
rect 1997 397 2006 410
rect 2022 397 2031 410
rect 1960 379 1994 390
rect 1997 379 2006 395
rect 2022 379 2031 395
rect 2038 390 2048 410
rect 2058 390 2072 410
rect 2073 397 2084 410
rect 2038 379 2072 390
rect 2073 379 2084 395
rect 2130 386 2146 402
rect 2153 400 2183 452
rect 2217 448 2218 455
rect 2202 440 2218 448
rect 2189 408 2202 427
rect 2217 408 2247 424
rect 2189 392 2263 408
rect 2189 390 2202 392
rect 2217 390 2251 392
rect 1854 368 1867 370
rect 1882 368 1916 370
rect 1854 352 1916 368
rect 1960 363 1976 366
rect 2038 363 2068 374
rect 2116 370 2162 386
rect 2189 374 2263 390
rect 2116 368 2150 370
rect 2115 352 2162 368
rect 2189 352 2202 374
rect 2217 352 2247 374
rect 2274 352 2275 368
rect 2290 352 2303 512
rect 2333 408 2346 512
rect 2391 490 2392 500
rect 2407 490 2420 500
rect 2391 486 2420 490
rect 2425 486 2455 512
rect 2473 498 2489 500
rect 2561 498 2614 512
rect 2562 496 2626 498
rect 2669 496 2684 512
rect 2733 509 2763 512
rect 2733 506 2769 509
rect 2699 498 2715 500
rect 2473 486 2488 490
rect 2391 484 2488 486
rect 2516 484 2684 496
rect 2700 486 2715 490
rect 2733 487 2772 506
rect 2791 500 2798 501
rect 2797 493 2798 500
rect 2781 490 2782 493
rect 2797 490 2810 493
rect 2733 486 2763 487
rect 2772 486 2778 487
rect 2781 486 2810 490
rect 2700 485 2810 486
rect 2700 484 2816 485
rect 2375 476 2426 484
rect 2375 464 2400 476
rect 2407 464 2426 476
rect 2457 476 2507 484
rect 2457 468 2473 476
rect 2480 474 2507 476
rect 2516 474 2737 484
rect 2480 464 2737 474
rect 2766 476 2816 484
rect 2766 467 2782 476
rect 2375 456 2426 464
rect 2473 456 2737 464
rect 2763 464 2782 467
rect 2789 464 2816 476
rect 2763 456 2816 464
rect 2391 448 2392 456
rect 2407 448 2420 456
rect 2391 440 2407 448
rect 2388 433 2407 436
rect 2388 424 2410 433
rect 2361 414 2410 424
rect 2361 408 2391 414
rect 2410 409 2415 414
rect 2333 392 2407 408
rect 2425 400 2455 456
rect 2490 446 2698 456
rect 2733 452 2778 456
rect 2781 455 2782 456
rect 2797 455 2810 456
rect 2516 416 2705 446
rect 2531 413 2705 416
rect 2524 410 2705 413
rect 2333 390 2346 392
rect 2361 390 2395 392
rect 2333 374 2407 390
rect 2434 386 2447 400
rect 2462 386 2478 402
rect 2524 397 2535 410
rect 2317 352 2318 368
rect 2333 352 2346 374
rect 2361 352 2391 374
rect 2434 370 2496 386
rect 2524 379 2535 395
rect 2540 390 2550 410
rect 2560 390 2574 410
rect 2577 397 2586 410
rect 2602 397 2611 410
rect 2540 379 2574 390
rect 2577 379 2586 395
rect 2602 379 2611 395
rect 2618 390 2628 410
rect 2638 390 2652 410
rect 2653 397 2664 410
rect 2618 379 2652 390
rect 2653 379 2664 395
rect 2710 386 2726 402
rect 2733 400 2763 452
rect 2797 448 2798 455
rect 2782 440 2798 448
rect 2769 408 2782 427
rect 2797 408 2827 424
rect 2769 392 2843 408
rect 2769 390 2782 392
rect 2797 390 2831 392
rect 2434 368 2447 370
rect 2462 368 2496 370
rect 2434 352 2496 368
rect 2540 363 2556 366
rect 2618 363 2648 374
rect 2696 370 2742 386
rect 2769 374 2843 390
rect 2696 368 2730 370
rect 2695 352 2742 368
rect 2769 352 2782 374
rect 2797 352 2827 374
rect 2854 352 2855 368
rect 2870 352 2883 512
rect 2913 408 2926 512
rect 2971 490 2972 500
rect 2987 490 3000 500
rect 2971 486 3000 490
rect 3005 486 3035 512
rect 3053 498 3069 500
rect 3141 498 3194 512
rect 3142 496 3206 498
rect 3249 496 3264 512
rect 3313 509 3343 512
rect 3313 506 3349 509
rect 3279 498 3295 500
rect 3053 486 3068 490
rect 2971 484 3068 486
rect 3096 484 3264 496
rect 3280 486 3295 490
rect 3313 487 3352 506
rect 3371 500 3378 501
rect 3377 493 3378 500
rect 3361 490 3362 493
rect 3377 490 3390 493
rect 3313 486 3343 487
rect 3352 486 3358 487
rect 3361 486 3390 490
rect 3280 485 3390 486
rect 3280 484 3396 485
rect 2955 476 3006 484
rect 2955 464 2980 476
rect 2987 464 3006 476
rect 3037 476 3087 484
rect 3037 468 3053 476
rect 3060 474 3087 476
rect 3096 474 3317 484
rect 3060 464 3317 474
rect 3346 476 3396 484
rect 3346 467 3362 476
rect 2955 456 3006 464
rect 3053 456 3317 464
rect 3343 464 3362 467
rect 3369 464 3396 476
rect 3343 456 3396 464
rect 2971 448 2972 456
rect 2987 448 3000 456
rect 2971 440 2987 448
rect 2968 433 2987 436
rect 2968 424 2990 433
rect 2941 414 2990 424
rect 2941 408 2971 414
rect 2990 409 2995 414
rect 2913 392 2987 408
rect 3005 400 3035 456
rect 3070 446 3278 456
rect 3313 452 3358 456
rect 3361 455 3362 456
rect 3377 455 3390 456
rect 3096 416 3285 446
rect 3111 413 3285 416
rect 3104 410 3285 413
rect 2913 390 2926 392
rect 2941 390 2975 392
rect 2913 374 2987 390
rect 3014 386 3027 400
rect 3042 386 3058 402
rect 3104 397 3115 410
rect 2897 352 2898 368
rect 2913 352 2926 374
rect 2941 352 2971 374
rect 3014 370 3076 386
rect 3104 379 3115 395
rect 3120 390 3130 410
rect 3140 390 3154 410
rect 3157 397 3166 410
rect 3182 397 3191 410
rect 3120 379 3154 390
rect 3157 379 3166 395
rect 3182 379 3191 395
rect 3198 390 3208 410
rect 3218 390 3232 410
rect 3233 397 3244 410
rect 3198 379 3232 390
rect 3233 379 3244 395
rect 3290 386 3306 402
rect 3313 400 3343 452
rect 3377 448 3378 455
rect 3362 440 3378 448
rect 3349 408 3362 427
rect 3377 408 3407 424
rect 3349 392 3423 408
rect 3349 390 3362 392
rect 3377 390 3411 392
rect 3014 368 3027 370
rect 3042 368 3076 370
rect 3014 352 3076 368
rect 3120 363 3136 366
rect 3198 363 3228 374
rect 3276 370 3322 386
rect 3349 374 3423 390
rect 3276 368 3310 370
rect 3275 352 3322 368
rect 3349 352 3362 374
rect 3377 352 3407 374
rect 3434 352 3435 368
rect 3450 352 3463 512
rect 5911 408 5924 512
rect 5969 490 5970 500
rect 5985 490 5998 500
rect 5969 486 5998 490
rect 6003 486 6033 512
rect 6051 498 6067 500
rect 6139 498 6192 512
rect 6140 496 6204 498
rect 6247 496 6262 512
rect 6311 509 6341 512
rect 6311 506 6347 509
rect 6277 498 6293 500
rect 6051 486 6066 490
rect 5969 484 6066 486
rect 6094 484 6262 496
rect 6278 486 6293 490
rect 6311 487 6350 506
rect 6369 500 6376 501
rect 6375 493 6376 500
rect 6359 490 6360 493
rect 6375 490 6388 493
rect 6311 486 6341 487
rect 6350 486 6356 487
rect 6359 486 6388 490
rect 6278 485 6388 486
rect 6278 484 6394 485
rect 5953 476 6004 484
rect 5953 464 5978 476
rect 5985 464 6004 476
rect 6035 476 6085 484
rect 6035 468 6051 476
rect 6058 474 6085 476
rect 6094 474 6315 484
rect 6058 464 6315 474
rect 6344 476 6394 484
rect 6344 467 6360 476
rect 5953 456 6004 464
rect 6051 456 6315 464
rect 6341 464 6360 467
rect 6367 464 6394 476
rect 6341 456 6394 464
rect 5969 448 5970 456
rect 5985 448 5998 456
rect 5969 440 5985 448
rect 5966 433 5985 436
rect 5966 424 5988 433
rect 5939 414 5988 424
rect 5939 408 5969 414
rect 5988 409 5993 414
rect 5911 392 5985 408
rect 6003 400 6033 456
rect 6068 446 6276 456
rect 6311 452 6356 456
rect 6359 455 6360 456
rect 6375 455 6388 456
rect 6094 416 6283 446
rect 6109 413 6283 416
rect 6102 410 6283 413
rect 5911 390 5924 392
rect 5939 390 5973 392
rect 5911 374 5985 390
rect 6012 386 6025 400
rect 6040 386 6056 402
rect 6102 397 6113 410
rect 5895 352 5896 368
rect 5911 352 5924 374
rect 5939 352 5969 374
rect 6012 370 6074 386
rect 6102 379 6113 395
rect 6118 390 6128 410
rect 6138 390 6152 410
rect 6155 397 6164 410
rect 6180 397 6189 410
rect 6118 379 6152 390
rect 6155 379 6164 395
rect 6180 379 6189 395
rect 6196 390 6206 410
rect 6216 390 6230 410
rect 6231 397 6242 410
rect 6196 379 6230 390
rect 6231 379 6242 395
rect 6288 386 6304 402
rect 6311 400 6341 452
rect 6375 448 6376 455
rect 6360 440 6376 448
rect 6347 408 6360 427
rect 6375 408 6405 424
rect 6347 392 6421 408
rect 6347 390 6360 392
rect 6375 390 6409 392
rect 6012 368 6025 370
rect 6040 368 6074 370
rect 6012 352 6074 368
rect 6118 363 6134 366
rect 6196 363 6226 374
rect 6274 370 6320 386
rect 6347 374 6421 390
rect 6274 368 6308 370
rect 6273 352 6320 368
rect 6347 352 6360 374
rect 6375 352 6405 374
rect 6432 352 6433 368
rect 6448 352 6461 512
rect 6491 408 6504 512
rect 6549 490 6550 500
rect 6565 490 6578 500
rect 6549 486 6578 490
rect 6583 486 6613 512
rect 6631 498 6647 500
rect 6719 498 6772 512
rect 6720 496 6784 498
rect 6827 496 6842 512
rect 6891 509 6921 512
rect 6891 506 6927 509
rect 6857 498 6873 500
rect 6631 486 6646 490
rect 6549 484 6646 486
rect 6674 484 6842 496
rect 6858 486 6873 490
rect 6891 487 6930 506
rect 6949 500 6956 501
rect 6955 493 6956 500
rect 6939 490 6940 493
rect 6955 490 6968 493
rect 6891 486 6921 487
rect 6930 486 6936 487
rect 6939 486 6968 490
rect 6858 485 6968 486
rect 6858 484 6974 485
rect 6533 476 6584 484
rect 6533 464 6558 476
rect 6565 464 6584 476
rect 6615 476 6665 484
rect 6615 468 6631 476
rect 6638 474 6665 476
rect 6674 474 6895 484
rect 6638 464 6895 474
rect 6924 476 6974 484
rect 6924 467 6940 476
rect 6533 456 6584 464
rect 6631 456 6895 464
rect 6921 464 6940 467
rect 6947 464 6974 476
rect 6921 456 6974 464
rect 6549 448 6550 456
rect 6565 448 6578 456
rect 6549 440 6565 448
rect 6546 433 6565 436
rect 6546 424 6568 433
rect 6519 414 6568 424
rect 6519 408 6549 414
rect 6568 409 6573 414
rect 6491 392 6565 408
rect 6583 400 6613 456
rect 6648 446 6856 456
rect 6891 452 6936 456
rect 6939 455 6940 456
rect 6955 455 6968 456
rect 6674 416 6863 446
rect 6689 413 6863 416
rect 6682 410 6863 413
rect 6491 390 6504 392
rect 6519 390 6553 392
rect 6491 374 6565 390
rect 6592 386 6605 400
rect 6620 386 6636 402
rect 6682 397 6693 410
rect 6475 352 6476 368
rect 6491 352 6504 374
rect 6519 352 6549 374
rect 6592 370 6654 386
rect 6682 379 6693 395
rect 6698 390 6708 410
rect 6718 390 6732 410
rect 6735 397 6744 410
rect 6760 397 6769 410
rect 6698 379 6732 390
rect 6735 379 6744 395
rect 6760 379 6769 395
rect 6776 390 6786 410
rect 6796 390 6810 410
rect 6811 397 6822 410
rect 6776 379 6810 390
rect 6811 379 6822 395
rect 6868 386 6884 402
rect 6891 400 6921 452
rect 6955 448 6956 455
rect 6940 440 6956 448
rect 6927 408 6940 427
rect 6955 408 6985 424
rect 6927 392 7001 408
rect 6927 390 6940 392
rect 6955 390 6989 392
rect 6592 368 6605 370
rect 6620 368 6654 370
rect 6592 352 6654 368
rect 6698 363 6714 366
rect 6776 363 6806 374
rect 6854 370 6900 386
rect 6927 374 7001 390
rect 6854 368 6888 370
rect 6853 352 6900 368
rect 6927 352 6940 374
rect 6955 352 6985 374
rect 7012 352 7013 368
rect 7028 352 7041 512
rect 7071 408 7084 512
rect 7129 490 7130 500
rect 7145 490 7158 500
rect 7129 486 7158 490
rect 7163 486 7193 512
rect 7211 498 7227 500
rect 7299 498 7352 512
rect 7300 496 7364 498
rect 7407 496 7422 512
rect 7471 509 7501 512
rect 7471 506 7507 509
rect 7437 498 7453 500
rect 7211 486 7226 490
rect 7129 484 7226 486
rect 7254 484 7422 496
rect 7438 486 7453 490
rect 7471 487 7510 506
rect 7529 500 7536 501
rect 7535 493 7536 500
rect 7519 490 7520 493
rect 7535 490 7548 493
rect 7471 486 7501 487
rect 7510 486 7516 487
rect 7519 486 7548 490
rect 7438 485 7548 486
rect 7438 484 7554 485
rect 7113 476 7164 484
rect 7113 464 7138 476
rect 7145 464 7164 476
rect 7195 476 7245 484
rect 7195 468 7211 476
rect 7218 474 7245 476
rect 7254 474 7475 484
rect 7218 464 7475 474
rect 7504 476 7554 484
rect 7504 467 7520 476
rect 7113 456 7164 464
rect 7211 456 7475 464
rect 7501 464 7520 467
rect 7527 464 7554 476
rect 7501 456 7554 464
rect 7129 448 7130 456
rect 7145 448 7158 456
rect 7129 440 7145 448
rect 7126 433 7145 436
rect 7126 424 7148 433
rect 7099 414 7148 424
rect 7099 408 7129 414
rect 7148 409 7153 414
rect 7071 392 7145 408
rect 7163 400 7193 456
rect 7228 446 7436 456
rect 7471 452 7516 456
rect 7519 455 7520 456
rect 7535 455 7548 456
rect 7254 416 7443 446
rect 7269 413 7443 416
rect 7262 410 7443 413
rect 7071 390 7084 392
rect 7099 390 7133 392
rect 7071 374 7145 390
rect 7172 386 7185 400
rect 7200 386 7216 402
rect 7262 397 7273 410
rect 7055 352 7056 368
rect 7071 352 7084 374
rect 7099 352 7129 374
rect 7172 370 7234 386
rect 7262 379 7273 395
rect 7278 390 7288 410
rect 7298 390 7312 410
rect 7315 397 7324 410
rect 7340 397 7349 410
rect 7278 379 7312 390
rect 7315 379 7324 395
rect 7340 379 7349 395
rect 7356 390 7366 410
rect 7376 390 7390 410
rect 7391 397 7402 410
rect 7356 379 7390 390
rect 7391 379 7402 395
rect 7448 386 7464 402
rect 7471 400 7501 452
rect 7535 448 7536 455
rect 7520 440 7536 448
rect 7507 408 7520 427
rect 7535 408 7565 424
rect 7507 392 7581 408
rect 7507 390 7520 392
rect 7535 390 7569 392
rect 7172 368 7185 370
rect 7200 368 7234 370
rect 7172 352 7234 368
rect 7278 363 7294 366
rect 7356 363 7386 374
rect 7434 370 7480 386
rect 7507 374 7581 390
rect 7434 368 7468 370
rect 7433 352 7480 368
rect 7507 352 7520 374
rect 7535 352 7565 374
rect 7592 352 7593 368
rect 7608 352 7621 512
rect 7651 408 7664 512
rect 7709 490 7710 500
rect 7725 490 7738 500
rect 7709 486 7738 490
rect 7743 486 7773 512
rect 7791 498 7807 500
rect 7879 498 7932 512
rect 7880 496 7944 498
rect 7987 496 8002 512
rect 8051 509 8081 512
rect 8051 506 8087 509
rect 8017 498 8033 500
rect 7791 486 7806 490
rect 7709 484 7806 486
rect 7834 484 8002 496
rect 8018 486 8033 490
rect 8051 487 8090 506
rect 8109 500 8116 501
rect 8115 493 8116 500
rect 8099 490 8100 493
rect 8115 490 8128 493
rect 8051 486 8081 487
rect 8090 486 8096 487
rect 8099 486 8128 490
rect 8018 485 8128 486
rect 8018 484 8134 485
rect 7693 476 7744 484
rect 7693 464 7718 476
rect 7725 464 7744 476
rect 7775 476 7825 484
rect 7775 468 7791 476
rect 7798 474 7825 476
rect 7834 474 8055 484
rect 7798 464 8055 474
rect 8084 476 8134 484
rect 8084 467 8100 476
rect 7693 456 7744 464
rect 7791 456 8055 464
rect 8081 464 8100 467
rect 8107 464 8134 476
rect 8081 456 8134 464
rect 7709 448 7710 456
rect 7725 448 7738 456
rect 7709 440 7725 448
rect 7706 433 7725 436
rect 7706 424 7728 433
rect 7679 414 7728 424
rect 7679 408 7709 414
rect 7728 409 7733 414
rect 7651 392 7725 408
rect 7743 400 7773 456
rect 7808 446 8016 456
rect 8051 452 8096 456
rect 8099 455 8100 456
rect 8115 455 8128 456
rect 7834 416 8023 446
rect 7849 413 8023 416
rect 7842 410 8023 413
rect 7651 390 7664 392
rect 7679 390 7713 392
rect 7651 374 7725 390
rect 7752 386 7765 400
rect 7780 386 7796 402
rect 7842 397 7853 410
rect 7635 352 7636 368
rect 7651 352 7664 374
rect 7679 352 7709 374
rect 7752 370 7814 386
rect 7842 379 7853 395
rect 7858 390 7868 410
rect 7878 390 7892 410
rect 7895 397 7904 410
rect 7920 397 7929 410
rect 7858 379 7892 390
rect 7895 379 7904 395
rect 7920 379 7929 395
rect 7936 390 7946 410
rect 7956 390 7970 410
rect 7971 397 7982 410
rect 7936 379 7970 390
rect 7971 379 7982 395
rect 8028 386 8044 402
rect 8051 400 8081 452
rect 8115 448 8116 455
rect 8100 440 8116 448
rect 8087 408 8100 427
rect 8115 408 8145 424
rect 8087 392 8161 408
rect 8087 390 8100 392
rect 8115 390 8149 392
rect 7752 368 7765 370
rect 7780 368 7814 370
rect 7752 352 7814 368
rect 7858 363 7874 366
rect 7936 363 7966 374
rect 8014 370 8060 386
rect 8087 374 8161 390
rect 8014 368 8048 370
rect 8013 352 8060 368
rect 8087 352 8100 374
rect 8115 352 8145 374
rect 8172 352 8173 368
rect 8188 352 8201 512
rect 8231 408 8244 512
rect 8289 490 8290 500
rect 8305 490 8318 500
rect 8289 486 8318 490
rect 8323 486 8353 512
rect 8371 498 8387 500
rect 8459 498 8512 512
rect 8460 496 8524 498
rect 8567 496 8582 512
rect 8631 509 8661 512
rect 8631 506 8667 509
rect 8597 498 8613 500
rect 8371 486 8386 490
rect 8289 484 8386 486
rect 8414 484 8582 496
rect 8598 486 8613 490
rect 8631 487 8670 506
rect 8689 500 8696 501
rect 8695 493 8696 500
rect 8679 490 8680 493
rect 8695 490 8708 493
rect 8631 486 8661 487
rect 8670 486 8676 487
rect 8679 486 8708 490
rect 8598 485 8708 486
rect 8598 484 8714 485
rect 8273 476 8324 484
rect 8273 464 8298 476
rect 8305 464 8324 476
rect 8355 476 8405 484
rect 8355 468 8371 476
rect 8378 474 8405 476
rect 8414 474 8635 484
rect 8378 464 8635 474
rect 8664 476 8714 484
rect 8664 467 8680 476
rect 8273 456 8324 464
rect 8371 456 8635 464
rect 8661 464 8680 467
rect 8687 464 8714 476
rect 8661 456 8714 464
rect 8289 448 8290 456
rect 8305 448 8318 456
rect 8289 440 8305 448
rect 8286 433 8305 436
rect 8286 424 8308 433
rect 8259 414 8308 424
rect 8259 408 8289 414
rect 8308 409 8313 414
rect 8231 392 8305 408
rect 8323 400 8353 456
rect 8388 446 8596 456
rect 8631 452 8676 456
rect 8679 455 8680 456
rect 8695 455 8708 456
rect 8414 416 8603 446
rect 8429 413 8603 416
rect 8422 410 8603 413
rect 8231 390 8244 392
rect 8259 390 8293 392
rect 8231 374 8305 390
rect 8332 386 8345 400
rect 8360 386 8376 402
rect 8422 397 8433 410
rect 8215 352 8216 368
rect 8231 352 8244 374
rect 8259 352 8289 374
rect 8332 370 8394 386
rect 8422 379 8433 395
rect 8438 390 8448 410
rect 8458 390 8472 410
rect 8475 397 8484 410
rect 8500 397 8509 410
rect 8438 379 8472 390
rect 8475 379 8484 395
rect 8500 379 8509 395
rect 8516 390 8526 410
rect 8536 390 8550 410
rect 8551 397 8562 410
rect 8516 379 8550 390
rect 8551 379 8562 395
rect 8608 386 8624 402
rect 8631 400 8661 452
rect 8695 448 8696 455
rect 8680 440 8696 448
rect 8667 408 8680 427
rect 8695 408 8725 424
rect 8667 392 8741 408
rect 8667 390 8680 392
rect 8695 390 8729 392
rect 8332 368 8345 370
rect 8360 368 8394 370
rect 8332 352 8394 368
rect 8438 363 8454 366
rect 8516 363 8546 374
rect 8594 370 8640 386
rect 8667 374 8741 390
rect 8594 368 8628 370
rect 8593 352 8640 368
rect 8667 352 8680 374
rect 8695 352 8725 374
rect 8752 352 8753 368
rect 8768 352 8781 512
rect 8811 408 8824 512
rect 8869 490 8870 500
rect 8885 490 8898 500
rect 8869 486 8898 490
rect 8903 486 8933 512
rect 8951 498 8967 500
rect 9039 498 9092 512
rect 9040 496 9104 498
rect 9147 496 9162 512
rect 9211 509 9241 512
rect 9211 506 9247 509
rect 9177 498 9193 500
rect 8951 486 8966 490
rect 8869 484 8966 486
rect 8994 484 9162 496
rect 9178 486 9193 490
rect 9211 487 9250 506
rect 9269 500 9276 501
rect 9275 493 9276 500
rect 9259 490 9260 493
rect 9275 490 9288 493
rect 9211 486 9241 487
rect 9250 486 9256 487
rect 9259 486 9288 490
rect 9178 485 9288 486
rect 9178 484 9294 485
rect 8853 476 8904 484
rect 8853 464 8878 476
rect 8885 464 8904 476
rect 8935 476 8985 484
rect 8935 468 8951 476
rect 8958 474 8985 476
rect 8994 474 9215 484
rect 8958 464 9215 474
rect 9244 476 9294 484
rect 9244 467 9260 476
rect 8853 456 8904 464
rect 8951 456 9215 464
rect 9241 464 9260 467
rect 9267 464 9294 476
rect 9241 456 9294 464
rect 8869 448 8870 456
rect 8885 448 8898 456
rect 8869 440 8885 448
rect 8866 433 8885 436
rect 8866 424 8888 433
rect 8839 414 8888 424
rect 8839 408 8869 414
rect 8888 409 8893 414
rect 8811 392 8885 408
rect 8903 400 8933 456
rect 8968 446 9176 456
rect 9211 452 9256 456
rect 9259 455 9260 456
rect 9275 455 9288 456
rect 8994 416 9183 446
rect 9009 413 9183 416
rect 9002 410 9183 413
rect 8811 390 8824 392
rect 8839 390 8873 392
rect 8811 374 8885 390
rect 8912 386 8925 400
rect 8940 386 8956 402
rect 9002 397 9013 410
rect 8795 352 8796 368
rect 8811 352 8824 374
rect 8839 352 8869 374
rect 8912 370 8974 386
rect 9002 379 9013 395
rect 9018 390 9028 410
rect 9038 390 9052 410
rect 9055 397 9064 410
rect 9080 397 9089 410
rect 9018 379 9052 390
rect 9055 379 9064 395
rect 9080 379 9089 395
rect 9096 390 9106 410
rect 9116 390 9130 410
rect 9131 397 9142 410
rect 9096 379 9130 390
rect 9131 379 9142 395
rect 9188 386 9204 402
rect 9211 400 9241 452
rect 9275 448 9276 455
rect 9260 440 9276 448
rect 9247 408 9260 427
rect 9275 408 9305 424
rect 9247 392 9321 408
rect 9247 390 9260 392
rect 9275 390 9309 392
rect 8912 368 8925 370
rect 8940 368 8974 370
rect 8912 352 8974 368
rect 9018 363 9034 366
rect 9096 363 9126 374
rect 9174 370 9220 386
rect 9247 374 9321 390
rect 9174 368 9208 370
rect 9173 352 9220 368
rect 9247 352 9260 374
rect 9275 352 9305 374
rect 9332 352 9333 368
rect 9348 352 9361 512
rect -9 344 32 352
rect -9 318 6 344
rect 13 318 32 344
rect 96 340 158 352
rect 170 340 245 352
rect 303 340 378 352
rect 390 340 421 352
rect 427 340 462 352
rect 96 338 258 340
rect -9 310 32 318
rect 114 314 127 338
rect 142 336 157 338
rect -3 300 -2 310
rect 13 300 26 310
rect 41 300 71 314
rect 114 300 157 314
rect 181 311 188 318
rect 191 314 258 338
rect 290 338 462 340
rect 260 316 288 320
rect 290 316 370 338
rect 391 336 406 338
rect 260 314 370 316
rect 191 310 370 314
rect 164 300 194 310
rect 196 300 349 310
rect 357 300 387 310
rect 391 300 421 314
rect 449 300 462 338
rect 534 344 569 352
rect 534 318 535 344
rect 542 318 569 344
rect 477 300 507 314
rect 534 310 569 318
rect 571 344 612 352
rect 571 318 586 344
rect 593 318 612 344
rect 676 340 738 352
rect 750 340 825 352
rect 883 340 958 352
rect 970 340 1001 352
rect 1007 340 1042 352
rect 676 338 838 340
rect 571 310 612 318
rect 694 314 707 338
rect 722 336 737 338
rect 534 300 535 310
rect 550 300 563 310
rect 577 300 578 310
rect 593 300 606 310
rect 621 300 651 314
rect 694 300 737 314
rect 761 311 768 318
rect 771 314 838 338
rect 870 338 1042 340
rect 840 316 868 320
rect 870 316 950 338
rect 971 336 986 338
rect 840 314 950 316
rect 771 310 950 314
rect 744 300 774 310
rect 776 300 929 310
rect 937 300 967 310
rect 971 300 1001 314
rect 1029 300 1042 338
rect 1114 344 1149 352
rect 1114 318 1115 344
rect 1122 318 1149 344
rect 1057 300 1087 314
rect 1114 310 1149 318
rect 1151 344 1192 352
rect 1151 318 1166 344
rect 1173 318 1192 344
rect 1256 340 1318 352
rect 1330 340 1405 352
rect 1463 340 1538 352
rect 1550 340 1581 352
rect 1587 340 1622 352
rect 1256 338 1418 340
rect 1151 310 1192 318
rect 1274 314 1287 338
rect 1302 336 1317 338
rect 1114 300 1115 310
rect 1130 300 1143 310
rect 1157 300 1158 310
rect 1173 300 1186 310
rect 1201 300 1231 314
rect 1274 300 1317 314
rect 1341 311 1348 318
rect 1351 314 1418 338
rect 1450 338 1622 340
rect 1420 316 1448 320
rect 1450 316 1530 338
rect 1551 336 1566 338
rect 1420 314 1530 316
rect 1351 310 1530 314
rect 1324 300 1354 310
rect 1356 300 1509 310
rect 1517 300 1547 310
rect 1551 300 1581 314
rect 1609 300 1622 338
rect 1694 344 1729 352
rect 1694 318 1695 344
rect 1702 318 1729 344
rect 1637 300 1667 314
rect 1694 310 1729 318
rect 1731 344 1772 352
rect 1731 318 1746 344
rect 1753 318 1772 344
rect 1836 340 1898 352
rect 1910 340 1985 352
rect 2043 340 2118 352
rect 2130 340 2161 352
rect 2167 340 2202 352
rect 1836 338 1998 340
rect 1731 310 1772 318
rect 1854 314 1867 338
rect 1882 336 1897 338
rect 1694 300 1695 310
rect 1710 300 1723 310
rect 1737 300 1738 310
rect 1753 300 1766 310
rect 1781 300 1811 314
rect 1854 300 1897 314
rect 1921 311 1928 318
rect 1931 314 1998 338
rect 2030 338 2202 340
rect 2000 316 2028 320
rect 2030 316 2110 338
rect 2131 336 2146 338
rect 2000 314 2110 316
rect 1931 310 2110 314
rect 1904 300 1934 310
rect 1936 300 2089 310
rect 2097 300 2127 310
rect 2131 300 2161 314
rect 2189 300 2202 338
rect 2274 344 2309 352
rect 2274 318 2275 344
rect 2282 318 2309 344
rect 2217 300 2247 314
rect 2274 310 2309 318
rect 2311 344 2352 352
rect 2311 318 2326 344
rect 2333 318 2352 344
rect 2416 340 2478 352
rect 2490 340 2565 352
rect 2623 340 2698 352
rect 2710 340 2741 352
rect 2747 340 2782 352
rect 2416 338 2578 340
rect 2311 310 2352 318
rect 2434 314 2447 338
rect 2462 336 2477 338
rect 2274 300 2275 310
rect 2290 300 2303 310
rect 2317 300 2318 310
rect 2333 300 2346 310
rect 2361 300 2391 314
rect 2434 300 2477 314
rect 2501 311 2508 318
rect 2511 314 2578 338
rect 2610 338 2782 340
rect 2580 316 2608 320
rect 2610 316 2690 338
rect 2711 336 2726 338
rect 2580 314 2690 316
rect 2511 310 2690 314
rect 2484 300 2514 310
rect 2516 300 2669 310
rect 2677 300 2707 310
rect 2711 300 2741 314
rect 2769 300 2782 338
rect 2854 344 2889 352
rect 2854 318 2855 344
rect 2862 318 2889 344
rect 2797 300 2827 314
rect 2854 310 2889 318
rect 2891 344 2932 352
rect 2891 318 2906 344
rect 2913 318 2932 344
rect 2996 340 3058 352
rect 3070 340 3145 352
rect 3203 340 3278 352
rect 3290 340 3321 352
rect 3327 340 3362 352
rect 2996 338 3158 340
rect 2891 310 2932 318
rect 3014 314 3027 338
rect 3042 336 3057 338
rect 2854 300 2855 310
rect 2870 300 2883 310
rect 2897 300 2898 310
rect 2913 300 2926 310
rect 2941 300 2971 314
rect 3014 300 3057 314
rect 3081 311 3088 318
rect 3091 314 3158 338
rect 3190 338 3362 340
rect 3160 316 3188 320
rect 3190 316 3270 338
rect 3291 336 3306 338
rect 3160 314 3270 316
rect 3091 310 3270 314
rect 3064 300 3094 310
rect 3096 300 3249 310
rect 3257 300 3287 310
rect 3291 300 3321 314
rect 3349 300 3362 338
rect 3434 344 3469 352
rect 3434 318 3435 344
rect 3442 318 3469 344
rect 3377 300 3407 314
rect 3434 310 3469 318
rect 3434 300 3435 310
rect 3450 300 3463 310
rect -3 294 3469 300
rect -2 286 3469 294
rect 5889 344 5930 352
rect 5889 318 5904 344
rect 5911 318 5930 344
rect 5994 340 6056 352
rect 6068 340 6143 352
rect 6201 340 6276 352
rect 6288 340 6319 352
rect 6325 340 6360 352
rect 5994 338 6156 340
rect 5889 310 5930 318
rect 6012 314 6025 338
rect 6040 336 6055 338
rect 5895 300 5896 310
rect 5911 300 5924 310
rect 5939 300 5969 314
rect 6012 300 6055 314
rect 6079 311 6086 318
rect 6089 314 6156 338
rect 6188 338 6360 340
rect 6158 316 6186 320
rect 6188 316 6268 338
rect 6289 336 6304 338
rect 6158 314 6268 316
rect 6089 310 6268 314
rect 6062 300 6092 310
rect 6094 300 6247 310
rect 6255 300 6285 310
rect 6289 300 6319 314
rect 6347 300 6360 338
rect 6432 344 6467 352
rect 6432 318 6433 344
rect 6440 318 6467 344
rect 6375 300 6405 314
rect 6432 310 6467 318
rect 6469 344 6510 352
rect 6469 318 6484 344
rect 6491 318 6510 344
rect 6574 340 6636 352
rect 6648 340 6723 352
rect 6781 340 6856 352
rect 6868 340 6899 352
rect 6905 340 6940 352
rect 6574 338 6736 340
rect 6469 310 6510 318
rect 6592 314 6605 338
rect 6620 336 6635 338
rect 6432 300 6433 310
rect 6448 300 6461 310
rect 6475 300 6476 310
rect 6491 300 6504 310
rect 6519 300 6549 314
rect 6592 300 6635 314
rect 6659 311 6666 318
rect 6669 314 6736 338
rect 6768 338 6940 340
rect 6738 316 6766 320
rect 6768 316 6848 338
rect 6869 336 6884 338
rect 6738 314 6848 316
rect 6669 310 6848 314
rect 6642 300 6672 310
rect 6674 300 6827 310
rect 6835 300 6865 310
rect 6869 300 6899 314
rect 6927 300 6940 338
rect 7012 344 7047 352
rect 7012 318 7013 344
rect 7020 318 7047 344
rect 6955 300 6985 314
rect 7012 310 7047 318
rect 7049 344 7090 352
rect 7049 318 7064 344
rect 7071 318 7090 344
rect 7154 340 7216 352
rect 7228 340 7303 352
rect 7361 340 7436 352
rect 7448 340 7479 352
rect 7485 340 7520 352
rect 7154 338 7316 340
rect 7049 310 7090 318
rect 7172 314 7185 338
rect 7200 336 7215 338
rect 7012 300 7013 310
rect 7028 300 7041 310
rect 7055 300 7056 310
rect 7071 300 7084 310
rect 7099 300 7129 314
rect 7172 300 7215 314
rect 7239 311 7246 318
rect 7249 314 7316 338
rect 7348 338 7520 340
rect 7318 316 7346 320
rect 7348 316 7428 338
rect 7449 336 7464 338
rect 7318 314 7428 316
rect 7249 310 7428 314
rect 7222 300 7252 310
rect 7254 300 7407 310
rect 7415 300 7445 310
rect 7449 300 7479 314
rect 7507 300 7520 338
rect 7592 344 7627 352
rect 7592 318 7593 344
rect 7600 318 7627 344
rect 7535 300 7565 314
rect 7592 310 7627 318
rect 7629 344 7670 352
rect 7629 318 7644 344
rect 7651 318 7670 344
rect 7734 340 7796 352
rect 7808 340 7883 352
rect 7941 340 8016 352
rect 8028 340 8059 352
rect 8065 340 8100 352
rect 7734 338 7896 340
rect 7629 310 7670 318
rect 7752 314 7765 338
rect 7780 336 7795 338
rect 7592 300 7593 310
rect 7608 300 7621 310
rect 7635 300 7636 310
rect 7651 300 7664 310
rect 7679 300 7709 314
rect 7752 300 7795 314
rect 7819 311 7826 318
rect 7829 314 7896 338
rect 7928 338 8100 340
rect 7898 316 7926 320
rect 7928 316 8008 338
rect 8029 336 8044 338
rect 7898 314 8008 316
rect 7829 310 8008 314
rect 7802 300 7832 310
rect 7834 300 7987 310
rect 7995 300 8025 310
rect 8029 300 8059 314
rect 8087 300 8100 338
rect 8172 344 8207 352
rect 8172 318 8173 344
rect 8180 318 8207 344
rect 8115 300 8145 314
rect 8172 310 8207 318
rect 8209 344 8250 352
rect 8209 318 8224 344
rect 8231 318 8250 344
rect 8314 340 8376 352
rect 8388 340 8463 352
rect 8521 340 8596 352
rect 8608 340 8639 352
rect 8645 340 8680 352
rect 8314 338 8476 340
rect 8209 310 8250 318
rect 8332 314 8345 338
rect 8360 336 8375 338
rect 8172 300 8173 310
rect 8188 300 8201 310
rect 8215 300 8216 310
rect 8231 300 8244 310
rect 8259 300 8289 314
rect 8332 300 8375 314
rect 8399 311 8406 318
rect 8409 314 8476 338
rect 8508 338 8680 340
rect 8478 316 8506 320
rect 8508 316 8588 338
rect 8609 336 8624 338
rect 8478 314 8588 316
rect 8409 310 8588 314
rect 8382 300 8412 310
rect 8414 300 8567 310
rect 8575 300 8605 310
rect 8609 300 8639 314
rect 8667 300 8680 338
rect 8752 344 8787 352
rect 8752 318 8753 344
rect 8760 318 8787 344
rect 8695 300 8725 314
rect 8752 310 8787 318
rect 8789 344 8830 352
rect 8789 318 8804 344
rect 8811 318 8830 344
rect 8894 340 8956 352
rect 8968 340 9043 352
rect 9101 340 9176 352
rect 9188 340 9219 352
rect 9225 340 9260 352
rect 8894 338 9056 340
rect 8789 310 8830 318
rect 8912 314 8925 338
rect 8940 336 8955 338
rect 8752 300 8753 310
rect 8768 300 8781 310
rect 8795 300 8796 310
rect 8811 300 8824 310
rect 8839 300 8869 314
rect 8912 300 8955 314
rect 8979 311 8986 318
rect 8989 314 9056 338
rect 9088 338 9260 340
rect 9058 316 9086 320
rect 9088 316 9168 338
rect 9189 336 9204 338
rect 9058 314 9168 316
rect 8989 310 9168 314
rect 8962 300 8992 310
rect 8994 300 9147 310
rect 9155 300 9185 310
rect 9189 300 9219 314
rect 9247 300 9260 338
rect 9332 344 9367 352
rect 9332 318 9333 344
rect 9340 318 9367 344
rect 9275 300 9305 314
rect 9332 310 9367 318
rect 9332 300 9333 310
rect 9348 300 9361 310
rect 5889 286 9361 300
rect 13 256 26 286
rect 41 268 71 286
rect 114 272 128 286
rect 164 272 384 286
rect 115 270 128 272
rect 81 258 96 270
rect 78 256 100 258
rect 105 256 135 270
rect 196 268 349 272
rect 178 256 370 268
rect 413 256 443 270
rect 449 256 462 286
rect 477 268 507 286
rect 550 256 563 286
rect 593 256 606 286
rect 621 268 651 286
rect 694 272 708 286
rect 744 272 964 286
rect 695 270 708 272
rect 661 258 676 270
rect 658 256 680 258
rect 685 256 715 270
rect 776 268 929 272
rect 758 256 950 268
rect 993 256 1023 270
rect 1029 256 1042 286
rect 1057 268 1087 286
rect 1130 256 1143 286
rect 1173 256 1186 286
rect 1201 268 1231 286
rect 1274 272 1288 286
rect 1324 272 1544 286
rect 1275 270 1288 272
rect 1241 258 1256 270
rect 1238 256 1260 258
rect 1265 256 1295 270
rect 1356 268 1509 272
rect 1338 256 1530 268
rect 1573 256 1603 270
rect 1609 256 1622 286
rect 1637 268 1667 286
rect 1710 256 1723 286
rect 1753 256 1766 286
rect 1781 268 1811 286
rect 1854 272 1868 286
rect 1904 272 2124 286
rect 1855 270 1868 272
rect 1821 258 1836 270
rect 1818 256 1840 258
rect 1845 256 1875 270
rect 1936 268 2089 272
rect 1918 256 2110 268
rect 2153 256 2183 270
rect 2189 256 2202 286
rect 2217 268 2247 286
rect 2290 256 2303 286
rect 2333 256 2346 286
rect 2361 268 2391 286
rect 2434 272 2448 286
rect 2484 272 2704 286
rect 2435 270 2448 272
rect 2401 258 2416 270
rect 2398 256 2420 258
rect 2425 256 2455 270
rect 2516 268 2669 272
rect 2498 256 2690 268
rect 2733 256 2763 270
rect 2769 256 2782 286
rect 2797 268 2827 286
rect 2870 256 2883 286
rect 2913 256 2926 286
rect 2941 268 2971 286
rect 3014 272 3028 286
rect 3064 272 3284 286
rect 3015 270 3028 272
rect 2981 258 2996 270
rect 2978 256 3000 258
rect 3005 256 3035 270
rect 3096 268 3249 272
rect 3078 256 3270 268
rect 3313 256 3343 270
rect 3349 256 3362 286
rect 3377 268 3407 286
rect 3450 256 3463 286
rect 5911 256 5924 286
rect 5939 268 5969 286
rect 6012 272 6026 286
rect 6062 272 6282 286
rect 6013 270 6026 272
rect 5979 258 5994 270
rect 5976 256 5998 258
rect 6003 256 6033 270
rect 6094 268 6247 272
rect 6076 256 6268 268
rect 6311 256 6341 270
rect 6347 256 6360 286
rect 6375 268 6405 286
rect 6448 256 6461 286
rect 6491 256 6504 286
rect 6519 268 6549 286
rect 6592 272 6606 286
rect 6642 272 6862 286
rect 6593 270 6606 272
rect 6559 258 6574 270
rect 6556 256 6578 258
rect 6583 256 6613 270
rect 6674 268 6827 272
rect 6656 256 6848 268
rect 6891 256 6921 270
rect 6927 256 6940 286
rect 6955 268 6985 286
rect 7028 256 7041 286
rect 7071 256 7084 286
rect 7099 268 7129 286
rect 7172 272 7186 286
rect 7222 272 7442 286
rect 7173 270 7186 272
rect 7139 258 7154 270
rect 7136 256 7158 258
rect 7163 256 7193 270
rect 7254 268 7407 272
rect 7236 256 7428 268
rect 7471 256 7501 270
rect 7507 256 7520 286
rect 7535 268 7565 286
rect 7608 256 7621 286
rect 7651 256 7664 286
rect 7679 268 7709 286
rect 7752 272 7766 286
rect 7802 272 8022 286
rect 7753 270 7766 272
rect 7719 258 7734 270
rect 7716 256 7738 258
rect 7743 256 7773 270
rect 7834 268 7987 272
rect 7816 256 8008 268
rect 8051 256 8081 270
rect 8087 256 8100 286
rect 8115 268 8145 286
rect 8188 256 8201 286
rect 8231 256 8244 286
rect 8259 268 8289 286
rect 8332 272 8346 286
rect 8382 272 8602 286
rect 8333 270 8346 272
rect 8299 258 8314 270
rect 8296 256 8318 258
rect 8323 256 8353 270
rect 8414 268 8567 272
rect 8396 256 8588 268
rect 8631 256 8661 270
rect 8667 256 8680 286
rect 8695 268 8725 286
rect 8768 256 8781 286
rect 8811 256 8824 286
rect 8839 268 8869 286
rect 8912 272 8926 286
rect 8962 272 9182 286
rect 8913 270 8926 272
rect 8879 258 8894 270
rect 8876 256 8898 258
rect 8903 256 8933 270
rect 8994 268 9147 272
rect 8976 256 9168 268
rect 9211 256 9241 270
rect 9247 256 9260 286
rect 9275 268 9305 286
rect 9348 256 9361 286
rect -2 242 3469 256
rect 5889 242 9361 256
rect 13 138 26 242
rect 71 220 72 230
rect 87 220 100 230
rect 71 216 100 220
rect 105 216 135 242
rect 153 228 169 230
rect 241 228 294 242
rect 242 226 306 228
rect 153 216 168 220
rect 71 214 168 216
rect 55 206 106 214
rect 55 194 80 206
rect 87 194 106 206
rect 137 206 187 214
rect 137 198 153 206
rect 160 204 187 206
rect 196 206 211 210
rect 258 206 290 226
rect 349 214 364 242
rect 413 239 443 242
rect 413 236 449 239
rect 379 228 395 230
rect 380 216 395 220
rect 413 217 452 236
rect 471 230 478 231
rect 477 223 478 230
rect 461 220 462 223
rect 477 220 490 223
rect 413 216 443 217
rect 452 216 458 217
rect 461 216 490 220
rect 380 215 490 216
rect 380 214 496 215
rect 349 206 417 214
rect 196 204 265 206
rect 283 204 417 206
rect 160 200 232 204
rect 160 198 285 200
rect 160 194 232 198
rect 55 186 106 194
rect 153 190 232 194
rect 313 190 417 204
rect 446 206 496 214
rect 446 197 462 206
rect 153 186 417 190
rect 443 194 462 197
rect 469 194 496 206
rect 443 186 496 194
rect 71 178 72 186
rect 87 178 100 186
rect 71 170 87 178
rect 68 163 87 166
rect 68 154 90 163
rect 41 144 90 154
rect 41 138 71 144
rect 90 139 95 144
rect 13 122 87 138
rect 105 130 135 186
rect 170 176 378 186
rect 413 182 458 186
rect 461 185 462 186
rect 477 185 490 186
rect 337 172 385 176
rect 220 150 250 159
rect 313 152 328 159
rect 349 150 385 172
rect 196 146 385 150
rect 211 143 385 146
rect 204 140 385 143
rect 13 120 26 122
rect 41 120 75 122
rect 13 104 87 120
rect 114 116 127 130
rect 142 116 158 132
rect 204 127 215 140
rect -3 82 -2 98
rect 13 82 26 104
rect 41 82 71 104
rect 114 100 176 116
rect 204 109 215 125
rect 220 120 230 140
rect 240 120 254 140
rect 257 127 266 140
rect 282 127 291 140
rect 220 109 254 120
rect 257 109 265 125
rect 282 109 291 125
rect 298 120 308 140
rect 318 120 332 140
rect 333 127 344 140
rect 298 109 332 120
rect 333 109 344 125
rect 390 116 406 132
rect 413 130 443 182
rect 477 178 478 185
rect 462 170 478 178
rect 449 138 462 157
rect 477 138 507 154
rect 449 122 523 138
rect 449 120 462 122
rect 477 120 511 122
rect 114 98 127 100
rect 142 98 176 100
rect 114 82 176 98
rect 220 93 233 96
rect 298 93 328 104
rect 376 100 422 116
rect 449 104 523 120
rect 376 98 410 100
rect 375 82 422 98
rect 449 82 462 104
rect 477 82 507 104
rect 534 82 535 98
rect 550 82 563 242
rect 593 138 606 242
rect 651 220 652 230
rect 667 220 680 230
rect 651 216 680 220
rect 685 216 715 242
rect 733 228 749 230
rect 821 228 874 242
rect 822 226 886 228
rect 733 216 748 220
rect 651 214 748 216
rect 635 206 686 214
rect 635 194 660 206
rect 667 194 686 206
rect 717 206 767 214
rect 717 198 733 206
rect 740 204 767 206
rect 776 206 791 210
rect 838 206 870 226
rect 929 214 944 242
rect 993 239 1023 242
rect 993 236 1029 239
rect 959 228 975 230
rect 960 216 975 220
rect 993 217 1032 236
rect 1051 230 1058 231
rect 1057 223 1058 230
rect 1041 220 1042 223
rect 1057 220 1070 223
rect 993 216 1023 217
rect 1032 216 1038 217
rect 1041 216 1070 220
rect 960 215 1070 216
rect 960 214 1076 215
rect 929 206 997 214
rect 776 204 845 206
rect 863 204 997 206
rect 740 200 812 204
rect 740 198 865 200
rect 740 194 812 198
rect 635 186 686 194
rect 733 190 812 194
rect 893 190 997 204
rect 1026 206 1076 214
rect 1026 197 1042 206
rect 733 186 997 190
rect 1023 194 1042 197
rect 1049 194 1076 206
rect 1023 186 1076 194
rect 651 178 652 186
rect 667 178 680 186
rect 651 170 667 178
rect 648 163 667 166
rect 648 154 670 163
rect 621 144 670 154
rect 621 138 651 144
rect 670 139 675 144
rect 593 122 667 138
rect 685 130 715 186
rect 750 176 958 186
rect 993 182 1038 186
rect 1041 185 1042 186
rect 1057 185 1070 186
rect 917 172 965 176
rect 800 150 830 159
rect 893 152 908 159
rect 929 150 965 172
rect 776 146 965 150
rect 791 143 965 146
rect 784 140 965 143
rect 593 120 606 122
rect 621 120 655 122
rect 593 104 667 120
rect 694 116 707 130
rect 722 116 738 132
rect 784 127 795 140
rect 577 82 578 98
rect 593 82 606 104
rect 621 82 651 104
rect 694 100 756 116
rect 784 109 795 125
rect 800 120 810 140
rect 820 120 834 140
rect 837 127 846 140
rect 862 127 871 140
rect 800 109 834 120
rect 837 109 845 125
rect 862 109 871 125
rect 878 120 888 140
rect 898 120 912 140
rect 913 127 924 140
rect 878 109 912 120
rect 913 109 924 125
rect 970 116 986 132
rect 993 130 1023 182
rect 1057 178 1058 185
rect 1042 170 1058 178
rect 1029 138 1042 157
rect 1057 138 1087 154
rect 1029 122 1103 138
rect 1029 120 1042 122
rect 1057 120 1091 122
rect 694 98 707 100
rect 722 98 756 100
rect 694 82 756 98
rect 800 93 813 96
rect 878 93 908 104
rect 956 100 1002 116
rect 1029 104 1103 120
rect 956 98 990 100
rect 955 82 1002 98
rect 1029 82 1042 104
rect 1057 82 1087 104
rect 1114 82 1115 98
rect 1130 82 1143 242
rect 1173 138 1186 242
rect 1231 220 1232 230
rect 1247 220 1260 230
rect 1231 216 1260 220
rect 1265 216 1295 242
rect 1313 228 1329 230
rect 1401 228 1454 242
rect 1402 226 1466 228
rect 1313 216 1328 220
rect 1231 214 1328 216
rect 1215 206 1266 214
rect 1215 194 1240 206
rect 1247 194 1266 206
rect 1297 206 1347 214
rect 1297 198 1313 206
rect 1320 204 1347 206
rect 1356 206 1371 210
rect 1418 206 1450 226
rect 1509 214 1524 242
rect 1573 239 1603 242
rect 1573 236 1609 239
rect 1539 228 1555 230
rect 1540 216 1555 220
rect 1573 217 1612 236
rect 1631 230 1638 231
rect 1637 223 1638 230
rect 1621 220 1622 223
rect 1637 220 1650 223
rect 1573 216 1603 217
rect 1612 216 1618 217
rect 1621 216 1650 220
rect 1540 215 1650 216
rect 1540 214 1656 215
rect 1509 206 1577 214
rect 1356 204 1425 206
rect 1443 204 1577 206
rect 1320 200 1392 204
rect 1320 198 1445 200
rect 1320 194 1392 198
rect 1215 186 1266 194
rect 1313 190 1392 194
rect 1473 190 1577 204
rect 1606 206 1656 214
rect 1606 197 1622 206
rect 1313 186 1577 190
rect 1603 194 1622 197
rect 1629 194 1656 206
rect 1603 186 1656 194
rect 1231 178 1232 186
rect 1247 178 1260 186
rect 1231 170 1247 178
rect 1228 163 1247 166
rect 1228 154 1250 163
rect 1201 144 1250 154
rect 1201 138 1231 144
rect 1250 139 1255 144
rect 1173 122 1247 138
rect 1265 130 1295 186
rect 1330 176 1538 186
rect 1573 182 1618 186
rect 1621 185 1622 186
rect 1637 185 1650 186
rect 1497 172 1545 176
rect 1380 150 1410 159
rect 1473 152 1488 159
rect 1509 150 1545 172
rect 1356 146 1545 150
rect 1371 143 1545 146
rect 1364 140 1545 143
rect 1173 120 1186 122
rect 1201 120 1235 122
rect 1173 104 1247 120
rect 1274 116 1287 130
rect 1302 116 1318 132
rect 1364 127 1375 140
rect 1157 82 1158 98
rect 1173 82 1186 104
rect 1201 82 1231 104
rect 1274 100 1336 116
rect 1364 109 1375 125
rect 1380 120 1390 140
rect 1400 120 1414 140
rect 1417 127 1426 140
rect 1442 127 1451 140
rect 1380 109 1414 120
rect 1417 109 1425 125
rect 1442 109 1451 125
rect 1458 120 1468 140
rect 1478 120 1492 140
rect 1493 127 1504 140
rect 1458 109 1492 120
rect 1493 109 1504 125
rect 1550 116 1566 132
rect 1573 130 1603 182
rect 1637 178 1638 185
rect 1622 170 1638 178
rect 1609 138 1622 157
rect 1637 138 1667 154
rect 1609 122 1683 138
rect 1609 120 1622 122
rect 1637 120 1671 122
rect 1274 98 1287 100
rect 1302 98 1336 100
rect 1274 82 1336 98
rect 1380 93 1393 96
rect 1458 93 1488 104
rect 1536 100 1582 116
rect 1609 104 1683 120
rect 1536 98 1570 100
rect 1535 82 1582 98
rect 1609 82 1622 104
rect 1637 82 1667 104
rect 1694 82 1695 98
rect 1710 82 1723 242
rect 1753 138 1766 242
rect 1811 220 1812 230
rect 1827 220 1840 230
rect 1811 216 1840 220
rect 1845 216 1875 242
rect 1893 228 1909 230
rect 1981 228 2034 242
rect 1982 226 2046 228
rect 1893 216 1908 220
rect 1811 214 1908 216
rect 1795 206 1846 214
rect 1795 194 1820 206
rect 1827 194 1846 206
rect 1877 206 1927 214
rect 1877 198 1893 206
rect 1900 204 1927 206
rect 1936 206 1951 210
rect 1998 206 2030 226
rect 2089 214 2104 242
rect 2153 239 2183 242
rect 2153 236 2189 239
rect 2119 228 2135 230
rect 2120 216 2135 220
rect 2153 217 2192 236
rect 2211 230 2218 231
rect 2217 223 2218 230
rect 2201 220 2202 223
rect 2217 220 2230 223
rect 2153 216 2183 217
rect 2192 216 2198 217
rect 2201 216 2230 220
rect 2120 215 2230 216
rect 2120 214 2236 215
rect 2089 206 2157 214
rect 1936 204 2005 206
rect 2023 204 2157 206
rect 1900 200 1972 204
rect 1900 198 2025 200
rect 1900 194 1972 198
rect 1795 186 1846 194
rect 1893 190 1972 194
rect 2053 190 2157 204
rect 2186 206 2236 214
rect 2186 197 2202 206
rect 1893 186 2157 190
rect 2183 194 2202 197
rect 2209 194 2236 206
rect 2183 186 2236 194
rect 1811 178 1812 186
rect 1827 178 1840 186
rect 1811 170 1827 178
rect 1808 163 1827 166
rect 1808 154 1830 163
rect 1781 144 1830 154
rect 1781 138 1811 144
rect 1830 139 1835 144
rect 1753 122 1827 138
rect 1845 130 1875 186
rect 1910 176 2118 186
rect 2153 182 2198 186
rect 2201 185 2202 186
rect 2217 185 2230 186
rect 2077 172 2125 176
rect 1960 150 1990 159
rect 2053 152 2068 159
rect 2089 150 2125 172
rect 1936 146 2125 150
rect 1951 143 2125 146
rect 1944 140 2125 143
rect 1753 120 1766 122
rect 1781 120 1815 122
rect 1753 104 1827 120
rect 1854 116 1867 130
rect 1882 116 1898 132
rect 1944 127 1955 140
rect 1737 82 1738 98
rect 1753 82 1766 104
rect 1781 82 1811 104
rect 1854 100 1916 116
rect 1944 109 1955 125
rect 1960 120 1970 140
rect 1980 120 1994 140
rect 1997 127 2006 140
rect 2022 127 2031 140
rect 1960 109 1994 120
rect 1997 109 2005 125
rect 2022 109 2031 125
rect 2038 120 2048 140
rect 2058 120 2072 140
rect 2073 127 2084 140
rect 2038 109 2072 120
rect 2073 109 2084 125
rect 2130 116 2146 132
rect 2153 130 2183 182
rect 2217 178 2218 185
rect 2202 170 2218 178
rect 2189 138 2202 157
rect 2217 138 2247 154
rect 2189 122 2263 138
rect 2189 120 2202 122
rect 2217 120 2251 122
rect 1854 98 1867 100
rect 1882 98 1916 100
rect 1854 82 1916 98
rect 1960 93 1973 96
rect 2038 93 2068 104
rect 2116 100 2162 116
rect 2189 104 2263 120
rect 2116 98 2150 100
rect 2115 82 2162 98
rect 2189 82 2202 104
rect 2217 82 2247 104
rect 2274 82 2275 98
rect 2290 82 2303 242
rect 2333 138 2346 242
rect 2391 220 2392 230
rect 2407 220 2420 230
rect 2391 216 2420 220
rect 2425 216 2455 242
rect 2473 228 2489 230
rect 2561 228 2614 242
rect 2562 226 2626 228
rect 2473 216 2488 220
rect 2391 214 2488 216
rect 2375 206 2426 214
rect 2375 194 2400 206
rect 2407 194 2426 206
rect 2457 206 2507 214
rect 2457 198 2473 206
rect 2480 204 2507 206
rect 2516 206 2531 210
rect 2578 206 2610 226
rect 2669 214 2684 242
rect 2733 239 2763 242
rect 2733 236 2769 239
rect 2699 228 2715 230
rect 2700 216 2715 220
rect 2733 217 2772 236
rect 2791 230 2798 231
rect 2797 223 2798 230
rect 2781 220 2782 223
rect 2797 220 2810 223
rect 2733 216 2763 217
rect 2772 216 2778 217
rect 2781 216 2810 220
rect 2700 215 2810 216
rect 2700 214 2816 215
rect 2669 206 2737 214
rect 2516 204 2585 206
rect 2603 204 2737 206
rect 2480 200 2552 204
rect 2480 198 2605 200
rect 2480 194 2552 198
rect 2375 186 2426 194
rect 2473 190 2552 194
rect 2633 190 2737 204
rect 2766 206 2816 214
rect 2766 197 2782 206
rect 2473 186 2737 190
rect 2763 194 2782 197
rect 2789 194 2816 206
rect 2763 186 2816 194
rect 2391 178 2392 186
rect 2407 178 2420 186
rect 2391 170 2407 178
rect 2388 163 2407 166
rect 2388 154 2410 163
rect 2361 144 2410 154
rect 2361 138 2391 144
rect 2410 139 2415 144
rect 2333 122 2407 138
rect 2425 130 2455 186
rect 2490 176 2698 186
rect 2733 182 2778 186
rect 2781 185 2782 186
rect 2797 185 2810 186
rect 2657 172 2705 176
rect 2540 150 2570 159
rect 2633 152 2648 159
rect 2669 150 2705 172
rect 2516 146 2705 150
rect 2531 143 2705 146
rect 2524 140 2705 143
rect 2333 120 2346 122
rect 2361 120 2395 122
rect 2333 104 2407 120
rect 2434 116 2447 130
rect 2462 116 2478 132
rect 2524 127 2535 140
rect 2317 82 2318 98
rect 2333 82 2346 104
rect 2361 82 2391 104
rect 2434 100 2496 116
rect 2524 109 2535 125
rect 2540 120 2550 140
rect 2560 120 2574 140
rect 2577 127 2586 140
rect 2602 127 2611 140
rect 2540 109 2574 120
rect 2577 109 2585 125
rect 2602 109 2611 125
rect 2618 120 2628 140
rect 2638 120 2652 140
rect 2653 127 2664 140
rect 2618 109 2652 120
rect 2653 109 2664 125
rect 2710 116 2726 132
rect 2733 130 2763 182
rect 2797 178 2798 185
rect 2782 170 2798 178
rect 2769 138 2782 157
rect 2797 138 2827 154
rect 2769 122 2843 138
rect 2769 120 2782 122
rect 2797 120 2831 122
rect 2434 98 2447 100
rect 2462 98 2496 100
rect 2434 82 2496 98
rect 2540 93 2553 96
rect 2618 93 2648 104
rect 2696 100 2742 116
rect 2769 104 2843 120
rect 2696 98 2730 100
rect 2695 82 2742 98
rect 2769 82 2782 104
rect 2797 82 2827 104
rect 2854 82 2855 98
rect 2870 82 2883 242
rect 2913 138 2926 242
rect 2971 220 2972 230
rect 2987 220 3000 230
rect 2971 216 3000 220
rect 3005 216 3035 242
rect 3053 228 3069 230
rect 3141 228 3194 242
rect 3142 226 3206 228
rect 3053 216 3068 220
rect 2971 214 3068 216
rect 2955 206 3006 214
rect 2955 194 2980 206
rect 2987 194 3006 206
rect 3037 206 3087 214
rect 3037 198 3053 206
rect 3060 204 3087 206
rect 3096 206 3111 210
rect 3158 206 3190 226
rect 3249 214 3264 242
rect 3313 239 3343 242
rect 3313 236 3349 239
rect 3279 228 3295 230
rect 3280 216 3295 220
rect 3313 217 3352 236
rect 3371 230 3378 231
rect 3377 223 3378 230
rect 3361 220 3362 223
rect 3377 220 3390 223
rect 3313 216 3343 217
rect 3352 216 3358 217
rect 3361 216 3390 220
rect 3280 215 3390 216
rect 3280 214 3396 215
rect 3249 206 3317 214
rect 3096 204 3165 206
rect 3183 204 3317 206
rect 3060 200 3132 204
rect 3060 198 3185 200
rect 3060 194 3132 198
rect 2955 186 3006 194
rect 3053 190 3132 194
rect 3213 190 3317 204
rect 3346 206 3396 214
rect 3346 197 3362 206
rect 3053 186 3317 190
rect 3343 194 3362 197
rect 3369 194 3396 206
rect 3343 186 3396 194
rect 2971 178 2972 186
rect 2987 178 3000 186
rect 2971 170 2987 178
rect 2968 163 2987 166
rect 2968 154 2990 163
rect 2941 144 2990 154
rect 2941 138 2971 144
rect 2990 139 2995 144
rect 2913 122 2987 138
rect 3005 130 3035 186
rect 3070 176 3278 186
rect 3313 182 3358 186
rect 3361 185 3362 186
rect 3377 185 3390 186
rect 3237 172 3285 176
rect 3120 150 3150 159
rect 3213 152 3228 159
rect 3249 150 3285 172
rect 3096 146 3285 150
rect 3111 143 3285 146
rect 3104 140 3285 143
rect 2913 120 2926 122
rect 2941 120 2975 122
rect 2913 104 2987 120
rect 3014 116 3027 130
rect 3042 116 3058 132
rect 3104 127 3115 140
rect 2897 82 2898 98
rect 2913 82 2926 104
rect 2941 82 2971 104
rect 3014 100 3076 116
rect 3104 109 3115 125
rect 3120 120 3130 140
rect 3140 120 3154 140
rect 3157 127 3166 140
rect 3182 127 3191 140
rect 3120 109 3154 120
rect 3157 109 3165 125
rect 3182 109 3191 125
rect 3198 120 3208 140
rect 3218 120 3232 140
rect 3233 127 3244 140
rect 3198 109 3232 120
rect 3233 109 3244 125
rect 3290 116 3306 132
rect 3313 130 3343 182
rect 3377 178 3378 185
rect 3362 170 3378 178
rect 3349 138 3362 157
rect 3377 138 3407 154
rect 3349 122 3423 138
rect 3349 120 3362 122
rect 3377 120 3411 122
rect 3014 98 3027 100
rect 3042 98 3076 100
rect 3014 82 3076 98
rect 3120 93 3133 96
rect 3198 93 3228 104
rect 3276 100 3322 116
rect 3349 104 3423 120
rect 3276 98 3310 100
rect 3275 82 3322 98
rect 3349 82 3362 104
rect 3377 82 3407 104
rect 3434 82 3435 98
rect 3450 82 3463 242
rect 5911 138 5924 242
rect 5969 220 5970 230
rect 5985 220 5998 230
rect 5969 216 5998 220
rect 6003 216 6033 242
rect 6051 228 6067 230
rect 6139 228 6192 242
rect 6140 226 6204 228
rect 6051 216 6066 220
rect 5969 214 6066 216
rect 5953 206 6004 214
rect 5953 194 5978 206
rect 5985 194 6004 206
rect 6035 206 6085 214
rect 6035 198 6051 206
rect 6058 204 6085 206
rect 6094 206 6109 210
rect 6156 206 6188 226
rect 6247 214 6262 242
rect 6311 239 6341 242
rect 6311 236 6347 239
rect 6277 228 6293 230
rect 6278 216 6293 220
rect 6311 217 6350 236
rect 6369 230 6376 231
rect 6375 223 6376 230
rect 6359 220 6360 223
rect 6375 220 6388 223
rect 6311 216 6341 217
rect 6350 216 6356 217
rect 6359 216 6388 220
rect 6278 215 6388 216
rect 6278 214 6394 215
rect 6247 206 6315 214
rect 6094 204 6163 206
rect 6181 204 6315 206
rect 6058 200 6130 204
rect 6058 198 6183 200
rect 6058 194 6130 198
rect 5953 186 6004 194
rect 6051 190 6130 194
rect 6211 190 6315 204
rect 6344 206 6394 214
rect 6344 197 6360 206
rect 6051 186 6315 190
rect 6341 194 6360 197
rect 6367 194 6394 206
rect 6341 186 6394 194
rect 5969 178 5970 186
rect 5985 178 5998 186
rect 5969 170 5985 178
rect 5966 163 5985 166
rect 5966 154 5988 163
rect 5939 144 5988 154
rect 5939 138 5969 144
rect 5988 139 5993 144
rect 5911 122 5985 138
rect 6003 130 6033 186
rect 6068 176 6276 186
rect 6311 182 6356 186
rect 6359 185 6360 186
rect 6375 185 6388 186
rect 6235 172 6283 176
rect 6118 150 6148 159
rect 6211 152 6226 159
rect 6247 150 6283 172
rect 6094 146 6283 150
rect 6109 143 6283 146
rect 6102 140 6283 143
rect 5911 120 5924 122
rect 5939 120 5973 122
rect 5911 104 5985 120
rect 6012 116 6025 130
rect 6040 116 6056 132
rect 6102 127 6113 140
rect 5895 82 5896 98
rect 5911 82 5924 104
rect 5939 82 5969 104
rect 6012 100 6074 116
rect 6102 109 6113 125
rect 6118 120 6128 140
rect 6138 120 6152 140
rect 6155 127 6164 140
rect 6180 127 6189 140
rect 6118 109 6152 120
rect 6155 109 6163 125
rect 6180 109 6189 125
rect 6196 120 6206 140
rect 6216 120 6230 140
rect 6231 127 6242 140
rect 6196 109 6230 120
rect 6231 109 6242 125
rect 6288 116 6304 132
rect 6311 130 6341 182
rect 6375 178 6376 185
rect 6360 170 6376 178
rect 6347 138 6360 157
rect 6375 138 6405 154
rect 6347 122 6421 138
rect 6347 120 6360 122
rect 6375 120 6409 122
rect 6012 98 6025 100
rect 6040 98 6074 100
rect 6012 82 6074 98
rect 6118 93 6131 96
rect 6196 93 6226 104
rect 6274 100 6320 116
rect 6347 104 6421 120
rect 6274 98 6308 100
rect 6273 82 6320 98
rect 6347 82 6360 104
rect 6375 82 6405 104
rect 6432 82 6433 98
rect 6448 82 6461 242
rect 6491 138 6504 242
rect 6549 220 6550 230
rect 6565 220 6578 230
rect 6549 216 6578 220
rect 6583 216 6613 242
rect 6631 228 6647 230
rect 6719 228 6772 242
rect 6720 226 6784 228
rect 6631 216 6646 220
rect 6549 214 6646 216
rect 6533 206 6584 214
rect 6533 194 6558 206
rect 6565 194 6584 206
rect 6615 206 6665 214
rect 6615 198 6631 206
rect 6638 204 6665 206
rect 6674 206 6689 210
rect 6736 206 6768 226
rect 6827 214 6842 242
rect 6891 239 6921 242
rect 6891 236 6927 239
rect 6857 228 6873 230
rect 6858 216 6873 220
rect 6891 217 6930 236
rect 6949 230 6956 231
rect 6955 223 6956 230
rect 6939 220 6940 223
rect 6955 220 6968 223
rect 6891 216 6921 217
rect 6930 216 6936 217
rect 6939 216 6968 220
rect 6858 215 6968 216
rect 6858 214 6974 215
rect 6827 206 6895 214
rect 6674 204 6743 206
rect 6761 204 6895 206
rect 6638 200 6710 204
rect 6638 198 6763 200
rect 6638 194 6710 198
rect 6533 186 6584 194
rect 6631 190 6710 194
rect 6791 190 6895 204
rect 6924 206 6974 214
rect 6924 197 6940 206
rect 6631 186 6895 190
rect 6921 194 6940 197
rect 6947 194 6974 206
rect 6921 186 6974 194
rect 6549 178 6550 186
rect 6565 178 6578 186
rect 6549 170 6565 178
rect 6546 163 6565 166
rect 6546 154 6568 163
rect 6519 144 6568 154
rect 6519 138 6549 144
rect 6568 139 6573 144
rect 6491 122 6565 138
rect 6583 130 6613 186
rect 6648 176 6856 186
rect 6891 182 6936 186
rect 6939 185 6940 186
rect 6955 185 6968 186
rect 6815 172 6863 176
rect 6698 150 6728 159
rect 6791 152 6806 159
rect 6827 150 6863 172
rect 6674 146 6863 150
rect 6689 143 6863 146
rect 6682 140 6863 143
rect 6491 120 6504 122
rect 6519 120 6553 122
rect 6491 104 6565 120
rect 6592 116 6605 130
rect 6620 116 6636 132
rect 6682 127 6693 140
rect 6475 82 6476 98
rect 6491 82 6504 104
rect 6519 82 6549 104
rect 6592 100 6654 116
rect 6682 109 6693 125
rect 6698 120 6708 140
rect 6718 120 6732 140
rect 6735 127 6744 140
rect 6760 127 6769 140
rect 6698 109 6732 120
rect 6735 109 6743 125
rect 6760 109 6769 125
rect 6776 120 6786 140
rect 6796 120 6810 140
rect 6811 127 6822 140
rect 6776 109 6810 120
rect 6811 109 6822 125
rect 6868 116 6884 132
rect 6891 130 6921 182
rect 6955 178 6956 185
rect 6940 170 6956 178
rect 6927 138 6940 157
rect 6955 138 6985 154
rect 6927 122 7001 138
rect 6927 120 6940 122
rect 6955 120 6989 122
rect 6592 98 6605 100
rect 6620 98 6654 100
rect 6592 82 6654 98
rect 6698 93 6711 96
rect 6776 93 6806 104
rect 6854 100 6900 116
rect 6927 104 7001 120
rect 6854 98 6888 100
rect 6853 82 6900 98
rect 6927 82 6940 104
rect 6955 82 6985 104
rect 7012 82 7013 98
rect 7028 82 7041 242
rect 7071 138 7084 242
rect 7129 220 7130 230
rect 7145 220 7158 230
rect 7129 216 7158 220
rect 7163 216 7193 242
rect 7211 228 7227 230
rect 7299 228 7352 242
rect 7300 226 7364 228
rect 7211 216 7226 220
rect 7129 214 7226 216
rect 7113 206 7164 214
rect 7113 194 7138 206
rect 7145 194 7164 206
rect 7195 206 7245 214
rect 7195 198 7211 206
rect 7218 204 7245 206
rect 7254 206 7269 210
rect 7316 206 7348 226
rect 7407 214 7422 242
rect 7471 239 7501 242
rect 7471 236 7507 239
rect 7437 228 7453 230
rect 7438 216 7453 220
rect 7471 217 7510 236
rect 7529 230 7536 231
rect 7535 223 7536 230
rect 7519 220 7520 223
rect 7535 220 7548 223
rect 7471 216 7501 217
rect 7510 216 7516 217
rect 7519 216 7548 220
rect 7438 215 7548 216
rect 7438 214 7554 215
rect 7407 206 7475 214
rect 7254 204 7323 206
rect 7341 204 7475 206
rect 7218 200 7290 204
rect 7218 198 7343 200
rect 7218 194 7290 198
rect 7113 186 7164 194
rect 7211 190 7290 194
rect 7371 190 7475 204
rect 7504 206 7554 214
rect 7504 197 7520 206
rect 7211 186 7475 190
rect 7501 194 7520 197
rect 7527 194 7554 206
rect 7501 186 7554 194
rect 7129 178 7130 186
rect 7145 178 7158 186
rect 7129 170 7145 178
rect 7126 163 7145 166
rect 7126 154 7148 163
rect 7099 144 7148 154
rect 7099 138 7129 144
rect 7148 139 7153 144
rect 7071 122 7145 138
rect 7163 130 7193 186
rect 7228 176 7436 186
rect 7471 182 7516 186
rect 7519 185 7520 186
rect 7535 185 7548 186
rect 7395 172 7443 176
rect 7278 150 7308 159
rect 7371 152 7386 159
rect 7407 150 7443 172
rect 7254 146 7443 150
rect 7269 143 7443 146
rect 7262 140 7443 143
rect 7071 120 7084 122
rect 7099 120 7133 122
rect 7071 104 7145 120
rect 7172 116 7185 130
rect 7200 116 7216 132
rect 7262 127 7273 140
rect 7055 82 7056 98
rect 7071 82 7084 104
rect 7099 82 7129 104
rect 7172 100 7234 116
rect 7262 109 7273 125
rect 7278 120 7288 140
rect 7298 120 7312 140
rect 7315 127 7324 140
rect 7340 127 7349 140
rect 7278 109 7312 120
rect 7315 109 7323 125
rect 7340 109 7349 125
rect 7356 120 7366 140
rect 7376 120 7390 140
rect 7391 127 7402 140
rect 7356 109 7390 120
rect 7391 109 7402 125
rect 7448 116 7464 132
rect 7471 130 7501 182
rect 7535 178 7536 185
rect 7520 170 7536 178
rect 7507 138 7520 157
rect 7535 138 7565 154
rect 7507 122 7581 138
rect 7507 120 7520 122
rect 7535 120 7569 122
rect 7172 98 7185 100
rect 7200 98 7234 100
rect 7172 82 7234 98
rect 7278 93 7291 96
rect 7356 93 7386 104
rect 7434 100 7480 116
rect 7507 104 7581 120
rect 7434 98 7468 100
rect 7433 82 7480 98
rect 7507 82 7520 104
rect 7535 82 7565 104
rect 7592 82 7593 98
rect 7608 82 7621 242
rect 7651 138 7664 242
rect 7709 220 7710 230
rect 7725 220 7738 230
rect 7709 216 7738 220
rect 7743 216 7773 242
rect 7791 228 7807 230
rect 7879 228 7932 242
rect 7880 226 7944 228
rect 7791 216 7806 220
rect 7709 214 7806 216
rect 7693 206 7744 214
rect 7693 194 7718 206
rect 7725 194 7744 206
rect 7775 206 7825 214
rect 7775 198 7791 206
rect 7798 204 7825 206
rect 7834 206 7849 210
rect 7896 206 7928 226
rect 7987 214 8002 242
rect 8051 239 8081 242
rect 8051 236 8087 239
rect 8017 228 8033 230
rect 8018 216 8033 220
rect 8051 217 8090 236
rect 8109 230 8116 231
rect 8115 223 8116 230
rect 8099 220 8100 223
rect 8115 220 8128 223
rect 8051 216 8081 217
rect 8090 216 8096 217
rect 8099 216 8128 220
rect 8018 215 8128 216
rect 8018 214 8134 215
rect 7987 206 8055 214
rect 7834 204 7903 206
rect 7921 204 8055 206
rect 7798 200 7870 204
rect 7798 198 7923 200
rect 7798 194 7870 198
rect 7693 186 7744 194
rect 7791 190 7870 194
rect 7951 190 8055 204
rect 8084 206 8134 214
rect 8084 197 8100 206
rect 7791 186 8055 190
rect 8081 194 8100 197
rect 8107 194 8134 206
rect 8081 186 8134 194
rect 7709 178 7710 186
rect 7725 178 7738 186
rect 7709 170 7725 178
rect 7706 163 7725 166
rect 7706 154 7728 163
rect 7679 144 7728 154
rect 7679 138 7709 144
rect 7728 139 7733 144
rect 7651 122 7725 138
rect 7743 130 7773 186
rect 7808 176 8016 186
rect 8051 182 8096 186
rect 8099 185 8100 186
rect 8115 185 8128 186
rect 7975 172 8023 176
rect 7858 150 7888 159
rect 7951 152 7966 159
rect 7987 150 8023 172
rect 7834 146 8023 150
rect 7849 143 8023 146
rect 7842 140 8023 143
rect 7651 120 7664 122
rect 7679 120 7713 122
rect 7651 104 7725 120
rect 7752 116 7765 130
rect 7780 116 7796 132
rect 7842 127 7853 140
rect 7635 82 7636 98
rect 7651 82 7664 104
rect 7679 82 7709 104
rect 7752 100 7814 116
rect 7842 109 7853 125
rect 7858 120 7868 140
rect 7878 120 7892 140
rect 7895 127 7904 140
rect 7920 127 7929 140
rect 7858 109 7892 120
rect 7895 109 7903 125
rect 7920 109 7929 125
rect 7936 120 7946 140
rect 7956 120 7970 140
rect 7971 127 7982 140
rect 7936 109 7970 120
rect 7971 109 7982 125
rect 8028 116 8044 132
rect 8051 130 8081 182
rect 8115 178 8116 185
rect 8100 170 8116 178
rect 8087 138 8100 157
rect 8115 138 8145 154
rect 8087 122 8161 138
rect 8087 120 8100 122
rect 8115 120 8149 122
rect 7752 98 7765 100
rect 7780 98 7814 100
rect 7752 82 7814 98
rect 7858 93 7871 96
rect 7936 93 7966 104
rect 8014 100 8060 116
rect 8087 104 8161 120
rect 8014 98 8048 100
rect 8013 82 8060 98
rect 8087 82 8100 104
rect 8115 82 8145 104
rect 8172 82 8173 98
rect 8188 82 8201 242
rect 8231 138 8244 242
rect 8289 220 8290 230
rect 8305 220 8318 230
rect 8289 216 8318 220
rect 8323 216 8353 242
rect 8371 228 8387 230
rect 8459 228 8512 242
rect 8460 226 8524 228
rect 8371 216 8386 220
rect 8289 214 8386 216
rect 8273 206 8324 214
rect 8273 194 8298 206
rect 8305 194 8324 206
rect 8355 206 8405 214
rect 8355 198 8371 206
rect 8378 204 8405 206
rect 8414 206 8429 210
rect 8476 206 8508 226
rect 8567 214 8582 242
rect 8631 239 8661 242
rect 8631 236 8667 239
rect 8597 228 8613 230
rect 8598 216 8613 220
rect 8631 217 8670 236
rect 8689 230 8696 231
rect 8695 223 8696 230
rect 8679 220 8680 223
rect 8695 220 8708 223
rect 8631 216 8661 217
rect 8670 216 8676 217
rect 8679 216 8708 220
rect 8598 215 8708 216
rect 8598 214 8714 215
rect 8567 206 8635 214
rect 8414 204 8483 206
rect 8501 204 8635 206
rect 8378 200 8450 204
rect 8378 198 8503 200
rect 8378 194 8450 198
rect 8273 186 8324 194
rect 8371 190 8450 194
rect 8531 190 8635 204
rect 8664 206 8714 214
rect 8664 197 8680 206
rect 8371 186 8635 190
rect 8661 194 8680 197
rect 8687 194 8714 206
rect 8661 186 8714 194
rect 8289 178 8290 186
rect 8305 178 8318 186
rect 8289 170 8305 178
rect 8286 163 8305 166
rect 8286 154 8308 163
rect 8259 144 8308 154
rect 8259 138 8289 144
rect 8308 139 8313 144
rect 8231 122 8305 138
rect 8323 130 8353 186
rect 8388 176 8596 186
rect 8631 182 8676 186
rect 8679 185 8680 186
rect 8695 185 8708 186
rect 8555 172 8603 176
rect 8438 150 8468 159
rect 8531 152 8546 159
rect 8567 150 8603 172
rect 8414 146 8603 150
rect 8429 143 8603 146
rect 8422 140 8603 143
rect 8231 120 8244 122
rect 8259 120 8293 122
rect 8231 104 8305 120
rect 8332 116 8345 130
rect 8360 116 8376 132
rect 8422 127 8433 140
rect 8215 82 8216 98
rect 8231 82 8244 104
rect 8259 82 8289 104
rect 8332 100 8394 116
rect 8422 109 8433 125
rect 8438 120 8448 140
rect 8458 120 8472 140
rect 8475 127 8484 140
rect 8500 127 8509 140
rect 8438 109 8472 120
rect 8475 109 8483 125
rect 8500 109 8509 125
rect 8516 120 8526 140
rect 8536 120 8550 140
rect 8551 127 8562 140
rect 8516 109 8550 120
rect 8551 109 8562 125
rect 8608 116 8624 132
rect 8631 130 8661 182
rect 8695 178 8696 185
rect 8680 170 8696 178
rect 8667 138 8680 157
rect 8695 138 8725 154
rect 8667 122 8741 138
rect 8667 120 8680 122
rect 8695 120 8729 122
rect 8332 98 8345 100
rect 8360 98 8394 100
rect 8332 82 8394 98
rect 8438 93 8451 96
rect 8516 93 8546 104
rect 8594 100 8640 116
rect 8667 104 8741 120
rect 8594 98 8628 100
rect 8593 82 8640 98
rect 8667 82 8680 104
rect 8695 82 8725 104
rect 8752 82 8753 98
rect 8768 82 8781 242
rect 8811 138 8824 242
rect 8869 220 8870 230
rect 8885 220 8898 230
rect 8869 216 8898 220
rect 8903 216 8933 242
rect 8951 228 8967 230
rect 9039 228 9092 242
rect 9040 226 9104 228
rect 8951 216 8966 220
rect 8869 214 8966 216
rect 8853 206 8904 214
rect 8853 194 8878 206
rect 8885 194 8904 206
rect 8935 206 8985 214
rect 8935 198 8951 206
rect 8958 204 8985 206
rect 8994 206 9009 210
rect 9056 206 9088 226
rect 9147 214 9162 242
rect 9211 239 9241 242
rect 9211 236 9247 239
rect 9177 228 9193 230
rect 9178 216 9193 220
rect 9211 217 9250 236
rect 9269 230 9276 231
rect 9275 223 9276 230
rect 9259 220 9260 223
rect 9275 220 9288 223
rect 9211 216 9241 217
rect 9250 216 9256 217
rect 9259 216 9288 220
rect 9178 215 9288 216
rect 9178 214 9294 215
rect 9147 206 9215 214
rect 8994 204 9063 206
rect 9081 204 9215 206
rect 8958 200 9030 204
rect 8958 198 9083 200
rect 8958 194 9030 198
rect 8853 186 8904 194
rect 8951 190 9030 194
rect 9111 190 9215 204
rect 9244 206 9294 214
rect 9244 197 9260 206
rect 8951 186 9215 190
rect 9241 194 9260 197
rect 9267 194 9294 206
rect 9241 186 9294 194
rect 8869 178 8870 186
rect 8885 178 8898 186
rect 8869 170 8885 178
rect 8866 163 8885 166
rect 8866 154 8888 163
rect 8839 144 8888 154
rect 8839 138 8869 144
rect 8888 139 8893 144
rect 8811 122 8885 138
rect 8903 130 8933 186
rect 8968 176 9176 186
rect 9211 182 9256 186
rect 9259 185 9260 186
rect 9275 185 9288 186
rect 9135 172 9183 176
rect 9018 150 9048 159
rect 9111 152 9126 159
rect 9147 150 9183 172
rect 8994 146 9183 150
rect 9009 143 9183 146
rect 9002 140 9183 143
rect 8811 120 8824 122
rect 8839 120 8873 122
rect 8811 104 8885 120
rect 8912 116 8925 130
rect 8940 116 8956 132
rect 9002 127 9013 140
rect 8795 82 8796 98
rect 8811 82 8824 104
rect 8839 82 8869 104
rect 8912 100 8974 116
rect 9002 109 9013 125
rect 9018 120 9028 140
rect 9038 120 9052 140
rect 9055 127 9064 140
rect 9080 127 9089 140
rect 9018 109 9052 120
rect 9055 109 9063 125
rect 9080 109 9089 125
rect 9096 120 9106 140
rect 9116 120 9130 140
rect 9131 127 9142 140
rect 9096 109 9130 120
rect 9131 109 9142 125
rect 9188 116 9204 132
rect 9211 130 9241 182
rect 9275 178 9276 185
rect 9260 170 9276 178
rect 9247 138 9260 157
rect 9275 138 9305 154
rect 9247 122 9321 138
rect 9247 120 9260 122
rect 9275 120 9309 122
rect 8912 98 8925 100
rect 8940 98 8974 100
rect 8912 82 8974 98
rect 9018 93 9031 96
rect 9096 93 9126 104
rect 9174 100 9220 116
rect 9247 104 9321 120
rect 9174 98 9208 100
rect 9173 82 9220 98
rect 9247 82 9260 104
rect 9275 82 9305 104
rect 9332 82 9333 98
rect 9348 82 9361 242
rect -9 74 32 82
rect -9 48 6 74
rect 13 48 32 74
rect 96 70 158 82
rect 170 70 245 82
rect 303 70 378 82
rect 390 70 421 82
rect 427 70 462 82
rect 96 68 258 70
rect -9 40 32 48
rect 114 40 127 68
rect 142 66 157 68
rect 181 41 188 48
rect 191 40 258 68
rect 290 68 462 70
rect 260 46 288 50
rect 290 46 370 68
rect 391 66 406 68
rect 260 44 370 46
rect 260 40 288 44
rect 290 40 370 44
rect -3 30 -2 40
rect 13 30 26 40
rect 41 30 71 40
rect 114 30 157 40
rect 164 30 172 40
rect 191 32 194 40
rect 258 32 290 40
rect 191 30 357 32
rect 376 30 387 40
rect 391 30 421 40
rect 449 30 462 68
rect 534 74 569 82
rect 534 48 535 74
rect 542 48 569 74
rect 534 40 569 48
rect 571 74 612 82
rect 571 48 586 74
rect 593 48 612 74
rect 676 70 738 82
rect 750 70 825 82
rect 883 70 958 82
rect 970 70 1001 82
rect 1007 70 1042 82
rect 676 68 838 70
rect 571 40 612 48
rect 694 40 707 68
rect 722 66 737 68
rect 761 41 768 48
rect 771 40 838 68
rect 870 68 1042 70
rect 840 46 868 50
rect 870 46 950 68
rect 971 66 986 68
rect 840 44 950 46
rect 840 40 868 44
rect 870 40 950 44
rect 477 30 507 40
rect 534 30 535 40
rect 550 30 563 40
rect 577 30 578 40
rect 593 30 606 40
rect 621 30 651 40
rect 694 30 737 40
rect 744 30 752 40
rect 771 32 774 40
rect 838 32 870 40
rect 771 30 937 32
rect 956 30 967 40
rect 971 30 1001 40
rect 1029 30 1042 68
rect 1114 74 1149 82
rect 1114 48 1115 74
rect 1122 48 1149 74
rect 1114 40 1149 48
rect 1151 74 1192 82
rect 1151 48 1166 74
rect 1173 48 1192 74
rect 1256 70 1318 82
rect 1330 70 1405 82
rect 1463 70 1538 82
rect 1550 70 1581 82
rect 1587 70 1622 82
rect 1256 68 1418 70
rect 1151 40 1192 48
rect 1274 40 1287 68
rect 1302 66 1317 68
rect 1341 41 1348 48
rect 1351 40 1418 68
rect 1450 68 1622 70
rect 1420 46 1448 50
rect 1450 46 1530 68
rect 1551 66 1566 68
rect 1420 44 1530 46
rect 1420 40 1448 44
rect 1450 40 1530 44
rect 1057 30 1087 40
rect 1114 30 1115 40
rect 1130 30 1143 40
rect 1157 30 1158 40
rect 1173 30 1186 40
rect 1201 30 1231 40
rect 1274 30 1317 40
rect 1324 30 1332 40
rect 1351 32 1354 40
rect 1418 32 1450 40
rect 1351 30 1517 32
rect 1536 30 1547 40
rect 1551 30 1581 40
rect 1609 30 1622 68
rect 1694 74 1729 82
rect 1694 48 1695 74
rect 1702 48 1729 74
rect 1694 40 1729 48
rect 1731 74 1772 82
rect 1731 48 1746 74
rect 1753 48 1772 74
rect 1836 70 1898 82
rect 1910 70 1985 82
rect 2043 70 2118 82
rect 2130 70 2161 82
rect 2167 70 2202 82
rect 1836 68 1998 70
rect 1731 40 1772 48
rect 1854 40 1867 68
rect 1882 66 1897 68
rect 1921 41 1928 48
rect 1931 40 1998 68
rect 2030 68 2202 70
rect 2000 46 2028 50
rect 2030 46 2110 68
rect 2131 66 2146 68
rect 2000 44 2110 46
rect 2000 40 2028 44
rect 2030 40 2110 44
rect 1637 30 1667 40
rect 1694 30 1695 40
rect 1710 30 1723 40
rect 1737 30 1738 40
rect 1753 30 1766 40
rect 1781 30 1811 40
rect 1854 30 1897 40
rect 1904 30 1912 40
rect 1931 32 1934 40
rect 1998 32 2030 40
rect 1931 30 2097 32
rect 2116 30 2127 40
rect 2131 30 2161 40
rect 2189 30 2202 68
rect 2274 74 2309 82
rect 2274 48 2275 74
rect 2282 48 2309 74
rect 2274 40 2309 48
rect 2311 74 2352 82
rect 2311 48 2326 74
rect 2333 48 2352 74
rect 2416 70 2478 82
rect 2490 70 2565 82
rect 2623 70 2698 82
rect 2710 70 2741 82
rect 2747 70 2782 82
rect 2416 68 2578 70
rect 2311 40 2352 48
rect 2434 40 2447 68
rect 2462 66 2477 68
rect 2501 41 2508 48
rect 2511 40 2578 68
rect 2610 68 2782 70
rect 2580 46 2608 50
rect 2610 46 2690 68
rect 2711 66 2726 68
rect 2580 44 2690 46
rect 2580 40 2608 44
rect 2610 40 2690 44
rect 2217 30 2247 40
rect 2274 30 2275 40
rect 2290 30 2303 40
rect 2317 30 2318 40
rect 2333 30 2346 40
rect 2361 30 2391 40
rect 2434 30 2477 40
rect 2484 30 2492 40
rect 2511 32 2514 40
rect 2578 32 2610 40
rect 2511 30 2677 32
rect 2696 30 2707 40
rect 2711 30 2741 40
rect 2769 30 2782 68
rect 2854 74 2889 82
rect 2854 48 2855 74
rect 2862 48 2889 74
rect 2854 40 2889 48
rect 2891 74 2932 82
rect 2891 48 2906 74
rect 2913 48 2932 74
rect 2996 70 3058 82
rect 3070 70 3145 82
rect 3203 70 3278 82
rect 3290 70 3321 82
rect 3327 70 3362 82
rect 2996 68 3158 70
rect 2891 40 2932 48
rect 3014 40 3027 68
rect 3042 66 3057 68
rect 3081 41 3088 48
rect 3091 40 3158 68
rect 3190 68 3362 70
rect 3160 46 3188 50
rect 3190 46 3270 68
rect 3291 66 3306 68
rect 3160 44 3270 46
rect 3160 40 3188 44
rect 3190 40 3270 44
rect 2797 30 2827 40
rect 2854 30 2855 40
rect 2870 30 2883 40
rect 2897 30 2898 40
rect 2913 30 2926 40
rect 2941 30 2971 40
rect 3014 30 3057 40
rect 3064 30 3072 40
rect 3091 32 3094 40
rect 3158 32 3190 40
rect 3091 30 3257 32
rect 3276 30 3287 40
rect 3291 30 3321 40
rect 3349 30 3362 68
rect 3434 74 3469 82
rect 3434 48 3435 74
rect 3442 48 3469 74
rect 3434 40 3469 48
rect 3377 30 3407 40
rect 3434 30 3435 40
rect 3450 30 3463 40
rect -3 24 3469 30
rect -2 16 3469 24
rect 5889 74 5930 82
rect 5889 48 5904 74
rect 5911 48 5930 74
rect 5994 70 6056 82
rect 6068 70 6143 82
rect 6201 70 6276 82
rect 6288 70 6319 82
rect 6325 70 6360 82
rect 5994 68 6156 70
rect 5889 40 5930 48
rect 6012 40 6025 68
rect 6040 66 6055 68
rect 6079 41 6086 48
rect 6089 40 6156 68
rect 6188 68 6360 70
rect 6158 46 6186 50
rect 6188 46 6268 68
rect 6289 66 6304 68
rect 6158 44 6268 46
rect 6158 40 6186 44
rect 6188 40 6268 44
rect 5895 30 5896 40
rect 5911 30 5924 40
rect 5939 30 5969 40
rect 6012 30 6055 40
rect 6062 30 6070 40
rect 6089 32 6092 40
rect 6156 32 6188 40
rect 6089 30 6255 32
rect 6274 30 6285 40
rect 6289 30 6319 40
rect 6347 30 6360 68
rect 6432 74 6467 82
rect 6432 48 6433 74
rect 6440 48 6467 74
rect 6432 40 6467 48
rect 6469 74 6510 82
rect 6469 48 6484 74
rect 6491 48 6510 74
rect 6574 70 6636 82
rect 6648 70 6723 82
rect 6781 70 6856 82
rect 6868 70 6899 82
rect 6905 70 6940 82
rect 6574 68 6736 70
rect 6469 40 6510 48
rect 6592 40 6605 68
rect 6620 66 6635 68
rect 6659 41 6666 48
rect 6669 40 6736 68
rect 6768 68 6940 70
rect 6738 46 6766 50
rect 6768 46 6848 68
rect 6869 66 6884 68
rect 6738 44 6848 46
rect 6738 40 6766 44
rect 6768 40 6848 44
rect 6375 30 6405 40
rect 6432 30 6433 40
rect 6448 30 6461 40
rect 6475 30 6476 40
rect 6491 30 6504 40
rect 6519 30 6549 40
rect 6592 30 6635 40
rect 6642 30 6650 40
rect 6669 32 6672 40
rect 6736 32 6768 40
rect 6669 30 6835 32
rect 6854 30 6865 40
rect 6869 30 6899 40
rect 6927 30 6940 68
rect 7012 74 7047 82
rect 7012 48 7013 74
rect 7020 48 7047 74
rect 7012 40 7047 48
rect 7049 74 7090 82
rect 7049 48 7064 74
rect 7071 48 7090 74
rect 7154 70 7216 82
rect 7228 70 7303 82
rect 7361 70 7436 82
rect 7448 70 7479 82
rect 7485 70 7520 82
rect 7154 68 7316 70
rect 7049 40 7090 48
rect 7172 40 7185 68
rect 7200 66 7215 68
rect 7239 41 7246 48
rect 7249 40 7316 68
rect 7348 68 7520 70
rect 7318 46 7346 50
rect 7348 46 7428 68
rect 7449 66 7464 68
rect 7318 44 7428 46
rect 7318 40 7346 44
rect 7348 40 7428 44
rect 6955 30 6985 40
rect 7012 30 7013 40
rect 7028 30 7041 40
rect 7055 30 7056 40
rect 7071 30 7084 40
rect 7099 30 7129 40
rect 7172 30 7215 40
rect 7222 30 7230 40
rect 7249 32 7252 40
rect 7316 32 7348 40
rect 7249 30 7415 32
rect 7434 30 7445 40
rect 7449 30 7479 40
rect 7507 30 7520 68
rect 7592 74 7627 82
rect 7592 48 7593 74
rect 7600 48 7627 74
rect 7592 40 7627 48
rect 7629 74 7670 82
rect 7629 48 7644 74
rect 7651 48 7670 74
rect 7734 70 7796 82
rect 7808 70 7883 82
rect 7941 70 8016 82
rect 8028 70 8059 82
rect 8065 70 8100 82
rect 7734 68 7896 70
rect 7629 40 7670 48
rect 7752 40 7765 68
rect 7780 66 7795 68
rect 7819 41 7826 48
rect 7829 40 7896 68
rect 7928 68 8100 70
rect 7898 46 7926 50
rect 7928 46 8008 68
rect 8029 66 8044 68
rect 7898 44 8008 46
rect 7898 40 7926 44
rect 7928 40 8008 44
rect 7535 30 7565 40
rect 7592 30 7593 40
rect 7608 30 7621 40
rect 7635 30 7636 40
rect 7651 30 7664 40
rect 7679 30 7709 40
rect 7752 30 7795 40
rect 7802 30 7810 40
rect 7829 32 7832 40
rect 7896 32 7928 40
rect 7829 30 7995 32
rect 8014 30 8025 40
rect 8029 30 8059 40
rect 8087 30 8100 68
rect 8172 74 8207 82
rect 8172 48 8173 74
rect 8180 48 8207 74
rect 8172 40 8207 48
rect 8209 74 8250 82
rect 8209 48 8224 74
rect 8231 48 8250 74
rect 8314 70 8376 82
rect 8388 70 8463 82
rect 8521 70 8596 82
rect 8608 70 8639 82
rect 8645 70 8680 82
rect 8314 68 8476 70
rect 8209 40 8250 48
rect 8332 40 8345 68
rect 8360 66 8375 68
rect 8399 41 8406 48
rect 8409 40 8476 68
rect 8508 68 8680 70
rect 8478 46 8506 50
rect 8508 46 8588 68
rect 8609 66 8624 68
rect 8478 44 8588 46
rect 8478 40 8506 44
rect 8508 40 8588 44
rect 8115 30 8145 40
rect 8172 30 8173 40
rect 8188 30 8201 40
rect 8215 30 8216 40
rect 8231 30 8244 40
rect 8259 30 8289 40
rect 8332 30 8375 40
rect 8382 30 8390 40
rect 8409 32 8412 40
rect 8476 32 8508 40
rect 8409 30 8575 32
rect 8594 30 8605 40
rect 8609 30 8639 40
rect 8667 30 8680 68
rect 8752 74 8787 82
rect 8752 48 8753 74
rect 8760 48 8787 74
rect 8752 40 8787 48
rect 8789 74 8830 82
rect 8789 48 8804 74
rect 8811 48 8830 74
rect 8894 70 8956 82
rect 8968 70 9043 82
rect 9101 70 9176 82
rect 9188 70 9219 82
rect 9225 70 9260 82
rect 8894 68 9056 70
rect 8789 40 8830 48
rect 8912 40 8925 68
rect 8940 66 8955 68
rect 8979 41 8986 48
rect 8989 40 9056 68
rect 9088 68 9260 70
rect 9058 46 9086 50
rect 9088 46 9168 68
rect 9189 66 9204 68
rect 9058 44 9168 46
rect 9058 40 9086 44
rect 9088 40 9168 44
rect 8695 30 8725 40
rect 8752 30 8753 40
rect 8768 30 8781 40
rect 8795 30 8796 40
rect 8811 30 8824 40
rect 8839 30 8869 40
rect 8912 30 8955 40
rect 8962 30 8970 40
rect 8989 32 8992 40
rect 9056 32 9088 40
rect 8989 30 9155 32
rect 9174 30 9185 40
rect 9189 30 9219 40
rect 9247 30 9260 68
rect 9332 74 9367 82
rect 9332 48 9333 74
rect 9340 48 9367 74
rect 9332 40 9367 48
rect 9275 30 9305 40
rect 9332 30 9333 40
rect 9348 30 9361 40
rect 5889 16 9361 30
rect 13 2 26 16
rect 41 -2 71 16
rect 114 2 127 16
rect 164 3 172 16
rect 205 3 343 16
rect 376 3 384 16
rect 241 2 292 3
rect 449 2 462 16
rect 242 0 306 2
rect 477 -2 507 16
rect 550 2 563 16
rect 593 2 606 16
rect 621 -2 651 16
rect 694 2 707 16
rect 744 3 752 16
rect 785 3 923 16
rect 956 3 964 16
rect 821 2 872 3
rect 1029 2 1042 16
rect 822 0 886 2
rect 1057 -2 1087 16
rect 1130 2 1143 16
rect 1173 2 1186 16
rect 1201 -2 1231 16
rect 1274 2 1287 16
rect 1324 3 1332 16
rect 1365 3 1503 16
rect 1536 3 1544 16
rect 1401 2 1452 3
rect 1609 2 1622 16
rect 1402 0 1466 2
rect 1637 -2 1667 16
rect 1710 2 1723 16
rect 1753 2 1766 16
rect 1781 -2 1811 16
rect 1854 2 1867 16
rect 1904 3 1912 16
rect 1945 3 2083 16
rect 2116 3 2124 16
rect 1981 2 2032 3
rect 2189 2 2202 16
rect 1982 0 2046 2
rect 2217 -2 2247 16
rect 2290 2 2303 16
rect 2333 2 2346 16
rect 2361 -2 2391 16
rect 2434 2 2447 16
rect 2484 3 2492 16
rect 2525 3 2663 16
rect 2696 3 2704 16
rect 2561 2 2612 3
rect 2769 2 2782 16
rect 2562 0 2626 2
rect 2797 -2 2827 16
rect 2870 2 2883 16
rect 2913 2 2926 16
rect 2941 -2 2971 16
rect 3014 2 3027 16
rect 3064 3 3072 16
rect 3105 3 3243 16
rect 3276 3 3284 16
rect 3141 2 3192 3
rect 3349 2 3362 16
rect 3142 0 3206 2
rect 3377 -2 3407 16
rect 3450 2 3463 16
rect 5911 2 5924 16
rect 5939 -2 5969 16
rect 6012 2 6025 16
rect 6062 3 6070 16
rect 6103 3 6241 16
rect 6274 3 6282 16
rect 6139 2 6190 3
rect 6347 2 6360 16
rect 6140 0 6204 2
rect 6375 -2 6405 16
rect 6448 2 6461 16
rect 6491 2 6504 16
rect 6519 -2 6549 16
rect 6592 2 6605 16
rect 6642 3 6650 16
rect 6683 3 6821 16
rect 6854 3 6862 16
rect 6719 2 6770 3
rect 6927 2 6940 16
rect 6720 0 6784 2
rect 6955 -2 6985 16
rect 7028 2 7041 16
rect 7071 2 7084 16
rect 7099 -2 7129 16
rect 7172 2 7185 16
rect 7222 3 7230 16
rect 7263 3 7401 16
rect 7434 3 7442 16
rect 7299 2 7350 3
rect 7507 2 7520 16
rect 7300 0 7364 2
rect 7535 -2 7565 16
rect 7608 2 7621 16
rect 7651 2 7664 16
rect 7679 -2 7709 16
rect 7752 2 7765 16
rect 7802 3 7810 16
rect 7843 3 7981 16
rect 8014 3 8022 16
rect 7879 2 7930 3
rect 8087 2 8100 16
rect 7880 0 7944 2
rect 8115 -2 8145 16
rect 8188 2 8201 16
rect 8231 2 8244 16
rect 8259 -2 8289 16
rect 8332 2 8345 16
rect 8382 3 8390 16
rect 8423 3 8561 16
rect 8594 3 8602 16
rect 8459 2 8510 3
rect 8667 2 8680 16
rect 8460 0 8524 2
rect 8695 -2 8725 16
rect 8768 2 8781 16
rect 8811 2 8824 16
rect 8839 -2 8869 16
rect 8912 2 8925 16
rect 8962 3 8970 16
rect 9003 3 9141 16
rect 9174 3 9182 16
rect 9039 2 9090 3
rect 9247 2 9260 16
rect 9040 0 9104 2
rect 9275 -2 9305 16
rect 9348 2 9361 16
<< error_s >>
rect 3493 2146 3506 2162
rect 3595 2160 3608 2162
rect 3561 2146 3576 2160
rect 3585 2146 3615 2160
rect 3676 2158 3829 2204
rect 3658 2146 3850 2158
rect 3893 2146 3923 2160
rect 3929 2146 3942 2162
rect 4030 2146 4043 2162
rect 4073 2146 4086 2162
rect 4175 2160 4188 2162
rect 4141 2146 4156 2160
rect 4165 2146 4195 2160
rect 4256 2158 4409 2204
rect 4238 2146 4430 2158
rect 4473 2146 4503 2160
rect 4509 2146 4522 2162
rect 4610 2146 4623 2162
rect 4751 2146 4764 2162
rect 4853 2160 4866 2162
rect 4819 2146 4834 2160
rect 4843 2146 4873 2160
rect 4934 2158 5087 2204
rect 4916 2146 5108 2158
rect 5151 2146 5181 2160
rect 5187 2146 5200 2162
rect 5288 2146 5301 2162
rect 5331 2146 5344 2162
rect 5433 2160 5446 2162
rect 5399 2146 5414 2160
rect 5423 2146 5453 2160
rect 5514 2158 5667 2204
rect 5496 2146 5688 2158
rect 5731 2146 5761 2160
rect 5767 2146 5780 2162
rect 5868 2146 5881 2162
rect 3469 2132 4623 2146
rect 4736 2132 5889 2146
rect 3493 2028 3506 2132
rect 3551 2110 3552 2120
rect 3567 2110 3580 2120
rect 3551 2106 3580 2110
rect 3585 2106 3615 2132
rect 3633 2118 3649 2120
rect 3721 2118 3774 2132
rect 3722 2116 3786 2118
rect 3829 2116 3844 2132
rect 3893 2129 3923 2132
rect 3893 2126 3929 2129
rect 3859 2118 3875 2120
rect 3633 2106 3648 2110
rect 3551 2104 3648 2106
rect 3676 2104 3844 2116
rect 3860 2106 3875 2110
rect 3893 2107 3932 2126
rect 3951 2120 3958 2121
rect 3957 2113 3958 2120
rect 3941 2110 3942 2113
rect 3957 2110 3970 2113
rect 3893 2106 3923 2107
rect 3932 2106 3938 2107
rect 3941 2106 3970 2110
rect 3860 2105 3970 2106
rect 3860 2104 3976 2105
rect 3535 2096 3586 2104
rect 3535 2084 3560 2096
rect 3567 2084 3586 2096
rect 3617 2096 3667 2104
rect 3617 2088 3633 2096
rect 3640 2094 3667 2096
rect 3676 2094 3897 2104
rect 3640 2084 3897 2094
rect 3926 2096 3976 2104
rect 3926 2087 3942 2096
rect 3535 2076 3586 2084
rect 3633 2076 3897 2084
rect 3923 2084 3942 2087
rect 3949 2084 3976 2096
rect 3923 2076 3976 2084
rect 3551 2068 3552 2076
rect 3567 2068 3580 2076
rect 3551 2060 3567 2068
rect 3548 2053 3567 2056
rect 3548 2044 3570 2053
rect 3521 2034 3570 2044
rect 3521 2028 3551 2034
rect 3570 2029 3575 2034
rect 3493 2012 3567 2028
rect 3585 2020 3615 2076
rect 3650 2066 3858 2076
rect 3893 2072 3938 2076
rect 3941 2075 3942 2076
rect 3957 2075 3970 2076
rect 3676 2036 3865 2066
rect 3691 2033 3865 2036
rect 3684 2030 3865 2033
rect 3493 2010 3506 2012
rect 3521 2010 3555 2012
rect 3493 1994 3567 2010
rect 3594 2006 3607 2020
rect 3622 2006 3638 2022
rect 3684 2017 3695 2030
rect 3477 1972 3478 1988
rect 3493 1972 3506 1994
rect 3521 1972 3551 1994
rect 3594 1990 3656 2006
rect 3684 1999 3695 2015
rect 3700 2010 3710 2030
rect 3720 2010 3734 2030
rect 3737 2017 3746 2030
rect 3762 2017 3771 2030
rect 3700 1999 3734 2010
rect 3737 1999 3746 2015
rect 3762 1999 3771 2015
rect 3778 2010 3788 2030
rect 3798 2010 3812 2030
rect 3813 2017 3824 2030
rect 3778 1999 3812 2010
rect 3813 1999 3824 2015
rect 3870 2006 3886 2022
rect 3893 2020 3923 2072
rect 3957 2068 3958 2075
rect 3942 2060 3958 2068
rect 3929 2028 3942 2047
rect 3957 2028 3987 2044
rect 3929 2012 4003 2028
rect 3929 2010 3942 2012
rect 3957 2010 3991 2012
rect 3594 1988 3607 1990
rect 3622 1988 3656 1990
rect 3594 1972 3656 1988
rect 3700 1983 3716 1986
rect 3778 1983 3808 1994
rect 3856 1990 3902 2006
rect 3929 1994 4003 2010
rect 3856 1988 3890 1990
rect 3855 1972 3902 1988
rect 3929 1972 3942 1994
rect 3957 1972 3987 1994
rect 4014 1972 4015 1988
rect 4030 1972 4043 2132
rect 4073 2028 4086 2132
rect 4131 2110 4132 2120
rect 4147 2110 4160 2120
rect 4131 2106 4160 2110
rect 4165 2106 4195 2132
rect 4213 2118 4229 2120
rect 4301 2118 4354 2132
rect 4302 2116 4366 2118
rect 4409 2116 4424 2132
rect 4473 2129 4503 2132
rect 4473 2126 4509 2129
rect 4439 2118 4455 2120
rect 4213 2106 4228 2110
rect 4131 2104 4228 2106
rect 4256 2104 4424 2116
rect 4440 2106 4455 2110
rect 4473 2107 4512 2126
rect 4531 2120 4538 2121
rect 4537 2113 4538 2120
rect 4521 2110 4522 2113
rect 4537 2110 4550 2113
rect 4473 2106 4503 2107
rect 4512 2106 4518 2107
rect 4521 2106 4550 2110
rect 4440 2105 4550 2106
rect 4440 2104 4556 2105
rect 4115 2096 4166 2104
rect 4115 2084 4140 2096
rect 4147 2084 4166 2096
rect 4197 2096 4247 2104
rect 4197 2088 4213 2096
rect 4220 2094 4247 2096
rect 4256 2094 4477 2104
rect 4220 2084 4477 2094
rect 4506 2096 4556 2104
rect 4506 2087 4522 2096
rect 4115 2076 4166 2084
rect 4213 2076 4477 2084
rect 4503 2084 4522 2087
rect 4529 2084 4556 2096
rect 4503 2076 4556 2084
rect 4131 2068 4132 2076
rect 4147 2068 4160 2076
rect 4131 2060 4147 2068
rect 4128 2053 4147 2056
rect 4128 2044 4150 2053
rect 4101 2034 4150 2044
rect 4101 2028 4131 2034
rect 4150 2029 4155 2034
rect 4073 2012 4147 2028
rect 4165 2020 4195 2076
rect 4230 2066 4438 2076
rect 4473 2072 4518 2076
rect 4521 2075 4522 2076
rect 4537 2075 4550 2076
rect 4256 2036 4445 2066
rect 4271 2033 4445 2036
rect 4264 2030 4445 2033
rect 4073 2010 4086 2012
rect 4101 2010 4135 2012
rect 4073 1994 4147 2010
rect 4174 2006 4187 2020
rect 4202 2006 4218 2022
rect 4264 2017 4275 2030
rect 4057 1972 4058 1988
rect 4073 1972 4086 1994
rect 4101 1972 4131 1994
rect 4174 1990 4236 2006
rect 4264 1999 4275 2015
rect 4280 2010 4290 2030
rect 4300 2010 4314 2030
rect 4317 2017 4326 2030
rect 4342 2017 4351 2030
rect 4280 1999 4314 2010
rect 4317 1999 4326 2015
rect 4342 1999 4351 2015
rect 4358 2010 4368 2030
rect 4378 2010 4392 2030
rect 4393 2017 4404 2030
rect 4358 1999 4392 2010
rect 4393 1999 4404 2015
rect 4450 2006 4466 2022
rect 4473 2020 4503 2072
rect 4537 2068 4538 2075
rect 4522 2060 4538 2068
rect 4509 2028 4522 2047
rect 4537 2028 4567 2044
rect 4509 2012 4583 2028
rect 4509 2010 4522 2012
rect 4537 2010 4571 2012
rect 4174 1988 4187 1990
rect 4202 1988 4236 1990
rect 4174 1972 4236 1988
rect 4280 1983 4296 1986
rect 4358 1983 4388 1994
rect 4436 1990 4482 2006
rect 4509 1994 4583 2010
rect 4436 1988 4470 1990
rect 4435 1972 4482 1988
rect 4509 1972 4522 1994
rect 4537 1972 4567 1994
rect 4594 1972 4595 1988
rect 4610 1972 4623 2132
rect 4751 2028 4764 2132
rect 4809 2110 4810 2120
rect 4825 2110 4838 2120
rect 4809 2106 4838 2110
rect 4843 2106 4873 2132
rect 4891 2118 4907 2120
rect 4979 2118 5032 2132
rect 4980 2116 5044 2118
rect 5087 2116 5102 2132
rect 5151 2129 5181 2132
rect 5151 2126 5187 2129
rect 5117 2118 5133 2120
rect 4891 2106 4906 2110
rect 4809 2104 4906 2106
rect 4934 2104 5102 2116
rect 5118 2106 5133 2110
rect 5151 2107 5190 2126
rect 5209 2120 5216 2121
rect 5215 2113 5216 2120
rect 5199 2110 5200 2113
rect 5215 2110 5228 2113
rect 5151 2106 5181 2107
rect 5190 2106 5196 2107
rect 5199 2106 5228 2110
rect 5118 2105 5228 2106
rect 5118 2104 5234 2105
rect 4793 2096 4844 2104
rect 4793 2084 4818 2096
rect 4825 2084 4844 2096
rect 4875 2096 4925 2104
rect 4875 2088 4891 2096
rect 4898 2094 4925 2096
rect 4934 2094 5155 2104
rect 4898 2084 5155 2094
rect 5184 2096 5234 2104
rect 5184 2087 5200 2096
rect 4793 2076 4844 2084
rect 4891 2076 5155 2084
rect 5181 2084 5200 2087
rect 5207 2084 5234 2096
rect 5181 2076 5234 2084
rect 4809 2068 4810 2076
rect 4825 2068 4838 2076
rect 4809 2060 4825 2068
rect 4806 2053 4825 2056
rect 4806 2044 4828 2053
rect 4779 2034 4828 2044
rect 4779 2028 4809 2034
rect 4828 2029 4833 2034
rect 4751 2012 4825 2028
rect 4843 2020 4873 2076
rect 4908 2066 5116 2076
rect 5151 2072 5196 2076
rect 5199 2075 5200 2076
rect 5215 2075 5228 2076
rect 4934 2036 5123 2066
rect 4949 2033 5123 2036
rect 4942 2030 5123 2033
rect 4751 2010 4764 2012
rect 4779 2010 4813 2012
rect 4751 1994 4825 2010
rect 4852 2006 4865 2020
rect 4880 2006 4896 2022
rect 4942 2017 4953 2030
rect 4735 1972 4736 1988
rect 4751 1972 4764 1994
rect 4779 1972 4809 1994
rect 4852 1990 4914 2006
rect 4942 1999 4953 2015
rect 4958 2010 4968 2030
rect 4978 2010 4992 2030
rect 4995 2017 5004 2030
rect 5020 2017 5029 2030
rect 4958 1999 4992 2010
rect 4995 1999 5004 2015
rect 5020 1999 5029 2015
rect 5036 2010 5046 2030
rect 5056 2010 5070 2030
rect 5071 2017 5082 2030
rect 5036 1999 5070 2010
rect 5071 1999 5082 2015
rect 5128 2006 5144 2022
rect 5151 2020 5181 2072
rect 5215 2068 5216 2075
rect 5200 2060 5216 2068
rect 5187 2028 5200 2047
rect 5215 2028 5245 2044
rect 5187 2012 5261 2028
rect 5187 2010 5200 2012
rect 5215 2010 5249 2012
rect 4852 1988 4865 1990
rect 4880 1988 4914 1990
rect 4852 1972 4914 1988
rect 4958 1983 4974 1986
rect 5036 1983 5066 1994
rect 5114 1990 5160 2006
rect 5187 1994 5261 2010
rect 5114 1988 5148 1990
rect 5113 1972 5160 1988
rect 5187 1972 5200 1994
rect 5215 1972 5245 1994
rect 5272 1972 5273 1988
rect 5288 1972 5301 2132
rect 5331 2028 5344 2132
rect 5389 2110 5390 2120
rect 5405 2110 5418 2120
rect 5389 2106 5418 2110
rect 5423 2106 5453 2132
rect 5471 2118 5487 2120
rect 5559 2118 5612 2132
rect 5560 2116 5624 2118
rect 5667 2116 5682 2132
rect 5731 2129 5761 2132
rect 5731 2126 5767 2129
rect 5697 2118 5713 2120
rect 5471 2106 5486 2110
rect 5389 2104 5486 2106
rect 5514 2104 5682 2116
rect 5698 2106 5713 2110
rect 5731 2107 5770 2126
rect 5789 2120 5796 2121
rect 5795 2113 5796 2120
rect 5779 2110 5780 2113
rect 5795 2110 5808 2113
rect 5731 2106 5761 2107
rect 5770 2106 5776 2107
rect 5779 2106 5808 2110
rect 5698 2105 5808 2106
rect 5698 2104 5814 2105
rect 5373 2096 5424 2104
rect 5373 2084 5398 2096
rect 5405 2084 5424 2096
rect 5455 2096 5505 2104
rect 5455 2088 5471 2096
rect 5478 2094 5505 2096
rect 5514 2094 5735 2104
rect 5478 2084 5735 2094
rect 5764 2096 5814 2104
rect 5764 2087 5780 2096
rect 5373 2076 5424 2084
rect 5471 2076 5735 2084
rect 5761 2084 5780 2087
rect 5787 2084 5814 2096
rect 5761 2076 5814 2084
rect 5389 2068 5390 2076
rect 5405 2068 5418 2076
rect 5389 2060 5405 2068
rect 5386 2053 5405 2056
rect 5386 2044 5408 2053
rect 5359 2034 5408 2044
rect 5359 2028 5389 2034
rect 5408 2029 5413 2034
rect 5331 2012 5405 2028
rect 5423 2020 5453 2076
rect 5488 2066 5696 2076
rect 5731 2072 5776 2076
rect 5779 2075 5780 2076
rect 5795 2075 5808 2076
rect 5514 2036 5703 2066
rect 5529 2033 5703 2036
rect 5522 2030 5703 2033
rect 5331 2010 5344 2012
rect 5359 2010 5393 2012
rect 5331 1994 5405 2010
rect 5432 2006 5445 2020
rect 5460 2006 5476 2022
rect 5522 2017 5533 2030
rect 5315 1972 5316 1988
rect 5331 1972 5344 1994
rect 5359 1972 5389 1994
rect 5432 1990 5494 2006
rect 5522 1999 5533 2015
rect 5538 2010 5548 2030
rect 5558 2010 5572 2030
rect 5575 2017 5584 2030
rect 5600 2017 5609 2030
rect 5538 1999 5572 2010
rect 5575 1999 5584 2015
rect 5600 1999 5609 2015
rect 5616 2010 5626 2030
rect 5636 2010 5650 2030
rect 5651 2017 5662 2030
rect 5616 1999 5650 2010
rect 5651 1999 5662 2015
rect 5708 2006 5724 2022
rect 5731 2020 5761 2072
rect 5795 2068 5796 2075
rect 5780 2060 5796 2068
rect 5767 2028 5780 2047
rect 5795 2028 5825 2044
rect 5767 2012 5841 2028
rect 5767 2010 5780 2012
rect 5795 2010 5829 2012
rect 5432 1988 5445 1990
rect 5460 1988 5494 1990
rect 5432 1972 5494 1988
rect 5538 1983 5554 1986
rect 5616 1983 5646 1994
rect 5694 1990 5740 2006
rect 5767 1994 5841 2010
rect 5694 1988 5728 1990
rect 5693 1972 5740 1988
rect 5767 1972 5780 1994
rect 5795 1972 5825 1994
rect 5852 1972 5853 1988
rect 5868 1972 5881 2132
rect 3471 1964 3512 1972
rect 3471 1938 3486 1964
rect 3493 1938 3512 1964
rect 3576 1960 3638 1972
rect 3650 1960 3725 1972
rect 3783 1960 3858 1972
rect 3870 1960 3901 1972
rect 3907 1960 3942 1972
rect 3576 1958 3738 1960
rect 3471 1930 3512 1938
rect 3594 1934 3607 1958
rect 3622 1956 3637 1958
rect 3477 1920 3478 1930
rect 3493 1920 3506 1930
rect 3521 1920 3551 1934
rect 3594 1920 3637 1934
rect 3661 1931 3668 1938
rect 3671 1934 3738 1958
rect 3770 1958 3942 1960
rect 3740 1936 3768 1940
rect 3770 1936 3850 1958
rect 3871 1956 3886 1958
rect 3740 1934 3850 1936
rect 3671 1930 3850 1934
rect 3644 1920 3674 1930
rect 3676 1920 3829 1930
rect 3837 1920 3867 1930
rect 3871 1920 3901 1934
rect 3929 1920 3942 1958
rect 4014 1964 4049 1972
rect 4014 1938 4015 1964
rect 4022 1938 4049 1964
rect 3957 1920 3987 1934
rect 4014 1930 4049 1938
rect 4051 1964 4092 1972
rect 4051 1938 4066 1964
rect 4073 1938 4092 1964
rect 4156 1960 4218 1972
rect 4230 1960 4305 1972
rect 4363 1960 4438 1972
rect 4450 1960 4481 1972
rect 4487 1960 4522 1972
rect 4156 1958 4318 1960
rect 4051 1930 4092 1938
rect 4174 1934 4187 1958
rect 4202 1956 4217 1958
rect 4014 1920 4015 1930
rect 4030 1920 4043 1930
rect 4057 1920 4058 1930
rect 4073 1920 4086 1930
rect 4101 1920 4131 1934
rect 4174 1920 4217 1934
rect 4241 1931 4248 1938
rect 4251 1934 4318 1958
rect 4350 1958 4522 1960
rect 4320 1936 4348 1940
rect 4350 1936 4430 1958
rect 4451 1956 4466 1958
rect 4320 1934 4430 1936
rect 4251 1930 4430 1934
rect 4224 1920 4254 1930
rect 4256 1920 4409 1930
rect 4417 1920 4447 1930
rect 4451 1920 4481 1934
rect 4509 1920 4522 1958
rect 4594 1964 4629 1972
rect 4594 1938 4595 1964
rect 4602 1938 4629 1964
rect 4537 1920 4567 1934
rect 4594 1930 4629 1938
rect 4729 1964 4770 1972
rect 4729 1938 4744 1964
rect 4751 1938 4770 1964
rect 4834 1960 4896 1972
rect 4908 1960 4983 1972
rect 5041 1960 5116 1972
rect 5128 1960 5159 1972
rect 5165 1960 5200 1972
rect 4834 1958 4996 1960
rect 4729 1930 4770 1938
rect 4852 1934 4865 1958
rect 4880 1956 4895 1958
rect 4594 1920 4595 1930
rect 4610 1920 4623 1930
rect 3469 1906 4623 1920
rect 4735 1920 4736 1930
rect 4751 1920 4764 1930
rect 4779 1920 4809 1934
rect 4852 1920 4895 1934
rect 4919 1931 4926 1938
rect 4929 1934 4996 1958
rect 5028 1958 5200 1960
rect 4998 1936 5026 1940
rect 5028 1936 5108 1958
rect 5129 1956 5144 1958
rect 4998 1934 5108 1936
rect 4929 1930 5108 1934
rect 4902 1920 4932 1930
rect 4934 1920 5087 1930
rect 5095 1920 5125 1930
rect 5129 1920 5159 1934
rect 5187 1920 5200 1958
rect 5272 1964 5307 1972
rect 5272 1938 5273 1964
rect 5280 1938 5307 1964
rect 5215 1920 5245 1934
rect 5272 1930 5307 1938
rect 5309 1964 5350 1972
rect 5309 1938 5324 1964
rect 5331 1938 5350 1964
rect 5414 1960 5476 1972
rect 5488 1960 5563 1972
rect 5621 1960 5696 1972
rect 5708 1960 5739 1972
rect 5745 1960 5780 1972
rect 5414 1958 5576 1960
rect 5309 1930 5350 1938
rect 5432 1934 5445 1958
rect 5460 1956 5475 1958
rect 5272 1920 5273 1930
rect 5288 1920 5301 1930
rect 5315 1920 5316 1930
rect 5331 1920 5344 1930
rect 5359 1920 5389 1934
rect 5432 1920 5475 1934
rect 5499 1931 5506 1938
rect 5509 1934 5576 1958
rect 5608 1958 5780 1960
rect 5578 1936 5606 1940
rect 5608 1936 5688 1958
rect 5709 1956 5724 1958
rect 5578 1934 5688 1936
rect 5509 1930 5688 1934
rect 5482 1920 5512 1930
rect 5514 1920 5667 1930
rect 5675 1920 5705 1930
rect 5709 1920 5739 1934
rect 5767 1920 5780 1958
rect 5852 1964 5887 1972
rect 5852 1938 5853 1964
rect 5860 1938 5887 1964
rect 5795 1920 5825 1934
rect 5852 1930 5887 1938
rect 5852 1920 5853 1930
rect 5868 1920 5881 1930
rect 4735 1914 5889 1920
rect 4736 1906 5889 1914
rect 3493 1876 3506 1906
rect 3521 1888 3551 1906
rect 3594 1892 3608 1906
rect 3644 1892 3864 1906
rect 3595 1890 3608 1892
rect 3561 1878 3576 1890
rect 3558 1876 3580 1878
rect 3585 1876 3615 1890
rect 3676 1888 3829 1892
rect 3658 1876 3850 1888
rect 3893 1876 3923 1890
rect 3929 1876 3942 1906
rect 3957 1888 3987 1906
rect 4030 1876 4043 1906
rect 4073 1876 4086 1906
rect 4101 1888 4131 1906
rect 4174 1892 4188 1906
rect 4224 1892 4444 1906
rect 4175 1890 4188 1892
rect 4141 1878 4156 1890
rect 4138 1876 4160 1878
rect 4165 1876 4195 1890
rect 4256 1888 4409 1892
rect 4238 1876 4430 1888
rect 4473 1876 4503 1890
rect 4509 1876 4522 1906
rect 4537 1888 4567 1906
rect 4610 1876 4623 1906
rect 4751 1876 4764 1906
rect 4779 1888 4809 1906
rect 4852 1892 4866 1906
rect 4902 1892 5122 1906
rect 4853 1890 4866 1892
rect 4819 1878 4834 1890
rect 4816 1876 4838 1878
rect 4843 1876 4873 1890
rect 4934 1888 5087 1892
rect 4916 1876 5108 1888
rect 5151 1876 5181 1890
rect 5187 1876 5200 1906
rect 5215 1888 5245 1906
rect 5288 1876 5301 1906
rect 5331 1876 5344 1906
rect 5359 1888 5389 1906
rect 5432 1892 5446 1906
rect 5482 1892 5702 1906
rect 5433 1890 5446 1892
rect 5399 1878 5414 1890
rect 5396 1876 5418 1878
rect 5423 1876 5453 1890
rect 5514 1888 5667 1892
rect 5496 1876 5688 1888
rect 5731 1876 5761 1890
rect 5767 1876 5780 1906
rect 5795 1888 5825 1906
rect 5868 1876 5881 1906
rect 3469 1862 4623 1876
rect 4736 1862 5889 1876
rect 3493 1758 3506 1862
rect 3551 1840 3552 1850
rect 3567 1840 3580 1850
rect 3551 1836 3580 1840
rect 3585 1836 3615 1862
rect 3633 1848 3649 1850
rect 3721 1848 3774 1862
rect 3722 1846 3786 1848
rect 3829 1846 3844 1862
rect 3893 1859 3923 1862
rect 3893 1856 3929 1859
rect 3859 1848 3875 1850
rect 3633 1836 3648 1840
rect 3551 1834 3648 1836
rect 3676 1834 3844 1846
rect 3860 1836 3875 1840
rect 3893 1837 3932 1856
rect 3951 1850 3958 1851
rect 3957 1843 3958 1850
rect 3941 1840 3942 1843
rect 3957 1840 3970 1843
rect 3893 1836 3923 1837
rect 3932 1836 3938 1837
rect 3941 1836 3970 1840
rect 3860 1835 3970 1836
rect 3860 1834 3976 1835
rect 3535 1826 3586 1834
rect 3535 1814 3560 1826
rect 3567 1814 3586 1826
rect 3617 1826 3667 1834
rect 3617 1818 3633 1826
rect 3640 1824 3667 1826
rect 3676 1824 3897 1834
rect 3640 1814 3897 1824
rect 3926 1826 3976 1834
rect 3926 1817 3942 1826
rect 3535 1806 3586 1814
rect 3633 1806 3897 1814
rect 3923 1814 3942 1817
rect 3949 1814 3976 1826
rect 3923 1806 3976 1814
rect 3551 1798 3552 1806
rect 3567 1798 3580 1806
rect 3551 1790 3567 1798
rect 3548 1783 3567 1786
rect 3548 1774 3570 1783
rect 3521 1764 3570 1774
rect 3521 1758 3551 1764
rect 3570 1759 3575 1764
rect 3493 1742 3567 1758
rect 3585 1750 3615 1806
rect 3650 1796 3858 1806
rect 3893 1802 3938 1806
rect 3941 1805 3942 1806
rect 3957 1805 3970 1806
rect 3676 1766 3865 1796
rect 3691 1763 3865 1766
rect 3684 1760 3865 1763
rect 3493 1740 3506 1742
rect 3521 1740 3555 1742
rect 3493 1724 3567 1740
rect 3594 1736 3607 1750
rect 3622 1736 3638 1752
rect 3684 1747 3695 1760
rect 3477 1702 3478 1718
rect 3493 1702 3506 1724
rect 3521 1702 3551 1724
rect 3594 1720 3656 1736
rect 3684 1729 3695 1745
rect 3700 1740 3710 1760
rect 3720 1740 3734 1760
rect 3737 1747 3746 1760
rect 3762 1747 3771 1760
rect 3700 1729 3734 1740
rect 3737 1729 3746 1745
rect 3762 1729 3771 1745
rect 3778 1740 3788 1760
rect 3798 1740 3812 1760
rect 3813 1747 3824 1760
rect 3778 1729 3812 1740
rect 3813 1729 3824 1745
rect 3870 1736 3886 1752
rect 3893 1750 3923 1802
rect 3957 1798 3958 1805
rect 3942 1790 3958 1798
rect 3929 1758 3942 1777
rect 3957 1758 3987 1774
rect 3929 1742 4003 1758
rect 3929 1740 3942 1742
rect 3957 1740 3991 1742
rect 3594 1718 3607 1720
rect 3622 1718 3656 1720
rect 3594 1702 3656 1718
rect 3700 1713 3716 1716
rect 3778 1713 3808 1724
rect 3856 1720 3902 1736
rect 3929 1724 4003 1740
rect 3856 1718 3890 1720
rect 3855 1702 3902 1718
rect 3929 1702 3942 1724
rect 3957 1702 3987 1724
rect 4014 1702 4015 1718
rect 4030 1702 4043 1862
rect 4073 1758 4086 1862
rect 4131 1840 4132 1850
rect 4147 1840 4160 1850
rect 4131 1836 4160 1840
rect 4165 1836 4195 1862
rect 4213 1848 4229 1850
rect 4301 1848 4354 1862
rect 4302 1846 4366 1848
rect 4409 1846 4424 1862
rect 4473 1859 4503 1862
rect 4473 1856 4509 1859
rect 4439 1848 4455 1850
rect 4213 1836 4228 1840
rect 4131 1834 4228 1836
rect 4256 1834 4424 1846
rect 4440 1836 4455 1840
rect 4473 1837 4512 1856
rect 4531 1850 4538 1851
rect 4537 1843 4538 1850
rect 4521 1840 4522 1843
rect 4537 1840 4550 1843
rect 4473 1836 4503 1837
rect 4512 1836 4518 1837
rect 4521 1836 4550 1840
rect 4440 1835 4550 1836
rect 4440 1834 4556 1835
rect 4115 1826 4166 1834
rect 4115 1814 4140 1826
rect 4147 1814 4166 1826
rect 4197 1826 4247 1834
rect 4197 1818 4213 1826
rect 4220 1824 4247 1826
rect 4256 1824 4477 1834
rect 4220 1814 4477 1824
rect 4506 1826 4556 1834
rect 4506 1817 4522 1826
rect 4115 1806 4166 1814
rect 4213 1806 4477 1814
rect 4503 1814 4522 1817
rect 4529 1814 4556 1826
rect 4503 1806 4556 1814
rect 4131 1798 4132 1806
rect 4147 1798 4160 1806
rect 4131 1790 4147 1798
rect 4128 1783 4147 1786
rect 4128 1774 4150 1783
rect 4101 1764 4150 1774
rect 4101 1758 4131 1764
rect 4150 1759 4155 1764
rect 4073 1742 4147 1758
rect 4165 1750 4195 1806
rect 4230 1796 4438 1806
rect 4473 1802 4518 1806
rect 4521 1805 4522 1806
rect 4537 1805 4550 1806
rect 4256 1766 4445 1796
rect 4271 1763 4445 1766
rect 4264 1760 4445 1763
rect 4073 1740 4086 1742
rect 4101 1740 4135 1742
rect 4073 1724 4147 1740
rect 4174 1736 4187 1750
rect 4202 1736 4218 1752
rect 4264 1747 4275 1760
rect 4057 1702 4058 1718
rect 4073 1702 4086 1724
rect 4101 1702 4131 1724
rect 4174 1720 4236 1736
rect 4264 1729 4275 1745
rect 4280 1740 4290 1760
rect 4300 1740 4314 1760
rect 4317 1747 4326 1760
rect 4342 1747 4351 1760
rect 4280 1729 4314 1740
rect 4317 1729 4326 1745
rect 4342 1729 4351 1745
rect 4358 1740 4368 1760
rect 4378 1740 4392 1760
rect 4393 1747 4404 1760
rect 4358 1729 4392 1740
rect 4393 1729 4404 1745
rect 4450 1736 4466 1752
rect 4473 1750 4503 1802
rect 4537 1798 4538 1805
rect 4522 1790 4538 1798
rect 4509 1758 4522 1777
rect 4537 1758 4567 1774
rect 4509 1742 4583 1758
rect 4509 1740 4522 1742
rect 4537 1740 4571 1742
rect 4174 1718 4187 1720
rect 4202 1718 4236 1720
rect 4174 1702 4236 1718
rect 4280 1713 4296 1716
rect 4358 1713 4388 1724
rect 4436 1720 4482 1736
rect 4509 1724 4583 1740
rect 4436 1718 4470 1720
rect 4435 1702 4482 1718
rect 4509 1702 4522 1724
rect 4537 1702 4567 1724
rect 4594 1702 4595 1718
rect 4610 1702 4623 1862
rect 4751 1758 4764 1862
rect 4809 1840 4810 1850
rect 4825 1840 4838 1850
rect 4809 1836 4838 1840
rect 4843 1836 4873 1862
rect 4891 1848 4907 1850
rect 4979 1848 5032 1862
rect 4980 1846 5044 1848
rect 5087 1846 5102 1862
rect 5151 1859 5181 1862
rect 5151 1856 5187 1859
rect 5117 1848 5133 1850
rect 4891 1836 4906 1840
rect 4809 1834 4906 1836
rect 4934 1834 5102 1846
rect 5118 1836 5133 1840
rect 5151 1837 5190 1856
rect 5209 1850 5216 1851
rect 5215 1843 5216 1850
rect 5199 1840 5200 1843
rect 5215 1840 5228 1843
rect 5151 1836 5181 1837
rect 5190 1836 5196 1837
rect 5199 1836 5228 1840
rect 5118 1835 5228 1836
rect 5118 1834 5234 1835
rect 4793 1826 4844 1834
rect 4793 1814 4818 1826
rect 4825 1814 4844 1826
rect 4875 1826 4925 1834
rect 4875 1818 4891 1826
rect 4898 1824 4925 1826
rect 4934 1824 5155 1834
rect 4898 1814 5155 1824
rect 5184 1826 5234 1834
rect 5184 1817 5200 1826
rect 4793 1806 4844 1814
rect 4891 1806 5155 1814
rect 5181 1814 5200 1817
rect 5207 1814 5234 1826
rect 5181 1806 5234 1814
rect 4809 1798 4810 1806
rect 4825 1798 4838 1806
rect 4809 1790 4825 1798
rect 4806 1783 4825 1786
rect 4806 1774 4828 1783
rect 4779 1764 4828 1774
rect 4779 1758 4809 1764
rect 4828 1759 4833 1764
rect 4751 1742 4825 1758
rect 4843 1750 4873 1806
rect 4908 1796 5116 1806
rect 5151 1802 5196 1806
rect 5199 1805 5200 1806
rect 5215 1805 5228 1806
rect 4934 1766 5123 1796
rect 4949 1763 5123 1766
rect 4942 1760 5123 1763
rect 4751 1740 4764 1742
rect 4779 1740 4813 1742
rect 4751 1724 4825 1740
rect 4852 1736 4865 1750
rect 4880 1736 4896 1752
rect 4942 1747 4953 1760
rect 4735 1702 4736 1718
rect 4751 1702 4764 1724
rect 4779 1702 4809 1724
rect 4852 1720 4914 1736
rect 4942 1729 4953 1745
rect 4958 1740 4968 1760
rect 4978 1740 4992 1760
rect 4995 1747 5004 1760
rect 5020 1747 5029 1760
rect 4958 1729 4992 1740
rect 4995 1729 5004 1745
rect 5020 1729 5029 1745
rect 5036 1740 5046 1760
rect 5056 1740 5070 1760
rect 5071 1747 5082 1760
rect 5036 1729 5070 1740
rect 5071 1729 5082 1745
rect 5128 1736 5144 1752
rect 5151 1750 5181 1802
rect 5215 1798 5216 1805
rect 5200 1790 5216 1798
rect 5187 1758 5200 1777
rect 5215 1758 5245 1774
rect 5187 1742 5261 1758
rect 5187 1740 5200 1742
rect 5215 1740 5249 1742
rect 4852 1718 4865 1720
rect 4880 1718 4914 1720
rect 4852 1702 4914 1718
rect 4958 1713 4974 1716
rect 5036 1713 5066 1724
rect 5114 1720 5160 1736
rect 5187 1724 5261 1740
rect 5114 1718 5148 1720
rect 5113 1702 5160 1718
rect 5187 1702 5200 1724
rect 5215 1702 5245 1724
rect 5272 1702 5273 1718
rect 5288 1702 5301 1862
rect 5331 1758 5344 1862
rect 5389 1840 5390 1850
rect 5405 1840 5418 1850
rect 5389 1836 5418 1840
rect 5423 1836 5453 1862
rect 5471 1848 5487 1850
rect 5559 1848 5612 1862
rect 5560 1846 5624 1848
rect 5667 1846 5682 1862
rect 5731 1859 5761 1862
rect 5731 1856 5767 1859
rect 5697 1848 5713 1850
rect 5471 1836 5486 1840
rect 5389 1834 5486 1836
rect 5514 1834 5682 1846
rect 5698 1836 5713 1840
rect 5731 1837 5770 1856
rect 5789 1850 5796 1851
rect 5795 1843 5796 1850
rect 5779 1840 5780 1843
rect 5795 1840 5808 1843
rect 5731 1836 5761 1837
rect 5770 1836 5776 1837
rect 5779 1836 5808 1840
rect 5698 1835 5808 1836
rect 5698 1834 5814 1835
rect 5373 1826 5424 1834
rect 5373 1814 5398 1826
rect 5405 1814 5424 1826
rect 5455 1826 5505 1834
rect 5455 1818 5471 1826
rect 5478 1824 5505 1826
rect 5514 1824 5735 1834
rect 5478 1814 5735 1824
rect 5764 1826 5814 1834
rect 5764 1817 5780 1826
rect 5373 1806 5424 1814
rect 5471 1806 5735 1814
rect 5761 1814 5780 1817
rect 5787 1814 5814 1826
rect 5761 1806 5814 1814
rect 5389 1798 5390 1806
rect 5405 1798 5418 1806
rect 5389 1790 5405 1798
rect 5386 1783 5405 1786
rect 5386 1774 5408 1783
rect 5359 1764 5408 1774
rect 5359 1758 5389 1764
rect 5408 1759 5413 1764
rect 5331 1742 5405 1758
rect 5423 1750 5453 1806
rect 5488 1796 5696 1806
rect 5731 1802 5776 1806
rect 5779 1805 5780 1806
rect 5795 1805 5808 1806
rect 5514 1766 5703 1796
rect 5529 1763 5703 1766
rect 5522 1760 5703 1763
rect 5331 1740 5344 1742
rect 5359 1740 5393 1742
rect 5331 1724 5405 1740
rect 5432 1736 5445 1750
rect 5460 1736 5476 1752
rect 5522 1747 5533 1760
rect 5315 1702 5316 1718
rect 5331 1702 5344 1724
rect 5359 1702 5389 1724
rect 5432 1720 5494 1736
rect 5522 1729 5533 1745
rect 5538 1740 5548 1760
rect 5558 1740 5572 1760
rect 5575 1747 5584 1760
rect 5600 1747 5609 1760
rect 5538 1729 5572 1740
rect 5575 1729 5584 1745
rect 5600 1729 5609 1745
rect 5616 1740 5626 1760
rect 5636 1740 5650 1760
rect 5651 1747 5662 1760
rect 5616 1729 5650 1740
rect 5651 1729 5662 1745
rect 5708 1736 5724 1752
rect 5731 1750 5761 1802
rect 5795 1798 5796 1805
rect 5780 1790 5796 1798
rect 5767 1758 5780 1777
rect 5795 1758 5825 1774
rect 5767 1742 5841 1758
rect 5767 1740 5780 1742
rect 5795 1740 5829 1742
rect 5432 1718 5445 1720
rect 5460 1718 5494 1720
rect 5432 1702 5494 1718
rect 5538 1713 5554 1716
rect 5616 1713 5646 1724
rect 5694 1720 5740 1736
rect 5767 1724 5841 1740
rect 5694 1718 5728 1720
rect 5693 1702 5740 1718
rect 5767 1702 5780 1724
rect 5795 1702 5825 1724
rect 5852 1702 5853 1718
rect 5868 1702 5881 1862
rect 3471 1694 3512 1702
rect 3471 1668 3486 1694
rect 3493 1668 3512 1694
rect 3576 1690 3638 1702
rect 3650 1690 3725 1702
rect 3783 1690 3858 1702
rect 3870 1690 3901 1702
rect 3907 1690 3942 1702
rect 3576 1688 3738 1690
rect 3471 1660 3512 1668
rect 3594 1664 3607 1688
rect 3622 1686 3637 1688
rect 3477 1650 3478 1660
rect 3493 1650 3506 1660
rect 3521 1650 3551 1664
rect 3594 1650 3637 1664
rect 3661 1661 3668 1668
rect 3671 1664 3738 1688
rect 3770 1688 3942 1690
rect 3740 1666 3768 1670
rect 3770 1666 3850 1688
rect 3871 1686 3886 1688
rect 3740 1664 3850 1666
rect 3671 1660 3850 1664
rect 3644 1650 3674 1660
rect 3676 1650 3829 1660
rect 3837 1650 3867 1660
rect 3871 1650 3901 1664
rect 3929 1650 3942 1688
rect 4014 1694 4049 1702
rect 4014 1668 4015 1694
rect 4022 1668 4049 1694
rect 3957 1650 3987 1664
rect 4014 1660 4049 1668
rect 4051 1694 4092 1702
rect 4051 1668 4066 1694
rect 4073 1668 4092 1694
rect 4156 1690 4218 1702
rect 4230 1690 4305 1702
rect 4363 1690 4438 1702
rect 4450 1690 4481 1702
rect 4487 1690 4522 1702
rect 4156 1688 4318 1690
rect 4051 1660 4092 1668
rect 4174 1664 4187 1688
rect 4202 1686 4217 1688
rect 4014 1650 4015 1660
rect 4030 1650 4043 1660
rect 4057 1650 4058 1660
rect 4073 1650 4086 1660
rect 4101 1650 4131 1664
rect 4174 1650 4217 1664
rect 4241 1661 4248 1668
rect 4251 1664 4318 1688
rect 4350 1688 4522 1690
rect 4320 1666 4348 1670
rect 4350 1666 4430 1688
rect 4451 1686 4466 1688
rect 4320 1664 4430 1666
rect 4251 1660 4430 1664
rect 4224 1650 4254 1660
rect 4256 1650 4409 1660
rect 4417 1650 4447 1660
rect 4451 1650 4481 1664
rect 4509 1650 4522 1688
rect 4594 1694 4629 1702
rect 4594 1668 4595 1694
rect 4602 1668 4629 1694
rect 4537 1650 4567 1664
rect 4594 1660 4629 1668
rect 4729 1694 4770 1702
rect 4729 1668 4744 1694
rect 4751 1668 4770 1694
rect 4834 1690 4896 1702
rect 4908 1690 4983 1702
rect 5041 1690 5116 1702
rect 5128 1690 5159 1702
rect 5165 1690 5200 1702
rect 4834 1688 4996 1690
rect 4729 1660 4770 1668
rect 4852 1664 4865 1688
rect 4880 1686 4895 1688
rect 4594 1650 4595 1660
rect 4610 1650 4623 1660
rect 3469 1636 4623 1650
rect 4735 1650 4736 1660
rect 4751 1650 4764 1660
rect 4779 1650 4809 1664
rect 4852 1650 4895 1664
rect 4919 1661 4926 1668
rect 4929 1664 4996 1688
rect 5028 1688 5200 1690
rect 4998 1666 5026 1670
rect 5028 1666 5108 1688
rect 5129 1686 5144 1688
rect 4998 1664 5108 1666
rect 4929 1660 5108 1664
rect 4902 1650 4932 1660
rect 4934 1650 5087 1660
rect 5095 1650 5125 1660
rect 5129 1650 5159 1664
rect 5187 1650 5200 1688
rect 5272 1694 5307 1702
rect 5272 1668 5273 1694
rect 5280 1668 5307 1694
rect 5215 1650 5245 1664
rect 5272 1660 5307 1668
rect 5309 1694 5350 1702
rect 5309 1668 5324 1694
rect 5331 1668 5350 1694
rect 5414 1690 5476 1702
rect 5488 1690 5563 1702
rect 5621 1690 5696 1702
rect 5708 1690 5739 1702
rect 5745 1690 5780 1702
rect 5414 1688 5576 1690
rect 5309 1660 5350 1668
rect 5432 1664 5445 1688
rect 5460 1686 5475 1688
rect 5272 1650 5273 1660
rect 5288 1650 5301 1660
rect 5315 1650 5316 1660
rect 5331 1650 5344 1660
rect 5359 1650 5389 1664
rect 5432 1650 5475 1664
rect 5499 1661 5506 1668
rect 5509 1664 5576 1688
rect 5608 1688 5780 1690
rect 5578 1666 5606 1670
rect 5608 1666 5688 1688
rect 5709 1686 5724 1688
rect 5578 1664 5688 1666
rect 5509 1660 5688 1664
rect 5482 1650 5512 1660
rect 5514 1650 5667 1660
rect 5675 1650 5705 1660
rect 5709 1650 5739 1664
rect 5767 1650 5780 1688
rect 5852 1694 5887 1702
rect 5852 1668 5853 1694
rect 5860 1668 5887 1694
rect 5795 1650 5825 1664
rect 5852 1660 5887 1668
rect 5852 1650 5853 1660
rect 5868 1650 5881 1660
rect 4735 1644 5889 1650
rect 4736 1636 5889 1644
rect 3493 1606 3506 1636
rect 3521 1618 3551 1636
rect 3594 1622 3608 1636
rect 3644 1622 3864 1636
rect 3595 1620 3608 1622
rect 3561 1608 3576 1620
rect 3558 1606 3580 1608
rect 3585 1606 3615 1620
rect 3676 1618 3829 1622
rect 3658 1606 3850 1618
rect 3893 1606 3923 1620
rect 3929 1606 3942 1636
rect 3957 1618 3987 1636
rect 4030 1606 4043 1636
rect 4073 1606 4086 1636
rect 4101 1618 4131 1636
rect 4174 1622 4188 1636
rect 4224 1622 4444 1636
rect 4175 1620 4188 1622
rect 4141 1608 4156 1620
rect 4138 1606 4160 1608
rect 4165 1606 4195 1620
rect 4256 1618 4409 1622
rect 4238 1606 4430 1618
rect 4473 1606 4503 1620
rect 4509 1606 4522 1636
rect 4537 1618 4567 1636
rect 4610 1606 4623 1636
rect 4751 1606 4764 1636
rect 4779 1618 4809 1636
rect 4852 1622 4866 1636
rect 4902 1622 5122 1636
rect 4853 1620 4866 1622
rect 4819 1608 4834 1620
rect 4816 1606 4838 1608
rect 4843 1606 4873 1620
rect 4934 1618 5087 1622
rect 4916 1606 5108 1618
rect 5151 1606 5181 1620
rect 5187 1606 5200 1636
rect 5215 1618 5245 1636
rect 5288 1606 5301 1636
rect 5331 1606 5344 1636
rect 5359 1618 5389 1636
rect 5432 1622 5446 1636
rect 5482 1622 5702 1636
rect 5433 1620 5446 1622
rect 5399 1608 5414 1620
rect 5396 1606 5418 1608
rect 5423 1606 5453 1620
rect 5514 1618 5667 1622
rect 5496 1606 5688 1618
rect 5731 1606 5761 1620
rect 5767 1606 5780 1636
rect 5795 1618 5825 1636
rect 5868 1606 5881 1636
rect 3469 1592 4623 1606
rect 4736 1592 5889 1606
rect 3493 1488 3506 1592
rect 3551 1570 3552 1580
rect 3567 1570 3580 1580
rect 3551 1566 3580 1570
rect 3585 1566 3615 1592
rect 3633 1578 3649 1580
rect 3721 1578 3774 1592
rect 3722 1576 3786 1578
rect 3829 1576 3844 1592
rect 3893 1589 3923 1592
rect 3893 1586 3929 1589
rect 3859 1578 3875 1580
rect 3633 1566 3648 1570
rect 3551 1564 3648 1566
rect 3676 1564 3844 1576
rect 3860 1566 3875 1570
rect 3893 1567 3932 1586
rect 3951 1580 3958 1581
rect 3957 1573 3958 1580
rect 3941 1570 3942 1573
rect 3957 1570 3970 1573
rect 3893 1566 3923 1567
rect 3932 1566 3938 1567
rect 3941 1566 3970 1570
rect 3860 1565 3970 1566
rect 3860 1564 3976 1565
rect 3535 1556 3586 1564
rect 3535 1544 3560 1556
rect 3567 1544 3586 1556
rect 3617 1556 3667 1564
rect 3617 1548 3633 1556
rect 3640 1554 3667 1556
rect 3676 1554 3897 1564
rect 3640 1544 3897 1554
rect 3926 1556 3976 1564
rect 3926 1547 3942 1556
rect 3535 1536 3586 1544
rect 3633 1536 3897 1544
rect 3923 1544 3942 1547
rect 3949 1544 3976 1556
rect 3923 1536 3976 1544
rect 3551 1528 3552 1536
rect 3567 1528 3580 1536
rect 3551 1520 3567 1528
rect 3548 1513 3567 1516
rect 3548 1504 3570 1513
rect 3521 1494 3570 1504
rect 3521 1488 3551 1494
rect 3570 1489 3575 1494
rect 3493 1472 3567 1488
rect 3585 1480 3615 1536
rect 3650 1526 3858 1536
rect 3893 1532 3938 1536
rect 3941 1535 3942 1536
rect 3957 1535 3970 1536
rect 3676 1496 3865 1526
rect 3691 1493 3865 1496
rect 3684 1490 3865 1493
rect 3493 1470 3506 1472
rect 3521 1470 3555 1472
rect 3493 1454 3567 1470
rect 3594 1466 3607 1480
rect 3622 1466 3638 1482
rect 3684 1477 3695 1490
rect 3477 1432 3478 1448
rect 3493 1432 3506 1454
rect 3521 1432 3551 1454
rect 3594 1450 3656 1466
rect 3684 1459 3695 1475
rect 3700 1470 3710 1490
rect 3720 1470 3734 1490
rect 3737 1477 3746 1490
rect 3762 1477 3771 1490
rect 3700 1459 3734 1470
rect 3737 1459 3746 1475
rect 3762 1459 3771 1475
rect 3778 1470 3788 1490
rect 3798 1470 3812 1490
rect 3813 1477 3824 1490
rect 3778 1459 3812 1470
rect 3813 1459 3824 1475
rect 3870 1466 3886 1482
rect 3893 1480 3923 1532
rect 3957 1528 3958 1535
rect 3942 1520 3958 1528
rect 3929 1488 3942 1507
rect 3957 1488 3987 1504
rect 3929 1472 4003 1488
rect 3929 1470 3942 1472
rect 3957 1470 3991 1472
rect 3594 1448 3607 1450
rect 3622 1448 3656 1450
rect 3594 1432 3656 1448
rect 3700 1443 3716 1446
rect 3778 1443 3808 1454
rect 3856 1450 3902 1466
rect 3929 1454 4003 1470
rect 3856 1448 3890 1450
rect 3855 1432 3902 1448
rect 3929 1432 3942 1454
rect 3957 1432 3987 1454
rect 4014 1432 4015 1448
rect 4030 1432 4043 1592
rect 4073 1488 4086 1592
rect 4131 1570 4132 1580
rect 4147 1570 4160 1580
rect 4131 1566 4160 1570
rect 4165 1566 4195 1592
rect 4213 1578 4229 1580
rect 4301 1578 4354 1592
rect 4302 1576 4366 1578
rect 4409 1576 4424 1592
rect 4473 1589 4503 1592
rect 4473 1586 4509 1589
rect 4439 1578 4455 1580
rect 4213 1566 4228 1570
rect 4131 1564 4228 1566
rect 4256 1564 4424 1576
rect 4440 1566 4455 1570
rect 4473 1567 4512 1586
rect 4531 1580 4538 1581
rect 4537 1573 4538 1580
rect 4521 1570 4522 1573
rect 4537 1570 4550 1573
rect 4473 1566 4503 1567
rect 4512 1566 4518 1567
rect 4521 1566 4550 1570
rect 4440 1565 4550 1566
rect 4440 1564 4556 1565
rect 4115 1556 4166 1564
rect 4115 1544 4140 1556
rect 4147 1544 4166 1556
rect 4197 1556 4247 1564
rect 4197 1548 4213 1556
rect 4220 1554 4247 1556
rect 4256 1554 4477 1564
rect 4220 1544 4477 1554
rect 4506 1556 4556 1564
rect 4506 1547 4522 1556
rect 4115 1536 4166 1544
rect 4213 1536 4477 1544
rect 4503 1544 4522 1547
rect 4529 1544 4556 1556
rect 4503 1536 4556 1544
rect 4131 1528 4132 1536
rect 4147 1528 4160 1536
rect 4131 1520 4147 1528
rect 4128 1513 4147 1516
rect 4128 1504 4150 1513
rect 4101 1494 4150 1504
rect 4101 1488 4131 1494
rect 4150 1489 4155 1494
rect 4073 1472 4147 1488
rect 4165 1480 4195 1536
rect 4230 1526 4438 1536
rect 4473 1532 4518 1536
rect 4521 1535 4522 1536
rect 4537 1535 4550 1536
rect 4256 1496 4445 1526
rect 4271 1493 4445 1496
rect 4264 1490 4445 1493
rect 4073 1470 4086 1472
rect 4101 1470 4135 1472
rect 4073 1454 4147 1470
rect 4174 1466 4187 1480
rect 4202 1466 4218 1482
rect 4264 1477 4275 1490
rect 4057 1432 4058 1448
rect 4073 1432 4086 1454
rect 4101 1432 4131 1454
rect 4174 1450 4236 1466
rect 4264 1459 4275 1475
rect 4280 1470 4290 1490
rect 4300 1470 4314 1490
rect 4317 1477 4326 1490
rect 4342 1477 4351 1490
rect 4280 1459 4314 1470
rect 4317 1459 4326 1475
rect 4342 1459 4351 1475
rect 4358 1470 4368 1490
rect 4378 1470 4392 1490
rect 4393 1477 4404 1490
rect 4358 1459 4392 1470
rect 4393 1459 4404 1475
rect 4450 1466 4466 1482
rect 4473 1480 4503 1532
rect 4537 1528 4538 1535
rect 4522 1520 4538 1528
rect 4509 1488 4522 1507
rect 4537 1488 4567 1504
rect 4509 1472 4583 1488
rect 4509 1470 4522 1472
rect 4537 1470 4571 1472
rect 4174 1448 4187 1450
rect 4202 1448 4236 1450
rect 4174 1432 4236 1448
rect 4280 1443 4296 1446
rect 4358 1443 4388 1454
rect 4436 1450 4482 1466
rect 4509 1454 4583 1470
rect 4436 1448 4470 1450
rect 4435 1432 4482 1448
rect 4509 1432 4522 1454
rect 4537 1432 4567 1454
rect 4594 1432 4595 1448
rect 4610 1432 4623 1592
rect 4751 1488 4764 1592
rect 4809 1570 4810 1580
rect 4825 1570 4838 1580
rect 4809 1566 4838 1570
rect 4843 1566 4873 1592
rect 4891 1578 4907 1580
rect 4979 1578 5032 1592
rect 4980 1576 5044 1578
rect 5087 1576 5102 1592
rect 5151 1589 5181 1592
rect 5151 1586 5187 1589
rect 5117 1578 5133 1580
rect 4891 1566 4906 1570
rect 4809 1564 4906 1566
rect 4934 1564 5102 1576
rect 5118 1566 5133 1570
rect 5151 1567 5190 1586
rect 5209 1580 5216 1581
rect 5215 1573 5216 1580
rect 5199 1570 5200 1573
rect 5215 1570 5228 1573
rect 5151 1566 5181 1567
rect 5190 1566 5196 1567
rect 5199 1566 5228 1570
rect 5118 1565 5228 1566
rect 5118 1564 5234 1565
rect 4793 1556 4844 1564
rect 4793 1544 4818 1556
rect 4825 1544 4844 1556
rect 4875 1556 4925 1564
rect 4875 1548 4891 1556
rect 4898 1554 4925 1556
rect 4934 1554 5155 1564
rect 4898 1544 5155 1554
rect 5184 1556 5234 1564
rect 5184 1547 5200 1556
rect 4793 1536 4844 1544
rect 4891 1536 5155 1544
rect 5181 1544 5200 1547
rect 5207 1544 5234 1556
rect 5181 1536 5234 1544
rect 4809 1528 4810 1536
rect 4825 1528 4838 1536
rect 4809 1520 4825 1528
rect 4806 1513 4825 1516
rect 4806 1504 4828 1513
rect 4779 1494 4828 1504
rect 4779 1488 4809 1494
rect 4828 1489 4833 1494
rect 4751 1472 4825 1488
rect 4843 1480 4873 1536
rect 4908 1526 5116 1536
rect 5151 1532 5196 1536
rect 5199 1535 5200 1536
rect 5215 1535 5228 1536
rect 4934 1496 5123 1526
rect 4949 1493 5123 1496
rect 4942 1490 5123 1493
rect 4751 1470 4764 1472
rect 4779 1470 4813 1472
rect 4751 1454 4825 1470
rect 4852 1466 4865 1480
rect 4880 1466 4896 1482
rect 4942 1477 4953 1490
rect 4735 1432 4736 1448
rect 4751 1432 4764 1454
rect 4779 1432 4809 1454
rect 4852 1450 4914 1466
rect 4942 1459 4953 1475
rect 4958 1470 4968 1490
rect 4978 1470 4992 1490
rect 4995 1477 5004 1490
rect 5020 1477 5029 1490
rect 4958 1459 4992 1470
rect 4995 1459 5004 1475
rect 5020 1459 5029 1475
rect 5036 1470 5046 1490
rect 5056 1470 5070 1490
rect 5071 1477 5082 1490
rect 5036 1459 5070 1470
rect 5071 1459 5082 1475
rect 5128 1466 5144 1482
rect 5151 1480 5181 1532
rect 5215 1528 5216 1535
rect 5200 1520 5216 1528
rect 5187 1488 5200 1507
rect 5215 1488 5245 1504
rect 5187 1472 5261 1488
rect 5187 1470 5200 1472
rect 5215 1470 5249 1472
rect 4852 1448 4865 1450
rect 4880 1448 4914 1450
rect 4852 1432 4914 1448
rect 4958 1443 4974 1446
rect 5036 1443 5066 1454
rect 5114 1450 5160 1466
rect 5187 1454 5261 1470
rect 5114 1448 5148 1450
rect 5113 1432 5160 1448
rect 5187 1432 5200 1454
rect 5215 1432 5245 1454
rect 5272 1432 5273 1448
rect 5288 1432 5301 1592
rect 5331 1488 5344 1592
rect 5389 1570 5390 1580
rect 5405 1570 5418 1580
rect 5389 1566 5418 1570
rect 5423 1566 5453 1592
rect 5471 1578 5487 1580
rect 5559 1578 5612 1592
rect 5560 1576 5624 1578
rect 5667 1576 5682 1592
rect 5731 1589 5761 1592
rect 5731 1586 5767 1589
rect 5697 1578 5713 1580
rect 5471 1566 5486 1570
rect 5389 1564 5486 1566
rect 5514 1564 5682 1576
rect 5698 1566 5713 1570
rect 5731 1567 5770 1586
rect 5789 1580 5796 1581
rect 5795 1573 5796 1580
rect 5779 1570 5780 1573
rect 5795 1570 5808 1573
rect 5731 1566 5761 1567
rect 5770 1566 5776 1567
rect 5779 1566 5808 1570
rect 5698 1565 5808 1566
rect 5698 1564 5814 1565
rect 5373 1556 5424 1564
rect 5373 1544 5398 1556
rect 5405 1544 5424 1556
rect 5455 1556 5505 1564
rect 5455 1548 5471 1556
rect 5478 1554 5505 1556
rect 5514 1554 5735 1564
rect 5478 1544 5735 1554
rect 5764 1556 5814 1564
rect 5764 1547 5780 1556
rect 5373 1536 5424 1544
rect 5471 1536 5735 1544
rect 5761 1544 5780 1547
rect 5787 1544 5814 1556
rect 5761 1536 5814 1544
rect 5389 1528 5390 1536
rect 5405 1528 5418 1536
rect 5389 1520 5405 1528
rect 5386 1513 5405 1516
rect 5386 1504 5408 1513
rect 5359 1494 5408 1504
rect 5359 1488 5389 1494
rect 5408 1489 5413 1494
rect 5331 1472 5405 1488
rect 5423 1480 5453 1536
rect 5488 1526 5696 1536
rect 5731 1532 5776 1536
rect 5779 1535 5780 1536
rect 5795 1535 5808 1536
rect 5514 1496 5703 1526
rect 5529 1493 5703 1496
rect 5522 1490 5703 1493
rect 5331 1470 5344 1472
rect 5359 1470 5393 1472
rect 5331 1454 5405 1470
rect 5432 1466 5445 1480
rect 5460 1466 5476 1482
rect 5522 1477 5533 1490
rect 5315 1432 5316 1448
rect 5331 1432 5344 1454
rect 5359 1432 5389 1454
rect 5432 1450 5494 1466
rect 5522 1459 5533 1475
rect 5538 1470 5548 1490
rect 5558 1470 5572 1490
rect 5575 1477 5584 1490
rect 5600 1477 5609 1490
rect 5538 1459 5572 1470
rect 5575 1459 5584 1475
rect 5600 1459 5609 1475
rect 5616 1470 5626 1490
rect 5636 1470 5650 1490
rect 5651 1477 5662 1490
rect 5616 1459 5650 1470
rect 5651 1459 5662 1475
rect 5708 1466 5724 1482
rect 5731 1480 5761 1532
rect 5795 1528 5796 1535
rect 5780 1520 5796 1528
rect 5767 1488 5780 1507
rect 5795 1488 5825 1504
rect 5767 1472 5841 1488
rect 5767 1470 5780 1472
rect 5795 1470 5829 1472
rect 5432 1448 5445 1450
rect 5460 1448 5494 1450
rect 5432 1432 5494 1448
rect 5538 1443 5554 1446
rect 5616 1443 5646 1454
rect 5694 1450 5740 1466
rect 5767 1454 5841 1470
rect 5694 1448 5728 1450
rect 5693 1432 5740 1448
rect 5767 1432 5780 1454
rect 5795 1432 5825 1454
rect 5852 1432 5853 1448
rect 5868 1432 5881 1592
rect 3471 1424 3512 1432
rect 3471 1398 3486 1424
rect 3493 1398 3512 1424
rect 3576 1420 3638 1432
rect 3650 1420 3725 1432
rect 3783 1420 3858 1432
rect 3870 1420 3901 1432
rect 3907 1420 3942 1432
rect 3576 1418 3738 1420
rect 3471 1390 3512 1398
rect 3594 1394 3607 1418
rect 3622 1416 3637 1418
rect 3477 1380 3478 1390
rect 3493 1380 3506 1390
rect 3521 1380 3551 1394
rect 3594 1380 3637 1394
rect 3661 1391 3668 1398
rect 3671 1394 3738 1418
rect 3770 1418 3942 1420
rect 3740 1396 3768 1400
rect 3770 1396 3850 1418
rect 3871 1416 3886 1418
rect 3740 1394 3850 1396
rect 3671 1390 3850 1394
rect 3644 1380 3674 1390
rect 3676 1380 3829 1390
rect 3837 1380 3867 1390
rect 3871 1380 3901 1394
rect 3929 1380 3942 1418
rect 4014 1424 4049 1432
rect 4014 1398 4015 1424
rect 4022 1398 4049 1424
rect 3957 1380 3987 1394
rect 4014 1390 4049 1398
rect 4051 1424 4092 1432
rect 4051 1398 4066 1424
rect 4073 1398 4092 1424
rect 4156 1420 4218 1432
rect 4230 1420 4305 1432
rect 4363 1420 4438 1432
rect 4450 1420 4481 1432
rect 4487 1420 4522 1432
rect 4156 1418 4318 1420
rect 4051 1390 4092 1398
rect 4174 1394 4187 1418
rect 4202 1416 4217 1418
rect 4014 1380 4015 1390
rect 4030 1380 4043 1390
rect 4057 1380 4058 1390
rect 4073 1380 4086 1390
rect 4101 1380 4131 1394
rect 4174 1380 4217 1394
rect 4241 1391 4248 1398
rect 4251 1394 4318 1418
rect 4350 1418 4522 1420
rect 4320 1396 4348 1400
rect 4350 1396 4430 1418
rect 4451 1416 4466 1418
rect 4320 1394 4430 1396
rect 4251 1390 4430 1394
rect 4224 1380 4254 1390
rect 4256 1380 4409 1390
rect 4417 1380 4447 1390
rect 4451 1380 4481 1394
rect 4509 1380 4522 1418
rect 4594 1424 4629 1432
rect 4594 1398 4595 1424
rect 4602 1398 4629 1424
rect 4537 1380 4567 1394
rect 4594 1390 4629 1398
rect 4729 1424 4770 1432
rect 4729 1398 4744 1424
rect 4751 1398 4770 1424
rect 4834 1420 4896 1432
rect 4908 1420 4983 1432
rect 5041 1420 5116 1432
rect 5128 1420 5159 1432
rect 5165 1420 5200 1432
rect 4834 1418 4996 1420
rect 4729 1390 4770 1398
rect 4852 1394 4865 1418
rect 4880 1416 4895 1418
rect 4594 1380 4595 1390
rect 4610 1380 4623 1390
rect 3469 1366 4623 1380
rect 4735 1380 4736 1390
rect 4751 1380 4764 1390
rect 4779 1380 4809 1394
rect 4852 1380 4895 1394
rect 4919 1391 4926 1398
rect 4929 1394 4996 1418
rect 5028 1418 5200 1420
rect 4998 1396 5026 1400
rect 5028 1396 5108 1418
rect 5129 1416 5144 1418
rect 4998 1394 5108 1396
rect 4929 1390 5108 1394
rect 4902 1380 4932 1390
rect 4934 1380 5087 1390
rect 5095 1380 5125 1390
rect 5129 1380 5159 1394
rect 5187 1380 5200 1418
rect 5272 1424 5307 1432
rect 5272 1398 5273 1424
rect 5280 1398 5307 1424
rect 5215 1380 5245 1394
rect 5272 1390 5307 1398
rect 5309 1424 5350 1432
rect 5309 1398 5324 1424
rect 5331 1398 5350 1424
rect 5414 1420 5476 1432
rect 5488 1420 5563 1432
rect 5621 1420 5696 1432
rect 5708 1420 5739 1432
rect 5745 1420 5780 1432
rect 5414 1418 5576 1420
rect 5309 1390 5350 1398
rect 5432 1394 5445 1418
rect 5460 1416 5475 1418
rect 5272 1380 5273 1390
rect 5288 1380 5301 1390
rect 5315 1380 5316 1390
rect 5331 1380 5344 1390
rect 5359 1380 5389 1394
rect 5432 1380 5475 1394
rect 5499 1391 5506 1398
rect 5509 1394 5576 1418
rect 5608 1418 5780 1420
rect 5578 1396 5606 1400
rect 5608 1396 5688 1418
rect 5709 1416 5724 1418
rect 5578 1394 5688 1396
rect 5509 1390 5688 1394
rect 5482 1380 5512 1390
rect 5514 1380 5667 1390
rect 5675 1380 5705 1390
rect 5709 1380 5739 1394
rect 5767 1380 5780 1418
rect 5852 1424 5887 1432
rect 5852 1398 5853 1424
rect 5860 1398 5887 1424
rect 5795 1380 5825 1394
rect 5852 1390 5887 1398
rect 5852 1380 5853 1390
rect 5868 1380 5881 1390
rect 4735 1374 5889 1380
rect 4736 1366 5889 1374
rect 3493 1336 3506 1366
rect 3521 1348 3551 1366
rect 3594 1352 3608 1366
rect 3644 1352 3864 1366
rect 3595 1350 3608 1352
rect 3561 1338 3576 1350
rect 3558 1336 3580 1338
rect 3585 1336 3615 1350
rect 3676 1348 3829 1352
rect 3658 1336 3850 1348
rect 3893 1336 3923 1350
rect 3929 1336 3942 1366
rect 3957 1348 3987 1366
rect 4030 1336 4043 1366
rect 4073 1336 4086 1366
rect 4101 1348 4131 1366
rect 4174 1352 4188 1366
rect 4224 1352 4444 1366
rect 4175 1350 4188 1352
rect 4141 1338 4156 1350
rect 4138 1336 4160 1338
rect 4165 1336 4195 1350
rect 4256 1348 4409 1352
rect 4238 1336 4430 1348
rect 4473 1336 4503 1350
rect 4509 1336 4522 1366
rect 4537 1348 4567 1366
rect 4610 1336 4623 1366
rect 4751 1336 4764 1366
rect 4779 1348 4809 1366
rect 4852 1352 4866 1366
rect 4902 1352 5122 1366
rect 4853 1350 4866 1352
rect 4819 1338 4834 1350
rect 4816 1336 4838 1338
rect 4843 1336 4873 1350
rect 4934 1348 5087 1352
rect 4916 1336 5108 1348
rect 5151 1336 5181 1350
rect 5187 1336 5200 1366
rect 5215 1348 5245 1366
rect 5288 1336 5301 1366
rect 5331 1336 5344 1366
rect 5359 1348 5389 1366
rect 5432 1352 5446 1366
rect 5482 1352 5702 1366
rect 5433 1350 5446 1352
rect 5399 1338 5414 1350
rect 5396 1336 5418 1338
rect 5423 1336 5453 1350
rect 5514 1348 5667 1352
rect 5496 1336 5688 1348
rect 5731 1336 5761 1350
rect 5767 1336 5780 1366
rect 5795 1348 5825 1366
rect 5868 1336 5881 1366
rect 3469 1322 4623 1336
rect 4736 1322 5889 1336
rect 3493 1218 3506 1322
rect 3551 1300 3552 1310
rect 3567 1300 3580 1310
rect 3551 1296 3580 1300
rect 3585 1296 3615 1322
rect 3633 1308 3649 1310
rect 3721 1308 3774 1322
rect 3722 1306 3786 1308
rect 3829 1306 3844 1322
rect 3893 1319 3923 1322
rect 3893 1316 3929 1319
rect 3859 1308 3875 1310
rect 3633 1296 3648 1300
rect 3551 1294 3648 1296
rect 3676 1294 3844 1306
rect 3860 1296 3875 1300
rect 3893 1297 3932 1316
rect 3951 1310 3958 1311
rect 3957 1303 3958 1310
rect 3941 1300 3942 1303
rect 3957 1300 3970 1303
rect 3893 1296 3923 1297
rect 3932 1296 3938 1297
rect 3941 1296 3970 1300
rect 3860 1295 3970 1296
rect 3860 1294 3976 1295
rect 3535 1286 3586 1294
rect 3535 1274 3560 1286
rect 3567 1274 3586 1286
rect 3617 1286 3667 1294
rect 3617 1278 3633 1286
rect 3640 1284 3667 1286
rect 3676 1284 3897 1294
rect 3640 1274 3897 1284
rect 3926 1286 3976 1294
rect 3926 1277 3942 1286
rect 3535 1266 3586 1274
rect 3633 1266 3897 1274
rect 3923 1274 3942 1277
rect 3949 1274 3976 1286
rect 3923 1266 3976 1274
rect 3551 1258 3552 1266
rect 3567 1258 3580 1266
rect 3551 1250 3567 1258
rect 3548 1243 3567 1246
rect 3548 1234 3570 1243
rect 3521 1224 3570 1234
rect 3521 1218 3551 1224
rect 3570 1219 3575 1224
rect 3493 1202 3567 1218
rect 3585 1210 3615 1266
rect 3650 1256 3858 1266
rect 3893 1262 3938 1266
rect 3941 1265 3942 1266
rect 3957 1265 3970 1266
rect 3676 1226 3865 1256
rect 3691 1223 3865 1226
rect 3684 1220 3865 1223
rect 3493 1200 3506 1202
rect 3521 1200 3555 1202
rect 3493 1184 3567 1200
rect 3594 1196 3607 1210
rect 3622 1196 3638 1212
rect 3684 1207 3695 1220
rect 3477 1162 3478 1178
rect 3493 1162 3506 1184
rect 3521 1162 3551 1184
rect 3594 1180 3656 1196
rect 3684 1189 3695 1205
rect 3700 1200 3710 1220
rect 3720 1200 3734 1220
rect 3737 1207 3746 1220
rect 3762 1207 3771 1220
rect 3700 1189 3734 1200
rect 3737 1189 3746 1205
rect 3762 1189 3771 1205
rect 3778 1200 3788 1220
rect 3798 1200 3812 1220
rect 3813 1207 3824 1220
rect 3778 1189 3812 1200
rect 3813 1189 3824 1205
rect 3870 1196 3886 1212
rect 3893 1210 3923 1262
rect 3957 1258 3958 1265
rect 3942 1250 3958 1258
rect 3929 1218 3942 1237
rect 3957 1218 3987 1234
rect 3929 1202 4003 1218
rect 3929 1200 3942 1202
rect 3957 1200 3991 1202
rect 3594 1178 3607 1180
rect 3622 1178 3656 1180
rect 3594 1162 3656 1178
rect 3700 1173 3716 1176
rect 3778 1173 3808 1184
rect 3856 1180 3902 1196
rect 3929 1184 4003 1200
rect 3856 1178 3890 1180
rect 3855 1162 3902 1178
rect 3929 1162 3942 1184
rect 3957 1162 3987 1184
rect 4014 1162 4015 1178
rect 4030 1162 4043 1322
rect 4073 1218 4086 1322
rect 4131 1300 4132 1310
rect 4147 1300 4160 1310
rect 4131 1296 4160 1300
rect 4165 1296 4195 1322
rect 4213 1308 4229 1310
rect 4301 1308 4354 1322
rect 4302 1306 4366 1308
rect 4409 1306 4424 1322
rect 4473 1319 4503 1322
rect 4473 1316 4509 1319
rect 4439 1308 4455 1310
rect 4213 1296 4228 1300
rect 4131 1294 4228 1296
rect 4256 1294 4424 1306
rect 4440 1296 4455 1300
rect 4473 1297 4512 1316
rect 4531 1310 4538 1311
rect 4537 1303 4538 1310
rect 4521 1300 4522 1303
rect 4537 1300 4550 1303
rect 4473 1296 4503 1297
rect 4512 1296 4518 1297
rect 4521 1296 4550 1300
rect 4440 1295 4550 1296
rect 4440 1294 4556 1295
rect 4115 1286 4166 1294
rect 4115 1274 4140 1286
rect 4147 1274 4166 1286
rect 4197 1286 4247 1294
rect 4197 1278 4213 1286
rect 4220 1284 4247 1286
rect 4256 1284 4477 1294
rect 4220 1274 4477 1284
rect 4506 1286 4556 1294
rect 4506 1277 4522 1286
rect 4115 1266 4166 1274
rect 4213 1266 4477 1274
rect 4503 1274 4522 1277
rect 4529 1274 4556 1286
rect 4503 1266 4556 1274
rect 4131 1258 4132 1266
rect 4147 1258 4160 1266
rect 4131 1250 4147 1258
rect 4128 1243 4147 1246
rect 4128 1234 4150 1243
rect 4101 1224 4150 1234
rect 4101 1218 4131 1224
rect 4150 1219 4155 1224
rect 4073 1202 4147 1218
rect 4165 1210 4195 1266
rect 4230 1256 4438 1266
rect 4473 1262 4518 1266
rect 4521 1265 4522 1266
rect 4537 1265 4550 1266
rect 4256 1226 4445 1256
rect 4271 1223 4445 1226
rect 4264 1220 4445 1223
rect 4073 1200 4086 1202
rect 4101 1200 4135 1202
rect 4073 1184 4147 1200
rect 4174 1196 4187 1210
rect 4202 1196 4218 1212
rect 4264 1207 4275 1220
rect 4057 1162 4058 1178
rect 4073 1162 4086 1184
rect 4101 1162 4131 1184
rect 4174 1180 4236 1196
rect 4264 1189 4275 1205
rect 4280 1200 4290 1220
rect 4300 1200 4314 1220
rect 4317 1207 4326 1220
rect 4342 1207 4351 1220
rect 4280 1189 4314 1200
rect 4317 1189 4326 1205
rect 4342 1189 4351 1205
rect 4358 1200 4368 1220
rect 4378 1200 4392 1220
rect 4393 1207 4404 1220
rect 4358 1189 4392 1200
rect 4393 1189 4404 1205
rect 4450 1196 4466 1212
rect 4473 1210 4503 1262
rect 4537 1258 4538 1265
rect 4522 1250 4538 1258
rect 4509 1218 4522 1237
rect 4537 1218 4567 1234
rect 4509 1202 4583 1218
rect 4509 1200 4522 1202
rect 4537 1200 4571 1202
rect 4174 1178 4187 1180
rect 4202 1178 4236 1180
rect 4174 1162 4236 1178
rect 4280 1173 4296 1176
rect 4358 1173 4388 1184
rect 4436 1180 4482 1196
rect 4509 1184 4583 1200
rect 4436 1178 4470 1180
rect 4435 1162 4482 1178
rect 4509 1162 4522 1184
rect 4537 1162 4567 1184
rect 4594 1162 4595 1178
rect 4610 1162 4623 1322
rect 4751 1218 4764 1322
rect 4809 1300 4810 1310
rect 4825 1300 4838 1310
rect 4809 1296 4838 1300
rect 4843 1296 4873 1322
rect 4891 1308 4907 1310
rect 4979 1308 5032 1322
rect 4980 1306 5044 1308
rect 5087 1306 5102 1322
rect 5151 1319 5181 1322
rect 5151 1316 5187 1319
rect 5117 1308 5133 1310
rect 4891 1296 4906 1300
rect 4809 1294 4906 1296
rect 4934 1294 5102 1306
rect 5118 1296 5133 1300
rect 5151 1297 5190 1316
rect 5209 1310 5216 1311
rect 5215 1303 5216 1310
rect 5199 1300 5200 1303
rect 5215 1300 5228 1303
rect 5151 1296 5181 1297
rect 5190 1296 5196 1297
rect 5199 1296 5228 1300
rect 5118 1295 5228 1296
rect 5118 1294 5234 1295
rect 4793 1286 4844 1294
rect 4793 1274 4818 1286
rect 4825 1274 4844 1286
rect 4875 1286 4925 1294
rect 4875 1278 4891 1286
rect 4898 1284 4925 1286
rect 4934 1284 5155 1294
rect 4898 1274 5155 1284
rect 5184 1286 5234 1294
rect 5184 1277 5200 1286
rect 4793 1266 4844 1274
rect 4891 1266 5155 1274
rect 5181 1274 5200 1277
rect 5207 1274 5234 1286
rect 5181 1266 5234 1274
rect 4809 1258 4810 1266
rect 4825 1258 4838 1266
rect 4809 1250 4825 1258
rect 4806 1243 4825 1246
rect 4806 1234 4828 1243
rect 4779 1224 4828 1234
rect 4779 1218 4809 1224
rect 4828 1219 4833 1224
rect 4751 1202 4825 1218
rect 4843 1210 4873 1266
rect 4908 1256 5116 1266
rect 5151 1262 5196 1266
rect 5199 1265 5200 1266
rect 5215 1265 5228 1266
rect 4934 1226 5123 1256
rect 4949 1223 5123 1226
rect 4942 1220 5123 1223
rect 4751 1200 4764 1202
rect 4779 1200 4813 1202
rect 4751 1184 4825 1200
rect 4852 1196 4865 1210
rect 4880 1196 4896 1212
rect 4942 1207 4953 1220
rect 4735 1162 4736 1178
rect 4751 1162 4764 1184
rect 4779 1162 4809 1184
rect 4852 1180 4914 1196
rect 4942 1189 4953 1205
rect 4958 1200 4968 1220
rect 4978 1200 4992 1220
rect 4995 1207 5004 1220
rect 5020 1207 5029 1220
rect 4958 1189 4992 1200
rect 4995 1189 5004 1205
rect 5020 1189 5029 1205
rect 5036 1200 5046 1220
rect 5056 1200 5070 1220
rect 5071 1207 5082 1220
rect 5036 1189 5070 1200
rect 5071 1189 5082 1205
rect 5128 1196 5144 1212
rect 5151 1210 5181 1262
rect 5215 1258 5216 1265
rect 5200 1250 5216 1258
rect 5187 1218 5200 1237
rect 5215 1218 5245 1234
rect 5187 1202 5261 1218
rect 5187 1200 5200 1202
rect 5215 1200 5249 1202
rect 4852 1178 4865 1180
rect 4880 1178 4914 1180
rect 4852 1162 4914 1178
rect 4958 1173 4974 1176
rect 5036 1173 5066 1184
rect 5114 1180 5160 1196
rect 5187 1184 5261 1200
rect 5114 1178 5148 1180
rect 5113 1162 5160 1178
rect 5187 1162 5200 1184
rect 5215 1162 5245 1184
rect 5272 1162 5273 1178
rect 5288 1162 5301 1322
rect 5331 1218 5344 1322
rect 5389 1300 5390 1310
rect 5405 1300 5418 1310
rect 5389 1296 5418 1300
rect 5423 1296 5453 1322
rect 5471 1308 5487 1310
rect 5559 1308 5612 1322
rect 5560 1306 5624 1308
rect 5667 1306 5682 1322
rect 5731 1319 5761 1322
rect 5731 1316 5767 1319
rect 5697 1308 5713 1310
rect 5471 1296 5486 1300
rect 5389 1294 5486 1296
rect 5514 1294 5682 1306
rect 5698 1296 5713 1300
rect 5731 1297 5770 1316
rect 5789 1310 5796 1311
rect 5795 1303 5796 1310
rect 5779 1300 5780 1303
rect 5795 1300 5808 1303
rect 5731 1296 5761 1297
rect 5770 1296 5776 1297
rect 5779 1296 5808 1300
rect 5698 1295 5808 1296
rect 5698 1294 5814 1295
rect 5373 1286 5424 1294
rect 5373 1274 5398 1286
rect 5405 1274 5424 1286
rect 5455 1286 5505 1294
rect 5455 1278 5471 1286
rect 5478 1284 5505 1286
rect 5514 1284 5735 1294
rect 5478 1274 5735 1284
rect 5764 1286 5814 1294
rect 5764 1277 5780 1286
rect 5373 1266 5424 1274
rect 5471 1266 5735 1274
rect 5761 1274 5780 1277
rect 5787 1274 5814 1286
rect 5761 1266 5814 1274
rect 5389 1258 5390 1266
rect 5405 1258 5418 1266
rect 5389 1250 5405 1258
rect 5386 1243 5405 1246
rect 5386 1234 5408 1243
rect 5359 1224 5408 1234
rect 5359 1218 5389 1224
rect 5408 1219 5413 1224
rect 5331 1202 5405 1218
rect 5423 1210 5453 1266
rect 5488 1256 5696 1266
rect 5731 1262 5776 1266
rect 5779 1265 5780 1266
rect 5795 1265 5808 1266
rect 5514 1226 5703 1256
rect 5529 1223 5703 1226
rect 5522 1220 5703 1223
rect 5331 1200 5344 1202
rect 5359 1200 5393 1202
rect 5331 1184 5405 1200
rect 5432 1196 5445 1210
rect 5460 1196 5476 1212
rect 5522 1207 5533 1220
rect 5315 1162 5316 1178
rect 5331 1162 5344 1184
rect 5359 1162 5389 1184
rect 5432 1180 5494 1196
rect 5522 1189 5533 1205
rect 5538 1200 5548 1220
rect 5558 1200 5572 1220
rect 5575 1207 5584 1220
rect 5600 1207 5609 1220
rect 5538 1189 5572 1200
rect 5575 1189 5584 1205
rect 5600 1189 5609 1205
rect 5616 1200 5626 1220
rect 5636 1200 5650 1220
rect 5651 1207 5662 1220
rect 5616 1189 5650 1200
rect 5651 1189 5662 1205
rect 5708 1196 5724 1212
rect 5731 1210 5761 1262
rect 5795 1258 5796 1265
rect 5780 1250 5796 1258
rect 5767 1218 5780 1237
rect 5795 1218 5825 1234
rect 5767 1202 5841 1218
rect 5767 1200 5780 1202
rect 5795 1200 5829 1202
rect 5432 1178 5445 1180
rect 5460 1178 5494 1180
rect 5432 1162 5494 1178
rect 5538 1173 5554 1176
rect 5616 1173 5646 1184
rect 5694 1180 5740 1196
rect 5767 1184 5841 1200
rect 5694 1178 5728 1180
rect 5693 1162 5740 1178
rect 5767 1162 5780 1184
rect 5795 1162 5825 1184
rect 5852 1162 5853 1178
rect 5868 1162 5881 1322
rect 3471 1154 3512 1162
rect 3471 1128 3486 1154
rect 3493 1128 3512 1154
rect 3576 1150 3638 1162
rect 3650 1150 3725 1162
rect 3783 1150 3858 1162
rect 3870 1150 3901 1162
rect 3907 1150 3942 1162
rect 3576 1148 3738 1150
rect 3471 1120 3512 1128
rect 3594 1124 3607 1148
rect 3622 1146 3637 1148
rect 3477 1110 3478 1120
rect 3493 1110 3506 1120
rect 3521 1110 3551 1124
rect 3594 1110 3637 1124
rect 3661 1121 3668 1128
rect 3671 1124 3738 1148
rect 3770 1148 3942 1150
rect 3740 1126 3768 1130
rect 3770 1126 3850 1148
rect 3871 1146 3886 1148
rect 3740 1124 3850 1126
rect 3671 1120 3850 1124
rect 3644 1110 3674 1120
rect 3676 1110 3829 1120
rect 3837 1110 3867 1120
rect 3871 1110 3901 1124
rect 3929 1110 3942 1148
rect 4014 1154 4049 1162
rect 4014 1128 4015 1154
rect 4022 1128 4049 1154
rect 3957 1110 3987 1124
rect 4014 1120 4049 1128
rect 4051 1154 4092 1162
rect 4051 1128 4066 1154
rect 4073 1128 4092 1154
rect 4156 1150 4218 1162
rect 4230 1150 4305 1162
rect 4363 1150 4438 1162
rect 4450 1150 4481 1162
rect 4487 1150 4522 1162
rect 4156 1148 4318 1150
rect 4051 1120 4092 1128
rect 4174 1124 4187 1148
rect 4202 1146 4217 1148
rect 4014 1110 4015 1120
rect 4030 1110 4043 1120
rect 4057 1110 4058 1120
rect 4073 1110 4086 1120
rect 4101 1110 4131 1124
rect 4174 1110 4217 1124
rect 4241 1121 4248 1128
rect 4251 1124 4318 1148
rect 4350 1148 4522 1150
rect 4320 1126 4348 1130
rect 4350 1126 4430 1148
rect 4451 1146 4466 1148
rect 4320 1124 4430 1126
rect 4251 1120 4430 1124
rect 4224 1110 4254 1120
rect 4256 1110 4409 1120
rect 4417 1110 4447 1120
rect 4451 1110 4481 1124
rect 4509 1110 4522 1148
rect 4594 1154 4629 1162
rect 4594 1128 4595 1154
rect 4602 1128 4629 1154
rect 4537 1110 4567 1124
rect 4594 1120 4629 1128
rect 4729 1154 4770 1162
rect 4729 1128 4744 1154
rect 4751 1128 4770 1154
rect 4834 1150 4896 1162
rect 4908 1150 4983 1162
rect 5041 1150 5116 1162
rect 5128 1150 5159 1162
rect 5165 1150 5200 1162
rect 4834 1148 4996 1150
rect 4729 1120 4770 1128
rect 4852 1124 4865 1148
rect 4880 1146 4895 1148
rect 4594 1110 4595 1120
rect 4610 1110 4623 1120
rect 3469 1096 4623 1110
rect 4735 1110 4736 1120
rect 4751 1110 4764 1120
rect 4779 1110 4809 1124
rect 4852 1110 4895 1124
rect 4919 1121 4926 1128
rect 4929 1124 4996 1148
rect 5028 1148 5200 1150
rect 4998 1126 5026 1130
rect 5028 1126 5108 1148
rect 5129 1146 5144 1148
rect 4998 1124 5108 1126
rect 4929 1120 5108 1124
rect 4902 1110 4932 1120
rect 4934 1110 5087 1120
rect 5095 1110 5125 1120
rect 5129 1110 5159 1124
rect 5187 1110 5200 1148
rect 5272 1154 5307 1162
rect 5272 1128 5273 1154
rect 5280 1128 5307 1154
rect 5215 1110 5245 1124
rect 5272 1120 5307 1128
rect 5309 1154 5350 1162
rect 5309 1128 5324 1154
rect 5331 1128 5350 1154
rect 5414 1150 5476 1162
rect 5488 1150 5563 1162
rect 5621 1150 5696 1162
rect 5708 1150 5739 1162
rect 5745 1150 5780 1162
rect 5414 1148 5576 1150
rect 5309 1120 5350 1128
rect 5432 1124 5445 1148
rect 5460 1146 5475 1148
rect 5272 1110 5273 1120
rect 5288 1110 5301 1120
rect 5315 1110 5316 1120
rect 5331 1110 5344 1120
rect 5359 1110 5389 1124
rect 5432 1110 5475 1124
rect 5499 1121 5506 1128
rect 5509 1124 5576 1148
rect 5608 1148 5780 1150
rect 5578 1126 5606 1130
rect 5608 1126 5688 1148
rect 5709 1146 5724 1148
rect 5578 1124 5688 1126
rect 5509 1120 5688 1124
rect 5482 1110 5512 1120
rect 5514 1110 5667 1120
rect 5675 1110 5705 1120
rect 5709 1110 5739 1124
rect 5767 1110 5780 1148
rect 5852 1154 5887 1162
rect 5852 1128 5853 1154
rect 5860 1128 5887 1154
rect 5795 1110 5825 1124
rect 5852 1120 5887 1128
rect 5852 1110 5853 1120
rect 5868 1110 5881 1120
rect 4735 1104 5889 1110
rect 4736 1096 5889 1104
rect 3493 1066 3506 1096
rect 3521 1078 3551 1096
rect 3594 1082 3608 1096
rect 3644 1082 3864 1096
rect 3595 1080 3608 1082
rect 3561 1068 3576 1080
rect 3558 1066 3580 1068
rect 3585 1066 3615 1080
rect 3676 1078 3829 1082
rect 3658 1066 3850 1078
rect 3893 1066 3923 1080
rect 3929 1066 3942 1096
rect 3957 1078 3987 1096
rect 4030 1066 4043 1096
rect 4073 1066 4086 1096
rect 4101 1078 4131 1096
rect 4174 1082 4188 1096
rect 4224 1082 4444 1096
rect 4175 1080 4188 1082
rect 4141 1068 4156 1080
rect 4138 1066 4160 1068
rect 4165 1066 4195 1080
rect 4256 1078 4409 1082
rect 4238 1066 4430 1078
rect 4473 1066 4503 1080
rect 4509 1066 4522 1096
rect 4537 1078 4567 1096
rect 4610 1066 4623 1096
rect 4751 1066 4764 1096
rect 4779 1078 4809 1096
rect 4852 1082 4866 1096
rect 4902 1082 5122 1096
rect 4853 1080 4866 1082
rect 4819 1068 4834 1080
rect 4816 1066 4838 1068
rect 4843 1066 4873 1080
rect 4934 1078 5087 1082
rect 4916 1066 5108 1078
rect 5151 1066 5181 1080
rect 5187 1066 5200 1096
rect 5215 1078 5245 1096
rect 5288 1066 5301 1096
rect 5331 1066 5344 1096
rect 5359 1078 5389 1096
rect 5432 1082 5446 1096
rect 5482 1082 5702 1096
rect 5433 1080 5446 1082
rect 5399 1068 5414 1080
rect 5396 1066 5418 1068
rect 5423 1066 5453 1080
rect 5514 1078 5667 1082
rect 5496 1066 5688 1078
rect 5731 1066 5761 1080
rect 5767 1066 5780 1096
rect 5795 1078 5825 1096
rect 5868 1066 5881 1096
rect 3469 1052 4623 1066
rect 4736 1052 5889 1066
rect 3493 948 3506 1052
rect 3551 1030 3552 1040
rect 3567 1030 3580 1040
rect 3551 1026 3580 1030
rect 3585 1026 3615 1052
rect 3633 1038 3649 1040
rect 3721 1038 3774 1052
rect 3722 1036 3786 1038
rect 3829 1036 3844 1052
rect 3893 1049 3923 1052
rect 3893 1046 3929 1049
rect 3859 1038 3875 1040
rect 3633 1026 3648 1030
rect 3551 1024 3648 1026
rect 3676 1024 3844 1036
rect 3860 1026 3875 1030
rect 3893 1027 3932 1046
rect 3951 1040 3958 1041
rect 3957 1033 3958 1040
rect 3941 1030 3942 1033
rect 3957 1030 3970 1033
rect 3893 1026 3923 1027
rect 3932 1026 3938 1027
rect 3941 1026 3970 1030
rect 3860 1025 3970 1026
rect 3860 1024 3976 1025
rect 3535 1016 3586 1024
rect 3535 1004 3560 1016
rect 3567 1004 3586 1016
rect 3617 1016 3667 1024
rect 3617 1008 3633 1016
rect 3640 1014 3667 1016
rect 3676 1014 3897 1024
rect 3640 1004 3897 1014
rect 3926 1016 3976 1024
rect 3926 1007 3942 1016
rect 3535 996 3586 1004
rect 3633 996 3897 1004
rect 3923 1004 3942 1007
rect 3949 1004 3976 1016
rect 3923 996 3976 1004
rect 3551 988 3552 996
rect 3567 988 3580 996
rect 3551 980 3567 988
rect 3548 973 3567 976
rect 3548 964 3570 973
rect 3521 954 3570 964
rect 3521 948 3551 954
rect 3570 949 3575 954
rect 3493 932 3567 948
rect 3585 940 3615 996
rect 3650 986 3858 996
rect 3893 992 3938 996
rect 3941 995 3942 996
rect 3957 995 3970 996
rect 3676 956 3865 986
rect 3691 953 3865 956
rect 3684 950 3865 953
rect 3493 930 3506 932
rect 3521 930 3555 932
rect 3493 914 3567 930
rect 3594 926 3607 940
rect 3622 926 3638 942
rect 3684 937 3695 950
rect 3477 892 3478 908
rect 3493 892 3506 914
rect 3521 892 3551 914
rect 3594 910 3656 926
rect 3684 919 3695 935
rect 3700 930 3710 950
rect 3720 930 3734 950
rect 3737 937 3746 950
rect 3762 937 3771 950
rect 3700 919 3734 930
rect 3737 919 3746 935
rect 3762 919 3771 935
rect 3778 930 3788 950
rect 3798 930 3812 950
rect 3813 937 3824 950
rect 3778 919 3812 930
rect 3813 919 3824 935
rect 3870 926 3886 942
rect 3893 940 3923 992
rect 3957 988 3958 995
rect 3942 980 3958 988
rect 3929 948 3942 967
rect 3957 948 3987 964
rect 3929 932 4003 948
rect 3929 930 3942 932
rect 3957 930 3991 932
rect 3594 908 3607 910
rect 3622 908 3656 910
rect 3594 892 3656 908
rect 3700 903 3716 906
rect 3778 903 3808 914
rect 3856 910 3902 926
rect 3929 914 4003 930
rect 3856 908 3890 910
rect 3855 892 3902 908
rect 3929 892 3942 914
rect 3957 892 3987 914
rect 4014 892 4015 908
rect 4030 892 4043 1052
rect 4073 948 4086 1052
rect 4131 1030 4132 1040
rect 4147 1030 4160 1040
rect 4131 1026 4160 1030
rect 4165 1026 4195 1052
rect 4213 1038 4229 1040
rect 4301 1038 4354 1052
rect 4302 1036 4366 1038
rect 4409 1036 4424 1052
rect 4473 1049 4503 1052
rect 4473 1046 4509 1049
rect 4439 1038 4455 1040
rect 4213 1026 4228 1030
rect 4131 1024 4228 1026
rect 4256 1024 4424 1036
rect 4440 1026 4455 1030
rect 4473 1027 4512 1046
rect 4531 1040 4538 1041
rect 4537 1033 4538 1040
rect 4521 1030 4522 1033
rect 4537 1030 4550 1033
rect 4473 1026 4503 1027
rect 4512 1026 4518 1027
rect 4521 1026 4550 1030
rect 4440 1025 4550 1026
rect 4440 1024 4556 1025
rect 4115 1016 4166 1024
rect 4115 1004 4140 1016
rect 4147 1004 4166 1016
rect 4197 1016 4247 1024
rect 4197 1008 4213 1016
rect 4220 1014 4247 1016
rect 4256 1014 4477 1024
rect 4220 1004 4477 1014
rect 4506 1016 4556 1024
rect 4506 1007 4522 1016
rect 4115 996 4166 1004
rect 4213 996 4477 1004
rect 4503 1004 4522 1007
rect 4529 1004 4556 1016
rect 4503 996 4556 1004
rect 4131 988 4132 996
rect 4147 988 4160 996
rect 4131 980 4147 988
rect 4128 973 4147 976
rect 4128 964 4150 973
rect 4101 954 4150 964
rect 4101 948 4131 954
rect 4150 949 4155 954
rect 4073 932 4147 948
rect 4165 940 4195 996
rect 4230 986 4438 996
rect 4473 992 4518 996
rect 4521 995 4522 996
rect 4537 995 4550 996
rect 4256 956 4445 986
rect 4271 953 4445 956
rect 4264 950 4445 953
rect 4073 930 4086 932
rect 4101 930 4135 932
rect 4073 914 4147 930
rect 4174 926 4187 940
rect 4202 926 4218 942
rect 4264 937 4275 950
rect 4057 892 4058 908
rect 4073 892 4086 914
rect 4101 892 4131 914
rect 4174 910 4236 926
rect 4264 919 4275 935
rect 4280 930 4290 950
rect 4300 930 4314 950
rect 4317 937 4326 950
rect 4342 937 4351 950
rect 4280 919 4314 930
rect 4317 919 4326 935
rect 4342 919 4351 935
rect 4358 930 4368 950
rect 4378 930 4392 950
rect 4393 937 4404 950
rect 4358 919 4392 930
rect 4393 919 4404 935
rect 4450 926 4466 942
rect 4473 940 4503 992
rect 4537 988 4538 995
rect 4522 980 4538 988
rect 4509 948 4522 967
rect 4537 948 4567 964
rect 4509 932 4583 948
rect 4509 930 4522 932
rect 4537 930 4571 932
rect 4174 908 4187 910
rect 4202 908 4236 910
rect 4174 892 4236 908
rect 4280 903 4296 906
rect 4358 903 4388 914
rect 4436 910 4482 926
rect 4509 914 4583 930
rect 4436 908 4470 910
rect 4435 892 4482 908
rect 4509 892 4522 914
rect 4537 892 4567 914
rect 4594 892 4595 908
rect 4610 892 4623 1052
rect 4751 948 4764 1052
rect 4809 1030 4810 1040
rect 4825 1030 4838 1040
rect 4809 1026 4838 1030
rect 4843 1026 4873 1052
rect 4891 1038 4907 1040
rect 4979 1038 5032 1052
rect 4980 1036 5044 1038
rect 5087 1036 5102 1052
rect 5151 1049 5181 1052
rect 5151 1046 5187 1049
rect 5117 1038 5133 1040
rect 4891 1026 4906 1030
rect 4809 1024 4906 1026
rect 4934 1024 5102 1036
rect 5118 1026 5133 1030
rect 5151 1027 5190 1046
rect 5209 1040 5216 1041
rect 5215 1033 5216 1040
rect 5199 1030 5200 1033
rect 5215 1030 5228 1033
rect 5151 1026 5181 1027
rect 5190 1026 5196 1027
rect 5199 1026 5228 1030
rect 5118 1025 5228 1026
rect 5118 1024 5234 1025
rect 4793 1016 4844 1024
rect 4793 1004 4818 1016
rect 4825 1004 4844 1016
rect 4875 1016 4925 1024
rect 4875 1008 4891 1016
rect 4898 1014 4925 1016
rect 4934 1014 5155 1024
rect 4898 1004 5155 1014
rect 5184 1016 5234 1024
rect 5184 1007 5200 1016
rect 4793 996 4844 1004
rect 4891 996 5155 1004
rect 5181 1004 5200 1007
rect 5207 1004 5234 1016
rect 5181 996 5234 1004
rect 4809 988 4810 996
rect 4825 988 4838 996
rect 4809 980 4825 988
rect 4806 973 4825 976
rect 4806 964 4828 973
rect 4779 954 4828 964
rect 4779 948 4809 954
rect 4828 949 4833 954
rect 4751 932 4825 948
rect 4843 940 4873 996
rect 4908 986 5116 996
rect 5151 992 5196 996
rect 5199 995 5200 996
rect 5215 995 5228 996
rect 4934 956 5123 986
rect 4949 953 5123 956
rect 4942 950 5123 953
rect 4751 930 4764 932
rect 4779 930 4813 932
rect 4751 914 4825 930
rect 4852 926 4865 940
rect 4880 926 4896 942
rect 4942 937 4953 950
rect 4735 892 4736 908
rect 4751 892 4764 914
rect 4779 892 4809 914
rect 4852 910 4914 926
rect 4942 919 4953 935
rect 4958 930 4968 950
rect 4978 930 4992 950
rect 4995 937 5004 950
rect 5020 937 5029 950
rect 4958 919 4992 930
rect 4995 919 5004 935
rect 5020 919 5029 935
rect 5036 930 5046 950
rect 5056 930 5070 950
rect 5071 937 5082 950
rect 5036 919 5070 930
rect 5071 919 5082 935
rect 5128 926 5144 942
rect 5151 940 5181 992
rect 5215 988 5216 995
rect 5200 980 5216 988
rect 5187 948 5200 967
rect 5215 948 5245 964
rect 5187 932 5261 948
rect 5187 930 5200 932
rect 5215 930 5249 932
rect 4852 908 4865 910
rect 4880 908 4914 910
rect 4852 892 4914 908
rect 4958 903 4974 906
rect 5036 903 5066 914
rect 5114 910 5160 926
rect 5187 914 5261 930
rect 5114 908 5148 910
rect 5113 892 5160 908
rect 5187 892 5200 914
rect 5215 892 5245 914
rect 5272 892 5273 908
rect 5288 892 5301 1052
rect 5331 948 5344 1052
rect 5389 1030 5390 1040
rect 5405 1030 5418 1040
rect 5389 1026 5418 1030
rect 5423 1026 5453 1052
rect 5471 1038 5487 1040
rect 5559 1038 5612 1052
rect 5560 1036 5624 1038
rect 5667 1036 5682 1052
rect 5731 1049 5761 1052
rect 5731 1046 5767 1049
rect 5697 1038 5713 1040
rect 5471 1026 5486 1030
rect 5389 1024 5486 1026
rect 5514 1024 5682 1036
rect 5698 1026 5713 1030
rect 5731 1027 5770 1046
rect 5789 1040 5796 1041
rect 5795 1033 5796 1040
rect 5779 1030 5780 1033
rect 5795 1030 5808 1033
rect 5731 1026 5761 1027
rect 5770 1026 5776 1027
rect 5779 1026 5808 1030
rect 5698 1025 5808 1026
rect 5698 1024 5814 1025
rect 5373 1016 5424 1024
rect 5373 1004 5398 1016
rect 5405 1004 5424 1016
rect 5455 1016 5505 1024
rect 5455 1008 5471 1016
rect 5478 1014 5505 1016
rect 5514 1014 5735 1024
rect 5478 1004 5735 1014
rect 5764 1016 5814 1024
rect 5764 1007 5780 1016
rect 5373 996 5424 1004
rect 5471 996 5735 1004
rect 5761 1004 5780 1007
rect 5787 1004 5814 1016
rect 5761 996 5814 1004
rect 5389 988 5390 996
rect 5405 988 5418 996
rect 5389 980 5405 988
rect 5386 973 5405 976
rect 5386 964 5408 973
rect 5359 954 5408 964
rect 5359 948 5389 954
rect 5408 949 5413 954
rect 5331 932 5405 948
rect 5423 940 5453 996
rect 5488 986 5696 996
rect 5731 992 5776 996
rect 5779 995 5780 996
rect 5795 995 5808 996
rect 5514 956 5703 986
rect 5529 953 5703 956
rect 5522 950 5703 953
rect 5331 930 5344 932
rect 5359 930 5393 932
rect 5331 914 5405 930
rect 5432 926 5445 940
rect 5460 926 5476 942
rect 5522 937 5533 950
rect 5315 892 5316 908
rect 5331 892 5344 914
rect 5359 892 5389 914
rect 5432 910 5494 926
rect 5522 919 5533 935
rect 5538 930 5548 950
rect 5558 930 5572 950
rect 5575 937 5584 950
rect 5600 937 5609 950
rect 5538 919 5572 930
rect 5575 919 5584 935
rect 5600 919 5609 935
rect 5616 930 5626 950
rect 5636 930 5650 950
rect 5651 937 5662 950
rect 5616 919 5650 930
rect 5651 919 5662 935
rect 5708 926 5724 942
rect 5731 940 5761 992
rect 5795 988 5796 995
rect 5780 980 5796 988
rect 5767 948 5780 967
rect 5795 948 5825 964
rect 5767 932 5841 948
rect 5767 930 5780 932
rect 5795 930 5829 932
rect 5432 908 5445 910
rect 5460 908 5494 910
rect 5432 892 5494 908
rect 5538 903 5554 906
rect 5616 903 5646 914
rect 5694 910 5740 926
rect 5767 914 5841 930
rect 5694 908 5728 910
rect 5693 892 5740 908
rect 5767 892 5780 914
rect 5795 892 5825 914
rect 5852 892 5853 908
rect 5868 892 5881 1052
rect 3471 884 3512 892
rect 3471 858 3486 884
rect 3493 858 3512 884
rect 3576 880 3638 892
rect 3650 880 3725 892
rect 3783 880 3858 892
rect 3870 880 3901 892
rect 3907 880 3942 892
rect 3576 878 3738 880
rect 3471 850 3512 858
rect 3594 854 3607 878
rect 3622 876 3637 878
rect 3477 840 3478 850
rect 3493 840 3506 850
rect 3521 840 3551 854
rect 3594 840 3637 854
rect 3661 851 3668 858
rect 3671 854 3738 878
rect 3770 878 3942 880
rect 3740 856 3768 860
rect 3770 856 3850 878
rect 3871 876 3886 878
rect 3740 854 3850 856
rect 3671 850 3850 854
rect 3644 840 3674 850
rect 3676 840 3829 850
rect 3837 840 3867 850
rect 3871 840 3901 854
rect 3929 840 3942 878
rect 4014 884 4049 892
rect 4014 858 4015 884
rect 4022 858 4049 884
rect 3957 840 3987 854
rect 4014 850 4049 858
rect 4051 884 4092 892
rect 4051 858 4066 884
rect 4073 858 4092 884
rect 4156 880 4218 892
rect 4230 880 4305 892
rect 4363 880 4438 892
rect 4450 880 4481 892
rect 4487 880 4522 892
rect 4156 878 4318 880
rect 4051 850 4092 858
rect 4174 854 4187 878
rect 4202 876 4217 878
rect 4014 840 4015 850
rect 4030 840 4043 850
rect 4057 840 4058 850
rect 4073 840 4086 850
rect 4101 840 4131 854
rect 4174 840 4217 854
rect 4241 851 4248 858
rect 4251 854 4318 878
rect 4350 878 4522 880
rect 4320 856 4348 860
rect 4350 856 4430 878
rect 4451 876 4466 878
rect 4320 854 4430 856
rect 4251 850 4430 854
rect 4224 840 4254 850
rect 4256 840 4409 850
rect 4417 840 4447 850
rect 4451 840 4481 854
rect 4509 840 4522 878
rect 4594 884 4629 892
rect 4594 858 4595 884
rect 4602 858 4629 884
rect 4537 840 4567 854
rect 4594 850 4629 858
rect 4729 884 4770 892
rect 4729 858 4744 884
rect 4751 858 4770 884
rect 4834 880 4896 892
rect 4908 880 4983 892
rect 5041 880 5116 892
rect 5128 880 5159 892
rect 5165 880 5200 892
rect 4834 878 4996 880
rect 4729 850 4770 858
rect 4852 854 4865 878
rect 4880 876 4895 878
rect 4594 840 4595 850
rect 4610 840 4623 850
rect 3469 826 4623 840
rect 4735 840 4736 850
rect 4751 840 4764 850
rect 4779 840 4809 854
rect 4852 840 4895 854
rect 4919 851 4926 858
rect 4929 854 4996 878
rect 5028 878 5200 880
rect 4998 856 5026 860
rect 5028 856 5108 878
rect 5129 876 5144 878
rect 4998 854 5108 856
rect 4929 850 5108 854
rect 4902 840 4932 850
rect 4934 840 5087 850
rect 5095 840 5125 850
rect 5129 840 5159 854
rect 5187 840 5200 878
rect 5272 884 5307 892
rect 5272 858 5273 884
rect 5280 858 5307 884
rect 5215 840 5245 854
rect 5272 850 5307 858
rect 5309 884 5350 892
rect 5309 858 5324 884
rect 5331 858 5350 884
rect 5414 880 5476 892
rect 5488 880 5563 892
rect 5621 880 5696 892
rect 5708 880 5739 892
rect 5745 880 5780 892
rect 5414 878 5576 880
rect 5309 850 5350 858
rect 5432 854 5445 878
rect 5460 876 5475 878
rect 5272 840 5273 850
rect 5288 840 5301 850
rect 5315 840 5316 850
rect 5331 840 5344 850
rect 5359 840 5389 854
rect 5432 840 5475 854
rect 5499 851 5506 858
rect 5509 854 5576 878
rect 5608 878 5780 880
rect 5578 856 5606 860
rect 5608 856 5688 878
rect 5709 876 5724 878
rect 5578 854 5688 856
rect 5509 850 5688 854
rect 5482 840 5512 850
rect 5514 840 5667 850
rect 5675 840 5705 850
rect 5709 840 5739 854
rect 5767 840 5780 878
rect 5852 884 5887 892
rect 5852 858 5853 884
rect 5860 858 5887 884
rect 5795 840 5825 854
rect 5852 850 5887 858
rect 5852 840 5853 850
rect 5868 840 5881 850
rect 4735 834 5889 840
rect 4736 826 5889 834
rect 3493 796 3506 826
rect 3521 808 3551 826
rect 3594 812 3608 826
rect 3644 812 3864 826
rect 3595 810 3608 812
rect 3561 798 3576 810
rect 3558 796 3580 798
rect 3585 796 3615 810
rect 3676 808 3829 812
rect 3658 796 3850 808
rect 3893 796 3923 810
rect 3929 796 3942 826
rect 3957 808 3987 826
rect 4030 796 4043 826
rect 4073 796 4086 826
rect 4101 808 4131 826
rect 4174 812 4188 826
rect 4224 812 4444 826
rect 4175 810 4188 812
rect 4141 798 4156 810
rect 4138 796 4160 798
rect 4165 796 4195 810
rect 4256 808 4409 812
rect 4238 796 4430 808
rect 4473 796 4503 810
rect 4509 796 4522 826
rect 4537 808 4567 826
rect 4610 796 4623 826
rect 4751 796 4764 826
rect 4779 808 4809 826
rect 4852 812 4866 826
rect 4902 812 5122 826
rect 4853 810 4866 812
rect 4819 798 4834 810
rect 4816 796 4838 798
rect 4843 796 4873 810
rect 4934 808 5087 812
rect 4916 796 5108 808
rect 5151 796 5181 810
rect 5187 796 5200 826
rect 5215 808 5245 826
rect 5288 796 5301 826
rect 5331 796 5344 826
rect 5359 808 5389 826
rect 5432 812 5446 826
rect 5482 812 5702 826
rect 5433 810 5446 812
rect 5399 798 5414 810
rect 5396 796 5418 798
rect 5423 796 5453 810
rect 5514 808 5667 812
rect 5496 796 5688 808
rect 5731 796 5761 810
rect 5767 796 5780 826
rect 5795 808 5825 826
rect 5868 796 5881 826
rect 3469 782 4623 796
rect 4736 782 5889 796
rect 3493 678 3506 782
rect 3551 760 3552 770
rect 3567 760 3580 770
rect 3551 756 3580 760
rect 3585 756 3615 782
rect 3633 768 3649 770
rect 3721 768 3774 782
rect 3722 766 3786 768
rect 3829 766 3844 782
rect 3893 779 3923 782
rect 3893 776 3929 779
rect 3859 768 3875 770
rect 3633 756 3648 760
rect 3551 754 3648 756
rect 3676 754 3844 766
rect 3860 756 3875 760
rect 3893 757 3932 776
rect 3951 770 3958 771
rect 3957 763 3958 770
rect 3941 760 3942 763
rect 3957 760 3970 763
rect 3893 756 3923 757
rect 3932 756 3938 757
rect 3941 756 3970 760
rect 3860 755 3970 756
rect 3860 754 3976 755
rect 3535 746 3586 754
rect 3535 734 3560 746
rect 3567 734 3586 746
rect 3617 746 3667 754
rect 3617 738 3633 746
rect 3640 744 3667 746
rect 3676 744 3897 754
rect 3640 734 3897 744
rect 3926 746 3976 754
rect 3926 737 3942 746
rect 3535 726 3586 734
rect 3633 726 3897 734
rect 3923 734 3942 737
rect 3949 734 3976 746
rect 3923 726 3976 734
rect 3551 718 3552 726
rect 3567 718 3580 726
rect 3551 710 3567 718
rect 3548 703 3567 706
rect 3548 694 3570 703
rect 3521 684 3570 694
rect 3521 678 3551 684
rect 3570 679 3575 684
rect 3493 662 3567 678
rect 3585 670 3615 726
rect 3650 716 3858 726
rect 3893 722 3938 726
rect 3941 725 3942 726
rect 3957 725 3970 726
rect 3676 686 3865 716
rect 3691 683 3865 686
rect 3684 680 3865 683
rect 3493 660 3506 662
rect 3521 660 3555 662
rect 3493 644 3567 660
rect 3594 656 3607 670
rect 3622 656 3638 672
rect 3684 667 3695 680
rect 3477 622 3478 638
rect 3493 622 3506 644
rect 3521 622 3551 644
rect 3594 640 3656 656
rect 3684 649 3695 665
rect 3700 660 3710 680
rect 3720 660 3734 680
rect 3737 667 3746 680
rect 3762 667 3771 680
rect 3700 649 3734 660
rect 3737 649 3746 665
rect 3762 649 3771 665
rect 3778 660 3788 680
rect 3798 660 3812 680
rect 3813 667 3824 680
rect 3778 649 3812 660
rect 3813 649 3824 665
rect 3870 656 3886 672
rect 3893 670 3923 722
rect 3957 718 3958 725
rect 3942 710 3958 718
rect 3929 678 3942 697
rect 3957 678 3987 694
rect 3929 662 4003 678
rect 3929 660 3942 662
rect 3957 660 3991 662
rect 3594 638 3607 640
rect 3622 638 3656 640
rect 3594 622 3656 638
rect 3700 633 3716 636
rect 3778 633 3808 644
rect 3856 640 3902 656
rect 3929 644 4003 660
rect 3856 638 3890 640
rect 3855 622 3902 638
rect 3929 622 3942 644
rect 3957 622 3987 644
rect 4014 622 4015 638
rect 4030 622 4043 782
rect 4073 678 4086 782
rect 4131 760 4132 770
rect 4147 760 4160 770
rect 4131 756 4160 760
rect 4165 756 4195 782
rect 4213 768 4229 770
rect 4301 768 4354 782
rect 4302 766 4366 768
rect 4409 766 4424 782
rect 4473 779 4503 782
rect 4473 776 4509 779
rect 4439 768 4455 770
rect 4213 756 4228 760
rect 4131 754 4228 756
rect 4256 754 4424 766
rect 4440 756 4455 760
rect 4473 757 4512 776
rect 4531 770 4538 771
rect 4537 763 4538 770
rect 4521 760 4522 763
rect 4537 760 4550 763
rect 4473 756 4503 757
rect 4512 756 4518 757
rect 4521 756 4550 760
rect 4440 755 4550 756
rect 4440 754 4556 755
rect 4115 746 4166 754
rect 4115 734 4140 746
rect 4147 734 4166 746
rect 4197 746 4247 754
rect 4197 738 4213 746
rect 4220 744 4247 746
rect 4256 744 4477 754
rect 4220 734 4477 744
rect 4506 746 4556 754
rect 4506 737 4522 746
rect 4115 726 4166 734
rect 4213 726 4477 734
rect 4503 734 4522 737
rect 4529 734 4556 746
rect 4503 726 4556 734
rect 4131 718 4132 726
rect 4147 718 4160 726
rect 4131 710 4147 718
rect 4128 703 4147 706
rect 4128 694 4150 703
rect 4101 684 4150 694
rect 4101 678 4131 684
rect 4150 679 4155 684
rect 4073 662 4147 678
rect 4165 670 4195 726
rect 4230 716 4438 726
rect 4473 722 4518 726
rect 4521 725 4522 726
rect 4537 725 4550 726
rect 4256 686 4445 716
rect 4271 683 4445 686
rect 4264 680 4445 683
rect 4073 660 4086 662
rect 4101 660 4135 662
rect 4073 644 4147 660
rect 4174 656 4187 670
rect 4202 656 4218 672
rect 4264 667 4275 680
rect 4057 622 4058 638
rect 4073 622 4086 644
rect 4101 622 4131 644
rect 4174 640 4236 656
rect 4264 649 4275 665
rect 4280 660 4290 680
rect 4300 660 4314 680
rect 4317 667 4326 680
rect 4342 667 4351 680
rect 4280 649 4314 660
rect 4317 649 4326 665
rect 4342 649 4351 665
rect 4358 660 4368 680
rect 4378 660 4392 680
rect 4393 667 4404 680
rect 4358 649 4392 660
rect 4393 649 4404 665
rect 4450 656 4466 672
rect 4473 670 4503 722
rect 4537 718 4538 725
rect 4522 710 4538 718
rect 4509 678 4522 697
rect 4537 678 4567 694
rect 4509 662 4583 678
rect 4509 660 4522 662
rect 4537 660 4571 662
rect 4174 638 4187 640
rect 4202 638 4236 640
rect 4174 622 4236 638
rect 4280 633 4296 636
rect 4358 633 4388 644
rect 4436 640 4482 656
rect 4509 644 4583 660
rect 4436 638 4470 640
rect 4435 622 4482 638
rect 4509 622 4522 644
rect 4537 622 4567 644
rect 4594 622 4595 638
rect 4610 622 4623 782
rect 4751 678 4764 782
rect 4809 760 4810 770
rect 4825 760 4838 770
rect 4809 756 4838 760
rect 4843 756 4873 782
rect 4891 768 4907 770
rect 4979 768 5032 782
rect 4980 766 5044 768
rect 5087 766 5102 782
rect 5151 779 5181 782
rect 5151 776 5187 779
rect 5117 768 5133 770
rect 4891 756 4906 760
rect 4809 754 4906 756
rect 4934 754 5102 766
rect 5118 756 5133 760
rect 5151 757 5190 776
rect 5209 770 5216 771
rect 5215 763 5216 770
rect 5199 760 5200 763
rect 5215 760 5228 763
rect 5151 756 5181 757
rect 5190 756 5196 757
rect 5199 756 5228 760
rect 5118 755 5228 756
rect 5118 754 5234 755
rect 4793 746 4844 754
rect 4793 734 4818 746
rect 4825 734 4844 746
rect 4875 746 4925 754
rect 4875 738 4891 746
rect 4898 744 4925 746
rect 4934 744 5155 754
rect 4898 734 5155 744
rect 5184 746 5234 754
rect 5184 737 5200 746
rect 4793 726 4844 734
rect 4891 726 5155 734
rect 5181 734 5200 737
rect 5207 734 5234 746
rect 5181 726 5234 734
rect 4809 718 4810 726
rect 4825 718 4838 726
rect 4809 710 4825 718
rect 4806 703 4825 706
rect 4806 694 4828 703
rect 4779 684 4828 694
rect 4779 678 4809 684
rect 4828 679 4833 684
rect 4751 662 4825 678
rect 4843 670 4873 726
rect 4908 716 5116 726
rect 5151 722 5196 726
rect 5199 725 5200 726
rect 5215 725 5228 726
rect 4934 686 5123 716
rect 4949 683 5123 686
rect 4942 680 5123 683
rect 4751 660 4764 662
rect 4779 660 4813 662
rect 4751 644 4825 660
rect 4852 656 4865 670
rect 4880 656 4896 672
rect 4942 667 4953 680
rect 4735 622 4736 638
rect 4751 622 4764 644
rect 4779 622 4809 644
rect 4852 640 4914 656
rect 4942 649 4953 665
rect 4958 660 4968 680
rect 4978 660 4992 680
rect 4995 667 5004 680
rect 5020 667 5029 680
rect 4958 649 4992 660
rect 4995 649 5004 665
rect 5020 649 5029 665
rect 5036 660 5046 680
rect 5056 660 5070 680
rect 5071 667 5082 680
rect 5036 649 5070 660
rect 5071 649 5082 665
rect 5128 656 5144 672
rect 5151 670 5181 722
rect 5215 718 5216 725
rect 5200 710 5216 718
rect 5187 678 5200 697
rect 5215 678 5245 694
rect 5187 662 5261 678
rect 5187 660 5200 662
rect 5215 660 5249 662
rect 4852 638 4865 640
rect 4880 638 4914 640
rect 4852 622 4914 638
rect 4958 633 4974 636
rect 5036 633 5066 644
rect 5114 640 5160 656
rect 5187 644 5261 660
rect 5114 638 5148 640
rect 5113 622 5160 638
rect 5187 622 5200 644
rect 5215 622 5245 644
rect 5272 622 5273 638
rect 5288 622 5301 782
rect 5331 678 5344 782
rect 5389 760 5390 770
rect 5405 760 5418 770
rect 5389 756 5418 760
rect 5423 756 5453 782
rect 5471 768 5487 770
rect 5559 768 5612 782
rect 5560 766 5624 768
rect 5667 766 5682 782
rect 5731 779 5761 782
rect 5731 776 5767 779
rect 5697 768 5713 770
rect 5471 756 5486 760
rect 5389 754 5486 756
rect 5514 754 5682 766
rect 5698 756 5713 760
rect 5731 757 5770 776
rect 5789 770 5796 771
rect 5795 763 5796 770
rect 5779 760 5780 763
rect 5795 760 5808 763
rect 5731 756 5761 757
rect 5770 756 5776 757
rect 5779 756 5808 760
rect 5698 755 5808 756
rect 5698 754 5814 755
rect 5373 746 5424 754
rect 5373 734 5398 746
rect 5405 734 5424 746
rect 5455 746 5505 754
rect 5455 738 5471 746
rect 5478 744 5505 746
rect 5514 744 5735 754
rect 5478 734 5735 744
rect 5764 746 5814 754
rect 5764 737 5780 746
rect 5373 726 5424 734
rect 5471 726 5735 734
rect 5761 734 5780 737
rect 5787 734 5814 746
rect 5761 726 5814 734
rect 5389 718 5390 726
rect 5405 718 5418 726
rect 5389 710 5405 718
rect 5386 703 5405 706
rect 5386 694 5408 703
rect 5359 684 5408 694
rect 5359 678 5389 684
rect 5408 679 5413 684
rect 5331 662 5405 678
rect 5423 670 5453 726
rect 5488 716 5696 726
rect 5731 722 5776 726
rect 5779 725 5780 726
rect 5795 725 5808 726
rect 5514 686 5703 716
rect 5529 683 5703 686
rect 5522 680 5703 683
rect 5331 660 5344 662
rect 5359 660 5393 662
rect 5331 644 5405 660
rect 5432 656 5445 670
rect 5460 656 5476 672
rect 5522 667 5533 680
rect 5315 622 5316 638
rect 5331 622 5344 644
rect 5359 622 5389 644
rect 5432 640 5494 656
rect 5522 649 5533 665
rect 5538 660 5548 680
rect 5558 660 5572 680
rect 5575 667 5584 680
rect 5600 667 5609 680
rect 5538 649 5572 660
rect 5575 649 5584 665
rect 5600 649 5609 665
rect 5616 660 5626 680
rect 5636 660 5650 680
rect 5651 667 5662 680
rect 5616 649 5650 660
rect 5651 649 5662 665
rect 5708 656 5724 672
rect 5731 670 5761 722
rect 5795 718 5796 725
rect 5780 710 5796 718
rect 5767 678 5780 697
rect 5795 678 5825 694
rect 5767 662 5841 678
rect 5767 660 5780 662
rect 5795 660 5829 662
rect 5432 638 5445 640
rect 5460 638 5494 640
rect 5432 622 5494 638
rect 5538 633 5554 636
rect 5616 633 5646 644
rect 5694 640 5740 656
rect 5767 644 5841 660
rect 5694 638 5728 640
rect 5693 622 5740 638
rect 5767 622 5780 644
rect 5795 622 5825 644
rect 5852 622 5853 638
rect 5868 622 5881 782
rect 3471 614 3512 622
rect 3471 588 3486 614
rect 3493 588 3512 614
rect 3576 610 3638 622
rect 3650 610 3725 622
rect 3783 610 3858 622
rect 3870 610 3901 622
rect 3907 610 3942 622
rect 3576 608 3738 610
rect 3471 580 3512 588
rect 3594 584 3607 608
rect 3622 606 3637 608
rect 3477 570 3478 580
rect 3493 570 3506 580
rect 3521 570 3551 584
rect 3594 570 3637 584
rect 3661 581 3668 588
rect 3671 584 3738 608
rect 3770 608 3942 610
rect 3740 586 3768 590
rect 3770 586 3850 608
rect 3871 606 3886 608
rect 3740 584 3850 586
rect 3671 580 3850 584
rect 3644 570 3674 580
rect 3676 570 3829 580
rect 3837 570 3867 580
rect 3871 570 3901 584
rect 3929 570 3942 608
rect 4014 614 4049 622
rect 4014 588 4015 614
rect 4022 588 4049 614
rect 3957 570 3987 584
rect 4014 580 4049 588
rect 4051 614 4092 622
rect 4051 588 4066 614
rect 4073 588 4092 614
rect 4156 610 4218 622
rect 4230 610 4305 622
rect 4363 610 4438 622
rect 4450 610 4481 622
rect 4487 610 4522 622
rect 4156 608 4318 610
rect 4051 580 4092 588
rect 4174 584 4187 608
rect 4202 606 4217 608
rect 4014 570 4015 580
rect 4030 570 4043 580
rect 4057 570 4058 580
rect 4073 570 4086 580
rect 4101 570 4131 584
rect 4174 570 4217 584
rect 4241 581 4248 588
rect 4251 584 4318 608
rect 4350 608 4522 610
rect 4320 586 4348 590
rect 4350 586 4430 608
rect 4451 606 4466 608
rect 4320 584 4430 586
rect 4251 580 4430 584
rect 4224 570 4254 580
rect 4256 570 4409 580
rect 4417 570 4447 580
rect 4451 570 4481 584
rect 4509 570 4522 608
rect 4594 614 4629 622
rect 4594 588 4595 614
rect 4602 588 4629 614
rect 4537 570 4567 584
rect 4594 580 4629 588
rect 4729 614 4770 622
rect 4729 588 4744 614
rect 4751 588 4770 614
rect 4834 610 4896 622
rect 4908 610 4983 622
rect 5041 610 5116 622
rect 5128 610 5159 622
rect 5165 610 5200 622
rect 4834 608 4996 610
rect 4729 580 4770 588
rect 4852 584 4865 608
rect 4880 606 4895 608
rect 4594 570 4595 580
rect 4610 570 4623 580
rect 3469 556 4623 570
rect 4735 570 4736 580
rect 4751 570 4764 580
rect 4779 570 4809 584
rect 4852 570 4895 584
rect 4919 581 4926 588
rect 4929 584 4996 608
rect 5028 608 5200 610
rect 4998 586 5026 590
rect 5028 586 5108 608
rect 5129 606 5144 608
rect 4998 584 5108 586
rect 4929 580 5108 584
rect 4902 570 4932 580
rect 4934 570 5087 580
rect 5095 570 5125 580
rect 5129 570 5159 584
rect 5187 570 5200 608
rect 5272 614 5307 622
rect 5272 588 5273 614
rect 5280 588 5307 614
rect 5215 570 5245 584
rect 5272 580 5307 588
rect 5309 614 5350 622
rect 5309 588 5324 614
rect 5331 588 5350 614
rect 5414 610 5476 622
rect 5488 610 5563 622
rect 5621 610 5696 622
rect 5708 610 5739 622
rect 5745 610 5780 622
rect 5414 608 5576 610
rect 5309 580 5350 588
rect 5432 584 5445 608
rect 5460 606 5475 608
rect 5272 570 5273 580
rect 5288 570 5301 580
rect 5315 570 5316 580
rect 5331 570 5344 580
rect 5359 570 5389 584
rect 5432 570 5475 584
rect 5499 581 5506 588
rect 5509 584 5576 608
rect 5608 608 5780 610
rect 5578 586 5606 590
rect 5608 586 5688 608
rect 5709 606 5724 608
rect 5578 584 5688 586
rect 5509 580 5688 584
rect 5482 570 5512 580
rect 5514 570 5667 580
rect 5675 570 5705 580
rect 5709 570 5739 584
rect 5767 570 5780 608
rect 5852 614 5887 622
rect 5852 588 5853 614
rect 5860 588 5887 614
rect 5795 570 5825 584
rect 5852 580 5887 588
rect 5852 570 5853 580
rect 5868 570 5881 580
rect 4735 564 5889 570
rect 4736 556 5889 564
rect 3493 526 3506 556
rect 3521 538 3551 556
rect 3594 542 3608 556
rect 3644 542 3864 556
rect 3595 540 3608 542
rect 3561 528 3576 540
rect 3558 526 3580 528
rect 3585 526 3615 540
rect 3676 538 3829 542
rect 3658 526 3850 538
rect 3893 526 3923 540
rect 3929 526 3942 556
rect 3957 538 3987 556
rect 4030 526 4043 556
rect 4073 526 4086 556
rect 4101 538 4131 556
rect 4174 542 4188 556
rect 4224 542 4444 556
rect 4175 540 4188 542
rect 4141 528 4156 540
rect 4138 526 4160 528
rect 4165 526 4195 540
rect 4256 538 4409 542
rect 4238 526 4430 538
rect 4473 526 4503 540
rect 4509 526 4522 556
rect 4537 538 4567 556
rect 4610 526 4623 556
rect 4751 526 4764 556
rect 4779 538 4809 556
rect 4852 542 4866 556
rect 4902 542 5122 556
rect 4853 540 4866 542
rect 4819 528 4834 540
rect 4816 526 4838 528
rect 4843 526 4873 540
rect 4934 538 5087 542
rect 4916 526 5108 538
rect 5151 526 5181 540
rect 5187 526 5200 556
rect 5215 538 5245 556
rect 5288 526 5301 556
rect 5331 526 5344 556
rect 5359 538 5389 556
rect 5432 542 5446 556
rect 5482 542 5702 556
rect 5433 540 5446 542
rect 5399 528 5414 540
rect 5396 526 5418 528
rect 5423 526 5453 540
rect 5514 538 5667 542
rect 5496 526 5688 538
rect 5731 526 5761 540
rect 5767 526 5780 556
rect 5795 538 5825 556
rect 5868 526 5881 556
rect 3469 512 4623 526
rect 4736 512 5889 526
rect 3493 408 3506 512
rect 3551 490 3552 500
rect 3567 490 3580 500
rect 3551 486 3580 490
rect 3585 486 3615 512
rect 3633 498 3649 500
rect 3721 498 3774 512
rect 3722 496 3786 498
rect 3829 496 3844 512
rect 3893 509 3923 512
rect 3893 506 3929 509
rect 3859 498 3875 500
rect 3633 486 3648 490
rect 3551 484 3648 486
rect 3676 484 3844 496
rect 3860 486 3875 490
rect 3893 487 3932 506
rect 3951 500 3958 501
rect 3957 493 3958 500
rect 3941 490 3942 493
rect 3957 490 3970 493
rect 3893 486 3923 487
rect 3932 486 3938 487
rect 3941 486 3970 490
rect 3860 485 3970 486
rect 3860 484 3976 485
rect 3535 476 3586 484
rect 3535 464 3560 476
rect 3567 464 3586 476
rect 3617 476 3667 484
rect 3617 468 3633 476
rect 3640 474 3667 476
rect 3676 474 3897 484
rect 3640 464 3897 474
rect 3926 476 3976 484
rect 3926 467 3942 476
rect 3535 456 3586 464
rect 3633 456 3897 464
rect 3923 464 3942 467
rect 3949 464 3976 476
rect 3923 456 3976 464
rect 3551 448 3552 456
rect 3567 448 3580 456
rect 3551 440 3567 448
rect 3548 433 3567 436
rect 3548 424 3570 433
rect 3521 414 3570 424
rect 3521 408 3551 414
rect 3570 409 3575 414
rect 3493 392 3567 408
rect 3585 400 3615 456
rect 3650 446 3858 456
rect 3893 452 3938 456
rect 3941 455 3942 456
rect 3957 455 3970 456
rect 3676 416 3865 446
rect 3691 413 3865 416
rect 3684 410 3865 413
rect 3493 390 3506 392
rect 3521 390 3555 392
rect 3493 374 3567 390
rect 3594 386 3607 400
rect 3622 386 3638 402
rect 3684 397 3695 410
rect 3477 352 3478 368
rect 3493 352 3506 374
rect 3521 352 3551 374
rect 3594 370 3656 386
rect 3684 379 3695 395
rect 3700 390 3710 410
rect 3720 390 3734 410
rect 3737 397 3746 410
rect 3762 397 3771 410
rect 3700 379 3734 390
rect 3737 379 3746 395
rect 3762 379 3771 395
rect 3778 390 3788 410
rect 3798 390 3812 410
rect 3813 397 3824 410
rect 3778 379 3812 390
rect 3813 379 3824 395
rect 3870 386 3886 402
rect 3893 400 3923 452
rect 3957 448 3958 455
rect 3942 440 3958 448
rect 3929 408 3942 427
rect 3957 408 3987 424
rect 3929 392 4003 408
rect 3929 390 3942 392
rect 3957 390 3991 392
rect 3594 368 3607 370
rect 3622 368 3656 370
rect 3594 352 3656 368
rect 3700 363 3716 366
rect 3778 363 3808 374
rect 3856 370 3902 386
rect 3929 374 4003 390
rect 3856 368 3890 370
rect 3855 352 3902 368
rect 3929 352 3942 374
rect 3957 352 3987 374
rect 4014 352 4015 368
rect 4030 352 4043 512
rect 4073 408 4086 512
rect 4131 490 4132 500
rect 4147 490 4160 500
rect 4131 486 4160 490
rect 4165 486 4195 512
rect 4213 498 4229 500
rect 4301 498 4354 512
rect 4302 496 4366 498
rect 4409 496 4424 512
rect 4473 509 4503 512
rect 4473 506 4509 509
rect 4439 498 4455 500
rect 4213 486 4228 490
rect 4131 484 4228 486
rect 4256 484 4424 496
rect 4440 486 4455 490
rect 4473 487 4512 506
rect 4531 500 4538 501
rect 4537 493 4538 500
rect 4521 490 4522 493
rect 4537 490 4550 493
rect 4473 486 4503 487
rect 4512 486 4518 487
rect 4521 486 4550 490
rect 4440 485 4550 486
rect 4440 484 4556 485
rect 4115 476 4166 484
rect 4115 464 4140 476
rect 4147 464 4166 476
rect 4197 476 4247 484
rect 4197 468 4213 476
rect 4220 474 4247 476
rect 4256 474 4477 484
rect 4220 464 4477 474
rect 4506 476 4556 484
rect 4506 467 4522 476
rect 4115 456 4166 464
rect 4213 456 4477 464
rect 4503 464 4522 467
rect 4529 464 4556 476
rect 4503 456 4556 464
rect 4131 448 4132 456
rect 4147 448 4160 456
rect 4131 440 4147 448
rect 4128 433 4147 436
rect 4128 424 4150 433
rect 4101 414 4150 424
rect 4101 408 4131 414
rect 4150 409 4155 414
rect 4073 392 4147 408
rect 4165 400 4195 456
rect 4230 446 4438 456
rect 4473 452 4518 456
rect 4521 455 4522 456
rect 4537 455 4550 456
rect 4256 416 4445 446
rect 4271 413 4445 416
rect 4264 410 4445 413
rect 4073 390 4086 392
rect 4101 390 4135 392
rect 4073 374 4147 390
rect 4174 386 4187 400
rect 4202 386 4218 402
rect 4264 397 4275 410
rect 4057 352 4058 368
rect 4073 352 4086 374
rect 4101 352 4131 374
rect 4174 370 4236 386
rect 4264 379 4275 395
rect 4280 390 4290 410
rect 4300 390 4314 410
rect 4317 397 4326 410
rect 4342 397 4351 410
rect 4280 379 4314 390
rect 4317 379 4326 395
rect 4342 379 4351 395
rect 4358 390 4368 410
rect 4378 390 4392 410
rect 4393 397 4404 410
rect 4358 379 4392 390
rect 4393 379 4404 395
rect 4450 386 4466 402
rect 4473 400 4503 452
rect 4537 448 4538 455
rect 4522 440 4538 448
rect 4509 408 4522 427
rect 4537 408 4567 424
rect 4509 392 4583 408
rect 4509 390 4522 392
rect 4537 390 4571 392
rect 4174 368 4187 370
rect 4202 368 4236 370
rect 4174 352 4236 368
rect 4280 363 4296 366
rect 4358 363 4388 374
rect 4436 370 4482 386
rect 4509 374 4583 390
rect 4436 368 4470 370
rect 4435 352 4482 368
rect 4509 352 4522 374
rect 4537 352 4567 374
rect 4594 352 4595 368
rect 4610 352 4623 512
rect 4751 408 4764 512
rect 4809 490 4810 500
rect 4825 490 4838 500
rect 4809 486 4838 490
rect 4843 486 4873 512
rect 4891 498 4907 500
rect 4979 498 5032 512
rect 4980 496 5044 498
rect 5087 496 5102 512
rect 5151 509 5181 512
rect 5151 506 5187 509
rect 5117 498 5133 500
rect 4891 486 4906 490
rect 4809 484 4906 486
rect 4934 484 5102 496
rect 5118 486 5133 490
rect 5151 487 5190 506
rect 5209 500 5216 501
rect 5215 493 5216 500
rect 5199 490 5200 493
rect 5215 490 5228 493
rect 5151 486 5181 487
rect 5190 486 5196 487
rect 5199 486 5228 490
rect 5118 485 5228 486
rect 5118 484 5234 485
rect 4793 476 4844 484
rect 4793 464 4818 476
rect 4825 464 4844 476
rect 4875 476 4925 484
rect 4875 468 4891 476
rect 4898 474 4925 476
rect 4934 474 5155 484
rect 4898 464 5155 474
rect 5184 476 5234 484
rect 5184 467 5200 476
rect 4793 456 4844 464
rect 4891 456 5155 464
rect 5181 464 5200 467
rect 5207 464 5234 476
rect 5181 456 5234 464
rect 4809 448 4810 456
rect 4825 448 4838 456
rect 4809 440 4825 448
rect 4806 433 4825 436
rect 4806 424 4828 433
rect 4779 414 4828 424
rect 4779 408 4809 414
rect 4828 409 4833 414
rect 4751 392 4825 408
rect 4843 400 4873 456
rect 4908 446 5116 456
rect 5151 452 5196 456
rect 5199 455 5200 456
rect 5215 455 5228 456
rect 4934 416 5123 446
rect 4949 413 5123 416
rect 4942 410 5123 413
rect 4751 390 4764 392
rect 4779 390 4813 392
rect 4751 374 4825 390
rect 4852 386 4865 400
rect 4880 386 4896 402
rect 4942 397 4953 410
rect 4735 352 4736 368
rect 4751 352 4764 374
rect 4779 352 4809 374
rect 4852 370 4914 386
rect 4942 379 4953 395
rect 4958 390 4968 410
rect 4978 390 4992 410
rect 4995 397 5004 410
rect 5020 397 5029 410
rect 4958 379 4992 390
rect 4995 379 5004 395
rect 5020 379 5029 395
rect 5036 390 5046 410
rect 5056 390 5070 410
rect 5071 397 5082 410
rect 5036 379 5070 390
rect 5071 379 5082 395
rect 5128 386 5144 402
rect 5151 400 5181 452
rect 5215 448 5216 455
rect 5200 440 5216 448
rect 5187 408 5200 427
rect 5215 408 5245 424
rect 5187 392 5261 408
rect 5187 390 5200 392
rect 5215 390 5249 392
rect 4852 368 4865 370
rect 4880 368 4914 370
rect 4852 352 4914 368
rect 4958 363 4974 366
rect 5036 363 5066 374
rect 5114 370 5160 386
rect 5187 374 5261 390
rect 5114 368 5148 370
rect 5113 352 5160 368
rect 5187 352 5200 374
rect 5215 352 5245 374
rect 5272 352 5273 368
rect 5288 352 5301 512
rect 5331 408 5344 512
rect 5389 490 5390 500
rect 5405 490 5418 500
rect 5389 486 5418 490
rect 5423 486 5453 512
rect 5471 498 5487 500
rect 5559 498 5612 512
rect 5560 496 5624 498
rect 5667 496 5682 512
rect 5731 509 5761 512
rect 5731 506 5767 509
rect 5697 498 5713 500
rect 5471 486 5486 490
rect 5389 484 5486 486
rect 5514 484 5682 496
rect 5698 486 5713 490
rect 5731 487 5770 506
rect 5789 500 5796 501
rect 5795 493 5796 500
rect 5779 490 5780 493
rect 5795 490 5808 493
rect 5731 486 5761 487
rect 5770 486 5776 487
rect 5779 486 5808 490
rect 5698 485 5808 486
rect 5698 484 5814 485
rect 5373 476 5424 484
rect 5373 464 5398 476
rect 5405 464 5424 476
rect 5455 476 5505 484
rect 5455 468 5471 476
rect 5478 474 5505 476
rect 5514 474 5735 484
rect 5478 464 5735 474
rect 5764 476 5814 484
rect 5764 467 5780 476
rect 5373 456 5424 464
rect 5471 456 5735 464
rect 5761 464 5780 467
rect 5787 464 5814 476
rect 5761 456 5814 464
rect 5389 448 5390 456
rect 5405 448 5418 456
rect 5389 440 5405 448
rect 5386 433 5405 436
rect 5386 424 5408 433
rect 5359 414 5408 424
rect 5359 408 5389 414
rect 5408 409 5413 414
rect 5331 392 5405 408
rect 5423 400 5453 456
rect 5488 446 5696 456
rect 5731 452 5776 456
rect 5779 455 5780 456
rect 5795 455 5808 456
rect 5514 416 5703 446
rect 5529 413 5703 416
rect 5522 410 5703 413
rect 5331 390 5344 392
rect 5359 390 5393 392
rect 5331 374 5405 390
rect 5432 386 5445 400
rect 5460 386 5476 402
rect 5522 397 5533 410
rect 5315 352 5316 368
rect 5331 352 5344 374
rect 5359 352 5389 374
rect 5432 370 5494 386
rect 5522 379 5533 395
rect 5538 390 5548 410
rect 5558 390 5572 410
rect 5575 397 5584 410
rect 5600 397 5609 410
rect 5538 379 5572 390
rect 5575 379 5584 395
rect 5600 379 5609 395
rect 5616 390 5626 410
rect 5636 390 5650 410
rect 5651 397 5662 410
rect 5616 379 5650 390
rect 5651 379 5662 395
rect 5708 386 5724 402
rect 5731 400 5761 452
rect 5795 448 5796 455
rect 5780 440 5796 448
rect 5767 408 5780 427
rect 5795 408 5825 424
rect 5767 392 5841 408
rect 5767 390 5780 392
rect 5795 390 5829 392
rect 5432 368 5445 370
rect 5460 368 5494 370
rect 5432 352 5494 368
rect 5538 363 5554 366
rect 5616 363 5646 374
rect 5694 370 5740 386
rect 5767 374 5841 390
rect 5694 368 5728 370
rect 5693 352 5740 368
rect 5767 352 5780 374
rect 5795 352 5825 374
rect 5852 352 5853 368
rect 5868 352 5881 512
rect 3471 344 3512 352
rect 3471 318 3486 344
rect 3493 318 3512 344
rect 3576 340 3638 352
rect 3650 340 3725 352
rect 3783 340 3858 352
rect 3870 340 3901 352
rect 3907 340 3942 352
rect 3576 338 3738 340
rect 3471 310 3512 318
rect 3594 314 3607 338
rect 3622 336 3637 338
rect 3477 300 3478 310
rect 3493 300 3506 310
rect 3521 300 3551 314
rect 3594 300 3637 314
rect 3661 311 3668 318
rect 3671 314 3738 338
rect 3770 338 3942 340
rect 3740 316 3768 320
rect 3770 316 3850 338
rect 3871 336 3886 338
rect 3740 314 3850 316
rect 3671 310 3850 314
rect 3644 300 3674 310
rect 3676 300 3829 310
rect 3837 300 3867 310
rect 3871 300 3901 314
rect 3929 300 3942 338
rect 4014 344 4049 352
rect 4014 318 4015 344
rect 4022 318 4049 344
rect 3957 300 3987 314
rect 4014 310 4049 318
rect 4051 344 4092 352
rect 4051 318 4066 344
rect 4073 318 4092 344
rect 4156 340 4218 352
rect 4230 340 4305 352
rect 4363 340 4438 352
rect 4450 340 4481 352
rect 4487 340 4522 352
rect 4156 338 4318 340
rect 4051 310 4092 318
rect 4174 314 4187 338
rect 4202 336 4217 338
rect 4014 300 4015 310
rect 4030 300 4043 310
rect 4057 300 4058 310
rect 4073 300 4086 310
rect 4101 300 4131 314
rect 4174 300 4217 314
rect 4241 311 4248 318
rect 4251 314 4318 338
rect 4350 338 4522 340
rect 4320 316 4348 320
rect 4350 316 4430 338
rect 4451 336 4466 338
rect 4320 314 4430 316
rect 4251 310 4430 314
rect 4224 300 4254 310
rect 4256 300 4409 310
rect 4417 300 4447 310
rect 4451 300 4481 314
rect 4509 300 4522 338
rect 4594 344 4629 352
rect 4594 318 4595 344
rect 4602 318 4629 344
rect 4537 300 4567 314
rect 4594 310 4629 318
rect 4729 344 4770 352
rect 4729 318 4744 344
rect 4751 318 4770 344
rect 4834 340 4896 352
rect 4908 340 4983 352
rect 5041 340 5116 352
rect 5128 340 5159 352
rect 5165 340 5200 352
rect 4834 338 4996 340
rect 4729 310 4770 318
rect 4852 314 4865 338
rect 4880 336 4895 338
rect 4594 300 4595 310
rect 4610 300 4623 310
rect 3469 286 4623 300
rect 4735 300 4736 310
rect 4751 300 4764 310
rect 4779 300 4809 314
rect 4852 300 4895 314
rect 4919 311 4926 318
rect 4929 314 4996 338
rect 5028 338 5200 340
rect 4998 316 5026 320
rect 5028 316 5108 338
rect 5129 336 5144 338
rect 4998 314 5108 316
rect 4929 310 5108 314
rect 4902 300 4932 310
rect 4934 300 5087 310
rect 5095 300 5125 310
rect 5129 300 5159 314
rect 5187 300 5200 338
rect 5272 344 5307 352
rect 5272 318 5273 344
rect 5280 318 5307 344
rect 5215 300 5245 314
rect 5272 310 5307 318
rect 5309 344 5350 352
rect 5309 318 5324 344
rect 5331 318 5350 344
rect 5414 340 5476 352
rect 5488 340 5563 352
rect 5621 340 5696 352
rect 5708 340 5739 352
rect 5745 340 5780 352
rect 5414 338 5576 340
rect 5309 310 5350 318
rect 5432 314 5445 338
rect 5460 336 5475 338
rect 5272 300 5273 310
rect 5288 300 5301 310
rect 5315 300 5316 310
rect 5331 300 5344 310
rect 5359 300 5389 314
rect 5432 300 5475 314
rect 5499 311 5506 318
rect 5509 314 5576 338
rect 5608 338 5780 340
rect 5578 316 5606 320
rect 5608 316 5688 338
rect 5709 336 5724 338
rect 5578 314 5688 316
rect 5509 310 5688 314
rect 5482 300 5512 310
rect 5514 300 5667 310
rect 5675 300 5705 310
rect 5709 300 5739 314
rect 5767 300 5780 338
rect 5852 344 5887 352
rect 5852 318 5853 344
rect 5860 318 5887 344
rect 5795 300 5825 314
rect 5852 310 5887 318
rect 5852 300 5853 310
rect 5868 300 5881 310
rect 4735 294 5889 300
rect 4736 286 5889 294
rect 3493 256 3506 286
rect 3521 268 3551 286
rect 3594 272 3608 286
rect 3644 272 3864 286
rect 3595 270 3608 272
rect 3561 258 3576 270
rect 3558 256 3580 258
rect 3585 256 3615 270
rect 3676 268 3829 272
rect 3658 256 3850 268
rect 3893 256 3923 270
rect 3929 256 3942 286
rect 3957 268 3987 286
rect 4030 256 4043 286
rect 4073 256 4086 286
rect 4101 268 4131 286
rect 4174 272 4188 286
rect 4224 272 4444 286
rect 4175 270 4188 272
rect 4141 258 4156 270
rect 4138 256 4160 258
rect 4165 256 4195 270
rect 4256 268 4409 272
rect 4238 256 4430 268
rect 4473 256 4503 270
rect 4509 256 4522 286
rect 4537 268 4567 286
rect 4610 256 4623 286
rect 4751 256 4764 286
rect 4779 268 4809 286
rect 4852 272 4866 286
rect 4902 272 5122 286
rect 4853 270 4866 272
rect 4819 258 4834 270
rect 4816 256 4838 258
rect 4843 256 4873 270
rect 4934 268 5087 272
rect 4916 256 5108 268
rect 5151 256 5181 270
rect 5187 256 5200 286
rect 5215 268 5245 286
rect 5288 256 5301 286
rect 5331 256 5344 286
rect 5359 268 5389 286
rect 5432 272 5446 286
rect 5482 272 5702 286
rect 5433 270 5446 272
rect 5399 258 5414 270
rect 5396 256 5418 258
rect 5423 256 5453 270
rect 5514 268 5667 272
rect 5496 256 5688 268
rect 5731 256 5761 270
rect 5767 256 5780 286
rect 5795 268 5825 286
rect 5868 256 5881 286
rect 3469 242 4623 256
rect 4736 242 5889 256
rect 3493 138 3506 242
rect 3551 220 3552 230
rect 3567 220 3580 230
rect 3551 216 3580 220
rect 3585 216 3615 242
rect 3633 228 3649 230
rect 3721 228 3774 242
rect 3722 226 3786 228
rect 3633 216 3648 220
rect 3551 214 3648 216
rect 3535 206 3586 214
rect 3535 194 3560 206
rect 3567 194 3586 206
rect 3617 206 3667 214
rect 3617 198 3633 206
rect 3640 204 3667 206
rect 3676 206 3691 210
rect 3738 206 3770 226
rect 3829 214 3844 242
rect 3893 239 3923 242
rect 3893 236 3929 239
rect 3859 228 3875 230
rect 3860 216 3875 220
rect 3893 217 3932 236
rect 3951 230 3958 231
rect 3957 223 3958 230
rect 3941 220 3942 223
rect 3957 220 3970 223
rect 3893 216 3923 217
rect 3932 216 3938 217
rect 3941 216 3970 220
rect 3860 215 3970 216
rect 3860 214 3976 215
rect 3829 206 3897 214
rect 3676 204 3745 206
rect 3763 204 3897 206
rect 3640 200 3712 204
rect 3640 198 3765 200
rect 3640 194 3712 198
rect 3535 186 3586 194
rect 3633 190 3712 194
rect 3793 190 3897 204
rect 3926 206 3976 214
rect 3926 197 3942 206
rect 3633 186 3897 190
rect 3923 194 3942 197
rect 3949 194 3976 206
rect 3923 186 3976 194
rect 3551 178 3552 186
rect 3567 178 3580 186
rect 3551 170 3567 178
rect 3548 163 3567 166
rect 3548 154 3570 163
rect 3521 144 3570 154
rect 3521 138 3551 144
rect 3570 139 3575 144
rect 3493 122 3567 138
rect 3585 130 3615 186
rect 3650 176 3858 186
rect 3893 182 3938 186
rect 3941 185 3942 186
rect 3957 185 3970 186
rect 3817 172 3865 176
rect 3700 150 3730 159
rect 3793 152 3808 159
rect 3829 150 3865 172
rect 3676 146 3865 150
rect 3691 143 3865 146
rect 3684 140 3865 143
rect 3493 120 3506 122
rect 3521 120 3555 122
rect 3493 104 3567 120
rect 3594 116 3607 130
rect 3622 116 3638 132
rect 3684 127 3695 140
rect 3477 82 3478 98
rect 3493 82 3506 104
rect 3521 82 3551 104
rect 3594 100 3656 116
rect 3684 109 3695 125
rect 3700 120 3710 140
rect 3720 120 3734 140
rect 3737 127 3746 140
rect 3762 127 3771 140
rect 3700 109 3734 120
rect 3737 109 3745 125
rect 3762 109 3771 125
rect 3778 120 3788 140
rect 3798 120 3812 140
rect 3813 127 3824 140
rect 3778 109 3812 120
rect 3813 109 3824 125
rect 3870 116 3886 132
rect 3893 130 3923 182
rect 3957 178 3958 185
rect 3942 170 3958 178
rect 3929 138 3942 157
rect 3957 138 3987 154
rect 3929 122 4003 138
rect 3929 120 3942 122
rect 3957 120 3991 122
rect 3594 98 3607 100
rect 3622 98 3656 100
rect 3594 82 3656 98
rect 3700 93 3713 96
rect 3778 93 3808 104
rect 3856 100 3902 116
rect 3929 104 4003 120
rect 3856 98 3890 100
rect 3855 82 3902 98
rect 3929 82 3942 104
rect 3957 82 3987 104
rect 4014 82 4015 98
rect 4030 82 4043 242
rect 4073 138 4086 242
rect 4131 220 4132 230
rect 4147 220 4160 230
rect 4131 216 4160 220
rect 4165 216 4195 242
rect 4213 228 4229 230
rect 4301 228 4354 242
rect 4302 226 4366 228
rect 4213 216 4228 220
rect 4131 214 4228 216
rect 4115 206 4166 214
rect 4115 194 4140 206
rect 4147 194 4166 206
rect 4197 206 4247 214
rect 4197 198 4213 206
rect 4220 204 4247 206
rect 4256 206 4271 210
rect 4318 206 4350 226
rect 4409 214 4424 242
rect 4473 239 4503 242
rect 4473 236 4509 239
rect 4439 228 4455 230
rect 4440 216 4455 220
rect 4473 217 4512 236
rect 4531 230 4538 231
rect 4537 223 4538 230
rect 4521 220 4522 223
rect 4537 220 4550 223
rect 4473 216 4503 217
rect 4512 216 4518 217
rect 4521 216 4550 220
rect 4440 215 4550 216
rect 4440 214 4556 215
rect 4409 206 4477 214
rect 4256 204 4325 206
rect 4343 204 4477 206
rect 4220 200 4292 204
rect 4220 198 4345 200
rect 4220 194 4292 198
rect 4115 186 4166 194
rect 4213 190 4292 194
rect 4373 190 4477 204
rect 4506 206 4556 214
rect 4506 197 4522 206
rect 4213 186 4477 190
rect 4503 194 4522 197
rect 4529 194 4556 206
rect 4503 186 4556 194
rect 4131 178 4132 186
rect 4147 178 4160 186
rect 4131 170 4147 178
rect 4128 163 4147 166
rect 4128 154 4150 163
rect 4101 144 4150 154
rect 4101 138 4131 144
rect 4150 139 4155 144
rect 4073 122 4147 138
rect 4165 130 4195 186
rect 4230 176 4438 186
rect 4473 182 4518 186
rect 4521 185 4522 186
rect 4537 185 4550 186
rect 4397 172 4445 176
rect 4280 150 4310 159
rect 4373 152 4388 159
rect 4409 150 4445 172
rect 4256 146 4445 150
rect 4271 143 4445 146
rect 4264 140 4445 143
rect 4073 120 4086 122
rect 4101 120 4135 122
rect 4073 104 4147 120
rect 4174 116 4187 130
rect 4202 116 4218 132
rect 4264 127 4275 140
rect 4057 82 4058 98
rect 4073 82 4086 104
rect 4101 82 4131 104
rect 4174 100 4236 116
rect 4264 109 4275 125
rect 4280 120 4290 140
rect 4300 120 4314 140
rect 4317 127 4326 140
rect 4342 127 4351 140
rect 4280 109 4314 120
rect 4317 109 4325 125
rect 4342 109 4351 125
rect 4358 120 4368 140
rect 4378 120 4392 140
rect 4393 127 4404 140
rect 4358 109 4392 120
rect 4393 109 4404 125
rect 4450 116 4466 132
rect 4473 130 4503 182
rect 4537 178 4538 185
rect 4522 170 4538 178
rect 4509 138 4522 157
rect 4537 138 4567 154
rect 4509 122 4583 138
rect 4509 120 4522 122
rect 4537 120 4571 122
rect 4174 98 4187 100
rect 4202 98 4236 100
rect 4174 82 4236 98
rect 4280 93 4293 96
rect 4358 93 4388 104
rect 4436 100 4482 116
rect 4509 104 4583 120
rect 4436 98 4470 100
rect 4435 82 4482 98
rect 4509 82 4522 104
rect 4537 82 4567 104
rect 4594 82 4595 98
rect 4610 82 4623 242
rect 4751 138 4764 242
rect 4809 220 4810 230
rect 4825 220 4838 230
rect 4809 216 4838 220
rect 4843 216 4873 242
rect 4891 228 4907 230
rect 4979 228 5032 242
rect 4980 226 5044 228
rect 4891 216 4906 220
rect 4809 214 4906 216
rect 4793 206 4844 214
rect 4793 194 4818 206
rect 4825 194 4844 206
rect 4875 206 4925 214
rect 4875 198 4891 206
rect 4898 204 4925 206
rect 4934 206 4949 210
rect 4996 206 5028 226
rect 5087 214 5102 242
rect 5151 239 5181 242
rect 5151 236 5187 239
rect 5117 228 5133 230
rect 5118 216 5133 220
rect 5151 217 5190 236
rect 5209 230 5216 231
rect 5215 223 5216 230
rect 5199 220 5200 223
rect 5215 220 5228 223
rect 5151 216 5181 217
rect 5190 216 5196 217
rect 5199 216 5228 220
rect 5118 215 5228 216
rect 5118 214 5234 215
rect 5087 206 5155 214
rect 4934 204 5003 206
rect 5021 204 5155 206
rect 4898 200 4970 204
rect 4898 198 5023 200
rect 4898 194 4970 198
rect 4793 186 4844 194
rect 4891 190 4970 194
rect 5051 190 5155 204
rect 5184 206 5234 214
rect 5184 197 5200 206
rect 4891 186 5155 190
rect 5181 194 5200 197
rect 5207 194 5234 206
rect 5181 186 5234 194
rect 4809 178 4810 186
rect 4825 178 4838 186
rect 4809 170 4825 178
rect 4806 163 4825 166
rect 4806 154 4828 163
rect 4779 144 4828 154
rect 4779 138 4809 144
rect 4828 139 4833 144
rect 4751 122 4825 138
rect 4843 130 4873 186
rect 4908 176 5116 186
rect 5151 182 5196 186
rect 5199 185 5200 186
rect 5215 185 5228 186
rect 5075 172 5123 176
rect 4958 150 4988 159
rect 5051 152 5066 159
rect 5087 150 5123 172
rect 4934 146 5123 150
rect 4949 143 5123 146
rect 4942 140 5123 143
rect 4751 120 4764 122
rect 4779 120 4813 122
rect 4751 104 4825 120
rect 4852 116 4865 130
rect 4880 116 4896 132
rect 4942 127 4953 140
rect 4735 82 4736 98
rect 4751 82 4764 104
rect 4779 82 4809 104
rect 4852 100 4914 116
rect 4942 109 4953 125
rect 4958 120 4968 140
rect 4978 120 4992 140
rect 4995 127 5004 140
rect 5020 127 5029 140
rect 4958 109 4992 120
rect 4995 109 5003 125
rect 5020 109 5029 125
rect 5036 120 5046 140
rect 5056 120 5070 140
rect 5071 127 5082 140
rect 5036 109 5070 120
rect 5071 109 5082 125
rect 5128 116 5144 132
rect 5151 130 5181 182
rect 5215 178 5216 185
rect 5200 170 5216 178
rect 5187 138 5200 157
rect 5215 138 5245 154
rect 5187 122 5261 138
rect 5187 120 5200 122
rect 5215 120 5249 122
rect 4852 98 4865 100
rect 4880 98 4914 100
rect 4852 82 4914 98
rect 4958 93 4971 96
rect 5036 93 5066 104
rect 5114 100 5160 116
rect 5187 104 5261 120
rect 5114 98 5148 100
rect 5113 82 5160 98
rect 5187 82 5200 104
rect 5215 82 5245 104
rect 5272 82 5273 98
rect 5288 82 5301 242
rect 5331 138 5344 242
rect 5389 220 5390 230
rect 5405 220 5418 230
rect 5389 216 5418 220
rect 5423 216 5453 242
rect 5471 228 5487 230
rect 5559 228 5612 242
rect 5560 226 5624 228
rect 5471 216 5486 220
rect 5389 214 5486 216
rect 5373 206 5424 214
rect 5373 194 5398 206
rect 5405 194 5424 206
rect 5455 206 5505 214
rect 5455 198 5471 206
rect 5478 204 5505 206
rect 5514 206 5529 210
rect 5576 206 5608 226
rect 5667 214 5682 242
rect 5731 239 5761 242
rect 5731 236 5767 239
rect 5697 228 5713 230
rect 5698 216 5713 220
rect 5731 217 5770 236
rect 5789 230 5796 231
rect 5795 223 5796 230
rect 5779 220 5780 223
rect 5795 220 5808 223
rect 5731 216 5761 217
rect 5770 216 5776 217
rect 5779 216 5808 220
rect 5698 215 5808 216
rect 5698 214 5814 215
rect 5667 206 5735 214
rect 5514 204 5583 206
rect 5601 204 5735 206
rect 5478 200 5550 204
rect 5478 198 5603 200
rect 5478 194 5550 198
rect 5373 186 5424 194
rect 5471 190 5550 194
rect 5631 190 5735 204
rect 5764 206 5814 214
rect 5764 197 5780 206
rect 5471 186 5735 190
rect 5761 194 5780 197
rect 5787 194 5814 206
rect 5761 186 5814 194
rect 5389 178 5390 186
rect 5405 178 5418 186
rect 5389 170 5405 178
rect 5386 163 5405 166
rect 5386 154 5408 163
rect 5359 144 5408 154
rect 5359 138 5389 144
rect 5408 139 5413 144
rect 5331 122 5405 138
rect 5423 130 5453 186
rect 5488 176 5696 186
rect 5731 182 5776 186
rect 5779 185 5780 186
rect 5795 185 5808 186
rect 5655 172 5703 176
rect 5538 150 5568 159
rect 5631 152 5646 159
rect 5667 150 5703 172
rect 5514 146 5703 150
rect 5529 143 5703 146
rect 5522 140 5703 143
rect 5331 120 5344 122
rect 5359 120 5393 122
rect 5331 104 5405 120
rect 5432 116 5445 130
rect 5460 116 5476 132
rect 5522 127 5533 140
rect 5315 82 5316 98
rect 5331 82 5344 104
rect 5359 82 5389 104
rect 5432 100 5494 116
rect 5522 109 5533 125
rect 5538 120 5548 140
rect 5558 120 5572 140
rect 5575 127 5584 140
rect 5600 127 5609 140
rect 5538 109 5572 120
rect 5575 109 5583 125
rect 5600 109 5609 125
rect 5616 120 5626 140
rect 5636 120 5650 140
rect 5651 127 5662 140
rect 5616 109 5650 120
rect 5651 109 5662 125
rect 5708 116 5724 132
rect 5731 130 5761 182
rect 5795 178 5796 185
rect 5780 170 5796 178
rect 5767 138 5780 157
rect 5795 138 5825 154
rect 5767 122 5841 138
rect 5767 120 5780 122
rect 5795 120 5829 122
rect 5432 98 5445 100
rect 5460 98 5494 100
rect 5432 82 5494 98
rect 5538 93 5551 96
rect 5616 93 5646 104
rect 5694 100 5740 116
rect 5767 104 5841 120
rect 5694 98 5728 100
rect 5693 82 5740 98
rect 5767 82 5780 104
rect 5795 82 5825 104
rect 5852 82 5853 98
rect 5868 82 5881 242
rect 3471 74 3512 82
rect 3471 48 3486 74
rect 3493 48 3512 74
rect 3576 70 3638 82
rect 3650 70 3725 82
rect 3783 70 3858 82
rect 3870 70 3901 82
rect 3907 70 3942 82
rect 3576 68 3738 70
rect 3471 40 3512 48
rect 3594 40 3607 68
rect 3622 66 3637 68
rect 3661 41 3668 48
rect 3671 40 3738 68
rect 3770 68 3942 70
rect 3740 46 3768 50
rect 3770 46 3850 68
rect 3871 66 3886 68
rect 3740 44 3850 46
rect 3740 40 3768 44
rect 3770 40 3850 44
rect 3477 30 3478 40
rect 3493 30 3506 40
rect 3521 30 3551 40
rect 3594 30 3637 40
rect 3644 30 3652 40
rect 3671 32 3674 40
rect 3738 32 3770 40
rect 3671 30 3837 32
rect 3856 30 3867 40
rect 3871 30 3901 40
rect 3929 30 3942 68
rect 4014 74 4049 82
rect 4014 48 4015 74
rect 4022 48 4049 74
rect 4014 40 4049 48
rect 4051 74 4092 82
rect 4051 48 4066 74
rect 4073 48 4092 74
rect 4156 70 4218 82
rect 4230 70 4305 82
rect 4363 70 4438 82
rect 4450 70 4481 82
rect 4487 70 4522 82
rect 4156 68 4318 70
rect 4051 40 4092 48
rect 4174 40 4187 68
rect 4202 66 4217 68
rect 4241 41 4248 48
rect 4251 40 4318 68
rect 4350 68 4522 70
rect 4320 46 4348 50
rect 4350 46 4430 68
rect 4451 66 4466 68
rect 4320 44 4430 46
rect 4320 40 4348 44
rect 4350 40 4430 44
rect 3957 30 3987 40
rect 4014 30 4015 40
rect 4030 30 4043 40
rect 4057 30 4058 40
rect 4073 30 4086 40
rect 4101 30 4131 40
rect 4174 30 4217 40
rect 4224 30 4232 40
rect 4251 32 4254 40
rect 4318 32 4350 40
rect 4251 30 4417 32
rect 4436 30 4447 40
rect 4451 30 4481 40
rect 4509 30 4522 68
rect 4594 74 4629 82
rect 4594 48 4595 74
rect 4602 48 4629 74
rect 4594 40 4629 48
rect 4729 74 4770 82
rect 4729 48 4744 74
rect 4751 48 4770 74
rect 4834 70 4896 82
rect 4908 70 4983 82
rect 5041 70 5116 82
rect 5128 70 5159 82
rect 5165 70 5200 82
rect 4834 68 4996 70
rect 4729 40 4770 48
rect 4852 40 4865 68
rect 4880 66 4895 68
rect 4919 41 4926 48
rect 4929 40 4996 68
rect 5028 68 5200 70
rect 4998 46 5026 50
rect 5028 46 5108 68
rect 5129 66 5144 68
rect 4998 44 5108 46
rect 4998 40 5026 44
rect 5028 40 5108 44
rect 4537 30 4567 40
rect 4594 30 4595 40
rect 4610 30 4623 40
rect 3469 16 4623 30
rect 4735 30 4736 40
rect 4751 30 4764 40
rect 4779 30 4809 40
rect 4852 30 4895 40
rect 4902 30 4910 40
rect 4929 32 4932 40
rect 4996 32 5028 40
rect 4929 30 5095 32
rect 5114 30 5125 40
rect 5129 30 5159 40
rect 5187 30 5200 68
rect 5272 74 5307 82
rect 5272 48 5273 74
rect 5280 48 5307 74
rect 5272 40 5307 48
rect 5309 74 5350 82
rect 5309 48 5324 74
rect 5331 48 5350 74
rect 5414 70 5476 82
rect 5488 70 5563 82
rect 5621 70 5696 82
rect 5708 70 5739 82
rect 5745 70 5780 82
rect 5414 68 5576 70
rect 5309 40 5350 48
rect 5432 40 5445 68
rect 5460 66 5475 68
rect 5499 41 5506 48
rect 5509 40 5576 68
rect 5608 68 5780 70
rect 5578 46 5606 50
rect 5608 46 5688 68
rect 5709 66 5724 68
rect 5578 44 5688 46
rect 5578 40 5606 44
rect 5608 40 5688 44
rect 5215 30 5245 40
rect 5272 30 5273 40
rect 5288 30 5301 40
rect 5315 30 5316 40
rect 5331 30 5344 40
rect 5359 30 5389 40
rect 5432 30 5475 40
rect 5482 30 5490 40
rect 5509 32 5512 40
rect 5576 32 5608 40
rect 5509 30 5675 32
rect 5694 30 5705 40
rect 5709 30 5739 40
rect 5767 30 5780 68
rect 5852 74 5887 82
rect 5852 48 5853 74
rect 5860 48 5887 74
rect 5852 40 5887 48
rect 5795 30 5825 40
rect 5852 30 5853 40
rect 5868 30 5881 40
rect 4735 24 5889 30
rect 4736 16 5889 24
rect 3493 2 3506 16
rect 3521 -2 3551 16
rect 3594 2 3607 16
rect 3644 3 3652 16
rect 3685 3 3823 16
rect 3856 3 3864 16
rect 3721 2 3772 3
rect 3929 2 3942 16
rect 3722 0 3786 2
rect 3957 -2 3987 16
rect 4030 2 4043 16
rect 4073 2 4086 16
rect 4101 -2 4131 16
rect 4174 2 4187 16
rect 4224 3 4232 16
rect 4265 3 4403 16
rect 4436 3 4444 16
rect 4301 2 4352 3
rect 4509 2 4522 16
rect 4302 0 4366 2
rect 4537 -2 4567 16
rect 4610 2 4623 16
rect 4751 2 4764 16
rect 4779 -2 4809 16
rect 4852 2 4865 16
rect 4902 3 4910 16
rect 4943 3 5081 16
rect 5114 3 5122 16
rect 4979 2 5030 3
rect 5187 2 5200 16
rect 4980 0 5044 2
rect 5215 -2 5245 16
rect 5288 2 5301 16
rect 5331 2 5344 16
rect 5359 -2 5389 16
rect 5432 2 5445 16
rect 5482 3 5490 16
rect 5523 3 5661 16
rect 5694 3 5702 16
rect 5559 2 5610 3
rect 5767 2 5780 16
rect 5560 0 5624 2
rect 5795 -2 5825 16
rect 5868 2 5881 16
use 10T_8x8_magic  10T_8x8_magic_0
timestamp 1666997038
transform 1 0 -2 0 1 1082
box -7 -1098 4631 1122
use 10T_8x8_magic  10T_8x8_magic_1
timestamp 1666997038
transform 1 0 4736 0 1 1082
box -7 -1098 4631 1122
<< end >>
