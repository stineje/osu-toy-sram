magic
tech sky130A
magscale 1 2
timestamp 1668975772
<< error_s >>
rect -478 1828 -465 1844
rect -410 1828 -395 1842
rect -376 1830 -363 1892
rect -295 1840 -142 1886
rect -313 1828 -121 1840
rect -42 1828 -29 1892
rect 53 1828 72 1844
rect 87 1828 93 1844
rect 102 1828 115 1844
rect 170 1828 185 1842
rect 204 1830 217 1892
rect 285 1840 438 1886
rect 267 1828 459 1840
rect 538 1828 551 1892
rect 633 1828 652 1844
rect 667 1828 673 1844
rect 682 1828 695 1844
rect 750 1828 765 1842
rect 784 1830 797 1892
rect 865 1840 1018 1886
rect 847 1828 1039 1840
rect 1118 1828 1131 1892
rect 1213 1828 1232 1844
rect 1247 1828 1253 1844
rect 1262 1828 1275 1844
rect 1330 1828 1345 1842
rect 1364 1830 1377 1892
rect 1445 1840 1598 1886
rect 1427 1828 1619 1840
rect 1698 1828 1711 1892
rect 1793 1828 1812 1844
rect 1827 1828 1833 1844
rect 1842 1828 1855 1844
rect 1910 1828 1925 1842
rect 1944 1830 1957 1892
rect 2025 1840 2178 1886
rect 2007 1828 2199 1840
rect 2278 1828 2291 1892
rect 2373 1828 2392 1844
rect 2407 1828 2413 1844
rect 2422 1828 2435 1844
rect 2490 1828 2505 1842
rect 2524 1830 2537 1892
rect 2605 1840 2758 1886
rect 2587 1828 2779 1840
rect 2858 1828 2871 1892
rect 2953 1828 2972 1844
rect 2987 1828 2993 1844
rect 3002 1828 3015 1844
rect 3070 1828 3085 1842
rect 3104 1830 3117 1892
rect 3185 1840 3338 1886
rect 3167 1828 3359 1840
rect 3438 1828 3451 1892
rect 3533 1828 3552 1844
rect 3567 1828 3573 1844
rect 3582 1828 3595 1844
rect 3650 1828 3665 1842
rect 3684 1830 3697 1892
rect 3765 1840 3918 1886
rect 3747 1828 3939 1840
rect 4018 1828 4031 1892
rect 4113 1828 4132 1844
rect 4147 1828 4153 1844
rect 4162 1828 4175 1844
rect 4230 1828 4245 1842
rect 4264 1830 4277 1892
rect 4345 1840 4498 1886
rect 4327 1828 4519 1840
rect 4598 1828 4611 1892
rect 4693 1828 4712 1844
rect 4727 1828 4733 1844
rect 4742 1828 4755 1844
rect 4810 1828 4825 1842
rect 4844 1830 4857 1892
rect 4925 1840 5078 1886
rect 4907 1828 5099 1840
rect 5178 1828 5191 1892
rect 5273 1828 5292 1844
rect 5307 1828 5313 1844
rect 5322 1828 5335 1844
rect 5390 1828 5405 1842
rect 5424 1830 5437 1892
rect 5505 1840 5658 1886
rect 5487 1828 5679 1840
rect 5758 1828 5771 1892
rect 5853 1828 5872 1844
rect 5887 1828 5893 1844
rect 5902 1828 5915 1844
rect 5970 1828 5985 1842
rect 6004 1830 6017 1892
rect 6085 1840 6238 1886
rect 6067 1828 6259 1840
rect 6338 1828 6351 1892
rect 6439 1828 6452 1844
rect -541 1814 6452 1828
rect -478 1744 -465 1814
rect -420 1798 -403 1802
rect -399 1800 -391 1802
rect -401 1798 -391 1800
rect -420 1788 -391 1798
rect -338 1788 -322 1802
rect -284 1798 -278 1800
rect -271 1798 -163 1814
rect -156 1798 -150 1800
rect -142 1798 -127 1814
rect -61 1808 -42 1811
rect -420 1786 -322 1788
rect -295 1786 -127 1798
rect -112 1788 -96 1802
rect -61 1789 -39 1808
rect -29 1802 -13 1803
rect -30 1800 -13 1802
rect -29 1795 -13 1800
rect -39 1788 -33 1789
rect -30 1788 -1 1795
rect -112 1787 -1 1788
rect -112 1786 5 1787
rect -436 1778 -385 1786
rect -338 1778 -304 1786
rect -436 1766 -411 1778
rect -404 1766 -385 1778
rect -331 1776 -304 1778
rect -295 1776 -74 1786
rect -39 1783 -33 1786
rect -331 1772 -74 1776
rect -436 1758 -385 1766
rect -338 1758 -74 1772
rect -30 1778 5 1786
rect -484 1710 -465 1744
rect -420 1750 -391 1758
rect -420 1744 -403 1750
rect -420 1742 -386 1744
rect -338 1742 -322 1758
rect -321 1748 -113 1758
rect -112 1748 -96 1758
rect -48 1754 -33 1769
rect -30 1766 -29 1778
rect -22 1766 5 1778
rect -30 1758 5 1766
rect -30 1757 -1 1758
rect -310 1744 -96 1748
rect -295 1742 -96 1744
rect -61 1744 -48 1754
rect -30 1744 -13 1757
rect -61 1742 -13 1744
rect -419 1738 -386 1742
rect -423 1736 -386 1738
rect -423 1735 -356 1736
rect -423 1730 -392 1735
rect -386 1730 -356 1735
rect -423 1726 -356 1730
rect -450 1723 -356 1726
rect -450 1716 -401 1723
rect -450 1710 -420 1716
rect -401 1711 -396 1716
rect -484 1694 -404 1710
rect -392 1702 -356 1723
rect -295 1718 -106 1742
rect -61 1741 -14 1742
rect -48 1736 -14 1741
rect -280 1715 -106 1718
rect -287 1712 -106 1715
rect -78 1735 -14 1736
rect -484 1692 -465 1694
rect -450 1692 -416 1694
rect -484 1676 -404 1692
rect -484 1670 -465 1676
rect -494 1654 -465 1670
rect -450 1660 -420 1676
rect -392 1654 -386 1702
rect -383 1696 -364 1702
rect -349 1696 -319 1704
rect -383 1688 -319 1696
rect -383 1672 -303 1688
rect -287 1681 -225 1712
rect -209 1681 -147 1712
rect -78 1710 -29 1735
rect -14 1710 16 1728
rect -115 1696 -85 1704
rect -78 1702 32 1710
rect -115 1688 -70 1696
rect -383 1670 -364 1672
rect -349 1670 -303 1672
rect -383 1654 -303 1670
rect -276 1668 -241 1681
rect -200 1678 -163 1681
rect -200 1676 -158 1678
rect -271 1665 -241 1668
rect -262 1661 -255 1665
rect -255 1660 -254 1661
rect -296 1654 -286 1660
rect -500 1646 -459 1654
rect -500 1620 -485 1646
rect -478 1620 -459 1646
rect -395 1642 -364 1654
rect -349 1642 -246 1654
rect -234 1644 -208 1670
rect -193 1665 -163 1676
rect -131 1672 -69 1688
rect -131 1670 -85 1672
rect -131 1654 -69 1670
rect -57 1654 -51 1702
rect -48 1694 32 1702
rect -48 1692 -29 1694
rect -14 1692 20 1694
rect -48 1677 32 1692
rect -48 1676 38 1677
rect -48 1654 -29 1676
rect -14 1660 16 1676
rect 44 1670 50 1744
rect 53 1670 72 1814
rect 87 1670 93 1814
rect 102 1744 115 1814
rect 160 1798 177 1802
rect 181 1800 189 1802
rect 179 1798 189 1800
rect 160 1788 189 1798
rect 242 1788 258 1802
rect 296 1798 302 1800
rect 309 1798 417 1814
rect 424 1798 430 1800
rect 438 1798 453 1814
rect 519 1808 538 1811
rect 160 1786 258 1788
rect 285 1786 453 1798
rect 468 1788 484 1802
rect 519 1789 541 1808
rect 551 1802 567 1803
rect 550 1800 567 1802
rect 551 1795 567 1800
rect 541 1788 547 1789
rect 550 1788 579 1795
rect 468 1787 579 1788
rect 468 1786 585 1787
rect 144 1778 195 1786
rect 242 1778 276 1786
rect 144 1766 169 1778
rect 176 1766 195 1778
rect 249 1776 276 1778
rect 285 1776 506 1786
rect 541 1783 547 1786
rect 249 1772 506 1776
rect 144 1758 195 1766
rect 242 1758 506 1772
rect 550 1778 585 1786
rect 96 1710 115 1744
rect 160 1750 189 1758
rect 160 1744 177 1750
rect 160 1742 194 1744
rect 242 1742 258 1758
rect 259 1748 467 1758
rect 468 1748 484 1758
rect 532 1754 547 1769
rect 550 1766 551 1778
rect 558 1766 585 1778
rect 550 1758 585 1766
rect 550 1757 579 1758
rect 270 1744 484 1748
rect 285 1742 484 1744
rect 519 1744 532 1754
rect 550 1744 567 1757
rect 519 1742 567 1744
rect 161 1738 194 1742
rect 157 1736 194 1738
rect 157 1735 224 1736
rect 157 1730 188 1735
rect 194 1730 224 1735
rect 157 1726 224 1730
rect 130 1723 224 1726
rect 130 1716 179 1723
rect 130 1710 160 1716
rect 179 1711 184 1716
rect 96 1694 176 1710
rect 188 1702 224 1723
rect 285 1718 474 1742
rect 519 1741 566 1742
rect 532 1736 566 1741
rect 606 1736 622 1738
rect 300 1715 474 1718
rect 293 1712 474 1715
rect 502 1735 566 1736
rect 96 1692 115 1694
rect 130 1692 164 1694
rect 96 1676 176 1692
rect 96 1670 115 1676
rect -188 1644 -85 1654
rect -234 1642 -85 1644
rect -64 1642 -29 1654
rect -395 1640 -233 1642
rect -383 1620 -364 1640
rect -349 1638 -319 1640
rect -500 1612 -459 1620
rect -377 1616 -364 1620
rect -312 1624 -233 1640
rect -201 1640 -29 1642
rect -201 1624 -122 1640
rect -115 1638 -85 1640
rect -494 1602 -465 1612
rect -450 1602 -420 1616
rect -377 1602 -334 1616
rect -312 1612 -122 1624
rect -57 1620 -51 1640
rect -327 1602 -297 1612
rect -296 1602 -138 1612
rect -134 1602 -104 1612
rect -100 1602 -70 1616
rect -42 1602 -29 1640
rect 43 1654 72 1670
rect 86 1654 115 1670
rect 130 1660 160 1676
rect 188 1654 194 1702
rect 197 1696 216 1702
rect 231 1696 261 1704
rect 197 1688 261 1696
rect 197 1672 277 1688
rect 293 1681 355 1712
rect 371 1681 433 1712
rect 502 1710 551 1735
rect 596 1726 622 1736
rect 566 1710 622 1726
rect 465 1696 495 1704
rect 502 1702 612 1710
rect 465 1688 510 1696
rect 197 1670 216 1672
rect 231 1670 277 1672
rect 197 1654 277 1670
rect 304 1668 339 1681
rect 380 1678 417 1681
rect 380 1676 422 1678
rect 309 1665 339 1668
rect 318 1661 325 1665
rect 325 1660 326 1661
rect 284 1654 294 1660
rect 43 1646 78 1654
rect 43 1620 44 1646
rect 51 1620 78 1646
rect -14 1602 16 1616
rect 43 1612 78 1620
rect 80 1646 121 1654
rect 80 1620 95 1646
rect 102 1620 121 1646
rect 185 1642 216 1654
rect 231 1642 334 1654
rect 346 1644 372 1670
rect 387 1665 417 1676
rect 449 1672 511 1688
rect 449 1670 495 1672
rect 449 1654 511 1670
rect 523 1654 529 1702
rect 532 1694 612 1702
rect 532 1692 551 1694
rect 566 1692 600 1694
rect 532 1676 612 1692
rect 532 1654 551 1676
rect 566 1660 596 1676
rect 624 1670 630 1744
rect 633 1670 652 1814
rect 667 1670 673 1814
rect 682 1744 695 1814
rect 740 1798 757 1802
rect 761 1800 769 1802
rect 759 1798 769 1800
rect 740 1788 769 1798
rect 822 1788 838 1802
rect 876 1798 882 1800
rect 889 1798 997 1814
rect 1004 1798 1010 1800
rect 1018 1798 1033 1814
rect 1099 1808 1118 1811
rect 740 1786 838 1788
rect 865 1786 1033 1798
rect 1048 1788 1064 1802
rect 1099 1789 1121 1808
rect 1131 1802 1147 1803
rect 1130 1800 1147 1802
rect 1131 1795 1147 1800
rect 1121 1788 1127 1789
rect 1130 1788 1159 1795
rect 1048 1787 1159 1788
rect 1048 1786 1165 1787
rect 724 1778 775 1786
rect 822 1778 856 1786
rect 724 1766 749 1778
rect 756 1766 775 1778
rect 829 1776 856 1778
rect 865 1776 1086 1786
rect 1121 1783 1127 1786
rect 829 1772 1086 1776
rect 724 1758 775 1766
rect 822 1758 1086 1772
rect 1130 1778 1165 1786
rect 676 1710 695 1744
rect 740 1750 769 1758
rect 740 1744 757 1750
rect 740 1742 774 1744
rect 822 1742 838 1758
rect 839 1748 1047 1758
rect 1048 1748 1064 1758
rect 1112 1754 1127 1769
rect 1130 1766 1131 1778
rect 1138 1766 1165 1778
rect 1130 1758 1165 1766
rect 1130 1757 1159 1758
rect 850 1744 1064 1748
rect 865 1742 1064 1744
rect 1099 1744 1112 1754
rect 1130 1744 1147 1757
rect 1099 1742 1147 1744
rect 741 1738 774 1742
rect 737 1736 774 1738
rect 737 1735 804 1736
rect 737 1730 768 1735
rect 774 1730 804 1735
rect 737 1726 804 1730
rect 710 1723 804 1726
rect 710 1716 759 1723
rect 710 1710 740 1716
rect 759 1711 764 1716
rect 676 1694 756 1710
rect 768 1702 804 1723
rect 865 1718 1054 1742
rect 1099 1741 1146 1742
rect 1112 1736 1146 1741
rect 880 1715 1054 1718
rect 873 1712 1054 1715
rect 1082 1735 1146 1736
rect 676 1692 695 1694
rect 710 1692 744 1694
rect 676 1676 756 1692
rect 676 1670 695 1676
rect 392 1644 495 1654
rect 346 1642 495 1644
rect 516 1642 551 1654
rect 185 1640 347 1642
rect 197 1620 216 1640
rect 231 1638 261 1640
rect 80 1612 121 1620
rect 203 1616 216 1620
rect 268 1624 347 1640
rect 379 1640 551 1642
rect 379 1624 458 1640
rect 465 1638 495 1640
rect 43 1602 72 1612
rect 86 1602 115 1612
rect 130 1602 160 1616
rect 203 1602 246 1616
rect 268 1612 458 1624
rect 523 1620 529 1640
rect 253 1602 283 1612
rect 284 1602 442 1612
rect 446 1602 476 1612
rect 480 1602 510 1616
rect 538 1602 551 1640
rect 623 1654 652 1670
rect 666 1654 695 1670
rect 710 1660 740 1676
rect 768 1654 774 1702
rect 777 1696 796 1702
rect 811 1696 841 1704
rect 777 1688 841 1696
rect 777 1672 857 1688
rect 873 1681 935 1712
rect 951 1681 1013 1712
rect 1082 1710 1131 1735
rect 1146 1710 1176 1728
rect 1045 1696 1075 1704
rect 1082 1702 1192 1710
rect 1045 1688 1090 1696
rect 777 1670 796 1672
rect 811 1670 857 1672
rect 777 1654 857 1670
rect 884 1668 919 1681
rect 960 1678 997 1681
rect 960 1676 1002 1678
rect 889 1665 919 1668
rect 898 1661 905 1665
rect 905 1660 906 1661
rect 864 1654 874 1660
rect 623 1646 658 1654
rect 623 1620 624 1646
rect 631 1620 658 1646
rect 566 1602 596 1616
rect 623 1612 658 1620
rect 660 1646 701 1654
rect 660 1620 675 1646
rect 682 1620 701 1646
rect 765 1642 796 1654
rect 811 1642 914 1654
rect 926 1644 952 1670
rect 967 1665 997 1676
rect 1029 1672 1091 1688
rect 1029 1670 1075 1672
rect 1029 1654 1091 1670
rect 1103 1654 1109 1702
rect 1112 1694 1192 1702
rect 1112 1692 1131 1694
rect 1146 1692 1180 1694
rect 1112 1677 1192 1692
rect 1112 1676 1198 1677
rect 1112 1654 1131 1676
rect 1146 1660 1176 1676
rect 1204 1670 1210 1744
rect 1213 1670 1232 1814
rect 1247 1670 1253 1814
rect 1262 1744 1275 1814
rect 1320 1798 1337 1802
rect 1341 1800 1349 1802
rect 1339 1798 1349 1800
rect 1320 1788 1349 1798
rect 1402 1788 1418 1802
rect 1456 1798 1462 1800
rect 1469 1798 1577 1814
rect 1584 1798 1590 1800
rect 1598 1798 1613 1814
rect 1679 1808 1698 1811
rect 1320 1786 1418 1788
rect 1445 1786 1613 1798
rect 1628 1788 1644 1802
rect 1679 1789 1701 1808
rect 1711 1802 1727 1803
rect 1710 1800 1727 1802
rect 1711 1795 1727 1800
rect 1701 1788 1707 1789
rect 1710 1788 1739 1795
rect 1628 1787 1739 1788
rect 1628 1786 1745 1787
rect 1304 1778 1355 1786
rect 1402 1778 1436 1786
rect 1304 1766 1329 1778
rect 1336 1766 1355 1778
rect 1409 1776 1436 1778
rect 1445 1776 1666 1786
rect 1701 1783 1707 1786
rect 1409 1772 1666 1776
rect 1304 1758 1355 1766
rect 1402 1758 1666 1772
rect 1710 1778 1745 1786
rect 1256 1710 1275 1744
rect 1320 1750 1349 1758
rect 1320 1744 1337 1750
rect 1320 1742 1354 1744
rect 1402 1742 1418 1758
rect 1419 1748 1627 1758
rect 1628 1748 1644 1758
rect 1692 1754 1707 1769
rect 1710 1766 1711 1778
rect 1718 1766 1745 1778
rect 1710 1758 1745 1766
rect 1710 1757 1739 1758
rect 1430 1744 1644 1748
rect 1445 1742 1644 1744
rect 1679 1744 1692 1754
rect 1710 1744 1727 1757
rect 1679 1742 1727 1744
rect 1321 1738 1354 1742
rect 1317 1736 1354 1738
rect 1317 1735 1384 1736
rect 1317 1730 1348 1735
rect 1354 1730 1384 1735
rect 1317 1726 1384 1730
rect 1290 1723 1384 1726
rect 1290 1716 1339 1723
rect 1290 1710 1320 1716
rect 1339 1711 1344 1716
rect 1256 1694 1336 1710
rect 1348 1702 1384 1723
rect 1445 1718 1634 1742
rect 1679 1741 1726 1742
rect 1692 1736 1726 1741
rect 1766 1736 1782 1738
rect 1460 1715 1634 1718
rect 1453 1712 1634 1715
rect 1662 1735 1726 1736
rect 1256 1692 1275 1694
rect 1290 1692 1324 1694
rect 1256 1676 1336 1692
rect 1256 1670 1275 1676
rect 972 1644 1075 1654
rect 926 1642 1075 1644
rect 1096 1642 1131 1654
rect 765 1640 927 1642
rect 777 1620 796 1640
rect 811 1638 841 1640
rect 660 1612 701 1620
rect 783 1616 796 1620
rect 848 1624 927 1640
rect 959 1640 1131 1642
rect 959 1624 1038 1640
rect 1045 1638 1075 1640
rect 623 1602 652 1612
rect 666 1602 695 1612
rect 710 1602 740 1616
rect 783 1602 826 1616
rect 848 1612 1038 1624
rect 1103 1620 1109 1640
rect 833 1602 863 1612
rect 864 1602 1022 1612
rect 1026 1602 1056 1612
rect 1060 1602 1090 1616
rect 1118 1602 1131 1640
rect 1203 1654 1232 1670
rect 1246 1654 1275 1670
rect 1290 1660 1320 1676
rect 1348 1654 1354 1702
rect 1357 1696 1376 1702
rect 1391 1696 1421 1704
rect 1357 1688 1421 1696
rect 1357 1672 1437 1688
rect 1453 1681 1515 1712
rect 1531 1681 1593 1712
rect 1662 1710 1711 1735
rect 1756 1726 1782 1736
rect 1726 1710 1782 1726
rect 1625 1696 1655 1704
rect 1662 1702 1772 1710
rect 1625 1688 1670 1696
rect 1357 1670 1376 1672
rect 1391 1670 1437 1672
rect 1357 1654 1437 1670
rect 1464 1668 1499 1681
rect 1540 1678 1577 1681
rect 1540 1676 1582 1678
rect 1469 1665 1499 1668
rect 1478 1661 1485 1665
rect 1485 1660 1486 1661
rect 1444 1654 1454 1660
rect 1203 1646 1238 1654
rect 1203 1620 1204 1646
rect 1211 1620 1238 1646
rect 1146 1602 1176 1616
rect 1203 1612 1238 1620
rect 1240 1646 1281 1654
rect 1240 1620 1255 1646
rect 1262 1620 1281 1646
rect 1345 1642 1376 1654
rect 1391 1642 1494 1654
rect 1506 1644 1532 1670
rect 1547 1665 1577 1676
rect 1609 1672 1671 1688
rect 1609 1670 1655 1672
rect 1609 1654 1671 1670
rect 1683 1654 1689 1702
rect 1692 1694 1772 1702
rect 1692 1692 1711 1694
rect 1726 1692 1760 1694
rect 1692 1676 1772 1692
rect 1692 1654 1711 1676
rect 1726 1660 1756 1676
rect 1784 1670 1790 1744
rect 1793 1670 1812 1814
rect 1827 1670 1833 1814
rect 1842 1744 1855 1814
rect 1900 1798 1917 1802
rect 1921 1800 1929 1802
rect 1919 1798 1929 1800
rect 1900 1788 1929 1798
rect 1982 1788 1998 1802
rect 2036 1798 2042 1800
rect 2049 1798 2157 1814
rect 2164 1798 2170 1800
rect 2178 1798 2193 1814
rect 2259 1808 2278 1811
rect 1900 1786 1998 1788
rect 2025 1786 2193 1798
rect 2208 1788 2224 1802
rect 2259 1789 2281 1808
rect 2291 1802 2307 1803
rect 2290 1800 2307 1802
rect 2291 1795 2307 1800
rect 2281 1788 2287 1789
rect 2290 1788 2319 1795
rect 2208 1787 2319 1788
rect 2208 1786 2325 1787
rect 1884 1778 1935 1786
rect 1982 1778 2016 1786
rect 1884 1766 1909 1778
rect 1916 1766 1935 1778
rect 1989 1776 2016 1778
rect 2025 1776 2246 1786
rect 2281 1783 2287 1786
rect 1989 1772 2246 1776
rect 1884 1758 1935 1766
rect 1982 1758 2246 1772
rect 2290 1778 2325 1786
rect 1836 1710 1855 1744
rect 1900 1750 1929 1758
rect 1900 1744 1917 1750
rect 1900 1742 1934 1744
rect 1982 1742 1998 1758
rect 1999 1748 2207 1758
rect 2208 1748 2224 1758
rect 2272 1754 2287 1769
rect 2290 1766 2291 1778
rect 2298 1766 2325 1778
rect 2290 1758 2325 1766
rect 2290 1757 2319 1758
rect 2010 1744 2224 1748
rect 2025 1742 2224 1744
rect 2259 1744 2272 1754
rect 2290 1744 2307 1757
rect 2259 1742 2307 1744
rect 1901 1738 1934 1742
rect 1897 1736 1934 1738
rect 1897 1735 1964 1736
rect 1897 1730 1928 1735
rect 1934 1730 1964 1735
rect 1897 1726 1964 1730
rect 1870 1723 1964 1726
rect 1870 1716 1919 1723
rect 1870 1710 1900 1716
rect 1919 1711 1924 1716
rect 1836 1694 1916 1710
rect 1928 1702 1964 1723
rect 2025 1718 2214 1742
rect 2259 1741 2306 1742
rect 2272 1736 2306 1741
rect 2040 1715 2214 1718
rect 2033 1712 2214 1715
rect 2242 1735 2306 1736
rect 1836 1692 1855 1694
rect 1870 1692 1904 1694
rect 1836 1676 1916 1692
rect 1836 1670 1855 1676
rect 1552 1644 1655 1654
rect 1506 1642 1655 1644
rect 1676 1642 1711 1654
rect 1345 1640 1507 1642
rect 1357 1620 1376 1640
rect 1391 1638 1421 1640
rect 1240 1612 1281 1620
rect 1363 1616 1376 1620
rect 1428 1624 1507 1640
rect 1539 1640 1711 1642
rect 1539 1624 1618 1640
rect 1625 1638 1655 1640
rect 1203 1602 1232 1612
rect 1246 1602 1275 1612
rect 1290 1602 1320 1616
rect 1363 1602 1406 1616
rect 1428 1612 1618 1624
rect 1683 1620 1689 1640
rect 1413 1602 1443 1612
rect 1444 1602 1602 1612
rect 1606 1602 1636 1612
rect 1640 1602 1670 1616
rect 1698 1602 1711 1640
rect 1783 1654 1812 1670
rect 1826 1654 1855 1670
rect 1870 1660 1900 1676
rect 1928 1654 1934 1702
rect 1937 1696 1956 1702
rect 1971 1696 2001 1704
rect 1937 1688 2001 1696
rect 1937 1672 2017 1688
rect 2033 1681 2095 1712
rect 2111 1681 2173 1712
rect 2242 1710 2291 1735
rect 2306 1710 2336 1728
rect 2205 1696 2235 1704
rect 2242 1702 2352 1710
rect 2205 1688 2250 1696
rect 1937 1670 1956 1672
rect 1971 1670 2017 1672
rect 1937 1654 2017 1670
rect 2044 1668 2079 1681
rect 2120 1678 2157 1681
rect 2120 1676 2162 1678
rect 2049 1665 2079 1668
rect 2058 1661 2065 1665
rect 2065 1660 2066 1661
rect 2024 1654 2034 1660
rect 1783 1646 1818 1654
rect 1783 1620 1784 1646
rect 1791 1620 1818 1646
rect 1726 1602 1756 1616
rect 1783 1612 1818 1620
rect 1820 1646 1861 1654
rect 1820 1620 1835 1646
rect 1842 1620 1861 1646
rect 1925 1642 1956 1654
rect 1971 1642 2074 1654
rect 2086 1644 2112 1670
rect 2127 1665 2157 1676
rect 2189 1672 2251 1688
rect 2189 1670 2235 1672
rect 2189 1654 2251 1670
rect 2263 1654 2269 1702
rect 2272 1694 2352 1702
rect 2272 1692 2291 1694
rect 2306 1692 2340 1694
rect 2272 1677 2352 1692
rect 2272 1676 2358 1677
rect 2272 1654 2291 1676
rect 2306 1660 2336 1676
rect 2364 1670 2370 1744
rect 2373 1670 2392 1814
rect 2407 1670 2413 1814
rect 2422 1744 2435 1814
rect 2480 1798 2497 1802
rect 2501 1800 2509 1802
rect 2499 1798 2509 1800
rect 2480 1788 2509 1798
rect 2562 1788 2578 1802
rect 2616 1798 2622 1800
rect 2629 1798 2737 1814
rect 2744 1798 2750 1800
rect 2758 1798 2773 1814
rect 2839 1808 2858 1811
rect 2480 1786 2578 1788
rect 2605 1786 2773 1798
rect 2788 1788 2804 1802
rect 2839 1789 2861 1808
rect 2871 1802 2887 1803
rect 2870 1800 2887 1802
rect 2871 1795 2887 1800
rect 2861 1788 2867 1789
rect 2870 1788 2899 1795
rect 2788 1787 2899 1788
rect 2788 1786 2905 1787
rect 2464 1778 2515 1786
rect 2562 1778 2596 1786
rect 2464 1766 2489 1778
rect 2496 1766 2515 1778
rect 2569 1776 2596 1778
rect 2605 1776 2826 1786
rect 2861 1783 2867 1786
rect 2569 1772 2826 1776
rect 2464 1758 2515 1766
rect 2562 1758 2826 1772
rect 2870 1778 2905 1786
rect 2416 1710 2435 1744
rect 2480 1750 2509 1758
rect 2480 1744 2497 1750
rect 2480 1742 2514 1744
rect 2562 1742 2578 1758
rect 2579 1748 2787 1758
rect 2788 1748 2804 1758
rect 2852 1754 2867 1769
rect 2870 1766 2871 1778
rect 2878 1766 2905 1778
rect 2870 1758 2905 1766
rect 2870 1757 2899 1758
rect 2590 1744 2804 1748
rect 2605 1742 2804 1744
rect 2839 1744 2852 1754
rect 2870 1744 2887 1757
rect 2839 1742 2887 1744
rect 2481 1738 2514 1742
rect 2477 1736 2514 1738
rect 2477 1735 2544 1736
rect 2477 1730 2508 1735
rect 2514 1730 2544 1735
rect 2477 1726 2544 1730
rect 2450 1723 2544 1726
rect 2450 1716 2499 1723
rect 2450 1710 2480 1716
rect 2499 1711 2504 1716
rect 2416 1694 2496 1710
rect 2508 1702 2544 1723
rect 2605 1718 2794 1742
rect 2839 1741 2886 1742
rect 2852 1736 2886 1741
rect 2926 1736 2942 1738
rect 2620 1715 2794 1718
rect 2613 1712 2794 1715
rect 2822 1735 2886 1736
rect 2416 1692 2435 1694
rect 2450 1692 2484 1694
rect 2416 1676 2496 1692
rect 2416 1670 2435 1676
rect 2132 1644 2235 1654
rect 2086 1642 2235 1644
rect 2256 1642 2291 1654
rect 1925 1640 2087 1642
rect 1937 1620 1956 1640
rect 1971 1638 2001 1640
rect 1820 1612 1861 1620
rect 1943 1616 1956 1620
rect 2008 1624 2087 1640
rect 2119 1640 2291 1642
rect 2119 1624 2198 1640
rect 2205 1638 2235 1640
rect 1783 1602 1812 1612
rect 1826 1602 1855 1612
rect 1870 1602 1900 1616
rect 1943 1602 1986 1616
rect 2008 1612 2198 1624
rect 2263 1620 2269 1640
rect 1993 1602 2023 1612
rect 2024 1602 2182 1612
rect 2186 1602 2216 1612
rect 2220 1602 2250 1616
rect 2278 1602 2291 1640
rect 2363 1654 2392 1670
rect 2406 1654 2435 1670
rect 2450 1660 2480 1676
rect 2508 1654 2514 1702
rect 2517 1696 2536 1702
rect 2551 1696 2581 1704
rect 2517 1688 2581 1696
rect 2517 1672 2597 1688
rect 2613 1681 2675 1712
rect 2691 1681 2753 1712
rect 2822 1710 2871 1735
rect 2916 1726 2942 1736
rect 2886 1710 2942 1726
rect 2785 1696 2815 1704
rect 2822 1702 2932 1710
rect 2785 1688 2830 1696
rect 2517 1670 2536 1672
rect 2551 1670 2597 1672
rect 2517 1654 2597 1670
rect 2624 1668 2659 1681
rect 2700 1678 2737 1681
rect 2700 1676 2742 1678
rect 2629 1665 2659 1668
rect 2638 1661 2645 1665
rect 2645 1660 2646 1661
rect 2604 1654 2614 1660
rect 2363 1646 2398 1654
rect 2363 1620 2364 1646
rect 2371 1620 2398 1646
rect 2306 1602 2336 1616
rect 2363 1612 2398 1620
rect 2400 1646 2441 1654
rect 2400 1620 2415 1646
rect 2422 1620 2441 1646
rect 2505 1642 2536 1654
rect 2551 1642 2654 1654
rect 2666 1644 2692 1670
rect 2707 1665 2737 1676
rect 2769 1672 2831 1688
rect 2769 1670 2815 1672
rect 2769 1654 2831 1670
rect 2843 1654 2849 1702
rect 2852 1694 2932 1702
rect 2852 1692 2871 1694
rect 2886 1692 2920 1694
rect 2852 1676 2932 1692
rect 2852 1654 2871 1676
rect 2886 1660 2916 1676
rect 2944 1670 2950 1744
rect 2953 1670 2972 1814
rect 2987 1670 2993 1814
rect 3002 1744 3015 1814
rect 3060 1798 3077 1802
rect 3081 1800 3089 1802
rect 3079 1798 3089 1800
rect 3060 1788 3089 1798
rect 3142 1788 3158 1802
rect 3196 1798 3202 1800
rect 3209 1798 3317 1814
rect 3324 1798 3330 1800
rect 3338 1798 3353 1814
rect 3419 1808 3438 1811
rect 3060 1786 3158 1788
rect 3185 1786 3353 1798
rect 3368 1788 3384 1802
rect 3419 1789 3441 1808
rect 3451 1802 3467 1803
rect 3450 1800 3467 1802
rect 3451 1795 3467 1800
rect 3441 1788 3447 1789
rect 3450 1788 3479 1795
rect 3368 1787 3479 1788
rect 3368 1786 3485 1787
rect 3044 1778 3095 1786
rect 3142 1778 3176 1786
rect 3044 1766 3069 1778
rect 3076 1766 3095 1778
rect 3149 1776 3176 1778
rect 3185 1776 3406 1786
rect 3441 1783 3447 1786
rect 3149 1772 3406 1776
rect 3044 1758 3095 1766
rect 3142 1758 3406 1772
rect 3450 1778 3485 1786
rect 2996 1710 3015 1744
rect 3060 1750 3089 1758
rect 3060 1744 3077 1750
rect 3060 1742 3094 1744
rect 3142 1742 3158 1758
rect 3159 1748 3367 1758
rect 3368 1748 3384 1758
rect 3432 1754 3447 1769
rect 3450 1766 3451 1778
rect 3458 1766 3485 1778
rect 3450 1758 3485 1766
rect 3450 1757 3479 1758
rect 3170 1744 3384 1748
rect 3185 1742 3384 1744
rect 3419 1744 3432 1754
rect 3450 1744 3467 1757
rect 3419 1742 3467 1744
rect 3061 1738 3094 1742
rect 3057 1736 3094 1738
rect 3057 1735 3124 1736
rect 3057 1730 3088 1735
rect 3094 1730 3124 1735
rect 3057 1726 3124 1730
rect 3030 1723 3124 1726
rect 3030 1716 3079 1723
rect 3030 1710 3060 1716
rect 3079 1711 3084 1716
rect 2996 1694 3076 1710
rect 3088 1702 3124 1723
rect 3185 1718 3374 1742
rect 3419 1741 3466 1742
rect 3432 1736 3466 1741
rect 3200 1715 3374 1718
rect 3193 1712 3374 1715
rect 3402 1735 3466 1736
rect 2996 1692 3015 1694
rect 3030 1692 3064 1694
rect 2996 1676 3076 1692
rect 2996 1670 3015 1676
rect 2712 1644 2815 1654
rect 2666 1642 2815 1644
rect 2836 1642 2871 1654
rect 2505 1640 2667 1642
rect 2517 1620 2536 1640
rect 2551 1638 2581 1640
rect 2400 1612 2441 1620
rect 2523 1616 2536 1620
rect 2588 1624 2667 1640
rect 2699 1640 2871 1642
rect 2699 1624 2778 1640
rect 2785 1638 2815 1640
rect 2363 1602 2392 1612
rect 2406 1602 2435 1612
rect 2450 1602 2480 1616
rect 2523 1602 2566 1616
rect 2588 1612 2778 1624
rect 2843 1620 2849 1640
rect 2573 1602 2603 1612
rect 2604 1602 2762 1612
rect 2766 1602 2796 1612
rect 2800 1602 2830 1616
rect 2858 1602 2871 1640
rect 2943 1654 2972 1670
rect 2986 1654 3015 1670
rect 3030 1660 3060 1676
rect 3088 1654 3094 1702
rect 3097 1696 3116 1702
rect 3131 1696 3161 1704
rect 3097 1688 3161 1696
rect 3097 1672 3177 1688
rect 3193 1681 3255 1712
rect 3271 1681 3333 1712
rect 3402 1710 3451 1735
rect 3466 1710 3496 1728
rect 3365 1696 3395 1704
rect 3402 1702 3512 1710
rect 3365 1688 3410 1696
rect 3097 1670 3116 1672
rect 3131 1670 3177 1672
rect 3097 1654 3177 1670
rect 3204 1668 3239 1681
rect 3280 1678 3317 1681
rect 3280 1676 3322 1678
rect 3209 1665 3239 1668
rect 3218 1661 3225 1665
rect 3225 1660 3226 1661
rect 3184 1654 3194 1660
rect 2943 1646 2978 1654
rect 2943 1620 2944 1646
rect 2951 1620 2978 1646
rect 2886 1602 2916 1616
rect 2943 1612 2978 1620
rect 2980 1646 3021 1654
rect 2980 1620 2995 1646
rect 3002 1620 3021 1646
rect 3085 1642 3116 1654
rect 3131 1642 3234 1654
rect 3246 1644 3272 1670
rect 3287 1665 3317 1676
rect 3349 1672 3411 1688
rect 3349 1670 3395 1672
rect 3349 1654 3411 1670
rect 3423 1654 3429 1702
rect 3432 1694 3512 1702
rect 3432 1692 3451 1694
rect 3466 1692 3500 1694
rect 3432 1677 3512 1692
rect 3432 1676 3518 1677
rect 3432 1654 3451 1676
rect 3466 1660 3496 1676
rect 3524 1670 3530 1744
rect 3533 1670 3552 1814
rect 3567 1670 3573 1814
rect 3582 1744 3595 1814
rect 3640 1798 3657 1802
rect 3661 1800 3669 1802
rect 3659 1798 3669 1800
rect 3640 1788 3669 1798
rect 3722 1788 3738 1802
rect 3776 1798 3782 1800
rect 3789 1798 3897 1814
rect 3904 1798 3910 1800
rect 3918 1798 3933 1814
rect 3999 1808 4018 1811
rect 3640 1786 3738 1788
rect 3765 1786 3933 1798
rect 3948 1788 3964 1802
rect 3999 1789 4021 1808
rect 4031 1802 4047 1803
rect 4030 1800 4047 1802
rect 4031 1795 4047 1800
rect 4021 1788 4027 1789
rect 4030 1788 4059 1795
rect 3948 1787 4059 1788
rect 3948 1786 4065 1787
rect 3624 1778 3675 1786
rect 3722 1778 3756 1786
rect 3624 1766 3649 1778
rect 3656 1766 3675 1778
rect 3729 1776 3756 1778
rect 3765 1776 3986 1786
rect 4021 1783 4027 1786
rect 3729 1772 3986 1776
rect 3624 1758 3675 1766
rect 3722 1758 3986 1772
rect 4030 1778 4065 1786
rect 3576 1710 3595 1744
rect 3640 1750 3669 1758
rect 3640 1744 3657 1750
rect 3640 1742 3674 1744
rect 3722 1742 3738 1758
rect 3739 1748 3947 1758
rect 3948 1748 3964 1758
rect 4012 1754 4027 1769
rect 4030 1766 4031 1778
rect 4038 1766 4065 1778
rect 4030 1758 4065 1766
rect 4030 1757 4059 1758
rect 3750 1744 3964 1748
rect 3765 1742 3964 1744
rect 3999 1744 4012 1754
rect 4030 1744 4047 1757
rect 3999 1742 4047 1744
rect 3641 1738 3674 1742
rect 3637 1736 3674 1738
rect 3637 1735 3704 1736
rect 3637 1730 3668 1735
rect 3674 1730 3704 1735
rect 3637 1726 3704 1730
rect 3610 1723 3704 1726
rect 3610 1716 3659 1723
rect 3610 1710 3640 1716
rect 3659 1711 3664 1716
rect 3576 1694 3656 1710
rect 3668 1702 3704 1723
rect 3765 1718 3954 1742
rect 3999 1741 4046 1742
rect 4012 1736 4046 1741
rect 4086 1736 4102 1738
rect 3780 1715 3954 1718
rect 3773 1712 3954 1715
rect 3982 1735 4046 1736
rect 3576 1692 3595 1694
rect 3610 1692 3644 1694
rect 3576 1676 3656 1692
rect 3576 1670 3595 1676
rect 3292 1644 3395 1654
rect 3246 1642 3395 1644
rect 3416 1642 3451 1654
rect 3085 1640 3247 1642
rect 3097 1620 3116 1640
rect 3131 1638 3161 1640
rect 2980 1612 3021 1620
rect 3103 1616 3116 1620
rect 3168 1624 3247 1640
rect 3279 1640 3451 1642
rect 3279 1624 3358 1640
rect 3365 1638 3395 1640
rect 2943 1602 2972 1612
rect 2986 1602 3015 1612
rect 3030 1602 3060 1616
rect 3103 1602 3146 1616
rect 3168 1612 3358 1624
rect 3423 1620 3429 1640
rect 3153 1602 3183 1612
rect 3184 1602 3342 1612
rect 3346 1602 3376 1612
rect 3380 1602 3410 1616
rect 3438 1602 3451 1640
rect 3523 1654 3552 1670
rect 3566 1654 3595 1670
rect 3610 1660 3640 1676
rect 3668 1654 3674 1702
rect 3677 1696 3696 1702
rect 3711 1696 3741 1704
rect 3677 1688 3741 1696
rect 3677 1672 3757 1688
rect 3773 1681 3835 1712
rect 3851 1681 3913 1712
rect 3982 1710 4031 1735
rect 4076 1726 4102 1736
rect 4046 1710 4102 1726
rect 3945 1696 3975 1704
rect 3982 1702 4092 1710
rect 3945 1688 3990 1696
rect 3677 1670 3696 1672
rect 3711 1670 3757 1672
rect 3677 1654 3757 1670
rect 3784 1668 3819 1681
rect 3860 1678 3897 1681
rect 3860 1676 3902 1678
rect 3789 1665 3819 1668
rect 3798 1661 3805 1665
rect 3805 1660 3806 1661
rect 3764 1654 3774 1660
rect 3523 1646 3558 1654
rect 3523 1620 3524 1646
rect 3531 1620 3558 1646
rect 3466 1602 3496 1616
rect 3523 1612 3558 1620
rect 3560 1646 3601 1654
rect 3560 1620 3575 1646
rect 3582 1620 3601 1646
rect 3665 1642 3696 1654
rect 3711 1642 3814 1654
rect 3826 1644 3852 1670
rect 3867 1665 3897 1676
rect 3929 1672 3991 1688
rect 3929 1670 3975 1672
rect 3929 1654 3991 1670
rect 4003 1654 4009 1702
rect 4012 1694 4092 1702
rect 4012 1692 4031 1694
rect 4046 1692 4080 1694
rect 4012 1676 4092 1692
rect 4012 1654 4031 1676
rect 4046 1660 4076 1676
rect 4104 1670 4110 1744
rect 4113 1670 4132 1814
rect 4147 1670 4153 1814
rect 4162 1744 4175 1814
rect 4220 1798 4237 1802
rect 4241 1800 4249 1802
rect 4239 1798 4249 1800
rect 4220 1788 4249 1798
rect 4302 1788 4318 1802
rect 4356 1798 4362 1800
rect 4369 1798 4477 1814
rect 4484 1798 4490 1800
rect 4498 1798 4513 1814
rect 4579 1808 4598 1811
rect 4220 1786 4318 1788
rect 4345 1786 4513 1798
rect 4528 1788 4544 1802
rect 4579 1789 4601 1808
rect 4611 1802 4627 1803
rect 4610 1800 4627 1802
rect 4611 1795 4627 1800
rect 4601 1788 4607 1789
rect 4610 1788 4639 1795
rect 4528 1787 4639 1788
rect 4528 1786 4645 1787
rect 4204 1778 4255 1786
rect 4302 1778 4336 1786
rect 4204 1766 4229 1778
rect 4236 1766 4255 1778
rect 4309 1776 4336 1778
rect 4345 1776 4566 1786
rect 4601 1783 4607 1786
rect 4309 1772 4566 1776
rect 4204 1758 4255 1766
rect 4302 1758 4566 1772
rect 4610 1778 4645 1786
rect 4156 1710 4175 1744
rect 4220 1750 4249 1758
rect 4220 1744 4237 1750
rect 4220 1742 4254 1744
rect 4302 1742 4318 1758
rect 4319 1748 4527 1758
rect 4528 1748 4544 1758
rect 4592 1754 4607 1769
rect 4610 1766 4611 1778
rect 4618 1766 4645 1778
rect 4610 1758 4645 1766
rect 4610 1757 4639 1758
rect 4330 1744 4544 1748
rect 4345 1742 4544 1744
rect 4579 1744 4592 1754
rect 4610 1744 4627 1757
rect 4579 1742 4627 1744
rect 4221 1738 4254 1742
rect 4217 1736 4254 1738
rect 4217 1735 4284 1736
rect 4217 1730 4248 1735
rect 4254 1730 4284 1735
rect 4217 1726 4284 1730
rect 4190 1723 4284 1726
rect 4190 1716 4239 1723
rect 4190 1710 4220 1716
rect 4239 1711 4244 1716
rect 4156 1694 4236 1710
rect 4248 1702 4284 1723
rect 4345 1718 4534 1742
rect 4579 1741 4626 1742
rect 4592 1736 4626 1741
rect 4360 1715 4534 1718
rect 4353 1712 4534 1715
rect 4562 1735 4626 1736
rect 4156 1692 4175 1694
rect 4190 1692 4224 1694
rect 4156 1676 4236 1692
rect 4156 1670 4175 1676
rect 3872 1644 3975 1654
rect 3826 1642 3975 1644
rect 3996 1642 4031 1654
rect 3665 1640 3827 1642
rect 3677 1620 3696 1640
rect 3711 1638 3741 1640
rect 3560 1612 3601 1620
rect 3683 1616 3696 1620
rect 3748 1624 3827 1640
rect 3859 1640 4031 1642
rect 3859 1624 3938 1640
rect 3945 1638 3975 1640
rect 3523 1602 3552 1612
rect 3566 1602 3595 1612
rect 3610 1602 3640 1616
rect 3683 1602 3726 1616
rect 3748 1612 3938 1624
rect 4003 1620 4009 1640
rect 3733 1602 3763 1612
rect 3764 1602 3922 1612
rect 3926 1602 3956 1612
rect 3960 1602 3990 1616
rect 4018 1602 4031 1640
rect 4103 1654 4132 1670
rect 4146 1654 4175 1670
rect 4190 1660 4220 1676
rect 4248 1654 4254 1702
rect 4257 1696 4276 1702
rect 4291 1696 4321 1704
rect 4257 1688 4321 1696
rect 4257 1672 4337 1688
rect 4353 1681 4415 1712
rect 4431 1681 4493 1712
rect 4562 1710 4611 1735
rect 4626 1710 4656 1728
rect 4525 1696 4555 1704
rect 4562 1702 4672 1710
rect 4525 1688 4570 1696
rect 4257 1670 4276 1672
rect 4291 1670 4337 1672
rect 4257 1654 4337 1670
rect 4364 1668 4399 1681
rect 4440 1678 4477 1681
rect 4440 1676 4482 1678
rect 4369 1665 4399 1668
rect 4378 1661 4385 1665
rect 4385 1660 4386 1661
rect 4344 1654 4354 1660
rect 4103 1646 4138 1654
rect 4103 1620 4104 1646
rect 4111 1620 4138 1646
rect 4046 1602 4076 1616
rect 4103 1612 4138 1620
rect 4140 1646 4181 1654
rect 4140 1620 4155 1646
rect 4162 1620 4181 1646
rect 4245 1642 4276 1654
rect 4291 1642 4394 1654
rect 4406 1644 4432 1670
rect 4447 1665 4477 1676
rect 4509 1672 4571 1688
rect 4509 1670 4555 1672
rect 4509 1654 4571 1670
rect 4583 1654 4589 1702
rect 4592 1694 4672 1702
rect 4592 1692 4611 1694
rect 4626 1692 4660 1694
rect 4592 1677 4672 1692
rect 4592 1676 4678 1677
rect 4592 1654 4611 1676
rect 4626 1660 4656 1676
rect 4684 1670 4690 1744
rect 4693 1670 4712 1814
rect 4727 1670 4733 1814
rect 4742 1744 4755 1814
rect 4800 1798 4817 1802
rect 4821 1800 4829 1802
rect 4819 1798 4829 1800
rect 4800 1788 4829 1798
rect 4882 1788 4898 1802
rect 4936 1798 4942 1800
rect 4949 1798 5057 1814
rect 5064 1798 5070 1800
rect 5078 1798 5093 1814
rect 5159 1808 5178 1811
rect 4800 1786 4898 1788
rect 4925 1786 5093 1798
rect 5108 1788 5124 1802
rect 5159 1789 5181 1808
rect 5191 1802 5207 1803
rect 5190 1800 5207 1802
rect 5191 1795 5207 1800
rect 5181 1788 5187 1789
rect 5190 1788 5219 1795
rect 5108 1787 5219 1788
rect 5108 1786 5225 1787
rect 4784 1778 4835 1786
rect 4882 1778 4916 1786
rect 4784 1766 4809 1778
rect 4816 1766 4835 1778
rect 4889 1776 4916 1778
rect 4925 1776 5146 1786
rect 5181 1783 5187 1786
rect 4889 1772 5146 1776
rect 4784 1758 4835 1766
rect 4882 1758 5146 1772
rect 5190 1778 5225 1786
rect 4736 1710 4755 1744
rect 4800 1750 4829 1758
rect 4800 1744 4817 1750
rect 4800 1742 4834 1744
rect 4882 1742 4898 1758
rect 4899 1748 5107 1758
rect 5108 1748 5124 1758
rect 5172 1754 5187 1769
rect 5190 1766 5191 1778
rect 5198 1766 5225 1778
rect 5190 1758 5225 1766
rect 5190 1757 5219 1758
rect 4910 1744 5124 1748
rect 4925 1742 5124 1744
rect 5159 1744 5172 1754
rect 5190 1744 5207 1757
rect 5159 1742 5207 1744
rect 4801 1738 4834 1742
rect 4797 1736 4834 1738
rect 4797 1735 4864 1736
rect 4797 1730 4828 1735
rect 4834 1730 4864 1735
rect 4797 1726 4864 1730
rect 4770 1723 4864 1726
rect 4770 1716 4819 1723
rect 4770 1710 4800 1716
rect 4819 1711 4824 1716
rect 4736 1694 4816 1710
rect 4828 1702 4864 1723
rect 4925 1718 5114 1742
rect 5159 1741 5206 1742
rect 5172 1736 5206 1741
rect 5246 1736 5262 1738
rect 4940 1715 5114 1718
rect 4933 1712 5114 1715
rect 5142 1735 5206 1736
rect 4736 1692 4755 1694
rect 4770 1692 4804 1694
rect 4736 1676 4816 1692
rect 4736 1670 4755 1676
rect 4452 1644 4555 1654
rect 4406 1642 4555 1644
rect 4576 1642 4611 1654
rect 4245 1640 4407 1642
rect 4257 1620 4276 1640
rect 4291 1638 4321 1640
rect 4140 1612 4181 1620
rect 4263 1616 4276 1620
rect 4328 1624 4407 1640
rect 4439 1640 4611 1642
rect 4439 1624 4518 1640
rect 4525 1638 4555 1640
rect 4103 1602 4132 1612
rect 4146 1602 4175 1612
rect 4190 1602 4220 1616
rect 4263 1602 4306 1616
rect 4328 1612 4518 1624
rect 4583 1620 4589 1640
rect 4313 1602 4343 1612
rect 4344 1602 4502 1612
rect 4506 1602 4536 1612
rect 4540 1602 4570 1616
rect 4598 1602 4611 1640
rect 4683 1654 4712 1670
rect 4726 1654 4755 1670
rect 4770 1660 4800 1676
rect 4828 1654 4834 1702
rect 4837 1696 4856 1702
rect 4871 1696 4901 1704
rect 4837 1688 4901 1696
rect 4837 1672 4917 1688
rect 4933 1681 4995 1712
rect 5011 1681 5073 1712
rect 5142 1710 5191 1735
rect 5236 1726 5262 1736
rect 5206 1710 5262 1726
rect 5105 1696 5135 1704
rect 5142 1702 5252 1710
rect 5105 1688 5150 1696
rect 4837 1670 4856 1672
rect 4871 1670 4917 1672
rect 4837 1654 4917 1670
rect 4944 1668 4979 1681
rect 5020 1678 5057 1681
rect 5020 1676 5062 1678
rect 4949 1665 4979 1668
rect 4958 1661 4965 1665
rect 4965 1660 4966 1661
rect 4924 1654 4934 1660
rect 4683 1646 4718 1654
rect 4683 1620 4684 1646
rect 4691 1620 4718 1646
rect 4626 1602 4656 1616
rect 4683 1612 4718 1620
rect 4720 1646 4761 1654
rect 4720 1620 4735 1646
rect 4742 1620 4761 1646
rect 4825 1642 4856 1654
rect 4871 1642 4974 1654
rect 4986 1644 5012 1670
rect 5027 1665 5057 1676
rect 5089 1672 5151 1688
rect 5089 1670 5135 1672
rect 5089 1654 5151 1670
rect 5163 1654 5169 1702
rect 5172 1694 5252 1702
rect 5172 1692 5191 1694
rect 5206 1692 5240 1694
rect 5172 1676 5252 1692
rect 5172 1654 5191 1676
rect 5206 1660 5236 1676
rect 5264 1670 5270 1744
rect 5273 1670 5292 1814
rect 5307 1670 5313 1814
rect 5322 1744 5335 1814
rect 5380 1798 5397 1802
rect 5401 1800 5409 1802
rect 5399 1798 5409 1800
rect 5380 1788 5409 1798
rect 5462 1788 5478 1802
rect 5516 1798 5522 1800
rect 5529 1798 5637 1814
rect 5644 1798 5650 1800
rect 5658 1798 5673 1814
rect 5739 1808 5758 1811
rect 5380 1786 5478 1788
rect 5505 1786 5673 1798
rect 5688 1788 5704 1802
rect 5739 1789 5761 1808
rect 5771 1802 5787 1803
rect 5770 1800 5787 1802
rect 5771 1795 5787 1800
rect 5761 1788 5767 1789
rect 5770 1788 5799 1795
rect 5688 1787 5799 1788
rect 5688 1786 5805 1787
rect 5364 1778 5415 1786
rect 5462 1778 5496 1786
rect 5364 1766 5389 1778
rect 5396 1766 5415 1778
rect 5469 1776 5496 1778
rect 5505 1776 5726 1786
rect 5761 1783 5767 1786
rect 5469 1772 5726 1776
rect 5364 1758 5415 1766
rect 5462 1758 5726 1772
rect 5770 1778 5805 1786
rect 5316 1710 5335 1744
rect 5380 1750 5409 1758
rect 5380 1744 5397 1750
rect 5380 1742 5414 1744
rect 5462 1742 5478 1758
rect 5479 1748 5687 1758
rect 5688 1748 5704 1758
rect 5752 1754 5767 1769
rect 5770 1766 5771 1778
rect 5778 1766 5805 1778
rect 5770 1758 5805 1766
rect 5770 1757 5799 1758
rect 5490 1744 5704 1748
rect 5505 1742 5704 1744
rect 5739 1744 5752 1754
rect 5770 1744 5787 1757
rect 5739 1742 5787 1744
rect 5381 1738 5414 1742
rect 5377 1736 5414 1738
rect 5377 1735 5444 1736
rect 5377 1730 5408 1735
rect 5414 1730 5444 1735
rect 5377 1726 5444 1730
rect 5350 1723 5444 1726
rect 5350 1716 5399 1723
rect 5350 1710 5380 1716
rect 5399 1711 5404 1716
rect 5316 1694 5396 1710
rect 5408 1702 5444 1723
rect 5505 1718 5694 1742
rect 5739 1741 5786 1742
rect 5752 1736 5786 1741
rect 5520 1715 5694 1718
rect 5513 1712 5694 1715
rect 5722 1735 5786 1736
rect 5316 1692 5335 1694
rect 5350 1692 5384 1694
rect 5316 1676 5396 1692
rect 5316 1670 5335 1676
rect 5032 1644 5135 1654
rect 4986 1642 5135 1644
rect 5156 1642 5191 1654
rect 4825 1640 4987 1642
rect 4837 1620 4856 1640
rect 4871 1638 4901 1640
rect 4720 1612 4761 1620
rect 4843 1616 4856 1620
rect 4908 1624 4987 1640
rect 5019 1640 5191 1642
rect 5019 1624 5098 1640
rect 5105 1638 5135 1640
rect 4683 1602 4712 1612
rect 4726 1602 4755 1612
rect 4770 1602 4800 1616
rect 4843 1602 4886 1616
rect 4908 1612 5098 1624
rect 5163 1620 5169 1640
rect 4893 1602 4923 1612
rect 4924 1602 5082 1612
rect 5086 1602 5116 1612
rect 5120 1602 5150 1616
rect 5178 1602 5191 1640
rect 5263 1654 5292 1670
rect 5306 1654 5335 1670
rect 5350 1660 5380 1676
rect 5408 1654 5414 1702
rect 5417 1696 5436 1702
rect 5451 1696 5481 1704
rect 5417 1688 5481 1696
rect 5417 1672 5497 1688
rect 5513 1681 5575 1712
rect 5591 1681 5653 1712
rect 5722 1710 5771 1735
rect 5786 1710 5816 1728
rect 5685 1696 5715 1704
rect 5722 1702 5832 1710
rect 5685 1688 5730 1696
rect 5417 1670 5436 1672
rect 5451 1670 5497 1672
rect 5417 1654 5497 1670
rect 5524 1668 5559 1681
rect 5600 1678 5637 1681
rect 5600 1676 5642 1678
rect 5529 1665 5559 1668
rect 5538 1661 5545 1665
rect 5545 1660 5546 1661
rect 5504 1654 5514 1660
rect 5263 1646 5298 1654
rect 5263 1620 5264 1646
rect 5271 1620 5298 1646
rect 5206 1602 5236 1616
rect 5263 1612 5298 1620
rect 5300 1646 5341 1654
rect 5300 1620 5315 1646
rect 5322 1620 5341 1646
rect 5405 1642 5436 1654
rect 5451 1642 5554 1654
rect 5566 1644 5592 1670
rect 5607 1665 5637 1676
rect 5669 1672 5731 1688
rect 5669 1670 5715 1672
rect 5669 1654 5731 1670
rect 5743 1654 5749 1702
rect 5752 1694 5832 1702
rect 5752 1692 5771 1694
rect 5786 1692 5820 1694
rect 5752 1677 5832 1692
rect 5752 1676 5838 1677
rect 5752 1654 5771 1676
rect 5786 1660 5816 1676
rect 5844 1670 5850 1744
rect 5853 1670 5872 1814
rect 5887 1670 5893 1814
rect 5902 1744 5915 1814
rect 5960 1798 5977 1802
rect 5981 1800 5989 1802
rect 5979 1798 5989 1800
rect 5960 1788 5989 1798
rect 6042 1788 6058 1802
rect 6096 1798 6102 1800
rect 6109 1798 6217 1814
rect 6224 1798 6230 1800
rect 6238 1798 6253 1814
rect 6319 1808 6338 1811
rect 5960 1786 6058 1788
rect 6085 1786 6253 1798
rect 6268 1788 6284 1802
rect 6319 1789 6341 1808
rect 6351 1802 6367 1803
rect 6350 1800 6367 1802
rect 6351 1795 6367 1800
rect 6341 1788 6347 1789
rect 6350 1788 6379 1795
rect 6268 1787 6379 1788
rect 6268 1786 6385 1787
rect 5944 1778 5995 1786
rect 6042 1778 6076 1786
rect 5944 1766 5969 1778
rect 5976 1766 5995 1778
rect 6049 1776 6076 1778
rect 6085 1776 6306 1786
rect 6341 1783 6347 1786
rect 6049 1772 6306 1776
rect 5944 1758 5995 1766
rect 6042 1758 6306 1772
rect 6350 1778 6385 1786
rect 5896 1710 5915 1744
rect 5960 1750 5989 1758
rect 5960 1744 5977 1750
rect 5960 1742 5994 1744
rect 6042 1742 6058 1758
rect 6059 1748 6267 1758
rect 6268 1748 6284 1758
rect 6332 1754 6347 1769
rect 6350 1766 6351 1778
rect 6358 1766 6385 1778
rect 6350 1758 6385 1766
rect 6350 1757 6379 1758
rect 6070 1744 6284 1748
rect 6085 1742 6284 1744
rect 6319 1744 6332 1754
rect 6350 1744 6367 1757
rect 6319 1742 6367 1744
rect 5961 1738 5994 1742
rect 5957 1736 5994 1738
rect 5957 1735 6024 1736
rect 5957 1730 5988 1735
rect 5994 1730 6024 1735
rect 5957 1726 6024 1730
rect 5930 1723 6024 1726
rect 5930 1716 5979 1723
rect 5930 1710 5960 1716
rect 5979 1711 5984 1716
rect 5896 1694 5976 1710
rect 5988 1702 6024 1723
rect 6085 1718 6274 1742
rect 6319 1741 6366 1742
rect 6332 1736 6366 1741
rect 6100 1715 6274 1718
rect 6093 1712 6274 1715
rect 6302 1735 6366 1736
rect 5896 1692 5915 1694
rect 5930 1692 5964 1694
rect 5896 1676 5976 1692
rect 5896 1670 5915 1676
rect 5612 1644 5715 1654
rect 5566 1642 5715 1644
rect 5736 1642 5771 1654
rect 5405 1640 5567 1642
rect 5417 1620 5436 1640
rect 5451 1638 5481 1640
rect 5300 1612 5341 1620
rect 5423 1616 5436 1620
rect 5488 1624 5567 1640
rect 5599 1640 5771 1642
rect 5599 1624 5678 1640
rect 5685 1638 5715 1640
rect 5263 1602 5292 1612
rect 5306 1602 5335 1612
rect 5350 1602 5380 1616
rect 5423 1602 5466 1616
rect 5488 1612 5678 1624
rect 5743 1620 5749 1640
rect 5473 1602 5503 1612
rect 5504 1602 5662 1612
rect 5666 1602 5696 1612
rect 5700 1602 5730 1616
rect 5758 1602 5771 1640
rect 5843 1654 5872 1670
rect 5886 1654 5915 1670
rect 5930 1660 5960 1676
rect 5988 1654 5994 1702
rect 5997 1696 6016 1702
rect 6031 1696 6061 1704
rect 5997 1688 6061 1696
rect 5997 1672 6077 1688
rect 6093 1681 6155 1712
rect 6171 1681 6233 1712
rect 6302 1710 6351 1735
rect 6366 1710 6396 1726
rect 6265 1696 6295 1704
rect 6302 1702 6412 1710
rect 6265 1688 6310 1696
rect 5997 1670 6016 1672
rect 6031 1670 6077 1672
rect 5997 1654 6077 1670
rect 6104 1668 6139 1681
rect 6180 1678 6217 1681
rect 6180 1676 6222 1678
rect 6109 1665 6139 1668
rect 6118 1661 6125 1665
rect 6125 1660 6126 1661
rect 6084 1654 6094 1660
rect 5843 1646 5878 1654
rect 5843 1620 5844 1646
rect 5851 1620 5878 1646
rect 5786 1602 5816 1616
rect 5843 1612 5878 1620
rect 5880 1646 5921 1654
rect 5880 1620 5895 1646
rect 5902 1620 5921 1646
rect 5985 1642 6016 1654
rect 6031 1642 6134 1654
rect 6146 1644 6172 1670
rect 6187 1665 6217 1676
rect 6249 1672 6311 1688
rect 6249 1670 6295 1672
rect 6249 1654 6311 1670
rect 6323 1654 6329 1702
rect 6332 1694 6412 1702
rect 6332 1692 6351 1694
rect 6366 1692 6400 1694
rect 6332 1676 6412 1692
rect 6332 1654 6351 1676
rect 6366 1660 6396 1676
rect 6424 1670 6430 1744
rect 6439 1670 6452 1814
rect 6192 1644 6295 1654
rect 6146 1642 6295 1644
rect 6316 1642 6351 1654
rect 5985 1640 6147 1642
rect 5997 1620 6016 1640
rect 6031 1638 6061 1640
rect 5880 1612 5921 1620
rect 6003 1616 6016 1620
rect 6068 1624 6147 1640
rect 6179 1640 6351 1642
rect 6179 1624 6258 1640
rect 6265 1638 6295 1640
rect 5843 1602 5872 1612
rect 5886 1602 5915 1612
rect 5930 1602 5960 1616
rect 6003 1602 6046 1616
rect 6068 1612 6258 1624
rect 6323 1620 6329 1640
rect 6053 1602 6083 1612
rect 6084 1602 6242 1612
rect 6246 1602 6276 1612
rect 6280 1602 6310 1616
rect 6338 1602 6351 1640
rect 6423 1654 6452 1670
rect 6423 1646 6458 1654
rect 6423 1620 6424 1646
rect 6431 1620 6458 1646
rect 6366 1602 6396 1616
rect 6423 1612 6458 1620
rect 6423 1602 6452 1612
rect -541 1588 6452 1602
rect -478 1558 -465 1588
rect -450 1574 -420 1588
rect -377 1574 -334 1588
rect -327 1574 -107 1588
rect -100 1574 -70 1588
rect -410 1560 -395 1572
rect -376 1560 -363 1574
rect -295 1570 -142 1574
rect -413 1558 -391 1560
rect -313 1558 -121 1570
rect -42 1558 -29 1588
rect -14 1574 16 1588
rect 53 1558 72 1588
rect 87 1558 93 1588
rect 102 1558 115 1588
rect 130 1574 160 1588
rect 203 1574 246 1588
rect 253 1574 473 1588
rect 480 1574 510 1588
rect 170 1560 185 1572
rect 204 1560 217 1574
rect 285 1570 438 1574
rect 167 1558 189 1560
rect 267 1558 459 1570
rect 538 1558 551 1588
rect 566 1574 596 1588
rect 633 1558 652 1588
rect 667 1558 673 1588
rect 682 1558 695 1588
rect 710 1574 740 1588
rect 783 1574 826 1588
rect 833 1574 1053 1588
rect 1060 1574 1090 1588
rect 750 1560 765 1572
rect 784 1560 797 1574
rect 865 1570 1018 1574
rect 747 1558 769 1560
rect 847 1558 1039 1570
rect 1118 1558 1131 1588
rect 1146 1574 1176 1588
rect 1213 1558 1232 1588
rect 1247 1558 1253 1588
rect 1262 1558 1275 1588
rect 1290 1574 1320 1588
rect 1363 1574 1406 1588
rect 1413 1574 1633 1588
rect 1640 1574 1670 1588
rect 1330 1560 1345 1572
rect 1364 1560 1377 1574
rect 1445 1570 1598 1574
rect 1327 1558 1349 1560
rect 1427 1558 1619 1570
rect 1698 1558 1711 1588
rect 1726 1574 1756 1588
rect 1793 1558 1812 1588
rect 1827 1558 1833 1588
rect 1842 1558 1855 1588
rect 1870 1574 1900 1588
rect 1943 1574 1986 1588
rect 1993 1574 2213 1588
rect 2220 1574 2250 1588
rect 1910 1560 1925 1572
rect 1944 1560 1957 1574
rect 2025 1570 2178 1574
rect 1907 1558 1929 1560
rect 2007 1558 2199 1570
rect 2278 1558 2291 1588
rect 2306 1574 2336 1588
rect 2373 1558 2392 1588
rect 2407 1558 2413 1588
rect 2422 1558 2435 1588
rect 2450 1574 2480 1588
rect 2523 1574 2566 1588
rect 2573 1574 2793 1588
rect 2800 1574 2830 1588
rect 2490 1560 2505 1572
rect 2524 1560 2537 1574
rect 2605 1570 2758 1574
rect 2487 1558 2509 1560
rect 2587 1558 2779 1570
rect 2858 1558 2871 1588
rect 2886 1574 2916 1588
rect 2953 1558 2972 1588
rect 2987 1558 2993 1588
rect 3002 1558 3015 1588
rect 3030 1574 3060 1588
rect 3103 1574 3146 1588
rect 3153 1574 3373 1588
rect 3380 1574 3410 1588
rect 3070 1560 3085 1572
rect 3104 1560 3117 1574
rect 3185 1570 3338 1574
rect 3067 1558 3089 1560
rect 3167 1558 3359 1570
rect 3438 1558 3451 1588
rect 3466 1574 3496 1588
rect 3533 1558 3552 1588
rect 3567 1558 3573 1588
rect 3582 1558 3595 1588
rect 3610 1574 3640 1588
rect 3683 1574 3726 1588
rect 3733 1574 3953 1588
rect 3960 1574 3990 1588
rect 3650 1560 3665 1572
rect 3684 1560 3697 1574
rect 3765 1570 3918 1574
rect 3647 1558 3669 1560
rect 3747 1558 3939 1570
rect 4018 1558 4031 1588
rect 4046 1574 4076 1588
rect 4113 1558 4132 1588
rect 4147 1558 4153 1588
rect 4162 1558 4175 1588
rect 4190 1574 4220 1588
rect 4263 1574 4306 1588
rect 4313 1574 4533 1588
rect 4540 1574 4570 1588
rect 4230 1560 4245 1572
rect 4264 1560 4277 1574
rect 4345 1570 4498 1574
rect 4227 1558 4249 1560
rect 4327 1558 4519 1570
rect 4598 1558 4611 1588
rect 4626 1574 4656 1588
rect 4693 1558 4712 1588
rect 4727 1558 4733 1588
rect 4742 1558 4755 1588
rect 4770 1574 4800 1588
rect 4843 1574 4886 1588
rect 4893 1574 5113 1588
rect 5120 1574 5150 1588
rect 4810 1560 4825 1572
rect 4844 1560 4857 1574
rect 4925 1570 5078 1574
rect 4807 1558 4829 1560
rect 4907 1558 5099 1570
rect 5178 1558 5191 1588
rect 5206 1574 5236 1588
rect 5273 1558 5292 1588
rect 5307 1558 5313 1588
rect 5322 1558 5335 1588
rect 5350 1574 5380 1588
rect 5423 1574 5466 1588
rect 5473 1574 5693 1588
rect 5700 1574 5730 1588
rect 5390 1560 5405 1572
rect 5424 1560 5437 1574
rect 5505 1570 5658 1574
rect 5387 1558 5409 1560
rect 5487 1558 5679 1570
rect 5758 1558 5771 1588
rect 5786 1574 5816 1588
rect 5853 1558 5872 1588
rect 5887 1558 5893 1588
rect 5902 1558 5915 1588
rect 5930 1574 5960 1588
rect 6003 1574 6046 1588
rect 6053 1574 6273 1588
rect 6280 1574 6310 1588
rect 5970 1560 5985 1572
rect 6004 1560 6017 1574
rect 6085 1570 6238 1574
rect 5967 1558 5989 1560
rect 6067 1558 6259 1570
rect 6338 1558 6351 1588
rect 6366 1574 6396 1588
rect 6439 1558 6452 1588
rect -541 1544 6452 1558
rect -478 1474 -465 1544
rect -413 1540 -391 1544
rect -420 1528 -403 1532
rect -399 1530 -391 1532
rect -401 1528 -391 1530
rect -420 1518 -391 1528
rect -338 1518 -322 1532
rect -284 1528 -278 1530
rect -271 1528 -163 1544
rect -156 1528 -150 1530
rect -142 1528 -127 1544
rect -61 1538 -42 1541
rect -420 1516 -322 1518
rect -295 1516 -127 1528
rect -112 1518 -96 1532
rect -61 1519 -39 1538
rect -29 1532 -13 1533
rect -30 1530 -13 1532
rect -29 1525 -13 1530
rect -39 1518 -33 1519
rect -30 1518 -1 1525
rect -112 1517 -1 1518
rect -112 1516 5 1517
rect -436 1508 -385 1516
rect -338 1508 -304 1516
rect -436 1496 -411 1508
rect -404 1496 -385 1508
rect -331 1506 -304 1508
rect -295 1506 -74 1516
rect -39 1513 -33 1516
rect -331 1502 -74 1506
rect -436 1488 -385 1496
rect -338 1488 -74 1502
rect -30 1508 5 1516
rect -484 1440 -465 1474
rect -420 1480 -391 1488
rect -420 1474 -403 1480
rect -420 1472 -386 1474
rect -338 1472 -322 1488
rect -321 1478 -113 1488
rect -112 1478 -96 1488
rect -48 1484 -33 1499
rect -30 1496 -29 1508
rect -22 1496 5 1508
rect -30 1488 5 1496
rect -30 1487 -1 1488
rect -310 1474 -96 1478
rect -295 1472 -96 1474
rect -61 1474 -48 1484
rect -30 1474 -13 1487
rect -61 1472 -13 1474
rect -419 1468 -386 1472
rect -423 1466 -386 1468
rect -423 1465 -356 1466
rect -423 1460 -392 1465
rect -386 1460 -356 1465
rect -423 1456 -356 1460
rect -450 1453 -356 1456
rect -450 1446 -401 1453
rect -450 1440 -420 1446
rect -401 1441 -396 1446
rect -484 1424 -404 1440
rect -392 1432 -356 1453
rect -295 1448 -106 1472
rect -61 1471 -14 1472
rect -48 1466 -14 1471
rect -280 1445 -106 1448
rect -287 1442 -106 1445
rect -78 1465 -14 1466
rect -484 1422 -465 1424
rect -450 1422 -416 1424
rect -484 1406 -404 1422
rect -484 1400 -465 1406
rect -494 1384 -465 1400
rect -450 1390 -420 1406
rect -392 1384 -386 1432
rect -383 1426 -364 1432
rect -349 1426 -319 1434
rect -383 1418 -319 1426
rect -383 1402 -303 1418
rect -287 1411 -225 1442
rect -209 1411 -147 1442
rect -78 1440 -29 1465
rect -14 1440 16 1458
rect -115 1426 -85 1434
rect -78 1432 32 1440
rect -115 1418 -70 1426
rect -383 1400 -364 1402
rect -349 1400 -303 1402
rect -383 1384 -303 1400
rect -276 1398 -241 1411
rect -200 1408 -163 1411
rect -200 1406 -158 1408
rect -271 1395 -241 1398
rect -262 1391 -255 1395
rect -255 1390 -254 1391
rect -296 1384 -286 1390
rect -500 1376 -459 1384
rect -500 1350 -485 1376
rect -478 1350 -459 1376
rect -395 1372 -364 1384
rect -349 1372 -246 1384
rect -234 1374 -208 1400
rect -193 1395 -163 1406
rect -131 1402 -69 1418
rect -131 1400 -85 1402
rect -131 1384 -69 1400
rect -57 1384 -51 1432
rect -48 1424 32 1432
rect -48 1422 -29 1424
rect -14 1422 20 1424
rect -48 1407 32 1422
rect -48 1406 38 1407
rect -48 1384 -29 1406
rect -14 1390 16 1406
rect 44 1400 50 1474
rect 53 1400 72 1544
rect 87 1400 93 1544
rect 102 1474 115 1544
rect 167 1540 189 1544
rect 160 1528 177 1532
rect 181 1530 189 1532
rect 179 1528 189 1530
rect 160 1518 189 1528
rect 242 1518 258 1532
rect 296 1528 302 1530
rect 309 1528 417 1544
rect 424 1528 430 1530
rect 438 1528 453 1544
rect 519 1538 538 1541
rect 160 1516 258 1518
rect 285 1516 453 1528
rect 468 1518 484 1532
rect 519 1519 541 1538
rect 551 1532 567 1533
rect 550 1530 567 1532
rect 551 1525 567 1530
rect 541 1518 547 1519
rect 550 1518 579 1525
rect 468 1517 579 1518
rect 468 1516 585 1517
rect 144 1508 195 1516
rect 242 1508 276 1516
rect 144 1496 169 1508
rect 176 1496 195 1508
rect 249 1506 276 1508
rect 285 1506 506 1516
rect 541 1513 547 1516
rect 249 1502 506 1506
rect 144 1488 195 1496
rect 242 1488 506 1502
rect 550 1508 585 1516
rect 96 1440 115 1474
rect 160 1480 189 1488
rect 160 1474 177 1480
rect 160 1472 194 1474
rect 242 1472 258 1488
rect 259 1478 467 1488
rect 468 1478 484 1488
rect 532 1484 547 1499
rect 550 1496 551 1508
rect 558 1496 585 1508
rect 550 1488 585 1496
rect 550 1487 579 1488
rect 270 1474 484 1478
rect 285 1472 484 1474
rect 519 1474 532 1484
rect 550 1474 567 1487
rect 519 1472 567 1474
rect 161 1468 194 1472
rect 157 1466 194 1468
rect 157 1465 224 1466
rect 157 1460 188 1465
rect 194 1460 224 1465
rect 157 1456 224 1460
rect 130 1453 224 1456
rect 130 1446 179 1453
rect 130 1440 160 1446
rect 179 1441 184 1446
rect 96 1424 176 1440
rect 188 1432 224 1453
rect 285 1448 474 1472
rect 519 1471 566 1472
rect 532 1466 566 1471
rect 606 1466 622 1468
rect 300 1445 474 1448
rect 293 1442 474 1445
rect 502 1465 566 1466
rect 96 1422 115 1424
rect 130 1422 164 1424
rect 96 1406 176 1422
rect 96 1400 115 1406
rect -188 1374 -85 1384
rect -234 1372 -85 1374
rect -64 1372 -29 1384
rect -395 1370 -233 1372
rect -383 1352 -364 1370
rect -349 1368 -319 1370
rect -500 1342 -459 1350
rect -376 1346 -364 1352
rect -312 1352 -233 1370
rect -201 1370 -29 1372
rect -201 1354 -122 1370
rect -115 1368 -85 1370
rect -226 1352 -122 1354
rect -494 1332 -465 1342
rect -450 1332 -420 1346
rect -376 1332 -334 1346
rect -312 1342 -122 1352
rect -57 1350 -51 1370
rect -327 1332 -297 1342
rect -296 1332 -138 1342
rect -134 1332 -104 1342
rect -100 1332 -70 1346
rect -42 1332 -29 1370
rect 43 1384 72 1400
rect 86 1384 115 1400
rect 130 1390 160 1406
rect 188 1384 194 1432
rect 197 1426 216 1432
rect 231 1426 261 1434
rect 197 1418 261 1426
rect 197 1402 277 1418
rect 293 1411 355 1442
rect 371 1411 433 1442
rect 502 1440 551 1465
rect 596 1456 622 1466
rect 566 1440 622 1456
rect 465 1426 495 1434
rect 502 1432 612 1440
rect 465 1418 510 1426
rect 197 1400 216 1402
rect 231 1400 277 1402
rect 197 1384 277 1400
rect 304 1398 339 1411
rect 380 1408 417 1411
rect 380 1406 422 1408
rect 309 1395 339 1398
rect 318 1391 325 1395
rect 325 1390 326 1391
rect 284 1384 294 1390
rect 43 1376 78 1384
rect 43 1350 44 1376
rect 51 1350 78 1376
rect -14 1332 16 1346
rect 43 1342 78 1350
rect 80 1376 121 1384
rect 80 1350 95 1376
rect 102 1350 121 1376
rect 185 1372 216 1384
rect 231 1372 334 1384
rect 346 1374 372 1400
rect 387 1395 417 1406
rect 449 1402 511 1418
rect 449 1400 495 1402
rect 449 1384 511 1400
rect 523 1384 529 1432
rect 532 1424 612 1432
rect 532 1422 551 1424
rect 566 1422 600 1424
rect 532 1406 612 1422
rect 532 1384 551 1406
rect 566 1390 596 1406
rect 624 1400 630 1474
rect 633 1400 652 1544
rect 667 1400 673 1544
rect 682 1474 695 1544
rect 747 1540 769 1544
rect 740 1528 757 1532
rect 761 1530 769 1532
rect 759 1528 769 1530
rect 740 1518 769 1528
rect 822 1518 838 1532
rect 876 1528 882 1530
rect 889 1528 997 1544
rect 1004 1528 1010 1530
rect 1018 1528 1033 1544
rect 1099 1538 1118 1541
rect 740 1516 838 1518
rect 865 1516 1033 1528
rect 1048 1518 1064 1532
rect 1099 1519 1121 1538
rect 1131 1532 1147 1533
rect 1130 1530 1147 1532
rect 1131 1525 1147 1530
rect 1121 1518 1127 1519
rect 1130 1518 1159 1525
rect 1048 1517 1159 1518
rect 1048 1516 1165 1517
rect 724 1508 775 1516
rect 822 1508 856 1516
rect 724 1496 749 1508
rect 756 1496 775 1508
rect 829 1506 856 1508
rect 865 1506 1086 1516
rect 1121 1513 1127 1516
rect 829 1502 1086 1506
rect 724 1488 775 1496
rect 822 1488 1086 1502
rect 1130 1508 1165 1516
rect 676 1440 695 1474
rect 740 1480 769 1488
rect 740 1474 757 1480
rect 740 1472 774 1474
rect 822 1472 838 1488
rect 839 1478 1047 1488
rect 1048 1478 1064 1488
rect 1112 1484 1127 1499
rect 1130 1496 1131 1508
rect 1138 1496 1165 1508
rect 1130 1488 1165 1496
rect 1130 1487 1159 1488
rect 850 1474 1064 1478
rect 865 1472 1064 1474
rect 1099 1474 1112 1484
rect 1130 1474 1147 1487
rect 1099 1472 1147 1474
rect 741 1468 774 1472
rect 737 1466 774 1468
rect 737 1465 804 1466
rect 737 1460 768 1465
rect 774 1460 804 1465
rect 737 1456 804 1460
rect 710 1453 804 1456
rect 710 1446 759 1453
rect 710 1440 740 1446
rect 759 1441 764 1446
rect 676 1424 756 1440
rect 768 1432 804 1453
rect 865 1448 1054 1472
rect 1099 1471 1146 1472
rect 1112 1466 1146 1471
rect 880 1445 1054 1448
rect 873 1442 1054 1445
rect 1082 1465 1146 1466
rect 676 1422 695 1424
rect 710 1422 744 1424
rect 676 1406 756 1422
rect 676 1400 695 1406
rect 392 1374 495 1384
rect 346 1372 495 1374
rect 516 1372 551 1384
rect 185 1370 347 1372
rect 197 1352 216 1370
rect 231 1368 261 1370
rect 80 1342 121 1350
rect 204 1346 216 1352
rect 268 1352 347 1370
rect 379 1370 551 1372
rect 379 1354 458 1370
rect 465 1368 495 1370
rect 354 1352 458 1354
rect 43 1332 72 1342
rect 86 1332 115 1342
rect 130 1332 160 1346
rect 204 1332 246 1346
rect 268 1342 458 1352
rect 523 1350 529 1370
rect 253 1332 283 1342
rect 284 1332 442 1342
rect 446 1332 476 1342
rect 480 1332 510 1346
rect 538 1332 551 1370
rect 623 1384 652 1400
rect 666 1384 695 1400
rect 710 1390 740 1406
rect 768 1384 774 1432
rect 777 1426 796 1432
rect 811 1426 841 1434
rect 777 1418 841 1426
rect 777 1402 857 1418
rect 873 1411 935 1442
rect 951 1411 1013 1442
rect 1082 1440 1131 1465
rect 1146 1440 1176 1458
rect 1045 1426 1075 1434
rect 1082 1432 1192 1440
rect 1045 1418 1090 1426
rect 777 1400 796 1402
rect 811 1400 857 1402
rect 777 1384 857 1400
rect 884 1398 919 1411
rect 960 1408 997 1411
rect 960 1406 1002 1408
rect 889 1395 919 1398
rect 898 1391 905 1395
rect 905 1390 906 1391
rect 864 1384 874 1390
rect 623 1376 658 1384
rect 623 1350 624 1376
rect 631 1350 658 1376
rect 566 1332 596 1346
rect 623 1342 658 1350
rect 660 1376 701 1384
rect 660 1350 675 1376
rect 682 1350 701 1376
rect 765 1372 796 1384
rect 811 1372 914 1384
rect 926 1374 952 1400
rect 967 1395 997 1406
rect 1029 1402 1091 1418
rect 1029 1400 1075 1402
rect 1029 1384 1091 1400
rect 1103 1384 1109 1432
rect 1112 1424 1192 1432
rect 1112 1422 1131 1424
rect 1146 1422 1180 1424
rect 1112 1407 1192 1422
rect 1112 1406 1198 1407
rect 1112 1384 1131 1406
rect 1146 1390 1176 1406
rect 1204 1400 1210 1474
rect 1213 1400 1232 1544
rect 1247 1400 1253 1544
rect 1262 1474 1275 1544
rect 1327 1540 1349 1544
rect 1320 1528 1337 1532
rect 1341 1530 1349 1532
rect 1339 1528 1349 1530
rect 1320 1518 1349 1528
rect 1402 1518 1418 1532
rect 1456 1528 1462 1530
rect 1469 1528 1577 1544
rect 1584 1528 1590 1530
rect 1598 1528 1613 1544
rect 1679 1538 1698 1541
rect 1320 1516 1418 1518
rect 1445 1516 1613 1528
rect 1628 1518 1644 1532
rect 1679 1519 1701 1538
rect 1711 1532 1727 1533
rect 1710 1530 1727 1532
rect 1711 1525 1727 1530
rect 1701 1518 1707 1519
rect 1710 1518 1739 1525
rect 1628 1517 1739 1518
rect 1628 1516 1745 1517
rect 1304 1508 1355 1516
rect 1402 1508 1436 1516
rect 1304 1496 1329 1508
rect 1336 1496 1355 1508
rect 1409 1506 1436 1508
rect 1445 1506 1666 1516
rect 1701 1513 1707 1516
rect 1409 1502 1666 1506
rect 1304 1488 1355 1496
rect 1402 1488 1666 1502
rect 1710 1508 1745 1516
rect 1256 1440 1275 1474
rect 1320 1480 1349 1488
rect 1320 1474 1337 1480
rect 1320 1472 1354 1474
rect 1402 1472 1418 1488
rect 1419 1478 1627 1488
rect 1628 1478 1644 1488
rect 1692 1484 1707 1499
rect 1710 1496 1711 1508
rect 1718 1496 1745 1508
rect 1710 1488 1745 1496
rect 1710 1487 1739 1488
rect 1430 1474 1644 1478
rect 1445 1472 1644 1474
rect 1679 1474 1692 1484
rect 1710 1474 1727 1487
rect 1679 1472 1727 1474
rect 1321 1468 1354 1472
rect 1317 1466 1354 1468
rect 1317 1465 1384 1466
rect 1317 1460 1348 1465
rect 1354 1460 1384 1465
rect 1317 1456 1384 1460
rect 1290 1453 1384 1456
rect 1290 1446 1339 1453
rect 1290 1440 1320 1446
rect 1339 1441 1344 1446
rect 1256 1424 1336 1440
rect 1348 1432 1384 1453
rect 1445 1448 1634 1472
rect 1679 1471 1726 1472
rect 1692 1466 1726 1471
rect 1766 1466 1782 1468
rect 1460 1445 1634 1448
rect 1453 1442 1634 1445
rect 1662 1465 1726 1466
rect 1256 1422 1275 1424
rect 1290 1422 1324 1424
rect 1256 1406 1336 1422
rect 1256 1400 1275 1406
rect 972 1374 1075 1384
rect 926 1372 1075 1374
rect 1096 1372 1131 1384
rect 765 1370 927 1372
rect 777 1352 796 1370
rect 811 1368 841 1370
rect 660 1342 701 1350
rect 784 1346 796 1352
rect 848 1352 927 1370
rect 959 1370 1131 1372
rect 959 1354 1038 1370
rect 1045 1368 1075 1370
rect 934 1352 1038 1354
rect 623 1332 652 1342
rect 666 1332 695 1342
rect 710 1332 740 1346
rect 784 1332 826 1346
rect 848 1342 1038 1352
rect 1103 1350 1109 1370
rect 833 1332 863 1342
rect 864 1332 1022 1342
rect 1026 1332 1056 1342
rect 1060 1332 1090 1346
rect 1118 1332 1131 1370
rect 1203 1384 1232 1400
rect 1246 1384 1275 1400
rect 1290 1390 1320 1406
rect 1348 1384 1354 1432
rect 1357 1426 1376 1432
rect 1391 1426 1421 1434
rect 1357 1418 1421 1426
rect 1357 1402 1437 1418
rect 1453 1411 1515 1442
rect 1531 1411 1593 1442
rect 1662 1440 1711 1465
rect 1756 1456 1782 1466
rect 1726 1440 1782 1456
rect 1625 1426 1655 1434
rect 1662 1432 1772 1440
rect 1625 1418 1670 1426
rect 1357 1400 1376 1402
rect 1391 1400 1437 1402
rect 1357 1384 1437 1400
rect 1464 1398 1499 1411
rect 1540 1408 1577 1411
rect 1540 1406 1582 1408
rect 1469 1395 1499 1398
rect 1478 1391 1485 1395
rect 1485 1390 1486 1391
rect 1444 1384 1454 1390
rect 1203 1376 1238 1384
rect 1203 1350 1204 1376
rect 1211 1350 1238 1376
rect 1146 1332 1176 1346
rect 1203 1342 1238 1350
rect 1240 1376 1281 1384
rect 1240 1350 1255 1376
rect 1262 1350 1281 1376
rect 1345 1372 1376 1384
rect 1391 1372 1494 1384
rect 1506 1374 1532 1400
rect 1547 1395 1577 1406
rect 1609 1402 1671 1418
rect 1609 1400 1655 1402
rect 1609 1384 1671 1400
rect 1683 1384 1689 1432
rect 1692 1424 1772 1432
rect 1692 1422 1711 1424
rect 1726 1422 1760 1424
rect 1692 1406 1772 1422
rect 1692 1384 1711 1406
rect 1726 1390 1756 1406
rect 1784 1400 1790 1474
rect 1793 1400 1812 1544
rect 1827 1400 1833 1544
rect 1842 1474 1855 1544
rect 1907 1540 1929 1544
rect 1900 1528 1917 1532
rect 1921 1530 1929 1532
rect 1919 1528 1929 1530
rect 1900 1518 1929 1528
rect 1982 1518 1998 1532
rect 2036 1528 2042 1530
rect 2049 1528 2157 1544
rect 2164 1528 2170 1530
rect 2178 1528 2193 1544
rect 2259 1538 2278 1541
rect 1900 1516 1998 1518
rect 2025 1516 2193 1528
rect 2208 1518 2224 1532
rect 2259 1519 2281 1538
rect 2291 1532 2307 1533
rect 2290 1530 2307 1532
rect 2291 1525 2307 1530
rect 2281 1518 2287 1519
rect 2290 1518 2319 1525
rect 2208 1517 2319 1518
rect 2208 1516 2325 1517
rect 1884 1508 1935 1516
rect 1982 1508 2016 1516
rect 1884 1496 1909 1508
rect 1916 1496 1935 1508
rect 1989 1506 2016 1508
rect 2025 1506 2246 1516
rect 2281 1513 2287 1516
rect 1989 1502 2246 1506
rect 1884 1488 1935 1496
rect 1982 1488 2246 1502
rect 2290 1508 2325 1516
rect 1836 1440 1855 1474
rect 1900 1480 1929 1488
rect 1900 1474 1917 1480
rect 1900 1472 1934 1474
rect 1982 1472 1998 1488
rect 1999 1478 2207 1488
rect 2208 1478 2224 1488
rect 2272 1484 2287 1499
rect 2290 1496 2291 1508
rect 2298 1496 2325 1508
rect 2290 1488 2325 1496
rect 2290 1487 2319 1488
rect 2010 1474 2224 1478
rect 2025 1472 2224 1474
rect 2259 1474 2272 1484
rect 2290 1474 2307 1487
rect 2259 1472 2307 1474
rect 1901 1468 1934 1472
rect 1897 1466 1934 1468
rect 1897 1465 1964 1466
rect 1897 1460 1928 1465
rect 1934 1460 1964 1465
rect 1897 1456 1964 1460
rect 1870 1453 1964 1456
rect 1870 1446 1919 1453
rect 1870 1440 1900 1446
rect 1919 1441 1924 1446
rect 1836 1424 1916 1440
rect 1928 1432 1964 1453
rect 2025 1448 2214 1472
rect 2259 1471 2306 1472
rect 2272 1466 2306 1471
rect 2040 1445 2214 1448
rect 2033 1442 2214 1445
rect 2242 1465 2306 1466
rect 1836 1422 1855 1424
rect 1870 1422 1904 1424
rect 1836 1406 1916 1422
rect 1836 1400 1855 1406
rect 1552 1374 1655 1384
rect 1506 1372 1655 1374
rect 1676 1372 1711 1384
rect 1345 1370 1507 1372
rect 1357 1352 1376 1370
rect 1391 1368 1421 1370
rect 1240 1342 1281 1350
rect 1364 1346 1376 1352
rect 1428 1352 1507 1370
rect 1539 1370 1711 1372
rect 1539 1354 1618 1370
rect 1625 1368 1655 1370
rect 1514 1352 1618 1354
rect 1203 1332 1232 1342
rect 1246 1332 1275 1342
rect 1290 1332 1320 1346
rect 1364 1332 1406 1346
rect 1428 1342 1618 1352
rect 1683 1350 1689 1370
rect 1413 1332 1443 1342
rect 1444 1332 1602 1342
rect 1606 1332 1636 1342
rect 1640 1332 1670 1346
rect 1698 1332 1711 1370
rect 1783 1384 1812 1400
rect 1826 1384 1855 1400
rect 1870 1390 1900 1406
rect 1928 1384 1934 1432
rect 1937 1426 1956 1432
rect 1971 1426 2001 1434
rect 1937 1418 2001 1426
rect 1937 1402 2017 1418
rect 2033 1411 2095 1442
rect 2111 1411 2173 1442
rect 2242 1440 2291 1465
rect 2306 1440 2336 1458
rect 2205 1426 2235 1434
rect 2242 1432 2352 1440
rect 2205 1418 2250 1426
rect 1937 1400 1956 1402
rect 1971 1400 2017 1402
rect 1937 1384 2017 1400
rect 2044 1398 2079 1411
rect 2120 1408 2157 1411
rect 2120 1406 2162 1408
rect 2049 1395 2079 1398
rect 2058 1391 2065 1395
rect 2065 1390 2066 1391
rect 2024 1384 2034 1390
rect 1783 1376 1818 1384
rect 1783 1350 1784 1376
rect 1791 1350 1818 1376
rect 1726 1332 1756 1346
rect 1783 1342 1818 1350
rect 1820 1376 1861 1384
rect 1820 1350 1835 1376
rect 1842 1350 1861 1376
rect 1925 1372 1956 1384
rect 1971 1372 2074 1384
rect 2086 1374 2112 1400
rect 2127 1395 2157 1406
rect 2189 1402 2251 1418
rect 2189 1400 2235 1402
rect 2189 1384 2251 1400
rect 2263 1384 2269 1432
rect 2272 1424 2352 1432
rect 2272 1422 2291 1424
rect 2306 1422 2340 1424
rect 2272 1407 2352 1422
rect 2272 1406 2358 1407
rect 2272 1384 2291 1406
rect 2306 1390 2336 1406
rect 2364 1400 2370 1474
rect 2373 1400 2392 1544
rect 2407 1400 2413 1544
rect 2422 1474 2435 1544
rect 2487 1540 2509 1544
rect 2480 1528 2497 1532
rect 2501 1530 2509 1532
rect 2499 1528 2509 1530
rect 2480 1518 2509 1528
rect 2562 1518 2578 1532
rect 2616 1528 2622 1530
rect 2629 1528 2737 1544
rect 2744 1528 2750 1530
rect 2758 1528 2773 1544
rect 2839 1538 2858 1541
rect 2480 1516 2578 1518
rect 2605 1516 2773 1528
rect 2788 1518 2804 1532
rect 2839 1519 2861 1538
rect 2871 1532 2887 1533
rect 2870 1530 2887 1532
rect 2871 1525 2887 1530
rect 2861 1518 2867 1519
rect 2870 1518 2899 1525
rect 2788 1517 2899 1518
rect 2788 1516 2905 1517
rect 2464 1508 2515 1516
rect 2562 1508 2596 1516
rect 2464 1496 2489 1508
rect 2496 1496 2515 1508
rect 2569 1506 2596 1508
rect 2605 1506 2826 1516
rect 2861 1513 2867 1516
rect 2569 1502 2826 1506
rect 2464 1488 2515 1496
rect 2562 1488 2826 1502
rect 2870 1508 2905 1516
rect 2416 1440 2435 1474
rect 2480 1480 2509 1488
rect 2480 1474 2497 1480
rect 2480 1472 2514 1474
rect 2562 1472 2578 1488
rect 2579 1478 2787 1488
rect 2788 1478 2804 1488
rect 2852 1484 2867 1499
rect 2870 1496 2871 1508
rect 2878 1496 2905 1508
rect 2870 1488 2905 1496
rect 2870 1487 2899 1488
rect 2590 1474 2804 1478
rect 2605 1472 2804 1474
rect 2839 1474 2852 1484
rect 2870 1474 2887 1487
rect 2839 1472 2887 1474
rect 2481 1468 2514 1472
rect 2477 1466 2514 1468
rect 2477 1465 2544 1466
rect 2477 1460 2508 1465
rect 2514 1460 2544 1465
rect 2477 1456 2544 1460
rect 2450 1453 2544 1456
rect 2450 1446 2499 1453
rect 2450 1440 2480 1446
rect 2499 1441 2504 1446
rect 2416 1424 2496 1440
rect 2508 1432 2544 1453
rect 2605 1448 2794 1472
rect 2839 1471 2886 1472
rect 2852 1466 2886 1471
rect 2926 1466 2942 1468
rect 2620 1445 2794 1448
rect 2613 1442 2794 1445
rect 2822 1465 2886 1466
rect 2416 1422 2435 1424
rect 2450 1422 2484 1424
rect 2416 1406 2496 1422
rect 2416 1400 2435 1406
rect 2132 1374 2235 1384
rect 2086 1372 2235 1374
rect 2256 1372 2291 1384
rect 1925 1370 2087 1372
rect 1937 1352 1956 1370
rect 1971 1368 2001 1370
rect 1820 1342 1861 1350
rect 1944 1346 1956 1352
rect 2008 1354 2087 1370
rect 2119 1370 2291 1372
rect 2119 1354 2198 1370
rect 2205 1368 2235 1370
rect 1783 1332 1812 1342
rect 1826 1332 1855 1342
rect 1870 1332 1900 1346
rect 1944 1332 1986 1346
rect 2008 1342 2198 1354
rect 2263 1350 2269 1370
rect 1993 1332 2023 1342
rect 2024 1332 2182 1342
rect 2186 1332 2216 1342
rect 2220 1332 2250 1346
rect 2278 1332 2291 1370
rect 2363 1384 2392 1400
rect 2406 1384 2435 1400
rect 2450 1390 2480 1406
rect 2508 1384 2514 1432
rect 2517 1426 2536 1432
rect 2551 1426 2581 1434
rect 2517 1418 2581 1426
rect 2517 1402 2597 1418
rect 2613 1411 2675 1442
rect 2691 1411 2753 1442
rect 2822 1440 2871 1465
rect 2916 1456 2942 1466
rect 2886 1440 2942 1456
rect 2785 1426 2815 1434
rect 2822 1432 2932 1440
rect 2785 1418 2830 1426
rect 2517 1400 2536 1402
rect 2551 1400 2597 1402
rect 2517 1384 2597 1400
rect 2624 1398 2659 1411
rect 2700 1408 2737 1411
rect 2700 1406 2742 1408
rect 2629 1395 2659 1398
rect 2638 1391 2645 1395
rect 2645 1390 2646 1391
rect 2604 1384 2614 1390
rect 2363 1376 2398 1384
rect 2363 1350 2364 1376
rect 2371 1350 2398 1376
rect 2306 1332 2336 1346
rect 2363 1342 2398 1350
rect 2400 1376 2441 1384
rect 2400 1350 2415 1376
rect 2422 1350 2441 1376
rect 2505 1372 2536 1384
rect 2551 1372 2654 1384
rect 2666 1374 2692 1400
rect 2707 1395 2737 1406
rect 2769 1402 2831 1418
rect 2769 1400 2815 1402
rect 2769 1384 2831 1400
rect 2843 1384 2849 1432
rect 2852 1424 2932 1432
rect 2852 1422 2871 1424
rect 2886 1422 2920 1424
rect 2852 1406 2932 1422
rect 2852 1384 2871 1406
rect 2886 1390 2916 1406
rect 2944 1400 2950 1474
rect 2953 1400 2972 1544
rect 2987 1400 2993 1544
rect 3002 1474 3015 1544
rect 3067 1540 3089 1544
rect 3060 1528 3077 1532
rect 3081 1530 3089 1532
rect 3079 1528 3089 1530
rect 3060 1518 3089 1528
rect 3142 1518 3158 1532
rect 3196 1528 3202 1530
rect 3209 1528 3317 1544
rect 3324 1528 3330 1530
rect 3338 1528 3353 1544
rect 3419 1538 3438 1541
rect 3060 1516 3158 1518
rect 3185 1516 3353 1528
rect 3368 1518 3384 1532
rect 3419 1519 3441 1538
rect 3451 1532 3467 1533
rect 3450 1530 3467 1532
rect 3451 1525 3467 1530
rect 3441 1518 3447 1519
rect 3450 1518 3479 1525
rect 3368 1517 3479 1518
rect 3368 1516 3485 1517
rect 3044 1508 3095 1516
rect 3142 1508 3176 1516
rect 3044 1496 3069 1508
rect 3076 1496 3095 1508
rect 3149 1506 3176 1508
rect 3185 1506 3406 1516
rect 3441 1513 3447 1516
rect 3149 1502 3406 1506
rect 3044 1488 3095 1496
rect 3142 1488 3406 1502
rect 3450 1508 3485 1516
rect 2996 1440 3015 1474
rect 3060 1480 3089 1488
rect 3060 1474 3077 1480
rect 3060 1472 3094 1474
rect 3142 1472 3158 1488
rect 3159 1478 3367 1488
rect 3368 1478 3384 1488
rect 3432 1484 3447 1499
rect 3450 1496 3451 1508
rect 3458 1496 3485 1508
rect 3450 1488 3485 1496
rect 3450 1487 3479 1488
rect 3170 1474 3384 1478
rect 3185 1472 3384 1474
rect 3419 1474 3432 1484
rect 3450 1474 3467 1487
rect 3419 1472 3467 1474
rect 3061 1468 3094 1472
rect 3057 1466 3094 1468
rect 3057 1465 3124 1466
rect 3057 1460 3088 1465
rect 3094 1460 3124 1465
rect 3057 1456 3124 1460
rect 3030 1453 3124 1456
rect 3030 1446 3079 1453
rect 3030 1440 3060 1446
rect 3079 1441 3084 1446
rect 2996 1424 3076 1440
rect 3088 1432 3124 1453
rect 3185 1448 3374 1472
rect 3419 1471 3466 1472
rect 3432 1466 3466 1471
rect 3200 1445 3374 1448
rect 3193 1442 3374 1445
rect 3402 1465 3466 1466
rect 2996 1422 3015 1424
rect 3030 1422 3064 1424
rect 2996 1406 3076 1422
rect 2996 1400 3015 1406
rect 2712 1374 2815 1384
rect 2666 1372 2815 1374
rect 2836 1372 2871 1384
rect 2505 1370 2667 1372
rect 2517 1352 2536 1370
rect 2551 1368 2581 1370
rect 2400 1342 2441 1350
rect 2524 1346 2536 1352
rect 2588 1354 2667 1370
rect 2699 1370 2871 1372
rect 2699 1354 2778 1370
rect 2785 1368 2815 1370
rect 2363 1332 2392 1342
rect 2406 1332 2435 1342
rect 2450 1332 2480 1346
rect 2524 1332 2566 1346
rect 2588 1342 2778 1354
rect 2843 1350 2849 1370
rect 2573 1332 2603 1342
rect 2604 1332 2762 1342
rect 2766 1332 2796 1342
rect 2800 1332 2830 1346
rect 2858 1332 2871 1370
rect 2943 1384 2972 1400
rect 2986 1384 3015 1400
rect 3030 1390 3060 1406
rect 3088 1384 3094 1432
rect 3097 1426 3116 1432
rect 3131 1426 3161 1434
rect 3097 1418 3161 1426
rect 3097 1402 3177 1418
rect 3193 1411 3255 1442
rect 3271 1411 3333 1442
rect 3402 1440 3451 1465
rect 3466 1440 3496 1458
rect 3365 1426 3395 1434
rect 3402 1432 3512 1440
rect 3365 1418 3410 1426
rect 3097 1400 3116 1402
rect 3131 1400 3177 1402
rect 3097 1384 3177 1400
rect 3204 1398 3239 1411
rect 3280 1408 3317 1411
rect 3280 1406 3322 1408
rect 3209 1395 3239 1398
rect 3218 1391 3225 1395
rect 3225 1390 3226 1391
rect 3184 1384 3194 1390
rect 2943 1376 2978 1384
rect 2943 1350 2944 1376
rect 2951 1350 2978 1376
rect 2886 1332 2916 1346
rect 2943 1342 2978 1350
rect 2980 1376 3021 1384
rect 2980 1350 2995 1376
rect 3002 1350 3021 1376
rect 3085 1372 3116 1384
rect 3131 1372 3234 1384
rect 3246 1374 3272 1400
rect 3287 1395 3317 1406
rect 3349 1402 3411 1418
rect 3349 1400 3395 1402
rect 3349 1384 3411 1400
rect 3423 1384 3429 1432
rect 3432 1424 3512 1432
rect 3432 1422 3451 1424
rect 3466 1422 3500 1424
rect 3432 1407 3512 1422
rect 3432 1406 3518 1407
rect 3432 1384 3451 1406
rect 3466 1390 3496 1406
rect 3524 1400 3530 1474
rect 3533 1400 3552 1544
rect 3567 1400 3573 1544
rect 3582 1474 3595 1544
rect 3647 1540 3669 1544
rect 3640 1528 3657 1532
rect 3661 1530 3669 1532
rect 3659 1528 3669 1530
rect 3640 1518 3669 1528
rect 3722 1518 3738 1532
rect 3776 1528 3782 1530
rect 3789 1528 3897 1544
rect 3904 1528 3910 1530
rect 3918 1528 3933 1544
rect 3999 1538 4018 1541
rect 3640 1516 3738 1518
rect 3765 1516 3933 1528
rect 3948 1518 3964 1532
rect 3999 1519 4021 1538
rect 4031 1532 4047 1533
rect 4030 1530 4047 1532
rect 4031 1525 4047 1530
rect 4021 1518 4027 1519
rect 4030 1518 4059 1525
rect 3948 1517 4059 1518
rect 3948 1516 4065 1517
rect 3624 1508 3675 1516
rect 3722 1508 3756 1516
rect 3624 1496 3649 1508
rect 3656 1496 3675 1508
rect 3729 1506 3756 1508
rect 3765 1506 3986 1516
rect 4021 1513 4027 1516
rect 3729 1502 3986 1506
rect 3624 1488 3675 1496
rect 3722 1488 3986 1502
rect 4030 1508 4065 1516
rect 3576 1440 3595 1474
rect 3640 1480 3669 1488
rect 3640 1474 3657 1480
rect 3640 1472 3674 1474
rect 3722 1472 3738 1488
rect 3739 1478 3947 1488
rect 3948 1478 3964 1488
rect 4012 1484 4027 1499
rect 4030 1496 4031 1508
rect 4038 1496 4065 1508
rect 4030 1488 4065 1496
rect 4030 1487 4059 1488
rect 3750 1474 3964 1478
rect 3765 1472 3964 1474
rect 3999 1474 4012 1484
rect 4030 1474 4047 1487
rect 3999 1472 4047 1474
rect 3641 1468 3674 1472
rect 3637 1466 3674 1468
rect 3637 1465 3704 1466
rect 3637 1460 3668 1465
rect 3674 1460 3704 1465
rect 3637 1456 3704 1460
rect 3610 1453 3704 1456
rect 3610 1446 3659 1453
rect 3610 1440 3640 1446
rect 3659 1441 3664 1446
rect 3576 1424 3656 1440
rect 3668 1432 3704 1453
rect 3765 1448 3954 1472
rect 3999 1471 4046 1472
rect 4012 1466 4046 1471
rect 4086 1466 4102 1468
rect 3780 1445 3954 1448
rect 3773 1442 3954 1445
rect 3982 1465 4046 1466
rect 3576 1422 3595 1424
rect 3610 1422 3644 1424
rect 3576 1406 3656 1422
rect 3576 1400 3595 1406
rect 3292 1374 3395 1384
rect 3246 1372 3395 1374
rect 3416 1372 3451 1384
rect 3085 1370 3247 1372
rect 3097 1352 3116 1370
rect 3131 1368 3161 1370
rect 2980 1342 3021 1350
rect 3104 1346 3116 1352
rect 3168 1354 3247 1370
rect 3279 1370 3451 1372
rect 3279 1354 3358 1370
rect 3365 1368 3395 1370
rect 2943 1332 2972 1342
rect 2986 1332 3015 1342
rect 3030 1332 3060 1346
rect 3104 1332 3146 1346
rect 3168 1342 3358 1354
rect 3423 1350 3429 1370
rect 3153 1332 3183 1342
rect 3184 1332 3342 1342
rect 3346 1332 3376 1342
rect 3380 1332 3410 1346
rect 3438 1332 3451 1370
rect 3523 1384 3552 1400
rect 3566 1384 3595 1400
rect 3610 1390 3640 1406
rect 3668 1384 3674 1432
rect 3677 1426 3696 1432
rect 3711 1426 3741 1434
rect 3677 1418 3741 1426
rect 3677 1402 3757 1418
rect 3773 1411 3835 1442
rect 3851 1411 3913 1442
rect 3982 1440 4031 1465
rect 4076 1456 4102 1466
rect 4046 1440 4102 1456
rect 3945 1426 3975 1434
rect 3982 1432 4092 1440
rect 3945 1418 3990 1426
rect 3677 1400 3696 1402
rect 3711 1400 3757 1402
rect 3677 1384 3757 1400
rect 3784 1398 3819 1411
rect 3860 1408 3897 1411
rect 3860 1406 3902 1408
rect 3789 1395 3819 1398
rect 3798 1391 3805 1395
rect 3805 1390 3806 1391
rect 3764 1384 3774 1390
rect 3523 1376 3558 1384
rect 3523 1350 3524 1376
rect 3531 1350 3558 1376
rect 3466 1332 3496 1346
rect 3523 1342 3558 1350
rect 3560 1376 3601 1384
rect 3560 1350 3575 1376
rect 3582 1350 3601 1376
rect 3665 1372 3696 1384
rect 3711 1372 3814 1384
rect 3826 1374 3852 1400
rect 3867 1395 3897 1406
rect 3929 1402 3991 1418
rect 3929 1400 3975 1402
rect 3929 1384 3991 1400
rect 4003 1384 4009 1432
rect 4012 1424 4092 1432
rect 4012 1422 4031 1424
rect 4046 1422 4080 1424
rect 4012 1406 4092 1422
rect 4012 1384 4031 1406
rect 4046 1390 4076 1406
rect 4104 1400 4110 1474
rect 4113 1400 4132 1544
rect 4147 1400 4153 1544
rect 4162 1474 4175 1544
rect 4227 1540 4249 1544
rect 4220 1528 4237 1532
rect 4241 1530 4249 1532
rect 4239 1528 4249 1530
rect 4220 1518 4249 1528
rect 4302 1518 4318 1532
rect 4356 1528 4362 1530
rect 4369 1528 4477 1544
rect 4484 1528 4490 1530
rect 4498 1528 4513 1544
rect 4579 1538 4598 1541
rect 4220 1516 4318 1518
rect 4345 1516 4513 1528
rect 4528 1518 4544 1532
rect 4579 1519 4601 1538
rect 4611 1532 4627 1533
rect 4610 1530 4627 1532
rect 4611 1525 4627 1530
rect 4601 1518 4607 1519
rect 4610 1518 4639 1525
rect 4528 1517 4639 1518
rect 4528 1516 4645 1517
rect 4204 1508 4255 1516
rect 4302 1508 4336 1516
rect 4204 1496 4229 1508
rect 4236 1496 4255 1508
rect 4309 1506 4336 1508
rect 4345 1506 4566 1516
rect 4601 1513 4607 1516
rect 4309 1502 4566 1506
rect 4204 1488 4255 1496
rect 4302 1488 4566 1502
rect 4610 1508 4645 1516
rect 4156 1440 4175 1474
rect 4220 1480 4249 1488
rect 4220 1474 4237 1480
rect 4220 1472 4254 1474
rect 4302 1472 4318 1488
rect 4319 1478 4527 1488
rect 4528 1478 4544 1488
rect 4592 1484 4607 1499
rect 4610 1496 4611 1508
rect 4618 1496 4645 1508
rect 4610 1488 4645 1496
rect 4610 1487 4639 1488
rect 4330 1474 4544 1478
rect 4345 1472 4544 1474
rect 4579 1474 4592 1484
rect 4610 1474 4627 1487
rect 4579 1472 4627 1474
rect 4221 1468 4254 1472
rect 4217 1466 4254 1468
rect 4217 1465 4284 1466
rect 4217 1460 4248 1465
rect 4254 1460 4284 1465
rect 4217 1456 4284 1460
rect 4190 1453 4284 1456
rect 4190 1446 4239 1453
rect 4190 1440 4220 1446
rect 4239 1441 4244 1446
rect 4156 1424 4236 1440
rect 4248 1432 4284 1453
rect 4345 1448 4534 1472
rect 4579 1471 4626 1472
rect 4592 1466 4626 1471
rect 4360 1445 4534 1448
rect 4353 1442 4534 1445
rect 4562 1465 4626 1466
rect 4156 1422 4175 1424
rect 4190 1422 4224 1424
rect 4156 1406 4236 1422
rect 4156 1400 4175 1406
rect 3872 1374 3975 1384
rect 3826 1372 3975 1374
rect 3996 1372 4031 1384
rect 3665 1370 3827 1372
rect 3677 1352 3696 1370
rect 3711 1368 3741 1370
rect 3560 1342 3601 1350
rect 3684 1346 3696 1352
rect 3748 1354 3827 1370
rect 3859 1370 4031 1372
rect 3859 1354 3938 1370
rect 3945 1368 3975 1370
rect 3523 1332 3552 1342
rect 3566 1332 3595 1342
rect 3610 1332 3640 1346
rect 3684 1332 3726 1346
rect 3748 1342 3938 1354
rect 4003 1350 4009 1370
rect 3733 1332 3763 1342
rect 3764 1332 3922 1342
rect 3926 1332 3956 1342
rect 3960 1332 3990 1346
rect 4018 1332 4031 1370
rect 4103 1384 4132 1400
rect 4146 1384 4175 1400
rect 4190 1390 4220 1406
rect 4248 1384 4254 1432
rect 4257 1426 4276 1432
rect 4291 1426 4321 1434
rect 4257 1418 4321 1426
rect 4257 1402 4337 1418
rect 4353 1411 4415 1442
rect 4431 1411 4493 1442
rect 4562 1440 4611 1465
rect 4626 1440 4656 1458
rect 4525 1426 4555 1434
rect 4562 1432 4672 1440
rect 4525 1418 4570 1426
rect 4257 1400 4276 1402
rect 4291 1400 4337 1402
rect 4257 1384 4337 1400
rect 4364 1398 4399 1411
rect 4440 1408 4477 1411
rect 4440 1406 4482 1408
rect 4369 1395 4399 1398
rect 4378 1391 4385 1395
rect 4385 1390 4386 1391
rect 4344 1384 4354 1390
rect 4103 1376 4138 1384
rect 4103 1350 4104 1376
rect 4111 1350 4138 1376
rect 4046 1332 4076 1346
rect 4103 1342 4138 1350
rect 4140 1376 4181 1384
rect 4140 1350 4155 1376
rect 4162 1350 4181 1376
rect 4245 1372 4276 1384
rect 4291 1372 4394 1384
rect 4406 1374 4432 1400
rect 4447 1395 4477 1406
rect 4509 1402 4571 1418
rect 4509 1400 4555 1402
rect 4509 1384 4571 1400
rect 4583 1384 4589 1432
rect 4592 1424 4672 1432
rect 4592 1422 4611 1424
rect 4626 1422 4660 1424
rect 4592 1407 4672 1422
rect 4592 1406 4678 1407
rect 4592 1384 4611 1406
rect 4626 1390 4656 1406
rect 4684 1400 4690 1474
rect 4693 1400 4712 1544
rect 4727 1400 4733 1544
rect 4742 1474 4755 1544
rect 4807 1540 4829 1544
rect 4800 1528 4817 1532
rect 4821 1530 4829 1532
rect 4819 1528 4829 1530
rect 4800 1518 4829 1528
rect 4882 1518 4898 1532
rect 4936 1528 4942 1530
rect 4949 1528 5057 1544
rect 5064 1528 5070 1530
rect 5078 1528 5093 1544
rect 5159 1538 5178 1541
rect 4800 1516 4898 1518
rect 4925 1516 5093 1528
rect 5108 1518 5124 1532
rect 5159 1519 5181 1538
rect 5191 1532 5207 1533
rect 5190 1530 5207 1532
rect 5191 1525 5207 1530
rect 5181 1518 5187 1519
rect 5190 1518 5219 1525
rect 5108 1517 5219 1518
rect 5108 1516 5225 1517
rect 4784 1508 4835 1516
rect 4882 1508 4916 1516
rect 4784 1496 4809 1508
rect 4816 1496 4835 1508
rect 4889 1506 4916 1508
rect 4925 1506 5146 1516
rect 5181 1513 5187 1516
rect 4889 1502 5146 1506
rect 4784 1488 4835 1496
rect 4882 1488 5146 1502
rect 5190 1508 5225 1516
rect 4736 1440 4755 1474
rect 4800 1480 4829 1488
rect 4800 1474 4817 1480
rect 4800 1472 4834 1474
rect 4882 1472 4898 1488
rect 4899 1478 5107 1488
rect 5108 1478 5124 1488
rect 5172 1484 5187 1499
rect 5190 1496 5191 1508
rect 5198 1496 5225 1508
rect 5190 1488 5225 1496
rect 5190 1487 5219 1488
rect 4910 1474 5124 1478
rect 4925 1472 5124 1474
rect 5159 1474 5172 1484
rect 5190 1474 5207 1487
rect 5159 1472 5207 1474
rect 4801 1468 4834 1472
rect 4797 1466 4834 1468
rect 4797 1465 4864 1466
rect 4797 1460 4828 1465
rect 4834 1460 4864 1465
rect 4797 1456 4864 1460
rect 4770 1453 4864 1456
rect 4770 1446 4819 1453
rect 4770 1440 4800 1446
rect 4819 1441 4824 1446
rect 4736 1424 4816 1440
rect 4828 1432 4864 1453
rect 4925 1448 5114 1472
rect 5159 1471 5206 1472
rect 5172 1466 5206 1471
rect 5246 1466 5262 1468
rect 4940 1445 5114 1448
rect 4933 1442 5114 1445
rect 5142 1465 5206 1466
rect 4736 1422 4755 1424
rect 4770 1422 4804 1424
rect 4736 1406 4816 1422
rect 4736 1400 4755 1406
rect 4452 1374 4555 1384
rect 4406 1372 4555 1374
rect 4576 1372 4611 1384
rect 4245 1370 4407 1372
rect 4257 1352 4276 1370
rect 4291 1368 4321 1370
rect 4140 1342 4181 1350
rect 4264 1346 4276 1352
rect 4328 1354 4407 1370
rect 4439 1370 4611 1372
rect 4439 1354 4518 1370
rect 4525 1368 4555 1370
rect 4103 1332 4132 1342
rect 4146 1332 4175 1342
rect 4190 1332 4220 1346
rect 4264 1332 4306 1346
rect 4328 1342 4518 1354
rect 4583 1350 4589 1370
rect 4313 1332 4343 1342
rect 4344 1332 4502 1342
rect 4506 1332 4536 1342
rect 4540 1332 4570 1346
rect 4598 1332 4611 1370
rect 4683 1384 4712 1400
rect 4726 1384 4755 1400
rect 4770 1390 4800 1406
rect 4828 1384 4834 1432
rect 4837 1426 4856 1432
rect 4871 1426 4901 1434
rect 4837 1418 4901 1426
rect 4837 1402 4917 1418
rect 4933 1411 4995 1442
rect 5011 1411 5073 1442
rect 5142 1440 5191 1465
rect 5236 1456 5262 1466
rect 5206 1440 5262 1456
rect 5105 1426 5135 1434
rect 5142 1432 5252 1440
rect 5105 1418 5150 1426
rect 4837 1400 4856 1402
rect 4871 1400 4917 1402
rect 4837 1384 4917 1400
rect 4944 1398 4979 1411
rect 5020 1408 5057 1411
rect 5020 1406 5062 1408
rect 4949 1395 4979 1398
rect 4958 1391 4965 1395
rect 4965 1390 4966 1391
rect 4924 1384 4934 1390
rect 4683 1376 4718 1384
rect 4683 1350 4684 1376
rect 4691 1350 4718 1376
rect 4626 1332 4656 1346
rect 4683 1342 4718 1350
rect 4720 1376 4761 1384
rect 4720 1350 4735 1376
rect 4742 1350 4761 1376
rect 4825 1372 4856 1384
rect 4871 1372 4974 1384
rect 4986 1374 5012 1400
rect 5027 1395 5057 1406
rect 5089 1402 5151 1418
rect 5089 1400 5135 1402
rect 5089 1384 5151 1400
rect 5163 1384 5169 1432
rect 5172 1424 5252 1432
rect 5172 1422 5191 1424
rect 5206 1422 5240 1424
rect 5172 1406 5252 1422
rect 5172 1384 5191 1406
rect 5206 1390 5236 1406
rect 5264 1400 5270 1474
rect 5273 1400 5292 1544
rect 5307 1400 5313 1544
rect 5322 1474 5335 1544
rect 5387 1540 5409 1544
rect 5380 1528 5397 1532
rect 5401 1530 5409 1532
rect 5399 1528 5409 1530
rect 5380 1518 5409 1528
rect 5462 1518 5478 1532
rect 5516 1528 5522 1530
rect 5529 1528 5637 1544
rect 5644 1528 5650 1530
rect 5658 1528 5673 1544
rect 5739 1538 5758 1541
rect 5380 1516 5478 1518
rect 5505 1516 5673 1528
rect 5688 1518 5704 1532
rect 5739 1519 5761 1538
rect 5771 1532 5787 1533
rect 5770 1530 5787 1532
rect 5771 1525 5787 1530
rect 5761 1518 5767 1519
rect 5770 1518 5799 1525
rect 5688 1517 5799 1518
rect 5688 1516 5805 1517
rect 5364 1508 5415 1516
rect 5462 1508 5496 1516
rect 5364 1496 5389 1508
rect 5396 1496 5415 1508
rect 5469 1506 5496 1508
rect 5505 1506 5726 1516
rect 5761 1513 5767 1516
rect 5469 1502 5726 1506
rect 5364 1488 5415 1496
rect 5462 1488 5726 1502
rect 5770 1508 5805 1516
rect 5316 1440 5335 1474
rect 5380 1480 5409 1488
rect 5380 1474 5397 1480
rect 5380 1472 5414 1474
rect 5462 1472 5478 1488
rect 5479 1478 5687 1488
rect 5688 1478 5704 1488
rect 5752 1484 5767 1499
rect 5770 1496 5771 1508
rect 5778 1496 5805 1508
rect 5770 1488 5805 1496
rect 5770 1487 5799 1488
rect 5490 1474 5704 1478
rect 5505 1472 5704 1474
rect 5739 1474 5752 1484
rect 5770 1474 5787 1487
rect 5739 1472 5787 1474
rect 5381 1468 5414 1472
rect 5377 1466 5414 1468
rect 5377 1465 5444 1466
rect 5377 1460 5408 1465
rect 5414 1460 5444 1465
rect 5377 1456 5444 1460
rect 5350 1453 5444 1456
rect 5350 1446 5399 1453
rect 5350 1440 5380 1446
rect 5399 1441 5404 1446
rect 5316 1424 5396 1440
rect 5408 1432 5444 1453
rect 5505 1448 5694 1472
rect 5739 1471 5786 1472
rect 5752 1466 5786 1471
rect 5520 1445 5694 1448
rect 5513 1442 5694 1445
rect 5722 1465 5786 1466
rect 5316 1422 5335 1424
rect 5350 1422 5384 1424
rect 5316 1406 5396 1422
rect 5316 1400 5335 1406
rect 5032 1374 5135 1384
rect 4986 1372 5135 1374
rect 5156 1372 5191 1384
rect 4825 1370 4987 1372
rect 4837 1352 4856 1370
rect 4871 1368 4901 1370
rect 4720 1342 4761 1350
rect 4844 1346 4856 1352
rect 4908 1354 4987 1370
rect 5019 1370 5191 1372
rect 5019 1354 5098 1370
rect 5105 1368 5135 1370
rect 4683 1332 4712 1342
rect 4726 1332 4755 1342
rect 4770 1332 4800 1346
rect 4844 1332 4886 1346
rect 4908 1342 5098 1354
rect 5163 1350 5169 1370
rect 4893 1332 4923 1342
rect 4924 1332 5082 1342
rect 5086 1332 5116 1342
rect 5120 1332 5150 1346
rect 5178 1332 5191 1370
rect 5263 1384 5292 1400
rect 5306 1384 5335 1400
rect 5350 1390 5380 1406
rect 5408 1384 5414 1432
rect 5417 1426 5436 1432
rect 5451 1426 5481 1434
rect 5417 1418 5481 1426
rect 5417 1402 5497 1418
rect 5513 1411 5575 1442
rect 5591 1411 5653 1442
rect 5722 1440 5771 1465
rect 5786 1440 5816 1458
rect 5685 1426 5715 1434
rect 5722 1432 5832 1440
rect 5685 1418 5730 1426
rect 5417 1400 5436 1402
rect 5451 1400 5497 1402
rect 5417 1384 5497 1400
rect 5524 1398 5559 1411
rect 5600 1408 5637 1411
rect 5600 1406 5642 1408
rect 5529 1395 5559 1398
rect 5538 1391 5545 1395
rect 5545 1390 5546 1391
rect 5504 1384 5514 1390
rect 5263 1376 5298 1384
rect 5263 1350 5264 1376
rect 5271 1350 5298 1376
rect 5206 1332 5236 1346
rect 5263 1342 5298 1350
rect 5300 1376 5341 1384
rect 5300 1350 5315 1376
rect 5322 1350 5341 1376
rect 5405 1372 5436 1384
rect 5451 1372 5554 1384
rect 5566 1374 5592 1400
rect 5607 1395 5637 1406
rect 5669 1402 5731 1418
rect 5669 1400 5715 1402
rect 5669 1384 5731 1400
rect 5743 1384 5749 1432
rect 5752 1424 5832 1432
rect 5752 1422 5771 1424
rect 5786 1422 5820 1424
rect 5752 1407 5832 1422
rect 5752 1406 5838 1407
rect 5752 1384 5771 1406
rect 5786 1390 5816 1406
rect 5844 1400 5850 1474
rect 5853 1400 5872 1544
rect 5887 1400 5893 1544
rect 5902 1474 5915 1544
rect 5967 1540 5989 1544
rect 5960 1528 5977 1532
rect 5981 1530 5989 1532
rect 5979 1528 5989 1530
rect 5960 1518 5989 1528
rect 6042 1518 6058 1532
rect 6096 1528 6102 1530
rect 6109 1528 6217 1544
rect 6224 1528 6230 1530
rect 6238 1528 6253 1544
rect 6319 1538 6338 1541
rect 5960 1516 6058 1518
rect 6085 1516 6253 1528
rect 6268 1518 6284 1532
rect 6319 1519 6341 1538
rect 6351 1532 6367 1533
rect 6350 1530 6367 1532
rect 6351 1525 6367 1530
rect 6341 1518 6347 1519
rect 6350 1518 6379 1525
rect 6268 1517 6379 1518
rect 6268 1516 6385 1517
rect 5944 1508 5995 1516
rect 6042 1508 6076 1516
rect 5944 1496 5969 1508
rect 5976 1496 5995 1508
rect 6049 1506 6076 1508
rect 6085 1506 6306 1516
rect 6341 1513 6347 1516
rect 6049 1502 6306 1506
rect 5944 1488 5995 1496
rect 6042 1488 6306 1502
rect 6350 1508 6385 1516
rect 5896 1440 5915 1474
rect 5960 1480 5989 1488
rect 5960 1474 5977 1480
rect 5960 1472 5994 1474
rect 6042 1472 6058 1488
rect 6059 1478 6267 1488
rect 6268 1478 6284 1488
rect 6332 1484 6347 1499
rect 6350 1496 6351 1508
rect 6358 1496 6385 1508
rect 6350 1488 6385 1496
rect 6350 1487 6379 1488
rect 6070 1474 6284 1478
rect 6085 1472 6284 1474
rect 6319 1474 6332 1484
rect 6350 1474 6367 1487
rect 6319 1472 6367 1474
rect 5961 1468 5994 1472
rect 5957 1466 5994 1468
rect 5957 1465 6024 1466
rect 5957 1460 5988 1465
rect 5994 1460 6024 1465
rect 5957 1456 6024 1460
rect 5930 1453 6024 1456
rect 5930 1446 5979 1453
rect 5930 1440 5960 1446
rect 5979 1441 5984 1446
rect 5896 1424 5976 1440
rect 5988 1432 6024 1453
rect 6085 1448 6274 1472
rect 6319 1471 6366 1472
rect 6332 1466 6366 1471
rect 6100 1445 6274 1448
rect 6093 1442 6274 1445
rect 6302 1465 6366 1466
rect 5896 1422 5915 1424
rect 5930 1422 5964 1424
rect 5896 1406 5976 1422
rect 5896 1400 5915 1406
rect 5612 1374 5715 1384
rect 5566 1372 5715 1374
rect 5736 1372 5771 1384
rect 5405 1370 5567 1372
rect 5417 1352 5436 1370
rect 5451 1368 5481 1370
rect 5300 1342 5341 1350
rect 5424 1346 5436 1352
rect 5488 1354 5567 1370
rect 5599 1370 5771 1372
rect 5599 1354 5678 1370
rect 5685 1368 5715 1370
rect 5263 1332 5292 1342
rect 5306 1332 5335 1342
rect 5350 1332 5380 1346
rect 5424 1332 5466 1346
rect 5488 1342 5678 1354
rect 5743 1350 5749 1370
rect 5473 1332 5503 1342
rect 5504 1332 5662 1342
rect 5666 1332 5696 1342
rect 5700 1332 5730 1346
rect 5758 1332 5771 1370
rect 5843 1384 5872 1400
rect 5886 1384 5915 1400
rect 5930 1390 5960 1406
rect 5988 1384 5994 1432
rect 5997 1426 6016 1432
rect 6031 1426 6061 1434
rect 5997 1418 6061 1426
rect 5997 1402 6077 1418
rect 6093 1411 6155 1442
rect 6171 1411 6233 1442
rect 6302 1440 6351 1465
rect 6366 1440 6396 1456
rect 6265 1426 6295 1434
rect 6302 1432 6412 1440
rect 6265 1418 6310 1426
rect 5997 1400 6016 1402
rect 6031 1400 6077 1402
rect 5997 1384 6077 1400
rect 6104 1398 6139 1411
rect 6180 1408 6217 1411
rect 6180 1406 6222 1408
rect 6109 1395 6139 1398
rect 6118 1391 6125 1395
rect 6125 1390 6126 1391
rect 6084 1384 6094 1390
rect 5843 1376 5878 1384
rect 5843 1350 5844 1376
rect 5851 1350 5878 1376
rect 5786 1332 5816 1346
rect 5843 1342 5878 1350
rect 5880 1376 5921 1384
rect 5880 1350 5895 1376
rect 5902 1350 5921 1376
rect 5985 1372 6016 1384
rect 6031 1372 6134 1384
rect 6146 1374 6172 1400
rect 6187 1395 6217 1406
rect 6249 1402 6311 1418
rect 6249 1400 6295 1402
rect 6249 1384 6311 1400
rect 6323 1384 6329 1432
rect 6332 1424 6412 1432
rect 6332 1422 6351 1424
rect 6366 1422 6400 1424
rect 6332 1406 6412 1422
rect 6332 1384 6351 1406
rect 6366 1390 6396 1406
rect 6424 1400 6430 1474
rect 6439 1400 6452 1544
rect 6192 1374 6295 1384
rect 6146 1372 6295 1374
rect 6316 1372 6351 1384
rect 5985 1370 6147 1372
rect 5997 1352 6016 1370
rect 6031 1368 6061 1370
rect 5880 1342 5921 1350
rect 6004 1346 6016 1352
rect 6068 1354 6147 1370
rect 6179 1370 6351 1372
rect 6179 1354 6258 1370
rect 6265 1368 6295 1370
rect 5843 1332 5872 1342
rect 5886 1332 5915 1342
rect 5930 1332 5960 1346
rect 6004 1332 6046 1346
rect 6068 1342 6258 1354
rect 6323 1350 6329 1370
rect 6053 1332 6083 1342
rect 6084 1332 6242 1342
rect 6246 1332 6276 1342
rect 6280 1332 6310 1346
rect 6338 1332 6351 1370
rect 6423 1384 6452 1400
rect 6423 1376 6458 1384
rect 6423 1350 6424 1376
rect 6431 1350 6458 1376
rect 6366 1332 6396 1346
rect 6423 1342 6458 1350
rect 6423 1332 6452 1342
rect -541 1318 6452 1332
rect -478 1288 -465 1318
rect -450 1304 -420 1318
rect -376 1304 -334 1318
rect -327 1304 -107 1318
rect -100 1304 -70 1318
rect -410 1290 -395 1302
rect -376 1290 -363 1304
rect -295 1300 -142 1304
rect -413 1288 -391 1290
rect -313 1288 -121 1300
rect -42 1288 -29 1318
rect -14 1304 16 1318
rect 53 1288 72 1318
rect 87 1288 93 1318
rect 102 1288 115 1318
rect 130 1304 160 1318
rect 204 1304 246 1318
rect 253 1304 473 1318
rect 480 1304 510 1318
rect 170 1290 185 1302
rect 204 1290 217 1304
rect 285 1300 438 1304
rect 167 1288 189 1290
rect 267 1288 459 1300
rect 538 1288 551 1318
rect 566 1304 596 1318
rect 633 1288 652 1318
rect 667 1288 673 1318
rect 682 1288 695 1318
rect 710 1304 740 1318
rect 784 1304 826 1318
rect 833 1304 1053 1318
rect 1060 1304 1090 1318
rect 750 1290 765 1302
rect 784 1290 797 1304
rect 865 1300 1018 1304
rect 747 1288 769 1290
rect 847 1288 1039 1300
rect 1118 1288 1131 1318
rect 1146 1304 1176 1318
rect 1213 1288 1232 1318
rect 1247 1288 1253 1318
rect 1262 1288 1275 1318
rect 1290 1304 1320 1318
rect 1364 1304 1406 1318
rect 1413 1304 1633 1318
rect 1640 1304 1670 1318
rect 1330 1290 1345 1302
rect 1364 1290 1377 1304
rect 1445 1300 1598 1304
rect 1327 1288 1349 1290
rect 1427 1288 1619 1300
rect 1698 1288 1711 1318
rect 1726 1304 1756 1318
rect 1793 1288 1812 1318
rect 1827 1288 1833 1318
rect 1842 1288 1855 1318
rect 1870 1304 1900 1318
rect 1944 1304 1986 1318
rect 1993 1304 2213 1318
rect 2220 1304 2250 1318
rect 1910 1290 1925 1302
rect 1944 1290 1957 1304
rect 2025 1300 2178 1304
rect 1907 1288 1929 1290
rect 2007 1288 2199 1300
rect 2278 1288 2291 1318
rect 2306 1304 2336 1318
rect 2373 1288 2392 1318
rect 2407 1288 2413 1318
rect 2422 1288 2435 1318
rect 2450 1304 2480 1318
rect 2524 1304 2566 1318
rect 2573 1304 2793 1318
rect 2800 1304 2830 1318
rect 2490 1290 2505 1302
rect 2524 1290 2537 1304
rect 2605 1300 2758 1304
rect 2487 1288 2509 1290
rect 2587 1288 2779 1300
rect 2858 1288 2871 1318
rect 2886 1304 2916 1318
rect 2953 1288 2972 1318
rect 2987 1288 2993 1318
rect 3002 1288 3015 1318
rect 3030 1304 3060 1318
rect 3104 1304 3146 1318
rect 3153 1304 3373 1318
rect 3380 1304 3410 1318
rect 3070 1290 3085 1302
rect 3104 1290 3117 1304
rect 3185 1300 3338 1304
rect 3067 1288 3089 1290
rect 3167 1288 3359 1300
rect 3438 1288 3451 1318
rect 3466 1304 3496 1318
rect 3533 1288 3552 1318
rect 3567 1288 3573 1318
rect 3582 1288 3595 1318
rect 3610 1304 3640 1318
rect 3684 1304 3726 1318
rect 3733 1304 3953 1318
rect 3960 1304 3990 1318
rect 3650 1290 3665 1302
rect 3684 1290 3697 1304
rect 3765 1300 3918 1304
rect 3647 1288 3669 1290
rect 3747 1288 3939 1300
rect 4018 1288 4031 1318
rect 4046 1304 4076 1318
rect 4113 1288 4132 1318
rect 4147 1288 4153 1318
rect 4162 1288 4175 1318
rect 4190 1304 4220 1318
rect 4264 1304 4306 1318
rect 4313 1304 4533 1318
rect 4540 1304 4570 1318
rect 4230 1290 4245 1302
rect 4264 1290 4277 1304
rect 4345 1300 4498 1304
rect 4227 1288 4249 1290
rect 4327 1288 4519 1300
rect 4598 1288 4611 1318
rect 4626 1304 4656 1318
rect 4693 1288 4712 1318
rect 4727 1288 4733 1318
rect 4742 1288 4755 1318
rect 4770 1304 4800 1318
rect 4844 1304 4886 1318
rect 4893 1304 5113 1318
rect 5120 1304 5150 1318
rect 4810 1290 4825 1302
rect 4844 1290 4857 1304
rect 4925 1300 5078 1304
rect 4807 1288 4829 1290
rect 4907 1288 5099 1300
rect 5178 1288 5191 1318
rect 5206 1304 5236 1318
rect 5273 1288 5292 1318
rect 5307 1288 5313 1318
rect 5322 1288 5335 1318
rect 5350 1304 5380 1318
rect 5424 1304 5466 1318
rect 5473 1304 5693 1318
rect 5700 1304 5730 1318
rect 5390 1290 5405 1302
rect 5424 1290 5437 1304
rect 5505 1300 5658 1304
rect 5387 1288 5409 1290
rect 5487 1288 5679 1300
rect 5758 1288 5771 1318
rect 5786 1304 5816 1318
rect 5853 1288 5872 1318
rect 5887 1288 5893 1318
rect 5902 1288 5915 1318
rect 5930 1304 5960 1318
rect 6004 1304 6046 1318
rect 6053 1304 6273 1318
rect 6280 1304 6310 1318
rect 5970 1290 5985 1302
rect 6004 1290 6017 1304
rect 6085 1300 6238 1304
rect 5967 1288 5989 1290
rect 6067 1288 6259 1300
rect 6338 1288 6351 1318
rect 6366 1304 6396 1318
rect 6439 1288 6452 1318
rect -541 1274 6452 1288
rect -478 1204 -465 1274
rect -413 1270 -391 1274
rect -420 1258 -403 1262
rect -399 1260 -391 1262
rect -401 1258 -391 1260
rect -420 1248 -391 1258
rect -338 1248 -322 1262
rect -284 1258 -278 1260
rect -271 1258 -163 1274
rect -156 1258 -150 1260
rect -142 1258 -127 1274
rect -61 1268 -42 1271
rect -420 1246 -322 1248
rect -295 1246 -127 1258
rect -112 1248 -96 1262
rect -61 1249 -39 1268
rect -29 1262 -13 1263
rect -30 1260 -13 1262
rect -29 1255 -13 1260
rect -39 1248 -33 1249
rect -30 1248 -1 1255
rect -112 1247 -1 1248
rect -112 1246 5 1247
rect -436 1238 -385 1246
rect -338 1238 -304 1246
rect -436 1226 -411 1238
rect -404 1226 -385 1238
rect -331 1236 -304 1238
rect -295 1236 -74 1246
rect -39 1243 -33 1246
rect -331 1232 -74 1236
rect -436 1218 -385 1226
rect -338 1218 -74 1232
rect -30 1238 5 1246
rect -484 1170 -465 1204
rect -420 1210 -391 1218
rect -420 1204 -403 1210
rect -420 1202 -386 1204
rect -338 1202 -322 1218
rect -321 1208 -113 1218
rect -112 1208 -96 1218
rect -48 1214 -33 1229
rect -30 1226 -29 1238
rect -22 1226 5 1238
rect -30 1218 5 1226
rect -30 1217 -1 1218
rect -310 1204 -96 1208
rect -295 1202 -96 1204
rect -61 1204 -48 1214
rect -30 1204 -13 1217
rect -61 1202 -13 1204
rect -419 1198 -386 1202
rect -423 1196 -386 1198
rect -423 1195 -356 1196
rect -423 1190 -392 1195
rect -386 1190 -356 1195
rect -423 1186 -356 1190
rect -450 1183 -356 1186
rect -450 1176 -401 1183
rect -450 1170 -420 1176
rect -401 1171 -396 1176
rect -484 1154 -404 1170
rect -392 1162 -356 1183
rect -295 1178 -106 1202
rect -61 1201 -14 1202
rect -48 1196 -14 1201
rect -280 1175 -106 1178
rect -287 1172 -106 1175
rect -78 1195 -14 1196
rect -484 1152 -465 1154
rect -450 1152 -416 1154
rect -484 1136 -404 1152
rect -484 1130 -465 1136
rect -494 1114 -465 1130
rect -450 1120 -420 1136
rect -392 1114 -386 1162
rect -383 1156 -364 1162
rect -349 1156 -319 1164
rect -383 1148 -319 1156
rect -383 1132 -303 1148
rect -287 1141 -225 1172
rect -209 1141 -147 1172
rect -78 1170 -29 1195
rect -14 1170 16 1188
rect -115 1156 -85 1164
rect -78 1162 32 1170
rect -115 1148 -70 1156
rect -383 1130 -364 1132
rect -349 1130 -303 1132
rect -383 1114 -303 1130
rect -276 1128 -241 1141
rect -200 1138 -163 1141
rect -200 1136 -158 1138
rect -271 1125 -241 1128
rect -262 1121 -255 1125
rect -255 1120 -254 1121
rect -296 1114 -286 1120
rect -500 1106 -459 1114
rect -500 1080 -485 1106
rect -478 1080 -459 1106
rect -395 1102 -364 1114
rect -349 1102 -246 1114
rect -234 1104 -208 1130
rect -193 1125 -163 1136
rect -131 1132 -69 1148
rect -131 1130 -85 1132
rect -131 1114 -69 1130
rect -57 1114 -51 1162
rect -48 1154 32 1162
rect -48 1152 -29 1154
rect -14 1152 20 1154
rect -48 1137 32 1152
rect -48 1136 38 1137
rect -48 1114 -29 1136
rect -14 1120 16 1136
rect 44 1130 50 1204
rect 53 1130 72 1274
rect 87 1130 93 1274
rect 102 1204 115 1274
rect 167 1270 189 1274
rect 160 1258 177 1262
rect 181 1260 189 1262
rect 179 1258 189 1260
rect 160 1248 189 1258
rect 242 1248 258 1262
rect 296 1258 302 1260
rect 309 1258 417 1274
rect 424 1258 430 1260
rect 438 1258 453 1274
rect 519 1268 538 1271
rect 160 1246 258 1248
rect 285 1246 453 1258
rect 468 1248 484 1262
rect 519 1249 541 1268
rect 551 1262 567 1263
rect 550 1260 567 1262
rect 551 1255 567 1260
rect 541 1248 547 1249
rect 550 1248 579 1255
rect 468 1247 579 1248
rect 468 1246 585 1247
rect 144 1238 195 1246
rect 242 1238 276 1246
rect 144 1226 169 1238
rect 176 1226 195 1238
rect 249 1236 276 1238
rect 285 1236 506 1246
rect 541 1243 547 1246
rect 249 1232 506 1236
rect 144 1218 195 1226
rect 242 1218 506 1232
rect 550 1238 585 1246
rect 96 1170 115 1204
rect 160 1210 189 1218
rect 160 1204 177 1210
rect 160 1202 194 1204
rect 242 1202 258 1218
rect 259 1208 467 1218
rect 468 1208 484 1218
rect 532 1214 547 1229
rect 550 1226 551 1238
rect 558 1226 585 1238
rect 550 1218 585 1226
rect 550 1217 579 1218
rect 270 1204 484 1208
rect 285 1202 484 1204
rect 519 1204 532 1214
rect 550 1204 567 1217
rect 519 1202 567 1204
rect 161 1198 194 1202
rect 157 1196 194 1198
rect 157 1195 224 1196
rect 157 1190 188 1195
rect 194 1190 224 1195
rect 157 1186 224 1190
rect 130 1183 224 1186
rect 130 1176 179 1183
rect 130 1170 160 1176
rect 179 1171 184 1176
rect 96 1154 176 1170
rect 188 1162 224 1183
rect 285 1178 474 1202
rect 519 1201 566 1202
rect 532 1196 566 1201
rect 606 1196 622 1198
rect 300 1175 474 1178
rect 293 1172 474 1175
rect 502 1195 566 1196
rect 96 1152 115 1154
rect 130 1152 164 1154
rect 96 1136 176 1152
rect 96 1130 115 1136
rect -188 1104 -85 1114
rect -234 1102 -85 1104
rect -64 1102 -29 1114
rect -395 1100 -233 1102
rect -383 1080 -364 1100
rect -349 1098 -319 1100
rect -500 1072 -459 1080
rect -377 1076 -364 1080
rect -312 1084 -233 1100
rect -201 1100 -29 1102
rect -201 1084 -122 1100
rect -115 1098 -85 1100
rect -494 1062 -465 1072
rect -450 1062 -420 1076
rect -377 1062 -334 1076
rect -312 1072 -122 1084
rect -57 1080 -51 1100
rect -327 1062 -297 1072
rect -296 1062 -138 1072
rect -134 1062 -104 1072
rect -100 1062 -70 1076
rect -42 1062 -29 1100
rect 43 1114 72 1130
rect 86 1114 115 1130
rect 130 1120 160 1136
rect 188 1114 194 1162
rect 197 1156 216 1162
rect 231 1156 261 1164
rect 197 1148 261 1156
rect 197 1132 277 1148
rect 293 1141 355 1172
rect 371 1141 433 1172
rect 502 1170 551 1195
rect 596 1186 622 1196
rect 566 1170 622 1186
rect 465 1156 495 1164
rect 502 1162 612 1170
rect 465 1148 510 1156
rect 197 1130 216 1132
rect 231 1130 277 1132
rect 197 1114 277 1130
rect 304 1128 339 1141
rect 380 1138 417 1141
rect 380 1136 422 1138
rect 309 1125 339 1128
rect 318 1121 325 1125
rect 325 1120 326 1121
rect 284 1114 294 1120
rect 43 1106 78 1114
rect 43 1080 44 1106
rect 51 1080 78 1106
rect -14 1062 16 1076
rect 43 1072 78 1080
rect 80 1106 121 1114
rect 80 1080 95 1106
rect 102 1080 121 1106
rect 185 1102 216 1114
rect 231 1102 334 1114
rect 346 1104 372 1130
rect 387 1125 417 1136
rect 449 1132 511 1148
rect 449 1130 495 1132
rect 449 1114 511 1130
rect 523 1114 529 1162
rect 532 1154 612 1162
rect 532 1152 551 1154
rect 566 1152 600 1154
rect 532 1136 612 1152
rect 532 1114 551 1136
rect 566 1120 596 1136
rect 624 1130 630 1204
rect 633 1130 652 1274
rect 667 1130 673 1274
rect 682 1204 695 1274
rect 747 1270 769 1274
rect 740 1258 757 1262
rect 761 1260 769 1262
rect 759 1258 769 1260
rect 740 1248 769 1258
rect 822 1248 838 1262
rect 876 1258 882 1260
rect 889 1258 997 1274
rect 1004 1258 1010 1260
rect 1018 1258 1033 1274
rect 1099 1268 1118 1271
rect 740 1246 838 1248
rect 865 1246 1033 1258
rect 1048 1248 1064 1262
rect 1099 1249 1121 1268
rect 1131 1262 1147 1263
rect 1130 1260 1147 1262
rect 1131 1255 1147 1260
rect 1121 1248 1127 1249
rect 1130 1248 1159 1255
rect 1048 1247 1159 1248
rect 1048 1246 1165 1247
rect 724 1238 775 1246
rect 822 1238 856 1246
rect 724 1226 749 1238
rect 756 1226 775 1238
rect 829 1236 856 1238
rect 865 1236 1086 1246
rect 1121 1243 1127 1246
rect 829 1232 1086 1236
rect 724 1218 775 1226
rect 822 1218 1086 1232
rect 1130 1238 1165 1246
rect 676 1170 695 1204
rect 740 1210 769 1218
rect 740 1204 757 1210
rect 740 1202 774 1204
rect 822 1202 838 1218
rect 839 1208 1047 1218
rect 1048 1208 1064 1218
rect 1112 1214 1127 1229
rect 1130 1226 1131 1238
rect 1138 1226 1165 1238
rect 1130 1218 1165 1226
rect 1130 1217 1159 1218
rect 850 1204 1064 1208
rect 865 1202 1064 1204
rect 1099 1204 1112 1214
rect 1130 1204 1147 1217
rect 1099 1202 1147 1204
rect 741 1198 774 1202
rect 737 1196 774 1198
rect 737 1195 804 1196
rect 737 1190 768 1195
rect 774 1190 804 1195
rect 737 1186 804 1190
rect 710 1183 804 1186
rect 710 1176 759 1183
rect 710 1170 740 1176
rect 759 1171 764 1176
rect 676 1154 756 1170
rect 768 1162 804 1183
rect 865 1178 1054 1202
rect 1099 1201 1146 1202
rect 1112 1196 1146 1201
rect 880 1175 1054 1178
rect 873 1172 1054 1175
rect 1082 1195 1146 1196
rect 676 1152 695 1154
rect 710 1152 744 1154
rect 676 1136 756 1152
rect 676 1130 695 1136
rect 392 1104 495 1114
rect 346 1102 495 1104
rect 516 1102 551 1114
rect 185 1100 347 1102
rect 197 1080 216 1100
rect 231 1098 261 1100
rect 80 1072 121 1080
rect 203 1076 216 1080
rect 268 1084 347 1100
rect 379 1100 551 1102
rect 379 1084 458 1100
rect 465 1098 495 1100
rect 43 1062 72 1072
rect 86 1062 115 1072
rect 130 1062 160 1076
rect 203 1062 246 1076
rect 268 1072 458 1084
rect 523 1080 529 1100
rect 253 1062 283 1072
rect 284 1062 442 1072
rect 446 1062 476 1072
rect 480 1062 510 1076
rect 538 1062 551 1100
rect 623 1114 652 1130
rect 666 1114 695 1130
rect 710 1120 740 1136
rect 768 1114 774 1162
rect 777 1156 796 1162
rect 811 1156 841 1164
rect 777 1148 841 1156
rect 777 1132 857 1148
rect 873 1141 935 1172
rect 951 1141 1013 1172
rect 1082 1170 1131 1195
rect 1146 1170 1176 1188
rect 1045 1156 1075 1164
rect 1082 1162 1192 1170
rect 1045 1148 1090 1156
rect 777 1130 796 1132
rect 811 1130 857 1132
rect 777 1114 857 1130
rect 884 1128 919 1141
rect 960 1138 997 1141
rect 960 1136 1002 1138
rect 889 1125 919 1128
rect 898 1121 905 1125
rect 905 1120 906 1121
rect 864 1114 874 1120
rect 623 1106 658 1114
rect 623 1080 624 1106
rect 631 1080 658 1106
rect 566 1062 596 1076
rect 623 1072 658 1080
rect 660 1106 701 1114
rect 660 1080 675 1106
rect 682 1080 701 1106
rect 765 1102 796 1114
rect 811 1102 914 1114
rect 926 1104 952 1130
rect 967 1125 997 1136
rect 1029 1132 1091 1148
rect 1029 1130 1075 1132
rect 1029 1114 1091 1130
rect 1103 1114 1109 1162
rect 1112 1154 1192 1162
rect 1112 1152 1131 1154
rect 1146 1152 1180 1154
rect 1112 1137 1192 1152
rect 1112 1136 1198 1137
rect 1112 1114 1131 1136
rect 1146 1120 1176 1136
rect 1204 1130 1210 1204
rect 1213 1130 1232 1274
rect 1247 1130 1253 1274
rect 1262 1204 1275 1274
rect 1327 1270 1349 1274
rect 1320 1258 1337 1262
rect 1341 1260 1349 1262
rect 1339 1258 1349 1260
rect 1320 1248 1349 1258
rect 1402 1248 1418 1262
rect 1456 1258 1462 1260
rect 1469 1258 1577 1274
rect 1584 1258 1590 1260
rect 1598 1258 1613 1274
rect 1679 1268 1698 1271
rect 1320 1246 1418 1248
rect 1445 1246 1613 1258
rect 1628 1248 1644 1262
rect 1679 1249 1701 1268
rect 1711 1262 1727 1263
rect 1710 1260 1727 1262
rect 1711 1255 1727 1260
rect 1701 1248 1707 1249
rect 1710 1248 1739 1255
rect 1628 1247 1739 1248
rect 1628 1246 1745 1247
rect 1304 1238 1355 1246
rect 1402 1238 1436 1246
rect 1304 1226 1329 1238
rect 1336 1226 1355 1238
rect 1409 1236 1436 1238
rect 1445 1236 1666 1246
rect 1701 1243 1707 1246
rect 1409 1232 1666 1236
rect 1304 1218 1355 1226
rect 1402 1218 1666 1232
rect 1710 1238 1745 1246
rect 1256 1170 1275 1204
rect 1320 1210 1349 1218
rect 1320 1204 1337 1210
rect 1320 1202 1354 1204
rect 1402 1202 1418 1218
rect 1419 1208 1627 1218
rect 1628 1208 1644 1218
rect 1692 1214 1707 1229
rect 1710 1226 1711 1238
rect 1718 1226 1745 1238
rect 1710 1218 1745 1226
rect 1710 1217 1739 1218
rect 1430 1204 1644 1208
rect 1445 1202 1644 1204
rect 1679 1204 1692 1214
rect 1710 1204 1727 1217
rect 1679 1202 1727 1204
rect 1321 1198 1354 1202
rect 1317 1196 1354 1198
rect 1317 1195 1384 1196
rect 1317 1190 1348 1195
rect 1354 1190 1384 1195
rect 1317 1186 1384 1190
rect 1290 1183 1384 1186
rect 1290 1176 1339 1183
rect 1290 1170 1320 1176
rect 1339 1171 1344 1176
rect 1256 1154 1336 1170
rect 1348 1162 1384 1183
rect 1445 1178 1634 1202
rect 1679 1201 1726 1202
rect 1692 1196 1726 1201
rect 1766 1196 1782 1198
rect 1460 1175 1634 1178
rect 1453 1172 1634 1175
rect 1662 1195 1726 1196
rect 1256 1152 1275 1154
rect 1290 1152 1324 1154
rect 1256 1136 1336 1152
rect 1256 1130 1275 1136
rect 972 1104 1075 1114
rect 926 1102 1075 1104
rect 1096 1102 1131 1114
rect 765 1100 927 1102
rect 777 1080 796 1100
rect 811 1098 841 1100
rect 660 1072 701 1080
rect 783 1076 796 1080
rect 848 1084 927 1100
rect 959 1100 1131 1102
rect 959 1084 1038 1100
rect 1045 1098 1075 1100
rect 623 1062 652 1072
rect 666 1062 695 1072
rect 710 1062 740 1076
rect 783 1062 826 1076
rect 848 1072 1038 1084
rect 1103 1080 1109 1100
rect 833 1062 863 1072
rect 864 1062 1022 1072
rect 1026 1062 1056 1072
rect 1060 1062 1090 1076
rect 1118 1062 1131 1100
rect 1203 1114 1232 1130
rect 1246 1114 1275 1130
rect 1290 1120 1320 1136
rect 1348 1114 1354 1162
rect 1357 1156 1376 1162
rect 1391 1156 1421 1164
rect 1357 1148 1421 1156
rect 1357 1132 1437 1148
rect 1453 1141 1515 1172
rect 1531 1141 1593 1172
rect 1662 1170 1711 1195
rect 1756 1186 1782 1196
rect 1726 1170 1782 1186
rect 1625 1156 1655 1164
rect 1662 1162 1772 1170
rect 1625 1148 1670 1156
rect 1357 1130 1376 1132
rect 1391 1130 1437 1132
rect 1357 1114 1437 1130
rect 1464 1128 1499 1141
rect 1540 1138 1577 1141
rect 1540 1136 1582 1138
rect 1469 1125 1499 1128
rect 1478 1121 1485 1125
rect 1485 1120 1486 1121
rect 1444 1114 1454 1120
rect 1203 1106 1238 1114
rect 1203 1080 1204 1106
rect 1211 1080 1238 1106
rect 1146 1062 1176 1076
rect 1203 1072 1238 1080
rect 1240 1106 1281 1114
rect 1240 1080 1255 1106
rect 1262 1080 1281 1106
rect 1345 1102 1376 1114
rect 1391 1102 1494 1114
rect 1506 1104 1532 1130
rect 1547 1125 1577 1136
rect 1609 1132 1671 1148
rect 1609 1130 1655 1132
rect 1609 1114 1671 1130
rect 1683 1114 1689 1162
rect 1692 1154 1772 1162
rect 1692 1152 1711 1154
rect 1726 1152 1760 1154
rect 1692 1136 1772 1152
rect 1692 1114 1711 1136
rect 1726 1120 1756 1136
rect 1784 1130 1790 1204
rect 1793 1130 1812 1274
rect 1827 1130 1833 1274
rect 1842 1204 1855 1274
rect 1907 1270 1929 1274
rect 1900 1258 1917 1262
rect 1921 1260 1929 1262
rect 1919 1258 1929 1260
rect 1900 1248 1929 1258
rect 1982 1248 1998 1262
rect 2036 1258 2042 1260
rect 2049 1258 2157 1274
rect 2164 1258 2170 1260
rect 2178 1258 2193 1274
rect 2259 1268 2278 1271
rect 1900 1246 1998 1248
rect 2025 1246 2193 1258
rect 2208 1248 2224 1262
rect 2259 1249 2281 1268
rect 2291 1262 2307 1263
rect 2290 1256 2307 1262
rect 2291 1255 2307 1256
rect 2281 1248 2287 1249
rect 2290 1248 2319 1255
rect 2208 1247 2319 1248
rect 2208 1246 2325 1247
rect 1884 1238 1935 1246
rect 1982 1238 2016 1246
rect 1884 1226 1909 1238
rect 1916 1226 1935 1238
rect 1989 1236 2016 1238
rect 2025 1236 2246 1246
rect 2281 1243 2287 1246
rect 1989 1232 2246 1236
rect 1884 1218 1935 1226
rect 1982 1218 2246 1232
rect 2290 1238 2325 1246
rect 1836 1170 1855 1204
rect 1900 1210 1929 1218
rect 1900 1204 1917 1210
rect 1900 1202 1934 1204
rect 1982 1202 1998 1218
rect 1999 1208 2207 1218
rect 2208 1208 2224 1218
rect 2272 1214 2287 1229
rect 2290 1226 2291 1238
rect 2298 1226 2325 1238
rect 2290 1218 2325 1226
rect 2290 1217 2319 1218
rect 2010 1204 2224 1208
rect 2025 1202 2224 1204
rect 2259 1204 2272 1214
rect 2290 1204 2307 1217
rect 2259 1202 2307 1204
rect 1901 1198 1934 1202
rect 1897 1196 1934 1198
rect 1897 1195 1964 1196
rect 1897 1190 1928 1195
rect 1934 1190 1964 1195
rect 1897 1186 1964 1190
rect 1870 1183 1964 1186
rect 1870 1176 1919 1183
rect 1870 1170 1900 1176
rect 1919 1171 1924 1176
rect 1836 1154 1916 1170
rect 1928 1162 1964 1183
rect 2025 1178 2214 1202
rect 2259 1201 2306 1202
rect 2272 1196 2306 1201
rect 2040 1175 2214 1178
rect 2033 1172 2214 1175
rect 2242 1195 2306 1196
rect 1836 1152 1855 1154
rect 1870 1152 1904 1154
rect 1836 1136 1916 1152
rect 1836 1130 1855 1136
rect 1552 1104 1655 1114
rect 1506 1102 1655 1104
rect 1676 1102 1711 1114
rect 1345 1100 1507 1102
rect 1357 1080 1376 1100
rect 1391 1098 1421 1100
rect 1240 1072 1281 1080
rect 1363 1076 1376 1080
rect 1428 1084 1507 1100
rect 1539 1100 1711 1102
rect 1539 1084 1618 1100
rect 1625 1098 1655 1100
rect 1203 1062 1232 1072
rect 1246 1062 1275 1072
rect 1290 1062 1320 1076
rect 1363 1062 1406 1076
rect 1428 1072 1618 1084
rect 1683 1080 1689 1100
rect 1413 1062 1443 1072
rect 1444 1062 1602 1072
rect 1606 1062 1636 1072
rect 1640 1062 1670 1076
rect 1698 1062 1711 1100
rect 1783 1114 1812 1130
rect 1826 1114 1855 1130
rect 1870 1120 1900 1136
rect 1928 1114 1934 1162
rect 1937 1156 1956 1162
rect 1971 1156 2001 1164
rect 1937 1148 2001 1156
rect 1937 1132 2017 1148
rect 2033 1141 2095 1172
rect 2111 1141 2173 1172
rect 2242 1170 2291 1195
rect 2306 1170 2336 1188
rect 2205 1156 2235 1164
rect 2242 1162 2352 1170
rect 2205 1148 2250 1156
rect 1937 1130 1956 1132
rect 1971 1130 2017 1132
rect 1937 1114 2017 1130
rect 2044 1128 2079 1141
rect 2120 1138 2157 1141
rect 2120 1136 2162 1138
rect 2049 1125 2079 1128
rect 2058 1121 2065 1125
rect 2065 1120 2066 1121
rect 2024 1114 2034 1120
rect 1783 1106 1818 1114
rect 1783 1080 1784 1106
rect 1791 1080 1818 1106
rect 1726 1062 1756 1076
rect 1783 1072 1818 1080
rect 1820 1106 1861 1114
rect 1820 1080 1835 1106
rect 1842 1080 1861 1106
rect 1925 1102 1956 1114
rect 1971 1102 2074 1114
rect 2086 1104 2112 1130
rect 2127 1125 2157 1136
rect 2189 1132 2251 1148
rect 2189 1130 2235 1132
rect 2189 1114 2251 1130
rect 2263 1114 2269 1162
rect 2272 1154 2352 1162
rect 2272 1152 2291 1154
rect 2306 1152 2340 1154
rect 2272 1137 2352 1152
rect 2272 1136 2358 1137
rect 2272 1114 2291 1136
rect 2306 1120 2336 1136
rect 2364 1130 2370 1204
rect 2373 1130 2392 1274
rect 2407 1130 2413 1274
rect 2422 1204 2435 1274
rect 2487 1270 2509 1274
rect 2480 1258 2497 1262
rect 2501 1260 2509 1262
rect 2499 1258 2509 1260
rect 2480 1248 2509 1258
rect 2562 1248 2578 1262
rect 2616 1258 2622 1260
rect 2629 1258 2737 1274
rect 2744 1258 2750 1260
rect 2758 1258 2773 1274
rect 2839 1268 2858 1271
rect 2480 1246 2578 1248
rect 2605 1246 2773 1258
rect 2788 1248 2804 1262
rect 2839 1249 2861 1268
rect 2871 1262 2887 1263
rect 2870 1256 2887 1262
rect 2871 1255 2887 1256
rect 2861 1248 2867 1249
rect 2870 1248 2899 1255
rect 2788 1247 2899 1248
rect 2788 1246 2905 1247
rect 2464 1238 2515 1246
rect 2562 1238 2596 1246
rect 2464 1226 2489 1238
rect 2496 1226 2515 1238
rect 2569 1236 2596 1238
rect 2605 1236 2826 1246
rect 2861 1243 2867 1246
rect 2569 1232 2826 1236
rect 2464 1218 2515 1226
rect 2562 1218 2826 1232
rect 2870 1238 2905 1246
rect 2416 1170 2435 1204
rect 2480 1210 2509 1218
rect 2480 1204 2497 1210
rect 2480 1202 2514 1204
rect 2562 1202 2578 1218
rect 2579 1208 2787 1218
rect 2788 1208 2804 1218
rect 2852 1214 2867 1229
rect 2870 1226 2871 1238
rect 2878 1226 2905 1238
rect 2870 1218 2905 1226
rect 2870 1217 2899 1218
rect 2590 1204 2804 1208
rect 2605 1202 2804 1204
rect 2839 1204 2852 1214
rect 2870 1204 2887 1217
rect 2839 1202 2887 1204
rect 2481 1198 2514 1202
rect 2477 1196 2514 1198
rect 2477 1195 2544 1196
rect 2477 1190 2508 1195
rect 2514 1190 2544 1195
rect 2477 1186 2544 1190
rect 2450 1183 2544 1186
rect 2450 1176 2499 1183
rect 2450 1170 2480 1176
rect 2499 1171 2504 1176
rect 2416 1154 2496 1170
rect 2508 1162 2544 1183
rect 2605 1178 2794 1202
rect 2839 1201 2886 1202
rect 2852 1196 2886 1201
rect 2926 1196 2942 1198
rect 2620 1175 2794 1178
rect 2613 1172 2794 1175
rect 2822 1195 2886 1196
rect 2416 1152 2435 1154
rect 2450 1152 2484 1154
rect 2416 1136 2496 1152
rect 2416 1130 2435 1136
rect 2132 1104 2235 1114
rect 2086 1102 2235 1104
rect 2256 1102 2291 1114
rect 1925 1100 2087 1102
rect 1937 1080 1956 1100
rect 1971 1098 2001 1100
rect 1820 1072 1861 1080
rect 1943 1076 1956 1080
rect 2008 1084 2087 1100
rect 2119 1100 2291 1102
rect 2119 1084 2198 1100
rect 2205 1098 2235 1100
rect 1783 1062 1812 1072
rect 1826 1062 1855 1072
rect 1870 1062 1900 1076
rect 1943 1062 1986 1076
rect 2008 1072 2198 1084
rect 2263 1080 2269 1100
rect 1993 1062 2023 1072
rect 2024 1062 2182 1072
rect 2186 1062 2216 1072
rect 2220 1062 2250 1076
rect 2278 1062 2291 1100
rect 2363 1114 2392 1130
rect 2406 1114 2435 1130
rect 2450 1120 2480 1136
rect 2508 1114 2514 1162
rect 2517 1156 2536 1162
rect 2551 1156 2581 1164
rect 2517 1148 2581 1156
rect 2517 1132 2597 1148
rect 2613 1141 2675 1172
rect 2691 1141 2753 1172
rect 2822 1170 2871 1195
rect 2916 1186 2942 1196
rect 2886 1170 2942 1186
rect 2785 1156 2815 1164
rect 2822 1162 2932 1170
rect 2785 1148 2830 1156
rect 2517 1130 2536 1132
rect 2551 1130 2597 1132
rect 2517 1114 2597 1130
rect 2624 1128 2659 1141
rect 2700 1138 2737 1141
rect 2700 1136 2742 1138
rect 2629 1125 2659 1128
rect 2638 1121 2645 1125
rect 2645 1120 2646 1121
rect 2604 1114 2614 1120
rect 2363 1106 2398 1114
rect 2363 1080 2364 1106
rect 2371 1080 2398 1106
rect 2306 1062 2336 1076
rect 2363 1072 2398 1080
rect 2400 1106 2441 1114
rect 2400 1080 2415 1106
rect 2422 1080 2441 1106
rect 2505 1102 2536 1114
rect 2551 1102 2654 1114
rect 2666 1104 2692 1130
rect 2707 1125 2737 1136
rect 2769 1132 2831 1148
rect 2769 1130 2815 1132
rect 2769 1114 2831 1130
rect 2843 1114 2849 1162
rect 2852 1154 2932 1162
rect 2852 1152 2871 1154
rect 2886 1152 2920 1154
rect 2852 1136 2932 1152
rect 2852 1114 2871 1136
rect 2886 1120 2916 1136
rect 2944 1130 2950 1204
rect 2953 1130 2972 1274
rect 2987 1130 2993 1274
rect 3002 1204 3015 1274
rect 3067 1270 3089 1274
rect 3060 1258 3077 1262
rect 3081 1260 3089 1262
rect 3079 1258 3089 1260
rect 3060 1248 3089 1258
rect 3142 1248 3158 1262
rect 3196 1258 3202 1260
rect 3209 1258 3317 1274
rect 3324 1258 3330 1260
rect 3338 1258 3353 1274
rect 3419 1268 3438 1271
rect 3060 1246 3158 1248
rect 3185 1246 3353 1258
rect 3368 1248 3384 1262
rect 3419 1249 3441 1268
rect 3451 1262 3467 1263
rect 3450 1256 3467 1262
rect 3451 1255 3467 1256
rect 3441 1248 3447 1249
rect 3450 1248 3479 1255
rect 3368 1247 3479 1248
rect 3368 1246 3485 1247
rect 3044 1238 3095 1246
rect 3142 1238 3176 1246
rect 3044 1226 3069 1238
rect 3076 1226 3095 1238
rect 3149 1236 3176 1238
rect 3185 1236 3406 1246
rect 3441 1243 3447 1246
rect 3149 1232 3406 1236
rect 3044 1218 3095 1226
rect 3142 1218 3406 1232
rect 3450 1238 3485 1246
rect 2996 1170 3015 1204
rect 3060 1210 3089 1218
rect 3060 1204 3077 1210
rect 3060 1202 3094 1204
rect 3142 1202 3158 1218
rect 3159 1208 3367 1218
rect 3368 1208 3384 1218
rect 3432 1214 3447 1229
rect 3450 1226 3451 1238
rect 3458 1226 3485 1238
rect 3450 1218 3485 1226
rect 3450 1217 3479 1218
rect 3170 1204 3384 1208
rect 3185 1202 3384 1204
rect 3419 1204 3432 1214
rect 3450 1204 3467 1217
rect 3419 1202 3467 1204
rect 3061 1198 3094 1202
rect 3057 1196 3094 1198
rect 3057 1195 3124 1196
rect 3057 1190 3088 1195
rect 3094 1190 3124 1195
rect 3057 1186 3124 1190
rect 3030 1183 3124 1186
rect 3030 1176 3079 1183
rect 3030 1170 3060 1176
rect 3079 1171 3084 1176
rect 2996 1154 3076 1170
rect 3088 1162 3124 1183
rect 3185 1178 3374 1202
rect 3419 1201 3466 1202
rect 3432 1196 3466 1201
rect 3200 1175 3374 1178
rect 3193 1172 3374 1175
rect 3402 1195 3466 1196
rect 2996 1152 3015 1154
rect 3030 1152 3064 1154
rect 2996 1136 3076 1152
rect 2996 1130 3015 1136
rect 2712 1104 2815 1114
rect 2666 1102 2815 1104
rect 2836 1102 2871 1114
rect 2505 1100 2667 1102
rect 2517 1080 2536 1100
rect 2551 1098 2581 1100
rect 2400 1072 2441 1080
rect 2523 1076 2536 1080
rect 2588 1084 2667 1100
rect 2699 1100 2871 1102
rect 2699 1084 2778 1100
rect 2785 1098 2815 1100
rect 2363 1062 2392 1072
rect 2406 1062 2435 1072
rect 2450 1062 2480 1076
rect 2523 1062 2566 1076
rect 2588 1072 2778 1084
rect 2843 1080 2849 1100
rect 2573 1062 2603 1072
rect 2604 1062 2762 1072
rect 2766 1062 2796 1072
rect 2800 1062 2830 1076
rect 2858 1062 2871 1100
rect 2943 1114 2972 1130
rect 2986 1114 3015 1130
rect 3030 1120 3060 1136
rect 3088 1114 3094 1162
rect 3097 1156 3116 1162
rect 3131 1156 3161 1164
rect 3097 1148 3161 1156
rect 3097 1132 3177 1148
rect 3193 1141 3255 1172
rect 3271 1141 3333 1172
rect 3402 1170 3451 1195
rect 3466 1170 3496 1188
rect 3365 1156 3395 1164
rect 3402 1162 3512 1170
rect 3365 1148 3410 1156
rect 3097 1130 3116 1132
rect 3131 1130 3177 1132
rect 3097 1114 3177 1130
rect 3204 1128 3239 1141
rect 3280 1138 3317 1141
rect 3280 1136 3322 1138
rect 3209 1125 3239 1128
rect 3218 1121 3225 1125
rect 3225 1120 3226 1121
rect 3184 1114 3194 1120
rect 2943 1106 2978 1114
rect 2943 1080 2944 1106
rect 2951 1080 2978 1106
rect 2886 1062 2916 1076
rect 2943 1072 2978 1080
rect 2980 1106 3021 1114
rect 2980 1080 2995 1106
rect 3002 1080 3021 1106
rect 3085 1102 3116 1114
rect 3131 1102 3234 1114
rect 3246 1104 3272 1130
rect 3287 1125 3317 1136
rect 3349 1132 3411 1148
rect 3349 1130 3395 1132
rect 3349 1114 3411 1130
rect 3423 1114 3429 1162
rect 3432 1154 3512 1162
rect 3432 1152 3451 1154
rect 3466 1152 3500 1154
rect 3432 1137 3512 1152
rect 3432 1136 3518 1137
rect 3432 1114 3451 1136
rect 3466 1120 3496 1136
rect 3524 1130 3530 1204
rect 3533 1130 3552 1274
rect 3567 1130 3573 1274
rect 3582 1204 3595 1274
rect 3647 1270 3669 1274
rect 3640 1258 3657 1262
rect 3661 1260 3669 1262
rect 3659 1258 3669 1260
rect 3640 1248 3669 1258
rect 3722 1248 3738 1262
rect 3776 1258 3782 1260
rect 3789 1258 3897 1274
rect 3904 1258 3910 1260
rect 3918 1258 3933 1274
rect 3999 1268 4018 1271
rect 3640 1246 3738 1248
rect 3765 1246 3933 1258
rect 3948 1248 3964 1262
rect 3999 1249 4021 1268
rect 4031 1262 4047 1263
rect 4030 1256 4047 1262
rect 4031 1255 4047 1256
rect 4021 1248 4027 1249
rect 4030 1248 4059 1255
rect 3948 1247 4059 1248
rect 3948 1246 4065 1247
rect 3624 1238 3675 1246
rect 3722 1238 3756 1246
rect 3624 1226 3649 1238
rect 3656 1226 3675 1238
rect 3729 1236 3756 1238
rect 3765 1236 3986 1246
rect 4021 1243 4027 1246
rect 3729 1232 3986 1236
rect 3624 1218 3675 1226
rect 3722 1218 3986 1232
rect 4030 1238 4065 1246
rect 3576 1170 3595 1204
rect 3640 1210 3669 1218
rect 3640 1204 3657 1210
rect 3640 1202 3674 1204
rect 3722 1202 3738 1218
rect 3739 1208 3947 1218
rect 3948 1208 3964 1218
rect 4012 1214 4027 1229
rect 4030 1226 4031 1238
rect 4038 1226 4065 1238
rect 4030 1218 4065 1226
rect 4030 1217 4059 1218
rect 3750 1204 3964 1208
rect 3765 1202 3964 1204
rect 3999 1204 4012 1214
rect 4030 1204 4047 1217
rect 3999 1202 4047 1204
rect 3641 1198 3674 1202
rect 3637 1196 3674 1198
rect 3637 1195 3704 1196
rect 3637 1190 3668 1195
rect 3674 1190 3704 1195
rect 3637 1186 3704 1190
rect 3610 1183 3704 1186
rect 3610 1176 3659 1183
rect 3610 1170 3640 1176
rect 3659 1171 3664 1176
rect 3576 1154 3656 1170
rect 3668 1162 3704 1183
rect 3765 1178 3954 1202
rect 3999 1201 4046 1202
rect 4012 1196 4046 1201
rect 4086 1196 4102 1198
rect 3780 1175 3954 1178
rect 3773 1172 3954 1175
rect 3982 1195 4046 1196
rect 3576 1152 3595 1154
rect 3610 1152 3644 1154
rect 3576 1136 3656 1152
rect 3576 1130 3595 1136
rect 3292 1104 3395 1114
rect 3246 1102 3395 1104
rect 3416 1102 3451 1114
rect 3085 1100 3247 1102
rect 3097 1080 3116 1100
rect 3131 1098 3161 1100
rect 2980 1072 3021 1080
rect 3103 1076 3116 1080
rect 3168 1084 3247 1100
rect 3279 1100 3451 1102
rect 3279 1084 3358 1100
rect 3365 1098 3395 1100
rect 2943 1062 2972 1072
rect 2986 1062 3015 1072
rect 3030 1062 3060 1076
rect 3103 1062 3146 1076
rect 3168 1072 3358 1084
rect 3423 1080 3429 1100
rect 3153 1062 3183 1072
rect 3184 1062 3342 1072
rect 3346 1062 3376 1072
rect 3380 1062 3410 1076
rect 3438 1062 3451 1100
rect 3523 1114 3552 1130
rect 3566 1114 3595 1130
rect 3610 1120 3640 1136
rect 3668 1114 3674 1162
rect 3677 1156 3696 1162
rect 3711 1156 3741 1164
rect 3677 1148 3741 1156
rect 3677 1132 3757 1148
rect 3773 1141 3835 1172
rect 3851 1141 3913 1172
rect 3982 1170 4031 1195
rect 4076 1186 4102 1196
rect 4046 1170 4102 1186
rect 3945 1156 3975 1164
rect 3982 1162 4092 1170
rect 3945 1148 3990 1156
rect 3677 1130 3696 1132
rect 3711 1130 3757 1132
rect 3677 1114 3757 1130
rect 3784 1128 3819 1141
rect 3860 1138 3897 1141
rect 3860 1136 3902 1138
rect 3789 1125 3819 1128
rect 3798 1121 3805 1125
rect 3805 1120 3806 1121
rect 3764 1114 3774 1120
rect 3523 1106 3558 1114
rect 3523 1080 3524 1106
rect 3531 1080 3558 1106
rect 3466 1062 3496 1076
rect 3523 1072 3558 1080
rect 3560 1106 3601 1114
rect 3560 1080 3575 1106
rect 3582 1080 3601 1106
rect 3665 1102 3696 1114
rect 3711 1102 3814 1114
rect 3826 1104 3852 1130
rect 3867 1125 3897 1136
rect 3929 1132 3991 1148
rect 3929 1130 3975 1132
rect 3929 1114 3991 1130
rect 4003 1114 4009 1162
rect 4012 1154 4092 1162
rect 4012 1152 4031 1154
rect 4046 1152 4080 1154
rect 4012 1136 4092 1152
rect 4012 1114 4031 1136
rect 4046 1120 4076 1136
rect 4104 1130 4110 1204
rect 4113 1130 4132 1274
rect 4147 1130 4153 1274
rect 4162 1204 4175 1274
rect 4227 1270 4249 1274
rect 4220 1258 4237 1262
rect 4241 1260 4249 1262
rect 4239 1258 4249 1260
rect 4220 1248 4249 1258
rect 4302 1248 4318 1262
rect 4356 1258 4362 1260
rect 4369 1258 4477 1274
rect 4484 1258 4490 1260
rect 4498 1258 4513 1274
rect 4579 1268 4598 1271
rect 4220 1246 4318 1248
rect 4345 1246 4513 1258
rect 4528 1248 4544 1262
rect 4579 1249 4601 1268
rect 4611 1262 4627 1263
rect 4610 1256 4627 1262
rect 4611 1255 4627 1256
rect 4601 1248 4607 1249
rect 4610 1248 4639 1255
rect 4528 1247 4639 1248
rect 4528 1246 4645 1247
rect 4204 1238 4255 1246
rect 4302 1238 4336 1246
rect 4204 1226 4229 1238
rect 4236 1226 4255 1238
rect 4309 1236 4336 1238
rect 4345 1236 4566 1246
rect 4601 1243 4607 1246
rect 4309 1232 4566 1236
rect 4204 1218 4255 1226
rect 4302 1218 4566 1232
rect 4610 1238 4645 1246
rect 4156 1170 4175 1204
rect 4220 1210 4249 1218
rect 4220 1204 4237 1210
rect 4220 1202 4254 1204
rect 4302 1202 4318 1218
rect 4319 1208 4527 1218
rect 4528 1208 4544 1218
rect 4592 1214 4607 1229
rect 4610 1226 4611 1238
rect 4618 1226 4645 1238
rect 4610 1218 4645 1226
rect 4610 1217 4639 1218
rect 4330 1204 4544 1208
rect 4345 1202 4544 1204
rect 4579 1204 4592 1214
rect 4610 1204 4627 1217
rect 4579 1202 4627 1204
rect 4221 1198 4254 1202
rect 4217 1196 4254 1198
rect 4217 1195 4284 1196
rect 4217 1190 4248 1195
rect 4254 1190 4284 1195
rect 4217 1186 4284 1190
rect 4190 1183 4284 1186
rect 4190 1176 4239 1183
rect 4190 1170 4220 1176
rect 4239 1171 4244 1176
rect 4156 1154 4236 1170
rect 4248 1162 4284 1183
rect 4345 1178 4534 1202
rect 4579 1201 4626 1202
rect 4592 1196 4626 1201
rect 4360 1175 4534 1178
rect 4353 1172 4534 1175
rect 4562 1195 4626 1196
rect 4156 1152 4175 1154
rect 4190 1152 4224 1154
rect 4156 1136 4236 1152
rect 4156 1130 4175 1136
rect 3872 1104 3975 1114
rect 3826 1102 3975 1104
rect 3996 1102 4031 1114
rect 3665 1100 3827 1102
rect 3677 1080 3696 1100
rect 3711 1098 3741 1100
rect 3560 1072 3601 1080
rect 3683 1076 3696 1080
rect 3748 1084 3827 1100
rect 3859 1100 4031 1102
rect 3859 1084 3938 1100
rect 3945 1098 3975 1100
rect 3523 1062 3552 1072
rect 3566 1062 3595 1072
rect 3610 1062 3640 1076
rect 3683 1062 3726 1076
rect 3748 1072 3938 1084
rect 4003 1080 4009 1100
rect 3733 1062 3763 1072
rect 3764 1062 3922 1072
rect 3926 1062 3956 1072
rect 3960 1062 3990 1076
rect 4018 1062 4031 1100
rect 4103 1114 4132 1130
rect 4146 1114 4175 1130
rect 4190 1120 4220 1136
rect 4248 1114 4254 1162
rect 4257 1156 4276 1162
rect 4291 1156 4321 1164
rect 4257 1148 4321 1156
rect 4257 1132 4337 1148
rect 4353 1141 4415 1172
rect 4431 1141 4493 1172
rect 4562 1170 4611 1195
rect 4626 1170 4656 1188
rect 4525 1156 4555 1164
rect 4562 1162 4672 1170
rect 4525 1148 4570 1156
rect 4257 1130 4276 1132
rect 4291 1130 4337 1132
rect 4257 1114 4337 1130
rect 4364 1128 4399 1141
rect 4440 1138 4477 1141
rect 4440 1136 4482 1138
rect 4369 1125 4399 1128
rect 4378 1121 4385 1125
rect 4385 1120 4386 1121
rect 4344 1114 4354 1120
rect 4103 1106 4138 1114
rect 4103 1080 4104 1106
rect 4111 1080 4138 1106
rect 4046 1062 4076 1076
rect 4103 1072 4138 1080
rect 4140 1106 4181 1114
rect 4140 1080 4155 1106
rect 4162 1080 4181 1106
rect 4245 1102 4276 1114
rect 4291 1102 4394 1114
rect 4406 1104 4432 1130
rect 4447 1125 4477 1136
rect 4509 1132 4571 1148
rect 4509 1130 4555 1132
rect 4509 1114 4571 1130
rect 4583 1114 4589 1162
rect 4592 1154 4672 1162
rect 4592 1152 4611 1154
rect 4626 1152 4660 1154
rect 4592 1137 4672 1152
rect 4592 1136 4678 1137
rect 4592 1114 4611 1136
rect 4626 1120 4656 1136
rect 4684 1130 4690 1204
rect 4693 1130 4712 1274
rect 4727 1130 4733 1274
rect 4742 1204 4755 1274
rect 4807 1270 4829 1274
rect 4800 1258 4817 1262
rect 4821 1260 4829 1262
rect 4819 1258 4829 1260
rect 4800 1248 4829 1258
rect 4882 1248 4898 1262
rect 4936 1258 4942 1260
rect 4949 1258 5057 1274
rect 5064 1258 5070 1260
rect 5078 1258 5093 1274
rect 5159 1268 5178 1271
rect 4800 1246 4898 1248
rect 4925 1246 5093 1258
rect 5108 1248 5124 1262
rect 5159 1249 5181 1268
rect 5191 1262 5207 1263
rect 5190 1256 5207 1262
rect 5191 1255 5207 1256
rect 5181 1248 5187 1249
rect 5190 1248 5219 1255
rect 5108 1247 5219 1248
rect 5108 1246 5225 1247
rect 4784 1238 4835 1246
rect 4882 1238 4916 1246
rect 4784 1226 4809 1238
rect 4816 1226 4835 1238
rect 4889 1236 4916 1238
rect 4925 1236 5146 1246
rect 5181 1243 5187 1246
rect 4889 1232 5146 1236
rect 4784 1218 4835 1226
rect 4882 1218 5146 1232
rect 5190 1238 5225 1246
rect 4736 1170 4755 1204
rect 4800 1210 4829 1218
rect 4800 1204 4817 1210
rect 4800 1202 4834 1204
rect 4882 1202 4898 1218
rect 4899 1208 5107 1218
rect 5108 1208 5124 1218
rect 5172 1214 5187 1229
rect 5190 1226 5191 1238
rect 5198 1226 5225 1238
rect 5190 1218 5225 1226
rect 5190 1217 5219 1218
rect 4910 1204 5124 1208
rect 4925 1202 5124 1204
rect 5159 1204 5172 1214
rect 5190 1204 5207 1217
rect 5159 1202 5207 1204
rect 4801 1198 4834 1202
rect 4797 1196 4834 1198
rect 4797 1195 4864 1196
rect 4797 1190 4828 1195
rect 4834 1190 4864 1195
rect 4797 1186 4864 1190
rect 4770 1183 4864 1186
rect 4770 1176 4819 1183
rect 4770 1170 4800 1176
rect 4819 1171 4824 1176
rect 4736 1154 4816 1170
rect 4828 1162 4864 1183
rect 4925 1178 5114 1202
rect 5159 1201 5206 1202
rect 5172 1196 5206 1201
rect 5246 1196 5262 1198
rect 4940 1175 5114 1178
rect 4933 1172 5114 1175
rect 5142 1195 5206 1196
rect 4736 1152 4755 1154
rect 4770 1152 4804 1154
rect 4736 1136 4816 1152
rect 4736 1130 4755 1136
rect 4452 1104 4555 1114
rect 4406 1102 4555 1104
rect 4576 1102 4611 1114
rect 4245 1100 4407 1102
rect 4257 1080 4276 1100
rect 4291 1098 4321 1100
rect 4140 1072 4181 1080
rect 4263 1076 4276 1080
rect 4328 1084 4407 1100
rect 4439 1100 4611 1102
rect 4439 1084 4518 1100
rect 4525 1098 4555 1100
rect 4103 1062 4132 1072
rect 4146 1062 4175 1072
rect 4190 1062 4220 1076
rect 4263 1062 4306 1076
rect 4328 1072 4518 1084
rect 4583 1080 4589 1100
rect 4313 1062 4343 1072
rect 4344 1062 4502 1072
rect 4506 1062 4536 1072
rect 4540 1062 4570 1076
rect 4598 1062 4611 1100
rect 4683 1114 4712 1130
rect 4726 1114 4755 1130
rect 4770 1120 4800 1136
rect 4828 1114 4834 1162
rect 4837 1156 4856 1162
rect 4871 1156 4901 1164
rect 4837 1148 4901 1156
rect 4837 1132 4917 1148
rect 4933 1141 4995 1172
rect 5011 1141 5073 1172
rect 5142 1170 5191 1195
rect 5236 1186 5262 1196
rect 5206 1170 5262 1186
rect 5105 1156 5135 1164
rect 5142 1162 5252 1170
rect 5105 1148 5150 1156
rect 4837 1130 4856 1132
rect 4871 1130 4917 1132
rect 4837 1114 4917 1130
rect 4944 1128 4979 1141
rect 5020 1138 5057 1141
rect 5020 1136 5062 1138
rect 4949 1125 4979 1128
rect 4958 1121 4965 1125
rect 4965 1120 4966 1121
rect 4924 1114 4934 1120
rect 4683 1106 4718 1114
rect 4683 1080 4684 1106
rect 4691 1080 4718 1106
rect 4626 1062 4656 1076
rect 4683 1072 4718 1080
rect 4720 1106 4761 1114
rect 4720 1080 4735 1106
rect 4742 1080 4761 1106
rect 4825 1102 4856 1114
rect 4871 1102 4974 1114
rect 4986 1104 5012 1130
rect 5027 1125 5057 1136
rect 5089 1132 5151 1148
rect 5089 1130 5135 1132
rect 5089 1114 5151 1130
rect 5163 1114 5169 1162
rect 5172 1154 5252 1162
rect 5172 1152 5191 1154
rect 5206 1152 5240 1154
rect 5172 1136 5252 1152
rect 5172 1114 5191 1136
rect 5206 1120 5236 1136
rect 5264 1130 5270 1204
rect 5273 1130 5292 1274
rect 5307 1130 5313 1274
rect 5322 1204 5335 1274
rect 5387 1270 5409 1274
rect 5380 1258 5397 1262
rect 5401 1260 5409 1262
rect 5399 1258 5409 1260
rect 5380 1248 5409 1258
rect 5462 1248 5478 1262
rect 5516 1258 5522 1260
rect 5529 1258 5637 1274
rect 5644 1258 5650 1260
rect 5658 1258 5673 1274
rect 5739 1268 5758 1271
rect 5380 1246 5478 1248
rect 5505 1246 5673 1258
rect 5688 1248 5704 1262
rect 5739 1249 5761 1268
rect 5771 1262 5787 1263
rect 5770 1256 5787 1262
rect 5771 1255 5787 1256
rect 5761 1248 5767 1249
rect 5770 1248 5799 1255
rect 5688 1247 5799 1248
rect 5688 1246 5805 1247
rect 5364 1238 5415 1246
rect 5462 1238 5496 1246
rect 5364 1226 5389 1238
rect 5396 1226 5415 1238
rect 5469 1236 5496 1238
rect 5505 1236 5726 1246
rect 5761 1243 5767 1246
rect 5469 1232 5726 1236
rect 5364 1218 5415 1226
rect 5462 1218 5726 1232
rect 5770 1238 5805 1246
rect 5316 1170 5335 1204
rect 5380 1210 5409 1218
rect 5380 1204 5397 1210
rect 5380 1202 5414 1204
rect 5462 1202 5478 1218
rect 5479 1208 5687 1218
rect 5688 1208 5704 1218
rect 5752 1214 5767 1229
rect 5770 1226 5771 1238
rect 5778 1226 5805 1238
rect 5770 1218 5805 1226
rect 5770 1217 5799 1218
rect 5490 1204 5704 1208
rect 5505 1202 5704 1204
rect 5739 1204 5752 1214
rect 5770 1204 5787 1217
rect 5739 1202 5787 1204
rect 5381 1198 5414 1202
rect 5377 1196 5414 1198
rect 5377 1195 5444 1196
rect 5377 1190 5408 1195
rect 5414 1190 5444 1195
rect 5377 1186 5444 1190
rect 5350 1183 5444 1186
rect 5350 1176 5399 1183
rect 5350 1170 5380 1176
rect 5399 1171 5404 1176
rect 5316 1154 5396 1170
rect 5408 1162 5444 1183
rect 5505 1178 5694 1202
rect 5739 1201 5786 1202
rect 5752 1196 5786 1201
rect 5520 1175 5694 1178
rect 5513 1172 5694 1175
rect 5722 1195 5786 1196
rect 5316 1152 5335 1154
rect 5350 1152 5384 1154
rect 5316 1136 5396 1152
rect 5316 1130 5335 1136
rect 5032 1104 5135 1114
rect 4986 1102 5135 1104
rect 5156 1102 5191 1114
rect 4825 1100 4987 1102
rect 4837 1080 4856 1100
rect 4871 1098 4901 1100
rect 4720 1072 4761 1080
rect 4843 1076 4856 1080
rect 4908 1084 4987 1100
rect 5019 1100 5191 1102
rect 5019 1084 5098 1100
rect 5105 1098 5135 1100
rect 4683 1062 4712 1072
rect 4726 1062 4755 1072
rect 4770 1062 4800 1076
rect 4843 1062 4886 1076
rect 4908 1072 5098 1084
rect 5163 1080 5169 1100
rect 4893 1062 4923 1072
rect 4924 1062 5082 1072
rect 5086 1062 5116 1072
rect 5120 1062 5150 1076
rect 5178 1062 5191 1100
rect 5263 1114 5292 1130
rect 5306 1114 5335 1130
rect 5350 1120 5380 1136
rect 5408 1114 5414 1162
rect 5417 1156 5436 1162
rect 5451 1156 5481 1164
rect 5417 1148 5481 1156
rect 5417 1132 5497 1148
rect 5513 1141 5575 1172
rect 5591 1141 5653 1172
rect 5722 1170 5771 1195
rect 5786 1170 5816 1188
rect 5685 1156 5715 1164
rect 5722 1162 5832 1170
rect 5685 1148 5730 1156
rect 5417 1130 5436 1132
rect 5451 1130 5497 1132
rect 5417 1114 5497 1130
rect 5524 1128 5559 1141
rect 5600 1138 5637 1141
rect 5600 1136 5642 1138
rect 5529 1125 5559 1128
rect 5538 1121 5545 1125
rect 5545 1120 5546 1121
rect 5504 1114 5514 1120
rect 5263 1106 5298 1114
rect 5263 1080 5264 1106
rect 5271 1080 5298 1106
rect 5206 1062 5236 1076
rect 5263 1072 5298 1080
rect 5300 1106 5341 1114
rect 5300 1080 5315 1106
rect 5322 1080 5341 1106
rect 5405 1102 5436 1114
rect 5451 1102 5554 1114
rect 5566 1104 5592 1130
rect 5607 1125 5637 1136
rect 5669 1132 5731 1148
rect 5669 1130 5715 1132
rect 5669 1114 5731 1130
rect 5743 1114 5749 1162
rect 5752 1154 5832 1162
rect 5752 1152 5771 1154
rect 5786 1152 5820 1154
rect 5752 1137 5832 1152
rect 5752 1136 5838 1137
rect 5752 1114 5771 1136
rect 5786 1120 5816 1136
rect 5844 1130 5850 1204
rect 5853 1130 5872 1274
rect 5887 1130 5893 1274
rect 5902 1204 5915 1274
rect 5967 1270 5989 1274
rect 5960 1258 5977 1262
rect 5981 1260 5989 1262
rect 5979 1258 5989 1260
rect 5960 1248 5989 1258
rect 6042 1248 6058 1262
rect 6096 1258 6102 1260
rect 6109 1258 6217 1274
rect 6224 1258 6230 1260
rect 6238 1258 6253 1274
rect 6319 1268 6338 1271
rect 5960 1246 6058 1248
rect 6085 1246 6253 1258
rect 6268 1248 6284 1262
rect 6319 1249 6341 1268
rect 6351 1262 6367 1263
rect 6350 1256 6367 1262
rect 6351 1255 6367 1256
rect 6341 1248 6347 1249
rect 6350 1248 6379 1255
rect 6268 1247 6379 1248
rect 6268 1246 6385 1247
rect 5944 1238 5995 1246
rect 6042 1238 6076 1246
rect 5944 1226 5969 1238
rect 5976 1226 5995 1238
rect 6049 1236 6076 1238
rect 6085 1236 6306 1246
rect 6341 1243 6347 1246
rect 6049 1232 6306 1236
rect 5944 1218 5995 1226
rect 6042 1218 6306 1232
rect 6350 1238 6385 1246
rect 5896 1170 5915 1204
rect 5960 1210 5989 1218
rect 5960 1204 5977 1210
rect 5960 1202 5994 1204
rect 6042 1202 6058 1218
rect 6059 1208 6267 1218
rect 6268 1208 6284 1218
rect 6332 1214 6347 1229
rect 6350 1226 6351 1238
rect 6358 1226 6385 1238
rect 6350 1218 6385 1226
rect 6350 1217 6379 1218
rect 6070 1204 6284 1208
rect 6085 1202 6284 1204
rect 6319 1204 6332 1214
rect 6350 1204 6367 1217
rect 6319 1202 6367 1204
rect 5961 1198 5994 1202
rect 5957 1196 5994 1198
rect 5957 1195 6024 1196
rect 5957 1190 5988 1195
rect 5994 1190 6024 1195
rect 5957 1186 6024 1190
rect 5930 1183 6024 1186
rect 5930 1176 5979 1183
rect 5930 1170 5960 1176
rect 5979 1171 5984 1176
rect 5896 1154 5976 1170
rect 5988 1162 6024 1183
rect 6085 1178 6274 1202
rect 6319 1201 6366 1202
rect 6332 1196 6366 1201
rect 6100 1175 6274 1178
rect 6093 1172 6274 1175
rect 6302 1195 6366 1196
rect 5896 1152 5915 1154
rect 5930 1152 5964 1154
rect 5896 1136 5976 1152
rect 5896 1130 5915 1136
rect 5612 1104 5715 1114
rect 5566 1102 5715 1104
rect 5736 1102 5771 1114
rect 5405 1100 5567 1102
rect 5417 1080 5436 1100
rect 5451 1098 5481 1100
rect 5300 1072 5341 1080
rect 5423 1076 5436 1080
rect 5488 1084 5567 1100
rect 5599 1100 5771 1102
rect 5599 1084 5678 1100
rect 5685 1098 5715 1100
rect 5263 1062 5292 1072
rect 5306 1062 5335 1072
rect 5350 1062 5380 1076
rect 5423 1062 5466 1076
rect 5488 1072 5678 1084
rect 5743 1080 5749 1100
rect 5473 1062 5503 1072
rect 5504 1062 5662 1072
rect 5666 1062 5696 1072
rect 5700 1062 5730 1076
rect 5758 1062 5771 1100
rect 5843 1114 5872 1130
rect 5886 1114 5915 1130
rect 5930 1120 5960 1136
rect 5988 1114 5994 1162
rect 5997 1156 6016 1162
rect 6031 1156 6061 1164
rect 5997 1148 6061 1156
rect 5997 1132 6077 1148
rect 6093 1141 6155 1172
rect 6171 1141 6233 1172
rect 6302 1170 6351 1195
rect 6366 1170 6396 1186
rect 6265 1156 6295 1164
rect 6302 1162 6412 1170
rect 6265 1148 6310 1156
rect 5997 1130 6016 1132
rect 6031 1130 6077 1132
rect 5997 1114 6077 1130
rect 6104 1128 6139 1141
rect 6180 1138 6217 1141
rect 6180 1136 6222 1138
rect 6109 1125 6139 1128
rect 6118 1121 6125 1125
rect 6125 1120 6126 1121
rect 6084 1114 6094 1120
rect 5843 1106 5878 1114
rect 5843 1080 5844 1106
rect 5851 1080 5878 1106
rect 5786 1062 5816 1076
rect 5843 1072 5878 1080
rect 5880 1106 5921 1114
rect 5880 1080 5895 1106
rect 5902 1080 5921 1106
rect 5985 1102 6016 1114
rect 6031 1102 6134 1114
rect 6146 1104 6172 1130
rect 6187 1125 6217 1136
rect 6249 1132 6311 1148
rect 6249 1130 6295 1132
rect 6249 1114 6311 1130
rect 6323 1114 6329 1162
rect 6332 1154 6412 1162
rect 6332 1152 6351 1154
rect 6366 1152 6400 1154
rect 6332 1136 6412 1152
rect 6332 1114 6351 1136
rect 6366 1120 6396 1136
rect 6424 1130 6430 1204
rect 6439 1130 6452 1274
rect 6192 1104 6295 1114
rect 6146 1102 6295 1104
rect 6316 1102 6351 1114
rect 5985 1100 6147 1102
rect 5997 1080 6016 1100
rect 6031 1098 6061 1100
rect 5880 1072 5921 1080
rect 6003 1076 6016 1080
rect 6068 1084 6147 1100
rect 6179 1100 6351 1102
rect 6179 1084 6258 1100
rect 6265 1098 6295 1100
rect 5843 1062 5872 1072
rect 5886 1062 5915 1072
rect 5930 1062 5960 1076
rect 6003 1062 6046 1076
rect 6068 1072 6258 1084
rect 6323 1080 6329 1100
rect 6053 1062 6083 1072
rect 6084 1062 6242 1072
rect 6246 1062 6276 1072
rect 6280 1062 6310 1076
rect 6338 1062 6351 1100
rect 6423 1114 6452 1130
rect 6423 1106 6458 1114
rect 6423 1080 6424 1106
rect 6431 1080 6458 1106
rect 6366 1062 6396 1076
rect 6423 1072 6458 1080
rect 6423 1062 6452 1072
rect -541 1048 6452 1062
rect -478 1018 -465 1048
rect -450 1034 -420 1048
rect -377 1034 -334 1048
rect -327 1034 -107 1048
rect -100 1034 -70 1048
rect -410 1020 -395 1032
rect -376 1020 -363 1034
rect -295 1030 -142 1034
rect -413 1018 -391 1020
rect -313 1018 -121 1030
rect -42 1018 -29 1048
rect -14 1034 16 1048
rect 53 1018 72 1048
rect 87 1018 93 1048
rect 102 1018 115 1048
rect 130 1034 160 1048
rect 203 1034 246 1048
rect 253 1034 473 1048
rect 480 1034 510 1048
rect 170 1020 185 1032
rect 204 1020 217 1034
rect 285 1030 438 1034
rect 167 1018 189 1020
rect 267 1018 459 1030
rect 538 1018 551 1048
rect 566 1034 596 1048
rect 633 1018 652 1048
rect 667 1018 673 1048
rect 682 1018 695 1048
rect 710 1034 740 1048
rect 783 1034 826 1048
rect 833 1034 1053 1048
rect 1060 1034 1090 1048
rect 750 1020 765 1032
rect 784 1020 797 1034
rect 865 1030 1018 1034
rect 747 1018 769 1020
rect 847 1018 1039 1030
rect 1118 1018 1131 1048
rect 1146 1034 1176 1048
rect 1213 1018 1232 1048
rect 1247 1018 1253 1048
rect 1262 1018 1275 1048
rect 1290 1034 1320 1048
rect 1363 1034 1406 1048
rect 1413 1034 1633 1048
rect 1640 1034 1670 1048
rect 1330 1020 1345 1032
rect 1364 1020 1377 1034
rect 1445 1030 1598 1034
rect 1327 1018 1349 1020
rect 1427 1018 1619 1030
rect 1698 1018 1711 1048
rect 1726 1034 1756 1048
rect 1793 1018 1812 1048
rect 1827 1018 1833 1048
rect 1842 1018 1855 1048
rect 1870 1034 1900 1048
rect 1943 1034 1986 1048
rect 1993 1034 2213 1048
rect 2220 1034 2250 1048
rect 1910 1020 1925 1032
rect 1944 1020 1957 1034
rect 2025 1030 2178 1034
rect 1907 1018 1929 1020
rect 2007 1018 2199 1030
rect 2278 1018 2291 1048
rect 2306 1034 2336 1048
rect 2373 1018 2392 1048
rect 2407 1018 2413 1048
rect 2422 1018 2435 1048
rect 2450 1034 2480 1048
rect 2523 1034 2566 1048
rect 2573 1034 2793 1048
rect 2800 1034 2830 1048
rect 2490 1020 2505 1032
rect 2524 1020 2537 1034
rect 2605 1030 2758 1034
rect 2487 1018 2509 1020
rect 2587 1018 2779 1030
rect 2858 1018 2871 1048
rect 2886 1034 2916 1048
rect 2953 1018 2972 1048
rect 2987 1018 2993 1048
rect 3002 1018 3015 1048
rect 3030 1034 3060 1048
rect 3103 1034 3146 1048
rect 3153 1034 3373 1048
rect 3380 1034 3410 1048
rect 3070 1020 3085 1032
rect 3104 1020 3117 1034
rect 3185 1030 3338 1034
rect 3067 1018 3089 1020
rect 3167 1018 3359 1030
rect 3438 1018 3451 1048
rect 3466 1034 3496 1048
rect 3533 1018 3552 1048
rect 3567 1018 3573 1048
rect 3582 1018 3595 1048
rect 3610 1034 3640 1048
rect 3683 1034 3726 1048
rect 3733 1034 3953 1048
rect 3960 1034 3990 1048
rect 3650 1020 3665 1032
rect 3684 1020 3697 1034
rect 3765 1030 3918 1034
rect 3647 1018 3669 1020
rect 3747 1018 3939 1030
rect 4018 1018 4031 1048
rect 4046 1034 4076 1048
rect 4113 1018 4132 1048
rect 4147 1018 4153 1048
rect 4162 1018 4175 1048
rect 4190 1034 4220 1048
rect 4263 1034 4306 1048
rect 4313 1034 4533 1048
rect 4540 1034 4570 1048
rect 4230 1020 4245 1032
rect 4264 1020 4277 1034
rect 4345 1030 4498 1034
rect 4227 1018 4249 1020
rect 4327 1018 4519 1030
rect 4598 1018 4611 1048
rect 4626 1034 4656 1048
rect 4693 1018 4712 1048
rect 4727 1018 4733 1048
rect 4742 1018 4755 1048
rect 4770 1034 4800 1048
rect 4843 1034 4886 1048
rect 4893 1034 5113 1048
rect 5120 1034 5150 1048
rect 4810 1020 4825 1032
rect 4844 1020 4857 1034
rect 4925 1030 5078 1034
rect 4807 1018 4829 1020
rect 4907 1018 5099 1030
rect 5178 1018 5191 1048
rect 5206 1034 5236 1048
rect 5273 1018 5292 1048
rect 5307 1018 5313 1048
rect 5322 1018 5335 1048
rect 5350 1034 5380 1048
rect 5423 1034 5466 1048
rect 5473 1034 5693 1048
rect 5700 1034 5730 1048
rect 5390 1020 5405 1032
rect 5424 1020 5437 1034
rect 5505 1030 5658 1034
rect 5387 1018 5409 1020
rect 5487 1018 5679 1030
rect 5758 1018 5771 1048
rect 5786 1034 5816 1048
rect 5853 1018 5872 1048
rect 5887 1018 5893 1048
rect 5902 1018 5915 1048
rect 5930 1034 5960 1048
rect 6003 1034 6046 1048
rect 6053 1034 6273 1048
rect 6280 1034 6310 1048
rect 5970 1020 5985 1032
rect 6004 1020 6017 1034
rect 6085 1030 6238 1034
rect 5967 1018 5989 1020
rect 6067 1018 6259 1030
rect 6338 1018 6351 1048
rect 6366 1034 6396 1048
rect 6439 1018 6452 1048
rect -541 1004 6452 1018
rect -478 934 -465 1004
rect -413 1000 -391 1004
rect -420 988 -403 992
rect -399 990 -391 992
rect -401 988 -391 990
rect -420 978 -391 988
rect -338 978 -322 992
rect -284 988 -278 990
rect -271 988 -163 1004
rect -156 988 -150 990
rect -142 988 -127 1004
rect -61 998 -42 1001
rect -420 976 -322 978
rect -295 976 -127 988
rect -112 978 -96 992
rect -61 979 -39 998
rect -29 992 -13 993
rect -30 990 -13 992
rect -29 985 -13 990
rect -39 978 -33 979
rect -30 978 -1 985
rect -112 977 -1 978
rect -112 976 5 977
rect -436 968 -385 976
rect -338 968 -304 976
rect -436 956 -411 968
rect -404 956 -385 968
rect -331 966 -304 968
rect -295 966 -74 976
rect -39 973 -33 976
rect -331 962 -74 966
rect -436 948 -385 956
rect -338 948 -74 962
rect -30 968 5 976
rect -484 900 -465 934
rect -420 940 -391 948
rect -420 934 -403 940
rect -420 932 -386 934
rect -338 932 -322 948
rect -321 938 -113 948
rect -112 938 -96 948
rect -48 944 -33 959
rect -30 956 -29 968
rect -22 956 5 968
rect -30 948 5 956
rect -30 947 -1 948
rect -310 934 -96 938
rect -295 932 -96 934
rect -61 934 -48 944
rect -30 934 -13 947
rect -61 932 -13 934
rect -419 928 -386 932
rect -423 926 -386 928
rect -423 925 -356 926
rect -423 920 -392 925
rect -386 920 -356 925
rect -423 916 -356 920
rect -450 913 -356 916
rect -450 906 -401 913
rect -450 900 -420 906
rect -401 901 -396 906
rect -484 884 -404 900
rect -392 892 -356 913
rect -295 908 -106 932
rect -61 931 -14 932
rect -48 926 -14 931
rect -280 905 -106 908
rect -287 902 -106 905
rect -78 925 -14 926
rect -484 882 -465 884
rect -450 882 -416 884
rect -484 866 -404 882
rect -484 860 -465 866
rect -494 844 -465 860
rect -450 850 -420 866
rect -392 844 -386 892
rect -383 886 -364 892
rect -349 886 -319 894
rect -383 878 -319 886
rect -383 862 -303 878
rect -287 871 -225 902
rect -209 871 -147 902
rect -78 900 -29 925
rect -14 900 16 918
rect -115 886 -85 894
rect -78 892 32 900
rect -115 878 -70 886
rect -383 860 -364 862
rect -349 860 -303 862
rect -383 844 -303 860
rect -276 858 -241 871
rect -200 868 -163 871
rect -200 866 -158 868
rect -271 855 -241 858
rect -262 851 -255 855
rect -255 850 -254 851
rect -296 844 -286 850
rect -500 836 -459 844
rect -500 810 -485 836
rect -478 810 -459 836
rect -395 832 -364 844
rect -349 832 -246 844
rect -234 834 -208 860
rect -193 855 -163 866
rect -131 862 -69 878
rect -131 860 -85 862
rect -131 844 -69 860
rect -57 844 -51 892
rect -48 884 32 892
rect -48 882 -29 884
rect -14 882 20 884
rect -48 867 32 882
rect -48 866 38 867
rect -48 844 -29 866
rect -14 850 16 866
rect 44 860 50 934
rect 53 860 72 1004
rect 87 860 93 1004
rect 102 934 115 1004
rect 167 1000 189 1004
rect 160 988 177 992
rect 181 990 189 992
rect 179 988 189 990
rect 160 978 189 988
rect 242 978 258 992
rect 296 988 302 990
rect 309 988 417 1004
rect 424 988 430 990
rect 438 988 453 1004
rect 519 998 538 1001
rect 160 976 258 978
rect 285 976 453 988
rect 468 978 484 992
rect 519 979 541 998
rect 551 992 567 993
rect 550 990 567 992
rect 551 985 567 990
rect 541 978 547 979
rect 550 978 579 985
rect 468 977 579 978
rect 468 976 585 977
rect 144 968 195 976
rect 242 968 276 976
rect 144 956 169 968
rect 176 956 195 968
rect 249 966 276 968
rect 285 966 506 976
rect 541 973 547 976
rect 249 962 506 966
rect 144 948 195 956
rect 242 948 506 962
rect 550 968 585 976
rect 96 900 115 934
rect 160 940 189 948
rect 160 934 177 940
rect 160 932 194 934
rect 242 932 258 948
rect 259 938 467 948
rect 468 938 484 948
rect 532 944 547 959
rect 550 956 551 968
rect 558 956 585 968
rect 550 948 585 956
rect 550 947 579 948
rect 270 934 484 938
rect 285 932 484 934
rect 519 934 532 944
rect 550 934 567 947
rect 519 932 567 934
rect 161 928 194 932
rect 157 926 194 928
rect 157 925 224 926
rect 157 920 188 925
rect 194 920 224 925
rect 157 916 224 920
rect 130 913 224 916
rect 130 906 179 913
rect 130 900 160 906
rect 179 901 184 906
rect 96 884 176 900
rect 188 892 224 913
rect 285 908 474 932
rect 519 931 566 932
rect 532 926 566 931
rect 606 926 622 928
rect 300 905 474 908
rect 293 902 474 905
rect 502 925 566 926
rect 96 882 115 884
rect 130 882 164 884
rect 96 866 176 882
rect 96 860 115 866
rect -188 834 -85 844
rect -234 832 -85 834
rect -64 832 -29 844
rect -395 830 -233 832
rect -383 812 -364 830
rect -349 828 -319 830
rect -500 802 -459 810
rect -376 806 -364 812
rect -312 812 -233 830
rect -201 830 -29 832
rect -201 814 -122 830
rect -115 828 -85 830
rect -226 812 -122 814
rect -494 792 -465 802
rect -450 792 -420 806
rect -376 792 -334 806
rect -312 802 -122 812
rect -57 810 -51 830
rect -327 792 -297 802
rect -296 792 -138 802
rect -134 792 -104 802
rect -100 792 -70 806
rect -42 792 -29 830
rect 43 844 72 860
rect 86 844 115 860
rect 130 850 160 866
rect 188 844 194 892
rect 197 886 216 892
rect 231 886 261 894
rect 197 878 261 886
rect 197 862 277 878
rect 293 871 355 902
rect 371 871 433 902
rect 502 900 551 925
rect 596 916 622 926
rect 566 900 622 916
rect 465 886 495 894
rect 502 892 612 900
rect 465 878 510 886
rect 197 860 216 862
rect 231 860 277 862
rect 197 844 277 860
rect 304 858 339 871
rect 380 868 417 871
rect 380 866 422 868
rect 309 855 339 858
rect 318 851 325 855
rect 325 850 326 851
rect 284 844 294 850
rect 43 836 78 844
rect 43 810 44 836
rect 51 810 78 836
rect -14 792 16 806
rect 43 802 78 810
rect 80 836 121 844
rect 80 810 95 836
rect 102 810 121 836
rect 185 832 216 844
rect 231 832 334 844
rect 346 834 372 860
rect 387 855 417 866
rect 449 862 511 878
rect 449 860 495 862
rect 449 844 511 860
rect 523 844 529 892
rect 532 884 612 892
rect 532 882 551 884
rect 566 882 600 884
rect 532 866 612 882
rect 532 844 551 866
rect 566 850 596 866
rect 624 860 630 934
rect 633 860 652 1004
rect 667 860 673 1004
rect 682 934 695 1004
rect 747 1000 769 1004
rect 740 988 757 992
rect 761 990 769 992
rect 759 988 769 990
rect 740 978 769 988
rect 822 978 838 992
rect 876 988 882 990
rect 889 988 997 1004
rect 1004 988 1010 990
rect 1018 988 1033 1004
rect 1099 998 1118 1001
rect 740 976 838 978
rect 865 976 1033 988
rect 1048 978 1064 992
rect 1099 979 1121 998
rect 1131 992 1147 993
rect 1130 990 1147 992
rect 1131 985 1147 990
rect 1121 978 1127 979
rect 1130 978 1159 985
rect 1048 977 1159 978
rect 1048 976 1165 977
rect 724 968 775 976
rect 822 968 856 976
rect 724 956 749 968
rect 756 956 775 968
rect 829 966 856 968
rect 865 966 1086 976
rect 1121 973 1127 976
rect 829 962 1086 966
rect 724 948 775 956
rect 822 948 1086 962
rect 1130 968 1165 976
rect 676 900 695 934
rect 740 940 769 948
rect 740 934 757 940
rect 740 932 774 934
rect 822 932 838 948
rect 839 938 1047 948
rect 1048 938 1064 948
rect 1112 944 1127 959
rect 1130 956 1131 968
rect 1138 956 1165 968
rect 1130 948 1165 956
rect 1130 947 1159 948
rect 850 934 1064 938
rect 865 932 1064 934
rect 1099 934 1112 944
rect 1130 934 1147 947
rect 1099 932 1147 934
rect 741 928 774 932
rect 737 926 774 928
rect 737 925 804 926
rect 737 920 768 925
rect 774 920 804 925
rect 737 916 804 920
rect 710 913 804 916
rect 710 906 759 913
rect 710 900 740 906
rect 759 901 764 906
rect 676 884 756 900
rect 768 892 804 913
rect 865 908 1054 932
rect 1099 931 1146 932
rect 1112 926 1146 931
rect 880 905 1054 908
rect 873 902 1054 905
rect 1082 925 1146 926
rect 676 882 695 884
rect 710 882 744 884
rect 676 866 756 882
rect 676 860 695 866
rect 392 834 495 844
rect 346 832 495 834
rect 516 832 551 844
rect 185 830 347 832
rect 197 812 216 830
rect 231 828 261 830
rect 80 802 121 810
rect 204 806 216 812
rect 268 812 347 830
rect 379 830 551 832
rect 379 814 458 830
rect 465 828 495 830
rect 354 812 458 814
rect 43 792 72 802
rect 86 792 115 802
rect 130 792 160 806
rect 204 792 246 806
rect 268 802 458 812
rect 523 810 529 830
rect 253 792 283 802
rect 284 792 442 802
rect 446 792 476 802
rect 480 792 510 806
rect 538 792 551 830
rect 623 844 652 860
rect 666 844 695 860
rect 710 850 740 866
rect 768 844 774 892
rect 777 886 796 892
rect 811 886 841 894
rect 777 878 841 886
rect 777 862 857 878
rect 873 871 935 902
rect 951 871 1013 902
rect 1082 900 1131 925
rect 1146 900 1176 918
rect 1045 886 1075 894
rect 1082 892 1192 900
rect 1045 878 1090 886
rect 777 860 796 862
rect 811 860 857 862
rect 777 844 857 860
rect 884 858 919 871
rect 960 868 997 871
rect 960 866 1002 868
rect 889 855 919 858
rect 898 851 905 855
rect 905 850 906 851
rect 864 844 874 850
rect 623 836 658 844
rect 623 810 624 836
rect 631 810 658 836
rect 566 792 596 806
rect 623 802 658 810
rect 660 836 701 844
rect 660 810 675 836
rect 682 810 701 836
rect 765 832 796 844
rect 811 832 914 844
rect 926 834 952 860
rect 967 855 997 866
rect 1029 862 1091 878
rect 1029 860 1075 862
rect 1029 844 1091 860
rect 1103 844 1109 892
rect 1112 884 1192 892
rect 1112 882 1131 884
rect 1146 882 1180 884
rect 1112 867 1192 882
rect 1112 866 1198 867
rect 1112 844 1131 866
rect 1146 850 1176 866
rect 1204 860 1210 934
rect 1213 860 1232 1004
rect 1247 860 1253 1004
rect 1262 934 1275 1004
rect 1327 1000 1349 1004
rect 1320 988 1337 992
rect 1341 990 1349 992
rect 1339 988 1349 990
rect 1320 978 1349 988
rect 1402 978 1418 992
rect 1456 988 1462 990
rect 1469 988 1577 1004
rect 1584 988 1590 990
rect 1598 988 1613 1004
rect 1679 998 1698 1001
rect 1320 976 1418 978
rect 1445 976 1613 988
rect 1628 978 1644 992
rect 1679 979 1701 998
rect 1711 992 1727 993
rect 1710 990 1727 992
rect 1711 985 1727 990
rect 1701 978 1707 979
rect 1710 978 1739 985
rect 1628 977 1739 978
rect 1628 976 1745 977
rect 1304 968 1355 976
rect 1402 968 1436 976
rect 1304 956 1329 968
rect 1336 956 1355 968
rect 1409 966 1436 968
rect 1445 966 1666 976
rect 1701 973 1707 976
rect 1409 962 1666 966
rect 1304 948 1355 956
rect 1402 948 1666 962
rect 1710 968 1745 976
rect 1256 900 1275 934
rect 1320 940 1349 948
rect 1320 934 1337 940
rect 1320 932 1354 934
rect 1402 932 1418 948
rect 1419 938 1627 948
rect 1628 938 1644 948
rect 1692 944 1707 959
rect 1710 956 1711 968
rect 1718 956 1745 968
rect 1710 948 1745 956
rect 1710 947 1739 948
rect 1430 934 1644 938
rect 1445 932 1644 934
rect 1679 934 1692 944
rect 1710 934 1727 947
rect 1679 932 1727 934
rect 1321 928 1354 932
rect 1317 926 1354 928
rect 1317 925 1384 926
rect 1317 920 1348 925
rect 1354 920 1384 925
rect 1317 916 1384 920
rect 1290 913 1384 916
rect 1290 906 1339 913
rect 1290 900 1320 906
rect 1339 901 1344 906
rect 1256 884 1336 900
rect 1348 892 1384 913
rect 1445 908 1634 932
rect 1679 931 1726 932
rect 1692 926 1726 931
rect 1766 926 1782 928
rect 1460 905 1634 908
rect 1453 902 1634 905
rect 1662 925 1726 926
rect 1256 882 1275 884
rect 1290 882 1324 884
rect 1256 866 1336 882
rect 1256 860 1275 866
rect 972 834 1075 844
rect 926 832 1075 834
rect 1096 832 1131 844
rect 765 830 927 832
rect 777 812 796 830
rect 811 828 841 830
rect 660 802 701 810
rect 784 806 796 812
rect 848 812 927 830
rect 959 830 1131 832
rect 959 814 1038 830
rect 1045 828 1075 830
rect 934 812 1038 814
rect 623 792 652 802
rect 666 792 695 802
rect 710 792 740 806
rect 784 792 826 806
rect 848 802 1038 812
rect 1103 810 1109 830
rect 833 792 863 802
rect 864 792 1022 802
rect 1026 792 1056 802
rect 1060 792 1090 806
rect 1118 792 1131 830
rect 1203 844 1232 860
rect 1246 844 1275 860
rect 1290 850 1320 866
rect 1348 844 1354 892
rect 1357 886 1376 892
rect 1391 886 1421 894
rect 1357 878 1421 886
rect 1357 862 1437 878
rect 1453 871 1515 902
rect 1531 871 1593 902
rect 1662 900 1711 925
rect 1756 916 1782 926
rect 1726 900 1782 916
rect 1625 886 1655 894
rect 1662 892 1772 900
rect 1625 878 1670 886
rect 1357 860 1376 862
rect 1391 860 1437 862
rect 1357 844 1437 860
rect 1464 858 1499 871
rect 1540 868 1577 871
rect 1540 866 1582 868
rect 1469 855 1499 858
rect 1478 851 1485 855
rect 1485 850 1486 851
rect 1444 844 1454 850
rect 1203 836 1238 844
rect 1203 810 1204 836
rect 1211 810 1238 836
rect 1146 792 1176 806
rect 1203 802 1238 810
rect 1240 836 1281 844
rect 1240 810 1255 836
rect 1262 810 1281 836
rect 1345 832 1376 844
rect 1391 832 1494 844
rect 1506 834 1532 860
rect 1547 855 1577 866
rect 1609 862 1671 878
rect 1609 860 1655 862
rect 1609 844 1671 860
rect 1683 844 1689 892
rect 1692 884 1772 892
rect 1692 882 1711 884
rect 1726 882 1760 884
rect 1692 866 1772 882
rect 1692 844 1711 866
rect 1726 850 1756 866
rect 1784 860 1790 934
rect 1793 860 1812 1004
rect 1827 860 1833 1004
rect 1842 934 1855 1004
rect 1907 1000 1929 1004
rect 1900 988 1917 992
rect 1921 990 1929 992
rect 1919 988 1929 990
rect 1900 978 1929 988
rect 1982 978 1998 992
rect 2036 988 2042 990
rect 2049 988 2157 1004
rect 2164 988 2170 990
rect 2178 988 2193 1004
rect 2259 998 2278 1001
rect 1900 976 1998 978
rect 2025 976 2193 988
rect 2208 978 2224 992
rect 2259 979 2281 998
rect 2291 992 2307 993
rect 2290 990 2307 992
rect 2291 985 2307 990
rect 2281 978 2287 979
rect 2290 978 2319 985
rect 2208 977 2319 978
rect 2208 976 2325 977
rect 1884 968 1935 976
rect 1982 968 2016 976
rect 1884 956 1909 968
rect 1916 956 1935 968
rect 1989 966 2016 968
rect 2025 966 2246 976
rect 2281 973 2287 976
rect 1989 962 2246 966
rect 1884 948 1935 956
rect 1982 948 2246 962
rect 2290 968 2325 976
rect 1836 900 1855 934
rect 1900 940 1929 948
rect 1900 934 1917 940
rect 1900 932 1934 934
rect 1982 932 1998 948
rect 1999 938 2207 948
rect 2208 938 2224 948
rect 2272 944 2287 959
rect 2290 956 2291 968
rect 2298 956 2325 968
rect 2290 948 2325 956
rect 2290 947 2319 948
rect 2010 934 2224 938
rect 2025 932 2224 934
rect 2259 934 2272 944
rect 2290 934 2307 947
rect 2259 932 2307 934
rect 1901 928 1934 932
rect 1897 926 1934 928
rect 1897 925 1964 926
rect 1897 920 1928 925
rect 1934 920 1964 925
rect 1897 916 1964 920
rect 1870 913 1964 916
rect 1870 906 1919 913
rect 1870 900 1900 906
rect 1919 901 1924 906
rect 1836 884 1916 900
rect 1928 892 1964 913
rect 2025 908 2214 932
rect 2259 931 2306 932
rect 2272 926 2306 931
rect 2040 905 2214 908
rect 2033 902 2214 905
rect 2242 925 2306 926
rect 1836 882 1855 884
rect 1870 882 1904 884
rect 1836 866 1916 882
rect 1836 860 1855 866
rect 1552 834 1655 844
rect 1506 832 1655 834
rect 1676 832 1711 844
rect 1345 830 1507 832
rect 1357 812 1376 830
rect 1391 828 1421 830
rect 1240 802 1281 810
rect 1364 806 1376 812
rect 1428 812 1507 830
rect 1539 830 1711 832
rect 1539 814 1618 830
rect 1625 828 1655 830
rect 1514 812 1618 814
rect 1203 792 1232 802
rect 1246 792 1275 802
rect 1290 792 1320 806
rect 1364 792 1406 806
rect 1428 802 1618 812
rect 1683 810 1689 830
rect 1413 792 1443 802
rect 1444 792 1602 802
rect 1606 792 1636 802
rect 1640 792 1670 806
rect 1698 792 1711 830
rect 1783 844 1812 860
rect 1826 844 1855 860
rect 1870 850 1900 866
rect 1928 844 1934 892
rect 1937 886 1956 892
rect 1971 886 2001 894
rect 1937 878 2001 886
rect 1937 862 2017 878
rect 2033 871 2095 902
rect 2111 871 2173 902
rect 2242 900 2291 925
rect 2306 900 2336 918
rect 2205 886 2235 894
rect 2242 892 2352 900
rect 2205 878 2250 886
rect 1937 860 1956 862
rect 1971 860 2017 862
rect 1937 844 2017 860
rect 2044 858 2079 871
rect 2120 868 2157 871
rect 2120 866 2162 868
rect 2049 855 2079 858
rect 2058 851 2065 855
rect 2065 850 2066 851
rect 2024 844 2034 850
rect 1783 836 1818 844
rect 1783 810 1784 836
rect 1791 810 1818 836
rect 1726 792 1756 806
rect 1783 802 1818 810
rect 1820 836 1861 844
rect 1820 810 1835 836
rect 1842 810 1861 836
rect 1925 832 1956 844
rect 1971 832 2074 844
rect 2086 834 2112 860
rect 2127 855 2157 866
rect 2189 862 2251 878
rect 2189 860 2235 862
rect 2189 844 2251 860
rect 2263 844 2269 892
rect 2272 884 2352 892
rect 2272 882 2291 884
rect 2306 882 2340 884
rect 2272 867 2352 882
rect 2272 866 2358 867
rect 2272 844 2291 866
rect 2306 850 2336 866
rect 2364 860 2370 934
rect 2373 860 2392 1004
rect 2407 860 2413 1004
rect 2422 934 2435 1004
rect 2487 1000 2509 1004
rect 2480 988 2497 992
rect 2501 990 2509 992
rect 2499 988 2509 990
rect 2480 978 2509 988
rect 2562 978 2578 992
rect 2616 988 2622 990
rect 2629 988 2737 1004
rect 2744 988 2750 990
rect 2758 988 2773 1004
rect 2839 998 2858 1001
rect 2480 976 2578 978
rect 2605 976 2773 988
rect 2788 978 2804 992
rect 2839 979 2861 998
rect 2871 992 2887 993
rect 2870 990 2887 992
rect 2871 985 2887 990
rect 2861 978 2867 979
rect 2870 978 2899 985
rect 2788 977 2899 978
rect 2788 976 2905 977
rect 2464 968 2515 976
rect 2562 968 2596 976
rect 2464 956 2489 968
rect 2496 956 2515 968
rect 2569 966 2596 968
rect 2605 966 2826 976
rect 2861 973 2867 976
rect 2569 962 2826 966
rect 2464 948 2515 956
rect 2562 948 2826 962
rect 2870 968 2905 976
rect 2416 900 2435 934
rect 2480 940 2509 948
rect 2480 934 2497 940
rect 2480 932 2514 934
rect 2562 932 2578 948
rect 2579 938 2787 948
rect 2788 938 2804 948
rect 2852 944 2867 959
rect 2870 956 2871 968
rect 2878 956 2905 968
rect 2870 948 2905 956
rect 2870 947 2899 948
rect 2590 934 2804 938
rect 2605 932 2804 934
rect 2839 934 2852 944
rect 2870 934 2887 947
rect 2839 932 2887 934
rect 2481 928 2514 932
rect 2477 926 2514 928
rect 2477 925 2544 926
rect 2477 920 2508 925
rect 2514 920 2544 925
rect 2477 916 2544 920
rect 2450 913 2544 916
rect 2450 906 2499 913
rect 2450 900 2480 906
rect 2499 901 2504 906
rect 2416 884 2496 900
rect 2508 892 2544 913
rect 2605 908 2794 932
rect 2839 931 2886 932
rect 2852 926 2886 931
rect 2926 926 2942 928
rect 2620 905 2794 908
rect 2613 902 2794 905
rect 2822 925 2886 926
rect 2416 882 2435 884
rect 2450 882 2484 884
rect 2416 866 2496 882
rect 2416 860 2435 866
rect 2132 834 2235 844
rect 2086 832 2235 834
rect 2256 832 2291 844
rect 1925 830 2087 832
rect 1937 812 1956 830
rect 1971 828 2001 830
rect 1820 802 1861 810
rect 1944 806 1956 812
rect 2008 812 2087 830
rect 2119 830 2291 832
rect 2119 814 2198 830
rect 2205 828 2235 830
rect 2094 812 2198 814
rect 1783 792 1812 802
rect 1826 792 1855 802
rect 1870 792 1900 806
rect 1944 792 1986 806
rect 2008 802 2198 812
rect 2263 810 2269 830
rect 1993 792 2023 802
rect 2024 792 2182 802
rect 2186 792 2216 802
rect 2220 792 2250 806
rect 2278 792 2291 830
rect 2363 844 2392 860
rect 2406 844 2435 860
rect 2450 850 2480 866
rect 2508 844 2514 892
rect 2517 886 2536 892
rect 2551 886 2581 894
rect 2517 878 2581 886
rect 2517 862 2597 878
rect 2613 871 2675 902
rect 2691 871 2753 902
rect 2822 900 2871 925
rect 2916 916 2942 926
rect 2886 900 2942 916
rect 2785 886 2815 894
rect 2822 892 2932 900
rect 2785 878 2830 886
rect 2517 860 2536 862
rect 2551 860 2597 862
rect 2517 844 2597 860
rect 2624 858 2659 871
rect 2700 868 2737 871
rect 2700 866 2742 868
rect 2629 855 2659 858
rect 2638 851 2645 855
rect 2645 850 2646 851
rect 2604 844 2614 850
rect 2363 836 2398 844
rect 2363 810 2364 836
rect 2371 810 2398 836
rect 2306 792 2336 806
rect 2363 802 2398 810
rect 2400 836 2441 844
rect 2400 810 2415 836
rect 2422 810 2441 836
rect 2505 832 2536 844
rect 2551 832 2654 844
rect 2666 834 2692 860
rect 2707 855 2737 866
rect 2769 862 2831 878
rect 2769 860 2815 862
rect 2769 844 2831 860
rect 2843 844 2849 892
rect 2852 884 2932 892
rect 2852 882 2871 884
rect 2886 882 2920 884
rect 2852 866 2932 882
rect 2852 844 2871 866
rect 2886 850 2916 866
rect 2944 860 2950 934
rect 2953 860 2972 1004
rect 2987 860 2993 1004
rect 3002 934 3015 1004
rect 3067 1000 3089 1004
rect 3060 988 3077 992
rect 3081 990 3089 992
rect 3079 988 3089 990
rect 3060 978 3089 988
rect 3142 978 3158 992
rect 3196 988 3202 990
rect 3209 988 3317 1004
rect 3324 988 3330 990
rect 3338 988 3353 1004
rect 3419 998 3438 1001
rect 3060 976 3158 978
rect 3185 976 3353 988
rect 3368 978 3384 992
rect 3419 979 3441 998
rect 3451 992 3467 993
rect 3450 990 3467 992
rect 3451 985 3467 990
rect 3441 978 3447 979
rect 3450 978 3479 985
rect 3368 977 3479 978
rect 3368 976 3485 977
rect 3044 968 3095 976
rect 3142 968 3176 976
rect 3044 956 3069 968
rect 3076 956 3095 968
rect 3149 966 3176 968
rect 3185 966 3406 976
rect 3441 973 3447 976
rect 3149 962 3406 966
rect 3044 948 3095 956
rect 3142 948 3406 962
rect 3450 968 3485 976
rect 2996 900 3015 934
rect 3060 940 3089 948
rect 3060 934 3077 940
rect 3060 932 3094 934
rect 3142 932 3158 948
rect 3159 938 3367 948
rect 3368 938 3384 948
rect 3432 944 3447 959
rect 3450 956 3451 968
rect 3458 956 3485 968
rect 3450 948 3485 956
rect 3450 947 3479 948
rect 3170 934 3384 938
rect 3185 932 3384 934
rect 3419 934 3432 944
rect 3450 934 3467 947
rect 3419 932 3467 934
rect 3061 928 3094 932
rect 3057 926 3094 928
rect 3057 925 3124 926
rect 3057 920 3088 925
rect 3094 920 3124 925
rect 3057 916 3124 920
rect 3030 913 3124 916
rect 3030 906 3079 913
rect 3030 900 3060 906
rect 3079 901 3084 906
rect 2996 884 3076 900
rect 3088 892 3124 913
rect 3185 908 3374 932
rect 3419 931 3466 932
rect 3432 926 3466 931
rect 3200 905 3374 908
rect 3193 902 3374 905
rect 3402 925 3466 926
rect 2996 882 3015 884
rect 3030 882 3064 884
rect 2996 866 3076 882
rect 2996 860 3015 866
rect 2712 834 2815 844
rect 2666 832 2815 834
rect 2836 832 2871 844
rect 2505 830 2667 832
rect 2517 812 2536 830
rect 2551 828 2581 830
rect 2400 802 2441 810
rect 2524 806 2536 812
rect 2588 812 2667 830
rect 2699 830 2871 832
rect 2699 814 2778 830
rect 2785 828 2815 830
rect 2674 812 2778 814
rect 2363 792 2392 802
rect 2406 792 2435 802
rect 2450 792 2480 806
rect 2524 792 2566 806
rect 2588 802 2778 812
rect 2843 810 2849 830
rect 2573 792 2603 802
rect 2604 792 2762 802
rect 2766 792 2796 802
rect 2800 792 2830 806
rect 2858 792 2871 830
rect 2943 844 2972 860
rect 2986 844 3015 860
rect 3030 850 3060 866
rect 3088 844 3094 892
rect 3097 886 3116 892
rect 3131 886 3161 894
rect 3097 878 3161 886
rect 3097 862 3177 878
rect 3193 871 3255 902
rect 3271 871 3333 902
rect 3402 900 3451 925
rect 3466 900 3496 918
rect 3365 886 3395 894
rect 3402 892 3512 900
rect 3365 878 3410 886
rect 3097 860 3116 862
rect 3131 860 3177 862
rect 3097 844 3177 860
rect 3204 858 3239 871
rect 3280 868 3317 871
rect 3280 866 3322 868
rect 3209 855 3239 858
rect 3218 851 3225 855
rect 3225 850 3226 851
rect 3184 844 3194 850
rect 2943 836 2978 844
rect 2943 810 2944 836
rect 2951 810 2978 836
rect 2886 792 2916 806
rect 2943 802 2978 810
rect 2980 836 3021 844
rect 2980 810 2995 836
rect 3002 810 3021 836
rect 3085 832 3116 844
rect 3131 832 3234 844
rect 3246 834 3272 860
rect 3287 855 3317 866
rect 3349 862 3411 878
rect 3349 860 3395 862
rect 3349 844 3411 860
rect 3423 844 3429 892
rect 3432 884 3512 892
rect 3432 882 3451 884
rect 3466 882 3500 884
rect 3432 867 3512 882
rect 3432 866 3518 867
rect 3432 844 3451 866
rect 3466 850 3496 866
rect 3524 860 3530 934
rect 3533 860 3552 1004
rect 3567 860 3573 1004
rect 3582 934 3595 1004
rect 3647 1000 3669 1004
rect 3640 988 3657 992
rect 3661 990 3669 992
rect 3659 988 3669 990
rect 3640 978 3669 988
rect 3722 978 3738 992
rect 3776 988 3782 990
rect 3789 988 3897 1004
rect 3904 988 3910 990
rect 3918 988 3933 1004
rect 3999 998 4018 1001
rect 3640 976 3738 978
rect 3765 976 3933 988
rect 3948 978 3964 992
rect 3999 979 4021 998
rect 4031 992 4047 993
rect 4030 990 4047 992
rect 4031 985 4047 990
rect 4021 978 4027 979
rect 4030 978 4059 985
rect 3948 977 4059 978
rect 3948 976 4065 977
rect 3624 968 3675 976
rect 3722 968 3756 976
rect 3624 956 3649 968
rect 3656 956 3675 968
rect 3729 966 3756 968
rect 3765 966 3986 976
rect 4021 973 4027 976
rect 3729 962 3986 966
rect 3624 948 3675 956
rect 3722 948 3986 962
rect 4030 968 4065 976
rect 3576 900 3595 934
rect 3640 940 3669 948
rect 3640 934 3657 940
rect 3640 932 3674 934
rect 3722 932 3738 948
rect 3739 938 3947 948
rect 3948 938 3964 948
rect 4012 944 4027 959
rect 4030 956 4031 968
rect 4038 956 4065 968
rect 4030 948 4065 956
rect 4030 947 4059 948
rect 3750 934 3964 938
rect 3765 932 3964 934
rect 3999 934 4012 944
rect 4030 934 4047 947
rect 3999 932 4047 934
rect 3641 928 3674 932
rect 3637 926 3674 928
rect 3637 925 3704 926
rect 3637 920 3668 925
rect 3674 920 3704 925
rect 3637 916 3704 920
rect 3610 913 3704 916
rect 3610 906 3659 913
rect 3610 900 3640 906
rect 3659 901 3664 906
rect 3576 884 3656 900
rect 3668 892 3704 913
rect 3765 908 3954 932
rect 3999 931 4046 932
rect 4012 926 4046 931
rect 4086 926 4102 928
rect 3780 905 3954 908
rect 3773 902 3954 905
rect 3982 925 4046 926
rect 3576 882 3595 884
rect 3610 882 3644 884
rect 3576 866 3656 882
rect 3576 860 3595 866
rect 3292 834 3395 844
rect 3246 832 3395 834
rect 3416 832 3451 844
rect 3085 830 3247 832
rect 3097 812 3116 830
rect 3131 828 3161 830
rect 2980 802 3021 810
rect 3104 806 3116 812
rect 3168 812 3247 830
rect 3279 830 3451 832
rect 3279 814 3358 830
rect 3365 828 3395 830
rect 3254 812 3358 814
rect 2943 792 2972 802
rect 2986 792 3015 802
rect 3030 792 3060 806
rect 3104 792 3146 806
rect 3168 802 3358 812
rect 3423 810 3429 830
rect 3153 792 3183 802
rect 3184 792 3342 802
rect 3346 792 3376 802
rect 3380 792 3410 806
rect 3438 792 3451 830
rect 3523 844 3552 860
rect 3566 844 3595 860
rect 3610 850 3640 866
rect 3668 844 3674 892
rect 3677 886 3696 892
rect 3711 886 3741 894
rect 3677 878 3741 886
rect 3677 862 3757 878
rect 3773 871 3835 902
rect 3851 871 3913 902
rect 3982 900 4031 925
rect 4076 916 4102 926
rect 4046 900 4102 916
rect 3945 886 3975 894
rect 3982 892 4092 900
rect 3945 878 3990 886
rect 3677 860 3696 862
rect 3711 860 3757 862
rect 3677 844 3757 860
rect 3784 858 3819 871
rect 3860 868 3897 871
rect 3860 866 3902 868
rect 3789 855 3819 858
rect 3798 851 3805 855
rect 3805 850 3806 851
rect 3764 844 3774 850
rect 3523 836 3558 844
rect 3523 810 3524 836
rect 3531 810 3558 836
rect 3466 792 3496 806
rect 3523 802 3558 810
rect 3560 836 3601 844
rect 3560 810 3575 836
rect 3582 810 3601 836
rect 3665 832 3696 844
rect 3711 832 3814 844
rect 3826 834 3852 860
rect 3867 855 3897 866
rect 3929 862 3991 878
rect 3929 860 3975 862
rect 3929 844 3991 860
rect 4003 844 4009 892
rect 4012 884 4092 892
rect 4012 882 4031 884
rect 4046 882 4080 884
rect 4012 866 4092 882
rect 4012 844 4031 866
rect 4046 850 4076 866
rect 4104 860 4110 934
rect 4113 860 4132 1004
rect 4147 860 4153 1004
rect 4162 934 4175 1004
rect 4227 1000 4249 1004
rect 4220 988 4237 992
rect 4241 990 4249 992
rect 4239 988 4249 990
rect 4220 978 4249 988
rect 4302 978 4318 992
rect 4356 988 4362 990
rect 4369 988 4477 1004
rect 4484 988 4490 990
rect 4498 988 4513 1004
rect 4579 998 4598 1001
rect 4220 976 4318 978
rect 4345 976 4513 988
rect 4528 978 4544 992
rect 4579 979 4601 998
rect 4611 992 4627 993
rect 4610 990 4627 992
rect 4611 985 4627 990
rect 4601 978 4607 979
rect 4610 978 4639 985
rect 4528 977 4639 978
rect 4528 976 4645 977
rect 4204 968 4255 976
rect 4302 968 4336 976
rect 4204 956 4229 968
rect 4236 956 4255 968
rect 4309 966 4336 968
rect 4345 966 4566 976
rect 4601 973 4607 976
rect 4309 962 4566 966
rect 4204 948 4255 956
rect 4302 948 4566 962
rect 4610 968 4645 976
rect 4156 900 4175 934
rect 4220 940 4249 948
rect 4220 934 4237 940
rect 4220 932 4254 934
rect 4302 932 4318 948
rect 4319 938 4527 948
rect 4528 938 4544 948
rect 4592 944 4607 959
rect 4610 956 4611 968
rect 4618 956 4645 968
rect 4610 948 4645 956
rect 4610 947 4639 948
rect 4330 934 4544 938
rect 4345 932 4544 934
rect 4579 934 4592 944
rect 4610 934 4627 947
rect 4579 932 4627 934
rect 4221 928 4254 932
rect 4217 926 4254 928
rect 4217 925 4284 926
rect 4217 920 4248 925
rect 4254 920 4284 925
rect 4217 916 4284 920
rect 4190 913 4284 916
rect 4190 906 4239 913
rect 4190 900 4220 906
rect 4239 901 4244 906
rect 4156 884 4236 900
rect 4248 892 4284 913
rect 4345 908 4534 932
rect 4579 931 4626 932
rect 4592 926 4626 931
rect 4360 905 4534 908
rect 4353 902 4534 905
rect 4562 925 4626 926
rect 4156 882 4175 884
rect 4190 882 4224 884
rect 4156 866 4236 882
rect 4156 860 4175 866
rect 3872 834 3975 844
rect 3826 832 3975 834
rect 3996 832 4031 844
rect 3665 830 3827 832
rect 3677 812 3696 830
rect 3711 828 3741 830
rect 3560 802 3601 810
rect 3684 806 3696 812
rect 3748 812 3827 830
rect 3859 830 4031 832
rect 3859 814 3938 830
rect 3945 828 3975 830
rect 3834 812 3938 814
rect 3523 792 3552 802
rect 3566 792 3595 802
rect 3610 792 3640 806
rect 3684 792 3726 806
rect 3748 802 3938 812
rect 4003 810 4009 830
rect 3733 792 3763 802
rect 3764 792 3922 802
rect 3926 792 3956 802
rect 3960 792 3990 806
rect 4018 792 4031 830
rect 4103 844 4132 860
rect 4146 844 4175 860
rect 4190 850 4220 866
rect 4248 844 4254 892
rect 4257 886 4276 892
rect 4291 886 4321 894
rect 4257 878 4321 886
rect 4257 862 4337 878
rect 4353 871 4415 902
rect 4431 871 4493 902
rect 4562 900 4611 925
rect 4626 900 4656 918
rect 4525 886 4555 894
rect 4562 892 4672 900
rect 4525 878 4570 886
rect 4257 860 4276 862
rect 4291 860 4337 862
rect 4257 844 4337 860
rect 4364 858 4399 871
rect 4440 868 4477 871
rect 4440 866 4482 868
rect 4369 855 4399 858
rect 4378 851 4385 855
rect 4385 850 4386 851
rect 4344 844 4354 850
rect 4103 836 4138 844
rect 4103 810 4104 836
rect 4111 810 4138 836
rect 4046 792 4076 806
rect 4103 802 4138 810
rect 4140 836 4181 844
rect 4140 810 4155 836
rect 4162 810 4181 836
rect 4245 832 4276 844
rect 4291 832 4394 844
rect 4406 834 4432 860
rect 4447 855 4477 866
rect 4509 862 4571 878
rect 4509 860 4555 862
rect 4509 844 4571 860
rect 4583 844 4589 892
rect 4592 884 4672 892
rect 4592 882 4611 884
rect 4626 882 4660 884
rect 4592 867 4672 882
rect 4592 866 4678 867
rect 4592 844 4611 866
rect 4626 850 4656 866
rect 4684 860 4690 934
rect 4693 860 4712 1004
rect 4727 860 4733 1004
rect 4742 934 4755 1004
rect 4807 1000 4829 1004
rect 4800 988 4817 992
rect 4821 990 4829 992
rect 4819 988 4829 990
rect 4800 978 4829 988
rect 4882 978 4898 992
rect 4936 988 4942 990
rect 4949 988 5057 1004
rect 5064 988 5070 990
rect 5078 988 5093 1004
rect 5159 998 5178 1001
rect 4800 976 4898 978
rect 4925 976 5093 988
rect 5108 978 5124 992
rect 5159 979 5181 998
rect 5191 992 5207 993
rect 5190 990 5207 992
rect 5191 985 5207 990
rect 5181 978 5187 979
rect 5190 978 5219 985
rect 5108 977 5219 978
rect 5108 976 5225 977
rect 4784 968 4835 976
rect 4882 968 4916 976
rect 4784 956 4809 968
rect 4816 956 4835 968
rect 4889 966 4916 968
rect 4925 966 5146 976
rect 5181 973 5187 976
rect 4889 962 5146 966
rect 4784 948 4835 956
rect 4882 948 5146 962
rect 5190 968 5225 976
rect 4736 900 4755 934
rect 4800 940 4829 948
rect 4800 934 4817 940
rect 4800 932 4834 934
rect 4882 932 4898 948
rect 4899 938 5107 948
rect 5108 938 5124 948
rect 5172 944 5187 959
rect 5190 956 5191 968
rect 5198 956 5225 968
rect 5190 948 5225 956
rect 5190 947 5219 948
rect 4910 934 5124 938
rect 4925 932 5124 934
rect 5159 934 5172 944
rect 5190 934 5207 947
rect 5159 932 5207 934
rect 4801 928 4834 932
rect 4797 926 4834 928
rect 4797 925 4864 926
rect 4797 920 4828 925
rect 4834 920 4864 925
rect 4797 916 4864 920
rect 4770 913 4864 916
rect 4770 906 4819 913
rect 4770 900 4800 906
rect 4819 901 4824 906
rect 4736 884 4816 900
rect 4828 892 4864 913
rect 4925 908 5114 932
rect 5159 931 5206 932
rect 5172 926 5206 931
rect 5246 926 5262 928
rect 4940 905 5114 908
rect 4933 902 5114 905
rect 5142 925 5206 926
rect 4736 882 4755 884
rect 4770 882 4804 884
rect 4736 866 4816 882
rect 4736 860 4755 866
rect 4452 834 4555 844
rect 4406 832 4555 834
rect 4576 832 4611 844
rect 4245 830 4407 832
rect 4257 812 4276 830
rect 4291 828 4321 830
rect 4140 802 4181 810
rect 4264 806 4276 812
rect 4328 812 4407 830
rect 4439 830 4611 832
rect 4439 814 4518 830
rect 4525 828 4555 830
rect 4414 812 4518 814
rect 4103 792 4132 802
rect 4146 792 4175 802
rect 4190 792 4220 806
rect 4264 792 4306 806
rect 4328 802 4518 812
rect 4583 810 4589 830
rect 4313 792 4343 802
rect 4344 792 4502 802
rect 4506 792 4536 802
rect 4540 792 4570 806
rect 4598 792 4611 830
rect 4683 844 4712 860
rect 4726 844 4755 860
rect 4770 850 4800 866
rect 4828 844 4834 892
rect 4837 886 4856 892
rect 4871 886 4901 894
rect 4837 878 4901 886
rect 4837 862 4917 878
rect 4933 871 4995 902
rect 5011 871 5073 902
rect 5142 900 5191 925
rect 5236 916 5262 926
rect 5206 900 5262 916
rect 5105 886 5135 894
rect 5142 892 5252 900
rect 5105 878 5150 886
rect 4837 860 4856 862
rect 4871 860 4917 862
rect 4837 844 4917 860
rect 4944 858 4979 871
rect 5020 868 5057 871
rect 5020 866 5062 868
rect 4949 855 4979 858
rect 4958 851 4965 855
rect 4965 850 4966 851
rect 4924 844 4934 850
rect 4683 836 4718 844
rect 4683 810 4684 836
rect 4691 810 4718 836
rect 4626 792 4656 806
rect 4683 802 4718 810
rect 4720 836 4761 844
rect 4720 810 4735 836
rect 4742 810 4761 836
rect 4825 832 4856 844
rect 4871 832 4974 844
rect 4986 834 5012 860
rect 5027 855 5057 866
rect 5089 862 5151 878
rect 5089 860 5135 862
rect 5089 844 5151 860
rect 5163 844 5169 892
rect 5172 884 5252 892
rect 5172 882 5191 884
rect 5206 882 5240 884
rect 5172 866 5252 882
rect 5172 844 5191 866
rect 5206 850 5236 866
rect 5264 860 5270 934
rect 5273 860 5292 1004
rect 5307 860 5313 1004
rect 5322 934 5335 1004
rect 5387 1000 5409 1004
rect 5380 988 5397 992
rect 5401 990 5409 992
rect 5399 988 5409 990
rect 5380 978 5409 988
rect 5462 978 5478 992
rect 5516 988 5522 990
rect 5529 988 5637 1004
rect 5644 988 5650 990
rect 5658 988 5673 1004
rect 5739 998 5758 1001
rect 5380 976 5478 978
rect 5505 976 5673 988
rect 5688 978 5704 992
rect 5739 979 5761 998
rect 5771 992 5787 993
rect 5770 990 5787 992
rect 5771 985 5787 990
rect 5761 978 5767 979
rect 5770 978 5799 985
rect 5688 977 5799 978
rect 5688 976 5805 977
rect 5364 968 5415 976
rect 5462 968 5496 976
rect 5364 956 5389 968
rect 5396 956 5415 968
rect 5469 966 5496 968
rect 5505 966 5726 976
rect 5761 973 5767 976
rect 5469 962 5726 966
rect 5364 948 5415 956
rect 5462 948 5726 962
rect 5770 968 5805 976
rect 5316 900 5335 934
rect 5380 940 5409 948
rect 5380 934 5397 940
rect 5380 932 5414 934
rect 5462 932 5478 948
rect 5479 938 5687 948
rect 5688 938 5704 948
rect 5752 944 5767 959
rect 5770 956 5771 968
rect 5778 956 5805 968
rect 5770 948 5805 956
rect 5770 947 5799 948
rect 5490 934 5704 938
rect 5505 932 5704 934
rect 5739 934 5752 944
rect 5770 934 5787 947
rect 5739 932 5787 934
rect 5381 928 5414 932
rect 5377 926 5414 928
rect 5377 925 5444 926
rect 5377 920 5408 925
rect 5414 920 5444 925
rect 5377 916 5444 920
rect 5350 913 5444 916
rect 5350 906 5399 913
rect 5350 900 5380 906
rect 5399 901 5404 906
rect 5316 884 5396 900
rect 5408 892 5444 913
rect 5505 908 5694 932
rect 5739 931 5786 932
rect 5752 926 5786 931
rect 5520 905 5694 908
rect 5513 902 5694 905
rect 5722 925 5786 926
rect 5316 882 5335 884
rect 5350 882 5384 884
rect 5316 866 5396 882
rect 5316 860 5335 866
rect 5032 834 5135 844
rect 4986 832 5135 834
rect 5156 832 5191 844
rect 4825 830 4987 832
rect 4837 812 4856 830
rect 4871 828 4901 830
rect 4720 802 4761 810
rect 4844 806 4856 812
rect 4908 812 4987 830
rect 5019 830 5191 832
rect 5019 814 5098 830
rect 5105 828 5135 830
rect 4994 812 5098 814
rect 4683 792 4712 802
rect 4726 792 4755 802
rect 4770 792 4800 806
rect 4844 792 4886 806
rect 4908 802 5098 812
rect 5163 810 5169 830
rect 4893 792 4923 802
rect 4924 792 5082 802
rect 5086 792 5116 802
rect 5120 792 5150 806
rect 5178 792 5191 830
rect 5263 844 5292 860
rect 5306 844 5335 860
rect 5350 850 5380 866
rect 5408 844 5414 892
rect 5417 886 5436 892
rect 5451 886 5481 894
rect 5417 878 5481 886
rect 5417 862 5497 878
rect 5513 871 5575 902
rect 5591 871 5653 902
rect 5722 900 5771 925
rect 5786 900 5816 918
rect 5685 886 5715 894
rect 5722 892 5832 900
rect 5685 878 5730 886
rect 5417 860 5436 862
rect 5451 860 5497 862
rect 5417 844 5497 860
rect 5524 858 5559 871
rect 5600 868 5637 871
rect 5600 866 5642 868
rect 5529 855 5559 858
rect 5538 851 5545 855
rect 5545 850 5546 851
rect 5504 844 5514 850
rect 5263 836 5298 844
rect 5263 810 5264 836
rect 5271 810 5298 836
rect 5206 792 5236 806
rect 5263 802 5298 810
rect 5300 836 5341 844
rect 5300 810 5315 836
rect 5322 810 5341 836
rect 5405 832 5436 844
rect 5451 832 5554 844
rect 5566 834 5592 860
rect 5607 855 5637 866
rect 5669 862 5731 878
rect 5669 860 5715 862
rect 5669 844 5731 860
rect 5743 844 5749 892
rect 5752 884 5832 892
rect 5752 882 5771 884
rect 5786 882 5820 884
rect 5752 867 5832 882
rect 5752 866 5838 867
rect 5752 844 5771 866
rect 5786 850 5816 866
rect 5844 860 5850 934
rect 5853 860 5872 1004
rect 5887 860 5893 1004
rect 5902 934 5915 1004
rect 5967 1000 5989 1004
rect 5960 988 5977 992
rect 5981 990 5989 992
rect 5979 988 5989 990
rect 5960 978 5989 988
rect 6042 978 6058 992
rect 6096 988 6102 990
rect 6109 988 6217 1004
rect 6224 988 6230 990
rect 6238 988 6253 1004
rect 6319 998 6338 1001
rect 5960 976 6058 978
rect 6085 976 6253 988
rect 6268 978 6284 992
rect 6319 979 6341 998
rect 6351 992 6367 993
rect 6350 990 6367 992
rect 6351 985 6367 990
rect 6341 978 6347 979
rect 6350 978 6379 985
rect 6268 977 6379 978
rect 6268 976 6385 977
rect 5944 968 5995 976
rect 6042 968 6076 976
rect 5944 956 5969 968
rect 5976 956 5995 968
rect 6049 966 6076 968
rect 6085 966 6306 976
rect 6341 973 6347 976
rect 6049 962 6306 966
rect 5944 948 5995 956
rect 6042 948 6306 962
rect 6350 968 6385 976
rect 5896 900 5915 934
rect 5960 940 5989 948
rect 5960 934 5977 940
rect 5960 932 5994 934
rect 6042 932 6058 948
rect 6059 938 6267 948
rect 6268 938 6284 948
rect 6332 944 6347 959
rect 6350 956 6351 968
rect 6358 956 6385 968
rect 6350 948 6385 956
rect 6350 947 6379 948
rect 6070 934 6284 938
rect 6085 932 6284 934
rect 6319 934 6332 944
rect 6350 934 6367 947
rect 6319 932 6367 934
rect 5961 928 5994 932
rect 5957 926 5994 928
rect 5957 925 6024 926
rect 5957 920 5988 925
rect 5994 920 6024 925
rect 5957 916 6024 920
rect 5930 913 6024 916
rect 5930 906 5979 913
rect 5930 900 5960 906
rect 5979 901 5984 906
rect 5896 884 5976 900
rect 5988 892 6024 913
rect 6085 908 6274 932
rect 6319 931 6366 932
rect 6332 926 6366 931
rect 6100 905 6274 908
rect 6093 902 6274 905
rect 6302 925 6366 926
rect 5896 882 5915 884
rect 5930 882 5964 884
rect 5896 866 5976 882
rect 5896 860 5915 866
rect 5612 834 5715 844
rect 5566 832 5715 834
rect 5736 832 5771 844
rect 5405 830 5567 832
rect 5417 812 5436 830
rect 5451 828 5481 830
rect 5300 802 5341 810
rect 5424 806 5436 812
rect 5488 812 5567 830
rect 5599 830 5771 832
rect 5599 814 5678 830
rect 5685 828 5715 830
rect 5574 812 5678 814
rect 5263 792 5292 802
rect 5306 792 5335 802
rect 5350 792 5380 806
rect 5424 792 5466 806
rect 5488 802 5678 812
rect 5743 810 5749 830
rect 5473 792 5503 802
rect 5504 792 5662 802
rect 5666 792 5696 802
rect 5700 792 5730 806
rect 5758 792 5771 830
rect 5843 844 5872 860
rect 5886 844 5915 860
rect 5930 850 5960 866
rect 5988 844 5994 892
rect 5997 886 6016 892
rect 6031 886 6061 894
rect 5997 878 6061 886
rect 5997 862 6077 878
rect 6093 871 6155 902
rect 6171 871 6233 902
rect 6302 900 6351 925
rect 6366 900 6396 916
rect 6265 886 6295 894
rect 6302 892 6412 900
rect 6265 878 6310 886
rect 5997 860 6016 862
rect 6031 860 6077 862
rect 5997 844 6077 860
rect 6104 858 6139 871
rect 6180 868 6217 871
rect 6180 866 6222 868
rect 6109 855 6139 858
rect 6118 851 6125 855
rect 6125 850 6126 851
rect 6084 844 6094 850
rect 5843 836 5878 844
rect 5843 810 5844 836
rect 5851 810 5878 836
rect 5786 792 5816 806
rect 5843 802 5878 810
rect 5880 836 5921 844
rect 5880 810 5895 836
rect 5902 810 5921 836
rect 5985 832 6016 844
rect 6031 832 6134 844
rect 6146 834 6172 860
rect 6187 855 6217 866
rect 6249 862 6311 878
rect 6249 860 6295 862
rect 6249 844 6311 860
rect 6323 844 6329 892
rect 6332 884 6412 892
rect 6332 882 6351 884
rect 6366 882 6400 884
rect 6332 866 6412 882
rect 6332 844 6351 866
rect 6366 850 6396 866
rect 6424 860 6430 934
rect 6439 860 6452 1004
rect 6192 834 6295 844
rect 6146 832 6295 834
rect 6316 832 6351 844
rect 5985 830 6147 832
rect 5997 812 6016 830
rect 6031 828 6061 830
rect 5880 802 5921 810
rect 6004 806 6016 812
rect 6068 812 6147 830
rect 6179 830 6351 832
rect 6179 814 6258 830
rect 6265 828 6295 830
rect 6154 812 6258 814
rect 5843 792 5872 802
rect 5886 792 5915 802
rect 5930 792 5960 806
rect 6004 792 6046 806
rect 6068 802 6258 812
rect 6323 810 6329 830
rect 6053 792 6083 802
rect 6084 792 6242 802
rect 6246 792 6276 802
rect 6280 792 6310 806
rect 6338 792 6351 830
rect 6423 844 6452 860
rect 6423 836 6458 844
rect 6423 810 6424 836
rect 6431 810 6458 836
rect 6366 792 6396 806
rect 6423 802 6458 810
rect 6423 792 6452 802
rect -541 778 6452 792
rect -478 748 -465 778
rect -450 764 -420 778
rect -376 764 -334 778
rect -327 764 -107 778
rect -100 764 -70 778
rect -410 750 -395 762
rect -376 750 -363 764
rect -295 760 -142 764
rect -413 748 -391 750
rect -313 748 -121 760
rect -42 748 -29 778
rect -14 764 16 778
rect 53 748 72 778
rect 87 748 93 778
rect 102 748 115 778
rect 130 764 160 778
rect 204 764 246 778
rect 253 764 473 778
rect 480 764 510 778
rect 170 750 185 762
rect 204 750 217 764
rect 285 760 438 764
rect 167 748 189 750
rect 267 748 459 760
rect 538 748 551 778
rect 566 764 596 778
rect 633 748 652 778
rect 667 748 673 778
rect 682 748 695 778
rect 710 764 740 778
rect 784 764 826 778
rect 833 764 1053 778
rect 1060 764 1090 778
rect 750 750 765 762
rect 784 750 797 764
rect 865 760 1018 764
rect 747 748 769 750
rect 847 748 1039 760
rect 1118 748 1131 778
rect 1146 764 1176 778
rect 1213 748 1232 778
rect 1247 748 1253 778
rect 1262 748 1275 778
rect 1290 764 1320 778
rect 1364 764 1406 778
rect 1413 764 1633 778
rect 1640 764 1670 778
rect 1330 750 1345 762
rect 1364 750 1377 764
rect 1445 760 1598 764
rect 1327 748 1349 750
rect 1427 748 1619 760
rect 1698 748 1711 778
rect 1726 764 1756 778
rect 1793 748 1812 778
rect 1827 748 1833 778
rect 1842 748 1855 778
rect 1870 764 1900 778
rect 1944 764 1986 778
rect 1993 764 2213 778
rect 2220 764 2250 778
rect 1910 750 1925 762
rect 1944 750 1957 764
rect 2025 760 2178 764
rect 1907 748 1929 750
rect 2007 748 2199 760
rect 2278 748 2291 778
rect 2306 764 2336 778
rect 2373 748 2392 778
rect 2407 748 2413 778
rect 2422 748 2435 778
rect 2450 764 2480 778
rect 2524 764 2566 778
rect 2573 764 2793 778
rect 2800 764 2830 778
rect 2490 750 2505 762
rect 2524 750 2537 764
rect 2605 760 2758 764
rect 2487 748 2509 750
rect 2587 748 2779 760
rect 2858 748 2871 778
rect 2886 764 2916 778
rect 2953 748 2972 778
rect 2987 748 2993 778
rect 3002 748 3015 778
rect 3030 764 3060 778
rect 3104 764 3146 778
rect 3153 764 3373 778
rect 3380 764 3410 778
rect 3070 750 3085 762
rect 3104 750 3117 764
rect 3185 760 3338 764
rect 3067 748 3089 750
rect 3167 748 3359 760
rect 3438 748 3451 778
rect 3466 764 3496 778
rect 3533 748 3552 778
rect 3567 748 3573 778
rect 3582 748 3595 778
rect 3610 764 3640 778
rect 3684 764 3726 778
rect 3733 764 3953 778
rect 3960 764 3990 778
rect 3650 750 3665 762
rect 3684 750 3697 764
rect 3765 760 3918 764
rect 3647 748 3669 750
rect 3747 748 3939 760
rect 4018 748 4031 778
rect 4046 764 4076 778
rect 4113 748 4132 778
rect 4147 748 4153 778
rect 4162 748 4175 778
rect 4190 764 4220 778
rect 4264 764 4306 778
rect 4313 764 4533 778
rect 4540 764 4570 778
rect 4230 750 4245 762
rect 4264 750 4277 764
rect 4345 760 4498 764
rect 4227 748 4249 750
rect 4327 748 4519 760
rect 4598 748 4611 778
rect 4626 764 4656 778
rect 4693 748 4712 778
rect 4727 748 4733 778
rect 4742 748 4755 778
rect 4770 764 4800 778
rect 4844 764 4886 778
rect 4893 764 5113 778
rect 5120 764 5150 778
rect 4810 750 4825 762
rect 4844 750 4857 764
rect 4925 760 5078 764
rect 4807 748 4829 750
rect 4907 748 5099 760
rect 5178 748 5191 778
rect 5206 764 5236 778
rect 5273 748 5292 778
rect 5307 748 5313 778
rect 5322 748 5335 778
rect 5350 764 5380 778
rect 5424 764 5466 778
rect 5473 764 5693 778
rect 5700 764 5730 778
rect 5390 750 5405 762
rect 5424 750 5437 764
rect 5505 760 5658 764
rect 5387 748 5409 750
rect 5487 748 5679 760
rect 5758 748 5771 778
rect 5786 764 5816 778
rect 5853 748 5872 778
rect 5887 748 5893 778
rect 5902 748 5915 778
rect 5930 764 5960 778
rect 6004 764 6046 778
rect 6053 764 6273 778
rect 6280 764 6310 778
rect 5970 750 5985 762
rect 6004 750 6017 764
rect 6085 760 6238 764
rect 5967 748 5989 750
rect 6067 748 6259 760
rect 6338 748 6351 778
rect 6366 764 6396 778
rect 6439 748 6452 778
rect -541 734 6452 748
rect -478 664 -465 734
rect -413 730 -391 734
rect -420 718 -403 722
rect -399 720 -391 722
rect -401 718 -391 720
rect -420 708 -391 718
rect -338 708 -322 722
rect -284 718 -278 720
rect -271 718 -163 734
rect -156 718 -150 720
rect -142 718 -127 734
rect -61 728 -42 731
rect -420 706 -322 708
rect -295 706 -127 718
rect -112 708 -96 722
rect -61 709 -39 728
rect -29 722 -13 723
rect -30 720 -13 722
rect -29 715 -13 720
rect -39 708 -33 709
rect -30 708 -1 715
rect -112 707 -1 708
rect -112 706 5 707
rect -436 698 -385 706
rect -338 698 -304 706
rect -436 686 -411 698
rect -404 686 -385 698
rect -331 696 -304 698
rect -295 696 -74 706
rect -39 703 -33 706
rect -331 692 -74 696
rect -436 678 -385 686
rect -338 678 -74 692
rect -30 698 5 706
rect -484 630 -465 664
rect -420 670 -391 678
rect -420 664 -403 670
rect -420 662 -386 664
rect -338 662 -322 678
rect -321 668 -113 678
rect -112 668 -96 678
rect -48 674 -33 689
rect -30 686 -29 698
rect -22 686 5 698
rect -30 678 5 686
rect -30 677 -1 678
rect -310 664 -96 668
rect -295 662 -96 664
rect -61 664 -48 674
rect -30 664 -13 677
rect -61 662 -13 664
rect -419 658 -386 662
rect -423 656 -386 658
rect -423 655 -356 656
rect -423 650 -392 655
rect -386 650 -356 655
rect -423 646 -356 650
rect -450 643 -356 646
rect -450 636 -401 643
rect -450 630 -420 636
rect -401 631 -396 636
rect -484 614 -404 630
rect -392 622 -356 643
rect -295 638 -106 662
rect -61 661 -14 662
rect -48 656 -14 661
rect -280 635 -106 638
rect -287 632 -106 635
rect -78 655 -14 656
rect -484 612 -465 614
rect -450 612 -416 614
rect -484 596 -404 612
rect -484 590 -465 596
rect -494 574 -465 590
rect -450 580 -420 596
rect -392 574 -386 622
rect -383 616 -364 622
rect -349 616 -319 624
rect -383 608 -319 616
rect -383 592 -303 608
rect -287 601 -225 632
rect -209 601 -147 632
rect -78 630 -29 655
rect -14 630 16 648
rect -115 616 -85 624
rect -78 622 32 630
rect -115 608 -70 616
rect -383 590 -364 592
rect -349 590 -303 592
rect -383 574 -303 590
rect -276 588 -241 601
rect -200 598 -163 601
rect -200 596 -158 598
rect -271 585 -241 588
rect -262 581 -255 585
rect -255 580 -254 581
rect -296 574 -286 580
rect -500 566 -459 574
rect -500 540 -485 566
rect -478 540 -459 566
rect -395 562 -364 574
rect -349 562 -246 574
rect -234 564 -208 590
rect -193 585 -163 596
rect -131 592 -69 608
rect -131 590 -85 592
rect -131 574 -69 590
rect -57 574 -51 622
rect -48 614 32 622
rect -48 612 -29 614
rect -14 612 20 614
rect -48 597 32 612
rect -48 596 38 597
rect -48 574 -29 596
rect -14 580 16 596
rect 44 590 50 664
rect 53 590 72 734
rect 87 590 93 734
rect 102 664 115 734
rect 167 730 189 734
rect 160 718 177 722
rect 181 720 189 722
rect 179 718 189 720
rect 160 708 189 718
rect 242 708 258 722
rect 296 718 302 720
rect 309 718 417 734
rect 424 718 430 720
rect 438 718 453 734
rect 519 728 538 731
rect 160 706 258 708
rect 285 706 453 718
rect 468 708 484 722
rect 519 709 541 728
rect 551 722 567 723
rect 550 720 567 722
rect 551 715 567 720
rect 541 708 547 709
rect 550 708 579 715
rect 468 707 579 708
rect 468 706 585 707
rect 144 698 195 706
rect 242 698 276 706
rect 144 686 169 698
rect 176 686 195 698
rect 249 696 276 698
rect 285 696 506 706
rect 541 703 547 706
rect 249 692 506 696
rect 144 678 195 686
rect 242 678 506 692
rect 550 698 585 706
rect 96 630 115 664
rect 160 670 189 678
rect 160 664 177 670
rect 160 662 194 664
rect 242 662 258 678
rect 259 668 467 678
rect 468 668 484 678
rect 532 674 547 689
rect 550 686 551 698
rect 558 686 585 698
rect 550 678 585 686
rect 550 677 579 678
rect 270 664 484 668
rect 285 662 484 664
rect 519 664 532 674
rect 550 664 567 677
rect 519 662 567 664
rect 161 658 194 662
rect 157 656 194 658
rect 157 655 224 656
rect 157 650 188 655
rect 194 650 224 655
rect 157 646 224 650
rect 130 643 224 646
rect 130 636 179 643
rect 130 630 160 636
rect 179 631 184 636
rect 96 614 176 630
rect 188 622 224 643
rect 285 638 474 662
rect 519 661 566 662
rect 532 656 566 661
rect 606 656 622 658
rect 300 635 474 638
rect 293 632 474 635
rect 502 655 566 656
rect 96 612 115 614
rect 130 612 164 614
rect 96 596 176 612
rect 96 590 115 596
rect -188 564 -85 574
rect -234 562 -85 564
rect -64 562 -29 574
rect -395 560 -233 562
rect -383 540 -364 560
rect -349 558 -319 560
rect -500 532 -459 540
rect -377 536 -364 540
rect -312 544 -233 560
rect -201 560 -29 562
rect -201 544 -122 560
rect -115 558 -85 560
rect -494 522 -465 532
rect -450 522 -420 536
rect -377 522 -334 536
rect -312 532 -122 544
rect -57 540 -51 560
rect -327 522 -297 532
rect -296 522 -138 532
rect -134 522 -104 532
rect -100 522 -70 536
rect -42 522 -29 560
rect 43 574 72 590
rect 86 574 115 590
rect 130 580 160 596
rect 188 574 194 622
rect 197 616 216 622
rect 231 616 261 624
rect 197 608 261 616
rect 197 592 277 608
rect 293 601 355 632
rect 371 601 433 632
rect 502 630 551 655
rect 596 646 622 656
rect 566 630 622 646
rect 465 616 495 624
rect 502 622 612 630
rect 465 608 510 616
rect 197 590 216 592
rect 231 590 277 592
rect 197 574 277 590
rect 304 588 339 601
rect 380 598 417 601
rect 380 596 422 598
rect 309 585 339 588
rect 318 581 325 585
rect 325 580 326 581
rect 284 574 294 580
rect 43 566 78 574
rect 43 540 44 566
rect 51 540 78 566
rect -14 522 16 536
rect 43 532 78 540
rect 80 566 121 574
rect 80 540 95 566
rect 102 540 121 566
rect 185 562 216 574
rect 231 562 334 574
rect 346 564 372 590
rect 387 585 417 596
rect 449 592 511 608
rect 449 590 495 592
rect 449 574 511 590
rect 523 574 529 622
rect 532 614 612 622
rect 532 612 551 614
rect 566 612 600 614
rect 532 596 612 612
rect 532 574 551 596
rect 566 580 596 596
rect 624 590 630 664
rect 633 590 652 734
rect 667 590 673 734
rect 682 664 695 734
rect 747 730 769 734
rect 740 718 757 722
rect 761 720 769 722
rect 759 718 769 720
rect 740 708 769 718
rect 822 708 838 722
rect 876 718 882 720
rect 889 718 997 734
rect 1004 718 1010 720
rect 1018 718 1033 734
rect 1099 728 1118 731
rect 740 706 838 708
rect 865 706 1033 718
rect 1048 708 1064 722
rect 1099 709 1121 728
rect 1131 722 1147 723
rect 1130 720 1147 722
rect 1131 715 1147 720
rect 1121 708 1127 709
rect 1130 708 1159 715
rect 1048 707 1159 708
rect 1048 706 1165 707
rect 724 698 775 706
rect 822 698 856 706
rect 724 686 749 698
rect 756 686 775 698
rect 829 696 856 698
rect 865 696 1086 706
rect 1121 703 1127 706
rect 829 692 1086 696
rect 724 678 775 686
rect 822 678 1086 692
rect 1130 698 1165 706
rect 676 630 695 664
rect 740 670 769 678
rect 740 664 757 670
rect 740 662 774 664
rect 822 662 838 678
rect 839 668 1047 678
rect 1048 668 1064 678
rect 1112 674 1127 689
rect 1130 686 1131 698
rect 1138 686 1165 698
rect 1130 678 1165 686
rect 1130 677 1159 678
rect 850 664 1064 668
rect 865 662 1064 664
rect 1099 664 1112 674
rect 1130 664 1147 677
rect 1099 662 1147 664
rect 741 658 774 662
rect 737 656 774 658
rect 737 655 804 656
rect 737 650 768 655
rect 774 650 804 655
rect 737 646 804 650
rect 710 643 804 646
rect 710 636 759 643
rect 710 630 740 636
rect 759 631 764 636
rect 676 614 756 630
rect 768 622 804 643
rect 865 638 1054 662
rect 1099 661 1146 662
rect 1112 656 1146 661
rect 880 635 1054 638
rect 873 632 1054 635
rect 1082 655 1146 656
rect 676 612 695 614
rect 710 612 744 614
rect 676 596 756 612
rect 676 590 695 596
rect 392 564 495 574
rect 346 562 495 564
rect 516 562 551 574
rect 185 560 347 562
rect 197 540 216 560
rect 231 558 261 560
rect 80 532 121 540
rect 203 536 216 540
rect 268 544 347 560
rect 379 560 551 562
rect 379 544 458 560
rect 465 558 495 560
rect 43 522 72 532
rect 86 522 115 532
rect 130 522 160 536
rect 203 522 246 536
rect 268 532 458 544
rect 523 540 529 560
rect 253 522 283 532
rect 284 522 442 532
rect 446 522 476 532
rect 480 522 510 536
rect 538 522 551 560
rect 623 574 652 590
rect 666 574 695 590
rect 710 580 740 596
rect 768 574 774 622
rect 777 616 796 622
rect 811 616 841 624
rect 777 608 841 616
rect 777 592 857 608
rect 873 601 935 632
rect 951 601 1013 632
rect 1082 630 1131 655
rect 1146 630 1176 648
rect 1045 616 1075 624
rect 1082 622 1192 630
rect 1045 608 1090 616
rect 777 590 796 592
rect 811 590 857 592
rect 777 574 857 590
rect 884 588 919 601
rect 960 598 997 601
rect 960 596 1002 598
rect 889 585 919 588
rect 898 581 905 585
rect 905 580 906 581
rect 864 574 874 580
rect 623 566 658 574
rect 623 540 624 566
rect 631 540 658 566
rect 566 522 596 536
rect 623 532 658 540
rect 660 566 701 574
rect 660 540 675 566
rect 682 540 701 566
rect 765 562 796 574
rect 811 562 914 574
rect 926 564 952 590
rect 967 585 997 596
rect 1029 592 1091 608
rect 1029 590 1075 592
rect 1029 574 1091 590
rect 1103 574 1109 622
rect 1112 614 1192 622
rect 1112 612 1131 614
rect 1146 612 1180 614
rect 1112 597 1192 612
rect 1112 596 1198 597
rect 1112 574 1131 596
rect 1146 580 1176 596
rect 1204 590 1210 664
rect 1213 590 1232 734
rect 1247 590 1253 734
rect 1262 664 1275 734
rect 1327 730 1349 734
rect 1320 718 1337 722
rect 1341 720 1349 722
rect 1339 718 1349 720
rect 1320 708 1349 718
rect 1402 708 1418 722
rect 1456 718 1462 720
rect 1469 718 1577 734
rect 1584 718 1590 720
rect 1598 718 1613 734
rect 1679 728 1698 731
rect 1320 706 1418 708
rect 1445 706 1613 718
rect 1628 708 1644 722
rect 1679 709 1701 728
rect 1711 722 1727 723
rect 1710 720 1727 722
rect 1711 715 1727 720
rect 1701 708 1707 709
rect 1710 708 1739 715
rect 1628 707 1739 708
rect 1628 706 1745 707
rect 1304 698 1355 706
rect 1402 698 1436 706
rect 1304 686 1329 698
rect 1336 686 1355 698
rect 1409 696 1436 698
rect 1445 696 1666 706
rect 1701 703 1707 706
rect 1409 692 1666 696
rect 1304 678 1355 686
rect 1402 678 1666 692
rect 1710 698 1745 706
rect 1256 630 1275 664
rect 1320 670 1349 678
rect 1320 664 1337 670
rect 1320 662 1354 664
rect 1402 662 1418 678
rect 1419 668 1627 678
rect 1628 668 1644 678
rect 1692 674 1707 689
rect 1710 686 1711 698
rect 1718 686 1745 698
rect 1710 678 1745 686
rect 1710 677 1739 678
rect 1430 664 1644 668
rect 1445 662 1644 664
rect 1679 664 1692 674
rect 1710 664 1727 677
rect 1679 662 1727 664
rect 1321 658 1354 662
rect 1317 656 1354 658
rect 1317 655 1384 656
rect 1317 650 1348 655
rect 1354 650 1384 655
rect 1317 646 1384 650
rect 1290 643 1384 646
rect 1290 636 1339 643
rect 1290 630 1320 636
rect 1339 631 1344 636
rect 1256 614 1336 630
rect 1348 622 1384 643
rect 1445 638 1634 662
rect 1679 661 1726 662
rect 1692 656 1726 661
rect 1766 656 1782 658
rect 1460 635 1634 638
rect 1453 632 1634 635
rect 1662 655 1726 656
rect 1256 612 1275 614
rect 1290 612 1324 614
rect 1256 596 1336 612
rect 1256 590 1275 596
rect 972 564 1075 574
rect 926 562 1075 564
rect 1096 562 1131 574
rect 765 560 927 562
rect 777 540 796 560
rect 811 558 841 560
rect 660 532 701 540
rect 783 536 796 540
rect 848 544 927 560
rect 959 560 1131 562
rect 959 544 1038 560
rect 1045 558 1075 560
rect 623 522 652 532
rect 666 522 695 532
rect 710 522 740 536
rect 783 522 826 536
rect 848 532 1038 544
rect 1103 540 1109 560
rect 833 522 863 532
rect 864 522 1022 532
rect 1026 522 1056 532
rect 1060 522 1090 536
rect 1118 522 1131 560
rect 1203 574 1232 590
rect 1246 574 1275 590
rect 1290 580 1320 596
rect 1348 574 1354 622
rect 1357 616 1376 622
rect 1391 616 1421 624
rect 1357 608 1421 616
rect 1357 592 1437 608
rect 1453 601 1515 632
rect 1531 601 1593 632
rect 1662 630 1711 655
rect 1756 646 1782 656
rect 1726 630 1782 646
rect 1625 616 1655 624
rect 1662 622 1772 630
rect 1625 608 1670 616
rect 1357 590 1376 592
rect 1391 590 1437 592
rect 1357 574 1437 590
rect 1464 588 1499 601
rect 1540 598 1577 601
rect 1540 596 1582 598
rect 1469 585 1499 588
rect 1478 581 1485 585
rect 1485 580 1486 581
rect 1444 574 1454 580
rect 1203 566 1238 574
rect 1203 540 1204 566
rect 1211 540 1238 566
rect 1146 522 1176 536
rect 1203 532 1238 540
rect 1240 566 1281 574
rect 1240 540 1255 566
rect 1262 540 1281 566
rect 1345 562 1376 574
rect 1391 562 1494 574
rect 1506 564 1532 590
rect 1547 585 1577 596
rect 1609 592 1671 608
rect 1609 590 1655 592
rect 1609 574 1671 590
rect 1683 574 1689 622
rect 1692 614 1772 622
rect 1692 612 1711 614
rect 1726 612 1760 614
rect 1692 596 1772 612
rect 1692 574 1711 596
rect 1726 580 1756 596
rect 1784 590 1790 664
rect 1793 590 1812 734
rect 1827 590 1833 734
rect 1842 664 1855 734
rect 1907 730 1929 734
rect 1900 718 1917 722
rect 1921 720 1929 722
rect 1919 718 1929 720
rect 1900 708 1929 718
rect 1982 708 1998 722
rect 2036 718 2042 720
rect 2049 718 2157 734
rect 2164 718 2170 720
rect 2178 718 2193 734
rect 2259 728 2278 731
rect 1900 706 1998 708
rect 2025 706 2193 718
rect 2208 708 2224 722
rect 2259 709 2281 728
rect 2291 722 2307 723
rect 2290 720 2307 722
rect 2291 715 2307 720
rect 2281 708 2287 709
rect 2290 708 2319 715
rect 2208 707 2319 708
rect 2208 706 2325 707
rect 1884 698 1935 706
rect 1982 698 2016 706
rect 1884 686 1909 698
rect 1916 686 1935 698
rect 1989 696 2016 698
rect 2025 696 2246 706
rect 2281 703 2287 706
rect 1989 692 2246 696
rect 1884 678 1935 686
rect 1982 678 2246 692
rect 2290 698 2325 706
rect 1836 630 1855 664
rect 1900 670 1929 678
rect 1900 664 1917 670
rect 1900 662 1934 664
rect 1982 662 1998 678
rect 1999 668 2207 678
rect 2208 668 2224 678
rect 2272 674 2287 689
rect 2290 686 2291 698
rect 2298 686 2325 698
rect 2290 678 2325 686
rect 2290 677 2319 678
rect 2010 664 2224 668
rect 2025 662 2224 664
rect 2259 664 2272 674
rect 2290 664 2307 677
rect 2259 662 2307 664
rect 1901 658 1934 662
rect 1897 656 1934 658
rect 1897 655 1964 656
rect 1897 650 1928 655
rect 1934 650 1964 655
rect 1897 646 1964 650
rect 1870 643 1964 646
rect 1870 636 1919 643
rect 1870 630 1900 636
rect 1919 631 1924 636
rect 1836 614 1916 630
rect 1928 622 1964 643
rect 2025 638 2214 662
rect 2259 661 2306 662
rect 2272 656 2306 661
rect 2040 635 2214 638
rect 2033 632 2214 635
rect 2242 655 2306 656
rect 1836 612 1855 614
rect 1870 612 1904 614
rect 1836 596 1916 612
rect 1836 590 1855 596
rect 1552 564 1655 574
rect 1506 562 1655 564
rect 1676 562 1711 574
rect 1345 560 1507 562
rect 1357 540 1376 560
rect 1391 558 1421 560
rect 1240 532 1281 540
rect 1363 536 1376 540
rect 1428 544 1507 560
rect 1539 560 1711 562
rect 1539 544 1618 560
rect 1625 558 1655 560
rect 1203 522 1232 532
rect 1246 522 1275 532
rect 1290 522 1320 536
rect 1363 522 1406 536
rect 1428 532 1618 544
rect 1683 540 1689 560
rect 1413 522 1443 532
rect 1444 522 1602 532
rect 1606 522 1636 532
rect 1640 522 1670 536
rect 1698 522 1711 560
rect 1783 574 1812 590
rect 1826 574 1855 590
rect 1870 580 1900 596
rect 1928 574 1934 622
rect 1937 616 1956 622
rect 1971 616 2001 624
rect 1937 608 2001 616
rect 1937 592 2017 608
rect 2033 601 2095 632
rect 2111 601 2173 632
rect 2242 630 2291 655
rect 2306 630 2336 648
rect 2205 616 2235 624
rect 2242 622 2352 630
rect 2205 608 2250 616
rect 1937 590 1956 592
rect 1971 590 2017 592
rect 1937 574 2017 590
rect 2044 588 2079 601
rect 2120 598 2157 601
rect 2120 596 2162 598
rect 2049 585 2079 588
rect 2058 581 2065 585
rect 2065 580 2066 581
rect 2024 574 2034 580
rect 1783 566 1818 574
rect 1783 540 1784 566
rect 1791 540 1818 566
rect 1726 522 1756 536
rect 1783 532 1818 540
rect 1820 566 1861 574
rect 1820 540 1835 566
rect 1842 540 1861 566
rect 1925 562 1956 574
rect 1971 562 2074 574
rect 2086 564 2112 590
rect 2127 585 2157 596
rect 2189 592 2251 608
rect 2189 590 2235 592
rect 2189 574 2251 590
rect 2263 574 2269 622
rect 2272 614 2352 622
rect 2272 612 2291 614
rect 2306 612 2340 614
rect 2272 597 2352 612
rect 2272 596 2358 597
rect 2272 574 2291 596
rect 2306 580 2336 596
rect 2364 590 2370 664
rect 2373 590 2392 734
rect 2407 590 2413 734
rect 2422 664 2435 734
rect 2487 730 2509 734
rect 2480 718 2497 722
rect 2501 720 2509 722
rect 2499 718 2509 720
rect 2480 708 2509 718
rect 2562 708 2578 722
rect 2616 718 2622 720
rect 2629 718 2737 734
rect 2744 718 2750 720
rect 2758 718 2773 734
rect 2839 728 2858 731
rect 2480 706 2578 708
rect 2605 706 2773 718
rect 2788 708 2804 722
rect 2839 709 2861 728
rect 2871 722 2887 723
rect 2870 720 2887 722
rect 2871 715 2887 720
rect 2861 708 2867 709
rect 2870 708 2899 715
rect 2788 707 2899 708
rect 2788 706 2905 707
rect 2464 698 2515 706
rect 2562 698 2596 706
rect 2464 686 2489 698
rect 2496 686 2515 698
rect 2569 696 2596 698
rect 2605 696 2826 706
rect 2861 703 2867 706
rect 2569 692 2826 696
rect 2464 678 2515 686
rect 2562 678 2826 692
rect 2870 698 2905 706
rect 2416 630 2435 664
rect 2480 670 2509 678
rect 2480 664 2497 670
rect 2480 662 2514 664
rect 2562 662 2578 678
rect 2579 668 2787 678
rect 2788 668 2804 678
rect 2852 674 2867 689
rect 2870 686 2871 698
rect 2878 686 2905 698
rect 2870 678 2905 686
rect 2870 677 2899 678
rect 2590 664 2804 668
rect 2605 662 2804 664
rect 2839 664 2852 674
rect 2870 664 2887 677
rect 2839 662 2887 664
rect 2481 658 2514 662
rect 2477 656 2514 658
rect 2477 655 2544 656
rect 2477 650 2508 655
rect 2514 650 2544 655
rect 2477 646 2544 650
rect 2450 643 2544 646
rect 2450 636 2499 643
rect 2450 630 2480 636
rect 2499 631 2504 636
rect 2416 614 2496 630
rect 2508 622 2544 643
rect 2605 638 2794 662
rect 2839 661 2886 662
rect 2852 656 2886 661
rect 2926 656 2942 658
rect 2620 635 2794 638
rect 2613 632 2794 635
rect 2822 655 2886 656
rect 2416 612 2435 614
rect 2450 612 2484 614
rect 2416 596 2496 612
rect 2416 590 2435 596
rect 2132 564 2235 574
rect 2086 562 2235 564
rect 2256 562 2291 574
rect 1925 560 2087 562
rect 1937 540 1956 560
rect 1971 558 2001 560
rect 1820 532 1861 540
rect 1943 536 1956 540
rect 2008 544 2087 560
rect 2119 560 2291 562
rect 2119 544 2198 560
rect 2205 558 2235 560
rect 1783 522 1812 532
rect 1826 522 1855 532
rect 1870 522 1900 536
rect 1943 522 1986 536
rect 2008 532 2198 544
rect 2263 540 2269 560
rect 1993 522 2023 532
rect 2024 522 2182 532
rect 2186 522 2216 532
rect 2220 522 2250 536
rect 2278 522 2291 560
rect 2363 574 2392 590
rect 2406 574 2435 590
rect 2450 580 2480 596
rect 2508 574 2514 622
rect 2517 616 2536 622
rect 2551 616 2581 624
rect 2517 608 2581 616
rect 2517 592 2597 608
rect 2613 601 2675 632
rect 2691 601 2753 632
rect 2822 630 2871 655
rect 2916 646 2942 656
rect 2886 630 2942 646
rect 2785 616 2815 624
rect 2822 622 2932 630
rect 2785 608 2830 616
rect 2517 590 2536 592
rect 2551 590 2597 592
rect 2517 574 2597 590
rect 2624 588 2659 601
rect 2700 598 2737 601
rect 2700 596 2742 598
rect 2629 585 2659 588
rect 2638 581 2645 585
rect 2645 580 2646 581
rect 2604 574 2614 580
rect 2363 566 2398 574
rect 2363 540 2364 566
rect 2371 540 2398 566
rect 2306 522 2336 536
rect 2363 532 2398 540
rect 2400 566 2441 574
rect 2400 540 2415 566
rect 2422 540 2441 566
rect 2505 562 2536 574
rect 2551 562 2654 574
rect 2666 564 2692 590
rect 2707 585 2737 596
rect 2769 592 2831 608
rect 2769 590 2815 592
rect 2769 574 2831 590
rect 2843 574 2849 622
rect 2852 614 2932 622
rect 2852 612 2871 614
rect 2886 612 2920 614
rect 2852 596 2932 612
rect 2852 574 2871 596
rect 2886 580 2916 596
rect 2944 590 2950 664
rect 2953 590 2972 734
rect 2987 590 2993 734
rect 3002 664 3015 734
rect 3067 730 3089 734
rect 3060 718 3077 722
rect 3081 720 3089 722
rect 3079 718 3089 720
rect 3060 708 3089 718
rect 3142 708 3158 722
rect 3196 718 3202 720
rect 3209 718 3317 734
rect 3324 718 3330 720
rect 3338 718 3353 734
rect 3419 728 3438 731
rect 3060 706 3158 708
rect 3185 706 3353 718
rect 3368 708 3384 722
rect 3419 709 3441 728
rect 3451 722 3467 723
rect 3450 720 3467 722
rect 3451 715 3467 720
rect 3441 708 3447 709
rect 3450 708 3479 715
rect 3368 707 3479 708
rect 3368 706 3485 707
rect 3044 698 3095 706
rect 3142 698 3176 706
rect 3044 686 3069 698
rect 3076 686 3095 698
rect 3149 696 3176 698
rect 3185 696 3406 706
rect 3441 703 3447 706
rect 3149 692 3406 696
rect 3044 678 3095 686
rect 3142 678 3406 692
rect 3450 698 3485 706
rect 2996 630 3015 664
rect 3060 670 3089 678
rect 3060 664 3077 670
rect 3060 662 3094 664
rect 3142 662 3158 678
rect 3159 668 3367 678
rect 3368 668 3384 678
rect 3432 674 3447 689
rect 3450 686 3451 698
rect 3458 686 3485 698
rect 3450 678 3485 686
rect 3450 677 3479 678
rect 3170 664 3384 668
rect 3185 662 3384 664
rect 3419 664 3432 674
rect 3450 664 3467 677
rect 3419 662 3467 664
rect 3061 658 3094 662
rect 3057 656 3094 658
rect 3057 655 3124 656
rect 3057 650 3088 655
rect 3094 650 3124 655
rect 3057 646 3124 650
rect 3030 643 3124 646
rect 3030 636 3079 643
rect 3030 630 3060 636
rect 3079 631 3084 636
rect 2996 614 3076 630
rect 3088 622 3124 643
rect 3185 638 3374 662
rect 3419 661 3466 662
rect 3432 656 3466 661
rect 3200 635 3374 638
rect 3193 632 3374 635
rect 3402 655 3466 656
rect 2996 612 3015 614
rect 3030 612 3064 614
rect 2996 596 3076 612
rect 2996 590 3015 596
rect 2712 564 2815 574
rect 2666 562 2815 564
rect 2836 562 2871 574
rect 2505 560 2667 562
rect 2517 540 2536 560
rect 2551 558 2581 560
rect 2400 532 2441 540
rect 2523 536 2536 540
rect 2588 544 2667 560
rect 2699 560 2871 562
rect 2699 544 2778 560
rect 2785 558 2815 560
rect 2363 522 2392 532
rect 2406 522 2435 532
rect 2450 522 2480 536
rect 2523 522 2566 536
rect 2588 532 2778 544
rect 2843 540 2849 560
rect 2573 522 2603 532
rect 2604 522 2762 532
rect 2766 522 2796 532
rect 2800 522 2830 536
rect 2858 522 2871 560
rect 2943 574 2972 590
rect 2986 574 3015 590
rect 3030 580 3060 596
rect 3088 574 3094 622
rect 3097 616 3116 622
rect 3131 616 3161 624
rect 3097 608 3161 616
rect 3097 592 3177 608
rect 3193 601 3255 632
rect 3271 601 3333 632
rect 3402 630 3451 655
rect 3466 630 3496 648
rect 3365 616 3395 624
rect 3402 622 3512 630
rect 3365 608 3410 616
rect 3097 590 3116 592
rect 3131 590 3177 592
rect 3097 574 3177 590
rect 3204 588 3239 601
rect 3280 598 3317 601
rect 3280 596 3322 598
rect 3209 585 3239 588
rect 3218 581 3225 585
rect 3225 580 3226 581
rect 3184 574 3194 580
rect 2943 566 2978 574
rect 2943 540 2944 566
rect 2951 540 2978 566
rect 2886 522 2916 536
rect 2943 532 2978 540
rect 2980 566 3021 574
rect 2980 540 2995 566
rect 3002 540 3021 566
rect 3085 562 3116 574
rect 3131 562 3234 574
rect 3246 564 3272 590
rect 3287 585 3317 596
rect 3349 592 3411 608
rect 3349 590 3395 592
rect 3349 574 3411 590
rect 3423 574 3429 622
rect 3432 614 3512 622
rect 3432 612 3451 614
rect 3466 612 3500 614
rect 3432 597 3512 612
rect 3432 596 3518 597
rect 3432 574 3451 596
rect 3466 580 3496 596
rect 3524 590 3530 664
rect 3533 590 3552 734
rect 3567 590 3573 734
rect 3582 664 3595 734
rect 3647 730 3669 734
rect 3640 718 3657 722
rect 3661 720 3669 722
rect 3659 718 3669 720
rect 3640 708 3669 718
rect 3722 708 3738 722
rect 3776 718 3782 720
rect 3789 718 3897 734
rect 3904 718 3910 720
rect 3918 718 3933 734
rect 3999 728 4018 731
rect 3640 706 3738 708
rect 3765 706 3933 718
rect 3948 708 3964 722
rect 3999 709 4021 728
rect 4031 722 4047 723
rect 4030 720 4047 722
rect 4031 715 4047 720
rect 4021 708 4027 709
rect 4030 708 4059 715
rect 3948 707 4059 708
rect 3948 706 4065 707
rect 3624 698 3675 706
rect 3722 698 3756 706
rect 3624 686 3649 698
rect 3656 686 3675 698
rect 3729 696 3756 698
rect 3765 696 3986 706
rect 4021 703 4027 706
rect 3729 692 3986 696
rect 3624 678 3675 686
rect 3722 678 3986 692
rect 4030 698 4065 706
rect 3576 630 3595 664
rect 3640 670 3669 678
rect 3640 664 3657 670
rect 3640 662 3674 664
rect 3722 662 3738 678
rect 3739 668 3947 678
rect 3948 668 3964 678
rect 4012 674 4027 689
rect 4030 686 4031 698
rect 4038 686 4065 698
rect 4030 678 4065 686
rect 4030 677 4059 678
rect 3750 664 3964 668
rect 3765 662 3964 664
rect 3999 664 4012 674
rect 4030 664 4047 677
rect 3999 662 4047 664
rect 3641 658 3674 662
rect 3637 656 3674 658
rect 3637 655 3704 656
rect 3637 650 3668 655
rect 3674 650 3704 655
rect 3637 646 3704 650
rect 3610 643 3704 646
rect 3610 636 3659 643
rect 3610 630 3640 636
rect 3659 631 3664 636
rect 3576 614 3656 630
rect 3668 622 3704 643
rect 3765 638 3954 662
rect 3999 661 4046 662
rect 4012 656 4046 661
rect 4086 656 4102 658
rect 3780 635 3954 638
rect 3773 632 3954 635
rect 3982 655 4046 656
rect 3576 612 3595 614
rect 3610 612 3644 614
rect 3576 596 3656 612
rect 3576 590 3595 596
rect 3292 564 3395 574
rect 3246 562 3395 564
rect 3416 562 3451 574
rect 3085 560 3247 562
rect 3097 540 3116 560
rect 3131 558 3161 560
rect 2980 532 3021 540
rect 3103 536 3116 540
rect 3168 544 3247 560
rect 3279 560 3451 562
rect 3279 544 3358 560
rect 3365 558 3395 560
rect 2943 522 2972 532
rect 2986 522 3015 532
rect 3030 522 3060 536
rect 3103 522 3146 536
rect 3168 532 3358 544
rect 3423 540 3429 560
rect 3153 522 3183 532
rect 3184 522 3342 532
rect 3346 522 3376 532
rect 3380 522 3410 536
rect 3438 522 3451 560
rect 3523 574 3552 590
rect 3566 574 3595 590
rect 3610 580 3640 596
rect 3668 574 3674 622
rect 3677 616 3696 622
rect 3711 616 3741 624
rect 3677 608 3741 616
rect 3677 592 3757 608
rect 3773 601 3835 632
rect 3851 601 3913 632
rect 3982 630 4031 655
rect 4076 646 4102 656
rect 4046 630 4102 646
rect 3945 616 3975 624
rect 3982 622 4092 630
rect 3945 608 3990 616
rect 3677 590 3696 592
rect 3711 590 3757 592
rect 3677 574 3757 590
rect 3784 588 3819 601
rect 3860 598 3897 601
rect 3860 596 3902 598
rect 3789 585 3819 588
rect 3798 581 3805 585
rect 3805 580 3806 581
rect 3764 574 3774 580
rect 3523 566 3558 574
rect 3523 540 3524 566
rect 3531 540 3558 566
rect 3466 522 3496 536
rect 3523 532 3558 540
rect 3560 566 3601 574
rect 3560 540 3575 566
rect 3582 540 3601 566
rect 3665 562 3696 574
rect 3711 562 3814 574
rect 3826 564 3852 590
rect 3867 585 3897 596
rect 3929 592 3991 608
rect 3929 590 3975 592
rect 3929 574 3991 590
rect 4003 574 4009 622
rect 4012 614 4092 622
rect 4012 612 4031 614
rect 4046 612 4080 614
rect 4012 596 4092 612
rect 4012 574 4031 596
rect 4046 580 4076 596
rect 4104 590 4110 664
rect 4113 590 4132 734
rect 4147 590 4153 734
rect 4162 664 4175 734
rect 4227 730 4249 734
rect 4220 718 4237 722
rect 4241 720 4249 722
rect 4239 718 4249 720
rect 4220 708 4249 718
rect 4302 708 4318 722
rect 4356 718 4362 720
rect 4369 718 4477 734
rect 4484 718 4490 720
rect 4498 718 4513 734
rect 4579 728 4598 731
rect 4220 706 4318 708
rect 4345 706 4513 718
rect 4528 708 4544 722
rect 4579 709 4601 728
rect 4611 722 4627 723
rect 4610 720 4627 722
rect 4611 715 4627 720
rect 4601 708 4607 709
rect 4610 708 4639 715
rect 4528 707 4639 708
rect 4528 706 4645 707
rect 4204 698 4255 706
rect 4302 698 4336 706
rect 4204 686 4229 698
rect 4236 686 4255 698
rect 4309 696 4336 698
rect 4345 696 4566 706
rect 4601 703 4607 706
rect 4309 692 4566 696
rect 4204 678 4255 686
rect 4302 678 4566 692
rect 4610 698 4645 706
rect 4156 630 4175 664
rect 4220 670 4249 678
rect 4220 664 4237 670
rect 4220 662 4254 664
rect 4302 662 4318 678
rect 4319 668 4527 678
rect 4528 668 4544 678
rect 4592 674 4607 689
rect 4610 686 4611 698
rect 4618 686 4645 698
rect 4610 678 4645 686
rect 4610 677 4639 678
rect 4330 664 4544 668
rect 4345 662 4544 664
rect 4579 664 4592 674
rect 4610 664 4627 677
rect 4579 662 4627 664
rect 4221 658 4254 662
rect 4217 656 4254 658
rect 4217 655 4284 656
rect 4217 650 4248 655
rect 4254 650 4284 655
rect 4217 646 4284 650
rect 4190 643 4284 646
rect 4190 636 4239 643
rect 4190 630 4220 636
rect 4239 631 4244 636
rect 4156 614 4236 630
rect 4248 622 4284 643
rect 4345 638 4534 662
rect 4579 661 4626 662
rect 4592 656 4626 661
rect 4360 635 4534 638
rect 4353 632 4534 635
rect 4562 655 4626 656
rect 4156 612 4175 614
rect 4190 612 4224 614
rect 4156 596 4236 612
rect 4156 590 4175 596
rect 3872 564 3975 574
rect 3826 562 3975 564
rect 3996 562 4031 574
rect 3665 560 3827 562
rect 3677 540 3696 560
rect 3711 558 3741 560
rect 3560 532 3601 540
rect 3683 536 3696 540
rect 3748 544 3827 560
rect 3859 560 4031 562
rect 3859 544 3938 560
rect 3945 558 3975 560
rect 3523 522 3552 532
rect 3566 522 3595 532
rect 3610 522 3640 536
rect 3683 522 3726 536
rect 3748 532 3938 544
rect 4003 540 4009 560
rect 3733 522 3763 532
rect 3764 522 3922 532
rect 3926 522 3956 532
rect 3960 522 3990 536
rect 4018 522 4031 560
rect 4103 574 4132 590
rect 4146 574 4175 590
rect 4190 580 4220 596
rect 4248 574 4254 622
rect 4257 616 4276 622
rect 4291 616 4321 624
rect 4257 608 4321 616
rect 4257 592 4337 608
rect 4353 601 4415 632
rect 4431 601 4493 632
rect 4562 630 4611 655
rect 4626 630 4656 648
rect 4525 616 4555 624
rect 4562 622 4672 630
rect 4525 608 4570 616
rect 4257 590 4276 592
rect 4291 590 4337 592
rect 4257 574 4337 590
rect 4364 588 4399 601
rect 4440 598 4477 601
rect 4440 596 4482 598
rect 4369 585 4399 588
rect 4378 581 4385 585
rect 4385 580 4386 581
rect 4344 574 4354 580
rect 4103 566 4138 574
rect 4103 540 4104 566
rect 4111 540 4138 566
rect 4046 522 4076 536
rect 4103 532 4138 540
rect 4140 566 4181 574
rect 4140 540 4155 566
rect 4162 540 4181 566
rect 4245 562 4276 574
rect 4291 562 4394 574
rect 4406 564 4432 590
rect 4447 585 4477 596
rect 4509 592 4571 608
rect 4509 590 4555 592
rect 4509 574 4571 590
rect 4583 574 4589 622
rect 4592 614 4672 622
rect 4592 612 4611 614
rect 4626 612 4660 614
rect 4592 597 4672 612
rect 4592 596 4678 597
rect 4592 574 4611 596
rect 4626 580 4656 596
rect 4684 590 4690 664
rect 4693 590 4712 734
rect 4727 590 4733 734
rect 4742 664 4755 734
rect 4807 730 4829 734
rect 4800 718 4817 722
rect 4821 720 4829 722
rect 4819 718 4829 720
rect 4800 708 4829 718
rect 4882 708 4898 722
rect 4936 718 4942 720
rect 4949 718 5057 734
rect 5064 718 5070 720
rect 5078 718 5093 734
rect 5159 728 5178 731
rect 4800 706 4898 708
rect 4925 706 5093 718
rect 5108 708 5124 722
rect 5159 709 5181 728
rect 5191 722 5207 723
rect 5190 720 5207 722
rect 5191 715 5207 720
rect 5181 708 5187 709
rect 5190 708 5219 715
rect 5108 707 5219 708
rect 5108 706 5225 707
rect 4784 698 4835 706
rect 4882 698 4916 706
rect 4784 686 4809 698
rect 4816 686 4835 698
rect 4889 696 4916 698
rect 4925 696 5146 706
rect 5181 703 5187 706
rect 4889 692 5146 696
rect 4784 678 4835 686
rect 4882 678 5146 692
rect 5190 698 5225 706
rect 4736 630 4755 664
rect 4800 670 4829 678
rect 4800 664 4817 670
rect 4800 662 4834 664
rect 4882 662 4898 678
rect 4899 668 5107 678
rect 5108 668 5124 678
rect 5172 674 5187 689
rect 5190 686 5191 698
rect 5198 686 5225 698
rect 5190 678 5225 686
rect 5190 677 5219 678
rect 4910 664 5124 668
rect 4925 662 5124 664
rect 5159 664 5172 674
rect 5190 664 5207 677
rect 5159 662 5207 664
rect 4801 658 4834 662
rect 4797 656 4834 658
rect 4797 655 4864 656
rect 4797 650 4828 655
rect 4834 650 4864 655
rect 4797 646 4864 650
rect 4770 643 4864 646
rect 4770 636 4819 643
rect 4770 630 4800 636
rect 4819 631 4824 636
rect 4736 614 4816 630
rect 4828 622 4864 643
rect 4925 638 5114 662
rect 5159 661 5206 662
rect 5172 656 5206 661
rect 5246 656 5262 658
rect 4940 635 5114 638
rect 4933 632 5114 635
rect 5142 655 5206 656
rect 4736 612 4755 614
rect 4770 612 4804 614
rect 4736 596 4816 612
rect 4736 590 4755 596
rect 4452 564 4555 574
rect 4406 562 4555 564
rect 4576 562 4611 574
rect 4245 560 4407 562
rect 4257 540 4276 560
rect 4291 558 4321 560
rect 4140 532 4181 540
rect 4263 536 4276 540
rect 4328 544 4407 560
rect 4439 560 4611 562
rect 4439 544 4518 560
rect 4525 558 4555 560
rect 4103 522 4132 532
rect 4146 522 4175 532
rect 4190 522 4220 536
rect 4263 522 4306 536
rect 4328 532 4518 544
rect 4583 540 4589 560
rect 4313 522 4343 532
rect 4344 522 4502 532
rect 4506 522 4536 532
rect 4540 522 4570 536
rect 4598 522 4611 560
rect 4683 574 4712 590
rect 4726 574 4755 590
rect 4770 580 4800 596
rect 4828 574 4834 622
rect 4837 616 4856 622
rect 4871 616 4901 624
rect 4837 608 4901 616
rect 4837 592 4917 608
rect 4933 601 4995 632
rect 5011 601 5073 632
rect 5142 630 5191 655
rect 5236 646 5262 656
rect 5206 630 5262 646
rect 5105 616 5135 624
rect 5142 622 5252 630
rect 5105 608 5150 616
rect 4837 590 4856 592
rect 4871 590 4917 592
rect 4837 574 4917 590
rect 4944 588 4979 601
rect 5020 598 5057 601
rect 5020 596 5062 598
rect 4949 585 4979 588
rect 4958 581 4965 585
rect 4965 580 4966 581
rect 4924 574 4934 580
rect 4683 566 4718 574
rect 4683 540 4684 566
rect 4691 540 4718 566
rect 4626 522 4656 536
rect 4683 532 4718 540
rect 4720 566 4761 574
rect 4720 540 4735 566
rect 4742 540 4761 566
rect 4825 562 4856 574
rect 4871 562 4974 574
rect 4986 564 5012 590
rect 5027 585 5057 596
rect 5089 592 5151 608
rect 5089 590 5135 592
rect 5089 574 5151 590
rect 5163 574 5169 622
rect 5172 614 5252 622
rect 5172 612 5191 614
rect 5206 612 5240 614
rect 5172 596 5252 612
rect 5172 574 5191 596
rect 5206 580 5236 596
rect 5264 590 5270 664
rect 5273 590 5292 734
rect 5307 590 5313 734
rect 5322 664 5335 734
rect 5387 730 5409 734
rect 5380 718 5397 722
rect 5401 720 5409 722
rect 5399 718 5409 720
rect 5380 708 5409 718
rect 5462 708 5478 722
rect 5516 718 5522 720
rect 5529 718 5637 734
rect 5644 718 5650 720
rect 5658 718 5673 734
rect 5739 728 5758 731
rect 5380 706 5478 708
rect 5505 706 5673 718
rect 5688 708 5704 722
rect 5739 709 5761 728
rect 5771 722 5787 723
rect 5770 720 5787 722
rect 5771 715 5787 720
rect 5761 708 5767 709
rect 5770 708 5799 715
rect 5688 707 5799 708
rect 5688 706 5805 707
rect 5364 698 5415 706
rect 5462 698 5496 706
rect 5364 686 5389 698
rect 5396 686 5415 698
rect 5469 696 5496 698
rect 5505 696 5726 706
rect 5761 703 5767 706
rect 5469 692 5726 696
rect 5364 678 5415 686
rect 5462 678 5726 692
rect 5770 698 5805 706
rect 5316 630 5335 664
rect 5380 670 5409 678
rect 5380 664 5397 670
rect 5380 662 5414 664
rect 5462 662 5478 678
rect 5479 668 5687 678
rect 5688 668 5704 678
rect 5752 674 5767 689
rect 5770 686 5771 698
rect 5778 686 5805 698
rect 5770 678 5805 686
rect 5770 677 5799 678
rect 5490 664 5704 668
rect 5505 662 5704 664
rect 5739 664 5752 674
rect 5770 664 5787 677
rect 5739 662 5787 664
rect 5381 658 5414 662
rect 5377 656 5414 658
rect 5377 655 5444 656
rect 5377 650 5408 655
rect 5414 650 5444 655
rect 5377 646 5444 650
rect 5350 643 5444 646
rect 5350 636 5399 643
rect 5350 630 5380 636
rect 5399 631 5404 636
rect 5316 614 5396 630
rect 5408 622 5444 643
rect 5505 638 5694 662
rect 5739 661 5786 662
rect 5752 656 5786 661
rect 5520 635 5694 638
rect 5513 632 5694 635
rect 5722 655 5786 656
rect 5316 612 5335 614
rect 5350 612 5384 614
rect 5316 596 5396 612
rect 5316 590 5335 596
rect 5032 564 5135 574
rect 4986 562 5135 564
rect 5156 562 5191 574
rect 4825 560 4987 562
rect 4837 540 4856 560
rect 4871 558 4901 560
rect 4720 532 4761 540
rect 4843 536 4856 540
rect 4908 544 4987 560
rect 5019 560 5191 562
rect 5019 544 5098 560
rect 5105 558 5135 560
rect 4683 522 4712 532
rect 4726 522 4755 532
rect 4770 522 4800 536
rect 4843 522 4886 536
rect 4908 532 5098 544
rect 5163 540 5169 560
rect 4893 522 4923 532
rect 4924 522 5082 532
rect 5086 522 5116 532
rect 5120 522 5150 536
rect 5178 522 5191 560
rect 5263 574 5292 590
rect 5306 574 5335 590
rect 5350 580 5380 596
rect 5408 574 5414 622
rect 5417 616 5436 622
rect 5451 616 5481 624
rect 5417 608 5481 616
rect 5417 592 5497 608
rect 5513 601 5575 632
rect 5591 601 5653 632
rect 5722 630 5771 655
rect 5786 630 5816 648
rect 5685 616 5715 624
rect 5722 622 5832 630
rect 5685 608 5730 616
rect 5417 590 5436 592
rect 5451 590 5497 592
rect 5417 574 5497 590
rect 5524 588 5559 601
rect 5600 598 5637 601
rect 5600 596 5642 598
rect 5529 585 5559 588
rect 5538 581 5545 585
rect 5545 580 5546 581
rect 5504 574 5514 580
rect 5263 566 5298 574
rect 5263 540 5264 566
rect 5271 540 5298 566
rect 5206 522 5236 536
rect 5263 532 5298 540
rect 5300 566 5341 574
rect 5300 540 5315 566
rect 5322 540 5341 566
rect 5405 562 5436 574
rect 5451 562 5554 574
rect 5566 564 5592 590
rect 5607 585 5637 596
rect 5669 592 5731 608
rect 5669 590 5715 592
rect 5669 574 5731 590
rect 5743 574 5749 622
rect 5752 614 5832 622
rect 5752 612 5771 614
rect 5786 612 5820 614
rect 5752 597 5832 612
rect 5752 596 5838 597
rect 5752 574 5771 596
rect 5786 580 5816 596
rect 5844 590 5850 664
rect 5853 590 5872 734
rect 5887 590 5893 734
rect 5902 664 5915 734
rect 5967 730 5989 734
rect 5960 718 5977 722
rect 5981 720 5989 722
rect 5979 718 5989 720
rect 5960 708 5989 718
rect 6042 708 6058 722
rect 6096 718 6102 720
rect 6109 718 6217 734
rect 6224 718 6230 720
rect 6238 718 6253 734
rect 6319 728 6338 731
rect 5960 706 6058 708
rect 6085 706 6253 718
rect 6268 708 6284 722
rect 6319 709 6341 728
rect 6351 722 6367 723
rect 6350 720 6367 722
rect 6351 715 6367 720
rect 6341 708 6347 709
rect 6350 708 6379 715
rect 6268 707 6379 708
rect 6268 706 6385 707
rect 5944 698 5995 706
rect 6042 698 6076 706
rect 5944 686 5969 698
rect 5976 686 5995 698
rect 6049 696 6076 698
rect 6085 696 6306 706
rect 6341 703 6347 706
rect 6049 692 6306 696
rect 5944 678 5995 686
rect 6042 678 6306 692
rect 6350 698 6385 706
rect 5896 630 5915 664
rect 5960 670 5989 678
rect 5960 664 5977 670
rect 5960 662 5994 664
rect 6042 662 6058 678
rect 6059 668 6267 678
rect 6268 668 6284 678
rect 6332 674 6347 689
rect 6350 686 6351 698
rect 6358 686 6385 698
rect 6350 678 6385 686
rect 6350 677 6379 678
rect 6070 664 6284 668
rect 6085 662 6284 664
rect 6319 664 6332 674
rect 6350 664 6367 677
rect 6319 662 6367 664
rect 5961 658 5994 662
rect 5957 656 5994 658
rect 5957 655 6024 656
rect 5957 650 5988 655
rect 5994 650 6024 655
rect 5957 646 6024 650
rect 5930 643 6024 646
rect 5930 636 5979 643
rect 5930 630 5960 636
rect 5979 631 5984 636
rect 5896 614 5976 630
rect 5988 622 6024 643
rect 6085 638 6274 662
rect 6319 661 6366 662
rect 6332 656 6366 661
rect 6100 635 6274 638
rect 6093 632 6274 635
rect 6302 655 6366 656
rect 5896 612 5915 614
rect 5930 612 5964 614
rect 5896 596 5976 612
rect 5896 590 5915 596
rect 5612 564 5715 574
rect 5566 562 5715 564
rect 5736 562 5771 574
rect 5405 560 5567 562
rect 5417 540 5436 560
rect 5451 558 5481 560
rect 5300 532 5341 540
rect 5423 536 5436 540
rect 5488 544 5567 560
rect 5599 560 5771 562
rect 5599 544 5678 560
rect 5685 558 5715 560
rect 5263 522 5292 532
rect 5306 522 5335 532
rect 5350 522 5380 536
rect 5423 522 5466 536
rect 5488 532 5678 544
rect 5743 540 5749 560
rect 5473 522 5503 532
rect 5504 522 5662 532
rect 5666 522 5696 532
rect 5700 522 5730 536
rect 5758 522 5771 560
rect 5843 574 5872 590
rect 5886 574 5915 590
rect 5930 580 5960 596
rect 5988 574 5994 622
rect 5997 616 6016 622
rect 6031 616 6061 624
rect 5997 608 6061 616
rect 5997 592 6077 608
rect 6093 601 6155 632
rect 6171 601 6233 632
rect 6302 630 6351 655
rect 6366 630 6396 646
rect 6265 616 6295 624
rect 6302 622 6412 630
rect 6265 608 6310 616
rect 5997 590 6016 592
rect 6031 590 6077 592
rect 5997 574 6077 590
rect 6104 588 6139 601
rect 6180 598 6217 601
rect 6180 596 6222 598
rect 6109 585 6139 588
rect 6118 581 6125 585
rect 6125 580 6126 581
rect 6084 574 6094 580
rect 5843 566 5878 574
rect 5843 540 5844 566
rect 5851 540 5878 566
rect 5786 522 5816 536
rect 5843 532 5878 540
rect 5880 566 5921 574
rect 5880 540 5895 566
rect 5902 540 5921 566
rect 5985 562 6016 574
rect 6031 562 6134 574
rect 6146 564 6172 590
rect 6187 585 6217 596
rect 6249 592 6311 608
rect 6249 590 6295 592
rect 6249 574 6311 590
rect 6323 574 6329 622
rect 6332 614 6412 622
rect 6332 612 6351 614
rect 6366 612 6400 614
rect 6332 596 6412 612
rect 6332 574 6351 596
rect 6366 580 6396 596
rect 6424 590 6430 664
rect 6439 590 6452 734
rect 6192 564 6295 574
rect 6146 562 6295 564
rect 6316 562 6351 574
rect 5985 560 6147 562
rect 5997 540 6016 560
rect 6031 558 6061 560
rect 5880 532 5921 540
rect 6003 536 6016 540
rect 6068 544 6147 560
rect 6179 560 6351 562
rect 6179 544 6258 560
rect 6265 558 6295 560
rect 5843 522 5872 532
rect 5886 522 5915 532
rect 5930 522 5960 536
rect 6003 522 6046 536
rect 6068 532 6258 544
rect 6323 540 6329 560
rect 6053 522 6083 532
rect 6084 522 6242 532
rect 6246 522 6276 532
rect 6280 522 6310 536
rect 6338 522 6351 560
rect 6423 574 6452 590
rect 6423 566 6458 574
rect 6423 540 6424 566
rect 6431 540 6458 566
rect 6366 522 6396 536
rect 6423 532 6458 540
rect 6423 522 6452 532
rect -541 508 6452 522
rect -478 478 -465 508
rect -450 494 -420 508
rect -377 494 -334 508
rect -327 494 -107 508
rect -100 494 -70 508
rect -410 480 -395 492
rect -376 480 -363 494
rect -295 490 -142 494
rect -413 478 -391 480
rect -313 478 -121 490
rect -42 478 -29 508
rect -14 494 16 508
rect 53 478 72 508
rect 87 478 93 508
rect 102 478 115 508
rect 130 494 160 508
rect 203 494 246 508
rect 253 494 473 508
rect 480 494 510 508
rect 170 480 185 492
rect 204 480 217 494
rect 285 490 438 494
rect 167 478 189 480
rect 267 478 459 490
rect 538 478 551 508
rect 566 494 596 508
rect 633 478 652 508
rect 667 478 673 508
rect 682 478 695 508
rect 710 494 740 508
rect 783 494 826 508
rect 833 494 1053 508
rect 1060 494 1090 508
rect 750 480 765 492
rect 784 480 797 494
rect 865 490 1018 494
rect 747 478 769 480
rect 847 478 1039 490
rect 1118 478 1131 508
rect 1146 494 1176 508
rect 1213 478 1232 508
rect 1247 478 1253 508
rect 1262 478 1275 508
rect 1290 494 1320 508
rect 1363 494 1406 508
rect 1413 494 1633 508
rect 1640 494 1670 508
rect 1330 480 1345 492
rect 1364 480 1377 494
rect 1445 490 1598 494
rect 1327 478 1349 480
rect 1427 478 1619 490
rect 1698 478 1711 508
rect 1726 494 1756 508
rect 1793 478 1812 508
rect 1827 478 1833 508
rect 1842 478 1855 508
rect 1870 494 1900 508
rect 1943 494 1986 508
rect 1993 494 2213 508
rect 2220 494 2250 508
rect 1910 480 1925 492
rect 1944 480 1957 494
rect 2025 490 2178 494
rect 1907 478 1929 480
rect 2007 478 2199 490
rect 2278 478 2291 508
rect 2306 494 2336 508
rect 2373 478 2392 508
rect 2407 478 2413 508
rect 2422 478 2435 508
rect 2450 494 2480 508
rect 2523 494 2566 508
rect 2573 494 2793 508
rect 2800 494 2830 508
rect 2490 480 2505 492
rect 2524 480 2537 494
rect 2605 490 2758 494
rect 2487 478 2509 480
rect 2587 478 2779 490
rect 2858 478 2871 508
rect 2886 494 2916 508
rect 2953 478 2972 508
rect 2987 478 2993 508
rect 3002 478 3015 508
rect 3030 494 3060 508
rect 3103 494 3146 508
rect 3153 494 3373 508
rect 3380 494 3410 508
rect 3070 480 3085 492
rect 3104 480 3117 494
rect 3185 490 3338 494
rect 3067 478 3089 480
rect 3167 478 3359 490
rect 3438 478 3451 508
rect 3466 494 3496 508
rect 3533 478 3552 508
rect 3567 478 3573 508
rect 3582 478 3595 508
rect 3610 494 3640 508
rect 3683 494 3726 508
rect 3733 494 3953 508
rect 3960 494 3990 508
rect 3650 480 3665 492
rect 3684 480 3697 494
rect 3765 490 3918 494
rect 3647 478 3669 480
rect 3747 478 3939 490
rect 4018 478 4031 508
rect 4046 494 4076 508
rect 4113 478 4132 508
rect 4147 478 4153 508
rect 4162 478 4175 508
rect 4190 494 4220 508
rect 4263 494 4306 508
rect 4313 494 4533 508
rect 4540 494 4570 508
rect 4230 480 4245 492
rect 4264 480 4277 494
rect 4345 490 4498 494
rect 4227 478 4249 480
rect 4327 478 4519 490
rect 4598 478 4611 508
rect 4626 494 4656 508
rect 4693 478 4712 508
rect 4727 478 4733 508
rect 4742 478 4755 508
rect 4770 494 4800 508
rect 4843 494 4886 508
rect 4893 494 5113 508
rect 5120 494 5150 508
rect 4810 480 4825 492
rect 4844 480 4857 494
rect 4925 490 5078 494
rect 4807 478 4829 480
rect 4907 478 5099 490
rect 5178 478 5191 508
rect 5206 494 5236 508
rect 5273 478 5292 508
rect 5307 478 5313 508
rect 5322 478 5335 508
rect 5350 494 5380 508
rect 5423 494 5466 508
rect 5473 494 5693 508
rect 5700 494 5730 508
rect 5390 480 5405 492
rect 5424 480 5437 494
rect 5505 490 5658 494
rect 5387 478 5409 480
rect 5487 478 5679 490
rect 5758 478 5771 508
rect 5786 494 5816 508
rect 5853 478 5872 508
rect 5887 478 5893 508
rect 5902 478 5915 508
rect 5930 494 5960 508
rect 6003 494 6046 508
rect 6053 494 6273 508
rect 6280 494 6310 508
rect 5970 480 5985 492
rect 6004 480 6017 494
rect 6085 490 6238 494
rect 5967 478 5989 480
rect 6067 478 6259 490
rect 6338 478 6351 508
rect 6366 494 6396 508
rect 6439 478 6452 508
rect -541 464 6452 478
rect -478 394 -465 464
rect -413 460 -391 464
rect -420 448 -403 452
rect -399 450 -391 452
rect -401 448 -391 450
rect -420 438 -391 448
rect -338 438 -322 452
rect -284 448 -278 450
rect -271 448 -163 464
rect -156 448 -150 450
rect -142 448 -127 464
rect -61 458 -42 461
rect -420 436 -322 438
rect -295 436 -127 448
rect -112 438 -96 452
rect -61 439 -39 458
rect -29 452 -13 453
rect -30 450 -13 452
rect -29 445 -13 450
rect -39 438 -33 439
rect -30 438 -1 445
rect -112 437 -1 438
rect -112 436 5 437
rect -436 428 -385 436
rect -338 428 -304 436
rect -436 416 -411 428
rect -404 416 -385 428
rect -331 426 -304 428
rect -295 426 -74 436
rect -39 433 -33 436
rect -331 422 -74 426
rect -436 408 -385 416
rect -338 408 -74 422
rect -30 428 5 436
rect -484 360 -465 394
rect -420 400 -391 408
rect -420 394 -403 400
rect -420 392 -386 394
rect -338 392 -322 408
rect -321 398 -113 408
rect -112 398 -96 408
rect -48 404 -33 419
rect -30 416 -29 428
rect -22 416 5 428
rect -30 408 5 416
rect -30 407 -1 408
rect -310 394 -96 398
rect -295 392 -96 394
rect -61 394 -48 404
rect -30 394 -13 407
rect -61 392 -13 394
rect -419 388 -386 392
rect -423 386 -386 388
rect -423 385 -356 386
rect -423 380 -392 385
rect -386 380 -356 385
rect -423 376 -356 380
rect -450 373 -356 376
rect -450 366 -401 373
rect -450 360 -420 366
rect -401 361 -396 366
rect -484 344 -404 360
rect -392 352 -356 373
rect -295 368 -106 392
rect -61 391 -14 392
rect -48 386 -14 391
rect -280 365 -106 368
rect -287 362 -106 365
rect -78 385 -14 386
rect -484 342 -465 344
rect -450 342 -416 344
rect -484 326 -404 342
rect -484 320 -465 326
rect -494 304 -465 320
rect -450 310 -420 326
rect -392 304 -386 352
rect -383 346 -364 352
rect -349 346 -319 354
rect -383 338 -319 346
rect -383 322 -303 338
rect -287 331 -225 362
rect -209 331 -147 362
rect -78 360 -29 385
rect -14 360 16 378
rect -115 346 -85 354
rect -78 352 32 360
rect -115 338 -70 346
rect -383 320 -364 322
rect -349 320 -303 322
rect -383 304 -303 320
rect -276 318 -241 331
rect -200 328 -163 331
rect -200 326 -158 328
rect -271 315 -241 318
rect -262 311 -255 315
rect -255 310 -254 311
rect -296 304 -286 310
rect -500 296 -459 304
rect -500 270 -485 296
rect -478 270 -459 296
rect -395 292 -364 304
rect -349 292 -246 304
rect -234 294 -208 320
rect -193 315 -163 326
rect -131 322 -69 338
rect -131 320 -85 322
rect -131 304 -69 320
rect -57 304 -51 352
rect -48 344 32 352
rect -48 342 -29 344
rect -14 342 20 344
rect -48 327 32 342
rect -48 326 38 327
rect -48 304 -29 326
rect -14 310 16 326
rect 44 320 50 394
rect 53 320 72 464
rect 87 320 93 464
rect 102 394 115 464
rect 167 460 189 464
rect 160 448 177 452
rect 181 450 189 452
rect 179 448 189 450
rect 160 438 189 448
rect 242 438 258 452
rect 296 448 302 450
rect 309 448 417 464
rect 424 448 430 450
rect 438 448 453 464
rect 519 458 538 461
rect 160 436 258 438
rect 285 436 453 448
rect 468 438 484 452
rect 519 439 541 458
rect 551 452 567 453
rect 550 450 567 452
rect 551 445 567 450
rect 541 438 547 439
rect 550 438 579 445
rect 468 437 579 438
rect 468 436 585 437
rect 144 428 195 436
rect 242 428 276 436
rect 144 416 169 428
rect 176 416 195 428
rect 249 426 276 428
rect 285 426 506 436
rect 541 433 547 436
rect 249 422 506 426
rect 144 408 195 416
rect 242 408 506 422
rect 550 428 585 436
rect 96 360 115 394
rect 160 400 189 408
rect 160 394 177 400
rect 160 392 194 394
rect 242 392 258 408
rect 259 398 467 408
rect 468 398 484 408
rect 532 404 547 419
rect 550 416 551 428
rect 558 416 585 428
rect 550 408 585 416
rect 550 407 579 408
rect 270 394 484 398
rect 285 392 484 394
rect 519 394 532 404
rect 550 394 567 407
rect 519 392 567 394
rect 161 388 194 392
rect 157 386 194 388
rect 157 385 224 386
rect 157 380 188 385
rect 194 380 224 385
rect 157 376 224 380
rect 130 373 224 376
rect 130 366 179 373
rect 130 360 160 366
rect 179 361 184 366
rect 96 344 176 360
rect 188 352 224 373
rect 285 368 474 392
rect 519 391 566 392
rect 532 386 566 391
rect 606 386 622 388
rect 300 365 474 368
rect 293 362 474 365
rect 502 385 566 386
rect 96 342 115 344
rect 130 342 164 344
rect 96 326 176 342
rect 96 320 115 326
rect -188 294 -85 304
rect -234 292 -85 294
rect -64 292 -29 304
rect -395 290 -233 292
rect -383 272 -364 290
rect -349 288 -319 290
rect -500 262 -459 270
rect -376 266 -364 272
rect -312 274 -233 290
rect -201 290 -29 292
rect -201 274 -122 290
rect -115 288 -85 290
rect -494 252 -465 262
rect -450 252 -420 266
rect -376 252 -334 266
rect -312 262 -122 274
rect -57 270 -51 290
rect -327 252 -297 262
rect -296 252 -138 262
rect -134 252 -104 262
rect -100 252 -70 266
rect -42 252 -29 290
rect 43 304 72 320
rect 86 304 115 320
rect 130 310 160 326
rect 188 304 194 352
rect 197 346 216 352
rect 231 346 261 354
rect 197 338 261 346
rect 197 322 277 338
rect 293 331 355 362
rect 371 331 433 362
rect 502 360 551 385
rect 596 376 622 386
rect 566 360 622 376
rect 465 346 495 354
rect 502 352 612 360
rect 465 338 510 346
rect 197 320 216 322
rect 231 320 277 322
rect 197 304 277 320
rect 304 318 339 331
rect 380 328 417 331
rect 380 326 422 328
rect 309 315 339 318
rect 318 311 325 315
rect 325 310 326 311
rect 284 304 294 310
rect 43 296 78 304
rect 43 270 44 296
rect 51 270 78 296
rect -14 252 16 266
rect 43 262 78 270
rect 80 296 121 304
rect 80 270 95 296
rect 102 270 121 296
rect 185 292 216 304
rect 231 292 334 304
rect 346 294 372 320
rect 387 315 417 326
rect 449 322 511 338
rect 449 320 495 322
rect 449 304 511 320
rect 523 304 529 352
rect 532 344 612 352
rect 532 342 551 344
rect 566 342 600 344
rect 532 326 612 342
rect 532 304 551 326
rect 566 310 596 326
rect 624 320 630 394
rect 633 320 652 464
rect 667 320 673 464
rect 682 394 695 464
rect 747 460 769 464
rect 740 448 757 452
rect 761 450 769 452
rect 759 448 769 450
rect 740 438 769 448
rect 822 438 838 452
rect 876 448 882 450
rect 889 448 997 464
rect 1004 448 1010 450
rect 1018 448 1033 464
rect 1099 458 1118 461
rect 740 436 838 438
rect 865 436 1033 448
rect 1048 438 1064 452
rect 1099 439 1121 458
rect 1131 452 1147 453
rect 1130 450 1147 452
rect 1131 445 1147 450
rect 1121 438 1127 439
rect 1130 438 1159 445
rect 1048 437 1159 438
rect 1048 436 1165 437
rect 724 428 775 436
rect 822 428 856 436
rect 724 416 749 428
rect 756 416 775 428
rect 829 426 856 428
rect 865 426 1086 436
rect 1121 433 1127 436
rect 829 422 1086 426
rect 724 408 775 416
rect 822 408 1086 422
rect 1130 428 1165 436
rect 676 360 695 394
rect 740 400 769 408
rect 740 394 757 400
rect 740 392 774 394
rect 822 392 838 408
rect 839 398 1047 408
rect 1048 398 1064 408
rect 1112 404 1127 419
rect 1130 416 1131 428
rect 1138 416 1165 428
rect 1130 408 1165 416
rect 1130 407 1159 408
rect 850 394 1064 398
rect 865 392 1064 394
rect 1099 394 1112 404
rect 1130 394 1147 407
rect 1099 392 1147 394
rect 741 388 774 392
rect 737 386 774 388
rect 737 385 804 386
rect 737 380 768 385
rect 774 380 804 385
rect 737 376 804 380
rect 710 373 804 376
rect 710 366 759 373
rect 710 360 740 366
rect 759 361 764 366
rect 676 344 756 360
rect 768 352 804 373
rect 865 368 1054 392
rect 1099 391 1146 392
rect 1112 386 1146 391
rect 880 365 1054 368
rect 873 362 1054 365
rect 1082 385 1146 386
rect 676 342 695 344
rect 710 342 744 344
rect 676 326 756 342
rect 676 320 695 326
rect 392 294 495 304
rect 346 292 495 294
rect 516 292 551 304
rect 185 290 347 292
rect 197 272 216 290
rect 231 288 261 290
rect 80 262 121 270
rect 204 266 216 272
rect 268 274 347 290
rect 379 290 551 292
rect 379 274 458 290
rect 465 288 495 290
rect 43 252 72 262
rect 86 252 115 262
rect 130 252 160 266
rect 204 252 246 266
rect 268 262 458 274
rect 523 270 529 290
rect 253 252 283 262
rect 284 252 442 262
rect 446 252 476 262
rect 480 252 510 266
rect 538 252 551 290
rect 623 304 652 320
rect 666 304 695 320
rect 710 310 740 326
rect 768 304 774 352
rect 777 346 796 352
rect 811 346 841 354
rect 777 338 841 346
rect 777 322 857 338
rect 873 331 935 362
rect 951 331 1013 362
rect 1082 360 1131 385
rect 1146 360 1176 378
rect 1045 346 1075 354
rect 1082 352 1192 360
rect 1045 338 1090 346
rect 777 320 796 322
rect 811 320 857 322
rect 777 304 857 320
rect 884 318 919 331
rect 960 328 997 331
rect 960 326 1002 328
rect 889 315 919 318
rect 898 311 905 315
rect 905 310 906 311
rect 864 304 874 310
rect 623 296 658 304
rect 623 270 624 296
rect 631 270 658 296
rect 566 252 596 266
rect 623 262 658 270
rect 660 296 701 304
rect 660 270 675 296
rect 682 270 701 296
rect 765 292 796 304
rect 811 292 914 304
rect 926 294 952 320
rect 967 315 997 326
rect 1029 322 1091 338
rect 1029 320 1075 322
rect 1029 304 1091 320
rect 1103 304 1109 352
rect 1112 344 1192 352
rect 1112 342 1131 344
rect 1146 342 1180 344
rect 1112 327 1192 342
rect 1112 326 1198 327
rect 1112 304 1131 326
rect 1146 310 1176 326
rect 1204 320 1210 394
rect 1213 320 1232 464
rect 1247 320 1253 464
rect 1262 394 1275 464
rect 1327 460 1349 464
rect 1320 448 1337 452
rect 1341 450 1349 452
rect 1339 448 1349 450
rect 1320 438 1349 448
rect 1402 438 1418 452
rect 1456 448 1462 450
rect 1469 448 1577 464
rect 1584 448 1590 450
rect 1598 448 1613 464
rect 1679 458 1698 461
rect 1320 436 1418 438
rect 1445 436 1613 448
rect 1628 438 1644 452
rect 1679 439 1701 458
rect 1711 452 1727 453
rect 1710 450 1727 452
rect 1711 445 1727 450
rect 1701 438 1707 439
rect 1710 438 1739 445
rect 1628 437 1739 438
rect 1628 436 1745 437
rect 1304 428 1355 436
rect 1402 428 1436 436
rect 1304 416 1329 428
rect 1336 416 1355 428
rect 1409 426 1436 428
rect 1445 426 1666 436
rect 1701 433 1707 436
rect 1409 422 1666 426
rect 1304 408 1355 416
rect 1402 408 1666 422
rect 1710 428 1745 436
rect 1256 360 1275 394
rect 1320 400 1349 408
rect 1320 394 1337 400
rect 1320 392 1354 394
rect 1402 392 1418 408
rect 1419 398 1627 408
rect 1628 398 1644 408
rect 1692 404 1707 419
rect 1710 416 1711 428
rect 1718 416 1745 428
rect 1710 408 1745 416
rect 1710 407 1739 408
rect 1430 394 1644 398
rect 1445 392 1644 394
rect 1679 394 1692 404
rect 1710 394 1727 407
rect 1679 392 1727 394
rect 1321 388 1354 392
rect 1317 386 1354 388
rect 1317 385 1384 386
rect 1317 380 1348 385
rect 1354 380 1384 385
rect 1317 376 1384 380
rect 1290 373 1384 376
rect 1290 366 1339 373
rect 1290 360 1320 366
rect 1339 361 1344 366
rect 1256 344 1336 360
rect 1348 352 1384 373
rect 1445 368 1634 392
rect 1679 391 1726 392
rect 1692 386 1726 391
rect 1766 386 1782 388
rect 1460 365 1634 368
rect 1453 362 1634 365
rect 1662 385 1726 386
rect 1256 342 1275 344
rect 1290 342 1324 344
rect 1256 326 1336 342
rect 1256 320 1275 326
rect 972 294 1075 304
rect 926 292 1075 294
rect 1096 292 1131 304
rect 765 290 927 292
rect 777 272 796 290
rect 811 288 841 290
rect 660 262 701 270
rect 784 266 796 272
rect 848 272 927 290
rect 959 290 1131 292
rect 959 274 1038 290
rect 1045 288 1075 290
rect 934 272 1038 274
rect 623 252 652 262
rect 666 252 695 262
rect 710 252 740 266
rect 784 252 826 266
rect 848 262 1038 272
rect 1103 270 1109 290
rect 833 252 863 262
rect 864 252 1022 262
rect 1026 252 1056 262
rect 1060 252 1090 266
rect 1118 252 1131 290
rect 1203 304 1232 320
rect 1246 304 1275 320
rect 1290 310 1320 326
rect 1348 304 1354 352
rect 1357 346 1376 352
rect 1391 346 1421 354
rect 1357 338 1421 346
rect 1357 322 1437 338
rect 1453 331 1515 362
rect 1531 331 1593 362
rect 1662 360 1711 385
rect 1756 376 1782 386
rect 1726 360 1782 376
rect 1625 346 1655 354
rect 1662 352 1772 360
rect 1625 338 1670 346
rect 1357 320 1376 322
rect 1391 320 1437 322
rect 1357 304 1437 320
rect 1464 318 1499 331
rect 1540 328 1577 331
rect 1540 326 1582 328
rect 1469 315 1499 318
rect 1478 311 1485 315
rect 1485 310 1486 311
rect 1444 304 1454 310
rect 1203 296 1238 304
rect 1203 270 1204 296
rect 1211 270 1238 296
rect 1146 252 1176 266
rect 1203 262 1238 270
rect 1240 296 1281 304
rect 1240 270 1255 296
rect 1262 270 1281 296
rect 1345 292 1376 304
rect 1391 292 1494 304
rect 1506 294 1532 320
rect 1547 315 1577 326
rect 1609 322 1671 338
rect 1609 320 1655 322
rect 1609 304 1671 320
rect 1683 304 1689 352
rect 1692 344 1772 352
rect 1692 342 1711 344
rect 1726 342 1760 344
rect 1692 326 1772 342
rect 1692 304 1711 326
rect 1726 310 1756 326
rect 1784 320 1790 394
rect 1793 320 1812 464
rect 1827 320 1833 464
rect 1842 394 1855 464
rect 1907 460 1929 464
rect 1900 448 1917 452
rect 1921 450 1929 452
rect 1919 448 1929 450
rect 1900 438 1929 448
rect 1982 438 1998 452
rect 2036 448 2042 450
rect 2049 448 2157 464
rect 2164 448 2170 450
rect 2178 448 2193 464
rect 2259 458 2278 461
rect 1900 436 1998 438
rect 2025 436 2193 448
rect 2208 438 2224 452
rect 2259 439 2281 458
rect 2291 452 2307 453
rect 2290 450 2307 452
rect 2291 445 2307 450
rect 2281 438 2287 439
rect 2290 438 2319 445
rect 2208 437 2319 438
rect 2208 436 2325 437
rect 1884 428 1935 436
rect 1982 428 2016 436
rect 1884 416 1909 428
rect 1916 416 1935 428
rect 1989 426 2016 428
rect 2025 426 2246 436
rect 2281 433 2287 436
rect 1989 422 2246 426
rect 1884 408 1935 416
rect 1982 408 2246 422
rect 2290 428 2325 436
rect 1836 360 1855 394
rect 1900 400 1929 408
rect 1900 394 1917 400
rect 1900 392 1934 394
rect 1982 392 1998 408
rect 1999 398 2207 408
rect 2208 398 2224 408
rect 2272 404 2287 419
rect 2290 416 2291 428
rect 2298 416 2325 428
rect 2290 408 2325 416
rect 2290 407 2319 408
rect 2010 394 2224 398
rect 2025 392 2224 394
rect 2259 394 2272 404
rect 2290 394 2307 407
rect 2259 392 2307 394
rect 1901 388 1934 392
rect 1897 386 1934 388
rect 1897 385 1964 386
rect 1897 380 1928 385
rect 1934 380 1964 385
rect 1897 376 1964 380
rect 1870 373 1964 376
rect 1870 366 1919 373
rect 1870 360 1900 366
rect 1919 361 1924 366
rect 1836 344 1916 360
rect 1928 352 1964 373
rect 2025 368 2214 392
rect 2259 391 2306 392
rect 2272 386 2306 391
rect 2040 365 2214 368
rect 2033 362 2214 365
rect 2242 385 2306 386
rect 1836 342 1855 344
rect 1870 342 1904 344
rect 1836 326 1916 342
rect 1836 320 1855 326
rect 1552 294 1655 304
rect 1506 292 1655 294
rect 1676 292 1711 304
rect 1345 290 1507 292
rect 1357 272 1376 290
rect 1391 288 1421 290
rect 1240 262 1281 270
rect 1364 266 1376 272
rect 1428 272 1507 290
rect 1539 290 1711 292
rect 1539 274 1618 290
rect 1625 288 1655 290
rect 1514 272 1618 274
rect 1203 252 1232 262
rect 1246 252 1275 262
rect 1290 252 1320 266
rect 1364 252 1406 266
rect 1428 262 1618 272
rect 1683 270 1689 290
rect 1413 252 1443 262
rect 1444 252 1602 262
rect 1606 252 1636 262
rect 1640 252 1670 266
rect 1698 252 1711 290
rect 1783 304 1812 320
rect 1826 304 1855 320
rect 1870 310 1900 326
rect 1928 304 1934 352
rect 1937 346 1956 352
rect 1971 346 2001 354
rect 1937 338 2001 346
rect 1937 322 2017 338
rect 2033 331 2095 362
rect 2111 331 2173 362
rect 2242 360 2291 385
rect 2306 360 2336 378
rect 2205 346 2235 354
rect 2242 352 2352 360
rect 2205 338 2250 346
rect 1937 320 1956 322
rect 1971 320 2017 322
rect 1937 304 2017 320
rect 2044 318 2079 331
rect 2120 328 2157 331
rect 2120 326 2162 328
rect 2049 315 2079 318
rect 2058 311 2065 315
rect 2065 310 2066 311
rect 2024 304 2034 310
rect 1783 296 1818 304
rect 1783 270 1784 296
rect 1791 270 1818 296
rect 1726 252 1756 266
rect 1783 262 1818 270
rect 1820 296 1861 304
rect 1820 270 1835 296
rect 1842 270 1861 296
rect 1925 292 1956 304
rect 1971 292 2074 304
rect 2086 294 2112 320
rect 2127 315 2157 326
rect 2189 322 2251 338
rect 2189 320 2235 322
rect 2189 304 2251 320
rect 2263 304 2269 352
rect 2272 344 2352 352
rect 2272 342 2291 344
rect 2306 342 2340 344
rect 2272 327 2352 342
rect 2272 326 2358 327
rect 2272 304 2291 326
rect 2306 310 2336 326
rect 2364 320 2370 394
rect 2373 320 2392 464
rect 2407 320 2413 464
rect 2422 394 2435 464
rect 2487 460 2509 464
rect 2480 448 2497 452
rect 2501 450 2509 452
rect 2499 448 2509 450
rect 2480 438 2509 448
rect 2562 438 2578 452
rect 2616 448 2622 450
rect 2629 448 2737 464
rect 2744 448 2750 450
rect 2758 448 2773 464
rect 2839 458 2858 461
rect 2480 436 2578 438
rect 2605 436 2773 448
rect 2788 438 2804 452
rect 2839 439 2861 458
rect 2871 452 2887 453
rect 2870 450 2887 452
rect 2871 445 2887 450
rect 2861 438 2867 439
rect 2870 438 2899 445
rect 2788 437 2899 438
rect 2788 436 2905 437
rect 2464 428 2515 436
rect 2562 428 2596 436
rect 2464 416 2489 428
rect 2496 416 2515 428
rect 2569 426 2596 428
rect 2605 426 2826 436
rect 2861 433 2867 436
rect 2569 422 2826 426
rect 2464 408 2515 416
rect 2562 408 2826 422
rect 2870 428 2905 436
rect 2416 360 2435 394
rect 2480 400 2509 408
rect 2480 394 2497 400
rect 2480 392 2514 394
rect 2562 392 2578 408
rect 2579 398 2787 408
rect 2788 398 2804 408
rect 2852 404 2867 419
rect 2870 416 2871 428
rect 2878 416 2905 428
rect 2870 408 2905 416
rect 2870 407 2899 408
rect 2590 394 2804 398
rect 2605 392 2804 394
rect 2839 394 2852 404
rect 2870 394 2887 407
rect 2839 392 2887 394
rect 2481 388 2514 392
rect 2477 386 2514 388
rect 2477 385 2544 386
rect 2477 380 2508 385
rect 2514 380 2544 385
rect 2477 376 2544 380
rect 2450 373 2544 376
rect 2450 366 2499 373
rect 2450 360 2480 366
rect 2499 361 2504 366
rect 2416 344 2496 360
rect 2508 352 2544 373
rect 2605 368 2794 392
rect 2839 391 2886 392
rect 2852 386 2886 391
rect 2926 386 2942 388
rect 2620 365 2794 368
rect 2613 362 2794 365
rect 2822 385 2886 386
rect 2416 342 2435 344
rect 2450 342 2484 344
rect 2416 326 2496 342
rect 2416 320 2435 326
rect 2132 294 2235 304
rect 2086 292 2235 294
rect 2256 292 2291 304
rect 1925 290 2087 292
rect 1937 272 1956 290
rect 1971 288 2001 290
rect 1820 262 1861 270
rect 1944 266 1956 272
rect 2008 274 2087 290
rect 2119 290 2291 292
rect 2119 274 2198 290
rect 2205 288 2235 290
rect 1783 252 1812 262
rect 1826 252 1855 262
rect 1870 252 1900 266
rect 1944 252 1986 266
rect 2008 262 2198 274
rect 2263 270 2269 290
rect 1993 252 2023 262
rect 2024 252 2182 262
rect 2186 252 2216 262
rect 2220 252 2250 266
rect 2278 252 2291 290
rect 2363 304 2392 320
rect 2406 304 2435 320
rect 2450 310 2480 326
rect 2508 304 2514 352
rect 2517 346 2536 352
rect 2551 346 2581 354
rect 2517 338 2581 346
rect 2517 322 2597 338
rect 2613 331 2675 362
rect 2691 331 2753 362
rect 2822 360 2871 385
rect 2916 376 2942 386
rect 2886 360 2942 376
rect 2785 346 2815 354
rect 2822 352 2932 360
rect 2785 338 2830 346
rect 2517 320 2536 322
rect 2551 320 2597 322
rect 2517 304 2597 320
rect 2624 318 2659 331
rect 2700 328 2737 331
rect 2700 326 2742 328
rect 2629 315 2659 318
rect 2638 311 2645 315
rect 2645 310 2646 311
rect 2604 304 2614 310
rect 2363 296 2398 304
rect 2363 270 2364 296
rect 2371 270 2398 296
rect 2306 252 2336 266
rect 2363 262 2398 270
rect 2400 296 2441 304
rect 2400 270 2415 296
rect 2422 270 2441 296
rect 2505 292 2536 304
rect 2551 292 2654 304
rect 2666 294 2692 320
rect 2707 315 2737 326
rect 2769 322 2831 338
rect 2769 320 2815 322
rect 2769 304 2831 320
rect 2843 304 2849 352
rect 2852 344 2932 352
rect 2852 342 2871 344
rect 2886 342 2920 344
rect 2852 326 2932 342
rect 2852 304 2871 326
rect 2886 310 2916 326
rect 2944 320 2950 394
rect 2953 320 2972 464
rect 2987 320 2993 464
rect 3002 394 3015 464
rect 3067 460 3089 464
rect 3060 448 3077 452
rect 3081 450 3089 452
rect 3079 448 3089 450
rect 3060 438 3089 448
rect 3142 438 3158 452
rect 3196 448 3202 450
rect 3209 448 3317 464
rect 3324 448 3330 450
rect 3338 448 3353 464
rect 3419 458 3438 461
rect 3060 436 3158 438
rect 3185 436 3353 448
rect 3368 438 3384 452
rect 3419 439 3441 458
rect 3451 452 3467 453
rect 3450 450 3467 452
rect 3451 445 3467 450
rect 3441 438 3447 439
rect 3450 438 3479 445
rect 3368 437 3479 438
rect 3368 436 3485 437
rect 3044 428 3095 436
rect 3142 428 3176 436
rect 3044 416 3069 428
rect 3076 416 3095 428
rect 3149 426 3176 428
rect 3185 426 3406 436
rect 3441 433 3447 436
rect 3149 422 3406 426
rect 3044 408 3095 416
rect 3142 408 3406 422
rect 3450 428 3485 436
rect 2996 360 3015 394
rect 3060 400 3089 408
rect 3060 394 3077 400
rect 3060 392 3094 394
rect 3142 392 3158 408
rect 3159 398 3367 408
rect 3368 398 3384 408
rect 3432 404 3447 419
rect 3450 416 3451 428
rect 3458 416 3485 428
rect 3450 408 3485 416
rect 3450 407 3479 408
rect 3170 394 3384 398
rect 3185 392 3384 394
rect 3419 394 3432 404
rect 3450 394 3467 407
rect 3419 392 3467 394
rect 3061 388 3094 392
rect 3057 386 3094 388
rect 3057 385 3124 386
rect 3057 380 3088 385
rect 3094 380 3124 385
rect 3057 376 3124 380
rect 3030 373 3124 376
rect 3030 366 3079 373
rect 3030 360 3060 366
rect 3079 361 3084 366
rect 2996 344 3076 360
rect 3088 352 3124 373
rect 3185 368 3374 392
rect 3419 391 3466 392
rect 3432 386 3466 391
rect 3200 365 3374 368
rect 3193 362 3374 365
rect 3402 385 3466 386
rect 2996 342 3015 344
rect 3030 342 3064 344
rect 2996 326 3076 342
rect 2996 320 3015 326
rect 2712 294 2815 304
rect 2666 292 2815 294
rect 2836 292 2871 304
rect 2505 290 2667 292
rect 2517 272 2536 290
rect 2551 288 2581 290
rect 2400 262 2441 270
rect 2524 266 2536 272
rect 2588 274 2667 290
rect 2699 290 2871 292
rect 2699 274 2778 290
rect 2785 288 2815 290
rect 2363 252 2392 262
rect 2406 252 2435 262
rect 2450 252 2480 266
rect 2524 252 2566 266
rect 2588 262 2778 274
rect 2843 270 2849 290
rect 2573 252 2603 262
rect 2604 252 2762 262
rect 2766 252 2796 262
rect 2800 252 2830 266
rect 2858 252 2871 290
rect 2943 304 2972 320
rect 2986 304 3015 320
rect 3030 310 3060 326
rect 3088 304 3094 352
rect 3097 346 3116 352
rect 3131 346 3161 354
rect 3097 338 3161 346
rect 3097 322 3177 338
rect 3193 331 3255 362
rect 3271 331 3333 362
rect 3402 360 3451 385
rect 3466 360 3496 378
rect 3365 346 3395 354
rect 3402 352 3512 360
rect 3365 338 3410 346
rect 3097 320 3116 322
rect 3131 320 3177 322
rect 3097 304 3177 320
rect 3204 318 3239 331
rect 3280 328 3317 331
rect 3280 326 3322 328
rect 3209 315 3239 318
rect 3218 311 3225 315
rect 3225 310 3226 311
rect 3184 304 3194 310
rect 2943 296 2978 304
rect 2943 270 2944 296
rect 2951 270 2978 296
rect 2886 252 2916 266
rect 2943 262 2978 270
rect 2980 296 3021 304
rect 2980 270 2995 296
rect 3002 270 3021 296
rect 3085 292 3116 304
rect 3131 292 3234 304
rect 3246 294 3272 320
rect 3287 315 3317 326
rect 3349 322 3411 338
rect 3349 320 3395 322
rect 3349 304 3411 320
rect 3423 304 3429 352
rect 3432 344 3512 352
rect 3432 342 3451 344
rect 3466 342 3500 344
rect 3432 327 3512 342
rect 3432 326 3518 327
rect 3432 304 3451 326
rect 3466 310 3496 326
rect 3524 320 3530 394
rect 3533 320 3552 464
rect 3567 320 3573 464
rect 3582 394 3595 464
rect 3647 460 3669 464
rect 3640 448 3657 452
rect 3661 450 3669 452
rect 3659 448 3669 450
rect 3640 438 3669 448
rect 3722 438 3738 452
rect 3776 448 3782 450
rect 3789 448 3897 464
rect 3904 448 3910 450
rect 3918 448 3933 464
rect 3999 458 4018 461
rect 3640 436 3738 438
rect 3765 436 3933 448
rect 3948 438 3964 452
rect 3999 439 4021 458
rect 4031 452 4047 453
rect 4030 450 4047 452
rect 4031 445 4047 450
rect 4021 438 4027 439
rect 4030 438 4059 445
rect 3948 437 4059 438
rect 3948 436 4065 437
rect 3624 428 3675 436
rect 3722 428 3756 436
rect 3624 416 3649 428
rect 3656 416 3675 428
rect 3729 426 3756 428
rect 3765 426 3986 436
rect 4021 433 4027 436
rect 3729 422 3986 426
rect 3624 408 3675 416
rect 3722 408 3986 422
rect 4030 428 4065 436
rect 3576 360 3595 394
rect 3640 400 3669 408
rect 3640 394 3657 400
rect 3640 392 3674 394
rect 3722 392 3738 408
rect 3739 398 3947 408
rect 3948 398 3964 408
rect 4012 404 4027 419
rect 4030 416 4031 428
rect 4038 416 4065 428
rect 4030 408 4065 416
rect 4030 407 4059 408
rect 3750 394 3964 398
rect 3765 392 3964 394
rect 3999 394 4012 404
rect 4030 394 4047 407
rect 3999 392 4047 394
rect 3641 388 3674 392
rect 3637 386 3674 388
rect 3637 385 3704 386
rect 3637 380 3668 385
rect 3674 380 3704 385
rect 3637 376 3704 380
rect 3610 373 3704 376
rect 3610 366 3659 373
rect 3610 360 3640 366
rect 3659 361 3664 366
rect 3576 344 3656 360
rect 3668 352 3704 373
rect 3765 368 3954 392
rect 3999 391 4046 392
rect 4012 386 4046 391
rect 4086 386 4102 388
rect 3780 365 3954 368
rect 3773 362 3954 365
rect 3982 385 4046 386
rect 3576 342 3595 344
rect 3610 342 3644 344
rect 3576 326 3656 342
rect 3576 320 3595 326
rect 3292 294 3395 304
rect 3246 292 3395 294
rect 3416 292 3451 304
rect 3085 290 3247 292
rect 3097 272 3116 290
rect 3131 288 3161 290
rect 2980 262 3021 270
rect 3104 266 3116 272
rect 3168 274 3247 290
rect 3279 290 3451 292
rect 3279 274 3358 290
rect 3365 288 3395 290
rect 2943 252 2972 262
rect 2986 252 3015 262
rect 3030 252 3060 266
rect 3104 252 3146 266
rect 3168 262 3358 274
rect 3423 270 3429 290
rect 3153 252 3183 262
rect 3184 252 3342 262
rect 3346 252 3376 262
rect 3380 252 3410 266
rect 3438 252 3451 290
rect 3523 304 3552 320
rect 3566 304 3595 320
rect 3610 310 3640 326
rect 3668 304 3674 352
rect 3677 346 3696 352
rect 3711 346 3741 354
rect 3677 338 3741 346
rect 3677 322 3757 338
rect 3773 331 3835 362
rect 3851 331 3913 362
rect 3982 360 4031 385
rect 4076 376 4102 386
rect 4046 360 4102 376
rect 3945 346 3975 354
rect 3982 352 4092 360
rect 3945 338 3990 346
rect 3677 320 3696 322
rect 3711 320 3757 322
rect 3677 304 3757 320
rect 3784 318 3819 331
rect 3860 328 3897 331
rect 3860 326 3902 328
rect 3789 315 3819 318
rect 3798 311 3805 315
rect 3805 310 3806 311
rect 3764 304 3774 310
rect 3523 296 3558 304
rect 3523 270 3524 296
rect 3531 270 3558 296
rect 3466 252 3496 266
rect 3523 262 3558 270
rect 3560 296 3601 304
rect 3560 270 3575 296
rect 3582 270 3601 296
rect 3665 292 3696 304
rect 3711 292 3814 304
rect 3826 294 3852 320
rect 3867 315 3897 326
rect 3929 322 3991 338
rect 3929 320 3975 322
rect 3929 304 3991 320
rect 4003 304 4009 352
rect 4012 344 4092 352
rect 4012 342 4031 344
rect 4046 342 4080 344
rect 4012 326 4092 342
rect 4012 304 4031 326
rect 4046 310 4076 326
rect 4104 320 4110 394
rect 4113 320 4132 464
rect 4147 320 4153 464
rect 4162 394 4175 464
rect 4227 460 4249 464
rect 4220 448 4237 452
rect 4241 450 4249 452
rect 4239 448 4249 450
rect 4220 438 4249 448
rect 4302 438 4318 452
rect 4356 448 4362 450
rect 4369 448 4477 464
rect 4484 448 4490 450
rect 4498 448 4513 464
rect 4579 458 4598 461
rect 4220 436 4318 438
rect 4345 436 4513 448
rect 4528 438 4544 452
rect 4579 439 4601 458
rect 4611 452 4627 453
rect 4610 450 4627 452
rect 4611 445 4627 450
rect 4601 438 4607 439
rect 4610 438 4639 445
rect 4528 437 4639 438
rect 4528 436 4645 437
rect 4204 428 4255 436
rect 4302 428 4336 436
rect 4204 416 4229 428
rect 4236 416 4255 428
rect 4309 426 4336 428
rect 4345 426 4566 436
rect 4601 433 4607 436
rect 4309 422 4566 426
rect 4204 408 4255 416
rect 4302 408 4566 422
rect 4610 428 4645 436
rect 4156 360 4175 394
rect 4220 400 4249 408
rect 4220 394 4237 400
rect 4220 392 4254 394
rect 4302 392 4318 408
rect 4319 398 4527 408
rect 4528 398 4544 408
rect 4592 404 4607 419
rect 4610 416 4611 428
rect 4618 416 4645 428
rect 4610 408 4645 416
rect 4610 407 4639 408
rect 4330 394 4544 398
rect 4345 392 4544 394
rect 4579 394 4592 404
rect 4610 394 4627 407
rect 4579 392 4627 394
rect 4221 388 4254 392
rect 4217 386 4254 388
rect 4217 385 4284 386
rect 4217 380 4248 385
rect 4254 380 4284 385
rect 4217 376 4284 380
rect 4190 373 4284 376
rect 4190 366 4239 373
rect 4190 360 4220 366
rect 4239 361 4244 366
rect 4156 344 4236 360
rect 4248 352 4284 373
rect 4345 368 4534 392
rect 4579 391 4626 392
rect 4592 386 4626 391
rect 4360 365 4534 368
rect 4353 362 4534 365
rect 4562 385 4626 386
rect 4156 342 4175 344
rect 4190 342 4224 344
rect 4156 326 4236 342
rect 4156 320 4175 326
rect 3872 294 3975 304
rect 3826 292 3975 294
rect 3996 292 4031 304
rect 3665 290 3827 292
rect 3677 272 3696 290
rect 3711 288 3741 290
rect 3560 262 3601 270
rect 3684 266 3696 272
rect 3748 274 3827 290
rect 3859 290 4031 292
rect 3859 274 3938 290
rect 3945 288 3975 290
rect 3523 252 3552 262
rect 3566 252 3595 262
rect 3610 252 3640 266
rect 3684 252 3726 266
rect 3748 262 3938 274
rect 4003 270 4009 290
rect 3733 252 3763 262
rect 3764 252 3922 262
rect 3926 252 3956 262
rect 3960 252 3990 266
rect 4018 252 4031 290
rect 4103 304 4132 320
rect 4146 304 4175 320
rect 4190 310 4220 326
rect 4248 304 4254 352
rect 4257 346 4276 352
rect 4291 346 4321 354
rect 4257 338 4321 346
rect 4257 322 4337 338
rect 4353 331 4415 362
rect 4431 331 4493 362
rect 4562 360 4611 385
rect 4626 360 4656 378
rect 4525 346 4555 354
rect 4562 352 4672 360
rect 4525 338 4570 346
rect 4257 320 4276 322
rect 4291 320 4337 322
rect 4257 304 4337 320
rect 4364 318 4399 331
rect 4440 328 4477 331
rect 4440 326 4482 328
rect 4369 315 4399 318
rect 4378 311 4385 315
rect 4385 310 4386 311
rect 4344 304 4354 310
rect 4103 296 4138 304
rect 4103 270 4104 296
rect 4111 270 4138 296
rect 4046 252 4076 266
rect 4103 262 4138 270
rect 4140 296 4181 304
rect 4140 270 4155 296
rect 4162 270 4181 296
rect 4245 292 4276 304
rect 4291 292 4394 304
rect 4406 294 4432 320
rect 4447 315 4477 326
rect 4509 322 4571 338
rect 4509 320 4555 322
rect 4509 304 4571 320
rect 4583 304 4589 352
rect 4592 344 4672 352
rect 4592 342 4611 344
rect 4626 342 4660 344
rect 4592 327 4672 342
rect 4592 326 4678 327
rect 4592 304 4611 326
rect 4626 310 4656 326
rect 4684 320 4690 394
rect 4693 320 4712 464
rect 4727 320 4733 464
rect 4742 394 4755 464
rect 4807 460 4829 464
rect 4800 448 4817 452
rect 4821 450 4829 452
rect 4819 448 4829 450
rect 4800 438 4829 448
rect 4882 438 4898 452
rect 4936 448 4942 450
rect 4949 448 5057 464
rect 5064 448 5070 450
rect 5078 448 5093 464
rect 5159 458 5178 461
rect 4800 436 4898 438
rect 4925 436 5093 448
rect 5108 438 5124 452
rect 5159 439 5181 458
rect 5191 452 5207 453
rect 5190 450 5207 452
rect 5191 445 5207 450
rect 5181 438 5187 439
rect 5190 438 5219 445
rect 5108 437 5219 438
rect 5108 436 5225 437
rect 4784 428 4835 436
rect 4882 428 4916 436
rect 4784 416 4809 428
rect 4816 416 4835 428
rect 4889 426 4916 428
rect 4925 426 5146 436
rect 5181 433 5187 436
rect 4889 422 5146 426
rect 4784 408 4835 416
rect 4882 408 5146 422
rect 5190 428 5225 436
rect 4736 360 4755 394
rect 4800 400 4829 408
rect 4800 394 4817 400
rect 4800 392 4834 394
rect 4882 392 4898 408
rect 4899 398 5107 408
rect 5108 398 5124 408
rect 5172 404 5187 419
rect 5190 416 5191 428
rect 5198 416 5225 428
rect 5190 408 5225 416
rect 5190 407 5219 408
rect 4910 394 5124 398
rect 4925 392 5124 394
rect 5159 394 5172 404
rect 5190 394 5207 407
rect 5159 392 5207 394
rect 4801 388 4834 392
rect 4797 386 4834 388
rect 4797 385 4864 386
rect 4797 380 4828 385
rect 4834 380 4864 385
rect 4797 376 4864 380
rect 4770 373 4864 376
rect 4770 366 4819 373
rect 4770 360 4800 366
rect 4819 361 4824 366
rect 4736 344 4816 360
rect 4828 352 4864 373
rect 4925 368 5114 392
rect 5159 391 5206 392
rect 5172 386 5206 391
rect 5246 386 5262 388
rect 4940 365 5114 368
rect 4933 362 5114 365
rect 5142 385 5206 386
rect 4736 342 4755 344
rect 4770 342 4804 344
rect 4736 326 4816 342
rect 4736 320 4755 326
rect 4452 294 4555 304
rect 4406 292 4555 294
rect 4576 292 4611 304
rect 4245 290 4407 292
rect 4257 272 4276 290
rect 4291 288 4321 290
rect 4140 262 4181 270
rect 4264 266 4276 272
rect 4328 274 4407 290
rect 4439 290 4611 292
rect 4439 274 4518 290
rect 4525 288 4555 290
rect 4103 252 4132 262
rect 4146 252 4175 262
rect 4190 252 4220 266
rect 4264 252 4306 266
rect 4328 262 4518 274
rect 4583 270 4589 290
rect 4313 252 4343 262
rect 4344 252 4502 262
rect 4506 252 4536 262
rect 4540 252 4570 266
rect 4598 252 4611 290
rect 4683 304 4712 320
rect 4726 304 4755 320
rect 4770 310 4800 326
rect 4828 304 4834 352
rect 4837 346 4856 352
rect 4871 346 4901 354
rect 4837 338 4901 346
rect 4837 322 4917 338
rect 4933 331 4995 362
rect 5011 331 5073 362
rect 5142 360 5191 385
rect 5236 376 5262 386
rect 5206 360 5262 376
rect 5105 346 5135 354
rect 5142 352 5252 360
rect 5105 338 5150 346
rect 4837 320 4856 322
rect 4871 320 4917 322
rect 4837 304 4917 320
rect 4944 318 4979 331
rect 5020 328 5057 331
rect 5020 326 5062 328
rect 4949 315 4979 318
rect 4958 311 4965 315
rect 4965 310 4966 311
rect 4924 304 4934 310
rect 4683 296 4718 304
rect 4683 270 4684 296
rect 4691 270 4718 296
rect 4626 252 4656 266
rect 4683 262 4718 270
rect 4720 296 4761 304
rect 4720 270 4735 296
rect 4742 270 4761 296
rect 4825 292 4856 304
rect 4871 292 4974 304
rect 4986 294 5012 320
rect 5027 315 5057 326
rect 5089 322 5151 338
rect 5089 320 5135 322
rect 5089 304 5151 320
rect 5163 304 5169 352
rect 5172 344 5252 352
rect 5172 342 5191 344
rect 5206 342 5240 344
rect 5172 326 5252 342
rect 5172 304 5191 326
rect 5206 310 5236 326
rect 5264 320 5270 394
rect 5273 320 5292 464
rect 5307 320 5313 464
rect 5322 394 5335 464
rect 5387 460 5409 464
rect 5380 448 5397 452
rect 5401 450 5409 452
rect 5399 448 5409 450
rect 5380 438 5409 448
rect 5462 438 5478 452
rect 5516 448 5522 450
rect 5529 448 5637 464
rect 5644 448 5650 450
rect 5658 448 5673 464
rect 5739 458 5758 461
rect 5380 436 5478 438
rect 5505 436 5673 448
rect 5688 438 5704 452
rect 5739 439 5761 458
rect 5771 452 5787 453
rect 5770 450 5787 452
rect 5771 445 5787 450
rect 5761 438 5767 439
rect 5770 438 5799 445
rect 5688 437 5799 438
rect 5688 436 5805 437
rect 5364 428 5415 436
rect 5462 428 5496 436
rect 5364 416 5389 428
rect 5396 416 5415 428
rect 5469 426 5496 428
rect 5505 426 5726 436
rect 5761 433 5767 436
rect 5469 422 5726 426
rect 5364 408 5415 416
rect 5462 408 5726 422
rect 5770 428 5805 436
rect 5316 360 5335 394
rect 5380 400 5409 408
rect 5380 394 5397 400
rect 5380 392 5414 394
rect 5462 392 5478 408
rect 5479 398 5687 408
rect 5688 398 5704 408
rect 5752 404 5767 419
rect 5770 416 5771 428
rect 5778 416 5805 428
rect 5770 408 5805 416
rect 5770 407 5799 408
rect 5490 394 5704 398
rect 5505 392 5704 394
rect 5739 394 5752 404
rect 5770 394 5787 407
rect 5739 392 5787 394
rect 5381 388 5414 392
rect 5377 386 5414 388
rect 5377 385 5444 386
rect 5377 380 5408 385
rect 5414 380 5444 385
rect 5377 376 5444 380
rect 5350 373 5444 376
rect 5350 366 5399 373
rect 5350 360 5380 366
rect 5399 361 5404 366
rect 5316 344 5396 360
rect 5408 352 5444 373
rect 5505 368 5694 392
rect 5739 391 5786 392
rect 5752 386 5786 391
rect 5520 365 5694 368
rect 5513 362 5694 365
rect 5722 385 5786 386
rect 5316 342 5335 344
rect 5350 342 5384 344
rect 5316 326 5396 342
rect 5316 320 5335 326
rect 5032 294 5135 304
rect 4986 292 5135 294
rect 5156 292 5191 304
rect 4825 290 4987 292
rect 4837 272 4856 290
rect 4871 288 4901 290
rect 4720 262 4761 270
rect 4844 266 4856 272
rect 4908 274 4987 290
rect 5019 290 5191 292
rect 5019 274 5098 290
rect 5105 288 5135 290
rect 4683 252 4712 262
rect 4726 252 4755 262
rect 4770 252 4800 266
rect 4844 252 4886 266
rect 4908 262 5098 274
rect 5163 270 5169 290
rect 4893 252 4923 262
rect 4924 252 5082 262
rect 5086 252 5116 262
rect 5120 252 5150 266
rect 5178 252 5191 290
rect 5263 304 5292 320
rect 5306 304 5335 320
rect 5350 310 5380 326
rect 5408 304 5414 352
rect 5417 346 5436 352
rect 5451 346 5481 354
rect 5417 338 5481 346
rect 5417 322 5497 338
rect 5513 331 5575 362
rect 5591 331 5653 362
rect 5722 360 5771 385
rect 5786 360 5816 378
rect 5685 346 5715 354
rect 5722 352 5832 360
rect 5685 338 5730 346
rect 5417 320 5436 322
rect 5451 320 5497 322
rect 5417 304 5497 320
rect 5524 318 5559 331
rect 5600 328 5637 331
rect 5600 326 5642 328
rect 5529 315 5559 318
rect 5538 311 5545 315
rect 5545 310 5546 311
rect 5504 304 5514 310
rect 5263 296 5298 304
rect 5263 270 5264 296
rect 5271 270 5298 296
rect 5206 252 5236 266
rect 5263 262 5298 270
rect 5300 296 5341 304
rect 5300 270 5315 296
rect 5322 270 5341 296
rect 5405 292 5436 304
rect 5451 292 5554 304
rect 5566 294 5592 320
rect 5607 315 5637 326
rect 5669 322 5731 338
rect 5669 320 5715 322
rect 5669 304 5731 320
rect 5743 304 5749 352
rect 5752 344 5832 352
rect 5752 342 5771 344
rect 5786 342 5820 344
rect 5752 327 5832 342
rect 5752 326 5838 327
rect 5752 304 5771 326
rect 5786 310 5816 326
rect 5844 320 5850 394
rect 5853 320 5872 464
rect 5887 320 5893 464
rect 5902 394 5915 464
rect 5967 460 5989 464
rect 5960 448 5977 452
rect 5981 450 5989 452
rect 5979 448 5989 450
rect 5960 438 5989 448
rect 6042 438 6058 452
rect 6096 448 6102 450
rect 6109 448 6217 464
rect 6224 448 6230 450
rect 6238 448 6253 464
rect 6319 458 6338 461
rect 5960 436 6058 438
rect 6085 436 6253 448
rect 6268 438 6284 452
rect 6319 439 6341 458
rect 6351 452 6367 453
rect 6350 450 6367 452
rect 6351 445 6367 450
rect 6341 438 6347 439
rect 6350 438 6379 445
rect 6268 437 6379 438
rect 6268 436 6385 437
rect 5944 428 5995 436
rect 6042 428 6076 436
rect 5944 416 5969 428
rect 5976 416 5995 428
rect 6049 426 6076 428
rect 6085 426 6306 436
rect 6341 433 6347 436
rect 6049 422 6306 426
rect 5944 408 5995 416
rect 6042 408 6306 422
rect 6350 428 6385 436
rect 5896 360 5915 394
rect 5960 400 5989 408
rect 5960 394 5977 400
rect 5960 392 5994 394
rect 6042 392 6058 408
rect 6059 398 6267 408
rect 6268 398 6284 408
rect 6332 404 6347 419
rect 6350 416 6351 428
rect 6358 416 6385 428
rect 6350 408 6385 416
rect 6350 407 6379 408
rect 6070 394 6284 398
rect 6085 392 6284 394
rect 6319 394 6332 404
rect 6350 394 6367 407
rect 6319 392 6367 394
rect 5961 388 5994 392
rect 5957 386 5994 388
rect 5957 385 6024 386
rect 5957 380 5988 385
rect 5994 380 6024 385
rect 5957 376 6024 380
rect 5930 373 6024 376
rect 5930 366 5979 373
rect 5930 360 5960 366
rect 5979 361 5984 366
rect 5896 344 5976 360
rect 5988 352 6024 373
rect 6085 368 6274 392
rect 6319 391 6366 392
rect 6332 386 6366 391
rect 6100 365 6274 368
rect 6093 362 6274 365
rect 6302 385 6366 386
rect 5896 342 5915 344
rect 5930 342 5964 344
rect 5896 326 5976 342
rect 5896 320 5915 326
rect 5612 294 5715 304
rect 5566 292 5715 294
rect 5736 292 5771 304
rect 5405 290 5567 292
rect 5417 272 5436 290
rect 5451 288 5481 290
rect 5300 262 5341 270
rect 5424 266 5436 272
rect 5488 274 5567 290
rect 5599 290 5771 292
rect 5599 274 5678 290
rect 5685 288 5715 290
rect 5263 252 5292 262
rect 5306 252 5335 262
rect 5350 252 5380 266
rect 5424 252 5466 266
rect 5488 262 5678 274
rect 5743 270 5749 290
rect 5473 252 5503 262
rect 5504 252 5662 262
rect 5666 252 5696 262
rect 5700 252 5730 266
rect 5758 252 5771 290
rect 5843 304 5872 320
rect 5886 304 5915 320
rect 5930 310 5960 326
rect 5988 304 5994 352
rect 5997 346 6016 352
rect 6031 346 6061 354
rect 5997 338 6061 346
rect 5997 322 6077 338
rect 6093 331 6155 362
rect 6171 331 6233 362
rect 6302 360 6351 385
rect 6366 360 6396 376
rect 6265 346 6295 354
rect 6302 352 6412 360
rect 6265 338 6310 346
rect 5997 320 6016 322
rect 6031 320 6077 322
rect 5997 304 6077 320
rect 6104 318 6139 331
rect 6180 328 6217 331
rect 6180 326 6222 328
rect 6109 315 6139 318
rect 6118 311 6125 315
rect 6125 310 6126 311
rect 6084 304 6094 310
rect 5843 296 5878 304
rect 5843 270 5844 296
rect 5851 270 5878 296
rect 5786 252 5816 266
rect 5843 262 5878 270
rect 5880 296 5921 304
rect 5880 270 5895 296
rect 5902 270 5921 296
rect 5985 292 6016 304
rect 6031 292 6134 304
rect 6146 294 6172 320
rect 6187 315 6217 326
rect 6249 322 6311 338
rect 6249 320 6295 322
rect 6249 304 6311 320
rect 6323 304 6329 352
rect 6332 344 6412 352
rect 6332 342 6351 344
rect 6366 342 6400 344
rect 6332 326 6412 342
rect 6332 304 6351 326
rect 6366 310 6396 326
rect 6424 320 6430 394
rect 6439 320 6452 464
rect 6192 294 6295 304
rect 6146 292 6295 294
rect 6316 292 6351 304
rect 5985 290 6147 292
rect 5997 272 6016 290
rect 6031 288 6061 290
rect 5880 262 5921 270
rect 6004 266 6016 272
rect 6068 274 6147 290
rect 6179 290 6351 292
rect 6179 274 6258 290
rect 6265 288 6295 290
rect 5843 252 5872 262
rect 5886 252 5915 262
rect 5930 252 5960 266
rect 6004 252 6046 266
rect 6068 262 6258 274
rect 6323 270 6329 290
rect 6053 252 6083 262
rect 6084 252 6242 262
rect 6246 252 6276 262
rect 6280 252 6310 266
rect 6338 252 6351 290
rect 6423 304 6452 320
rect 6423 296 6458 304
rect 6423 270 6424 296
rect 6431 270 6458 296
rect 6366 252 6396 266
rect 6423 262 6458 270
rect 6423 252 6452 262
rect -541 238 6452 252
rect -478 208 -465 238
rect -450 224 -420 238
rect -376 224 -334 238
rect -327 224 -107 238
rect -100 224 -70 238
rect -410 210 -395 222
rect -376 210 -363 224
rect -295 220 -142 224
rect -413 208 -391 210
rect -313 208 -121 220
rect -42 208 -29 238
rect -14 224 16 238
rect 53 208 72 238
rect 87 208 93 238
rect 102 208 115 238
rect 130 224 160 238
rect 204 224 246 238
rect 253 224 473 238
rect 480 224 510 238
rect 170 210 185 222
rect 204 210 217 224
rect 285 220 438 224
rect 167 208 189 210
rect 267 208 459 220
rect 538 208 551 238
rect 566 224 596 238
rect 633 208 652 238
rect 667 208 673 238
rect 682 208 695 238
rect 710 224 740 238
rect 784 224 826 238
rect 833 224 1053 238
rect 1060 224 1090 238
rect 750 210 765 222
rect 784 210 797 224
rect 865 220 1018 224
rect 747 208 769 210
rect 847 208 1039 220
rect 1118 208 1131 238
rect 1146 224 1176 238
rect 1213 208 1232 238
rect 1247 208 1253 238
rect 1262 208 1275 238
rect 1290 224 1320 238
rect 1364 224 1406 238
rect 1413 224 1633 238
rect 1640 224 1670 238
rect 1330 210 1345 222
rect 1364 210 1377 224
rect 1445 220 1598 224
rect 1327 208 1349 210
rect 1427 208 1619 220
rect 1698 208 1711 238
rect 1726 224 1756 238
rect 1793 208 1812 238
rect 1827 208 1833 238
rect 1842 208 1855 238
rect 1870 224 1900 238
rect 1944 224 1986 238
rect 1993 224 2213 238
rect 2220 224 2250 238
rect 1910 210 1925 222
rect 1944 210 1957 224
rect 2025 220 2178 224
rect 1907 208 1929 210
rect 2007 208 2199 220
rect 2278 208 2291 238
rect 2306 224 2336 238
rect 2373 208 2392 238
rect 2407 208 2413 238
rect 2422 208 2435 238
rect 2450 224 2480 238
rect 2524 224 2566 238
rect 2573 224 2793 238
rect 2800 224 2830 238
rect 2490 210 2505 222
rect 2524 210 2537 224
rect 2605 220 2758 224
rect 2487 208 2509 210
rect 2587 208 2779 220
rect 2858 208 2871 238
rect 2886 224 2916 238
rect 2953 208 2972 238
rect 2987 208 2993 238
rect 3002 208 3015 238
rect 3030 224 3060 238
rect 3104 224 3146 238
rect 3153 224 3373 238
rect 3380 224 3410 238
rect 3070 210 3085 222
rect 3104 210 3117 224
rect 3185 220 3338 224
rect 3067 208 3089 210
rect 3167 208 3359 220
rect 3438 208 3451 238
rect 3466 224 3496 238
rect 3533 208 3552 238
rect 3567 208 3573 238
rect 3582 208 3595 238
rect 3610 224 3640 238
rect 3684 224 3726 238
rect 3733 224 3953 238
rect 3960 224 3990 238
rect 3650 210 3665 222
rect 3684 210 3697 224
rect 3765 220 3918 224
rect 3647 208 3669 210
rect 3747 208 3939 220
rect 4018 208 4031 238
rect 4046 224 4076 238
rect 4113 208 4132 238
rect 4147 208 4153 238
rect 4162 208 4175 238
rect 4190 224 4220 238
rect 4264 224 4306 238
rect 4313 224 4533 238
rect 4540 224 4570 238
rect 4230 210 4245 222
rect 4264 210 4277 224
rect 4345 220 4498 224
rect 4227 208 4249 210
rect 4327 208 4519 220
rect 4598 208 4611 238
rect 4626 224 4656 238
rect 4693 208 4712 238
rect 4727 208 4733 238
rect 4742 208 4755 238
rect 4770 224 4800 238
rect 4844 224 4886 238
rect 4893 224 5113 238
rect 5120 224 5150 238
rect 4810 210 4825 222
rect 4844 210 4857 224
rect 4925 220 5078 224
rect 4807 208 4829 210
rect 4907 208 5099 220
rect 5178 208 5191 238
rect 5206 224 5236 238
rect 5273 208 5292 238
rect 5307 208 5313 238
rect 5322 208 5335 238
rect 5350 224 5380 238
rect 5424 224 5466 238
rect 5473 224 5693 238
rect 5700 224 5730 238
rect 5390 210 5405 222
rect 5424 210 5437 224
rect 5505 220 5658 224
rect 5387 208 5409 210
rect 5487 208 5679 220
rect 5758 208 5771 238
rect 5786 224 5816 238
rect 5853 208 5872 238
rect 5887 208 5893 238
rect 5902 208 5915 238
rect 5930 224 5960 238
rect 6004 224 6046 238
rect 6053 224 6273 238
rect 6280 224 6310 238
rect 5970 210 5985 222
rect 6004 210 6017 224
rect 6085 220 6238 224
rect 5967 208 5989 210
rect 6067 208 6259 220
rect 6338 208 6351 238
rect 6366 224 6396 238
rect 6439 208 6452 238
rect -541 194 6452 208
rect -478 124 -465 194
rect -413 190 -391 194
rect -420 178 -403 182
rect -399 180 -391 182
rect -401 178 -391 180
rect -420 168 -391 178
rect -338 168 -322 182
rect -284 178 -278 180
rect -271 178 -163 194
rect -156 178 -150 180
rect -142 178 -127 194
rect -61 188 -42 191
rect -420 166 -322 168
rect -295 166 -127 178
rect -112 168 -96 182
rect -61 169 -39 188
rect -29 182 -13 183
rect -30 176 -13 182
rect -29 175 -13 176
rect -39 168 -33 169
rect -30 168 -1 175
rect -112 167 -1 168
rect -112 166 5 167
rect -436 158 -385 166
rect -338 158 -304 166
rect -436 146 -411 158
rect -404 146 -385 158
rect -331 156 -304 158
rect -295 156 -74 166
rect -39 163 -33 166
rect -331 152 -74 156
rect -436 138 -385 146
rect -338 138 -74 152
rect -30 158 5 166
rect -484 90 -465 124
rect -420 130 -391 138
rect -420 124 -403 130
rect -420 122 -386 124
rect -338 122 -322 138
rect -321 128 -113 138
rect -112 128 -96 138
rect -48 134 -33 149
rect -30 146 -29 158
rect -22 146 5 158
rect -30 138 5 146
rect -30 137 -1 138
rect -310 124 -96 128
rect -295 122 -96 124
rect -61 124 -48 134
rect -30 124 -13 137
rect -61 122 -13 124
rect -419 118 -386 122
rect -423 116 -386 118
rect -423 115 -356 116
rect -423 110 -392 115
rect -386 110 -356 115
rect -423 106 -356 110
rect -450 103 -356 106
rect -450 96 -401 103
rect -450 90 -420 96
rect -401 91 -396 96
rect -484 74 -404 90
rect -392 82 -356 103
rect -295 98 -106 122
rect -61 121 -14 122
rect -48 116 -14 121
rect -280 95 -106 98
rect -287 92 -106 95
rect -78 115 -14 116
rect -484 72 -465 74
rect -450 72 -416 74
rect -484 56 -404 72
rect -484 50 -465 56
rect -494 34 -465 50
rect -450 40 -420 56
rect -392 34 -386 82
rect -383 76 -364 82
rect -349 76 -319 84
rect -383 68 -319 76
rect -383 52 -303 68
rect -287 61 -225 92
rect -209 61 -147 92
rect -78 90 -29 115
rect -14 90 16 108
rect -115 76 -85 84
rect -78 82 32 90
rect -115 68 -70 76
rect -383 50 -364 52
rect -349 50 -303 52
rect -383 34 -303 50
rect -276 48 -241 61
rect -200 58 -163 61
rect -200 56 -158 58
rect -271 45 -241 48
rect -262 41 -255 45
rect -255 40 -254 41
rect -296 34 -286 40
rect -500 26 -459 34
rect -500 0 -485 26
rect -478 0 -459 26
rect -395 22 -364 34
rect -349 22 -246 34
rect -234 24 -208 50
rect -193 45 -163 56
rect -131 52 -69 68
rect -131 50 -85 52
rect -131 34 -69 50
rect -57 34 -51 82
rect -48 74 32 82
rect -48 72 -29 74
rect -14 72 20 74
rect -48 57 32 72
rect -48 56 38 57
rect -48 34 -29 56
rect -14 40 16 56
rect 44 50 50 124
rect 53 50 72 194
rect 87 50 93 194
rect 102 124 115 194
rect 167 190 189 194
rect 160 178 177 182
rect 181 180 189 182
rect 179 178 189 180
rect 160 168 189 178
rect 242 168 258 182
rect 296 178 302 180
rect 309 178 417 194
rect 424 178 430 180
rect 438 178 453 194
rect 519 188 538 191
rect 160 166 258 168
rect 285 166 453 178
rect 468 168 484 182
rect 519 169 541 188
rect 551 182 567 183
rect 550 176 567 182
rect 551 175 567 176
rect 541 168 547 169
rect 550 168 579 175
rect 468 167 579 168
rect 468 166 585 167
rect 144 158 195 166
rect 242 158 276 166
rect 144 146 169 158
rect 176 146 195 158
rect 249 156 276 158
rect 285 156 506 166
rect 541 163 547 166
rect 249 152 506 156
rect 144 138 195 146
rect 242 138 506 152
rect 550 158 585 166
rect 96 90 115 124
rect 160 130 189 138
rect 160 124 177 130
rect 160 122 194 124
rect 242 122 258 138
rect 259 128 467 138
rect 468 128 484 138
rect 532 134 547 149
rect 550 146 551 158
rect 558 146 585 158
rect 550 138 585 146
rect 550 137 579 138
rect 270 124 484 128
rect 285 122 484 124
rect 519 124 532 134
rect 550 124 567 137
rect 519 122 567 124
rect 161 118 194 122
rect 157 116 194 118
rect 157 115 224 116
rect 157 110 188 115
rect 194 110 224 115
rect 157 106 224 110
rect 130 103 224 106
rect 130 96 179 103
rect 130 90 160 96
rect 179 91 184 96
rect 96 74 176 90
rect 188 82 224 103
rect 285 98 474 122
rect 519 121 566 122
rect 532 116 566 121
rect 606 116 622 118
rect 300 95 474 98
rect 293 92 474 95
rect 502 115 566 116
rect 96 72 115 74
rect 130 72 164 74
rect 96 56 176 72
rect 96 50 115 56
rect -188 24 -85 34
rect -234 22 -85 24
rect -64 22 -29 34
rect -395 20 -233 22
rect -383 0 -364 20
rect -349 18 -319 20
rect -500 -8 -459 0
rect -377 -4 -364 0
rect -312 4 -233 20
rect -201 20 -29 22
rect -201 4 -122 20
rect -115 18 -85 20
rect -494 -18 -465 -8
rect -450 -18 -420 -4
rect -377 -18 -334 -4
rect -312 -8 -122 4
rect -57 0 -51 20
rect -327 -18 -297 -8
rect -296 -18 -138 -8
rect -134 -18 -104 -8
rect -100 -18 -70 -4
rect -42 -18 -29 20
rect 43 34 72 50
rect 86 34 115 50
rect 130 40 160 56
rect 188 34 194 82
rect 197 76 216 82
rect 231 76 261 84
rect 197 68 261 76
rect 197 52 277 68
rect 293 61 355 92
rect 371 61 433 92
rect 502 90 551 115
rect 596 106 622 116
rect 566 90 622 106
rect 465 76 495 84
rect 502 82 612 90
rect 465 68 510 76
rect 197 50 216 52
rect 231 50 277 52
rect 197 34 277 50
rect 304 48 339 61
rect 380 58 417 61
rect 380 56 422 58
rect 309 45 339 48
rect 318 41 325 45
rect 325 40 326 41
rect 284 34 294 40
rect 43 26 78 34
rect 43 0 44 26
rect 51 0 78 26
rect -14 -18 16 -4
rect 43 -8 78 0
rect 80 26 121 34
rect 80 0 95 26
rect 102 0 121 26
rect 185 22 216 34
rect 231 22 334 34
rect 346 24 372 50
rect 387 45 417 56
rect 449 52 511 68
rect 449 50 495 52
rect 449 34 511 50
rect 523 34 529 82
rect 532 74 612 82
rect 532 72 551 74
rect 566 72 600 74
rect 532 56 612 72
rect 532 34 551 56
rect 566 40 596 56
rect 624 50 630 124
rect 633 50 652 194
rect 667 50 673 194
rect 682 124 695 194
rect 747 190 769 194
rect 740 178 757 182
rect 761 180 769 182
rect 759 178 769 180
rect 740 168 769 178
rect 822 168 838 182
rect 876 178 882 180
rect 889 178 997 194
rect 1004 178 1010 180
rect 1018 178 1033 194
rect 1099 188 1118 191
rect 740 166 838 168
rect 865 166 1033 178
rect 1048 168 1064 182
rect 1099 169 1121 188
rect 1131 182 1147 183
rect 1130 180 1147 182
rect 1131 175 1147 180
rect 1121 168 1127 169
rect 1130 168 1159 175
rect 1048 167 1159 168
rect 1048 166 1165 167
rect 724 158 775 166
rect 822 158 856 166
rect 724 146 749 158
rect 756 146 775 158
rect 829 156 856 158
rect 865 156 1086 166
rect 1121 163 1127 166
rect 829 152 1086 156
rect 724 138 775 146
rect 822 138 1086 152
rect 1130 158 1165 166
rect 676 90 695 124
rect 740 130 769 138
rect 740 124 757 130
rect 740 122 774 124
rect 822 122 838 138
rect 839 128 1047 138
rect 1048 128 1064 138
rect 1112 134 1127 149
rect 1130 146 1131 158
rect 1138 146 1165 158
rect 1130 138 1165 146
rect 1130 137 1159 138
rect 850 124 1064 128
rect 865 122 1064 124
rect 1099 124 1112 134
rect 1130 124 1147 137
rect 1099 122 1147 124
rect 741 118 774 122
rect 737 116 774 118
rect 737 115 804 116
rect 737 110 768 115
rect 774 110 804 115
rect 737 106 804 110
rect 710 103 804 106
rect 710 96 759 103
rect 710 90 740 96
rect 759 91 764 96
rect 676 74 756 90
rect 768 82 804 103
rect 865 98 1054 122
rect 1099 121 1146 122
rect 1112 116 1146 121
rect 880 95 1054 98
rect 873 92 1054 95
rect 1082 115 1146 116
rect 676 72 695 74
rect 710 72 744 74
rect 676 56 756 72
rect 676 50 695 56
rect 392 24 495 34
rect 346 22 495 24
rect 516 22 551 34
rect 185 20 347 22
rect 197 0 216 20
rect 231 18 261 20
rect 80 -8 121 0
rect 203 -4 216 0
rect 268 4 347 20
rect 379 20 551 22
rect 379 4 458 20
rect 465 18 495 20
rect 43 -18 72 -8
rect 86 -18 115 -8
rect 130 -18 160 -4
rect 203 -18 246 -4
rect 268 -8 458 4
rect 523 0 529 20
rect 253 -18 283 -8
rect 284 -18 442 -8
rect 446 -18 476 -8
rect 480 -18 510 -4
rect 538 -18 551 20
rect 623 34 652 50
rect 666 34 695 50
rect 710 40 740 56
rect 768 34 774 82
rect 777 76 796 82
rect 811 76 841 84
rect 777 68 841 76
rect 777 52 857 68
rect 873 61 935 92
rect 951 61 1013 92
rect 1082 90 1131 115
rect 1146 90 1176 108
rect 1045 76 1075 84
rect 1082 82 1192 90
rect 1045 68 1090 76
rect 777 50 796 52
rect 811 50 857 52
rect 777 34 857 50
rect 884 48 919 61
rect 960 58 997 61
rect 960 56 1002 58
rect 889 45 919 48
rect 898 41 905 45
rect 905 40 906 41
rect 864 34 874 40
rect 623 26 658 34
rect 623 0 624 26
rect 631 0 658 26
rect 566 -18 596 -4
rect 623 -8 658 0
rect 660 26 701 34
rect 660 0 675 26
rect 682 0 701 26
rect 765 22 796 34
rect 811 22 914 34
rect 926 24 952 50
rect 967 45 997 56
rect 1029 52 1091 68
rect 1029 50 1075 52
rect 1029 34 1091 50
rect 1103 34 1109 82
rect 1112 74 1192 82
rect 1112 72 1131 74
rect 1146 72 1180 74
rect 1112 57 1192 72
rect 1112 56 1198 57
rect 1112 34 1131 56
rect 1146 40 1176 56
rect 1204 50 1210 124
rect 1213 50 1232 194
rect 1247 50 1253 194
rect 1262 124 1275 194
rect 1327 190 1349 194
rect 1320 178 1337 182
rect 1341 180 1349 182
rect 1339 178 1349 180
rect 1320 168 1349 178
rect 1402 168 1418 182
rect 1456 178 1462 180
rect 1469 178 1577 194
rect 1584 178 1590 180
rect 1598 178 1613 194
rect 1679 188 1698 191
rect 1320 166 1418 168
rect 1445 166 1613 178
rect 1628 168 1644 182
rect 1679 169 1701 188
rect 1711 182 1727 183
rect 1710 180 1727 182
rect 1711 175 1727 180
rect 1701 168 1707 169
rect 1710 168 1739 175
rect 1628 167 1739 168
rect 1628 166 1745 167
rect 1304 158 1355 166
rect 1402 158 1436 166
rect 1304 146 1329 158
rect 1336 146 1355 158
rect 1409 156 1436 158
rect 1445 156 1666 166
rect 1701 163 1707 166
rect 1409 152 1666 156
rect 1304 138 1355 146
rect 1402 138 1666 152
rect 1710 158 1745 166
rect 1256 90 1275 124
rect 1320 130 1349 138
rect 1320 124 1337 130
rect 1320 122 1354 124
rect 1402 122 1418 138
rect 1419 128 1627 138
rect 1628 128 1644 138
rect 1692 134 1707 149
rect 1710 146 1711 158
rect 1718 146 1745 158
rect 1710 138 1745 146
rect 1710 137 1739 138
rect 1430 124 1644 128
rect 1445 122 1644 124
rect 1679 124 1692 134
rect 1710 124 1727 137
rect 1679 122 1727 124
rect 1321 118 1354 122
rect 1317 116 1354 118
rect 1317 115 1384 116
rect 1317 110 1348 115
rect 1354 110 1384 115
rect 1317 106 1384 110
rect 1290 103 1384 106
rect 1290 96 1339 103
rect 1290 90 1320 96
rect 1339 91 1344 96
rect 1256 74 1336 90
rect 1348 82 1384 103
rect 1445 98 1634 122
rect 1679 121 1726 122
rect 1692 116 1726 121
rect 1766 116 1782 118
rect 1460 95 1634 98
rect 1453 92 1634 95
rect 1662 115 1726 116
rect 1256 72 1275 74
rect 1290 72 1324 74
rect 1256 56 1336 72
rect 1256 50 1275 56
rect 972 24 1075 34
rect 926 22 1075 24
rect 1096 22 1131 34
rect 765 20 927 22
rect 777 0 796 20
rect 811 18 841 20
rect 660 -8 701 0
rect 783 -4 796 0
rect 848 4 927 20
rect 959 20 1131 22
rect 959 4 1038 20
rect 1045 18 1075 20
rect 623 -18 652 -8
rect 666 -18 695 -8
rect 710 -18 740 -4
rect 783 -18 826 -4
rect 848 -8 1038 4
rect 1103 0 1109 20
rect 833 -18 863 -8
rect 864 -18 1022 -8
rect 1026 -18 1056 -8
rect 1060 -18 1090 -4
rect 1118 -18 1131 20
rect 1203 34 1232 50
rect 1246 34 1275 50
rect 1290 40 1320 56
rect 1348 34 1354 82
rect 1357 76 1376 82
rect 1391 76 1421 84
rect 1357 68 1421 76
rect 1357 52 1437 68
rect 1453 61 1515 92
rect 1531 61 1593 92
rect 1662 90 1711 115
rect 1756 106 1782 116
rect 1726 90 1782 106
rect 1625 76 1655 84
rect 1662 82 1772 90
rect 1625 68 1670 76
rect 1357 50 1376 52
rect 1391 50 1437 52
rect 1357 34 1437 50
rect 1464 48 1499 61
rect 1540 58 1577 61
rect 1540 56 1582 58
rect 1469 45 1499 48
rect 1478 41 1485 45
rect 1485 40 1486 41
rect 1444 34 1454 40
rect 1203 26 1238 34
rect 1203 0 1204 26
rect 1211 0 1238 26
rect 1146 -18 1176 -4
rect 1203 -8 1238 0
rect 1240 26 1281 34
rect 1240 0 1255 26
rect 1262 0 1281 26
rect 1345 22 1376 34
rect 1391 22 1494 34
rect 1506 24 1532 50
rect 1547 45 1577 56
rect 1609 52 1671 68
rect 1609 50 1655 52
rect 1609 34 1671 50
rect 1683 34 1689 82
rect 1692 74 1772 82
rect 1692 72 1711 74
rect 1726 72 1760 74
rect 1692 56 1772 72
rect 1692 34 1711 56
rect 1726 40 1756 56
rect 1784 50 1790 124
rect 1793 50 1812 194
rect 1827 50 1833 194
rect 1842 124 1855 194
rect 1907 190 1929 194
rect 1900 178 1917 182
rect 1921 180 1929 182
rect 1919 178 1929 180
rect 1900 168 1929 178
rect 1982 168 1998 182
rect 2036 178 2042 180
rect 2049 178 2157 194
rect 2164 178 2170 180
rect 2178 178 2193 194
rect 2259 188 2278 191
rect 1900 166 1998 168
rect 2025 166 2193 178
rect 2208 168 2224 182
rect 2259 169 2281 188
rect 2291 182 2307 183
rect 2290 176 2307 182
rect 2291 175 2307 176
rect 2281 168 2287 169
rect 2290 168 2319 175
rect 2208 167 2319 168
rect 2208 166 2325 167
rect 1884 158 1935 166
rect 1982 158 2016 166
rect 1884 146 1909 158
rect 1916 146 1935 158
rect 1989 156 2016 158
rect 2025 156 2246 166
rect 2281 163 2287 166
rect 1989 152 2246 156
rect 1884 138 1935 146
rect 1982 138 2246 152
rect 2290 158 2325 166
rect 1836 90 1855 124
rect 1900 130 1929 138
rect 1900 124 1917 130
rect 1900 122 1934 124
rect 1982 122 1998 138
rect 1999 128 2207 138
rect 2208 128 2224 138
rect 2272 134 2287 149
rect 2290 146 2291 158
rect 2298 146 2325 158
rect 2290 138 2325 146
rect 2290 137 2319 138
rect 2010 124 2224 128
rect 2025 122 2224 124
rect 2259 124 2272 134
rect 2290 124 2307 137
rect 2259 122 2307 124
rect 1901 118 1934 122
rect 1897 116 1934 118
rect 1897 115 1964 116
rect 1897 110 1928 115
rect 1934 110 1964 115
rect 1897 106 1964 110
rect 1870 103 1964 106
rect 1870 96 1919 103
rect 1870 90 1900 96
rect 1919 91 1924 96
rect 1836 74 1916 90
rect 1928 82 1964 103
rect 2025 98 2214 122
rect 2259 121 2306 122
rect 2272 116 2306 121
rect 2040 95 2214 98
rect 2033 92 2214 95
rect 2242 115 2306 116
rect 1836 72 1855 74
rect 1870 72 1904 74
rect 1836 56 1916 72
rect 1836 50 1855 56
rect 1552 24 1655 34
rect 1506 22 1655 24
rect 1676 22 1711 34
rect 1345 20 1507 22
rect 1357 0 1376 20
rect 1391 18 1421 20
rect 1240 -8 1281 0
rect 1363 -4 1376 0
rect 1428 4 1507 20
rect 1539 20 1711 22
rect 1539 4 1618 20
rect 1625 18 1655 20
rect 1203 -18 1232 -8
rect 1246 -18 1275 -8
rect 1290 -18 1320 -4
rect 1363 -18 1406 -4
rect 1428 -8 1618 4
rect 1683 0 1689 20
rect 1413 -18 1443 -8
rect 1444 -18 1602 -8
rect 1606 -18 1636 -8
rect 1640 -18 1670 -4
rect 1698 -18 1711 20
rect 1783 34 1812 50
rect 1826 34 1855 50
rect 1870 40 1900 56
rect 1928 34 1934 82
rect 1937 76 1956 82
rect 1971 76 2001 84
rect 1937 68 2001 76
rect 1937 52 2017 68
rect 2033 61 2095 92
rect 2111 61 2173 92
rect 2242 90 2291 115
rect 2306 90 2336 108
rect 2205 76 2235 84
rect 2242 82 2352 90
rect 2205 68 2250 76
rect 1937 50 1956 52
rect 1971 50 2017 52
rect 1937 34 2017 50
rect 2044 48 2079 61
rect 2120 58 2157 61
rect 2120 56 2162 58
rect 2049 45 2079 48
rect 2058 41 2065 45
rect 2065 40 2066 41
rect 2024 34 2034 40
rect 1783 26 1818 34
rect 1783 0 1784 26
rect 1791 0 1818 26
rect 1726 -18 1756 -4
rect 1783 -8 1818 0
rect 1820 26 1861 34
rect 1820 0 1835 26
rect 1842 0 1861 26
rect 1925 22 1956 34
rect 1971 22 2074 34
rect 2086 24 2112 50
rect 2127 45 2157 56
rect 2189 52 2251 68
rect 2189 50 2235 52
rect 2189 34 2251 50
rect 2263 34 2269 82
rect 2272 74 2352 82
rect 2272 72 2291 74
rect 2306 72 2340 74
rect 2272 57 2352 72
rect 2272 56 2358 57
rect 2272 34 2291 56
rect 2306 40 2336 56
rect 2364 50 2370 124
rect 2373 50 2392 194
rect 2407 50 2413 194
rect 2422 124 2435 194
rect 2487 190 2509 194
rect 2480 178 2497 182
rect 2501 180 2509 182
rect 2499 178 2509 180
rect 2480 168 2509 178
rect 2562 168 2578 182
rect 2616 178 2622 180
rect 2629 178 2737 194
rect 2744 178 2750 180
rect 2758 178 2773 194
rect 2839 188 2858 191
rect 2480 166 2578 168
rect 2605 166 2773 178
rect 2788 168 2804 182
rect 2839 169 2861 188
rect 2871 182 2887 183
rect 2870 176 2887 182
rect 2871 175 2887 176
rect 2861 168 2867 169
rect 2870 168 2899 175
rect 2788 167 2899 168
rect 2788 166 2905 167
rect 2464 158 2515 166
rect 2562 158 2596 166
rect 2464 146 2489 158
rect 2496 146 2515 158
rect 2569 156 2596 158
rect 2605 156 2826 166
rect 2861 163 2867 166
rect 2569 152 2826 156
rect 2464 138 2515 146
rect 2562 138 2826 152
rect 2870 158 2905 166
rect 2416 90 2435 124
rect 2480 130 2509 138
rect 2480 124 2497 130
rect 2480 122 2514 124
rect 2562 122 2578 138
rect 2579 128 2787 138
rect 2788 128 2804 138
rect 2852 134 2867 149
rect 2870 146 2871 158
rect 2878 146 2905 158
rect 2870 138 2905 146
rect 2870 137 2899 138
rect 2590 124 2804 128
rect 2605 122 2804 124
rect 2839 124 2852 134
rect 2870 124 2887 137
rect 2839 122 2887 124
rect 2481 118 2514 122
rect 2477 116 2514 118
rect 2477 115 2544 116
rect 2477 110 2508 115
rect 2514 110 2544 115
rect 2477 106 2544 110
rect 2450 103 2544 106
rect 2450 96 2499 103
rect 2450 90 2480 96
rect 2499 91 2504 96
rect 2416 74 2496 90
rect 2508 82 2544 103
rect 2605 98 2794 122
rect 2839 121 2886 122
rect 2852 116 2886 121
rect 2926 116 2942 118
rect 2620 95 2794 98
rect 2613 92 2794 95
rect 2822 115 2886 116
rect 2416 72 2435 74
rect 2450 72 2484 74
rect 2416 56 2496 72
rect 2416 50 2435 56
rect 2132 24 2235 34
rect 2086 22 2235 24
rect 2256 22 2291 34
rect 1925 20 2087 22
rect 1937 0 1956 20
rect 1971 18 2001 20
rect 1820 -8 1861 0
rect 1943 -4 1956 0
rect 2008 4 2087 20
rect 2119 20 2291 22
rect 2119 4 2198 20
rect 2205 18 2235 20
rect 1783 -18 1812 -8
rect 1826 -18 1855 -8
rect 1870 -18 1900 -4
rect 1943 -18 1986 -4
rect 2008 -8 2198 4
rect 2263 0 2269 20
rect 1993 -18 2023 -8
rect 2024 -18 2182 -8
rect 2186 -18 2216 -8
rect 2220 -18 2250 -4
rect 2278 -18 2291 20
rect 2363 34 2392 50
rect 2406 34 2435 50
rect 2450 40 2480 56
rect 2508 34 2514 82
rect 2517 76 2536 82
rect 2551 76 2581 84
rect 2517 68 2581 76
rect 2517 52 2597 68
rect 2613 61 2675 92
rect 2691 61 2753 92
rect 2822 90 2871 115
rect 2916 106 2942 116
rect 2886 90 2942 106
rect 2785 76 2815 84
rect 2822 82 2932 90
rect 2785 68 2830 76
rect 2517 50 2536 52
rect 2551 50 2597 52
rect 2517 34 2597 50
rect 2624 48 2659 61
rect 2700 58 2737 61
rect 2700 56 2742 58
rect 2629 45 2659 48
rect 2638 41 2645 45
rect 2645 40 2646 41
rect 2604 34 2614 40
rect 2363 26 2398 34
rect 2363 0 2364 26
rect 2371 0 2398 26
rect 2306 -18 2336 -4
rect 2363 -8 2398 0
rect 2400 26 2441 34
rect 2400 0 2415 26
rect 2422 0 2441 26
rect 2505 22 2536 34
rect 2551 22 2654 34
rect 2666 24 2692 50
rect 2707 45 2737 56
rect 2769 52 2831 68
rect 2769 50 2815 52
rect 2769 34 2831 50
rect 2843 34 2849 82
rect 2852 74 2932 82
rect 2852 72 2871 74
rect 2886 72 2920 74
rect 2852 56 2932 72
rect 2852 34 2871 56
rect 2886 40 2916 56
rect 2944 50 2950 124
rect 2953 50 2972 194
rect 2987 50 2993 194
rect 3002 124 3015 194
rect 3067 190 3089 194
rect 3060 178 3077 182
rect 3081 180 3089 182
rect 3079 178 3089 180
rect 3060 168 3089 178
rect 3142 168 3158 182
rect 3196 178 3202 180
rect 3209 178 3317 194
rect 3324 178 3330 180
rect 3338 178 3353 194
rect 3419 188 3438 191
rect 3060 166 3158 168
rect 3185 166 3353 178
rect 3368 168 3384 182
rect 3419 169 3441 188
rect 3451 182 3467 183
rect 3450 176 3467 182
rect 3451 175 3467 176
rect 3441 168 3447 169
rect 3450 168 3479 175
rect 3368 167 3479 168
rect 3368 166 3485 167
rect 3044 158 3095 166
rect 3142 158 3176 166
rect 3044 146 3069 158
rect 3076 146 3095 158
rect 3149 156 3176 158
rect 3185 156 3406 166
rect 3441 163 3447 166
rect 3149 152 3406 156
rect 3044 138 3095 146
rect 3142 138 3406 152
rect 3450 158 3485 166
rect 2996 90 3015 124
rect 3060 130 3089 138
rect 3060 124 3077 130
rect 3060 122 3094 124
rect 3142 122 3158 138
rect 3159 128 3367 138
rect 3368 128 3384 138
rect 3432 134 3447 149
rect 3450 146 3451 158
rect 3458 146 3485 158
rect 3450 138 3485 146
rect 3450 137 3479 138
rect 3170 124 3384 128
rect 3185 122 3384 124
rect 3419 124 3432 134
rect 3450 124 3467 137
rect 3419 122 3467 124
rect 3061 118 3094 122
rect 3057 116 3094 118
rect 3057 115 3124 116
rect 3057 110 3088 115
rect 3094 110 3124 115
rect 3057 106 3124 110
rect 3030 103 3124 106
rect 3030 96 3079 103
rect 3030 90 3060 96
rect 3079 91 3084 96
rect 2996 74 3076 90
rect 3088 82 3124 103
rect 3185 98 3374 122
rect 3419 121 3466 122
rect 3432 116 3466 121
rect 3200 95 3374 98
rect 3193 92 3374 95
rect 3402 115 3466 116
rect 2996 72 3015 74
rect 3030 72 3064 74
rect 2996 56 3076 72
rect 2996 50 3015 56
rect 2712 24 2815 34
rect 2666 22 2815 24
rect 2836 22 2871 34
rect 2505 20 2667 22
rect 2517 0 2536 20
rect 2551 18 2581 20
rect 2400 -8 2441 0
rect 2523 -4 2536 0
rect 2588 4 2667 20
rect 2699 20 2871 22
rect 2699 4 2778 20
rect 2785 18 2815 20
rect 2363 -18 2392 -8
rect 2406 -18 2435 -8
rect 2450 -18 2480 -4
rect 2523 -18 2566 -4
rect 2588 -8 2778 4
rect 2843 0 2849 20
rect 2573 -18 2603 -8
rect 2604 -18 2762 -8
rect 2766 -18 2796 -8
rect 2800 -18 2830 -4
rect 2858 -18 2871 20
rect 2943 34 2972 50
rect 2986 34 3015 50
rect 3030 40 3060 56
rect 3088 34 3094 82
rect 3097 76 3116 82
rect 3131 76 3161 84
rect 3097 68 3161 76
rect 3097 52 3177 68
rect 3193 61 3255 92
rect 3271 61 3333 92
rect 3402 90 3451 115
rect 3466 90 3496 108
rect 3365 76 3395 84
rect 3402 82 3512 90
rect 3365 68 3410 76
rect 3097 50 3116 52
rect 3131 50 3177 52
rect 3097 34 3177 50
rect 3204 48 3239 61
rect 3280 58 3317 61
rect 3280 56 3322 58
rect 3209 45 3239 48
rect 3218 41 3225 45
rect 3225 40 3226 41
rect 3184 34 3194 40
rect 2943 26 2978 34
rect 2943 0 2944 26
rect 2951 0 2978 26
rect 2886 -18 2916 -4
rect 2943 -8 2978 0
rect 2980 26 3021 34
rect 2980 0 2995 26
rect 3002 0 3021 26
rect 3085 22 3116 34
rect 3131 22 3234 34
rect 3246 24 3272 50
rect 3287 45 3317 56
rect 3349 52 3411 68
rect 3349 50 3395 52
rect 3349 34 3411 50
rect 3423 34 3429 82
rect 3432 74 3512 82
rect 3432 72 3451 74
rect 3466 72 3500 74
rect 3432 57 3512 72
rect 3432 56 3518 57
rect 3432 34 3451 56
rect 3466 40 3496 56
rect 3524 50 3530 124
rect 3533 50 3552 194
rect 3567 50 3573 194
rect 3582 124 3595 194
rect 3647 190 3669 194
rect 3640 178 3657 182
rect 3661 180 3669 182
rect 3659 178 3669 180
rect 3640 168 3669 178
rect 3722 168 3738 182
rect 3776 178 3782 180
rect 3789 178 3897 194
rect 3904 178 3910 180
rect 3918 178 3933 194
rect 3999 188 4018 191
rect 3640 166 3738 168
rect 3765 166 3933 178
rect 3948 168 3964 182
rect 3999 169 4021 188
rect 4031 182 4047 183
rect 4030 176 4047 182
rect 4031 175 4047 176
rect 4021 168 4027 169
rect 4030 168 4059 175
rect 3948 167 4059 168
rect 3948 166 4065 167
rect 3624 158 3675 166
rect 3722 158 3756 166
rect 3624 146 3649 158
rect 3656 146 3675 158
rect 3729 156 3756 158
rect 3765 156 3986 166
rect 4021 163 4027 166
rect 3729 152 3986 156
rect 3624 138 3675 146
rect 3722 138 3986 152
rect 4030 158 4065 166
rect 3576 90 3595 124
rect 3640 130 3669 138
rect 3640 124 3657 130
rect 3640 122 3674 124
rect 3722 122 3738 138
rect 3739 128 3947 138
rect 3948 128 3964 138
rect 4012 134 4027 149
rect 4030 146 4031 158
rect 4038 146 4065 158
rect 4030 138 4065 146
rect 4030 137 4059 138
rect 3750 124 3964 128
rect 3765 122 3964 124
rect 3999 124 4012 134
rect 4030 124 4047 137
rect 3999 122 4047 124
rect 3641 118 3674 122
rect 3637 116 3674 118
rect 3637 115 3704 116
rect 3637 110 3668 115
rect 3674 110 3704 115
rect 3637 106 3704 110
rect 3610 103 3704 106
rect 3610 96 3659 103
rect 3610 90 3640 96
rect 3659 91 3664 96
rect 3576 74 3656 90
rect 3668 82 3704 103
rect 3765 98 3954 122
rect 3999 121 4046 122
rect 4012 116 4046 121
rect 4086 116 4102 118
rect 3780 95 3954 98
rect 3773 92 3954 95
rect 3982 115 4046 116
rect 3576 72 3595 74
rect 3610 72 3644 74
rect 3576 56 3656 72
rect 3576 50 3595 56
rect 3292 24 3395 34
rect 3246 22 3395 24
rect 3416 22 3451 34
rect 3085 20 3247 22
rect 3097 0 3116 20
rect 3131 18 3161 20
rect 2980 -8 3021 0
rect 3103 -4 3116 0
rect 3168 4 3247 20
rect 3279 20 3451 22
rect 3279 4 3358 20
rect 3365 18 3395 20
rect 2943 -18 2972 -8
rect 2986 -18 3015 -8
rect 3030 -18 3060 -4
rect 3103 -18 3146 -4
rect 3168 -8 3358 4
rect 3423 0 3429 20
rect 3153 -18 3183 -8
rect 3184 -18 3342 -8
rect 3346 -18 3376 -8
rect 3380 -18 3410 -4
rect 3438 -18 3451 20
rect 3523 34 3552 50
rect 3566 34 3595 50
rect 3610 40 3640 56
rect 3668 34 3674 82
rect 3677 76 3696 82
rect 3711 76 3741 84
rect 3677 68 3741 76
rect 3677 52 3757 68
rect 3773 61 3835 92
rect 3851 61 3913 92
rect 3982 90 4031 115
rect 4076 106 4102 116
rect 4046 90 4102 106
rect 3945 76 3975 84
rect 3982 82 4092 90
rect 3945 68 3990 76
rect 3677 50 3696 52
rect 3711 50 3757 52
rect 3677 34 3757 50
rect 3784 48 3819 61
rect 3860 58 3897 61
rect 3860 56 3902 58
rect 3789 45 3819 48
rect 3798 41 3805 45
rect 3805 40 3806 41
rect 3764 34 3774 40
rect 3523 26 3558 34
rect 3523 0 3524 26
rect 3531 0 3558 26
rect 3466 -18 3496 -4
rect 3523 -8 3558 0
rect 3560 26 3601 34
rect 3560 0 3575 26
rect 3582 0 3601 26
rect 3665 22 3696 34
rect 3711 22 3814 34
rect 3826 24 3852 50
rect 3867 45 3897 56
rect 3929 52 3991 68
rect 3929 50 3975 52
rect 3929 34 3991 50
rect 4003 34 4009 82
rect 4012 74 4092 82
rect 4012 72 4031 74
rect 4046 72 4080 74
rect 4012 56 4092 72
rect 4012 34 4031 56
rect 4046 40 4076 56
rect 4104 50 4110 124
rect 4113 50 4132 194
rect 4147 50 4153 194
rect 4162 124 4175 194
rect 4227 190 4249 194
rect 4220 178 4237 182
rect 4241 180 4249 182
rect 4239 178 4249 180
rect 4220 168 4249 178
rect 4302 168 4318 182
rect 4356 178 4362 180
rect 4369 178 4477 194
rect 4484 178 4490 180
rect 4498 178 4513 194
rect 4579 188 4598 191
rect 4220 166 4318 168
rect 4345 166 4513 178
rect 4528 168 4544 182
rect 4579 169 4601 188
rect 4611 182 4627 183
rect 4610 176 4627 182
rect 4611 175 4627 176
rect 4601 168 4607 169
rect 4610 168 4639 175
rect 4528 167 4639 168
rect 4528 166 4645 167
rect 4204 158 4255 166
rect 4302 158 4336 166
rect 4204 146 4229 158
rect 4236 146 4255 158
rect 4309 156 4336 158
rect 4345 156 4566 166
rect 4601 163 4607 166
rect 4309 152 4566 156
rect 4204 138 4255 146
rect 4302 138 4566 152
rect 4610 158 4645 166
rect 4156 90 4175 124
rect 4220 130 4249 138
rect 4220 124 4237 130
rect 4220 122 4254 124
rect 4302 122 4318 138
rect 4319 128 4527 138
rect 4528 128 4544 138
rect 4592 134 4607 149
rect 4610 146 4611 158
rect 4618 146 4645 158
rect 4610 138 4645 146
rect 4610 137 4639 138
rect 4330 124 4544 128
rect 4345 122 4544 124
rect 4579 124 4592 134
rect 4610 124 4627 137
rect 4579 122 4627 124
rect 4221 118 4254 122
rect 4217 116 4254 118
rect 4217 115 4284 116
rect 4217 110 4248 115
rect 4254 110 4284 115
rect 4217 106 4284 110
rect 4190 103 4284 106
rect 4190 96 4239 103
rect 4190 90 4220 96
rect 4239 91 4244 96
rect 4156 74 4236 90
rect 4248 82 4284 103
rect 4345 98 4534 122
rect 4579 121 4626 122
rect 4592 116 4626 121
rect 4360 95 4534 98
rect 4353 92 4534 95
rect 4562 115 4626 116
rect 4156 72 4175 74
rect 4190 72 4224 74
rect 4156 56 4236 72
rect 4156 50 4175 56
rect 3872 24 3975 34
rect 3826 22 3975 24
rect 3996 22 4031 34
rect 3665 20 3827 22
rect 3677 0 3696 20
rect 3711 18 3741 20
rect 3560 -8 3601 0
rect 3683 -4 3696 0
rect 3748 4 3827 20
rect 3859 20 4031 22
rect 3859 4 3938 20
rect 3945 18 3975 20
rect 3523 -18 3552 -8
rect 3566 -18 3595 -8
rect 3610 -18 3640 -4
rect 3683 -18 3726 -4
rect 3748 -8 3938 4
rect 4003 0 4009 20
rect 3733 -18 3763 -8
rect 3764 -18 3922 -8
rect 3926 -18 3956 -8
rect 3960 -18 3990 -4
rect 4018 -18 4031 20
rect 4103 34 4132 50
rect 4146 34 4175 50
rect 4190 40 4220 56
rect 4248 34 4254 82
rect 4257 76 4276 82
rect 4291 76 4321 84
rect 4257 68 4321 76
rect 4257 52 4337 68
rect 4353 61 4415 92
rect 4431 61 4493 92
rect 4562 90 4611 115
rect 4626 90 4656 108
rect 4525 76 4555 84
rect 4562 82 4672 90
rect 4525 68 4570 76
rect 4257 50 4276 52
rect 4291 50 4337 52
rect 4257 34 4337 50
rect 4364 48 4399 61
rect 4440 58 4477 61
rect 4440 56 4482 58
rect 4369 45 4399 48
rect 4378 41 4385 45
rect 4385 40 4386 41
rect 4344 34 4354 40
rect 4103 26 4138 34
rect 4103 0 4104 26
rect 4111 0 4138 26
rect 4046 -18 4076 -4
rect 4103 -8 4138 0
rect 4140 26 4181 34
rect 4140 0 4155 26
rect 4162 0 4181 26
rect 4245 22 4276 34
rect 4291 22 4394 34
rect 4406 24 4432 50
rect 4447 45 4477 56
rect 4509 52 4571 68
rect 4509 50 4555 52
rect 4509 34 4571 50
rect 4583 34 4589 82
rect 4592 74 4672 82
rect 4592 72 4611 74
rect 4626 72 4660 74
rect 4592 57 4672 72
rect 4592 56 4678 57
rect 4592 34 4611 56
rect 4626 40 4656 56
rect 4684 50 4690 124
rect 4693 50 4712 194
rect 4727 50 4733 194
rect 4742 124 4755 194
rect 4807 190 4829 194
rect 4800 178 4817 182
rect 4821 180 4829 182
rect 4819 178 4829 180
rect 4800 168 4829 178
rect 4882 168 4898 182
rect 4936 178 4942 180
rect 4949 178 5057 194
rect 5064 178 5070 180
rect 5078 178 5093 194
rect 5159 188 5178 191
rect 4800 166 4898 168
rect 4925 166 5093 178
rect 5108 168 5124 182
rect 5159 169 5181 188
rect 5191 182 5207 183
rect 5190 176 5207 182
rect 5191 175 5207 176
rect 5181 168 5187 169
rect 5190 168 5219 175
rect 5108 167 5219 168
rect 5108 166 5225 167
rect 4784 158 4835 166
rect 4882 158 4916 166
rect 4784 146 4809 158
rect 4816 146 4835 158
rect 4889 156 4916 158
rect 4925 156 5146 166
rect 5181 163 5187 166
rect 4889 152 5146 156
rect 4784 138 4835 146
rect 4882 138 5146 152
rect 5190 158 5225 166
rect 4736 90 4755 124
rect 4800 130 4829 138
rect 4800 124 4817 130
rect 4800 122 4834 124
rect 4882 122 4898 138
rect 4899 128 5107 138
rect 5108 128 5124 138
rect 5172 134 5187 149
rect 5190 146 5191 158
rect 5198 146 5225 158
rect 5190 138 5225 146
rect 5190 137 5219 138
rect 4910 124 5124 128
rect 4925 122 5124 124
rect 5159 124 5172 134
rect 5190 124 5207 137
rect 5159 122 5207 124
rect 4801 118 4834 122
rect 4797 116 4834 118
rect 4797 115 4864 116
rect 4797 110 4828 115
rect 4834 110 4864 115
rect 4797 106 4864 110
rect 4770 103 4864 106
rect 4770 96 4819 103
rect 4770 90 4800 96
rect 4819 91 4824 96
rect 4736 74 4816 90
rect 4828 82 4864 103
rect 4925 98 5114 122
rect 5159 121 5206 122
rect 5172 116 5206 121
rect 5246 116 5262 118
rect 4940 95 5114 98
rect 4933 92 5114 95
rect 5142 115 5206 116
rect 4736 72 4755 74
rect 4770 72 4804 74
rect 4736 56 4816 72
rect 4736 50 4755 56
rect 4452 24 4555 34
rect 4406 22 4555 24
rect 4576 22 4611 34
rect 4245 20 4407 22
rect 4257 0 4276 20
rect 4291 18 4321 20
rect 4140 -8 4181 0
rect 4263 -4 4276 0
rect 4328 4 4407 20
rect 4439 20 4611 22
rect 4439 4 4518 20
rect 4525 18 4555 20
rect 4103 -18 4132 -8
rect 4146 -18 4175 -8
rect 4190 -18 4220 -4
rect 4263 -18 4306 -4
rect 4328 -8 4518 4
rect 4583 0 4589 20
rect 4313 -18 4343 -8
rect 4344 -18 4502 -8
rect 4506 -18 4536 -8
rect 4540 -18 4570 -4
rect 4598 -18 4611 20
rect 4683 34 4712 50
rect 4726 34 4755 50
rect 4770 40 4800 56
rect 4828 34 4834 82
rect 4837 76 4856 82
rect 4871 76 4901 84
rect 4837 68 4901 76
rect 4837 52 4917 68
rect 4933 61 4995 92
rect 5011 61 5073 92
rect 5142 90 5191 115
rect 5236 106 5262 116
rect 5206 90 5262 106
rect 5105 76 5135 84
rect 5142 82 5252 90
rect 5105 68 5150 76
rect 4837 50 4856 52
rect 4871 50 4917 52
rect 4837 34 4917 50
rect 4944 48 4979 61
rect 5020 58 5057 61
rect 5020 56 5062 58
rect 4949 45 4979 48
rect 4958 41 4965 45
rect 4965 40 4966 41
rect 4924 34 4934 40
rect 4683 26 4718 34
rect 4683 0 4684 26
rect 4691 0 4718 26
rect 4626 -18 4656 -4
rect 4683 -8 4718 0
rect 4720 26 4761 34
rect 4720 0 4735 26
rect 4742 0 4761 26
rect 4825 22 4856 34
rect 4871 22 4974 34
rect 4986 24 5012 50
rect 5027 45 5057 56
rect 5089 52 5151 68
rect 5089 50 5135 52
rect 5089 34 5151 50
rect 5163 34 5169 82
rect 5172 74 5252 82
rect 5172 72 5191 74
rect 5206 72 5240 74
rect 5172 56 5252 72
rect 5172 34 5191 56
rect 5206 40 5236 56
rect 5264 50 5270 124
rect 5273 50 5292 194
rect 5307 50 5313 194
rect 5322 124 5335 194
rect 5387 190 5409 194
rect 5380 178 5397 182
rect 5401 180 5409 182
rect 5399 178 5409 180
rect 5380 168 5409 178
rect 5462 168 5478 182
rect 5516 178 5522 180
rect 5529 178 5637 194
rect 5644 178 5650 180
rect 5658 178 5673 194
rect 5739 188 5758 191
rect 5380 166 5478 168
rect 5505 166 5673 178
rect 5688 168 5704 182
rect 5739 169 5761 188
rect 5771 182 5787 183
rect 5770 176 5787 182
rect 5771 175 5787 176
rect 5761 168 5767 169
rect 5770 168 5799 175
rect 5688 167 5799 168
rect 5688 166 5805 167
rect 5364 158 5415 166
rect 5462 158 5496 166
rect 5364 146 5389 158
rect 5396 146 5415 158
rect 5469 156 5496 158
rect 5505 156 5726 166
rect 5761 163 5767 166
rect 5469 152 5726 156
rect 5364 138 5415 146
rect 5462 138 5726 152
rect 5770 158 5805 166
rect 5316 90 5335 124
rect 5380 130 5409 138
rect 5380 124 5397 130
rect 5380 122 5414 124
rect 5462 122 5478 138
rect 5479 128 5687 138
rect 5688 128 5704 138
rect 5752 134 5767 149
rect 5770 146 5771 158
rect 5778 146 5805 158
rect 5770 138 5805 146
rect 5770 137 5799 138
rect 5490 124 5704 128
rect 5505 122 5704 124
rect 5739 124 5752 134
rect 5770 124 5787 137
rect 5739 122 5787 124
rect 5381 118 5414 122
rect 5377 116 5414 118
rect 5377 115 5444 116
rect 5377 110 5408 115
rect 5414 110 5444 115
rect 5377 106 5444 110
rect 5350 103 5444 106
rect 5350 96 5399 103
rect 5350 90 5380 96
rect 5399 91 5404 96
rect 5316 74 5396 90
rect 5408 82 5444 103
rect 5505 98 5694 122
rect 5739 121 5786 122
rect 5752 116 5786 121
rect 5520 95 5694 98
rect 5513 92 5694 95
rect 5722 115 5786 116
rect 5316 72 5335 74
rect 5350 72 5384 74
rect 5316 56 5396 72
rect 5316 50 5335 56
rect 5032 24 5135 34
rect 4986 22 5135 24
rect 5156 22 5191 34
rect 4825 20 4987 22
rect 4837 0 4856 20
rect 4871 18 4901 20
rect 4720 -8 4761 0
rect 4843 -4 4856 0
rect 4908 4 4987 20
rect 5019 20 5191 22
rect 5019 4 5098 20
rect 5105 18 5135 20
rect 4683 -18 4712 -8
rect 4726 -18 4755 -8
rect 4770 -18 4800 -4
rect 4843 -18 4886 -4
rect 4908 -8 5098 4
rect 5163 0 5169 20
rect 4893 -18 4923 -8
rect 4924 -18 5082 -8
rect 5086 -18 5116 -8
rect 5120 -18 5150 -4
rect 5178 -18 5191 20
rect 5263 34 5292 50
rect 5306 34 5335 50
rect 5350 40 5380 56
rect 5408 34 5414 82
rect 5417 76 5436 82
rect 5451 76 5481 84
rect 5417 68 5481 76
rect 5417 52 5497 68
rect 5513 61 5575 92
rect 5591 61 5653 92
rect 5722 90 5771 115
rect 5786 90 5816 108
rect 5685 76 5715 84
rect 5722 82 5832 90
rect 5685 68 5730 76
rect 5417 50 5436 52
rect 5451 50 5497 52
rect 5417 34 5497 50
rect 5524 48 5559 61
rect 5600 58 5637 61
rect 5600 56 5642 58
rect 5529 45 5559 48
rect 5538 41 5545 45
rect 5545 40 5546 41
rect 5504 34 5514 40
rect 5263 26 5298 34
rect 5263 0 5264 26
rect 5271 0 5298 26
rect 5206 -18 5236 -4
rect 5263 -8 5298 0
rect 5300 26 5341 34
rect 5300 0 5315 26
rect 5322 0 5341 26
rect 5405 22 5436 34
rect 5451 22 5554 34
rect 5566 24 5592 50
rect 5607 45 5637 56
rect 5669 52 5731 68
rect 5669 50 5715 52
rect 5669 34 5731 50
rect 5743 34 5749 82
rect 5752 74 5832 82
rect 5752 72 5771 74
rect 5786 72 5820 74
rect 5752 57 5832 72
rect 5752 56 5838 57
rect 5752 34 5771 56
rect 5786 40 5816 56
rect 5844 50 5850 124
rect 5853 50 5872 194
rect 5887 50 5893 194
rect 5902 124 5915 194
rect 5967 190 5989 194
rect 5960 178 5977 182
rect 5981 180 5989 182
rect 5979 178 5989 180
rect 5960 168 5989 178
rect 6042 168 6058 182
rect 6096 178 6102 180
rect 6109 178 6217 194
rect 6224 178 6230 180
rect 6238 178 6253 194
rect 6319 188 6338 191
rect 5960 166 6058 168
rect 6085 166 6253 178
rect 6268 168 6284 182
rect 6319 169 6341 188
rect 6351 182 6367 183
rect 6350 176 6367 182
rect 6351 175 6367 176
rect 6341 168 6347 169
rect 6350 168 6379 175
rect 6268 167 6379 168
rect 6268 166 6385 167
rect 5944 158 5995 166
rect 6042 158 6076 166
rect 5944 146 5969 158
rect 5976 146 5995 158
rect 6049 156 6076 158
rect 6085 156 6306 166
rect 6341 163 6347 166
rect 6049 152 6306 156
rect 5944 138 5995 146
rect 6042 138 6306 152
rect 6350 158 6385 166
rect 5896 90 5915 124
rect 5960 130 5989 138
rect 5960 124 5977 130
rect 5960 122 5994 124
rect 6042 122 6058 138
rect 6059 128 6267 138
rect 6268 128 6284 138
rect 6332 134 6347 149
rect 6350 146 6351 158
rect 6358 146 6385 158
rect 6350 138 6385 146
rect 6350 137 6379 138
rect 6070 124 6284 128
rect 6085 122 6284 124
rect 6319 124 6332 134
rect 6350 124 6367 137
rect 6319 122 6367 124
rect 5961 118 5994 122
rect 5957 116 5994 118
rect 5957 115 6024 116
rect 5957 110 5988 115
rect 5994 110 6024 115
rect 5957 106 6024 110
rect 5930 103 6024 106
rect 5930 96 5979 103
rect 5930 90 5960 96
rect 5979 91 5984 96
rect 5896 74 5976 90
rect 5988 82 6024 103
rect 6085 98 6274 122
rect 6319 121 6366 122
rect 6332 116 6366 121
rect 6100 95 6274 98
rect 6093 92 6274 95
rect 6302 115 6366 116
rect 5896 72 5915 74
rect 5930 72 5964 74
rect 5896 56 5976 72
rect 5896 50 5915 56
rect 5612 24 5715 34
rect 5566 22 5715 24
rect 5736 22 5771 34
rect 5405 20 5567 22
rect 5417 0 5436 20
rect 5451 18 5481 20
rect 5300 -8 5341 0
rect 5423 -4 5436 0
rect 5488 4 5567 20
rect 5599 20 5771 22
rect 5599 4 5678 20
rect 5685 18 5715 20
rect 5263 -18 5292 -8
rect 5306 -18 5335 -8
rect 5350 -18 5380 -4
rect 5423 -18 5466 -4
rect 5488 -8 5678 4
rect 5743 0 5749 20
rect 5473 -18 5503 -8
rect 5504 -18 5662 -8
rect 5666 -18 5696 -8
rect 5700 -18 5730 -4
rect 5758 -18 5771 20
rect 5843 34 5872 50
rect 5886 34 5915 50
rect 5930 40 5960 56
rect 5988 34 5994 82
rect 5997 76 6016 82
rect 6031 76 6061 84
rect 5997 68 6061 76
rect 5997 52 6077 68
rect 6093 61 6155 92
rect 6171 61 6233 92
rect 6302 90 6351 115
rect 6366 90 6396 106
rect 6265 76 6295 84
rect 6302 82 6412 90
rect 6265 68 6310 76
rect 5997 50 6016 52
rect 6031 50 6077 52
rect 5997 34 6077 50
rect 6104 48 6139 61
rect 6180 58 6217 61
rect 6180 56 6222 58
rect 6109 45 6139 48
rect 6118 41 6125 45
rect 6125 40 6126 41
rect 6084 34 6094 40
rect 5843 26 5878 34
rect 5843 0 5844 26
rect 5851 0 5878 26
rect 5786 -18 5816 -4
rect 5843 -8 5878 0
rect 5880 26 5921 34
rect 5880 0 5895 26
rect 5902 0 5921 26
rect 5985 22 6016 34
rect 6031 22 6134 34
rect 6146 24 6172 50
rect 6187 45 6217 56
rect 6249 52 6311 68
rect 6249 50 6295 52
rect 6249 34 6311 50
rect 6323 34 6329 82
rect 6332 74 6412 82
rect 6332 72 6351 74
rect 6366 72 6400 74
rect 6332 56 6412 72
rect 6332 34 6351 56
rect 6366 40 6396 56
rect 6424 50 6430 124
rect 6439 50 6452 194
rect 6192 24 6295 34
rect 6146 22 6295 24
rect 6316 22 6351 34
rect 5985 20 6147 22
rect 5997 0 6016 20
rect 6031 18 6061 20
rect 5880 -8 5921 0
rect 6003 -4 6016 0
rect 6068 4 6147 20
rect 6179 20 6351 22
rect 6179 4 6258 20
rect 6265 18 6295 20
rect 5843 -18 5872 -8
rect 5886 -18 5915 -8
rect 5930 -18 5960 -4
rect 6003 -18 6046 -4
rect 6068 -8 6258 4
rect 6323 0 6329 20
rect 6053 -18 6083 -8
rect 6084 -18 6242 -8
rect 6246 -18 6276 -8
rect 6280 -18 6310 -4
rect 6338 -18 6351 20
rect 6423 34 6452 50
rect 6423 26 6458 34
rect 6423 0 6424 26
rect 6431 0 6458 26
rect 6366 -18 6396 -4
rect 6423 -8 6458 0
rect 6423 -18 6452 -8
rect -541 -32 6452 -18
rect -478 -62 -465 -32
rect -450 -46 -420 -32
rect -377 -46 -334 -32
rect -327 -46 -107 -32
rect -100 -46 -70 -32
rect -410 -60 -395 -48
rect -376 -60 -363 -46
rect -295 -50 -142 -46
rect -413 -62 -391 -60
rect -313 -62 -121 -50
rect -42 -62 -29 -32
rect -14 -46 16 -32
rect 53 -62 72 -32
rect 87 -62 93 -32
rect 102 -62 115 -32
rect 130 -46 160 -32
rect 203 -46 246 -32
rect 253 -46 473 -32
rect 480 -46 510 -32
rect 170 -60 185 -48
rect 204 -60 217 -46
rect 285 -50 438 -46
rect 167 -62 189 -60
rect 267 -62 459 -50
rect 538 -62 551 -32
rect 566 -46 596 -32
rect 633 -62 652 -32
rect 667 -62 673 -32
rect 682 -62 695 -32
rect 710 -46 740 -32
rect 783 -46 826 -32
rect 833 -46 1053 -32
rect 1060 -46 1090 -32
rect 750 -60 765 -48
rect 784 -60 797 -46
rect 865 -50 1018 -46
rect 747 -62 769 -60
rect 847 -62 1039 -50
rect 1118 -62 1131 -32
rect 1146 -46 1176 -32
rect 1213 -62 1232 -32
rect 1247 -62 1253 -32
rect 1262 -62 1275 -32
rect 1290 -46 1320 -32
rect 1363 -46 1406 -32
rect 1413 -46 1633 -32
rect 1640 -46 1670 -32
rect 1330 -60 1345 -48
rect 1364 -60 1377 -46
rect 1445 -50 1598 -46
rect 1327 -62 1349 -60
rect 1427 -62 1619 -50
rect 1698 -62 1711 -32
rect 1726 -46 1756 -32
rect 1793 -62 1812 -32
rect 1827 -62 1833 -32
rect 1842 -62 1855 -32
rect 1870 -46 1900 -32
rect 1943 -46 1986 -32
rect 1993 -46 2213 -32
rect 2220 -46 2250 -32
rect 1910 -60 1925 -48
rect 1944 -60 1957 -46
rect 2025 -50 2178 -46
rect 1907 -62 1929 -60
rect 2007 -62 2199 -50
rect 2278 -62 2291 -32
rect 2306 -46 2336 -32
rect 2373 -62 2392 -32
rect 2407 -62 2413 -32
rect 2422 -62 2435 -32
rect 2450 -46 2480 -32
rect 2523 -46 2566 -32
rect 2573 -46 2793 -32
rect 2800 -46 2830 -32
rect 2490 -60 2505 -48
rect 2524 -60 2537 -46
rect 2605 -50 2758 -46
rect 2487 -62 2509 -60
rect 2587 -62 2779 -50
rect 2858 -62 2871 -32
rect 2886 -46 2916 -32
rect 2953 -62 2972 -32
rect 2987 -62 2993 -32
rect 3002 -62 3015 -32
rect 3030 -46 3060 -32
rect 3103 -46 3146 -32
rect 3153 -46 3373 -32
rect 3380 -46 3410 -32
rect 3070 -60 3085 -48
rect 3104 -60 3117 -46
rect 3185 -50 3338 -46
rect 3067 -62 3089 -60
rect 3167 -62 3359 -50
rect 3438 -62 3451 -32
rect 3466 -46 3496 -32
rect 3533 -62 3552 -32
rect 3567 -62 3573 -32
rect 3582 -62 3595 -32
rect 3610 -46 3640 -32
rect 3683 -46 3726 -32
rect 3733 -46 3953 -32
rect 3960 -46 3990 -32
rect 3650 -60 3665 -48
rect 3684 -60 3697 -46
rect 3765 -50 3918 -46
rect 3647 -62 3669 -60
rect 3747 -62 3939 -50
rect 4018 -62 4031 -32
rect 4046 -46 4076 -32
rect 4113 -62 4132 -32
rect 4147 -62 4153 -32
rect 4162 -62 4175 -32
rect 4190 -46 4220 -32
rect 4263 -46 4306 -32
rect 4313 -46 4533 -32
rect 4540 -46 4570 -32
rect 4230 -60 4245 -48
rect 4264 -60 4277 -46
rect 4345 -50 4498 -46
rect 4227 -62 4249 -60
rect 4327 -62 4519 -50
rect 4598 -62 4611 -32
rect 4626 -46 4656 -32
rect 4693 -62 4712 -32
rect 4727 -62 4733 -32
rect 4742 -62 4755 -32
rect 4770 -46 4800 -32
rect 4843 -46 4886 -32
rect 4893 -46 5113 -32
rect 5120 -46 5150 -32
rect 4810 -60 4825 -48
rect 4844 -60 4857 -46
rect 4925 -50 5078 -46
rect 4807 -62 4829 -60
rect 4907 -62 5099 -50
rect 5178 -62 5191 -32
rect 5206 -46 5236 -32
rect 5273 -62 5292 -32
rect 5307 -62 5313 -32
rect 5322 -62 5335 -32
rect 5350 -46 5380 -32
rect 5423 -46 5466 -32
rect 5473 -46 5693 -32
rect 5700 -46 5730 -32
rect 5390 -60 5405 -48
rect 5424 -60 5437 -46
rect 5505 -50 5658 -46
rect 5387 -62 5409 -60
rect 5487 -62 5679 -50
rect 5758 -62 5771 -32
rect 5786 -46 5816 -32
rect 5853 -62 5872 -32
rect 5887 -62 5893 -32
rect 5902 -62 5915 -32
rect 5930 -46 5960 -32
rect 6003 -46 6046 -32
rect 6053 -46 6273 -32
rect 6280 -46 6310 -32
rect 5970 -60 5985 -48
rect 6004 -60 6017 -46
rect 6085 -50 6238 -46
rect 5967 -62 5989 -60
rect 6067 -62 6259 -50
rect 6338 -62 6351 -32
rect 6366 -46 6396 -32
rect 6439 -62 6452 -32
rect -541 -76 6452 -62
rect -478 -146 -465 -76
rect -413 -80 -391 -76
rect -420 -92 -403 -88
rect -399 -90 -391 -88
rect -401 -92 -391 -90
rect -420 -102 -391 -92
rect -338 -102 -322 -88
rect -284 -92 -278 -90
rect -271 -92 -163 -76
rect -156 -92 -150 -90
rect -142 -92 -127 -76
rect -61 -82 -42 -79
rect -420 -104 -322 -102
rect -295 -104 -127 -92
rect -112 -102 -96 -88
rect -61 -101 -39 -82
rect -29 -88 -13 -87
rect -30 -90 -13 -88
rect -29 -95 -13 -90
rect -39 -102 -33 -101
rect -30 -102 -1 -95
rect -112 -103 -1 -102
rect -112 -104 5 -103
rect -436 -112 -385 -104
rect -338 -112 -304 -104
rect -436 -124 -411 -112
rect -404 -124 -385 -112
rect -331 -114 -304 -112
rect -295 -114 -74 -104
rect -39 -107 -33 -104
rect -331 -118 -74 -114
rect -436 -132 -385 -124
rect -338 -132 -74 -118
rect -30 -112 5 -104
rect -484 -180 -465 -146
rect -420 -140 -391 -132
rect -420 -146 -403 -140
rect -420 -148 -386 -146
rect -338 -148 -322 -132
rect -321 -142 -113 -132
rect -112 -142 -96 -132
rect -48 -136 -33 -121
rect -30 -124 -29 -112
rect -22 -124 5 -112
rect -30 -132 5 -124
rect -30 -133 -1 -132
rect -310 -146 -96 -142
rect -295 -148 -96 -146
rect -61 -146 -48 -136
rect -30 -146 -13 -133
rect -61 -148 -13 -146
rect -419 -152 -386 -148
rect -423 -154 -386 -152
rect -423 -155 -356 -154
rect -423 -160 -392 -155
rect -386 -160 -356 -155
rect -423 -164 -356 -160
rect -450 -167 -356 -164
rect -450 -174 -401 -167
rect -450 -180 -420 -174
rect -401 -179 -396 -174
rect -484 -196 -404 -180
rect -392 -188 -356 -167
rect -295 -172 -106 -148
rect -61 -149 -14 -148
rect -48 -154 -14 -149
rect -280 -175 -106 -172
rect -287 -178 -106 -175
rect -78 -155 -14 -154
rect -484 -198 -465 -196
rect -450 -198 -416 -196
rect -484 -214 -404 -198
rect -484 -220 -465 -214
rect -494 -236 -465 -220
rect -450 -230 -420 -214
rect -392 -236 -386 -188
rect -383 -194 -364 -188
rect -349 -194 -319 -186
rect -383 -202 -319 -194
rect -383 -218 -303 -202
rect -287 -209 -225 -178
rect -209 -209 -147 -178
rect -78 -180 -29 -155
rect -14 -180 16 -162
rect -115 -194 -85 -186
rect -78 -188 32 -180
rect -115 -202 -70 -194
rect -383 -220 -364 -218
rect -349 -220 -303 -218
rect -383 -236 -303 -220
rect -276 -222 -241 -209
rect -200 -212 -163 -209
rect -200 -214 -158 -212
rect -271 -225 -241 -222
rect -262 -229 -255 -225
rect -255 -230 -254 -229
rect -296 -236 -286 -230
rect -500 -244 -459 -236
rect -500 -270 -485 -244
rect -478 -270 -459 -244
rect -395 -248 -364 -236
rect -349 -248 -246 -236
rect -234 -246 -208 -220
rect -193 -225 -163 -214
rect -131 -218 -69 -202
rect -131 -220 -85 -218
rect -131 -236 -69 -220
rect -57 -236 -51 -188
rect -48 -196 32 -188
rect -48 -198 -29 -196
rect -14 -198 20 -196
rect -48 -213 32 -198
rect -48 -214 38 -213
rect -48 -236 -29 -214
rect -14 -230 16 -214
rect 44 -220 50 -146
rect 53 -220 72 -76
rect 87 -220 93 -76
rect 102 -146 115 -76
rect 167 -80 189 -76
rect 160 -92 177 -88
rect 181 -90 189 -88
rect 179 -92 189 -90
rect 160 -102 189 -92
rect 242 -102 258 -88
rect 296 -92 302 -90
rect 309 -92 417 -76
rect 424 -92 430 -90
rect 438 -92 453 -76
rect 519 -82 538 -79
rect 160 -104 258 -102
rect 285 -104 453 -92
rect 468 -102 484 -88
rect 519 -101 541 -82
rect 551 -88 567 -87
rect 550 -90 567 -88
rect 551 -95 567 -90
rect 541 -102 547 -101
rect 550 -102 579 -95
rect 468 -103 579 -102
rect 468 -104 585 -103
rect 144 -112 195 -104
rect 242 -112 276 -104
rect 144 -124 169 -112
rect 176 -124 195 -112
rect 249 -114 276 -112
rect 285 -114 506 -104
rect 541 -107 547 -104
rect 249 -118 506 -114
rect 144 -132 195 -124
rect 242 -132 506 -118
rect 550 -112 585 -104
rect 96 -180 115 -146
rect 160 -140 189 -132
rect 160 -146 177 -140
rect 160 -148 194 -146
rect 242 -148 258 -132
rect 259 -142 467 -132
rect 468 -142 484 -132
rect 532 -136 547 -121
rect 550 -124 551 -112
rect 558 -124 585 -112
rect 550 -132 585 -124
rect 550 -133 579 -132
rect 270 -146 484 -142
rect 285 -148 484 -146
rect 519 -146 532 -136
rect 550 -146 567 -133
rect 519 -148 567 -146
rect 161 -152 194 -148
rect 157 -154 194 -152
rect 157 -155 224 -154
rect 157 -160 188 -155
rect 194 -160 224 -155
rect 157 -164 224 -160
rect 130 -167 224 -164
rect 130 -174 179 -167
rect 130 -180 160 -174
rect 179 -179 184 -174
rect 96 -196 176 -180
rect 188 -188 224 -167
rect 285 -172 474 -148
rect 519 -149 566 -148
rect 532 -154 566 -149
rect 606 -154 622 -152
rect 300 -175 474 -172
rect 293 -178 474 -175
rect 502 -155 566 -154
rect 96 -198 115 -196
rect 130 -198 164 -196
rect 96 -214 176 -198
rect 96 -220 115 -214
rect -188 -246 -85 -236
rect -234 -248 -85 -246
rect -64 -248 -29 -236
rect -395 -250 -233 -248
rect -383 -268 -364 -250
rect -349 -252 -319 -250
rect -500 -278 -459 -270
rect -376 -274 -364 -268
rect -312 -268 -233 -250
rect -201 -250 -29 -248
rect -201 -266 -122 -250
rect -115 -252 -85 -250
rect -226 -268 -122 -266
rect -494 -288 -465 -278
rect -450 -288 -420 -274
rect -376 -288 -334 -274
rect -312 -278 -122 -268
rect -57 -270 -51 -250
rect -327 -288 -297 -278
rect -296 -288 -138 -278
rect -134 -288 -104 -278
rect -100 -288 -70 -274
rect -42 -288 -29 -250
rect 43 -236 72 -220
rect 86 -236 115 -220
rect 130 -230 160 -214
rect 188 -236 194 -188
rect 197 -194 216 -188
rect 231 -194 261 -186
rect 197 -202 261 -194
rect 197 -218 277 -202
rect 293 -209 355 -178
rect 371 -209 433 -178
rect 502 -180 551 -155
rect 596 -164 622 -154
rect 566 -180 622 -164
rect 465 -194 495 -186
rect 502 -188 612 -180
rect 465 -202 510 -194
rect 197 -220 216 -218
rect 231 -220 277 -218
rect 197 -236 277 -220
rect 304 -222 339 -209
rect 380 -212 417 -209
rect 380 -214 422 -212
rect 309 -225 339 -222
rect 318 -229 325 -225
rect 325 -230 326 -229
rect 284 -236 294 -230
rect 43 -244 78 -236
rect 43 -270 44 -244
rect 51 -270 78 -244
rect -14 -288 16 -274
rect 43 -278 78 -270
rect 80 -244 121 -236
rect 80 -270 95 -244
rect 102 -270 121 -244
rect 185 -248 216 -236
rect 231 -248 334 -236
rect 346 -246 372 -220
rect 387 -225 417 -214
rect 449 -218 511 -202
rect 449 -220 495 -218
rect 449 -236 511 -220
rect 523 -236 529 -188
rect 532 -196 612 -188
rect 532 -198 551 -196
rect 566 -198 600 -196
rect 532 -214 612 -198
rect 532 -236 551 -214
rect 566 -230 596 -214
rect 624 -220 630 -146
rect 633 -220 652 -76
rect 667 -220 673 -76
rect 682 -146 695 -76
rect 747 -80 769 -76
rect 740 -92 757 -88
rect 761 -90 769 -88
rect 759 -92 769 -90
rect 740 -102 769 -92
rect 822 -102 838 -88
rect 876 -92 882 -90
rect 889 -92 997 -76
rect 1004 -92 1010 -90
rect 1018 -92 1033 -76
rect 1099 -82 1118 -79
rect 740 -104 838 -102
rect 865 -104 1033 -92
rect 1048 -102 1064 -88
rect 1099 -101 1121 -82
rect 1131 -88 1147 -87
rect 1130 -90 1147 -88
rect 1131 -95 1147 -90
rect 1121 -102 1127 -101
rect 1130 -102 1159 -95
rect 1048 -103 1159 -102
rect 1048 -104 1165 -103
rect 724 -112 775 -104
rect 822 -112 856 -104
rect 724 -124 749 -112
rect 756 -124 775 -112
rect 829 -114 856 -112
rect 865 -114 1086 -104
rect 1121 -107 1127 -104
rect 829 -118 1086 -114
rect 724 -132 775 -124
rect 822 -132 1086 -118
rect 1130 -112 1165 -104
rect 676 -180 695 -146
rect 740 -140 769 -132
rect 740 -146 757 -140
rect 740 -148 774 -146
rect 822 -148 838 -132
rect 839 -142 1047 -132
rect 1048 -142 1064 -132
rect 1112 -136 1127 -121
rect 1130 -124 1131 -112
rect 1138 -124 1165 -112
rect 1130 -132 1165 -124
rect 1130 -133 1159 -132
rect 850 -146 1064 -142
rect 865 -148 1064 -146
rect 1099 -146 1112 -136
rect 1130 -146 1147 -133
rect 1099 -148 1147 -146
rect 741 -152 774 -148
rect 737 -154 774 -152
rect 737 -155 804 -154
rect 737 -160 768 -155
rect 774 -160 804 -155
rect 737 -164 804 -160
rect 710 -167 804 -164
rect 710 -174 759 -167
rect 710 -180 740 -174
rect 759 -179 764 -174
rect 676 -196 756 -180
rect 768 -188 804 -167
rect 865 -172 1054 -148
rect 1099 -149 1146 -148
rect 1112 -154 1146 -149
rect 880 -175 1054 -172
rect 873 -178 1054 -175
rect 1082 -155 1146 -154
rect 676 -198 695 -196
rect 710 -198 744 -196
rect 676 -214 756 -198
rect 676 -220 695 -214
rect 392 -246 495 -236
rect 346 -248 495 -246
rect 516 -248 551 -236
rect 185 -250 347 -248
rect 197 -268 216 -250
rect 231 -252 261 -250
rect 80 -278 121 -270
rect 204 -274 216 -268
rect 268 -268 347 -250
rect 379 -250 551 -248
rect 379 -266 458 -250
rect 465 -252 495 -250
rect 354 -268 458 -266
rect 43 -288 72 -278
rect 86 -288 115 -278
rect 130 -288 160 -274
rect 204 -288 246 -274
rect 268 -278 458 -268
rect 523 -270 529 -250
rect 253 -288 283 -278
rect 284 -288 442 -278
rect 446 -288 476 -278
rect 480 -288 510 -274
rect 538 -288 551 -250
rect 623 -236 652 -220
rect 666 -236 695 -220
rect 710 -230 740 -214
rect 768 -236 774 -188
rect 777 -194 796 -188
rect 811 -194 841 -186
rect 777 -202 841 -194
rect 777 -218 857 -202
rect 873 -209 935 -178
rect 951 -209 1013 -178
rect 1082 -180 1131 -155
rect 1146 -180 1176 -162
rect 1045 -194 1075 -186
rect 1082 -188 1192 -180
rect 1045 -202 1090 -194
rect 777 -220 796 -218
rect 811 -220 857 -218
rect 777 -236 857 -220
rect 884 -222 919 -209
rect 960 -212 997 -209
rect 960 -214 1002 -212
rect 889 -225 919 -222
rect 898 -229 905 -225
rect 905 -230 906 -229
rect 864 -236 874 -230
rect 623 -244 658 -236
rect 623 -270 624 -244
rect 631 -270 658 -244
rect 566 -288 596 -274
rect 623 -278 658 -270
rect 660 -244 701 -236
rect 660 -270 675 -244
rect 682 -270 701 -244
rect 765 -248 796 -236
rect 811 -248 914 -236
rect 926 -246 952 -220
rect 967 -225 997 -214
rect 1029 -218 1091 -202
rect 1029 -220 1075 -218
rect 1029 -236 1091 -220
rect 1103 -236 1109 -188
rect 1112 -196 1192 -188
rect 1112 -198 1131 -196
rect 1146 -198 1180 -196
rect 1112 -213 1192 -198
rect 1112 -214 1198 -213
rect 1112 -236 1131 -214
rect 1146 -230 1176 -214
rect 1204 -220 1210 -146
rect 1213 -220 1232 -76
rect 1247 -220 1253 -76
rect 1262 -146 1275 -76
rect 1327 -80 1349 -76
rect 1320 -92 1337 -88
rect 1341 -90 1349 -88
rect 1339 -92 1349 -90
rect 1320 -102 1349 -92
rect 1402 -102 1418 -88
rect 1456 -92 1462 -90
rect 1469 -92 1577 -76
rect 1584 -92 1590 -90
rect 1598 -92 1613 -76
rect 1679 -82 1698 -79
rect 1320 -104 1418 -102
rect 1445 -104 1613 -92
rect 1628 -102 1644 -88
rect 1679 -101 1701 -82
rect 1711 -88 1727 -87
rect 1710 -90 1727 -88
rect 1711 -95 1727 -90
rect 1701 -102 1707 -101
rect 1710 -102 1739 -95
rect 1628 -103 1739 -102
rect 1628 -104 1745 -103
rect 1304 -112 1355 -104
rect 1402 -112 1436 -104
rect 1304 -124 1329 -112
rect 1336 -124 1355 -112
rect 1409 -114 1436 -112
rect 1445 -114 1666 -104
rect 1701 -107 1707 -104
rect 1409 -118 1666 -114
rect 1304 -132 1355 -124
rect 1402 -132 1666 -118
rect 1710 -112 1745 -104
rect 1256 -180 1275 -146
rect 1320 -140 1349 -132
rect 1320 -146 1337 -140
rect 1320 -148 1354 -146
rect 1402 -148 1418 -132
rect 1419 -142 1627 -132
rect 1628 -142 1644 -132
rect 1692 -136 1707 -121
rect 1710 -124 1711 -112
rect 1718 -124 1745 -112
rect 1710 -132 1745 -124
rect 1710 -133 1739 -132
rect 1430 -146 1644 -142
rect 1445 -148 1644 -146
rect 1679 -146 1692 -136
rect 1710 -146 1727 -133
rect 1679 -148 1727 -146
rect 1321 -152 1354 -148
rect 1317 -154 1354 -152
rect 1317 -155 1384 -154
rect 1317 -160 1348 -155
rect 1354 -160 1384 -155
rect 1317 -164 1384 -160
rect 1290 -167 1384 -164
rect 1290 -174 1339 -167
rect 1290 -180 1320 -174
rect 1339 -179 1344 -174
rect 1256 -196 1336 -180
rect 1348 -188 1384 -167
rect 1445 -172 1634 -148
rect 1679 -149 1726 -148
rect 1692 -154 1726 -149
rect 1766 -154 1782 -152
rect 1460 -175 1634 -172
rect 1453 -178 1634 -175
rect 1662 -155 1726 -154
rect 1256 -198 1275 -196
rect 1290 -198 1324 -196
rect 1256 -214 1336 -198
rect 1256 -220 1275 -214
rect 972 -246 1075 -236
rect 926 -248 1075 -246
rect 1096 -248 1131 -236
rect 765 -250 927 -248
rect 777 -268 796 -250
rect 811 -252 841 -250
rect 660 -278 701 -270
rect 784 -274 796 -268
rect 848 -268 927 -250
rect 959 -250 1131 -248
rect 959 -266 1038 -250
rect 1045 -252 1075 -250
rect 934 -268 1038 -266
rect 623 -288 652 -278
rect 666 -288 695 -278
rect 710 -288 740 -274
rect 784 -288 826 -274
rect 848 -278 1038 -268
rect 1103 -270 1109 -250
rect 833 -288 863 -278
rect 864 -288 1022 -278
rect 1026 -288 1056 -278
rect 1060 -288 1090 -274
rect 1118 -288 1131 -250
rect 1203 -236 1232 -220
rect 1246 -236 1275 -220
rect 1290 -230 1320 -214
rect 1348 -236 1354 -188
rect 1357 -194 1376 -188
rect 1391 -194 1421 -186
rect 1357 -202 1421 -194
rect 1357 -218 1437 -202
rect 1453 -209 1515 -178
rect 1531 -209 1593 -178
rect 1662 -180 1711 -155
rect 1756 -164 1782 -154
rect 1726 -180 1782 -164
rect 1625 -194 1655 -186
rect 1662 -188 1772 -180
rect 1625 -202 1670 -194
rect 1357 -220 1376 -218
rect 1391 -220 1437 -218
rect 1357 -236 1437 -220
rect 1464 -222 1499 -209
rect 1540 -212 1577 -209
rect 1540 -214 1582 -212
rect 1469 -225 1499 -222
rect 1478 -229 1485 -225
rect 1485 -230 1486 -229
rect 1444 -236 1454 -230
rect 1203 -244 1238 -236
rect 1203 -270 1204 -244
rect 1211 -270 1238 -244
rect 1146 -288 1176 -274
rect 1203 -278 1238 -270
rect 1240 -244 1281 -236
rect 1240 -270 1255 -244
rect 1262 -270 1281 -244
rect 1345 -248 1376 -236
rect 1391 -248 1494 -236
rect 1506 -246 1532 -220
rect 1547 -225 1577 -214
rect 1609 -218 1671 -202
rect 1609 -220 1655 -218
rect 1609 -236 1671 -220
rect 1683 -236 1689 -188
rect 1692 -196 1772 -188
rect 1692 -198 1711 -196
rect 1726 -198 1760 -196
rect 1692 -214 1772 -198
rect 1692 -236 1711 -214
rect 1726 -230 1756 -214
rect 1784 -220 1790 -146
rect 1793 -220 1812 -76
rect 1827 -220 1833 -76
rect 1842 -146 1855 -76
rect 1907 -80 1929 -76
rect 1900 -92 1917 -88
rect 1921 -90 1929 -88
rect 1919 -92 1929 -90
rect 1900 -102 1929 -92
rect 1982 -102 1998 -88
rect 2036 -92 2042 -90
rect 2049 -92 2157 -76
rect 2164 -92 2170 -90
rect 2178 -92 2193 -76
rect 2259 -82 2278 -79
rect 1900 -104 1998 -102
rect 2025 -104 2193 -92
rect 2208 -102 2224 -88
rect 2259 -101 2281 -82
rect 2291 -88 2307 -87
rect 2290 -90 2307 -88
rect 2291 -95 2307 -90
rect 2281 -102 2287 -101
rect 2290 -102 2319 -95
rect 2208 -103 2319 -102
rect 2208 -104 2325 -103
rect 1884 -112 1935 -104
rect 1982 -112 2016 -104
rect 1884 -124 1909 -112
rect 1916 -124 1935 -112
rect 1989 -114 2016 -112
rect 2025 -114 2246 -104
rect 2281 -107 2287 -104
rect 1989 -118 2246 -114
rect 1884 -132 1935 -124
rect 1982 -132 2246 -118
rect 2290 -112 2325 -104
rect 1836 -180 1855 -146
rect 1900 -140 1929 -132
rect 1900 -146 1917 -140
rect 1900 -148 1934 -146
rect 1982 -148 1998 -132
rect 1999 -142 2207 -132
rect 2208 -142 2224 -132
rect 2272 -136 2287 -121
rect 2290 -124 2291 -112
rect 2298 -124 2325 -112
rect 2290 -132 2325 -124
rect 2290 -133 2319 -132
rect 2010 -146 2224 -142
rect 2025 -148 2224 -146
rect 2259 -146 2272 -136
rect 2290 -146 2307 -133
rect 2259 -148 2307 -146
rect 1901 -152 1934 -148
rect 1897 -154 1934 -152
rect 1897 -155 1964 -154
rect 1897 -160 1928 -155
rect 1934 -160 1964 -155
rect 1897 -164 1964 -160
rect 1870 -167 1964 -164
rect 1870 -174 1919 -167
rect 1870 -180 1900 -174
rect 1919 -179 1924 -174
rect 1836 -196 1916 -180
rect 1928 -188 1964 -167
rect 2025 -172 2214 -148
rect 2259 -149 2306 -148
rect 2272 -154 2306 -149
rect 2040 -175 2214 -172
rect 2033 -178 2214 -175
rect 2242 -155 2306 -154
rect 1836 -198 1855 -196
rect 1870 -198 1904 -196
rect 1836 -214 1916 -198
rect 1836 -220 1855 -214
rect 1552 -246 1655 -236
rect 1506 -248 1655 -246
rect 1676 -248 1711 -236
rect 1345 -250 1507 -248
rect 1357 -268 1376 -250
rect 1391 -252 1421 -250
rect 1240 -278 1281 -270
rect 1364 -274 1376 -268
rect 1428 -268 1507 -250
rect 1539 -250 1711 -248
rect 1539 -266 1618 -250
rect 1625 -252 1655 -250
rect 1514 -268 1618 -266
rect 1203 -288 1232 -278
rect 1246 -288 1275 -278
rect 1290 -288 1320 -274
rect 1364 -288 1406 -274
rect 1428 -278 1618 -268
rect 1683 -270 1689 -250
rect 1413 -288 1443 -278
rect 1444 -288 1602 -278
rect 1606 -288 1636 -278
rect 1640 -288 1670 -274
rect 1698 -288 1711 -250
rect 1783 -236 1812 -220
rect 1826 -236 1855 -220
rect 1870 -230 1900 -214
rect 1928 -236 1934 -188
rect 1937 -194 1956 -188
rect 1971 -194 2001 -186
rect 1937 -202 2001 -194
rect 1937 -218 2017 -202
rect 2033 -209 2095 -178
rect 2111 -209 2173 -178
rect 2242 -180 2291 -155
rect 2306 -180 2336 -162
rect 2205 -194 2235 -186
rect 2242 -188 2352 -180
rect 2205 -202 2250 -194
rect 1937 -220 1956 -218
rect 1971 -220 2017 -218
rect 1937 -236 2017 -220
rect 2044 -222 2079 -209
rect 2120 -212 2157 -209
rect 2120 -214 2162 -212
rect 2049 -225 2079 -222
rect 2058 -229 2065 -225
rect 2065 -230 2066 -229
rect 2024 -236 2034 -230
rect 1783 -244 1818 -236
rect 1783 -270 1784 -244
rect 1791 -270 1818 -244
rect 1726 -288 1756 -274
rect 1783 -278 1818 -270
rect 1820 -244 1861 -236
rect 1820 -270 1835 -244
rect 1842 -270 1861 -244
rect 1925 -248 1956 -236
rect 1971 -248 2074 -236
rect 2086 -246 2112 -220
rect 2127 -225 2157 -214
rect 2189 -218 2251 -202
rect 2189 -220 2235 -218
rect 2189 -236 2251 -220
rect 2263 -236 2269 -188
rect 2272 -196 2352 -188
rect 2272 -198 2291 -196
rect 2306 -198 2340 -196
rect 2272 -213 2352 -198
rect 2272 -214 2358 -213
rect 2272 -236 2291 -214
rect 2306 -230 2336 -214
rect 2364 -220 2370 -146
rect 2373 -220 2392 -76
rect 2407 -220 2413 -76
rect 2422 -146 2435 -76
rect 2487 -80 2509 -76
rect 2480 -92 2497 -88
rect 2501 -90 2509 -88
rect 2499 -92 2509 -90
rect 2480 -102 2509 -92
rect 2562 -102 2578 -88
rect 2616 -92 2622 -90
rect 2629 -92 2737 -76
rect 2744 -92 2750 -90
rect 2758 -92 2773 -76
rect 2839 -82 2858 -79
rect 2480 -104 2578 -102
rect 2605 -104 2773 -92
rect 2788 -102 2804 -88
rect 2839 -101 2861 -82
rect 2871 -88 2887 -87
rect 2870 -90 2887 -88
rect 2871 -95 2887 -90
rect 2861 -102 2867 -101
rect 2870 -102 2899 -95
rect 2788 -103 2899 -102
rect 2788 -104 2905 -103
rect 2464 -112 2515 -104
rect 2562 -112 2596 -104
rect 2464 -124 2489 -112
rect 2496 -124 2515 -112
rect 2569 -114 2596 -112
rect 2605 -114 2826 -104
rect 2861 -107 2867 -104
rect 2569 -118 2826 -114
rect 2464 -132 2515 -124
rect 2562 -132 2826 -118
rect 2870 -112 2905 -104
rect 2416 -180 2435 -146
rect 2480 -140 2509 -132
rect 2480 -146 2497 -140
rect 2480 -148 2514 -146
rect 2562 -148 2578 -132
rect 2579 -142 2787 -132
rect 2788 -142 2804 -132
rect 2852 -136 2867 -121
rect 2870 -124 2871 -112
rect 2878 -124 2905 -112
rect 2870 -132 2905 -124
rect 2870 -133 2899 -132
rect 2590 -146 2804 -142
rect 2605 -148 2804 -146
rect 2839 -146 2852 -136
rect 2870 -146 2887 -133
rect 2839 -148 2887 -146
rect 2481 -152 2514 -148
rect 2477 -154 2514 -152
rect 2477 -155 2544 -154
rect 2477 -160 2508 -155
rect 2514 -160 2544 -155
rect 2477 -164 2544 -160
rect 2450 -167 2544 -164
rect 2450 -174 2499 -167
rect 2450 -180 2480 -174
rect 2499 -179 2504 -174
rect 2416 -196 2496 -180
rect 2508 -188 2544 -167
rect 2605 -172 2794 -148
rect 2839 -149 2886 -148
rect 2852 -154 2886 -149
rect 2926 -154 2942 -152
rect 2620 -175 2794 -172
rect 2613 -178 2794 -175
rect 2822 -155 2886 -154
rect 2416 -198 2435 -196
rect 2450 -198 2484 -196
rect 2416 -214 2496 -198
rect 2416 -220 2435 -214
rect 2132 -246 2235 -236
rect 2086 -248 2235 -246
rect 2256 -248 2291 -236
rect 1925 -250 2087 -248
rect 1937 -268 1956 -250
rect 1971 -252 2001 -250
rect 1820 -278 1861 -270
rect 1944 -274 1956 -268
rect 2008 -266 2087 -250
rect 2119 -250 2291 -248
rect 2119 -266 2198 -250
rect 2205 -252 2235 -250
rect 1783 -288 1812 -278
rect 1826 -288 1855 -278
rect 1870 -288 1900 -274
rect 1944 -288 1986 -274
rect 2008 -278 2198 -266
rect 2263 -270 2269 -250
rect 1993 -288 2023 -278
rect 2024 -288 2182 -278
rect 2186 -288 2216 -278
rect 2220 -288 2250 -274
rect 2278 -288 2291 -250
rect 2363 -236 2392 -220
rect 2406 -236 2435 -220
rect 2450 -230 2480 -214
rect 2508 -236 2514 -188
rect 2517 -194 2536 -188
rect 2551 -194 2581 -186
rect 2517 -202 2581 -194
rect 2517 -218 2597 -202
rect 2613 -209 2675 -178
rect 2691 -209 2753 -178
rect 2822 -180 2871 -155
rect 2916 -164 2942 -154
rect 2886 -180 2942 -164
rect 2785 -194 2815 -186
rect 2822 -188 2932 -180
rect 2785 -202 2830 -194
rect 2517 -220 2536 -218
rect 2551 -220 2597 -218
rect 2517 -236 2597 -220
rect 2624 -222 2659 -209
rect 2700 -212 2737 -209
rect 2700 -214 2742 -212
rect 2629 -225 2659 -222
rect 2638 -229 2645 -225
rect 2645 -230 2646 -229
rect 2604 -236 2614 -230
rect 2363 -244 2398 -236
rect 2363 -270 2364 -244
rect 2371 -270 2398 -244
rect 2306 -288 2336 -274
rect 2363 -278 2398 -270
rect 2400 -244 2441 -236
rect 2400 -270 2415 -244
rect 2422 -270 2441 -244
rect 2505 -248 2536 -236
rect 2551 -248 2654 -236
rect 2666 -246 2692 -220
rect 2707 -225 2737 -214
rect 2769 -218 2831 -202
rect 2769 -220 2815 -218
rect 2769 -236 2831 -220
rect 2843 -236 2849 -188
rect 2852 -196 2932 -188
rect 2852 -198 2871 -196
rect 2886 -198 2920 -196
rect 2852 -214 2932 -198
rect 2852 -236 2871 -214
rect 2886 -230 2916 -214
rect 2944 -220 2950 -146
rect 2953 -220 2972 -76
rect 2987 -220 2993 -76
rect 3002 -146 3015 -76
rect 3067 -80 3089 -76
rect 3060 -92 3077 -88
rect 3081 -90 3089 -88
rect 3079 -92 3089 -90
rect 3060 -102 3089 -92
rect 3142 -102 3158 -88
rect 3196 -92 3202 -90
rect 3209 -92 3317 -76
rect 3324 -92 3330 -90
rect 3338 -92 3353 -76
rect 3419 -82 3438 -79
rect 3060 -104 3158 -102
rect 3185 -104 3353 -92
rect 3368 -102 3384 -88
rect 3419 -101 3441 -82
rect 3451 -88 3467 -87
rect 3450 -90 3467 -88
rect 3451 -95 3467 -90
rect 3441 -102 3447 -101
rect 3450 -102 3479 -95
rect 3368 -103 3479 -102
rect 3368 -104 3485 -103
rect 3044 -112 3095 -104
rect 3142 -112 3176 -104
rect 3044 -124 3069 -112
rect 3076 -124 3095 -112
rect 3149 -114 3176 -112
rect 3185 -114 3406 -104
rect 3441 -107 3447 -104
rect 3149 -118 3406 -114
rect 3044 -132 3095 -124
rect 3142 -132 3406 -118
rect 3450 -112 3485 -104
rect 2996 -180 3015 -146
rect 3060 -140 3089 -132
rect 3060 -146 3077 -140
rect 3060 -148 3094 -146
rect 3142 -148 3158 -132
rect 3159 -142 3367 -132
rect 3368 -142 3384 -132
rect 3432 -136 3447 -121
rect 3450 -124 3451 -112
rect 3458 -124 3485 -112
rect 3450 -132 3485 -124
rect 3450 -133 3479 -132
rect 3170 -146 3384 -142
rect 3185 -148 3384 -146
rect 3419 -146 3432 -136
rect 3450 -146 3467 -133
rect 3419 -148 3467 -146
rect 3061 -152 3094 -148
rect 3057 -154 3094 -152
rect 3057 -155 3124 -154
rect 3057 -160 3088 -155
rect 3094 -160 3124 -155
rect 3057 -164 3124 -160
rect 3030 -167 3124 -164
rect 3030 -174 3079 -167
rect 3030 -180 3060 -174
rect 3079 -179 3084 -174
rect 2996 -196 3076 -180
rect 3088 -188 3124 -167
rect 3185 -172 3374 -148
rect 3419 -149 3466 -148
rect 3432 -154 3466 -149
rect 3200 -175 3374 -172
rect 3193 -178 3374 -175
rect 3402 -155 3466 -154
rect 2996 -198 3015 -196
rect 3030 -198 3064 -196
rect 2996 -214 3076 -198
rect 2996 -220 3015 -214
rect 2712 -246 2815 -236
rect 2666 -248 2815 -246
rect 2836 -248 2871 -236
rect 2505 -250 2667 -248
rect 2517 -268 2536 -250
rect 2551 -252 2581 -250
rect 2400 -278 2441 -270
rect 2524 -274 2536 -268
rect 2588 -266 2667 -250
rect 2699 -250 2871 -248
rect 2699 -266 2778 -250
rect 2785 -252 2815 -250
rect 2363 -288 2392 -278
rect 2406 -288 2435 -278
rect 2450 -288 2480 -274
rect 2524 -288 2566 -274
rect 2588 -278 2778 -266
rect 2843 -270 2849 -250
rect 2573 -288 2603 -278
rect 2604 -288 2762 -278
rect 2766 -288 2796 -278
rect 2800 -288 2830 -274
rect 2858 -288 2871 -250
rect 2943 -236 2972 -220
rect 2986 -236 3015 -220
rect 3030 -230 3060 -214
rect 3088 -236 3094 -188
rect 3097 -194 3116 -188
rect 3131 -194 3161 -186
rect 3097 -202 3161 -194
rect 3097 -218 3177 -202
rect 3193 -209 3255 -178
rect 3271 -209 3333 -178
rect 3402 -180 3451 -155
rect 3466 -180 3496 -162
rect 3365 -194 3395 -186
rect 3402 -188 3512 -180
rect 3365 -202 3410 -194
rect 3097 -220 3116 -218
rect 3131 -220 3177 -218
rect 3097 -236 3177 -220
rect 3204 -222 3239 -209
rect 3280 -212 3317 -209
rect 3280 -214 3322 -212
rect 3209 -225 3239 -222
rect 3218 -229 3225 -225
rect 3225 -230 3226 -229
rect 3184 -236 3194 -230
rect 2943 -244 2978 -236
rect 2943 -270 2944 -244
rect 2951 -270 2978 -244
rect 2886 -288 2916 -274
rect 2943 -278 2978 -270
rect 2980 -244 3021 -236
rect 2980 -270 2995 -244
rect 3002 -270 3021 -244
rect 3085 -248 3116 -236
rect 3131 -248 3234 -236
rect 3246 -246 3272 -220
rect 3287 -225 3317 -214
rect 3349 -218 3411 -202
rect 3349 -220 3395 -218
rect 3349 -236 3411 -220
rect 3423 -236 3429 -188
rect 3432 -196 3512 -188
rect 3432 -198 3451 -196
rect 3466 -198 3500 -196
rect 3432 -213 3512 -198
rect 3432 -214 3518 -213
rect 3432 -236 3451 -214
rect 3466 -230 3496 -214
rect 3524 -220 3530 -146
rect 3533 -220 3552 -76
rect 3567 -220 3573 -76
rect 3582 -146 3595 -76
rect 3647 -80 3669 -76
rect 3640 -92 3657 -88
rect 3661 -90 3669 -88
rect 3659 -92 3669 -90
rect 3640 -102 3669 -92
rect 3722 -102 3738 -88
rect 3776 -92 3782 -90
rect 3789 -92 3897 -76
rect 3904 -92 3910 -90
rect 3918 -92 3933 -76
rect 3999 -82 4018 -79
rect 3640 -104 3738 -102
rect 3765 -104 3933 -92
rect 3948 -102 3964 -88
rect 3999 -101 4021 -82
rect 4031 -88 4047 -87
rect 4030 -90 4047 -88
rect 4031 -95 4047 -90
rect 4021 -102 4027 -101
rect 4030 -102 4059 -95
rect 3948 -103 4059 -102
rect 3948 -104 4065 -103
rect 3624 -112 3675 -104
rect 3722 -112 3756 -104
rect 3624 -124 3649 -112
rect 3656 -124 3675 -112
rect 3729 -114 3756 -112
rect 3765 -114 3986 -104
rect 4021 -107 4027 -104
rect 3729 -118 3986 -114
rect 3624 -132 3675 -124
rect 3722 -132 3986 -118
rect 4030 -112 4065 -104
rect 3576 -180 3595 -146
rect 3640 -140 3669 -132
rect 3640 -146 3657 -140
rect 3640 -148 3674 -146
rect 3722 -148 3738 -132
rect 3739 -142 3947 -132
rect 3948 -142 3964 -132
rect 4012 -136 4027 -121
rect 4030 -124 4031 -112
rect 4038 -124 4065 -112
rect 4030 -132 4065 -124
rect 4030 -133 4059 -132
rect 3750 -146 3964 -142
rect 3765 -148 3964 -146
rect 3999 -146 4012 -136
rect 4030 -146 4047 -133
rect 3999 -148 4047 -146
rect 3641 -152 3674 -148
rect 3637 -154 3674 -152
rect 3637 -155 3704 -154
rect 3637 -160 3668 -155
rect 3674 -160 3704 -155
rect 3637 -164 3704 -160
rect 3610 -167 3704 -164
rect 3610 -174 3659 -167
rect 3610 -180 3640 -174
rect 3659 -179 3664 -174
rect 3576 -196 3656 -180
rect 3668 -188 3704 -167
rect 3765 -172 3954 -148
rect 3999 -149 4046 -148
rect 4012 -154 4046 -149
rect 4086 -154 4102 -152
rect 3780 -175 3954 -172
rect 3773 -178 3954 -175
rect 3982 -155 4046 -154
rect 3576 -198 3595 -196
rect 3610 -198 3644 -196
rect 3576 -214 3656 -198
rect 3576 -220 3595 -214
rect 3292 -246 3395 -236
rect 3246 -248 3395 -246
rect 3416 -248 3451 -236
rect 3085 -250 3247 -248
rect 3097 -268 3116 -250
rect 3131 -252 3161 -250
rect 2980 -278 3021 -270
rect 3104 -274 3116 -268
rect 3168 -266 3247 -250
rect 3279 -250 3451 -248
rect 3279 -266 3358 -250
rect 3365 -252 3395 -250
rect 2943 -288 2972 -278
rect 2986 -288 3015 -278
rect 3030 -288 3060 -274
rect 3104 -288 3146 -274
rect 3168 -278 3358 -266
rect 3423 -270 3429 -250
rect 3153 -288 3183 -278
rect 3184 -288 3342 -278
rect 3346 -288 3376 -278
rect 3380 -288 3410 -274
rect 3438 -288 3451 -250
rect 3523 -236 3552 -220
rect 3566 -236 3595 -220
rect 3610 -230 3640 -214
rect 3668 -236 3674 -188
rect 3677 -194 3696 -188
rect 3711 -194 3741 -186
rect 3677 -202 3741 -194
rect 3677 -218 3757 -202
rect 3773 -209 3835 -178
rect 3851 -209 3913 -178
rect 3982 -180 4031 -155
rect 4076 -164 4102 -154
rect 4046 -180 4102 -164
rect 3945 -194 3975 -186
rect 3982 -188 4092 -180
rect 3945 -202 3990 -194
rect 3677 -220 3696 -218
rect 3711 -220 3757 -218
rect 3677 -236 3757 -220
rect 3784 -222 3819 -209
rect 3860 -212 3897 -209
rect 3860 -214 3902 -212
rect 3789 -225 3819 -222
rect 3798 -229 3805 -225
rect 3805 -230 3806 -229
rect 3764 -236 3774 -230
rect 3523 -244 3558 -236
rect 3523 -270 3524 -244
rect 3531 -270 3558 -244
rect 3466 -288 3496 -274
rect 3523 -278 3558 -270
rect 3560 -244 3601 -236
rect 3560 -270 3575 -244
rect 3582 -270 3601 -244
rect 3665 -248 3696 -236
rect 3711 -248 3814 -236
rect 3826 -246 3852 -220
rect 3867 -225 3897 -214
rect 3929 -218 3991 -202
rect 3929 -220 3975 -218
rect 3929 -236 3991 -220
rect 4003 -236 4009 -188
rect 4012 -196 4092 -188
rect 4012 -198 4031 -196
rect 4046 -198 4080 -196
rect 4012 -214 4092 -198
rect 4012 -236 4031 -214
rect 4046 -230 4076 -214
rect 4104 -220 4110 -146
rect 4113 -220 4132 -76
rect 4147 -220 4153 -76
rect 4162 -146 4175 -76
rect 4227 -80 4249 -76
rect 4220 -92 4237 -88
rect 4241 -90 4249 -88
rect 4239 -92 4249 -90
rect 4220 -102 4249 -92
rect 4302 -102 4318 -88
rect 4356 -92 4362 -90
rect 4369 -92 4477 -76
rect 4484 -92 4490 -90
rect 4498 -92 4513 -76
rect 4579 -82 4598 -79
rect 4220 -104 4318 -102
rect 4345 -104 4513 -92
rect 4528 -102 4544 -88
rect 4579 -101 4601 -82
rect 4611 -88 4627 -87
rect 4610 -90 4627 -88
rect 4611 -95 4627 -90
rect 4601 -102 4607 -101
rect 4610 -102 4639 -95
rect 4528 -103 4639 -102
rect 4528 -104 4645 -103
rect 4204 -112 4255 -104
rect 4302 -112 4336 -104
rect 4204 -124 4229 -112
rect 4236 -124 4255 -112
rect 4309 -114 4336 -112
rect 4345 -114 4566 -104
rect 4601 -107 4607 -104
rect 4309 -118 4566 -114
rect 4204 -132 4255 -124
rect 4302 -132 4566 -118
rect 4610 -112 4645 -104
rect 4156 -180 4175 -146
rect 4220 -140 4249 -132
rect 4220 -146 4237 -140
rect 4220 -148 4254 -146
rect 4302 -148 4318 -132
rect 4319 -142 4527 -132
rect 4528 -142 4544 -132
rect 4592 -136 4607 -121
rect 4610 -124 4611 -112
rect 4618 -124 4645 -112
rect 4610 -132 4645 -124
rect 4610 -133 4639 -132
rect 4330 -146 4544 -142
rect 4345 -148 4544 -146
rect 4579 -146 4592 -136
rect 4610 -146 4627 -133
rect 4579 -148 4627 -146
rect 4221 -152 4254 -148
rect 4217 -154 4254 -152
rect 4217 -155 4284 -154
rect 4217 -160 4248 -155
rect 4254 -160 4284 -155
rect 4217 -164 4284 -160
rect 4190 -167 4284 -164
rect 4190 -174 4239 -167
rect 4190 -180 4220 -174
rect 4239 -179 4244 -174
rect 4156 -196 4236 -180
rect 4248 -188 4284 -167
rect 4345 -172 4534 -148
rect 4579 -149 4626 -148
rect 4592 -154 4626 -149
rect 4360 -175 4534 -172
rect 4353 -178 4534 -175
rect 4562 -155 4626 -154
rect 4156 -198 4175 -196
rect 4190 -198 4224 -196
rect 4156 -214 4236 -198
rect 4156 -220 4175 -214
rect 3872 -246 3975 -236
rect 3826 -248 3975 -246
rect 3996 -248 4031 -236
rect 3665 -250 3827 -248
rect 3677 -268 3696 -250
rect 3711 -252 3741 -250
rect 3560 -278 3601 -270
rect 3684 -274 3696 -268
rect 3748 -266 3827 -250
rect 3859 -250 4031 -248
rect 3859 -266 3938 -250
rect 3945 -252 3975 -250
rect 3523 -288 3552 -278
rect 3566 -288 3595 -278
rect 3610 -288 3640 -274
rect 3684 -288 3726 -274
rect 3748 -278 3938 -266
rect 4003 -270 4009 -250
rect 3733 -288 3763 -278
rect 3764 -288 3922 -278
rect 3926 -288 3956 -278
rect 3960 -288 3990 -274
rect 4018 -288 4031 -250
rect 4103 -236 4132 -220
rect 4146 -236 4175 -220
rect 4190 -230 4220 -214
rect 4248 -236 4254 -188
rect 4257 -194 4276 -188
rect 4291 -194 4321 -186
rect 4257 -202 4321 -194
rect 4257 -218 4337 -202
rect 4353 -209 4415 -178
rect 4431 -209 4493 -178
rect 4562 -180 4611 -155
rect 4626 -180 4656 -162
rect 4525 -194 4555 -186
rect 4562 -188 4672 -180
rect 4525 -202 4570 -194
rect 4257 -220 4276 -218
rect 4291 -220 4337 -218
rect 4257 -236 4337 -220
rect 4364 -222 4399 -209
rect 4440 -212 4477 -209
rect 4440 -214 4482 -212
rect 4369 -225 4399 -222
rect 4378 -229 4385 -225
rect 4385 -230 4386 -229
rect 4344 -236 4354 -230
rect 4103 -244 4138 -236
rect 4103 -270 4104 -244
rect 4111 -270 4138 -244
rect 4046 -288 4076 -274
rect 4103 -278 4138 -270
rect 4140 -244 4181 -236
rect 4140 -270 4155 -244
rect 4162 -270 4181 -244
rect 4245 -248 4276 -236
rect 4291 -248 4394 -236
rect 4406 -246 4432 -220
rect 4447 -225 4477 -214
rect 4509 -218 4571 -202
rect 4509 -220 4555 -218
rect 4509 -236 4571 -220
rect 4583 -236 4589 -188
rect 4592 -196 4672 -188
rect 4592 -198 4611 -196
rect 4626 -198 4660 -196
rect 4592 -213 4672 -198
rect 4592 -214 4678 -213
rect 4592 -236 4611 -214
rect 4626 -230 4656 -214
rect 4684 -220 4690 -146
rect 4693 -220 4712 -76
rect 4727 -220 4733 -76
rect 4742 -146 4755 -76
rect 4807 -80 4829 -76
rect 4800 -92 4817 -88
rect 4821 -90 4829 -88
rect 4819 -92 4829 -90
rect 4800 -102 4829 -92
rect 4882 -102 4898 -88
rect 4936 -92 4942 -90
rect 4949 -92 5057 -76
rect 5064 -92 5070 -90
rect 5078 -92 5093 -76
rect 5159 -82 5178 -79
rect 4800 -104 4898 -102
rect 4925 -104 5093 -92
rect 5108 -102 5124 -88
rect 5159 -101 5181 -82
rect 5191 -88 5207 -87
rect 5190 -90 5207 -88
rect 5191 -95 5207 -90
rect 5181 -102 5187 -101
rect 5190 -102 5219 -95
rect 5108 -103 5219 -102
rect 5108 -104 5225 -103
rect 4784 -112 4835 -104
rect 4882 -112 4916 -104
rect 4784 -124 4809 -112
rect 4816 -124 4835 -112
rect 4889 -114 4916 -112
rect 4925 -114 5146 -104
rect 5181 -107 5187 -104
rect 4889 -118 5146 -114
rect 4784 -132 4835 -124
rect 4882 -132 5146 -118
rect 5190 -112 5225 -104
rect 4736 -180 4755 -146
rect 4800 -140 4829 -132
rect 4800 -146 4817 -140
rect 4800 -148 4834 -146
rect 4882 -148 4898 -132
rect 4899 -142 5107 -132
rect 5108 -142 5124 -132
rect 5172 -136 5187 -121
rect 5190 -124 5191 -112
rect 5198 -124 5225 -112
rect 5190 -132 5225 -124
rect 5190 -133 5219 -132
rect 4910 -146 5124 -142
rect 4925 -148 5124 -146
rect 5159 -146 5172 -136
rect 5190 -146 5207 -133
rect 5159 -148 5207 -146
rect 4801 -152 4834 -148
rect 4797 -154 4834 -152
rect 4797 -155 4864 -154
rect 4797 -160 4828 -155
rect 4834 -160 4864 -155
rect 4797 -164 4864 -160
rect 4770 -167 4864 -164
rect 4770 -174 4819 -167
rect 4770 -180 4800 -174
rect 4819 -179 4824 -174
rect 4736 -196 4816 -180
rect 4828 -188 4864 -167
rect 4925 -172 5114 -148
rect 5159 -149 5206 -148
rect 5172 -154 5206 -149
rect 5246 -154 5262 -152
rect 4940 -175 5114 -172
rect 4933 -178 5114 -175
rect 5142 -155 5206 -154
rect 4736 -198 4755 -196
rect 4770 -198 4804 -196
rect 4736 -214 4816 -198
rect 4736 -220 4755 -214
rect 4452 -246 4555 -236
rect 4406 -248 4555 -246
rect 4576 -248 4611 -236
rect 4245 -250 4407 -248
rect 4257 -268 4276 -250
rect 4291 -252 4321 -250
rect 4140 -278 4181 -270
rect 4264 -274 4276 -268
rect 4328 -266 4407 -250
rect 4439 -250 4611 -248
rect 4439 -266 4518 -250
rect 4525 -252 4555 -250
rect 4103 -288 4132 -278
rect 4146 -288 4175 -278
rect 4190 -288 4220 -274
rect 4264 -288 4306 -274
rect 4328 -278 4518 -266
rect 4583 -270 4589 -250
rect 4313 -288 4343 -278
rect 4344 -288 4502 -278
rect 4506 -288 4536 -278
rect 4540 -288 4570 -274
rect 4598 -288 4611 -250
rect 4683 -236 4712 -220
rect 4726 -236 4755 -220
rect 4770 -230 4800 -214
rect 4828 -236 4834 -188
rect 4837 -194 4856 -188
rect 4871 -194 4901 -186
rect 4837 -202 4901 -194
rect 4837 -218 4917 -202
rect 4933 -209 4995 -178
rect 5011 -209 5073 -178
rect 5142 -180 5191 -155
rect 5236 -164 5262 -154
rect 5206 -180 5262 -164
rect 5105 -194 5135 -186
rect 5142 -188 5252 -180
rect 5105 -202 5150 -194
rect 4837 -220 4856 -218
rect 4871 -220 4917 -218
rect 4837 -236 4917 -220
rect 4944 -222 4979 -209
rect 5020 -212 5057 -209
rect 5020 -214 5062 -212
rect 4949 -225 4979 -222
rect 4958 -229 4965 -225
rect 4965 -230 4966 -229
rect 4924 -236 4934 -230
rect 4683 -244 4718 -236
rect 4683 -270 4684 -244
rect 4691 -270 4718 -244
rect 4626 -288 4656 -274
rect 4683 -278 4718 -270
rect 4720 -244 4761 -236
rect 4720 -270 4735 -244
rect 4742 -270 4761 -244
rect 4825 -248 4856 -236
rect 4871 -248 4974 -236
rect 4986 -246 5012 -220
rect 5027 -225 5057 -214
rect 5089 -218 5151 -202
rect 5089 -220 5135 -218
rect 5089 -236 5151 -220
rect 5163 -236 5169 -188
rect 5172 -196 5252 -188
rect 5172 -198 5191 -196
rect 5206 -198 5240 -196
rect 5172 -214 5252 -198
rect 5172 -236 5191 -214
rect 5206 -230 5236 -214
rect 5264 -220 5270 -146
rect 5273 -220 5292 -76
rect 5307 -220 5313 -76
rect 5322 -146 5335 -76
rect 5387 -80 5409 -76
rect 5380 -92 5397 -88
rect 5401 -90 5409 -88
rect 5399 -92 5409 -90
rect 5380 -102 5409 -92
rect 5462 -102 5478 -88
rect 5516 -92 5522 -90
rect 5529 -92 5637 -76
rect 5644 -92 5650 -90
rect 5658 -92 5673 -76
rect 5739 -82 5758 -79
rect 5380 -104 5478 -102
rect 5505 -104 5673 -92
rect 5688 -102 5704 -88
rect 5739 -101 5761 -82
rect 5771 -88 5787 -87
rect 5770 -90 5787 -88
rect 5771 -95 5787 -90
rect 5761 -102 5767 -101
rect 5770 -102 5799 -95
rect 5688 -103 5799 -102
rect 5688 -104 5805 -103
rect 5364 -112 5415 -104
rect 5462 -112 5496 -104
rect 5364 -124 5389 -112
rect 5396 -124 5415 -112
rect 5469 -114 5496 -112
rect 5505 -114 5726 -104
rect 5761 -107 5767 -104
rect 5469 -118 5726 -114
rect 5364 -132 5415 -124
rect 5462 -132 5726 -118
rect 5770 -112 5805 -104
rect 5316 -180 5335 -146
rect 5380 -140 5409 -132
rect 5380 -146 5397 -140
rect 5380 -148 5414 -146
rect 5462 -148 5478 -132
rect 5479 -142 5687 -132
rect 5688 -142 5704 -132
rect 5752 -136 5767 -121
rect 5770 -124 5771 -112
rect 5778 -124 5805 -112
rect 5770 -132 5805 -124
rect 5770 -133 5799 -132
rect 5490 -146 5704 -142
rect 5505 -148 5704 -146
rect 5739 -146 5752 -136
rect 5770 -146 5787 -133
rect 5739 -148 5787 -146
rect 5381 -152 5414 -148
rect 5377 -154 5414 -152
rect 5377 -155 5444 -154
rect 5377 -160 5408 -155
rect 5414 -160 5444 -155
rect 5377 -164 5444 -160
rect 5350 -167 5444 -164
rect 5350 -174 5399 -167
rect 5350 -180 5380 -174
rect 5399 -179 5404 -174
rect 5316 -196 5396 -180
rect 5408 -188 5444 -167
rect 5505 -172 5694 -148
rect 5739 -149 5786 -148
rect 5752 -154 5786 -149
rect 5520 -175 5694 -172
rect 5513 -178 5694 -175
rect 5722 -155 5786 -154
rect 5316 -198 5335 -196
rect 5350 -198 5384 -196
rect 5316 -214 5396 -198
rect 5316 -220 5335 -214
rect 5032 -246 5135 -236
rect 4986 -248 5135 -246
rect 5156 -248 5191 -236
rect 4825 -250 4987 -248
rect 4837 -268 4856 -250
rect 4871 -252 4901 -250
rect 4720 -278 4761 -270
rect 4844 -274 4856 -268
rect 4908 -266 4987 -250
rect 5019 -250 5191 -248
rect 5019 -266 5098 -250
rect 5105 -252 5135 -250
rect 4683 -288 4712 -278
rect 4726 -288 4755 -278
rect 4770 -288 4800 -274
rect 4844 -288 4886 -274
rect 4908 -278 5098 -266
rect 5163 -270 5169 -250
rect 4893 -288 4923 -278
rect 4924 -288 5082 -278
rect 5086 -288 5116 -278
rect 5120 -288 5150 -274
rect 5178 -288 5191 -250
rect 5263 -236 5292 -220
rect 5306 -236 5335 -220
rect 5350 -230 5380 -214
rect 5408 -236 5414 -188
rect 5417 -194 5436 -188
rect 5451 -194 5481 -186
rect 5417 -202 5481 -194
rect 5417 -218 5497 -202
rect 5513 -209 5575 -178
rect 5591 -209 5653 -178
rect 5722 -180 5771 -155
rect 5786 -180 5816 -162
rect 5685 -194 5715 -186
rect 5722 -188 5832 -180
rect 5685 -202 5730 -194
rect 5417 -220 5436 -218
rect 5451 -220 5497 -218
rect 5417 -236 5497 -220
rect 5524 -222 5559 -209
rect 5600 -212 5637 -209
rect 5600 -214 5642 -212
rect 5529 -225 5559 -222
rect 5538 -229 5545 -225
rect 5545 -230 5546 -229
rect 5504 -236 5514 -230
rect 5263 -244 5298 -236
rect 5263 -270 5264 -244
rect 5271 -270 5298 -244
rect 5206 -288 5236 -274
rect 5263 -278 5298 -270
rect 5300 -244 5341 -236
rect 5300 -270 5315 -244
rect 5322 -270 5341 -244
rect 5405 -248 5436 -236
rect 5451 -248 5554 -236
rect 5566 -246 5592 -220
rect 5607 -225 5637 -214
rect 5669 -218 5731 -202
rect 5669 -220 5715 -218
rect 5669 -236 5731 -220
rect 5743 -236 5749 -188
rect 5752 -196 5832 -188
rect 5752 -198 5771 -196
rect 5786 -198 5820 -196
rect 5752 -213 5832 -198
rect 5752 -214 5838 -213
rect 5752 -236 5771 -214
rect 5786 -230 5816 -214
rect 5844 -220 5850 -146
rect 5853 -220 5872 -76
rect 5887 -220 5893 -76
rect 5902 -146 5915 -76
rect 5967 -80 5989 -76
rect 5960 -92 5977 -88
rect 5981 -90 5989 -88
rect 5979 -92 5989 -90
rect 5960 -102 5989 -92
rect 6042 -102 6058 -88
rect 6096 -92 6102 -90
rect 6109 -92 6217 -76
rect 6224 -92 6230 -90
rect 6238 -92 6253 -76
rect 6319 -82 6338 -79
rect 5960 -104 6058 -102
rect 6085 -104 6253 -92
rect 6268 -102 6284 -88
rect 6319 -101 6341 -82
rect 6351 -88 6367 -87
rect 6350 -90 6367 -88
rect 6351 -95 6367 -90
rect 6341 -102 6347 -101
rect 6350 -102 6379 -95
rect 6268 -103 6379 -102
rect 6268 -104 6385 -103
rect 5944 -112 5995 -104
rect 6042 -112 6076 -104
rect 5944 -124 5969 -112
rect 5976 -124 5995 -112
rect 6049 -114 6076 -112
rect 6085 -114 6306 -104
rect 6341 -107 6347 -104
rect 6049 -118 6306 -114
rect 5944 -132 5995 -124
rect 6042 -132 6306 -118
rect 6350 -112 6385 -104
rect 5896 -180 5915 -146
rect 5960 -140 5989 -132
rect 5960 -146 5977 -140
rect 5960 -148 5994 -146
rect 6042 -148 6058 -132
rect 6059 -142 6267 -132
rect 6268 -142 6284 -132
rect 6332 -136 6347 -121
rect 6350 -124 6351 -112
rect 6358 -124 6385 -112
rect 6350 -132 6385 -124
rect 6350 -133 6379 -132
rect 6070 -146 6284 -142
rect 6085 -148 6284 -146
rect 6319 -146 6332 -136
rect 6350 -146 6367 -133
rect 6319 -148 6367 -146
rect 5961 -152 5994 -148
rect 5957 -154 5994 -152
rect 5957 -155 6024 -154
rect 5957 -160 5988 -155
rect 5994 -160 6024 -155
rect 5957 -164 6024 -160
rect 5930 -167 6024 -164
rect 5930 -174 5979 -167
rect 5930 -180 5960 -174
rect 5979 -179 5984 -174
rect 5896 -196 5976 -180
rect 5988 -188 6024 -167
rect 6085 -172 6274 -148
rect 6319 -149 6366 -148
rect 6332 -154 6366 -149
rect 6100 -175 6274 -172
rect 6093 -178 6274 -175
rect 6302 -155 6366 -154
rect 5896 -198 5915 -196
rect 5930 -198 5964 -196
rect 5896 -214 5976 -198
rect 5896 -220 5915 -214
rect 5612 -246 5715 -236
rect 5566 -248 5715 -246
rect 5736 -248 5771 -236
rect 5405 -250 5567 -248
rect 5417 -268 5436 -250
rect 5451 -252 5481 -250
rect 5300 -278 5341 -270
rect 5424 -274 5436 -268
rect 5488 -268 5567 -250
rect 5599 -250 5771 -248
rect 5599 -266 5678 -250
rect 5685 -252 5715 -250
rect 5574 -268 5678 -266
rect 5263 -288 5292 -278
rect 5306 -288 5335 -278
rect 5350 -288 5380 -274
rect 5424 -288 5466 -274
rect 5488 -278 5678 -268
rect 5743 -270 5749 -250
rect 5473 -288 5503 -278
rect 5504 -288 5662 -278
rect 5666 -288 5696 -278
rect 5700 -288 5730 -274
rect 5758 -288 5771 -250
rect 5843 -236 5872 -220
rect 5886 -236 5915 -220
rect 5930 -230 5960 -214
rect 5988 -236 5994 -188
rect 5997 -194 6016 -188
rect 6031 -194 6061 -186
rect 5997 -202 6061 -194
rect 5997 -218 6077 -202
rect 6093 -209 6155 -178
rect 6171 -209 6233 -178
rect 6302 -180 6351 -155
rect 6366 -180 6396 -164
rect 6265 -194 6295 -186
rect 6302 -188 6412 -180
rect 6265 -202 6310 -194
rect 5997 -220 6016 -218
rect 6031 -220 6077 -218
rect 5997 -236 6077 -220
rect 6104 -222 6139 -209
rect 6180 -212 6217 -209
rect 6180 -214 6222 -212
rect 6109 -225 6139 -222
rect 6118 -229 6125 -225
rect 6125 -230 6126 -229
rect 6084 -236 6094 -230
rect 5843 -244 5878 -236
rect 5843 -270 5844 -244
rect 5851 -270 5878 -244
rect 5786 -288 5816 -274
rect 5843 -278 5878 -270
rect 5880 -244 5921 -236
rect 5880 -270 5895 -244
rect 5902 -270 5921 -244
rect 5985 -248 6016 -236
rect 6031 -248 6134 -236
rect 6146 -246 6172 -220
rect 6187 -225 6217 -214
rect 6249 -218 6311 -202
rect 6249 -220 6295 -218
rect 6249 -236 6311 -220
rect 6323 -236 6329 -188
rect 6332 -196 6412 -188
rect 6332 -198 6351 -196
rect 6366 -198 6400 -196
rect 6332 -214 6412 -198
rect 6332 -236 6351 -214
rect 6366 -230 6396 -214
rect 6424 -220 6430 -146
rect 6439 -220 6452 -76
rect 6192 -246 6295 -236
rect 6146 -248 6295 -246
rect 6316 -248 6351 -236
rect 5985 -250 6147 -248
rect 5997 -268 6016 -250
rect 6031 -252 6061 -250
rect 5880 -278 5921 -270
rect 6004 -274 6016 -268
rect 6068 -268 6147 -250
rect 6179 -250 6351 -248
rect 6179 -266 6258 -250
rect 6265 -252 6295 -250
rect 6154 -268 6258 -266
rect 5843 -288 5872 -278
rect 5886 -288 5915 -278
rect 5930 -288 5960 -274
rect 6004 -288 6046 -274
rect 6068 -278 6258 -268
rect 6323 -270 6329 -250
rect 6053 -288 6083 -278
rect 6084 -288 6242 -278
rect 6246 -288 6276 -278
rect 6280 -288 6310 -274
rect 6338 -288 6351 -250
rect 6423 -236 6452 -220
rect 6423 -244 6458 -236
rect 6423 -270 6424 -244
rect 6431 -270 6458 -244
rect 6366 -288 6396 -274
rect 6423 -278 6458 -270
rect 6423 -288 6452 -278
rect -541 -302 6452 -288
rect -478 -332 -465 -302
rect -450 -316 -420 -302
rect -376 -316 -334 -302
rect -327 -316 -107 -302
rect -100 -316 -70 -302
rect -410 -330 -395 -318
rect -376 -330 -363 -316
rect -295 -320 -142 -316
rect -413 -332 -391 -330
rect -313 -332 -121 -320
rect -42 -332 -29 -302
rect -14 -316 16 -302
rect 53 -332 72 -302
rect 87 -332 93 -302
rect 102 -332 115 -302
rect 130 -316 160 -302
rect 204 -316 246 -302
rect 253 -316 473 -302
rect 480 -316 510 -302
rect 170 -330 185 -318
rect 204 -330 217 -316
rect 285 -320 438 -316
rect 167 -332 189 -330
rect 267 -332 459 -320
rect 538 -332 551 -302
rect 566 -316 596 -302
rect 633 -332 652 -302
rect 667 -332 673 -302
rect 682 -332 695 -302
rect 710 -316 740 -302
rect 784 -316 826 -302
rect 833 -316 1053 -302
rect 1060 -316 1090 -302
rect 750 -330 765 -318
rect 784 -330 797 -316
rect 865 -320 1018 -316
rect 747 -332 769 -330
rect 847 -332 1039 -320
rect 1118 -332 1131 -302
rect 1146 -316 1176 -302
rect 1213 -332 1232 -302
rect 1247 -332 1253 -302
rect 1262 -332 1275 -302
rect 1290 -316 1320 -302
rect 1364 -316 1406 -302
rect 1413 -316 1633 -302
rect 1640 -316 1670 -302
rect 1330 -330 1345 -318
rect 1364 -330 1377 -316
rect 1445 -320 1598 -316
rect 1327 -332 1349 -330
rect 1427 -332 1619 -320
rect 1698 -332 1711 -302
rect 1726 -316 1756 -302
rect 1793 -332 1812 -302
rect 1827 -332 1833 -302
rect 1842 -332 1855 -302
rect 1870 -316 1900 -302
rect 1944 -316 1986 -302
rect 1993 -316 2213 -302
rect 2220 -316 2250 -302
rect 1910 -330 1925 -318
rect 1944 -330 1957 -316
rect 2025 -320 2178 -316
rect 1907 -332 1929 -330
rect 2007 -332 2199 -320
rect 2278 -332 2291 -302
rect 2306 -316 2336 -302
rect 2373 -332 2392 -302
rect 2407 -332 2413 -302
rect 2422 -332 2435 -302
rect 2450 -316 2480 -302
rect 2524 -316 2566 -302
rect 2573 -316 2793 -302
rect 2800 -316 2830 -302
rect 2490 -330 2505 -318
rect 2524 -330 2537 -316
rect 2605 -320 2758 -316
rect 2487 -332 2509 -330
rect 2587 -332 2779 -320
rect 2858 -332 2871 -302
rect 2886 -316 2916 -302
rect 2953 -332 2972 -302
rect 2987 -332 2993 -302
rect 3002 -332 3015 -302
rect 3030 -316 3060 -302
rect 3104 -316 3146 -302
rect 3153 -316 3373 -302
rect 3380 -316 3410 -302
rect 3070 -330 3085 -318
rect 3104 -330 3117 -316
rect 3185 -320 3338 -316
rect 3067 -332 3089 -330
rect 3167 -332 3359 -320
rect 3438 -332 3451 -302
rect 3466 -316 3496 -302
rect 3533 -332 3552 -302
rect 3567 -332 3573 -302
rect 3582 -332 3595 -302
rect 3610 -316 3640 -302
rect 3684 -316 3726 -302
rect 3733 -316 3953 -302
rect 3960 -316 3990 -302
rect 3650 -330 3665 -318
rect 3684 -330 3697 -316
rect 3765 -320 3918 -316
rect 3647 -332 3669 -330
rect 3747 -332 3939 -320
rect 4018 -332 4031 -302
rect 4046 -316 4076 -302
rect 4113 -332 4132 -302
rect 4147 -332 4153 -302
rect 4162 -332 4175 -302
rect 4190 -316 4220 -302
rect 4264 -316 4306 -302
rect 4313 -316 4533 -302
rect 4540 -316 4570 -302
rect 4230 -330 4245 -318
rect 4264 -330 4277 -316
rect 4345 -320 4498 -316
rect 4227 -332 4249 -330
rect 4327 -332 4519 -320
rect 4598 -332 4611 -302
rect 4626 -316 4656 -302
rect 4693 -332 4712 -302
rect 4727 -332 4733 -302
rect 4742 -332 4755 -302
rect 4770 -316 4800 -302
rect 4844 -316 4886 -302
rect 4893 -316 5113 -302
rect 5120 -316 5150 -302
rect 4810 -330 4825 -318
rect 4844 -330 4857 -316
rect 4925 -320 5078 -316
rect 4807 -332 4829 -330
rect 4907 -332 5099 -320
rect 5178 -332 5191 -302
rect 5206 -316 5236 -302
rect 5273 -332 5292 -302
rect 5307 -332 5313 -302
rect 5322 -332 5335 -302
rect 5350 -316 5380 -302
rect 5424 -316 5466 -302
rect 5473 -316 5693 -302
rect 5700 -316 5730 -302
rect 5390 -330 5405 -318
rect 5424 -330 5437 -316
rect 5505 -320 5658 -316
rect 5387 -332 5409 -330
rect 5487 -332 5679 -320
rect 5758 -332 5771 -302
rect 5786 -316 5816 -302
rect 5853 -332 5872 -302
rect 5887 -332 5893 -302
rect 5902 -332 5915 -302
rect 5930 -316 5960 -302
rect 6004 -316 6046 -302
rect 6053 -316 6273 -302
rect 6280 -316 6310 -302
rect 5970 -330 5985 -318
rect 6004 -330 6017 -316
rect 6085 -320 6238 -316
rect 5967 -332 5989 -330
rect 6067 -332 6259 -320
rect 6338 -332 6351 -302
rect 6366 -316 6396 -302
rect 6439 -332 6452 -302
rect -541 -346 6452 -332
rect -478 -416 -465 -346
rect -413 -350 -391 -346
rect -420 -362 -403 -358
rect -399 -360 -391 -358
rect -401 -362 -391 -360
rect -420 -372 -391 -362
rect -338 -372 -322 -358
rect -284 -362 -278 -360
rect -271 -362 -163 -346
rect -156 -362 -150 -360
rect -142 -362 -127 -346
rect -61 -352 -42 -349
rect -420 -374 -322 -372
rect -295 -374 -127 -362
rect -112 -372 -96 -358
rect -61 -371 -39 -352
rect -29 -358 -13 -357
rect -30 -360 -13 -358
rect -29 -365 -13 -360
rect -39 -372 -33 -371
rect -30 -372 -1 -365
rect -112 -373 -1 -372
rect -112 -374 5 -373
rect -436 -382 -385 -374
rect -338 -382 -304 -374
rect -436 -394 -411 -382
rect -404 -394 -385 -382
rect -331 -384 -304 -382
rect -295 -384 -74 -374
rect -39 -377 -33 -374
rect -331 -388 -74 -384
rect -436 -402 -385 -394
rect -338 -402 -74 -388
rect -30 -382 5 -374
rect -484 -450 -465 -416
rect -420 -410 -391 -402
rect -420 -416 -403 -410
rect -420 -418 -386 -416
rect -338 -418 -322 -402
rect -321 -412 -113 -402
rect -112 -412 -96 -402
rect -48 -406 -33 -391
rect -30 -394 -29 -382
rect -22 -394 5 -382
rect -30 -402 5 -394
rect -30 -403 -1 -402
rect -310 -416 -96 -412
rect -295 -418 -96 -416
rect -61 -416 -48 -406
rect -30 -416 -13 -403
rect -61 -418 -13 -416
rect -419 -422 -386 -418
rect -423 -424 -386 -422
rect -423 -425 -356 -424
rect -423 -430 -392 -425
rect -386 -430 -356 -425
rect -423 -434 -356 -430
rect -450 -437 -356 -434
rect -450 -444 -401 -437
rect -450 -450 -420 -444
rect -401 -449 -396 -444
rect -484 -466 -404 -450
rect -392 -458 -356 -437
rect -295 -442 -106 -418
rect -61 -419 -14 -418
rect -48 -424 -14 -419
rect -280 -445 -106 -442
rect -287 -448 -106 -445
rect -78 -425 -14 -424
rect -484 -468 -465 -466
rect -450 -468 -416 -466
rect -484 -484 -404 -468
rect -484 -490 -465 -484
rect -494 -506 -465 -490
rect -450 -500 -420 -484
rect -392 -506 -386 -458
rect -383 -464 -364 -458
rect -349 -464 -319 -456
rect -383 -472 -319 -464
rect -383 -488 -303 -472
rect -287 -479 -225 -448
rect -209 -479 -147 -448
rect -78 -450 -29 -425
rect -14 -450 16 -432
rect -115 -464 -85 -456
rect -78 -458 32 -450
rect -115 -472 -70 -464
rect -383 -490 -364 -488
rect -349 -490 -303 -488
rect -383 -506 -303 -490
rect -276 -492 -241 -479
rect -200 -482 -163 -479
rect -200 -484 -158 -482
rect -271 -495 -241 -492
rect -262 -499 -255 -495
rect -255 -500 -254 -499
rect -296 -506 -286 -500
rect -500 -514 -459 -506
rect -500 -540 -485 -514
rect -478 -540 -459 -514
rect -395 -518 -364 -506
rect -349 -518 -246 -506
rect -234 -516 -208 -490
rect -193 -495 -163 -484
rect -131 -488 -69 -472
rect -131 -490 -85 -488
rect -131 -506 -69 -490
rect -57 -506 -51 -458
rect -48 -466 32 -458
rect -48 -468 -29 -466
rect -14 -468 20 -466
rect -48 -483 32 -468
rect -48 -484 38 -483
rect -48 -506 -29 -484
rect -14 -500 16 -484
rect 44 -490 50 -416
rect 53 -490 72 -346
rect 87 -490 93 -346
rect 102 -416 115 -346
rect 167 -350 189 -346
rect 160 -362 177 -358
rect 181 -360 189 -358
rect 179 -362 189 -360
rect 160 -372 189 -362
rect 242 -372 258 -358
rect 296 -362 302 -360
rect 309 -362 417 -346
rect 424 -362 430 -360
rect 438 -362 453 -346
rect 519 -352 538 -349
rect 160 -374 258 -372
rect 285 -374 453 -362
rect 468 -372 484 -358
rect 519 -371 541 -352
rect 551 -358 567 -357
rect 550 -360 567 -358
rect 551 -365 567 -360
rect 541 -372 547 -371
rect 550 -372 579 -365
rect 468 -373 579 -372
rect 468 -374 585 -373
rect 144 -382 195 -374
rect 242 -382 276 -374
rect 144 -394 169 -382
rect 176 -394 195 -382
rect 249 -384 276 -382
rect 285 -384 506 -374
rect 541 -377 547 -374
rect 249 -388 506 -384
rect 144 -402 195 -394
rect 242 -402 506 -388
rect 550 -382 585 -374
rect 96 -450 115 -416
rect 160 -410 189 -402
rect 160 -416 177 -410
rect 160 -418 194 -416
rect 242 -418 258 -402
rect 259 -412 467 -402
rect 468 -412 484 -402
rect 532 -406 547 -391
rect 550 -394 551 -382
rect 558 -394 585 -382
rect 550 -402 585 -394
rect 550 -403 579 -402
rect 270 -416 484 -412
rect 285 -418 484 -416
rect 519 -416 532 -406
rect 550 -416 567 -403
rect 519 -418 567 -416
rect 161 -422 194 -418
rect 157 -424 194 -422
rect 157 -425 224 -424
rect 157 -430 188 -425
rect 194 -430 224 -425
rect 157 -434 224 -430
rect 130 -437 224 -434
rect 130 -444 179 -437
rect 130 -450 160 -444
rect 179 -449 184 -444
rect 96 -466 176 -450
rect 188 -458 224 -437
rect 285 -442 474 -418
rect 519 -419 566 -418
rect 532 -424 566 -419
rect 606 -424 622 -422
rect 300 -445 474 -442
rect 293 -448 474 -445
rect 502 -425 566 -424
rect 96 -468 115 -466
rect 130 -468 164 -466
rect 96 -484 176 -468
rect 96 -490 115 -484
rect -188 -516 -85 -506
rect -234 -518 -85 -516
rect -64 -518 -29 -506
rect -395 -520 -233 -518
rect -383 -540 -364 -520
rect -349 -522 -319 -520
rect -500 -548 -459 -540
rect -377 -544 -364 -540
rect -312 -536 -233 -520
rect -201 -520 -29 -518
rect -201 -536 -122 -520
rect -115 -522 -85 -520
rect -494 -558 -465 -548
rect -450 -558 -420 -544
rect -377 -558 -334 -544
rect -312 -548 -122 -536
rect -57 -540 -51 -520
rect -327 -558 -297 -548
rect -296 -558 -138 -548
rect -134 -558 -104 -548
rect -100 -558 -70 -544
rect -42 -558 -29 -520
rect 43 -506 72 -490
rect 86 -506 115 -490
rect 130 -500 160 -484
rect 188 -506 194 -458
rect 197 -464 216 -458
rect 231 -464 261 -456
rect 197 -472 261 -464
rect 197 -488 277 -472
rect 293 -479 355 -448
rect 371 -479 433 -448
rect 502 -450 551 -425
rect 596 -434 622 -424
rect 566 -450 622 -434
rect 465 -464 495 -456
rect 502 -458 612 -450
rect 465 -472 510 -464
rect 197 -490 216 -488
rect 231 -490 277 -488
rect 197 -506 277 -490
rect 304 -492 339 -479
rect 380 -482 417 -479
rect 380 -484 422 -482
rect 309 -495 339 -492
rect 318 -499 325 -495
rect 325 -500 326 -499
rect 284 -506 294 -500
rect 43 -514 78 -506
rect 43 -540 44 -514
rect 51 -540 78 -514
rect -14 -558 16 -544
rect 43 -548 78 -540
rect 80 -514 121 -506
rect 80 -540 95 -514
rect 102 -540 121 -514
rect 185 -518 216 -506
rect 231 -518 334 -506
rect 346 -516 372 -490
rect 387 -495 417 -484
rect 449 -488 511 -472
rect 449 -490 495 -488
rect 449 -506 511 -490
rect 523 -506 529 -458
rect 532 -466 612 -458
rect 532 -468 551 -466
rect 566 -468 600 -466
rect 532 -484 612 -468
rect 532 -506 551 -484
rect 566 -500 596 -484
rect 624 -490 630 -416
rect 633 -490 652 -346
rect 667 -490 673 -346
rect 682 -416 695 -346
rect 747 -350 769 -346
rect 740 -362 757 -358
rect 761 -360 769 -358
rect 759 -362 769 -360
rect 740 -372 769 -362
rect 822 -372 838 -358
rect 876 -362 882 -360
rect 889 -362 997 -346
rect 1004 -362 1010 -360
rect 1018 -362 1033 -346
rect 1099 -352 1118 -349
rect 740 -374 838 -372
rect 865 -374 1033 -362
rect 1048 -372 1064 -358
rect 1099 -371 1121 -352
rect 1131 -358 1147 -357
rect 1130 -360 1147 -358
rect 1131 -365 1147 -360
rect 1121 -372 1127 -371
rect 1130 -372 1159 -365
rect 1048 -373 1159 -372
rect 1048 -374 1165 -373
rect 724 -382 775 -374
rect 822 -382 856 -374
rect 724 -394 749 -382
rect 756 -394 775 -382
rect 829 -384 856 -382
rect 865 -384 1086 -374
rect 1121 -377 1127 -374
rect 829 -388 1086 -384
rect 724 -402 775 -394
rect 822 -402 1086 -388
rect 1130 -382 1165 -374
rect 676 -450 695 -416
rect 740 -410 769 -402
rect 740 -416 757 -410
rect 740 -418 774 -416
rect 822 -418 838 -402
rect 839 -412 1047 -402
rect 1048 -412 1064 -402
rect 1112 -406 1127 -391
rect 1130 -394 1131 -382
rect 1138 -394 1165 -382
rect 1130 -402 1165 -394
rect 1130 -403 1159 -402
rect 850 -416 1064 -412
rect 865 -418 1064 -416
rect 1099 -416 1112 -406
rect 1130 -416 1147 -403
rect 1099 -418 1147 -416
rect 741 -422 774 -418
rect 737 -424 774 -422
rect 737 -425 804 -424
rect 737 -430 768 -425
rect 774 -430 804 -425
rect 737 -434 804 -430
rect 710 -437 804 -434
rect 710 -444 759 -437
rect 710 -450 740 -444
rect 759 -449 764 -444
rect 676 -466 756 -450
rect 768 -458 804 -437
rect 865 -442 1054 -418
rect 1099 -419 1146 -418
rect 1112 -424 1146 -419
rect 880 -445 1054 -442
rect 873 -448 1054 -445
rect 1082 -425 1146 -424
rect 676 -468 695 -466
rect 710 -468 744 -466
rect 676 -484 756 -468
rect 676 -490 695 -484
rect 392 -516 495 -506
rect 346 -518 495 -516
rect 516 -518 551 -506
rect 185 -520 347 -518
rect 197 -540 216 -520
rect 231 -522 261 -520
rect 80 -548 121 -540
rect 203 -544 216 -540
rect 268 -536 347 -520
rect 379 -520 551 -518
rect 379 -536 458 -520
rect 465 -522 495 -520
rect 43 -558 72 -548
rect 86 -558 115 -548
rect 130 -558 160 -544
rect 203 -558 246 -544
rect 268 -548 458 -536
rect 523 -540 529 -520
rect 253 -558 283 -548
rect 284 -558 442 -548
rect 446 -558 476 -548
rect 480 -558 510 -544
rect 538 -558 551 -520
rect 623 -506 652 -490
rect 666 -506 695 -490
rect 710 -500 740 -484
rect 768 -506 774 -458
rect 777 -464 796 -458
rect 811 -464 841 -456
rect 777 -472 841 -464
rect 777 -488 857 -472
rect 873 -479 935 -448
rect 951 -479 1013 -448
rect 1082 -450 1131 -425
rect 1146 -450 1176 -432
rect 1045 -464 1075 -456
rect 1082 -458 1192 -450
rect 1045 -472 1090 -464
rect 777 -490 796 -488
rect 811 -490 857 -488
rect 777 -506 857 -490
rect 884 -492 919 -479
rect 960 -482 997 -479
rect 960 -484 1002 -482
rect 889 -495 919 -492
rect 898 -499 905 -495
rect 905 -500 906 -499
rect 864 -506 874 -500
rect 623 -514 658 -506
rect 623 -540 624 -514
rect 631 -540 658 -514
rect 566 -558 596 -544
rect 623 -548 658 -540
rect 660 -514 701 -506
rect 660 -540 675 -514
rect 682 -540 701 -514
rect 765 -518 796 -506
rect 811 -518 914 -506
rect 926 -516 952 -490
rect 967 -495 997 -484
rect 1029 -488 1091 -472
rect 1029 -490 1075 -488
rect 1029 -506 1091 -490
rect 1103 -506 1109 -458
rect 1112 -466 1192 -458
rect 1112 -468 1131 -466
rect 1146 -468 1180 -466
rect 1112 -483 1192 -468
rect 1112 -484 1198 -483
rect 1112 -506 1131 -484
rect 1146 -500 1176 -484
rect 1204 -490 1210 -416
rect 1213 -490 1232 -346
rect 1247 -490 1253 -346
rect 1262 -416 1275 -346
rect 1327 -350 1349 -346
rect 1320 -362 1337 -358
rect 1341 -360 1349 -358
rect 1339 -362 1349 -360
rect 1320 -372 1349 -362
rect 1402 -372 1418 -358
rect 1456 -362 1462 -360
rect 1469 -362 1577 -346
rect 1584 -362 1590 -360
rect 1598 -362 1613 -346
rect 1679 -352 1698 -349
rect 1320 -374 1418 -372
rect 1445 -374 1613 -362
rect 1628 -372 1644 -358
rect 1679 -371 1701 -352
rect 1711 -358 1727 -357
rect 1710 -360 1727 -358
rect 1711 -365 1727 -360
rect 1701 -372 1707 -371
rect 1710 -372 1739 -365
rect 1628 -373 1739 -372
rect 1628 -374 1745 -373
rect 1304 -382 1355 -374
rect 1402 -382 1436 -374
rect 1304 -394 1329 -382
rect 1336 -394 1355 -382
rect 1409 -384 1436 -382
rect 1445 -384 1666 -374
rect 1701 -377 1707 -374
rect 1409 -388 1666 -384
rect 1304 -402 1355 -394
rect 1402 -402 1666 -388
rect 1710 -382 1745 -374
rect 1256 -450 1275 -416
rect 1320 -410 1349 -402
rect 1320 -416 1337 -410
rect 1320 -418 1354 -416
rect 1402 -418 1418 -402
rect 1419 -412 1627 -402
rect 1628 -412 1644 -402
rect 1692 -406 1707 -391
rect 1710 -394 1711 -382
rect 1718 -394 1745 -382
rect 1710 -402 1745 -394
rect 1710 -403 1739 -402
rect 1430 -416 1644 -412
rect 1445 -418 1644 -416
rect 1679 -416 1692 -406
rect 1710 -416 1727 -403
rect 1679 -418 1727 -416
rect 1321 -422 1354 -418
rect 1317 -424 1354 -422
rect 1317 -425 1384 -424
rect 1317 -430 1348 -425
rect 1354 -430 1384 -425
rect 1317 -434 1384 -430
rect 1290 -437 1384 -434
rect 1290 -444 1339 -437
rect 1290 -450 1320 -444
rect 1339 -449 1344 -444
rect 1256 -466 1336 -450
rect 1348 -458 1384 -437
rect 1445 -442 1634 -418
rect 1679 -419 1726 -418
rect 1692 -424 1726 -419
rect 1766 -424 1782 -422
rect 1460 -445 1634 -442
rect 1453 -448 1634 -445
rect 1662 -425 1726 -424
rect 1256 -468 1275 -466
rect 1290 -468 1324 -466
rect 1256 -484 1336 -468
rect 1256 -490 1275 -484
rect 972 -516 1075 -506
rect 926 -518 1075 -516
rect 1096 -518 1131 -506
rect 765 -520 927 -518
rect 777 -540 796 -520
rect 811 -522 841 -520
rect 660 -548 701 -540
rect 783 -544 796 -540
rect 848 -536 927 -520
rect 959 -520 1131 -518
rect 959 -536 1038 -520
rect 1045 -522 1075 -520
rect 623 -558 652 -548
rect 666 -558 695 -548
rect 710 -558 740 -544
rect 783 -558 826 -544
rect 848 -548 1038 -536
rect 1103 -540 1109 -520
rect 833 -558 863 -548
rect 864 -558 1022 -548
rect 1026 -558 1056 -548
rect 1060 -558 1090 -544
rect 1118 -558 1131 -520
rect 1203 -506 1232 -490
rect 1246 -506 1275 -490
rect 1290 -500 1320 -484
rect 1348 -506 1354 -458
rect 1357 -464 1376 -458
rect 1391 -464 1421 -456
rect 1357 -472 1421 -464
rect 1357 -488 1437 -472
rect 1453 -479 1515 -448
rect 1531 -479 1593 -448
rect 1662 -450 1711 -425
rect 1756 -434 1782 -424
rect 1726 -450 1782 -434
rect 1625 -464 1655 -456
rect 1662 -458 1772 -450
rect 1625 -472 1670 -464
rect 1357 -490 1376 -488
rect 1391 -490 1437 -488
rect 1357 -506 1437 -490
rect 1464 -492 1499 -479
rect 1540 -482 1577 -479
rect 1540 -484 1582 -482
rect 1469 -495 1499 -492
rect 1478 -499 1485 -495
rect 1485 -500 1486 -499
rect 1444 -506 1454 -500
rect 1203 -514 1238 -506
rect 1203 -540 1204 -514
rect 1211 -540 1238 -514
rect 1146 -558 1176 -544
rect 1203 -548 1238 -540
rect 1240 -514 1281 -506
rect 1240 -540 1255 -514
rect 1262 -540 1281 -514
rect 1345 -518 1376 -506
rect 1391 -518 1494 -506
rect 1506 -516 1532 -490
rect 1547 -495 1577 -484
rect 1609 -488 1671 -472
rect 1609 -490 1655 -488
rect 1609 -506 1671 -490
rect 1683 -506 1689 -458
rect 1692 -466 1772 -458
rect 1692 -468 1711 -466
rect 1726 -468 1760 -466
rect 1692 -484 1772 -468
rect 1692 -506 1711 -484
rect 1726 -500 1756 -484
rect 1784 -490 1790 -416
rect 1793 -490 1812 -346
rect 1827 -490 1833 -346
rect 1842 -416 1855 -346
rect 1907 -350 1929 -346
rect 1900 -362 1917 -358
rect 1921 -360 1929 -358
rect 1919 -362 1929 -360
rect 1900 -372 1929 -362
rect 1982 -372 1998 -358
rect 2036 -362 2042 -360
rect 2049 -362 2157 -346
rect 2164 -362 2170 -360
rect 2178 -362 2193 -346
rect 2259 -352 2278 -349
rect 1900 -374 1998 -372
rect 2025 -374 2193 -362
rect 2208 -372 2224 -358
rect 2259 -371 2281 -352
rect 2291 -358 2307 -357
rect 2290 -364 2307 -358
rect 2291 -365 2307 -364
rect 2281 -372 2287 -371
rect 2290 -372 2319 -365
rect 2208 -373 2319 -372
rect 2208 -374 2325 -373
rect 1884 -382 1935 -374
rect 1982 -382 2016 -374
rect 1884 -394 1909 -382
rect 1916 -394 1935 -382
rect 1989 -384 2016 -382
rect 2025 -384 2246 -374
rect 2281 -377 2287 -374
rect 1989 -388 2246 -384
rect 1884 -402 1935 -394
rect 1982 -402 2246 -388
rect 2290 -382 2325 -374
rect 1836 -450 1855 -416
rect 1900 -410 1929 -402
rect 1900 -416 1917 -410
rect 1900 -418 1934 -416
rect 1982 -418 1998 -402
rect 1999 -412 2207 -402
rect 2208 -412 2224 -402
rect 2272 -406 2287 -391
rect 2290 -394 2291 -382
rect 2298 -394 2325 -382
rect 2290 -402 2325 -394
rect 2290 -403 2319 -402
rect 2010 -416 2224 -412
rect 2025 -418 2224 -416
rect 2259 -416 2272 -406
rect 2290 -416 2307 -403
rect 2259 -418 2307 -416
rect 1901 -422 1934 -418
rect 1897 -424 1934 -422
rect 1897 -425 1964 -424
rect 1897 -430 1928 -425
rect 1934 -430 1964 -425
rect 1897 -434 1964 -430
rect 1870 -437 1964 -434
rect 1870 -444 1919 -437
rect 1870 -450 1900 -444
rect 1919 -449 1924 -444
rect 1836 -466 1916 -450
rect 1928 -458 1964 -437
rect 2025 -442 2214 -418
rect 2259 -419 2306 -418
rect 2272 -424 2306 -419
rect 2040 -445 2214 -442
rect 2033 -448 2214 -445
rect 2242 -425 2306 -424
rect 1836 -468 1855 -466
rect 1870 -468 1904 -466
rect 1836 -484 1916 -468
rect 1836 -490 1855 -484
rect 1552 -516 1655 -506
rect 1506 -518 1655 -516
rect 1676 -518 1711 -506
rect 1345 -520 1507 -518
rect 1357 -540 1376 -520
rect 1391 -522 1421 -520
rect 1240 -548 1281 -540
rect 1363 -544 1376 -540
rect 1428 -536 1507 -520
rect 1539 -520 1711 -518
rect 1539 -536 1618 -520
rect 1625 -522 1655 -520
rect 1203 -558 1232 -548
rect 1246 -558 1275 -548
rect 1290 -558 1320 -544
rect 1363 -558 1406 -544
rect 1428 -548 1618 -536
rect 1683 -540 1689 -520
rect 1413 -558 1443 -548
rect 1444 -558 1602 -548
rect 1606 -558 1636 -548
rect 1640 -558 1670 -544
rect 1698 -558 1711 -520
rect 1783 -506 1812 -490
rect 1826 -506 1855 -490
rect 1870 -500 1900 -484
rect 1928 -506 1934 -458
rect 1937 -464 1956 -458
rect 1971 -464 2001 -456
rect 1937 -472 2001 -464
rect 1937 -488 2017 -472
rect 2033 -479 2095 -448
rect 2111 -479 2173 -448
rect 2242 -450 2291 -425
rect 2306 -450 2336 -432
rect 2205 -464 2235 -456
rect 2242 -458 2352 -450
rect 2205 -472 2250 -464
rect 1937 -490 1956 -488
rect 1971 -490 2017 -488
rect 1937 -506 2017 -490
rect 2044 -492 2079 -479
rect 2120 -482 2157 -479
rect 2120 -484 2162 -482
rect 2049 -495 2079 -492
rect 2058 -499 2065 -495
rect 2065 -500 2066 -499
rect 2024 -506 2034 -500
rect 1783 -514 1818 -506
rect 1783 -540 1784 -514
rect 1791 -540 1818 -514
rect 1726 -558 1756 -544
rect 1783 -548 1818 -540
rect 1820 -514 1861 -506
rect 1820 -540 1835 -514
rect 1842 -540 1861 -514
rect 1925 -518 1956 -506
rect 1971 -518 2074 -506
rect 2086 -516 2112 -490
rect 2127 -495 2157 -484
rect 2189 -488 2251 -472
rect 2189 -490 2235 -488
rect 2189 -506 2251 -490
rect 2263 -506 2269 -458
rect 2272 -466 2352 -458
rect 2272 -468 2291 -466
rect 2306 -468 2340 -466
rect 2272 -483 2352 -468
rect 2272 -484 2358 -483
rect 2272 -506 2291 -484
rect 2306 -500 2336 -484
rect 2364 -490 2370 -416
rect 2373 -490 2392 -346
rect 2407 -490 2413 -346
rect 2422 -416 2435 -346
rect 2487 -350 2509 -346
rect 2480 -362 2497 -358
rect 2501 -360 2509 -358
rect 2499 -362 2509 -360
rect 2480 -372 2509 -362
rect 2562 -372 2578 -358
rect 2616 -362 2622 -360
rect 2629 -362 2737 -346
rect 2744 -362 2750 -360
rect 2758 -362 2773 -346
rect 2839 -352 2858 -349
rect 2480 -374 2578 -372
rect 2605 -374 2773 -362
rect 2788 -372 2804 -358
rect 2839 -371 2861 -352
rect 2871 -358 2887 -357
rect 2870 -364 2887 -358
rect 2871 -365 2887 -364
rect 2861 -372 2867 -371
rect 2870 -372 2899 -365
rect 2788 -373 2899 -372
rect 2788 -374 2905 -373
rect 2464 -382 2515 -374
rect 2562 -382 2596 -374
rect 2464 -394 2489 -382
rect 2496 -394 2515 -382
rect 2569 -384 2596 -382
rect 2605 -384 2826 -374
rect 2861 -377 2867 -374
rect 2569 -388 2826 -384
rect 2464 -402 2515 -394
rect 2562 -402 2826 -388
rect 2870 -382 2905 -374
rect 2416 -450 2435 -416
rect 2480 -410 2509 -402
rect 2480 -416 2497 -410
rect 2480 -418 2514 -416
rect 2562 -418 2578 -402
rect 2579 -412 2787 -402
rect 2788 -412 2804 -402
rect 2852 -406 2867 -391
rect 2870 -394 2871 -382
rect 2878 -394 2905 -382
rect 2870 -402 2905 -394
rect 2870 -403 2899 -402
rect 2590 -416 2804 -412
rect 2605 -418 2804 -416
rect 2839 -416 2852 -406
rect 2870 -416 2887 -403
rect 2839 -418 2887 -416
rect 2481 -422 2514 -418
rect 2477 -424 2514 -422
rect 2477 -425 2544 -424
rect 2477 -430 2508 -425
rect 2514 -430 2544 -425
rect 2477 -434 2544 -430
rect 2450 -437 2544 -434
rect 2450 -444 2499 -437
rect 2450 -450 2480 -444
rect 2499 -449 2504 -444
rect 2416 -466 2496 -450
rect 2508 -458 2544 -437
rect 2605 -442 2794 -418
rect 2839 -419 2886 -418
rect 2852 -424 2886 -419
rect 2926 -424 2942 -422
rect 2620 -445 2794 -442
rect 2613 -448 2794 -445
rect 2822 -425 2886 -424
rect 2416 -468 2435 -466
rect 2450 -468 2484 -466
rect 2416 -484 2496 -468
rect 2416 -490 2435 -484
rect 2132 -516 2235 -506
rect 2086 -518 2235 -516
rect 2256 -518 2291 -506
rect 1925 -520 2087 -518
rect 1937 -540 1956 -520
rect 1971 -522 2001 -520
rect 1820 -548 1861 -540
rect 1943 -544 1956 -540
rect 2008 -536 2087 -520
rect 2119 -520 2291 -518
rect 2119 -536 2198 -520
rect 2205 -522 2235 -520
rect 1783 -558 1812 -548
rect 1826 -558 1855 -548
rect 1870 -558 1900 -544
rect 1943 -558 1986 -544
rect 2008 -548 2198 -536
rect 2263 -540 2269 -520
rect 1993 -558 2023 -548
rect 2024 -558 2182 -548
rect 2186 -558 2216 -548
rect 2220 -558 2250 -544
rect 2278 -558 2291 -520
rect 2363 -506 2392 -490
rect 2406 -506 2435 -490
rect 2450 -500 2480 -484
rect 2508 -506 2514 -458
rect 2517 -464 2536 -458
rect 2551 -464 2581 -456
rect 2517 -472 2581 -464
rect 2517 -488 2597 -472
rect 2613 -479 2675 -448
rect 2691 -479 2753 -448
rect 2822 -450 2871 -425
rect 2916 -434 2942 -424
rect 2886 -450 2942 -434
rect 2785 -464 2815 -456
rect 2822 -458 2932 -450
rect 2785 -472 2830 -464
rect 2517 -490 2536 -488
rect 2551 -490 2597 -488
rect 2517 -506 2597 -490
rect 2624 -492 2659 -479
rect 2700 -482 2737 -479
rect 2700 -484 2742 -482
rect 2629 -495 2659 -492
rect 2638 -499 2645 -495
rect 2645 -500 2646 -499
rect 2604 -506 2614 -500
rect 2363 -514 2398 -506
rect 2363 -540 2364 -514
rect 2371 -540 2398 -514
rect 2306 -558 2336 -544
rect 2363 -548 2398 -540
rect 2400 -514 2441 -506
rect 2400 -540 2415 -514
rect 2422 -540 2441 -514
rect 2505 -518 2536 -506
rect 2551 -518 2654 -506
rect 2666 -516 2692 -490
rect 2707 -495 2737 -484
rect 2769 -488 2831 -472
rect 2769 -490 2815 -488
rect 2769 -506 2831 -490
rect 2843 -506 2849 -458
rect 2852 -466 2932 -458
rect 2852 -468 2871 -466
rect 2886 -468 2920 -466
rect 2852 -484 2932 -468
rect 2852 -506 2871 -484
rect 2886 -500 2916 -484
rect 2944 -490 2950 -416
rect 2953 -490 2972 -346
rect 2987 -490 2993 -346
rect 3002 -416 3015 -346
rect 3067 -350 3089 -346
rect 3060 -362 3077 -358
rect 3081 -360 3089 -358
rect 3079 -362 3089 -360
rect 3060 -372 3089 -362
rect 3142 -372 3158 -358
rect 3196 -362 3202 -360
rect 3209 -362 3317 -346
rect 3324 -362 3330 -360
rect 3338 -362 3353 -346
rect 3419 -352 3438 -349
rect 3060 -374 3158 -372
rect 3185 -374 3353 -362
rect 3368 -372 3384 -358
rect 3419 -371 3441 -352
rect 3451 -358 3467 -357
rect 3450 -364 3467 -358
rect 3451 -365 3467 -364
rect 3441 -372 3447 -371
rect 3450 -372 3479 -365
rect 3368 -373 3479 -372
rect 3368 -374 3485 -373
rect 3044 -382 3095 -374
rect 3142 -382 3176 -374
rect 3044 -394 3069 -382
rect 3076 -394 3095 -382
rect 3149 -384 3176 -382
rect 3185 -384 3406 -374
rect 3441 -377 3447 -374
rect 3149 -388 3406 -384
rect 3044 -402 3095 -394
rect 3142 -402 3406 -388
rect 3450 -382 3485 -374
rect 2996 -450 3015 -416
rect 3060 -410 3089 -402
rect 3060 -416 3077 -410
rect 3060 -418 3094 -416
rect 3142 -418 3158 -402
rect 3159 -412 3367 -402
rect 3368 -412 3384 -402
rect 3432 -406 3447 -391
rect 3450 -394 3451 -382
rect 3458 -394 3485 -382
rect 3450 -402 3485 -394
rect 3450 -403 3479 -402
rect 3170 -416 3384 -412
rect 3185 -418 3384 -416
rect 3419 -416 3432 -406
rect 3450 -416 3467 -403
rect 3419 -418 3467 -416
rect 3061 -422 3094 -418
rect 3057 -424 3094 -422
rect 3057 -425 3124 -424
rect 3057 -430 3088 -425
rect 3094 -430 3124 -425
rect 3057 -434 3124 -430
rect 3030 -437 3124 -434
rect 3030 -444 3079 -437
rect 3030 -450 3060 -444
rect 3079 -449 3084 -444
rect 2996 -466 3076 -450
rect 3088 -458 3124 -437
rect 3185 -442 3374 -418
rect 3419 -419 3466 -418
rect 3432 -424 3466 -419
rect 3200 -445 3374 -442
rect 3193 -448 3374 -445
rect 3402 -425 3466 -424
rect 2996 -468 3015 -466
rect 3030 -468 3064 -466
rect 2996 -484 3076 -468
rect 2996 -490 3015 -484
rect 2712 -516 2815 -506
rect 2666 -518 2815 -516
rect 2836 -518 2871 -506
rect 2505 -520 2667 -518
rect 2517 -540 2536 -520
rect 2551 -522 2581 -520
rect 2400 -548 2441 -540
rect 2523 -544 2536 -540
rect 2588 -536 2667 -520
rect 2699 -520 2871 -518
rect 2699 -536 2778 -520
rect 2785 -522 2815 -520
rect 2363 -558 2392 -548
rect 2406 -558 2435 -548
rect 2450 -558 2480 -544
rect 2523 -558 2566 -544
rect 2588 -548 2778 -536
rect 2843 -540 2849 -520
rect 2573 -558 2603 -548
rect 2604 -558 2762 -548
rect 2766 -558 2796 -548
rect 2800 -558 2830 -544
rect 2858 -558 2871 -520
rect 2943 -506 2972 -490
rect 2986 -506 3015 -490
rect 3030 -500 3060 -484
rect 3088 -506 3094 -458
rect 3097 -464 3116 -458
rect 3131 -464 3161 -456
rect 3097 -472 3161 -464
rect 3097 -488 3177 -472
rect 3193 -479 3255 -448
rect 3271 -479 3333 -448
rect 3402 -450 3451 -425
rect 3466 -450 3496 -432
rect 3365 -464 3395 -456
rect 3402 -458 3512 -450
rect 3365 -472 3410 -464
rect 3097 -490 3116 -488
rect 3131 -490 3177 -488
rect 3097 -506 3177 -490
rect 3204 -492 3239 -479
rect 3280 -482 3317 -479
rect 3280 -484 3322 -482
rect 3209 -495 3239 -492
rect 3218 -499 3225 -495
rect 3225 -500 3226 -499
rect 3184 -506 3194 -500
rect 2943 -514 2978 -506
rect 2943 -540 2944 -514
rect 2951 -540 2978 -514
rect 2886 -558 2916 -544
rect 2943 -548 2978 -540
rect 2980 -514 3021 -506
rect 2980 -540 2995 -514
rect 3002 -540 3021 -514
rect 3085 -518 3116 -506
rect 3131 -518 3234 -506
rect 3246 -516 3272 -490
rect 3287 -495 3317 -484
rect 3349 -488 3411 -472
rect 3349 -490 3395 -488
rect 3349 -506 3411 -490
rect 3423 -506 3429 -458
rect 3432 -466 3512 -458
rect 3432 -468 3451 -466
rect 3466 -468 3500 -466
rect 3432 -483 3512 -468
rect 3432 -484 3518 -483
rect 3432 -506 3451 -484
rect 3466 -500 3496 -484
rect 3524 -490 3530 -416
rect 3533 -490 3552 -346
rect 3567 -490 3573 -346
rect 3582 -416 3595 -346
rect 3647 -350 3669 -346
rect 3640 -362 3657 -358
rect 3661 -360 3669 -358
rect 3659 -362 3669 -360
rect 3640 -372 3669 -362
rect 3722 -372 3738 -358
rect 3776 -362 3782 -360
rect 3789 -362 3897 -346
rect 3904 -362 3910 -360
rect 3918 -362 3933 -346
rect 3999 -352 4018 -349
rect 3640 -374 3738 -372
rect 3765 -374 3933 -362
rect 3948 -372 3964 -358
rect 3999 -371 4021 -352
rect 4031 -358 4047 -357
rect 4030 -364 4047 -358
rect 4031 -365 4047 -364
rect 4021 -372 4027 -371
rect 4030 -372 4059 -365
rect 3948 -373 4059 -372
rect 3948 -374 4065 -373
rect 3624 -382 3675 -374
rect 3722 -382 3756 -374
rect 3624 -394 3649 -382
rect 3656 -394 3675 -382
rect 3729 -384 3756 -382
rect 3765 -384 3986 -374
rect 4021 -377 4027 -374
rect 3729 -388 3986 -384
rect 3624 -402 3675 -394
rect 3722 -402 3986 -388
rect 4030 -382 4065 -374
rect 3576 -450 3595 -416
rect 3640 -410 3669 -402
rect 3640 -416 3657 -410
rect 3640 -418 3674 -416
rect 3722 -418 3738 -402
rect 3739 -412 3947 -402
rect 3948 -412 3964 -402
rect 4012 -406 4027 -391
rect 4030 -394 4031 -382
rect 4038 -394 4065 -382
rect 4030 -402 4065 -394
rect 4030 -403 4059 -402
rect 3750 -416 3964 -412
rect 3765 -418 3964 -416
rect 3999 -416 4012 -406
rect 4030 -416 4047 -403
rect 3999 -418 4047 -416
rect 3641 -422 3674 -418
rect 3637 -424 3674 -422
rect 3637 -425 3704 -424
rect 3637 -430 3668 -425
rect 3674 -430 3704 -425
rect 3637 -434 3704 -430
rect 3610 -437 3704 -434
rect 3610 -444 3659 -437
rect 3610 -450 3640 -444
rect 3659 -449 3664 -444
rect 3576 -466 3656 -450
rect 3668 -458 3704 -437
rect 3765 -442 3954 -418
rect 3999 -419 4046 -418
rect 4012 -424 4046 -419
rect 4086 -424 4102 -422
rect 3780 -445 3954 -442
rect 3773 -448 3954 -445
rect 3982 -425 4046 -424
rect 3576 -468 3595 -466
rect 3610 -468 3644 -466
rect 3576 -484 3656 -468
rect 3576 -490 3595 -484
rect 3292 -516 3395 -506
rect 3246 -518 3395 -516
rect 3416 -518 3451 -506
rect 3085 -520 3247 -518
rect 3097 -540 3116 -520
rect 3131 -522 3161 -520
rect 2980 -548 3021 -540
rect 3103 -544 3116 -540
rect 3168 -536 3247 -520
rect 3279 -520 3451 -518
rect 3279 -536 3358 -520
rect 3365 -522 3395 -520
rect 2943 -558 2972 -548
rect 2986 -558 3015 -548
rect 3030 -558 3060 -544
rect 3103 -558 3146 -544
rect 3168 -548 3358 -536
rect 3423 -540 3429 -520
rect 3153 -558 3183 -548
rect 3184 -558 3342 -548
rect 3346 -558 3376 -548
rect 3380 -558 3410 -544
rect 3438 -558 3451 -520
rect 3523 -506 3552 -490
rect 3566 -506 3595 -490
rect 3610 -500 3640 -484
rect 3668 -506 3674 -458
rect 3677 -464 3696 -458
rect 3711 -464 3741 -456
rect 3677 -472 3741 -464
rect 3677 -488 3757 -472
rect 3773 -479 3835 -448
rect 3851 -479 3913 -448
rect 3982 -450 4031 -425
rect 4076 -434 4102 -424
rect 4046 -450 4102 -434
rect 3945 -464 3975 -456
rect 3982 -458 4092 -450
rect 3945 -472 3990 -464
rect 3677 -490 3696 -488
rect 3711 -490 3757 -488
rect 3677 -506 3757 -490
rect 3784 -492 3819 -479
rect 3860 -482 3897 -479
rect 3860 -484 3902 -482
rect 3789 -495 3819 -492
rect 3798 -499 3805 -495
rect 3805 -500 3806 -499
rect 3764 -506 3774 -500
rect 3523 -514 3558 -506
rect 3523 -540 3524 -514
rect 3531 -540 3558 -514
rect 3466 -558 3496 -544
rect 3523 -548 3558 -540
rect 3560 -514 3601 -506
rect 3560 -540 3575 -514
rect 3582 -540 3601 -514
rect 3665 -518 3696 -506
rect 3711 -518 3814 -506
rect 3826 -516 3852 -490
rect 3867 -495 3897 -484
rect 3929 -488 3991 -472
rect 3929 -490 3975 -488
rect 3929 -506 3991 -490
rect 4003 -506 4009 -458
rect 4012 -466 4092 -458
rect 4012 -468 4031 -466
rect 4046 -468 4080 -466
rect 4012 -484 4092 -468
rect 4012 -506 4031 -484
rect 4046 -500 4076 -484
rect 4104 -490 4110 -416
rect 4113 -490 4132 -346
rect 4147 -490 4153 -346
rect 4162 -416 4175 -346
rect 4227 -350 4249 -346
rect 4220 -362 4237 -358
rect 4241 -360 4249 -358
rect 4239 -362 4249 -360
rect 4220 -372 4249 -362
rect 4302 -372 4318 -358
rect 4356 -362 4362 -360
rect 4369 -362 4477 -346
rect 4484 -362 4490 -360
rect 4498 -362 4513 -346
rect 4579 -352 4598 -349
rect 4220 -374 4318 -372
rect 4345 -374 4513 -362
rect 4528 -372 4544 -358
rect 4579 -371 4601 -352
rect 4611 -358 4627 -357
rect 4610 -364 4627 -358
rect 4611 -365 4627 -364
rect 4601 -372 4607 -371
rect 4610 -372 4639 -365
rect 4528 -373 4639 -372
rect 4528 -374 4645 -373
rect 4204 -382 4255 -374
rect 4302 -382 4336 -374
rect 4204 -394 4229 -382
rect 4236 -394 4255 -382
rect 4309 -384 4336 -382
rect 4345 -384 4566 -374
rect 4601 -377 4607 -374
rect 4309 -388 4566 -384
rect 4204 -402 4255 -394
rect 4302 -402 4566 -388
rect 4610 -382 4645 -374
rect 4156 -450 4175 -416
rect 4220 -410 4249 -402
rect 4220 -416 4237 -410
rect 4220 -418 4254 -416
rect 4302 -418 4318 -402
rect 4319 -412 4527 -402
rect 4528 -412 4544 -402
rect 4592 -406 4607 -391
rect 4610 -394 4611 -382
rect 4618 -394 4645 -382
rect 4610 -402 4645 -394
rect 4610 -403 4639 -402
rect 4330 -416 4544 -412
rect 4345 -418 4544 -416
rect 4579 -416 4592 -406
rect 4610 -416 4627 -403
rect 4579 -418 4627 -416
rect 4221 -422 4254 -418
rect 4217 -424 4254 -422
rect 4217 -425 4284 -424
rect 4217 -430 4248 -425
rect 4254 -430 4284 -425
rect 4217 -434 4284 -430
rect 4190 -437 4284 -434
rect 4190 -444 4239 -437
rect 4190 -450 4220 -444
rect 4239 -449 4244 -444
rect 4156 -466 4236 -450
rect 4248 -458 4284 -437
rect 4345 -442 4534 -418
rect 4579 -419 4626 -418
rect 4592 -424 4626 -419
rect 4360 -445 4534 -442
rect 4353 -448 4534 -445
rect 4562 -425 4626 -424
rect 4156 -468 4175 -466
rect 4190 -468 4224 -466
rect 4156 -484 4236 -468
rect 4156 -490 4175 -484
rect 3872 -516 3975 -506
rect 3826 -518 3975 -516
rect 3996 -518 4031 -506
rect 3665 -520 3827 -518
rect 3677 -540 3696 -520
rect 3711 -522 3741 -520
rect 3560 -548 3601 -540
rect 3683 -544 3696 -540
rect 3748 -536 3827 -520
rect 3859 -520 4031 -518
rect 3859 -536 3938 -520
rect 3945 -522 3975 -520
rect 3523 -558 3552 -548
rect 3566 -558 3595 -548
rect 3610 -558 3640 -544
rect 3683 -558 3726 -544
rect 3748 -548 3938 -536
rect 4003 -540 4009 -520
rect 3733 -558 3763 -548
rect 3764 -558 3922 -548
rect 3926 -558 3956 -548
rect 3960 -558 3990 -544
rect 4018 -558 4031 -520
rect 4103 -506 4132 -490
rect 4146 -506 4175 -490
rect 4190 -500 4220 -484
rect 4248 -506 4254 -458
rect 4257 -464 4276 -458
rect 4291 -464 4321 -456
rect 4257 -472 4321 -464
rect 4257 -488 4337 -472
rect 4353 -479 4415 -448
rect 4431 -479 4493 -448
rect 4562 -450 4611 -425
rect 4626 -450 4656 -432
rect 4525 -464 4555 -456
rect 4562 -458 4672 -450
rect 4525 -472 4570 -464
rect 4257 -490 4276 -488
rect 4291 -490 4337 -488
rect 4257 -506 4337 -490
rect 4364 -492 4399 -479
rect 4440 -482 4477 -479
rect 4440 -484 4482 -482
rect 4369 -495 4399 -492
rect 4378 -499 4385 -495
rect 4385 -500 4386 -499
rect 4344 -506 4354 -500
rect 4103 -514 4138 -506
rect 4103 -540 4104 -514
rect 4111 -540 4138 -514
rect 4046 -558 4076 -544
rect 4103 -548 4138 -540
rect 4140 -514 4181 -506
rect 4140 -540 4155 -514
rect 4162 -540 4181 -514
rect 4245 -518 4276 -506
rect 4291 -518 4394 -506
rect 4406 -516 4432 -490
rect 4447 -495 4477 -484
rect 4509 -488 4571 -472
rect 4509 -490 4555 -488
rect 4509 -506 4571 -490
rect 4583 -506 4589 -458
rect 4592 -466 4672 -458
rect 4592 -468 4611 -466
rect 4626 -468 4660 -466
rect 4592 -483 4672 -468
rect 4592 -484 4678 -483
rect 4592 -506 4611 -484
rect 4626 -500 4656 -484
rect 4684 -490 4690 -416
rect 4693 -490 4712 -346
rect 4727 -490 4733 -346
rect 4742 -416 4755 -346
rect 4807 -350 4829 -346
rect 4800 -362 4817 -358
rect 4821 -360 4829 -358
rect 4819 -362 4829 -360
rect 4800 -372 4829 -362
rect 4882 -372 4898 -358
rect 4936 -362 4942 -360
rect 4949 -362 5057 -346
rect 5064 -362 5070 -360
rect 5078 -362 5093 -346
rect 5159 -352 5178 -349
rect 4800 -374 4898 -372
rect 4925 -374 5093 -362
rect 5108 -372 5124 -358
rect 5159 -371 5181 -352
rect 5191 -358 5207 -357
rect 5190 -364 5207 -358
rect 5191 -365 5207 -364
rect 5181 -372 5187 -371
rect 5190 -372 5219 -365
rect 5108 -373 5219 -372
rect 5108 -374 5225 -373
rect 4784 -382 4835 -374
rect 4882 -382 4916 -374
rect 4784 -394 4809 -382
rect 4816 -394 4835 -382
rect 4889 -384 4916 -382
rect 4925 -384 5146 -374
rect 5181 -377 5187 -374
rect 4889 -388 5146 -384
rect 4784 -402 4835 -394
rect 4882 -402 5146 -388
rect 5190 -382 5225 -374
rect 4736 -450 4755 -416
rect 4800 -410 4829 -402
rect 4800 -416 4817 -410
rect 4800 -418 4834 -416
rect 4882 -418 4898 -402
rect 4899 -412 5107 -402
rect 5108 -412 5124 -402
rect 5172 -406 5187 -391
rect 5190 -394 5191 -382
rect 5198 -394 5225 -382
rect 5190 -402 5225 -394
rect 5190 -403 5219 -402
rect 4910 -416 5124 -412
rect 4925 -418 5124 -416
rect 5159 -416 5172 -406
rect 5190 -416 5207 -403
rect 5159 -418 5207 -416
rect 4801 -422 4834 -418
rect 4797 -424 4834 -422
rect 4797 -425 4864 -424
rect 4797 -430 4828 -425
rect 4834 -430 4864 -425
rect 4797 -434 4864 -430
rect 4770 -437 4864 -434
rect 4770 -444 4819 -437
rect 4770 -450 4800 -444
rect 4819 -449 4824 -444
rect 4736 -466 4816 -450
rect 4828 -458 4864 -437
rect 4925 -442 5114 -418
rect 5159 -419 5206 -418
rect 5172 -424 5206 -419
rect 5246 -424 5262 -422
rect 4940 -445 5114 -442
rect 4933 -448 5114 -445
rect 5142 -425 5206 -424
rect 4736 -468 4755 -466
rect 4770 -468 4804 -466
rect 4736 -484 4816 -468
rect 4736 -490 4755 -484
rect 4452 -516 4555 -506
rect 4406 -518 4555 -516
rect 4576 -518 4611 -506
rect 4245 -520 4407 -518
rect 4257 -540 4276 -520
rect 4291 -522 4321 -520
rect 4140 -548 4181 -540
rect 4263 -544 4276 -540
rect 4328 -536 4407 -520
rect 4439 -520 4611 -518
rect 4439 -536 4518 -520
rect 4525 -522 4555 -520
rect 4103 -558 4132 -548
rect 4146 -558 4175 -548
rect 4190 -558 4220 -544
rect 4263 -558 4306 -544
rect 4328 -548 4518 -536
rect 4583 -540 4589 -520
rect 4313 -558 4343 -548
rect 4344 -558 4502 -548
rect 4506 -558 4536 -548
rect 4540 -558 4570 -544
rect 4598 -558 4611 -520
rect 4683 -506 4712 -490
rect 4726 -506 4755 -490
rect 4770 -500 4800 -484
rect 4828 -506 4834 -458
rect 4837 -464 4856 -458
rect 4871 -464 4901 -456
rect 4837 -472 4901 -464
rect 4837 -488 4917 -472
rect 4933 -479 4995 -448
rect 5011 -479 5073 -448
rect 5142 -450 5191 -425
rect 5236 -434 5262 -424
rect 5206 -450 5262 -434
rect 5105 -464 5135 -456
rect 5142 -458 5252 -450
rect 5105 -472 5150 -464
rect 4837 -490 4856 -488
rect 4871 -490 4917 -488
rect 4837 -506 4917 -490
rect 4944 -492 4979 -479
rect 5020 -482 5057 -479
rect 5020 -484 5062 -482
rect 4949 -495 4979 -492
rect 4958 -499 4965 -495
rect 4965 -500 4966 -499
rect 4924 -506 4934 -500
rect 4683 -514 4718 -506
rect 4683 -540 4684 -514
rect 4691 -540 4718 -514
rect 4626 -558 4656 -544
rect 4683 -548 4718 -540
rect 4720 -514 4761 -506
rect 4720 -540 4735 -514
rect 4742 -540 4761 -514
rect 4825 -518 4856 -506
rect 4871 -518 4974 -506
rect 4986 -516 5012 -490
rect 5027 -495 5057 -484
rect 5089 -488 5151 -472
rect 5089 -490 5135 -488
rect 5089 -506 5151 -490
rect 5163 -506 5169 -458
rect 5172 -466 5252 -458
rect 5172 -468 5191 -466
rect 5206 -468 5240 -466
rect 5172 -484 5252 -468
rect 5172 -506 5191 -484
rect 5206 -500 5236 -484
rect 5264 -490 5270 -416
rect 5273 -490 5292 -346
rect 5307 -490 5313 -346
rect 5322 -416 5335 -346
rect 5387 -350 5409 -346
rect 5380 -362 5397 -358
rect 5401 -360 5409 -358
rect 5399 -362 5409 -360
rect 5380 -372 5409 -362
rect 5462 -372 5478 -358
rect 5516 -362 5522 -360
rect 5529 -362 5637 -346
rect 5644 -362 5650 -360
rect 5658 -362 5673 -346
rect 5739 -352 5758 -349
rect 5380 -374 5478 -372
rect 5505 -374 5673 -362
rect 5688 -372 5704 -358
rect 5739 -371 5761 -352
rect 5771 -358 5787 -357
rect 5770 -360 5787 -358
rect 5771 -365 5787 -360
rect 5761 -372 5767 -371
rect 5770 -372 5799 -365
rect 5688 -373 5799 -372
rect 5688 -374 5805 -373
rect 5364 -382 5415 -374
rect 5462 -382 5496 -374
rect 5364 -394 5389 -382
rect 5396 -394 5415 -382
rect 5469 -384 5496 -382
rect 5505 -384 5726 -374
rect 5761 -377 5767 -374
rect 5469 -388 5726 -384
rect 5364 -402 5415 -394
rect 5462 -402 5726 -388
rect 5770 -382 5805 -374
rect 5316 -450 5335 -416
rect 5380 -410 5409 -402
rect 5380 -416 5397 -410
rect 5380 -418 5414 -416
rect 5462 -418 5478 -402
rect 5479 -412 5687 -402
rect 5688 -412 5704 -402
rect 5752 -406 5767 -391
rect 5770 -394 5771 -382
rect 5778 -394 5805 -382
rect 5770 -402 5805 -394
rect 5770 -403 5799 -402
rect 5490 -416 5704 -412
rect 5505 -418 5704 -416
rect 5739 -416 5752 -406
rect 5770 -416 5787 -403
rect 5739 -418 5787 -416
rect 5381 -422 5414 -418
rect 5377 -424 5414 -422
rect 5377 -425 5444 -424
rect 5377 -430 5408 -425
rect 5414 -430 5444 -425
rect 5377 -434 5444 -430
rect 5350 -437 5444 -434
rect 5350 -444 5399 -437
rect 5350 -450 5380 -444
rect 5399 -449 5404 -444
rect 5316 -466 5396 -450
rect 5408 -458 5444 -437
rect 5505 -442 5694 -418
rect 5739 -419 5786 -418
rect 5752 -424 5786 -419
rect 5520 -445 5694 -442
rect 5513 -448 5694 -445
rect 5722 -425 5786 -424
rect 5316 -468 5335 -466
rect 5350 -468 5384 -466
rect 5316 -484 5396 -468
rect 5316 -490 5335 -484
rect 5032 -516 5135 -506
rect 4986 -518 5135 -516
rect 5156 -518 5191 -506
rect 4825 -520 4987 -518
rect 4837 -540 4856 -520
rect 4871 -522 4901 -520
rect 4720 -548 4761 -540
rect 4843 -544 4856 -540
rect 4908 -536 4987 -520
rect 5019 -520 5191 -518
rect 5019 -536 5098 -520
rect 5105 -522 5135 -520
rect 4683 -558 4712 -548
rect 4726 -558 4755 -548
rect 4770 -558 4800 -544
rect 4843 -558 4886 -544
rect 4908 -548 5098 -536
rect 5163 -540 5169 -520
rect 4893 -558 4923 -548
rect 4924 -558 5082 -548
rect 5086 -558 5116 -548
rect 5120 -558 5150 -544
rect 5178 -558 5191 -520
rect 5263 -506 5292 -490
rect 5306 -506 5335 -490
rect 5350 -500 5380 -484
rect 5408 -506 5414 -458
rect 5417 -464 5436 -458
rect 5451 -464 5481 -456
rect 5417 -472 5481 -464
rect 5417 -488 5497 -472
rect 5513 -479 5575 -448
rect 5591 -479 5653 -448
rect 5722 -450 5771 -425
rect 5786 -450 5816 -432
rect 5685 -464 5715 -456
rect 5722 -458 5832 -450
rect 5685 -472 5730 -464
rect 5417 -490 5436 -488
rect 5451 -490 5497 -488
rect 5417 -506 5497 -490
rect 5524 -492 5559 -479
rect 5600 -482 5637 -479
rect 5600 -484 5642 -482
rect 5529 -495 5559 -492
rect 5538 -499 5545 -495
rect 5545 -500 5546 -499
rect 5504 -506 5514 -500
rect 5263 -514 5298 -506
rect 5263 -540 5264 -514
rect 5271 -540 5298 -514
rect 5206 -558 5236 -544
rect 5263 -548 5298 -540
rect 5300 -514 5341 -506
rect 5300 -540 5315 -514
rect 5322 -540 5341 -514
rect 5405 -518 5436 -506
rect 5451 -518 5554 -506
rect 5566 -516 5592 -490
rect 5607 -495 5637 -484
rect 5669 -488 5731 -472
rect 5669 -490 5715 -488
rect 5669 -506 5731 -490
rect 5743 -506 5749 -458
rect 5752 -466 5832 -458
rect 5752 -468 5771 -466
rect 5786 -468 5820 -466
rect 5752 -483 5832 -468
rect 5752 -484 5838 -483
rect 5752 -506 5771 -484
rect 5786 -500 5816 -484
rect 5844 -490 5850 -416
rect 5853 -490 5872 -346
rect 5887 -490 5893 -346
rect 5902 -416 5915 -346
rect 5967 -350 5989 -346
rect 5960 -362 5977 -358
rect 5981 -360 5989 -358
rect 5979 -362 5989 -360
rect 5960 -372 5989 -362
rect 6042 -372 6058 -358
rect 6096 -362 6102 -360
rect 6109 -362 6217 -346
rect 6224 -362 6230 -360
rect 6238 -362 6253 -346
rect 6319 -352 6338 -349
rect 5960 -374 6058 -372
rect 6085 -374 6253 -362
rect 6268 -372 6284 -358
rect 6319 -371 6341 -352
rect 6351 -358 6367 -357
rect 6350 -360 6367 -358
rect 6351 -365 6367 -360
rect 6341 -372 6347 -371
rect 6350 -372 6379 -365
rect 6268 -373 6379 -372
rect 6268 -374 6385 -373
rect 5944 -382 5995 -374
rect 6042 -382 6076 -374
rect 5944 -394 5969 -382
rect 5976 -394 5995 -382
rect 6049 -384 6076 -382
rect 6085 -384 6306 -374
rect 6341 -377 6347 -374
rect 6049 -388 6306 -384
rect 5944 -402 5995 -394
rect 6042 -402 6306 -388
rect 6350 -382 6385 -374
rect 5896 -450 5915 -416
rect 5960 -410 5989 -402
rect 5960 -416 5977 -410
rect 5960 -418 5994 -416
rect 6042 -418 6058 -402
rect 6059 -412 6267 -402
rect 6268 -412 6284 -402
rect 6332 -406 6347 -391
rect 6350 -394 6351 -382
rect 6358 -394 6385 -382
rect 6350 -402 6385 -394
rect 6350 -403 6379 -402
rect 6070 -416 6284 -412
rect 6085 -418 6284 -416
rect 6319 -416 6332 -406
rect 6350 -416 6367 -403
rect 6319 -418 6367 -416
rect 5961 -422 5994 -418
rect 5957 -424 5994 -422
rect 5957 -425 6024 -424
rect 5957 -430 5988 -425
rect 5994 -430 6024 -425
rect 5957 -434 6024 -430
rect 5930 -437 6024 -434
rect 5930 -444 5979 -437
rect 5930 -450 5960 -444
rect 5979 -449 5984 -444
rect 5896 -466 5976 -450
rect 5988 -458 6024 -437
rect 6085 -442 6274 -418
rect 6319 -419 6366 -418
rect 6332 -424 6366 -419
rect 6100 -445 6274 -442
rect 6093 -448 6274 -445
rect 6302 -425 6366 -424
rect 5896 -468 5915 -466
rect 5930 -468 5964 -466
rect 5896 -484 5976 -468
rect 5896 -490 5915 -484
rect 5612 -516 5715 -506
rect 5566 -518 5715 -516
rect 5736 -518 5771 -506
rect 5405 -520 5567 -518
rect 5417 -540 5436 -520
rect 5451 -522 5481 -520
rect 5300 -548 5341 -540
rect 5423 -544 5436 -540
rect 5488 -536 5567 -520
rect 5599 -520 5771 -518
rect 5599 -536 5678 -520
rect 5685 -522 5715 -520
rect 5263 -558 5292 -548
rect 5306 -558 5335 -548
rect 5350 -558 5380 -544
rect 5423 -558 5466 -544
rect 5488 -548 5678 -536
rect 5743 -540 5749 -520
rect 5473 -558 5503 -548
rect 5504 -558 5662 -548
rect 5666 -558 5696 -548
rect 5700 -558 5730 -544
rect 5758 -558 5771 -520
rect 5843 -506 5872 -490
rect 5886 -506 5915 -490
rect 5930 -500 5960 -484
rect 5988 -506 5994 -458
rect 5997 -464 6016 -458
rect 6031 -464 6061 -456
rect 5997 -472 6061 -464
rect 5997 -488 6077 -472
rect 6093 -479 6155 -448
rect 6171 -479 6233 -448
rect 6302 -450 6351 -425
rect 6366 -450 6396 -434
rect 6265 -464 6295 -456
rect 6302 -458 6412 -450
rect 6265 -472 6310 -464
rect 5997 -490 6016 -488
rect 6031 -490 6077 -488
rect 5997 -506 6077 -490
rect 6104 -492 6139 -479
rect 6180 -482 6217 -479
rect 6180 -484 6222 -482
rect 6109 -495 6139 -492
rect 6118 -499 6125 -495
rect 6125 -500 6126 -499
rect 6084 -506 6094 -500
rect 5843 -514 5878 -506
rect 5843 -540 5844 -514
rect 5851 -540 5878 -514
rect 5786 -558 5816 -544
rect 5843 -548 5878 -540
rect 5880 -514 5921 -506
rect 5880 -540 5895 -514
rect 5902 -540 5921 -514
rect 5985 -518 6016 -506
rect 6031 -518 6134 -506
rect 6146 -516 6172 -490
rect 6187 -495 6217 -484
rect 6249 -488 6311 -472
rect 6249 -490 6295 -488
rect 6249 -506 6311 -490
rect 6323 -506 6329 -458
rect 6332 -466 6412 -458
rect 6332 -468 6351 -466
rect 6366 -468 6400 -466
rect 6332 -484 6412 -468
rect 6332 -506 6351 -484
rect 6366 -500 6396 -484
rect 6424 -490 6430 -416
rect 6439 -490 6452 -346
rect 6192 -516 6295 -506
rect 6146 -518 6295 -516
rect 6316 -518 6351 -506
rect 5985 -520 6147 -518
rect 5997 -540 6016 -520
rect 6031 -522 6061 -520
rect 5880 -548 5921 -540
rect 6003 -544 6016 -540
rect 6068 -536 6147 -520
rect 6179 -520 6351 -518
rect 6179 -536 6258 -520
rect 6265 -522 6295 -520
rect 5843 -558 5872 -548
rect 5886 -558 5915 -548
rect 5930 -558 5960 -544
rect 6003 -558 6046 -544
rect 6068 -548 6258 -536
rect 6323 -540 6329 -520
rect 6053 -558 6083 -548
rect 6084 -558 6242 -548
rect 6246 -558 6276 -548
rect 6280 -558 6310 -544
rect 6338 -558 6351 -520
rect 6423 -506 6452 -490
rect 6423 -514 6458 -506
rect 6423 -540 6424 -514
rect 6431 -540 6458 -514
rect 6366 -558 6396 -544
rect 6423 -548 6458 -540
rect 6423 -558 6452 -548
rect -541 -572 6452 -558
rect -478 -602 -465 -572
rect -450 -586 -420 -572
rect -377 -586 -334 -572
rect -327 -586 -107 -572
rect -100 -586 -70 -572
rect -410 -600 -395 -588
rect -376 -600 -363 -586
rect -295 -590 -142 -586
rect -413 -602 -391 -600
rect -313 -602 -121 -590
rect -42 -602 -29 -572
rect -14 -586 16 -572
rect 53 -602 72 -572
rect 87 -602 93 -572
rect 102 -602 115 -572
rect 130 -586 160 -572
rect 203 -586 246 -572
rect 253 -586 473 -572
rect 480 -586 510 -572
rect 170 -600 185 -588
rect 204 -600 217 -586
rect 285 -590 438 -586
rect 167 -602 189 -600
rect 267 -602 459 -590
rect 538 -602 551 -572
rect 566 -586 596 -572
rect 633 -602 652 -572
rect 667 -602 673 -572
rect 682 -602 695 -572
rect 710 -586 740 -572
rect 783 -586 826 -572
rect 833 -586 1053 -572
rect 1060 -586 1090 -572
rect 750 -600 765 -588
rect 784 -600 797 -586
rect 865 -590 1018 -586
rect 747 -602 769 -600
rect 847 -602 1039 -590
rect 1118 -602 1131 -572
rect 1146 -586 1176 -572
rect 1213 -602 1232 -572
rect 1247 -602 1253 -572
rect 1262 -602 1275 -572
rect 1290 -586 1320 -572
rect 1363 -586 1406 -572
rect 1413 -586 1633 -572
rect 1640 -586 1670 -572
rect 1330 -600 1345 -588
rect 1364 -600 1377 -586
rect 1445 -590 1598 -586
rect 1327 -602 1349 -600
rect 1427 -602 1619 -590
rect 1698 -602 1711 -572
rect 1726 -586 1756 -572
rect 1793 -602 1812 -572
rect 1827 -602 1833 -572
rect 1842 -602 1855 -572
rect 1870 -586 1900 -572
rect 1943 -586 1986 -572
rect 1993 -586 2213 -572
rect 2220 -586 2250 -572
rect 1910 -600 1925 -588
rect 1944 -600 1957 -586
rect 2025 -590 2178 -586
rect 1907 -602 1929 -600
rect 2007 -602 2199 -590
rect 2278 -602 2291 -572
rect 2306 -586 2336 -572
rect 2373 -602 2392 -572
rect 2407 -602 2413 -572
rect 2422 -602 2435 -572
rect 2450 -586 2480 -572
rect 2523 -586 2566 -572
rect 2573 -586 2793 -572
rect 2800 -586 2830 -572
rect 2490 -600 2505 -588
rect 2524 -600 2537 -586
rect 2605 -590 2758 -586
rect 2487 -602 2509 -600
rect 2587 -602 2779 -590
rect 2858 -602 2871 -572
rect 2886 -586 2916 -572
rect 2953 -602 2972 -572
rect 2987 -602 2993 -572
rect 3002 -602 3015 -572
rect 3030 -586 3060 -572
rect 3103 -586 3146 -572
rect 3153 -586 3373 -572
rect 3380 -586 3410 -572
rect 3070 -600 3085 -588
rect 3104 -600 3117 -586
rect 3185 -590 3338 -586
rect 3067 -602 3089 -600
rect 3167 -602 3359 -590
rect 3438 -602 3451 -572
rect 3466 -586 3496 -572
rect 3533 -602 3552 -572
rect 3567 -602 3573 -572
rect 3582 -602 3595 -572
rect 3610 -586 3640 -572
rect 3683 -586 3726 -572
rect 3733 -586 3953 -572
rect 3960 -586 3990 -572
rect 3650 -600 3665 -588
rect 3684 -600 3697 -586
rect 3765 -590 3918 -586
rect 3647 -602 3669 -600
rect 3747 -602 3939 -590
rect 4018 -602 4031 -572
rect 4046 -586 4076 -572
rect 4113 -602 4132 -572
rect 4147 -602 4153 -572
rect 4162 -602 4175 -572
rect 4190 -586 4220 -572
rect 4263 -586 4306 -572
rect 4313 -586 4533 -572
rect 4540 -586 4570 -572
rect 4230 -600 4245 -588
rect 4264 -600 4277 -586
rect 4345 -590 4498 -586
rect 4227 -602 4249 -600
rect 4327 -602 4519 -590
rect 4598 -602 4611 -572
rect 4626 -586 4656 -572
rect 4693 -602 4712 -572
rect 4727 -602 4733 -572
rect 4742 -602 4755 -572
rect 4770 -586 4800 -572
rect 4843 -586 4886 -572
rect 4893 -586 5113 -572
rect 5120 -586 5150 -572
rect 4810 -600 4825 -588
rect 4844 -600 4857 -586
rect 4925 -590 5078 -586
rect 4807 -602 4829 -600
rect 4907 -602 5099 -590
rect 5178 -602 5191 -572
rect 5206 -586 5236 -572
rect 5273 -602 5292 -572
rect 5307 -602 5313 -572
rect 5322 -602 5335 -572
rect 5350 -586 5380 -572
rect 5423 -586 5466 -572
rect 5473 -586 5693 -572
rect 5700 -586 5730 -572
rect 5390 -600 5405 -588
rect 5424 -600 5437 -586
rect 5505 -590 5658 -586
rect 5387 -602 5409 -600
rect 5487 -602 5679 -590
rect 5758 -602 5771 -572
rect 5786 -586 5816 -572
rect 5853 -602 5872 -572
rect 5887 -602 5893 -572
rect 5902 -602 5915 -572
rect 5930 -586 5960 -572
rect 6003 -586 6046 -572
rect 6053 -586 6273 -572
rect 6280 -586 6310 -572
rect 5970 -600 5985 -588
rect 6004 -600 6017 -586
rect 6085 -590 6238 -586
rect 5967 -602 5989 -600
rect 6067 -602 6259 -590
rect 6338 -602 6351 -572
rect 6366 -586 6396 -572
rect 6439 -602 6452 -572
rect -541 -616 6452 -602
rect -478 -686 -465 -616
rect -413 -620 -391 -616
rect -420 -632 -403 -628
rect -399 -630 -391 -628
rect -401 -632 -391 -630
rect -420 -642 -391 -632
rect -338 -642 -322 -628
rect -284 -632 -278 -630
rect -271 -632 -163 -616
rect -156 -632 -150 -630
rect -142 -632 -127 -616
rect -61 -622 -42 -619
rect -420 -644 -322 -642
rect -295 -644 -127 -632
rect -112 -642 -96 -628
rect -61 -641 -39 -622
rect -29 -628 -13 -627
rect -30 -630 -13 -628
rect -29 -635 -13 -630
rect -39 -642 -33 -641
rect -30 -642 -1 -635
rect -112 -643 -1 -642
rect -112 -644 5 -643
rect -436 -652 -385 -644
rect -338 -652 -304 -644
rect -436 -664 -411 -652
rect -404 -664 -385 -652
rect -331 -654 -304 -652
rect -295 -654 -74 -644
rect -39 -647 -33 -644
rect -331 -658 -74 -654
rect -436 -672 -385 -664
rect -338 -672 -74 -658
rect -30 -652 5 -644
rect -484 -720 -465 -686
rect -420 -680 -391 -672
rect -420 -686 -403 -680
rect -420 -688 -386 -686
rect -338 -688 -322 -672
rect -321 -682 -113 -672
rect -112 -682 -96 -672
rect -48 -676 -33 -661
rect -30 -664 -29 -652
rect -22 -664 5 -652
rect -30 -672 5 -664
rect -30 -673 -1 -672
rect -310 -686 -96 -682
rect -295 -688 -96 -686
rect -61 -686 -48 -676
rect -30 -686 -13 -673
rect -61 -688 -13 -686
rect -419 -692 -386 -688
rect -423 -694 -386 -692
rect -423 -695 -356 -694
rect -423 -700 -392 -695
rect -386 -700 -356 -695
rect -423 -704 -356 -700
rect -450 -707 -356 -704
rect -450 -714 -401 -707
rect -450 -720 -420 -714
rect -401 -719 -396 -714
rect -484 -736 -404 -720
rect -392 -728 -356 -707
rect -295 -712 -106 -688
rect -61 -689 -14 -688
rect -48 -694 -14 -689
rect -280 -715 -106 -712
rect -287 -718 -106 -715
rect -78 -695 -14 -694
rect -484 -738 -465 -736
rect -450 -738 -416 -736
rect -484 -754 -404 -738
rect -484 -760 -465 -754
rect -494 -776 -465 -760
rect -450 -770 -420 -754
rect -392 -776 -386 -728
rect -383 -734 -364 -728
rect -349 -734 -319 -726
rect -383 -742 -319 -734
rect -383 -758 -303 -742
rect -287 -749 -225 -718
rect -209 -749 -147 -718
rect -78 -720 -29 -695
rect -14 -720 16 -702
rect -115 -734 -85 -726
rect -78 -728 32 -720
rect -115 -742 -70 -734
rect -383 -760 -364 -758
rect -349 -760 -303 -758
rect -383 -776 -303 -760
rect -276 -762 -241 -749
rect -200 -752 -163 -749
rect -200 -754 -158 -752
rect -271 -765 -241 -762
rect -262 -769 -255 -765
rect -255 -770 -254 -769
rect -296 -776 -286 -770
rect -500 -784 -459 -776
rect -500 -810 -485 -784
rect -478 -810 -459 -784
rect -395 -788 -364 -776
rect -349 -788 -246 -776
rect -234 -786 -208 -760
rect -193 -765 -163 -754
rect -131 -758 -69 -742
rect -131 -760 -85 -758
rect -131 -776 -69 -760
rect -57 -776 -51 -728
rect -48 -736 32 -728
rect -48 -738 -29 -736
rect -14 -738 20 -736
rect -48 -753 32 -738
rect -48 -754 38 -753
rect -48 -776 -29 -754
rect -14 -770 16 -754
rect 44 -760 50 -686
rect 53 -760 72 -616
rect 87 -760 93 -616
rect 102 -686 115 -616
rect 167 -620 189 -616
rect 160 -632 177 -628
rect 181 -630 189 -628
rect 179 -632 189 -630
rect 160 -642 189 -632
rect 242 -642 258 -628
rect 296 -632 302 -630
rect 309 -632 417 -616
rect 424 -632 430 -630
rect 438 -632 453 -616
rect 519 -622 538 -619
rect 160 -644 258 -642
rect 285 -644 453 -632
rect 468 -642 484 -628
rect 519 -641 541 -622
rect 551 -628 567 -627
rect 550 -630 567 -628
rect 551 -635 567 -630
rect 541 -642 547 -641
rect 550 -642 579 -635
rect 468 -643 579 -642
rect 468 -644 585 -643
rect 144 -652 195 -644
rect 242 -652 276 -644
rect 144 -664 169 -652
rect 176 -664 195 -652
rect 249 -654 276 -652
rect 285 -654 506 -644
rect 541 -647 547 -644
rect 249 -658 506 -654
rect 144 -672 195 -664
rect 242 -672 506 -658
rect 550 -652 585 -644
rect 96 -720 115 -686
rect 160 -680 189 -672
rect 160 -686 177 -680
rect 160 -688 194 -686
rect 242 -688 258 -672
rect 259 -682 467 -672
rect 468 -682 484 -672
rect 532 -676 547 -661
rect 550 -664 551 -652
rect 558 -664 585 -652
rect 550 -672 585 -664
rect 550 -673 579 -672
rect 270 -686 484 -682
rect 285 -688 484 -686
rect 519 -686 532 -676
rect 550 -686 567 -673
rect 519 -688 567 -686
rect 161 -692 194 -688
rect 157 -694 194 -692
rect 157 -695 224 -694
rect 157 -700 188 -695
rect 194 -700 224 -695
rect 157 -704 224 -700
rect 130 -707 224 -704
rect 130 -714 179 -707
rect 130 -720 160 -714
rect 179 -719 184 -714
rect 96 -736 176 -720
rect 188 -728 224 -707
rect 285 -712 474 -688
rect 519 -689 566 -688
rect 532 -694 566 -689
rect 606 -694 622 -692
rect 300 -715 474 -712
rect 293 -718 474 -715
rect 502 -695 566 -694
rect 96 -738 115 -736
rect 130 -738 164 -736
rect 96 -754 176 -738
rect 96 -760 115 -754
rect -188 -786 -85 -776
rect -234 -788 -85 -786
rect -64 -788 -29 -776
rect -395 -790 -233 -788
rect -383 -808 -364 -790
rect -349 -792 -319 -790
rect -500 -818 -459 -810
rect -376 -814 -364 -808
rect -312 -808 -233 -790
rect -201 -790 -29 -788
rect -201 -806 -122 -790
rect -115 -792 -85 -790
rect -226 -808 -122 -806
rect -494 -828 -465 -818
rect -450 -828 -420 -814
rect -376 -828 -334 -814
rect -312 -818 -122 -808
rect -57 -810 -51 -790
rect -327 -828 -297 -818
rect -296 -828 -138 -818
rect -134 -828 -104 -818
rect -100 -828 -70 -814
rect -42 -828 -29 -790
rect 43 -776 72 -760
rect 86 -776 115 -760
rect 130 -770 160 -754
rect 188 -776 194 -728
rect 197 -734 216 -728
rect 231 -734 261 -726
rect 197 -742 261 -734
rect 197 -758 277 -742
rect 293 -749 355 -718
rect 371 -749 433 -718
rect 502 -720 551 -695
rect 596 -704 622 -694
rect 566 -720 622 -704
rect 465 -734 495 -726
rect 502 -728 612 -720
rect 465 -742 510 -734
rect 197 -760 216 -758
rect 231 -760 277 -758
rect 197 -776 277 -760
rect 304 -762 339 -749
rect 380 -752 417 -749
rect 380 -754 422 -752
rect 309 -765 339 -762
rect 318 -769 325 -765
rect 325 -770 326 -769
rect 284 -776 294 -770
rect 43 -784 78 -776
rect 43 -810 44 -784
rect 51 -810 78 -784
rect -14 -828 16 -814
rect 43 -818 78 -810
rect 80 -784 121 -776
rect 80 -810 95 -784
rect 102 -810 121 -784
rect 185 -788 216 -776
rect 231 -788 334 -776
rect 346 -786 372 -760
rect 387 -765 417 -754
rect 449 -758 511 -742
rect 449 -760 495 -758
rect 449 -776 511 -760
rect 523 -776 529 -728
rect 532 -736 612 -728
rect 532 -738 551 -736
rect 566 -738 600 -736
rect 532 -754 612 -738
rect 532 -776 551 -754
rect 566 -770 596 -754
rect 624 -760 630 -686
rect 633 -760 652 -616
rect 667 -760 673 -616
rect 682 -686 695 -616
rect 747 -620 769 -616
rect 740 -632 757 -628
rect 761 -630 769 -628
rect 759 -632 769 -630
rect 740 -642 769 -632
rect 822 -642 838 -628
rect 876 -632 882 -630
rect 889 -632 997 -616
rect 1004 -632 1010 -630
rect 1018 -632 1033 -616
rect 1099 -622 1118 -619
rect 740 -644 838 -642
rect 865 -644 1033 -632
rect 1048 -642 1064 -628
rect 1099 -641 1121 -622
rect 1131 -628 1147 -627
rect 1130 -630 1147 -628
rect 1131 -635 1147 -630
rect 1121 -642 1127 -641
rect 1130 -642 1159 -635
rect 1048 -643 1159 -642
rect 1048 -644 1165 -643
rect 724 -652 775 -644
rect 822 -652 856 -644
rect 724 -664 749 -652
rect 756 -664 775 -652
rect 829 -654 856 -652
rect 865 -654 1086 -644
rect 1121 -647 1127 -644
rect 829 -658 1086 -654
rect 724 -672 775 -664
rect 822 -672 1086 -658
rect 1130 -652 1165 -644
rect 676 -720 695 -686
rect 740 -680 769 -672
rect 740 -686 757 -680
rect 740 -688 774 -686
rect 822 -688 838 -672
rect 839 -682 1047 -672
rect 1048 -682 1064 -672
rect 1112 -676 1127 -661
rect 1130 -664 1131 -652
rect 1138 -664 1165 -652
rect 1130 -672 1165 -664
rect 1130 -673 1159 -672
rect 850 -686 1064 -682
rect 865 -688 1064 -686
rect 1099 -686 1112 -676
rect 1130 -686 1147 -673
rect 1099 -688 1147 -686
rect 741 -692 774 -688
rect 737 -694 774 -692
rect 737 -695 804 -694
rect 737 -700 768 -695
rect 774 -700 804 -695
rect 737 -704 804 -700
rect 710 -707 804 -704
rect 710 -714 759 -707
rect 710 -720 740 -714
rect 759 -719 764 -714
rect 676 -736 756 -720
rect 768 -728 804 -707
rect 865 -712 1054 -688
rect 1099 -689 1146 -688
rect 1112 -694 1146 -689
rect 880 -715 1054 -712
rect 873 -718 1054 -715
rect 1082 -695 1146 -694
rect 676 -738 695 -736
rect 710 -738 744 -736
rect 676 -754 756 -738
rect 676 -760 695 -754
rect 392 -786 495 -776
rect 346 -788 495 -786
rect 516 -788 551 -776
rect 185 -790 347 -788
rect 197 -808 216 -790
rect 231 -792 261 -790
rect 80 -818 121 -810
rect 204 -814 216 -808
rect 268 -808 347 -790
rect 379 -790 551 -788
rect 379 -806 458 -790
rect 465 -792 495 -790
rect 354 -808 458 -806
rect 43 -828 72 -818
rect 86 -828 115 -818
rect 130 -828 160 -814
rect 204 -828 246 -814
rect 268 -818 458 -808
rect 523 -810 529 -790
rect 253 -828 283 -818
rect 284 -828 442 -818
rect 446 -828 476 -818
rect 480 -828 510 -814
rect 538 -828 551 -790
rect 623 -776 652 -760
rect 666 -776 695 -760
rect 710 -770 740 -754
rect 768 -776 774 -728
rect 777 -734 796 -728
rect 811 -734 841 -726
rect 777 -742 841 -734
rect 777 -758 857 -742
rect 873 -749 935 -718
rect 951 -749 1013 -718
rect 1082 -720 1131 -695
rect 1146 -720 1176 -702
rect 1045 -734 1075 -726
rect 1082 -728 1192 -720
rect 1045 -742 1090 -734
rect 777 -760 796 -758
rect 811 -760 857 -758
rect 777 -776 857 -760
rect 884 -762 919 -749
rect 960 -752 997 -749
rect 960 -754 1002 -752
rect 889 -765 919 -762
rect 898 -769 905 -765
rect 905 -770 906 -769
rect 864 -776 874 -770
rect 623 -784 658 -776
rect 623 -810 624 -784
rect 631 -810 658 -784
rect 566 -828 596 -814
rect 623 -818 658 -810
rect 660 -784 701 -776
rect 660 -810 675 -784
rect 682 -810 701 -784
rect 765 -788 796 -776
rect 811 -788 914 -776
rect 926 -786 952 -760
rect 967 -765 997 -754
rect 1029 -758 1091 -742
rect 1029 -760 1075 -758
rect 1029 -776 1091 -760
rect 1103 -776 1109 -728
rect 1112 -736 1192 -728
rect 1112 -738 1131 -736
rect 1146 -738 1180 -736
rect 1112 -753 1192 -738
rect 1112 -754 1198 -753
rect 1112 -776 1131 -754
rect 1146 -770 1176 -754
rect 1204 -760 1210 -686
rect 1213 -760 1232 -616
rect 1247 -760 1253 -616
rect 1262 -686 1275 -616
rect 1327 -620 1349 -616
rect 1320 -632 1337 -628
rect 1341 -630 1349 -628
rect 1339 -632 1349 -630
rect 1320 -642 1349 -632
rect 1402 -642 1418 -628
rect 1456 -632 1462 -630
rect 1469 -632 1577 -616
rect 1584 -632 1590 -630
rect 1598 -632 1613 -616
rect 1679 -622 1698 -619
rect 1320 -644 1418 -642
rect 1445 -644 1613 -632
rect 1628 -642 1644 -628
rect 1679 -641 1701 -622
rect 1711 -628 1727 -627
rect 1710 -630 1727 -628
rect 1711 -635 1727 -630
rect 1701 -642 1707 -641
rect 1710 -642 1739 -635
rect 1628 -643 1739 -642
rect 1628 -644 1745 -643
rect 1304 -652 1355 -644
rect 1402 -652 1436 -644
rect 1304 -664 1329 -652
rect 1336 -664 1355 -652
rect 1409 -654 1436 -652
rect 1445 -654 1666 -644
rect 1701 -647 1707 -644
rect 1409 -658 1666 -654
rect 1304 -672 1355 -664
rect 1402 -672 1666 -658
rect 1710 -652 1745 -644
rect 1256 -720 1275 -686
rect 1320 -680 1349 -672
rect 1320 -686 1337 -680
rect 1320 -688 1354 -686
rect 1402 -688 1418 -672
rect 1419 -682 1627 -672
rect 1628 -682 1644 -672
rect 1692 -676 1707 -661
rect 1710 -664 1711 -652
rect 1718 -664 1745 -652
rect 1710 -672 1745 -664
rect 1710 -673 1739 -672
rect 1430 -686 1644 -682
rect 1445 -688 1644 -686
rect 1679 -686 1692 -676
rect 1710 -686 1727 -673
rect 1679 -688 1727 -686
rect 1321 -692 1354 -688
rect 1317 -694 1354 -692
rect 1317 -695 1384 -694
rect 1317 -700 1348 -695
rect 1354 -700 1384 -695
rect 1317 -704 1384 -700
rect 1290 -707 1384 -704
rect 1290 -714 1339 -707
rect 1290 -720 1320 -714
rect 1339 -719 1344 -714
rect 1256 -736 1336 -720
rect 1348 -728 1384 -707
rect 1445 -712 1634 -688
rect 1679 -689 1726 -688
rect 1692 -694 1726 -689
rect 1766 -694 1782 -692
rect 1460 -715 1634 -712
rect 1453 -718 1634 -715
rect 1662 -695 1726 -694
rect 1256 -738 1275 -736
rect 1290 -738 1324 -736
rect 1256 -754 1336 -738
rect 1256 -760 1275 -754
rect 972 -786 1075 -776
rect 926 -788 1075 -786
rect 1096 -788 1131 -776
rect 765 -790 927 -788
rect 777 -808 796 -790
rect 811 -792 841 -790
rect 660 -818 701 -810
rect 784 -814 796 -808
rect 848 -808 927 -790
rect 959 -790 1131 -788
rect 959 -806 1038 -790
rect 1045 -792 1075 -790
rect 934 -808 1038 -806
rect 623 -828 652 -818
rect 666 -828 695 -818
rect 710 -828 740 -814
rect 784 -828 826 -814
rect 848 -818 1038 -808
rect 1103 -810 1109 -790
rect 833 -828 863 -818
rect 864 -828 1022 -818
rect 1026 -828 1056 -818
rect 1060 -828 1090 -814
rect 1118 -828 1131 -790
rect 1203 -776 1232 -760
rect 1246 -776 1275 -760
rect 1290 -770 1320 -754
rect 1348 -776 1354 -728
rect 1357 -734 1376 -728
rect 1391 -734 1421 -726
rect 1357 -742 1421 -734
rect 1357 -758 1437 -742
rect 1453 -749 1515 -718
rect 1531 -749 1593 -718
rect 1662 -720 1711 -695
rect 1756 -704 1782 -694
rect 1726 -720 1782 -704
rect 1625 -734 1655 -726
rect 1662 -728 1772 -720
rect 1625 -742 1670 -734
rect 1357 -760 1376 -758
rect 1391 -760 1437 -758
rect 1357 -776 1437 -760
rect 1464 -762 1499 -749
rect 1540 -752 1577 -749
rect 1540 -754 1582 -752
rect 1469 -765 1499 -762
rect 1478 -769 1485 -765
rect 1485 -770 1486 -769
rect 1444 -776 1454 -770
rect 1203 -784 1238 -776
rect 1203 -810 1204 -784
rect 1211 -810 1238 -784
rect 1146 -828 1176 -814
rect 1203 -818 1238 -810
rect 1240 -784 1281 -776
rect 1240 -810 1255 -784
rect 1262 -810 1281 -784
rect 1345 -788 1376 -776
rect 1391 -788 1494 -776
rect 1506 -786 1532 -760
rect 1547 -765 1577 -754
rect 1609 -758 1671 -742
rect 1609 -760 1655 -758
rect 1609 -776 1671 -760
rect 1683 -776 1689 -728
rect 1692 -736 1772 -728
rect 1692 -738 1711 -736
rect 1726 -738 1760 -736
rect 1692 -754 1772 -738
rect 1692 -776 1711 -754
rect 1726 -770 1756 -754
rect 1784 -760 1790 -686
rect 1793 -760 1812 -616
rect 1827 -760 1833 -616
rect 1842 -686 1855 -616
rect 1907 -620 1929 -616
rect 1900 -632 1917 -628
rect 1921 -630 1929 -628
rect 1919 -632 1929 -630
rect 1900 -642 1929 -632
rect 1982 -642 1998 -628
rect 2036 -632 2042 -630
rect 2049 -632 2157 -616
rect 2164 -632 2170 -630
rect 2178 -632 2193 -616
rect 2259 -622 2278 -619
rect 1900 -644 1998 -642
rect 2025 -644 2193 -632
rect 2208 -642 2224 -628
rect 2259 -641 2281 -622
rect 2291 -628 2307 -627
rect 2290 -630 2307 -628
rect 2291 -635 2307 -630
rect 2281 -642 2287 -641
rect 2290 -642 2319 -635
rect 2208 -643 2319 -642
rect 2208 -644 2325 -643
rect 1884 -652 1935 -644
rect 1982 -652 2016 -644
rect 1884 -664 1909 -652
rect 1916 -664 1935 -652
rect 1989 -654 2016 -652
rect 2025 -654 2246 -644
rect 2281 -647 2287 -644
rect 1989 -658 2246 -654
rect 1884 -672 1935 -664
rect 1982 -672 2246 -658
rect 2290 -652 2325 -644
rect 1836 -720 1855 -686
rect 1900 -680 1929 -672
rect 1900 -686 1917 -680
rect 1900 -688 1934 -686
rect 1982 -688 1998 -672
rect 1999 -682 2207 -672
rect 2208 -682 2224 -672
rect 2272 -676 2287 -661
rect 2290 -664 2291 -652
rect 2298 -664 2325 -652
rect 2290 -672 2325 -664
rect 2290 -673 2319 -672
rect 2010 -686 2224 -682
rect 2025 -688 2224 -686
rect 2259 -686 2272 -676
rect 2290 -686 2307 -673
rect 2259 -688 2307 -686
rect 1901 -692 1934 -688
rect 1897 -694 1934 -692
rect 1897 -695 1964 -694
rect 1897 -700 1928 -695
rect 1934 -700 1964 -695
rect 1897 -704 1964 -700
rect 1870 -707 1964 -704
rect 1870 -714 1919 -707
rect 1870 -720 1900 -714
rect 1919 -719 1924 -714
rect 1836 -736 1916 -720
rect 1928 -728 1964 -707
rect 2025 -712 2214 -688
rect 2259 -689 2306 -688
rect 2272 -694 2306 -689
rect 2040 -715 2214 -712
rect 2033 -718 2214 -715
rect 2242 -695 2306 -694
rect 1836 -738 1855 -736
rect 1870 -738 1904 -736
rect 1836 -754 1916 -738
rect 1836 -760 1855 -754
rect 1552 -786 1655 -776
rect 1506 -788 1655 -786
rect 1676 -788 1711 -776
rect 1345 -790 1507 -788
rect 1357 -808 1376 -790
rect 1391 -792 1421 -790
rect 1240 -818 1281 -810
rect 1364 -814 1376 -808
rect 1428 -808 1507 -790
rect 1539 -790 1711 -788
rect 1539 -806 1618 -790
rect 1625 -792 1655 -790
rect 1514 -808 1618 -806
rect 1203 -828 1232 -818
rect 1246 -828 1275 -818
rect 1290 -828 1320 -814
rect 1364 -828 1406 -814
rect 1428 -818 1618 -808
rect 1683 -810 1689 -790
rect 1413 -828 1443 -818
rect 1444 -828 1602 -818
rect 1606 -828 1636 -818
rect 1640 -828 1670 -814
rect 1698 -828 1711 -790
rect 1783 -776 1812 -760
rect 1826 -776 1855 -760
rect 1870 -770 1900 -754
rect 1928 -776 1934 -728
rect 1937 -734 1956 -728
rect 1971 -734 2001 -726
rect 1937 -742 2001 -734
rect 1937 -758 2017 -742
rect 2033 -749 2095 -718
rect 2111 -749 2173 -718
rect 2242 -720 2291 -695
rect 2306 -720 2336 -702
rect 2205 -734 2235 -726
rect 2242 -728 2352 -720
rect 2205 -742 2250 -734
rect 1937 -760 1956 -758
rect 1971 -760 2017 -758
rect 1937 -776 2017 -760
rect 2044 -762 2079 -749
rect 2120 -752 2157 -749
rect 2120 -754 2162 -752
rect 2049 -765 2079 -762
rect 2058 -769 2065 -765
rect 2065 -770 2066 -769
rect 2024 -776 2034 -770
rect 1783 -784 1818 -776
rect 1783 -810 1784 -784
rect 1791 -810 1818 -784
rect 1726 -828 1756 -814
rect 1783 -818 1818 -810
rect 1820 -784 1861 -776
rect 1820 -810 1835 -784
rect 1842 -810 1861 -784
rect 1925 -788 1956 -776
rect 1971 -788 2074 -776
rect 2086 -786 2112 -760
rect 2127 -765 2157 -754
rect 2189 -758 2251 -742
rect 2189 -760 2235 -758
rect 2189 -776 2251 -760
rect 2263 -776 2269 -728
rect 2272 -736 2352 -728
rect 2272 -738 2291 -736
rect 2306 -738 2340 -736
rect 2272 -753 2352 -738
rect 2272 -754 2358 -753
rect 2272 -776 2291 -754
rect 2306 -770 2336 -754
rect 2364 -760 2370 -686
rect 2373 -760 2392 -616
rect 2407 -760 2413 -616
rect 2422 -686 2435 -616
rect 2487 -620 2509 -616
rect 2480 -632 2497 -628
rect 2501 -630 2509 -628
rect 2499 -632 2509 -630
rect 2480 -642 2509 -632
rect 2562 -642 2578 -628
rect 2616 -632 2622 -630
rect 2629 -632 2737 -616
rect 2744 -632 2750 -630
rect 2758 -632 2773 -616
rect 2839 -622 2858 -619
rect 2480 -644 2578 -642
rect 2605 -644 2773 -632
rect 2788 -642 2804 -628
rect 2839 -641 2861 -622
rect 2871 -628 2887 -627
rect 2870 -630 2887 -628
rect 2871 -635 2887 -630
rect 2861 -642 2867 -641
rect 2870 -642 2899 -635
rect 2788 -643 2899 -642
rect 2788 -644 2905 -643
rect 2464 -652 2515 -644
rect 2562 -652 2596 -644
rect 2464 -664 2489 -652
rect 2496 -664 2515 -652
rect 2569 -654 2596 -652
rect 2605 -654 2826 -644
rect 2861 -647 2867 -644
rect 2569 -658 2826 -654
rect 2464 -672 2515 -664
rect 2562 -672 2826 -658
rect 2870 -652 2905 -644
rect 2416 -720 2435 -686
rect 2480 -680 2509 -672
rect 2480 -686 2497 -680
rect 2480 -688 2514 -686
rect 2562 -688 2578 -672
rect 2579 -682 2787 -672
rect 2788 -682 2804 -672
rect 2852 -676 2867 -661
rect 2870 -664 2871 -652
rect 2878 -664 2905 -652
rect 2870 -672 2905 -664
rect 2870 -673 2899 -672
rect 2590 -686 2804 -682
rect 2605 -688 2804 -686
rect 2839 -686 2852 -676
rect 2870 -686 2887 -673
rect 2839 -688 2887 -686
rect 2481 -692 2514 -688
rect 2477 -694 2514 -692
rect 2477 -695 2544 -694
rect 2477 -700 2508 -695
rect 2514 -700 2544 -695
rect 2477 -704 2544 -700
rect 2450 -707 2544 -704
rect 2450 -714 2499 -707
rect 2450 -720 2480 -714
rect 2499 -719 2504 -714
rect 2416 -736 2496 -720
rect 2508 -728 2544 -707
rect 2605 -712 2794 -688
rect 2839 -689 2886 -688
rect 2852 -694 2886 -689
rect 2926 -694 2942 -692
rect 2620 -715 2794 -712
rect 2613 -718 2794 -715
rect 2822 -695 2886 -694
rect 2416 -738 2435 -736
rect 2450 -738 2484 -736
rect 2416 -754 2496 -738
rect 2416 -760 2435 -754
rect 2132 -786 2235 -776
rect 2086 -788 2235 -786
rect 2256 -788 2291 -776
rect 1925 -790 2087 -788
rect 1937 -808 1956 -790
rect 1971 -792 2001 -790
rect 1820 -818 1861 -810
rect 1944 -814 1956 -808
rect 2008 -808 2087 -790
rect 2119 -790 2291 -788
rect 2119 -806 2198 -790
rect 2205 -792 2235 -790
rect 2094 -808 2198 -806
rect 1783 -828 1812 -818
rect 1826 -828 1855 -818
rect 1870 -828 1900 -814
rect 1944 -828 1986 -814
rect 2008 -818 2198 -808
rect 2263 -810 2269 -790
rect 1993 -828 2023 -818
rect 2024 -828 2182 -818
rect 2186 -828 2216 -818
rect 2220 -828 2250 -814
rect 2278 -828 2291 -790
rect 2363 -776 2392 -760
rect 2406 -776 2435 -760
rect 2450 -770 2480 -754
rect 2508 -776 2514 -728
rect 2517 -734 2536 -728
rect 2551 -734 2581 -726
rect 2517 -742 2581 -734
rect 2517 -758 2597 -742
rect 2613 -749 2675 -718
rect 2691 -749 2753 -718
rect 2822 -720 2871 -695
rect 2916 -704 2942 -694
rect 2886 -720 2942 -704
rect 2785 -734 2815 -726
rect 2822 -728 2932 -720
rect 2785 -742 2830 -734
rect 2517 -760 2536 -758
rect 2551 -760 2597 -758
rect 2517 -776 2597 -760
rect 2624 -762 2659 -749
rect 2700 -752 2737 -749
rect 2700 -754 2742 -752
rect 2629 -765 2659 -762
rect 2638 -769 2645 -765
rect 2645 -770 2646 -769
rect 2604 -776 2614 -770
rect 2363 -784 2398 -776
rect 2363 -810 2364 -784
rect 2371 -810 2398 -784
rect 2306 -828 2336 -814
rect 2363 -818 2398 -810
rect 2400 -784 2441 -776
rect 2400 -810 2415 -784
rect 2422 -810 2441 -784
rect 2505 -788 2536 -776
rect 2551 -788 2654 -776
rect 2666 -786 2692 -760
rect 2707 -765 2737 -754
rect 2769 -758 2831 -742
rect 2769 -760 2815 -758
rect 2769 -776 2831 -760
rect 2843 -776 2849 -728
rect 2852 -736 2932 -728
rect 2852 -738 2871 -736
rect 2886 -738 2920 -736
rect 2852 -754 2932 -738
rect 2852 -776 2871 -754
rect 2886 -770 2916 -754
rect 2944 -760 2950 -686
rect 2953 -760 2972 -616
rect 2987 -760 2993 -616
rect 3002 -686 3015 -616
rect 3067 -620 3089 -616
rect 3060 -632 3077 -628
rect 3081 -630 3089 -628
rect 3079 -632 3089 -630
rect 3060 -642 3089 -632
rect 3142 -642 3158 -628
rect 3196 -632 3202 -630
rect 3209 -632 3317 -616
rect 3324 -632 3330 -630
rect 3338 -632 3353 -616
rect 3419 -622 3438 -619
rect 3060 -644 3158 -642
rect 3185 -644 3353 -632
rect 3368 -642 3384 -628
rect 3419 -641 3441 -622
rect 3451 -628 3467 -627
rect 3450 -630 3467 -628
rect 3451 -635 3467 -630
rect 3441 -642 3447 -641
rect 3450 -642 3479 -635
rect 3368 -643 3479 -642
rect 3368 -644 3485 -643
rect 3044 -652 3095 -644
rect 3142 -652 3176 -644
rect 3044 -664 3069 -652
rect 3076 -664 3095 -652
rect 3149 -654 3176 -652
rect 3185 -654 3406 -644
rect 3441 -647 3447 -644
rect 3149 -658 3406 -654
rect 3044 -672 3095 -664
rect 3142 -672 3406 -658
rect 3450 -652 3485 -644
rect 2996 -720 3015 -686
rect 3060 -680 3089 -672
rect 3060 -686 3077 -680
rect 3060 -688 3094 -686
rect 3142 -688 3158 -672
rect 3159 -682 3367 -672
rect 3368 -682 3384 -672
rect 3432 -676 3447 -661
rect 3450 -664 3451 -652
rect 3458 -664 3485 -652
rect 3450 -672 3485 -664
rect 3450 -673 3479 -672
rect 3170 -686 3384 -682
rect 3185 -688 3384 -686
rect 3419 -686 3432 -676
rect 3450 -686 3467 -673
rect 3419 -688 3467 -686
rect 3061 -692 3094 -688
rect 3057 -694 3094 -692
rect 3057 -695 3124 -694
rect 3057 -700 3088 -695
rect 3094 -700 3124 -695
rect 3057 -704 3124 -700
rect 3030 -707 3124 -704
rect 3030 -714 3079 -707
rect 3030 -720 3060 -714
rect 3079 -719 3084 -714
rect 2996 -736 3076 -720
rect 3088 -728 3124 -707
rect 3185 -712 3374 -688
rect 3419 -689 3466 -688
rect 3432 -694 3466 -689
rect 3200 -715 3374 -712
rect 3193 -718 3374 -715
rect 3402 -695 3466 -694
rect 2996 -738 3015 -736
rect 3030 -738 3064 -736
rect 2996 -754 3076 -738
rect 2996 -760 3015 -754
rect 2712 -786 2815 -776
rect 2666 -788 2815 -786
rect 2836 -788 2871 -776
rect 2505 -790 2667 -788
rect 2517 -808 2536 -790
rect 2551 -792 2581 -790
rect 2400 -818 2441 -810
rect 2524 -814 2536 -808
rect 2588 -808 2667 -790
rect 2699 -790 2871 -788
rect 2699 -806 2778 -790
rect 2785 -792 2815 -790
rect 2674 -808 2778 -806
rect 2363 -828 2392 -818
rect 2406 -828 2435 -818
rect 2450 -828 2480 -814
rect 2524 -828 2566 -814
rect 2588 -818 2778 -808
rect 2843 -810 2849 -790
rect 2573 -828 2603 -818
rect 2604 -828 2762 -818
rect 2766 -828 2796 -818
rect 2800 -828 2830 -814
rect 2858 -828 2871 -790
rect 2943 -776 2972 -760
rect 2986 -776 3015 -760
rect 3030 -770 3060 -754
rect 3088 -776 3094 -728
rect 3097 -734 3116 -728
rect 3131 -734 3161 -726
rect 3097 -742 3161 -734
rect 3097 -758 3177 -742
rect 3193 -749 3255 -718
rect 3271 -749 3333 -718
rect 3402 -720 3451 -695
rect 3466 -720 3496 -702
rect 3365 -734 3395 -726
rect 3402 -728 3512 -720
rect 3365 -742 3410 -734
rect 3097 -760 3116 -758
rect 3131 -760 3177 -758
rect 3097 -776 3177 -760
rect 3204 -762 3239 -749
rect 3280 -752 3317 -749
rect 3280 -754 3322 -752
rect 3209 -765 3239 -762
rect 3218 -769 3225 -765
rect 3225 -770 3226 -769
rect 3184 -776 3194 -770
rect 2943 -784 2978 -776
rect 2943 -810 2944 -784
rect 2951 -810 2978 -784
rect 2886 -828 2916 -814
rect 2943 -818 2978 -810
rect 2980 -784 3021 -776
rect 2980 -810 2995 -784
rect 3002 -810 3021 -784
rect 3085 -788 3116 -776
rect 3131 -788 3234 -776
rect 3246 -786 3272 -760
rect 3287 -765 3317 -754
rect 3349 -758 3411 -742
rect 3349 -760 3395 -758
rect 3349 -776 3411 -760
rect 3423 -776 3429 -728
rect 3432 -736 3512 -728
rect 3432 -738 3451 -736
rect 3466 -738 3500 -736
rect 3432 -753 3512 -738
rect 3432 -754 3518 -753
rect 3432 -776 3451 -754
rect 3466 -770 3496 -754
rect 3524 -760 3530 -686
rect 3533 -760 3552 -616
rect 3567 -760 3573 -616
rect 3582 -686 3595 -616
rect 3647 -620 3669 -616
rect 3640 -632 3657 -628
rect 3661 -630 3669 -628
rect 3659 -632 3669 -630
rect 3640 -642 3669 -632
rect 3722 -642 3738 -628
rect 3776 -632 3782 -630
rect 3789 -632 3897 -616
rect 3904 -632 3910 -630
rect 3918 -632 3933 -616
rect 3999 -622 4018 -619
rect 3640 -644 3738 -642
rect 3765 -644 3933 -632
rect 3948 -642 3964 -628
rect 3999 -641 4021 -622
rect 4031 -628 4047 -627
rect 4030 -630 4047 -628
rect 4031 -635 4047 -630
rect 4021 -642 4027 -641
rect 4030 -642 4059 -635
rect 3948 -643 4059 -642
rect 3948 -644 4065 -643
rect 3624 -652 3675 -644
rect 3722 -652 3756 -644
rect 3624 -664 3649 -652
rect 3656 -664 3675 -652
rect 3729 -654 3756 -652
rect 3765 -654 3986 -644
rect 4021 -647 4027 -644
rect 3729 -658 3986 -654
rect 3624 -672 3675 -664
rect 3722 -672 3986 -658
rect 4030 -652 4065 -644
rect 3576 -720 3595 -686
rect 3640 -680 3669 -672
rect 3640 -686 3657 -680
rect 3640 -688 3674 -686
rect 3722 -688 3738 -672
rect 3739 -682 3947 -672
rect 3948 -682 3964 -672
rect 4012 -676 4027 -661
rect 4030 -664 4031 -652
rect 4038 -664 4065 -652
rect 4030 -672 4065 -664
rect 4030 -673 4059 -672
rect 3750 -686 3964 -682
rect 3765 -688 3964 -686
rect 3999 -686 4012 -676
rect 4030 -686 4047 -673
rect 3999 -688 4047 -686
rect 3641 -692 3674 -688
rect 3637 -694 3674 -692
rect 3637 -695 3704 -694
rect 3637 -700 3668 -695
rect 3674 -700 3704 -695
rect 3637 -704 3704 -700
rect 3610 -707 3704 -704
rect 3610 -714 3659 -707
rect 3610 -720 3640 -714
rect 3659 -719 3664 -714
rect 3576 -736 3656 -720
rect 3668 -728 3704 -707
rect 3765 -712 3954 -688
rect 3999 -689 4046 -688
rect 4012 -694 4046 -689
rect 4086 -694 4102 -692
rect 3780 -715 3954 -712
rect 3773 -718 3954 -715
rect 3982 -695 4046 -694
rect 3576 -738 3595 -736
rect 3610 -738 3644 -736
rect 3576 -754 3656 -738
rect 3576 -760 3595 -754
rect 3292 -786 3395 -776
rect 3246 -788 3395 -786
rect 3416 -788 3451 -776
rect 3085 -790 3247 -788
rect 3097 -808 3116 -790
rect 3131 -792 3161 -790
rect 2980 -818 3021 -810
rect 3104 -814 3116 -808
rect 3168 -808 3247 -790
rect 3279 -790 3451 -788
rect 3279 -806 3358 -790
rect 3365 -792 3395 -790
rect 3254 -808 3358 -806
rect 2943 -828 2972 -818
rect 2986 -828 3015 -818
rect 3030 -828 3060 -814
rect 3104 -828 3146 -814
rect 3168 -818 3358 -808
rect 3423 -810 3429 -790
rect 3153 -828 3183 -818
rect 3184 -828 3342 -818
rect 3346 -828 3376 -818
rect 3380 -828 3410 -814
rect 3438 -828 3451 -790
rect 3523 -776 3552 -760
rect 3566 -776 3595 -760
rect 3610 -770 3640 -754
rect 3668 -776 3674 -728
rect 3677 -734 3696 -728
rect 3711 -734 3741 -726
rect 3677 -742 3741 -734
rect 3677 -758 3757 -742
rect 3773 -749 3835 -718
rect 3851 -749 3913 -718
rect 3982 -720 4031 -695
rect 4076 -704 4102 -694
rect 4046 -720 4102 -704
rect 3945 -734 3975 -726
rect 3982 -728 4092 -720
rect 3945 -742 3990 -734
rect 3677 -760 3696 -758
rect 3711 -760 3757 -758
rect 3677 -776 3757 -760
rect 3784 -762 3819 -749
rect 3860 -752 3897 -749
rect 3860 -754 3902 -752
rect 3789 -765 3819 -762
rect 3798 -769 3805 -765
rect 3805 -770 3806 -769
rect 3764 -776 3774 -770
rect 3523 -784 3558 -776
rect 3523 -810 3524 -784
rect 3531 -810 3558 -784
rect 3466 -828 3496 -814
rect 3523 -818 3558 -810
rect 3560 -784 3601 -776
rect 3560 -810 3575 -784
rect 3582 -810 3601 -784
rect 3665 -788 3696 -776
rect 3711 -788 3814 -776
rect 3826 -786 3852 -760
rect 3867 -765 3897 -754
rect 3929 -758 3991 -742
rect 3929 -760 3975 -758
rect 3929 -776 3991 -760
rect 4003 -776 4009 -728
rect 4012 -736 4092 -728
rect 4012 -738 4031 -736
rect 4046 -738 4080 -736
rect 4012 -754 4092 -738
rect 4012 -776 4031 -754
rect 4046 -770 4076 -754
rect 4104 -760 4110 -686
rect 4113 -760 4132 -616
rect 4147 -760 4153 -616
rect 4162 -686 4175 -616
rect 4227 -620 4249 -616
rect 4220 -632 4237 -628
rect 4241 -630 4249 -628
rect 4239 -632 4249 -630
rect 4220 -642 4249 -632
rect 4302 -642 4318 -628
rect 4356 -632 4362 -630
rect 4369 -632 4477 -616
rect 4484 -632 4490 -630
rect 4498 -632 4513 -616
rect 4579 -622 4598 -619
rect 4220 -644 4318 -642
rect 4345 -644 4513 -632
rect 4528 -642 4544 -628
rect 4579 -641 4601 -622
rect 4611 -628 4627 -627
rect 4610 -630 4627 -628
rect 4611 -635 4627 -630
rect 4601 -642 4607 -641
rect 4610 -642 4639 -635
rect 4528 -643 4639 -642
rect 4528 -644 4645 -643
rect 4204 -652 4255 -644
rect 4302 -652 4336 -644
rect 4204 -664 4229 -652
rect 4236 -664 4255 -652
rect 4309 -654 4336 -652
rect 4345 -654 4566 -644
rect 4601 -647 4607 -644
rect 4309 -658 4566 -654
rect 4204 -672 4255 -664
rect 4302 -672 4566 -658
rect 4610 -652 4645 -644
rect 4156 -720 4175 -686
rect 4220 -680 4249 -672
rect 4220 -686 4237 -680
rect 4220 -688 4254 -686
rect 4302 -688 4318 -672
rect 4319 -682 4527 -672
rect 4528 -682 4544 -672
rect 4592 -676 4607 -661
rect 4610 -664 4611 -652
rect 4618 -664 4645 -652
rect 4610 -672 4645 -664
rect 4610 -673 4639 -672
rect 4330 -686 4544 -682
rect 4345 -688 4544 -686
rect 4579 -686 4592 -676
rect 4610 -686 4627 -673
rect 4579 -688 4627 -686
rect 4221 -692 4254 -688
rect 4217 -694 4254 -692
rect 4217 -695 4284 -694
rect 4217 -700 4248 -695
rect 4254 -700 4284 -695
rect 4217 -704 4284 -700
rect 4190 -707 4284 -704
rect 4190 -714 4239 -707
rect 4190 -720 4220 -714
rect 4239 -719 4244 -714
rect 4156 -736 4236 -720
rect 4248 -728 4284 -707
rect 4345 -712 4534 -688
rect 4579 -689 4626 -688
rect 4592 -694 4626 -689
rect 4360 -715 4534 -712
rect 4353 -718 4534 -715
rect 4562 -695 4626 -694
rect 4156 -738 4175 -736
rect 4190 -738 4224 -736
rect 4156 -754 4236 -738
rect 4156 -760 4175 -754
rect 3872 -786 3975 -776
rect 3826 -788 3975 -786
rect 3996 -788 4031 -776
rect 3665 -790 3827 -788
rect 3677 -808 3696 -790
rect 3711 -792 3741 -790
rect 3560 -818 3601 -810
rect 3684 -814 3696 -808
rect 3748 -808 3827 -790
rect 3859 -790 4031 -788
rect 3859 -806 3938 -790
rect 3945 -792 3975 -790
rect 3834 -808 3938 -806
rect 3523 -828 3552 -818
rect 3566 -828 3595 -818
rect 3610 -828 3640 -814
rect 3684 -828 3726 -814
rect 3748 -818 3938 -808
rect 4003 -810 4009 -790
rect 3733 -828 3763 -818
rect 3764 -828 3922 -818
rect 3926 -828 3956 -818
rect 3960 -828 3990 -814
rect 4018 -828 4031 -790
rect 4103 -776 4132 -760
rect 4146 -776 4175 -760
rect 4190 -770 4220 -754
rect 4248 -776 4254 -728
rect 4257 -734 4276 -728
rect 4291 -734 4321 -726
rect 4257 -742 4321 -734
rect 4257 -758 4337 -742
rect 4353 -749 4415 -718
rect 4431 -749 4493 -718
rect 4562 -720 4611 -695
rect 4626 -720 4656 -702
rect 4525 -734 4555 -726
rect 4562 -728 4672 -720
rect 4525 -742 4570 -734
rect 4257 -760 4276 -758
rect 4291 -760 4337 -758
rect 4257 -776 4337 -760
rect 4364 -762 4399 -749
rect 4440 -752 4477 -749
rect 4440 -754 4482 -752
rect 4369 -765 4399 -762
rect 4378 -769 4385 -765
rect 4385 -770 4386 -769
rect 4344 -776 4354 -770
rect 4103 -784 4138 -776
rect 4103 -810 4104 -784
rect 4111 -810 4138 -784
rect 4046 -828 4076 -814
rect 4103 -818 4138 -810
rect 4140 -784 4181 -776
rect 4140 -810 4155 -784
rect 4162 -810 4181 -784
rect 4245 -788 4276 -776
rect 4291 -788 4394 -776
rect 4406 -786 4432 -760
rect 4447 -765 4477 -754
rect 4509 -758 4571 -742
rect 4509 -760 4555 -758
rect 4509 -776 4571 -760
rect 4583 -776 4589 -728
rect 4592 -736 4672 -728
rect 4592 -738 4611 -736
rect 4626 -738 4660 -736
rect 4592 -753 4672 -738
rect 4592 -754 4678 -753
rect 4592 -776 4611 -754
rect 4626 -770 4656 -754
rect 4684 -760 4690 -686
rect 4693 -760 4712 -616
rect 4727 -760 4733 -616
rect 4742 -686 4755 -616
rect 4807 -620 4829 -616
rect 4800 -632 4817 -628
rect 4821 -630 4829 -628
rect 4819 -632 4829 -630
rect 4800 -642 4829 -632
rect 4882 -642 4898 -628
rect 4936 -632 4942 -630
rect 4949 -632 5057 -616
rect 5064 -632 5070 -630
rect 5078 -632 5093 -616
rect 5159 -622 5178 -619
rect 4800 -644 4898 -642
rect 4925 -644 5093 -632
rect 5108 -642 5124 -628
rect 5159 -641 5181 -622
rect 5191 -628 5207 -627
rect 5190 -630 5207 -628
rect 5191 -635 5207 -630
rect 5181 -642 5187 -641
rect 5190 -642 5219 -635
rect 5108 -643 5219 -642
rect 5108 -644 5225 -643
rect 4784 -652 4835 -644
rect 4882 -652 4916 -644
rect 4784 -664 4809 -652
rect 4816 -664 4835 -652
rect 4889 -654 4916 -652
rect 4925 -654 5146 -644
rect 5181 -647 5187 -644
rect 4889 -658 5146 -654
rect 4784 -672 4835 -664
rect 4882 -672 5146 -658
rect 5190 -652 5225 -644
rect 4736 -720 4755 -686
rect 4800 -680 4829 -672
rect 4800 -686 4817 -680
rect 4800 -688 4834 -686
rect 4882 -688 4898 -672
rect 4899 -682 5107 -672
rect 5108 -682 5124 -672
rect 5172 -676 5187 -661
rect 5190 -664 5191 -652
rect 5198 -664 5225 -652
rect 5190 -672 5225 -664
rect 5190 -673 5219 -672
rect 4910 -686 5124 -682
rect 4925 -688 5124 -686
rect 5159 -686 5172 -676
rect 5190 -686 5207 -673
rect 5159 -688 5207 -686
rect 4801 -692 4834 -688
rect 4797 -694 4834 -692
rect 4797 -695 4864 -694
rect 4797 -700 4828 -695
rect 4834 -700 4864 -695
rect 4797 -704 4864 -700
rect 4770 -707 4864 -704
rect 4770 -714 4819 -707
rect 4770 -720 4800 -714
rect 4819 -719 4824 -714
rect 4736 -736 4816 -720
rect 4828 -728 4864 -707
rect 4925 -712 5114 -688
rect 5159 -689 5206 -688
rect 5172 -694 5206 -689
rect 5246 -694 5262 -692
rect 4940 -715 5114 -712
rect 4933 -718 5114 -715
rect 5142 -695 5206 -694
rect 4736 -738 4755 -736
rect 4770 -738 4804 -736
rect 4736 -754 4816 -738
rect 4736 -760 4755 -754
rect 4452 -786 4555 -776
rect 4406 -788 4555 -786
rect 4576 -788 4611 -776
rect 4245 -790 4407 -788
rect 4257 -808 4276 -790
rect 4291 -792 4321 -790
rect 4140 -818 4181 -810
rect 4264 -814 4276 -808
rect 4328 -808 4407 -790
rect 4439 -790 4611 -788
rect 4439 -806 4518 -790
rect 4525 -792 4555 -790
rect 4414 -808 4518 -806
rect 4103 -828 4132 -818
rect 4146 -828 4175 -818
rect 4190 -828 4220 -814
rect 4264 -828 4306 -814
rect 4328 -818 4518 -808
rect 4583 -810 4589 -790
rect 4313 -828 4343 -818
rect 4344 -828 4502 -818
rect 4506 -828 4536 -818
rect 4540 -828 4570 -814
rect 4598 -828 4611 -790
rect 4683 -776 4712 -760
rect 4726 -776 4755 -760
rect 4770 -770 4800 -754
rect 4828 -776 4834 -728
rect 4837 -734 4856 -728
rect 4871 -734 4901 -726
rect 4837 -742 4901 -734
rect 4837 -758 4917 -742
rect 4933 -749 4995 -718
rect 5011 -749 5073 -718
rect 5142 -720 5191 -695
rect 5236 -704 5262 -694
rect 5206 -720 5262 -704
rect 5105 -734 5135 -726
rect 5142 -728 5252 -720
rect 5105 -742 5150 -734
rect 4837 -760 4856 -758
rect 4871 -760 4917 -758
rect 4837 -776 4917 -760
rect 4944 -762 4979 -749
rect 5020 -752 5057 -749
rect 5020 -754 5062 -752
rect 4949 -765 4979 -762
rect 4958 -769 4965 -765
rect 4965 -770 4966 -769
rect 4924 -776 4934 -770
rect 4683 -784 4718 -776
rect 4683 -810 4684 -784
rect 4691 -810 4718 -784
rect 4626 -828 4656 -814
rect 4683 -818 4718 -810
rect 4720 -784 4761 -776
rect 4720 -810 4735 -784
rect 4742 -810 4761 -784
rect 4825 -788 4856 -776
rect 4871 -788 4974 -776
rect 4986 -786 5012 -760
rect 5027 -765 5057 -754
rect 5089 -758 5151 -742
rect 5089 -760 5135 -758
rect 5089 -776 5151 -760
rect 5163 -776 5169 -728
rect 5172 -736 5252 -728
rect 5172 -738 5191 -736
rect 5206 -738 5240 -736
rect 5172 -754 5252 -738
rect 5172 -776 5191 -754
rect 5206 -770 5236 -754
rect 5264 -760 5270 -686
rect 5273 -760 5292 -616
rect 5307 -760 5313 -616
rect 5322 -686 5335 -616
rect 5387 -620 5409 -616
rect 5380 -632 5397 -628
rect 5401 -630 5409 -628
rect 5399 -632 5409 -630
rect 5380 -642 5409 -632
rect 5462 -642 5478 -628
rect 5516 -632 5522 -630
rect 5529 -632 5637 -616
rect 5644 -632 5650 -630
rect 5658 -632 5673 -616
rect 5739 -622 5758 -619
rect 5380 -644 5478 -642
rect 5505 -644 5673 -632
rect 5688 -642 5704 -628
rect 5739 -641 5761 -622
rect 5771 -628 5787 -627
rect 5770 -630 5787 -628
rect 5771 -635 5787 -630
rect 5761 -642 5767 -641
rect 5770 -642 5799 -635
rect 5688 -643 5799 -642
rect 5688 -644 5805 -643
rect 5364 -652 5415 -644
rect 5462 -652 5496 -644
rect 5364 -664 5389 -652
rect 5396 -664 5415 -652
rect 5469 -654 5496 -652
rect 5505 -654 5726 -644
rect 5761 -647 5767 -644
rect 5469 -658 5726 -654
rect 5364 -672 5415 -664
rect 5462 -672 5726 -658
rect 5770 -652 5805 -644
rect 5316 -720 5335 -686
rect 5380 -680 5409 -672
rect 5380 -686 5397 -680
rect 5380 -688 5414 -686
rect 5462 -688 5478 -672
rect 5479 -682 5687 -672
rect 5688 -682 5704 -672
rect 5752 -676 5767 -661
rect 5770 -664 5771 -652
rect 5778 -664 5805 -652
rect 5770 -672 5805 -664
rect 5770 -673 5799 -672
rect 5490 -686 5704 -682
rect 5505 -688 5704 -686
rect 5739 -686 5752 -676
rect 5770 -686 5787 -673
rect 5739 -688 5787 -686
rect 5381 -692 5414 -688
rect 5377 -694 5414 -692
rect 5377 -695 5444 -694
rect 5377 -700 5408 -695
rect 5414 -700 5444 -695
rect 5377 -704 5444 -700
rect 5350 -707 5444 -704
rect 5350 -714 5399 -707
rect 5350 -720 5380 -714
rect 5399 -719 5404 -714
rect 5316 -736 5396 -720
rect 5408 -728 5444 -707
rect 5505 -712 5694 -688
rect 5739 -689 5786 -688
rect 5752 -694 5786 -689
rect 5520 -715 5694 -712
rect 5513 -718 5694 -715
rect 5722 -695 5786 -694
rect 5316 -738 5335 -736
rect 5350 -738 5384 -736
rect 5316 -754 5396 -738
rect 5316 -760 5335 -754
rect 5032 -786 5135 -776
rect 4986 -788 5135 -786
rect 5156 -788 5191 -776
rect 4825 -790 4987 -788
rect 4837 -808 4856 -790
rect 4871 -792 4901 -790
rect 4720 -818 4761 -810
rect 4844 -814 4856 -808
rect 4908 -808 4987 -790
rect 5019 -790 5191 -788
rect 5019 -806 5098 -790
rect 5105 -792 5135 -790
rect 4994 -808 5098 -806
rect 4683 -828 4712 -818
rect 4726 -828 4755 -818
rect 4770 -828 4800 -814
rect 4844 -828 4886 -814
rect 4908 -818 5098 -808
rect 5163 -810 5169 -790
rect 4893 -828 4923 -818
rect 4924 -828 5082 -818
rect 5086 -828 5116 -818
rect 5120 -828 5150 -814
rect 5178 -828 5191 -790
rect 5263 -776 5292 -760
rect 5306 -776 5335 -760
rect 5350 -770 5380 -754
rect 5408 -776 5414 -728
rect 5417 -734 5436 -728
rect 5451 -734 5481 -726
rect 5417 -742 5481 -734
rect 5417 -758 5497 -742
rect 5513 -749 5575 -718
rect 5591 -749 5653 -718
rect 5722 -720 5771 -695
rect 5786 -720 5816 -702
rect 5685 -734 5715 -726
rect 5722 -728 5832 -720
rect 5685 -742 5730 -734
rect 5417 -760 5436 -758
rect 5451 -760 5497 -758
rect 5417 -776 5497 -760
rect 5524 -762 5559 -749
rect 5600 -752 5637 -749
rect 5600 -754 5642 -752
rect 5529 -765 5559 -762
rect 5538 -769 5545 -765
rect 5545 -770 5546 -769
rect 5504 -776 5514 -770
rect 5263 -784 5298 -776
rect 5263 -810 5264 -784
rect 5271 -810 5298 -784
rect 5206 -828 5236 -814
rect 5263 -818 5298 -810
rect 5300 -784 5341 -776
rect 5300 -810 5315 -784
rect 5322 -810 5341 -784
rect 5405 -788 5436 -776
rect 5451 -788 5554 -776
rect 5566 -786 5592 -760
rect 5607 -765 5637 -754
rect 5669 -758 5731 -742
rect 5669 -760 5715 -758
rect 5669 -776 5731 -760
rect 5743 -776 5749 -728
rect 5752 -736 5832 -728
rect 5752 -738 5771 -736
rect 5786 -738 5820 -736
rect 5752 -753 5832 -738
rect 5752 -754 5838 -753
rect 5752 -776 5771 -754
rect 5786 -770 5816 -754
rect 5844 -760 5850 -686
rect 5853 -760 5872 -616
rect 5887 -760 5893 -616
rect 5902 -686 5915 -616
rect 5967 -620 5989 -616
rect 5960 -632 5977 -628
rect 5981 -630 5989 -628
rect 5979 -632 5989 -630
rect 5960 -642 5989 -632
rect 6042 -642 6058 -628
rect 6096 -632 6102 -630
rect 6109 -632 6217 -616
rect 6224 -632 6230 -630
rect 6238 -632 6253 -616
rect 6319 -622 6338 -619
rect 5960 -644 6058 -642
rect 6085 -644 6253 -632
rect 6268 -642 6284 -628
rect 6319 -641 6341 -622
rect 6351 -628 6367 -627
rect 6350 -630 6367 -628
rect 6351 -635 6367 -630
rect 6341 -642 6347 -641
rect 6350 -642 6379 -635
rect 6268 -643 6379 -642
rect 6268 -644 6385 -643
rect 5944 -652 5995 -644
rect 6042 -652 6076 -644
rect 5944 -664 5969 -652
rect 5976 -664 5995 -652
rect 6049 -654 6076 -652
rect 6085 -654 6306 -644
rect 6341 -647 6347 -644
rect 6049 -658 6306 -654
rect 5944 -672 5995 -664
rect 6042 -672 6306 -658
rect 6350 -652 6385 -644
rect 5896 -720 5915 -686
rect 5960 -680 5989 -672
rect 5960 -686 5977 -680
rect 5960 -688 5994 -686
rect 6042 -688 6058 -672
rect 6059 -682 6267 -672
rect 6268 -682 6284 -672
rect 6332 -676 6347 -661
rect 6350 -664 6351 -652
rect 6358 -664 6385 -652
rect 6350 -672 6385 -664
rect 6350 -673 6379 -672
rect 6070 -686 6284 -682
rect 6085 -688 6284 -686
rect 6319 -686 6332 -676
rect 6350 -686 6367 -673
rect 6319 -688 6367 -686
rect 5961 -692 5994 -688
rect 5957 -694 5994 -692
rect 5957 -695 6024 -694
rect 5957 -700 5988 -695
rect 5994 -700 6024 -695
rect 5957 -704 6024 -700
rect 5930 -707 6024 -704
rect 5930 -714 5979 -707
rect 5930 -720 5960 -714
rect 5979 -719 5984 -714
rect 5896 -736 5976 -720
rect 5988 -728 6024 -707
rect 6085 -712 6274 -688
rect 6319 -689 6366 -688
rect 6332 -694 6366 -689
rect 6100 -715 6274 -712
rect 6093 -718 6274 -715
rect 6302 -695 6366 -694
rect 5896 -738 5915 -736
rect 5930 -738 5964 -736
rect 5896 -754 5976 -738
rect 5896 -760 5915 -754
rect 5612 -786 5715 -776
rect 5566 -788 5715 -786
rect 5736 -788 5771 -776
rect 5405 -790 5567 -788
rect 5417 -808 5436 -790
rect 5451 -792 5481 -790
rect 5300 -818 5341 -810
rect 5424 -814 5436 -808
rect 5488 -808 5567 -790
rect 5599 -790 5771 -788
rect 5599 -806 5678 -790
rect 5685 -792 5715 -790
rect 5574 -808 5678 -806
rect 5263 -828 5292 -818
rect 5306 -828 5335 -818
rect 5350 -828 5380 -814
rect 5424 -828 5466 -814
rect 5488 -818 5678 -808
rect 5743 -810 5749 -790
rect 5473 -828 5503 -818
rect 5504 -828 5662 -818
rect 5666 -828 5696 -818
rect 5700 -828 5730 -814
rect 5758 -828 5771 -790
rect 5843 -776 5872 -760
rect 5886 -776 5915 -760
rect 5930 -770 5960 -754
rect 5988 -776 5994 -728
rect 5997 -734 6016 -728
rect 6031 -734 6061 -726
rect 5997 -742 6061 -734
rect 5997 -758 6077 -742
rect 6093 -749 6155 -718
rect 6171 -749 6233 -718
rect 6302 -720 6351 -695
rect 6366 -720 6396 -704
rect 6265 -734 6295 -726
rect 6302 -728 6412 -720
rect 6265 -742 6310 -734
rect 5997 -760 6016 -758
rect 6031 -760 6077 -758
rect 5997 -776 6077 -760
rect 6104 -762 6139 -749
rect 6180 -752 6217 -749
rect 6180 -754 6222 -752
rect 6109 -765 6139 -762
rect 6118 -769 6125 -765
rect 6125 -770 6126 -769
rect 6084 -776 6094 -770
rect 5843 -784 5878 -776
rect 5843 -810 5844 -784
rect 5851 -810 5878 -784
rect 5786 -828 5816 -814
rect 5843 -818 5878 -810
rect 5880 -784 5921 -776
rect 5880 -810 5895 -784
rect 5902 -810 5921 -784
rect 5985 -788 6016 -776
rect 6031 -788 6134 -776
rect 6146 -786 6172 -760
rect 6187 -765 6217 -754
rect 6249 -758 6311 -742
rect 6249 -760 6295 -758
rect 6249 -776 6311 -760
rect 6323 -776 6329 -728
rect 6332 -736 6412 -728
rect 6332 -738 6351 -736
rect 6366 -738 6400 -736
rect 6332 -754 6412 -738
rect 6332 -776 6351 -754
rect 6366 -770 6396 -754
rect 6424 -760 6430 -686
rect 6439 -760 6452 -616
rect 6192 -786 6295 -776
rect 6146 -788 6295 -786
rect 6316 -788 6351 -776
rect 5985 -790 6147 -788
rect 5997 -808 6016 -790
rect 6031 -792 6061 -790
rect 5880 -818 5921 -810
rect 6004 -814 6016 -808
rect 6068 -808 6147 -790
rect 6179 -790 6351 -788
rect 6179 -806 6258 -790
rect 6265 -792 6295 -790
rect 6154 -808 6258 -806
rect 5843 -828 5872 -818
rect 5886 -828 5915 -818
rect 5930 -828 5960 -814
rect 6004 -828 6046 -814
rect 6068 -818 6258 -808
rect 6323 -810 6329 -790
rect 6053 -828 6083 -818
rect 6084 -828 6242 -818
rect 6246 -828 6276 -818
rect 6280 -828 6310 -814
rect 6338 -828 6351 -790
rect 6423 -776 6452 -760
rect 6423 -784 6458 -776
rect 6423 -810 6424 -784
rect 6431 -810 6458 -784
rect 6366 -828 6396 -814
rect 6423 -818 6458 -810
rect 6423 -828 6452 -818
rect -541 -842 6452 -828
rect -478 -872 -465 -842
rect -450 -856 -420 -842
rect -376 -856 -334 -842
rect -327 -856 -107 -842
rect -100 -856 -70 -842
rect -410 -870 -395 -858
rect -376 -870 -363 -856
rect -295 -860 -142 -856
rect -413 -872 -391 -870
rect -313 -872 -121 -860
rect -42 -872 -29 -842
rect -14 -856 16 -842
rect 53 -872 72 -842
rect 87 -872 93 -842
rect 102 -872 115 -842
rect 130 -856 160 -842
rect 204 -856 246 -842
rect 253 -856 473 -842
rect 480 -856 510 -842
rect 170 -870 185 -858
rect 204 -870 217 -856
rect 285 -860 438 -856
rect 167 -872 189 -870
rect 267 -872 459 -860
rect 538 -872 551 -842
rect 566 -856 596 -842
rect 633 -872 652 -842
rect 667 -872 673 -842
rect 682 -872 695 -842
rect 710 -856 740 -842
rect 784 -856 826 -842
rect 833 -856 1053 -842
rect 1060 -856 1090 -842
rect 750 -870 765 -858
rect 784 -870 797 -856
rect 865 -860 1018 -856
rect 747 -872 769 -870
rect 847 -872 1039 -860
rect 1118 -872 1131 -842
rect 1146 -856 1176 -842
rect 1213 -872 1232 -842
rect 1247 -872 1253 -842
rect 1262 -872 1275 -842
rect 1290 -856 1320 -842
rect 1364 -856 1406 -842
rect 1413 -856 1633 -842
rect 1640 -856 1670 -842
rect 1330 -870 1345 -858
rect 1364 -870 1377 -856
rect 1445 -860 1598 -856
rect 1327 -872 1349 -870
rect 1427 -872 1619 -860
rect 1698 -872 1711 -842
rect 1726 -856 1756 -842
rect 1793 -872 1812 -842
rect 1827 -872 1833 -842
rect 1842 -872 1855 -842
rect 1870 -856 1900 -842
rect 1944 -856 1986 -842
rect 1993 -856 2213 -842
rect 2220 -856 2250 -842
rect 1910 -870 1925 -858
rect 1944 -870 1957 -856
rect 2025 -860 2178 -856
rect 1907 -872 1929 -870
rect 2007 -872 2199 -860
rect 2278 -872 2291 -842
rect 2306 -856 2336 -842
rect 2373 -872 2392 -842
rect 2407 -872 2413 -842
rect 2422 -872 2435 -842
rect 2450 -856 2480 -842
rect 2524 -856 2566 -842
rect 2573 -856 2793 -842
rect 2800 -856 2830 -842
rect 2490 -870 2505 -858
rect 2524 -870 2537 -856
rect 2605 -860 2758 -856
rect 2487 -872 2509 -870
rect 2587 -872 2779 -860
rect 2858 -872 2871 -842
rect 2886 -856 2916 -842
rect 2953 -872 2972 -842
rect 2987 -872 2993 -842
rect 3002 -872 3015 -842
rect 3030 -856 3060 -842
rect 3104 -856 3146 -842
rect 3153 -856 3373 -842
rect 3380 -856 3410 -842
rect 3070 -870 3085 -858
rect 3104 -870 3117 -856
rect 3185 -860 3338 -856
rect 3067 -872 3089 -870
rect 3167 -872 3359 -860
rect 3438 -872 3451 -842
rect 3466 -856 3496 -842
rect 3533 -872 3552 -842
rect 3567 -872 3573 -842
rect 3582 -872 3595 -842
rect 3610 -856 3640 -842
rect 3684 -856 3726 -842
rect 3733 -856 3953 -842
rect 3960 -856 3990 -842
rect 3650 -870 3665 -858
rect 3684 -870 3697 -856
rect 3765 -860 3918 -856
rect 3647 -872 3669 -870
rect 3747 -872 3939 -860
rect 4018 -872 4031 -842
rect 4046 -856 4076 -842
rect 4113 -872 4132 -842
rect 4147 -872 4153 -842
rect 4162 -872 4175 -842
rect 4190 -856 4220 -842
rect 4264 -856 4306 -842
rect 4313 -856 4533 -842
rect 4540 -856 4570 -842
rect 4230 -870 4245 -858
rect 4264 -870 4277 -856
rect 4345 -860 4498 -856
rect 4227 -872 4249 -870
rect 4327 -872 4519 -860
rect 4598 -872 4611 -842
rect 4626 -856 4656 -842
rect 4693 -872 4712 -842
rect 4727 -872 4733 -842
rect 4742 -872 4755 -842
rect 4770 -856 4800 -842
rect 4844 -856 4886 -842
rect 4893 -856 5113 -842
rect 5120 -856 5150 -842
rect 4810 -870 4825 -858
rect 4844 -870 4857 -856
rect 4925 -860 5078 -856
rect 4807 -872 4829 -870
rect 4907 -872 5099 -860
rect 5178 -872 5191 -842
rect 5206 -856 5236 -842
rect 5273 -872 5292 -842
rect 5307 -872 5313 -842
rect 5322 -872 5335 -842
rect 5350 -856 5380 -842
rect 5424 -856 5466 -842
rect 5473 -856 5693 -842
rect 5700 -856 5730 -842
rect 5390 -870 5405 -858
rect 5424 -870 5437 -856
rect 5505 -860 5658 -856
rect 5387 -872 5409 -870
rect 5487 -872 5679 -860
rect 5758 -872 5771 -842
rect 5786 -856 5816 -842
rect 5853 -872 5872 -842
rect 5887 -872 5893 -842
rect 5902 -872 5915 -842
rect 5930 -856 5960 -842
rect 6004 -856 6046 -842
rect 6053 -856 6273 -842
rect 6280 -856 6310 -842
rect 5970 -870 5985 -858
rect 6004 -870 6017 -856
rect 6085 -860 6238 -856
rect 5967 -872 5989 -870
rect 6067 -872 6259 -860
rect 6338 -872 6351 -842
rect 6366 -856 6396 -842
rect 6439 -872 6452 -842
rect -541 -886 6452 -872
rect -478 -956 -465 -886
rect -413 -890 -391 -886
rect -420 -902 -403 -898
rect -399 -900 -391 -898
rect -401 -902 -391 -900
rect -420 -912 -391 -902
rect -338 -912 -322 -898
rect -284 -902 -278 -900
rect -271 -902 -163 -886
rect -156 -902 -150 -900
rect -142 -902 -127 -886
rect -61 -892 -42 -889
rect -420 -914 -322 -912
rect -295 -914 -127 -902
rect -112 -912 -96 -898
rect -61 -911 -39 -892
rect -29 -898 -13 -897
rect -30 -900 -13 -898
rect -29 -905 -13 -900
rect -39 -912 -33 -911
rect -30 -912 -1 -905
rect -112 -913 -1 -912
rect -112 -914 5 -913
rect -436 -922 -385 -914
rect -338 -922 -304 -914
rect -436 -934 -411 -922
rect -404 -934 -385 -922
rect -331 -924 -304 -922
rect -295 -924 -74 -914
rect -39 -917 -33 -914
rect -331 -928 -74 -924
rect -436 -942 -385 -934
rect -338 -942 -74 -928
rect -30 -922 5 -914
rect -484 -990 -465 -956
rect -420 -950 -391 -942
rect -420 -956 -403 -950
rect -420 -958 -386 -956
rect -338 -958 -322 -942
rect -321 -952 -113 -942
rect -112 -952 -96 -942
rect -48 -946 -33 -931
rect -30 -934 -29 -922
rect -22 -934 5 -922
rect -30 -942 5 -934
rect -30 -943 -1 -942
rect -310 -956 -96 -952
rect -295 -958 -96 -956
rect -61 -956 -48 -946
rect -30 -956 -13 -943
rect -61 -958 -13 -956
rect -419 -962 -386 -958
rect -423 -964 -386 -962
rect -423 -965 -356 -964
rect -423 -970 -392 -965
rect -386 -970 -356 -965
rect -423 -974 -356 -970
rect -450 -977 -356 -974
rect -450 -984 -401 -977
rect -450 -990 -420 -984
rect -401 -989 -396 -984
rect -484 -1006 -404 -990
rect -392 -998 -356 -977
rect -295 -982 -106 -958
rect -61 -959 -14 -958
rect -48 -964 -14 -959
rect -280 -985 -106 -982
rect -287 -988 -106 -985
rect -78 -965 -14 -964
rect -484 -1008 -465 -1006
rect -450 -1008 -416 -1006
rect -484 -1024 -404 -1008
rect -484 -1030 -465 -1024
rect -494 -1046 -465 -1030
rect -450 -1040 -420 -1024
rect -392 -1046 -386 -998
rect -383 -1004 -364 -998
rect -349 -1004 -319 -996
rect -383 -1012 -319 -1004
rect -383 -1028 -303 -1012
rect -287 -1019 -225 -988
rect -209 -1019 -147 -988
rect -78 -990 -29 -965
rect -14 -990 16 -972
rect -115 -1004 -85 -996
rect -78 -998 32 -990
rect -115 -1012 -70 -1004
rect -383 -1030 -364 -1028
rect -349 -1030 -303 -1028
rect -383 -1046 -303 -1030
rect -276 -1032 -241 -1019
rect -200 -1022 -163 -1019
rect -200 -1024 -158 -1022
rect -271 -1035 -241 -1032
rect -262 -1039 -255 -1035
rect -255 -1040 -254 -1039
rect -296 -1046 -286 -1040
rect -500 -1054 -459 -1046
rect -500 -1080 -485 -1054
rect -478 -1080 -459 -1054
rect -395 -1058 -364 -1046
rect -349 -1058 -246 -1046
rect -234 -1056 -208 -1030
rect -193 -1035 -163 -1024
rect -131 -1028 -69 -1012
rect -131 -1030 -85 -1028
rect -131 -1046 -69 -1030
rect -57 -1046 -51 -998
rect -48 -1006 32 -998
rect -48 -1008 -29 -1006
rect -14 -1008 20 -1006
rect -48 -1023 32 -1008
rect -48 -1024 38 -1023
rect -48 -1046 -29 -1024
rect -14 -1040 16 -1024
rect 44 -1030 50 -956
rect 53 -1030 72 -886
rect 87 -1030 93 -886
rect 102 -956 115 -886
rect 167 -890 189 -886
rect 160 -902 177 -898
rect 181 -900 189 -898
rect 179 -902 189 -900
rect 160 -912 189 -902
rect 242 -912 258 -898
rect 296 -902 302 -900
rect 309 -902 417 -886
rect 424 -902 430 -900
rect 438 -902 453 -886
rect 519 -892 538 -889
rect 160 -914 258 -912
rect 285 -914 453 -902
rect 468 -912 484 -898
rect 519 -911 541 -892
rect 551 -898 567 -897
rect 550 -900 567 -898
rect 551 -905 567 -900
rect 541 -912 547 -911
rect 550 -912 579 -905
rect 468 -913 579 -912
rect 468 -914 585 -913
rect 144 -922 195 -914
rect 242 -922 276 -914
rect 144 -934 169 -922
rect 176 -934 195 -922
rect 249 -924 276 -922
rect 285 -924 506 -914
rect 541 -917 547 -914
rect 249 -928 506 -924
rect 144 -942 195 -934
rect 242 -942 506 -928
rect 550 -922 585 -914
rect 96 -990 115 -956
rect 160 -950 189 -942
rect 160 -956 177 -950
rect 160 -958 194 -956
rect 242 -958 258 -942
rect 259 -952 467 -942
rect 468 -952 484 -942
rect 532 -946 547 -931
rect 550 -934 551 -922
rect 558 -934 585 -922
rect 550 -942 585 -934
rect 550 -943 579 -942
rect 270 -956 484 -952
rect 285 -958 484 -956
rect 519 -956 532 -946
rect 550 -956 567 -943
rect 519 -958 567 -956
rect 161 -962 194 -958
rect 157 -964 194 -962
rect 157 -965 224 -964
rect 157 -970 188 -965
rect 194 -970 224 -965
rect 157 -974 224 -970
rect 130 -977 224 -974
rect 130 -984 179 -977
rect 130 -990 160 -984
rect 179 -989 184 -984
rect 96 -1006 176 -990
rect 188 -998 224 -977
rect 285 -982 474 -958
rect 519 -959 566 -958
rect 532 -964 566 -959
rect 606 -964 622 -962
rect 300 -985 474 -982
rect 293 -988 474 -985
rect 502 -965 566 -964
rect 96 -1008 115 -1006
rect 130 -1008 164 -1006
rect 96 -1024 176 -1008
rect 96 -1030 115 -1024
rect -188 -1056 -85 -1046
rect -234 -1058 -85 -1056
rect -64 -1058 -29 -1046
rect -395 -1060 -233 -1058
rect -383 -1080 -364 -1060
rect -349 -1062 -319 -1060
rect -500 -1088 -459 -1080
rect -377 -1084 -364 -1080
rect -312 -1076 -233 -1060
rect -201 -1060 -29 -1058
rect -201 -1076 -122 -1060
rect -115 -1062 -85 -1060
rect -494 -1098 -465 -1088
rect -450 -1098 -420 -1084
rect -377 -1098 -334 -1084
rect -312 -1088 -122 -1076
rect -57 -1080 -51 -1060
rect -327 -1098 -297 -1088
rect -296 -1098 -138 -1088
rect -134 -1098 -104 -1088
rect -100 -1098 -70 -1084
rect -42 -1098 -29 -1060
rect 43 -1046 72 -1030
rect 86 -1046 115 -1030
rect 130 -1040 160 -1024
rect 188 -1046 194 -998
rect 197 -1004 216 -998
rect 231 -1004 261 -996
rect 197 -1012 261 -1004
rect 197 -1028 277 -1012
rect 293 -1019 355 -988
rect 371 -1019 433 -988
rect 502 -990 551 -965
rect 596 -974 622 -964
rect 566 -990 622 -974
rect 465 -1004 495 -996
rect 502 -998 612 -990
rect 465 -1012 510 -1004
rect 197 -1030 216 -1028
rect 231 -1030 277 -1028
rect 197 -1046 277 -1030
rect 304 -1032 339 -1019
rect 380 -1022 417 -1019
rect 380 -1024 422 -1022
rect 309 -1035 339 -1032
rect 318 -1039 325 -1035
rect 325 -1040 326 -1039
rect 284 -1046 294 -1040
rect 43 -1054 78 -1046
rect 43 -1080 44 -1054
rect 51 -1080 78 -1054
rect -14 -1098 16 -1084
rect 43 -1088 78 -1080
rect 80 -1054 121 -1046
rect 80 -1080 95 -1054
rect 102 -1080 121 -1054
rect 185 -1058 216 -1046
rect 231 -1058 334 -1046
rect 346 -1056 372 -1030
rect 387 -1035 417 -1024
rect 449 -1028 511 -1012
rect 449 -1030 495 -1028
rect 449 -1046 511 -1030
rect 523 -1046 529 -998
rect 532 -1006 612 -998
rect 532 -1008 551 -1006
rect 566 -1008 600 -1006
rect 532 -1024 612 -1008
rect 532 -1046 551 -1024
rect 566 -1040 596 -1024
rect 624 -1030 630 -956
rect 633 -1030 652 -886
rect 667 -1030 673 -886
rect 682 -956 695 -886
rect 747 -890 769 -886
rect 740 -902 757 -898
rect 761 -900 769 -898
rect 759 -902 769 -900
rect 740 -912 769 -902
rect 822 -912 838 -898
rect 876 -902 882 -900
rect 889 -902 997 -886
rect 1004 -902 1010 -900
rect 1018 -902 1033 -886
rect 1099 -892 1118 -889
rect 740 -914 838 -912
rect 865 -914 1033 -902
rect 1048 -912 1064 -898
rect 1099 -911 1121 -892
rect 1131 -898 1147 -897
rect 1130 -900 1147 -898
rect 1131 -905 1147 -900
rect 1121 -912 1127 -911
rect 1130 -912 1159 -905
rect 1048 -913 1159 -912
rect 1048 -914 1165 -913
rect 724 -922 775 -914
rect 822 -922 856 -914
rect 724 -934 749 -922
rect 756 -934 775 -922
rect 829 -924 856 -922
rect 865 -924 1086 -914
rect 1121 -917 1127 -914
rect 829 -928 1086 -924
rect 724 -942 775 -934
rect 822 -942 1086 -928
rect 1130 -922 1165 -914
rect 676 -990 695 -956
rect 740 -950 769 -942
rect 740 -956 757 -950
rect 740 -958 774 -956
rect 822 -958 838 -942
rect 839 -952 1047 -942
rect 1048 -952 1064 -942
rect 1112 -946 1127 -931
rect 1130 -934 1131 -922
rect 1138 -934 1165 -922
rect 1130 -942 1165 -934
rect 1130 -943 1159 -942
rect 850 -956 1064 -952
rect 865 -958 1064 -956
rect 1099 -956 1112 -946
rect 1130 -956 1147 -943
rect 1099 -958 1147 -956
rect 741 -962 774 -958
rect 737 -964 774 -962
rect 737 -965 804 -964
rect 737 -970 768 -965
rect 774 -970 804 -965
rect 737 -974 804 -970
rect 710 -977 804 -974
rect 710 -984 759 -977
rect 710 -990 740 -984
rect 759 -989 764 -984
rect 676 -1006 756 -990
rect 768 -998 804 -977
rect 865 -982 1054 -958
rect 1099 -959 1146 -958
rect 1112 -964 1146 -959
rect 880 -985 1054 -982
rect 873 -988 1054 -985
rect 1082 -965 1146 -964
rect 676 -1008 695 -1006
rect 710 -1008 744 -1006
rect 676 -1024 756 -1008
rect 676 -1030 695 -1024
rect 392 -1056 495 -1046
rect 346 -1058 495 -1056
rect 516 -1058 551 -1046
rect 185 -1060 347 -1058
rect 197 -1080 216 -1060
rect 231 -1062 261 -1060
rect 80 -1088 121 -1080
rect 203 -1084 216 -1080
rect 268 -1076 347 -1060
rect 379 -1060 551 -1058
rect 379 -1076 458 -1060
rect 465 -1062 495 -1060
rect 43 -1098 72 -1088
rect 86 -1098 115 -1088
rect 130 -1098 160 -1084
rect 203 -1098 246 -1084
rect 268 -1088 458 -1076
rect 523 -1080 529 -1060
rect 253 -1098 283 -1088
rect 284 -1098 442 -1088
rect 446 -1098 476 -1088
rect 480 -1098 510 -1084
rect 538 -1098 551 -1060
rect 623 -1046 652 -1030
rect 666 -1046 695 -1030
rect 710 -1040 740 -1024
rect 768 -1046 774 -998
rect 777 -1004 796 -998
rect 811 -1004 841 -996
rect 777 -1012 841 -1004
rect 777 -1028 857 -1012
rect 873 -1019 935 -988
rect 951 -1019 1013 -988
rect 1082 -990 1131 -965
rect 1146 -990 1176 -972
rect 1045 -1004 1075 -996
rect 1082 -998 1192 -990
rect 1045 -1012 1090 -1004
rect 777 -1030 796 -1028
rect 811 -1030 857 -1028
rect 777 -1046 857 -1030
rect 884 -1032 919 -1019
rect 960 -1022 997 -1019
rect 960 -1024 1002 -1022
rect 889 -1035 919 -1032
rect 898 -1039 905 -1035
rect 905 -1040 906 -1039
rect 864 -1046 874 -1040
rect 623 -1054 658 -1046
rect 623 -1080 624 -1054
rect 631 -1080 658 -1054
rect 566 -1098 596 -1084
rect 623 -1088 658 -1080
rect 660 -1054 701 -1046
rect 660 -1080 675 -1054
rect 682 -1080 701 -1054
rect 765 -1058 796 -1046
rect 811 -1058 914 -1046
rect 926 -1056 952 -1030
rect 967 -1035 997 -1024
rect 1029 -1028 1091 -1012
rect 1029 -1030 1075 -1028
rect 1029 -1046 1091 -1030
rect 1103 -1046 1109 -998
rect 1112 -1006 1192 -998
rect 1112 -1008 1131 -1006
rect 1146 -1008 1180 -1006
rect 1112 -1023 1192 -1008
rect 1112 -1024 1198 -1023
rect 1112 -1046 1131 -1024
rect 1146 -1040 1176 -1024
rect 1204 -1030 1210 -956
rect 1213 -1030 1232 -886
rect 1247 -1030 1253 -886
rect 1262 -956 1275 -886
rect 1327 -890 1349 -886
rect 1320 -902 1337 -898
rect 1341 -900 1349 -898
rect 1339 -902 1349 -900
rect 1320 -912 1349 -902
rect 1402 -912 1418 -898
rect 1456 -902 1462 -900
rect 1469 -902 1577 -886
rect 1584 -902 1590 -900
rect 1598 -902 1613 -886
rect 1679 -892 1698 -889
rect 1320 -914 1418 -912
rect 1445 -914 1613 -902
rect 1628 -912 1644 -898
rect 1679 -911 1701 -892
rect 1711 -898 1727 -897
rect 1710 -900 1727 -898
rect 1711 -905 1727 -900
rect 1701 -912 1707 -911
rect 1710 -912 1739 -905
rect 1628 -913 1739 -912
rect 1628 -914 1745 -913
rect 1304 -922 1355 -914
rect 1402 -922 1436 -914
rect 1304 -934 1329 -922
rect 1336 -934 1355 -922
rect 1409 -924 1436 -922
rect 1445 -924 1666 -914
rect 1701 -917 1707 -914
rect 1409 -928 1666 -924
rect 1304 -942 1355 -934
rect 1402 -942 1666 -928
rect 1710 -922 1745 -914
rect 1256 -990 1275 -956
rect 1320 -950 1349 -942
rect 1320 -956 1337 -950
rect 1320 -958 1354 -956
rect 1402 -958 1418 -942
rect 1419 -952 1627 -942
rect 1628 -952 1644 -942
rect 1692 -946 1707 -931
rect 1710 -934 1711 -922
rect 1718 -934 1745 -922
rect 1710 -942 1745 -934
rect 1710 -943 1739 -942
rect 1430 -956 1644 -952
rect 1445 -958 1644 -956
rect 1679 -956 1692 -946
rect 1710 -956 1727 -943
rect 1679 -958 1727 -956
rect 1321 -962 1354 -958
rect 1317 -964 1354 -962
rect 1317 -965 1384 -964
rect 1317 -970 1348 -965
rect 1354 -970 1384 -965
rect 1317 -974 1384 -970
rect 1290 -977 1384 -974
rect 1290 -984 1339 -977
rect 1290 -990 1320 -984
rect 1339 -989 1344 -984
rect 1256 -1006 1336 -990
rect 1348 -998 1384 -977
rect 1445 -982 1634 -958
rect 1679 -959 1726 -958
rect 1692 -964 1726 -959
rect 1766 -964 1782 -962
rect 1460 -985 1634 -982
rect 1453 -988 1634 -985
rect 1662 -965 1726 -964
rect 1256 -1008 1275 -1006
rect 1290 -1008 1324 -1006
rect 1256 -1024 1336 -1008
rect 1256 -1030 1275 -1024
rect 972 -1056 1075 -1046
rect 926 -1058 1075 -1056
rect 1096 -1058 1131 -1046
rect 765 -1060 927 -1058
rect 777 -1080 796 -1060
rect 811 -1062 841 -1060
rect 660 -1088 701 -1080
rect 783 -1084 796 -1080
rect 848 -1076 927 -1060
rect 959 -1060 1131 -1058
rect 959 -1076 1038 -1060
rect 1045 -1062 1075 -1060
rect 623 -1098 652 -1088
rect 666 -1098 695 -1088
rect 710 -1098 740 -1084
rect 783 -1098 826 -1084
rect 848 -1088 1038 -1076
rect 1103 -1080 1109 -1060
rect 833 -1098 863 -1088
rect 864 -1098 1022 -1088
rect 1026 -1098 1056 -1088
rect 1060 -1098 1090 -1084
rect 1118 -1098 1131 -1060
rect 1203 -1046 1232 -1030
rect 1246 -1046 1275 -1030
rect 1290 -1040 1320 -1024
rect 1348 -1046 1354 -998
rect 1357 -1004 1376 -998
rect 1391 -1004 1421 -996
rect 1357 -1012 1421 -1004
rect 1357 -1028 1437 -1012
rect 1453 -1019 1515 -988
rect 1531 -1019 1593 -988
rect 1662 -990 1711 -965
rect 1756 -974 1782 -964
rect 1726 -990 1782 -974
rect 1625 -1004 1655 -996
rect 1662 -998 1772 -990
rect 1625 -1012 1670 -1004
rect 1357 -1030 1376 -1028
rect 1391 -1030 1437 -1028
rect 1357 -1046 1437 -1030
rect 1464 -1032 1499 -1019
rect 1540 -1022 1577 -1019
rect 1540 -1024 1582 -1022
rect 1469 -1035 1499 -1032
rect 1478 -1039 1485 -1035
rect 1485 -1040 1486 -1039
rect 1444 -1046 1454 -1040
rect 1203 -1054 1238 -1046
rect 1203 -1080 1204 -1054
rect 1211 -1080 1238 -1054
rect 1146 -1098 1176 -1084
rect 1203 -1088 1238 -1080
rect 1240 -1054 1281 -1046
rect 1240 -1080 1255 -1054
rect 1262 -1080 1281 -1054
rect 1345 -1058 1376 -1046
rect 1391 -1058 1494 -1046
rect 1506 -1056 1532 -1030
rect 1547 -1035 1577 -1024
rect 1609 -1028 1671 -1012
rect 1609 -1030 1655 -1028
rect 1609 -1046 1671 -1030
rect 1683 -1046 1689 -998
rect 1692 -1006 1772 -998
rect 1692 -1008 1711 -1006
rect 1726 -1008 1760 -1006
rect 1692 -1024 1772 -1008
rect 1692 -1046 1711 -1024
rect 1726 -1040 1756 -1024
rect 1784 -1030 1790 -956
rect 1793 -1030 1812 -886
rect 1827 -1030 1833 -886
rect 1842 -956 1855 -886
rect 1907 -890 1929 -886
rect 1900 -902 1917 -898
rect 1921 -900 1929 -898
rect 1919 -902 1929 -900
rect 1900 -912 1929 -902
rect 1982 -912 1998 -898
rect 2036 -902 2042 -900
rect 2049 -902 2157 -886
rect 2164 -902 2170 -900
rect 2178 -902 2193 -886
rect 2259 -892 2278 -889
rect 1900 -914 1998 -912
rect 2025 -914 2193 -902
rect 2208 -912 2224 -898
rect 2259 -911 2281 -892
rect 2291 -898 2307 -897
rect 2290 -900 2307 -898
rect 2291 -905 2307 -900
rect 2281 -912 2287 -911
rect 2290 -912 2319 -905
rect 2208 -913 2319 -912
rect 2208 -914 2325 -913
rect 1884 -922 1935 -914
rect 1982 -922 2016 -914
rect 1884 -934 1909 -922
rect 1916 -934 1935 -922
rect 1989 -924 2016 -922
rect 2025 -924 2246 -914
rect 2281 -917 2287 -914
rect 1989 -928 2246 -924
rect 1884 -942 1935 -934
rect 1982 -942 2246 -928
rect 2290 -922 2325 -914
rect 1836 -990 1855 -956
rect 1900 -950 1929 -942
rect 1900 -956 1917 -950
rect 1900 -958 1934 -956
rect 1982 -958 1998 -942
rect 1999 -952 2207 -942
rect 2208 -952 2224 -942
rect 2272 -946 2287 -931
rect 2290 -934 2291 -922
rect 2298 -934 2325 -922
rect 2290 -942 2325 -934
rect 2290 -943 2319 -942
rect 2010 -956 2224 -952
rect 2025 -958 2224 -956
rect 2259 -956 2272 -946
rect 2290 -956 2307 -943
rect 2259 -958 2307 -956
rect 1901 -962 1934 -958
rect 1897 -964 1934 -962
rect 1897 -965 1964 -964
rect 1897 -970 1928 -965
rect 1934 -970 1964 -965
rect 1897 -974 1964 -970
rect 1870 -977 1964 -974
rect 1870 -984 1919 -977
rect 1870 -990 1900 -984
rect 1919 -989 1924 -984
rect 1836 -1006 1916 -990
rect 1928 -998 1964 -977
rect 2025 -982 2214 -958
rect 2259 -959 2306 -958
rect 2272 -964 2306 -959
rect 2040 -985 2214 -982
rect 2033 -988 2214 -985
rect 2242 -965 2306 -964
rect 1836 -1008 1855 -1006
rect 1870 -1008 1904 -1006
rect 1836 -1024 1916 -1008
rect 1836 -1030 1855 -1024
rect 1552 -1056 1655 -1046
rect 1506 -1058 1655 -1056
rect 1676 -1058 1711 -1046
rect 1345 -1060 1507 -1058
rect 1357 -1080 1376 -1060
rect 1391 -1062 1421 -1060
rect 1240 -1088 1281 -1080
rect 1363 -1084 1376 -1080
rect 1428 -1076 1507 -1060
rect 1539 -1060 1711 -1058
rect 1539 -1076 1618 -1060
rect 1625 -1062 1655 -1060
rect 1203 -1098 1232 -1088
rect 1246 -1098 1275 -1088
rect 1290 -1098 1320 -1084
rect 1363 -1098 1406 -1084
rect 1428 -1088 1618 -1076
rect 1683 -1080 1689 -1060
rect 1413 -1098 1443 -1088
rect 1444 -1098 1602 -1088
rect 1606 -1098 1636 -1088
rect 1640 -1098 1670 -1084
rect 1698 -1098 1711 -1060
rect 1783 -1046 1812 -1030
rect 1826 -1046 1855 -1030
rect 1870 -1040 1900 -1024
rect 1928 -1046 1934 -998
rect 1937 -1004 1956 -998
rect 1971 -1004 2001 -996
rect 1937 -1012 2001 -1004
rect 1937 -1028 2017 -1012
rect 2033 -1019 2095 -988
rect 2111 -1019 2173 -988
rect 2242 -990 2291 -965
rect 2306 -990 2336 -972
rect 2205 -1004 2235 -996
rect 2242 -998 2352 -990
rect 2205 -1012 2250 -1004
rect 1937 -1030 1956 -1028
rect 1971 -1030 2017 -1028
rect 1937 -1046 2017 -1030
rect 2044 -1032 2079 -1019
rect 2120 -1022 2157 -1019
rect 2120 -1024 2162 -1022
rect 2049 -1035 2079 -1032
rect 2058 -1039 2065 -1035
rect 2065 -1040 2066 -1039
rect 2024 -1046 2034 -1040
rect 1783 -1054 1818 -1046
rect 1783 -1080 1784 -1054
rect 1791 -1080 1818 -1054
rect 1726 -1098 1756 -1084
rect 1783 -1088 1818 -1080
rect 1820 -1054 1861 -1046
rect 1820 -1080 1835 -1054
rect 1842 -1080 1861 -1054
rect 1925 -1058 1956 -1046
rect 1971 -1058 2074 -1046
rect 2086 -1056 2112 -1030
rect 2127 -1035 2157 -1024
rect 2189 -1028 2251 -1012
rect 2189 -1030 2235 -1028
rect 2189 -1046 2251 -1030
rect 2263 -1046 2269 -998
rect 2272 -1006 2352 -998
rect 2272 -1008 2291 -1006
rect 2306 -1008 2340 -1006
rect 2272 -1023 2352 -1008
rect 2272 -1024 2358 -1023
rect 2272 -1046 2291 -1024
rect 2306 -1040 2336 -1024
rect 2364 -1030 2370 -956
rect 2373 -1030 2392 -886
rect 2407 -1030 2413 -886
rect 2422 -956 2435 -886
rect 2487 -890 2509 -886
rect 2480 -902 2497 -898
rect 2501 -900 2509 -898
rect 2499 -902 2509 -900
rect 2480 -912 2509 -902
rect 2562 -912 2578 -898
rect 2616 -902 2622 -900
rect 2629 -902 2737 -886
rect 2744 -902 2750 -900
rect 2758 -902 2773 -886
rect 2839 -892 2858 -889
rect 2480 -914 2578 -912
rect 2605 -914 2773 -902
rect 2788 -912 2804 -898
rect 2839 -911 2861 -892
rect 2871 -898 2887 -897
rect 2870 -900 2887 -898
rect 2871 -905 2887 -900
rect 2861 -912 2867 -911
rect 2870 -912 2899 -905
rect 2788 -913 2899 -912
rect 2788 -914 2905 -913
rect 2464 -922 2515 -914
rect 2562 -922 2596 -914
rect 2464 -934 2489 -922
rect 2496 -934 2515 -922
rect 2569 -924 2596 -922
rect 2605 -924 2826 -914
rect 2861 -917 2867 -914
rect 2569 -928 2826 -924
rect 2464 -942 2515 -934
rect 2562 -942 2826 -928
rect 2870 -922 2905 -914
rect 2416 -990 2435 -956
rect 2480 -950 2509 -942
rect 2480 -956 2497 -950
rect 2480 -958 2514 -956
rect 2562 -958 2578 -942
rect 2579 -952 2787 -942
rect 2788 -952 2804 -942
rect 2852 -946 2867 -931
rect 2870 -934 2871 -922
rect 2878 -934 2905 -922
rect 2870 -942 2905 -934
rect 2870 -943 2899 -942
rect 2590 -956 2804 -952
rect 2605 -958 2804 -956
rect 2839 -956 2852 -946
rect 2870 -956 2887 -943
rect 2839 -958 2887 -956
rect 2481 -962 2514 -958
rect 2477 -964 2514 -962
rect 2477 -965 2544 -964
rect 2477 -970 2508 -965
rect 2514 -970 2544 -965
rect 2477 -974 2544 -970
rect 2450 -977 2544 -974
rect 2450 -984 2499 -977
rect 2450 -990 2480 -984
rect 2499 -989 2504 -984
rect 2416 -1006 2496 -990
rect 2508 -998 2544 -977
rect 2605 -982 2794 -958
rect 2839 -959 2886 -958
rect 2852 -964 2886 -959
rect 2926 -964 2942 -962
rect 2620 -985 2794 -982
rect 2613 -988 2794 -985
rect 2822 -965 2886 -964
rect 2416 -1008 2435 -1006
rect 2450 -1008 2484 -1006
rect 2416 -1024 2496 -1008
rect 2416 -1030 2435 -1024
rect 2132 -1056 2235 -1046
rect 2086 -1058 2235 -1056
rect 2256 -1058 2291 -1046
rect 1925 -1060 2087 -1058
rect 1937 -1080 1956 -1060
rect 1971 -1062 2001 -1060
rect 1820 -1088 1861 -1080
rect 1943 -1084 1956 -1080
rect 2008 -1076 2087 -1060
rect 2119 -1060 2291 -1058
rect 2119 -1076 2198 -1060
rect 2205 -1062 2235 -1060
rect 1783 -1098 1812 -1088
rect 1826 -1098 1855 -1088
rect 1870 -1098 1900 -1084
rect 1943 -1098 1986 -1084
rect 2008 -1088 2198 -1076
rect 2263 -1080 2269 -1060
rect 1993 -1098 2023 -1088
rect 2024 -1098 2182 -1088
rect 2186 -1098 2216 -1088
rect 2220 -1098 2250 -1084
rect 2278 -1098 2291 -1060
rect 2363 -1046 2392 -1030
rect 2406 -1046 2435 -1030
rect 2450 -1040 2480 -1024
rect 2508 -1046 2514 -998
rect 2517 -1004 2536 -998
rect 2551 -1004 2581 -996
rect 2517 -1012 2581 -1004
rect 2517 -1028 2597 -1012
rect 2613 -1019 2675 -988
rect 2691 -1019 2753 -988
rect 2822 -990 2871 -965
rect 2916 -974 2942 -964
rect 2886 -990 2942 -974
rect 2785 -1004 2815 -996
rect 2822 -998 2932 -990
rect 2785 -1012 2830 -1004
rect 2517 -1030 2536 -1028
rect 2551 -1030 2597 -1028
rect 2517 -1046 2597 -1030
rect 2624 -1032 2659 -1019
rect 2700 -1022 2737 -1019
rect 2700 -1024 2742 -1022
rect 2629 -1035 2659 -1032
rect 2638 -1039 2645 -1035
rect 2645 -1040 2646 -1039
rect 2604 -1046 2614 -1040
rect 2363 -1054 2398 -1046
rect 2363 -1080 2364 -1054
rect 2371 -1080 2398 -1054
rect 2306 -1098 2336 -1084
rect 2363 -1088 2398 -1080
rect 2400 -1054 2441 -1046
rect 2400 -1080 2415 -1054
rect 2422 -1080 2441 -1054
rect 2505 -1058 2536 -1046
rect 2551 -1058 2654 -1046
rect 2666 -1056 2692 -1030
rect 2707 -1035 2737 -1024
rect 2769 -1028 2831 -1012
rect 2769 -1030 2815 -1028
rect 2769 -1046 2831 -1030
rect 2843 -1046 2849 -998
rect 2852 -1006 2932 -998
rect 2852 -1008 2871 -1006
rect 2886 -1008 2920 -1006
rect 2852 -1024 2932 -1008
rect 2852 -1046 2871 -1024
rect 2886 -1040 2916 -1024
rect 2944 -1030 2950 -956
rect 2953 -1030 2972 -886
rect 2987 -1030 2993 -886
rect 3002 -956 3015 -886
rect 3067 -890 3089 -886
rect 3060 -902 3077 -898
rect 3081 -900 3089 -898
rect 3079 -902 3089 -900
rect 3060 -912 3089 -902
rect 3142 -912 3158 -898
rect 3196 -902 3202 -900
rect 3209 -902 3317 -886
rect 3324 -902 3330 -900
rect 3338 -902 3353 -886
rect 3419 -892 3438 -889
rect 3060 -914 3158 -912
rect 3185 -914 3353 -902
rect 3368 -912 3384 -898
rect 3419 -911 3441 -892
rect 3451 -898 3467 -897
rect 3450 -900 3467 -898
rect 3451 -905 3467 -900
rect 3441 -912 3447 -911
rect 3450 -912 3479 -905
rect 3368 -913 3479 -912
rect 3368 -914 3485 -913
rect 3044 -922 3095 -914
rect 3142 -922 3176 -914
rect 3044 -934 3069 -922
rect 3076 -934 3095 -922
rect 3149 -924 3176 -922
rect 3185 -924 3406 -914
rect 3441 -917 3447 -914
rect 3149 -928 3406 -924
rect 3044 -942 3095 -934
rect 3142 -942 3406 -928
rect 3450 -922 3485 -914
rect 2996 -990 3015 -956
rect 3060 -950 3089 -942
rect 3060 -956 3077 -950
rect 3060 -958 3094 -956
rect 3142 -958 3158 -942
rect 3159 -952 3367 -942
rect 3368 -952 3384 -942
rect 3432 -946 3447 -931
rect 3450 -934 3451 -922
rect 3458 -934 3485 -922
rect 3450 -942 3485 -934
rect 3450 -943 3479 -942
rect 3170 -956 3384 -952
rect 3185 -958 3384 -956
rect 3419 -956 3432 -946
rect 3450 -956 3467 -943
rect 3419 -958 3467 -956
rect 3061 -962 3094 -958
rect 3057 -964 3094 -962
rect 3057 -965 3124 -964
rect 3057 -970 3088 -965
rect 3094 -970 3124 -965
rect 3057 -974 3124 -970
rect 3030 -977 3124 -974
rect 3030 -984 3079 -977
rect 3030 -990 3060 -984
rect 3079 -989 3084 -984
rect 2996 -1006 3076 -990
rect 3088 -998 3124 -977
rect 3185 -982 3374 -958
rect 3419 -959 3466 -958
rect 3432 -964 3466 -959
rect 3200 -985 3374 -982
rect 3193 -988 3374 -985
rect 3402 -965 3466 -964
rect 2996 -1008 3015 -1006
rect 3030 -1008 3064 -1006
rect 2996 -1024 3076 -1008
rect 2996 -1030 3015 -1024
rect 2712 -1056 2815 -1046
rect 2666 -1058 2815 -1056
rect 2836 -1058 2871 -1046
rect 2505 -1060 2667 -1058
rect 2517 -1080 2536 -1060
rect 2551 -1062 2581 -1060
rect 2400 -1088 2441 -1080
rect 2523 -1084 2536 -1080
rect 2588 -1076 2667 -1060
rect 2699 -1060 2871 -1058
rect 2699 -1076 2778 -1060
rect 2785 -1062 2815 -1060
rect 2363 -1098 2392 -1088
rect 2406 -1098 2435 -1088
rect 2450 -1098 2480 -1084
rect 2523 -1098 2566 -1084
rect 2588 -1088 2778 -1076
rect 2843 -1080 2849 -1060
rect 2573 -1098 2603 -1088
rect 2604 -1098 2762 -1088
rect 2766 -1098 2796 -1088
rect 2800 -1098 2830 -1084
rect 2858 -1098 2871 -1060
rect 2943 -1046 2972 -1030
rect 2986 -1046 3015 -1030
rect 3030 -1040 3060 -1024
rect 3088 -1046 3094 -998
rect 3097 -1004 3116 -998
rect 3131 -1004 3161 -996
rect 3097 -1012 3161 -1004
rect 3097 -1028 3177 -1012
rect 3193 -1019 3255 -988
rect 3271 -1019 3333 -988
rect 3402 -990 3451 -965
rect 3466 -990 3496 -972
rect 3365 -1004 3395 -996
rect 3402 -998 3512 -990
rect 3365 -1012 3410 -1004
rect 3097 -1030 3116 -1028
rect 3131 -1030 3177 -1028
rect 3097 -1046 3177 -1030
rect 3204 -1032 3239 -1019
rect 3280 -1022 3317 -1019
rect 3280 -1024 3322 -1022
rect 3209 -1035 3239 -1032
rect 3218 -1039 3225 -1035
rect 3225 -1040 3226 -1039
rect 3184 -1046 3194 -1040
rect 2943 -1054 2978 -1046
rect 2943 -1080 2944 -1054
rect 2951 -1080 2978 -1054
rect 2886 -1098 2916 -1084
rect 2943 -1088 2978 -1080
rect 2980 -1054 3021 -1046
rect 2980 -1080 2995 -1054
rect 3002 -1080 3021 -1054
rect 3085 -1058 3116 -1046
rect 3131 -1058 3234 -1046
rect 3246 -1056 3272 -1030
rect 3287 -1035 3317 -1024
rect 3349 -1028 3411 -1012
rect 3349 -1030 3395 -1028
rect 3349 -1046 3411 -1030
rect 3423 -1046 3429 -998
rect 3432 -1006 3512 -998
rect 3432 -1008 3451 -1006
rect 3466 -1008 3500 -1006
rect 3432 -1023 3512 -1008
rect 3432 -1024 3518 -1023
rect 3432 -1046 3451 -1024
rect 3466 -1040 3496 -1024
rect 3524 -1030 3530 -956
rect 3533 -1030 3552 -886
rect 3567 -1030 3573 -886
rect 3582 -956 3595 -886
rect 3647 -890 3669 -886
rect 3640 -902 3657 -898
rect 3661 -900 3669 -898
rect 3659 -902 3669 -900
rect 3640 -912 3669 -902
rect 3722 -912 3738 -898
rect 3776 -902 3782 -900
rect 3789 -902 3897 -886
rect 3904 -902 3910 -900
rect 3918 -902 3933 -886
rect 3999 -892 4018 -889
rect 3640 -914 3738 -912
rect 3765 -914 3933 -902
rect 3948 -912 3964 -898
rect 3999 -911 4021 -892
rect 4031 -898 4047 -897
rect 4030 -900 4047 -898
rect 4031 -905 4047 -900
rect 4021 -912 4027 -911
rect 4030 -912 4059 -905
rect 3948 -913 4059 -912
rect 3948 -914 4065 -913
rect 3624 -922 3675 -914
rect 3722 -922 3756 -914
rect 3624 -934 3649 -922
rect 3656 -934 3675 -922
rect 3729 -924 3756 -922
rect 3765 -924 3986 -914
rect 4021 -917 4027 -914
rect 3729 -928 3986 -924
rect 3624 -942 3675 -934
rect 3722 -942 3986 -928
rect 4030 -922 4065 -914
rect 3576 -990 3595 -956
rect 3640 -950 3669 -942
rect 3640 -956 3657 -950
rect 3640 -958 3674 -956
rect 3722 -958 3738 -942
rect 3739 -952 3947 -942
rect 3948 -952 3964 -942
rect 4012 -946 4027 -931
rect 4030 -934 4031 -922
rect 4038 -934 4065 -922
rect 4030 -942 4065 -934
rect 4030 -943 4059 -942
rect 3750 -956 3964 -952
rect 3765 -958 3964 -956
rect 3999 -956 4012 -946
rect 4030 -956 4047 -943
rect 3999 -958 4047 -956
rect 3641 -962 3674 -958
rect 3637 -964 3674 -962
rect 3637 -965 3704 -964
rect 3637 -970 3668 -965
rect 3674 -970 3704 -965
rect 3637 -974 3704 -970
rect 3610 -977 3704 -974
rect 3610 -984 3659 -977
rect 3610 -990 3640 -984
rect 3659 -989 3664 -984
rect 3576 -1006 3656 -990
rect 3668 -998 3704 -977
rect 3765 -982 3954 -958
rect 3999 -959 4046 -958
rect 4012 -964 4046 -959
rect 4086 -964 4102 -962
rect 3780 -985 3954 -982
rect 3773 -988 3954 -985
rect 3982 -965 4046 -964
rect 3576 -1008 3595 -1006
rect 3610 -1008 3644 -1006
rect 3576 -1024 3656 -1008
rect 3576 -1030 3595 -1024
rect 3292 -1056 3395 -1046
rect 3246 -1058 3395 -1056
rect 3416 -1058 3451 -1046
rect 3085 -1060 3247 -1058
rect 3097 -1080 3116 -1060
rect 3131 -1062 3161 -1060
rect 2980 -1088 3021 -1080
rect 3103 -1084 3116 -1080
rect 3168 -1076 3247 -1060
rect 3279 -1060 3451 -1058
rect 3279 -1076 3358 -1060
rect 3365 -1062 3395 -1060
rect 2943 -1098 2972 -1088
rect 2986 -1098 3015 -1088
rect 3030 -1098 3060 -1084
rect 3103 -1098 3146 -1084
rect 3168 -1088 3358 -1076
rect 3423 -1080 3429 -1060
rect 3153 -1098 3183 -1088
rect 3184 -1098 3342 -1088
rect 3346 -1098 3376 -1088
rect 3380 -1098 3410 -1084
rect 3438 -1098 3451 -1060
rect 3523 -1046 3552 -1030
rect 3566 -1046 3595 -1030
rect 3610 -1040 3640 -1024
rect 3668 -1046 3674 -998
rect 3677 -1004 3696 -998
rect 3711 -1004 3741 -996
rect 3677 -1012 3741 -1004
rect 3677 -1028 3757 -1012
rect 3773 -1019 3835 -988
rect 3851 -1019 3913 -988
rect 3982 -990 4031 -965
rect 4076 -974 4102 -964
rect 4046 -990 4102 -974
rect 3945 -1004 3975 -996
rect 3982 -998 4092 -990
rect 3945 -1012 3990 -1004
rect 3677 -1030 3696 -1028
rect 3711 -1030 3757 -1028
rect 3677 -1046 3757 -1030
rect 3784 -1032 3819 -1019
rect 3860 -1022 3897 -1019
rect 3860 -1024 3902 -1022
rect 3789 -1035 3819 -1032
rect 3798 -1039 3805 -1035
rect 3805 -1040 3806 -1039
rect 3764 -1046 3774 -1040
rect 3523 -1054 3558 -1046
rect 3523 -1080 3524 -1054
rect 3531 -1080 3558 -1054
rect 3466 -1098 3496 -1084
rect 3523 -1088 3558 -1080
rect 3560 -1054 3601 -1046
rect 3560 -1080 3575 -1054
rect 3582 -1080 3601 -1054
rect 3665 -1058 3696 -1046
rect 3711 -1058 3814 -1046
rect 3826 -1056 3852 -1030
rect 3867 -1035 3897 -1024
rect 3929 -1028 3991 -1012
rect 3929 -1030 3975 -1028
rect 3929 -1046 3991 -1030
rect 4003 -1046 4009 -998
rect 4012 -1006 4092 -998
rect 4012 -1008 4031 -1006
rect 4046 -1008 4080 -1006
rect 4012 -1024 4092 -1008
rect 4012 -1046 4031 -1024
rect 4046 -1040 4076 -1024
rect 4104 -1030 4110 -956
rect 4113 -1030 4132 -886
rect 4147 -1030 4153 -886
rect 4162 -956 4175 -886
rect 4227 -890 4249 -886
rect 4220 -902 4237 -898
rect 4241 -900 4249 -898
rect 4239 -902 4249 -900
rect 4220 -912 4249 -902
rect 4302 -912 4318 -898
rect 4356 -902 4362 -900
rect 4369 -902 4477 -886
rect 4484 -902 4490 -900
rect 4498 -902 4513 -886
rect 4579 -892 4598 -889
rect 4220 -914 4318 -912
rect 4345 -914 4513 -902
rect 4528 -912 4544 -898
rect 4579 -911 4601 -892
rect 4611 -898 4627 -897
rect 4610 -900 4627 -898
rect 4611 -905 4627 -900
rect 4601 -912 4607 -911
rect 4610 -912 4639 -905
rect 4528 -913 4639 -912
rect 4528 -914 4645 -913
rect 4204 -922 4255 -914
rect 4302 -922 4336 -914
rect 4204 -934 4229 -922
rect 4236 -934 4255 -922
rect 4309 -924 4336 -922
rect 4345 -924 4566 -914
rect 4601 -917 4607 -914
rect 4309 -928 4566 -924
rect 4204 -942 4255 -934
rect 4302 -942 4566 -928
rect 4610 -922 4645 -914
rect 4156 -990 4175 -956
rect 4220 -950 4249 -942
rect 4220 -956 4237 -950
rect 4220 -958 4254 -956
rect 4302 -958 4318 -942
rect 4319 -952 4527 -942
rect 4528 -952 4544 -942
rect 4592 -946 4607 -931
rect 4610 -934 4611 -922
rect 4618 -934 4645 -922
rect 4610 -942 4645 -934
rect 4610 -943 4639 -942
rect 4330 -956 4544 -952
rect 4345 -958 4544 -956
rect 4579 -956 4592 -946
rect 4610 -956 4627 -943
rect 4579 -958 4627 -956
rect 4221 -962 4254 -958
rect 4217 -964 4254 -962
rect 4217 -965 4284 -964
rect 4217 -970 4248 -965
rect 4254 -970 4284 -965
rect 4217 -974 4284 -970
rect 4190 -977 4284 -974
rect 4190 -984 4239 -977
rect 4190 -990 4220 -984
rect 4239 -989 4244 -984
rect 4156 -1006 4236 -990
rect 4248 -998 4284 -977
rect 4345 -982 4534 -958
rect 4579 -959 4626 -958
rect 4592 -964 4626 -959
rect 4360 -985 4534 -982
rect 4353 -988 4534 -985
rect 4562 -965 4626 -964
rect 4156 -1008 4175 -1006
rect 4190 -1008 4224 -1006
rect 4156 -1024 4236 -1008
rect 4156 -1030 4175 -1024
rect 3872 -1056 3975 -1046
rect 3826 -1058 3975 -1056
rect 3996 -1058 4031 -1046
rect 3665 -1060 3827 -1058
rect 3677 -1080 3696 -1060
rect 3711 -1062 3741 -1060
rect 3560 -1088 3601 -1080
rect 3683 -1084 3696 -1080
rect 3748 -1076 3827 -1060
rect 3859 -1060 4031 -1058
rect 3859 -1076 3938 -1060
rect 3945 -1062 3975 -1060
rect 3523 -1098 3552 -1088
rect 3566 -1098 3595 -1088
rect 3610 -1098 3640 -1084
rect 3683 -1098 3726 -1084
rect 3748 -1088 3938 -1076
rect 4003 -1080 4009 -1060
rect 3733 -1098 3763 -1088
rect 3764 -1098 3922 -1088
rect 3926 -1098 3956 -1088
rect 3960 -1098 3990 -1084
rect 4018 -1098 4031 -1060
rect 4103 -1046 4132 -1030
rect 4146 -1046 4175 -1030
rect 4190 -1040 4220 -1024
rect 4248 -1046 4254 -998
rect 4257 -1004 4276 -998
rect 4291 -1004 4321 -996
rect 4257 -1012 4321 -1004
rect 4257 -1028 4337 -1012
rect 4353 -1019 4415 -988
rect 4431 -1019 4493 -988
rect 4562 -990 4611 -965
rect 4626 -990 4656 -972
rect 4525 -1004 4555 -996
rect 4562 -998 4672 -990
rect 4525 -1012 4570 -1004
rect 4257 -1030 4276 -1028
rect 4291 -1030 4337 -1028
rect 4257 -1046 4337 -1030
rect 4364 -1032 4399 -1019
rect 4440 -1022 4477 -1019
rect 4440 -1024 4482 -1022
rect 4369 -1035 4399 -1032
rect 4378 -1039 4385 -1035
rect 4385 -1040 4386 -1039
rect 4344 -1046 4354 -1040
rect 4103 -1054 4138 -1046
rect 4103 -1080 4104 -1054
rect 4111 -1080 4138 -1054
rect 4046 -1098 4076 -1084
rect 4103 -1088 4138 -1080
rect 4140 -1054 4181 -1046
rect 4140 -1080 4155 -1054
rect 4162 -1080 4181 -1054
rect 4245 -1058 4276 -1046
rect 4291 -1058 4394 -1046
rect 4406 -1056 4432 -1030
rect 4447 -1035 4477 -1024
rect 4509 -1028 4571 -1012
rect 4509 -1030 4555 -1028
rect 4509 -1046 4571 -1030
rect 4583 -1046 4589 -998
rect 4592 -1006 4672 -998
rect 4592 -1008 4611 -1006
rect 4626 -1008 4660 -1006
rect 4592 -1023 4672 -1008
rect 4592 -1024 4678 -1023
rect 4592 -1046 4611 -1024
rect 4626 -1040 4656 -1024
rect 4684 -1030 4690 -956
rect 4693 -1030 4712 -886
rect 4727 -1030 4733 -886
rect 4742 -956 4755 -886
rect 4807 -890 4829 -886
rect 4800 -902 4817 -898
rect 4821 -900 4829 -898
rect 4819 -902 4829 -900
rect 4800 -912 4829 -902
rect 4882 -912 4898 -898
rect 4936 -902 4942 -900
rect 4949 -902 5057 -886
rect 5064 -902 5070 -900
rect 5078 -902 5093 -886
rect 5159 -892 5178 -889
rect 4800 -914 4898 -912
rect 4925 -914 5093 -902
rect 5108 -912 5124 -898
rect 5159 -911 5181 -892
rect 5191 -898 5207 -897
rect 5190 -900 5207 -898
rect 5191 -905 5207 -900
rect 5181 -912 5187 -911
rect 5190 -912 5219 -905
rect 5108 -913 5219 -912
rect 5108 -914 5225 -913
rect 4784 -922 4835 -914
rect 4882 -922 4916 -914
rect 4784 -934 4809 -922
rect 4816 -934 4835 -922
rect 4889 -924 4916 -922
rect 4925 -924 5146 -914
rect 5181 -917 5187 -914
rect 4889 -928 5146 -924
rect 4784 -942 4835 -934
rect 4882 -942 5146 -928
rect 5190 -922 5225 -914
rect 4736 -990 4755 -956
rect 4800 -950 4829 -942
rect 4800 -956 4817 -950
rect 4800 -958 4834 -956
rect 4882 -958 4898 -942
rect 4899 -952 5107 -942
rect 5108 -952 5124 -942
rect 5172 -946 5187 -931
rect 5190 -934 5191 -922
rect 5198 -934 5225 -922
rect 5190 -942 5225 -934
rect 5190 -943 5219 -942
rect 4910 -956 5124 -952
rect 4925 -958 5124 -956
rect 5159 -956 5172 -946
rect 5190 -956 5207 -943
rect 5159 -958 5207 -956
rect 4801 -962 4834 -958
rect 4797 -964 4834 -962
rect 4797 -965 4864 -964
rect 4797 -970 4828 -965
rect 4834 -970 4864 -965
rect 4797 -974 4864 -970
rect 4770 -977 4864 -974
rect 4770 -984 4819 -977
rect 4770 -990 4800 -984
rect 4819 -989 4824 -984
rect 4736 -1006 4816 -990
rect 4828 -998 4864 -977
rect 4925 -982 5114 -958
rect 5159 -959 5206 -958
rect 5172 -964 5206 -959
rect 5246 -964 5262 -962
rect 4940 -985 5114 -982
rect 4933 -988 5114 -985
rect 5142 -965 5206 -964
rect 4736 -1008 4755 -1006
rect 4770 -1008 4804 -1006
rect 4736 -1024 4816 -1008
rect 4736 -1030 4755 -1024
rect 4452 -1056 4555 -1046
rect 4406 -1058 4555 -1056
rect 4576 -1058 4611 -1046
rect 4245 -1060 4407 -1058
rect 4257 -1080 4276 -1060
rect 4291 -1062 4321 -1060
rect 4140 -1088 4181 -1080
rect 4263 -1084 4276 -1080
rect 4328 -1076 4407 -1060
rect 4439 -1060 4611 -1058
rect 4439 -1076 4518 -1060
rect 4525 -1062 4555 -1060
rect 4103 -1098 4132 -1088
rect 4146 -1098 4175 -1088
rect 4190 -1098 4220 -1084
rect 4263 -1098 4306 -1084
rect 4328 -1088 4518 -1076
rect 4583 -1080 4589 -1060
rect 4313 -1098 4343 -1088
rect 4344 -1098 4502 -1088
rect 4506 -1098 4536 -1088
rect 4540 -1098 4570 -1084
rect 4598 -1098 4611 -1060
rect 4683 -1046 4712 -1030
rect 4726 -1046 4755 -1030
rect 4770 -1040 4800 -1024
rect 4828 -1046 4834 -998
rect 4837 -1004 4856 -998
rect 4871 -1004 4901 -996
rect 4837 -1012 4901 -1004
rect 4837 -1028 4917 -1012
rect 4933 -1019 4995 -988
rect 5011 -1019 5073 -988
rect 5142 -990 5191 -965
rect 5236 -974 5262 -964
rect 5206 -990 5262 -974
rect 5105 -1004 5135 -996
rect 5142 -998 5252 -990
rect 5105 -1012 5150 -1004
rect 4837 -1030 4856 -1028
rect 4871 -1030 4917 -1028
rect 4837 -1046 4917 -1030
rect 4944 -1032 4979 -1019
rect 5020 -1022 5057 -1019
rect 5020 -1024 5062 -1022
rect 4949 -1035 4979 -1032
rect 4958 -1039 4965 -1035
rect 4965 -1040 4966 -1039
rect 4924 -1046 4934 -1040
rect 4683 -1054 4718 -1046
rect 4683 -1080 4684 -1054
rect 4691 -1080 4718 -1054
rect 4626 -1098 4656 -1084
rect 4683 -1088 4718 -1080
rect 4720 -1054 4761 -1046
rect 4720 -1080 4735 -1054
rect 4742 -1080 4761 -1054
rect 4825 -1058 4856 -1046
rect 4871 -1058 4974 -1046
rect 4986 -1056 5012 -1030
rect 5027 -1035 5057 -1024
rect 5089 -1028 5151 -1012
rect 5089 -1030 5135 -1028
rect 5089 -1046 5151 -1030
rect 5163 -1046 5169 -998
rect 5172 -1006 5252 -998
rect 5172 -1008 5191 -1006
rect 5206 -1008 5240 -1006
rect 5172 -1024 5252 -1008
rect 5172 -1046 5191 -1024
rect 5206 -1040 5236 -1024
rect 5264 -1030 5270 -956
rect 5273 -1030 5292 -886
rect 5307 -1030 5313 -886
rect 5322 -956 5335 -886
rect 5387 -890 5409 -886
rect 5380 -902 5397 -898
rect 5401 -900 5409 -898
rect 5399 -902 5409 -900
rect 5380 -912 5409 -902
rect 5462 -912 5478 -898
rect 5516 -902 5522 -900
rect 5529 -902 5637 -886
rect 5644 -902 5650 -900
rect 5658 -902 5673 -886
rect 5739 -892 5758 -889
rect 5380 -914 5478 -912
rect 5505 -914 5673 -902
rect 5688 -912 5704 -898
rect 5739 -911 5761 -892
rect 5771 -898 5787 -897
rect 5770 -900 5787 -898
rect 5771 -905 5787 -900
rect 5761 -912 5767 -911
rect 5770 -912 5799 -905
rect 5688 -913 5799 -912
rect 5688 -914 5805 -913
rect 5364 -922 5415 -914
rect 5462 -922 5496 -914
rect 5364 -934 5389 -922
rect 5396 -934 5415 -922
rect 5469 -924 5496 -922
rect 5505 -924 5726 -914
rect 5761 -917 5767 -914
rect 5469 -928 5726 -924
rect 5364 -942 5415 -934
rect 5462 -942 5726 -928
rect 5770 -922 5805 -914
rect 5316 -990 5335 -956
rect 5380 -950 5409 -942
rect 5380 -956 5397 -950
rect 5380 -958 5414 -956
rect 5462 -958 5478 -942
rect 5479 -952 5687 -942
rect 5688 -952 5704 -942
rect 5752 -946 5767 -931
rect 5770 -934 5771 -922
rect 5778 -934 5805 -922
rect 5770 -942 5805 -934
rect 5770 -943 5799 -942
rect 5490 -956 5704 -952
rect 5505 -958 5704 -956
rect 5739 -956 5752 -946
rect 5770 -956 5787 -943
rect 5739 -958 5787 -956
rect 5381 -962 5414 -958
rect 5377 -964 5414 -962
rect 5377 -965 5444 -964
rect 5377 -970 5408 -965
rect 5414 -970 5444 -965
rect 5377 -974 5444 -970
rect 5350 -977 5444 -974
rect 5350 -984 5399 -977
rect 5350 -990 5380 -984
rect 5399 -989 5404 -984
rect 5316 -1006 5396 -990
rect 5408 -998 5444 -977
rect 5505 -982 5694 -958
rect 5739 -959 5786 -958
rect 5752 -964 5786 -959
rect 5520 -985 5694 -982
rect 5513 -988 5694 -985
rect 5722 -965 5786 -964
rect 5316 -1008 5335 -1006
rect 5350 -1008 5384 -1006
rect 5316 -1024 5396 -1008
rect 5316 -1030 5335 -1024
rect 5032 -1056 5135 -1046
rect 4986 -1058 5135 -1056
rect 5156 -1058 5191 -1046
rect 4825 -1060 4987 -1058
rect 4837 -1080 4856 -1060
rect 4871 -1062 4901 -1060
rect 4720 -1088 4761 -1080
rect 4843 -1084 4856 -1080
rect 4908 -1076 4987 -1060
rect 5019 -1060 5191 -1058
rect 5019 -1076 5098 -1060
rect 5105 -1062 5135 -1060
rect 4683 -1098 4712 -1088
rect 4726 -1098 4755 -1088
rect 4770 -1098 4800 -1084
rect 4843 -1098 4886 -1084
rect 4908 -1088 5098 -1076
rect 5163 -1080 5169 -1060
rect 4893 -1098 4923 -1088
rect 4924 -1098 5082 -1088
rect 5086 -1098 5116 -1088
rect 5120 -1098 5150 -1084
rect 5178 -1098 5191 -1060
rect 5263 -1046 5292 -1030
rect 5306 -1046 5335 -1030
rect 5350 -1040 5380 -1024
rect 5408 -1046 5414 -998
rect 5417 -1004 5436 -998
rect 5451 -1004 5481 -996
rect 5417 -1012 5481 -1004
rect 5417 -1028 5497 -1012
rect 5513 -1019 5575 -988
rect 5591 -1019 5653 -988
rect 5722 -990 5771 -965
rect 5786 -990 5816 -972
rect 5685 -1004 5715 -996
rect 5722 -998 5832 -990
rect 5685 -1012 5730 -1004
rect 5417 -1030 5436 -1028
rect 5451 -1030 5497 -1028
rect 5417 -1046 5497 -1030
rect 5524 -1032 5559 -1019
rect 5600 -1022 5637 -1019
rect 5600 -1024 5642 -1022
rect 5529 -1035 5559 -1032
rect 5538 -1039 5545 -1035
rect 5545 -1040 5546 -1039
rect 5504 -1046 5514 -1040
rect 5263 -1054 5298 -1046
rect 5263 -1080 5264 -1054
rect 5271 -1080 5298 -1054
rect 5206 -1098 5236 -1084
rect 5263 -1088 5298 -1080
rect 5300 -1054 5341 -1046
rect 5300 -1080 5315 -1054
rect 5322 -1080 5341 -1054
rect 5405 -1058 5436 -1046
rect 5451 -1058 5554 -1046
rect 5566 -1056 5592 -1030
rect 5607 -1035 5637 -1024
rect 5669 -1028 5731 -1012
rect 5669 -1030 5715 -1028
rect 5669 -1046 5731 -1030
rect 5743 -1046 5749 -998
rect 5752 -1006 5832 -998
rect 5752 -1008 5771 -1006
rect 5786 -1008 5820 -1006
rect 5752 -1023 5832 -1008
rect 5752 -1024 5838 -1023
rect 5752 -1046 5771 -1024
rect 5786 -1040 5816 -1024
rect 5844 -1030 5850 -956
rect 5853 -1030 5872 -886
rect 5887 -1030 5893 -886
rect 5902 -956 5915 -886
rect 5967 -890 5989 -886
rect 5960 -902 5977 -898
rect 5981 -900 5989 -898
rect 5979 -902 5989 -900
rect 5960 -912 5989 -902
rect 6042 -912 6058 -898
rect 6096 -902 6102 -900
rect 6109 -902 6217 -886
rect 6224 -902 6230 -900
rect 6238 -902 6253 -886
rect 6319 -892 6338 -889
rect 5960 -914 6058 -912
rect 6085 -914 6253 -902
rect 6268 -912 6284 -898
rect 6319 -911 6341 -892
rect 6351 -898 6367 -897
rect 6350 -900 6367 -898
rect 6351 -905 6367 -900
rect 6341 -912 6347 -911
rect 6350 -912 6379 -905
rect 6268 -913 6379 -912
rect 6268 -914 6385 -913
rect 5944 -922 5995 -914
rect 6042 -922 6076 -914
rect 5944 -934 5969 -922
rect 5976 -934 5995 -922
rect 6049 -924 6076 -922
rect 6085 -924 6306 -914
rect 6341 -917 6347 -914
rect 6049 -928 6306 -924
rect 5944 -942 5995 -934
rect 6042 -942 6306 -928
rect 6350 -922 6385 -914
rect 5896 -990 5915 -956
rect 5960 -950 5989 -942
rect 5960 -956 5977 -950
rect 5960 -958 5994 -956
rect 6042 -958 6058 -942
rect 6059 -952 6267 -942
rect 6268 -952 6284 -942
rect 6332 -946 6347 -931
rect 6350 -934 6351 -922
rect 6358 -934 6385 -922
rect 6350 -942 6385 -934
rect 6350 -943 6379 -942
rect 6070 -956 6284 -952
rect 6085 -958 6284 -956
rect 6319 -956 6332 -946
rect 6350 -956 6367 -943
rect 6319 -958 6367 -956
rect 5961 -962 5994 -958
rect 5957 -964 5994 -962
rect 5957 -965 6024 -964
rect 5957 -970 5988 -965
rect 5994 -970 6024 -965
rect 5957 -974 6024 -970
rect 5930 -977 6024 -974
rect 5930 -984 5979 -977
rect 5930 -990 5960 -984
rect 5979 -989 5984 -984
rect 5896 -1006 5976 -990
rect 5988 -998 6024 -977
rect 6085 -982 6274 -958
rect 6319 -959 6366 -958
rect 6332 -964 6366 -959
rect 6100 -985 6274 -982
rect 6093 -988 6274 -985
rect 6302 -965 6366 -964
rect 5896 -1008 5915 -1006
rect 5930 -1008 5964 -1006
rect 5896 -1024 5976 -1008
rect 5896 -1030 5915 -1024
rect 5612 -1056 5715 -1046
rect 5566 -1058 5715 -1056
rect 5736 -1058 5771 -1046
rect 5405 -1060 5567 -1058
rect 5417 -1080 5436 -1060
rect 5451 -1062 5481 -1060
rect 5300 -1088 5341 -1080
rect 5423 -1084 5436 -1080
rect 5488 -1076 5567 -1060
rect 5599 -1060 5771 -1058
rect 5599 -1076 5678 -1060
rect 5685 -1062 5715 -1060
rect 5263 -1098 5292 -1088
rect 5306 -1098 5335 -1088
rect 5350 -1098 5380 -1084
rect 5423 -1098 5466 -1084
rect 5488 -1088 5678 -1076
rect 5743 -1080 5749 -1060
rect 5473 -1098 5503 -1088
rect 5504 -1098 5662 -1088
rect 5666 -1098 5696 -1088
rect 5700 -1098 5730 -1084
rect 5758 -1098 5771 -1060
rect 5843 -1046 5872 -1030
rect 5886 -1046 5915 -1030
rect 5930 -1040 5960 -1024
rect 5988 -1046 5994 -998
rect 5997 -1004 6016 -998
rect 6031 -1004 6061 -996
rect 5997 -1012 6061 -1004
rect 5997 -1028 6077 -1012
rect 6093 -1019 6155 -988
rect 6171 -1019 6233 -988
rect 6302 -990 6351 -965
rect 6366 -990 6396 -974
rect 6265 -1004 6295 -996
rect 6302 -998 6412 -990
rect 6265 -1012 6310 -1004
rect 5997 -1030 6016 -1028
rect 6031 -1030 6077 -1028
rect 5997 -1046 6077 -1030
rect 6104 -1032 6139 -1019
rect 6180 -1022 6217 -1019
rect 6180 -1024 6222 -1022
rect 6109 -1035 6139 -1032
rect 6118 -1039 6125 -1035
rect 6125 -1040 6126 -1039
rect 6084 -1046 6094 -1040
rect 5843 -1054 5878 -1046
rect 5843 -1080 5844 -1054
rect 5851 -1080 5878 -1054
rect 5786 -1098 5816 -1084
rect 5843 -1088 5878 -1080
rect 5880 -1054 5921 -1046
rect 5880 -1080 5895 -1054
rect 5902 -1080 5921 -1054
rect 5985 -1058 6016 -1046
rect 6031 -1058 6134 -1046
rect 6146 -1056 6172 -1030
rect 6187 -1035 6217 -1024
rect 6249 -1028 6311 -1012
rect 6249 -1030 6295 -1028
rect 6249 -1046 6311 -1030
rect 6323 -1046 6329 -998
rect 6332 -1006 6412 -998
rect 6332 -1008 6351 -1006
rect 6366 -1008 6400 -1006
rect 6332 -1024 6412 -1008
rect 6332 -1046 6351 -1024
rect 6366 -1040 6396 -1024
rect 6424 -1030 6430 -956
rect 6439 -1030 6452 -886
rect 6192 -1056 6295 -1046
rect 6146 -1058 6295 -1056
rect 6316 -1058 6351 -1046
rect 5985 -1060 6147 -1058
rect 5997 -1080 6016 -1060
rect 6031 -1062 6061 -1060
rect 5880 -1088 5921 -1080
rect 6003 -1084 6016 -1080
rect 6068 -1076 6147 -1060
rect 6179 -1060 6351 -1058
rect 6179 -1076 6258 -1060
rect 6265 -1062 6295 -1060
rect 5843 -1098 5872 -1088
rect 5886 -1098 5915 -1088
rect 5930 -1098 5960 -1084
rect 6003 -1098 6046 -1084
rect 6068 -1088 6258 -1076
rect 6323 -1080 6329 -1060
rect 6053 -1098 6083 -1088
rect 6084 -1098 6242 -1088
rect 6246 -1098 6276 -1088
rect 6280 -1098 6310 -1084
rect 6338 -1098 6351 -1060
rect 6423 -1046 6452 -1030
rect 6423 -1054 6458 -1046
rect 6423 -1080 6424 -1054
rect 6431 -1080 6458 -1054
rect 6366 -1098 6396 -1084
rect 6423 -1088 6458 -1080
rect 6423 -1098 6452 -1088
rect -541 -1112 6452 -1098
rect -478 -1142 -465 -1112
rect -450 -1126 -420 -1112
rect -377 -1126 -334 -1112
rect -327 -1126 -107 -1112
rect -100 -1126 -70 -1112
rect -410 -1140 -395 -1128
rect -376 -1140 -363 -1126
rect -295 -1130 -142 -1126
rect -413 -1142 -391 -1140
rect -313 -1142 -121 -1130
rect -42 -1142 -29 -1112
rect -14 -1126 16 -1112
rect 53 -1142 72 -1112
rect 87 -1142 93 -1112
rect 102 -1142 115 -1112
rect 130 -1126 160 -1112
rect 203 -1126 246 -1112
rect 253 -1126 473 -1112
rect 480 -1126 510 -1112
rect 170 -1140 185 -1128
rect 204 -1140 217 -1126
rect 285 -1130 438 -1126
rect 167 -1142 189 -1140
rect 267 -1142 459 -1130
rect 538 -1142 551 -1112
rect 566 -1126 596 -1112
rect 633 -1142 652 -1112
rect 667 -1142 673 -1112
rect 682 -1142 695 -1112
rect 710 -1126 740 -1112
rect 783 -1126 826 -1112
rect 833 -1126 1053 -1112
rect 1060 -1126 1090 -1112
rect 750 -1140 765 -1128
rect 784 -1140 797 -1126
rect 865 -1130 1018 -1126
rect 747 -1142 769 -1140
rect 847 -1142 1039 -1130
rect 1118 -1142 1131 -1112
rect 1146 -1126 1176 -1112
rect 1213 -1142 1232 -1112
rect 1247 -1142 1253 -1112
rect 1262 -1142 1275 -1112
rect 1290 -1126 1320 -1112
rect 1363 -1126 1406 -1112
rect 1413 -1126 1633 -1112
rect 1640 -1126 1670 -1112
rect 1330 -1140 1345 -1128
rect 1364 -1140 1377 -1126
rect 1445 -1130 1598 -1126
rect 1327 -1142 1349 -1140
rect 1427 -1142 1619 -1130
rect 1698 -1142 1711 -1112
rect 1726 -1126 1756 -1112
rect 1793 -1142 1812 -1112
rect 1827 -1142 1833 -1112
rect 1842 -1142 1855 -1112
rect 1870 -1126 1900 -1112
rect 1943 -1126 1986 -1112
rect 1993 -1126 2213 -1112
rect 2220 -1126 2250 -1112
rect 1910 -1140 1925 -1128
rect 1944 -1140 1957 -1126
rect 2025 -1130 2178 -1126
rect 1907 -1142 1929 -1140
rect 2007 -1142 2199 -1130
rect 2278 -1142 2291 -1112
rect 2306 -1126 2336 -1112
rect 2373 -1142 2392 -1112
rect 2407 -1142 2413 -1112
rect 2422 -1142 2435 -1112
rect 2450 -1126 2480 -1112
rect 2523 -1126 2566 -1112
rect 2573 -1126 2793 -1112
rect 2800 -1126 2830 -1112
rect 2490 -1140 2505 -1128
rect 2524 -1140 2537 -1126
rect 2605 -1130 2758 -1126
rect 2487 -1142 2509 -1140
rect 2587 -1142 2779 -1130
rect 2858 -1142 2871 -1112
rect 2886 -1126 2916 -1112
rect 2953 -1142 2972 -1112
rect 2987 -1142 2993 -1112
rect 3002 -1142 3015 -1112
rect 3030 -1126 3060 -1112
rect 3103 -1126 3146 -1112
rect 3153 -1126 3373 -1112
rect 3380 -1126 3410 -1112
rect 3070 -1140 3085 -1128
rect 3104 -1140 3117 -1126
rect 3185 -1130 3338 -1126
rect 3067 -1142 3089 -1140
rect 3167 -1142 3359 -1130
rect 3438 -1142 3451 -1112
rect 3466 -1126 3496 -1112
rect 3533 -1142 3552 -1112
rect 3567 -1142 3573 -1112
rect 3582 -1142 3595 -1112
rect 3610 -1126 3640 -1112
rect 3683 -1126 3726 -1112
rect 3733 -1126 3953 -1112
rect 3960 -1126 3990 -1112
rect 3650 -1140 3665 -1128
rect 3684 -1140 3697 -1126
rect 3765 -1130 3918 -1126
rect 3647 -1142 3669 -1140
rect 3747 -1142 3939 -1130
rect 4018 -1142 4031 -1112
rect 4046 -1126 4076 -1112
rect 4113 -1142 4132 -1112
rect 4147 -1142 4153 -1112
rect 4162 -1142 4175 -1112
rect 4190 -1126 4220 -1112
rect 4263 -1126 4306 -1112
rect 4313 -1126 4533 -1112
rect 4540 -1126 4570 -1112
rect 4230 -1140 4245 -1128
rect 4264 -1140 4277 -1126
rect 4345 -1130 4498 -1126
rect 4227 -1142 4249 -1140
rect 4327 -1142 4519 -1130
rect 4598 -1142 4611 -1112
rect 4626 -1126 4656 -1112
rect 4693 -1142 4712 -1112
rect 4727 -1142 4733 -1112
rect 4742 -1142 4755 -1112
rect 4770 -1126 4800 -1112
rect 4843 -1126 4886 -1112
rect 4893 -1126 5113 -1112
rect 5120 -1126 5150 -1112
rect 4810 -1140 4825 -1128
rect 4844 -1140 4857 -1126
rect 4925 -1130 5078 -1126
rect 4807 -1142 4829 -1140
rect 4907 -1142 5099 -1130
rect 5178 -1142 5191 -1112
rect 5206 -1126 5236 -1112
rect 5273 -1142 5292 -1112
rect 5307 -1142 5313 -1112
rect 5322 -1142 5335 -1112
rect 5350 -1126 5380 -1112
rect 5423 -1126 5466 -1112
rect 5473 -1126 5693 -1112
rect 5700 -1126 5730 -1112
rect 5390 -1140 5405 -1128
rect 5424 -1140 5437 -1126
rect 5505 -1130 5658 -1126
rect 5387 -1142 5409 -1140
rect 5487 -1142 5679 -1130
rect 5758 -1142 5771 -1112
rect 5786 -1126 5816 -1112
rect 5853 -1142 5872 -1112
rect 5887 -1142 5893 -1112
rect 5902 -1142 5915 -1112
rect 5930 -1126 5960 -1112
rect 6003 -1126 6046 -1112
rect 6053 -1126 6273 -1112
rect 6280 -1126 6310 -1112
rect 5970 -1140 5985 -1128
rect 6004 -1140 6017 -1126
rect 6085 -1130 6238 -1126
rect 5967 -1142 5989 -1140
rect 6067 -1142 6259 -1130
rect 6338 -1142 6351 -1112
rect 6366 -1126 6396 -1112
rect 6439 -1142 6452 -1112
rect -541 -1156 6452 -1142
rect -478 -1226 -465 -1156
rect -413 -1160 -391 -1156
rect -420 -1172 -403 -1168
rect -399 -1170 -391 -1168
rect -401 -1172 -391 -1170
rect -420 -1182 -391 -1172
rect -338 -1182 -322 -1168
rect -284 -1172 -278 -1170
rect -271 -1172 -163 -1156
rect -156 -1172 -150 -1170
rect -142 -1172 -127 -1156
rect -61 -1162 -42 -1159
rect -420 -1184 -322 -1182
rect -295 -1184 -127 -1172
rect -112 -1182 -96 -1168
rect -61 -1181 -39 -1162
rect -29 -1168 -13 -1167
rect -30 -1170 -13 -1168
rect -29 -1175 -13 -1170
rect -39 -1182 -33 -1181
rect -30 -1182 -1 -1175
rect -112 -1183 -1 -1182
rect -112 -1184 5 -1183
rect -436 -1192 -385 -1184
rect -338 -1192 -304 -1184
rect -436 -1204 -411 -1192
rect -404 -1204 -385 -1192
rect -331 -1194 -304 -1192
rect -295 -1194 -74 -1184
rect -39 -1187 -33 -1184
rect -331 -1198 -74 -1194
rect -436 -1212 -385 -1204
rect -338 -1212 -74 -1198
rect -30 -1192 5 -1184
rect -484 -1260 -465 -1226
rect -420 -1220 -391 -1212
rect -420 -1226 -403 -1220
rect -420 -1228 -386 -1226
rect -338 -1228 -322 -1212
rect -321 -1222 -113 -1212
rect -112 -1222 -96 -1212
rect -48 -1216 -33 -1201
rect -30 -1204 -29 -1192
rect -22 -1204 5 -1192
rect -30 -1212 5 -1204
rect -30 -1213 -1 -1212
rect -310 -1226 -96 -1222
rect -295 -1228 -96 -1226
rect -61 -1226 -48 -1216
rect -30 -1226 -13 -1213
rect -61 -1228 -13 -1226
rect -419 -1232 -386 -1228
rect -423 -1234 -386 -1232
rect -423 -1235 -356 -1234
rect -423 -1240 -392 -1235
rect -386 -1240 -356 -1235
rect -423 -1244 -356 -1240
rect -450 -1247 -356 -1244
rect -450 -1254 -401 -1247
rect -450 -1260 -420 -1254
rect -401 -1259 -396 -1254
rect -484 -1276 -404 -1260
rect -392 -1268 -356 -1247
rect -295 -1252 -106 -1228
rect -61 -1229 -14 -1228
rect -48 -1234 -14 -1229
rect -280 -1255 -106 -1252
rect -287 -1258 -106 -1255
rect -78 -1235 -14 -1234
rect -484 -1278 -465 -1276
rect -450 -1278 -416 -1276
rect -484 -1294 -404 -1278
rect -484 -1300 -465 -1294
rect -494 -1316 -465 -1300
rect -450 -1310 -420 -1294
rect -392 -1316 -386 -1268
rect -383 -1274 -364 -1268
rect -349 -1274 -319 -1266
rect -383 -1282 -319 -1274
rect -383 -1298 -303 -1282
rect -287 -1289 -225 -1258
rect -209 -1289 -147 -1258
rect -78 -1260 -29 -1235
rect -14 -1260 16 -1242
rect -115 -1274 -85 -1266
rect -78 -1268 32 -1260
rect -115 -1282 -70 -1274
rect -383 -1300 -364 -1298
rect -349 -1300 -303 -1298
rect -383 -1316 -303 -1300
rect -276 -1302 -241 -1289
rect -200 -1292 -163 -1289
rect -200 -1294 -158 -1292
rect -271 -1305 -241 -1302
rect -262 -1309 -255 -1305
rect -255 -1310 -254 -1309
rect -296 -1316 -286 -1310
rect -500 -1324 -459 -1316
rect -500 -1350 -485 -1324
rect -478 -1350 -459 -1324
rect -395 -1328 -364 -1316
rect -349 -1328 -246 -1316
rect -234 -1326 -208 -1300
rect -193 -1305 -163 -1294
rect -131 -1298 -69 -1282
rect -131 -1300 -85 -1298
rect -131 -1316 -69 -1300
rect -57 -1316 -51 -1268
rect -48 -1276 32 -1268
rect -48 -1278 -29 -1276
rect -14 -1278 20 -1276
rect -48 -1293 32 -1278
rect -48 -1294 38 -1293
rect -48 -1316 -29 -1294
rect -14 -1310 16 -1294
rect 44 -1300 50 -1226
rect 53 -1300 72 -1156
rect 87 -1300 93 -1156
rect 102 -1226 115 -1156
rect 167 -1160 189 -1156
rect 160 -1172 177 -1168
rect 181 -1170 189 -1168
rect 179 -1172 189 -1170
rect 160 -1182 189 -1172
rect 242 -1182 258 -1168
rect 296 -1172 302 -1170
rect 309 -1172 417 -1156
rect 424 -1172 430 -1170
rect 438 -1172 453 -1156
rect 519 -1162 538 -1159
rect 160 -1184 258 -1182
rect 285 -1184 453 -1172
rect 468 -1182 484 -1168
rect 519 -1181 541 -1162
rect 551 -1168 567 -1167
rect 550 -1170 567 -1168
rect 551 -1175 567 -1170
rect 541 -1182 547 -1181
rect 550 -1182 579 -1175
rect 468 -1183 579 -1182
rect 468 -1184 585 -1183
rect 144 -1192 195 -1184
rect 242 -1192 276 -1184
rect 144 -1204 169 -1192
rect 176 -1204 195 -1192
rect 249 -1194 276 -1192
rect 285 -1194 506 -1184
rect 541 -1187 547 -1184
rect 249 -1198 506 -1194
rect 144 -1212 195 -1204
rect 242 -1212 506 -1198
rect 550 -1192 585 -1184
rect 96 -1260 115 -1226
rect 160 -1220 189 -1212
rect 160 -1226 177 -1220
rect 160 -1228 194 -1226
rect 242 -1228 258 -1212
rect 259 -1222 467 -1212
rect 468 -1222 484 -1212
rect 532 -1216 547 -1201
rect 550 -1204 551 -1192
rect 558 -1204 585 -1192
rect 550 -1212 585 -1204
rect 550 -1213 579 -1212
rect 270 -1226 484 -1222
rect 285 -1228 484 -1226
rect 519 -1226 532 -1216
rect 550 -1226 567 -1213
rect 519 -1228 567 -1226
rect 161 -1232 194 -1228
rect 157 -1234 194 -1232
rect 157 -1235 224 -1234
rect 157 -1240 188 -1235
rect 194 -1240 224 -1235
rect 157 -1244 224 -1240
rect 130 -1247 224 -1244
rect 130 -1254 179 -1247
rect 130 -1260 160 -1254
rect 179 -1259 184 -1254
rect 96 -1276 176 -1260
rect 188 -1268 224 -1247
rect 285 -1252 474 -1228
rect 519 -1229 566 -1228
rect 532 -1234 566 -1229
rect 606 -1234 622 -1232
rect 300 -1255 474 -1252
rect 293 -1258 474 -1255
rect 502 -1235 566 -1234
rect 96 -1278 115 -1276
rect 130 -1278 164 -1276
rect 96 -1294 176 -1278
rect 96 -1300 115 -1294
rect -188 -1326 -85 -1316
rect -234 -1328 -85 -1326
rect -64 -1328 -29 -1316
rect -395 -1330 -233 -1328
rect -383 -1348 -364 -1330
rect -349 -1332 -319 -1330
rect -500 -1358 -459 -1350
rect -376 -1354 -364 -1348
rect -312 -1346 -233 -1330
rect -201 -1330 -29 -1328
rect -201 -1346 -122 -1330
rect -115 -1332 -85 -1330
rect -494 -1368 -465 -1358
rect -450 -1368 -420 -1354
rect -376 -1368 -334 -1354
rect -312 -1358 -122 -1346
rect -57 -1350 -51 -1330
rect -327 -1368 -297 -1358
rect -296 -1368 -138 -1358
rect -134 -1368 -104 -1358
rect -100 -1368 -70 -1354
rect -42 -1368 -29 -1330
rect 43 -1316 72 -1300
rect 86 -1316 115 -1300
rect 130 -1310 160 -1294
rect 188 -1316 194 -1268
rect 197 -1274 216 -1268
rect 231 -1274 261 -1266
rect 197 -1282 261 -1274
rect 197 -1298 277 -1282
rect 293 -1289 355 -1258
rect 371 -1289 433 -1258
rect 502 -1260 551 -1235
rect 596 -1244 622 -1234
rect 566 -1260 622 -1244
rect 465 -1274 495 -1266
rect 502 -1268 612 -1260
rect 465 -1282 510 -1274
rect 197 -1300 216 -1298
rect 231 -1300 277 -1298
rect 197 -1316 277 -1300
rect 304 -1302 339 -1289
rect 380 -1292 417 -1289
rect 380 -1294 422 -1292
rect 309 -1305 339 -1302
rect 318 -1309 325 -1305
rect 325 -1310 326 -1309
rect 284 -1316 294 -1310
rect 43 -1324 78 -1316
rect 43 -1350 44 -1324
rect 51 -1350 78 -1324
rect -14 -1368 16 -1354
rect 43 -1358 78 -1350
rect 80 -1324 121 -1316
rect 80 -1350 95 -1324
rect 102 -1350 121 -1324
rect 185 -1328 216 -1316
rect 231 -1328 334 -1316
rect 346 -1326 372 -1300
rect 387 -1305 417 -1294
rect 449 -1298 511 -1282
rect 449 -1300 495 -1298
rect 449 -1316 511 -1300
rect 523 -1316 529 -1268
rect 532 -1276 612 -1268
rect 532 -1278 551 -1276
rect 566 -1278 600 -1276
rect 532 -1294 612 -1278
rect 532 -1316 551 -1294
rect 566 -1310 596 -1294
rect 624 -1300 630 -1226
rect 633 -1300 652 -1156
rect 667 -1300 673 -1156
rect 682 -1226 695 -1156
rect 747 -1160 769 -1156
rect 740 -1172 757 -1168
rect 761 -1170 769 -1168
rect 759 -1172 769 -1170
rect 740 -1182 769 -1172
rect 822 -1182 838 -1168
rect 876 -1172 882 -1170
rect 889 -1172 997 -1156
rect 1004 -1172 1010 -1170
rect 1018 -1172 1033 -1156
rect 1099 -1162 1118 -1159
rect 740 -1184 838 -1182
rect 865 -1184 1033 -1172
rect 1048 -1182 1064 -1168
rect 1099 -1181 1121 -1162
rect 1131 -1168 1147 -1167
rect 1130 -1170 1147 -1168
rect 1131 -1175 1147 -1170
rect 1121 -1182 1127 -1181
rect 1130 -1182 1159 -1175
rect 1048 -1183 1159 -1182
rect 1048 -1184 1165 -1183
rect 724 -1192 775 -1184
rect 822 -1192 856 -1184
rect 724 -1204 749 -1192
rect 756 -1204 775 -1192
rect 829 -1194 856 -1192
rect 865 -1194 1086 -1184
rect 1121 -1187 1127 -1184
rect 829 -1198 1086 -1194
rect 724 -1212 775 -1204
rect 822 -1212 1086 -1198
rect 1130 -1192 1165 -1184
rect 676 -1260 695 -1226
rect 740 -1220 769 -1212
rect 740 -1226 757 -1220
rect 740 -1228 774 -1226
rect 822 -1228 838 -1212
rect 839 -1222 1047 -1212
rect 1048 -1222 1064 -1212
rect 1112 -1216 1127 -1201
rect 1130 -1204 1131 -1192
rect 1138 -1204 1165 -1192
rect 1130 -1212 1165 -1204
rect 1130 -1213 1159 -1212
rect 850 -1226 1064 -1222
rect 865 -1228 1064 -1226
rect 1099 -1226 1112 -1216
rect 1130 -1226 1147 -1213
rect 1099 -1228 1147 -1226
rect 741 -1232 774 -1228
rect 737 -1234 774 -1232
rect 737 -1235 804 -1234
rect 737 -1240 768 -1235
rect 774 -1240 804 -1235
rect 737 -1244 804 -1240
rect 710 -1247 804 -1244
rect 710 -1254 759 -1247
rect 710 -1260 740 -1254
rect 759 -1259 764 -1254
rect 676 -1276 756 -1260
rect 768 -1268 804 -1247
rect 865 -1252 1054 -1228
rect 1099 -1229 1146 -1228
rect 1112 -1234 1146 -1229
rect 880 -1255 1054 -1252
rect 873 -1258 1054 -1255
rect 1082 -1235 1146 -1234
rect 676 -1278 695 -1276
rect 710 -1278 744 -1276
rect 676 -1294 756 -1278
rect 676 -1300 695 -1294
rect 392 -1326 495 -1316
rect 346 -1328 495 -1326
rect 516 -1328 551 -1316
rect 185 -1330 347 -1328
rect 197 -1348 216 -1330
rect 231 -1332 261 -1330
rect 80 -1358 121 -1350
rect 204 -1354 216 -1348
rect 268 -1346 347 -1330
rect 379 -1330 551 -1328
rect 379 -1346 458 -1330
rect 465 -1332 495 -1330
rect 43 -1368 72 -1358
rect 86 -1368 115 -1358
rect 130 -1368 160 -1354
rect 204 -1368 246 -1354
rect 268 -1358 458 -1346
rect 523 -1350 529 -1330
rect 253 -1368 283 -1358
rect 284 -1368 442 -1358
rect 446 -1368 476 -1358
rect 480 -1368 510 -1354
rect 538 -1368 551 -1330
rect 623 -1316 652 -1300
rect 666 -1316 695 -1300
rect 710 -1310 740 -1294
rect 768 -1316 774 -1268
rect 777 -1274 796 -1268
rect 811 -1274 841 -1266
rect 777 -1282 841 -1274
rect 777 -1298 857 -1282
rect 873 -1289 935 -1258
rect 951 -1289 1013 -1258
rect 1082 -1260 1131 -1235
rect 1146 -1260 1176 -1242
rect 1045 -1274 1075 -1266
rect 1082 -1268 1192 -1260
rect 1045 -1282 1090 -1274
rect 777 -1300 796 -1298
rect 811 -1300 857 -1298
rect 777 -1316 857 -1300
rect 884 -1302 919 -1289
rect 960 -1292 997 -1289
rect 960 -1294 1002 -1292
rect 889 -1305 919 -1302
rect 898 -1309 905 -1305
rect 905 -1310 906 -1309
rect 864 -1316 874 -1310
rect 623 -1324 658 -1316
rect 623 -1350 624 -1324
rect 631 -1350 658 -1324
rect 566 -1368 596 -1354
rect 623 -1358 658 -1350
rect 660 -1324 701 -1316
rect 660 -1350 675 -1324
rect 682 -1350 701 -1324
rect 765 -1328 796 -1316
rect 811 -1328 914 -1316
rect 926 -1326 952 -1300
rect 967 -1305 997 -1294
rect 1029 -1298 1091 -1282
rect 1029 -1300 1075 -1298
rect 1029 -1316 1091 -1300
rect 1103 -1316 1109 -1268
rect 1112 -1276 1192 -1268
rect 1112 -1278 1131 -1276
rect 1146 -1278 1180 -1276
rect 1112 -1293 1192 -1278
rect 1112 -1294 1198 -1293
rect 1112 -1316 1131 -1294
rect 1146 -1310 1176 -1294
rect 1204 -1300 1210 -1226
rect 1213 -1300 1232 -1156
rect 1247 -1300 1253 -1156
rect 1262 -1226 1275 -1156
rect 1327 -1160 1349 -1156
rect 1320 -1172 1337 -1168
rect 1341 -1170 1349 -1168
rect 1339 -1172 1349 -1170
rect 1320 -1182 1349 -1172
rect 1402 -1182 1418 -1168
rect 1456 -1172 1462 -1170
rect 1469 -1172 1577 -1156
rect 1584 -1172 1590 -1170
rect 1598 -1172 1613 -1156
rect 1679 -1162 1698 -1159
rect 1320 -1184 1418 -1182
rect 1445 -1184 1613 -1172
rect 1628 -1182 1644 -1168
rect 1679 -1181 1701 -1162
rect 1711 -1168 1727 -1167
rect 1710 -1170 1727 -1168
rect 1711 -1175 1727 -1170
rect 1701 -1182 1707 -1181
rect 1710 -1182 1739 -1175
rect 1628 -1183 1739 -1182
rect 1628 -1184 1745 -1183
rect 1304 -1192 1355 -1184
rect 1402 -1192 1436 -1184
rect 1304 -1204 1329 -1192
rect 1336 -1204 1355 -1192
rect 1409 -1194 1436 -1192
rect 1445 -1194 1666 -1184
rect 1701 -1187 1707 -1184
rect 1409 -1198 1666 -1194
rect 1304 -1212 1355 -1204
rect 1402 -1212 1666 -1198
rect 1710 -1192 1745 -1184
rect 1256 -1260 1275 -1226
rect 1320 -1220 1349 -1212
rect 1320 -1226 1337 -1220
rect 1320 -1228 1354 -1226
rect 1402 -1228 1418 -1212
rect 1419 -1222 1627 -1212
rect 1628 -1222 1644 -1212
rect 1692 -1216 1707 -1201
rect 1710 -1204 1711 -1192
rect 1718 -1204 1745 -1192
rect 1710 -1212 1745 -1204
rect 1710 -1213 1739 -1212
rect 1430 -1226 1644 -1222
rect 1445 -1228 1644 -1226
rect 1679 -1226 1692 -1216
rect 1710 -1226 1727 -1213
rect 1679 -1228 1727 -1226
rect 1321 -1232 1354 -1228
rect 1317 -1234 1354 -1232
rect 1317 -1235 1384 -1234
rect 1317 -1240 1348 -1235
rect 1354 -1240 1384 -1235
rect 1317 -1244 1384 -1240
rect 1290 -1247 1384 -1244
rect 1290 -1254 1339 -1247
rect 1290 -1260 1320 -1254
rect 1339 -1259 1344 -1254
rect 1256 -1276 1336 -1260
rect 1348 -1268 1384 -1247
rect 1445 -1252 1634 -1228
rect 1679 -1229 1726 -1228
rect 1692 -1234 1726 -1229
rect 1766 -1234 1782 -1232
rect 1460 -1255 1634 -1252
rect 1453 -1258 1634 -1255
rect 1662 -1235 1726 -1234
rect 1256 -1278 1275 -1276
rect 1290 -1278 1324 -1276
rect 1256 -1294 1336 -1278
rect 1256 -1300 1275 -1294
rect 972 -1326 1075 -1316
rect 926 -1328 1075 -1326
rect 1096 -1328 1131 -1316
rect 765 -1330 927 -1328
rect 777 -1348 796 -1330
rect 811 -1332 841 -1330
rect 660 -1358 701 -1350
rect 784 -1354 796 -1348
rect 848 -1348 927 -1330
rect 959 -1330 1131 -1328
rect 959 -1346 1038 -1330
rect 1045 -1332 1075 -1330
rect 934 -1348 1038 -1346
rect 623 -1368 652 -1358
rect 666 -1368 695 -1358
rect 710 -1368 740 -1354
rect 784 -1368 826 -1354
rect 848 -1358 1038 -1348
rect 1103 -1350 1109 -1330
rect 833 -1368 863 -1358
rect 864 -1368 1022 -1358
rect 1026 -1368 1056 -1358
rect 1060 -1368 1090 -1354
rect 1118 -1368 1131 -1330
rect 1203 -1316 1232 -1300
rect 1246 -1316 1275 -1300
rect 1290 -1310 1320 -1294
rect 1348 -1316 1354 -1268
rect 1357 -1274 1376 -1268
rect 1391 -1274 1421 -1266
rect 1357 -1282 1421 -1274
rect 1357 -1298 1437 -1282
rect 1453 -1289 1515 -1258
rect 1531 -1289 1593 -1258
rect 1662 -1260 1711 -1235
rect 1756 -1244 1782 -1234
rect 1726 -1260 1782 -1244
rect 1625 -1274 1655 -1266
rect 1662 -1268 1772 -1260
rect 1625 -1282 1670 -1274
rect 1357 -1300 1376 -1298
rect 1391 -1300 1437 -1298
rect 1357 -1316 1437 -1300
rect 1464 -1302 1499 -1289
rect 1540 -1292 1577 -1289
rect 1540 -1294 1582 -1292
rect 1469 -1305 1499 -1302
rect 1478 -1309 1485 -1305
rect 1485 -1310 1486 -1309
rect 1444 -1316 1454 -1310
rect 1203 -1324 1238 -1316
rect 1203 -1350 1204 -1324
rect 1211 -1350 1238 -1324
rect 1146 -1368 1176 -1354
rect 1203 -1358 1238 -1350
rect 1240 -1324 1281 -1316
rect 1240 -1350 1255 -1324
rect 1262 -1350 1281 -1324
rect 1345 -1328 1376 -1316
rect 1391 -1328 1494 -1316
rect 1506 -1326 1532 -1300
rect 1547 -1305 1577 -1294
rect 1609 -1298 1671 -1282
rect 1609 -1300 1655 -1298
rect 1609 -1316 1671 -1300
rect 1683 -1316 1689 -1268
rect 1692 -1276 1772 -1268
rect 1692 -1278 1711 -1276
rect 1726 -1278 1760 -1276
rect 1692 -1294 1772 -1278
rect 1692 -1316 1711 -1294
rect 1726 -1310 1756 -1294
rect 1784 -1300 1790 -1226
rect 1793 -1300 1812 -1156
rect 1827 -1300 1833 -1156
rect 1842 -1226 1855 -1156
rect 1907 -1160 1929 -1156
rect 1900 -1172 1917 -1168
rect 1921 -1170 1929 -1168
rect 1919 -1172 1929 -1170
rect 1900 -1182 1929 -1172
rect 1982 -1182 1998 -1168
rect 2036 -1172 2042 -1170
rect 2049 -1172 2157 -1156
rect 2164 -1172 2170 -1170
rect 2178 -1172 2193 -1156
rect 2259 -1162 2278 -1159
rect 1900 -1184 1998 -1182
rect 2025 -1184 2193 -1172
rect 2208 -1182 2224 -1168
rect 2259 -1181 2281 -1162
rect 2291 -1168 2307 -1167
rect 2290 -1170 2307 -1168
rect 2291 -1175 2307 -1170
rect 2281 -1182 2287 -1181
rect 2290 -1182 2319 -1175
rect 2208 -1183 2319 -1182
rect 2208 -1184 2325 -1183
rect 1884 -1192 1935 -1184
rect 1982 -1192 2016 -1184
rect 1884 -1204 1909 -1192
rect 1916 -1204 1935 -1192
rect 1989 -1194 2016 -1192
rect 2025 -1194 2246 -1184
rect 2281 -1187 2287 -1184
rect 1989 -1198 2246 -1194
rect 1884 -1212 1935 -1204
rect 1982 -1212 2246 -1198
rect 2290 -1192 2325 -1184
rect 1836 -1260 1855 -1226
rect 1900 -1220 1929 -1212
rect 1900 -1226 1917 -1220
rect 1900 -1228 1934 -1226
rect 1982 -1228 1998 -1212
rect 1999 -1222 2207 -1212
rect 2208 -1222 2224 -1212
rect 2272 -1216 2287 -1201
rect 2290 -1204 2291 -1192
rect 2298 -1204 2325 -1192
rect 2290 -1212 2325 -1204
rect 2290 -1213 2319 -1212
rect 2010 -1226 2224 -1222
rect 2025 -1228 2224 -1226
rect 2259 -1226 2272 -1216
rect 2290 -1226 2307 -1213
rect 2259 -1228 2307 -1226
rect 1901 -1232 1934 -1228
rect 1897 -1234 1934 -1232
rect 1897 -1235 1964 -1234
rect 1897 -1240 1928 -1235
rect 1934 -1240 1964 -1235
rect 1897 -1244 1964 -1240
rect 1870 -1247 1964 -1244
rect 1870 -1254 1919 -1247
rect 1870 -1260 1900 -1254
rect 1919 -1259 1924 -1254
rect 1836 -1276 1916 -1260
rect 1928 -1268 1964 -1247
rect 2025 -1252 2214 -1228
rect 2259 -1229 2306 -1228
rect 2272 -1234 2306 -1229
rect 2040 -1255 2214 -1252
rect 2033 -1258 2214 -1255
rect 2242 -1235 2306 -1234
rect 1836 -1278 1855 -1276
rect 1870 -1278 1904 -1276
rect 1836 -1294 1916 -1278
rect 1836 -1300 1855 -1294
rect 1552 -1326 1655 -1316
rect 1506 -1328 1655 -1326
rect 1676 -1328 1711 -1316
rect 1345 -1330 1507 -1328
rect 1357 -1348 1376 -1330
rect 1391 -1332 1421 -1330
rect 1240 -1358 1281 -1350
rect 1364 -1354 1376 -1348
rect 1428 -1348 1507 -1330
rect 1539 -1330 1711 -1328
rect 1539 -1346 1618 -1330
rect 1625 -1332 1655 -1330
rect 1514 -1348 1618 -1346
rect 1203 -1368 1232 -1358
rect 1246 -1368 1275 -1358
rect 1290 -1368 1320 -1354
rect 1364 -1368 1406 -1354
rect 1428 -1358 1618 -1348
rect 1683 -1350 1689 -1330
rect 1413 -1368 1443 -1358
rect 1444 -1368 1602 -1358
rect 1606 -1368 1636 -1358
rect 1640 -1368 1670 -1354
rect 1698 -1368 1711 -1330
rect 1783 -1316 1812 -1300
rect 1826 -1316 1855 -1300
rect 1870 -1310 1900 -1294
rect 1928 -1316 1934 -1268
rect 1937 -1274 1956 -1268
rect 1971 -1274 2001 -1266
rect 1937 -1282 2001 -1274
rect 1937 -1298 2017 -1282
rect 2033 -1289 2095 -1258
rect 2111 -1289 2173 -1258
rect 2242 -1260 2291 -1235
rect 2306 -1260 2336 -1242
rect 2205 -1274 2235 -1266
rect 2242 -1268 2352 -1260
rect 2205 -1282 2250 -1274
rect 1937 -1300 1956 -1298
rect 1971 -1300 2017 -1298
rect 1937 -1316 2017 -1300
rect 2044 -1302 2079 -1289
rect 2120 -1292 2157 -1289
rect 2120 -1294 2162 -1292
rect 2049 -1305 2079 -1302
rect 2058 -1309 2065 -1305
rect 2065 -1310 2066 -1309
rect 2024 -1316 2034 -1310
rect 1783 -1324 1818 -1316
rect 1783 -1350 1784 -1324
rect 1791 -1350 1818 -1324
rect 1726 -1368 1756 -1354
rect 1783 -1358 1818 -1350
rect 1820 -1324 1861 -1316
rect 1820 -1350 1835 -1324
rect 1842 -1350 1861 -1324
rect 1925 -1328 1956 -1316
rect 1971 -1328 2074 -1316
rect 2086 -1326 2112 -1300
rect 2127 -1305 2157 -1294
rect 2189 -1298 2251 -1282
rect 2189 -1300 2235 -1298
rect 2189 -1316 2251 -1300
rect 2263 -1316 2269 -1268
rect 2272 -1276 2352 -1268
rect 2272 -1278 2291 -1276
rect 2306 -1278 2340 -1276
rect 2272 -1293 2352 -1278
rect 2272 -1294 2358 -1293
rect 2272 -1316 2291 -1294
rect 2306 -1310 2336 -1294
rect 2364 -1300 2370 -1226
rect 2373 -1300 2392 -1156
rect 2407 -1300 2413 -1156
rect 2422 -1226 2435 -1156
rect 2487 -1160 2509 -1156
rect 2480 -1172 2497 -1168
rect 2501 -1170 2509 -1168
rect 2499 -1172 2509 -1170
rect 2480 -1182 2509 -1172
rect 2562 -1182 2578 -1168
rect 2616 -1172 2622 -1170
rect 2629 -1172 2737 -1156
rect 2744 -1172 2750 -1170
rect 2758 -1172 2773 -1156
rect 2839 -1162 2858 -1159
rect 2480 -1184 2578 -1182
rect 2605 -1184 2773 -1172
rect 2788 -1182 2804 -1168
rect 2839 -1181 2861 -1162
rect 2871 -1168 2887 -1167
rect 2870 -1170 2887 -1168
rect 2871 -1175 2887 -1170
rect 2861 -1182 2867 -1181
rect 2870 -1182 2899 -1175
rect 2788 -1183 2899 -1182
rect 2788 -1184 2905 -1183
rect 2464 -1192 2515 -1184
rect 2562 -1192 2596 -1184
rect 2464 -1204 2489 -1192
rect 2496 -1204 2515 -1192
rect 2569 -1194 2596 -1192
rect 2605 -1194 2826 -1184
rect 2861 -1187 2867 -1184
rect 2569 -1198 2826 -1194
rect 2464 -1212 2515 -1204
rect 2562 -1212 2826 -1198
rect 2870 -1192 2905 -1184
rect 2416 -1260 2435 -1226
rect 2480 -1220 2509 -1212
rect 2480 -1226 2497 -1220
rect 2480 -1228 2514 -1226
rect 2562 -1228 2578 -1212
rect 2579 -1222 2787 -1212
rect 2788 -1222 2804 -1212
rect 2852 -1216 2867 -1201
rect 2870 -1204 2871 -1192
rect 2878 -1204 2905 -1192
rect 2870 -1212 2905 -1204
rect 2870 -1213 2899 -1212
rect 2590 -1226 2804 -1222
rect 2605 -1228 2804 -1226
rect 2839 -1226 2852 -1216
rect 2870 -1226 2887 -1213
rect 2839 -1228 2887 -1226
rect 2481 -1232 2514 -1228
rect 2477 -1234 2514 -1232
rect 2477 -1235 2544 -1234
rect 2477 -1240 2508 -1235
rect 2514 -1240 2544 -1235
rect 2477 -1244 2544 -1240
rect 2450 -1247 2544 -1244
rect 2450 -1254 2499 -1247
rect 2450 -1260 2480 -1254
rect 2499 -1259 2504 -1254
rect 2416 -1276 2496 -1260
rect 2508 -1268 2544 -1247
rect 2605 -1252 2794 -1228
rect 2839 -1229 2886 -1228
rect 2852 -1234 2886 -1229
rect 2926 -1234 2942 -1232
rect 2620 -1255 2794 -1252
rect 2613 -1258 2794 -1255
rect 2822 -1235 2886 -1234
rect 2416 -1278 2435 -1276
rect 2450 -1278 2484 -1276
rect 2416 -1294 2496 -1278
rect 2416 -1300 2435 -1294
rect 2132 -1326 2235 -1316
rect 2086 -1328 2235 -1326
rect 2256 -1328 2291 -1316
rect 1925 -1330 2087 -1328
rect 1937 -1348 1956 -1330
rect 1971 -1332 2001 -1330
rect 1820 -1358 1861 -1350
rect 1944 -1354 1956 -1348
rect 2008 -1346 2087 -1330
rect 2119 -1330 2291 -1328
rect 2119 -1346 2198 -1330
rect 2205 -1332 2235 -1330
rect 1783 -1368 1812 -1358
rect 1826 -1368 1855 -1358
rect 1870 -1368 1900 -1354
rect 1944 -1368 1986 -1354
rect 2008 -1358 2198 -1346
rect 2263 -1350 2269 -1330
rect 1993 -1368 2023 -1358
rect 2024 -1368 2182 -1358
rect 2186 -1368 2216 -1358
rect 2220 -1368 2250 -1354
rect 2278 -1368 2291 -1330
rect 2363 -1316 2392 -1300
rect 2406 -1316 2435 -1300
rect 2450 -1310 2480 -1294
rect 2508 -1316 2514 -1268
rect 2517 -1274 2536 -1268
rect 2551 -1274 2581 -1266
rect 2517 -1282 2581 -1274
rect 2517 -1298 2597 -1282
rect 2613 -1289 2675 -1258
rect 2691 -1289 2753 -1258
rect 2822 -1260 2871 -1235
rect 2916 -1244 2942 -1234
rect 2886 -1260 2942 -1244
rect 2785 -1274 2815 -1266
rect 2822 -1268 2932 -1260
rect 2785 -1282 2830 -1274
rect 2517 -1300 2536 -1298
rect 2551 -1300 2597 -1298
rect 2517 -1316 2597 -1300
rect 2624 -1302 2659 -1289
rect 2700 -1292 2737 -1289
rect 2700 -1294 2742 -1292
rect 2629 -1305 2659 -1302
rect 2638 -1309 2645 -1305
rect 2645 -1310 2646 -1309
rect 2604 -1316 2614 -1310
rect 2363 -1324 2398 -1316
rect 2363 -1350 2364 -1324
rect 2371 -1350 2398 -1324
rect 2306 -1368 2336 -1354
rect 2363 -1358 2398 -1350
rect 2400 -1324 2441 -1316
rect 2400 -1350 2415 -1324
rect 2422 -1350 2441 -1324
rect 2505 -1328 2536 -1316
rect 2551 -1328 2654 -1316
rect 2666 -1326 2692 -1300
rect 2707 -1305 2737 -1294
rect 2769 -1298 2831 -1282
rect 2769 -1300 2815 -1298
rect 2769 -1316 2831 -1300
rect 2843 -1316 2849 -1268
rect 2852 -1276 2932 -1268
rect 2852 -1278 2871 -1276
rect 2886 -1278 2920 -1276
rect 2852 -1294 2932 -1278
rect 2852 -1316 2871 -1294
rect 2886 -1310 2916 -1294
rect 2944 -1300 2950 -1226
rect 2953 -1300 2972 -1156
rect 2987 -1300 2993 -1156
rect 3002 -1226 3015 -1156
rect 3067 -1160 3089 -1156
rect 3060 -1172 3077 -1168
rect 3081 -1170 3089 -1168
rect 3079 -1172 3089 -1170
rect 3060 -1182 3089 -1172
rect 3142 -1182 3158 -1168
rect 3196 -1172 3202 -1170
rect 3209 -1172 3317 -1156
rect 3324 -1172 3330 -1170
rect 3338 -1172 3353 -1156
rect 3419 -1162 3438 -1159
rect 3060 -1184 3158 -1182
rect 3185 -1184 3353 -1172
rect 3368 -1182 3384 -1168
rect 3419 -1181 3441 -1162
rect 3451 -1168 3467 -1167
rect 3450 -1170 3467 -1168
rect 3451 -1175 3467 -1170
rect 3441 -1182 3447 -1181
rect 3450 -1182 3479 -1175
rect 3368 -1183 3479 -1182
rect 3368 -1184 3485 -1183
rect 3044 -1192 3095 -1184
rect 3142 -1192 3176 -1184
rect 3044 -1204 3069 -1192
rect 3076 -1204 3095 -1192
rect 3149 -1194 3176 -1192
rect 3185 -1194 3406 -1184
rect 3441 -1187 3447 -1184
rect 3149 -1198 3406 -1194
rect 3044 -1212 3095 -1204
rect 3142 -1212 3406 -1198
rect 3450 -1192 3485 -1184
rect 2996 -1260 3015 -1226
rect 3060 -1220 3089 -1212
rect 3060 -1226 3077 -1220
rect 3060 -1228 3094 -1226
rect 3142 -1228 3158 -1212
rect 3159 -1222 3367 -1212
rect 3368 -1222 3384 -1212
rect 3432 -1216 3447 -1201
rect 3450 -1204 3451 -1192
rect 3458 -1204 3485 -1192
rect 3450 -1212 3485 -1204
rect 3450 -1213 3479 -1212
rect 3170 -1226 3384 -1222
rect 3185 -1228 3384 -1226
rect 3419 -1226 3432 -1216
rect 3450 -1226 3467 -1213
rect 3419 -1228 3467 -1226
rect 3061 -1232 3094 -1228
rect 3057 -1234 3094 -1232
rect 3057 -1235 3124 -1234
rect 3057 -1240 3088 -1235
rect 3094 -1240 3124 -1235
rect 3057 -1244 3124 -1240
rect 3030 -1247 3124 -1244
rect 3030 -1254 3079 -1247
rect 3030 -1260 3060 -1254
rect 3079 -1259 3084 -1254
rect 2996 -1276 3076 -1260
rect 3088 -1268 3124 -1247
rect 3185 -1252 3374 -1228
rect 3419 -1229 3466 -1228
rect 3432 -1234 3466 -1229
rect 3200 -1255 3374 -1252
rect 3193 -1258 3374 -1255
rect 3402 -1235 3466 -1234
rect 2996 -1278 3015 -1276
rect 3030 -1278 3064 -1276
rect 2996 -1294 3076 -1278
rect 2996 -1300 3015 -1294
rect 2712 -1326 2815 -1316
rect 2666 -1328 2815 -1326
rect 2836 -1328 2871 -1316
rect 2505 -1330 2667 -1328
rect 2517 -1348 2536 -1330
rect 2551 -1332 2581 -1330
rect 2400 -1358 2441 -1350
rect 2524 -1354 2536 -1348
rect 2588 -1346 2667 -1330
rect 2699 -1330 2871 -1328
rect 2699 -1346 2778 -1330
rect 2785 -1332 2815 -1330
rect 2363 -1368 2392 -1358
rect 2406 -1368 2435 -1358
rect 2450 -1368 2480 -1354
rect 2524 -1368 2566 -1354
rect 2588 -1358 2778 -1346
rect 2843 -1350 2849 -1330
rect 2573 -1368 2603 -1358
rect 2604 -1368 2762 -1358
rect 2766 -1368 2796 -1358
rect 2800 -1368 2830 -1354
rect 2858 -1368 2871 -1330
rect 2943 -1316 2972 -1300
rect 2986 -1316 3015 -1300
rect 3030 -1310 3060 -1294
rect 3088 -1316 3094 -1268
rect 3097 -1274 3116 -1268
rect 3131 -1274 3161 -1266
rect 3097 -1282 3161 -1274
rect 3097 -1298 3177 -1282
rect 3193 -1289 3255 -1258
rect 3271 -1289 3333 -1258
rect 3402 -1260 3451 -1235
rect 3466 -1260 3496 -1242
rect 3365 -1274 3395 -1266
rect 3402 -1268 3512 -1260
rect 3365 -1282 3410 -1274
rect 3097 -1300 3116 -1298
rect 3131 -1300 3177 -1298
rect 3097 -1316 3177 -1300
rect 3204 -1302 3239 -1289
rect 3280 -1292 3317 -1289
rect 3280 -1294 3322 -1292
rect 3209 -1305 3239 -1302
rect 3218 -1309 3225 -1305
rect 3225 -1310 3226 -1309
rect 3184 -1316 3194 -1310
rect 2943 -1324 2978 -1316
rect 2943 -1350 2944 -1324
rect 2951 -1350 2978 -1324
rect 2886 -1368 2916 -1354
rect 2943 -1358 2978 -1350
rect 2980 -1324 3021 -1316
rect 2980 -1350 2995 -1324
rect 3002 -1350 3021 -1324
rect 3085 -1328 3116 -1316
rect 3131 -1328 3234 -1316
rect 3246 -1326 3272 -1300
rect 3287 -1305 3317 -1294
rect 3349 -1298 3411 -1282
rect 3349 -1300 3395 -1298
rect 3349 -1316 3411 -1300
rect 3423 -1316 3429 -1268
rect 3432 -1276 3512 -1268
rect 3432 -1278 3451 -1276
rect 3466 -1278 3500 -1276
rect 3432 -1293 3512 -1278
rect 3432 -1294 3518 -1293
rect 3432 -1316 3451 -1294
rect 3466 -1310 3496 -1294
rect 3524 -1300 3530 -1226
rect 3533 -1300 3552 -1156
rect 3567 -1300 3573 -1156
rect 3582 -1226 3595 -1156
rect 3647 -1160 3669 -1156
rect 3640 -1172 3657 -1168
rect 3661 -1170 3669 -1168
rect 3659 -1172 3669 -1170
rect 3640 -1182 3669 -1172
rect 3722 -1182 3738 -1168
rect 3776 -1172 3782 -1170
rect 3789 -1172 3897 -1156
rect 3904 -1172 3910 -1170
rect 3918 -1172 3933 -1156
rect 3999 -1162 4018 -1159
rect 3640 -1184 3738 -1182
rect 3765 -1184 3933 -1172
rect 3948 -1182 3964 -1168
rect 3999 -1181 4021 -1162
rect 4031 -1168 4047 -1167
rect 4030 -1170 4047 -1168
rect 4031 -1175 4047 -1170
rect 4021 -1182 4027 -1181
rect 4030 -1182 4059 -1175
rect 3948 -1183 4059 -1182
rect 3948 -1184 4065 -1183
rect 3624 -1192 3675 -1184
rect 3722 -1192 3756 -1184
rect 3624 -1204 3649 -1192
rect 3656 -1204 3675 -1192
rect 3729 -1194 3756 -1192
rect 3765 -1194 3986 -1184
rect 4021 -1187 4027 -1184
rect 3729 -1198 3986 -1194
rect 3624 -1212 3675 -1204
rect 3722 -1212 3986 -1198
rect 4030 -1192 4065 -1184
rect 3576 -1260 3595 -1226
rect 3640 -1220 3669 -1212
rect 3640 -1226 3657 -1220
rect 3640 -1228 3674 -1226
rect 3722 -1228 3738 -1212
rect 3739 -1222 3947 -1212
rect 3948 -1222 3964 -1212
rect 4012 -1216 4027 -1201
rect 4030 -1204 4031 -1192
rect 4038 -1204 4065 -1192
rect 4030 -1212 4065 -1204
rect 4030 -1213 4059 -1212
rect 3750 -1226 3964 -1222
rect 3765 -1228 3964 -1226
rect 3999 -1226 4012 -1216
rect 4030 -1226 4047 -1213
rect 3999 -1228 4047 -1226
rect 3641 -1232 3674 -1228
rect 3637 -1234 3674 -1232
rect 3637 -1235 3704 -1234
rect 3637 -1240 3668 -1235
rect 3674 -1240 3704 -1235
rect 3637 -1244 3704 -1240
rect 3610 -1247 3704 -1244
rect 3610 -1254 3659 -1247
rect 3610 -1260 3640 -1254
rect 3659 -1259 3664 -1254
rect 3576 -1276 3656 -1260
rect 3668 -1268 3704 -1247
rect 3765 -1252 3954 -1228
rect 3999 -1229 4046 -1228
rect 4012 -1234 4046 -1229
rect 4086 -1234 4102 -1232
rect 3780 -1255 3954 -1252
rect 3773 -1258 3954 -1255
rect 3982 -1235 4046 -1234
rect 3576 -1278 3595 -1276
rect 3610 -1278 3644 -1276
rect 3576 -1294 3656 -1278
rect 3576 -1300 3595 -1294
rect 3292 -1326 3395 -1316
rect 3246 -1328 3395 -1326
rect 3416 -1328 3451 -1316
rect 3085 -1330 3247 -1328
rect 3097 -1348 3116 -1330
rect 3131 -1332 3161 -1330
rect 2980 -1358 3021 -1350
rect 3104 -1354 3116 -1348
rect 3168 -1346 3247 -1330
rect 3279 -1330 3451 -1328
rect 3279 -1346 3358 -1330
rect 3365 -1332 3395 -1330
rect 2943 -1368 2972 -1358
rect 2986 -1368 3015 -1358
rect 3030 -1368 3060 -1354
rect 3104 -1368 3146 -1354
rect 3168 -1358 3358 -1346
rect 3423 -1350 3429 -1330
rect 3153 -1368 3183 -1358
rect 3184 -1368 3342 -1358
rect 3346 -1368 3376 -1358
rect 3380 -1368 3410 -1354
rect 3438 -1368 3451 -1330
rect 3523 -1316 3552 -1300
rect 3566 -1316 3595 -1300
rect 3610 -1310 3640 -1294
rect 3668 -1316 3674 -1268
rect 3677 -1274 3696 -1268
rect 3711 -1274 3741 -1266
rect 3677 -1282 3741 -1274
rect 3677 -1298 3757 -1282
rect 3773 -1289 3835 -1258
rect 3851 -1289 3913 -1258
rect 3982 -1260 4031 -1235
rect 4076 -1244 4102 -1234
rect 4046 -1260 4102 -1244
rect 3945 -1274 3975 -1266
rect 3982 -1268 4092 -1260
rect 3945 -1282 3990 -1274
rect 3677 -1300 3696 -1298
rect 3711 -1300 3757 -1298
rect 3677 -1316 3757 -1300
rect 3784 -1302 3819 -1289
rect 3860 -1292 3897 -1289
rect 3860 -1294 3902 -1292
rect 3789 -1305 3819 -1302
rect 3798 -1309 3805 -1305
rect 3805 -1310 3806 -1309
rect 3764 -1316 3774 -1310
rect 3523 -1324 3558 -1316
rect 3523 -1350 3524 -1324
rect 3531 -1350 3558 -1324
rect 3466 -1368 3496 -1354
rect 3523 -1358 3558 -1350
rect 3560 -1324 3601 -1316
rect 3560 -1350 3575 -1324
rect 3582 -1350 3601 -1324
rect 3665 -1328 3696 -1316
rect 3711 -1328 3814 -1316
rect 3826 -1326 3852 -1300
rect 3867 -1305 3897 -1294
rect 3929 -1298 3991 -1282
rect 3929 -1300 3975 -1298
rect 3929 -1316 3991 -1300
rect 4003 -1316 4009 -1268
rect 4012 -1276 4092 -1268
rect 4012 -1278 4031 -1276
rect 4046 -1278 4080 -1276
rect 4012 -1294 4092 -1278
rect 4012 -1316 4031 -1294
rect 4046 -1310 4076 -1294
rect 4104 -1300 4110 -1226
rect 4113 -1300 4132 -1156
rect 4147 -1300 4153 -1156
rect 4162 -1226 4175 -1156
rect 4227 -1160 4249 -1156
rect 4220 -1172 4237 -1168
rect 4241 -1170 4249 -1168
rect 4239 -1172 4249 -1170
rect 4220 -1182 4249 -1172
rect 4302 -1182 4318 -1168
rect 4356 -1172 4362 -1170
rect 4369 -1172 4477 -1156
rect 4484 -1172 4490 -1170
rect 4498 -1172 4513 -1156
rect 4579 -1162 4598 -1159
rect 4220 -1184 4318 -1182
rect 4345 -1184 4513 -1172
rect 4528 -1182 4544 -1168
rect 4579 -1181 4601 -1162
rect 4611 -1168 4627 -1167
rect 4610 -1170 4627 -1168
rect 4611 -1175 4627 -1170
rect 4601 -1182 4607 -1181
rect 4610 -1182 4639 -1175
rect 4528 -1183 4639 -1182
rect 4528 -1184 4645 -1183
rect 4204 -1192 4255 -1184
rect 4302 -1192 4336 -1184
rect 4204 -1204 4229 -1192
rect 4236 -1204 4255 -1192
rect 4309 -1194 4336 -1192
rect 4345 -1194 4566 -1184
rect 4601 -1187 4607 -1184
rect 4309 -1198 4566 -1194
rect 4204 -1212 4255 -1204
rect 4302 -1212 4566 -1198
rect 4610 -1192 4645 -1184
rect 4156 -1260 4175 -1226
rect 4220 -1220 4249 -1212
rect 4220 -1226 4237 -1220
rect 4220 -1228 4254 -1226
rect 4302 -1228 4318 -1212
rect 4319 -1222 4527 -1212
rect 4528 -1222 4544 -1212
rect 4592 -1216 4607 -1201
rect 4610 -1204 4611 -1192
rect 4618 -1204 4645 -1192
rect 4610 -1212 4645 -1204
rect 4610 -1213 4639 -1212
rect 4330 -1226 4544 -1222
rect 4345 -1228 4544 -1226
rect 4579 -1226 4592 -1216
rect 4610 -1226 4627 -1213
rect 4579 -1228 4627 -1226
rect 4221 -1232 4254 -1228
rect 4217 -1234 4254 -1232
rect 4217 -1235 4284 -1234
rect 4217 -1240 4248 -1235
rect 4254 -1240 4284 -1235
rect 4217 -1244 4284 -1240
rect 4190 -1247 4284 -1244
rect 4190 -1254 4239 -1247
rect 4190 -1260 4220 -1254
rect 4239 -1259 4244 -1254
rect 4156 -1276 4236 -1260
rect 4248 -1268 4284 -1247
rect 4345 -1252 4534 -1228
rect 4579 -1229 4626 -1228
rect 4592 -1234 4626 -1229
rect 4360 -1255 4534 -1252
rect 4353 -1258 4534 -1255
rect 4562 -1235 4626 -1234
rect 4156 -1278 4175 -1276
rect 4190 -1278 4224 -1276
rect 4156 -1294 4236 -1278
rect 4156 -1300 4175 -1294
rect 3872 -1326 3975 -1316
rect 3826 -1328 3975 -1326
rect 3996 -1328 4031 -1316
rect 3665 -1330 3827 -1328
rect 3677 -1348 3696 -1330
rect 3711 -1332 3741 -1330
rect 3560 -1358 3601 -1350
rect 3684 -1354 3696 -1348
rect 3748 -1346 3827 -1330
rect 3859 -1330 4031 -1328
rect 3859 -1346 3938 -1330
rect 3945 -1332 3975 -1330
rect 3523 -1368 3552 -1358
rect 3566 -1368 3595 -1358
rect 3610 -1368 3640 -1354
rect 3684 -1368 3726 -1354
rect 3748 -1358 3938 -1346
rect 4003 -1350 4009 -1330
rect 3733 -1368 3763 -1358
rect 3764 -1368 3922 -1358
rect 3926 -1368 3956 -1358
rect 3960 -1368 3990 -1354
rect 4018 -1368 4031 -1330
rect 4103 -1316 4132 -1300
rect 4146 -1316 4175 -1300
rect 4190 -1310 4220 -1294
rect 4248 -1316 4254 -1268
rect 4257 -1274 4276 -1268
rect 4291 -1274 4321 -1266
rect 4257 -1282 4321 -1274
rect 4257 -1298 4337 -1282
rect 4353 -1289 4415 -1258
rect 4431 -1289 4493 -1258
rect 4562 -1260 4611 -1235
rect 4626 -1260 4656 -1242
rect 4525 -1274 4555 -1266
rect 4562 -1268 4672 -1260
rect 4525 -1282 4570 -1274
rect 4257 -1300 4276 -1298
rect 4291 -1300 4337 -1298
rect 4257 -1316 4337 -1300
rect 4364 -1302 4399 -1289
rect 4440 -1292 4477 -1289
rect 4440 -1294 4482 -1292
rect 4369 -1305 4399 -1302
rect 4378 -1309 4385 -1305
rect 4385 -1310 4386 -1309
rect 4344 -1316 4354 -1310
rect 4103 -1324 4138 -1316
rect 4103 -1350 4104 -1324
rect 4111 -1350 4138 -1324
rect 4046 -1368 4076 -1354
rect 4103 -1358 4138 -1350
rect 4140 -1324 4181 -1316
rect 4140 -1350 4155 -1324
rect 4162 -1350 4181 -1324
rect 4245 -1328 4276 -1316
rect 4291 -1328 4394 -1316
rect 4406 -1326 4432 -1300
rect 4447 -1305 4477 -1294
rect 4509 -1298 4571 -1282
rect 4509 -1300 4555 -1298
rect 4509 -1316 4571 -1300
rect 4583 -1316 4589 -1268
rect 4592 -1276 4672 -1268
rect 4592 -1278 4611 -1276
rect 4626 -1278 4660 -1276
rect 4592 -1293 4672 -1278
rect 4592 -1294 4678 -1293
rect 4592 -1316 4611 -1294
rect 4626 -1310 4656 -1294
rect 4684 -1300 4690 -1226
rect 4693 -1300 4712 -1156
rect 4727 -1300 4733 -1156
rect 4742 -1226 4755 -1156
rect 4807 -1160 4829 -1156
rect 4800 -1172 4817 -1168
rect 4821 -1170 4829 -1168
rect 4819 -1172 4829 -1170
rect 4800 -1182 4829 -1172
rect 4882 -1182 4898 -1168
rect 4936 -1172 4942 -1170
rect 4949 -1172 5057 -1156
rect 5064 -1172 5070 -1170
rect 5078 -1172 5093 -1156
rect 5159 -1162 5178 -1159
rect 4800 -1184 4898 -1182
rect 4925 -1184 5093 -1172
rect 5108 -1182 5124 -1168
rect 5159 -1181 5181 -1162
rect 5191 -1168 5207 -1167
rect 5190 -1170 5207 -1168
rect 5191 -1175 5207 -1170
rect 5181 -1182 5187 -1181
rect 5190 -1182 5219 -1175
rect 5108 -1183 5219 -1182
rect 5108 -1184 5225 -1183
rect 4784 -1192 4835 -1184
rect 4882 -1192 4916 -1184
rect 4784 -1204 4809 -1192
rect 4816 -1204 4835 -1192
rect 4889 -1194 4916 -1192
rect 4925 -1194 5146 -1184
rect 5181 -1187 5187 -1184
rect 4889 -1198 5146 -1194
rect 4784 -1212 4835 -1204
rect 4882 -1212 5146 -1198
rect 5190 -1192 5225 -1184
rect 4736 -1260 4755 -1226
rect 4800 -1220 4829 -1212
rect 4800 -1226 4817 -1220
rect 4800 -1228 4834 -1226
rect 4882 -1228 4898 -1212
rect 4899 -1222 5107 -1212
rect 5108 -1222 5124 -1212
rect 5172 -1216 5187 -1201
rect 5190 -1204 5191 -1192
rect 5198 -1204 5225 -1192
rect 5190 -1212 5225 -1204
rect 5190 -1213 5219 -1212
rect 4910 -1226 5124 -1222
rect 4925 -1228 5124 -1226
rect 5159 -1226 5172 -1216
rect 5190 -1226 5207 -1213
rect 5159 -1228 5207 -1226
rect 4801 -1232 4834 -1228
rect 4797 -1234 4834 -1232
rect 4797 -1235 4864 -1234
rect 4797 -1240 4828 -1235
rect 4834 -1240 4864 -1235
rect 4797 -1244 4864 -1240
rect 4770 -1247 4864 -1244
rect 4770 -1254 4819 -1247
rect 4770 -1260 4800 -1254
rect 4819 -1259 4824 -1254
rect 4736 -1276 4816 -1260
rect 4828 -1268 4864 -1247
rect 4925 -1252 5114 -1228
rect 5159 -1229 5206 -1228
rect 5172 -1234 5206 -1229
rect 5246 -1234 5262 -1232
rect 4940 -1255 5114 -1252
rect 4933 -1258 5114 -1255
rect 5142 -1235 5206 -1234
rect 4736 -1278 4755 -1276
rect 4770 -1278 4804 -1276
rect 4736 -1294 4816 -1278
rect 4736 -1300 4755 -1294
rect 4452 -1326 4555 -1316
rect 4406 -1328 4555 -1326
rect 4576 -1328 4611 -1316
rect 4245 -1330 4407 -1328
rect 4257 -1348 4276 -1330
rect 4291 -1332 4321 -1330
rect 4140 -1358 4181 -1350
rect 4264 -1354 4276 -1348
rect 4328 -1346 4407 -1330
rect 4439 -1330 4611 -1328
rect 4439 -1346 4518 -1330
rect 4525 -1332 4555 -1330
rect 4103 -1368 4132 -1358
rect 4146 -1368 4175 -1358
rect 4190 -1368 4220 -1354
rect 4264 -1368 4306 -1354
rect 4328 -1358 4518 -1346
rect 4583 -1350 4589 -1330
rect 4313 -1368 4343 -1358
rect 4344 -1368 4502 -1358
rect 4506 -1368 4536 -1358
rect 4540 -1368 4570 -1354
rect 4598 -1368 4611 -1330
rect 4683 -1316 4712 -1300
rect 4726 -1316 4755 -1300
rect 4770 -1310 4800 -1294
rect 4828 -1316 4834 -1268
rect 4837 -1274 4856 -1268
rect 4871 -1274 4901 -1266
rect 4837 -1282 4901 -1274
rect 4837 -1298 4917 -1282
rect 4933 -1289 4995 -1258
rect 5011 -1289 5073 -1258
rect 5142 -1260 5191 -1235
rect 5236 -1244 5262 -1234
rect 5206 -1260 5262 -1244
rect 5105 -1274 5135 -1266
rect 5142 -1268 5252 -1260
rect 5105 -1282 5150 -1274
rect 4837 -1300 4856 -1298
rect 4871 -1300 4917 -1298
rect 4837 -1316 4917 -1300
rect 4944 -1302 4979 -1289
rect 5020 -1292 5057 -1289
rect 5020 -1294 5062 -1292
rect 4949 -1305 4979 -1302
rect 4958 -1309 4965 -1305
rect 4965 -1310 4966 -1309
rect 4924 -1316 4934 -1310
rect 4683 -1324 4718 -1316
rect 4683 -1350 4684 -1324
rect 4691 -1350 4718 -1324
rect 4626 -1368 4656 -1354
rect 4683 -1358 4718 -1350
rect 4720 -1324 4761 -1316
rect 4720 -1350 4735 -1324
rect 4742 -1350 4761 -1324
rect 4825 -1328 4856 -1316
rect 4871 -1328 4974 -1316
rect 4986 -1326 5012 -1300
rect 5027 -1305 5057 -1294
rect 5089 -1298 5151 -1282
rect 5089 -1300 5135 -1298
rect 5089 -1316 5151 -1300
rect 5163 -1316 5169 -1268
rect 5172 -1276 5252 -1268
rect 5172 -1278 5191 -1276
rect 5206 -1278 5240 -1276
rect 5172 -1294 5252 -1278
rect 5172 -1316 5191 -1294
rect 5206 -1310 5236 -1294
rect 5264 -1300 5270 -1226
rect 5273 -1300 5292 -1156
rect 5307 -1300 5313 -1156
rect 5322 -1226 5335 -1156
rect 5387 -1160 5409 -1156
rect 5380 -1172 5397 -1168
rect 5401 -1170 5409 -1168
rect 5399 -1172 5409 -1170
rect 5380 -1182 5409 -1172
rect 5462 -1182 5478 -1168
rect 5516 -1172 5522 -1170
rect 5529 -1172 5637 -1156
rect 5644 -1172 5650 -1170
rect 5658 -1172 5673 -1156
rect 5739 -1162 5758 -1159
rect 5380 -1184 5478 -1182
rect 5505 -1184 5673 -1172
rect 5688 -1182 5704 -1168
rect 5739 -1181 5761 -1162
rect 5771 -1168 5787 -1167
rect 5770 -1170 5787 -1168
rect 5771 -1175 5787 -1170
rect 5761 -1182 5767 -1181
rect 5770 -1182 5799 -1175
rect 5688 -1183 5799 -1182
rect 5688 -1184 5805 -1183
rect 5364 -1192 5415 -1184
rect 5462 -1192 5496 -1184
rect 5364 -1204 5389 -1192
rect 5396 -1204 5415 -1192
rect 5469 -1194 5496 -1192
rect 5505 -1194 5726 -1184
rect 5761 -1187 5767 -1184
rect 5469 -1198 5726 -1194
rect 5364 -1212 5415 -1204
rect 5462 -1212 5726 -1198
rect 5770 -1192 5805 -1184
rect 5316 -1260 5335 -1226
rect 5380 -1220 5409 -1212
rect 5380 -1226 5397 -1220
rect 5380 -1228 5414 -1226
rect 5462 -1228 5478 -1212
rect 5479 -1222 5687 -1212
rect 5688 -1222 5704 -1212
rect 5752 -1216 5767 -1201
rect 5770 -1204 5771 -1192
rect 5778 -1204 5805 -1192
rect 5770 -1212 5805 -1204
rect 5770 -1213 5799 -1212
rect 5490 -1226 5704 -1222
rect 5505 -1228 5704 -1226
rect 5739 -1226 5752 -1216
rect 5770 -1226 5787 -1213
rect 5739 -1228 5787 -1226
rect 5381 -1232 5414 -1228
rect 5377 -1234 5414 -1232
rect 5377 -1235 5444 -1234
rect 5377 -1240 5408 -1235
rect 5414 -1240 5444 -1235
rect 5377 -1244 5444 -1240
rect 5350 -1247 5444 -1244
rect 5350 -1254 5399 -1247
rect 5350 -1260 5380 -1254
rect 5399 -1259 5404 -1254
rect 5316 -1276 5396 -1260
rect 5408 -1268 5444 -1247
rect 5505 -1252 5694 -1228
rect 5739 -1229 5786 -1228
rect 5752 -1234 5786 -1229
rect 5520 -1255 5694 -1252
rect 5513 -1258 5694 -1255
rect 5722 -1235 5786 -1234
rect 5316 -1278 5335 -1276
rect 5350 -1278 5384 -1276
rect 5316 -1294 5396 -1278
rect 5316 -1300 5335 -1294
rect 5032 -1326 5135 -1316
rect 4986 -1328 5135 -1326
rect 5156 -1328 5191 -1316
rect 4825 -1330 4987 -1328
rect 4837 -1348 4856 -1330
rect 4871 -1332 4901 -1330
rect 4720 -1358 4761 -1350
rect 4844 -1354 4856 -1348
rect 4908 -1346 4987 -1330
rect 5019 -1330 5191 -1328
rect 5019 -1346 5098 -1330
rect 5105 -1332 5135 -1330
rect 4683 -1368 4712 -1358
rect 4726 -1368 4755 -1358
rect 4770 -1368 4800 -1354
rect 4844 -1368 4886 -1354
rect 4908 -1358 5098 -1346
rect 5163 -1350 5169 -1330
rect 4893 -1368 4923 -1358
rect 4924 -1368 5082 -1358
rect 5086 -1368 5116 -1358
rect 5120 -1368 5150 -1354
rect 5178 -1368 5191 -1330
rect 5263 -1316 5292 -1300
rect 5306 -1316 5335 -1300
rect 5350 -1310 5380 -1294
rect 5408 -1316 5414 -1268
rect 5417 -1274 5436 -1268
rect 5451 -1274 5481 -1266
rect 5417 -1282 5481 -1274
rect 5417 -1298 5497 -1282
rect 5513 -1289 5575 -1258
rect 5591 -1289 5653 -1258
rect 5722 -1260 5771 -1235
rect 5786 -1260 5816 -1242
rect 5685 -1274 5715 -1266
rect 5722 -1268 5832 -1260
rect 5685 -1282 5730 -1274
rect 5417 -1300 5436 -1298
rect 5451 -1300 5497 -1298
rect 5417 -1316 5497 -1300
rect 5524 -1302 5559 -1289
rect 5600 -1292 5637 -1289
rect 5600 -1294 5642 -1292
rect 5529 -1305 5559 -1302
rect 5538 -1309 5545 -1305
rect 5545 -1310 5546 -1309
rect 5504 -1316 5514 -1310
rect 5263 -1324 5298 -1316
rect 5263 -1350 5264 -1324
rect 5271 -1350 5298 -1324
rect 5206 -1368 5236 -1354
rect 5263 -1358 5298 -1350
rect 5300 -1324 5341 -1316
rect 5300 -1350 5315 -1324
rect 5322 -1350 5341 -1324
rect 5405 -1328 5436 -1316
rect 5451 -1328 5554 -1316
rect 5566 -1326 5592 -1300
rect 5607 -1305 5637 -1294
rect 5669 -1298 5731 -1282
rect 5669 -1300 5715 -1298
rect 5669 -1316 5731 -1300
rect 5743 -1316 5749 -1268
rect 5752 -1276 5832 -1268
rect 5752 -1278 5771 -1276
rect 5786 -1278 5820 -1276
rect 5752 -1293 5832 -1278
rect 5752 -1294 5838 -1293
rect 5752 -1316 5771 -1294
rect 5786 -1310 5816 -1294
rect 5844 -1300 5850 -1226
rect 5853 -1300 5872 -1156
rect 5887 -1300 5893 -1156
rect 5902 -1226 5915 -1156
rect 5967 -1160 5989 -1156
rect 5960 -1172 5977 -1168
rect 5981 -1170 5989 -1168
rect 5979 -1172 5989 -1170
rect 5960 -1182 5989 -1172
rect 6042 -1182 6058 -1168
rect 6096 -1172 6102 -1170
rect 6109 -1172 6217 -1156
rect 6224 -1172 6230 -1170
rect 6238 -1172 6253 -1156
rect 6319 -1162 6338 -1159
rect 5960 -1184 6058 -1182
rect 6085 -1184 6253 -1172
rect 6268 -1182 6284 -1168
rect 6319 -1181 6341 -1162
rect 6351 -1168 6367 -1167
rect 6350 -1170 6367 -1168
rect 6351 -1175 6367 -1170
rect 6341 -1182 6347 -1181
rect 6350 -1182 6379 -1175
rect 6268 -1183 6379 -1182
rect 6268 -1184 6385 -1183
rect 5944 -1192 5995 -1184
rect 6042 -1192 6076 -1184
rect 5944 -1204 5969 -1192
rect 5976 -1204 5995 -1192
rect 6049 -1194 6076 -1192
rect 6085 -1194 6306 -1184
rect 6341 -1187 6347 -1184
rect 6049 -1198 6306 -1194
rect 5944 -1212 5995 -1204
rect 6042 -1212 6306 -1198
rect 6350 -1192 6385 -1184
rect 5896 -1260 5915 -1226
rect 5960 -1220 5989 -1212
rect 5960 -1226 5977 -1220
rect 5960 -1228 5994 -1226
rect 6042 -1228 6058 -1212
rect 6059 -1222 6267 -1212
rect 6268 -1222 6284 -1212
rect 6332 -1216 6347 -1201
rect 6350 -1204 6351 -1192
rect 6358 -1204 6385 -1192
rect 6350 -1212 6385 -1204
rect 6350 -1213 6379 -1212
rect 6070 -1226 6284 -1222
rect 6085 -1228 6284 -1226
rect 6319 -1226 6332 -1216
rect 6350 -1226 6367 -1213
rect 6319 -1228 6367 -1226
rect 5961 -1232 5994 -1228
rect 5957 -1234 5994 -1232
rect 5957 -1235 6024 -1234
rect 5957 -1240 5988 -1235
rect 5994 -1240 6024 -1235
rect 5957 -1244 6024 -1240
rect 5930 -1247 6024 -1244
rect 5930 -1254 5979 -1247
rect 5930 -1260 5960 -1254
rect 5979 -1259 5984 -1254
rect 5896 -1276 5976 -1260
rect 5988 -1268 6024 -1247
rect 6085 -1252 6274 -1228
rect 6319 -1229 6366 -1228
rect 6332 -1234 6366 -1229
rect 6100 -1255 6274 -1252
rect 6093 -1258 6274 -1255
rect 6302 -1235 6366 -1234
rect 5896 -1278 5915 -1276
rect 5930 -1278 5964 -1276
rect 5896 -1294 5976 -1278
rect 5896 -1300 5915 -1294
rect 5612 -1326 5715 -1316
rect 5566 -1328 5715 -1326
rect 5736 -1328 5771 -1316
rect 5405 -1330 5567 -1328
rect 5417 -1348 5436 -1330
rect 5451 -1332 5481 -1330
rect 5300 -1358 5341 -1350
rect 5424 -1354 5436 -1348
rect 5488 -1346 5567 -1330
rect 5599 -1330 5771 -1328
rect 5599 -1346 5678 -1330
rect 5685 -1332 5715 -1330
rect 5263 -1368 5292 -1358
rect 5306 -1368 5335 -1358
rect 5350 -1368 5380 -1354
rect 5424 -1368 5466 -1354
rect 5488 -1358 5678 -1346
rect 5743 -1350 5749 -1330
rect 5473 -1368 5503 -1358
rect 5504 -1368 5662 -1358
rect 5666 -1368 5696 -1358
rect 5700 -1368 5730 -1354
rect 5758 -1368 5771 -1330
rect 5843 -1316 5872 -1300
rect 5886 -1316 5915 -1300
rect 5930 -1310 5960 -1294
rect 5988 -1316 5994 -1268
rect 5997 -1274 6016 -1268
rect 6031 -1274 6061 -1266
rect 5997 -1282 6061 -1274
rect 5997 -1298 6077 -1282
rect 6093 -1289 6155 -1258
rect 6171 -1289 6233 -1258
rect 6302 -1260 6351 -1235
rect 6366 -1260 6396 -1244
rect 6265 -1274 6295 -1266
rect 6302 -1268 6412 -1260
rect 6265 -1282 6310 -1274
rect 5997 -1300 6016 -1298
rect 6031 -1300 6077 -1298
rect 5997 -1316 6077 -1300
rect 6104 -1302 6139 -1289
rect 6180 -1292 6217 -1289
rect 6180 -1294 6222 -1292
rect 6109 -1305 6139 -1302
rect 6118 -1309 6125 -1305
rect 6125 -1310 6126 -1309
rect 6084 -1316 6094 -1310
rect 5843 -1324 5878 -1316
rect 5843 -1350 5844 -1324
rect 5851 -1350 5878 -1324
rect 5786 -1368 5816 -1354
rect 5843 -1358 5878 -1350
rect 5880 -1324 5921 -1316
rect 5880 -1350 5895 -1324
rect 5902 -1350 5921 -1324
rect 5985 -1328 6016 -1316
rect 6031 -1328 6134 -1316
rect 6146 -1326 6172 -1300
rect 6187 -1305 6217 -1294
rect 6249 -1298 6311 -1282
rect 6249 -1300 6295 -1298
rect 6249 -1316 6311 -1300
rect 6323 -1316 6329 -1268
rect 6332 -1276 6412 -1268
rect 6332 -1278 6351 -1276
rect 6366 -1278 6400 -1276
rect 6332 -1294 6412 -1278
rect 6332 -1316 6351 -1294
rect 6366 -1310 6396 -1294
rect 6424 -1300 6430 -1226
rect 6439 -1300 6452 -1156
rect 6192 -1326 6295 -1316
rect 6146 -1328 6295 -1326
rect 6316 -1328 6351 -1316
rect 5985 -1330 6147 -1328
rect 5997 -1348 6016 -1330
rect 6031 -1332 6061 -1330
rect 5880 -1358 5921 -1350
rect 6004 -1354 6016 -1348
rect 6068 -1346 6147 -1330
rect 6179 -1330 6351 -1328
rect 6179 -1346 6258 -1330
rect 6265 -1332 6295 -1330
rect 5843 -1368 5872 -1358
rect 5886 -1368 5915 -1358
rect 5930 -1368 5960 -1354
rect 6004 -1368 6046 -1354
rect 6068 -1358 6258 -1346
rect 6323 -1350 6329 -1330
rect 6053 -1368 6083 -1358
rect 6084 -1368 6242 -1358
rect 6246 -1368 6276 -1358
rect 6280 -1368 6310 -1354
rect 6338 -1368 6351 -1330
rect 6423 -1316 6452 -1300
rect 6423 -1324 6458 -1316
rect 6423 -1350 6424 -1324
rect 6431 -1350 6458 -1324
rect 6366 -1368 6396 -1354
rect 6423 -1358 6458 -1350
rect 6423 -1368 6452 -1358
rect -541 -1382 6452 -1368
rect -478 -1412 -465 -1382
rect -450 -1396 -420 -1382
rect -376 -1396 -334 -1382
rect -327 -1396 -107 -1382
rect -100 -1396 -70 -1382
rect -410 -1410 -395 -1398
rect -376 -1410 -363 -1396
rect -295 -1400 -142 -1396
rect -413 -1412 -391 -1410
rect -313 -1412 -121 -1400
rect -42 -1412 -29 -1382
rect -14 -1396 16 -1382
rect 53 -1412 72 -1382
rect 87 -1412 93 -1382
rect 102 -1412 115 -1382
rect 130 -1396 160 -1382
rect 204 -1396 246 -1382
rect 253 -1396 473 -1382
rect 480 -1396 510 -1382
rect 170 -1410 185 -1398
rect 204 -1410 217 -1396
rect 285 -1400 438 -1396
rect 167 -1412 189 -1410
rect 267 -1412 459 -1400
rect 538 -1412 551 -1382
rect 566 -1396 596 -1382
rect 633 -1412 652 -1382
rect 667 -1412 673 -1382
rect 682 -1412 695 -1382
rect 710 -1396 740 -1382
rect 784 -1396 826 -1382
rect 833 -1396 1053 -1382
rect 1060 -1396 1090 -1382
rect 750 -1410 765 -1398
rect 784 -1410 797 -1396
rect 865 -1400 1018 -1396
rect 747 -1412 769 -1410
rect 847 -1412 1039 -1400
rect 1118 -1412 1131 -1382
rect 1146 -1396 1176 -1382
rect 1213 -1412 1232 -1382
rect 1247 -1412 1253 -1382
rect 1262 -1412 1275 -1382
rect 1290 -1396 1320 -1382
rect 1364 -1396 1406 -1382
rect 1413 -1396 1633 -1382
rect 1640 -1396 1670 -1382
rect 1330 -1410 1345 -1398
rect 1364 -1410 1377 -1396
rect 1445 -1400 1598 -1396
rect 1327 -1412 1349 -1410
rect 1427 -1412 1619 -1400
rect 1698 -1412 1711 -1382
rect 1726 -1396 1756 -1382
rect 1793 -1412 1812 -1382
rect 1827 -1412 1833 -1382
rect 1842 -1412 1855 -1382
rect 1870 -1396 1900 -1382
rect 1944 -1396 1986 -1382
rect 1993 -1396 2213 -1382
rect 2220 -1396 2250 -1382
rect 1910 -1410 1925 -1398
rect 1944 -1410 1957 -1396
rect 2025 -1400 2178 -1396
rect 1907 -1412 1929 -1410
rect 2007 -1412 2199 -1400
rect 2278 -1412 2291 -1382
rect 2306 -1396 2336 -1382
rect 2373 -1412 2392 -1382
rect 2407 -1412 2413 -1382
rect 2422 -1412 2435 -1382
rect 2450 -1396 2480 -1382
rect 2524 -1396 2566 -1382
rect 2573 -1396 2793 -1382
rect 2800 -1396 2830 -1382
rect 2490 -1410 2505 -1398
rect 2524 -1410 2537 -1396
rect 2605 -1400 2758 -1396
rect 2487 -1412 2509 -1410
rect 2587 -1412 2779 -1400
rect 2858 -1412 2871 -1382
rect 2886 -1396 2916 -1382
rect 2953 -1412 2972 -1382
rect 2987 -1412 2993 -1382
rect 3002 -1412 3015 -1382
rect 3030 -1396 3060 -1382
rect 3104 -1396 3146 -1382
rect 3153 -1396 3373 -1382
rect 3380 -1396 3410 -1382
rect 3070 -1410 3085 -1398
rect 3104 -1410 3117 -1396
rect 3185 -1400 3338 -1396
rect 3067 -1412 3089 -1410
rect 3167 -1412 3359 -1400
rect 3438 -1412 3451 -1382
rect 3466 -1396 3496 -1382
rect 3533 -1412 3552 -1382
rect 3567 -1412 3573 -1382
rect 3582 -1412 3595 -1382
rect 3610 -1396 3640 -1382
rect 3684 -1396 3726 -1382
rect 3733 -1396 3953 -1382
rect 3960 -1396 3990 -1382
rect 3650 -1410 3665 -1398
rect 3684 -1410 3697 -1396
rect 3765 -1400 3918 -1396
rect 3647 -1412 3669 -1410
rect 3747 -1412 3939 -1400
rect 4018 -1412 4031 -1382
rect 4046 -1396 4076 -1382
rect 4113 -1412 4132 -1382
rect 4147 -1412 4153 -1382
rect 4162 -1412 4175 -1382
rect 4190 -1396 4220 -1382
rect 4264 -1396 4306 -1382
rect 4313 -1396 4533 -1382
rect 4540 -1396 4570 -1382
rect 4230 -1410 4245 -1398
rect 4264 -1410 4277 -1396
rect 4345 -1400 4498 -1396
rect 4227 -1412 4249 -1410
rect 4327 -1412 4519 -1400
rect 4598 -1412 4611 -1382
rect 4626 -1396 4656 -1382
rect 4693 -1412 4712 -1382
rect 4727 -1412 4733 -1382
rect 4742 -1412 4755 -1382
rect 4770 -1396 4800 -1382
rect 4844 -1396 4886 -1382
rect 4893 -1396 5113 -1382
rect 5120 -1396 5150 -1382
rect 4810 -1410 4825 -1398
rect 4844 -1410 4857 -1396
rect 4925 -1400 5078 -1396
rect 4807 -1412 4829 -1410
rect 4907 -1412 5099 -1400
rect 5178 -1412 5191 -1382
rect 5206 -1396 5236 -1382
rect 5273 -1412 5292 -1382
rect 5307 -1412 5313 -1382
rect 5322 -1412 5335 -1382
rect 5350 -1396 5380 -1382
rect 5424 -1396 5466 -1382
rect 5473 -1396 5693 -1382
rect 5700 -1396 5730 -1382
rect 5390 -1410 5405 -1398
rect 5424 -1410 5437 -1396
rect 5505 -1400 5658 -1396
rect 5387 -1412 5409 -1410
rect 5487 -1412 5679 -1400
rect 5758 -1412 5771 -1382
rect 5786 -1396 5816 -1382
rect 5853 -1412 5872 -1382
rect 5887 -1412 5893 -1382
rect 5902 -1412 5915 -1382
rect 5930 -1396 5960 -1382
rect 6004 -1396 6046 -1382
rect 6053 -1396 6273 -1382
rect 6280 -1396 6310 -1382
rect 5970 -1410 5985 -1398
rect 6004 -1410 6017 -1396
rect 6085 -1400 6238 -1396
rect 5967 -1412 5989 -1410
rect 6067 -1412 6259 -1400
rect 6338 -1412 6351 -1382
rect 6366 -1396 6396 -1382
rect 6439 -1412 6452 -1382
rect -541 -1426 6452 -1412
rect -478 -1496 -465 -1426
rect -413 -1430 -391 -1426
rect -420 -1442 -403 -1438
rect -399 -1440 -391 -1438
rect -401 -1442 -391 -1440
rect -420 -1452 -391 -1442
rect -338 -1452 -322 -1438
rect -284 -1442 -278 -1440
rect -271 -1442 -163 -1426
rect -156 -1442 -150 -1440
rect -142 -1442 -127 -1426
rect -61 -1432 -42 -1429
rect -420 -1454 -322 -1452
rect -295 -1454 -127 -1442
rect -112 -1452 -96 -1438
rect -61 -1451 -39 -1432
rect -29 -1438 -13 -1437
rect -30 -1444 -13 -1438
rect -29 -1445 -13 -1444
rect -39 -1452 -33 -1451
rect -30 -1452 -1 -1445
rect -112 -1453 -1 -1452
rect -112 -1454 5 -1453
rect -436 -1462 -385 -1454
rect -338 -1462 -304 -1454
rect -436 -1474 -411 -1462
rect -404 -1474 -385 -1462
rect -331 -1464 -304 -1462
rect -295 -1464 -74 -1454
rect -39 -1457 -33 -1454
rect -331 -1468 -74 -1464
rect -436 -1482 -385 -1474
rect -338 -1482 -74 -1468
rect -30 -1462 5 -1454
rect -484 -1530 -465 -1496
rect -420 -1490 -391 -1482
rect -420 -1496 -403 -1490
rect -420 -1498 -386 -1496
rect -338 -1498 -322 -1482
rect -321 -1492 -113 -1482
rect -112 -1492 -96 -1482
rect -48 -1486 -33 -1471
rect -30 -1474 -29 -1462
rect -22 -1474 5 -1462
rect -30 -1482 5 -1474
rect -30 -1483 -1 -1482
rect -310 -1496 -96 -1492
rect -295 -1498 -96 -1496
rect -61 -1496 -48 -1486
rect -30 -1496 -13 -1483
rect -61 -1498 -13 -1496
rect -419 -1502 -386 -1498
rect -423 -1504 -386 -1502
rect -423 -1505 -356 -1504
rect -423 -1510 -392 -1505
rect -386 -1510 -356 -1505
rect -423 -1514 -356 -1510
rect -450 -1517 -356 -1514
rect -450 -1524 -401 -1517
rect -450 -1530 -420 -1524
rect -401 -1529 -396 -1524
rect -484 -1546 -404 -1530
rect -392 -1538 -356 -1517
rect -295 -1522 -106 -1498
rect -61 -1499 -14 -1498
rect -48 -1504 -14 -1499
rect -280 -1525 -106 -1522
rect -287 -1528 -106 -1525
rect -78 -1505 -14 -1504
rect -484 -1548 -465 -1546
rect -450 -1548 -416 -1546
rect -484 -1564 -404 -1548
rect -484 -1570 -465 -1564
rect -494 -1586 -465 -1570
rect -450 -1580 -420 -1564
rect -392 -1586 -386 -1538
rect -383 -1544 -364 -1538
rect -349 -1544 -319 -1536
rect -383 -1552 -319 -1544
rect -383 -1568 -303 -1552
rect -287 -1559 -225 -1528
rect -209 -1559 -147 -1528
rect -78 -1530 -29 -1505
rect -14 -1530 16 -1512
rect -115 -1544 -85 -1536
rect -78 -1538 32 -1530
rect -115 -1552 -70 -1544
rect -383 -1570 -364 -1568
rect -349 -1570 -303 -1568
rect -383 -1586 -303 -1570
rect -276 -1572 -241 -1559
rect -200 -1562 -163 -1559
rect -200 -1564 -158 -1562
rect -271 -1575 -241 -1572
rect -262 -1579 -255 -1575
rect -255 -1580 -254 -1579
rect -296 -1586 -286 -1580
rect -500 -1594 -459 -1586
rect -500 -1620 -485 -1594
rect -478 -1620 -459 -1594
rect -395 -1598 -364 -1586
rect -349 -1598 -246 -1586
rect -234 -1596 -208 -1570
rect -193 -1575 -163 -1564
rect -131 -1568 -69 -1552
rect -131 -1570 -85 -1568
rect -131 -1586 -69 -1570
rect -57 -1586 -51 -1538
rect -48 -1546 32 -1538
rect -48 -1548 -29 -1546
rect -14 -1548 20 -1546
rect -48 -1563 32 -1548
rect -48 -1564 38 -1563
rect -48 -1586 -29 -1564
rect -14 -1580 16 -1564
rect 44 -1570 50 -1496
rect 53 -1570 72 -1426
rect 87 -1570 93 -1426
rect 102 -1496 115 -1426
rect 167 -1430 189 -1426
rect 160 -1442 177 -1438
rect 181 -1440 189 -1438
rect 179 -1442 189 -1440
rect 160 -1452 189 -1442
rect 242 -1452 258 -1438
rect 296 -1442 302 -1440
rect 309 -1442 417 -1426
rect 424 -1442 430 -1440
rect 438 -1442 453 -1426
rect 519 -1432 538 -1429
rect 160 -1454 258 -1452
rect 285 -1454 453 -1442
rect 468 -1452 484 -1438
rect 519 -1451 541 -1432
rect 551 -1438 567 -1437
rect 550 -1444 567 -1438
rect 551 -1445 567 -1444
rect 541 -1452 547 -1451
rect 550 -1452 579 -1445
rect 468 -1453 579 -1452
rect 468 -1454 585 -1453
rect 144 -1462 195 -1454
rect 242 -1462 276 -1454
rect 144 -1474 169 -1462
rect 176 -1474 195 -1462
rect 249 -1464 276 -1462
rect 285 -1464 506 -1454
rect 541 -1457 547 -1454
rect 249 -1468 506 -1464
rect 144 -1482 195 -1474
rect 242 -1482 506 -1468
rect 550 -1462 585 -1454
rect 96 -1530 115 -1496
rect 160 -1490 189 -1482
rect 160 -1496 177 -1490
rect 160 -1498 194 -1496
rect 242 -1498 258 -1482
rect 259 -1492 467 -1482
rect 468 -1492 484 -1482
rect 532 -1486 547 -1471
rect 550 -1474 551 -1462
rect 558 -1474 585 -1462
rect 550 -1482 585 -1474
rect 550 -1483 579 -1482
rect 270 -1496 484 -1492
rect 285 -1498 484 -1496
rect 519 -1496 532 -1486
rect 550 -1496 567 -1483
rect 519 -1498 567 -1496
rect 161 -1502 194 -1498
rect 157 -1504 194 -1502
rect 157 -1505 224 -1504
rect 157 -1510 188 -1505
rect 194 -1510 224 -1505
rect 157 -1514 224 -1510
rect 130 -1517 224 -1514
rect 130 -1524 179 -1517
rect 130 -1530 160 -1524
rect 179 -1529 184 -1524
rect 96 -1546 176 -1530
rect 188 -1538 224 -1517
rect 285 -1522 474 -1498
rect 519 -1499 566 -1498
rect 532 -1504 566 -1499
rect 606 -1504 622 -1502
rect 300 -1525 474 -1522
rect 293 -1528 474 -1525
rect 502 -1505 566 -1504
rect 96 -1548 115 -1546
rect 130 -1548 164 -1546
rect 96 -1564 176 -1548
rect 96 -1570 115 -1564
rect -188 -1596 -85 -1586
rect -234 -1598 -85 -1596
rect -64 -1598 -29 -1586
rect -395 -1600 -233 -1598
rect -383 -1620 -364 -1600
rect -349 -1602 -319 -1600
rect -500 -1628 -459 -1620
rect -377 -1624 -364 -1620
rect -312 -1616 -233 -1600
rect -201 -1600 -29 -1598
rect -201 -1616 -122 -1600
rect -115 -1602 -85 -1600
rect -494 -1638 -465 -1628
rect -450 -1638 -420 -1624
rect -377 -1638 -334 -1624
rect -312 -1628 -122 -1616
rect -57 -1620 -51 -1600
rect -327 -1638 -297 -1628
rect -296 -1638 -138 -1628
rect -134 -1638 -104 -1628
rect -100 -1638 -70 -1624
rect -42 -1638 -29 -1600
rect 43 -1586 72 -1570
rect 86 -1586 115 -1570
rect 130 -1580 160 -1564
rect 188 -1586 194 -1538
rect 197 -1544 216 -1538
rect 231 -1544 261 -1536
rect 197 -1552 261 -1544
rect 197 -1568 277 -1552
rect 293 -1559 355 -1528
rect 371 -1559 433 -1528
rect 502 -1530 551 -1505
rect 596 -1514 622 -1504
rect 566 -1530 622 -1514
rect 465 -1544 495 -1536
rect 502 -1538 612 -1530
rect 465 -1552 510 -1544
rect 197 -1570 216 -1568
rect 231 -1570 277 -1568
rect 197 -1586 277 -1570
rect 304 -1572 339 -1559
rect 380 -1562 417 -1559
rect 380 -1564 422 -1562
rect 309 -1575 339 -1572
rect 318 -1579 325 -1575
rect 325 -1580 326 -1579
rect 284 -1586 294 -1580
rect 43 -1594 78 -1586
rect 43 -1620 44 -1594
rect 51 -1620 78 -1594
rect -14 -1638 16 -1624
rect 43 -1628 78 -1620
rect 80 -1594 121 -1586
rect 80 -1620 95 -1594
rect 102 -1620 121 -1594
rect 185 -1598 216 -1586
rect 231 -1598 334 -1586
rect 346 -1596 372 -1570
rect 387 -1575 417 -1564
rect 449 -1568 511 -1552
rect 449 -1570 495 -1568
rect 449 -1586 511 -1570
rect 523 -1586 529 -1538
rect 532 -1546 612 -1538
rect 532 -1548 551 -1546
rect 566 -1548 600 -1546
rect 532 -1564 612 -1548
rect 532 -1586 551 -1564
rect 566 -1580 596 -1564
rect 624 -1570 630 -1496
rect 633 -1570 652 -1426
rect 667 -1570 673 -1426
rect 682 -1496 695 -1426
rect 747 -1430 769 -1426
rect 740 -1442 757 -1438
rect 761 -1440 769 -1438
rect 759 -1442 769 -1440
rect 740 -1452 769 -1442
rect 822 -1452 838 -1438
rect 876 -1442 882 -1440
rect 889 -1442 997 -1426
rect 1004 -1442 1010 -1440
rect 1018 -1442 1033 -1426
rect 1099 -1432 1118 -1429
rect 740 -1454 838 -1452
rect 865 -1454 1033 -1442
rect 1048 -1452 1064 -1438
rect 1099 -1451 1121 -1432
rect 1131 -1438 1147 -1437
rect 1130 -1440 1147 -1438
rect 1131 -1445 1147 -1440
rect 1121 -1452 1127 -1451
rect 1130 -1452 1159 -1445
rect 1048 -1453 1159 -1452
rect 1048 -1454 1165 -1453
rect 724 -1462 775 -1454
rect 822 -1462 856 -1454
rect 724 -1474 749 -1462
rect 756 -1474 775 -1462
rect 829 -1464 856 -1462
rect 865 -1464 1086 -1454
rect 1121 -1457 1127 -1454
rect 829 -1468 1086 -1464
rect 724 -1482 775 -1474
rect 822 -1482 1086 -1468
rect 1130 -1462 1165 -1454
rect 676 -1530 695 -1496
rect 740 -1490 769 -1482
rect 740 -1496 757 -1490
rect 740 -1498 774 -1496
rect 822 -1498 838 -1482
rect 839 -1492 1047 -1482
rect 1048 -1492 1064 -1482
rect 1112 -1486 1127 -1471
rect 1130 -1474 1131 -1462
rect 1138 -1474 1165 -1462
rect 1130 -1482 1165 -1474
rect 1130 -1483 1159 -1482
rect 850 -1496 1064 -1492
rect 865 -1498 1064 -1496
rect 1099 -1496 1112 -1486
rect 1130 -1496 1147 -1483
rect 1099 -1498 1147 -1496
rect 741 -1502 774 -1498
rect 737 -1504 774 -1502
rect 737 -1505 804 -1504
rect 737 -1510 768 -1505
rect 774 -1510 804 -1505
rect 737 -1514 804 -1510
rect 710 -1517 804 -1514
rect 710 -1524 759 -1517
rect 710 -1530 740 -1524
rect 759 -1529 764 -1524
rect 676 -1546 756 -1530
rect 768 -1538 804 -1517
rect 865 -1522 1054 -1498
rect 1099 -1499 1146 -1498
rect 1112 -1504 1146 -1499
rect 880 -1525 1054 -1522
rect 873 -1528 1054 -1525
rect 1082 -1505 1146 -1504
rect 676 -1548 695 -1546
rect 710 -1548 744 -1546
rect 676 -1564 756 -1548
rect 676 -1570 695 -1564
rect 392 -1596 495 -1586
rect 346 -1598 495 -1596
rect 516 -1598 551 -1586
rect 185 -1600 347 -1598
rect 197 -1620 216 -1600
rect 231 -1602 261 -1600
rect 80 -1628 121 -1620
rect 203 -1624 216 -1620
rect 268 -1616 347 -1600
rect 379 -1600 551 -1598
rect 379 -1616 458 -1600
rect 465 -1602 495 -1600
rect 43 -1638 72 -1628
rect 86 -1638 115 -1628
rect 130 -1638 160 -1624
rect 203 -1638 246 -1624
rect 268 -1628 458 -1616
rect 523 -1620 529 -1600
rect 253 -1638 283 -1628
rect 284 -1638 442 -1628
rect 446 -1638 476 -1628
rect 480 -1638 510 -1624
rect 538 -1638 551 -1600
rect 623 -1586 652 -1570
rect 666 -1586 695 -1570
rect 710 -1580 740 -1564
rect 768 -1586 774 -1538
rect 777 -1544 796 -1538
rect 811 -1544 841 -1536
rect 777 -1552 841 -1544
rect 777 -1568 857 -1552
rect 873 -1559 935 -1528
rect 951 -1559 1013 -1528
rect 1082 -1530 1131 -1505
rect 1146 -1530 1176 -1512
rect 1045 -1544 1075 -1536
rect 1082 -1538 1192 -1530
rect 1045 -1552 1090 -1544
rect 777 -1570 796 -1568
rect 811 -1570 857 -1568
rect 777 -1586 857 -1570
rect 884 -1572 919 -1559
rect 960 -1562 997 -1559
rect 960 -1564 1002 -1562
rect 889 -1575 919 -1572
rect 898 -1579 905 -1575
rect 905 -1580 906 -1579
rect 864 -1586 874 -1580
rect 623 -1594 658 -1586
rect 623 -1620 624 -1594
rect 631 -1620 658 -1594
rect 566 -1638 596 -1624
rect 623 -1628 658 -1620
rect 660 -1594 701 -1586
rect 660 -1620 675 -1594
rect 682 -1620 701 -1594
rect 765 -1598 796 -1586
rect 811 -1598 914 -1586
rect 926 -1596 952 -1570
rect 967 -1575 997 -1564
rect 1029 -1568 1091 -1552
rect 1029 -1570 1075 -1568
rect 1029 -1586 1091 -1570
rect 1103 -1586 1109 -1538
rect 1112 -1546 1192 -1538
rect 1112 -1548 1131 -1546
rect 1146 -1548 1180 -1546
rect 1112 -1563 1192 -1548
rect 1112 -1564 1198 -1563
rect 1112 -1586 1131 -1564
rect 1146 -1580 1176 -1564
rect 1204 -1570 1210 -1496
rect 1213 -1570 1232 -1426
rect 1247 -1570 1253 -1426
rect 1262 -1496 1275 -1426
rect 1327 -1430 1349 -1426
rect 1320 -1442 1337 -1438
rect 1341 -1440 1349 -1438
rect 1339 -1442 1349 -1440
rect 1320 -1452 1349 -1442
rect 1402 -1452 1418 -1438
rect 1456 -1442 1462 -1440
rect 1469 -1442 1577 -1426
rect 1584 -1442 1590 -1440
rect 1598 -1442 1613 -1426
rect 1679 -1432 1698 -1429
rect 1320 -1454 1418 -1452
rect 1445 -1454 1613 -1442
rect 1628 -1452 1644 -1438
rect 1679 -1451 1701 -1432
rect 1711 -1438 1727 -1437
rect 1710 -1440 1727 -1438
rect 1711 -1445 1727 -1440
rect 1701 -1452 1707 -1451
rect 1710 -1452 1739 -1445
rect 1628 -1453 1739 -1452
rect 1628 -1454 1745 -1453
rect 1304 -1462 1355 -1454
rect 1402 -1462 1436 -1454
rect 1304 -1474 1329 -1462
rect 1336 -1474 1355 -1462
rect 1409 -1464 1436 -1462
rect 1445 -1464 1666 -1454
rect 1701 -1457 1707 -1454
rect 1409 -1468 1666 -1464
rect 1304 -1482 1355 -1474
rect 1402 -1482 1666 -1468
rect 1710 -1462 1745 -1454
rect 1256 -1530 1275 -1496
rect 1320 -1490 1349 -1482
rect 1320 -1496 1337 -1490
rect 1320 -1498 1354 -1496
rect 1402 -1498 1418 -1482
rect 1419 -1492 1627 -1482
rect 1628 -1492 1644 -1482
rect 1692 -1486 1707 -1471
rect 1710 -1474 1711 -1462
rect 1718 -1474 1745 -1462
rect 1710 -1482 1745 -1474
rect 1710 -1483 1739 -1482
rect 1430 -1496 1644 -1492
rect 1445 -1498 1644 -1496
rect 1679 -1496 1692 -1486
rect 1710 -1496 1727 -1483
rect 1679 -1498 1727 -1496
rect 1321 -1502 1354 -1498
rect 1317 -1504 1354 -1502
rect 1317 -1505 1384 -1504
rect 1317 -1510 1348 -1505
rect 1354 -1510 1384 -1505
rect 1317 -1514 1384 -1510
rect 1290 -1517 1384 -1514
rect 1290 -1524 1339 -1517
rect 1290 -1530 1320 -1524
rect 1339 -1529 1344 -1524
rect 1256 -1546 1336 -1530
rect 1348 -1538 1384 -1517
rect 1445 -1522 1634 -1498
rect 1679 -1499 1726 -1498
rect 1692 -1504 1726 -1499
rect 1766 -1504 1782 -1502
rect 1460 -1525 1634 -1522
rect 1453 -1528 1634 -1525
rect 1662 -1505 1726 -1504
rect 1256 -1548 1275 -1546
rect 1290 -1548 1324 -1546
rect 1256 -1564 1336 -1548
rect 1256 -1570 1275 -1564
rect 972 -1596 1075 -1586
rect 926 -1598 1075 -1596
rect 1096 -1598 1131 -1586
rect 765 -1600 927 -1598
rect 777 -1620 796 -1600
rect 811 -1602 841 -1600
rect 660 -1628 701 -1620
rect 783 -1624 796 -1620
rect 848 -1616 927 -1600
rect 959 -1600 1131 -1598
rect 959 -1616 1038 -1600
rect 1045 -1602 1075 -1600
rect 623 -1638 652 -1628
rect 666 -1638 695 -1628
rect 710 -1638 740 -1624
rect 783 -1638 826 -1624
rect 848 -1628 1038 -1616
rect 1103 -1620 1109 -1600
rect 833 -1638 863 -1628
rect 864 -1638 1022 -1628
rect 1026 -1638 1056 -1628
rect 1060 -1638 1090 -1624
rect 1118 -1638 1131 -1600
rect 1203 -1586 1232 -1570
rect 1246 -1586 1275 -1570
rect 1290 -1580 1320 -1564
rect 1348 -1586 1354 -1538
rect 1357 -1544 1376 -1538
rect 1391 -1544 1421 -1536
rect 1357 -1552 1421 -1544
rect 1357 -1568 1437 -1552
rect 1453 -1559 1515 -1528
rect 1531 -1559 1593 -1528
rect 1662 -1530 1711 -1505
rect 1756 -1514 1782 -1504
rect 1726 -1530 1782 -1514
rect 1625 -1544 1655 -1536
rect 1662 -1538 1772 -1530
rect 1625 -1552 1670 -1544
rect 1357 -1570 1376 -1568
rect 1391 -1570 1437 -1568
rect 1357 -1586 1437 -1570
rect 1464 -1572 1499 -1559
rect 1540 -1562 1577 -1559
rect 1540 -1564 1582 -1562
rect 1469 -1575 1499 -1572
rect 1478 -1579 1485 -1575
rect 1485 -1580 1486 -1579
rect 1444 -1586 1454 -1580
rect 1203 -1594 1238 -1586
rect 1203 -1620 1204 -1594
rect 1211 -1620 1238 -1594
rect 1146 -1638 1176 -1624
rect 1203 -1628 1238 -1620
rect 1240 -1594 1281 -1586
rect 1240 -1620 1255 -1594
rect 1262 -1620 1281 -1594
rect 1345 -1598 1376 -1586
rect 1391 -1598 1494 -1586
rect 1506 -1596 1532 -1570
rect 1547 -1575 1577 -1564
rect 1609 -1568 1671 -1552
rect 1609 -1570 1655 -1568
rect 1609 -1586 1671 -1570
rect 1683 -1586 1689 -1538
rect 1692 -1546 1772 -1538
rect 1692 -1548 1711 -1546
rect 1726 -1548 1760 -1546
rect 1692 -1564 1772 -1548
rect 1692 -1586 1711 -1564
rect 1726 -1580 1756 -1564
rect 1784 -1570 1790 -1496
rect 1793 -1570 1812 -1426
rect 1827 -1570 1833 -1426
rect 1842 -1496 1855 -1426
rect 1907 -1430 1929 -1426
rect 1900 -1442 1917 -1438
rect 1921 -1440 1929 -1438
rect 1919 -1442 1929 -1440
rect 1900 -1452 1929 -1442
rect 1982 -1452 1998 -1438
rect 2036 -1442 2042 -1440
rect 2049 -1442 2157 -1426
rect 2164 -1442 2170 -1440
rect 2178 -1442 2193 -1426
rect 2259 -1432 2278 -1429
rect 1900 -1454 1998 -1452
rect 2025 -1454 2193 -1442
rect 2208 -1452 2224 -1438
rect 2259 -1451 2281 -1432
rect 2291 -1438 2307 -1437
rect 2290 -1444 2307 -1438
rect 2291 -1445 2307 -1444
rect 2281 -1452 2287 -1451
rect 2290 -1452 2319 -1445
rect 2208 -1453 2319 -1452
rect 2208 -1454 2325 -1453
rect 1884 -1462 1935 -1454
rect 1982 -1462 2016 -1454
rect 1884 -1474 1909 -1462
rect 1916 -1474 1935 -1462
rect 1989 -1464 2016 -1462
rect 2025 -1464 2246 -1454
rect 2281 -1457 2287 -1454
rect 1989 -1468 2246 -1464
rect 1884 -1482 1935 -1474
rect 1982 -1482 2246 -1468
rect 2290 -1462 2325 -1454
rect 1836 -1530 1855 -1496
rect 1900 -1490 1929 -1482
rect 1900 -1496 1917 -1490
rect 1900 -1498 1934 -1496
rect 1982 -1498 1998 -1482
rect 1999 -1492 2207 -1482
rect 2208 -1492 2224 -1482
rect 2272 -1486 2287 -1471
rect 2290 -1474 2291 -1462
rect 2298 -1474 2325 -1462
rect 2290 -1482 2325 -1474
rect 2290 -1483 2319 -1482
rect 2010 -1496 2224 -1492
rect 2025 -1498 2224 -1496
rect 2259 -1496 2272 -1486
rect 2290 -1496 2307 -1483
rect 2259 -1498 2307 -1496
rect 1901 -1502 1934 -1498
rect 1897 -1504 1934 -1502
rect 1897 -1505 1964 -1504
rect 1897 -1510 1928 -1505
rect 1934 -1510 1964 -1505
rect 1897 -1514 1964 -1510
rect 1870 -1517 1964 -1514
rect 1870 -1524 1919 -1517
rect 1870 -1530 1900 -1524
rect 1919 -1529 1924 -1524
rect 1836 -1546 1916 -1530
rect 1928 -1538 1964 -1517
rect 2025 -1522 2214 -1498
rect 2259 -1499 2306 -1498
rect 2272 -1504 2306 -1499
rect 2040 -1525 2214 -1522
rect 2033 -1528 2214 -1525
rect 2242 -1505 2306 -1504
rect 1836 -1548 1855 -1546
rect 1870 -1548 1904 -1546
rect 1836 -1564 1916 -1548
rect 1836 -1570 1855 -1564
rect 1552 -1596 1655 -1586
rect 1506 -1598 1655 -1596
rect 1676 -1598 1711 -1586
rect 1345 -1600 1507 -1598
rect 1357 -1620 1376 -1600
rect 1391 -1602 1421 -1600
rect 1240 -1628 1281 -1620
rect 1363 -1624 1376 -1620
rect 1428 -1616 1507 -1600
rect 1539 -1600 1711 -1598
rect 1539 -1616 1618 -1600
rect 1625 -1602 1655 -1600
rect 1203 -1638 1232 -1628
rect 1246 -1638 1275 -1628
rect 1290 -1638 1320 -1624
rect 1363 -1638 1406 -1624
rect 1428 -1628 1618 -1616
rect 1683 -1620 1689 -1600
rect 1413 -1638 1443 -1628
rect 1444 -1638 1602 -1628
rect 1606 -1638 1636 -1628
rect 1640 -1638 1670 -1624
rect 1698 -1638 1711 -1600
rect 1783 -1586 1812 -1570
rect 1826 -1586 1855 -1570
rect 1870 -1580 1900 -1564
rect 1928 -1586 1934 -1538
rect 1937 -1544 1956 -1538
rect 1971 -1544 2001 -1536
rect 1937 -1552 2001 -1544
rect 1937 -1568 2017 -1552
rect 2033 -1559 2095 -1528
rect 2111 -1559 2173 -1528
rect 2242 -1530 2291 -1505
rect 2306 -1530 2336 -1512
rect 2205 -1544 2235 -1536
rect 2242 -1538 2352 -1530
rect 2205 -1552 2250 -1544
rect 1937 -1570 1956 -1568
rect 1971 -1570 2017 -1568
rect 1937 -1586 2017 -1570
rect 2044 -1572 2079 -1559
rect 2120 -1562 2157 -1559
rect 2120 -1564 2162 -1562
rect 2049 -1575 2079 -1572
rect 2058 -1579 2065 -1575
rect 2065 -1580 2066 -1579
rect 2024 -1586 2034 -1580
rect 1783 -1594 1818 -1586
rect 1783 -1620 1784 -1594
rect 1791 -1620 1818 -1594
rect 1726 -1638 1756 -1624
rect 1783 -1628 1818 -1620
rect 1820 -1594 1861 -1586
rect 1820 -1620 1835 -1594
rect 1842 -1620 1861 -1594
rect 1925 -1598 1956 -1586
rect 1971 -1598 2074 -1586
rect 2086 -1596 2112 -1570
rect 2127 -1575 2157 -1564
rect 2189 -1568 2251 -1552
rect 2189 -1570 2235 -1568
rect 2189 -1586 2251 -1570
rect 2263 -1586 2269 -1538
rect 2272 -1546 2352 -1538
rect 2272 -1548 2291 -1546
rect 2306 -1548 2340 -1546
rect 2272 -1563 2352 -1548
rect 2272 -1564 2358 -1563
rect 2272 -1586 2291 -1564
rect 2306 -1580 2336 -1564
rect 2364 -1570 2370 -1496
rect 2373 -1570 2392 -1426
rect 2407 -1570 2413 -1426
rect 2422 -1496 2435 -1426
rect 2487 -1430 2509 -1426
rect 2480 -1442 2497 -1438
rect 2501 -1440 2509 -1438
rect 2499 -1442 2509 -1440
rect 2480 -1452 2509 -1442
rect 2562 -1452 2578 -1438
rect 2616 -1442 2622 -1440
rect 2629 -1442 2737 -1426
rect 2744 -1442 2750 -1440
rect 2758 -1442 2773 -1426
rect 2839 -1432 2858 -1429
rect 2480 -1454 2578 -1452
rect 2605 -1454 2773 -1442
rect 2788 -1452 2804 -1438
rect 2839 -1451 2861 -1432
rect 2871 -1438 2887 -1437
rect 2870 -1444 2887 -1438
rect 2871 -1445 2887 -1444
rect 2861 -1452 2867 -1451
rect 2870 -1452 2899 -1445
rect 2788 -1453 2899 -1452
rect 2788 -1454 2905 -1453
rect 2464 -1462 2515 -1454
rect 2562 -1462 2596 -1454
rect 2464 -1474 2489 -1462
rect 2496 -1474 2515 -1462
rect 2569 -1464 2596 -1462
rect 2605 -1464 2826 -1454
rect 2861 -1457 2867 -1454
rect 2569 -1468 2826 -1464
rect 2464 -1482 2515 -1474
rect 2562 -1482 2826 -1468
rect 2870 -1462 2905 -1454
rect 2416 -1530 2435 -1496
rect 2480 -1490 2509 -1482
rect 2480 -1496 2497 -1490
rect 2480 -1498 2514 -1496
rect 2562 -1498 2578 -1482
rect 2579 -1492 2787 -1482
rect 2788 -1492 2804 -1482
rect 2852 -1486 2867 -1471
rect 2870 -1474 2871 -1462
rect 2878 -1474 2905 -1462
rect 2870 -1482 2905 -1474
rect 2870 -1483 2899 -1482
rect 2590 -1496 2804 -1492
rect 2605 -1498 2804 -1496
rect 2839 -1496 2852 -1486
rect 2870 -1496 2887 -1483
rect 2839 -1498 2887 -1496
rect 2481 -1502 2514 -1498
rect 2477 -1504 2514 -1502
rect 2477 -1505 2544 -1504
rect 2477 -1510 2508 -1505
rect 2514 -1510 2544 -1505
rect 2477 -1514 2544 -1510
rect 2450 -1517 2544 -1514
rect 2450 -1524 2499 -1517
rect 2450 -1530 2480 -1524
rect 2499 -1529 2504 -1524
rect 2416 -1546 2496 -1530
rect 2508 -1538 2544 -1517
rect 2605 -1522 2794 -1498
rect 2839 -1499 2886 -1498
rect 2852 -1504 2886 -1499
rect 2926 -1504 2942 -1502
rect 2620 -1525 2794 -1522
rect 2613 -1528 2794 -1525
rect 2822 -1505 2886 -1504
rect 2416 -1548 2435 -1546
rect 2450 -1548 2484 -1546
rect 2416 -1564 2496 -1548
rect 2416 -1570 2435 -1564
rect 2132 -1596 2235 -1586
rect 2086 -1598 2235 -1596
rect 2256 -1598 2291 -1586
rect 1925 -1600 2087 -1598
rect 1937 -1620 1956 -1600
rect 1971 -1602 2001 -1600
rect 1820 -1628 1861 -1620
rect 1943 -1624 1956 -1620
rect 2008 -1616 2087 -1600
rect 2119 -1600 2291 -1598
rect 2119 -1616 2198 -1600
rect 2205 -1602 2235 -1600
rect 1783 -1638 1812 -1628
rect 1826 -1638 1855 -1628
rect 1870 -1638 1900 -1624
rect 1943 -1638 1986 -1624
rect 2008 -1628 2198 -1616
rect 2263 -1620 2269 -1600
rect 1993 -1638 2023 -1628
rect 2024 -1638 2182 -1628
rect 2186 -1638 2216 -1628
rect 2220 -1638 2250 -1624
rect 2278 -1638 2291 -1600
rect 2363 -1586 2392 -1570
rect 2406 -1586 2435 -1570
rect 2450 -1580 2480 -1564
rect 2508 -1586 2514 -1538
rect 2517 -1544 2536 -1538
rect 2551 -1544 2581 -1536
rect 2517 -1552 2581 -1544
rect 2517 -1568 2597 -1552
rect 2613 -1559 2675 -1528
rect 2691 -1559 2753 -1528
rect 2822 -1530 2871 -1505
rect 2916 -1514 2942 -1504
rect 2886 -1530 2942 -1514
rect 2785 -1544 2815 -1536
rect 2822 -1538 2932 -1530
rect 2785 -1552 2830 -1544
rect 2517 -1570 2536 -1568
rect 2551 -1570 2597 -1568
rect 2517 -1586 2597 -1570
rect 2624 -1572 2659 -1559
rect 2700 -1562 2737 -1559
rect 2700 -1564 2742 -1562
rect 2629 -1575 2659 -1572
rect 2638 -1579 2645 -1575
rect 2645 -1580 2646 -1579
rect 2604 -1586 2614 -1580
rect 2363 -1594 2398 -1586
rect 2363 -1620 2364 -1594
rect 2371 -1620 2398 -1594
rect 2306 -1638 2336 -1624
rect 2363 -1628 2398 -1620
rect 2400 -1594 2441 -1586
rect 2400 -1620 2415 -1594
rect 2422 -1620 2441 -1594
rect 2505 -1598 2536 -1586
rect 2551 -1598 2654 -1586
rect 2666 -1596 2692 -1570
rect 2707 -1575 2737 -1564
rect 2769 -1568 2831 -1552
rect 2769 -1570 2815 -1568
rect 2769 -1586 2831 -1570
rect 2843 -1586 2849 -1538
rect 2852 -1546 2932 -1538
rect 2852 -1548 2871 -1546
rect 2886 -1548 2920 -1546
rect 2852 -1564 2932 -1548
rect 2852 -1586 2871 -1564
rect 2886 -1580 2916 -1564
rect 2944 -1570 2950 -1496
rect 2953 -1570 2972 -1426
rect 2987 -1570 2993 -1426
rect 3002 -1496 3015 -1426
rect 3067 -1430 3089 -1426
rect 3060 -1442 3077 -1438
rect 3081 -1440 3089 -1438
rect 3079 -1442 3089 -1440
rect 3060 -1452 3089 -1442
rect 3142 -1452 3158 -1438
rect 3196 -1442 3202 -1440
rect 3209 -1442 3317 -1426
rect 3324 -1442 3330 -1440
rect 3338 -1442 3353 -1426
rect 3419 -1432 3438 -1429
rect 3060 -1454 3158 -1452
rect 3185 -1454 3353 -1442
rect 3368 -1452 3384 -1438
rect 3419 -1451 3441 -1432
rect 3451 -1438 3467 -1437
rect 3450 -1444 3467 -1438
rect 3451 -1445 3467 -1444
rect 3441 -1452 3447 -1451
rect 3450 -1452 3479 -1445
rect 3368 -1453 3479 -1452
rect 3368 -1454 3485 -1453
rect 3044 -1462 3095 -1454
rect 3142 -1462 3176 -1454
rect 3044 -1474 3069 -1462
rect 3076 -1474 3095 -1462
rect 3149 -1464 3176 -1462
rect 3185 -1464 3406 -1454
rect 3441 -1457 3447 -1454
rect 3149 -1468 3406 -1464
rect 3044 -1482 3095 -1474
rect 3142 -1482 3406 -1468
rect 3450 -1462 3485 -1454
rect 2996 -1530 3015 -1496
rect 3060 -1490 3089 -1482
rect 3060 -1496 3077 -1490
rect 3060 -1498 3094 -1496
rect 3142 -1498 3158 -1482
rect 3159 -1492 3367 -1482
rect 3368 -1492 3384 -1482
rect 3432 -1486 3447 -1471
rect 3450 -1474 3451 -1462
rect 3458 -1474 3485 -1462
rect 3450 -1482 3485 -1474
rect 3450 -1483 3479 -1482
rect 3170 -1496 3384 -1492
rect 3185 -1498 3384 -1496
rect 3419 -1496 3432 -1486
rect 3450 -1496 3467 -1483
rect 3419 -1498 3467 -1496
rect 3061 -1502 3094 -1498
rect 3057 -1504 3094 -1502
rect 3057 -1505 3124 -1504
rect 3057 -1510 3088 -1505
rect 3094 -1510 3124 -1505
rect 3057 -1514 3124 -1510
rect 3030 -1517 3124 -1514
rect 3030 -1524 3079 -1517
rect 3030 -1530 3060 -1524
rect 3079 -1529 3084 -1524
rect 2996 -1546 3076 -1530
rect 3088 -1538 3124 -1517
rect 3185 -1522 3374 -1498
rect 3419 -1499 3466 -1498
rect 3432 -1504 3466 -1499
rect 3200 -1525 3374 -1522
rect 3193 -1528 3374 -1525
rect 3402 -1505 3466 -1504
rect 2996 -1548 3015 -1546
rect 3030 -1548 3064 -1546
rect 2996 -1564 3076 -1548
rect 2996 -1570 3015 -1564
rect 2712 -1596 2815 -1586
rect 2666 -1598 2815 -1596
rect 2836 -1598 2871 -1586
rect 2505 -1600 2667 -1598
rect 2517 -1620 2536 -1600
rect 2551 -1602 2581 -1600
rect 2400 -1628 2441 -1620
rect 2523 -1624 2536 -1620
rect 2588 -1616 2667 -1600
rect 2699 -1600 2871 -1598
rect 2699 -1616 2778 -1600
rect 2785 -1602 2815 -1600
rect 2363 -1638 2392 -1628
rect 2406 -1638 2435 -1628
rect 2450 -1638 2480 -1624
rect 2523 -1638 2566 -1624
rect 2588 -1628 2778 -1616
rect 2843 -1620 2849 -1600
rect 2573 -1638 2603 -1628
rect 2604 -1638 2762 -1628
rect 2766 -1638 2796 -1628
rect 2800 -1638 2830 -1624
rect 2858 -1638 2871 -1600
rect 2943 -1586 2972 -1570
rect 2986 -1586 3015 -1570
rect 3030 -1580 3060 -1564
rect 3088 -1586 3094 -1538
rect 3097 -1544 3116 -1538
rect 3131 -1544 3161 -1536
rect 3097 -1552 3161 -1544
rect 3097 -1568 3177 -1552
rect 3193 -1559 3255 -1528
rect 3271 -1559 3333 -1528
rect 3402 -1530 3451 -1505
rect 3466 -1530 3496 -1512
rect 3365 -1544 3395 -1536
rect 3402 -1538 3512 -1530
rect 3365 -1552 3410 -1544
rect 3097 -1570 3116 -1568
rect 3131 -1570 3177 -1568
rect 3097 -1586 3177 -1570
rect 3204 -1572 3239 -1559
rect 3280 -1562 3317 -1559
rect 3280 -1564 3322 -1562
rect 3209 -1575 3239 -1572
rect 3218 -1579 3225 -1575
rect 3225 -1580 3226 -1579
rect 3184 -1586 3194 -1580
rect 2943 -1594 2978 -1586
rect 2943 -1620 2944 -1594
rect 2951 -1620 2978 -1594
rect 2886 -1638 2916 -1624
rect 2943 -1628 2978 -1620
rect 2980 -1594 3021 -1586
rect 2980 -1620 2995 -1594
rect 3002 -1620 3021 -1594
rect 3085 -1598 3116 -1586
rect 3131 -1598 3234 -1586
rect 3246 -1596 3272 -1570
rect 3287 -1575 3317 -1564
rect 3349 -1568 3411 -1552
rect 3349 -1570 3395 -1568
rect 3349 -1586 3411 -1570
rect 3423 -1586 3429 -1538
rect 3432 -1546 3512 -1538
rect 3432 -1548 3451 -1546
rect 3466 -1548 3500 -1546
rect 3432 -1563 3512 -1548
rect 3432 -1564 3518 -1563
rect 3432 -1586 3451 -1564
rect 3466 -1580 3496 -1564
rect 3524 -1570 3530 -1496
rect 3533 -1570 3552 -1426
rect 3567 -1570 3573 -1426
rect 3582 -1496 3595 -1426
rect 3647 -1430 3669 -1426
rect 3640 -1442 3657 -1438
rect 3661 -1440 3669 -1438
rect 3659 -1442 3669 -1440
rect 3640 -1452 3669 -1442
rect 3722 -1452 3738 -1438
rect 3776 -1442 3782 -1440
rect 3789 -1442 3897 -1426
rect 3904 -1442 3910 -1440
rect 3918 -1442 3933 -1426
rect 3999 -1432 4018 -1429
rect 3640 -1454 3738 -1452
rect 3765 -1454 3933 -1442
rect 3948 -1452 3964 -1438
rect 3999 -1451 4021 -1432
rect 4031 -1438 4047 -1437
rect 4030 -1444 4047 -1438
rect 4031 -1445 4047 -1444
rect 4021 -1452 4027 -1451
rect 4030 -1452 4059 -1445
rect 3948 -1453 4059 -1452
rect 3948 -1454 4065 -1453
rect 3624 -1462 3675 -1454
rect 3722 -1462 3756 -1454
rect 3624 -1474 3649 -1462
rect 3656 -1474 3675 -1462
rect 3729 -1464 3756 -1462
rect 3765 -1464 3986 -1454
rect 4021 -1457 4027 -1454
rect 3729 -1468 3986 -1464
rect 3624 -1482 3675 -1474
rect 3722 -1482 3986 -1468
rect 4030 -1462 4065 -1454
rect 3576 -1530 3595 -1496
rect 3640 -1490 3669 -1482
rect 3640 -1496 3657 -1490
rect 3640 -1498 3674 -1496
rect 3722 -1498 3738 -1482
rect 3739 -1492 3947 -1482
rect 3948 -1492 3964 -1482
rect 4012 -1486 4027 -1471
rect 4030 -1474 4031 -1462
rect 4038 -1474 4065 -1462
rect 4030 -1482 4065 -1474
rect 4030 -1483 4059 -1482
rect 3750 -1496 3964 -1492
rect 3765 -1498 3964 -1496
rect 3999 -1496 4012 -1486
rect 4030 -1496 4047 -1483
rect 3999 -1498 4047 -1496
rect 3641 -1502 3674 -1498
rect 3637 -1504 3674 -1502
rect 3637 -1505 3704 -1504
rect 3637 -1510 3668 -1505
rect 3674 -1510 3704 -1505
rect 3637 -1514 3704 -1510
rect 3610 -1517 3704 -1514
rect 3610 -1524 3659 -1517
rect 3610 -1530 3640 -1524
rect 3659 -1529 3664 -1524
rect 3576 -1546 3656 -1530
rect 3668 -1538 3704 -1517
rect 3765 -1522 3954 -1498
rect 3999 -1499 4046 -1498
rect 4012 -1504 4046 -1499
rect 4086 -1504 4102 -1502
rect 3780 -1525 3954 -1522
rect 3773 -1528 3954 -1525
rect 3982 -1505 4046 -1504
rect 3576 -1548 3595 -1546
rect 3610 -1548 3644 -1546
rect 3576 -1564 3656 -1548
rect 3576 -1570 3595 -1564
rect 3292 -1596 3395 -1586
rect 3246 -1598 3395 -1596
rect 3416 -1598 3451 -1586
rect 3085 -1600 3247 -1598
rect 3097 -1620 3116 -1600
rect 3131 -1602 3161 -1600
rect 2980 -1628 3021 -1620
rect 3103 -1624 3116 -1620
rect 3168 -1616 3247 -1600
rect 3279 -1600 3451 -1598
rect 3279 -1616 3358 -1600
rect 3365 -1602 3395 -1600
rect 2943 -1638 2972 -1628
rect 2986 -1638 3015 -1628
rect 3030 -1638 3060 -1624
rect 3103 -1638 3146 -1624
rect 3168 -1628 3358 -1616
rect 3423 -1620 3429 -1600
rect 3153 -1638 3183 -1628
rect 3184 -1638 3342 -1628
rect 3346 -1638 3376 -1628
rect 3380 -1638 3410 -1624
rect 3438 -1638 3451 -1600
rect 3523 -1586 3552 -1570
rect 3566 -1586 3595 -1570
rect 3610 -1580 3640 -1564
rect 3668 -1586 3674 -1538
rect 3677 -1544 3696 -1538
rect 3711 -1544 3741 -1536
rect 3677 -1552 3741 -1544
rect 3677 -1568 3757 -1552
rect 3773 -1559 3835 -1528
rect 3851 -1559 3913 -1528
rect 3982 -1530 4031 -1505
rect 4076 -1514 4102 -1504
rect 4046 -1530 4102 -1514
rect 3945 -1544 3975 -1536
rect 3982 -1538 4092 -1530
rect 3945 -1552 3990 -1544
rect 3677 -1570 3696 -1568
rect 3711 -1570 3757 -1568
rect 3677 -1586 3757 -1570
rect 3784 -1572 3819 -1559
rect 3860 -1562 3897 -1559
rect 3860 -1564 3902 -1562
rect 3789 -1575 3819 -1572
rect 3798 -1579 3805 -1575
rect 3805 -1580 3806 -1579
rect 3764 -1586 3774 -1580
rect 3523 -1594 3558 -1586
rect 3523 -1620 3524 -1594
rect 3531 -1620 3558 -1594
rect 3466 -1638 3496 -1624
rect 3523 -1628 3558 -1620
rect 3560 -1594 3601 -1586
rect 3560 -1620 3575 -1594
rect 3582 -1620 3601 -1594
rect 3665 -1598 3696 -1586
rect 3711 -1598 3814 -1586
rect 3826 -1596 3852 -1570
rect 3867 -1575 3897 -1564
rect 3929 -1568 3991 -1552
rect 3929 -1570 3975 -1568
rect 3929 -1586 3991 -1570
rect 4003 -1586 4009 -1538
rect 4012 -1546 4092 -1538
rect 4012 -1548 4031 -1546
rect 4046 -1548 4080 -1546
rect 4012 -1564 4092 -1548
rect 4012 -1586 4031 -1564
rect 4046 -1580 4076 -1564
rect 4104 -1570 4110 -1496
rect 4113 -1570 4132 -1426
rect 4147 -1570 4153 -1426
rect 4162 -1496 4175 -1426
rect 4227 -1430 4249 -1426
rect 4220 -1442 4237 -1438
rect 4241 -1440 4249 -1438
rect 4239 -1442 4249 -1440
rect 4220 -1452 4249 -1442
rect 4302 -1452 4318 -1438
rect 4356 -1442 4362 -1440
rect 4369 -1442 4477 -1426
rect 4484 -1442 4490 -1440
rect 4498 -1442 4513 -1426
rect 4579 -1432 4598 -1429
rect 4220 -1454 4318 -1452
rect 4345 -1454 4513 -1442
rect 4528 -1452 4544 -1438
rect 4579 -1451 4601 -1432
rect 4611 -1438 4627 -1437
rect 4610 -1444 4627 -1438
rect 4611 -1445 4627 -1444
rect 4601 -1452 4607 -1451
rect 4610 -1452 4639 -1445
rect 4528 -1453 4639 -1452
rect 4528 -1454 4645 -1453
rect 4204 -1462 4255 -1454
rect 4302 -1462 4336 -1454
rect 4204 -1474 4229 -1462
rect 4236 -1474 4255 -1462
rect 4309 -1464 4336 -1462
rect 4345 -1464 4566 -1454
rect 4601 -1457 4607 -1454
rect 4309 -1468 4566 -1464
rect 4204 -1482 4255 -1474
rect 4302 -1482 4566 -1468
rect 4610 -1462 4645 -1454
rect 4156 -1530 4175 -1496
rect 4220 -1490 4249 -1482
rect 4220 -1496 4237 -1490
rect 4220 -1498 4254 -1496
rect 4302 -1498 4318 -1482
rect 4319 -1492 4527 -1482
rect 4528 -1492 4544 -1482
rect 4592 -1486 4607 -1471
rect 4610 -1474 4611 -1462
rect 4618 -1474 4645 -1462
rect 4610 -1482 4645 -1474
rect 4610 -1483 4639 -1482
rect 4330 -1496 4544 -1492
rect 4345 -1498 4544 -1496
rect 4579 -1496 4592 -1486
rect 4610 -1496 4627 -1483
rect 4579 -1498 4627 -1496
rect 4221 -1502 4254 -1498
rect 4217 -1504 4254 -1502
rect 4217 -1505 4284 -1504
rect 4217 -1510 4248 -1505
rect 4254 -1510 4284 -1505
rect 4217 -1514 4284 -1510
rect 4190 -1517 4284 -1514
rect 4190 -1524 4239 -1517
rect 4190 -1530 4220 -1524
rect 4239 -1529 4244 -1524
rect 4156 -1546 4236 -1530
rect 4248 -1538 4284 -1517
rect 4345 -1522 4534 -1498
rect 4579 -1499 4626 -1498
rect 4592 -1504 4626 -1499
rect 4360 -1525 4534 -1522
rect 4353 -1528 4534 -1525
rect 4562 -1505 4626 -1504
rect 4156 -1548 4175 -1546
rect 4190 -1548 4224 -1546
rect 4156 -1564 4236 -1548
rect 4156 -1570 4175 -1564
rect 3872 -1596 3975 -1586
rect 3826 -1598 3975 -1596
rect 3996 -1598 4031 -1586
rect 3665 -1600 3827 -1598
rect 3677 -1620 3696 -1600
rect 3711 -1602 3741 -1600
rect 3560 -1628 3601 -1620
rect 3683 -1624 3696 -1620
rect 3748 -1616 3827 -1600
rect 3859 -1600 4031 -1598
rect 3859 -1616 3938 -1600
rect 3945 -1602 3975 -1600
rect 3523 -1638 3552 -1628
rect 3566 -1638 3595 -1628
rect 3610 -1638 3640 -1624
rect 3683 -1638 3726 -1624
rect 3748 -1628 3938 -1616
rect 4003 -1620 4009 -1600
rect 3733 -1638 3763 -1628
rect 3764 -1638 3922 -1628
rect 3926 -1638 3956 -1628
rect 3960 -1638 3990 -1624
rect 4018 -1638 4031 -1600
rect 4103 -1586 4132 -1570
rect 4146 -1586 4175 -1570
rect 4190 -1580 4220 -1564
rect 4248 -1586 4254 -1538
rect 4257 -1544 4276 -1538
rect 4291 -1544 4321 -1536
rect 4257 -1552 4321 -1544
rect 4257 -1568 4337 -1552
rect 4353 -1559 4415 -1528
rect 4431 -1559 4493 -1528
rect 4562 -1530 4611 -1505
rect 4626 -1530 4656 -1512
rect 4525 -1544 4555 -1536
rect 4562 -1538 4672 -1530
rect 4525 -1552 4570 -1544
rect 4257 -1570 4276 -1568
rect 4291 -1570 4337 -1568
rect 4257 -1586 4337 -1570
rect 4364 -1572 4399 -1559
rect 4440 -1562 4477 -1559
rect 4440 -1564 4482 -1562
rect 4369 -1575 4399 -1572
rect 4378 -1579 4385 -1575
rect 4385 -1580 4386 -1579
rect 4344 -1586 4354 -1580
rect 4103 -1594 4138 -1586
rect 4103 -1620 4104 -1594
rect 4111 -1620 4138 -1594
rect 4046 -1638 4076 -1624
rect 4103 -1628 4138 -1620
rect 4140 -1594 4181 -1586
rect 4140 -1620 4155 -1594
rect 4162 -1620 4181 -1594
rect 4245 -1598 4276 -1586
rect 4291 -1598 4394 -1586
rect 4406 -1596 4432 -1570
rect 4447 -1575 4477 -1564
rect 4509 -1568 4571 -1552
rect 4509 -1570 4555 -1568
rect 4509 -1586 4571 -1570
rect 4583 -1586 4589 -1538
rect 4592 -1546 4672 -1538
rect 4592 -1548 4611 -1546
rect 4626 -1548 4660 -1546
rect 4592 -1563 4672 -1548
rect 4592 -1564 4678 -1563
rect 4592 -1586 4611 -1564
rect 4626 -1580 4656 -1564
rect 4684 -1570 4690 -1496
rect 4693 -1570 4712 -1426
rect 4727 -1570 4733 -1426
rect 4742 -1496 4755 -1426
rect 4807 -1430 4829 -1426
rect 4800 -1442 4817 -1438
rect 4821 -1440 4829 -1438
rect 4819 -1442 4829 -1440
rect 4800 -1452 4829 -1442
rect 4882 -1452 4898 -1438
rect 4936 -1442 4942 -1440
rect 4949 -1442 5057 -1426
rect 5064 -1442 5070 -1440
rect 5078 -1442 5093 -1426
rect 5159 -1432 5178 -1429
rect 4800 -1454 4898 -1452
rect 4925 -1454 5093 -1442
rect 5108 -1452 5124 -1438
rect 5159 -1451 5181 -1432
rect 5191 -1438 5207 -1437
rect 5190 -1444 5207 -1438
rect 5191 -1445 5207 -1444
rect 5181 -1452 5187 -1451
rect 5190 -1452 5219 -1445
rect 5108 -1453 5219 -1452
rect 5108 -1454 5225 -1453
rect 4784 -1462 4835 -1454
rect 4882 -1462 4916 -1454
rect 4784 -1474 4809 -1462
rect 4816 -1474 4835 -1462
rect 4889 -1464 4916 -1462
rect 4925 -1464 5146 -1454
rect 5181 -1457 5187 -1454
rect 4889 -1468 5146 -1464
rect 4784 -1482 4835 -1474
rect 4882 -1482 5146 -1468
rect 5190 -1462 5225 -1454
rect 4736 -1530 4755 -1496
rect 4800 -1490 4829 -1482
rect 4800 -1496 4817 -1490
rect 4800 -1498 4834 -1496
rect 4882 -1498 4898 -1482
rect 4899 -1492 5107 -1482
rect 5108 -1492 5124 -1482
rect 5172 -1486 5187 -1471
rect 5190 -1474 5191 -1462
rect 5198 -1474 5225 -1462
rect 5190 -1482 5225 -1474
rect 5190 -1483 5219 -1482
rect 4910 -1496 5124 -1492
rect 4925 -1498 5124 -1496
rect 5159 -1496 5172 -1486
rect 5190 -1496 5207 -1483
rect 5159 -1498 5207 -1496
rect 4801 -1502 4834 -1498
rect 4797 -1504 4834 -1502
rect 4797 -1505 4864 -1504
rect 4797 -1510 4828 -1505
rect 4834 -1510 4864 -1505
rect 4797 -1514 4864 -1510
rect 4770 -1517 4864 -1514
rect 4770 -1524 4819 -1517
rect 4770 -1530 4800 -1524
rect 4819 -1529 4824 -1524
rect 4736 -1546 4816 -1530
rect 4828 -1538 4864 -1517
rect 4925 -1522 5114 -1498
rect 5159 -1499 5206 -1498
rect 5172 -1504 5206 -1499
rect 5246 -1504 5262 -1502
rect 4940 -1525 5114 -1522
rect 4933 -1528 5114 -1525
rect 5142 -1505 5206 -1504
rect 4736 -1548 4755 -1546
rect 4770 -1548 4804 -1546
rect 4736 -1564 4816 -1548
rect 4736 -1570 4755 -1564
rect 4452 -1596 4555 -1586
rect 4406 -1598 4555 -1596
rect 4576 -1598 4611 -1586
rect 4245 -1600 4407 -1598
rect 4257 -1620 4276 -1600
rect 4291 -1602 4321 -1600
rect 4140 -1628 4181 -1620
rect 4263 -1624 4276 -1620
rect 4328 -1616 4407 -1600
rect 4439 -1600 4611 -1598
rect 4439 -1616 4518 -1600
rect 4525 -1602 4555 -1600
rect 4103 -1638 4132 -1628
rect 4146 -1638 4175 -1628
rect 4190 -1638 4220 -1624
rect 4263 -1638 4306 -1624
rect 4328 -1628 4518 -1616
rect 4583 -1620 4589 -1600
rect 4313 -1638 4343 -1628
rect 4344 -1638 4502 -1628
rect 4506 -1638 4536 -1628
rect 4540 -1638 4570 -1624
rect 4598 -1638 4611 -1600
rect 4683 -1586 4712 -1570
rect 4726 -1586 4755 -1570
rect 4770 -1580 4800 -1564
rect 4828 -1586 4834 -1538
rect 4837 -1544 4856 -1538
rect 4871 -1544 4901 -1536
rect 4837 -1552 4901 -1544
rect 4837 -1568 4917 -1552
rect 4933 -1559 4995 -1528
rect 5011 -1559 5073 -1528
rect 5142 -1530 5191 -1505
rect 5236 -1514 5262 -1504
rect 5206 -1530 5262 -1514
rect 5105 -1544 5135 -1536
rect 5142 -1538 5252 -1530
rect 5105 -1552 5150 -1544
rect 4837 -1570 4856 -1568
rect 4871 -1570 4917 -1568
rect 4837 -1586 4917 -1570
rect 4944 -1572 4979 -1559
rect 5020 -1562 5057 -1559
rect 5020 -1564 5062 -1562
rect 4949 -1575 4979 -1572
rect 4958 -1579 4965 -1575
rect 4965 -1580 4966 -1579
rect 4924 -1586 4934 -1580
rect 4683 -1594 4718 -1586
rect 4683 -1620 4684 -1594
rect 4691 -1620 4718 -1594
rect 4626 -1638 4656 -1624
rect 4683 -1628 4718 -1620
rect 4720 -1594 4761 -1586
rect 4720 -1620 4735 -1594
rect 4742 -1620 4761 -1594
rect 4825 -1598 4856 -1586
rect 4871 -1598 4974 -1586
rect 4986 -1596 5012 -1570
rect 5027 -1575 5057 -1564
rect 5089 -1568 5151 -1552
rect 5089 -1570 5135 -1568
rect 5089 -1586 5151 -1570
rect 5163 -1586 5169 -1538
rect 5172 -1546 5252 -1538
rect 5172 -1548 5191 -1546
rect 5206 -1548 5240 -1546
rect 5172 -1564 5252 -1548
rect 5172 -1586 5191 -1564
rect 5206 -1580 5236 -1564
rect 5264 -1570 5270 -1496
rect 5273 -1570 5292 -1426
rect 5307 -1570 5313 -1426
rect 5322 -1496 5335 -1426
rect 5387 -1430 5409 -1426
rect 5380 -1442 5397 -1438
rect 5401 -1440 5409 -1438
rect 5399 -1442 5409 -1440
rect 5380 -1452 5409 -1442
rect 5462 -1452 5478 -1438
rect 5516 -1442 5522 -1440
rect 5529 -1442 5637 -1426
rect 5644 -1442 5650 -1440
rect 5658 -1442 5673 -1426
rect 5739 -1432 5758 -1429
rect 5380 -1454 5478 -1452
rect 5505 -1454 5673 -1442
rect 5688 -1452 5704 -1438
rect 5739 -1451 5761 -1432
rect 5771 -1438 5787 -1437
rect 5770 -1444 5787 -1438
rect 5771 -1445 5787 -1444
rect 5761 -1452 5767 -1451
rect 5770 -1452 5799 -1445
rect 5688 -1453 5799 -1452
rect 5688 -1454 5805 -1453
rect 5364 -1462 5415 -1454
rect 5462 -1462 5496 -1454
rect 5364 -1474 5389 -1462
rect 5396 -1474 5415 -1462
rect 5469 -1464 5496 -1462
rect 5505 -1464 5726 -1454
rect 5761 -1457 5767 -1454
rect 5469 -1468 5726 -1464
rect 5364 -1482 5415 -1474
rect 5462 -1482 5726 -1468
rect 5770 -1462 5805 -1454
rect 5316 -1530 5335 -1496
rect 5380 -1490 5409 -1482
rect 5380 -1496 5397 -1490
rect 5380 -1498 5414 -1496
rect 5462 -1498 5478 -1482
rect 5479 -1492 5687 -1482
rect 5688 -1492 5704 -1482
rect 5752 -1486 5767 -1471
rect 5770 -1474 5771 -1462
rect 5778 -1474 5805 -1462
rect 5770 -1482 5805 -1474
rect 5770 -1483 5799 -1482
rect 5490 -1496 5704 -1492
rect 5505 -1498 5704 -1496
rect 5739 -1496 5752 -1486
rect 5770 -1496 5787 -1483
rect 5739 -1498 5787 -1496
rect 5381 -1502 5414 -1498
rect 5377 -1504 5414 -1502
rect 5377 -1505 5444 -1504
rect 5377 -1510 5408 -1505
rect 5414 -1510 5444 -1505
rect 5377 -1514 5444 -1510
rect 5350 -1517 5444 -1514
rect 5350 -1524 5399 -1517
rect 5350 -1530 5380 -1524
rect 5399 -1529 5404 -1524
rect 5316 -1546 5396 -1530
rect 5408 -1538 5444 -1517
rect 5505 -1522 5694 -1498
rect 5739 -1499 5786 -1498
rect 5752 -1504 5786 -1499
rect 5520 -1525 5694 -1522
rect 5513 -1528 5694 -1525
rect 5722 -1505 5786 -1504
rect 5316 -1548 5335 -1546
rect 5350 -1548 5384 -1546
rect 5316 -1564 5396 -1548
rect 5316 -1570 5335 -1564
rect 5032 -1596 5135 -1586
rect 4986 -1598 5135 -1596
rect 5156 -1598 5191 -1586
rect 4825 -1600 4987 -1598
rect 4837 -1620 4856 -1600
rect 4871 -1602 4901 -1600
rect 4720 -1628 4761 -1620
rect 4843 -1624 4856 -1620
rect 4908 -1616 4987 -1600
rect 5019 -1600 5191 -1598
rect 5019 -1616 5098 -1600
rect 5105 -1602 5135 -1600
rect 4683 -1638 4712 -1628
rect 4726 -1638 4755 -1628
rect 4770 -1638 4800 -1624
rect 4843 -1638 4886 -1624
rect 4908 -1628 5098 -1616
rect 5163 -1620 5169 -1600
rect 4893 -1638 4923 -1628
rect 4924 -1638 5082 -1628
rect 5086 -1638 5116 -1628
rect 5120 -1638 5150 -1624
rect 5178 -1638 5191 -1600
rect 5263 -1586 5292 -1570
rect 5306 -1586 5335 -1570
rect 5350 -1580 5380 -1564
rect 5408 -1586 5414 -1538
rect 5417 -1544 5436 -1538
rect 5451 -1544 5481 -1536
rect 5417 -1552 5481 -1544
rect 5417 -1568 5497 -1552
rect 5513 -1559 5575 -1528
rect 5591 -1559 5653 -1528
rect 5722 -1530 5771 -1505
rect 5786 -1530 5816 -1512
rect 5685 -1544 5715 -1536
rect 5722 -1538 5832 -1530
rect 5685 -1552 5730 -1544
rect 5417 -1570 5436 -1568
rect 5451 -1570 5497 -1568
rect 5417 -1586 5497 -1570
rect 5524 -1572 5559 -1559
rect 5600 -1562 5637 -1559
rect 5600 -1564 5642 -1562
rect 5529 -1575 5559 -1572
rect 5538 -1579 5545 -1575
rect 5545 -1580 5546 -1579
rect 5504 -1586 5514 -1580
rect 5263 -1594 5298 -1586
rect 5263 -1620 5264 -1594
rect 5271 -1620 5298 -1594
rect 5206 -1638 5236 -1624
rect 5263 -1628 5298 -1620
rect 5300 -1594 5341 -1586
rect 5300 -1620 5315 -1594
rect 5322 -1620 5341 -1594
rect 5405 -1598 5436 -1586
rect 5451 -1598 5554 -1586
rect 5566 -1596 5592 -1570
rect 5607 -1575 5637 -1564
rect 5669 -1568 5731 -1552
rect 5669 -1570 5715 -1568
rect 5669 -1586 5731 -1570
rect 5743 -1586 5749 -1538
rect 5752 -1546 5832 -1538
rect 5752 -1548 5771 -1546
rect 5786 -1548 5820 -1546
rect 5752 -1563 5832 -1548
rect 5752 -1564 5838 -1563
rect 5752 -1586 5771 -1564
rect 5786 -1580 5816 -1564
rect 5844 -1570 5850 -1496
rect 5853 -1570 5872 -1426
rect 5887 -1570 5893 -1426
rect 5902 -1496 5915 -1426
rect 5967 -1430 5989 -1426
rect 5960 -1442 5977 -1438
rect 5981 -1440 5989 -1438
rect 5979 -1442 5989 -1440
rect 5960 -1452 5989 -1442
rect 6042 -1452 6058 -1438
rect 6096 -1442 6102 -1440
rect 6109 -1442 6217 -1426
rect 6224 -1442 6230 -1440
rect 6238 -1442 6253 -1426
rect 6319 -1432 6338 -1429
rect 5960 -1454 6058 -1452
rect 6085 -1454 6253 -1442
rect 6268 -1452 6284 -1438
rect 6319 -1451 6341 -1432
rect 6351 -1438 6367 -1437
rect 6350 -1444 6367 -1438
rect 6351 -1445 6367 -1444
rect 6341 -1452 6347 -1451
rect 6350 -1452 6379 -1445
rect 6268 -1453 6379 -1452
rect 6268 -1454 6385 -1453
rect 5944 -1462 5995 -1454
rect 6042 -1462 6076 -1454
rect 5944 -1474 5969 -1462
rect 5976 -1474 5995 -1462
rect 6049 -1464 6076 -1462
rect 6085 -1464 6306 -1454
rect 6341 -1457 6347 -1454
rect 6049 -1468 6306 -1464
rect 5944 -1482 5995 -1474
rect 6042 -1482 6306 -1468
rect 6350 -1462 6385 -1454
rect 5896 -1530 5915 -1496
rect 5960 -1490 5989 -1482
rect 5960 -1496 5977 -1490
rect 5960 -1498 5994 -1496
rect 6042 -1498 6058 -1482
rect 6059 -1492 6267 -1482
rect 6268 -1492 6284 -1482
rect 6332 -1486 6347 -1471
rect 6350 -1474 6351 -1462
rect 6358 -1474 6385 -1462
rect 6350 -1482 6385 -1474
rect 6350 -1483 6379 -1482
rect 6070 -1496 6284 -1492
rect 6085 -1498 6284 -1496
rect 6319 -1496 6332 -1486
rect 6350 -1496 6367 -1483
rect 6319 -1498 6367 -1496
rect 5961 -1502 5994 -1498
rect 5957 -1504 5994 -1502
rect 5957 -1505 6024 -1504
rect 5957 -1510 5988 -1505
rect 5994 -1510 6024 -1505
rect 5957 -1514 6024 -1510
rect 5930 -1517 6024 -1514
rect 5930 -1524 5979 -1517
rect 5930 -1530 5960 -1524
rect 5979 -1529 5984 -1524
rect 5896 -1546 5976 -1530
rect 5988 -1538 6024 -1517
rect 6085 -1522 6274 -1498
rect 6319 -1499 6366 -1498
rect 6332 -1504 6366 -1499
rect 6100 -1525 6274 -1522
rect 6093 -1528 6274 -1525
rect 6302 -1505 6366 -1504
rect 5896 -1548 5915 -1546
rect 5930 -1548 5964 -1546
rect 5896 -1564 5976 -1548
rect 5896 -1570 5915 -1564
rect 5612 -1596 5715 -1586
rect 5566 -1598 5715 -1596
rect 5736 -1598 5771 -1586
rect 5405 -1600 5567 -1598
rect 5417 -1620 5436 -1600
rect 5451 -1602 5481 -1600
rect 5300 -1628 5341 -1620
rect 5423 -1624 5436 -1620
rect 5488 -1616 5567 -1600
rect 5599 -1600 5771 -1598
rect 5599 -1616 5678 -1600
rect 5685 -1602 5715 -1600
rect 5263 -1638 5292 -1628
rect 5306 -1638 5335 -1628
rect 5350 -1638 5380 -1624
rect 5423 -1638 5466 -1624
rect 5488 -1628 5678 -1616
rect 5743 -1620 5749 -1600
rect 5473 -1638 5503 -1628
rect 5504 -1638 5662 -1628
rect 5666 -1638 5696 -1628
rect 5700 -1638 5730 -1624
rect 5758 -1638 5771 -1600
rect 5843 -1586 5872 -1570
rect 5886 -1586 5915 -1570
rect 5930 -1580 5960 -1564
rect 5988 -1586 5994 -1538
rect 5997 -1544 6016 -1538
rect 6031 -1544 6061 -1536
rect 5997 -1552 6061 -1544
rect 5997 -1568 6077 -1552
rect 6093 -1559 6155 -1528
rect 6171 -1559 6233 -1528
rect 6302 -1530 6351 -1505
rect 6366 -1530 6396 -1514
rect 6265 -1544 6295 -1536
rect 6302 -1538 6412 -1530
rect 6265 -1552 6310 -1544
rect 5997 -1570 6016 -1568
rect 6031 -1570 6077 -1568
rect 5997 -1586 6077 -1570
rect 6104 -1572 6139 -1559
rect 6180 -1562 6217 -1559
rect 6180 -1564 6222 -1562
rect 6109 -1575 6139 -1572
rect 6118 -1579 6125 -1575
rect 6125 -1580 6126 -1579
rect 6084 -1586 6094 -1580
rect 5843 -1594 5878 -1586
rect 5843 -1620 5844 -1594
rect 5851 -1620 5878 -1594
rect 5786 -1638 5816 -1624
rect 5843 -1628 5878 -1620
rect 5880 -1594 5921 -1586
rect 5880 -1620 5895 -1594
rect 5902 -1620 5921 -1594
rect 5985 -1598 6016 -1586
rect 6031 -1598 6134 -1586
rect 6146 -1596 6172 -1570
rect 6187 -1575 6217 -1564
rect 6249 -1568 6311 -1552
rect 6249 -1570 6295 -1568
rect 6249 -1586 6311 -1570
rect 6323 -1586 6329 -1538
rect 6332 -1546 6412 -1538
rect 6332 -1548 6351 -1546
rect 6366 -1548 6400 -1546
rect 6332 -1564 6412 -1548
rect 6332 -1586 6351 -1564
rect 6366 -1580 6396 -1564
rect 6424 -1570 6430 -1496
rect 6439 -1570 6452 -1426
rect 6192 -1596 6295 -1586
rect 6146 -1598 6295 -1596
rect 6316 -1598 6351 -1586
rect 5985 -1600 6147 -1598
rect 5997 -1620 6016 -1600
rect 6031 -1602 6061 -1600
rect 5880 -1628 5921 -1620
rect 6003 -1624 6016 -1620
rect 6068 -1616 6147 -1600
rect 6179 -1600 6351 -1598
rect 6179 -1616 6258 -1600
rect 6265 -1602 6295 -1600
rect 5843 -1638 5872 -1628
rect 5886 -1638 5915 -1628
rect 5930 -1638 5960 -1624
rect 6003 -1638 6046 -1624
rect 6068 -1628 6258 -1616
rect 6323 -1620 6329 -1600
rect 6053 -1638 6083 -1628
rect 6084 -1638 6242 -1628
rect 6246 -1638 6276 -1628
rect 6280 -1638 6310 -1624
rect 6338 -1638 6351 -1600
rect 6423 -1586 6452 -1570
rect 6423 -1594 6458 -1586
rect 6423 -1620 6424 -1594
rect 6431 -1620 6458 -1594
rect 6366 -1638 6396 -1624
rect 6423 -1628 6458 -1620
rect 6423 -1638 6452 -1628
rect -541 -1652 6452 -1638
rect -478 -1682 -465 -1652
rect -450 -1666 -420 -1652
rect -377 -1666 -334 -1652
rect -327 -1666 -107 -1652
rect -100 -1666 -70 -1652
rect -410 -1680 -395 -1668
rect -376 -1680 -363 -1666
rect -295 -1670 -142 -1666
rect -413 -1682 -391 -1680
rect -313 -1682 -121 -1670
rect -42 -1682 -29 -1652
rect -14 -1666 16 -1652
rect 53 -1682 72 -1652
rect 87 -1682 93 -1652
rect 102 -1682 115 -1652
rect 130 -1666 160 -1652
rect 203 -1666 246 -1652
rect 253 -1666 473 -1652
rect 480 -1666 510 -1652
rect 170 -1680 185 -1668
rect 204 -1680 217 -1666
rect 285 -1670 438 -1666
rect 167 -1682 189 -1680
rect 267 -1682 459 -1670
rect 538 -1682 551 -1652
rect 566 -1666 596 -1652
rect 633 -1682 652 -1652
rect 667 -1682 673 -1652
rect 682 -1682 695 -1652
rect 710 -1666 740 -1652
rect 783 -1666 826 -1652
rect 833 -1666 1053 -1652
rect 1060 -1666 1090 -1652
rect 750 -1680 765 -1668
rect 784 -1680 797 -1666
rect 865 -1670 1018 -1666
rect 747 -1682 769 -1680
rect 847 -1682 1039 -1670
rect 1118 -1682 1131 -1652
rect 1146 -1666 1176 -1652
rect 1213 -1682 1232 -1652
rect 1247 -1682 1253 -1652
rect 1262 -1682 1275 -1652
rect 1290 -1666 1320 -1652
rect 1363 -1666 1406 -1652
rect 1413 -1666 1633 -1652
rect 1640 -1666 1670 -1652
rect 1330 -1680 1345 -1668
rect 1364 -1680 1377 -1666
rect 1445 -1670 1598 -1666
rect 1327 -1682 1349 -1680
rect 1427 -1682 1619 -1670
rect 1698 -1682 1711 -1652
rect 1726 -1666 1756 -1652
rect 1793 -1682 1812 -1652
rect 1827 -1682 1833 -1652
rect 1842 -1682 1855 -1652
rect 1870 -1666 1900 -1652
rect 1943 -1666 1986 -1652
rect 1993 -1666 2213 -1652
rect 2220 -1666 2250 -1652
rect 1910 -1680 1925 -1668
rect 1944 -1680 1957 -1666
rect 2025 -1670 2178 -1666
rect 1907 -1682 1929 -1680
rect 2007 -1682 2199 -1670
rect 2278 -1682 2291 -1652
rect 2306 -1666 2336 -1652
rect 2373 -1682 2392 -1652
rect 2407 -1682 2413 -1652
rect 2422 -1682 2435 -1652
rect 2450 -1666 2480 -1652
rect 2523 -1666 2566 -1652
rect 2573 -1666 2793 -1652
rect 2800 -1666 2830 -1652
rect 2490 -1680 2505 -1668
rect 2524 -1680 2537 -1666
rect 2605 -1670 2758 -1666
rect 2487 -1682 2509 -1680
rect 2587 -1682 2779 -1670
rect 2858 -1682 2871 -1652
rect 2886 -1666 2916 -1652
rect 2953 -1682 2972 -1652
rect 2987 -1682 2993 -1652
rect 3002 -1682 3015 -1652
rect 3030 -1666 3060 -1652
rect 3103 -1666 3146 -1652
rect 3153 -1666 3373 -1652
rect 3380 -1666 3410 -1652
rect 3070 -1680 3085 -1668
rect 3104 -1680 3117 -1666
rect 3185 -1670 3338 -1666
rect 3067 -1682 3089 -1680
rect 3167 -1682 3359 -1670
rect 3438 -1682 3451 -1652
rect 3466 -1666 3496 -1652
rect 3533 -1682 3552 -1652
rect 3567 -1682 3573 -1652
rect 3582 -1682 3595 -1652
rect 3610 -1666 3640 -1652
rect 3683 -1666 3726 -1652
rect 3733 -1666 3953 -1652
rect 3960 -1666 3990 -1652
rect 3650 -1680 3665 -1668
rect 3684 -1680 3697 -1666
rect 3765 -1670 3918 -1666
rect 3647 -1682 3669 -1680
rect 3747 -1682 3939 -1670
rect 4018 -1682 4031 -1652
rect 4046 -1666 4076 -1652
rect 4113 -1682 4132 -1652
rect 4147 -1682 4153 -1652
rect 4162 -1682 4175 -1652
rect 4190 -1666 4220 -1652
rect 4263 -1666 4306 -1652
rect 4313 -1666 4533 -1652
rect 4540 -1666 4570 -1652
rect 4230 -1680 4245 -1668
rect 4264 -1680 4277 -1666
rect 4345 -1670 4498 -1666
rect 4227 -1682 4249 -1680
rect 4327 -1682 4519 -1670
rect 4598 -1682 4611 -1652
rect 4626 -1666 4656 -1652
rect 4693 -1682 4712 -1652
rect 4727 -1682 4733 -1652
rect 4742 -1682 4755 -1652
rect 4770 -1666 4800 -1652
rect 4843 -1666 4886 -1652
rect 4893 -1666 5113 -1652
rect 5120 -1666 5150 -1652
rect 4810 -1680 4825 -1668
rect 4844 -1680 4857 -1666
rect 4925 -1670 5078 -1666
rect 4807 -1682 4829 -1680
rect 4907 -1682 5099 -1670
rect 5178 -1682 5191 -1652
rect 5206 -1666 5236 -1652
rect 5273 -1682 5292 -1652
rect 5307 -1682 5313 -1652
rect 5322 -1682 5335 -1652
rect 5350 -1666 5380 -1652
rect 5423 -1666 5466 -1652
rect 5473 -1666 5693 -1652
rect 5700 -1666 5730 -1652
rect 5390 -1680 5405 -1668
rect 5424 -1680 5437 -1666
rect 5505 -1670 5658 -1666
rect 5387 -1682 5409 -1680
rect 5487 -1682 5679 -1670
rect 5758 -1682 5771 -1652
rect 5786 -1666 5816 -1652
rect 5853 -1682 5872 -1652
rect 5887 -1682 5893 -1652
rect 5902 -1682 5915 -1652
rect 5930 -1666 5960 -1652
rect 6003 -1666 6046 -1652
rect 6053 -1666 6273 -1652
rect 6280 -1666 6310 -1652
rect 5970 -1680 5985 -1668
rect 6004 -1680 6017 -1666
rect 6085 -1670 6238 -1666
rect 5967 -1682 5989 -1680
rect 6067 -1682 6259 -1670
rect 6338 -1682 6351 -1652
rect 6366 -1666 6396 -1652
rect 6439 -1682 6452 -1652
rect -541 -1696 6452 -1682
rect -478 -1766 -465 -1696
rect -413 -1700 -391 -1696
rect -420 -1712 -403 -1708
rect -399 -1710 -391 -1708
rect -401 -1712 -391 -1710
rect -420 -1722 -391 -1712
rect -338 -1722 -322 -1708
rect -284 -1712 -278 -1710
rect -271 -1712 -163 -1696
rect -156 -1712 -150 -1710
rect -142 -1712 -127 -1696
rect -61 -1702 -42 -1699
rect -420 -1724 -322 -1722
rect -295 -1724 -127 -1712
rect -112 -1722 -96 -1708
rect -61 -1721 -39 -1702
rect -29 -1708 -13 -1707
rect -30 -1710 -13 -1708
rect -29 -1715 -13 -1710
rect -39 -1722 -33 -1721
rect -30 -1722 -1 -1715
rect -112 -1723 -1 -1722
rect -112 -1724 5 -1723
rect -436 -1732 -385 -1724
rect -338 -1732 -304 -1724
rect -436 -1744 -411 -1732
rect -404 -1744 -385 -1732
rect -331 -1734 -304 -1732
rect -295 -1734 -74 -1724
rect -39 -1727 -33 -1724
rect -331 -1738 -74 -1734
rect -436 -1752 -385 -1744
rect -338 -1752 -74 -1738
rect -30 -1732 5 -1724
rect -484 -1800 -465 -1766
rect -420 -1760 -391 -1752
rect -420 -1766 -403 -1760
rect -420 -1768 -386 -1766
rect -338 -1768 -322 -1752
rect -321 -1762 -113 -1752
rect -112 -1762 -96 -1752
rect -48 -1756 -33 -1741
rect -30 -1744 -29 -1732
rect -22 -1744 5 -1732
rect -30 -1752 5 -1744
rect -30 -1753 -1 -1752
rect -310 -1766 -96 -1762
rect -295 -1768 -96 -1766
rect -61 -1766 -48 -1756
rect -30 -1766 -13 -1753
rect -61 -1768 -13 -1766
rect -419 -1772 -386 -1768
rect -423 -1774 -386 -1772
rect -423 -1775 -356 -1774
rect -423 -1780 -392 -1775
rect -386 -1780 -356 -1775
rect -423 -1784 -356 -1780
rect -450 -1787 -356 -1784
rect -450 -1794 -401 -1787
rect -450 -1800 -420 -1794
rect -401 -1799 -396 -1794
rect -484 -1816 -404 -1800
rect -392 -1808 -356 -1787
rect -295 -1792 -106 -1768
rect -61 -1769 -14 -1768
rect -48 -1774 -14 -1769
rect -280 -1795 -106 -1792
rect -287 -1798 -106 -1795
rect -78 -1775 -14 -1774
rect -484 -1818 -465 -1816
rect -450 -1818 -416 -1816
rect -484 -1834 -404 -1818
rect -484 -1840 -465 -1834
rect -494 -1856 -465 -1840
rect -450 -1850 -420 -1834
rect -392 -1856 -386 -1808
rect -383 -1814 -364 -1808
rect -349 -1814 -319 -1806
rect -383 -1822 -319 -1814
rect -383 -1838 -303 -1822
rect -287 -1829 -225 -1798
rect -209 -1829 -147 -1798
rect -78 -1800 -29 -1775
rect -14 -1800 16 -1782
rect -115 -1814 -85 -1806
rect -78 -1808 32 -1800
rect -115 -1822 -70 -1814
rect -383 -1840 -364 -1838
rect -349 -1840 -303 -1838
rect -383 -1856 -303 -1840
rect -276 -1842 -241 -1829
rect -200 -1832 -163 -1829
rect -200 -1834 -158 -1832
rect -271 -1845 -241 -1842
rect -262 -1849 -255 -1845
rect -255 -1850 -254 -1849
rect -296 -1856 -286 -1850
rect -500 -1864 -459 -1856
rect -500 -1890 -485 -1864
rect -478 -1890 -459 -1864
rect -395 -1868 -364 -1856
rect -349 -1868 -246 -1856
rect -234 -1866 -208 -1840
rect -193 -1845 -163 -1834
rect -131 -1838 -69 -1822
rect -131 -1840 -85 -1838
rect -131 -1856 -69 -1840
rect -57 -1856 -51 -1808
rect -48 -1816 32 -1808
rect -48 -1818 -29 -1816
rect -14 -1818 20 -1816
rect -48 -1833 32 -1818
rect -48 -1834 38 -1833
rect -48 -1856 -29 -1834
rect -14 -1850 16 -1834
rect 44 -1840 50 -1766
rect 53 -1840 72 -1696
rect 87 -1840 93 -1696
rect 102 -1766 115 -1696
rect 167 -1700 189 -1696
rect 160 -1712 177 -1708
rect 181 -1710 189 -1708
rect 179 -1712 189 -1710
rect 160 -1722 189 -1712
rect 242 -1722 258 -1708
rect 296 -1712 302 -1710
rect 309 -1712 417 -1696
rect 424 -1712 430 -1710
rect 438 -1712 453 -1696
rect 519 -1702 538 -1699
rect 160 -1724 258 -1722
rect 285 -1724 453 -1712
rect 468 -1722 484 -1708
rect 519 -1721 541 -1702
rect 551 -1708 567 -1707
rect 550 -1710 567 -1708
rect 551 -1715 567 -1710
rect 541 -1722 547 -1721
rect 550 -1722 579 -1715
rect 468 -1723 579 -1722
rect 468 -1724 585 -1723
rect 144 -1732 195 -1724
rect 242 -1732 276 -1724
rect 144 -1744 169 -1732
rect 176 -1744 195 -1732
rect 249 -1734 276 -1732
rect 285 -1734 506 -1724
rect 541 -1727 547 -1724
rect 249 -1738 506 -1734
rect 144 -1752 195 -1744
rect 242 -1752 506 -1738
rect 550 -1732 585 -1724
rect 96 -1800 115 -1766
rect 160 -1760 189 -1752
rect 160 -1766 177 -1760
rect 160 -1768 194 -1766
rect 242 -1768 258 -1752
rect 259 -1762 467 -1752
rect 468 -1762 484 -1752
rect 532 -1756 547 -1741
rect 550 -1744 551 -1732
rect 558 -1744 585 -1732
rect 550 -1752 585 -1744
rect 550 -1753 579 -1752
rect 270 -1766 484 -1762
rect 285 -1768 484 -1766
rect 519 -1766 532 -1756
rect 550 -1766 567 -1753
rect 519 -1768 567 -1766
rect 161 -1772 194 -1768
rect 157 -1774 194 -1772
rect 157 -1775 224 -1774
rect 157 -1780 188 -1775
rect 194 -1780 224 -1775
rect 157 -1784 224 -1780
rect 130 -1787 224 -1784
rect 130 -1794 179 -1787
rect 130 -1800 160 -1794
rect 179 -1799 184 -1794
rect 96 -1816 176 -1800
rect 188 -1808 224 -1787
rect 285 -1792 474 -1768
rect 519 -1769 566 -1768
rect 532 -1774 566 -1769
rect 606 -1774 622 -1772
rect 300 -1795 474 -1792
rect 293 -1798 474 -1795
rect 502 -1775 566 -1774
rect 96 -1818 115 -1816
rect 130 -1818 164 -1816
rect 96 -1834 176 -1818
rect 96 -1840 115 -1834
rect -188 -1866 -85 -1856
rect -234 -1868 -85 -1866
rect -64 -1868 -29 -1856
rect -395 -1870 -233 -1868
rect -383 -1888 -364 -1870
rect -349 -1872 -319 -1870
rect -500 -1898 -459 -1890
rect -376 -1894 -364 -1888
rect -312 -1888 -233 -1870
rect -201 -1870 -29 -1868
rect -201 -1886 -122 -1870
rect -115 -1872 -85 -1870
rect -226 -1888 -122 -1886
rect -494 -1908 -465 -1898
rect -450 -1908 -420 -1894
rect -376 -1908 -334 -1894
rect -312 -1898 -122 -1888
rect -57 -1890 -51 -1870
rect -327 -1908 -297 -1898
rect -296 -1908 -138 -1898
rect -134 -1908 -104 -1898
rect -100 -1908 -70 -1894
rect -42 -1908 -29 -1870
rect 43 -1856 72 -1840
rect 86 -1856 115 -1840
rect 130 -1850 160 -1834
rect 188 -1856 194 -1808
rect 197 -1814 216 -1808
rect 231 -1814 261 -1806
rect 197 -1822 261 -1814
rect 197 -1838 277 -1822
rect 293 -1829 355 -1798
rect 371 -1829 433 -1798
rect 502 -1800 551 -1775
rect 596 -1784 622 -1774
rect 566 -1800 622 -1784
rect 465 -1814 495 -1806
rect 502 -1808 612 -1800
rect 465 -1822 510 -1814
rect 197 -1840 216 -1838
rect 231 -1840 277 -1838
rect 197 -1856 277 -1840
rect 304 -1842 339 -1829
rect 380 -1832 417 -1829
rect 380 -1834 422 -1832
rect 309 -1845 339 -1842
rect 318 -1849 325 -1845
rect 325 -1850 326 -1849
rect 284 -1856 294 -1850
rect 43 -1864 78 -1856
rect 43 -1890 44 -1864
rect 51 -1890 78 -1864
rect -14 -1908 16 -1894
rect 43 -1898 78 -1890
rect 80 -1864 121 -1856
rect 80 -1890 95 -1864
rect 102 -1890 121 -1864
rect 185 -1868 216 -1856
rect 231 -1868 334 -1856
rect 346 -1866 372 -1840
rect 387 -1845 417 -1834
rect 449 -1838 511 -1822
rect 449 -1840 495 -1838
rect 449 -1856 511 -1840
rect 523 -1856 529 -1808
rect 532 -1816 612 -1808
rect 532 -1818 551 -1816
rect 566 -1818 600 -1816
rect 532 -1834 612 -1818
rect 532 -1856 551 -1834
rect 566 -1850 596 -1834
rect 624 -1840 630 -1766
rect 633 -1840 652 -1696
rect 667 -1840 673 -1696
rect 682 -1766 695 -1696
rect 747 -1700 769 -1696
rect 740 -1712 757 -1708
rect 761 -1710 769 -1708
rect 759 -1712 769 -1710
rect 740 -1722 769 -1712
rect 822 -1722 838 -1708
rect 876 -1712 882 -1710
rect 889 -1712 997 -1696
rect 1004 -1712 1010 -1710
rect 1018 -1712 1033 -1696
rect 1099 -1702 1118 -1699
rect 740 -1724 838 -1722
rect 865 -1724 1033 -1712
rect 1048 -1722 1064 -1708
rect 1099 -1721 1121 -1702
rect 1131 -1708 1147 -1707
rect 1130 -1710 1147 -1708
rect 1131 -1715 1147 -1710
rect 1121 -1722 1127 -1721
rect 1130 -1722 1159 -1715
rect 1048 -1723 1159 -1722
rect 1048 -1724 1165 -1723
rect 724 -1732 775 -1724
rect 822 -1732 856 -1724
rect 724 -1744 749 -1732
rect 756 -1744 775 -1732
rect 829 -1734 856 -1732
rect 865 -1734 1086 -1724
rect 1121 -1727 1127 -1724
rect 829 -1738 1086 -1734
rect 724 -1752 775 -1744
rect 822 -1752 1086 -1738
rect 1130 -1732 1165 -1724
rect 676 -1800 695 -1766
rect 740 -1760 769 -1752
rect 740 -1766 757 -1760
rect 740 -1768 774 -1766
rect 822 -1768 838 -1752
rect 839 -1762 1047 -1752
rect 1048 -1762 1064 -1752
rect 1112 -1756 1127 -1741
rect 1130 -1744 1131 -1732
rect 1138 -1744 1165 -1732
rect 1130 -1752 1165 -1744
rect 1130 -1753 1159 -1752
rect 850 -1766 1064 -1762
rect 865 -1768 1064 -1766
rect 1099 -1766 1112 -1756
rect 1130 -1766 1147 -1753
rect 1099 -1768 1147 -1766
rect 741 -1772 774 -1768
rect 737 -1774 774 -1772
rect 737 -1775 804 -1774
rect 737 -1780 768 -1775
rect 774 -1780 804 -1775
rect 737 -1784 804 -1780
rect 710 -1787 804 -1784
rect 710 -1794 759 -1787
rect 710 -1800 740 -1794
rect 759 -1799 764 -1794
rect 676 -1816 756 -1800
rect 768 -1808 804 -1787
rect 865 -1792 1054 -1768
rect 1099 -1769 1146 -1768
rect 1112 -1774 1146 -1769
rect 880 -1795 1054 -1792
rect 873 -1798 1054 -1795
rect 1082 -1775 1146 -1774
rect 676 -1818 695 -1816
rect 710 -1818 744 -1816
rect 676 -1834 756 -1818
rect 676 -1840 695 -1834
rect 392 -1866 495 -1856
rect 346 -1868 495 -1866
rect 516 -1868 551 -1856
rect 185 -1870 347 -1868
rect 197 -1888 216 -1870
rect 231 -1872 261 -1870
rect 80 -1898 121 -1890
rect 204 -1894 216 -1888
rect 268 -1888 347 -1870
rect 379 -1870 551 -1868
rect 379 -1886 458 -1870
rect 465 -1872 495 -1870
rect 354 -1888 458 -1886
rect 43 -1908 72 -1898
rect 86 -1908 115 -1898
rect 130 -1908 160 -1894
rect 204 -1908 246 -1894
rect 268 -1898 458 -1888
rect 523 -1890 529 -1870
rect 253 -1908 283 -1898
rect 284 -1908 442 -1898
rect 446 -1908 476 -1898
rect 480 -1908 510 -1894
rect 538 -1908 551 -1870
rect 623 -1856 652 -1840
rect 666 -1856 695 -1840
rect 710 -1850 740 -1834
rect 768 -1856 774 -1808
rect 777 -1814 796 -1808
rect 811 -1814 841 -1806
rect 777 -1822 841 -1814
rect 777 -1838 857 -1822
rect 873 -1829 935 -1798
rect 951 -1829 1013 -1798
rect 1082 -1800 1131 -1775
rect 1146 -1800 1176 -1782
rect 1045 -1814 1075 -1806
rect 1082 -1808 1192 -1800
rect 1045 -1822 1090 -1814
rect 777 -1840 796 -1838
rect 811 -1840 857 -1838
rect 777 -1856 857 -1840
rect 884 -1842 919 -1829
rect 960 -1832 997 -1829
rect 960 -1834 1002 -1832
rect 889 -1845 919 -1842
rect 898 -1849 905 -1845
rect 905 -1850 906 -1849
rect 864 -1856 874 -1850
rect 623 -1864 658 -1856
rect 623 -1890 624 -1864
rect 631 -1890 658 -1864
rect 566 -1908 596 -1894
rect 623 -1898 658 -1890
rect 660 -1864 701 -1856
rect 660 -1890 675 -1864
rect 682 -1890 701 -1864
rect 765 -1868 796 -1856
rect 811 -1868 914 -1856
rect 926 -1866 952 -1840
rect 967 -1845 997 -1834
rect 1029 -1838 1091 -1822
rect 1029 -1840 1075 -1838
rect 1029 -1856 1091 -1840
rect 1103 -1856 1109 -1808
rect 1112 -1816 1192 -1808
rect 1112 -1818 1131 -1816
rect 1146 -1818 1180 -1816
rect 1112 -1833 1192 -1818
rect 1112 -1834 1198 -1833
rect 1112 -1856 1131 -1834
rect 1146 -1850 1176 -1834
rect 1204 -1840 1210 -1766
rect 1213 -1840 1232 -1696
rect 1247 -1840 1253 -1696
rect 1262 -1766 1275 -1696
rect 1327 -1700 1349 -1696
rect 1320 -1712 1337 -1708
rect 1341 -1710 1349 -1708
rect 1339 -1712 1349 -1710
rect 1320 -1722 1349 -1712
rect 1402 -1722 1418 -1708
rect 1456 -1712 1462 -1710
rect 1469 -1712 1577 -1696
rect 1584 -1712 1590 -1710
rect 1598 -1712 1613 -1696
rect 1679 -1702 1698 -1699
rect 1320 -1724 1418 -1722
rect 1445 -1724 1613 -1712
rect 1628 -1722 1644 -1708
rect 1679 -1721 1701 -1702
rect 1711 -1708 1727 -1707
rect 1710 -1710 1727 -1708
rect 1711 -1715 1727 -1710
rect 1701 -1722 1707 -1721
rect 1710 -1722 1739 -1715
rect 1628 -1723 1739 -1722
rect 1628 -1724 1745 -1723
rect 1304 -1732 1355 -1724
rect 1402 -1732 1436 -1724
rect 1304 -1744 1329 -1732
rect 1336 -1744 1355 -1732
rect 1409 -1734 1436 -1732
rect 1445 -1734 1666 -1724
rect 1701 -1727 1707 -1724
rect 1409 -1738 1666 -1734
rect 1304 -1752 1355 -1744
rect 1402 -1752 1666 -1738
rect 1710 -1732 1745 -1724
rect 1256 -1800 1275 -1766
rect 1320 -1760 1349 -1752
rect 1320 -1766 1337 -1760
rect 1320 -1768 1354 -1766
rect 1402 -1768 1418 -1752
rect 1419 -1762 1627 -1752
rect 1628 -1762 1644 -1752
rect 1692 -1756 1707 -1741
rect 1710 -1744 1711 -1732
rect 1718 -1744 1745 -1732
rect 1710 -1752 1745 -1744
rect 1710 -1753 1739 -1752
rect 1430 -1766 1644 -1762
rect 1445 -1768 1644 -1766
rect 1679 -1766 1692 -1756
rect 1710 -1766 1727 -1753
rect 1679 -1768 1727 -1766
rect 1321 -1772 1354 -1768
rect 1317 -1774 1354 -1772
rect 1317 -1775 1384 -1774
rect 1317 -1780 1348 -1775
rect 1354 -1780 1384 -1775
rect 1317 -1784 1384 -1780
rect 1290 -1787 1384 -1784
rect 1290 -1794 1339 -1787
rect 1290 -1800 1320 -1794
rect 1339 -1799 1344 -1794
rect 1256 -1816 1336 -1800
rect 1348 -1808 1384 -1787
rect 1445 -1792 1634 -1768
rect 1679 -1769 1726 -1768
rect 1692 -1774 1726 -1769
rect 1766 -1774 1782 -1772
rect 1460 -1795 1634 -1792
rect 1453 -1798 1634 -1795
rect 1662 -1775 1726 -1774
rect 1256 -1818 1275 -1816
rect 1290 -1818 1324 -1816
rect 1256 -1834 1336 -1818
rect 1256 -1840 1275 -1834
rect 972 -1866 1075 -1856
rect 926 -1868 1075 -1866
rect 1096 -1868 1131 -1856
rect 765 -1870 927 -1868
rect 777 -1888 796 -1870
rect 811 -1872 841 -1870
rect 660 -1898 701 -1890
rect 784 -1894 796 -1888
rect 848 -1888 927 -1870
rect 959 -1870 1131 -1868
rect 959 -1886 1038 -1870
rect 1045 -1872 1075 -1870
rect 934 -1888 1038 -1886
rect 623 -1908 652 -1898
rect 666 -1908 695 -1898
rect 710 -1908 740 -1894
rect 784 -1908 826 -1894
rect 848 -1898 1038 -1888
rect 1103 -1890 1109 -1870
rect 833 -1908 863 -1898
rect 864 -1908 1022 -1898
rect 1026 -1908 1056 -1898
rect 1060 -1908 1090 -1894
rect 1118 -1908 1131 -1870
rect 1203 -1856 1232 -1840
rect 1246 -1856 1275 -1840
rect 1290 -1850 1320 -1834
rect 1348 -1856 1354 -1808
rect 1357 -1814 1376 -1808
rect 1391 -1814 1421 -1806
rect 1357 -1822 1421 -1814
rect 1357 -1838 1437 -1822
rect 1453 -1829 1515 -1798
rect 1531 -1829 1593 -1798
rect 1662 -1800 1711 -1775
rect 1756 -1784 1782 -1774
rect 1726 -1800 1782 -1784
rect 1625 -1814 1655 -1806
rect 1662 -1808 1772 -1800
rect 1625 -1822 1670 -1814
rect 1357 -1840 1376 -1838
rect 1391 -1840 1437 -1838
rect 1357 -1856 1437 -1840
rect 1464 -1842 1499 -1829
rect 1540 -1832 1577 -1829
rect 1540 -1834 1582 -1832
rect 1469 -1845 1499 -1842
rect 1478 -1849 1485 -1845
rect 1485 -1850 1486 -1849
rect 1444 -1856 1454 -1850
rect 1203 -1864 1238 -1856
rect 1203 -1890 1204 -1864
rect 1211 -1890 1238 -1864
rect 1146 -1908 1176 -1894
rect 1203 -1898 1238 -1890
rect 1240 -1864 1281 -1856
rect 1240 -1890 1255 -1864
rect 1262 -1890 1281 -1864
rect 1345 -1868 1376 -1856
rect 1391 -1868 1494 -1856
rect 1506 -1866 1532 -1840
rect 1547 -1845 1577 -1834
rect 1609 -1838 1671 -1822
rect 1609 -1840 1655 -1838
rect 1609 -1856 1671 -1840
rect 1683 -1856 1689 -1808
rect 1692 -1816 1772 -1808
rect 1692 -1818 1711 -1816
rect 1726 -1818 1760 -1816
rect 1692 -1834 1772 -1818
rect 1692 -1856 1711 -1834
rect 1726 -1850 1756 -1834
rect 1784 -1840 1790 -1766
rect 1793 -1840 1812 -1696
rect 1827 -1840 1833 -1696
rect 1842 -1766 1855 -1696
rect 1907 -1700 1929 -1696
rect 1900 -1712 1917 -1708
rect 1921 -1710 1929 -1708
rect 1919 -1712 1929 -1710
rect 1900 -1722 1929 -1712
rect 1982 -1722 1998 -1708
rect 2036 -1712 2042 -1710
rect 2049 -1712 2157 -1696
rect 2164 -1712 2170 -1710
rect 2178 -1712 2193 -1696
rect 2259 -1702 2278 -1699
rect 1900 -1724 1998 -1722
rect 2025 -1724 2193 -1712
rect 2208 -1722 2224 -1708
rect 2259 -1721 2281 -1702
rect 2291 -1708 2307 -1707
rect 2290 -1710 2307 -1708
rect 2291 -1715 2307 -1710
rect 2281 -1722 2287 -1721
rect 2290 -1722 2319 -1715
rect 2208 -1723 2319 -1722
rect 2208 -1724 2325 -1723
rect 1884 -1732 1935 -1724
rect 1982 -1732 2016 -1724
rect 1884 -1744 1909 -1732
rect 1916 -1744 1935 -1732
rect 1989 -1734 2016 -1732
rect 2025 -1734 2246 -1724
rect 2281 -1727 2287 -1724
rect 1989 -1738 2246 -1734
rect 1884 -1752 1935 -1744
rect 1982 -1752 2246 -1738
rect 2290 -1732 2325 -1724
rect 1836 -1800 1855 -1766
rect 1900 -1760 1929 -1752
rect 1900 -1766 1917 -1760
rect 1900 -1768 1934 -1766
rect 1982 -1768 1998 -1752
rect 1999 -1762 2207 -1752
rect 2208 -1762 2224 -1752
rect 2272 -1756 2287 -1741
rect 2290 -1744 2291 -1732
rect 2298 -1744 2325 -1732
rect 2290 -1752 2325 -1744
rect 2290 -1753 2319 -1752
rect 2010 -1766 2224 -1762
rect 2025 -1768 2224 -1766
rect 2259 -1766 2272 -1756
rect 2290 -1766 2307 -1753
rect 2259 -1768 2307 -1766
rect 1901 -1772 1934 -1768
rect 1897 -1774 1934 -1772
rect 1897 -1775 1964 -1774
rect 1897 -1780 1928 -1775
rect 1934 -1780 1964 -1775
rect 1897 -1784 1964 -1780
rect 1870 -1787 1964 -1784
rect 1870 -1794 1919 -1787
rect 1870 -1800 1900 -1794
rect 1919 -1799 1924 -1794
rect 1836 -1816 1916 -1800
rect 1928 -1808 1964 -1787
rect 2025 -1792 2214 -1768
rect 2259 -1769 2306 -1768
rect 2272 -1774 2306 -1769
rect 2040 -1795 2214 -1792
rect 2033 -1798 2214 -1795
rect 2242 -1775 2306 -1774
rect 1836 -1818 1855 -1816
rect 1870 -1818 1904 -1816
rect 1836 -1834 1916 -1818
rect 1836 -1840 1855 -1834
rect 1552 -1866 1655 -1856
rect 1506 -1868 1655 -1866
rect 1676 -1868 1711 -1856
rect 1345 -1870 1507 -1868
rect 1357 -1888 1376 -1870
rect 1391 -1872 1421 -1870
rect 1240 -1898 1281 -1890
rect 1364 -1894 1376 -1888
rect 1428 -1888 1507 -1870
rect 1539 -1870 1711 -1868
rect 1539 -1886 1618 -1870
rect 1625 -1872 1655 -1870
rect 1514 -1888 1618 -1886
rect 1203 -1908 1232 -1898
rect 1246 -1908 1275 -1898
rect 1290 -1908 1320 -1894
rect 1364 -1908 1406 -1894
rect 1428 -1898 1618 -1888
rect 1683 -1890 1689 -1870
rect 1413 -1908 1443 -1898
rect 1444 -1908 1602 -1898
rect 1606 -1908 1636 -1898
rect 1640 -1908 1670 -1894
rect 1698 -1908 1711 -1870
rect 1783 -1856 1812 -1840
rect 1826 -1856 1855 -1840
rect 1870 -1850 1900 -1834
rect 1928 -1856 1934 -1808
rect 1937 -1814 1956 -1808
rect 1971 -1814 2001 -1806
rect 1937 -1822 2001 -1814
rect 1937 -1838 2017 -1822
rect 2033 -1829 2095 -1798
rect 2111 -1829 2173 -1798
rect 2242 -1800 2291 -1775
rect 2306 -1800 2336 -1782
rect 2205 -1814 2235 -1806
rect 2242 -1808 2352 -1800
rect 2205 -1822 2250 -1814
rect 1937 -1840 1956 -1838
rect 1971 -1840 2017 -1838
rect 1937 -1856 2017 -1840
rect 2044 -1842 2079 -1829
rect 2120 -1832 2157 -1829
rect 2120 -1834 2162 -1832
rect 2049 -1845 2079 -1842
rect 2058 -1849 2065 -1845
rect 2065 -1850 2066 -1849
rect 2024 -1856 2034 -1850
rect 1783 -1864 1818 -1856
rect 1783 -1890 1784 -1864
rect 1791 -1890 1818 -1864
rect 1726 -1908 1756 -1894
rect 1783 -1898 1818 -1890
rect 1820 -1864 1861 -1856
rect 1820 -1890 1835 -1864
rect 1842 -1890 1861 -1864
rect 1925 -1868 1956 -1856
rect 1971 -1868 2074 -1856
rect 2086 -1866 2112 -1840
rect 2127 -1845 2157 -1834
rect 2189 -1838 2251 -1822
rect 2189 -1840 2235 -1838
rect 2189 -1856 2251 -1840
rect 2263 -1856 2269 -1808
rect 2272 -1816 2352 -1808
rect 2272 -1818 2291 -1816
rect 2306 -1818 2340 -1816
rect 2272 -1833 2352 -1818
rect 2272 -1834 2358 -1833
rect 2272 -1856 2291 -1834
rect 2306 -1850 2336 -1834
rect 2364 -1840 2370 -1766
rect 2373 -1840 2392 -1696
rect 2407 -1840 2413 -1696
rect 2422 -1766 2435 -1696
rect 2487 -1700 2509 -1696
rect 2480 -1712 2497 -1708
rect 2501 -1710 2509 -1708
rect 2499 -1712 2509 -1710
rect 2480 -1722 2509 -1712
rect 2562 -1722 2578 -1708
rect 2616 -1712 2622 -1710
rect 2629 -1712 2737 -1696
rect 2744 -1712 2750 -1710
rect 2758 -1712 2773 -1696
rect 2839 -1702 2858 -1699
rect 2480 -1724 2578 -1722
rect 2605 -1724 2773 -1712
rect 2788 -1722 2804 -1708
rect 2839 -1721 2861 -1702
rect 2871 -1708 2887 -1707
rect 2870 -1710 2887 -1708
rect 2871 -1715 2887 -1710
rect 2861 -1722 2867 -1721
rect 2870 -1722 2899 -1715
rect 2788 -1723 2899 -1722
rect 2788 -1724 2905 -1723
rect 2464 -1732 2515 -1724
rect 2562 -1732 2596 -1724
rect 2464 -1744 2489 -1732
rect 2496 -1744 2515 -1732
rect 2569 -1734 2596 -1732
rect 2605 -1734 2826 -1724
rect 2861 -1727 2867 -1724
rect 2569 -1738 2826 -1734
rect 2464 -1752 2515 -1744
rect 2562 -1752 2826 -1738
rect 2870 -1732 2905 -1724
rect 2416 -1800 2435 -1766
rect 2480 -1760 2509 -1752
rect 2480 -1766 2497 -1760
rect 2480 -1768 2514 -1766
rect 2562 -1768 2578 -1752
rect 2579 -1762 2787 -1752
rect 2788 -1762 2804 -1752
rect 2852 -1756 2867 -1741
rect 2870 -1744 2871 -1732
rect 2878 -1744 2905 -1732
rect 2870 -1752 2905 -1744
rect 2870 -1753 2899 -1752
rect 2590 -1766 2804 -1762
rect 2605 -1768 2804 -1766
rect 2839 -1766 2852 -1756
rect 2870 -1766 2887 -1753
rect 2839 -1768 2887 -1766
rect 2481 -1772 2514 -1768
rect 2477 -1774 2514 -1772
rect 2477 -1775 2544 -1774
rect 2477 -1780 2508 -1775
rect 2514 -1780 2544 -1775
rect 2477 -1784 2544 -1780
rect 2450 -1787 2544 -1784
rect 2450 -1794 2499 -1787
rect 2450 -1800 2480 -1794
rect 2499 -1799 2504 -1794
rect 2416 -1816 2496 -1800
rect 2508 -1808 2544 -1787
rect 2605 -1792 2794 -1768
rect 2839 -1769 2886 -1768
rect 2852 -1774 2886 -1769
rect 2926 -1774 2942 -1772
rect 2620 -1795 2794 -1792
rect 2613 -1798 2794 -1795
rect 2822 -1775 2886 -1774
rect 2416 -1818 2435 -1816
rect 2450 -1818 2484 -1816
rect 2416 -1834 2496 -1818
rect 2416 -1840 2435 -1834
rect 2132 -1866 2235 -1856
rect 2086 -1868 2235 -1866
rect 2256 -1868 2291 -1856
rect 1925 -1870 2087 -1868
rect 1937 -1888 1956 -1870
rect 1971 -1872 2001 -1870
rect 1820 -1898 1861 -1890
rect 1944 -1894 1956 -1888
rect 2008 -1886 2087 -1870
rect 2119 -1870 2291 -1868
rect 2119 -1886 2198 -1870
rect 2205 -1872 2235 -1870
rect 1783 -1908 1812 -1898
rect 1826 -1908 1855 -1898
rect 1870 -1908 1900 -1894
rect 1944 -1908 1986 -1894
rect 2008 -1898 2198 -1886
rect 2263 -1890 2269 -1870
rect 1993 -1908 2023 -1898
rect 2024 -1908 2182 -1898
rect 2186 -1908 2216 -1898
rect 2220 -1908 2250 -1894
rect 2278 -1908 2291 -1870
rect 2363 -1856 2392 -1840
rect 2406 -1856 2435 -1840
rect 2450 -1850 2480 -1834
rect 2508 -1856 2514 -1808
rect 2517 -1814 2536 -1808
rect 2551 -1814 2581 -1806
rect 2517 -1822 2581 -1814
rect 2517 -1838 2597 -1822
rect 2613 -1829 2675 -1798
rect 2691 -1829 2753 -1798
rect 2822 -1800 2871 -1775
rect 2916 -1784 2942 -1774
rect 2886 -1800 2942 -1784
rect 2785 -1814 2815 -1806
rect 2822 -1808 2932 -1800
rect 2785 -1822 2830 -1814
rect 2517 -1840 2536 -1838
rect 2551 -1840 2597 -1838
rect 2517 -1856 2597 -1840
rect 2624 -1842 2659 -1829
rect 2700 -1832 2737 -1829
rect 2700 -1834 2742 -1832
rect 2629 -1845 2659 -1842
rect 2638 -1849 2645 -1845
rect 2645 -1850 2646 -1849
rect 2604 -1856 2614 -1850
rect 2363 -1864 2398 -1856
rect 2363 -1890 2364 -1864
rect 2371 -1890 2398 -1864
rect 2306 -1908 2336 -1894
rect 2363 -1898 2398 -1890
rect 2400 -1864 2441 -1856
rect 2400 -1890 2415 -1864
rect 2422 -1890 2441 -1864
rect 2505 -1868 2536 -1856
rect 2551 -1868 2654 -1856
rect 2666 -1866 2692 -1840
rect 2707 -1845 2737 -1834
rect 2769 -1838 2831 -1822
rect 2769 -1840 2815 -1838
rect 2769 -1856 2831 -1840
rect 2843 -1856 2849 -1808
rect 2852 -1816 2932 -1808
rect 2852 -1818 2871 -1816
rect 2886 -1818 2920 -1816
rect 2852 -1834 2932 -1818
rect 2852 -1856 2871 -1834
rect 2886 -1850 2916 -1834
rect 2944 -1840 2950 -1766
rect 2953 -1840 2972 -1696
rect 2987 -1840 2993 -1696
rect 3002 -1766 3015 -1696
rect 3067 -1700 3089 -1696
rect 3060 -1712 3077 -1708
rect 3081 -1710 3089 -1708
rect 3079 -1712 3089 -1710
rect 3060 -1722 3089 -1712
rect 3142 -1722 3158 -1708
rect 3196 -1712 3202 -1710
rect 3209 -1712 3317 -1696
rect 3324 -1712 3330 -1710
rect 3338 -1712 3353 -1696
rect 3419 -1702 3438 -1699
rect 3060 -1724 3158 -1722
rect 3185 -1724 3353 -1712
rect 3368 -1722 3384 -1708
rect 3419 -1721 3441 -1702
rect 3451 -1708 3467 -1707
rect 3450 -1710 3467 -1708
rect 3451 -1715 3467 -1710
rect 3441 -1722 3447 -1721
rect 3450 -1722 3479 -1715
rect 3368 -1723 3479 -1722
rect 3368 -1724 3485 -1723
rect 3044 -1732 3095 -1724
rect 3142 -1732 3176 -1724
rect 3044 -1744 3069 -1732
rect 3076 -1744 3095 -1732
rect 3149 -1734 3176 -1732
rect 3185 -1734 3406 -1724
rect 3441 -1727 3447 -1724
rect 3149 -1738 3406 -1734
rect 3044 -1752 3095 -1744
rect 3142 -1752 3406 -1738
rect 3450 -1732 3485 -1724
rect 2996 -1800 3015 -1766
rect 3060 -1760 3089 -1752
rect 3060 -1766 3077 -1760
rect 3060 -1768 3094 -1766
rect 3142 -1768 3158 -1752
rect 3159 -1762 3367 -1752
rect 3368 -1762 3384 -1752
rect 3432 -1756 3447 -1741
rect 3450 -1744 3451 -1732
rect 3458 -1744 3485 -1732
rect 3450 -1752 3485 -1744
rect 3450 -1753 3479 -1752
rect 3170 -1766 3384 -1762
rect 3185 -1768 3384 -1766
rect 3419 -1766 3432 -1756
rect 3450 -1766 3467 -1753
rect 3419 -1768 3467 -1766
rect 3061 -1772 3094 -1768
rect 3057 -1774 3094 -1772
rect 3057 -1775 3124 -1774
rect 3057 -1780 3088 -1775
rect 3094 -1780 3124 -1775
rect 3057 -1784 3124 -1780
rect 3030 -1787 3124 -1784
rect 3030 -1794 3079 -1787
rect 3030 -1800 3060 -1794
rect 3079 -1799 3084 -1794
rect 2996 -1816 3076 -1800
rect 3088 -1808 3124 -1787
rect 3185 -1792 3374 -1768
rect 3419 -1769 3466 -1768
rect 3432 -1774 3466 -1769
rect 3200 -1795 3374 -1792
rect 3193 -1798 3374 -1795
rect 3402 -1775 3466 -1774
rect 2996 -1818 3015 -1816
rect 3030 -1818 3064 -1816
rect 2996 -1834 3076 -1818
rect 2996 -1840 3015 -1834
rect 2712 -1866 2815 -1856
rect 2666 -1868 2815 -1866
rect 2836 -1868 2871 -1856
rect 2505 -1870 2667 -1868
rect 2517 -1888 2536 -1870
rect 2551 -1872 2581 -1870
rect 2400 -1898 2441 -1890
rect 2524 -1894 2536 -1888
rect 2588 -1886 2667 -1870
rect 2699 -1870 2871 -1868
rect 2699 -1886 2778 -1870
rect 2785 -1872 2815 -1870
rect 2363 -1908 2392 -1898
rect 2406 -1908 2435 -1898
rect 2450 -1908 2480 -1894
rect 2524 -1908 2566 -1894
rect 2588 -1898 2778 -1886
rect 2843 -1890 2849 -1870
rect 2573 -1908 2603 -1898
rect 2604 -1908 2762 -1898
rect 2766 -1908 2796 -1898
rect 2800 -1908 2830 -1894
rect 2858 -1908 2871 -1870
rect 2943 -1856 2972 -1840
rect 2986 -1856 3015 -1840
rect 3030 -1850 3060 -1834
rect 3088 -1856 3094 -1808
rect 3097 -1814 3116 -1808
rect 3131 -1814 3161 -1806
rect 3097 -1822 3161 -1814
rect 3097 -1838 3177 -1822
rect 3193 -1829 3255 -1798
rect 3271 -1829 3333 -1798
rect 3402 -1800 3451 -1775
rect 3466 -1800 3496 -1782
rect 3365 -1814 3395 -1806
rect 3402 -1808 3512 -1800
rect 3365 -1822 3410 -1814
rect 3097 -1840 3116 -1838
rect 3131 -1840 3177 -1838
rect 3097 -1856 3177 -1840
rect 3204 -1842 3239 -1829
rect 3280 -1832 3317 -1829
rect 3280 -1834 3322 -1832
rect 3209 -1845 3239 -1842
rect 3218 -1849 3225 -1845
rect 3225 -1850 3226 -1849
rect 3184 -1856 3194 -1850
rect 2943 -1864 2978 -1856
rect 2943 -1890 2944 -1864
rect 2951 -1890 2978 -1864
rect 2886 -1908 2916 -1894
rect 2943 -1898 2978 -1890
rect 2980 -1864 3021 -1856
rect 2980 -1890 2995 -1864
rect 3002 -1890 3021 -1864
rect 3085 -1868 3116 -1856
rect 3131 -1868 3234 -1856
rect 3246 -1866 3272 -1840
rect 3287 -1845 3317 -1834
rect 3349 -1838 3411 -1822
rect 3349 -1840 3395 -1838
rect 3349 -1856 3411 -1840
rect 3423 -1856 3429 -1808
rect 3432 -1816 3512 -1808
rect 3432 -1818 3451 -1816
rect 3466 -1818 3500 -1816
rect 3432 -1833 3512 -1818
rect 3432 -1834 3518 -1833
rect 3432 -1856 3451 -1834
rect 3466 -1850 3496 -1834
rect 3524 -1840 3530 -1766
rect 3533 -1840 3552 -1696
rect 3567 -1840 3573 -1696
rect 3582 -1766 3595 -1696
rect 3647 -1700 3669 -1696
rect 3640 -1712 3657 -1708
rect 3661 -1710 3669 -1708
rect 3659 -1712 3669 -1710
rect 3640 -1722 3669 -1712
rect 3722 -1722 3738 -1708
rect 3776 -1712 3782 -1710
rect 3789 -1712 3897 -1696
rect 3904 -1712 3910 -1710
rect 3918 -1712 3933 -1696
rect 3999 -1702 4018 -1699
rect 3640 -1724 3738 -1722
rect 3765 -1724 3933 -1712
rect 3948 -1722 3964 -1708
rect 3999 -1721 4021 -1702
rect 4031 -1708 4047 -1707
rect 4030 -1710 4047 -1708
rect 4031 -1715 4047 -1710
rect 4021 -1722 4027 -1721
rect 4030 -1722 4059 -1715
rect 3948 -1723 4059 -1722
rect 3948 -1724 4065 -1723
rect 3624 -1732 3675 -1724
rect 3722 -1732 3756 -1724
rect 3624 -1744 3649 -1732
rect 3656 -1744 3675 -1732
rect 3729 -1734 3756 -1732
rect 3765 -1734 3986 -1724
rect 4021 -1727 4027 -1724
rect 3729 -1738 3986 -1734
rect 3624 -1752 3675 -1744
rect 3722 -1752 3986 -1738
rect 4030 -1732 4065 -1724
rect 3576 -1800 3595 -1766
rect 3640 -1760 3669 -1752
rect 3640 -1766 3657 -1760
rect 3640 -1768 3674 -1766
rect 3722 -1768 3738 -1752
rect 3739 -1762 3947 -1752
rect 3948 -1762 3964 -1752
rect 4012 -1756 4027 -1741
rect 4030 -1744 4031 -1732
rect 4038 -1744 4065 -1732
rect 4030 -1752 4065 -1744
rect 4030 -1753 4059 -1752
rect 3750 -1766 3964 -1762
rect 3765 -1768 3964 -1766
rect 3999 -1766 4012 -1756
rect 4030 -1766 4047 -1753
rect 3999 -1768 4047 -1766
rect 3641 -1772 3674 -1768
rect 3637 -1774 3674 -1772
rect 3637 -1775 3704 -1774
rect 3637 -1780 3668 -1775
rect 3674 -1780 3704 -1775
rect 3637 -1784 3704 -1780
rect 3610 -1787 3704 -1784
rect 3610 -1794 3659 -1787
rect 3610 -1800 3640 -1794
rect 3659 -1799 3664 -1794
rect 3576 -1816 3656 -1800
rect 3668 -1808 3704 -1787
rect 3765 -1792 3954 -1768
rect 3999 -1769 4046 -1768
rect 4012 -1774 4046 -1769
rect 4086 -1774 4102 -1772
rect 3780 -1795 3954 -1792
rect 3773 -1798 3954 -1795
rect 3982 -1775 4046 -1774
rect 3576 -1818 3595 -1816
rect 3610 -1818 3644 -1816
rect 3576 -1834 3656 -1818
rect 3576 -1840 3595 -1834
rect 3292 -1866 3395 -1856
rect 3246 -1868 3395 -1866
rect 3416 -1868 3451 -1856
rect 3085 -1870 3247 -1868
rect 3097 -1888 3116 -1870
rect 3131 -1872 3161 -1870
rect 2980 -1898 3021 -1890
rect 3104 -1894 3116 -1888
rect 3168 -1886 3247 -1870
rect 3279 -1870 3451 -1868
rect 3279 -1886 3358 -1870
rect 3365 -1872 3395 -1870
rect 2943 -1908 2972 -1898
rect 2986 -1908 3015 -1898
rect 3030 -1908 3060 -1894
rect 3104 -1908 3146 -1894
rect 3168 -1898 3358 -1886
rect 3423 -1890 3429 -1870
rect 3153 -1908 3183 -1898
rect 3184 -1908 3342 -1898
rect 3346 -1908 3376 -1898
rect 3380 -1908 3410 -1894
rect 3438 -1908 3451 -1870
rect 3523 -1856 3552 -1840
rect 3566 -1856 3595 -1840
rect 3610 -1850 3640 -1834
rect 3668 -1856 3674 -1808
rect 3677 -1814 3696 -1808
rect 3711 -1814 3741 -1806
rect 3677 -1822 3741 -1814
rect 3677 -1838 3757 -1822
rect 3773 -1829 3835 -1798
rect 3851 -1829 3913 -1798
rect 3982 -1800 4031 -1775
rect 4076 -1784 4102 -1774
rect 4046 -1800 4102 -1784
rect 3945 -1814 3975 -1806
rect 3982 -1808 4092 -1800
rect 3945 -1822 3990 -1814
rect 3677 -1840 3696 -1838
rect 3711 -1840 3757 -1838
rect 3677 -1856 3757 -1840
rect 3784 -1842 3819 -1829
rect 3860 -1832 3897 -1829
rect 3860 -1834 3902 -1832
rect 3789 -1845 3819 -1842
rect 3798 -1849 3805 -1845
rect 3805 -1850 3806 -1849
rect 3764 -1856 3774 -1850
rect 3523 -1864 3558 -1856
rect 3523 -1890 3524 -1864
rect 3531 -1890 3558 -1864
rect 3466 -1908 3496 -1894
rect 3523 -1898 3558 -1890
rect 3560 -1864 3601 -1856
rect 3560 -1890 3575 -1864
rect 3582 -1890 3601 -1864
rect 3665 -1868 3696 -1856
rect 3711 -1868 3814 -1856
rect 3826 -1866 3852 -1840
rect 3867 -1845 3897 -1834
rect 3929 -1838 3991 -1822
rect 3929 -1840 3975 -1838
rect 3929 -1856 3991 -1840
rect 4003 -1856 4009 -1808
rect 4012 -1816 4092 -1808
rect 4012 -1818 4031 -1816
rect 4046 -1818 4080 -1816
rect 4012 -1834 4092 -1818
rect 4012 -1856 4031 -1834
rect 4046 -1850 4076 -1834
rect 4104 -1840 4110 -1766
rect 4113 -1840 4132 -1696
rect 4147 -1840 4153 -1696
rect 4162 -1766 4175 -1696
rect 4227 -1700 4249 -1696
rect 4220 -1712 4237 -1708
rect 4241 -1710 4249 -1708
rect 4239 -1712 4249 -1710
rect 4220 -1722 4249 -1712
rect 4302 -1722 4318 -1708
rect 4356 -1712 4362 -1710
rect 4369 -1712 4477 -1696
rect 4484 -1712 4490 -1710
rect 4498 -1712 4513 -1696
rect 4579 -1702 4598 -1699
rect 4220 -1724 4318 -1722
rect 4345 -1724 4513 -1712
rect 4528 -1722 4544 -1708
rect 4579 -1721 4601 -1702
rect 4611 -1708 4627 -1707
rect 4610 -1710 4627 -1708
rect 4611 -1715 4627 -1710
rect 4601 -1722 4607 -1721
rect 4610 -1722 4639 -1715
rect 4528 -1723 4639 -1722
rect 4528 -1724 4645 -1723
rect 4204 -1732 4255 -1724
rect 4302 -1732 4336 -1724
rect 4204 -1744 4229 -1732
rect 4236 -1744 4255 -1732
rect 4309 -1734 4336 -1732
rect 4345 -1734 4566 -1724
rect 4601 -1727 4607 -1724
rect 4309 -1738 4566 -1734
rect 4204 -1752 4255 -1744
rect 4302 -1752 4566 -1738
rect 4610 -1732 4645 -1724
rect 4156 -1800 4175 -1766
rect 4220 -1760 4249 -1752
rect 4220 -1766 4237 -1760
rect 4220 -1768 4254 -1766
rect 4302 -1768 4318 -1752
rect 4319 -1762 4527 -1752
rect 4528 -1762 4544 -1752
rect 4592 -1756 4607 -1741
rect 4610 -1744 4611 -1732
rect 4618 -1744 4645 -1732
rect 4610 -1752 4645 -1744
rect 4610 -1753 4639 -1752
rect 4330 -1766 4544 -1762
rect 4345 -1768 4544 -1766
rect 4579 -1766 4592 -1756
rect 4610 -1766 4627 -1753
rect 4579 -1768 4627 -1766
rect 4221 -1772 4254 -1768
rect 4217 -1774 4254 -1772
rect 4217 -1775 4284 -1774
rect 4217 -1780 4248 -1775
rect 4254 -1780 4284 -1775
rect 4217 -1784 4284 -1780
rect 4190 -1787 4284 -1784
rect 4190 -1794 4239 -1787
rect 4190 -1800 4220 -1794
rect 4239 -1799 4244 -1794
rect 4156 -1816 4236 -1800
rect 4248 -1808 4284 -1787
rect 4345 -1792 4534 -1768
rect 4579 -1769 4626 -1768
rect 4592 -1774 4626 -1769
rect 4360 -1795 4534 -1792
rect 4353 -1798 4534 -1795
rect 4562 -1775 4626 -1774
rect 4156 -1818 4175 -1816
rect 4190 -1818 4224 -1816
rect 4156 -1834 4236 -1818
rect 4156 -1840 4175 -1834
rect 3872 -1866 3975 -1856
rect 3826 -1868 3975 -1866
rect 3996 -1868 4031 -1856
rect 3665 -1870 3827 -1868
rect 3677 -1888 3696 -1870
rect 3711 -1872 3741 -1870
rect 3560 -1898 3601 -1890
rect 3684 -1894 3696 -1888
rect 3748 -1886 3827 -1870
rect 3859 -1870 4031 -1868
rect 3859 -1886 3938 -1870
rect 3945 -1872 3975 -1870
rect 3523 -1908 3552 -1898
rect 3566 -1908 3595 -1898
rect 3610 -1908 3640 -1894
rect 3684 -1908 3726 -1894
rect 3748 -1898 3938 -1886
rect 4003 -1890 4009 -1870
rect 3733 -1908 3763 -1898
rect 3764 -1908 3922 -1898
rect 3926 -1908 3956 -1898
rect 3960 -1908 3990 -1894
rect 4018 -1908 4031 -1870
rect 4103 -1856 4132 -1840
rect 4146 -1856 4175 -1840
rect 4190 -1850 4220 -1834
rect 4248 -1856 4254 -1808
rect 4257 -1814 4276 -1808
rect 4291 -1814 4321 -1806
rect 4257 -1822 4321 -1814
rect 4257 -1838 4337 -1822
rect 4353 -1829 4415 -1798
rect 4431 -1829 4493 -1798
rect 4562 -1800 4611 -1775
rect 4626 -1800 4656 -1782
rect 4525 -1814 4555 -1806
rect 4562 -1808 4672 -1800
rect 4525 -1822 4570 -1814
rect 4257 -1840 4276 -1838
rect 4291 -1840 4337 -1838
rect 4257 -1856 4337 -1840
rect 4364 -1842 4399 -1829
rect 4440 -1832 4477 -1829
rect 4440 -1834 4482 -1832
rect 4369 -1845 4399 -1842
rect 4378 -1849 4385 -1845
rect 4385 -1850 4386 -1849
rect 4344 -1856 4354 -1850
rect 4103 -1864 4138 -1856
rect 4103 -1890 4104 -1864
rect 4111 -1890 4138 -1864
rect 4046 -1908 4076 -1894
rect 4103 -1898 4138 -1890
rect 4140 -1864 4181 -1856
rect 4140 -1890 4155 -1864
rect 4162 -1890 4181 -1864
rect 4245 -1868 4276 -1856
rect 4291 -1868 4394 -1856
rect 4406 -1866 4432 -1840
rect 4447 -1845 4477 -1834
rect 4509 -1838 4571 -1822
rect 4509 -1840 4555 -1838
rect 4509 -1856 4571 -1840
rect 4583 -1856 4589 -1808
rect 4592 -1816 4672 -1808
rect 4592 -1818 4611 -1816
rect 4626 -1818 4660 -1816
rect 4592 -1833 4672 -1818
rect 4592 -1834 4678 -1833
rect 4592 -1856 4611 -1834
rect 4626 -1850 4656 -1834
rect 4684 -1840 4690 -1766
rect 4693 -1840 4712 -1696
rect 4727 -1840 4733 -1696
rect 4742 -1766 4755 -1696
rect 4807 -1700 4829 -1696
rect 4800 -1712 4817 -1708
rect 4821 -1710 4829 -1708
rect 4819 -1712 4829 -1710
rect 4800 -1722 4829 -1712
rect 4882 -1722 4898 -1708
rect 4936 -1712 4942 -1710
rect 4949 -1712 5057 -1696
rect 5064 -1712 5070 -1710
rect 5078 -1712 5093 -1696
rect 5159 -1702 5178 -1699
rect 4800 -1724 4898 -1722
rect 4925 -1724 5093 -1712
rect 5108 -1722 5124 -1708
rect 5159 -1721 5181 -1702
rect 5191 -1708 5207 -1707
rect 5190 -1710 5207 -1708
rect 5191 -1715 5207 -1710
rect 5181 -1722 5187 -1721
rect 5190 -1722 5219 -1715
rect 5108 -1723 5219 -1722
rect 5108 -1724 5225 -1723
rect 4784 -1732 4835 -1724
rect 4882 -1732 4916 -1724
rect 4784 -1744 4809 -1732
rect 4816 -1744 4835 -1732
rect 4889 -1734 4916 -1732
rect 4925 -1734 5146 -1724
rect 5181 -1727 5187 -1724
rect 4889 -1738 5146 -1734
rect 4784 -1752 4835 -1744
rect 4882 -1752 5146 -1738
rect 5190 -1732 5225 -1724
rect 4736 -1800 4755 -1766
rect 4800 -1760 4829 -1752
rect 4800 -1766 4817 -1760
rect 4800 -1768 4834 -1766
rect 4882 -1768 4898 -1752
rect 4899 -1762 5107 -1752
rect 5108 -1762 5124 -1752
rect 5172 -1756 5187 -1741
rect 5190 -1744 5191 -1732
rect 5198 -1744 5225 -1732
rect 5190 -1752 5225 -1744
rect 5190 -1753 5219 -1752
rect 4910 -1766 5124 -1762
rect 4925 -1768 5124 -1766
rect 5159 -1766 5172 -1756
rect 5190 -1766 5207 -1753
rect 5159 -1768 5207 -1766
rect 4801 -1772 4834 -1768
rect 4797 -1774 4834 -1772
rect 4797 -1775 4864 -1774
rect 4797 -1780 4828 -1775
rect 4834 -1780 4864 -1775
rect 4797 -1784 4864 -1780
rect 4770 -1787 4864 -1784
rect 4770 -1794 4819 -1787
rect 4770 -1800 4800 -1794
rect 4819 -1799 4824 -1794
rect 4736 -1816 4816 -1800
rect 4828 -1808 4864 -1787
rect 4925 -1792 5114 -1768
rect 5159 -1769 5206 -1768
rect 5172 -1774 5206 -1769
rect 5246 -1774 5262 -1772
rect 4940 -1795 5114 -1792
rect 4933 -1798 5114 -1795
rect 5142 -1775 5206 -1774
rect 4736 -1818 4755 -1816
rect 4770 -1818 4804 -1816
rect 4736 -1834 4816 -1818
rect 4736 -1840 4755 -1834
rect 4452 -1866 4555 -1856
rect 4406 -1868 4555 -1866
rect 4576 -1868 4611 -1856
rect 4245 -1870 4407 -1868
rect 4257 -1888 4276 -1870
rect 4291 -1872 4321 -1870
rect 4140 -1898 4181 -1890
rect 4264 -1894 4276 -1888
rect 4328 -1886 4407 -1870
rect 4439 -1870 4611 -1868
rect 4439 -1886 4518 -1870
rect 4525 -1872 4555 -1870
rect 4103 -1908 4132 -1898
rect 4146 -1908 4175 -1898
rect 4190 -1908 4220 -1894
rect 4264 -1908 4306 -1894
rect 4328 -1898 4518 -1886
rect 4583 -1890 4589 -1870
rect 4313 -1908 4343 -1898
rect 4344 -1908 4502 -1898
rect 4506 -1908 4536 -1898
rect 4540 -1908 4570 -1894
rect 4598 -1908 4611 -1870
rect 4683 -1856 4712 -1840
rect 4726 -1856 4755 -1840
rect 4770 -1850 4800 -1834
rect 4828 -1856 4834 -1808
rect 4837 -1814 4856 -1808
rect 4871 -1814 4901 -1806
rect 4837 -1822 4901 -1814
rect 4837 -1838 4917 -1822
rect 4933 -1829 4995 -1798
rect 5011 -1829 5073 -1798
rect 5142 -1800 5191 -1775
rect 5236 -1784 5262 -1774
rect 5206 -1800 5262 -1784
rect 5105 -1814 5135 -1806
rect 5142 -1808 5252 -1800
rect 5105 -1822 5150 -1814
rect 4837 -1840 4856 -1838
rect 4871 -1840 4917 -1838
rect 4837 -1856 4917 -1840
rect 4944 -1842 4979 -1829
rect 5020 -1832 5057 -1829
rect 5020 -1834 5062 -1832
rect 4949 -1845 4979 -1842
rect 4958 -1849 4965 -1845
rect 4965 -1850 4966 -1849
rect 4924 -1856 4934 -1850
rect 4683 -1864 4718 -1856
rect 4683 -1890 4684 -1864
rect 4691 -1890 4718 -1864
rect 4626 -1908 4656 -1894
rect 4683 -1898 4718 -1890
rect 4720 -1864 4761 -1856
rect 4720 -1890 4735 -1864
rect 4742 -1890 4761 -1864
rect 4825 -1868 4856 -1856
rect 4871 -1868 4974 -1856
rect 4986 -1866 5012 -1840
rect 5027 -1845 5057 -1834
rect 5089 -1838 5151 -1822
rect 5089 -1840 5135 -1838
rect 5089 -1856 5151 -1840
rect 5163 -1856 5169 -1808
rect 5172 -1816 5252 -1808
rect 5172 -1818 5191 -1816
rect 5206 -1818 5240 -1816
rect 5172 -1834 5252 -1818
rect 5172 -1856 5191 -1834
rect 5206 -1850 5236 -1834
rect 5264 -1840 5270 -1766
rect 5273 -1840 5292 -1696
rect 5307 -1840 5313 -1696
rect 5322 -1766 5335 -1696
rect 5387 -1700 5409 -1696
rect 5380 -1712 5397 -1708
rect 5401 -1710 5409 -1708
rect 5399 -1712 5409 -1710
rect 5380 -1722 5409 -1712
rect 5462 -1722 5478 -1708
rect 5516 -1712 5522 -1710
rect 5529 -1712 5637 -1696
rect 5644 -1712 5650 -1710
rect 5658 -1712 5673 -1696
rect 5739 -1702 5758 -1699
rect 5380 -1724 5478 -1722
rect 5505 -1724 5673 -1712
rect 5688 -1722 5704 -1708
rect 5739 -1721 5761 -1702
rect 5771 -1708 5787 -1707
rect 5770 -1710 5787 -1708
rect 5771 -1715 5787 -1710
rect 5761 -1722 5767 -1721
rect 5770 -1722 5799 -1715
rect 5688 -1723 5799 -1722
rect 5688 -1724 5805 -1723
rect 5364 -1732 5415 -1724
rect 5462 -1732 5496 -1724
rect 5364 -1744 5389 -1732
rect 5396 -1744 5415 -1732
rect 5469 -1734 5496 -1732
rect 5505 -1734 5726 -1724
rect 5761 -1727 5767 -1724
rect 5469 -1738 5726 -1734
rect 5364 -1752 5415 -1744
rect 5462 -1752 5726 -1738
rect 5770 -1732 5805 -1724
rect 5316 -1800 5335 -1766
rect 5380 -1760 5409 -1752
rect 5380 -1766 5397 -1760
rect 5380 -1768 5414 -1766
rect 5462 -1768 5478 -1752
rect 5479 -1762 5687 -1752
rect 5688 -1762 5704 -1752
rect 5752 -1756 5767 -1741
rect 5770 -1744 5771 -1732
rect 5778 -1744 5805 -1732
rect 5770 -1752 5805 -1744
rect 5770 -1753 5799 -1752
rect 5490 -1766 5704 -1762
rect 5505 -1768 5704 -1766
rect 5739 -1766 5752 -1756
rect 5770 -1766 5787 -1753
rect 5739 -1768 5787 -1766
rect 5381 -1772 5414 -1768
rect 5377 -1774 5414 -1772
rect 5377 -1775 5444 -1774
rect 5377 -1780 5408 -1775
rect 5414 -1780 5444 -1775
rect 5377 -1784 5444 -1780
rect 5350 -1787 5444 -1784
rect 5350 -1794 5399 -1787
rect 5350 -1800 5380 -1794
rect 5399 -1799 5404 -1794
rect 5316 -1816 5396 -1800
rect 5408 -1808 5444 -1787
rect 5505 -1792 5694 -1768
rect 5739 -1769 5786 -1768
rect 5752 -1774 5786 -1769
rect 5520 -1795 5694 -1792
rect 5513 -1798 5694 -1795
rect 5722 -1775 5786 -1774
rect 5316 -1818 5335 -1816
rect 5350 -1818 5384 -1816
rect 5316 -1834 5396 -1818
rect 5316 -1840 5335 -1834
rect 5032 -1866 5135 -1856
rect 4986 -1868 5135 -1866
rect 5156 -1868 5191 -1856
rect 4825 -1870 4987 -1868
rect 4837 -1888 4856 -1870
rect 4871 -1872 4901 -1870
rect 4720 -1898 4761 -1890
rect 4844 -1894 4856 -1888
rect 4908 -1886 4987 -1870
rect 5019 -1870 5191 -1868
rect 5019 -1886 5098 -1870
rect 5105 -1872 5135 -1870
rect 4683 -1908 4712 -1898
rect 4726 -1908 4755 -1898
rect 4770 -1908 4800 -1894
rect 4844 -1908 4886 -1894
rect 4908 -1898 5098 -1886
rect 5163 -1890 5169 -1870
rect 4893 -1908 4923 -1898
rect 4924 -1908 5082 -1898
rect 5086 -1908 5116 -1898
rect 5120 -1908 5150 -1894
rect 5178 -1908 5191 -1870
rect 5263 -1856 5292 -1840
rect 5306 -1856 5335 -1840
rect 5350 -1850 5380 -1834
rect 5408 -1856 5414 -1808
rect 5417 -1814 5436 -1808
rect 5451 -1814 5481 -1806
rect 5417 -1822 5481 -1814
rect 5417 -1838 5497 -1822
rect 5513 -1829 5575 -1798
rect 5591 -1829 5653 -1798
rect 5722 -1800 5771 -1775
rect 5786 -1800 5816 -1782
rect 5685 -1814 5715 -1806
rect 5722 -1808 5832 -1800
rect 5685 -1822 5730 -1814
rect 5417 -1840 5436 -1838
rect 5451 -1840 5497 -1838
rect 5417 -1856 5497 -1840
rect 5524 -1842 5559 -1829
rect 5600 -1832 5637 -1829
rect 5600 -1834 5642 -1832
rect 5529 -1845 5559 -1842
rect 5538 -1849 5545 -1845
rect 5545 -1850 5546 -1849
rect 5504 -1856 5514 -1850
rect 5263 -1864 5298 -1856
rect 5263 -1890 5264 -1864
rect 5271 -1890 5298 -1864
rect 5206 -1908 5236 -1894
rect 5263 -1898 5298 -1890
rect 5300 -1864 5341 -1856
rect 5300 -1890 5315 -1864
rect 5322 -1890 5341 -1864
rect 5405 -1868 5436 -1856
rect 5451 -1868 5554 -1856
rect 5566 -1866 5592 -1840
rect 5607 -1845 5637 -1834
rect 5669 -1838 5731 -1822
rect 5669 -1840 5715 -1838
rect 5669 -1856 5731 -1840
rect 5743 -1856 5749 -1808
rect 5752 -1816 5832 -1808
rect 5752 -1818 5771 -1816
rect 5786 -1818 5820 -1816
rect 5752 -1833 5832 -1818
rect 5752 -1834 5838 -1833
rect 5752 -1856 5771 -1834
rect 5786 -1850 5816 -1834
rect 5844 -1840 5850 -1766
rect 5853 -1840 5872 -1696
rect 5887 -1840 5893 -1696
rect 5902 -1766 5915 -1696
rect 5967 -1700 5989 -1696
rect 5960 -1712 5977 -1708
rect 5981 -1710 5989 -1708
rect 5979 -1712 5989 -1710
rect 5960 -1722 5989 -1712
rect 6042 -1722 6058 -1708
rect 6096 -1712 6102 -1710
rect 6109 -1712 6217 -1696
rect 6224 -1712 6230 -1710
rect 6238 -1712 6253 -1696
rect 6319 -1702 6338 -1699
rect 5960 -1724 6058 -1722
rect 6085 -1724 6253 -1712
rect 6268 -1722 6284 -1708
rect 6319 -1721 6341 -1702
rect 6351 -1708 6367 -1707
rect 6350 -1710 6367 -1708
rect 6351 -1715 6367 -1710
rect 6341 -1722 6347 -1721
rect 6350 -1722 6379 -1715
rect 6268 -1723 6379 -1722
rect 6268 -1724 6385 -1723
rect 5944 -1732 5995 -1724
rect 6042 -1732 6076 -1724
rect 5944 -1744 5969 -1732
rect 5976 -1744 5995 -1732
rect 6049 -1734 6076 -1732
rect 6085 -1734 6306 -1724
rect 6341 -1727 6347 -1724
rect 6049 -1738 6306 -1734
rect 5944 -1752 5995 -1744
rect 6042 -1752 6306 -1738
rect 6350 -1732 6385 -1724
rect 5896 -1800 5915 -1766
rect 5960 -1760 5989 -1752
rect 5960 -1766 5977 -1760
rect 5960 -1768 5994 -1766
rect 6042 -1768 6058 -1752
rect 6059 -1762 6267 -1752
rect 6268 -1762 6284 -1752
rect 6332 -1756 6347 -1741
rect 6350 -1744 6351 -1732
rect 6358 -1744 6385 -1732
rect 6350 -1752 6385 -1744
rect 6350 -1753 6379 -1752
rect 6070 -1766 6284 -1762
rect 6085 -1768 6284 -1766
rect 6319 -1766 6332 -1756
rect 6350 -1766 6367 -1753
rect 6319 -1768 6367 -1766
rect 5961 -1772 5994 -1768
rect 5957 -1774 5994 -1772
rect 5957 -1775 6024 -1774
rect 5957 -1780 5988 -1775
rect 5994 -1780 6024 -1775
rect 5957 -1784 6024 -1780
rect 5930 -1787 6024 -1784
rect 5930 -1794 5979 -1787
rect 5930 -1800 5960 -1794
rect 5979 -1799 5984 -1794
rect 5896 -1816 5976 -1800
rect 5988 -1808 6024 -1787
rect 6085 -1792 6274 -1768
rect 6319 -1769 6366 -1768
rect 6332 -1774 6366 -1769
rect 6100 -1795 6274 -1792
rect 6093 -1798 6274 -1795
rect 6302 -1775 6366 -1774
rect 5896 -1818 5915 -1816
rect 5930 -1818 5964 -1816
rect 5896 -1834 5976 -1818
rect 5896 -1840 5915 -1834
rect 5612 -1866 5715 -1856
rect 5566 -1868 5715 -1866
rect 5736 -1868 5771 -1856
rect 5405 -1870 5567 -1868
rect 5417 -1888 5436 -1870
rect 5451 -1872 5481 -1870
rect 5300 -1898 5341 -1890
rect 5424 -1894 5436 -1888
rect 5488 -1886 5567 -1870
rect 5599 -1870 5771 -1868
rect 5599 -1886 5678 -1870
rect 5685 -1872 5715 -1870
rect 5263 -1908 5292 -1898
rect 5306 -1908 5335 -1898
rect 5350 -1908 5380 -1894
rect 5424 -1908 5466 -1894
rect 5488 -1898 5678 -1886
rect 5743 -1890 5749 -1870
rect 5473 -1908 5503 -1898
rect 5504 -1908 5662 -1898
rect 5666 -1908 5696 -1898
rect 5700 -1908 5730 -1894
rect 5758 -1908 5771 -1870
rect 5843 -1856 5872 -1840
rect 5886 -1856 5915 -1840
rect 5930 -1850 5960 -1834
rect 5988 -1856 5994 -1808
rect 5997 -1814 6016 -1808
rect 6031 -1814 6061 -1806
rect 5997 -1822 6061 -1814
rect 5997 -1838 6077 -1822
rect 6093 -1829 6155 -1798
rect 6171 -1829 6233 -1798
rect 6302 -1800 6351 -1775
rect 6366 -1800 6396 -1784
rect 6265 -1814 6295 -1806
rect 6302 -1808 6412 -1800
rect 6265 -1822 6310 -1814
rect 5997 -1840 6016 -1838
rect 6031 -1840 6077 -1838
rect 5997 -1856 6077 -1840
rect 6104 -1842 6139 -1829
rect 6180 -1832 6217 -1829
rect 6180 -1834 6222 -1832
rect 6109 -1845 6139 -1842
rect 6118 -1849 6125 -1845
rect 6125 -1850 6126 -1849
rect 6084 -1856 6094 -1850
rect 5843 -1864 5878 -1856
rect 5843 -1890 5844 -1864
rect 5851 -1890 5878 -1864
rect 5786 -1908 5816 -1894
rect 5843 -1898 5878 -1890
rect 5880 -1864 5921 -1856
rect 5880 -1890 5895 -1864
rect 5902 -1890 5921 -1864
rect 5985 -1868 6016 -1856
rect 6031 -1868 6134 -1856
rect 6146 -1866 6172 -1840
rect 6187 -1845 6217 -1834
rect 6249 -1838 6311 -1822
rect 6249 -1840 6295 -1838
rect 6249 -1856 6311 -1840
rect 6323 -1856 6329 -1808
rect 6332 -1816 6412 -1808
rect 6332 -1818 6351 -1816
rect 6366 -1818 6400 -1816
rect 6332 -1834 6412 -1818
rect 6332 -1856 6351 -1834
rect 6366 -1850 6396 -1834
rect 6424 -1840 6430 -1766
rect 6439 -1840 6452 -1696
rect 6192 -1866 6295 -1856
rect 6146 -1868 6295 -1866
rect 6316 -1868 6351 -1856
rect 5985 -1870 6147 -1868
rect 5997 -1888 6016 -1870
rect 6031 -1872 6061 -1870
rect 5880 -1898 5921 -1890
rect 6004 -1894 6016 -1888
rect 6068 -1886 6147 -1870
rect 6179 -1870 6351 -1868
rect 6179 -1886 6258 -1870
rect 6265 -1872 6295 -1870
rect 5843 -1908 5872 -1898
rect 5886 -1908 5915 -1898
rect 5930 -1908 5960 -1894
rect 6004 -1908 6046 -1894
rect 6068 -1898 6258 -1886
rect 6323 -1890 6329 -1870
rect 6053 -1908 6083 -1898
rect 6084 -1908 6242 -1898
rect 6246 -1908 6276 -1898
rect 6280 -1908 6310 -1894
rect 6338 -1908 6351 -1870
rect 6423 -1856 6452 -1840
rect 6423 -1864 6458 -1856
rect 6423 -1890 6424 -1864
rect 6431 -1890 6458 -1864
rect 6366 -1908 6396 -1894
rect 6423 -1898 6458 -1890
rect 6423 -1908 6452 -1898
rect -541 -1922 6452 -1908
rect -478 -1952 -465 -1922
rect -450 -1936 -420 -1922
rect -376 -1936 -334 -1922
rect -327 -1936 -107 -1922
rect -100 -1936 -70 -1922
rect -410 -1950 -395 -1938
rect -376 -1950 -363 -1936
rect -295 -1940 -142 -1936
rect -413 -1952 -391 -1950
rect -313 -1952 -121 -1940
rect -42 -1952 -29 -1922
rect -14 -1936 16 -1922
rect 53 -1952 72 -1922
rect 87 -1952 93 -1922
rect 102 -1952 115 -1922
rect 130 -1936 160 -1922
rect 204 -1936 246 -1922
rect 253 -1936 473 -1922
rect 480 -1936 510 -1922
rect 170 -1950 185 -1938
rect 204 -1950 217 -1936
rect 285 -1940 438 -1936
rect 167 -1952 189 -1950
rect 267 -1952 459 -1940
rect 538 -1952 551 -1922
rect 566 -1936 596 -1922
rect 633 -1952 652 -1922
rect 667 -1952 673 -1922
rect 682 -1952 695 -1922
rect 710 -1936 740 -1922
rect 784 -1936 826 -1922
rect 833 -1936 1053 -1922
rect 1060 -1936 1090 -1922
rect 750 -1950 765 -1938
rect 784 -1950 797 -1936
rect 865 -1940 1018 -1936
rect 747 -1952 769 -1950
rect 847 -1952 1039 -1940
rect 1118 -1952 1131 -1922
rect 1146 -1936 1176 -1922
rect 1213 -1952 1232 -1922
rect 1247 -1952 1253 -1922
rect 1262 -1952 1275 -1922
rect 1290 -1936 1320 -1922
rect 1364 -1936 1406 -1922
rect 1413 -1936 1633 -1922
rect 1640 -1936 1670 -1922
rect 1330 -1950 1345 -1938
rect 1364 -1950 1377 -1936
rect 1445 -1940 1598 -1936
rect 1327 -1952 1349 -1950
rect 1427 -1952 1619 -1940
rect 1698 -1952 1711 -1922
rect 1726 -1936 1756 -1922
rect 1793 -1952 1812 -1922
rect 1827 -1952 1833 -1922
rect 1842 -1952 1855 -1922
rect 1870 -1936 1900 -1922
rect 1944 -1936 1986 -1922
rect 1993 -1936 2213 -1922
rect 2220 -1936 2250 -1922
rect 1910 -1950 1925 -1938
rect 1944 -1950 1957 -1936
rect 2025 -1940 2178 -1936
rect 1907 -1952 1929 -1950
rect 2007 -1952 2199 -1940
rect 2278 -1952 2291 -1922
rect 2306 -1936 2336 -1922
rect 2373 -1952 2392 -1922
rect 2407 -1952 2413 -1922
rect 2422 -1952 2435 -1922
rect 2450 -1936 2480 -1922
rect 2524 -1936 2566 -1922
rect 2573 -1936 2793 -1922
rect 2800 -1936 2830 -1922
rect 2490 -1950 2505 -1938
rect 2524 -1950 2537 -1936
rect 2605 -1940 2758 -1936
rect 2487 -1952 2509 -1950
rect 2587 -1952 2779 -1940
rect 2858 -1952 2871 -1922
rect 2886 -1936 2916 -1922
rect 2953 -1952 2972 -1922
rect 2987 -1952 2993 -1922
rect 3002 -1952 3015 -1922
rect 3030 -1936 3060 -1922
rect 3104 -1936 3146 -1922
rect 3153 -1936 3373 -1922
rect 3380 -1936 3410 -1922
rect 3070 -1950 3085 -1938
rect 3104 -1950 3117 -1936
rect 3185 -1940 3338 -1936
rect 3067 -1952 3089 -1950
rect 3167 -1952 3359 -1940
rect 3438 -1952 3451 -1922
rect 3466 -1936 3496 -1922
rect 3533 -1952 3552 -1922
rect 3567 -1952 3573 -1922
rect 3582 -1952 3595 -1922
rect 3610 -1936 3640 -1922
rect 3684 -1936 3726 -1922
rect 3733 -1936 3953 -1922
rect 3960 -1936 3990 -1922
rect 3650 -1950 3665 -1938
rect 3684 -1950 3697 -1936
rect 3765 -1940 3918 -1936
rect 3647 -1952 3669 -1950
rect 3747 -1952 3939 -1940
rect 4018 -1952 4031 -1922
rect 4046 -1936 4076 -1922
rect 4113 -1952 4132 -1922
rect 4147 -1952 4153 -1922
rect 4162 -1952 4175 -1922
rect 4190 -1936 4220 -1922
rect 4264 -1936 4306 -1922
rect 4313 -1936 4533 -1922
rect 4540 -1936 4570 -1922
rect 4230 -1950 4245 -1938
rect 4264 -1950 4277 -1936
rect 4345 -1940 4498 -1936
rect 4227 -1952 4249 -1950
rect 4327 -1952 4519 -1940
rect 4598 -1952 4611 -1922
rect 4626 -1936 4656 -1922
rect 4693 -1952 4712 -1922
rect 4727 -1952 4733 -1922
rect 4742 -1952 4755 -1922
rect 4770 -1936 4800 -1922
rect 4844 -1936 4886 -1922
rect 4893 -1936 5113 -1922
rect 5120 -1936 5150 -1922
rect 4810 -1950 4825 -1938
rect 4844 -1950 4857 -1936
rect 4925 -1940 5078 -1936
rect 4807 -1952 4829 -1950
rect 4907 -1952 5099 -1940
rect 5178 -1952 5191 -1922
rect 5206 -1936 5236 -1922
rect 5273 -1952 5292 -1922
rect 5307 -1952 5313 -1922
rect 5322 -1952 5335 -1922
rect 5350 -1936 5380 -1922
rect 5424 -1936 5466 -1922
rect 5473 -1936 5693 -1922
rect 5700 -1936 5730 -1922
rect 5390 -1950 5405 -1938
rect 5424 -1950 5437 -1936
rect 5505 -1940 5658 -1936
rect 5387 -1952 5409 -1950
rect 5487 -1952 5679 -1940
rect 5758 -1952 5771 -1922
rect 5786 -1936 5816 -1922
rect 5853 -1952 5872 -1922
rect 5887 -1952 5893 -1922
rect 5902 -1952 5915 -1922
rect 5930 -1936 5960 -1922
rect 6004 -1936 6046 -1922
rect 6053 -1936 6273 -1922
rect 6280 -1936 6310 -1922
rect 5970 -1950 5985 -1938
rect 6004 -1950 6017 -1936
rect 6085 -1940 6238 -1936
rect 5967 -1952 5989 -1950
rect 6067 -1952 6259 -1940
rect 6338 -1952 6351 -1922
rect 6366 -1936 6396 -1922
rect 6439 -1952 6452 -1922
rect -541 -1966 6452 -1952
rect -478 -2036 -465 -1966
rect -413 -1970 -391 -1966
rect -420 -1982 -403 -1978
rect -399 -1980 -391 -1978
rect -401 -1982 -391 -1980
rect -420 -1992 -391 -1982
rect -338 -1992 -322 -1978
rect -284 -1982 -278 -1980
rect -271 -1982 -163 -1966
rect -156 -1982 -150 -1980
rect -142 -1982 -127 -1966
rect -61 -1972 -42 -1969
rect -420 -1994 -322 -1992
rect -295 -1994 -127 -1982
rect -112 -1992 -96 -1978
rect -61 -1991 -39 -1972
rect -29 -1978 -13 -1977
rect -30 -1980 -13 -1978
rect -29 -1985 -13 -1980
rect -39 -1992 -33 -1991
rect -30 -1992 -1 -1985
rect -112 -1993 -1 -1992
rect -112 -1994 5 -1993
rect -436 -2002 -385 -1994
rect -338 -2002 -304 -1994
rect -436 -2014 -411 -2002
rect -404 -2014 -385 -2002
rect -331 -2004 -304 -2002
rect -295 -2004 -74 -1994
rect -39 -1997 -33 -1994
rect -331 -2008 -74 -2004
rect -436 -2022 -385 -2014
rect -338 -2022 -74 -2008
rect -30 -2002 5 -1994
rect -484 -2070 -465 -2036
rect -420 -2030 -391 -2022
rect -420 -2036 -403 -2030
rect -420 -2038 -386 -2036
rect -338 -2038 -322 -2022
rect -321 -2032 -113 -2022
rect -112 -2032 -96 -2022
rect -48 -2026 -33 -2011
rect -30 -2014 -29 -2002
rect -22 -2014 5 -2002
rect -30 -2022 5 -2014
rect -30 -2023 -1 -2022
rect -310 -2036 -96 -2032
rect -295 -2038 -96 -2036
rect -61 -2036 -48 -2026
rect -30 -2036 -13 -2023
rect -61 -2038 -13 -2036
rect -419 -2042 -386 -2038
rect -423 -2044 -386 -2042
rect -423 -2045 -356 -2044
rect -423 -2050 -392 -2045
rect -386 -2050 -356 -2045
rect -423 -2054 -356 -2050
rect -450 -2057 -356 -2054
rect -450 -2064 -401 -2057
rect -450 -2070 -420 -2064
rect -401 -2069 -396 -2064
rect -484 -2086 -404 -2070
rect -392 -2078 -356 -2057
rect -295 -2062 -106 -2038
rect -61 -2039 -14 -2038
rect -48 -2044 -14 -2039
rect -280 -2065 -106 -2062
rect -287 -2068 -106 -2065
rect -78 -2045 -14 -2044
rect -484 -2088 -465 -2086
rect -450 -2088 -416 -2086
rect -484 -2104 -404 -2088
rect -484 -2110 -465 -2104
rect -494 -2126 -465 -2110
rect -450 -2120 -420 -2104
rect -392 -2126 -386 -2078
rect -383 -2084 -364 -2078
rect -349 -2084 -319 -2076
rect -383 -2092 -319 -2084
rect -383 -2108 -303 -2092
rect -287 -2099 -225 -2068
rect -209 -2099 -147 -2068
rect -78 -2070 -29 -2045
rect -14 -2070 16 -2052
rect -115 -2084 -85 -2076
rect -78 -2078 32 -2070
rect -115 -2092 -70 -2084
rect -383 -2110 -364 -2108
rect -349 -2110 -303 -2108
rect -383 -2126 -303 -2110
rect -276 -2112 -241 -2099
rect -200 -2102 -163 -2099
rect -200 -2104 -158 -2102
rect -271 -2115 -241 -2112
rect -262 -2119 -255 -2115
rect -255 -2120 -254 -2119
rect -296 -2126 -286 -2120
rect -500 -2134 -459 -2126
rect -500 -2160 -485 -2134
rect -478 -2160 -459 -2134
rect -395 -2138 -364 -2126
rect -349 -2138 -246 -2126
rect -234 -2136 -208 -2110
rect -193 -2115 -163 -2104
rect -131 -2108 -69 -2092
rect -131 -2110 -85 -2108
rect -131 -2126 -69 -2110
rect -57 -2126 -51 -2078
rect -48 -2086 32 -2078
rect -48 -2088 -29 -2086
rect -14 -2088 20 -2086
rect -48 -2103 32 -2088
rect -48 -2104 38 -2103
rect -48 -2126 -29 -2104
rect -14 -2120 16 -2104
rect 44 -2110 50 -2036
rect 53 -2110 72 -1966
rect 87 -2110 93 -1966
rect 102 -2036 115 -1966
rect 167 -1970 189 -1966
rect 160 -1982 177 -1978
rect 181 -1980 189 -1978
rect 179 -1982 189 -1980
rect 160 -1992 189 -1982
rect 242 -1992 258 -1978
rect 296 -1982 302 -1980
rect 309 -1982 417 -1966
rect 424 -1982 430 -1980
rect 438 -1982 453 -1966
rect 519 -1972 538 -1969
rect 160 -1994 258 -1992
rect 285 -1994 453 -1982
rect 468 -1992 484 -1978
rect 519 -1991 541 -1972
rect 551 -1978 567 -1977
rect 550 -1980 567 -1978
rect 551 -1985 567 -1980
rect 541 -1992 547 -1991
rect 550 -1992 579 -1985
rect 468 -1993 579 -1992
rect 468 -1994 585 -1993
rect 144 -2002 195 -1994
rect 242 -2002 276 -1994
rect 144 -2014 169 -2002
rect 176 -2014 195 -2002
rect 249 -2004 276 -2002
rect 285 -2004 506 -1994
rect 541 -1997 547 -1994
rect 249 -2008 506 -2004
rect 144 -2022 195 -2014
rect 242 -2022 506 -2008
rect 550 -2002 585 -1994
rect 96 -2070 115 -2036
rect 160 -2030 189 -2022
rect 160 -2036 177 -2030
rect 160 -2038 194 -2036
rect 242 -2038 258 -2022
rect 259 -2032 467 -2022
rect 468 -2032 484 -2022
rect 532 -2026 547 -2011
rect 550 -2014 551 -2002
rect 558 -2014 585 -2002
rect 550 -2022 585 -2014
rect 550 -2023 579 -2022
rect 270 -2036 484 -2032
rect 285 -2038 484 -2036
rect 519 -2036 532 -2026
rect 550 -2036 567 -2023
rect 519 -2038 567 -2036
rect 161 -2042 194 -2038
rect 157 -2044 194 -2042
rect 157 -2045 224 -2044
rect 157 -2050 188 -2045
rect 194 -2050 224 -2045
rect 157 -2054 224 -2050
rect 130 -2057 224 -2054
rect 130 -2064 179 -2057
rect 130 -2070 160 -2064
rect 179 -2069 184 -2064
rect 96 -2086 176 -2070
rect 188 -2078 224 -2057
rect 285 -2062 474 -2038
rect 519 -2039 566 -2038
rect 532 -2044 566 -2039
rect 606 -2044 622 -2042
rect 300 -2065 474 -2062
rect 293 -2068 474 -2065
rect 502 -2045 566 -2044
rect 96 -2088 115 -2086
rect 130 -2088 164 -2086
rect 96 -2104 176 -2088
rect 96 -2110 115 -2104
rect -188 -2136 -85 -2126
rect -234 -2138 -85 -2136
rect -64 -2138 -29 -2126
rect -395 -2140 -233 -2138
rect -383 -2160 -364 -2140
rect -349 -2142 -319 -2140
rect -500 -2168 -459 -2160
rect -377 -2164 -364 -2160
rect -312 -2156 -233 -2140
rect -201 -2140 -29 -2138
rect -201 -2156 -122 -2140
rect -115 -2142 -85 -2140
rect -494 -2178 -465 -2168
rect -450 -2178 -420 -2164
rect -377 -2178 -334 -2164
rect -312 -2168 -122 -2156
rect -57 -2160 -51 -2140
rect -327 -2178 -297 -2168
rect -296 -2178 -138 -2168
rect -134 -2178 -104 -2168
rect -100 -2178 -70 -2164
rect -42 -2178 -29 -2140
rect 43 -2126 72 -2110
rect 86 -2126 115 -2110
rect 130 -2120 160 -2104
rect 188 -2126 194 -2078
rect 197 -2084 216 -2078
rect 231 -2084 261 -2076
rect 197 -2092 261 -2084
rect 197 -2108 277 -2092
rect 293 -2099 355 -2068
rect 371 -2099 433 -2068
rect 502 -2070 551 -2045
rect 596 -2054 622 -2044
rect 566 -2070 622 -2054
rect 465 -2084 495 -2076
rect 502 -2078 612 -2070
rect 465 -2092 510 -2084
rect 197 -2110 216 -2108
rect 231 -2110 277 -2108
rect 197 -2126 277 -2110
rect 304 -2112 339 -2099
rect 380 -2102 417 -2099
rect 380 -2104 422 -2102
rect 309 -2115 339 -2112
rect 318 -2119 325 -2115
rect 325 -2120 326 -2119
rect 284 -2126 294 -2120
rect 43 -2134 78 -2126
rect 43 -2160 44 -2134
rect 51 -2160 78 -2134
rect -14 -2178 16 -2164
rect 43 -2168 78 -2160
rect 80 -2134 121 -2126
rect 80 -2160 95 -2134
rect 102 -2160 121 -2134
rect 185 -2138 216 -2126
rect 231 -2138 334 -2126
rect 346 -2136 372 -2110
rect 387 -2115 417 -2104
rect 449 -2108 511 -2092
rect 449 -2110 495 -2108
rect 449 -2126 511 -2110
rect 523 -2126 529 -2078
rect 532 -2086 612 -2078
rect 532 -2088 551 -2086
rect 566 -2088 600 -2086
rect 532 -2104 612 -2088
rect 532 -2126 551 -2104
rect 566 -2120 596 -2104
rect 624 -2110 630 -2036
rect 633 -2110 652 -1966
rect 667 -2110 673 -1966
rect 682 -2036 695 -1966
rect 747 -1970 769 -1966
rect 740 -1982 757 -1978
rect 761 -1980 769 -1978
rect 759 -1982 769 -1980
rect 740 -1992 769 -1982
rect 822 -1992 838 -1978
rect 876 -1982 882 -1980
rect 889 -1982 997 -1966
rect 1004 -1982 1010 -1980
rect 1018 -1982 1033 -1966
rect 1099 -1972 1118 -1969
rect 740 -1994 838 -1992
rect 865 -1994 1033 -1982
rect 1048 -1992 1064 -1978
rect 1099 -1991 1121 -1972
rect 1131 -1978 1147 -1977
rect 1130 -1980 1147 -1978
rect 1131 -1985 1147 -1980
rect 1121 -1992 1127 -1991
rect 1130 -1992 1159 -1985
rect 1048 -1993 1159 -1992
rect 1048 -1994 1165 -1993
rect 724 -2002 775 -1994
rect 822 -2002 856 -1994
rect 724 -2014 749 -2002
rect 756 -2014 775 -2002
rect 829 -2004 856 -2002
rect 865 -2004 1086 -1994
rect 1121 -1997 1127 -1994
rect 829 -2008 1086 -2004
rect 724 -2022 775 -2014
rect 822 -2022 1086 -2008
rect 1130 -2002 1165 -1994
rect 676 -2070 695 -2036
rect 740 -2030 769 -2022
rect 740 -2036 757 -2030
rect 740 -2038 774 -2036
rect 822 -2038 838 -2022
rect 839 -2032 1047 -2022
rect 1048 -2032 1064 -2022
rect 1112 -2026 1127 -2011
rect 1130 -2014 1131 -2002
rect 1138 -2014 1165 -2002
rect 1130 -2022 1165 -2014
rect 1130 -2023 1159 -2022
rect 850 -2036 1064 -2032
rect 865 -2038 1064 -2036
rect 1099 -2036 1112 -2026
rect 1130 -2036 1147 -2023
rect 1099 -2038 1147 -2036
rect 741 -2042 774 -2038
rect 737 -2044 774 -2042
rect 737 -2045 804 -2044
rect 737 -2050 768 -2045
rect 774 -2050 804 -2045
rect 737 -2054 804 -2050
rect 710 -2057 804 -2054
rect 710 -2064 759 -2057
rect 710 -2070 740 -2064
rect 759 -2069 764 -2064
rect 676 -2086 756 -2070
rect 768 -2078 804 -2057
rect 865 -2062 1054 -2038
rect 1099 -2039 1146 -2038
rect 1112 -2044 1146 -2039
rect 880 -2065 1054 -2062
rect 873 -2068 1054 -2065
rect 1082 -2045 1146 -2044
rect 676 -2088 695 -2086
rect 710 -2088 744 -2086
rect 676 -2104 756 -2088
rect 676 -2110 695 -2104
rect 392 -2136 495 -2126
rect 346 -2138 495 -2136
rect 516 -2138 551 -2126
rect 185 -2140 347 -2138
rect 197 -2160 216 -2140
rect 231 -2142 261 -2140
rect 80 -2168 121 -2160
rect 203 -2164 216 -2160
rect 268 -2156 347 -2140
rect 379 -2140 551 -2138
rect 379 -2156 458 -2140
rect 465 -2142 495 -2140
rect 43 -2178 72 -2168
rect 86 -2178 115 -2168
rect 130 -2178 160 -2164
rect 203 -2178 246 -2164
rect 268 -2168 458 -2156
rect 523 -2160 529 -2140
rect 253 -2178 283 -2168
rect 284 -2178 442 -2168
rect 446 -2178 476 -2168
rect 480 -2178 510 -2164
rect 538 -2178 551 -2140
rect 623 -2126 652 -2110
rect 666 -2126 695 -2110
rect 710 -2120 740 -2104
rect 768 -2126 774 -2078
rect 777 -2084 796 -2078
rect 811 -2084 841 -2076
rect 777 -2092 841 -2084
rect 777 -2108 857 -2092
rect 873 -2099 935 -2068
rect 951 -2099 1013 -2068
rect 1082 -2070 1131 -2045
rect 1146 -2070 1176 -2052
rect 1045 -2084 1075 -2076
rect 1082 -2078 1192 -2070
rect 1045 -2092 1090 -2084
rect 777 -2110 796 -2108
rect 811 -2110 857 -2108
rect 777 -2126 857 -2110
rect 884 -2112 919 -2099
rect 960 -2102 997 -2099
rect 960 -2104 1002 -2102
rect 889 -2115 919 -2112
rect 898 -2119 905 -2115
rect 905 -2120 906 -2119
rect 864 -2126 874 -2120
rect 623 -2134 658 -2126
rect 623 -2160 624 -2134
rect 631 -2160 658 -2134
rect 566 -2178 596 -2164
rect 623 -2168 658 -2160
rect 660 -2134 701 -2126
rect 660 -2160 675 -2134
rect 682 -2160 701 -2134
rect 765 -2138 796 -2126
rect 811 -2138 914 -2126
rect 926 -2136 952 -2110
rect 967 -2115 997 -2104
rect 1029 -2108 1091 -2092
rect 1029 -2110 1075 -2108
rect 1029 -2126 1091 -2110
rect 1103 -2126 1109 -2078
rect 1112 -2086 1192 -2078
rect 1112 -2088 1131 -2086
rect 1146 -2088 1180 -2086
rect 1112 -2103 1192 -2088
rect 1112 -2104 1198 -2103
rect 1112 -2126 1131 -2104
rect 1146 -2120 1176 -2104
rect 1204 -2110 1210 -2036
rect 1213 -2110 1232 -1966
rect 1247 -2110 1253 -1966
rect 1262 -2036 1275 -1966
rect 1327 -1970 1349 -1966
rect 1320 -1982 1337 -1978
rect 1341 -1980 1349 -1978
rect 1339 -1982 1349 -1980
rect 1320 -1992 1349 -1982
rect 1402 -1992 1418 -1978
rect 1456 -1982 1462 -1980
rect 1469 -1982 1577 -1966
rect 1584 -1982 1590 -1980
rect 1598 -1982 1613 -1966
rect 1679 -1972 1698 -1969
rect 1320 -1994 1418 -1992
rect 1445 -1994 1613 -1982
rect 1628 -1992 1644 -1978
rect 1679 -1991 1701 -1972
rect 1711 -1978 1727 -1977
rect 1710 -1980 1727 -1978
rect 1711 -1985 1727 -1980
rect 1701 -1992 1707 -1991
rect 1710 -1992 1739 -1985
rect 1628 -1993 1739 -1992
rect 1628 -1994 1745 -1993
rect 1304 -2002 1355 -1994
rect 1402 -2002 1436 -1994
rect 1304 -2014 1329 -2002
rect 1336 -2014 1355 -2002
rect 1409 -2004 1436 -2002
rect 1445 -2004 1666 -1994
rect 1701 -1997 1707 -1994
rect 1409 -2008 1666 -2004
rect 1304 -2022 1355 -2014
rect 1402 -2022 1666 -2008
rect 1710 -2002 1745 -1994
rect 1256 -2070 1275 -2036
rect 1320 -2030 1349 -2022
rect 1320 -2036 1337 -2030
rect 1320 -2038 1354 -2036
rect 1402 -2038 1418 -2022
rect 1419 -2032 1627 -2022
rect 1628 -2032 1644 -2022
rect 1692 -2026 1707 -2011
rect 1710 -2014 1711 -2002
rect 1718 -2014 1745 -2002
rect 1710 -2022 1745 -2014
rect 1710 -2023 1739 -2022
rect 1430 -2036 1644 -2032
rect 1445 -2038 1644 -2036
rect 1679 -2036 1692 -2026
rect 1710 -2036 1727 -2023
rect 1679 -2038 1727 -2036
rect 1321 -2042 1354 -2038
rect 1317 -2044 1354 -2042
rect 1317 -2045 1384 -2044
rect 1317 -2050 1348 -2045
rect 1354 -2050 1384 -2045
rect 1317 -2054 1384 -2050
rect 1290 -2057 1384 -2054
rect 1290 -2064 1339 -2057
rect 1290 -2070 1320 -2064
rect 1339 -2069 1344 -2064
rect 1256 -2086 1336 -2070
rect 1348 -2078 1384 -2057
rect 1445 -2062 1634 -2038
rect 1679 -2039 1726 -2038
rect 1692 -2044 1726 -2039
rect 1766 -2044 1782 -2042
rect 1460 -2065 1634 -2062
rect 1453 -2068 1634 -2065
rect 1662 -2045 1726 -2044
rect 1256 -2088 1275 -2086
rect 1290 -2088 1324 -2086
rect 1256 -2104 1336 -2088
rect 1256 -2110 1275 -2104
rect 972 -2136 1075 -2126
rect 926 -2138 1075 -2136
rect 1096 -2138 1131 -2126
rect 765 -2140 927 -2138
rect 777 -2160 796 -2140
rect 811 -2142 841 -2140
rect 660 -2168 701 -2160
rect 783 -2164 796 -2160
rect 848 -2156 927 -2140
rect 959 -2140 1131 -2138
rect 959 -2156 1038 -2140
rect 1045 -2142 1075 -2140
rect 623 -2178 652 -2168
rect 666 -2178 695 -2168
rect 710 -2178 740 -2164
rect 783 -2178 826 -2164
rect 848 -2168 1038 -2156
rect 1103 -2160 1109 -2140
rect 833 -2178 863 -2168
rect 864 -2178 1022 -2168
rect 1026 -2178 1056 -2168
rect 1060 -2178 1090 -2164
rect 1118 -2178 1131 -2140
rect 1203 -2126 1232 -2110
rect 1246 -2126 1275 -2110
rect 1290 -2120 1320 -2104
rect 1348 -2126 1354 -2078
rect 1357 -2084 1376 -2078
rect 1391 -2084 1421 -2076
rect 1357 -2092 1421 -2084
rect 1357 -2108 1437 -2092
rect 1453 -2099 1515 -2068
rect 1531 -2099 1593 -2068
rect 1662 -2070 1711 -2045
rect 1756 -2054 1782 -2044
rect 1726 -2070 1782 -2054
rect 1625 -2084 1655 -2076
rect 1662 -2078 1772 -2070
rect 1625 -2092 1670 -2084
rect 1357 -2110 1376 -2108
rect 1391 -2110 1437 -2108
rect 1357 -2126 1437 -2110
rect 1464 -2112 1499 -2099
rect 1540 -2102 1577 -2099
rect 1540 -2104 1582 -2102
rect 1469 -2115 1499 -2112
rect 1478 -2119 1485 -2115
rect 1485 -2120 1486 -2119
rect 1444 -2126 1454 -2120
rect 1203 -2134 1238 -2126
rect 1203 -2160 1204 -2134
rect 1211 -2160 1238 -2134
rect 1146 -2178 1176 -2164
rect 1203 -2168 1238 -2160
rect 1240 -2134 1281 -2126
rect 1240 -2160 1255 -2134
rect 1262 -2160 1281 -2134
rect 1345 -2138 1376 -2126
rect 1391 -2138 1494 -2126
rect 1506 -2136 1532 -2110
rect 1547 -2115 1577 -2104
rect 1609 -2108 1671 -2092
rect 1609 -2110 1655 -2108
rect 1609 -2126 1671 -2110
rect 1683 -2126 1689 -2078
rect 1692 -2086 1772 -2078
rect 1692 -2088 1711 -2086
rect 1726 -2088 1760 -2086
rect 1692 -2104 1772 -2088
rect 1692 -2126 1711 -2104
rect 1726 -2120 1756 -2104
rect 1784 -2110 1790 -2036
rect 1793 -2110 1812 -1966
rect 1827 -2110 1833 -1966
rect 1842 -2036 1855 -1966
rect 1907 -1970 1929 -1966
rect 1900 -1982 1917 -1978
rect 1921 -1980 1929 -1978
rect 1919 -1982 1929 -1980
rect 1900 -1992 1929 -1982
rect 1982 -1992 1998 -1978
rect 2036 -1982 2042 -1980
rect 2049 -1982 2157 -1966
rect 2164 -1982 2170 -1980
rect 2178 -1982 2193 -1966
rect 2259 -1972 2278 -1969
rect 1900 -1994 1998 -1992
rect 2025 -1994 2193 -1982
rect 2208 -1992 2224 -1978
rect 2259 -1991 2281 -1972
rect 2291 -1978 2307 -1977
rect 2290 -1984 2307 -1978
rect 2291 -1985 2307 -1984
rect 2281 -1992 2287 -1991
rect 2290 -1992 2319 -1985
rect 2208 -1993 2319 -1992
rect 2208 -1994 2325 -1993
rect 1884 -2002 1935 -1994
rect 1982 -2002 2016 -1994
rect 1884 -2014 1909 -2002
rect 1916 -2014 1935 -2002
rect 1989 -2004 2016 -2002
rect 2025 -2004 2246 -1994
rect 2281 -1997 2287 -1994
rect 1989 -2008 2246 -2004
rect 1884 -2022 1935 -2014
rect 1982 -2022 2246 -2008
rect 2290 -2002 2325 -1994
rect 1836 -2070 1855 -2036
rect 1900 -2030 1929 -2022
rect 1900 -2036 1917 -2030
rect 1900 -2038 1934 -2036
rect 1982 -2038 1998 -2022
rect 1999 -2032 2207 -2022
rect 2208 -2032 2224 -2022
rect 2272 -2026 2287 -2011
rect 2290 -2014 2291 -2002
rect 2298 -2014 2325 -2002
rect 2290 -2022 2325 -2014
rect 2290 -2023 2319 -2022
rect 2010 -2036 2224 -2032
rect 2025 -2038 2224 -2036
rect 2259 -2036 2272 -2026
rect 2290 -2036 2307 -2023
rect 2259 -2038 2307 -2036
rect 1901 -2042 1934 -2038
rect 1897 -2044 1934 -2042
rect 1897 -2045 1964 -2044
rect 1897 -2050 1928 -2045
rect 1934 -2050 1964 -2045
rect 1897 -2054 1964 -2050
rect 1870 -2057 1964 -2054
rect 1870 -2064 1919 -2057
rect 1870 -2070 1900 -2064
rect 1919 -2069 1924 -2064
rect 1836 -2086 1916 -2070
rect 1928 -2078 1964 -2057
rect 2025 -2062 2214 -2038
rect 2259 -2039 2306 -2038
rect 2272 -2044 2306 -2039
rect 2040 -2065 2214 -2062
rect 2033 -2068 2214 -2065
rect 2242 -2045 2306 -2044
rect 1836 -2088 1855 -2086
rect 1870 -2088 1904 -2086
rect 1836 -2104 1916 -2088
rect 1836 -2110 1855 -2104
rect 1552 -2136 1655 -2126
rect 1506 -2138 1655 -2136
rect 1676 -2138 1711 -2126
rect 1345 -2140 1507 -2138
rect 1357 -2160 1376 -2140
rect 1391 -2142 1421 -2140
rect 1240 -2168 1281 -2160
rect 1363 -2164 1376 -2160
rect 1428 -2156 1507 -2140
rect 1539 -2140 1711 -2138
rect 1539 -2156 1618 -2140
rect 1625 -2142 1655 -2140
rect 1203 -2178 1232 -2168
rect 1246 -2178 1275 -2168
rect 1290 -2178 1320 -2164
rect 1363 -2178 1406 -2164
rect 1428 -2168 1618 -2156
rect 1683 -2160 1689 -2140
rect 1413 -2178 1443 -2168
rect 1444 -2178 1602 -2168
rect 1606 -2178 1636 -2168
rect 1640 -2178 1670 -2164
rect 1698 -2178 1711 -2140
rect 1783 -2126 1812 -2110
rect 1826 -2126 1855 -2110
rect 1870 -2120 1900 -2104
rect 1928 -2126 1934 -2078
rect 1937 -2084 1956 -2078
rect 1971 -2084 2001 -2076
rect 1937 -2092 2001 -2084
rect 1937 -2108 2017 -2092
rect 2033 -2099 2095 -2068
rect 2111 -2099 2173 -2068
rect 2242 -2070 2291 -2045
rect 2306 -2070 2336 -2052
rect 2205 -2084 2235 -2076
rect 2242 -2078 2352 -2070
rect 2205 -2092 2250 -2084
rect 1937 -2110 1956 -2108
rect 1971 -2110 2017 -2108
rect 1937 -2126 2017 -2110
rect 2044 -2112 2079 -2099
rect 2120 -2102 2157 -2099
rect 2120 -2104 2162 -2102
rect 2049 -2115 2079 -2112
rect 2058 -2119 2065 -2115
rect 2065 -2120 2066 -2119
rect 2024 -2126 2034 -2120
rect 1783 -2134 1818 -2126
rect 1783 -2160 1784 -2134
rect 1791 -2160 1818 -2134
rect 1726 -2178 1756 -2164
rect 1783 -2168 1818 -2160
rect 1820 -2134 1861 -2126
rect 1820 -2160 1835 -2134
rect 1842 -2160 1861 -2134
rect 1925 -2138 1956 -2126
rect 1971 -2138 2074 -2126
rect 2086 -2136 2112 -2110
rect 2127 -2115 2157 -2104
rect 2189 -2108 2251 -2092
rect 2189 -2110 2235 -2108
rect 2189 -2126 2251 -2110
rect 2263 -2126 2269 -2078
rect 2272 -2086 2352 -2078
rect 2272 -2088 2291 -2086
rect 2306 -2088 2340 -2086
rect 2272 -2103 2352 -2088
rect 2272 -2104 2358 -2103
rect 2272 -2126 2291 -2104
rect 2306 -2120 2336 -2104
rect 2364 -2110 2370 -2036
rect 2373 -2110 2392 -1966
rect 2407 -2110 2413 -1966
rect 2422 -2036 2435 -1966
rect 2487 -1970 2509 -1966
rect 2480 -1982 2497 -1978
rect 2501 -1980 2509 -1978
rect 2499 -1982 2509 -1980
rect 2480 -1992 2509 -1982
rect 2562 -1992 2578 -1978
rect 2616 -1982 2622 -1980
rect 2629 -1982 2737 -1966
rect 2744 -1982 2750 -1980
rect 2758 -1982 2773 -1966
rect 2839 -1972 2858 -1969
rect 2480 -1994 2578 -1992
rect 2605 -1994 2773 -1982
rect 2788 -1992 2804 -1978
rect 2839 -1991 2861 -1972
rect 2871 -1978 2887 -1977
rect 2870 -1984 2887 -1978
rect 2871 -1985 2887 -1984
rect 2861 -1992 2867 -1991
rect 2870 -1992 2899 -1985
rect 2788 -1993 2899 -1992
rect 2788 -1994 2905 -1993
rect 2464 -2002 2515 -1994
rect 2562 -2002 2596 -1994
rect 2464 -2014 2489 -2002
rect 2496 -2014 2515 -2002
rect 2569 -2004 2596 -2002
rect 2605 -2004 2826 -1994
rect 2861 -1997 2867 -1994
rect 2569 -2008 2826 -2004
rect 2464 -2022 2515 -2014
rect 2562 -2022 2826 -2008
rect 2870 -2002 2905 -1994
rect 2416 -2070 2435 -2036
rect 2480 -2030 2509 -2022
rect 2480 -2036 2497 -2030
rect 2480 -2038 2514 -2036
rect 2562 -2038 2578 -2022
rect 2579 -2032 2787 -2022
rect 2788 -2032 2804 -2022
rect 2852 -2026 2867 -2011
rect 2870 -2014 2871 -2002
rect 2878 -2014 2905 -2002
rect 2870 -2022 2905 -2014
rect 2870 -2023 2899 -2022
rect 2590 -2036 2804 -2032
rect 2605 -2038 2804 -2036
rect 2839 -2036 2852 -2026
rect 2870 -2036 2887 -2023
rect 2839 -2038 2887 -2036
rect 2481 -2042 2514 -2038
rect 2477 -2044 2514 -2042
rect 2477 -2045 2544 -2044
rect 2477 -2050 2508 -2045
rect 2514 -2050 2544 -2045
rect 2477 -2054 2544 -2050
rect 2450 -2057 2544 -2054
rect 2450 -2064 2499 -2057
rect 2450 -2070 2480 -2064
rect 2499 -2069 2504 -2064
rect 2416 -2086 2496 -2070
rect 2508 -2078 2544 -2057
rect 2605 -2062 2794 -2038
rect 2839 -2039 2886 -2038
rect 2852 -2044 2886 -2039
rect 2926 -2044 2942 -2042
rect 2620 -2065 2794 -2062
rect 2613 -2068 2794 -2065
rect 2822 -2045 2886 -2044
rect 2416 -2088 2435 -2086
rect 2450 -2088 2484 -2086
rect 2416 -2104 2496 -2088
rect 2416 -2110 2435 -2104
rect 2132 -2136 2235 -2126
rect 2086 -2138 2235 -2136
rect 2256 -2138 2291 -2126
rect 1925 -2140 2087 -2138
rect 1937 -2160 1956 -2140
rect 1971 -2142 2001 -2140
rect 1820 -2168 1861 -2160
rect 1943 -2164 1956 -2160
rect 2008 -2156 2087 -2140
rect 2119 -2140 2291 -2138
rect 2119 -2156 2198 -2140
rect 2205 -2142 2235 -2140
rect 1783 -2178 1812 -2168
rect 1826 -2178 1855 -2168
rect 1870 -2178 1900 -2164
rect 1943 -2178 1986 -2164
rect 2008 -2168 2198 -2156
rect 2263 -2160 2269 -2140
rect 1993 -2178 2023 -2168
rect 2024 -2178 2182 -2168
rect 2186 -2178 2216 -2168
rect 2220 -2178 2250 -2164
rect 2278 -2178 2291 -2140
rect 2363 -2126 2392 -2110
rect 2406 -2126 2435 -2110
rect 2450 -2120 2480 -2104
rect 2508 -2126 2514 -2078
rect 2517 -2084 2536 -2078
rect 2551 -2084 2581 -2076
rect 2517 -2092 2581 -2084
rect 2517 -2108 2597 -2092
rect 2613 -2099 2675 -2068
rect 2691 -2099 2753 -2068
rect 2822 -2070 2871 -2045
rect 2916 -2054 2942 -2044
rect 2886 -2070 2942 -2054
rect 2785 -2084 2815 -2076
rect 2822 -2078 2932 -2070
rect 2785 -2092 2830 -2084
rect 2517 -2110 2536 -2108
rect 2551 -2110 2597 -2108
rect 2517 -2126 2597 -2110
rect 2624 -2112 2659 -2099
rect 2700 -2102 2737 -2099
rect 2700 -2104 2742 -2102
rect 2629 -2115 2659 -2112
rect 2638 -2119 2645 -2115
rect 2645 -2120 2646 -2119
rect 2604 -2126 2614 -2120
rect 2363 -2134 2398 -2126
rect 2363 -2160 2364 -2134
rect 2371 -2160 2398 -2134
rect 2306 -2178 2336 -2164
rect 2363 -2168 2398 -2160
rect 2400 -2134 2441 -2126
rect 2400 -2160 2415 -2134
rect 2422 -2160 2441 -2134
rect 2505 -2138 2536 -2126
rect 2551 -2138 2654 -2126
rect 2666 -2136 2692 -2110
rect 2707 -2115 2737 -2104
rect 2769 -2108 2831 -2092
rect 2769 -2110 2815 -2108
rect 2769 -2126 2831 -2110
rect 2843 -2126 2849 -2078
rect 2852 -2086 2932 -2078
rect 2852 -2088 2871 -2086
rect 2886 -2088 2920 -2086
rect 2852 -2104 2932 -2088
rect 2852 -2126 2871 -2104
rect 2886 -2120 2916 -2104
rect 2944 -2110 2950 -2036
rect 2953 -2110 2972 -1966
rect 2987 -2110 2993 -1966
rect 3002 -2036 3015 -1966
rect 3067 -1970 3089 -1966
rect 3060 -1982 3077 -1978
rect 3081 -1980 3089 -1978
rect 3079 -1982 3089 -1980
rect 3060 -1992 3089 -1982
rect 3142 -1992 3158 -1978
rect 3196 -1982 3202 -1980
rect 3209 -1982 3317 -1966
rect 3324 -1982 3330 -1980
rect 3338 -1982 3353 -1966
rect 3419 -1972 3438 -1969
rect 3060 -1994 3158 -1992
rect 3185 -1994 3353 -1982
rect 3368 -1992 3384 -1978
rect 3419 -1991 3441 -1972
rect 3451 -1978 3467 -1977
rect 3450 -1984 3467 -1978
rect 3451 -1985 3467 -1984
rect 3441 -1992 3447 -1991
rect 3450 -1992 3479 -1985
rect 3368 -1993 3479 -1992
rect 3368 -1994 3485 -1993
rect 3044 -2002 3095 -1994
rect 3142 -2002 3176 -1994
rect 3044 -2014 3069 -2002
rect 3076 -2014 3095 -2002
rect 3149 -2004 3176 -2002
rect 3185 -2004 3406 -1994
rect 3441 -1997 3447 -1994
rect 3149 -2008 3406 -2004
rect 3044 -2022 3095 -2014
rect 3142 -2022 3406 -2008
rect 3450 -2002 3485 -1994
rect 2996 -2070 3015 -2036
rect 3060 -2030 3089 -2022
rect 3060 -2036 3077 -2030
rect 3060 -2038 3094 -2036
rect 3142 -2038 3158 -2022
rect 3159 -2032 3367 -2022
rect 3368 -2032 3384 -2022
rect 3432 -2026 3447 -2011
rect 3450 -2014 3451 -2002
rect 3458 -2014 3485 -2002
rect 3450 -2022 3485 -2014
rect 3450 -2023 3479 -2022
rect 3170 -2036 3384 -2032
rect 3185 -2038 3384 -2036
rect 3419 -2036 3432 -2026
rect 3450 -2036 3467 -2023
rect 3419 -2038 3467 -2036
rect 3061 -2042 3094 -2038
rect 3057 -2044 3094 -2042
rect 3057 -2045 3124 -2044
rect 3057 -2050 3088 -2045
rect 3094 -2050 3124 -2045
rect 3057 -2054 3124 -2050
rect 3030 -2057 3124 -2054
rect 3030 -2064 3079 -2057
rect 3030 -2070 3060 -2064
rect 3079 -2069 3084 -2064
rect 2996 -2086 3076 -2070
rect 3088 -2078 3124 -2057
rect 3185 -2062 3374 -2038
rect 3419 -2039 3466 -2038
rect 3432 -2044 3466 -2039
rect 3200 -2065 3374 -2062
rect 3193 -2068 3374 -2065
rect 3402 -2045 3466 -2044
rect 2996 -2088 3015 -2086
rect 3030 -2088 3064 -2086
rect 2996 -2104 3076 -2088
rect 2996 -2110 3015 -2104
rect 2712 -2136 2815 -2126
rect 2666 -2138 2815 -2136
rect 2836 -2138 2871 -2126
rect 2505 -2140 2667 -2138
rect 2517 -2160 2536 -2140
rect 2551 -2142 2581 -2140
rect 2400 -2168 2441 -2160
rect 2523 -2164 2536 -2160
rect 2588 -2156 2667 -2140
rect 2699 -2140 2871 -2138
rect 2699 -2156 2778 -2140
rect 2785 -2142 2815 -2140
rect 2363 -2178 2392 -2168
rect 2406 -2178 2435 -2168
rect 2450 -2178 2480 -2164
rect 2523 -2178 2566 -2164
rect 2588 -2168 2778 -2156
rect 2843 -2160 2849 -2140
rect 2573 -2178 2603 -2168
rect 2604 -2178 2762 -2168
rect 2766 -2178 2796 -2168
rect 2800 -2178 2830 -2164
rect 2858 -2178 2871 -2140
rect 2943 -2126 2972 -2110
rect 2986 -2126 3015 -2110
rect 3030 -2120 3060 -2104
rect 3088 -2126 3094 -2078
rect 3097 -2084 3116 -2078
rect 3131 -2084 3161 -2076
rect 3097 -2092 3161 -2084
rect 3097 -2108 3177 -2092
rect 3193 -2099 3255 -2068
rect 3271 -2099 3333 -2068
rect 3402 -2070 3451 -2045
rect 3466 -2070 3496 -2052
rect 3365 -2084 3395 -2076
rect 3402 -2078 3512 -2070
rect 3365 -2092 3410 -2084
rect 3097 -2110 3116 -2108
rect 3131 -2110 3177 -2108
rect 3097 -2126 3177 -2110
rect 3204 -2112 3239 -2099
rect 3280 -2102 3317 -2099
rect 3280 -2104 3322 -2102
rect 3209 -2115 3239 -2112
rect 3218 -2119 3225 -2115
rect 3225 -2120 3226 -2119
rect 3184 -2126 3194 -2120
rect 2943 -2134 2978 -2126
rect 2943 -2160 2944 -2134
rect 2951 -2160 2978 -2134
rect 2886 -2178 2916 -2164
rect 2943 -2168 2978 -2160
rect 2980 -2134 3021 -2126
rect 2980 -2160 2995 -2134
rect 3002 -2160 3021 -2134
rect 3085 -2138 3116 -2126
rect 3131 -2138 3234 -2126
rect 3246 -2136 3272 -2110
rect 3287 -2115 3317 -2104
rect 3349 -2108 3411 -2092
rect 3349 -2110 3395 -2108
rect 3349 -2126 3411 -2110
rect 3423 -2126 3429 -2078
rect 3432 -2086 3512 -2078
rect 3432 -2088 3451 -2086
rect 3466 -2088 3500 -2086
rect 3432 -2103 3512 -2088
rect 3432 -2104 3518 -2103
rect 3432 -2126 3451 -2104
rect 3466 -2120 3496 -2104
rect 3524 -2110 3530 -2036
rect 3533 -2110 3552 -1966
rect 3567 -2110 3573 -1966
rect 3582 -2036 3595 -1966
rect 3647 -1970 3669 -1966
rect 3640 -1982 3657 -1978
rect 3661 -1980 3669 -1978
rect 3659 -1982 3669 -1980
rect 3640 -1992 3669 -1982
rect 3722 -1992 3738 -1978
rect 3776 -1982 3782 -1980
rect 3789 -1982 3897 -1966
rect 3904 -1982 3910 -1980
rect 3918 -1982 3933 -1966
rect 3999 -1972 4018 -1969
rect 3640 -1994 3738 -1992
rect 3765 -1994 3933 -1982
rect 3948 -1992 3964 -1978
rect 3999 -1991 4021 -1972
rect 4031 -1978 4047 -1977
rect 4030 -1984 4047 -1978
rect 4031 -1985 4047 -1984
rect 4021 -1992 4027 -1991
rect 4030 -1992 4059 -1985
rect 3948 -1993 4059 -1992
rect 3948 -1994 4065 -1993
rect 3624 -2002 3675 -1994
rect 3722 -2002 3756 -1994
rect 3624 -2014 3649 -2002
rect 3656 -2014 3675 -2002
rect 3729 -2004 3756 -2002
rect 3765 -2004 3986 -1994
rect 4021 -1997 4027 -1994
rect 3729 -2008 3986 -2004
rect 3624 -2022 3675 -2014
rect 3722 -2022 3986 -2008
rect 4030 -2002 4065 -1994
rect 3576 -2070 3595 -2036
rect 3640 -2030 3669 -2022
rect 3640 -2036 3657 -2030
rect 3640 -2038 3674 -2036
rect 3722 -2038 3738 -2022
rect 3739 -2032 3947 -2022
rect 3948 -2032 3964 -2022
rect 4012 -2026 4027 -2011
rect 4030 -2014 4031 -2002
rect 4038 -2014 4065 -2002
rect 4030 -2022 4065 -2014
rect 4030 -2023 4059 -2022
rect 3750 -2036 3964 -2032
rect 3765 -2038 3964 -2036
rect 3999 -2036 4012 -2026
rect 4030 -2036 4047 -2023
rect 3999 -2038 4047 -2036
rect 3641 -2042 3674 -2038
rect 3637 -2044 3674 -2042
rect 3637 -2045 3704 -2044
rect 3637 -2050 3668 -2045
rect 3674 -2050 3704 -2045
rect 3637 -2054 3704 -2050
rect 3610 -2057 3704 -2054
rect 3610 -2064 3659 -2057
rect 3610 -2070 3640 -2064
rect 3659 -2069 3664 -2064
rect 3576 -2086 3656 -2070
rect 3668 -2078 3704 -2057
rect 3765 -2062 3954 -2038
rect 3999 -2039 4046 -2038
rect 4012 -2044 4046 -2039
rect 4086 -2044 4102 -2042
rect 3780 -2065 3954 -2062
rect 3773 -2068 3954 -2065
rect 3982 -2045 4046 -2044
rect 3576 -2088 3595 -2086
rect 3610 -2088 3644 -2086
rect 3576 -2104 3656 -2088
rect 3576 -2110 3595 -2104
rect 3292 -2136 3395 -2126
rect 3246 -2138 3395 -2136
rect 3416 -2138 3451 -2126
rect 3085 -2140 3247 -2138
rect 3097 -2160 3116 -2140
rect 3131 -2142 3161 -2140
rect 2980 -2168 3021 -2160
rect 3103 -2164 3116 -2160
rect 3168 -2156 3247 -2140
rect 3279 -2140 3451 -2138
rect 3279 -2156 3358 -2140
rect 3365 -2142 3395 -2140
rect 2943 -2178 2972 -2168
rect 2986 -2178 3015 -2168
rect 3030 -2178 3060 -2164
rect 3103 -2178 3146 -2164
rect 3168 -2168 3358 -2156
rect 3423 -2160 3429 -2140
rect 3153 -2178 3183 -2168
rect 3184 -2178 3342 -2168
rect 3346 -2178 3376 -2168
rect 3380 -2178 3410 -2164
rect 3438 -2178 3451 -2140
rect 3523 -2126 3552 -2110
rect 3566 -2126 3595 -2110
rect 3610 -2120 3640 -2104
rect 3668 -2126 3674 -2078
rect 3677 -2084 3696 -2078
rect 3711 -2084 3741 -2076
rect 3677 -2092 3741 -2084
rect 3677 -2108 3757 -2092
rect 3773 -2099 3835 -2068
rect 3851 -2099 3913 -2068
rect 3982 -2070 4031 -2045
rect 4076 -2054 4102 -2044
rect 4046 -2070 4102 -2054
rect 3945 -2084 3975 -2076
rect 3982 -2078 4092 -2070
rect 3945 -2092 3990 -2084
rect 3677 -2110 3696 -2108
rect 3711 -2110 3757 -2108
rect 3677 -2126 3757 -2110
rect 3784 -2112 3819 -2099
rect 3860 -2102 3897 -2099
rect 3860 -2104 3902 -2102
rect 3789 -2115 3819 -2112
rect 3798 -2119 3805 -2115
rect 3805 -2120 3806 -2119
rect 3764 -2126 3774 -2120
rect 3523 -2134 3558 -2126
rect 3523 -2160 3524 -2134
rect 3531 -2160 3558 -2134
rect 3466 -2178 3496 -2164
rect 3523 -2168 3558 -2160
rect 3560 -2134 3601 -2126
rect 3560 -2160 3575 -2134
rect 3582 -2160 3601 -2134
rect 3665 -2138 3696 -2126
rect 3711 -2138 3814 -2126
rect 3826 -2136 3852 -2110
rect 3867 -2115 3897 -2104
rect 3929 -2108 3991 -2092
rect 3929 -2110 3975 -2108
rect 3929 -2126 3991 -2110
rect 4003 -2126 4009 -2078
rect 4012 -2086 4092 -2078
rect 4012 -2088 4031 -2086
rect 4046 -2088 4080 -2086
rect 4012 -2104 4092 -2088
rect 4012 -2126 4031 -2104
rect 4046 -2120 4076 -2104
rect 4104 -2110 4110 -2036
rect 4113 -2110 4132 -1966
rect 4147 -2110 4153 -1966
rect 4162 -2036 4175 -1966
rect 4227 -1970 4249 -1966
rect 4220 -1982 4237 -1978
rect 4241 -1980 4249 -1978
rect 4239 -1982 4249 -1980
rect 4220 -1992 4249 -1982
rect 4302 -1992 4318 -1978
rect 4356 -1982 4362 -1980
rect 4369 -1982 4477 -1966
rect 4484 -1982 4490 -1980
rect 4498 -1982 4513 -1966
rect 4579 -1972 4598 -1969
rect 4220 -1994 4318 -1992
rect 4345 -1994 4513 -1982
rect 4528 -1992 4544 -1978
rect 4579 -1991 4601 -1972
rect 4611 -1978 4627 -1977
rect 4610 -1984 4627 -1978
rect 4611 -1985 4627 -1984
rect 4601 -1992 4607 -1991
rect 4610 -1992 4639 -1985
rect 4528 -1993 4639 -1992
rect 4528 -1994 4645 -1993
rect 4204 -2002 4255 -1994
rect 4302 -2002 4336 -1994
rect 4204 -2014 4229 -2002
rect 4236 -2014 4255 -2002
rect 4309 -2004 4336 -2002
rect 4345 -2004 4566 -1994
rect 4601 -1997 4607 -1994
rect 4309 -2008 4566 -2004
rect 4204 -2022 4255 -2014
rect 4302 -2022 4566 -2008
rect 4610 -2002 4645 -1994
rect 4156 -2070 4175 -2036
rect 4220 -2030 4249 -2022
rect 4220 -2036 4237 -2030
rect 4220 -2038 4254 -2036
rect 4302 -2038 4318 -2022
rect 4319 -2032 4527 -2022
rect 4528 -2032 4544 -2022
rect 4592 -2026 4607 -2011
rect 4610 -2014 4611 -2002
rect 4618 -2014 4645 -2002
rect 4610 -2022 4645 -2014
rect 4610 -2023 4639 -2022
rect 4330 -2036 4544 -2032
rect 4345 -2038 4544 -2036
rect 4579 -2036 4592 -2026
rect 4610 -2036 4627 -2023
rect 4579 -2038 4627 -2036
rect 4221 -2042 4254 -2038
rect 4217 -2044 4254 -2042
rect 4217 -2045 4284 -2044
rect 4217 -2050 4248 -2045
rect 4254 -2050 4284 -2045
rect 4217 -2054 4284 -2050
rect 4190 -2057 4284 -2054
rect 4190 -2064 4239 -2057
rect 4190 -2070 4220 -2064
rect 4239 -2069 4244 -2064
rect 4156 -2086 4236 -2070
rect 4248 -2078 4284 -2057
rect 4345 -2062 4534 -2038
rect 4579 -2039 4626 -2038
rect 4592 -2044 4626 -2039
rect 4360 -2065 4534 -2062
rect 4353 -2068 4534 -2065
rect 4562 -2045 4626 -2044
rect 4156 -2088 4175 -2086
rect 4190 -2088 4224 -2086
rect 4156 -2104 4236 -2088
rect 4156 -2110 4175 -2104
rect 3872 -2136 3975 -2126
rect 3826 -2138 3975 -2136
rect 3996 -2138 4031 -2126
rect 3665 -2140 3827 -2138
rect 3677 -2160 3696 -2140
rect 3711 -2142 3741 -2140
rect 3560 -2168 3601 -2160
rect 3683 -2164 3696 -2160
rect 3748 -2156 3827 -2140
rect 3859 -2140 4031 -2138
rect 3859 -2156 3938 -2140
rect 3945 -2142 3975 -2140
rect 3523 -2178 3552 -2168
rect 3566 -2178 3595 -2168
rect 3610 -2178 3640 -2164
rect 3683 -2178 3726 -2164
rect 3748 -2168 3938 -2156
rect 4003 -2160 4009 -2140
rect 3733 -2178 3763 -2168
rect 3764 -2178 3922 -2168
rect 3926 -2178 3956 -2168
rect 3960 -2178 3990 -2164
rect 4018 -2178 4031 -2140
rect 4103 -2126 4132 -2110
rect 4146 -2126 4175 -2110
rect 4190 -2120 4220 -2104
rect 4248 -2126 4254 -2078
rect 4257 -2084 4276 -2078
rect 4291 -2084 4321 -2076
rect 4257 -2092 4321 -2084
rect 4257 -2108 4337 -2092
rect 4353 -2099 4415 -2068
rect 4431 -2099 4493 -2068
rect 4562 -2070 4611 -2045
rect 4626 -2070 4656 -2052
rect 4525 -2084 4555 -2076
rect 4562 -2078 4672 -2070
rect 4525 -2092 4570 -2084
rect 4257 -2110 4276 -2108
rect 4291 -2110 4337 -2108
rect 4257 -2126 4337 -2110
rect 4364 -2112 4399 -2099
rect 4440 -2102 4477 -2099
rect 4440 -2104 4482 -2102
rect 4369 -2115 4399 -2112
rect 4378 -2119 4385 -2115
rect 4385 -2120 4386 -2119
rect 4344 -2126 4354 -2120
rect 4103 -2134 4138 -2126
rect 4103 -2160 4104 -2134
rect 4111 -2160 4138 -2134
rect 4046 -2178 4076 -2164
rect 4103 -2168 4138 -2160
rect 4140 -2134 4181 -2126
rect 4140 -2160 4155 -2134
rect 4162 -2160 4181 -2134
rect 4245 -2138 4276 -2126
rect 4291 -2138 4394 -2126
rect 4406 -2136 4432 -2110
rect 4447 -2115 4477 -2104
rect 4509 -2108 4571 -2092
rect 4509 -2110 4555 -2108
rect 4509 -2126 4571 -2110
rect 4583 -2126 4589 -2078
rect 4592 -2086 4672 -2078
rect 4592 -2088 4611 -2086
rect 4626 -2088 4660 -2086
rect 4592 -2103 4672 -2088
rect 4592 -2104 4678 -2103
rect 4592 -2126 4611 -2104
rect 4626 -2120 4656 -2104
rect 4684 -2110 4690 -2036
rect 4693 -2110 4712 -1966
rect 4727 -2110 4733 -1966
rect 4742 -2036 4755 -1966
rect 4807 -1970 4829 -1966
rect 4800 -1982 4817 -1978
rect 4821 -1980 4829 -1978
rect 4819 -1982 4829 -1980
rect 4800 -1992 4829 -1982
rect 4882 -1992 4898 -1978
rect 4936 -1982 4942 -1980
rect 4949 -1982 5057 -1966
rect 5064 -1982 5070 -1980
rect 5078 -1982 5093 -1966
rect 5159 -1972 5178 -1969
rect 4800 -1994 4898 -1992
rect 4925 -1994 5093 -1982
rect 5108 -1992 5124 -1978
rect 5159 -1991 5181 -1972
rect 5191 -1978 5207 -1977
rect 5190 -1984 5207 -1978
rect 5191 -1985 5207 -1984
rect 5181 -1992 5187 -1991
rect 5190 -1992 5219 -1985
rect 5108 -1993 5219 -1992
rect 5108 -1994 5225 -1993
rect 4784 -2002 4835 -1994
rect 4882 -2002 4916 -1994
rect 4784 -2014 4809 -2002
rect 4816 -2014 4835 -2002
rect 4889 -2004 4916 -2002
rect 4925 -2004 5146 -1994
rect 5181 -1997 5187 -1994
rect 4889 -2008 5146 -2004
rect 4784 -2022 4835 -2014
rect 4882 -2022 5146 -2008
rect 5190 -2002 5225 -1994
rect 4736 -2070 4755 -2036
rect 4800 -2030 4829 -2022
rect 4800 -2036 4817 -2030
rect 4800 -2038 4834 -2036
rect 4882 -2038 4898 -2022
rect 4899 -2032 5107 -2022
rect 5108 -2032 5124 -2022
rect 5172 -2026 5187 -2011
rect 5190 -2014 5191 -2002
rect 5198 -2014 5225 -2002
rect 5190 -2022 5225 -2014
rect 5190 -2023 5219 -2022
rect 4910 -2036 5124 -2032
rect 4925 -2038 5124 -2036
rect 5159 -2036 5172 -2026
rect 5190 -2036 5207 -2023
rect 5159 -2038 5207 -2036
rect 4801 -2042 4834 -2038
rect 4797 -2044 4834 -2042
rect 4797 -2045 4864 -2044
rect 4797 -2050 4828 -2045
rect 4834 -2050 4864 -2045
rect 4797 -2054 4864 -2050
rect 4770 -2057 4864 -2054
rect 4770 -2064 4819 -2057
rect 4770 -2070 4800 -2064
rect 4819 -2069 4824 -2064
rect 4736 -2086 4816 -2070
rect 4828 -2078 4864 -2057
rect 4925 -2062 5114 -2038
rect 5159 -2039 5206 -2038
rect 5172 -2044 5206 -2039
rect 5246 -2044 5262 -2042
rect 4940 -2065 5114 -2062
rect 4933 -2068 5114 -2065
rect 5142 -2045 5206 -2044
rect 4736 -2088 4755 -2086
rect 4770 -2088 4804 -2086
rect 4736 -2104 4816 -2088
rect 4736 -2110 4755 -2104
rect 4452 -2136 4555 -2126
rect 4406 -2138 4555 -2136
rect 4576 -2138 4611 -2126
rect 4245 -2140 4407 -2138
rect 4257 -2160 4276 -2140
rect 4291 -2142 4321 -2140
rect 4140 -2168 4181 -2160
rect 4263 -2164 4276 -2160
rect 4328 -2156 4407 -2140
rect 4439 -2140 4611 -2138
rect 4439 -2156 4518 -2140
rect 4525 -2142 4555 -2140
rect 4103 -2178 4132 -2168
rect 4146 -2178 4175 -2168
rect 4190 -2178 4220 -2164
rect 4263 -2178 4306 -2164
rect 4328 -2168 4518 -2156
rect 4583 -2160 4589 -2140
rect 4313 -2178 4343 -2168
rect 4344 -2178 4502 -2168
rect 4506 -2178 4536 -2168
rect 4540 -2178 4570 -2164
rect 4598 -2178 4611 -2140
rect 4683 -2126 4712 -2110
rect 4726 -2126 4755 -2110
rect 4770 -2120 4800 -2104
rect 4828 -2126 4834 -2078
rect 4837 -2084 4856 -2078
rect 4871 -2084 4901 -2076
rect 4837 -2092 4901 -2084
rect 4837 -2108 4917 -2092
rect 4933 -2099 4995 -2068
rect 5011 -2099 5073 -2068
rect 5142 -2070 5191 -2045
rect 5236 -2054 5262 -2044
rect 5206 -2070 5262 -2054
rect 5105 -2084 5135 -2076
rect 5142 -2078 5252 -2070
rect 5105 -2092 5150 -2084
rect 4837 -2110 4856 -2108
rect 4871 -2110 4917 -2108
rect 4837 -2126 4917 -2110
rect 4944 -2112 4979 -2099
rect 5020 -2102 5057 -2099
rect 5020 -2104 5062 -2102
rect 4949 -2115 4979 -2112
rect 4958 -2119 4965 -2115
rect 4965 -2120 4966 -2119
rect 4924 -2126 4934 -2120
rect 4683 -2134 4718 -2126
rect 4683 -2160 4684 -2134
rect 4691 -2160 4718 -2134
rect 4626 -2178 4656 -2164
rect 4683 -2168 4718 -2160
rect 4720 -2134 4761 -2126
rect 4720 -2160 4735 -2134
rect 4742 -2160 4761 -2134
rect 4825 -2138 4856 -2126
rect 4871 -2138 4974 -2126
rect 4986 -2136 5012 -2110
rect 5027 -2115 5057 -2104
rect 5089 -2108 5151 -2092
rect 5089 -2110 5135 -2108
rect 5089 -2126 5151 -2110
rect 5163 -2126 5169 -2078
rect 5172 -2086 5252 -2078
rect 5172 -2088 5191 -2086
rect 5206 -2088 5240 -2086
rect 5172 -2104 5252 -2088
rect 5172 -2126 5191 -2104
rect 5206 -2120 5236 -2104
rect 5264 -2110 5270 -2036
rect 5273 -2110 5292 -1966
rect 5307 -2110 5313 -1966
rect 5322 -2036 5335 -1966
rect 5387 -1970 5409 -1966
rect 5380 -1982 5397 -1978
rect 5401 -1980 5409 -1978
rect 5399 -1982 5409 -1980
rect 5380 -1992 5409 -1982
rect 5462 -1992 5478 -1978
rect 5516 -1982 5522 -1980
rect 5529 -1982 5637 -1966
rect 5644 -1982 5650 -1980
rect 5658 -1982 5673 -1966
rect 5739 -1972 5758 -1969
rect 5380 -1994 5478 -1992
rect 5505 -1994 5673 -1982
rect 5688 -1992 5704 -1978
rect 5739 -1991 5761 -1972
rect 5771 -1978 5787 -1977
rect 5770 -1984 5787 -1978
rect 5771 -1985 5787 -1984
rect 5761 -1992 5767 -1991
rect 5770 -1992 5799 -1985
rect 5688 -1993 5799 -1992
rect 5688 -1994 5805 -1993
rect 5364 -2002 5415 -1994
rect 5462 -2002 5496 -1994
rect 5364 -2014 5389 -2002
rect 5396 -2014 5415 -2002
rect 5469 -2004 5496 -2002
rect 5505 -2004 5726 -1994
rect 5761 -1997 5767 -1994
rect 5469 -2008 5726 -2004
rect 5364 -2022 5415 -2014
rect 5462 -2022 5726 -2008
rect 5770 -2002 5805 -1994
rect 5316 -2070 5335 -2036
rect 5380 -2030 5409 -2022
rect 5380 -2036 5397 -2030
rect 5380 -2038 5414 -2036
rect 5462 -2038 5478 -2022
rect 5479 -2032 5687 -2022
rect 5688 -2032 5704 -2022
rect 5752 -2026 5767 -2011
rect 5770 -2014 5771 -2002
rect 5778 -2014 5805 -2002
rect 5770 -2022 5805 -2014
rect 5770 -2023 5799 -2022
rect 5490 -2036 5704 -2032
rect 5505 -2038 5704 -2036
rect 5739 -2036 5752 -2026
rect 5770 -2036 5787 -2023
rect 5739 -2038 5787 -2036
rect 5381 -2042 5414 -2038
rect 5377 -2044 5414 -2042
rect 5377 -2045 5444 -2044
rect 5377 -2050 5408 -2045
rect 5414 -2050 5444 -2045
rect 5377 -2054 5444 -2050
rect 5350 -2057 5444 -2054
rect 5350 -2064 5399 -2057
rect 5350 -2070 5380 -2064
rect 5399 -2069 5404 -2064
rect 5316 -2086 5396 -2070
rect 5408 -2078 5444 -2057
rect 5505 -2062 5694 -2038
rect 5739 -2039 5786 -2038
rect 5752 -2044 5786 -2039
rect 5520 -2065 5694 -2062
rect 5513 -2068 5694 -2065
rect 5722 -2045 5786 -2044
rect 5316 -2088 5335 -2086
rect 5350 -2088 5384 -2086
rect 5316 -2104 5396 -2088
rect 5316 -2110 5335 -2104
rect 5032 -2136 5135 -2126
rect 4986 -2138 5135 -2136
rect 5156 -2138 5191 -2126
rect 4825 -2140 4987 -2138
rect 4837 -2160 4856 -2140
rect 4871 -2142 4901 -2140
rect 4720 -2168 4761 -2160
rect 4843 -2164 4856 -2160
rect 4908 -2156 4987 -2140
rect 5019 -2140 5191 -2138
rect 5019 -2156 5098 -2140
rect 5105 -2142 5135 -2140
rect 4683 -2178 4712 -2168
rect 4726 -2178 4755 -2168
rect 4770 -2178 4800 -2164
rect 4843 -2178 4886 -2164
rect 4908 -2168 5098 -2156
rect 5163 -2160 5169 -2140
rect 4893 -2178 4923 -2168
rect 4924 -2178 5082 -2168
rect 5086 -2178 5116 -2168
rect 5120 -2178 5150 -2164
rect 5178 -2178 5191 -2140
rect 5263 -2126 5292 -2110
rect 5306 -2126 5335 -2110
rect 5350 -2120 5380 -2104
rect 5408 -2126 5414 -2078
rect 5417 -2084 5436 -2078
rect 5451 -2084 5481 -2076
rect 5417 -2092 5481 -2084
rect 5417 -2108 5497 -2092
rect 5513 -2099 5575 -2068
rect 5591 -2099 5653 -2068
rect 5722 -2070 5771 -2045
rect 5786 -2070 5816 -2052
rect 5685 -2084 5715 -2076
rect 5722 -2078 5832 -2070
rect 5685 -2092 5730 -2084
rect 5417 -2110 5436 -2108
rect 5451 -2110 5497 -2108
rect 5417 -2126 5497 -2110
rect 5524 -2112 5559 -2099
rect 5600 -2102 5637 -2099
rect 5600 -2104 5642 -2102
rect 5529 -2115 5559 -2112
rect 5538 -2119 5545 -2115
rect 5545 -2120 5546 -2119
rect 5504 -2126 5514 -2120
rect 5263 -2134 5298 -2126
rect 5263 -2160 5264 -2134
rect 5271 -2160 5298 -2134
rect 5206 -2178 5236 -2164
rect 5263 -2168 5298 -2160
rect 5300 -2134 5341 -2126
rect 5300 -2160 5315 -2134
rect 5322 -2160 5341 -2134
rect 5405 -2138 5436 -2126
rect 5451 -2138 5554 -2126
rect 5566 -2136 5592 -2110
rect 5607 -2115 5637 -2104
rect 5669 -2108 5731 -2092
rect 5669 -2110 5715 -2108
rect 5669 -2126 5731 -2110
rect 5743 -2126 5749 -2078
rect 5752 -2086 5832 -2078
rect 5752 -2088 5771 -2086
rect 5786 -2088 5820 -2086
rect 5752 -2103 5832 -2088
rect 5752 -2104 5838 -2103
rect 5752 -2126 5771 -2104
rect 5786 -2120 5816 -2104
rect 5844 -2110 5850 -2036
rect 5853 -2110 5872 -1966
rect 5887 -2110 5893 -1966
rect 5902 -2036 5915 -1966
rect 5967 -1970 5989 -1966
rect 5960 -1982 5977 -1978
rect 5981 -1980 5989 -1978
rect 5979 -1982 5989 -1980
rect 5960 -1992 5989 -1982
rect 6042 -1992 6058 -1978
rect 6096 -1982 6102 -1980
rect 6109 -1982 6217 -1966
rect 6224 -1982 6230 -1980
rect 6238 -1982 6253 -1966
rect 6319 -1972 6338 -1969
rect 5960 -1994 6058 -1992
rect 6085 -1994 6253 -1982
rect 6268 -1992 6284 -1978
rect 6319 -1991 6341 -1972
rect 6351 -1978 6367 -1977
rect 6350 -1984 6367 -1978
rect 6351 -1985 6367 -1984
rect 6341 -1992 6347 -1991
rect 6350 -1992 6379 -1985
rect 6268 -1993 6379 -1992
rect 6268 -1994 6385 -1993
rect 5944 -2002 5995 -1994
rect 6042 -2002 6076 -1994
rect 5944 -2014 5969 -2002
rect 5976 -2014 5995 -2002
rect 6049 -2004 6076 -2002
rect 6085 -2004 6306 -1994
rect 6341 -1997 6347 -1994
rect 6049 -2008 6306 -2004
rect 5944 -2022 5995 -2014
rect 6042 -2022 6306 -2008
rect 6350 -2002 6385 -1994
rect 5896 -2070 5915 -2036
rect 5960 -2030 5989 -2022
rect 5960 -2036 5977 -2030
rect 5960 -2038 5994 -2036
rect 6042 -2038 6058 -2022
rect 6059 -2032 6267 -2022
rect 6268 -2032 6284 -2022
rect 6332 -2026 6347 -2011
rect 6350 -2014 6351 -2002
rect 6358 -2014 6385 -2002
rect 6350 -2022 6385 -2014
rect 6350 -2023 6379 -2022
rect 6070 -2036 6284 -2032
rect 6085 -2038 6284 -2036
rect 6319 -2036 6332 -2026
rect 6350 -2036 6367 -2023
rect 6319 -2038 6367 -2036
rect 5961 -2042 5994 -2038
rect 5957 -2044 5994 -2042
rect 5957 -2045 6024 -2044
rect 5957 -2050 5988 -2045
rect 5994 -2050 6024 -2045
rect 5957 -2054 6024 -2050
rect 5930 -2057 6024 -2054
rect 5930 -2064 5979 -2057
rect 5930 -2070 5960 -2064
rect 5979 -2069 5984 -2064
rect 5896 -2086 5976 -2070
rect 5988 -2078 6024 -2057
rect 6085 -2062 6274 -2038
rect 6319 -2039 6366 -2038
rect 6332 -2044 6366 -2039
rect 6100 -2065 6274 -2062
rect 6093 -2068 6274 -2065
rect 6302 -2045 6366 -2044
rect 5896 -2088 5915 -2086
rect 5930 -2088 5964 -2086
rect 5896 -2104 5976 -2088
rect 5896 -2110 5915 -2104
rect 5612 -2136 5715 -2126
rect 5566 -2138 5715 -2136
rect 5736 -2138 5771 -2126
rect 5405 -2140 5567 -2138
rect 5417 -2160 5436 -2140
rect 5451 -2142 5481 -2140
rect 5300 -2168 5341 -2160
rect 5423 -2164 5436 -2160
rect 5488 -2156 5567 -2140
rect 5599 -2140 5771 -2138
rect 5599 -2156 5678 -2140
rect 5685 -2142 5715 -2140
rect 5263 -2178 5292 -2168
rect 5306 -2178 5335 -2168
rect 5350 -2178 5380 -2164
rect 5423 -2178 5466 -2164
rect 5488 -2168 5678 -2156
rect 5743 -2160 5749 -2140
rect 5473 -2178 5503 -2168
rect 5504 -2178 5662 -2168
rect 5666 -2178 5696 -2168
rect 5700 -2178 5730 -2164
rect 5758 -2178 5771 -2140
rect 5843 -2126 5872 -2110
rect 5886 -2126 5915 -2110
rect 5930 -2120 5960 -2104
rect 5988 -2126 5994 -2078
rect 5997 -2084 6016 -2078
rect 6031 -2084 6061 -2076
rect 5997 -2092 6061 -2084
rect 5997 -2108 6077 -2092
rect 6093 -2099 6155 -2068
rect 6171 -2099 6233 -2068
rect 6302 -2070 6351 -2045
rect 6366 -2070 6396 -2054
rect 6265 -2084 6295 -2076
rect 6302 -2078 6412 -2070
rect 6265 -2092 6310 -2084
rect 5997 -2110 6016 -2108
rect 6031 -2110 6077 -2108
rect 5997 -2126 6077 -2110
rect 6104 -2112 6139 -2099
rect 6180 -2102 6217 -2099
rect 6180 -2104 6222 -2102
rect 6109 -2115 6139 -2112
rect 6118 -2119 6125 -2115
rect 6125 -2120 6126 -2119
rect 6084 -2126 6094 -2120
rect 5843 -2134 5878 -2126
rect 5843 -2160 5844 -2134
rect 5851 -2160 5878 -2134
rect 5786 -2178 5816 -2164
rect 5843 -2168 5878 -2160
rect 5880 -2134 5921 -2126
rect 5880 -2160 5895 -2134
rect 5902 -2160 5921 -2134
rect 5985 -2138 6016 -2126
rect 6031 -2138 6134 -2126
rect 6146 -2136 6172 -2110
rect 6187 -2115 6217 -2104
rect 6249 -2108 6311 -2092
rect 6249 -2110 6295 -2108
rect 6249 -2126 6311 -2110
rect 6323 -2126 6329 -2078
rect 6332 -2086 6412 -2078
rect 6332 -2088 6351 -2086
rect 6366 -2088 6400 -2086
rect 6332 -2104 6412 -2088
rect 6332 -2126 6351 -2104
rect 6366 -2120 6396 -2104
rect 6424 -2110 6430 -2036
rect 6439 -2110 6452 -1966
rect 6192 -2136 6295 -2126
rect 6146 -2138 6295 -2136
rect 6316 -2138 6351 -2126
rect 5985 -2140 6147 -2138
rect 5997 -2160 6016 -2140
rect 6031 -2142 6061 -2140
rect 5880 -2168 5921 -2160
rect 6003 -2164 6016 -2160
rect 6068 -2156 6147 -2140
rect 6179 -2140 6351 -2138
rect 6179 -2156 6258 -2140
rect 6265 -2142 6295 -2140
rect 5843 -2178 5872 -2168
rect 5886 -2178 5915 -2168
rect 5930 -2178 5960 -2164
rect 6003 -2178 6046 -2164
rect 6068 -2168 6258 -2156
rect 6323 -2160 6329 -2140
rect 6053 -2178 6083 -2168
rect 6084 -2178 6242 -2168
rect 6246 -2178 6276 -2168
rect 6280 -2178 6310 -2164
rect 6338 -2178 6351 -2140
rect 6423 -2126 6452 -2110
rect 6423 -2134 6458 -2126
rect 6423 -2160 6424 -2134
rect 6431 -2160 6458 -2134
rect 6366 -2178 6396 -2164
rect 6423 -2168 6458 -2160
rect 6423 -2178 6452 -2168
rect -541 -2192 6452 -2178
rect -478 -2222 -465 -2192
rect -450 -2206 -420 -2192
rect -377 -2206 -334 -2192
rect -327 -2206 -107 -2192
rect -100 -2206 -70 -2192
rect -410 -2220 -395 -2208
rect -376 -2220 -363 -2206
rect -295 -2210 -142 -2206
rect -413 -2222 -391 -2220
rect -313 -2222 -121 -2210
rect -42 -2222 -29 -2192
rect -14 -2206 16 -2192
rect 53 -2222 72 -2192
rect 87 -2222 93 -2192
rect 102 -2222 115 -2192
rect 130 -2206 160 -2192
rect 203 -2206 246 -2192
rect 253 -2206 473 -2192
rect 480 -2206 510 -2192
rect 170 -2220 185 -2208
rect 204 -2220 217 -2206
rect 285 -2210 438 -2206
rect 167 -2222 189 -2220
rect 267 -2222 459 -2210
rect 538 -2222 551 -2192
rect 566 -2206 596 -2192
rect 633 -2222 652 -2192
rect 667 -2222 673 -2192
rect 682 -2222 695 -2192
rect 710 -2206 740 -2192
rect 783 -2206 826 -2192
rect 833 -2206 1053 -2192
rect 1060 -2206 1090 -2192
rect 750 -2220 765 -2208
rect 784 -2220 797 -2206
rect 865 -2210 1018 -2206
rect 747 -2222 769 -2220
rect 847 -2222 1039 -2210
rect 1118 -2222 1131 -2192
rect 1146 -2206 1176 -2192
rect 1213 -2222 1232 -2192
rect 1247 -2222 1253 -2192
rect 1262 -2222 1275 -2192
rect 1290 -2206 1320 -2192
rect 1363 -2206 1406 -2192
rect 1413 -2206 1633 -2192
rect 1640 -2206 1670 -2192
rect 1330 -2220 1345 -2208
rect 1364 -2220 1377 -2206
rect 1445 -2210 1598 -2206
rect 1327 -2222 1349 -2220
rect 1427 -2222 1619 -2210
rect 1698 -2222 1711 -2192
rect 1726 -2206 1756 -2192
rect 1793 -2222 1812 -2192
rect 1827 -2222 1833 -2192
rect 1842 -2222 1855 -2192
rect 1870 -2206 1900 -2192
rect 1943 -2206 1986 -2192
rect 1993 -2206 2213 -2192
rect 2220 -2206 2250 -2192
rect 1910 -2220 1925 -2208
rect 1944 -2220 1957 -2206
rect 2025 -2210 2178 -2206
rect 1907 -2222 1929 -2220
rect 2007 -2222 2199 -2210
rect 2278 -2222 2291 -2192
rect 2306 -2206 2336 -2192
rect 2373 -2222 2392 -2192
rect 2407 -2222 2413 -2192
rect 2422 -2222 2435 -2192
rect 2450 -2206 2480 -2192
rect 2523 -2206 2566 -2192
rect 2573 -2206 2793 -2192
rect 2800 -2206 2830 -2192
rect 2490 -2220 2505 -2208
rect 2524 -2220 2537 -2206
rect 2605 -2210 2758 -2206
rect 2487 -2222 2509 -2220
rect 2587 -2222 2779 -2210
rect 2858 -2222 2871 -2192
rect 2886 -2206 2916 -2192
rect 2953 -2222 2972 -2192
rect 2987 -2222 2993 -2192
rect 3002 -2222 3015 -2192
rect 3030 -2206 3060 -2192
rect 3103 -2206 3146 -2192
rect 3153 -2206 3373 -2192
rect 3380 -2206 3410 -2192
rect 3070 -2220 3085 -2208
rect 3104 -2220 3117 -2206
rect 3185 -2210 3338 -2206
rect 3067 -2222 3089 -2220
rect 3167 -2222 3359 -2210
rect 3438 -2222 3451 -2192
rect 3466 -2206 3496 -2192
rect 3533 -2222 3552 -2192
rect 3567 -2222 3573 -2192
rect 3582 -2222 3595 -2192
rect 3610 -2206 3640 -2192
rect 3683 -2206 3726 -2192
rect 3733 -2206 3953 -2192
rect 3960 -2206 3990 -2192
rect 3650 -2220 3665 -2208
rect 3684 -2220 3697 -2206
rect 3765 -2210 3918 -2206
rect 3647 -2222 3669 -2220
rect 3747 -2222 3939 -2210
rect 4018 -2222 4031 -2192
rect 4046 -2206 4076 -2192
rect 4113 -2222 4132 -2192
rect 4147 -2222 4153 -2192
rect 4162 -2222 4175 -2192
rect 4190 -2206 4220 -2192
rect 4263 -2206 4306 -2192
rect 4313 -2206 4533 -2192
rect 4540 -2206 4570 -2192
rect 4230 -2220 4245 -2208
rect 4264 -2220 4277 -2206
rect 4345 -2210 4498 -2206
rect 4227 -2222 4249 -2220
rect 4327 -2222 4519 -2210
rect 4598 -2222 4611 -2192
rect 4626 -2206 4656 -2192
rect 4693 -2222 4712 -2192
rect 4727 -2222 4733 -2192
rect 4742 -2222 4755 -2192
rect 4770 -2206 4800 -2192
rect 4843 -2206 4886 -2192
rect 4893 -2206 5113 -2192
rect 5120 -2206 5150 -2192
rect 4810 -2220 4825 -2208
rect 4844 -2220 4857 -2206
rect 4925 -2210 5078 -2206
rect 4807 -2222 4829 -2220
rect 4907 -2222 5099 -2210
rect 5178 -2222 5191 -2192
rect 5206 -2206 5236 -2192
rect 5273 -2222 5292 -2192
rect 5307 -2222 5313 -2192
rect 5322 -2222 5335 -2192
rect 5350 -2206 5380 -2192
rect 5423 -2206 5466 -2192
rect 5473 -2206 5693 -2192
rect 5700 -2206 5730 -2192
rect 5390 -2220 5405 -2208
rect 5424 -2220 5437 -2206
rect 5505 -2210 5658 -2206
rect 5387 -2222 5409 -2220
rect 5487 -2222 5679 -2210
rect 5758 -2222 5771 -2192
rect 5786 -2206 5816 -2192
rect 5853 -2222 5872 -2192
rect 5887 -2222 5893 -2192
rect 5902 -2222 5915 -2192
rect 5930 -2206 5960 -2192
rect 6003 -2206 6046 -2192
rect 6053 -2206 6273 -2192
rect 6280 -2206 6310 -2192
rect 5970 -2220 5985 -2208
rect 6004 -2220 6017 -2206
rect 6085 -2210 6238 -2206
rect 5967 -2222 5989 -2220
rect 6067 -2222 6259 -2210
rect 6338 -2222 6351 -2192
rect 6366 -2206 6396 -2192
rect 6439 -2222 6452 -2192
rect -541 -2236 6452 -2222
rect -478 -2306 -465 -2236
rect -413 -2240 -391 -2236
rect -420 -2252 -403 -2248
rect -399 -2250 -391 -2248
rect -401 -2252 -391 -2250
rect -420 -2262 -391 -2252
rect -338 -2262 -322 -2248
rect -284 -2258 -278 -2250
rect -271 -2252 -163 -2236
rect -420 -2264 -322 -2262
rect -436 -2272 -385 -2264
rect -338 -2272 -304 -2264
rect -436 -2284 -411 -2272
rect -404 -2284 -385 -2272
rect -331 -2274 -304 -2272
rect -295 -2272 -278 -2258
rect -233 -2272 -201 -2252
rect -156 -2258 -150 -2250
rect -142 -2258 -127 -2236
rect -61 -2242 -42 -2239
rect -156 -2264 -127 -2258
rect -112 -2262 -96 -2248
rect -61 -2261 -39 -2242
rect -29 -2248 -13 -2247
rect -30 -2250 -13 -2248
rect -29 -2255 -13 -2250
rect -39 -2262 -33 -2261
rect -30 -2262 -1 -2255
rect -112 -2263 -1 -2262
rect -112 -2264 5 -2263
rect -156 -2272 -74 -2264
rect -39 -2267 -33 -2264
rect -295 -2274 -74 -2272
rect -331 -2278 -259 -2274
rect -231 -2276 -203 -2274
rect -178 -2278 -74 -2274
rect -436 -2292 -385 -2284
rect -338 -2286 -206 -2278
rect -201 -2286 -74 -2278
rect -30 -2272 5 -2264
rect -338 -2288 -259 -2286
rect -178 -2288 -74 -2286
rect -338 -2292 -241 -2288
rect -484 -2340 -465 -2306
rect -420 -2300 -391 -2292
rect -420 -2306 -403 -2300
rect -420 -2308 -386 -2306
rect -338 -2308 -322 -2292
rect -321 -2296 -241 -2292
rect -193 -2292 -74 -2288
rect -193 -2296 -113 -2292
rect -321 -2302 -113 -2296
rect -112 -2302 -96 -2292
rect -48 -2296 -33 -2281
rect -30 -2284 -29 -2272
rect -22 -2284 5 -2272
rect -30 -2292 5 -2284
rect -30 -2293 -1 -2292
rect -310 -2306 -206 -2302
rect -419 -2312 -386 -2308
rect -423 -2314 -386 -2312
rect -423 -2315 -356 -2314
rect -423 -2320 -392 -2315
rect -386 -2320 -356 -2315
rect -295 -2318 -280 -2306
rect -423 -2324 -356 -2320
rect -450 -2327 -356 -2324
rect -450 -2334 -401 -2327
rect -450 -2340 -420 -2334
rect -401 -2339 -396 -2334
rect -484 -2356 -404 -2340
rect -392 -2348 -356 -2327
rect -271 -2328 -241 -2319
rect -218 -2324 -200 -2306
rect -142 -2308 -96 -2302
rect -61 -2306 -48 -2296
rect -30 -2306 -13 -2293
rect -61 -2308 -13 -2306
rect -180 -2314 -178 -2312
rect -178 -2319 -166 -2314
rect -193 -2326 -163 -2319
rect -193 -2328 -162 -2326
rect -142 -2328 -106 -2308
rect -61 -2309 -14 -2308
rect -48 -2314 -14 -2309
rect -295 -2332 -106 -2328
rect -280 -2335 -106 -2332
rect -287 -2338 -106 -2335
rect -78 -2315 -14 -2314
rect -484 -2358 -465 -2356
rect -450 -2358 -416 -2356
rect -484 -2374 -404 -2358
rect -484 -2380 -465 -2374
rect -494 -2396 -465 -2380
rect -450 -2390 -420 -2374
rect -392 -2396 -386 -2348
rect -383 -2354 -364 -2348
rect -349 -2354 -319 -2346
rect -383 -2362 -319 -2354
rect -383 -2378 -303 -2362
rect -287 -2369 -225 -2338
rect -209 -2369 -147 -2338
rect -78 -2340 -29 -2315
rect -14 -2340 16 -2322
rect -115 -2354 -85 -2346
rect -78 -2348 32 -2340
rect -115 -2362 -70 -2354
rect -383 -2380 -364 -2378
rect -349 -2380 -303 -2378
rect -383 -2396 -303 -2380
rect -276 -2382 -241 -2369
rect -200 -2372 -163 -2369
rect -200 -2374 -158 -2372
rect -271 -2385 -241 -2382
rect -262 -2389 -255 -2385
rect -255 -2390 -254 -2389
rect -296 -2396 -286 -2390
rect -500 -2404 -459 -2396
rect -500 -2430 -485 -2404
rect -478 -2430 -459 -2404
rect -395 -2408 -364 -2396
rect -349 -2408 -246 -2396
rect -234 -2406 -208 -2380
rect -193 -2385 -163 -2374
rect -131 -2378 -69 -2362
rect -131 -2380 -85 -2378
rect -131 -2396 -69 -2380
rect -57 -2396 -51 -2348
rect -48 -2356 32 -2348
rect -48 -2358 -29 -2356
rect -14 -2358 20 -2356
rect -48 -2373 32 -2358
rect -48 -2374 38 -2373
rect -48 -2396 -29 -2374
rect -14 -2390 16 -2374
rect 44 -2380 50 -2306
rect 53 -2380 72 -2236
rect 87 -2380 93 -2236
rect 102 -2306 115 -2236
rect 167 -2240 189 -2236
rect 160 -2252 177 -2248
rect 181 -2250 189 -2248
rect 179 -2252 189 -2250
rect 160 -2262 189 -2252
rect 242 -2262 258 -2248
rect 296 -2258 302 -2250
rect 309 -2252 417 -2236
rect 160 -2264 258 -2262
rect 144 -2272 195 -2264
rect 242 -2272 276 -2264
rect 144 -2284 169 -2272
rect 176 -2284 195 -2272
rect 249 -2274 276 -2272
rect 285 -2272 302 -2258
rect 347 -2272 379 -2252
rect 424 -2258 430 -2250
rect 438 -2258 453 -2236
rect 519 -2242 538 -2239
rect 424 -2264 453 -2258
rect 468 -2262 484 -2248
rect 519 -2261 541 -2242
rect 551 -2248 567 -2247
rect 550 -2250 567 -2248
rect 551 -2255 567 -2250
rect 541 -2262 547 -2261
rect 550 -2262 579 -2255
rect 468 -2263 579 -2262
rect 468 -2264 585 -2263
rect 424 -2272 506 -2264
rect 541 -2267 547 -2264
rect 285 -2274 506 -2272
rect 249 -2278 321 -2274
rect 349 -2276 377 -2274
rect 402 -2278 506 -2274
rect 144 -2292 195 -2284
rect 242 -2286 374 -2278
rect 379 -2286 506 -2278
rect 550 -2272 585 -2264
rect 242 -2288 321 -2286
rect 402 -2288 506 -2286
rect 242 -2292 339 -2288
rect 96 -2340 115 -2306
rect 160 -2300 189 -2292
rect 160 -2306 177 -2300
rect 160 -2308 194 -2306
rect 242 -2308 258 -2292
rect 259 -2296 339 -2292
rect 387 -2292 506 -2288
rect 387 -2296 467 -2292
rect 259 -2302 467 -2296
rect 468 -2302 484 -2292
rect 532 -2296 547 -2281
rect 550 -2284 551 -2272
rect 558 -2284 585 -2272
rect 550 -2292 585 -2284
rect 550 -2293 579 -2292
rect 270 -2306 374 -2302
rect 161 -2312 194 -2308
rect 157 -2314 194 -2312
rect 157 -2315 224 -2314
rect 157 -2320 188 -2315
rect 194 -2320 224 -2315
rect 285 -2318 300 -2306
rect 157 -2324 224 -2320
rect 130 -2327 224 -2324
rect 130 -2334 179 -2327
rect 130 -2340 160 -2334
rect 179 -2339 184 -2334
rect 96 -2356 176 -2340
rect 188 -2348 224 -2327
rect 309 -2328 339 -2319
rect 362 -2324 380 -2306
rect 438 -2308 484 -2302
rect 519 -2306 532 -2296
rect 550 -2306 567 -2293
rect 519 -2308 567 -2306
rect 400 -2314 402 -2312
rect 402 -2319 414 -2314
rect 387 -2326 417 -2319
rect 387 -2328 418 -2326
rect 438 -2328 474 -2308
rect 519 -2309 566 -2308
rect 532 -2314 566 -2309
rect 606 -2314 622 -2312
rect 285 -2332 474 -2328
rect 300 -2335 474 -2332
rect 293 -2338 474 -2335
rect 502 -2315 566 -2314
rect 96 -2358 115 -2356
rect 130 -2358 164 -2356
rect 96 -2374 176 -2358
rect 96 -2380 115 -2374
rect -188 -2406 -85 -2396
rect -234 -2408 -85 -2406
rect -64 -2408 -29 -2396
rect -395 -2410 -233 -2408
rect -383 -2430 -364 -2410
rect -349 -2412 -319 -2410
rect -500 -2438 -459 -2430
rect -494 -2448 -465 -2438
rect -377 -2448 -364 -2430
rect -312 -2426 -233 -2410
rect -201 -2410 -29 -2408
rect -201 -2426 -122 -2410
rect -115 -2412 -85 -2410
rect -312 -2438 -122 -2426
rect -57 -2430 -51 -2410
rect -327 -2448 -319 -2438
rect -300 -2446 -297 -2438
rect -296 -2446 -278 -2438
rect -233 -2446 -201 -2438
rect -156 -2446 -138 -2438
rect -300 -2448 -134 -2446
rect -115 -2448 -104 -2438
rect -42 -2448 -29 -2410
rect 43 -2396 72 -2380
rect 86 -2396 115 -2380
rect 130 -2390 160 -2374
rect 188 -2396 194 -2348
rect 197 -2354 216 -2348
rect 231 -2354 261 -2346
rect 197 -2362 261 -2354
rect 197 -2378 277 -2362
rect 293 -2369 355 -2338
rect 371 -2369 433 -2338
rect 502 -2340 551 -2315
rect 596 -2324 622 -2314
rect 566 -2340 622 -2324
rect 465 -2354 495 -2346
rect 502 -2348 612 -2340
rect 465 -2362 510 -2354
rect 197 -2380 216 -2378
rect 231 -2380 277 -2378
rect 197 -2396 277 -2380
rect 304 -2382 339 -2369
rect 380 -2372 417 -2369
rect 380 -2374 422 -2372
rect 309 -2385 339 -2382
rect 318 -2389 325 -2385
rect 325 -2390 326 -2389
rect 284 -2396 294 -2390
rect 43 -2404 78 -2396
rect 43 -2430 44 -2404
rect 51 -2430 78 -2404
rect 43 -2438 78 -2430
rect 80 -2404 121 -2396
rect 80 -2430 95 -2404
rect 102 -2430 121 -2404
rect 185 -2408 216 -2396
rect 231 -2408 334 -2396
rect 346 -2406 372 -2380
rect 387 -2385 417 -2374
rect 449 -2378 511 -2362
rect 449 -2380 495 -2378
rect 449 -2396 511 -2380
rect 523 -2396 529 -2348
rect 532 -2356 612 -2348
rect 532 -2358 551 -2356
rect 566 -2358 600 -2356
rect 532 -2374 612 -2358
rect 532 -2396 551 -2374
rect 566 -2390 596 -2374
rect 624 -2380 630 -2306
rect 633 -2380 652 -2236
rect 667 -2380 673 -2236
rect 682 -2306 695 -2236
rect 747 -2240 769 -2236
rect 740 -2252 757 -2248
rect 761 -2250 769 -2248
rect 759 -2252 769 -2250
rect 740 -2262 769 -2252
rect 822 -2262 838 -2248
rect 876 -2258 882 -2250
rect 889 -2252 997 -2236
rect 740 -2264 838 -2262
rect 724 -2272 775 -2264
rect 822 -2272 856 -2264
rect 724 -2284 749 -2272
rect 756 -2284 775 -2272
rect 829 -2274 856 -2272
rect 865 -2272 882 -2258
rect 927 -2272 959 -2252
rect 1004 -2258 1010 -2250
rect 1018 -2258 1033 -2236
rect 1099 -2242 1118 -2239
rect 1004 -2264 1033 -2258
rect 1048 -2262 1064 -2248
rect 1099 -2261 1121 -2242
rect 1131 -2248 1147 -2247
rect 1130 -2250 1147 -2248
rect 1131 -2255 1147 -2250
rect 1121 -2262 1127 -2261
rect 1130 -2262 1159 -2255
rect 1048 -2263 1159 -2262
rect 1048 -2264 1165 -2263
rect 1004 -2272 1086 -2264
rect 1121 -2267 1127 -2264
rect 865 -2274 1086 -2272
rect 829 -2278 901 -2274
rect 929 -2276 957 -2274
rect 982 -2278 1086 -2274
rect 724 -2292 775 -2284
rect 822 -2286 954 -2278
rect 959 -2286 1086 -2278
rect 1130 -2272 1165 -2264
rect 822 -2288 901 -2286
rect 982 -2288 1086 -2286
rect 822 -2292 919 -2288
rect 676 -2340 695 -2306
rect 740 -2300 769 -2292
rect 740 -2306 757 -2300
rect 740 -2308 774 -2306
rect 822 -2308 838 -2292
rect 839 -2296 919 -2292
rect 967 -2292 1086 -2288
rect 967 -2296 1047 -2292
rect 839 -2302 1047 -2296
rect 1048 -2302 1064 -2292
rect 1112 -2296 1127 -2281
rect 1130 -2284 1131 -2272
rect 1138 -2284 1165 -2272
rect 1130 -2292 1165 -2284
rect 1130 -2293 1159 -2292
rect 850 -2306 954 -2302
rect 741 -2312 774 -2308
rect 737 -2314 774 -2312
rect 737 -2315 804 -2314
rect 737 -2320 768 -2315
rect 774 -2320 804 -2315
rect 865 -2318 880 -2306
rect 737 -2324 804 -2320
rect 710 -2327 804 -2324
rect 710 -2334 759 -2327
rect 710 -2340 740 -2334
rect 759 -2339 764 -2334
rect 676 -2356 756 -2340
rect 768 -2348 804 -2327
rect 889 -2328 919 -2319
rect 942 -2324 960 -2306
rect 1018 -2308 1064 -2302
rect 1099 -2306 1112 -2296
rect 1130 -2306 1147 -2293
rect 1099 -2308 1147 -2306
rect 980 -2314 982 -2312
rect 982 -2319 994 -2314
rect 967 -2326 997 -2319
rect 967 -2328 998 -2326
rect 1018 -2328 1054 -2308
rect 1099 -2309 1146 -2308
rect 1112 -2314 1146 -2309
rect 865 -2332 1054 -2328
rect 880 -2335 1054 -2332
rect 873 -2338 1054 -2335
rect 1082 -2315 1146 -2314
rect 676 -2358 695 -2356
rect 710 -2358 744 -2356
rect 676 -2374 756 -2358
rect 676 -2380 695 -2374
rect 392 -2406 495 -2396
rect 346 -2408 495 -2406
rect 516 -2408 551 -2396
rect 185 -2410 347 -2408
rect 197 -2430 216 -2410
rect 231 -2412 261 -2410
rect 80 -2438 121 -2430
rect 43 -2448 72 -2438
rect 86 -2448 115 -2438
rect 203 -2448 216 -2430
rect 268 -2426 347 -2410
rect 379 -2410 551 -2408
rect 379 -2426 458 -2410
rect 465 -2412 495 -2410
rect 268 -2438 458 -2426
rect 523 -2430 529 -2410
rect 253 -2448 261 -2438
rect 280 -2446 283 -2438
rect 284 -2446 302 -2438
rect 347 -2446 379 -2438
rect 424 -2446 442 -2438
rect 280 -2448 446 -2446
rect 465 -2448 476 -2438
rect 538 -2448 551 -2410
rect 623 -2396 652 -2380
rect 666 -2396 695 -2380
rect 710 -2390 740 -2374
rect 768 -2396 774 -2348
rect 777 -2354 796 -2348
rect 811 -2354 841 -2346
rect 777 -2362 841 -2354
rect 777 -2378 857 -2362
rect 873 -2369 935 -2338
rect 951 -2369 1013 -2338
rect 1082 -2340 1131 -2315
rect 1146 -2340 1176 -2322
rect 1045 -2354 1075 -2346
rect 1082 -2348 1192 -2340
rect 1045 -2362 1090 -2354
rect 777 -2380 796 -2378
rect 811 -2380 857 -2378
rect 777 -2396 857 -2380
rect 884 -2382 919 -2369
rect 960 -2372 997 -2369
rect 960 -2374 1002 -2372
rect 889 -2385 919 -2382
rect 898 -2389 905 -2385
rect 905 -2390 906 -2389
rect 864 -2396 874 -2390
rect 623 -2404 658 -2396
rect 623 -2430 624 -2404
rect 631 -2430 658 -2404
rect 623 -2438 658 -2430
rect 660 -2404 701 -2396
rect 660 -2430 675 -2404
rect 682 -2430 701 -2404
rect 765 -2408 796 -2396
rect 811 -2408 914 -2396
rect 926 -2406 952 -2380
rect 967 -2385 997 -2374
rect 1029 -2378 1091 -2362
rect 1029 -2380 1075 -2378
rect 1029 -2396 1091 -2380
rect 1103 -2396 1109 -2348
rect 1112 -2356 1192 -2348
rect 1112 -2358 1131 -2356
rect 1146 -2358 1180 -2356
rect 1112 -2373 1192 -2358
rect 1112 -2374 1198 -2373
rect 1112 -2396 1131 -2374
rect 1146 -2390 1176 -2374
rect 1204 -2380 1210 -2306
rect 1213 -2380 1232 -2236
rect 1247 -2380 1253 -2236
rect 1262 -2306 1275 -2236
rect 1327 -2240 1349 -2236
rect 1320 -2252 1337 -2248
rect 1341 -2250 1349 -2248
rect 1339 -2252 1349 -2250
rect 1320 -2262 1349 -2252
rect 1402 -2262 1418 -2248
rect 1456 -2258 1462 -2250
rect 1469 -2252 1577 -2236
rect 1320 -2264 1418 -2262
rect 1304 -2272 1355 -2264
rect 1402 -2272 1436 -2264
rect 1304 -2284 1329 -2272
rect 1336 -2284 1355 -2272
rect 1409 -2274 1436 -2272
rect 1445 -2272 1462 -2258
rect 1507 -2272 1539 -2252
rect 1584 -2258 1590 -2250
rect 1598 -2258 1613 -2236
rect 1679 -2242 1698 -2239
rect 1584 -2264 1613 -2258
rect 1628 -2262 1644 -2248
rect 1679 -2261 1701 -2242
rect 1711 -2248 1727 -2247
rect 1710 -2250 1727 -2248
rect 1711 -2255 1727 -2250
rect 1701 -2262 1707 -2261
rect 1710 -2262 1739 -2255
rect 1628 -2263 1739 -2262
rect 1628 -2264 1745 -2263
rect 1584 -2272 1666 -2264
rect 1701 -2267 1707 -2264
rect 1445 -2274 1666 -2272
rect 1409 -2278 1481 -2274
rect 1509 -2276 1537 -2274
rect 1562 -2278 1666 -2274
rect 1304 -2292 1355 -2284
rect 1402 -2286 1534 -2278
rect 1539 -2286 1666 -2278
rect 1710 -2272 1745 -2264
rect 1402 -2288 1481 -2286
rect 1562 -2288 1666 -2286
rect 1402 -2292 1499 -2288
rect 1256 -2340 1275 -2306
rect 1320 -2300 1349 -2292
rect 1320 -2306 1337 -2300
rect 1320 -2308 1354 -2306
rect 1402 -2308 1418 -2292
rect 1419 -2296 1499 -2292
rect 1547 -2292 1666 -2288
rect 1547 -2296 1627 -2292
rect 1419 -2302 1627 -2296
rect 1628 -2302 1644 -2292
rect 1692 -2296 1707 -2281
rect 1710 -2284 1711 -2272
rect 1718 -2284 1745 -2272
rect 1710 -2292 1745 -2284
rect 1710 -2293 1739 -2292
rect 1430 -2306 1534 -2302
rect 1321 -2312 1354 -2308
rect 1317 -2314 1354 -2312
rect 1317 -2315 1384 -2314
rect 1317 -2320 1348 -2315
rect 1354 -2320 1384 -2315
rect 1445 -2318 1460 -2306
rect 1317 -2324 1384 -2320
rect 1290 -2327 1384 -2324
rect 1290 -2334 1339 -2327
rect 1290 -2340 1320 -2334
rect 1339 -2339 1344 -2334
rect 1256 -2356 1336 -2340
rect 1348 -2348 1384 -2327
rect 1469 -2328 1499 -2319
rect 1522 -2324 1540 -2306
rect 1598 -2308 1644 -2302
rect 1679 -2306 1692 -2296
rect 1710 -2306 1727 -2293
rect 1679 -2308 1727 -2306
rect 1560 -2314 1562 -2312
rect 1562 -2319 1574 -2314
rect 1547 -2326 1577 -2319
rect 1547 -2328 1578 -2326
rect 1598 -2328 1634 -2308
rect 1679 -2309 1726 -2308
rect 1692 -2314 1726 -2309
rect 1766 -2314 1782 -2312
rect 1445 -2332 1634 -2328
rect 1460 -2335 1634 -2332
rect 1453 -2338 1634 -2335
rect 1662 -2315 1726 -2314
rect 1256 -2358 1275 -2356
rect 1290 -2358 1324 -2356
rect 1256 -2374 1336 -2358
rect 1256 -2380 1275 -2374
rect 972 -2406 1075 -2396
rect 926 -2408 1075 -2406
rect 1096 -2408 1131 -2396
rect 765 -2410 927 -2408
rect 777 -2430 796 -2410
rect 811 -2412 841 -2410
rect 660 -2438 701 -2430
rect 623 -2448 652 -2438
rect 666 -2448 695 -2438
rect 783 -2448 796 -2430
rect 848 -2426 927 -2410
rect 959 -2410 1131 -2408
rect 959 -2426 1038 -2410
rect 1045 -2412 1075 -2410
rect 848 -2438 1038 -2426
rect 1103 -2430 1109 -2410
rect 833 -2448 841 -2438
rect 860 -2446 863 -2438
rect 864 -2446 882 -2438
rect 927 -2446 959 -2438
rect 1004 -2446 1022 -2438
rect 860 -2448 1026 -2446
rect 1045 -2448 1056 -2438
rect 1118 -2448 1131 -2410
rect 1203 -2396 1232 -2380
rect 1246 -2396 1275 -2380
rect 1290 -2390 1320 -2374
rect 1348 -2396 1354 -2348
rect 1357 -2354 1376 -2348
rect 1391 -2354 1421 -2346
rect 1357 -2362 1421 -2354
rect 1357 -2378 1437 -2362
rect 1453 -2369 1515 -2338
rect 1531 -2369 1593 -2338
rect 1662 -2340 1711 -2315
rect 1756 -2324 1782 -2314
rect 1726 -2340 1782 -2324
rect 1625 -2354 1655 -2346
rect 1662 -2348 1772 -2340
rect 1625 -2362 1670 -2354
rect 1357 -2380 1376 -2378
rect 1391 -2380 1437 -2378
rect 1357 -2396 1437 -2380
rect 1464 -2382 1499 -2369
rect 1540 -2372 1577 -2369
rect 1540 -2374 1582 -2372
rect 1469 -2385 1499 -2382
rect 1478 -2389 1485 -2385
rect 1485 -2390 1486 -2389
rect 1444 -2396 1454 -2390
rect 1203 -2404 1238 -2396
rect 1203 -2430 1204 -2404
rect 1211 -2430 1238 -2404
rect 1203 -2438 1238 -2430
rect 1240 -2404 1281 -2396
rect 1240 -2430 1255 -2404
rect 1262 -2430 1281 -2404
rect 1345 -2408 1376 -2396
rect 1391 -2408 1494 -2396
rect 1506 -2406 1532 -2380
rect 1547 -2385 1577 -2374
rect 1609 -2378 1671 -2362
rect 1609 -2380 1655 -2378
rect 1609 -2396 1671 -2380
rect 1683 -2396 1689 -2348
rect 1692 -2356 1772 -2348
rect 1692 -2358 1711 -2356
rect 1726 -2358 1760 -2356
rect 1692 -2374 1772 -2358
rect 1692 -2396 1711 -2374
rect 1726 -2390 1756 -2374
rect 1784 -2380 1790 -2306
rect 1793 -2380 1812 -2236
rect 1827 -2380 1833 -2236
rect 1842 -2306 1855 -2236
rect 1907 -2240 1929 -2236
rect 1900 -2252 1917 -2248
rect 1921 -2250 1929 -2248
rect 1919 -2252 1929 -2250
rect 1900 -2262 1929 -2252
rect 1982 -2262 1998 -2248
rect 2036 -2258 2042 -2250
rect 2049 -2252 2157 -2236
rect 1900 -2264 1998 -2262
rect 1884 -2272 1935 -2264
rect 1982 -2272 2016 -2264
rect 1884 -2284 1909 -2272
rect 1916 -2284 1935 -2272
rect 1989 -2274 2016 -2272
rect 2025 -2272 2042 -2258
rect 2087 -2272 2119 -2252
rect 2164 -2258 2170 -2250
rect 2178 -2258 2193 -2236
rect 2259 -2242 2278 -2239
rect 2164 -2264 2193 -2258
rect 2208 -2262 2224 -2248
rect 2259 -2261 2281 -2242
rect 2291 -2248 2307 -2247
rect 2290 -2250 2307 -2248
rect 2291 -2255 2307 -2250
rect 2281 -2262 2287 -2261
rect 2290 -2262 2319 -2255
rect 2208 -2263 2319 -2262
rect 2208 -2264 2325 -2263
rect 2164 -2272 2246 -2264
rect 2281 -2267 2287 -2264
rect 2025 -2274 2246 -2272
rect 1989 -2278 2061 -2274
rect 2089 -2276 2117 -2274
rect 2142 -2278 2246 -2274
rect 1884 -2292 1935 -2284
rect 1982 -2286 2114 -2278
rect 2119 -2286 2246 -2278
rect 2290 -2272 2325 -2264
rect 1982 -2288 2061 -2286
rect 2142 -2288 2246 -2286
rect 1982 -2292 2079 -2288
rect 1836 -2340 1855 -2306
rect 1900 -2300 1929 -2292
rect 1900 -2306 1917 -2300
rect 1900 -2308 1934 -2306
rect 1982 -2308 1998 -2292
rect 1999 -2296 2079 -2292
rect 2127 -2292 2246 -2288
rect 2127 -2296 2207 -2292
rect 1999 -2302 2207 -2296
rect 2208 -2302 2224 -2292
rect 2272 -2296 2287 -2281
rect 2290 -2284 2291 -2272
rect 2298 -2284 2325 -2272
rect 2290 -2292 2325 -2284
rect 2290 -2293 2319 -2292
rect 2010 -2306 2114 -2302
rect 1901 -2312 1934 -2308
rect 1897 -2314 1934 -2312
rect 1897 -2315 1964 -2314
rect 1897 -2320 1928 -2315
rect 1934 -2320 1964 -2315
rect 2025 -2318 2040 -2306
rect 1897 -2324 1964 -2320
rect 1870 -2327 1964 -2324
rect 1870 -2334 1919 -2327
rect 1870 -2340 1900 -2334
rect 1919 -2339 1924 -2334
rect 1836 -2356 1916 -2340
rect 1928 -2348 1964 -2327
rect 2049 -2328 2079 -2319
rect 2102 -2324 2120 -2306
rect 2178 -2308 2224 -2302
rect 2259 -2306 2272 -2296
rect 2290 -2306 2307 -2293
rect 2259 -2308 2307 -2306
rect 2140 -2314 2142 -2312
rect 2142 -2319 2154 -2314
rect 2127 -2326 2157 -2319
rect 2127 -2328 2158 -2326
rect 2178 -2328 2214 -2308
rect 2259 -2309 2306 -2308
rect 2272 -2314 2306 -2309
rect 2025 -2332 2214 -2328
rect 2040 -2335 2214 -2332
rect 2033 -2338 2214 -2335
rect 2242 -2315 2306 -2314
rect 1836 -2358 1855 -2356
rect 1870 -2358 1904 -2356
rect 1836 -2374 1916 -2358
rect 1836 -2380 1855 -2374
rect 1552 -2406 1655 -2396
rect 1506 -2408 1655 -2406
rect 1676 -2408 1711 -2396
rect 1345 -2410 1507 -2408
rect 1357 -2430 1376 -2410
rect 1391 -2412 1421 -2410
rect 1240 -2438 1281 -2430
rect 1203 -2448 1232 -2438
rect 1246 -2448 1275 -2438
rect 1363 -2448 1376 -2430
rect 1428 -2426 1507 -2410
rect 1539 -2410 1711 -2408
rect 1539 -2426 1618 -2410
rect 1625 -2412 1655 -2410
rect 1428 -2438 1618 -2426
rect 1683 -2430 1689 -2410
rect 1413 -2448 1421 -2438
rect 1440 -2446 1443 -2438
rect 1444 -2446 1462 -2438
rect 1507 -2446 1539 -2438
rect 1584 -2446 1602 -2438
rect 1440 -2448 1606 -2446
rect 1625 -2448 1636 -2438
rect 1698 -2448 1711 -2410
rect 1783 -2396 1812 -2380
rect 1826 -2396 1855 -2380
rect 1870 -2390 1900 -2374
rect 1928 -2396 1934 -2348
rect 1937 -2354 1956 -2348
rect 1971 -2354 2001 -2346
rect 1937 -2362 2001 -2354
rect 1937 -2378 2017 -2362
rect 2033 -2369 2095 -2338
rect 2111 -2369 2173 -2338
rect 2242 -2340 2291 -2315
rect 2306 -2340 2336 -2322
rect 2205 -2354 2235 -2346
rect 2242 -2348 2352 -2340
rect 2205 -2362 2250 -2354
rect 1937 -2380 1956 -2378
rect 1971 -2380 2017 -2378
rect 1937 -2396 2017 -2380
rect 2044 -2382 2079 -2369
rect 2120 -2372 2157 -2369
rect 2120 -2374 2162 -2372
rect 2049 -2385 2079 -2382
rect 2058 -2389 2065 -2385
rect 2065 -2390 2066 -2389
rect 2024 -2396 2034 -2390
rect 1783 -2404 1818 -2396
rect 1783 -2430 1784 -2404
rect 1791 -2430 1818 -2404
rect 1783 -2438 1818 -2430
rect 1820 -2404 1861 -2396
rect 1820 -2430 1835 -2404
rect 1842 -2430 1861 -2404
rect 1925 -2408 1956 -2396
rect 1971 -2408 2074 -2396
rect 2086 -2406 2112 -2380
rect 2127 -2385 2157 -2374
rect 2189 -2378 2251 -2362
rect 2189 -2380 2235 -2378
rect 2189 -2396 2251 -2380
rect 2263 -2396 2269 -2348
rect 2272 -2356 2352 -2348
rect 2272 -2358 2291 -2356
rect 2306 -2358 2340 -2356
rect 2272 -2373 2352 -2358
rect 2272 -2374 2358 -2373
rect 2272 -2396 2291 -2374
rect 2306 -2390 2336 -2374
rect 2364 -2380 2370 -2306
rect 2373 -2380 2392 -2236
rect 2407 -2380 2413 -2236
rect 2422 -2306 2435 -2236
rect 2487 -2240 2509 -2236
rect 2480 -2252 2497 -2248
rect 2501 -2250 2509 -2248
rect 2499 -2252 2509 -2250
rect 2480 -2262 2509 -2252
rect 2562 -2262 2578 -2248
rect 2616 -2258 2622 -2250
rect 2629 -2252 2737 -2236
rect 2480 -2264 2578 -2262
rect 2464 -2272 2515 -2264
rect 2562 -2272 2596 -2264
rect 2464 -2284 2489 -2272
rect 2496 -2284 2515 -2272
rect 2569 -2274 2596 -2272
rect 2605 -2272 2622 -2258
rect 2667 -2272 2699 -2252
rect 2744 -2258 2750 -2250
rect 2758 -2258 2773 -2236
rect 2839 -2242 2858 -2239
rect 2744 -2264 2773 -2258
rect 2788 -2262 2804 -2248
rect 2839 -2261 2861 -2242
rect 2871 -2248 2887 -2247
rect 2870 -2250 2887 -2248
rect 2871 -2255 2887 -2250
rect 2861 -2262 2867 -2261
rect 2870 -2262 2899 -2255
rect 2788 -2263 2899 -2262
rect 2788 -2264 2905 -2263
rect 2744 -2272 2826 -2264
rect 2861 -2267 2867 -2264
rect 2605 -2274 2826 -2272
rect 2569 -2278 2641 -2274
rect 2669 -2276 2697 -2274
rect 2722 -2278 2826 -2274
rect 2464 -2292 2515 -2284
rect 2562 -2286 2694 -2278
rect 2699 -2286 2826 -2278
rect 2870 -2272 2905 -2264
rect 2562 -2288 2641 -2286
rect 2722 -2288 2826 -2286
rect 2562 -2292 2659 -2288
rect 2416 -2340 2435 -2306
rect 2480 -2300 2509 -2292
rect 2480 -2306 2497 -2300
rect 2480 -2308 2514 -2306
rect 2562 -2308 2578 -2292
rect 2579 -2296 2659 -2292
rect 2707 -2292 2826 -2288
rect 2707 -2296 2787 -2292
rect 2579 -2302 2787 -2296
rect 2788 -2302 2804 -2292
rect 2852 -2296 2867 -2281
rect 2870 -2284 2871 -2272
rect 2878 -2284 2905 -2272
rect 2870 -2292 2905 -2284
rect 2870 -2293 2899 -2292
rect 2590 -2306 2694 -2302
rect 2481 -2312 2514 -2308
rect 2477 -2314 2514 -2312
rect 2477 -2315 2544 -2314
rect 2477 -2320 2508 -2315
rect 2514 -2320 2544 -2315
rect 2605 -2318 2620 -2306
rect 2477 -2324 2544 -2320
rect 2450 -2327 2544 -2324
rect 2450 -2334 2499 -2327
rect 2450 -2340 2480 -2334
rect 2499 -2339 2504 -2334
rect 2416 -2356 2496 -2340
rect 2508 -2348 2544 -2327
rect 2629 -2328 2659 -2319
rect 2682 -2324 2700 -2306
rect 2758 -2308 2804 -2302
rect 2839 -2306 2852 -2296
rect 2870 -2306 2887 -2293
rect 2839 -2308 2887 -2306
rect 2720 -2314 2722 -2312
rect 2722 -2319 2734 -2314
rect 2707 -2326 2737 -2319
rect 2707 -2328 2738 -2326
rect 2758 -2328 2794 -2308
rect 2839 -2309 2886 -2308
rect 2852 -2314 2886 -2309
rect 2926 -2314 2942 -2312
rect 2605 -2332 2794 -2328
rect 2620 -2335 2794 -2332
rect 2613 -2338 2794 -2335
rect 2822 -2315 2886 -2314
rect 2416 -2358 2435 -2356
rect 2450 -2358 2484 -2356
rect 2416 -2374 2496 -2358
rect 2416 -2380 2435 -2374
rect 2132 -2406 2235 -2396
rect 2086 -2408 2235 -2406
rect 2256 -2408 2291 -2396
rect 1925 -2410 2087 -2408
rect 1937 -2430 1956 -2410
rect 1971 -2412 2001 -2410
rect 1820 -2438 1861 -2430
rect 1783 -2448 1812 -2438
rect 1826 -2448 1855 -2438
rect 1943 -2448 1956 -2430
rect 2008 -2426 2087 -2410
rect 2119 -2410 2291 -2408
rect 2119 -2426 2198 -2410
rect 2205 -2412 2235 -2410
rect 2008 -2438 2198 -2426
rect 2263 -2430 2269 -2410
rect 1993 -2448 2001 -2438
rect 2020 -2446 2023 -2438
rect 2024 -2446 2042 -2438
rect 2087 -2446 2119 -2438
rect 2164 -2446 2182 -2438
rect 2020 -2448 2186 -2446
rect 2205 -2448 2216 -2438
rect 2278 -2448 2291 -2410
rect 2363 -2396 2392 -2380
rect 2406 -2396 2435 -2380
rect 2450 -2390 2480 -2374
rect 2508 -2396 2514 -2348
rect 2517 -2354 2536 -2348
rect 2551 -2354 2581 -2346
rect 2517 -2362 2581 -2354
rect 2517 -2378 2597 -2362
rect 2613 -2369 2675 -2338
rect 2691 -2369 2753 -2338
rect 2822 -2340 2871 -2315
rect 2916 -2324 2942 -2314
rect 2886 -2340 2942 -2324
rect 2785 -2354 2815 -2346
rect 2822 -2348 2932 -2340
rect 2785 -2362 2830 -2354
rect 2517 -2380 2536 -2378
rect 2551 -2380 2597 -2378
rect 2517 -2396 2597 -2380
rect 2624 -2382 2659 -2369
rect 2700 -2372 2737 -2369
rect 2700 -2374 2742 -2372
rect 2629 -2385 2659 -2382
rect 2638 -2389 2645 -2385
rect 2645 -2390 2646 -2389
rect 2604 -2396 2614 -2390
rect 2363 -2404 2398 -2396
rect 2363 -2430 2364 -2404
rect 2371 -2430 2398 -2404
rect 2363 -2438 2398 -2430
rect 2400 -2404 2441 -2396
rect 2400 -2430 2415 -2404
rect 2422 -2430 2441 -2404
rect 2505 -2408 2536 -2396
rect 2551 -2408 2654 -2396
rect 2666 -2406 2692 -2380
rect 2707 -2385 2737 -2374
rect 2769 -2378 2831 -2362
rect 2769 -2380 2815 -2378
rect 2769 -2396 2831 -2380
rect 2843 -2396 2849 -2348
rect 2852 -2356 2932 -2348
rect 2852 -2358 2871 -2356
rect 2886 -2358 2920 -2356
rect 2852 -2374 2932 -2358
rect 2852 -2396 2871 -2374
rect 2886 -2390 2916 -2374
rect 2944 -2380 2950 -2306
rect 2953 -2380 2972 -2236
rect 2987 -2380 2993 -2236
rect 3002 -2306 3015 -2236
rect 3067 -2240 3089 -2236
rect 3060 -2252 3077 -2248
rect 3081 -2250 3089 -2248
rect 3079 -2252 3089 -2250
rect 3060 -2262 3089 -2252
rect 3142 -2262 3158 -2248
rect 3196 -2258 3202 -2250
rect 3209 -2252 3317 -2236
rect 3060 -2264 3158 -2262
rect 3044 -2272 3095 -2264
rect 3142 -2272 3176 -2264
rect 3044 -2284 3069 -2272
rect 3076 -2284 3095 -2272
rect 3149 -2274 3176 -2272
rect 3185 -2272 3202 -2258
rect 3247 -2272 3279 -2252
rect 3324 -2258 3330 -2250
rect 3338 -2258 3353 -2236
rect 3419 -2242 3438 -2239
rect 3324 -2264 3353 -2258
rect 3368 -2262 3384 -2248
rect 3419 -2261 3441 -2242
rect 3451 -2248 3467 -2247
rect 3450 -2250 3467 -2248
rect 3451 -2255 3467 -2250
rect 3441 -2262 3447 -2261
rect 3450 -2262 3479 -2255
rect 3368 -2263 3479 -2262
rect 3368 -2264 3485 -2263
rect 3324 -2272 3406 -2264
rect 3441 -2267 3447 -2264
rect 3185 -2274 3406 -2272
rect 3149 -2278 3221 -2274
rect 3249 -2276 3277 -2274
rect 3302 -2278 3406 -2274
rect 3044 -2292 3095 -2284
rect 3142 -2286 3274 -2278
rect 3279 -2286 3406 -2278
rect 3450 -2272 3485 -2264
rect 3142 -2288 3221 -2286
rect 3302 -2288 3406 -2286
rect 3142 -2292 3239 -2288
rect 2996 -2340 3015 -2306
rect 3060 -2300 3089 -2292
rect 3060 -2306 3077 -2300
rect 3060 -2308 3094 -2306
rect 3142 -2308 3158 -2292
rect 3159 -2296 3239 -2292
rect 3287 -2292 3406 -2288
rect 3287 -2296 3367 -2292
rect 3159 -2302 3367 -2296
rect 3368 -2302 3384 -2292
rect 3432 -2296 3447 -2281
rect 3450 -2284 3451 -2272
rect 3458 -2284 3485 -2272
rect 3450 -2292 3485 -2284
rect 3450 -2293 3479 -2292
rect 3170 -2306 3274 -2302
rect 3061 -2312 3094 -2308
rect 3057 -2314 3094 -2312
rect 3057 -2315 3124 -2314
rect 3057 -2320 3088 -2315
rect 3094 -2320 3124 -2315
rect 3185 -2318 3200 -2306
rect 3057 -2324 3124 -2320
rect 3030 -2327 3124 -2324
rect 3030 -2334 3079 -2327
rect 3030 -2340 3060 -2334
rect 3079 -2339 3084 -2334
rect 2996 -2356 3076 -2340
rect 3088 -2348 3124 -2327
rect 3209 -2328 3239 -2319
rect 3262 -2324 3280 -2306
rect 3338 -2308 3384 -2302
rect 3419 -2306 3432 -2296
rect 3450 -2306 3467 -2293
rect 3419 -2308 3467 -2306
rect 3300 -2314 3302 -2312
rect 3302 -2319 3314 -2314
rect 3287 -2326 3317 -2319
rect 3287 -2328 3318 -2326
rect 3338 -2328 3374 -2308
rect 3419 -2309 3466 -2308
rect 3432 -2314 3466 -2309
rect 3185 -2332 3374 -2328
rect 3200 -2335 3374 -2332
rect 3193 -2338 3374 -2335
rect 3402 -2315 3466 -2314
rect 2996 -2358 3015 -2356
rect 3030 -2358 3064 -2356
rect 2996 -2374 3076 -2358
rect 2996 -2380 3015 -2374
rect 2712 -2406 2815 -2396
rect 2666 -2408 2815 -2406
rect 2836 -2408 2871 -2396
rect 2505 -2410 2667 -2408
rect 2517 -2430 2536 -2410
rect 2551 -2412 2581 -2410
rect 2400 -2438 2441 -2430
rect 2363 -2448 2392 -2438
rect 2406 -2448 2435 -2438
rect 2523 -2448 2536 -2430
rect 2588 -2426 2667 -2410
rect 2699 -2410 2871 -2408
rect 2699 -2426 2778 -2410
rect 2785 -2412 2815 -2410
rect 2588 -2438 2778 -2426
rect 2843 -2430 2849 -2410
rect 2573 -2448 2581 -2438
rect 2600 -2446 2603 -2438
rect 2604 -2446 2622 -2438
rect 2667 -2446 2699 -2438
rect 2744 -2446 2762 -2438
rect 2600 -2448 2766 -2446
rect 2785 -2448 2796 -2438
rect 2858 -2448 2871 -2410
rect 2943 -2396 2972 -2380
rect 2986 -2396 3015 -2380
rect 3030 -2390 3060 -2374
rect 3088 -2396 3094 -2348
rect 3097 -2354 3116 -2348
rect 3131 -2354 3161 -2346
rect 3097 -2362 3161 -2354
rect 3097 -2378 3177 -2362
rect 3193 -2369 3255 -2338
rect 3271 -2369 3333 -2338
rect 3402 -2340 3451 -2315
rect 3466 -2340 3496 -2322
rect 3365 -2354 3395 -2346
rect 3402 -2348 3512 -2340
rect 3365 -2362 3410 -2354
rect 3097 -2380 3116 -2378
rect 3131 -2380 3177 -2378
rect 3097 -2396 3177 -2380
rect 3204 -2382 3239 -2369
rect 3280 -2372 3317 -2369
rect 3280 -2374 3322 -2372
rect 3209 -2385 3239 -2382
rect 3218 -2389 3225 -2385
rect 3225 -2390 3226 -2389
rect 3184 -2396 3194 -2390
rect 2943 -2404 2978 -2396
rect 2943 -2430 2944 -2404
rect 2951 -2430 2978 -2404
rect 2943 -2438 2978 -2430
rect 2980 -2404 3021 -2396
rect 2980 -2430 2995 -2404
rect 3002 -2430 3021 -2404
rect 3085 -2408 3116 -2396
rect 3131 -2408 3234 -2396
rect 3246 -2406 3272 -2380
rect 3287 -2385 3317 -2374
rect 3349 -2378 3411 -2362
rect 3349 -2380 3395 -2378
rect 3349 -2396 3411 -2380
rect 3423 -2396 3429 -2348
rect 3432 -2356 3512 -2348
rect 3432 -2358 3451 -2356
rect 3466 -2358 3500 -2356
rect 3432 -2373 3512 -2358
rect 3432 -2374 3518 -2373
rect 3432 -2396 3451 -2374
rect 3466 -2390 3496 -2374
rect 3524 -2380 3530 -2306
rect 3533 -2380 3552 -2236
rect 3567 -2380 3573 -2236
rect 3582 -2306 3595 -2236
rect 3647 -2240 3669 -2236
rect 3640 -2252 3657 -2248
rect 3661 -2250 3669 -2248
rect 3659 -2252 3669 -2250
rect 3640 -2262 3669 -2252
rect 3722 -2262 3738 -2248
rect 3776 -2258 3782 -2250
rect 3789 -2252 3897 -2236
rect 3640 -2264 3738 -2262
rect 3624 -2272 3675 -2264
rect 3722 -2272 3756 -2264
rect 3624 -2284 3649 -2272
rect 3656 -2284 3675 -2272
rect 3729 -2274 3756 -2272
rect 3765 -2272 3782 -2258
rect 3827 -2272 3859 -2252
rect 3904 -2258 3910 -2250
rect 3918 -2258 3933 -2236
rect 3999 -2242 4018 -2239
rect 3904 -2264 3933 -2258
rect 3948 -2262 3964 -2248
rect 3999 -2261 4021 -2242
rect 4031 -2248 4047 -2247
rect 4030 -2250 4047 -2248
rect 4031 -2255 4047 -2250
rect 4021 -2262 4027 -2261
rect 4030 -2262 4059 -2255
rect 3948 -2263 4059 -2262
rect 3948 -2264 4065 -2263
rect 3904 -2272 3986 -2264
rect 4021 -2267 4027 -2264
rect 3765 -2274 3986 -2272
rect 3729 -2278 3801 -2274
rect 3829 -2276 3857 -2274
rect 3882 -2278 3986 -2274
rect 3624 -2292 3675 -2284
rect 3722 -2286 3854 -2278
rect 3859 -2286 3986 -2278
rect 4030 -2272 4065 -2264
rect 3722 -2288 3801 -2286
rect 3882 -2288 3986 -2286
rect 3722 -2292 3819 -2288
rect 3576 -2340 3595 -2306
rect 3640 -2300 3669 -2292
rect 3640 -2306 3657 -2300
rect 3640 -2308 3674 -2306
rect 3722 -2308 3738 -2292
rect 3739 -2296 3819 -2292
rect 3867 -2292 3986 -2288
rect 3867 -2296 3947 -2292
rect 3739 -2302 3947 -2296
rect 3948 -2302 3964 -2292
rect 4012 -2296 4027 -2281
rect 4030 -2284 4031 -2272
rect 4038 -2284 4065 -2272
rect 4030 -2292 4065 -2284
rect 4030 -2293 4059 -2292
rect 3750 -2306 3854 -2302
rect 3641 -2312 3674 -2308
rect 3637 -2314 3674 -2312
rect 3637 -2315 3704 -2314
rect 3637 -2320 3668 -2315
rect 3674 -2320 3704 -2315
rect 3765 -2318 3780 -2306
rect 3637 -2324 3704 -2320
rect 3610 -2327 3704 -2324
rect 3610 -2334 3659 -2327
rect 3610 -2340 3640 -2334
rect 3659 -2339 3664 -2334
rect 3576 -2356 3656 -2340
rect 3668 -2348 3704 -2327
rect 3789 -2328 3819 -2319
rect 3842 -2324 3860 -2306
rect 3918 -2308 3964 -2302
rect 3999 -2306 4012 -2296
rect 4030 -2306 4047 -2293
rect 3999 -2308 4047 -2306
rect 3880 -2314 3882 -2312
rect 3882 -2319 3894 -2314
rect 3867 -2326 3897 -2319
rect 3867 -2328 3898 -2326
rect 3918 -2328 3954 -2308
rect 3999 -2309 4046 -2308
rect 4012 -2314 4046 -2309
rect 4086 -2314 4102 -2312
rect 3765 -2332 3954 -2328
rect 3780 -2335 3954 -2332
rect 3773 -2338 3954 -2335
rect 3982 -2315 4046 -2314
rect 3576 -2358 3595 -2356
rect 3610 -2358 3644 -2356
rect 3576 -2374 3656 -2358
rect 3576 -2380 3595 -2374
rect 3292 -2406 3395 -2396
rect 3246 -2408 3395 -2406
rect 3416 -2408 3451 -2396
rect 3085 -2410 3247 -2408
rect 3097 -2430 3116 -2410
rect 3131 -2412 3161 -2410
rect 2980 -2438 3021 -2430
rect 2943 -2448 2972 -2438
rect 2986 -2448 3015 -2438
rect 3103 -2448 3116 -2430
rect 3168 -2426 3247 -2410
rect 3279 -2410 3451 -2408
rect 3279 -2426 3358 -2410
rect 3365 -2412 3395 -2410
rect 3168 -2438 3358 -2426
rect 3423 -2430 3429 -2410
rect 3153 -2448 3161 -2438
rect 3180 -2446 3183 -2438
rect 3184 -2446 3202 -2438
rect 3247 -2446 3279 -2438
rect 3324 -2446 3342 -2438
rect 3180 -2448 3346 -2446
rect 3365 -2448 3376 -2438
rect 3438 -2448 3451 -2410
rect 3523 -2396 3552 -2380
rect 3566 -2396 3595 -2380
rect 3610 -2390 3640 -2374
rect 3668 -2396 3674 -2348
rect 3677 -2354 3696 -2348
rect 3711 -2354 3741 -2346
rect 3677 -2362 3741 -2354
rect 3677 -2378 3757 -2362
rect 3773 -2369 3835 -2338
rect 3851 -2369 3913 -2338
rect 3982 -2340 4031 -2315
rect 4076 -2324 4102 -2314
rect 4046 -2340 4102 -2324
rect 3945 -2354 3975 -2346
rect 3982 -2348 4092 -2340
rect 3945 -2362 3990 -2354
rect 3677 -2380 3696 -2378
rect 3711 -2380 3757 -2378
rect 3677 -2396 3757 -2380
rect 3784 -2382 3819 -2369
rect 3860 -2372 3897 -2369
rect 3860 -2374 3902 -2372
rect 3789 -2385 3819 -2382
rect 3798 -2389 3805 -2385
rect 3805 -2390 3806 -2389
rect 3764 -2396 3774 -2390
rect 3523 -2404 3558 -2396
rect 3523 -2430 3524 -2404
rect 3531 -2430 3558 -2404
rect 3523 -2438 3558 -2430
rect 3560 -2404 3601 -2396
rect 3560 -2430 3575 -2404
rect 3582 -2430 3601 -2404
rect 3665 -2408 3696 -2396
rect 3711 -2408 3814 -2396
rect 3826 -2406 3852 -2380
rect 3867 -2385 3897 -2374
rect 3929 -2378 3991 -2362
rect 3929 -2380 3975 -2378
rect 3929 -2396 3991 -2380
rect 4003 -2396 4009 -2348
rect 4012 -2356 4092 -2348
rect 4012 -2358 4031 -2356
rect 4046 -2358 4080 -2356
rect 4012 -2374 4092 -2358
rect 4012 -2396 4031 -2374
rect 4046 -2390 4076 -2374
rect 4104 -2380 4110 -2306
rect 4113 -2380 4132 -2236
rect 4147 -2380 4153 -2236
rect 4162 -2306 4175 -2236
rect 4227 -2240 4249 -2236
rect 4220 -2252 4237 -2248
rect 4241 -2250 4249 -2248
rect 4239 -2252 4249 -2250
rect 4220 -2262 4249 -2252
rect 4302 -2262 4318 -2248
rect 4356 -2258 4362 -2250
rect 4369 -2252 4477 -2236
rect 4220 -2264 4318 -2262
rect 4204 -2272 4255 -2264
rect 4302 -2272 4336 -2264
rect 4204 -2284 4229 -2272
rect 4236 -2284 4255 -2272
rect 4309 -2274 4336 -2272
rect 4345 -2272 4362 -2258
rect 4407 -2272 4439 -2252
rect 4484 -2258 4490 -2250
rect 4498 -2258 4513 -2236
rect 4579 -2242 4598 -2239
rect 4484 -2264 4513 -2258
rect 4528 -2262 4544 -2248
rect 4579 -2261 4601 -2242
rect 4611 -2248 4627 -2247
rect 4610 -2250 4627 -2248
rect 4611 -2255 4627 -2250
rect 4601 -2262 4607 -2261
rect 4610 -2262 4639 -2255
rect 4528 -2263 4639 -2262
rect 4528 -2264 4645 -2263
rect 4484 -2272 4566 -2264
rect 4601 -2267 4607 -2264
rect 4345 -2274 4566 -2272
rect 4309 -2278 4381 -2274
rect 4409 -2276 4437 -2274
rect 4462 -2278 4566 -2274
rect 4204 -2292 4255 -2284
rect 4302 -2286 4434 -2278
rect 4439 -2286 4566 -2278
rect 4610 -2272 4645 -2264
rect 4302 -2288 4381 -2286
rect 4462 -2288 4566 -2286
rect 4302 -2292 4399 -2288
rect 4156 -2340 4175 -2306
rect 4220 -2300 4249 -2292
rect 4220 -2306 4237 -2300
rect 4220 -2308 4254 -2306
rect 4302 -2308 4318 -2292
rect 4319 -2296 4399 -2292
rect 4447 -2292 4566 -2288
rect 4447 -2296 4527 -2292
rect 4319 -2302 4527 -2296
rect 4528 -2302 4544 -2292
rect 4592 -2296 4607 -2281
rect 4610 -2284 4611 -2272
rect 4618 -2284 4645 -2272
rect 4610 -2292 4645 -2284
rect 4610 -2293 4639 -2292
rect 4330 -2306 4434 -2302
rect 4221 -2312 4254 -2308
rect 4217 -2314 4254 -2312
rect 4217 -2315 4284 -2314
rect 4217 -2320 4248 -2315
rect 4254 -2320 4284 -2315
rect 4345 -2318 4360 -2306
rect 4217 -2324 4284 -2320
rect 4190 -2327 4284 -2324
rect 4190 -2334 4239 -2327
rect 4190 -2340 4220 -2334
rect 4239 -2339 4244 -2334
rect 4156 -2356 4236 -2340
rect 4248 -2348 4284 -2327
rect 4369 -2328 4399 -2319
rect 4422 -2324 4440 -2306
rect 4498 -2308 4544 -2302
rect 4579 -2306 4592 -2296
rect 4610 -2306 4627 -2293
rect 4579 -2308 4627 -2306
rect 4460 -2314 4462 -2312
rect 4462 -2319 4474 -2314
rect 4447 -2326 4477 -2319
rect 4447 -2328 4478 -2326
rect 4498 -2328 4534 -2308
rect 4579 -2309 4626 -2308
rect 4592 -2314 4626 -2309
rect 4345 -2332 4534 -2328
rect 4360 -2335 4534 -2332
rect 4353 -2338 4534 -2335
rect 4562 -2315 4626 -2314
rect 4156 -2358 4175 -2356
rect 4190 -2358 4224 -2356
rect 4156 -2374 4236 -2358
rect 4156 -2380 4175 -2374
rect 3872 -2406 3975 -2396
rect 3826 -2408 3975 -2406
rect 3996 -2408 4031 -2396
rect 3665 -2410 3827 -2408
rect 3677 -2430 3696 -2410
rect 3711 -2412 3741 -2410
rect 3560 -2438 3601 -2430
rect 3523 -2448 3552 -2438
rect 3566 -2448 3595 -2438
rect 3683 -2448 3696 -2430
rect 3748 -2426 3827 -2410
rect 3859 -2410 4031 -2408
rect 3859 -2426 3938 -2410
rect 3945 -2412 3975 -2410
rect 3748 -2438 3938 -2426
rect 4003 -2430 4009 -2410
rect 3733 -2448 3741 -2438
rect 3760 -2446 3763 -2438
rect 3764 -2446 3782 -2438
rect 3827 -2446 3859 -2438
rect 3904 -2446 3922 -2438
rect 3760 -2448 3926 -2446
rect 3945 -2448 3956 -2438
rect 4018 -2448 4031 -2410
rect 4103 -2396 4132 -2380
rect 4146 -2396 4175 -2380
rect 4190 -2390 4220 -2374
rect 4248 -2396 4254 -2348
rect 4257 -2354 4276 -2348
rect 4291 -2354 4321 -2346
rect 4257 -2362 4321 -2354
rect 4257 -2378 4337 -2362
rect 4353 -2369 4415 -2338
rect 4431 -2369 4493 -2338
rect 4562 -2340 4611 -2315
rect 4626 -2340 4656 -2322
rect 4525 -2354 4555 -2346
rect 4562 -2348 4672 -2340
rect 4525 -2362 4570 -2354
rect 4257 -2380 4276 -2378
rect 4291 -2380 4337 -2378
rect 4257 -2396 4337 -2380
rect 4364 -2382 4399 -2369
rect 4440 -2372 4477 -2369
rect 4440 -2374 4482 -2372
rect 4369 -2385 4399 -2382
rect 4378 -2389 4385 -2385
rect 4385 -2390 4386 -2389
rect 4344 -2396 4354 -2390
rect 4103 -2404 4138 -2396
rect 4103 -2430 4104 -2404
rect 4111 -2430 4138 -2404
rect 4103 -2438 4138 -2430
rect 4140 -2404 4181 -2396
rect 4140 -2430 4155 -2404
rect 4162 -2430 4181 -2404
rect 4245 -2408 4276 -2396
rect 4291 -2408 4394 -2396
rect 4406 -2406 4432 -2380
rect 4447 -2385 4477 -2374
rect 4509 -2378 4571 -2362
rect 4509 -2380 4555 -2378
rect 4509 -2396 4571 -2380
rect 4583 -2396 4589 -2348
rect 4592 -2356 4672 -2348
rect 4592 -2358 4611 -2356
rect 4626 -2358 4660 -2356
rect 4592 -2373 4672 -2358
rect 4592 -2374 4678 -2373
rect 4592 -2396 4611 -2374
rect 4626 -2390 4656 -2374
rect 4684 -2380 4690 -2306
rect 4693 -2380 4712 -2236
rect 4727 -2380 4733 -2236
rect 4742 -2306 4755 -2236
rect 4807 -2240 4829 -2236
rect 4800 -2252 4817 -2248
rect 4821 -2250 4829 -2248
rect 4819 -2252 4829 -2250
rect 4800 -2262 4829 -2252
rect 4882 -2262 4898 -2248
rect 4936 -2258 4942 -2250
rect 4949 -2252 5057 -2236
rect 4800 -2264 4898 -2262
rect 4784 -2272 4835 -2264
rect 4882 -2272 4916 -2264
rect 4784 -2284 4809 -2272
rect 4816 -2284 4835 -2272
rect 4889 -2274 4916 -2272
rect 4925 -2272 4942 -2258
rect 4987 -2272 5019 -2252
rect 5064 -2258 5070 -2250
rect 5078 -2258 5093 -2236
rect 5159 -2242 5178 -2239
rect 5064 -2264 5093 -2258
rect 5108 -2262 5124 -2248
rect 5159 -2261 5181 -2242
rect 5191 -2248 5207 -2247
rect 5190 -2250 5207 -2248
rect 5191 -2255 5207 -2250
rect 5181 -2262 5187 -2261
rect 5190 -2262 5219 -2255
rect 5108 -2263 5219 -2262
rect 5108 -2264 5225 -2263
rect 5064 -2272 5146 -2264
rect 5181 -2267 5187 -2264
rect 4925 -2274 5146 -2272
rect 4889 -2278 4961 -2274
rect 4989 -2276 5017 -2274
rect 5042 -2278 5146 -2274
rect 4784 -2292 4835 -2284
rect 4882 -2286 5014 -2278
rect 5019 -2286 5146 -2278
rect 5190 -2272 5225 -2264
rect 4882 -2288 4961 -2286
rect 5042 -2288 5146 -2286
rect 4882 -2292 4979 -2288
rect 4736 -2340 4755 -2306
rect 4800 -2300 4829 -2292
rect 4800 -2306 4817 -2300
rect 4800 -2308 4834 -2306
rect 4882 -2308 4898 -2292
rect 4899 -2296 4979 -2292
rect 5027 -2292 5146 -2288
rect 5027 -2296 5107 -2292
rect 4899 -2302 5107 -2296
rect 5108 -2302 5124 -2292
rect 5172 -2296 5187 -2281
rect 5190 -2284 5191 -2272
rect 5198 -2284 5225 -2272
rect 5190 -2292 5225 -2284
rect 5190 -2293 5219 -2292
rect 4910 -2306 5014 -2302
rect 4801 -2312 4834 -2308
rect 4797 -2314 4834 -2312
rect 4797 -2315 4864 -2314
rect 4797 -2320 4828 -2315
rect 4834 -2320 4864 -2315
rect 4925 -2318 4940 -2306
rect 4797 -2324 4864 -2320
rect 4770 -2327 4864 -2324
rect 4770 -2334 4819 -2327
rect 4770 -2340 4800 -2334
rect 4819 -2339 4824 -2334
rect 4736 -2356 4816 -2340
rect 4828 -2348 4864 -2327
rect 4949 -2328 4979 -2319
rect 5002 -2324 5020 -2306
rect 5078 -2308 5124 -2302
rect 5159 -2306 5172 -2296
rect 5190 -2306 5207 -2293
rect 5159 -2308 5207 -2306
rect 5040 -2314 5042 -2312
rect 5042 -2319 5054 -2314
rect 5027 -2326 5057 -2319
rect 5027 -2328 5058 -2326
rect 5078 -2328 5114 -2308
rect 5159 -2309 5206 -2308
rect 5172 -2314 5206 -2309
rect 5246 -2314 5262 -2312
rect 4925 -2332 5114 -2328
rect 4940 -2335 5114 -2332
rect 4933 -2338 5114 -2335
rect 5142 -2315 5206 -2314
rect 4736 -2358 4755 -2356
rect 4770 -2358 4804 -2356
rect 4736 -2374 4816 -2358
rect 4736 -2380 4755 -2374
rect 4452 -2406 4555 -2396
rect 4406 -2408 4555 -2406
rect 4576 -2408 4611 -2396
rect 4245 -2410 4407 -2408
rect 4257 -2430 4276 -2410
rect 4291 -2412 4321 -2410
rect 4140 -2438 4181 -2430
rect 4103 -2448 4132 -2438
rect 4146 -2448 4175 -2438
rect 4263 -2448 4276 -2430
rect 4328 -2426 4407 -2410
rect 4439 -2410 4611 -2408
rect 4439 -2426 4518 -2410
rect 4525 -2412 4555 -2410
rect 4328 -2438 4518 -2426
rect 4583 -2430 4589 -2410
rect 4313 -2448 4321 -2438
rect 4340 -2446 4343 -2438
rect 4344 -2446 4362 -2438
rect 4407 -2446 4439 -2438
rect 4484 -2446 4502 -2438
rect 4340 -2448 4506 -2446
rect 4525 -2448 4536 -2438
rect 4598 -2448 4611 -2410
rect 4683 -2396 4712 -2380
rect 4726 -2396 4755 -2380
rect 4770 -2390 4800 -2374
rect 4828 -2396 4834 -2348
rect 4837 -2354 4856 -2348
rect 4871 -2354 4901 -2346
rect 4837 -2362 4901 -2354
rect 4837 -2378 4917 -2362
rect 4933 -2369 4995 -2338
rect 5011 -2369 5073 -2338
rect 5142 -2340 5191 -2315
rect 5236 -2324 5262 -2314
rect 5206 -2340 5262 -2324
rect 5105 -2354 5135 -2346
rect 5142 -2348 5252 -2340
rect 5105 -2362 5150 -2354
rect 4837 -2380 4856 -2378
rect 4871 -2380 4917 -2378
rect 4837 -2396 4917 -2380
rect 4944 -2382 4979 -2369
rect 5020 -2372 5057 -2369
rect 5020 -2374 5062 -2372
rect 4949 -2385 4979 -2382
rect 4958 -2389 4965 -2385
rect 4965 -2390 4966 -2389
rect 4924 -2396 4934 -2390
rect 4683 -2404 4718 -2396
rect 4683 -2430 4684 -2404
rect 4691 -2430 4718 -2404
rect 4683 -2438 4718 -2430
rect 4720 -2404 4761 -2396
rect 4720 -2430 4735 -2404
rect 4742 -2430 4761 -2404
rect 4825 -2408 4856 -2396
rect 4871 -2408 4974 -2396
rect 4986 -2406 5012 -2380
rect 5027 -2385 5057 -2374
rect 5089 -2378 5151 -2362
rect 5089 -2380 5135 -2378
rect 5089 -2396 5151 -2380
rect 5163 -2396 5169 -2348
rect 5172 -2356 5252 -2348
rect 5172 -2358 5191 -2356
rect 5206 -2358 5240 -2356
rect 5172 -2374 5252 -2358
rect 5172 -2396 5191 -2374
rect 5206 -2390 5236 -2374
rect 5264 -2380 5270 -2306
rect 5273 -2380 5292 -2236
rect 5307 -2380 5313 -2236
rect 5322 -2306 5335 -2236
rect 5387 -2240 5409 -2236
rect 5380 -2252 5397 -2248
rect 5401 -2250 5409 -2248
rect 5399 -2252 5409 -2250
rect 5380 -2262 5409 -2252
rect 5462 -2262 5478 -2248
rect 5516 -2258 5522 -2250
rect 5529 -2252 5637 -2236
rect 5380 -2264 5478 -2262
rect 5364 -2272 5415 -2264
rect 5462 -2272 5496 -2264
rect 5364 -2284 5389 -2272
rect 5396 -2284 5415 -2272
rect 5469 -2274 5496 -2272
rect 5505 -2272 5522 -2258
rect 5567 -2272 5599 -2252
rect 5644 -2258 5650 -2250
rect 5658 -2258 5673 -2236
rect 5739 -2242 5758 -2239
rect 5644 -2264 5673 -2258
rect 5688 -2262 5704 -2248
rect 5739 -2261 5761 -2242
rect 5771 -2248 5787 -2247
rect 5770 -2250 5787 -2248
rect 5771 -2255 5787 -2250
rect 5761 -2262 5767 -2261
rect 5770 -2262 5799 -2255
rect 5688 -2263 5799 -2262
rect 5688 -2264 5805 -2263
rect 5644 -2272 5726 -2264
rect 5761 -2267 5767 -2264
rect 5505 -2274 5726 -2272
rect 5469 -2278 5541 -2274
rect 5569 -2276 5597 -2274
rect 5622 -2278 5726 -2274
rect 5364 -2292 5415 -2284
rect 5462 -2286 5594 -2278
rect 5599 -2286 5726 -2278
rect 5770 -2272 5805 -2264
rect 5462 -2288 5541 -2286
rect 5622 -2288 5726 -2286
rect 5462 -2292 5559 -2288
rect 5316 -2340 5335 -2306
rect 5380 -2300 5409 -2292
rect 5380 -2306 5397 -2300
rect 5380 -2308 5414 -2306
rect 5462 -2308 5478 -2292
rect 5479 -2296 5559 -2292
rect 5607 -2292 5726 -2288
rect 5607 -2296 5687 -2292
rect 5479 -2302 5687 -2296
rect 5688 -2302 5704 -2292
rect 5752 -2296 5767 -2281
rect 5770 -2284 5771 -2272
rect 5778 -2284 5805 -2272
rect 5770 -2292 5805 -2284
rect 5770 -2293 5799 -2292
rect 5490 -2306 5594 -2302
rect 5381 -2312 5414 -2308
rect 5377 -2314 5414 -2312
rect 5377 -2315 5444 -2314
rect 5377 -2320 5408 -2315
rect 5414 -2320 5444 -2315
rect 5505 -2318 5520 -2306
rect 5377 -2324 5444 -2320
rect 5350 -2327 5444 -2324
rect 5350 -2334 5399 -2327
rect 5350 -2340 5380 -2334
rect 5399 -2339 5404 -2334
rect 5316 -2356 5396 -2340
rect 5408 -2348 5444 -2327
rect 5529 -2328 5559 -2319
rect 5582 -2324 5600 -2306
rect 5658 -2308 5704 -2302
rect 5739 -2306 5752 -2296
rect 5770 -2306 5787 -2293
rect 5739 -2308 5787 -2306
rect 5620 -2314 5622 -2312
rect 5622 -2319 5634 -2314
rect 5607 -2326 5637 -2319
rect 5607 -2328 5638 -2326
rect 5658 -2328 5694 -2308
rect 5739 -2309 5786 -2308
rect 5752 -2314 5786 -2309
rect 5505 -2332 5694 -2328
rect 5520 -2335 5694 -2332
rect 5513 -2338 5694 -2335
rect 5722 -2315 5786 -2314
rect 5316 -2358 5335 -2356
rect 5350 -2358 5384 -2356
rect 5316 -2374 5396 -2358
rect 5316 -2380 5335 -2374
rect 5032 -2406 5135 -2396
rect 4986 -2408 5135 -2406
rect 5156 -2408 5191 -2396
rect 4825 -2410 4987 -2408
rect 4837 -2430 4856 -2410
rect 4871 -2412 4901 -2410
rect 4720 -2438 4761 -2430
rect 4683 -2448 4712 -2438
rect 4726 -2448 4755 -2438
rect 4843 -2448 4856 -2430
rect 4908 -2426 4987 -2410
rect 5019 -2410 5191 -2408
rect 5019 -2426 5098 -2410
rect 5105 -2412 5135 -2410
rect 4908 -2438 5098 -2426
rect 5163 -2430 5169 -2410
rect 4893 -2448 4901 -2438
rect 4920 -2446 4923 -2438
rect 4924 -2446 4942 -2438
rect 4987 -2446 5019 -2438
rect 5064 -2446 5082 -2438
rect 4920 -2448 5086 -2446
rect 5105 -2448 5116 -2438
rect 5178 -2448 5191 -2410
rect 5263 -2396 5292 -2380
rect 5306 -2396 5335 -2380
rect 5350 -2390 5380 -2374
rect 5408 -2396 5414 -2348
rect 5417 -2354 5436 -2348
rect 5451 -2354 5481 -2346
rect 5417 -2362 5481 -2354
rect 5417 -2378 5497 -2362
rect 5513 -2369 5575 -2338
rect 5591 -2369 5653 -2338
rect 5722 -2340 5771 -2315
rect 5786 -2340 5816 -2322
rect 5685 -2354 5715 -2346
rect 5722 -2348 5832 -2340
rect 5685 -2362 5730 -2354
rect 5417 -2380 5436 -2378
rect 5451 -2380 5497 -2378
rect 5417 -2396 5497 -2380
rect 5524 -2382 5559 -2369
rect 5600 -2372 5637 -2369
rect 5600 -2374 5642 -2372
rect 5529 -2385 5559 -2382
rect 5538 -2389 5545 -2385
rect 5545 -2390 5546 -2389
rect 5504 -2396 5514 -2390
rect 5263 -2404 5298 -2396
rect 5263 -2430 5264 -2404
rect 5271 -2430 5298 -2404
rect 5263 -2438 5298 -2430
rect 5300 -2404 5341 -2396
rect 5300 -2430 5315 -2404
rect 5322 -2430 5341 -2404
rect 5405 -2408 5436 -2396
rect 5451 -2408 5554 -2396
rect 5566 -2406 5592 -2380
rect 5607 -2385 5637 -2374
rect 5669 -2378 5731 -2362
rect 5669 -2380 5715 -2378
rect 5669 -2396 5731 -2380
rect 5743 -2396 5749 -2348
rect 5752 -2356 5832 -2348
rect 5752 -2358 5771 -2356
rect 5786 -2358 5820 -2356
rect 5752 -2373 5832 -2358
rect 5752 -2374 5838 -2373
rect 5752 -2396 5771 -2374
rect 5786 -2390 5816 -2374
rect 5844 -2380 5850 -2306
rect 5853 -2380 5872 -2236
rect 5887 -2380 5893 -2236
rect 5902 -2306 5915 -2236
rect 5967 -2240 5989 -2236
rect 5960 -2252 5977 -2248
rect 5981 -2250 5989 -2248
rect 5979 -2252 5989 -2250
rect 5960 -2262 5989 -2252
rect 6042 -2262 6058 -2248
rect 6096 -2258 6102 -2250
rect 6109 -2252 6217 -2236
rect 5960 -2264 6058 -2262
rect 5944 -2272 5995 -2264
rect 6042 -2272 6076 -2264
rect 5944 -2284 5969 -2272
rect 5976 -2284 5995 -2272
rect 6049 -2274 6076 -2272
rect 6085 -2272 6102 -2258
rect 6147 -2272 6179 -2252
rect 6224 -2258 6230 -2250
rect 6238 -2258 6253 -2236
rect 6319 -2242 6338 -2239
rect 6224 -2264 6253 -2258
rect 6268 -2262 6284 -2248
rect 6319 -2261 6341 -2242
rect 6351 -2248 6367 -2247
rect 6350 -2250 6367 -2248
rect 6351 -2255 6367 -2250
rect 6341 -2262 6347 -2261
rect 6350 -2262 6379 -2255
rect 6268 -2263 6379 -2262
rect 6268 -2264 6385 -2263
rect 6224 -2272 6306 -2264
rect 6341 -2267 6347 -2264
rect 6085 -2274 6306 -2272
rect 6049 -2278 6121 -2274
rect 6149 -2276 6177 -2274
rect 6202 -2278 6306 -2274
rect 5944 -2292 5995 -2284
rect 6042 -2286 6174 -2278
rect 6179 -2286 6306 -2278
rect 6350 -2272 6385 -2264
rect 6042 -2288 6121 -2286
rect 6202 -2288 6306 -2286
rect 6042 -2292 6139 -2288
rect 5896 -2340 5915 -2306
rect 5960 -2300 5989 -2292
rect 5960 -2306 5977 -2300
rect 5960 -2308 5994 -2306
rect 6042 -2308 6058 -2292
rect 6059 -2296 6139 -2292
rect 6187 -2292 6306 -2288
rect 6187 -2296 6267 -2292
rect 6059 -2302 6267 -2296
rect 6268 -2302 6284 -2292
rect 6332 -2296 6347 -2281
rect 6350 -2284 6351 -2272
rect 6358 -2284 6385 -2272
rect 6350 -2292 6385 -2284
rect 6350 -2293 6379 -2292
rect 6070 -2306 6174 -2302
rect 5961 -2312 5994 -2308
rect 5957 -2314 5994 -2312
rect 5957 -2315 6024 -2314
rect 5957 -2320 5988 -2315
rect 5994 -2320 6024 -2315
rect 6085 -2318 6100 -2306
rect 5957 -2324 6024 -2320
rect 5930 -2327 6024 -2324
rect 5930 -2334 5979 -2327
rect 5930 -2340 5960 -2334
rect 5979 -2339 5984 -2334
rect 5896 -2356 5976 -2340
rect 5988 -2348 6024 -2327
rect 6109 -2328 6139 -2319
rect 6162 -2324 6180 -2306
rect 6238 -2308 6284 -2302
rect 6319 -2306 6332 -2296
rect 6350 -2306 6367 -2293
rect 6319 -2308 6367 -2306
rect 6200 -2314 6202 -2312
rect 6202 -2319 6214 -2314
rect 6187 -2326 6217 -2319
rect 6187 -2328 6218 -2326
rect 6238 -2328 6274 -2308
rect 6319 -2309 6366 -2308
rect 6332 -2314 6366 -2309
rect 6085 -2332 6274 -2328
rect 6100 -2335 6274 -2332
rect 6093 -2338 6274 -2335
rect 6302 -2315 6366 -2314
rect 5896 -2358 5915 -2356
rect 5930 -2358 5964 -2356
rect 5896 -2374 5976 -2358
rect 5896 -2380 5915 -2374
rect 5612 -2406 5715 -2396
rect 5566 -2408 5715 -2406
rect 5736 -2408 5771 -2396
rect 5405 -2410 5567 -2408
rect 5417 -2430 5436 -2410
rect 5451 -2412 5481 -2410
rect 5300 -2438 5341 -2430
rect 5263 -2448 5292 -2438
rect 5306 -2448 5335 -2438
rect 5423 -2448 5436 -2430
rect 5488 -2426 5567 -2410
rect 5599 -2410 5771 -2408
rect 5599 -2426 5678 -2410
rect 5685 -2412 5715 -2410
rect 5488 -2438 5678 -2426
rect 5743 -2430 5749 -2410
rect 5473 -2448 5481 -2438
rect 5500 -2446 5503 -2438
rect 5504 -2446 5522 -2438
rect 5567 -2446 5599 -2438
rect 5644 -2446 5662 -2438
rect 5500 -2448 5666 -2446
rect 5685 -2448 5696 -2438
rect 5758 -2448 5771 -2410
rect 5843 -2396 5872 -2380
rect 5886 -2396 5915 -2380
rect 5930 -2390 5960 -2374
rect 5988 -2396 5994 -2348
rect 5997 -2354 6016 -2348
rect 6031 -2354 6061 -2346
rect 5997 -2362 6061 -2354
rect 5997 -2378 6077 -2362
rect 6093 -2369 6155 -2338
rect 6171 -2369 6233 -2338
rect 6302 -2340 6351 -2315
rect 6366 -2340 6396 -2324
rect 6265 -2354 6295 -2346
rect 6302 -2348 6412 -2340
rect 6265 -2362 6310 -2354
rect 5997 -2380 6016 -2378
rect 6031 -2380 6077 -2378
rect 5997 -2396 6077 -2380
rect 6104 -2382 6139 -2369
rect 6180 -2372 6217 -2369
rect 6180 -2374 6222 -2372
rect 6109 -2385 6139 -2382
rect 6118 -2389 6125 -2385
rect 6125 -2390 6126 -2389
rect 6084 -2396 6094 -2390
rect 5843 -2404 5878 -2396
rect 5843 -2430 5844 -2404
rect 5851 -2430 5878 -2404
rect 5843 -2438 5878 -2430
rect 5880 -2404 5921 -2396
rect 5880 -2430 5895 -2404
rect 5902 -2430 5921 -2404
rect 5985 -2408 6016 -2396
rect 6031 -2408 6134 -2396
rect 6146 -2406 6172 -2380
rect 6187 -2385 6217 -2374
rect 6249 -2378 6311 -2362
rect 6249 -2380 6295 -2378
rect 6249 -2396 6311 -2380
rect 6323 -2396 6329 -2348
rect 6332 -2356 6412 -2348
rect 6332 -2358 6351 -2356
rect 6366 -2358 6400 -2356
rect 6332 -2374 6412 -2358
rect 6332 -2396 6351 -2374
rect 6366 -2390 6396 -2374
rect 6424 -2380 6430 -2306
rect 6439 -2380 6452 -2236
rect 6192 -2406 6295 -2396
rect 6146 -2408 6295 -2406
rect 6316 -2408 6351 -2396
rect 5985 -2410 6147 -2408
rect 5997 -2430 6016 -2410
rect 6031 -2412 6061 -2410
rect 5880 -2438 5921 -2430
rect 5843 -2448 5872 -2438
rect 5886 -2448 5915 -2438
rect 6003 -2448 6016 -2430
rect 6068 -2426 6147 -2410
rect 6179 -2410 6351 -2408
rect 6179 -2426 6258 -2410
rect 6265 -2412 6295 -2410
rect 6068 -2438 6258 -2426
rect 6323 -2430 6329 -2410
rect 6053 -2448 6061 -2438
rect 6080 -2446 6083 -2438
rect 6084 -2446 6102 -2438
rect 6147 -2446 6179 -2438
rect 6224 -2446 6242 -2438
rect 6080 -2448 6246 -2446
rect 6265 -2448 6276 -2438
rect 6338 -2448 6351 -2410
rect 6423 -2396 6452 -2380
rect 6423 -2404 6458 -2396
rect 6423 -2430 6424 -2404
rect 6431 -2430 6458 -2404
rect 6423 -2438 6458 -2430
rect 6423 -2448 6452 -2438
rect -541 -2462 6452 -2448
rect -478 -2524 -465 -2462
rect -450 -2480 -420 -2462
rect -377 -2476 -334 -2462
rect -327 -2475 -319 -2462
rect -286 -2475 -148 -2462
rect -115 -2475 -107 -2462
rect -364 -2494 -334 -2476
rect -271 -2476 -163 -2475
rect -271 -2480 -241 -2476
rect -233 -2478 -201 -2476
rect -193 -2480 -163 -2476
rect -100 -2494 -70 -2462
rect -42 -2476 -29 -2462
rect -14 -2480 16 -2462
rect 53 -2524 72 -2462
rect 87 -2524 93 -2462
rect 102 -2524 115 -2462
rect 130 -2480 160 -2462
rect 203 -2476 246 -2462
rect 253 -2475 261 -2462
rect 294 -2475 432 -2462
rect 465 -2475 473 -2462
rect 216 -2494 246 -2476
rect 309 -2476 417 -2475
rect 309 -2480 339 -2476
rect 347 -2478 379 -2476
rect 387 -2480 417 -2476
rect 480 -2494 510 -2462
rect 538 -2476 551 -2462
rect 566 -2480 596 -2462
rect 633 -2524 652 -2462
rect 667 -2524 673 -2462
rect 682 -2524 695 -2462
rect 710 -2480 740 -2462
rect 783 -2476 826 -2462
rect 833 -2475 841 -2462
rect 874 -2475 1012 -2462
rect 1045 -2475 1053 -2462
rect 796 -2494 826 -2476
rect 889 -2476 997 -2475
rect 889 -2480 919 -2476
rect 927 -2478 959 -2476
rect 967 -2480 997 -2476
rect 1060 -2494 1090 -2462
rect 1118 -2476 1131 -2462
rect 1146 -2480 1176 -2462
rect 1213 -2524 1232 -2462
rect 1247 -2524 1253 -2462
rect 1262 -2524 1275 -2462
rect 1290 -2480 1320 -2462
rect 1363 -2476 1406 -2462
rect 1413 -2475 1421 -2462
rect 1454 -2475 1592 -2462
rect 1625 -2475 1633 -2462
rect 1376 -2494 1406 -2476
rect 1469 -2476 1577 -2475
rect 1469 -2480 1499 -2476
rect 1507 -2478 1539 -2476
rect 1547 -2480 1577 -2476
rect 1640 -2494 1670 -2462
rect 1698 -2476 1711 -2462
rect 1726 -2480 1756 -2462
rect 1793 -2524 1812 -2462
rect 1827 -2524 1833 -2462
rect 1842 -2524 1855 -2462
rect 1870 -2480 1900 -2462
rect 1943 -2476 1986 -2462
rect 1993 -2475 2001 -2462
rect 2034 -2475 2172 -2462
rect 2205 -2475 2213 -2462
rect 1956 -2494 1986 -2476
rect 2049 -2476 2157 -2475
rect 2049 -2480 2079 -2476
rect 2087 -2478 2119 -2476
rect 2127 -2480 2157 -2476
rect 2220 -2494 2250 -2462
rect 2278 -2476 2291 -2462
rect 2306 -2480 2336 -2462
rect 2373 -2524 2392 -2462
rect 2407 -2524 2413 -2462
rect 2422 -2524 2435 -2462
rect 2450 -2480 2480 -2462
rect 2523 -2476 2566 -2462
rect 2573 -2475 2581 -2462
rect 2614 -2475 2752 -2462
rect 2785 -2475 2793 -2462
rect 2536 -2494 2566 -2476
rect 2629 -2476 2737 -2475
rect 2629 -2480 2659 -2476
rect 2667 -2478 2699 -2476
rect 2707 -2480 2737 -2476
rect 2800 -2494 2830 -2462
rect 2858 -2476 2871 -2462
rect 2886 -2480 2916 -2462
rect 2953 -2524 2972 -2462
rect 2987 -2524 2993 -2462
rect 3002 -2524 3015 -2462
rect 3030 -2480 3060 -2462
rect 3103 -2476 3146 -2462
rect 3153 -2475 3161 -2462
rect 3194 -2475 3332 -2462
rect 3365 -2475 3373 -2462
rect 3116 -2494 3146 -2476
rect 3209 -2476 3317 -2475
rect 3209 -2480 3239 -2476
rect 3247 -2478 3279 -2476
rect 3287 -2480 3317 -2476
rect 3380 -2494 3410 -2462
rect 3438 -2476 3451 -2462
rect 3466 -2480 3496 -2462
rect 3533 -2524 3552 -2462
rect 3567 -2524 3573 -2462
rect 3582 -2524 3595 -2462
rect 3610 -2480 3640 -2462
rect 3683 -2476 3726 -2462
rect 3733 -2475 3741 -2462
rect 3774 -2475 3912 -2462
rect 3945 -2475 3953 -2462
rect 3696 -2494 3726 -2476
rect 3789 -2476 3897 -2475
rect 3789 -2480 3819 -2476
rect 3827 -2478 3859 -2476
rect 3867 -2480 3897 -2476
rect 3960 -2494 3990 -2462
rect 4018 -2476 4031 -2462
rect 4046 -2480 4076 -2462
rect 4113 -2524 4132 -2462
rect 4147 -2524 4153 -2462
rect 4162 -2524 4175 -2462
rect 4190 -2480 4220 -2462
rect 4263 -2476 4306 -2462
rect 4313 -2475 4321 -2462
rect 4354 -2475 4492 -2462
rect 4525 -2475 4533 -2462
rect 4276 -2494 4306 -2476
rect 4369 -2476 4477 -2475
rect 4369 -2480 4399 -2476
rect 4407 -2478 4439 -2476
rect 4447 -2480 4477 -2476
rect 4540 -2494 4570 -2462
rect 4598 -2476 4611 -2462
rect 4626 -2480 4656 -2462
rect 4693 -2524 4712 -2462
rect 4727 -2524 4733 -2462
rect 4742 -2524 4755 -2462
rect 4770 -2480 4800 -2462
rect 4843 -2476 4886 -2462
rect 4893 -2475 4901 -2462
rect 4934 -2475 5072 -2462
rect 5105 -2475 5113 -2462
rect 4856 -2494 4886 -2476
rect 4949 -2476 5057 -2475
rect 4949 -2480 4979 -2476
rect 4987 -2478 5019 -2476
rect 5027 -2480 5057 -2476
rect 5120 -2494 5150 -2462
rect 5178 -2476 5191 -2462
rect 5206 -2480 5236 -2462
rect 5273 -2524 5292 -2462
rect 5307 -2524 5313 -2462
rect 5322 -2524 5335 -2462
rect 5350 -2480 5380 -2462
rect 5423 -2476 5466 -2462
rect 5473 -2475 5481 -2462
rect 5514 -2475 5652 -2462
rect 5685 -2475 5693 -2462
rect 5436 -2494 5466 -2476
rect 5529 -2476 5637 -2475
rect 5529 -2480 5559 -2476
rect 5567 -2478 5599 -2476
rect 5607 -2480 5637 -2476
rect 5700 -2494 5730 -2462
rect 5758 -2476 5771 -2462
rect 5786 -2480 5816 -2462
rect 5853 -2524 5872 -2462
rect 5887 -2524 5893 -2462
rect 5902 -2524 5915 -2462
rect 5930 -2480 5960 -2462
rect 6003 -2476 6046 -2462
rect 6053 -2475 6061 -2462
rect 6094 -2475 6232 -2462
rect 6265 -2475 6273 -2462
rect 6016 -2494 6046 -2476
rect 6109 -2476 6217 -2475
rect 6109 -2480 6139 -2476
rect 6147 -2478 6179 -2476
rect 6187 -2480 6217 -2476
rect 6280 -2494 6310 -2462
rect 6338 -2476 6351 -2462
rect 6366 -2480 6396 -2462
rect 6439 -2524 6452 -2462
use 10T_4x4_magic  10T_4x4_magic_0
timestamp 1668471109
transform 1 0 -487 0 1 1570
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_1
timestamp 1668471109
transform 1 0 -487 0 1 1030
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_2
timestamp 1668471109
transform 1 0 -487 0 1 490
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_3
timestamp 1668471109
transform 1 0 673 0 1 -1670
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_4
timestamp 1668471109
transform 1 0 673 0 1 -2210
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_5
timestamp 1668471109
transform 1 0 673 0 1 -1130
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_6
timestamp 1668471109
transform 1 0 673 0 1 -590
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_7
timestamp 1668471109
transform 1 0 673 0 1 -50
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_8
timestamp 1668471109
transform 1 0 673 0 1 490
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_9
timestamp 1668471109
transform 1 0 -487 0 1 -50
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_10
timestamp 1668471109
transform 1 0 -487 0 1 -590
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_11
timestamp 1668471109
transform 1 0 -487 0 1 -1130
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_12
timestamp 1668471109
transform 1 0 673 0 1 1030
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_13
timestamp 1668471109
transform 1 0 -487 0 1 -1670
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_14
timestamp 1668471109
transform 1 0 -487 0 1 -2210
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_15
timestamp 1668471109
transform 1 0 673 0 1 1570
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_16
timestamp 1668471109
transform 1 0 1833 0 1 -1670
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_17
timestamp 1668471109
transform 1 0 1833 0 1 -2210
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_18
timestamp 1668471109
transform 1 0 2993 0 1 -1670
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_19
timestamp 1668471109
transform 1 0 2993 0 1 -2210
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_20
timestamp 1668471109
transform 1 0 1833 0 1 -1130
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_21
timestamp 1668471109
transform 1 0 2993 0 1 -1130
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_22
timestamp 1668471109
transform 1 0 1833 0 1 -590
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_23
timestamp 1668471109
transform 1 0 2993 0 1 -590
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_24
timestamp 1668471109
transform 1 0 1833 0 1 -50
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_25
timestamp 1668471109
transform 1 0 2993 0 1 -50
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_26
timestamp 1668471109
transform 1 0 1833 0 1 490
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_27
timestamp 1668471109
transform 1 0 2993 0 1 490
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_28
timestamp 1668471109
transform 1 0 1833 0 1 1570
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_29
timestamp 1668471109
transform 1 0 1833 0 1 1030
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_30
timestamp 1668471109
transform 1 0 2993 0 1 1570
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_31
timestamp 1668471109
transform 1 0 2993 0 1 1030
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_32
timestamp 1668471109
transform 1 0 4153 0 1 -1670
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_33
timestamp 1668471109
transform 1 0 4153 0 1 -2210
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_34
timestamp 1668471109
transform 1 0 5313 0 1 -1670
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_35
timestamp 1668471109
transform 1 0 5313 0 1 -2210
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_36
timestamp 1668471109
transform 1 0 4153 0 1 -1130
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_37
timestamp 1668471109
transform 1 0 4153 0 1 -590
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_38
timestamp 1668471109
transform 1 0 4153 0 1 -50
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_39
timestamp 1668471109
transform 1 0 5313 0 1 -1130
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_40
timestamp 1668471109
transform 1 0 5313 0 1 -590
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_41
timestamp 1668471109
transform 1 0 5313 0 1 -50
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_42
timestamp 1668471109
transform 1 0 4153 0 1 490
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_43
timestamp 1668471109
transform 1 0 4153 0 1 1570
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_44
timestamp 1668471109
transform 1 0 4153 0 1 1030
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_45
timestamp 1668471109
transform 1 0 5313 0 1 490
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_46
timestamp 1668471109
transform 1 0 5313 0 1 1570
box -54 -314 1153 322
use 10T_4x4_magic  10T_4x4_magic_47
timestamp 1668471109
transform 1 0 5313 0 1 1030
box -54 -314 1153 322
<< end >>
