*
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/models.all"

.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/tt_discrete.cor"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/ttcell.cor"

.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/npd.pm3"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/npass.pm3"
.include "/home/tdene/Public/skywater-src-nda/s8_spice_models/ppu.pm3"

*** Define power and ground
vvdd vdd 0 DC 1.8V
vgnd gnd 0 DC 0V

vin in gnd pulse 0 1.8V 0ns 750ps 750ps 14.8ns 30ns

M1000 out in vdd vdd ppu w=0.14 l=0.15
+  ad=0.3339 pd=3.05 as=0.3339 ps=3.05
*M1001 out in gnd gnd npass w=0.14 l=0.15
M1001 out in gnd gnd npd w=0.21 l=0.15
+  ad=0.1378 pd=1.57 as=0.1378 ps=1.57

C1 out gnd 100fF

.tran 1ns 45ns

.print DC V(in) V(out) 
.print tran V(in) V(out)
.probe V(in) V(out)
.op
.options probe post measout captab
.end

