* FILE: 12Tcell.sp

********************** begin header *****************************

* SPICE Header file for TSMC 3.3 0.35 process (scn4me_subm)

.OPTIONS post NOMOD probe measout captab 

**################################################
* Only Typical/Typical spice models included
.include '/programs/micromagic/mmi_local/ami05.mod'
**################################################

.param ln_min   =  0.4u
.param lp_min   =  0.4u

.PARAM vddp=3.30	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 25
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "12Tcell" generated by MMI_SUE5.6.37 on Fri Nov 12 
*+ 13:58:42 CST 2021.

* start main CELL 12Tcell
* .SUBCKT 12Tcell BL BR WWLA WWLB 
M_1 net_6 net_8 BL gnd n W='0.42*1u' L='0.15*1u' 
M_2 net_1 WWLA net_6 gnd n W='0.42*1u' L='0.15*1u' 
M_3 BR net_8 net_7 gnd n W='0.42*1u' L='0.15*1u' 
M_4 net_7 WWLB net_2 gnd n W='0.42*1u' L='0.15*1u' 
M_5 net_4 net_1 net_6 gnd n W='0.42*1u' L='0.15*1u' 
M_6 net_7 net_2 net_4 gnd n W='0.42*1u' L='0.15*1u' 
M_7 net_3 net_1 vdd vdd p W='0.42*1u' L='0.15*1u' 
M_8 vdd net_2 net_5 vdd p W='0.42*1u' L='0.15*1u' 
M_9 net_1 WWLA net_5 vdd p W='0.42*1u' L='0.15*1u' 
M_10 net_3 WWLB net_2 vdd p W='0.42*1u' L='0.15*1u' 
M_11 gnd net_2 net_1 gnd n W='0.42*1u' L='0.15*1u' 
M_12 net_2 net_1 gnd gnd n W='0.42*1u' L='0.15*1u' 
* .ENDS	$ 12Tcell

.GLOBAL gnd vdd

.END

