magic
tech sky130A
magscale 1 2
timestamp 1653511563
<< error_p >>
rect 38 376 66 388
rect 38 370 68 376
rect 14 357 90 370
rect 14 342 72 357
rect 22 341 82 342
rect 66 338 68 341
rect -18 334 38 338
rect 66 334 122 338
rect -18 308 122 334
rect 174 329 211 342
rect 152 316 226 329
rect 152 308 211 316
rect 66 292 68 308
rect 84 296 100 308
rect 102 296 118 308
rect 152 304 182 308
rect 203 304 211 308
rect 152 301 211 304
rect 161 300 221 301
rect 84 292 118 296
rect 174 292 211 300
rect 24 279 38 292
rect 66 282 258 292
rect 66 279 104 282
rect 0 276 104 279
rect 0 273 80 276
rect -12 271 80 273
rect -16 245 80 271
rect 84 275 104 276
rect 108 276 258 282
rect 108 275 118 276
rect 84 262 118 275
rect 127 262 258 276
rect 168 260 211 262
rect 168 257 213 260
rect 167 251 219 257
rect 240 251 266 254
rect -16 241 0 245
rect 14 242 80 245
rect 14 241 61 242
rect 66 241 80 242
rect 14 227 30 241
rect 1 191 30 227
rect 0 190 30 191
rect -2 174 30 190
rect 38 217 80 241
rect 144 236 266 251
rect 107 217 123 228
rect 125 221 141 228
rect 144 221 148 236
rect 166 221 170 236
rect 125 217 148 221
rect 38 174 68 217
rect 69 212 80 217
rect 138 216 148 217
rect 107 212 148 216
rect 174 212 211 236
rect 91 196 98 212
rect 107 202 157 212
rect 107 192 118 202
rect 138 192 157 202
rect 107 182 157 192
rect 174 200 204 212
rect 174 182 188 200
rect 138 175 148 182
rect -2 172 38 174
rect -16 167 38 172
rect -16 149 34 167
rect -16 142 38 149
rect -2 126 30 142
rect 0 125 30 126
rect 1 99 30 125
rect 38 129 68 142
rect 69 134 80 172
rect 107 166 123 175
rect 125 166 148 175
rect 174 174 180 182
rect 174 172 188 174
rect 107 141 123 150
rect 138 138 148 166
rect 172 142 188 172
rect 195 142 198 200
rect 202 174 204 200
rect 240 191 312 236
rect 226 190 312 191
rect 224 175 312 190
rect 223 174 312 175
rect 202 167 312 174
rect 204 149 312 167
rect 202 142 312 149
rect 174 138 188 142
rect 202 138 204 142
rect 223 141 312 142
rect 224 138 312 141
rect 38 99 80 129
rect 91 104 102 134
rect 107 124 312 138
rect 107 114 118 124
rect 138 114 312 124
rect 107 104 312 114
rect 138 99 312 104
rect 1 89 80 99
rect 14 70 80 89
rect 107 88 123 99
rect 125 88 312 99
rect 138 83 312 88
rect 14 69 89 70
rect 1 61 89 69
rect 38 58 89 61
rect 138 67 209 83
rect 38 54 107 58
rect 138 57 218 67
rect 138 54 202 57
rect 207 55 218 57
rect 24 51 38 54
rect 66 51 107 54
rect 16 40 107 51
rect 123 40 174 54
rect 16 28 174 40
rect 176 28 204 34
rect 207 28 258 54
rect 16 24 258 28
rect 66 9 68 24
rect 73 9 89 24
rect 91 9 107 24
rect 146 15 226 24
rect -18 -11 38 9
rect 66 -11 122 9
rect 146 8 182 15
rect 199 8 210 15
rect 146 0 210 8
rect 160 -1 220 0
rect -18 -21 122 -11
rect 12 -30 90 -21
rect 174 -26 207 -1
rect 12 -37 46 -30
rect 58 -37 72 -30
rect 12 -45 72 -37
rect 22 -46 82 -45
rect 38 -71 66 -46
<< nwell >>
rect 144 83 240 236
<< pwell >>
rect 12 263 92 357
rect 177 301 205 316
rect 12 257 106 263
rect 0 200 106 257
rect 179 245 207 260
rect -26 116 106 200
rect 0 61 106 116
rect 12 53 106 61
rect 175 57 206 67
rect 12 -45 92 53
rect 176 0 204 15
<< nmos >>
rect 38 308 66 338
rect 174 262 211 292
rect 174 24 207 54
rect 38 -21 66 9
<< npd >>
rect 38 182 80 212
rect 38 104 80 134
<< npass >>
rect 38 262 66 292
rect 38 24 66 54
<< ppu >>
rect 174 182 202 212
rect 174 104 202 134
<< ndiff >>
rect 38 338 66 342
rect 38 292 66 308
rect 174 301 177 316
rect 205 301 211 316
rect 174 292 211 301
rect 38 255 66 262
rect 0 241 66 255
rect 174 260 211 262
rect 174 245 179 260
rect 207 245 211 260
rect 174 243 211 245
rect 0 174 14 241
tri 61 220 71 230 se
rect 71 220 80 237
rect 38 212 80 220
rect 38 174 80 182
rect 14 142 80 174
rect 0 75 14 142
rect 38 134 80 142
rect 38 96 80 104
rect 70 79 80 96
rect 0 61 66 75
rect 38 54 66 61
rect 174 67 207 70
rect 174 57 175 67
rect 206 57 207 67
rect 174 54 207 57
rect 38 9 66 24
rect 174 15 207 24
rect 174 0 176 15
rect 204 0 207 15
rect 38 -30 66 -21
<< pdiff >>
rect 174 212 202 221
rect 174 174 202 182
rect 174 142 226 174
rect 174 134 202 142
rect 174 95 202 104
tri 174 83 186 95 nw
<< ndiffc >>
rect 38 342 66 357
rect 177 301 205 316
rect 179 245 207 260
rect 38 230 71 237
rect 38 220 61 230
tri 61 220 71 230 nw
rect 0 142 14 174
rect 38 79 70 96
rect 175 57 206 67
rect 176 0 204 15
rect 38 -45 66 -30
<< pdiffc >>
rect 174 221 202 236
rect 226 142 240 174
tri 174 83 186 95 se
rect 186 83 202 95
<< poly >>
rect 16 308 38 338
rect 66 308 84 338
rect 16 262 38 292
rect 66 262 84 292
rect 152 262 174 292
rect 211 262 270 292
rect 16 182 38 212
rect 80 182 107 212
rect 141 182 174 212
rect 202 182 224 212
rect 16 104 38 134
rect 80 104 107 134
rect 141 104 174 134
rect 202 104 224 134
rect 240 54 270 262
rect 16 24 38 54
rect 66 24 73 54
rect 146 24 174 54
rect 207 24 270 54
rect 16 -21 38 9
rect 66 -21 82 9
<< polycont >>
rect 84 262 118 292
rect 107 182 141 212
rect 107 104 141 134
rect 73 24 107 54
<< locali >>
rect 66 342 68 357
rect 15 255 67 260
rect 14 245 67 255
rect 174 245 179 255
rect 14 241 22 245
rect 39 242 67 245
rect 38 237 66 240
rect 174 236 202 245
rect 38 75 66 78
rect 14 65 66 75
rect 38 62 66 65
rect 174 67 202 83
rect 174 61 175 67
rect 66 -45 68 -30
<< corelocali >>
rect 14 342 38 357
rect 68 342 90 357
rect 152 301 177 316
rect 205 301 226 316
rect 14 262 84 273
rect 118 262 226 273
rect 14 260 226 262
rect 14 255 15 260
rect 67 255 179 260
rect 67 245 174 255
rect 207 245 226 260
rect 22 242 39 245
rect 67 242 71 245
rect 22 241 71 242
rect 14 240 71 241
rect 14 220 38 240
rect 66 237 71 240
tri 71 230 86 245 nw
rect 170 221 174 245
rect 202 221 226 245
rect 14 219 60 220
tri 60 219 61 220 nw
rect 170 219 226 221
rect 0 174 14 191
tri 63 182 98 217 se
rect 98 212 142 217
rect 98 182 107 212
rect 141 182 142 212
rect 0 125 14 142
tri 42 161 63 182 se
rect 63 175 142 182
rect 63 161 70 175
rect 42 97 70 161
tri 70 149 96 175 nw
tri 160 149 170 159 se
rect 170 149 198 219
rect 226 175 240 191
tri 152 141 160 149 se
rect 160 147 198 149
rect 160 141 170 147
rect 102 134 170 141
rect 102 104 107 134
rect 141 119 170 134
tri 170 119 198 147 nw
rect 226 125 240 141
rect 141 104 150 119
rect 102 99 150 104
tri 150 99 170 119 nw
rect 14 96 70 97
rect 14 79 38 96
tri 186 95 188 97 se
rect 188 95 226 97
rect 14 78 70 79
rect 14 75 38 78
rect 66 71 70 78
tri 162 71 174 83 se
rect 14 62 38 65
rect 66 62 174 71
rect 202 67 226 95
rect 14 61 174 62
rect 14 57 175 61
rect 206 57 226 67
rect 14 54 226 57
rect 14 43 73 54
rect 107 43 226 54
rect 146 0 176 15
rect 204 0 226 15
rect 12 -45 38 -30
rect 68 -45 90 -30
<< viali >>
rect 223 174 240 175
rect 223 142 226 174
rect 226 142 240 174
rect 223 141 240 142
<< labels >>
rlabel space 16 182 224 212 1 INV1
rlabel space 16 104 224 134 1 INV2
rlabel space 168 24 240 54 1 left_N
rlabel space 168 262 240 292 1 right_N
rlabel poly 240 24 270 292 1 WWl
rlabel space 146 0 226 15 1 WBL
rlabel space 152 301 232 316 1 WBLb
rlabel ndiffc 38 -45 66 -30 1 RBL0
rlabel nmos 38 -21 66 9 1 RWL0
rlabel ndiffc 38 342 66 357 1 RBL1
rlabel nmos 38 308 66 338 1 RWL1
<< end >>
