magic
tech sky130A
magscale 1 2
timestamp 1606864424
<< checkpaint >>
rect -1269 2461 1459 2601
rect -1760 -1129 6260 2461
rect -1269 -1260 1459 -1129
<< nwell >>
rect -9 485 199 897
<< nmos >>
rect 80 115 110 219
<< pmos >>
rect 80 521 110 773
<< ndiff >>
rect 27 171 80 219
rect 27 131 35 171
rect 69 131 80 171
rect 27 115 80 131
rect 110 171 163 219
rect 110 131 121 171
rect 155 131 163 171
rect 110 115 163 131
<< pdiff >>
rect 27 757 80 773
rect 27 697 35 757
rect 69 697 80 757
rect 27 521 80 697
rect 110 757 163 773
rect 110 561 121 757
rect 155 561 163 757
rect 110 521 163 561
<< ndiffc >>
rect 35 131 69 171
rect 121 131 155 171
<< pdiffc >>
rect 35 697 69 757
rect 121 561 155 757
<< psubdiff >>
rect 27 27 51 61
rect 85 27 109 61
<< nsubdiff >>
rect 27 827 51 861
rect 85 827 109 861
<< psubdiffcont >>
rect 51 27 85 61
<< nsubdiffcont >>
rect 51 827 85 861
<< poly >>
rect 80 773 110 799
rect 80 398 110 521
rect 80 382 134 398
rect 80 348 90 382
rect 124 348 134 382
rect 80 332 134 348
rect 80 219 110 332
rect 80 89 110 115
<< polycont >>
rect 90 348 124 382
<< locali >>
rect 0 867 198 888
rect 0 827 51 867
rect 85 827 198 867
rect 35 757 69 827
rect 35 681 69 697
rect 121 757 155 773
rect 47 382 81 553
rect 121 513 155 561
rect 47 348 90 382
rect 124 348 140 382
rect 35 171 69 187
rect 35 61 69 131
rect 121 171 155 183
rect 121 115 155 131
rect 0 21 51 61
rect 85 21 198 61
rect 0 0 198 21
<< viali >>
rect 51 861 85 867
rect 51 833 85 861
rect 47 553 81 587
rect 121 479 155 513
rect 121 183 155 217
rect 51 27 85 55
rect 51 21 85 27
<< metal1 >>
rect 0 867 198 888
rect 0 833 51 867
rect 85 833 198 867
rect 0 827 198 833
rect 35 587 93 593
rect 35 553 47 587
rect 81 553 127 587
rect 35 547 93 553
rect 109 513 167 519
rect 109 479 121 513
rect 155 479 167 513
rect 109 473 167 479
rect 121 223 155 473
rect 109 217 167 223
rect 109 183 121 217
rect 155 183 167 217
rect 109 177 167 183
rect 0 55 198 61
rect 0 21 51 55
rect 85 21 198 55
rect 0 0 198 21
<< labels >>
rlabel metal1 151 345 151 345 1 Y
port 1 n
rlabel viali 64 570 64 570 1 A
port 2 n
rlabel viali 68 48 68 48 1 gnd
rlabel viali 68 840 68 840 1 vdd
<< end >>
