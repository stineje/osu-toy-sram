VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO 10T_16x12_2r1w_magic_flattened
  CLASS CORE ;
  ORIGIN 0.455 0.275 ;
  FOREIGN 10T_16x12_2r1w_magic_flattened -0.455 -0.275 ;
  SIZE 35.215 BY 22.085 ;
  SYMMETRY X Y ;
  SITE 12T ;
  PIN RBL0_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_0
  PIN RBL0_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_1
  PIN RBL0_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_10
  PIN RBL0_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_11
  PIN RBL0_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_2
  PIN RBL0_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_3
  PIN RBL0_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_4
  PIN RBL0_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_5
  PIN RBL0_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_6
  PIN RBL0_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_7
  PIN RBL0_8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_8
  PIN RBL0_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL0_9
  PIN RBL1_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_0
  PIN RBL1_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_1
  PIN RBL1_10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_10
  PIN RBL1_11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_11
  PIN RBL1_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_2
  PIN RBL1_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_3
  PIN RBL1_4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_4
  PIN RBL1_5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_5
  PIN RBL1_6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_6
  PIN RBL1_7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_7
  PIN RBL1_8
    DIRECTION INPUT ;
    USE SIGNAL ;
  END RBL1_8
  PIN RBL1_9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
  END RBL1_9
  PIN WBL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_0
  PIN WBL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_1
  PIN WBL_10
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_10
  PIN WBL_11
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_11
  PIN WBL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_2
  PIN WBL_3
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_3
  PIN WBL_4
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_4
  PIN WBL_5
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_5
  PIN WBL_6
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_6
  PIN WBL_7
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_7
  PIN WBL_8
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_8
  PIN WBL_9
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBL_9
  PIN WBLb_0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_0
  PIN WBLb_1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_1
  PIN WBLb_10
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_10
  PIN WBLb_11
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_11
  PIN WBLb_2
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_2
  PIN WBLb_3
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_3
  PIN WBLb_4
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_4
  PIN WBLb_5
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_5
  PIN WBLb_6
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_6
  PIN WBLb_7
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_7
  PIN WBLb_8
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_8
  PIN WBLb_9
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WBLb_9
  PIN WWL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_0
  PIN WWL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_1
  PIN WWL_10
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_10
  PIN WWL_11
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_11
  PIN WWL_12
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_12
  PIN WWL_13
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_13
  PIN WWL_14
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_14
  PIN WWL_15
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_15
  PIN WWL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_2
  PIN WWL_3
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_3
  PIN WWL_4
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_4
  PIN WWL_5
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_5
  PIN WWL_6
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_6
  PIN WWL_7
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_7
  PIN WWL_8
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_8
  PIN WWL_9
    DIRECTION INPUT ;
    USE SIGNAL ;
  END WWL_9
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.455 -0.035 34.625 0.035 ;
        RECT -0.455 1.315 34.625 1.385 ;
        RECT -0.455 2.665 34.625 2.735 ;
        RECT -0.455 4.015 34.625 4.085 ;
        RECT -0.455 5.365 34.625 5.435 ;
        RECT -0.455 6.715 34.625 6.785 ;
        RECT -0.455 8.065 34.625 8.135 ;
        RECT -0.455 9.415 34.625 9.485 ;
        RECT -0.455 10.765 34.625 10.835 ;
        RECT -0.455 12.115 34.625 12.185 ;
        RECT -0.455 13.465 34.625 13.535 ;
        RECT -0.455 14.815 34.625 14.885 ;
        RECT -0.455 16.165 34.625 16.235 ;
        RECT -0.455 17.515 34.625 17.585 ;
        RECT -0.455 18.865 34.625 18.935 ;
        RECT -0.455 20.215 34.625 20.285 ;
    END
  END GND
  PIN RWL1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 0.475 34.76 0.67 ;
        RECT 34.53 0.62 34.71 0.715 ;
        RECT 34.6 0.55 34.76 0.67 ;
        RECT 34.67 0.495 34.71 0.715 ;
        RECT 34.46 0.69 34.67 0.77 ;
        RECT 34.41 0.75 34.6 0.84 ;
        RECT 34.17 0.775 34.53 0.91 ;
        RECT 34.21 0.775 34.46 0.945 ;
        RECT 34.03 0.75 34.26 0.8 ;
        RECT 34.03 0.705 34.21 0.8 ;
        RECT 34.17 0.775 34.46 0.925 ;
        RECT 33.96 0.65 34.17 0.73 ;
        RECT 34.1 0.775 34.53 0.87 ;
        RECT 33.91 0.58 34.1 0.67 ;
        RECT 31.7 0.55 34.03 0.645 ;
        RECT 31.77 0.51 34.03 0.645 ;
        RECT 31.77 0.495 33.96 0.645 ;
        RECT 31.81 0.475 33.96 0.645 ;
        RECT 31.63 0.62 31.86 0.67 ;
        RECT 31.63 0.62 31.81 0.715 ;
        RECT 31.56 0.69 31.77 0.77 ;
        RECT 31.51 0.75 31.7 0.84 ;
        RECT 31.27 0.775 31.63 0.91 ;
        RECT 31.31 0.775 31.56 0.945 ;
        RECT 31.13 0.75 31.36 0.8 ;
        RECT 31.13 0.705 31.31 0.8 ;
        RECT 31.27 0.775 31.56 0.925 ;
        RECT 31.06 0.65 31.27 0.73 ;
        RECT 31.2 0.775 31.63 0.87 ;
        RECT 31.01 0.58 31.2 0.67 ;
        RECT 28.725 0.51 31.13 0.645 ;
        RECT 28.725 0.475 31.06 0.645 ;
        RECT 28.74 0.475 28.96 0.65 ;
        RECT 28.74 0.475 28.95 0.69 ;
        RECT 28.3 0.775 28.74 0.87 ;
        RECT 28.61 0.75 28.81 0.83 ;
        RECT 28.73 0.65 28.74 0.87 ;
        RECT 28.37 0.775 28.73 0.91 ;
        RECT 28.66 0.69 28.88 0.76 ;
        RECT 28.41 0.775 28.66 0.945 ;
        RECT 28.23 0.75 28.46 0.8 ;
        RECT 28.23 0.705 28.41 0.8 ;
        RECT 28.37 0.775 28.66 0.925 ;
        RECT 28.16 0.65 28.37 0.73 ;
        RECT 28.11 0.58 28.3 0.67 ;
        RECT 25.9 0.55 28.23 0.645 ;
        RECT 25.97 0.51 28.23 0.645 ;
        RECT 25.97 0.495 28.16 0.645 ;
        RECT 26.01 0.475 28.16 0.645 ;
        RECT 25.83 0.62 26.06 0.67 ;
        RECT 25.83 0.62 26.01 0.715 ;
        RECT 25.76 0.69 25.97 0.77 ;
        RECT 25.71 0.75 25.9 0.84 ;
        RECT 25.47 0.775 25.83 0.91 ;
        RECT 25.51 0.775 25.76 0.945 ;
        RECT 25.33 0.75 25.56 0.8 ;
        RECT 25.33 0.705 25.51 0.8 ;
        RECT 25.47 0.775 25.76 0.925 ;
        RECT 25.26 0.65 25.47 0.73 ;
        RECT 25.4 0.775 25.83 0.87 ;
        RECT 25.21 0.58 25.4 0.67 ;
        RECT 22.925 0.51 25.33 0.645 ;
        RECT 22.925 0.475 25.26 0.645 ;
        RECT 22.94 0.475 23.16 0.65 ;
        RECT 22.94 0.475 23.15 0.69 ;
        RECT 22.5 0.775 22.94 0.87 ;
        RECT 22.81 0.75 23.01 0.83 ;
        RECT 22.93 0.65 22.94 0.87 ;
        RECT 22.57 0.775 22.93 0.91 ;
        RECT 22.86 0.69 23.08 0.76 ;
        RECT 22.61 0.775 22.86 0.945 ;
        RECT 22.43 0.75 22.66 0.8 ;
        RECT 22.43 0.705 22.61 0.8 ;
        RECT 22.57 0.775 22.86 0.925 ;
        RECT 22.36 0.65 22.57 0.73 ;
        RECT 22.31 0.58 22.5 0.67 ;
        RECT 20.1 0.55 22.43 0.645 ;
        RECT 20.17 0.51 22.43 0.645 ;
        RECT 20.17 0.495 22.36 0.645 ;
        RECT 20.21 0.475 22.36 0.645 ;
        RECT 20.03 0.62 20.26 0.67 ;
        RECT 20.03 0.62 20.21 0.715 ;
        RECT 19.96 0.69 20.17 0.77 ;
        RECT 19.91 0.75 20.1 0.84 ;
        RECT 19.67 0.775 20.03 0.91 ;
        RECT 19.71 0.775 19.96 0.945 ;
        RECT 19.53 0.75 19.76 0.8 ;
        RECT 19.53 0.705 19.71 0.8 ;
        RECT 19.67 0.775 19.96 0.925 ;
        RECT 19.46 0.65 19.67 0.73 ;
        RECT 19.6 0.775 20.03 0.87 ;
        RECT 19.41 0.58 19.6 0.67 ;
        RECT 17.125 0.51 19.53 0.645 ;
        RECT 17.125 0.475 19.46 0.645 ;
        RECT 17.14 0.475 17.36 0.65 ;
        RECT 17.14 0.475 17.35 0.69 ;
        RECT 16.7 0.775 17.14 0.87 ;
        RECT 17.01 0.75 17.21 0.83 ;
        RECT 17.13 0.65 17.14 0.87 ;
        RECT 16.77 0.775 17.13 0.91 ;
        RECT 17.06 0.69 17.28 0.76 ;
        RECT 16.81 0.775 17.06 0.945 ;
        RECT 16.63 0.75 16.86 0.8 ;
        RECT 16.63 0.705 16.81 0.8 ;
        RECT 16.77 0.775 17.06 0.925 ;
        RECT 16.56 0.65 16.77 0.73 ;
        RECT 16.51 0.58 16.7 0.67 ;
        RECT 14.3 0.55 16.63 0.645 ;
        RECT 14.37 0.51 16.63 0.645 ;
        RECT 14.37 0.495 16.56 0.645 ;
        RECT 14.41 0.475 16.56 0.645 ;
        RECT 14.23 0.62 14.46 0.67 ;
        RECT 14.23 0.62 14.41 0.715 ;
        RECT 14.16 0.69 14.37 0.77 ;
        RECT 14.11 0.75 14.3 0.84 ;
        RECT 13.87 0.775 14.23 0.91 ;
        RECT 13.91 0.775 14.16 0.945 ;
        RECT 13.73 0.75 13.96 0.8 ;
        RECT 13.73 0.705 13.91 0.8 ;
        RECT 13.87 0.775 14.16 0.925 ;
        RECT 13.66 0.65 13.87 0.73 ;
        RECT 13.8 0.775 14.23 0.87 ;
        RECT 13.61 0.58 13.8 0.67 ;
        RECT 11.325 0.51 13.73 0.645 ;
        RECT 11.325 0.475 13.66 0.645 ;
        RECT 11.34 0.475 11.56 0.65 ;
        RECT 11.34 0.475 11.55 0.69 ;
        RECT 10.9 0.775 11.34 0.87 ;
        RECT 11.21 0.75 11.41 0.83 ;
        RECT 11.33 0.65 11.34 0.87 ;
        RECT 10.97 0.775 11.33 0.91 ;
        RECT 11.26 0.69 11.48 0.76 ;
        RECT 11.01 0.775 11.26 0.945 ;
        RECT 10.83 0.75 11.06 0.8 ;
        RECT 10.83 0.705 11.01 0.8 ;
        RECT 10.97 0.775 11.26 0.925 ;
        RECT 10.76 0.65 10.97 0.73 ;
        RECT 10.71 0.58 10.9 0.67 ;
        RECT 8.5 0.55 10.83 0.645 ;
        RECT 8.57 0.51 10.83 0.645 ;
        RECT 8.57 0.495 10.76 0.645 ;
        RECT 8.61 0.475 10.76 0.645 ;
        RECT 8.43 0.62 8.66 0.67 ;
        RECT 8.43 0.62 8.61 0.715 ;
        RECT 8.36 0.69 8.57 0.77 ;
        RECT 8.31 0.75 8.5 0.84 ;
        RECT 8.07 0.775 8.43 0.91 ;
        RECT 8.11 0.775 8.36 0.945 ;
        RECT 7.93 0.75 8.16 0.8 ;
        RECT 7.93 0.705 8.11 0.8 ;
        RECT 8.07 0.775 8.36 0.925 ;
        RECT 7.86 0.65 8.07 0.73 ;
        RECT 8 0.775 8.43 0.87 ;
        RECT 7.81 0.58 8 0.67 ;
        RECT 5.525 0.51 7.93 0.645 ;
        RECT 5.525 0.475 7.86 0.645 ;
        RECT 5.54 0.475 5.76 0.65 ;
        RECT 5.54 0.475 5.75 0.69 ;
        RECT 5.1 0.775 5.54 0.87 ;
        RECT 5.41 0.75 5.61 0.83 ;
        RECT 5.53 0.65 5.54 0.87 ;
        RECT 5.17 0.775 5.53 0.91 ;
        RECT 5.46 0.69 5.68 0.76 ;
        RECT 5.21 0.775 5.46 0.945 ;
        RECT 5.03 0.75 5.26 0.8 ;
        RECT 5.03 0.705 5.21 0.8 ;
        RECT 5.17 0.775 5.46 0.925 ;
        RECT 4.96 0.65 5.17 0.73 ;
        RECT 4.91 0.58 5.1 0.67 ;
        RECT 2.7 0.55 5.03 0.645 ;
        RECT 2.77 0.51 5.03 0.645 ;
        RECT 2.77 0.495 4.96 0.645 ;
        RECT 2.81 0.475 4.96 0.645 ;
        RECT 2.63 0.62 2.86 0.67 ;
        RECT 2.63 0.62 2.81 0.715 ;
        RECT 2.56 0.69 2.77 0.77 ;
        RECT 2.51 0.75 2.7 0.84 ;
        RECT 2.27 0.775 2.63 0.91 ;
        RECT 2.31 0.775 2.56 0.945 ;
        RECT 2.13 0.75 2.36 0.8 ;
        RECT 2.13 0.705 2.31 0.8 ;
        RECT 2.27 0.775 2.56 0.925 ;
        RECT 2.06 0.65 2.27 0.73 ;
        RECT 2.2 0.775 2.63 0.87 ;
        RECT 2.01 0.58 2.2 0.67 ;
        RECT -0.455 0.51 2.13 0.645 ;
        RECT -0.455 0.475 2.06 0.645 ;
    END
  END RWL1_0
  PIN RWL1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 1.825 34.76 2.02 ;
        RECT 34.53 1.97 34.71 2.065 ;
        RECT 34.6 1.9 34.76 2.02 ;
        RECT 34.67 1.845 34.71 2.065 ;
        RECT 34.46 2.04 34.67 2.12 ;
        RECT 34.41 2.1 34.6 2.19 ;
        RECT 34.17 2.125 34.53 2.26 ;
        RECT 34.21 2.125 34.46 2.295 ;
        RECT 34.03 2.1 34.26 2.15 ;
        RECT 34.03 2.055 34.21 2.15 ;
        RECT 34.17 2.125 34.46 2.275 ;
        RECT 33.96 2 34.17 2.08 ;
        RECT 34.1 2.125 34.53 2.22 ;
        RECT 33.91 1.93 34.1 2.02 ;
        RECT 31.7 1.9 34.03 1.995 ;
        RECT 31.77 1.86 34.03 1.995 ;
        RECT 31.77 1.845 33.96 1.995 ;
        RECT 31.81 1.825 33.96 1.995 ;
        RECT 31.63 1.97 31.86 2.02 ;
        RECT 31.63 1.97 31.81 2.065 ;
        RECT 31.56 2.04 31.77 2.12 ;
        RECT 31.51 2.1 31.7 2.19 ;
        RECT 31.27 2.125 31.63 2.26 ;
        RECT 31.31 2.125 31.56 2.295 ;
        RECT 31.13 2.1 31.36 2.15 ;
        RECT 31.13 2.055 31.31 2.15 ;
        RECT 31.27 2.125 31.56 2.275 ;
        RECT 31.06 2 31.27 2.08 ;
        RECT 31.2 2.125 31.63 2.22 ;
        RECT 31.01 1.93 31.2 2.02 ;
        RECT 28.725 1.86 31.13 1.995 ;
        RECT 28.725 1.825 31.06 1.995 ;
        RECT 28.74 1.825 28.96 2 ;
        RECT 28.74 1.825 28.95 2.04 ;
        RECT 28.3 2.125 28.74 2.22 ;
        RECT 28.61 2.1 28.81 2.18 ;
        RECT 28.73 2 28.74 2.22 ;
        RECT 28.37 2.125 28.73 2.26 ;
        RECT 28.66 2.04 28.88 2.11 ;
        RECT 28.41 2.125 28.66 2.295 ;
        RECT 28.23 2.1 28.46 2.15 ;
        RECT 28.23 2.055 28.41 2.15 ;
        RECT 28.37 2.125 28.66 2.275 ;
        RECT 28.16 2 28.37 2.08 ;
        RECT 28.11 1.93 28.3 2.02 ;
        RECT 25.9 1.9 28.23 1.995 ;
        RECT 25.97 1.86 28.23 1.995 ;
        RECT 25.97 1.845 28.16 1.995 ;
        RECT 26.01 1.825 28.16 1.995 ;
        RECT 25.83 1.97 26.06 2.02 ;
        RECT 25.83 1.97 26.01 2.065 ;
        RECT 25.76 2.04 25.97 2.12 ;
        RECT 25.71 2.1 25.9 2.19 ;
        RECT 25.47 2.125 25.83 2.26 ;
        RECT 25.51 2.125 25.76 2.295 ;
        RECT 25.33 2.1 25.56 2.15 ;
        RECT 25.33 2.055 25.51 2.15 ;
        RECT 25.47 2.125 25.76 2.275 ;
        RECT 25.26 2 25.47 2.08 ;
        RECT 25.4 2.125 25.83 2.22 ;
        RECT 25.21 1.93 25.4 2.02 ;
        RECT 22.925 1.86 25.33 1.995 ;
        RECT 22.925 1.825 25.26 1.995 ;
        RECT 22.94 1.825 23.16 2 ;
        RECT 22.94 1.825 23.15 2.04 ;
        RECT 22.5 2.125 22.94 2.22 ;
        RECT 22.81 2.1 23.01 2.18 ;
        RECT 22.93 2 22.94 2.22 ;
        RECT 22.57 2.125 22.93 2.26 ;
        RECT 22.86 2.04 23.08 2.11 ;
        RECT 22.61 2.125 22.86 2.295 ;
        RECT 22.43 2.1 22.66 2.15 ;
        RECT 22.43 2.055 22.61 2.15 ;
        RECT 22.57 2.125 22.86 2.275 ;
        RECT 22.36 2 22.57 2.08 ;
        RECT 22.31 1.93 22.5 2.02 ;
        RECT 20.1 1.9 22.43 1.995 ;
        RECT 20.17 1.86 22.43 1.995 ;
        RECT 20.17 1.845 22.36 1.995 ;
        RECT 20.21 1.825 22.36 1.995 ;
        RECT 20.03 1.97 20.26 2.02 ;
        RECT 20.03 1.97 20.21 2.065 ;
        RECT 19.96 2.04 20.17 2.12 ;
        RECT 19.91 2.1 20.1 2.19 ;
        RECT 19.67 2.125 20.03 2.26 ;
        RECT 19.71 2.125 19.96 2.295 ;
        RECT 19.53 2.1 19.76 2.15 ;
        RECT 19.53 2.055 19.71 2.15 ;
        RECT 19.67 2.125 19.96 2.275 ;
        RECT 19.46 2 19.67 2.08 ;
        RECT 19.6 2.125 20.03 2.22 ;
        RECT 19.41 1.93 19.6 2.02 ;
        RECT 17.125 1.86 19.53 1.995 ;
        RECT 17.125 1.825 19.46 1.995 ;
        RECT 17.14 1.825 17.36 2 ;
        RECT 17.14 1.825 17.35 2.04 ;
        RECT 16.7 2.125 17.14 2.22 ;
        RECT 17.01 2.1 17.21 2.18 ;
        RECT 17.13 2 17.14 2.22 ;
        RECT 16.77 2.125 17.13 2.26 ;
        RECT 17.06 2.04 17.28 2.11 ;
        RECT 16.81 2.125 17.06 2.295 ;
        RECT 16.63 2.1 16.86 2.15 ;
        RECT 16.63 2.055 16.81 2.15 ;
        RECT 16.77 2.125 17.06 2.275 ;
        RECT 16.56 2 16.77 2.08 ;
        RECT 16.51 1.93 16.7 2.02 ;
        RECT 14.3 1.9 16.63 1.995 ;
        RECT 14.37 1.86 16.63 1.995 ;
        RECT 14.37 1.845 16.56 1.995 ;
        RECT 14.41 1.825 16.56 1.995 ;
        RECT 14.23 1.97 14.46 2.02 ;
        RECT 14.23 1.97 14.41 2.065 ;
        RECT 14.16 2.04 14.37 2.12 ;
        RECT 14.11 2.1 14.3 2.19 ;
        RECT 13.87 2.125 14.23 2.26 ;
        RECT 13.91 2.125 14.16 2.295 ;
        RECT 13.73 2.1 13.96 2.15 ;
        RECT 13.73 2.055 13.91 2.15 ;
        RECT 13.87 2.125 14.16 2.275 ;
        RECT 13.66 2 13.87 2.08 ;
        RECT 13.8 2.125 14.23 2.22 ;
        RECT 13.61 1.93 13.8 2.02 ;
        RECT 11.325 1.86 13.73 1.995 ;
        RECT 11.325 1.825 13.66 1.995 ;
        RECT 11.34 1.825 11.56 2 ;
        RECT 11.34 1.825 11.55 2.04 ;
        RECT 10.9 2.125 11.34 2.22 ;
        RECT 11.21 2.1 11.41 2.18 ;
        RECT 11.33 2 11.34 2.22 ;
        RECT 10.97 2.125 11.33 2.26 ;
        RECT 11.26 2.04 11.48 2.11 ;
        RECT 11.01 2.125 11.26 2.295 ;
        RECT 10.83 2.1 11.06 2.15 ;
        RECT 10.83 2.055 11.01 2.15 ;
        RECT 10.97 2.125 11.26 2.275 ;
        RECT 10.76 2 10.97 2.08 ;
        RECT 10.71 1.93 10.9 2.02 ;
        RECT 8.5 1.9 10.83 1.995 ;
        RECT 8.57 1.86 10.83 1.995 ;
        RECT 8.57 1.845 10.76 1.995 ;
        RECT 8.61 1.825 10.76 1.995 ;
        RECT 8.43 1.97 8.66 2.02 ;
        RECT 8.43 1.97 8.61 2.065 ;
        RECT 8.36 2.04 8.57 2.12 ;
        RECT 8.31 2.1 8.5 2.19 ;
        RECT 8.07 2.125 8.43 2.26 ;
        RECT 8.11 2.125 8.36 2.295 ;
        RECT 7.93 2.1 8.16 2.15 ;
        RECT 7.93 2.055 8.11 2.15 ;
        RECT 8.07 2.125 8.36 2.275 ;
        RECT 7.86 2 8.07 2.08 ;
        RECT 8 2.125 8.43 2.22 ;
        RECT 7.81 1.93 8 2.02 ;
        RECT 5.525 1.86 7.93 1.995 ;
        RECT 5.525 1.825 7.86 1.995 ;
        RECT 5.54 1.825 5.76 2 ;
        RECT 5.54 1.825 5.75 2.04 ;
        RECT 5.1 2.125 5.54 2.22 ;
        RECT 5.41 2.1 5.61 2.18 ;
        RECT 5.53 2 5.54 2.22 ;
        RECT 5.17 2.125 5.53 2.26 ;
        RECT 5.46 2.04 5.68 2.11 ;
        RECT 5.21 2.125 5.46 2.295 ;
        RECT 5.03 2.1 5.26 2.15 ;
        RECT 5.03 2.055 5.21 2.15 ;
        RECT 5.17 2.125 5.46 2.275 ;
        RECT 4.96 2 5.17 2.08 ;
        RECT 4.91 1.93 5.1 2.02 ;
        RECT 2.7 1.9 5.03 1.995 ;
        RECT 2.77 1.86 5.03 1.995 ;
        RECT 2.77 1.845 4.96 1.995 ;
        RECT 2.81 1.825 4.96 1.995 ;
        RECT 2.63 1.97 2.86 2.02 ;
        RECT 2.63 1.97 2.81 2.065 ;
        RECT 2.56 2.04 2.77 2.12 ;
        RECT 2.51 2.1 2.7 2.19 ;
        RECT 2.27 2.125 2.63 2.26 ;
        RECT 2.31 2.125 2.56 2.295 ;
        RECT 2.13 2.1 2.36 2.15 ;
        RECT 2.13 2.055 2.31 2.15 ;
        RECT 2.27 2.125 2.56 2.275 ;
        RECT 2.06 2 2.27 2.08 ;
        RECT 2.2 2.125 2.63 2.22 ;
        RECT 2.01 1.93 2.2 2.02 ;
        RECT -0.455 1.86 2.13 1.995 ;
        RECT -0.455 1.825 2.06 1.995 ;
    END
  END RWL1_1
  PIN RWL1_10
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 13.975 34.76 14.17 ;
        RECT 34.53 14.12 34.71 14.215 ;
        RECT 34.6 14.05 34.76 14.17 ;
        RECT 34.67 13.995 34.71 14.215 ;
        RECT 34.46 14.19 34.67 14.27 ;
        RECT 34.41 14.25 34.6 14.34 ;
        RECT 34.17 14.275 34.53 14.41 ;
        RECT 34.21 14.275 34.46 14.445 ;
        RECT 34.03 14.25 34.26 14.3 ;
        RECT 34.03 14.205 34.21 14.3 ;
        RECT 34.17 14.275 34.46 14.425 ;
        RECT 33.96 14.15 34.17 14.23 ;
        RECT 34.1 14.275 34.53 14.37 ;
        RECT 33.91 14.08 34.1 14.17 ;
        RECT 31.7 14.05 34.03 14.145 ;
        RECT 31.77 14.01 34.03 14.145 ;
        RECT 31.77 13.995 33.96 14.145 ;
        RECT 31.81 13.975 33.96 14.145 ;
        RECT 31.63 14.12 31.86 14.17 ;
        RECT 31.63 14.12 31.81 14.215 ;
        RECT 31.56 14.19 31.77 14.27 ;
        RECT 31.51 14.25 31.7 14.34 ;
        RECT 31.27 14.275 31.63 14.41 ;
        RECT 31.31 14.275 31.56 14.445 ;
        RECT 31.13 14.25 31.36 14.3 ;
        RECT 31.13 14.205 31.31 14.3 ;
        RECT 31.27 14.275 31.56 14.425 ;
        RECT 31.06 14.15 31.27 14.23 ;
        RECT 31.2 14.275 31.63 14.37 ;
        RECT 31.01 14.08 31.2 14.17 ;
        RECT 28.725 14.01 31.13 14.145 ;
        RECT 28.725 13.975 31.06 14.145 ;
        RECT 28.74 13.975 28.96 14.15 ;
        RECT 28.74 13.975 28.95 14.19 ;
        RECT 28.3 14.275 28.74 14.37 ;
        RECT 28.61 14.25 28.81 14.33 ;
        RECT 28.73 14.15 28.74 14.37 ;
        RECT 28.37 14.275 28.73 14.41 ;
        RECT 28.66 14.19 28.88 14.26 ;
        RECT 28.41 14.275 28.66 14.445 ;
        RECT 28.23 14.25 28.46 14.3 ;
        RECT 28.23 14.205 28.41 14.3 ;
        RECT 28.37 14.275 28.66 14.425 ;
        RECT 28.16 14.15 28.37 14.23 ;
        RECT 28.11 14.08 28.3 14.17 ;
        RECT 25.9 14.05 28.23 14.145 ;
        RECT 25.97 14.01 28.23 14.145 ;
        RECT 25.97 13.995 28.16 14.145 ;
        RECT 26.01 13.975 28.16 14.145 ;
        RECT 25.83 14.12 26.06 14.17 ;
        RECT 25.83 14.12 26.01 14.215 ;
        RECT 25.76 14.19 25.97 14.27 ;
        RECT 25.71 14.25 25.9 14.34 ;
        RECT 25.47 14.275 25.83 14.41 ;
        RECT 25.51 14.275 25.76 14.445 ;
        RECT 25.33 14.25 25.56 14.3 ;
        RECT 25.33 14.205 25.51 14.3 ;
        RECT 25.47 14.275 25.76 14.425 ;
        RECT 25.26 14.15 25.47 14.23 ;
        RECT 25.4 14.275 25.83 14.37 ;
        RECT 25.21 14.08 25.4 14.17 ;
        RECT 22.925 14.01 25.33 14.145 ;
        RECT 22.925 13.975 25.26 14.145 ;
        RECT 22.94 13.975 23.16 14.15 ;
        RECT 22.94 13.975 23.15 14.19 ;
        RECT 22.5 14.275 22.94 14.37 ;
        RECT 22.81 14.25 23.01 14.33 ;
        RECT 22.93 14.15 22.94 14.37 ;
        RECT 22.57 14.275 22.93 14.41 ;
        RECT 22.86 14.19 23.08 14.26 ;
        RECT 22.61 14.275 22.86 14.445 ;
        RECT 22.43 14.25 22.66 14.3 ;
        RECT 22.43 14.205 22.61 14.3 ;
        RECT 22.57 14.275 22.86 14.425 ;
        RECT 22.36 14.15 22.57 14.23 ;
        RECT 22.31 14.08 22.5 14.17 ;
        RECT 20.1 14.05 22.43 14.145 ;
        RECT 20.17 14.01 22.43 14.145 ;
        RECT 20.17 13.995 22.36 14.145 ;
        RECT 20.21 13.975 22.36 14.145 ;
        RECT 20.03 14.12 20.26 14.17 ;
        RECT 20.03 14.12 20.21 14.215 ;
        RECT 19.96 14.19 20.17 14.27 ;
        RECT 19.91 14.25 20.1 14.34 ;
        RECT 19.67 14.275 20.03 14.41 ;
        RECT 19.71 14.275 19.96 14.445 ;
        RECT 19.53 14.25 19.76 14.3 ;
        RECT 19.53 14.205 19.71 14.3 ;
        RECT 19.67 14.275 19.96 14.425 ;
        RECT 19.46 14.15 19.67 14.23 ;
        RECT 19.6 14.275 20.03 14.37 ;
        RECT 19.41 14.08 19.6 14.17 ;
        RECT 17.125 14.01 19.53 14.145 ;
        RECT 17.125 13.975 19.46 14.145 ;
        RECT 17.14 13.975 17.36 14.15 ;
        RECT 17.14 13.975 17.35 14.19 ;
        RECT 16.7 14.275 17.14 14.37 ;
        RECT 17.01 14.25 17.21 14.33 ;
        RECT 17.13 14.15 17.14 14.37 ;
        RECT 16.77 14.275 17.13 14.41 ;
        RECT 17.06 14.19 17.28 14.26 ;
        RECT 16.81 14.275 17.06 14.445 ;
        RECT 16.63 14.25 16.86 14.3 ;
        RECT 16.63 14.205 16.81 14.3 ;
        RECT 16.77 14.275 17.06 14.425 ;
        RECT 16.56 14.15 16.77 14.23 ;
        RECT 16.51 14.08 16.7 14.17 ;
        RECT 14.3 14.05 16.63 14.145 ;
        RECT 14.37 14.01 16.63 14.145 ;
        RECT 14.37 13.995 16.56 14.145 ;
        RECT 14.41 13.975 16.56 14.145 ;
        RECT 14.23 14.12 14.46 14.17 ;
        RECT 14.23 14.12 14.41 14.215 ;
        RECT 14.16 14.19 14.37 14.27 ;
        RECT 14.11 14.25 14.3 14.34 ;
        RECT 13.87 14.275 14.23 14.41 ;
        RECT 13.91 14.275 14.16 14.445 ;
        RECT 13.73 14.25 13.96 14.3 ;
        RECT 13.73 14.205 13.91 14.3 ;
        RECT 13.87 14.275 14.16 14.425 ;
        RECT 13.66 14.15 13.87 14.23 ;
        RECT 13.8 14.275 14.23 14.37 ;
        RECT 13.61 14.08 13.8 14.17 ;
        RECT 11.325 14.01 13.73 14.145 ;
        RECT 11.325 13.975 13.66 14.145 ;
        RECT 11.34 13.975 11.56 14.15 ;
        RECT 11.34 13.975 11.55 14.19 ;
        RECT 10.9 14.275 11.34 14.37 ;
        RECT 11.21 14.25 11.41 14.33 ;
        RECT 11.33 14.15 11.34 14.37 ;
        RECT 10.97 14.275 11.33 14.41 ;
        RECT 11.26 14.19 11.48 14.26 ;
        RECT 11.01 14.275 11.26 14.445 ;
        RECT 10.83 14.25 11.06 14.3 ;
        RECT 10.83 14.205 11.01 14.3 ;
        RECT 10.97 14.275 11.26 14.425 ;
        RECT 10.76 14.15 10.97 14.23 ;
        RECT 10.71 14.08 10.9 14.17 ;
        RECT 8.5 14.05 10.83 14.145 ;
        RECT 8.57 14.01 10.83 14.145 ;
        RECT 8.57 13.995 10.76 14.145 ;
        RECT 8.61 13.975 10.76 14.145 ;
        RECT 8.43 14.12 8.66 14.17 ;
        RECT 8.43 14.12 8.61 14.215 ;
        RECT 8.36 14.19 8.57 14.27 ;
        RECT 8.31 14.25 8.5 14.34 ;
        RECT 8.07 14.275 8.43 14.41 ;
        RECT 8.11 14.275 8.36 14.445 ;
        RECT 7.93 14.25 8.16 14.3 ;
        RECT 7.93 14.205 8.11 14.3 ;
        RECT 8.07 14.275 8.36 14.425 ;
        RECT 7.86 14.15 8.07 14.23 ;
        RECT 8 14.275 8.43 14.37 ;
        RECT 7.81 14.08 8 14.17 ;
        RECT 5.525 14.01 7.93 14.145 ;
        RECT 5.525 13.975 7.86 14.145 ;
        RECT 5.54 13.975 5.76 14.15 ;
        RECT 5.54 13.975 5.75 14.19 ;
        RECT 5.1 14.275 5.54 14.37 ;
        RECT 5.41 14.25 5.61 14.33 ;
        RECT 5.53 14.15 5.54 14.37 ;
        RECT 5.17 14.275 5.53 14.41 ;
        RECT 5.46 14.19 5.68 14.26 ;
        RECT 5.21 14.275 5.46 14.445 ;
        RECT 5.03 14.25 5.26 14.3 ;
        RECT 5.03 14.205 5.21 14.3 ;
        RECT 5.17 14.275 5.46 14.425 ;
        RECT 4.96 14.15 5.17 14.23 ;
        RECT 4.91 14.08 5.1 14.17 ;
        RECT 2.7 14.05 5.03 14.145 ;
        RECT 2.77 14.01 5.03 14.145 ;
        RECT 2.77 13.995 4.96 14.145 ;
        RECT 2.81 13.975 4.96 14.145 ;
        RECT 2.63 14.12 2.86 14.17 ;
        RECT 2.63 14.12 2.81 14.215 ;
        RECT 2.56 14.19 2.77 14.27 ;
        RECT 2.51 14.25 2.7 14.34 ;
        RECT 2.27 14.275 2.63 14.41 ;
        RECT 2.31 14.275 2.56 14.445 ;
        RECT 2.13 14.25 2.36 14.3 ;
        RECT 2.13 14.205 2.31 14.3 ;
        RECT 2.27 14.275 2.56 14.425 ;
        RECT 2.06 14.15 2.27 14.23 ;
        RECT 2.2 14.275 2.63 14.37 ;
        RECT 2.01 14.08 2.2 14.17 ;
        RECT -0.455 14.01 2.13 14.145 ;
        RECT -0.455 13.975 2.06 14.145 ;
    END
  END RWL1_10
  PIN RWL1_11
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 15.325 34.76 15.52 ;
        RECT 34.53 15.47 34.71 15.565 ;
        RECT 34.6 15.4 34.76 15.52 ;
        RECT 34.67 15.345 34.71 15.565 ;
        RECT 34.46 15.54 34.67 15.62 ;
        RECT 34.41 15.6 34.6 15.69 ;
        RECT 34.17 15.625 34.53 15.76 ;
        RECT 34.21 15.625 34.46 15.795 ;
        RECT 34.03 15.6 34.26 15.65 ;
        RECT 34.03 15.555 34.21 15.65 ;
        RECT 34.17 15.625 34.46 15.775 ;
        RECT 33.96 15.5 34.17 15.58 ;
        RECT 34.1 15.625 34.53 15.72 ;
        RECT 33.91 15.43 34.1 15.52 ;
        RECT 31.7 15.4 34.03 15.495 ;
        RECT 31.77 15.36 34.03 15.495 ;
        RECT 31.77 15.345 33.96 15.495 ;
        RECT 31.81 15.325 33.96 15.495 ;
        RECT 31.63 15.47 31.86 15.52 ;
        RECT 31.63 15.47 31.81 15.565 ;
        RECT 31.56 15.54 31.77 15.62 ;
        RECT 31.51 15.6 31.7 15.69 ;
        RECT 31.27 15.625 31.63 15.76 ;
        RECT 31.31 15.625 31.56 15.795 ;
        RECT 31.13 15.6 31.36 15.65 ;
        RECT 31.13 15.555 31.31 15.65 ;
        RECT 31.27 15.625 31.56 15.775 ;
        RECT 31.06 15.5 31.27 15.58 ;
        RECT 31.2 15.625 31.63 15.72 ;
        RECT 31.01 15.43 31.2 15.52 ;
        RECT 28.725 15.36 31.13 15.495 ;
        RECT 28.725 15.325 31.06 15.495 ;
        RECT 28.74 15.325 28.96 15.5 ;
        RECT 28.74 15.325 28.95 15.54 ;
        RECT 28.3 15.625 28.74 15.72 ;
        RECT 28.61 15.6 28.81 15.68 ;
        RECT 28.73 15.5 28.74 15.72 ;
        RECT 28.37 15.625 28.73 15.76 ;
        RECT 28.66 15.54 28.88 15.61 ;
        RECT 28.41 15.625 28.66 15.795 ;
        RECT 28.23 15.6 28.46 15.65 ;
        RECT 28.23 15.555 28.41 15.65 ;
        RECT 28.37 15.625 28.66 15.775 ;
        RECT 28.16 15.5 28.37 15.58 ;
        RECT 28.11 15.43 28.3 15.52 ;
        RECT 25.9 15.4 28.23 15.495 ;
        RECT 25.97 15.36 28.23 15.495 ;
        RECT 25.97 15.345 28.16 15.495 ;
        RECT 26.01 15.325 28.16 15.495 ;
        RECT 25.83 15.47 26.06 15.52 ;
        RECT 25.83 15.47 26.01 15.565 ;
        RECT 25.76 15.54 25.97 15.62 ;
        RECT 25.71 15.6 25.9 15.69 ;
        RECT 25.47 15.625 25.83 15.76 ;
        RECT 25.51 15.625 25.76 15.795 ;
        RECT 25.33 15.6 25.56 15.65 ;
        RECT 25.33 15.555 25.51 15.65 ;
        RECT 25.47 15.625 25.76 15.775 ;
        RECT 25.26 15.5 25.47 15.58 ;
        RECT 25.4 15.625 25.83 15.72 ;
        RECT 25.21 15.43 25.4 15.52 ;
        RECT 22.925 15.36 25.33 15.495 ;
        RECT 22.925 15.325 25.26 15.495 ;
        RECT 22.94 15.325 23.16 15.5 ;
        RECT 22.94 15.325 23.15 15.54 ;
        RECT 22.5 15.625 22.94 15.72 ;
        RECT 22.81 15.6 23.01 15.68 ;
        RECT 22.93 15.5 22.94 15.72 ;
        RECT 22.57 15.625 22.93 15.76 ;
        RECT 22.86 15.54 23.08 15.61 ;
        RECT 22.61 15.625 22.86 15.795 ;
        RECT 22.43 15.6 22.66 15.65 ;
        RECT 22.43 15.555 22.61 15.65 ;
        RECT 22.57 15.625 22.86 15.775 ;
        RECT 22.36 15.5 22.57 15.58 ;
        RECT 22.31 15.43 22.5 15.52 ;
        RECT 20.1 15.4 22.43 15.495 ;
        RECT 20.17 15.36 22.43 15.495 ;
        RECT 20.17 15.345 22.36 15.495 ;
        RECT 20.21 15.325 22.36 15.495 ;
        RECT 20.03 15.47 20.26 15.52 ;
        RECT 20.03 15.47 20.21 15.565 ;
        RECT 19.96 15.54 20.17 15.62 ;
        RECT 19.91 15.6 20.1 15.69 ;
        RECT 19.67 15.625 20.03 15.76 ;
        RECT 19.71 15.625 19.96 15.795 ;
        RECT 19.53 15.6 19.76 15.65 ;
        RECT 19.53 15.555 19.71 15.65 ;
        RECT 19.67 15.625 19.96 15.775 ;
        RECT 19.46 15.5 19.67 15.58 ;
        RECT 19.6 15.625 20.03 15.72 ;
        RECT 19.41 15.43 19.6 15.52 ;
        RECT 17.125 15.36 19.53 15.495 ;
        RECT 17.125 15.325 19.46 15.495 ;
        RECT 17.14 15.325 17.36 15.5 ;
        RECT 17.14 15.325 17.35 15.54 ;
        RECT 16.7 15.625 17.14 15.72 ;
        RECT 17.01 15.6 17.21 15.68 ;
        RECT 17.13 15.5 17.14 15.72 ;
        RECT 16.77 15.625 17.13 15.76 ;
        RECT 17.06 15.54 17.28 15.61 ;
        RECT 16.81 15.625 17.06 15.795 ;
        RECT 16.63 15.6 16.86 15.65 ;
        RECT 16.63 15.555 16.81 15.65 ;
        RECT 16.77 15.625 17.06 15.775 ;
        RECT 16.56 15.5 16.77 15.58 ;
        RECT 16.51 15.43 16.7 15.52 ;
        RECT 14.3 15.4 16.63 15.495 ;
        RECT 14.37 15.36 16.63 15.495 ;
        RECT 14.37 15.345 16.56 15.495 ;
        RECT 14.41 15.325 16.56 15.495 ;
        RECT 14.23 15.47 14.46 15.52 ;
        RECT 14.23 15.47 14.41 15.565 ;
        RECT 14.16 15.54 14.37 15.62 ;
        RECT 14.11 15.6 14.3 15.69 ;
        RECT 13.87 15.625 14.23 15.76 ;
        RECT 13.91 15.625 14.16 15.795 ;
        RECT 13.73 15.6 13.96 15.65 ;
        RECT 13.73 15.555 13.91 15.65 ;
        RECT 13.87 15.625 14.16 15.775 ;
        RECT 13.66 15.5 13.87 15.58 ;
        RECT 13.8 15.625 14.23 15.72 ;
        RECT 13.61 15.43 13.8 15.52 ;
        RECT 11.325 15.36 13.73 15.495 ;
        RECT 11.325 15.325 13.66 15.495 ;
        RECT 11.34 15.325 11.56 15.5 ;
        RECT 11.34 15.325 11.55 15.54 ;
        RECT 10.9 15.625 11.34 15.72 ;
        RECT 11.21 15.6 11.41 15.68 ;
        RECT 11.33 15.5 11.34 15.72 ;
        RECT 10.97 15.625 11.33 15.76 ;
        RECT 11.26 15.54 11.48 15.61 ;
        RECT 11.01 15.625 11.26 15.795 ;
        RECT 10.83 15.6 11.06 15.65 ;
        RECT 10.83 15.555 11.01 15.65 ;
        RECT 10.97 15.625 11.26 15.775 ;
        RECT 10.76 15.5 10.97 15.58 ;
        RECT 10.71 15.43 10.9 15.52 ;
        RECT 8.5 15.4 10.83 15.495 ;
        RECT 8.57 15.36 10.83 15.495 ;
        RECT 8.57 15.345 10.76 15.495 ;
        RECT 8.61 15.325 10.76 15.495 ;
        RECT 8.43 15.47 8.66 15.52 ;
        RECT 8.43 15.47 8.61 15.565 ;
        RECT 8.36 15.54 8.57 15.62 ;
        RECT 8.31 15.6 8.5 15.69 ;
        RECT 8.07 15.625 8.43 15.76 ;
        RECT 8.11 15.625 8.36 15.795 ;
        RECT 7.93 15.6 8.16 15.65 ;
        RECT 7.93 15.555 8.11 15.65 ;
        RECT 8.07 15.625 8.36 15.775 ;
        RECT 7.86 15.5 8.07 15.58 ;
        RECT 8 15.625 8.43 15.72 ;
        RECT 7.81 15.43 8 15.52 ;
        RECT 5.525 15.36 7.93 15.495 ;
        RECT 5.525 15.325 7.86 15.495 ;
        RECT 5.54 15.325 5.76 15.5 ;
        RECT 5.54 15.325 5.75 15.54 ;
        RECT 5.1 15.625 5.54 15.72 ;
        RECT 5.41 15.6 5.61 15.68 ;
        RECT 5.53 15.5 5.54 15.72 ;
        RECT 5.17 15.625 5.53 15.76 ;
        RECT 5.46 15.54 5.68 15.61 ;
        RECT 5.21 15.625 5.46 15.795 ;
        RECT 5.03 15.6 5.26 15.65 ;
        RECT 5.03 15.555 5.21 15.65 ;
        RECT 5.17 15.625 5.46 15.775 ;
        RECT 4.96 15.5 5.17 15.58 ;
        RECT 4.91 15.43 5.1 15.52 ;
        RECT 2.7 15.4 5.03 15.495 ;
        RECT 2.77 15.36 5.03 15.495 ;
        RECT 2.77 15.345 4.96 15.495 ;
        RECT 2.81 15.325 4.96 15.495 ;
        RECT 2.63 15.47 2.86 15.52 ;
        RECT 2.63 15.47 2.81 15.565 ;
        RECT 2.56 15.54 2.77 15.62 ;
        RECT 2.51 15.6 2.7 15.69 ;
        RECT 2.27 15.625 2.63 15.76 ;
        RECT 2.31 15.625 2.56 15.795 ;
        RECT 2.13 15.6 2.36 15.65 ;
        RECT 2.13 15.555 2.31 15.65 ;
        RECT 2.27 15.625 2.56 15.775 ;
        RECT 2.06 15.5 2.27 15.58 ;
        RECT 2.2 15.625 2.63 15.72 ;
        RECT 2.01 15.43 2.2 15.52 ;
        RECT -0.455 15.36 2.13 15.495 ;
        RECT -0.455 15.325 2.06 15.495 ;
    END
  END RWL1_11
  PIN RWL1_12
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 16.675 34.76 16.87 ;
        RECT 34.53 16.82 34.71 16.915 ;
        RECT 34.6 16.75 34.76 16.87 ;
        RECT 34.67 16.695 34.71 16.915 ;
        RECT 34.46 16.89 34.67 16.97 ;
        RECT 34.41 16.95 34.6 17.04 ;
        RECT 34.17 16.975 34.53 17.11 ;
        RECT 34.21 16.975 34.46 17.145 ;
        RECT 34.03 16.95 34.26 17 ;
        RECT 34.03 16.905 34.21 17 ;
        RECT 34.17 16.975 34.46 17.125 ;
        RECT 33.96 16.85 34.17 16.93 ;
        RECT 34.1 16.975 34.53 17.07 ;
        RECT 33.91 16.78 34.1 16.87 ;
        RECT 31.7 16.75 34.03 16.845 ;
        RECT 31.77 16.71 34.03 16.845 ;
        RECT 31.77 16.695 33.96 16.845 ;
        RECT 31.81 16.675 33.96 16.845 ;
        RECT 31.63 16.82 31.86 16.87 ;
        RECT 31.63 16.82 31.81 16.915 ;
        RECT 31.56 16.89 31.77 16.97 ;
        RECT 31.51 16.95 31.7 17.04 ;
        RECT 31.27 16.975 31.63 17.11 ;
        RECT 31.31 16.975 31.56 17.145 ;
        RECT 31.13 16.95 31.36 17 ;
        RECT 31.13 16.905 31.31 17 ;
        RECT 31.27 16.975 31.56 17.125 ;
        RECT 31.06 16.85 31.27 16.93 ;
        RECT 31.2 16.975 31.63 17.07 ;
        RECT 31.01 16.78 31.2 16.87 ;
        RECT 28.725 16.71 31.13 16.845 ;
        RECT 28.725 16.675 31.06 16.845 ;
        RECT 28.74 16.675 28.96 16.85 ;
        RECT 28.74 16.675 28.95 16.89 ;
        RECT 28.3 16.975 28.74 17.07 ;
        RECT 28.61 16.95 28.81 17.03 ;
        RECT 28.73 16.85 28.74 17.07 ;
        RECT 28.37 16.975 28.73 17.11 ;
        RECT 28.66 16.89 28.88 16.96 ;
        RECT 28.41 16.975 28.66 17.145 ;
        RECT 28.23 16.95 28.46 17 ;
        RECT 28.23 16.905 28.41 17 ;
        RECT 28.37 16.975 28.66 17.125 ;
        RECT 28.16 16.85 28.37 16.93 ;
        RECT 28.11 16.78 28.3 16.87 ;
        RECT 25.9 16.75 28.23 16.845 ;
        RECT 25.97 16.71 28.23 16.845 ;
        RECT 25.97 16.695 28.16 16.845 ;
        RECT 26.01 16.675 28.16 16.845 ;
        RECT 25.83 16.82 26.06 16.87 ;
        RECT 25.83 16.82 26.01 16.915 ;
        RECT 25.76 16.89 25.97 16.97 ;
        RECT 25.71 16.95 25.9 17.04 ;
        RECT 25.47 16.975 25.83 17.11 ;
        RECT 25.51 16.975 25.76 17.145 ;
        RECT 25.33 16.95 25.56 17 ;
        RECT 25.33 16.905 25.51 17 ;
        RECT 25.47 16.975 25.76 17.125 ;
        RECT 25.26 16.85 25.47 16.93 ;
        RECT 25.4 16.975 25.83 17.07 ;
        RECT 25.21 16.78 25.4 16.87 ;
        RECT 22.925 16.71 25.33 16.845 ;
        RECT 22.925 16.675 25.26 16.845 ;
        RECT 22.94 16.675 23.16 16.85 ;
        RECT 22.94 16.675 23.15 16.89 ;
        RECT 22.5 16.975 22.94 17.07 ;
        RECT 22.81 16.95 23.01 17.03 ;
        RECT 22.93 16.85 22.94 17.07 ;
        RECT 22.57 16.975 22.93 17.11 ;
        RECT 22.86 16.89 23.08 16.96 ;
        RECT 22.61 16.975 22.86 17.145 ;
        RECT 22.43 16.95 22.66 17 ;
        RECT 22.43 16.905 22.61 17 ;
        RECT 22.57 16.975 22.86 17.125 ;
        RECT 22.36 16.85 22.57 16.93 ;
        RECT 22.31 16.78 22.5 16.87 ;
        RECT 20.1 16.75 22.43 16.845 ;
        RECT 20.17 16.71 22.43 16.845 ;
        RECT 20.17 16.695 22.36 16.845 ;
        RECT 20.21 16.675 22.36 16.845 ;
        RECT 20.03 16.82 20.26 16.87 ;
        RECT 20.03 16.82 20.21 16.915 ;
        RECT 19.96 16.89 20.17 16.97 ;
        RECT 19.91 16.95 20.1 17.04 ;
        RECT 19.67 16.975 20.03 17.11 ;
        RECT 19.71 16.975 19.96 17.145 ;
        RECT 19.53 16.95 19.76 17 ;
        RECT 19.53 16.905 19.71 17 ;
        RECT 19.67 16.975 19.96 17.125 ;
        RECT 19.46 16.85 19.67 16.93 ;
        RECT 19.6 16.975 20.03 17.07 ;
        RECT 19.41 16.78 19.6 16.87 ;
        RECT 17.125 16.71 19.53 16.845 ;
        RECT 17.125 16.675 19.46 16.845 ;
        RECT 17.14 16.675 17.36 16.85 ;
        RECT 17.14 16.675 17.35 16.89 ;
        RECT 16.7 16.975 17.14 17.07 ;
        RECT 17.01 16.95 17.21 17.03 ;
        RECT 17.13 16.85 17.14 17.07 ;
        RECT 16.77 16.975 17.13 17.11 ;
        RECT 17.06 16.89 17.28 16.96 ;
        RECT 16.81 16.975 17.06 17.145 ;
        RECT 16.63 16.95 16.86 17 ;
        RECT 16.63 16.905 16.81 17 ;
        RECT 16.77 16.975 17.06 17.125 ;
        RECT 16.56 16.85 16.77 16.93 ;
        RECT 16.51 16.78 16.7 16.87 ;
        RECT 14.3 16.75 16.63 16.845 ;
        RECT 14.37 16.71 16.63 16.845 ;
        RECT 14.37 16.695 16.56 16.845 ;
        RECT 14.41 16.675 16.56 16.845 ;
        RECT 14.23 16.82 14.46 16.87 ;
        RECT 14.23 16.82 14.41 16.915 ;
        RECT 14.16 16.89 14.37 16.97 ;
        RECT 14.11 16.95 14.3 17.04 ;
        RECT 13.87 16.975 14.23 17.11 ;
        RECT 13.91 16.975 14.16 17.145 ;
        RECT 13.73 16.95 13.96 17 ;
        RECT 13.73 16.905 13.91 17 ;
        RECT 13.87 16.975 14.16 17.125 ;
        RECT 13.66 16.85 13.87 16.93 ;
        RECT 13.8 16.975 14.23 17.07 ;
        RECT 13.61 16.78 13.8 16.87 ;
        RECT 11.325 16.71 13.73 16.845 ;
        RECT 11.325 16.675 13.66 16.845 ;
        RECT 11.34 16.675 11.56 16.85 ;
        RECT 11.34 16.675 11.55 16.89 ;
        RECT 10.9 16.975 11.34 17.07 ;
        RECT 11.21 16.95 11.41 17.03 ;
        RECT 11.33 16.85 11.34 17.07 ;
        RECT 10.97 16.975 11.33 17.11 ;
        RECT 11.26 16.89 11.48 16.96 ;
        RECT 11.01 16.975 11.26 17.145 ;
        RECT 10.83 16.95 11.06 17 ;
        RECT 10.83 16.905 11.01 17 ;
        RECT 10.97 16.975 11.26 17.125 ;
        RECT 10.76 16.85 10.97 16.93 ;
        RECT 10.71 16.78 10.9 16.87 ;
        RECT 8.5 16.75 10.83 16.845 ;
        RECT 8.57 16.71 10.83 16.845 ;
        RECT 8.57 16.695 10.76 16.845 ;
        RECT 8.61 16.675 10.76 16.845 ;
        RECT 8.43 16.82 8.66 16.87 ;
        RECT 8.43 16.82 8.61 16.915 ;
        RECT 8.36 16.89 8.57 16.97 ;
        RECT 8.31 16.95 8.5 17.04 ;
        RECT 8.07 16.975 8.43 17.11 ;
        RECT 8.11 16.975 8.36 17.145 ;
        RECT 7.93 16.95 8.16 17 ;
        RECT 7.93 16.905 8.11 17 ;
        RECT 8.07 16.975 8.36 17.125 ;
        RECT 7.86 16.85 8.07 16.93 ;
        RECT 8 16.975 8.43 17.07 ;
        RECT 7.81 16.78 8 16.87 ;
        RECT 5.525 16.71 7.93 16.845 ;
        RECT 5.525 16.675 7.86 16.845 ;
        RECT 5.54 16.675 5.76 16.85 ;
        RECT 5.54 16.675 5.75 16.89 ;
        RECT 5.1 16.975 5.54 17.07 ;
        RECT 5.41 16.95 5.61 17.03 ;
        RECT 5.53 16.85 5.54 17.07 ;
        RECT 5.17 16.975 5.53 17.11 ;
        RECT 5.46 16.89 5.68 16.96 ;
        RECT 5.21 16.975 5.46 17.145 ;
        RECT 5.03 16.95 5.26 17 ;
        RECT 5.03 16.905 5.21 17 ;
        RECT 5.17 16.975 5.46 17.125 ;
        RECT 4.96 16.85 5.17 16.93 ;
        RECT 4.91 16.78 5.1 16.87 ;
        RECT 2.7 16.75 5.03 16.845 ;
        RECT 2.77 16.71 5.03 16.845 ;
        RECT 2.77 16.695 4.96 16.845 ;
        RECT 2.81 16.675 4.96 16.845 ;
        RECT 2.63 16.82 2.86 16.87 ;
        RECT 2.63 16.82 2.81 16.915 ;
        RECT 2.56 16.89 2.77 16.97 ;
        RECT 2.51 16.95 2.7 17.04 ;
        RECT 2.27 16.975 2.63 17.11 ;
        RECT 2.31 16.975 2.56 17.145 ;
        RECT 2.13 16.95 2.36 17 ;
        RECT 2.13 16.905 2.31 17 ;
        RECT 2.27 16.975 2.56 17.125 ;
        RECT 2.06 16.85 2.27 16.93 ;
        RECT 2.2 16.975 2.63 17.07 ;
        RECT 2.01 16.78 2.2 16.87 ;
        RECT -0.455 16.71 2.13 16.845 ;
        RECT -0.455 16.675 2.06 16.845 ;
    END
  END RWL1_12
  PIN RWL1_13
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 18.025 34.76 18.22 ;
        RECT 34.53 18.17 34.71 18.265 ;
        RECT 34.6 18.1 34.76 18.22 ;
        RECT 34.67 18.045 34.71 18.265 ;
        RECT 34.46 18.24 34.67 18.32 ;
        RECT 34.41 18.3 34.6 18.39 ;
        RECT 34.17 18.325 34.53 18.46 ;
        RECT 34.21 18.325 34.46 18.495 ;
        RECT 34.03 18.3 34.26 18.35 ;
        RECT 34.03 18.255 34.21 18.35 ;
        RECT 34.17 18.325 34.46 18.475 ;
        RECT 33.96 18.2 34.17 18.28 ;
        RECT 34.1 18.325 34.53 18.42 ;
        RECT 33.91 18.13 34.1 18.22 ;
        RECT 31.7 18.1 34.03 18.195 ;
        RECT 31.77 18.06 34.03 18.195 ;
        RECT 31.77 18.045 33.96 18.195 ;
        RECT 31.81 18.025 33.96 18.195 ;
        RECT 31.63 18.17 31.86 18.22 ;
        RECT 31.63 18.17 31.81 18.265 ;
        RECT 31.56 18.24 31.77 18.32 ;
        RECT 31.51 18.3 31.7 18.39 ;
        RECT 31.27 18.325 31.63 18.46 ;
        RECT 31.31 18.325 31.56 18.495 ;
        RECT 31.13 18.3 31.36 18.35 ;
        RECT 31.13 18.255 31.31 18.35 ;
        RECT 31.27 18.325 31.56 18.475 ;
        RECT 31.06 18.2 31.27 18.28 ;
        RECT 31.2 18.325 31.63 18.42 ;
        RECT 31.01 18.13 31.2 18.22 ;
        RECT 28.725 18.06 31.13 18.195 ;
        RECT 28.725 18.025 31.06 18.195 ;
        RECT 28.74 18.025 28.96 18.2 ;
        RECT 28.74 18.025 28.95 18.24 ;
        RECT 28.3 18.325 28.74 18.42 ;
        RECT 28.61 18.3 28.81 18.38 ;
        RECT 28.73 18.2 28.74 18.42 ;
        RECT 28.37 18.325 28.73 18.46 ;
        RECT 28.66 18.24 28.88 18.31 ;
        RECT 28.41 18.325 28.66 18.495 ;
        RECT 28.23 18.3 28.46 18.35 ;
        RECT 28.23 18.255 28.41 18.35 ;
        RECT 28.37 18.325 28.66 18.475 ;
        RECT 28.16 18.2 28.37 18.28 ;
        RECT 28.11 18.13 28.3 18.22 ;
        RECT 25.9 18.1 28.23 18.195 ;
        RECT 25.97 18.06 28.23 18.195 ;
        RECT 25.97 18.045 28.16 18.195 ;
        RECT 26.01 18.025 28.16 18.195 ;
        RECT 25.83 18.17 26.06 18.22 ;
        RECT 25.83 18.17 26.01 18.265 ;
        RECT 25.76 18.24 25.97 18.32 ;
        RECT 25.71 18.3 25.9 18.39 ;
        RECT 25.47 18.325 25.83 18.46 ;
        RECT 25.51 18.325 25.76 18.495 ;
        RECT 25.33 18.3 25.56 18.35 ;
        RECT 25.33 18.255 25.51 18.35 ;
        RECT 25.47 18.325 25.76 18.475 ;
        RECT 25.26 18.2 25.47 18.28 ;
        RECT 25.4 18.325 25.83 18.42 ;
        RECT 25.21 18.13 25.4 18.22 ;
        RECT 22.925 18.06 25.33 18.195 ;
        RECT 22.925 18.025 25.26 18.195 ;
        RECT 22.94 18.025 23.16 18.2 ;
        RECT 22.94 18.025 23.15 18.24 ;
        RECT 22.5 18.325 22.94 18.42 ;
        RECT 22.81 18.3 23.01 18.38 ;
        RECT 22.93 18.2 22.94 18.42 ;
        RECT 22.57 18.325 22.93 18.46 ;
        RECT 22.86 18.24 23.08 18.31 ;
        RECT 22.61 18.325 22.86 18.495 ;
        RECT 22.43 18.3 22.66 18.35 ;
        RECT 22.43 18.255 22.61 18.35 ;
        RECT 22.57 18.325 22.86 18.475 ;
        RECT 22.36 18.2 22.57 18.28 ;
        RECT 22.31 18.13 22.5 18.22 ;
        RECT 20.1 18.1 22.43 18.195 ;
        RECT 20.17 18.06 22.43 18.195 ;
        RECT 20.17 18.045 22.36 18.195 ;
        RECT 20.21 18.025 22.36 18.195 ;
        RECT 20.03 18.17 20.26 18.22 ;
        RECT 20.03 18.17 20.21 18.265 ;
        RECT 19.96 18.24 20.17 18.32 ;
        RECT 19.91 18.3 20.1 18.39 ;
        RECT 19.67 18.325 20.03 18.46 ;
        RECT 19.71 18.325 19.96 18.495 ;
        RECT 19.53 18.3 19.76 18.35 ;
        RECT 19.53 18.255 19.71 18.35 ;
        RECT 19.67 18.325 19.96 18.475 ;
        RECT 19.46 18.2 19.67 18.28 ;
        RECT 19.6 18.325 20.03 18.42 ;
        RECT 19.41 18.13 19.6 18.22 ;
        RECT 17.125 18.06 19.53 18.195 ;
        RECT 17.125 18.025 19.46 18.195 ;
        RECT 17.14 18.025 17.36 18.2 ;
        RECT 17.14 18.025 17.35 18.24 ;
        RECT 16.7 18.325 17.14 18.42 ;
        RECT 17.01 18.3 17.21 18.38 ;
        RECT 17.13 18.2 17.14 18.42 ;
        RECT 16.77 18.325 17.13 18.46 ;
        RECT 17.06 18.24 17.28 18.31 ;
        RECT 16.81 18.325 17.06 18.495 ;
        RECT 16.63 18.3 16.86 18.35 ;
        RECT 16.63 18.255 16.81 18.35 ;
        RECT 16.77 18.325 17.06 18.475 ;
        RECT 16.56 18.2 16.77 18.28 ;
        RECT 16.51 18.13 16.7 18.22 ;
        RECT 14.3 18.1 16.63 18.195 ;
        RECT 14.37 18.06 16.63 18.195 ;
        RECT 14.37 18.045 16.56 18.195 ;
        RECT 14.41 18.025 16.56 18.195 ;
        RECT 14.23 18.17 14.46 18.22 ;
        RECT 14.23 18.17 14.41 18.265 ;
        RECT 14.16 18.24 14.37 18.32 ;
        RECT 14.11 18.3 14.3 18.39 ;
        RECT 13.87 18.325 14.23 18.46 ;
        RECT 13.91 18.325 14.16 18.495 ;
        RECT 13.73 18.3 13.96 18.35 ;
        RECT 13.73 18.255 13.91 18.35 ;
        RECT 13.87 18.325 14.16 18.475 ;
        RECT 13.66 18.2 13.87 18.28 ;
        RECT 13.8 18.325 14.23 18.42 ;
        RECT 13.61 18.13 13.8 18.22 ;
        RECT 11.325 18.06 13.73 18.195 ;
        RECT 11.325 18.025 13.66 18.195 ;
        RECT 11.34 18.025 11.56 18.2 ;
        RECT 11.34 18.025 11.55 18.24 ;
        RECT 10.9 18.325 11.34 18.42 ;
        RECT 11.21 18.3 11.41 18.38 ;
        RECT 11.33 18.2 11.34 18.42 ;
        RECT 10.97 18.325 11.33 18.46 ;
        RECT 11.26 18.24 11.48 18.31 ;
        RECT 11.01 18.325 11.26 18.495 ;
        RECT 10.83 18.3 11.06 18.35 ;
        RECT 10.83 18.255 11.01 18.35 ;
        RECT 10.97 18.325 11.26 18.475 ;
        RECT 10.76 18.2 10.97 18.28 ;
        RECT 10.71 18.13 10.9 18.22 ;
        RECT 8.5 18.1 10.83 18.195 ;
        RECT 8.57 18.06 10.83 18.195 ;
        RECT 8.57 18.045 10.76 18.195 ;
        RECT 8.61 18.025 10.76 18.195 ;
        RECT 8.43 18.17 8.66 18.22 ;
        RECT 8.43 18.17 8.61 18.265 ;
        RECT 8.36 18.24 8.57 18.32 ;
        RECT 8.31 18.3 8.5 18.39 ;
        RECT 8.07 18.325 8.43 18.46 ;
        RECT 8.11 18.325 8.36 18.495 ;
        RECT 7.93 18.3 8.16 18.35 ;
        RECT 7.93 18.255 8.11 18.35 ;
        RECT 8.07 18.325 8.36 18.475 ;
        RECT 7.86 18.2 8.07 18.28 ;
        RECT 8 18.325 8.43 18.42 ;
        RECT 7.81 18.13 8 18.22 ;
        RECT 5.525 18.06 7.93 18.195 ;
        RECT 5.525 18.025 7.86 18.195 ;
        RECT 5.54 18.025 5.76 18.2 ;
        RECT 5.54 18.025 5.75 18.24 ;
        RECT 5.1 18.325 5.54 18.42 ;
        RECT 5.41 18.3 5.61 18.38 ;
        RECT 5.53 18.2 5.54 18.42 ;
        RECT 5.17 18.325 5.53 18.46 ;
        RECT 5.46 18.24 5.68 18.31 ;
        RECT 5.21 18.325 5.46 18.495 ;
        RECT 5.03 18.3 5.26 18.35 ;
        RECT 5.03 18.255 5.21 18.35 ;
        RECT 5.17 18.325 5.46 18.475 ;
        RECT 4.96 18.2 5.17 18.28 ;
        RECT 4.91 18.13 5.1 18.22 ;
        RECT 2.7 18.1 5.03 18.195 ;
        RECT 2.77 18.06 5.03 18.195 ;
        RECT 2.77 18.045 4.96 18.195 ;
        RECT 2.81 18.025 4.96 18.195 ;
        RECT 2.63 18.17 2.86 18.22 ;
        RECT 2.63 18.17 2.81 18.265 ;
        RECT 2.56 18.24 2.77 18.32 ;
        RECT 2.51 18.3 2.7 18.39 ;
        RECT 2.27 18.325 2.63 18.46 ;
        RECT 2.31 18.325 2.56 18.495 ;
        RECT 2.13 18.3 2.36 18.35 ;
        RECT 2.13 18.255 2.31 18.35 ;
        RECT 2.27 18.325 2.56 18.475 ;
        RECT 2.06 18.2 2.27 18.28 ;
        RECT 2.2 18.325 2.63 18.42 ;
        RECT 2.01 18.13 2.2 18.22 ;
        RECT -0.455 18.06 2.13 18.195 ;
        RECT -0.455 18.025 2.06 18.195 ;
    END
  END RWL1_13
  PIN RWL1_14
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 19.375 34.76 19.57 ;
        RECT 34.53 19.52 34.71 19.615 ;
        RECT 34.6 19.45 34.76 19.57 ;
        RECT 34.67 19.395 34.71 19.615 ;
        RECT 34.46 19.59 34.67 19.67 ;
        RECT 34.41 19.65 34.6 19.74 ;
        RECT 34.17 19.675 34.53 19.81 ;
        RECT 34.21 19.675 34.46 19.845 ;
        RECT 34.03 19.65 34.26 19.7 ;
        RECT 34.03 19.605 34.21 19.7 ;
        RECT 34.17 19.675 34.46 19.825 ;
        RECT 33.96 19.55 34.17 19.63 ;
        RECT 34.1 19.675 34.53 19.77 ;
        RECT 33.91 19.48 34.1 19.57 ;
        RECT 31.7 19.45 34.03 19.545 ;
        RECT 31.77 19.41 34.03 19.545 ;
        RECT 31.77 19.395 33.96 19.545 ;
        RECT 31.81 19.375 33.96 19.545 ;
        RECT 31.63 19.52 31.86 19.57 ;
        RECT 31.63 19.52 31.81 19.615 ;
        RECT 31.56 19.59 31.77 19.67 ;
        RECT 31.51 19.65 31.7 19.74 ;
        RECT 31.27 19.675 31.63 19.81 ;
        RECT 31.31 19.675 31.56 19.845 ;
        RECT 31.13 19.65 31.36 19.7 ;
        RECT 31.13 19.605 31.31 19.7 ;
        RECT 31.27 19.675 31.56 19.825 ;
        RECT 31.06 19.55 31.27 19.63 ;
        RECT 31.2 19.675 31.63 19.77 ;
        RECT 31.01 19.48 31.2 19.57 ;
        RECT 28.725 19.41 31.13 19.545 ;
        RECT 28.725 19.375 31.06 19.545 ;
        RECT 28.74 19.375 28.96 19.55 ;
        RECT 28.74 19.375 28.95 19.59 ;
        RECT 28.3 19.675 28.74 19.77 ;
        RECT 28.61 19.65 28.81 19.73 ;
        RECT 28.73 19.55 28.74 19.77 ;
        RECT 28.37 19.675 28.73 19.81 ;
        RECT 28.66 19.59 28.88 19.66 ;
        RECT 28.41 19.675 28.66 19.845 ;
        RECT 28.23 19.65 28.46 19.7 ;
        RECT 28.23 19.605 28.41 19.7 ;
        RECT 28.37 19.675 28.66 19.825 ;
        RECT 28.16 19.55 28.37 19.63 ;
        RECT 28.11 19.48 28.3 19.57 ;
        RECT 25.9 19.45 28.23 19.545 ;
        RECT 25.97 19.41 28.23 19.545 ;
        RECT 25.97 19.395 28.16 19.545 ;
        RECT 26.01 19.375 28.16 19.545 ;
        RECT 25.83 19.52 26.06 19.57 ;
        RECT 25.83 19.52 26.01 19.615 ;
        RECT 25.76 19.59 25.97 19.67 ;
        RECT 25.71 19.65 25.9 19.74 ;
        RECT 25.47 19.675 25.83 19.81 ;
        RECT 25.51 19.675 25.76 19.845 ;
        RECT 25.33 19.65 25.56 19.7 ;
        RECT 25.33 19.605 25.51 19.7 ;
        RECT 25.47 19.675 25.76 19.825 ;
        RECT 25.26 19.55 25.47 19.63 ;
        RECT 25.4 19.675 25.83 19.77 ;
        RECT 25.21 19.48 25.4 19.57 ;
        RECT 22.925 19.41 25.33 19.545 ;
        RECT 22.925 19.375 25.26 19.545 ;
        RECT 22.94 19.375 23.16 19.55 ;
        RECT 22.94 19.375 23.15 19.59 ;
        RECT 22.5 19.675 22.94 19.77 ;
        RECT 22.81 19.65 23.01 19.73 ;
        RECT 22.93 19.55 22.94 19.77 ;
        RECT 22.57 19.675 22.93 19.81 ;
        RECT 22.86 19.59 23.08 19.66 ;
        RECT 22.61 19.675 22.86 19.845 ;
        RECT 22.43 19.65 22.66 19.7 ;
        RECT 22.43 19.605 22.61 19.7 ;
        RECT 22.57 19.675 22.86 19.825 ;
        RECT 22.36 19.55 22.57 19.63 ;
        RECT 22.31 19.48 22.5 19.57 ;
        RECT 20.1 19.45 22.43 19.545 ;
        RECT 20.17 19.41 22.43 19.545 ;
        RECT 20.17 19.395 22.36 19.545 ;
        RECT 20.21 19.375 22.36 19.545 ;
        RECT 20.03 19.52 20.26 19.57 ;
        RECT 20.03 19.52 20.21 19.615 ;
        RECT 19.96 19.59 20.17 19.67 ;
        RECT 19.91 19.65 20.1 19.74 ;
        RECT 19.67 19.675 20.03 19.81 ;
        RECT 19.71 19.675 19.96 19.845 ;
        RECT 19.53 19.65 19.76 19.7 ;
        RECT 19.53 19.605 19.71 19.7 ;
        RECT 19.67 19.675 19.96 19.825 ;
        RECT 19.46 19.55 19.67 19.63 ;
        RECT 19.6 19.675 20.03 19.77 ;
        RECT 19.41 19.48 19.6 19.57 ;
        RECT 17.125 19.41 19.53 19.545 ;
        RECT 17.125 19.375 19.46 19.545 ;
        RECT 17.14 19.375 17.36 19.55 ;
        RECT 17.14 19.375 17.35 19.59 ;
        RECT 16.7 19.675 17.14 19.77 ;
        RECT 17.01 19.65 17.21 19.73 ;
        RECT 17.13 19.55 17.14 19.77 ;
        RECT 16.77 19.675 17.13 19.81 ;
        RECT 17.06 19.59 17.28 19.66 ;
        RECT 16.81 19.675 17.06 19.845 ;
        RECT 16.63 19.65 16.86 19.7 ;
        RECT 16.63 19.605 16.81 19.7 ;
        RECT 16.77 19.675 17.06 19.825 ;
        RECT 16.56 19.55 16.77 19.63 ;
        RECT 16.51 19.48 16.7 19.57 ;
        RECT 14.3 19.45 16.63 19.545 ;
        RECT 14.37 19.41 16.63 19.545 ;
        RECT 14.37 19.395 16.56 19.545 ;
        RECT 14.41 19.375 16.56 19.545 ;
        RECT 14.23 19.52 14.46 19.57 ;
        RECT 14.23 19.52 14.41 19.615 ;
        RECT 14.16 19.59 14.37 19.67 ;
        RECT 14.11 19.65 14.3 19.74 ;
        RECT 13.87 19.675 14.23 19.81 ;
        RECT 13.91 19.675 14.16 19.845 ;
        RECT 13.73 19.65 13.96 19.7 ;
        RECT 13.73 19.605 13.91 19.7 ;
        RECT 13.87 19.675 14.16 19.825 ;
        RECT 13.66 19.55 13.87 19.63 ;
        RECT 13.8 19.675 14.23 19.77 ;
        RECT 13.61 19.48 13.8 19.57 ;
        RECT 11.325 19.41 13.73 19.545 ;
        RECT 11.325 19.375 13.66 19.545 ;
        RECT 11.34 19.375 11.56 19.55 ;
        RECT 11.34 19.375 11.55 19.59 ;
        RECT 10.9 19.675 11.34 19.77 ;
        RECT 11.21 19.65 11.41 19.73 ;
        RECT 11.33 19.55 11.34 19.77 ;
        RECT 10.97 19.675 11.33 19.81 ;
        RECT 11.26 19.59 11.48 19.66 ;
        RECT 11.01 19.675 11.26 19.845 ;
        RECT 10.83 19.65 11.06 19.7 ;
        RECT 10.83 19.605 11.01 19.7 ;
        RECT 10.97 19.675 11.26 19.825 ;
        RECT 10.76 19.55 10.97 19.63 ;
        RECT 10.71 19.48 10.9 19.57 ;
        RECT 8.5 19.45 10.83 19.545 ;
        RECT 8.57 19.41 10.83 19.545 ;
        RECT 8.57 19.395 10.76 19.545 ;
        RECT 8.61 19.375 10.76 19.545 ;
        RECT 8.43 19.52 8.66 19.57 ;
        RECT 8.43 19.52 8.61 19.615 ;
        RECT 8.36 19.59 8.57 19.67 ;
        RECT 8.31 19.65 8.5 19.74 ;
        RECT 8.07 19.675 8.43 19.81 ;
        RECT 8.11 19.675 8.36 19.845 ;
        RECT 7.93 19.65 8.16 19.7 ;
        RECT 7.93 19.605 8.11 19.7 ;
        RECT 8.07 19.675 8.36 19.825 ;
        RECT 7.86 19.55 8.07 19.63 ;
        RECT 8 19.675 8.43 19.77 ;
        RECT 7.81 19.48 8 19.57 ;
        RECT 5.525 19.41 7.93 19.545 ;
        RECT 5.525 19.375 7.86 19.545 ;
        RECT 5.54 19.375 5.76 19.55 ;
        RECT 5.54 19.375 5.75 19.59 ;
        RECT 5.1 19.675 5.54 19.77 ;
        RECT 5.41 19.65 5.61 19.73 ;
        RECT 5.53 19.55 5.54 19.77 ;
        RECT 5.17 19.675 5.53 19.81 ;
        RECT 5.46 19.59 5.68 19.66 ;
        RECT 5.21 19.675 5.46 19.845 ;
        RECT 5.03 19.65 5.26 19.7 ;
        RECT 5.03 19.605 5.21 19.7 ;
        RECT 5.17 19.675 5.46 19.825 ;
        RECT 4.96 19.55 5.17 19.63 ;
        RECT 4.91 19.48 5.1 19.57 ;
        RECT 2.7 19.45 5.03 19.545 ;
        RECT 2.77 19.41 5.03 19.545 ;
        RECT 2.77 19.395 4.96 19.545 ;
        RECT 2.81 19.375 4.96 19.545 ;
        RECT 2.63 19.52 2.86 19.57 ;
        RECT 2.63 19.52 2.81 19.615 ;
        RECT 2.56 19.59 2.77 19.67 ;
        RECT 2.51 19.65 2.7 19.74 ;
        RECT 2.27 19.675 2.63 19.81 ;
        RECT 2.31 19.675 2.56 19.845 ;
        RECT 2.13 19.65 2.36 19.7 ;
        RECT 2.13 19.605 2.31 19.7 ;
        RECT 2.27 19.675 2.56 19.825 ;
        RECT 2.06 19.55 2.27 19.63 ;
        RECT 2.2 19.675 2.63 19.77 ;
        RECT 2.01 19.48 2.2 19.57 ;
        RECT -0.455 19.41 2.13 19.545 ;
        RECT -0.455 19.375 2.06 19.545 ;
    END
  END RWL1_14
  PIN RWL1_15
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 20.725 34.76 20.92 ;
        RECT 34.53 20.87 34.71 20.965 ;
        RECT 34.6 20.8 34.76 20.92 ;
        RECT 34.67 20.745 34.71 20.965 ;
        RECT 34.46 20.94 34.67 21.02 ;
        RECT 34.41 21 34.6 21.09 ;
        RECT 34.17 21.025 34.53 21.16 ;
        RECT 34.21 21.025 34.46 21.195 ;
        RECT 34.03 21 34.26 21.05 ;
        RECT 34.03 20.955 34.21 21.05 ;
        RECT 34.17 21.025 34.46 21.175 ;
        RECT 33.96 20.9 34.17 20.98 ;
        RECT 34.1 21.025 34.53 21.12 ;
        RECT 33.91 20.83 34.1 20.92 ;
        RECT 31.7 20.8 34.03 20.895 ;
        RECT 31.77 20.76 34.03 20.895 ;
        RECT 31.77 20.745 33.96 20.895 ;
        RECT 31.81 20.725 33.96 20.895 ;
        RECT 31.63 20.87 31.86 20.92 ;
        RECT 31.63 20.87 31.81 20.965 ;
        RECT 31.56 20.94 31.77 21.02 ;
        RECT 31.51 21 31.7 21.09 ;
        RECT 31.27 21.025 31.63 21.16 ;
        RECT 31.31 21.025 31.56 21.195 ;
        RECT 31.13 21 31.36 21.05 ;
        RECT 31.13 20.955 31.31 21.05 ;
        RECT 31.27 21.025 31.56 21.175 ;
        RECT 31.06 20.9 31.27 20.98 ;
        RECT 31.2 21.025 31.63 21.12 ;
        RECT 31.01 20.83 31.2 20.92 ;
        RECT 28.725 20.76 31.13 20.895 ;
        RECT 28.725 20.725 31.06 20.895 ;
        RECT 28.74 20.725 28.96 20.9 ;
        RECT 28.74 20.725 28.95 20.94 ;
        RECT 28.3 21.025 28.74 21.12 ;
        RECT 28.61 21 28.81 21.08 ;
        RECT 28.73 20.9 28.74 21.12 ;
        RECT 28.37 21.025 28.73 21.16 ;
        RECT 28.66 20.94 28.88 21.01 ;
        RECT 28.41 21.025 28.66 21.195 ;
        RECT 28.23 21 28.46 21.05 ;
        RECT 28.23 20.955 28.41 21.05 ;
        RECT 28.37 21.025 28.66 21.175 ;
        RECT 28.16 20.9 28.37 20.98 ;
        RECT 28.11 20.83 28.3 20.92 ;
        RECT 25.9 20.8 28.23 20.895 ;
        RECT 25.97 20.76 28.23 20.895 ;
        RECT 25.97 20.745 28.16 20.895 ;
        RECT 26.01 20.725 28.16 20.895 ;
        RECT 25.83 20.87 26.06 20.92 ;
        RECT 25.83 20.87 26.01 20.965 ;
        RECT 25.76 20.94 25.97 21.02 ;
        RECT 25.71 21 25.9 21.09 ;
        RECT 25.47 21.025 25.83 21.16 ;
        RECT 25.51 21.025 25.76 21.195 ;
        RECT 25.33 21 25.56 21.05 ;
        RECT 25.33 20.955 25.51 21.05 ;
        RECT 25.47 21.025 25.76 21.175 ;
        RECT 25.26 20.9 25.47 20.98 ;
        RECT 25.4 21.025 25.83 21.12 ;
        RECT 25.21 20.83 25.4 20.92 ;
        RECT 22.925 20.76 25.33 20.895 ;
        RECT 22.925 20.725 25.26 20.895 ;
        RECT 22.94 20.725 23.16 20.9 ;
        RECT 22.94 20.725 23.15 20.94 ;
        RECT 22.5 21.025 22.94 21.12 ;
        RECT 22.81 21 23.01 21.08 ;
        RECT 22.93 20.9 22.94 21.12 ;
        RECT 22.57 21.025 22.93 21.16 ;
        RECT 22.86 20.94 23.08 21.01 ;
        RECT 22.61 21.025 22.86 21.195 ;
        RECT 22.43 21 22.66 21.05 ;
        RECT 22.43 20.955 22.61 21.05 ;
        RECT 22.57 21.025 22.86 21.175 ;
        RECT 22.36 20.9 22.57 20.98 ;
        RECT 22.31 20.83 22.5 20.92 ;
        RECT 20.1 20.8 22.43 20.895 ;
        RECT 20.17 20.76 22.43 20.895 ;
        RECT 20.17 20.745 22.36 20.895 ;
        RECT 20.21 20.725 22.36 20.895 ;
        RECT 20.03 20.87 20.26 20.92 ;
        RECT 20.03 20.87 20.21 20.965 ;
        RECT 19.96 20.94 20.17 21.02 ;
        RECT 19.91 21 20.1 21.09 ;
        RECT 19.67 21.025 20.03 21.16 ;
        RECT 19.71 21.025 19.96 21.195 ;
        RECT 19.53 21 19.76 21.05 ;
        RECT 19.53 20.955 19.71 21.05 ;
        RECT 19.67 21.025 19.96 21.175 ;
        RECT 19.46 20.9 19.67 20.98 ;
        RECT 19.6 21.025 20.03 21.12 ;
        RECT 19.41 20.83 19.6 20.92 ;
        RECT 17.125 20.76 19.53 20.895 ;
        RECT 17.125 20.725 19.46 20.895 ;
        RECT 17.14 20.725 17.36 20.9 ;
        RECT 17.14 20.725 17.35 20.94 ;
        RECT 16.7 21.025 17.14 21.12 ;
        RECT 17.01 21 17.21 21.08 ;
        RECT 17.13 20.9 17.14 21.12 ;
        RECT 16.77 21.025 17.13 21.16 ;
        RECT 17.06 20.94 17.28 21.01 ;
        RECT 16.81 21.025 17.06 21.195 ;
        RECT 16.63 21 16.86 21.05 ;
        RECT 16.63 20.955 16.81 21.05 ;
        RECT 16.77 21.025 17.06 21.175 ;
        RECT 16.56 20.9 16.77 20.98 ;
        RECT 16.51 20.83 16.7 20.92 ;
        RECT 14.3 20.8 16.63 20.895 ;
        RECT 14.37 20.76 16.63 20.895 ;
        RECT 14.37 20.745 16.56 20.895 ;
        RECT 14.41 20.725 16.56 20.895 ;
        RECT 14.23 20.87 14.46 20.92 ;
        RECT 14.23 20.87 14.41 20.965 ;
        RECT 14.16 20.94 14.37 21.02 ;
        RECT 14.11 21 14.3 21.09 ;
        RECT 13.87 21.025 14.23 21.16 ;
        RECT 13.91 21.025 14.16 21.195 ;
        RECT 13.73 21 13.96 21.05 ;
        RECT 13.73 20.955 13.91 21.05 ;
        RECT 13.87 21.025 14.16 21.175 ;
        RECT 13.66 20.9 13.87 20.98 ;
        RECT 13.8 21.025 14.23 21.12 ;
        RECT 13.61 20.83 13.8 20.92 ;
        RECT 11.325 20.76 13.73 20.895 ;
        RECT 11.325 20.725 13.66 20.895 ;
        RECT 11.34 20.725 11.56 20.9 ;
        RECT 11.34 20.725 11.55 20.94 ;
        RECT 10.9 21.025 11.34 21.12 ;
        RECT 11.21 21 11.41 21.08 ;
        RECT 11.33 20.9 11.34 21.12 ;
        RECT 10.97 21.025 11.33 21.16 ;
        RECT 11.26 20.94 11.48 21.01 ;
        RECT 11.01 21.025 11.26 21.195 ;
        RECT 10.83 21 11.06 21.05 ;
        RECT 10.83 20.955 11.01 21.05 ;
        RECT 10.97 21.025 11.26 21.175 ;
        RECT 10.76 20.9 10.97 20.98 ;
        RECT 10.71 20.83 10.9 20.92 ;
        RECT 8.5 20.8 10.83 20.895 ;
        RECT 8.57 20.76 10.83 20.895 ;
        RECT 8.57 20.745 10.76 20.895 ;
        RECT 8.61 20.725 10.76 20.895 ;
        RECT 8.43 20.87 8.66 20.92 ;
        RECT 8.43 20.87 8.61 20.965 ;
        RECT 8.36 20.94 8.57 21.02 ;
        RECT 8.31 21 8.5 21.09 ;
        RECT 8.07 21.025 8.43 21.16 ;
        RECT 8.11 21.025 8.36 21.195 ;
        RECT 7.93 21 8.16 21.05 ;
        RECT 7.93 20.955 8.11 21.05 ;
        RECT 8.07 21.025 8.36 21.175 ;
        RECT 7.86 20.9 8.07 20.98 ;
        RECT 8 21.025 8.43 21.12 ;
        RECT 7.81 20.83 8 20.92 ;
        RECT 5.525 20.76 7.93 20.895 ;
        RECT 5.525 20.725 7.86 20.895 ;
        RECT 5.54 20.725 5.76 20.9 ;
        RECT 5.54 20.725 5.75 20.94 ;
        RECT 5.1 21.025 5.54 21.12 ;
        RECT 5.41 21 5.61 21.08 ;
        RECT 5.53 20.9 5.54 21.12 ;
        RECT 5.17 21.025 5.53 21.16 ;
        RECT 5.46 20.94 5.68 21.01 ;
        RECT 5.21 21.025 5.46 21.195 ;
        RECT 5.03 21 5.26 21.05 ;
        RECT 5.03 20.955 5.21 21.05 ;
        RECT 5.17 21.025 5.46 21.175 ;
        RECT 4.96 20.9 5.17 20.98 ;
        RECT 4.91 20.83 5.1 20.92 ;
        RECT 2.7 20.8 5.03 20.895 ;
        RECT 2.77 20.76 5.03 20.895 ;
        RECT 2.77 20.745 4.96 20.895 ;
        RECT 2.81 20.725 4.96 20.895 ;
        RECT 2.63 20.87 2.86 20.92 ;
        RECT 2.63 20.87 2.81 20.965 ;
        RECT 2.56 20.94 2.77 21.02 ;
        RECT 2.51 21 2.7 21.09 ;
        RECT 2.27 21.025 2.63 21.16 ;
        RECT 2.31 21.025 2.56 21.195 ;
        RECT 2.13 21 2.36 21.05 ;
        RECT 2.13 20.955 2.31 21.05 ;
        RECT 2.27 21.025 2.56 21.175 ;
        RECT 2.06 20.9 2.27 20.98 ;
        RECT 2.2 21.025 2.63 21.12 ;
        RECT 2.01 20.83 2.2 20.92 ;
        RECT -0.455 20.76 2.13 20.895 ;
        RECT -0.455 20.725 2.06 20.895 ;
    END
  END RWL1_15
  PIN RWL1_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 3.175 34.76 3.37 ;
        RECT 34.53 3.32 34.71 3.415 ;
        RECT 34.6 3.25 34.76 3.37 ;
        RECT 34.67 3.195 34.71 3.415 ;
        RECT 34.46 3.39 34.67 3.47 ;
        RECT 34.41 3.45 34.6 3.54 ;
        RECT 34.17 3.475 34.53 3.61 ;
        RECT 34.21 3.475 34.46 3.645 ;
        RECT 34.03 3.45 34.26 3.5 ;
        RECT 34.03 3.405 34.21 3.5 ;
        RECT 34.17 3.475 34.46 3.625 ;
        RECT 33.96 3.35 34.17 3.43 ;
        RECT 34.1 3.475 34.53 3.57 ;
        RECT 33.91 3.28 34.1 3.37 ;
        RECT 31.7 3.25 34.03 3.345 ;
        RECT 31.77 3.21 34.03 3.345 ;
        RECT 31.77 3.195 33.96 3.345 ;
        RECT 31.81 3.175 33.96 3.345 ;
        RECT 31.63 3.32 31.86 3.37 ;
        RECT 31.63 3.32 31.81 3.415 ;
        RECT 31.56 3.39 31.77 3.47 ;
        RECT 31.51 3.45 31.7 3.54 ;
        RECT 31.27 3.475 31.63 3.61 ;
        RECT 31.31 3.475 31.56 3.645 ;
        RECT 31.13 3.45 31.36 3.5 ;
        RECT 31.13 3.405 31.31 3.5 ;
        RECT 31.27 3.475 31.56 3.625 ;
        RECT 31.06 3.35 31.27 3.43 ;
        RECT 31.2 3.475 31.63 3.57 ;
        RECT 31.01 3.28 31.2 3.37 ;
        RECT 28.725 3.21 31.13 3.345 ;
        RECT 28.725 3.175 31.06 3.345 ;
        RECT 28.74 3.175 28.96 3.35 ;
        RECT 28.74 3.175 28.95 3.39 ;
        RECT 28.3 3.475 28.74 3.57 ;
        RECT 28.61 3.45 28.81 3.53 ;
        RECT 28.73 3.35 28.74 3.57 ;
        RECT 28.37 3.475 28.73 3.61 ;
        RECT 28.66 3.39 28.88 3.46 ;
        RECT 28.41 3.475 28.66 3.645 ;
        RECT 28.23 3.45 28.46 3.5 ;
        RECT 28.23 3.405 28.41 3.5 ;
        RECT 28.37 3.475 28.66 3.625 ;
        RECT 28.16 3.35 28.37 3.43 ;
        RECT 28.11 3.28 28.3 3.37 ;
        RECT 25.9 3.25 28.23 3.345 ;
        RECT 25.97 3.21 28.23 3.345 ;
        RECT 25.97 3.195 28.16 3.345 ;
        RECT 26.01 3.175 28.16 3.345 ;
        RECT 25.83 3.32 26.06 3.37 ;
        RECT 25.83 3.32 26.01 3.415 ;
        RECT 25.76 3.39 25.97 3.47 ;
        RECT 25.71 3.45 25.9 3.54 ;
        RECT 25.47 3.475 25.83 3.61 ;
        RECT 25.51 3.475 25.76 3.645 ;
        RECT 25.33 3.45 25.56 3.5 ;
        RECT 25.33 3.405 25.51 3.5 ;
        RECT 25.47 3.475 25.76 3.625 ;
        RECT 25.26 3.35 25.47 3.43 ;
        RECT 25.4 3.475 25.83 3.57 ;
        RECT 25.21 3.28 25.4 3.37 ;
        RECT 22.925 3.21 25.33 3.345 ;
        RECT 22.925 3.175 25.26 3.345 ;
        RECT 22.94 3.175 23.16 3.35 ;
        RECT 22.94 3.175 23.15 3.39 ;
        RECT 22.5 3.475 22.94 3.57 ;
        RECT 22.81 3.45 23.01 3.53 ;
        RECT 22.93 3.35 22.94 3.57 ;
        RECT 22.57 3.475 22.93 3.61 ;
        RECT 22.86 3.39 23.08 3.46 ;
        RECT 22.61 3.475 22.86 3.645 ;
        RECT 22.43 3.45 22.66 3.5 ;
        RECT 22.43 3.405 22.61 3.5 ;
        RECT 22.57 3.475 22.86 3.625 ;
        RECT 22.36 3.35 22.57 3.43 ;
        RECT 22.31 3.28 22.5 3.37 ;
        RECT 20.1 3.25 22.43 3.345 ;
        RECT 20.17 3.21 22.43 3.345 ;
        RECT 20.17 3.195 22.36 3.345 ;
        RECT 20.21 3.175 22.36 3.345 ;
        RECT 20.03 3.32 20.26 3.37 ;
        RECT 20.03 3.32 20.21 3.415 ;
        RECT 19.96 3.39 20.17 3.47 ;
        RECT 19.91 3.45 20.1 3.54 ;
        RECT 19.67 3.475 20.03 3.61 ;
        RECT 19.71 3.475 19.96 3.645 ;
        RECT 19.53 3.45 19.76 3.5 ;
        RECT 19.53 3.405 19.71 3.5 ;
        RECT 19.67 3.475 19.96 3.625 ;
        RECT 19.46 3.35 19.67 3.43 ;
        RECT 19.6 3.475 20.03 3.57 ;
        RECT 19.41 3.28 19.6 3.37 ;
        RECT 17.125 3.21 19.53 3.345 ;
        RECT 17.125 3.175 19.46 3.345 ;
        RECT 17.14 3.175 17.36 3.35 ;
        RECT 17.14 3.175 17.35 3.39 ;
        RECT 16.7 3.475 17.14 3.57 ;
        RECT 17.01 3.45 17.21 3.53 ;
        RECT 17.13 3.35 17.14 3.57 ;
        RECT 16.77 3.475 17.13 3.61 ;
        RECT 17.06 3.39 17.28 3.46 ;
        RECT 16.81 3.475 17.06 3.645 ;
        RECT 16.63 3.45 16.86 3.5 ;
        RECT 16.63 3.405 16.81 3.5 ;
        RECT 16.77 3.475 17.06 3.625 ;
        RECT 16.56 3.35 16.77 3.43 ;
        RECT 16.51 3.28 16.7 3.37 ;
        RECT 14.3 3.25 16.63 3.345 ;
        RECT 14.37 3.21 16.63 3.345 ;
        RECT 14.37 3.195 16.56 3.345 ;
        RECT 14.41 3.175 16.56 3.345 ;
        RECT 14.23 3.32 14.46 3.37 ;
        RECT 14.23 3.32 14.41 3.415 ;
        RECT 14.16 3.39 14.37 3.47 ;
        RECT 14.11 3.45 14.3 3.54 ;
        RECT 13.87 3.475 14.23 3.61 ;
        RECT 13.91 3.475 14.16 3.645 ;
        RECT 13.73 3.45 13.96 3.5 ;
        RECT 13.73 3.405 13.91 3.5 ;
        RECT 13.87 3.475 14.16 3.625 ;
        RECT 13.66 3.35 13.87 3.43 ;
        RECT 13.8 3.475 14.23 3.57 ;
        RECT 13.61 3.28 13.8 3.37 ;
        RECT 11.325 3.21 13.73 3.345 ;
        RECT 11.325 3.175 13.66 3.345 ;
        RECT 11.34 3.175 11.56 3.35 ;
        RECT 11.34 3.175 11.55 3.39 ;
        RECT 10.9 3.475 11.34 3.57 ;
        RECT 11.21 3.45 11.41 3.53 ;
        RECT 11.33 3.35 11.34 3.57 ;
        RECT 10.97 3.475 11.33 3.61 ;
        RECT 11.26 3.39 11.48 3.46 ;
        RECT 11.01 3.475 11.26 3.645 ;
        RECT 10.83 3.45 11.06 3.5 ;
        RECT 10.83 3.405 11.01 3.5 ;
        RECT 10.97 3.475 11.26 3.625 ;
        RECT 10.76 3.35 10.97 3.43 ;
        RECT 10.71 3.28 10.9 3.37 ;
        RECT 8.5 3.25 10.83 3.345 ;
        RECT 8.57 3.21 10.83 3.345 ;
        RECT 8.57 3.195 10.76 3.345 ;
        RECT 8.61 3.175 10.76 3.345 ;
        RECT 8.43 3.32 8.66 3.37 ;
        RECT 8.43 3.32 8.61 3.415 ;
        RECT 8.36 3.39 8.57 3.47 ;
        RECT 8.31 3.45 8.5 3.54 ;
        RECT 8.07 3.475 8.43 3.61 ;
        RECT 8.11 3.475 8.36 3.645 ;
        RECT 7.93 3.45 8.16 3.5 ;
        RECT 7.93 3.405 8.11 3.5 ;
        RECT 8.07 3.475 8.36 3.625 ;
        RECT 7.86 3.35 8.07 3.43 ;
        RECT 8 3.475 8.43 3.57 ;
        RECT 7.81 3.28 8 3.37 ;
        RECT 5.525 3.21 7.93 3.345 ;
        RECT 5.525 3.175 7.86 3.345 ;
        RECT 5.54 3.175 5.76 3.35 ;
        RECT 5.54 3.175 5.75 3.39 ;
        RECT 5.1 3.475 5.54 3.57 ;
        RECT 5.41 3.45 5.61 3.53 ;
        RECT 5.53 3.35 5.54 3.57 ;
        RECT 5.17 3.475 5.53 3.61 ;
        RECT 5.46 3.39 5.68 3.46 ;
        RECT 5.21 3.475 5.46 3.645 ;
        RECT 5.03 3.45 5.26 3.5 ;
        RECT 5.03 3.405 5.21 3.5 ;
        RECT 5.17 3.475 5.46 3.625 ;
        RECT 4.96 3.35 5.17 3.43 ;
        RECT 4.91 3.28 5.1 3.37 ;
        RECT 2.7 3.25 5.03 3.345 ;
        RECT 2.77 3.21 5.03 3.345 ;
        RECT 2.77 3.195 4.96 3.345 ;
        RECT 2.81 3.175 4.96 3.345 ;
        RECT 2.63 3.32 2.86 3.37 ;
        RECT 2.63 3.32 2.81 3.415 ;
        RECT 2.56 3.39 2.77 3.47 ;
        RECT 2.51 3.45 2.7 3.54 ;
        RECT 2.27 3.475 2.63 3.61 ;
        RECT 2.31 3.475 2.56 3.645 ;
        RECT 2.13 3.45 2.36 3.5 ;
        RECT 2.13 3.405 2.31 3.5 ;
        RECT 2.27 3.475 2.56 3.625 ;
        RECT 2.06 3.35 2.27 3.43 ;
        RECT 2.2 3.475 2.63 3.57 ;
        RECT 2.01 3.28 2.2 3.37 ;
        RECT -0.455 3.21 2.13 3.345 ;
        RECT -0.455 3.175 2.06 3.345 ;
    END
  END RWL1_2
  PIN RWL1_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 4.525 34.76 4.72 ;
        RECT 34.53 4.67 34.71 4.765 ;
        RECT 34.6 4.6 34.76 4.72 ;
        RECT 34.67 4.545 34.71 4.765 ;
        RECT 34.46 4.74 34.67 4.82 ;
        RECT 34.41 4.8 34.6 4.89 ;
        RECT 34.17 4.825 34.53 4.96 ;
        RECT 34.21 4.825 34.46 4.995 ;
        RECT 34.03 4.8 34.26 4.85 ;
        RECT 34.03 4.755 34.21 4.85 ;
        RECT 34.17 4.825 34.46 4.975 ;
        RECT 33.96 4.7 34.17 4.78 ;
        RECT 34.1 4.825 34.53 4.92 ;
        RECT 33.91 4.63 34.1 4.72 ;
        RECT 31.7 4.6 34.03 4.695 ;
        RECT 31.77 4.56 34.03 4.695 ;
        RECT 31.77 4.545 33.96 4.695 ;
        RECT 31.81 4.525 33.96 4.695 ;
        RECT 31.63 4.67 31.86 4.72 ;
        RECT 31.63 4.67 31.81 4.765 ;
        RECT 31.56 4.74 31.77 4.82 ;
        RECT 31.51 4.8 31.7 4.89 ;
        RECT 31.27 4.825 31.63 4.96 ;
        RECT 31.31 4.825 31.56 4.995 ;
        RECT 31.13 4.8 31.36 4.85 ;
        RECT 31.13 4.755 31.31 4.85 ;
        RECT 31.27 4.825 31.56 4.975 ;
        RECT 31.06 4.7 31.27 4.78 ;
        RECT 31.2 4.825 31.63 4.92 ;
        RECT 31.01 4.63 31.2 4.72 ;
        RECT 28.725 4.56 31.13 4.695 ;
        RECT 28.725 4.525 31.06 4.695 ;
        RECT 28.74 4.525 28.96 4.7 ;
        RECT 28.74 4.525 28.95 4.74 ;
        RECT 28.3 4.825 28.74 4.92 ;
        RECT 28.61 4.8 28.81 4.88 ;
        RECT 28.73 4.7 28.74 4.92 ;
        RECT 28.37 4.825 28.73 4.96 ;
        RECT 28.66 4.74 28.88 4.81 ;
        RECT 28.41 4.825 28.66 4.995 ;
        RECT 28.23 4.8 28.46 4.85 ;
        RECT 28.23 4.755 28.41 4.85 ;
        RECT 28.37 4.825 28.66 4.975 ;
        RECT 28.16 4.7 28.37 4.78 ;
        RECT 28.11 4.63 28.3 4.72 ;
        RECT 25.9 4.6 28.23 4.695 ;
        RECT 25.97 4.56 28.23 4.695 ;
        RECT 25.97 4.545 28.16 4.695 ;
        RECT 26.01 4.525 28.16 4.695 ;
        RECT 25.83 4.67 26.06 4.72 ;
        RECT 25.83 4.67 26.01 4.765 ;
        RECT 25.76 4.74 25.97 4.82 ;
        RECT 25.71 4.8 25.9 4.89 ;
        RECT 25.47 4.825 25.83 4.96 ;
        RECT 25.51 4.825 25.76 4.995 ;
        RECT 25.33 4.8 25.56 4.85 ;
        RECT 25.33 4.755 25.51 4.85 ;
        RECT 25.47 4.825 25.76 4.975 ;
        RECT 25.26 4.7 25.47 4.78 ;
        RECT 25.4 4.825 25.83 4.92 ;
        RECT 25.21 4.63 25.4 4.72 ;
        RECT 22.925 4.56 25.33 4.695 ;
        RECT 22.925 4.525 25.26 4.695 ;
        RECT 22.94 4.525 23.16 4.7 ;
        RECT 22.94 4.525 23.15 4.74 ;
        RECT 22.5 4.825 22.94 4.92 ;
        RECT 22.81 4.8 23.01 4.88 ;
        RECT 22.93 4.7 22.94 4.92 ;
        RECT 22.57 4.825 22.93 4.96 ;
        RECT 22.86 4.74 23.08 4.81 ;
        RECT 22.61 4.825 22.86 4.995 ;
        RECT 22.43 4.8 22.66 4.85 ;
        RECT 22.43 4.755 22.61 4.85 ;
        RECT 22.57 4.825 22.86 4.975 ;
        RECT 22.36 4.7 22.57 4.78 ;
        RECT 22.31 4.63 22.5 4.72 ;
        RECT 20.1 4.6 22.43 4.695 ;
        RECT 20.17 4.56 22.43 4.695 ;
        RECT 20.17 4.545 22.36 4.695 ;
        RECT 20.21 4.525 22.36 4.695 ;
        RECT 20.03 4.67 20.26 4.72 ;
        RECT 20.03 4.67 20.21 4.765 ;
        RECT 19.96 4.74 20.17 4.82 ;
        RECT 19.91 4.8 20.1 4.89 ;
        RECT 19.67 4.825 20.03 4.96 ;
        RECT 19.71 4.825 19.96 4.995 ;
        RECT 19.53 4.8 19.76 4.85 ;
        RECT 19.53 4.755 19.71 4.85 ;
        RECT 19.67 4.825 19.96 4.975 ;
        RECT 19.46 4.7 19.67 4.78 ;
        RECT 19.6 4.825 20.03 4.92 ;
        RECT 19.41 4.63 19.6 4.72 ;
        RECT 17.125 4.56 19.53 4.695 ;
        RECT 17.125 4.525 19.46 4.695 ;
        RECT 17.14 4.525 17.36 4.7 ;
        RECT 17.14 4.525 17.35 4.74 ;
        RECT 16.7 4.825 17.14 4.92 ;
        RECT 17.01 4.8 17.21 4.88 ;
        RECT 17.13 4.7 17.14 4.92 ;
        RECT 16.77 4.825 17.13 4.96 ;
        RECT 17.06 4.74 17.28 4.81 ;
        RECT 16.81 4.825 17.06 4.995 ;
        RECT 16.63 4.8 16.86 4.85 ;
        RECT 16.63 4.755 16.81 4.85 ;
        RECT 16.77 4.825 17.06 4.975 ;
        RECT 16.56 4.7 16.77 4.78 ;
        RECT 16.51 4.63 16.7 4.72 ;
        RECT 14.3 4.6 16.63 4.695 ;
        RECT 14.37 4.56 16.63 4.695 ;
        RECT 14.37 4.545 16.56 4.695 ;
        RECT 14.41 4.525 16.56 4.695 ;
        RECT 14.23 4.67 14.46 4.72 ;
        RECT 14.23 4.67 14.41 4.765 ;
        RECT 14.16 4.74 14.37 4.82 ;
        RECT 14.11 4.8 14.3 4.89 ;
        RECT 13.87 4.825 14.23 4.96 ;
        RECT 13.91 4.825 14.16 4.995 ;
        RECT 13.73 4.8 13.96 4.85 ;
        RECT 13.73 4.755 13.91 4.85 ;
        RECT 13.87 4.825 14.16 4.975 ;
        RECT 13.66 4.7 13.87 4.78 ;
        RECT 13.8 4.825 14.23 4.92 ;
        RECT 13.61 4.63 13.8 4.72 ;
        RECT 11.325 4.56 13.73 4.695 ;
        RECT 11.325 4.525 13.66 4.695 ;
        RECT 11.34 4.525 11.56 4.7 ;
        RECT 11.34 4.525 11.55 4.74 ;
        RECT 10.9 4.825 11.34 4.92 ;
        RECT 11.21 4.8 11.41 4.88 ;
        RECT 11.33 4.7 11.34 4.92 ;
        RECT 10.97 4.825 11.33 4.96 ;
        RECT 11.26 4.74 11.48 4.81 ;
        RECT 11.01 4.825 11.26 4.995 ;
        RECT 10.83 4.8 11.06 4.85 ;
        RECT 10.83 4.755 11.01 4.85 ;
        RECT 10.97 4.825 11.26 4.975 ;
        RECT 10.76 4.7 10.97 4.78 ;
        RECT 10.71 4.63 10.9 4.72 ;
        RECT 8.5 4.6 10.83 4.695 ;
        RECT 8.57 4.56 10.83 4.695 ;
        RECT 8.57 4.545 10.76 4.695 ;
        RECT 8.61 4.525 10.76 4.695 ;
        RECT 8.43 4.67 8.66 4.72 ;
        RECT 8.43 4.67 8.61 4.765 ;
        RECT 8.36 4.74 8.57 4.82 ;
        RECT 8.31 4.8 8.5 4.89 ;
        RECT 8.07 4.825 8.43 4.96 ;
        RECT 8.11 4.825 8.36 4.995 ;
        RECT 7.93 4.8 8.16 4.85 ;
        RECT 7.93 4.755 8.11 4.85 ;
        RECT 8.07 4.825 8.36 4.975 ;
        RECT 7.86 4.7 8.07 4.78 ;
        RECT 8 4.825 8.43 4.92 ;
        RECT 7.81 4.63 8 4.72 ;
        RECT 5.525 4.56 7.93 4.695 ;
        RECT 5.525 4.525 7.86 4.695 ;
        RECT 5.54 4.525 5.76 4.7 ;
        RECT 5.54 4.525 5.75 4.74 ;
        RECT 5.1 4.825 5.54 4.92 ;
        RECT 5.41 4.8 5.61 4.88 ;
        RECT 5.53 4.7 5.54 4.92 ;
        RECT 5.17 4.825 5.53 4.96 ;
        RECT 5.46 4.74 5.68 4.81 ;
        RECT 5.21 4.825 5.46 4.995 ;
        RECT 5.03 4.8 5.26 4.85 ;
        RECT 5.03 4.755 5.21 4.85 ;
        RECT 5.17 4.825 5.46 4.975 ;
        RECT 4.96 4.7 5.17 4.78 ;
        RECT 4.91 4.63 5.1 4.72 ;
        RECT 2.7 4.6 5.03 4.695 ;
        RECT 2.77 4.56 5.03 4.695 ;
        RECT 2.77 4.545 4.96 4.695 ;
        RECT 2.81 4.525 4.96 4.695 ;
        RECT 2.63 4.67 2.86 4.72 ;
        RECT 2.63 4.67 2.81 4.765 ;
        RECT 2.56 4.74 2.77 4.82 ;
        RECT 2.51 4.8 2.7 4.89 ;
        RECT 2.27 4.825 2.63 4.96 ;
        RECT 2.31 4.825 2.56 4.995 ;
        RECT 2.13 4.8 2.36 4.85 ;
        RECT 2.13 4.755 2.31 4.85 ;
        RECT 2.27 4.825 2.56 4.975 ;
        RECT 2.06 4.7 2.27 4.78 ;
        RECT 2.2 4.825 2.63 4.92 ;
        RECT 2.01 4.63 2.2 4.72 ;
        RECT -0.455 4.56 2.13 4.695 ;
        RECT -0.455 4.525 2.06 4.695 ;
    END
  END RWL1_3
  PIN RWL1_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 5.875 34.76 6.07 ;
        RECT 34.53 6.02 34.71 6.115 ;
        RECT 34.6 5.95 34.76 6.07 ;
        RECT 34.67 5.895 34.71 6.115 ;
        RECT 34.46 6.09 34.67 6.17 ;
        RECT 34.41 6.15 34.6 6.24 ;
        RECT 34.17 6.175 34.53 6.31 ;
        RECT 34.21 6.175 34.46 6.345 ;
        RECT 34.03 6.15 34.26 6.2 ;
        RECT 34.03 6.105 34.21 6.2 ;
        RECT 34.17 6.175 34.46 6.325 ;
        RECT 33.96 6.05 34.17 6.13 ;
        RECT 34.1 6.175 34.53 6.27 ;
        RECT 33.91 5.98 34.1 6.07 ;
        RECT 31.7 5.95 34.03 6.045 ;
        RECT 31.77 5.91 34.03 6.045 ;
        RECT 31.77 5.895 33.96 6.045 ;
        RECT 31.81 5.875 33.96 6.045 ;
        RECT 31.63 6.02 31.86 6.07 ;
        RECT 31.63 6.02 31.81 6.115 ;
        RECT 31.56 6.09 31.77 6.17 ;
        RECT 31.51 6.15 31.7 6.24 ;
        RECT 31.27 6.175 31.63 6.31 ;
        RECT 31.31 6.175 31.56 6.345 ;
        RECT 31.13 6.15 31.36 6.2 ;
        RECT 31.13 6.105 31.31 6.2 ;
        RECT 31.27 6.175 31.56 6.325 ;
        RECT 31.06 6.05 31.27 6.13 ;
        RECT 31.2 6.175 31.63 6.27 ;
        RECT 31.01 5.98 31.2 6.07 ;
        RECT 28.725 5.91 31.13 6.045 ;
        RECT 28.725 5.875 31.06 6.045 ;
        RECT 28.74 5.875 28.96 6.05 ;
        RECT 28.74 5.875 28.95 6.09 ;
        RECT 28.3 6.175 28.74 6.27 ;
        RECT 28.61 6.15 28.81 6.23 ;
        RECT 28.73 6.05 28.74 6.27 ;
        RECT 28.37 6.175 28.73 6.31 ;
        RECT 28.66 6.09 28.88 6.16 ;
        RECT 28.41 6.175 28.66 6.345 ;
        RECT 28.23 6.15 28.46 6.2 ;
        RECT 28.23 6.105 28.41 6.2 ;
        RECT 28.37 6.175 28.66 6.325 ;
        RECT 28.16 6.05 28.37 6.13 ;
        RECT 28.11 5.98 28.3 6.07 ;
        RECT 25.9 5.95 28.23 6.045 ;
        RECT 25.97 5.91 28.23 6.045 ;
        RECT 25.97 5.895 28.16 6.045 ;
        RECT 26.01 5.875 28.16 6.045 ;
        RECT 25.83 6.02 26.06 6.07 ;
        RECT 25.83 6.02 26.01 6.115 ;
        RECT 25.76 6.09 25.97 6.17 ;
        RECT 25.71 6.15 25.9 6.24 ;
        RECT 25.47 6.175 25.83 6.31 ;
        RECT 25.51 6.175 25.76 6.345 ;
        RECT 25.33 6.15 25.56 6.2 ;
        RECT 25.33 6.105 25.51 6.2 ;
        RECT 25.47 6.175 25.76 6.325 ;
        RECT 25.26 6.05 25.47 6.13 ;
        RECT 25.4 6.175 25.83 6.27 ;
        RECT 25.21 5.98 25.4 6.07 ;
        RECT 22.925 5.91 25.33 6.045 ;
        RECT 22.925 5.875 25.26 6.045 ;
        RECT 22.94 5.875 23.16 6.05 ;
        RECT 22.94 5.875 23.15 6.09 ;
        RECT 22.5 6.175 22.94 6.27 ;
        RECT 22.81 6.15 23.01 6.23 ;
        RECT 22.93 6.05 22.94 6.27 ;
        RECT 22.57 6.175 22.93 6.31 ;
        RECT 22.86 6.09 23.08 6.16 ;
        RECT 22.61 6.175 22.86 6.345 ;
        RECT 22.43 6.15 22.66 6.2 ;
        RECT 22.43 6.105 22.61 6.2 ;
        RECT 22.57 6.175 22.86 6.325 ;
        RECT 22.36 6.05 22.57 6.13 ;
        RECT 22.31 5.98 22.5 6.07 ;
        RECT 20.1 5.95 22.43 6.045 ;
        RECT 20.17 5.91 22.43 6.045 ;
        RECT 20.17 5.895 22.36 6.045 ;
        RECT 20.21 5.875 22.36 6.045 ;
        RECT 20.03 6.02 20.26 6.07 ;
        RECT 20.03 6.02 20.21 6.115 ;
        RECT 19.96 6.09 20.17 6.17 ;
        RECT 19.91 6.15 20.1 6.24 ;
        RECT 19.67 6.175 20.03 6.31 ;
        RECT 19.71 6.175 19.96 6.345 ;
        RECT 19.53 6.15 19.76 6.2 ;
        RECT 19.53 6.105 19.71 6.2 ;
        RECT 19.67 6.175 19.96 6.325 ;
        RECT 19.46 6.05 19.67 6.13 ;
        RECT 19.6 6.175 20.03 6.27 ;
        RECT 19.41 5.98 19.6 6.07 ;
        RECT 17.125 5.91 19.53 6.045 ;
        RECT 17.125 5.875 19.46 6.045 ;
        RECT 17.14 5.875 17.36 6.05 ;
        RECT 17.14 5.875 17.35 6.09 ;
        RECT 16.7 6.175 17.14 6.27 ;
        RECT 17.01 6.15 17.21 6.23 ;
        RECT 17.13 6.05 17.14 6.27 ;
        RECT 16.77 6.175 17.13 6.31 ;
        RECT 17.06 6.09 17.28 6.16 ;
        RECT 16.81 6.175 17.06 6.345 ;
        RECT 16.63 6.15 16.86 6.2 ;
        RECT 16.63 6.105 16.81 6.2 ;
        RECT 16.77 6.175 17.06 6.325 ;
        RECT 16.56 6.05 16.77 6.13 ;
        RECT 16.51 5.98 16.7 6.07 ;
        RECT 14.3 5.95 16.63 6.045 ;
        RECT 14.37 5.91 16.63 6.045 ;
        RECT 14.37 5.895 16.56 6.045 ;
        RECT 14.41 5.875 16.56 6.045 ;
        RECT 14.23 6.02 14.46 6.07 ;
        RECT 14.23 6.02 14.41 6.115 ;
        RECT 14.16 6.09 14.37 6.17 ;
        RECT 14.11 6.15 14.3 6.24 ;
        RECT 13.87 6.175 14.23 6.31 ;
        RECT 13.91 6.175 14.16 6.345 ;
        RECT 13.73 6.15 13.96 6.2 ;
        RECT 13.73 6.105 13.91 6.2 ;
        RECT 13.87 6.175 14.16 6.325 ;
        RECT 13.66 6.05 13.87 6.13 ;
        RECT 13.8 6.175 14.23 6.27 ;
        RECT 13.61 5.98 13.8 6.07 ;
        RECT 11.325 5.91 13.73 6.045 ;
        RECT 11.325 5.875 13.66 6.045 ;
        RECT 11.34 5.875 11.56 6.05 ;
        RECT 11.34 5.875 11.55 6.09 ;
        RECT 10.9 6.175 11.34 6.27 ;
        RECT 11.21 6.15 11.41 6.23 ;
        RECT 11.33 6.05 11.34 6.27 ;
        RECT 10.97 6.175 11.33 6.31 ;
        RECT 11.26 6.09 11.48 6.16 ;
        RECT 11.01 6.175 11.26 6.345 ;
        RECT 10.83 6.15 11.06 6.2 ;
        RECT 10.83 6.105 11.01 6.2 ;
        RECT 10.97 6.175 11.26 6.325 ;
        RECT 10.76 6.05 10.97 6.13 ;
        RECT 10.71 5.98 10.9 6.07 ;
        RECT 8.5 5.95 10.83 6.045 ;
        RECT 8.57 5.91 10.83 6.045 ;
        RECT 8.57 5.895 10.76 6.045 ;
        RECT 8.61 5.875 10.76 6.045 ;
        RECT 8.43 6.02 8.66 6.07 ;
        RECT 8.43 6.02 8.61 6.115 ;
        RECT 8.36 6.09 8.57 6.17 ;
        RECT 8.31 6.15 8.5 6.24 ;
        RECT 8.07 6.175 8.43 6.31 ;
        RECT 8.11 6.175 8.36 6.345 ;
        RECT 7.93 6.15 8.16 6.2 ;
        RECT 7.93 6.105 8.11 6.2 ;
        RECT 8.07 6.175 8.36 6.325 ;
        RECT 7.86 6.05 8.07 6.13 ;
        RECT 8 6.175 8.43 6.27 ;
        RECT 7.81 5.98 8 6.07 ;
        RECT 5.525 5.91 7.93 6.045 ;
        RECT 5.525 5.875 7.86 6.045 ;
        RECT 5.54 5.875 5.76 6.05 ;
        RECT 5.54 5.875 5.75 6.09 ;
        RECT 5.1 6.175 5.54 6.27 ;
        RECT 5.41 6.15 5.61 6.23 ;
        RECT 5.53 6.05 5.54 6.27 ;
        RECT 5.17 6.175 5.53 6.31 ;
        RECT 5.46 6.09 5.68 6.16 ;
        RECT 5.21 6.175 5.46 6.345 ;
        RECT 5.03 6.15 5.26 6.2 ;
        RECT 5.03 6.105 5.21 6.2 ;
        RECT 5.17 6.175 5.46 6.325 ;
        RECT 4.96 6.05 5.17 6.13 ;
        RECT 4.91 5.98 5.1 6.07 ;
        RECT 2.7 5.95 5.03 6.045 ;
        RECT 2.77 5.91 5.03 6.045 ;
        RECT 2.77 5.895 4.96 6.045 ;
        RECT 2.81 5.875 4.96 6.045 ;
        RECT 2.63 6.02 2.86 6.07 ;
        RECT 2.63 6.02 2.81 6.115 ;
        RECT 2.56 6.09 2.77 6.17 ;
        RECT 2.51 6.15 2.7 6.24 ;
        RECT 2.27 6.175 2.63 6.31 ;
        RECT 2.31 6.175 2.56 6.345 ;
        RECT 2.13 6.15 2.36 6.2 ;
        RECT 2.13 6.105 2.31 6.2 ;
        RECT 2.27 6.175 2.56 6.325 ;
        RECT 2.06 6.05 2.27 6.13 ;
        RECT 2.2 6.175 2.63 6.27 ;
        RECT 2.01 5.98 2.2 6.07 ;
        RECT -0.455 5.91 2.13 6.045 ;
        RECT -0.455 5.875 2.06 6.045 ;
    END
  END RWL1_4
  PIN RWL1_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 7.225 34.76 7.42 ;
        RECT 34.53 7.37 34.71 7.465 ;
        RECT 34.6 7.3 34.76 7.42 ;
        RECT 34.67 7.245 34.71 7.465 ;
        RECT 34.46 7.44 34.67 7.52 ;
        RECT 34.41 7.5 34.6 7.59 ;
        RECT 34.17 7.525 34.53 7.66 ;
        RECT 34.21 7.525 34.46 7.695 ;
        RECT 34.03 7.5 34.26 7.55 ;
        RECT 34.03 7.455 34.21 7.55 ;
        RECT 34.17 7.525 34.46 7.675 ;
        RECT 33.96 7.4 34.17 7.48 ;
        RECT 34.1 7.525 34.53 7.62 ;
        RECT 33.91 7.33 34.1 7.42 ;
        RECT 31.7 7.3 34.03 7.395 ;
        RECT 31.77 7.26 34.03 7.395 ;
        RECT 31.77 7.245 33.96 7.395 ;
        RECT 31.81 7.225 33.96 7.395 ;
        RECT 31.63 7.37 31.86 7.42 ;
        RECT 31.63 7.37 31.81 7.465 ;
        RECT 31.56 7.44 31.77 7.52 ;
        RECT 31.51 7.5 31.7 7.59 ;
        RECT 31.27 7.525 31.63 7.66 ;
        RECT 31.31 7.525 31.56 7.695 ;
        RECT 31.13 7.5 31.36 7.55 ;
        RECT 31.13 7.455 31.31 7.55 ;
        RECT 31.27 7.525 31.56 7.675 ;
        RECT 31.06 7.4 31.27 7.48 ;
        RECT 31.2 7.525 31.63 7.62 ;
        RECT 31.01 7.33 31.2 7.42 ;
        RECT 28.725 7.26 31.13 7.395 ;
        RECT 28.725 7.225 31.06 7.395 ;
        RECT 28.74 7.225 28.96 7.4 ;
        RECT 28.74 7.225 28.95 7.44 ;
        RECT 28.3 7.525 28.74 7.62 ;
        RECT 28.61 7.5 28.81 7.58 ;
        RECT 28.73 7.4 28.74 7.62 ;
        RECT 28.37 7.525 28.73 7.66 ;
        RECT 28.66 7.44 28.88 7.51 ;
        RECT 28.41 7.525 28.66 7.695 ;
        RECT 28.23 7.5 28.46 7.55 ;
        RECT 28.23 7.455 28.41 7.55 ;
        RECT 28.37 7.525 28.66 7.675 ;
        RECT 28.16 7.4 28.37 7.48 ;
        RECT 28.11 7.33 28.3 7.42 ;
        RECT 25.9 7.3 28.23 7.395 ;
        RECT 25.97 7.26 28.23 7.395 ;
        RECT 25.97 7.245 28.16 7.395 ;
        RECT 26.01 7.225 28.16 7.395 ;
        RECT 25.83 7.37 26.06 7.42 ;
        RECT 25.83 7.37 26.01 7.465 ;
        RECT 25.76 7.44 25.97 7.52 ;
        RECT 25.71 7.5 25.9 7.59 ;
        RECT 25.47 7.525 25.83 7.66 ;
        RECT 25.51 7.525 25.76 7.695 ;
        RECT 25.33 7.5 25.56 7.55 ;
        RECT 25.33 7.455 25.51 7.55 ;
        RECT 25.47 7.525 25.76 7.675 ;
        RECT 25.26 7.4 25.47 7.48 ;
        RECT 25.4 7.525 25.83 7.62 ;
        RECT 25.21 7.33 25.4 7.42 ;
        RECT 22.925 7.26 25.33 7.395 ;
        RECT 22.925 7.225 25.26 7.395 ;
        RECT 22.94 7.225 23.16 7.4 ;
        RECT 22.94 7.225 23.15 7.44 ;
        RECT 22.5 7.525 22.94 7.62 ;
        RECT 22.81 7.5 23.01 7.58 ;
        RECT 22.93 7.4 22.94 7.62 ;
        RECT 22.57 7.525 22.93 7.66 ;
        RECT 22.86 7.44 23.08 7.51 ;
        RECT 22.61 7.525 22.86 7.695 ;
        RECT 22.43 7.5 22.66 7.55 ;
        RECT 22.43 7.455 22.61 7.55 ;
        RECT 22.57 7.525 22.86 7.675 ;
        RECT 22.36 7.4 22.57 7.48 ;
        RECT 22.31 7.33 22.5 7.42 ;
        RECT 20.1 7.3 22.43 7.395 ;
        RECT 20.17 7.26 22.43 7.395 ;
        RECT 20.17 7.245 22.36 7.395 ;
        RECT 20.21 7.225 22.36 7.395 ;
        RECT 20.03 7.37 20.26 7.42 ;
        RECT 20.03 7.37 20.21 7.465 ;
        RECT 19.96 7.44 20.17 7.52 ;
        RECT 19.91 7.5 20.1 7.59 ;
        RECT 19.67 7.525 20.03 7.66 ;
        RECT 19.71 7.525 19.96 7.695 ;
        RECT 19.53 7.5 19.76 7.55 ;
        RECT 19.53 7.455 19.71 7.55 ;
        RECT 19.67 7.525 19.96 7.675 ;
        RECT 19.46 7.4 19.67 7.48 ;
        RECT 19.6 7.525 20.03 7.62 ;
        RECT 19.41 7.33 19.6 7.42 ;
        RECT 17.125 7.26 19.53 7.395 ;
        RECT 17.125 7.225 19.46 7.395 ;
        RECT 17.14 7.225 17.36 7.4 ;
        RECT 17.14 7.225 17.35 7.44 ;
        RECT 16.7 7.525 17.14 7.62 ;
        RECT 17.01 7.5 17.21 7.58 ;
        RECT 17.13 7.4 17.14 7.62 ;
        RECT 16.77 7.525 17.13 7.66 ;
        RECT 17.06 7.44 17.28 7.51 ;
        RECT 16.81 7.525 17.06 7.695 ;
        RECT 16.63 7.5 16.86 7.55 ;
        RECT 16.63 7.455 16.81 7.55 ;
        RECT 16.77 7.525 17.06 7.675 ;
        RECT 16.56 7.4 16.77 7.48 ;
        RECT 16.51 7.33 16.7 7.42 ;
        RECT 14.3 7.3 16.63 7.395 ;
        RECT 14.37 7.26 16.63 7.395 ;
        RECT 14.37 7.245 16.56 7.395 ;
        RECT 14.41 7.225 16.56 7.395 ;
        RECT 14.23 7.37 14.46 7.42 ;
        RECT 14.23 7.37 14.41 7.465 ;
        RECT 14.16 7.44 14.37 7.52 ;
        RECT 14.11 7.5 14.3 7.59 ;
        RECT 13.87 7.525 14.23 7.66 ;
        RECT 13.91 7.525 14.16 7.695 ;
        RECT 13.73 7.5 13.96 7.55 ;
        RECT 13.73 7.455 13.91 7.55 ;
        RECT 13.87 7.525 14.16 7.675 ;
        RECT 13.66 7.4 13.87 7.48 ;
        RECT 13.8 7.525 14.23 7.62 ;
        RECT 13.61 7.33 13.8 7.42 ;
        RECT 11.325 7.26 13.73 7.395 ;
        RECT 11.325 7.225 13.66 7.395 ;
        RECT 11.34 7.225 11.56 7.4 ;
        RECT 11.34 7.225 11.55 7.44 ;
        RECT 10.9 7.525 11.34 7.62 ;
        RECT 11.21 7.5 11.41 7.58 ;
        RECT 11.33 7.4 11.34 7.62 ;
        RECT 10.97 7.525 11.33 7.66 ;
        RECT 11.26 7.44 11.48 7.51 ;
        RECT 11.01 7.525 11.26 7.695 ;
        RECT 10.83 7.5 11.06 7.55 ;
        RECT 10.83 7.455 11.01 7.55 ;
        RECT 10.97 7.525 11.26 7.675 ;
        RECT 10.76 7.4 10.97 7.48 ;
        RECT 10.71 7.33 10.9 7.42 ;
        RECT 8.5 7.3 10.83 7.395 ;
        RECT 8.57 7.26 10.83 7.395 ;
        RECT 8.57 7.245 10.76 7.395 ;
        RECT 8.61 7.225 10.76 7.395 ;
        RECT 8.43 7.37 8.66 7.42 ;
        RECT 8.43 7.37 8.61 7.465 ;
        RECT 8.36 7.44 8.57 7.52 ;
        RECT 8.31 7.5 8.5 7.59 ;
        RECT 8.07 7.525 8.43 7.66 ;
        RECT 8.11 7.525 8.36 7.695 ;
        RECT 7.93 7.5 8.16 7.55 ;
        RECT 7.93 7.455 8.11 7.55 ;
        RECT 8.07 7.525 8.36 7.675 ;
        RECT 7.86 7.4 8.07 7.48 ;
        RECT 8 7.525 8.43 7.62 ;
        RECT 7.81 7.33 8 7.42 ;
        RECT 5.525 7.26 7.93 7.395 ;
        RECT 5.525 7.225 7.86 7.395 ;
        RECT 5.54 7.225 5.76 7.4 ;
        RECT 5.54 7.225 5.75 7.44 ;
        RECT 5.1 7.525 5.54 7.62 ;
        RECT 5.41 7.5 5.61 7.58 ;
        RECT 5.53 7.4 5.54 7.62 ;
        RECT 5.17 7.525 5.53 7.66 ;
        RECT 5.46 7.44 5.68 7.51 ;
        RECT 5.21 7.525 5.46 7.695 ;
        RECT 5.03 7.5 5.26 7.55 ;
        RECT 5.03 7.455 5.21 7.55 ;
        RECT 5.17 7.525 5.46 7.675 ;
        RECT 4.96 7.4 5.17 7.48 ;
        RECT 4.91 7.33 5.1 7.42 ;
        RECT 2.7 7.3 5.03 7.395 ;
        RECT 2.77 7.26 5.03 7.395 ;
        RECT 2.77 7.245 4.96 7.395 ;
        RECT 2.81 7.225 4.96 7.395 ;
        RECT 2.63 7.37 2.86 7.42 ;
        RECT 2.63 7.37 2.81 7.465 ;
        RECT 2.56 7.44 2.77 7.52 ;
        RECT 2.51 7.5 2.7 7.59 ;
        RECT 2.27 7.525 2.63 7.66 ;
        RECT 2.31 7.525 2.56 7.695 ;
        RECT 2.13 7.5 2.36 7.55 ;
        RECT 2.13 7.455 2.31 7.55 ;
        RECT 2.27 7.525 2.56 7.675 ;
        RECT 2.06 7.4 2.27 7.48 ;
        RECT 2.2 7.525 2.63 7.62 ;
        RECT 2.01 7.33 2.2 7.42 ;
        RECT -0.455 7.26 2.13 7.395 ;
        RECT -0.455 7.225 2.06 7.395 ;
    END
  END RWL1_5
  PIN RWL1_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 8.575 34.76 8.77 ;
        RECT 34.53 8.72 34.71 8.815 ;
        RECT 34.6 8.65 34.76 8.77 ;
        RECT 34.67 8.595 34.71 8.815 ;
        RECT 34.46 8.79 34.67 8.87 ;
        RECT 34.41 8.85 34.6 8.94 ;
        RECT 34.17 8.875 34.53 9.01 ;
        RECT 34.21 8.875 34.46 9.045 ;
        RECT 34.03 8.85 34.26 8.9 ;
        RECT 34.03 8.805 34.21 8.9 ;
        RECT 34.17 8.875 34.46 9.025 ;
        RECT 33.96 8.75 34.17 8.83 ;
        RECT 34.1 8.875 34.53 8.97 ;
        RECT 33.91 8.68 34.1 8.77 ;
        RECT 31.7 8.65 34.03 8.745 ;
        RECT 31.77 8.61 34.03 8.745 ;
        RECT 31.77 8.595 33.96 8.745 ;
        RECT 31.81 8.575 33.96 8.745 ;
        RECT 31.63 8.72 31.86 8.77 ;
        RECT 31.63 8.72 31.81 8.815 ;
        RECT 31.56 8.79 31.77 8.87 ;
        RECT 31.51 8.85 31.7 8.94 ;
        RECT 31.27 8.875 31.63 9.01 ;
        RECT 31.31 8.875 31.56 9.045 ;
        RECT 31.13 8.85 31.36 8.9 ;
        RECT 31.13 8.805 31.31 8.9 ;
        RECT 31.27 8.875 31.56 9.025 ;
        RECT 31.06 8.75 31.27 8.83 ;
        RECT 31.2 8.875 31.63 8.97 ;
        RECT 31.01 8.68 31.2 8.77 ;
        RECT 28.725 8.61 31.13 8.745 ;
        RECT 28.725 8.575 31.06 8.745 ;
        RECT 28.74 8.575 28.96 8.75 ;
        RECT 28.74 8.575 28.95 8.79 ;
        RECT 28.3 8.875 28.74 8.97 ;
        RECT 28.61 8.85 28.81 8.93 ;
        RECT 28.73 8.75 28.74 8.97 ;
        RECT 28.37 8.875 28.73 9.01 ;
        RECT 28.66 8.79 28.88 8.86 ;
        RECT 28.41 8.875 28.66 9.045 ;
        RECT 28.23 8.85 28.46 8.9 ;
        RECT 28.23 8.805 28.41 8.9 ;
        RECT 28.37 8.875 28.66 9.025 ;
        RECT 28.16 8.75 28.37 8.83 ;
        RECT 28.11 8.68 28.3 8.77 ;
        RECT 25.9 8.65 28.23 8.745 ;
        RECT 25.97 8.61 28.23 8.745 ;
        RECT 25.97 8.595 28.16 8.745 ;
        RECT 26.01 8.575 28.16 8.745 ;
        RECT 25.83 8.72 26.06 8.77 ;
        RECT 25.83 8.72 26.01 8.815 ;
        RECT 25.76 8.79 25.97 8.87 ;
        RECT 25.71 8.85 25.9 8.94 ;
        RECT 25.47 8.875 25.83 9.01 ;
        RECT 25.51 8.875 25.76 9.045 ;
        RECT 25.33 8.85 25.56 8.9 ;
        RECT 25.33 8.805 25.51 8.9 ;
        RECT 25.47 8.875 25.76 9.025 ;
        RECT 25.26 8.75 25.47 8.83 ;
        RECT 25.4 8.875 25.83 8.97 ;
        RECT 25.21 8.68 25.4 8.77 ;
        RECT 22.925 8.61 25.33 8.745 ;
        RECT 22.925 8.575 25.26 8.745 ;
        RECT 22.94 8.575 23.16 8.75 ;
        RECT 22.94 8.575 23.15 8.79 ;
        RECT 22.5 8.875 22.94 8.97 ;
        RECT 22.81 8.85 23.01 8.93 ;
        RECT 22.93 8.75 22.94 8.97 ;
        RECT 22.57 8.875 22.93 9.01 ;
        RECT 22.86 8.79 23.08 8.86 ;
        RECT 22.61 8.875 22.86 9.045 ;
        RECT 22.43 8.85 22.66 8.9 ;
        RECT 22.43 8.805 22.61 8.9 ;
        RECT 22.57 8.875 22.86 9.025 ;
        RECT 22.36 8.75 22.57 8.83 ;
        RECT 22.31 8.68 22.5 8.77 ;
        RECT 20.1 8.65 22.43 8.745 ;
        RECT 20.17 8.61 22.43 8.745 ;
        RECT 20.17 8.595 22.36 8.745 ;
        RECT 20.21 8.575 22.36 8.745 ;
        RECT 20.03 8.72 20.26 8.77 ;
        RECT 20.03 8.72 20.21 8.815 ;
        RECT 19.96 8.79 20.17 8.87 ;
        RECT 19.91 8.85 20.1 8.94 ;
        RECT 19.67 8.875 20.03 9.01 ;
        RECT 19.71 8.875 19.96 9.045 ;
        RECT 19.53 8.85 19.76 8.9 ;
        RECT 19.53 8.805 19.71 8.9 ;
        RECT 19.67 8.875 19.96 9.025 ;
        RECT 19.46 8.75 19.67 8.83 ;
        RECT 19.6 8.875 20.03 8.97 ;
        RECT 19.41 8.68 19.6 8.77 ;
        RECT 17.125 8.61 19.53 8.745 ;
        RECT 17.125 8.575 19.46 8.745 ;
        RECT 17.14 8.575 17.36 8.75 ;
        RECT 17.14 8.575 17.35 8.79 ;
        RECT 16.7 8.875 17.14 8.97 ;
        RECT 17.01 8.85 17.21 8.93 ;
        RECT 17.13 8.75 17.14 8.97 ;
        RECT 16.77 8.875 17.13 9.01 ;
        RECT 17.06 8.79 17.28 8.86 ;
        RECT 16.81 8.875 17.06 9.045 ;
        RECT 16.63 8.85 16.86 8.9 ;
        RECT 16.63 8.805 16.81 8.9 ;
        RECT 16.77 8.875 17.06 9.025 ;
        RECT 16.56 8.75 16.77 8.83 ;
        RECT 16.51 8.68 16.7 8.77 ;
        RECT 14.3 8.65 16.63 8.745 ;
        RECT 14.37 8.61 16.63 8.745 ;
        RECT 14.37 8.595 16.56 8.745 ;
        RECT 14.41 8.575 16.56 8.745 ;
        RECT 14.23 8.72 14.46 8.77 ;
        RECT 14.23 8.72 14.41 8.815 ;
        RECT 14.16 8.79 14.37 8.87 ;
        RECT 14.11 8.85 14.3 8.94 ;
        RECT 13.87 8.875 14.23 9.01 ;
        RECT 13.91 8.875 14.16 9.045 ;
        RECT 13.73 8.85 13.96 8.9 ;
        RECT 13.73 8.805 13.91 8.9 ;
        RECT 13.87 8.875 14.16 9.025 ;
        RECT 13.66 8.75 13.87 8.83 ;
        RECT 13.8 8.875 14.23 8.97 ;
        RECT 13.61 8.68 13.8 8.77 ;
        RECT 11.325 8.61 13.73 8.745 ;
        RECT 11.325 8.575 13.66 8.745 ;
        RECT 11.34 8.575 11.56 8.75 ;
        RECT 11.34 8.575 11.55 8.79 ;
        RECT 10.9 8.875 11.34 8.97 ;
        RECT 11.21 8.85 11.41 8.93 ;
        RECT 11.33 8.75 11.34 8.97 ;
        RECT 10.97 8.875 11.33 9.01 ;
        RECT 11.26 8.79 11.48 8.86 ;
        RECT 11.01 8.875 11.26 9.045 ;
        RECT 10.83 8.85 11.06 8.9 ;
        RECT 10.83 8.805 11.01 8.9 ;
        RECT 10.97 8.875 11.26 9.025 ;
        RECT 10.76 8.75 10.97 8.83 ;
        RECT 10.71 8.68 10.9 8.77 ;
        RECT 8.5 8.65 10.83 8.745 ;
        RECT 8.57 8.61 10.83 8.745 ;
        RECT 8.57 8.595 10.76 8.745 ;
        RECT 8.61 8.575 10.76 8.745 ;
        RECT 8.43 8.72 8.66 8.77 ;
        RECT 8.43 8.72 8.61 8.815 ;
        RECT 8.36 8.79 8.57 8.87 ;
        RECT 8.31 8.85 8.5 8.94 ;
        RECT 8.07 8.875 8.43 9.01 ;
        RECT 8.11 8.875 8.36 9.045 ;
        RECT 7.93 8.85 8.16 8.9 ;
        RECT 7.93 8.805 8.11 8.9 ;
        RECT 8.07 8.875 8.36 9.025 ;
        RECT 7.86 8.75 8.07 8.83 ;
        RECT 8 8.875 8.43 8.97 ;
        RECT 7.81 8.68 8 8.77 ;
        RECT 5.525 8.61 7.93 8.745 ;
        RECT 5.525 8.575 7.86 8.745 ;
        RECT 5.54 8.575 5.76 8.75 ;
        RECT 5.54 8.575 5.75 8.79 ;
        RECT 5.1 8.875 5.54 8.97 ;
        RECT 5.41 8.85 5.61 8.93 ;
        RECT 5.53 8.75 5.54 8.97 ;
        RECT 5.17 8.875 5.53 9.01 ;
        RECT 5.46 8.79 5.68 8.86 ;
        RECT 5.21 8.875 5.46 9.045 ;
        RECT 5.03 8.85 5.26 8.9 ;
        RECT 5.03 8.805 5.21 8.9 ;
        RECT 5.17 8.875 5.46 9.025 ;
        RECT 4.96 8.75 5.17 8.83 ;
        RECT 4.91 8.68 5.1 8.77 ;
        RECT 2.7 8.65 5.03 8.745 ;
        RECT 2.77 8.61 5.03 8.745 ;
        RECT 2.77 8.595 4.96 8.745 ;
        RECT 2.81 8.575 4.96 8.745 ;
        RECT 2.63 8.72 2.86 8.77 ;
        RECT 2.63 8.72 2.81 8.815 ;
        RECT 2.56 8.79 2.77 8.87 ;
        RECT 2.51 8.85 2.7 8.94 ;
        RECT 2.27 8.875 2.63 9.01 ;
        RECT 2.31 8.875 2.56 9.045 ;
        RECT 2.13 8.85 2.36 8.9 ;
        RECT 2.13 8.805 2.31 8.9 ;
        RECT 2.27 8.875 2.56 9.025 ;
        RECT 2.06 8.75 2.27 8.83 ;
        RECT 2.2 8.875 2.63 8.97 ;
        RECT 2.01 8.68 2.2 8.77 ;
        RECT -0.455 8.61 2.13 8.745 ;
        RECT -0.455 8.575 2.06 8.745 ;
    END
  END RWL1_6
  PIN RWL1_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 9.925 34.76 10.12 ;
        RECT 34.53 10.07 34.71 10.165 ;
        RECT 34.6 10 34.76 10.12 ;
        RECT 34.67 9.945 34.71 10.165 ;
        RECT 34.46 10.14 34.67 10.22 ;
        RECT 34.41 10.2 34.6 10.29 ;
        RECT 34.17 10.225 34.53 10.36 ;
        RECT 34.21 10.225 34.46 10.395 ;
        RECT 34.03 10.2 34.26 10.25 ;
        RECT 34.03 10.155 34.21 10.25 ;
        RECT 34.17 10.225 34.46 10.375 ;
        RECT 33.96 10.1 34.17 10.18 ;
        RECT 34.1 10.225 34.53 10.32 ;
        RECT 33.91 10.03 34.1 10.12 ;
        RECT 31.7 10 34.03 10.095 ;
        RECT 31.77 9.96 34.03 10.095 ;
        RECT 31.77 9.945 33.96 10.095 ;
        RECT 31.81 9.925 33.96 10.095 ;
        RECT 31.63 10.07 31.86 10.12 ;
        RECT 31.63 10.07 31.81 10.165 ;
        RECT 31.56 10.14 31.77 10.22 ;
        RECT 31.51 10.2 31.7 10.29 ;
        RECT 31.27 10.225 31.63 10.36 ;
        RECT 31.31 10.225 31.56 10.395 ;
        RECT 31.13 10.2 31.36 10.25 ;
        RECT 31.13 10.155 31.31 10.25 ;
        RECT 31.27 10.225 31.56 10.375 ;
        RECT 31.06 10.1 31.27 10.18 ;
        RECT 31.2 10.225 31.63 10.32 ;
        RECT 31.01 10.03 31.2 10.12 ;
        RECT 28.725 9.96 31.13 10.095 ;
        RECT 28.725 9.925 31.06 10.095 ;
        RECT 28.74 9.925 28.96 10.1 ;
        RECT 28.74 9.925 28.95 10.14 ;
        RECT 28.3 10.225 28.74 10.32 ;
        RECT 28.61 10.2 28.81 10.28 ;
        RECT 28.73 10.1 28.74 10.32 ;
        RECT 28.37 10.225 28.73 10.36 ;
        RECT 28.66 10.14 28.88 10.21 ;
        RECT 28.41 10.225 28.66 10.395 ;
        RECT 28.23 10.2 28.46 10.25 ;
        RECT 28.23 10.155 28.41 10.25 ;
        RECT 28.37 10.225 28.66 10.375 ;
        RECT 28.16 10.1 28.37 10.18 ;
        RECT 28.11 10.03 28.3 10.12 ;
        RECT 25.9 10 28.23 10.095 ;
        RECT 25.97 9.96 28.23 10.095 ;
        RECT 25.97 9.945 28.16 10.095 ;
        RECT 26.01 9.925 28.16 10.095 ;
        RECT 25.83 10.07 26.06 10.12 ;
        RECT 25.83 10.07 26.01 10.165 ;
        RECT 25.76 10.14 25.97 10.22 ;
        RECT 25.71 10.2 25.9 10.29 ;
        RECT 25.47 10.225 25.83 10.36 ;
        RECT 25.51 10.225 25.76 10.395 ;
        RECT 25.33 10.2 25.56 10.25 ;
        RECT 25.33 10.155 25.51 10.25 ;
        RECT 25.47 10.225 25.76 10.375 ;
        RECT 25.26 10.1 25.47 10.18 ;
        RECT 25.4 10.225 25.83 10.32 ;
        RECT 25.21 10.03 25.4 10.12 ;
        RECT 22.925 9.96 25.33 10.095 ;
        RECT 22.925 9.925 25.26 10.095 ;
        RECT 22.94 9.925 23.16 10.1 ;
        RECT 22.94 9.925 23.15 10.14 ;
        RECT 22.5 10.225 22.94 10.32 ;
        RECT 22.81 10.2 23.01 10.28 ;
        RECT 22.93 10.1 22.94 10.32 ;
        RECT 22.57 10.225 22.93 10.36 ;
        RECT 22.86 10.14 23.08 10.21 ;
        RECT 22.61 10.225 22.86 10.395 ;
        RECT 22.43 10.2 22.66 10.25 ;
        RECT 22.43 10.155 22.61 10.25 ;
        RECT 22.57 10.225 22.86 10.375 ;
        RECT 22.36 10.1 22.57 10.18 ;
        RECT 22.31 10.03 22.5 10.12 ;
        RECT 20.1 10 22.43 10.095 ;
        RECT 20.17 9.96 22.43 10.095 ;
        RECT 20.17 9.945 22.36 10.095 ;
        RECT 20.21 9.925 22.36 10.095 ;
        RECT 20.03 10.07 20.26 10.12 ;
        RECT 20.03 10.07 20.21 10.165 ;
        RECT 19.96 10.14 20.17 10.22 ;
        RECT 19.91 10.2 20.1 10.29 ;
        RECT 19.67 10.225 20.03 10.36 ;
        RECT 19.71 10.225 19.96 10.395 ;
        RECT 19.53 10.2 19.76 10.25 ;
        RECT 19.53 10.155 19.71 10.25 ;
        RECT 19.67 10.225 19.96 10.375 ;
        RECT 19.46 10.1 19.67 10.18 ;
        RECT 19.6 10.225 20.03 10.32 ;
        RECT 19.41 10.03 19.6 10.12 ;
        RECT 17.125 9.96 19.53 10.095 ;
        RECT 17.125 9.925 19.46 10.095 ;
        RECT 17.14 9.925 17.36 10.1 ;
        RECT 17.14 9.925 17.35 10.14 ;
        RECT 16.7 10.225 17.14 10.32 ;
        RECT 17.01 10.2 17.21 10.28 ;
        RECT 17.13 10.1 17.14 10.32 ;
        RECT 16.77 10.225 17.13 10.36 ;
        RECT 17.06 10.14 17.28 10.21 ;
        RECT 16.81 10.225 17.06 10.395 ;
        RECT 16.63 10.2 16.86 10.25 ;
        RECT 16.63 10.155 16.81 10.25 ;
        RECT 16.77 10.225 17.06 10.375 ;
        RECT 16.56 10.1 16.77 10.18 ;
        RECT 16.51 10.03 16.7 10.12 ;
        RECT 14.3 10 16.63 10.095 ;
        RECT 14.37 9.96 16.63 10.095 ;
        RECT 14.37 9.945 16.56 10.095 ;
        RECT 14.41 9.925 16.56 10.095 ;
        RECT 14.23 10.07 14.46 10.12 ;
        RECT 14.23 10.07 14.41 10.165 ;
        RECT 14.16 10.14 14.37 10.22 ;
        RECT 14.11 10.2 14.3 10.29 ;
        RECT 13.87 10.225 14.23 10.36 ;
        RECT 13.91 10.225 14.16 10.395 ;
        RECT 13.73 10.2 13.96 10.25 ;
        RECT 13.73 10.155 13.91 10.25 ;
        RECT 13.87 10.225 14.16 10.375 ;
        RECT 13.66 10.1 13.87 10.18 ;
        RECT 13.8 10.225 14.23 10.32 ;
        RECT 13.61 10.03 13.8 10.12 ;
        RECT 11.325 9.96 13.73 10.095 ;
        RECT 11.325 9.925 13.66 10.095 ;
        RECT 11.34 9.925 11.56 10.1 ;
        RECT 11.34 9.925 11.55 10.14 ;
        RECT 10.9 10.225 11.34 10.32 ;
        RECT 11.21 10.2 11.41 10.28 ;
        RECT 11.33 10.1 11.34 10.32 ;
        RECT 10.97 10.225 11.33 10.36 ;
        RECT 11.26 10.14 11.48 10.21 ;
        RECT 11.01 10.225 11.26 10.395 ;
        RECT 10.83 10.2 11.06 10.25 ;
        RECT 10.83 10.155 11.01 10.25 ;
        RECT 10.97 10.225 11.26 10.375 ;
        RECT 10.76 10.1 10.97 10.18 ;
        RECT 10.71 10.03 10.9 10.12 ;
        RECT 8.5 10 10.83 10.095 ;
        RECT 8.57 9.96 10.83 10.095 ;
        RECT 8.57 9.945 10.76 10.095 ;
        RECT 8.61 9.925 10.76 10.095 ;
        RECT 8.43 10.07 8.66 10.12 ;
        RECT 8.43 10.07 8.61 10.165 ;
        RECT 8.36 10.14 8.57 10.22 ;
        RECT 8.31 10.2 8.5 10.29 ;
        RECT 8.07 10.225 8.43 10.36 ;
        RECT 8.11 10.225 8.36 10.395 ;
        RECT 7.93 10.2 8.16 10.25 ;
        RECT 7.93 10.155 8.11 10.25 ;
        RECT 8.07 10.225 8.36 10.375 ;
        RECT 7.86 10.1 8.07 10.18 ;
        RECT 8 10.225 8.43 10.32 ;
        RECT 7.81 10.03 8 10.12 ;
        RECT 5.525 9.96 7.93 10.095 ;
        RECT 5.525 9.925 7.86 10.095 ;
        RECT 5.54 9.925 5.76 10.1 ;
        RECT 5.54 9.925 5.75 10.14 ;
        RECT 5.1 10.225 5.54 10.32 ;
        RECT 5.41 10.2 5.61 10.28 ;
        RECT 5.53 10.1 5.54 10.32 ;
        RECT 5.17 10.225 5.53 10.36 ;
        RECT 5.46 10.14 5.68 10.21 ;
        RECT 5.21 10.225 5.46 10.395 ;
        RECT 5.03 10.2 5.26 10.25 ;
        RECT 5.03 10.155 5.21 10.25 ;
        RECT 5.17 10.225 5.46 10.375 ;
        RECT 4.96 10.1 5.17 10.18 ;
        RECT 4.91 10.03 5.1 10.12 ;
        RECT 2.7 10 5.03 10.095 ;
        RECT 2.77 9.96 5.03 10.095 ;
        RECT 2.77 9.945 4.96 10.095 ;
        RECT 2.81 9.925 4.96 10.095 ;
        RECT 2.63 10.07 2.86 10.12 ;
        RECT 2.63 10.07 2.81 10.165 ;
        RECT 2.56 10.14 2.77 10.22 ;
        RECT 2.51 10.2 2.7 10.29 ;
        RECT 2.27 10.225 2.63 10.36 ;
        RECT 2.31 10.225 2.56 10.395 ;
        RECT 2.13 10.2 2.36 10.25 ;
        RECT 2.13 10.155 2.31 10.25 ;
        RECT 2.27 10.225 2.56 10.375 ;
        RECT 2.06 10.1 2.27 10.18 ;
        RECT 2.2 10.225 2.63 10.32 ;
        RECT 2.01 10.03 2.2 10.12 ;
        RECT -0.455 9.96 2.13 10.095 ;
        RECT -0.455 9.925 2.06 10.095 ;
    END
  END RWL1_7
  PIN RWL1_8
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 11.275 34.76 11.47 ;
        RECT 34.53 11.42 34.71 11.515 ;
        RECT 34.6 11.35 34.76 11.47 ;
        RECT 34.67 11.295 34.71 11.515 ;
        RECT 34.46 11.49 34.67 11.57 ;
        RECT 34.41 11.55 34.6 11.64 ;
        RECT 34.17 11.575 34.53 11.71 ;
        RECT 34.21 11.575 34.46 11.745 ;
        RECT 34.03 11.55 34.26 11.6 ;
        RECT 34.03 11.505 34.21 11.6 ;
        RECT 34.17 11.575 34.46 11.725 ;
        RECT 33.96 11.45 34.17 11.53 ;
        RECT 34.1 11.575 34.53 11.67 ;
        RECT 33.91 11.38 34.1 11.47 ;
        RECT 31.7 11.35 34.03 11.445 ;
        RECT 31.77 11.31 34.03 11.445 ;
        RECT 31.77 11.295 33.96 11.445 ;
        RECT 31.81 11.275 33.96 11.445 ;
        RECT 31.63 11.42 31.86 11.47 ;
        RECT 31.63 11.42 31.81 11.515 ;
        RECT 31.56 11.49 31.77 11.57 ;
        RECT 31.51 11.55 31.7 11.64 ;
        RECT 31.27 11.575 31.63 11.71 ;
        RECT 31.31 11.575 31.56 11.745 ;
        RECT 31.13 11.55 31.36 11.6 ;
        RECT 31.13 11.505 31.31 11.6 ;
        RECT 31.27 11.575 31.56 11.725 ;
        RECT 31.06 11.45 31.27 11.53 ;
        RECT 31.2 11.575 31.63 11.67 ;
        RECT 31.01 11.38 31.2 11.47 ;
        RECT 28.725 11.31 31.13 11.445 ;
        RECT 28.725 11.275 31.06 11.445 ;
        RECT 28.74 11.275 28.96 11.45 ;
        RECT 28.74 11.275 28.95 11.49 ;
        RECT 28.3 11.575 28.74 11.67 ;
        RECT 28.61 11.55 28.81 11.63 ;
        RECT 28.73 11.45 28.74 11.67 ;
        RECT 28.37 11.575 28.73 11.71 ;
        RECT 28.66 11.49 28.88 11.56 ;
        RECT 28.41 11.575 28.66 11.745 ;
        RECT 28.23 11.55 28.46 11.6 ;
        RECT 28.23 11.505 28.41 11.6 ;
        RECT 28.37 11.575 28.66 11.725 ;
        RECT 28.16 11.45 28.37 11.53 ;
        RECT 28.11 11.38 28.3 11.47 ;
        RECT 25.9 11.35 28.23 11.445 ;
        RECT 25.97 11.31 28.23 11.445 ;
        RECT 25.97 11.295 28.16 11.445 ;
        RECT 26.01 11.275 28.16 11.445 ;
        RECT 25.83 11.42 26.06 11.47 ;
        RECT 25.83 11.42 26.01 11.515 ;
        RECT 25.76 11.49 25.97 11.57 ;
        RECT 25.71 11.55 25.9 11.64 ;
        RECT 25.47 11.575 25.83 11.71 ;
        RECT 25.51 11.575 25.76 11.745 ;
        RECT 25.33 11.55 25.56 11.6 ;
        RECT 25.33 11.505 25.51 11.6 ;
        RECT 25.47 11.575 25.76 11.725 ;
        RECT 25.26 11.45 25.47 11.53 ;
        RECT 25.4 11.575 25.83 11.67 ;
        RECT 25.21 11.38 25.4 11.47 ;
        RECT 22.925 11.31 25.33 11.445 ;
        RECT 22.925 11.275 25.26 11.445 ;
        RECT 22.94 11.275 23.16 11.45 ;
        RECT 22.94 11.275 23.15 11.49 ;
        RECT 22.5 11.575 22.94 11.67 ;
        RECT 22.81 11.55 23.01 11.63 ;
        RECT 22.93 11.45 22.94 11.67 ;
        RECT 22.57 11.575 22.93 11.71 ;
        RECT 22.86 11.49 23.08 11.56 ;
        RECT 22.61 11.575 22.86 11.745 ;
        RECT 22.43 11.55 22.66 11.6 ;
        RECT 22.43 11.505 22.61 11.6 ;
        RECT 22.57 11.575 22.86 11.725 ;
        RECT 22.36 11.45 22.57 11.53 ;
        RECT 22.31 11.38 22.5 11.47 ;
        RECT 20.1 11.35 22.43 11.445 ;
        RECT 20.17 11.31 22.43 11.445 ;
        RECT 20.17 11.295 22.36 11.445 ;
        RECT 20.21 11.275 22.36 11.445 ;
        RECT 20.03 11.42 20.26 11.47 ;
        RECT 20.03 11.42 20.21 11.515 ;
        RECT 19.96 11.49 20.17 11.57 ;
        RECT 19.91 11.55 20.1 11.64 ;
        RECT 19.67 11.575 20.03 11.71 ;
        RECT 19.71 11.575 19.96 11.745 ;
        RECT 19.53 11.55 19.76 11.6 ;
        RECT 19.53 11.505 19.71 11.6 ;
        RECT 19.67 11.575 19.96 11.725 ;
        RECT 19.46 11.45 19.67 11.53 ;
        RECT 19.6 11.575 20.03 11.67 ;
        RECT 19.41 11.38 19.6 11.47 ;
        RECT 17.125 11.31 19.53 11.445 ;
        RECT 17.125 11.275 19.46 11.445 ;
        RECT 17.14 11.275 17.36 11.45 ;
        RECT 17.14 11.275 17.35 11.49 ;
        RECT 16.7 11.575 17.14 11.67 ;
        RECT 17.01 11.55 17.21 11.63 ;
        RECT 17.13 11.45 17.14 11.67 ;
        RECT 16.77 11.575 17.13 11.71 ;
        RECT 17.06 11.49 17.28 11.56 ;
        RECT 16.81 11.575 17.06 11.745 ;
        RECT 16.63 11.55 16.86 11.6 ;
        RECT 16.63 11.505 16.81 11.6 ;
        RECT 16.77 11.575 17.06 11.725 ;
        RECT 16.56 11.45 16.77 11.53 ;
        RECT 16.51 11.38 16.7 11.47 ;
        RECT 14.3 11.35 16.63 11.445 ;
        RECT 14.37 11.31 16.63 11.445 ;
        RECT 14.37 11.295 16.56 11.445 ;
        RECT 14.41 11.275 16.56 11.445 ;
        RECT 14.23 11.42 14.46 11.47 ;
        RECT 14.23 11.42 14.41 11.515 ;
        RECT 14.16 11.49 14.37 11.57 ;
        RECT 14.11 11.55 14.3 11.64 ;
        RECT 13.87 11.575 14.23 11.71 ;
        RECT 13.91 11.575 14.16 11.745 ;
        RECT 13.73 11.55 13.96 11.6 ;
        RECT 13.73 11.505 13.91 11.6 ;
        RECT 13.87 11.575 14.16 11.725 ;
        RECT 13.66 11.45 13.87 11.53 ;
        RECT 13.8 11.575 14.23 11.67 ;
        RECT 13.61 11.38 13.8 11.47 ;
        RECT 11.325 11.31 13.73 11.445 ;
        RECT 11.325 11.275 13.66 11.445 ;
        RECT 11.34 11.275 11.56 11.45 ;
        RECT 11.34 11.275 11.55 11.49 ;
        RECT 10.9 11.575 11.34 11.67 ;
        RECT 11.21 11.55 11.41 11.63 ;
        RECT 11.33 11.45 11.34 11.67 ;
        RECT 10.97 11.575 11.33 11.71 ;
        RECT 11.26 11.49 11.48 11.56 ;
        RECT 11.01 11.575 11.26 11.745 ;
        RECT 10.83 11.55 11.06 11.6 ;
        RECT 10.83 11.505 11.01 11.6 ;
        RECT 10.97 11.575 11.26 11.725 ;
        RECT 10.76 11.45 10.97 11.53 ;
        RECT 10.71 11.38 10.9 11.47 ;
        RECT 8.5 11.35 10.83 11.445 ;
        RECT 8.57 11.31 10.83 11.445 ;
        RECT 8.57 11.295 10.76 11.445 ;
        RECT 8.61 11.275 10.76 11.445 ;
        RECT 8.43 11.42 8.66 11.47 ;
        RECT 8.43 11.42 8.61 11.515 ;
        RECT 8.36 11.49 8.57 11.57 ;
        RECT 8.31 11.55 8.5 11.64 ;
        RECT 8.07 11.575 8.43 11.71 ;
        RECT 8.11 11.575 8.36 11.745 ;
        RECT 7.93 11.55 8.16 11.6 ;
        RECT 7.93 11.505 8.11 11.6 ;
        RECT 8.07 11.575 8.36 11.725 ;
        RECT 7.86 11.45 8.07 11.53 ;
        RECT 8 11.575 8.43 11.67 ;
        RECT 7.81 11.38 8 11.47 ;
        RECT 5.525 11.31 7.93 11.445 ;
        RECT 5.525 11.275 7.86 11.445 ;
        RECT 5.54 11.275 5.76 11.45 ;
        RECT 5.54 11.275 5.75 11.49 ;
        RECT 5.1 11.575 5.54 11.67 ;
        RECT 5.41 11.55 5.61 11.63 ;
        RECT 5.53 11.45 5.54 11.67 ;
        RECT 5.17 11.575 5.53 11.71 ;
        RECT 5.46 11.49 5.68 11.56 ;
        RECT 5.21 11.575 5.46 11.745 ;
        RECT 5.03 11.55 5.26 11.6 ;
        RECT 5.03 11.505 5.21 11.6 ;
        RECT 5.17 11.575 5.46 11.725 ;
        RECT 4.96 11.45 5.17 11.53 ;
        RECT 4.91 11.38 5.1 11.47 ;
        RECT 2.7 11.35 5.03 11.445 ;
        RECT 2.77 11.31 5.03 11.445 ;
        RECT 2.77 11.295 4.96 11.445 ;
        RECT 2.81 11.275 4.96 11.445 ;
        RECT 2.63 11.42 2.86 11.47 ;
        RECT 2.63 11.42 2.81 11.515 ;
        RECT 2.56 11.49 2.77 11.57 ;
        RECT 2.51 11.55 2.7 11.64 ;
        RECT 2.27 11.575 2.63 11.71 ;
        RECT 2.31 11.575 2.56 11.745 ;
        RECT 2.13 11.55 2.36 11.6 ;
        RECT 2.13 11.505 2.31 11.6 ;
        RECT 2.27 11.575 2.56 11.725 ;
        RECT 2.06 11.45 2.27 11.53 ;
        RECT 2.2 11.575 2.63 11.67 ;
        RECT 2.01 11.38 2.2 11.47 ;
        RECT -0.455 11.31 2.13 11.445 ;
        RECT -0.455 11.275 2.06 11.445 ;
    END
  END RWL1_8
  PIN RWL1_9
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 34.71 12.625 34.76 12.82 ;
        RECT 34.53 12.77 34.71 12.865 ;
        RECT 34.6 12.7 34.76 12.82 ;
        RECT 34.67 12.645 34.71 12.865 ;
        RECT 34.46 12.84 34.67 12.92 ;
        RECT 34.41 12.9 34.6 12.99 ;
        RECT 34.17 12.925 34.53 13.06 ;
        RECT 34.21 12.925 34.46 13.095 ;
        RECT 34.03 12.9 34.26 12.95 ;
        RECT 34.03 12.855 34.21 12.95 ;
        RECT 34.17 12.925 34.46 13.075 ;
        RECT 33.96 12.8 34.17 12.88 ;
        RECT 34.1 12.925 34.53 13.02 ;
        RECT 33.91 12.73 34.1 12.82 ;
        RECT 31.7 12.7 34.03 12.795 ;
        RECT 31.77 12.66 34.03 12.795 ;
        RECT 31.77 12.645 33.96 12.795 ;
        RECT 31.81 12.625 33.96 12.795 ;
        RECT 31.63 12.77 31.86 12.82 ;
        RECT 31.63 12.77 31.81 12.865 ;
        RECT 31.56 12.84 31.77 12.92 ;
        RECT 31.51 12.9 31.7 12.99 ;
        RECT 31.27 12.925 31.63 13.06 ;
        RECT 31.31 12.925 31.56 13.095 ;
        RECT 31.13 12.9 31.36 12.95 ;
        RECT 31.13 12.855 31.31 12.95 ;
        RECT 31.27 12.925 31.56 13.075 ;
        RECT 31.06 12.8 31.27 12.88 ;
        RECT 31.2 12.925 31.63 13.02 ;
        RECT 31.01 12.73 31.2 12.82 ;
        RECT 28.725 12.66 31.13 12.795 ;
        RECT 28.725 12.625 31.06 12.795 ;
        RECT 28.74 12.625 28.96 12.8 ;
        RECT 28.74 12.625 28.95 12.84 ;
        RECT 28.3 12.925 28.74 13.02 ;
        RECT 28.61 12.9 28.81 12.98 ;
        RECT 28.73 12.8 28.74 13.02 ;
        RECT 28.37 12.925 28.73 13.06 ;
        RECT 28.66 12.84 28.88 12.91 ;
        RECT 28.41 12.925 28.66 13.095 ;
        RECT 28.23 12.9 28.46 12.95 ;
        RECT 28.23 12.855 28.41 12.95 ;
        RECT 28.37 12.925 28.66 13.075 ;
        RECT 28.16 12.8 28.37 12.88 ;
        RECT 28.11 12.73 28.3 12.82 ;
        RECT 25.9 12.7 28.23 12.795 ;
        RECT 25.97 12.66 28.23 12.795 ;
        RECT 25.97 12.645 28.16 12.795 ;
        RECT 26.01 12.625 28.16 12.795 ;
        RECT 25.83 12.77 26.06 12.82 ;
        RECT 25.83 12.77 26.01 12.865 ;
        RECT 25.76 12.84 25.97 12.92 ;
        RECT 25.71 12.9 25.9 12.99 ;
        RECT 25.47 12.925 25.83 13.06 ;
        RECT 25.51 12.925 25.76 13.095 ;
        RECT 25.33 12.9 25.56 12.95 ;
        RECT 25.33 12.855 25.51 12.95 ;
        RECT 25.47 12.925 25.76 13.075 ;
        RECT 25.26 12.8 25.47 12.88 ;
        RECT 25.4 12.925 25.83 13.02 ;
        RECT 25.21 12.73 25.4 12.82 ;
        RECT 22.925 12.66 25.33 12.795 ;
        RECT 22.925 12.625 25.26 12.795 ;
        RECT 22.94 12.625 23.16 12.8 ;
        RECT 22.94 12.625 23.15 12.84 ;
        RECT 22.5 12.925 22.94 13.02 ;
        RECT 22.81 12.9 23.01 12.98 ;
        RECT 22.93 12.8 22.94 13.02 ;
        RECT 22.57 12.925 22.93 13.06 ;
        RECT 22.86 12.84 23.08 12.91 ;
        RECT 22.61 12.925 22.86 13.095 ;
        RECT 22.43 12.9 22.66 12.95 ;
        RECT 22.43 12.855 22.61 12.95 ;
        RECT 22.57 12.925 22.86 13.075 ;
        RECT 22.36 12.8 22.57 12.88 ;
        RECT 22.31 12.73 22.5 12.82 ;
        RECT 20.1 12.7 22.43 12.795 ;
        RECT 20.17 12.66 22.43 12.795 ;
        RECT 20.17 12.645 22.36 12.795 ;
        RECT 20.21 12.625 22.36 12.795 ;
        RECT 20.03 12.77 20.26 12.82 ;
        RECT 20.03 12.77 20.21 12.865 ;
        RECT 19.96 12.84 20.17 12.92 ;
        RECT 19.91 12.9 20.1 12.99 ;
        RECT 19.67 12.925 20.03 13.06 ;
        RECT 19.71 12.925 19.96 13.095 ;
        RECT 19.53 12.9 19.76 12.95 ;
        RECT 19.53 12.855 19.71 12.95 ;
        RECT 19.67 12.925 19.96 13.075 ;
        RECT 19.46 12.8 19.67 12.88 ;
        RECT 19.6 12.925 20.03 13.02 ;
        RECT 19.41 12.73 19.6 12.82 ;
        RECT 17.125 12.66 19.53 12.795 ;
        RECT 17.125 12.625 19.46 12.795 ;
        RECT 17.14 12.625 17.36 12.8 ;
        RECT 17.14 12.625 17.35 12.84 ;
        RECT 16.7 12.925 17.14 13.02 ;
        RECT 17.01 12.9 17.21 12.98 ;
        RECT 17.13 12.8 17.14 13.02 ;
        RECT 16.77 12.925 17.13 13.06 ;
        RECT 17.06 12.84 17.28 12.91 ;
        RECT 16.81 12.925 17.06 13.095 ;
        RECT 16.63 12.9 16.86 12.95 ;
        RECT 16.63 12.855 16.81 12.95 ;
        RECT 16.77 12.925 17.06 13.075 ;
        RECT 16.56 12.8 16.77 12.88 ;
        RECT 16.51 12.73 16.7 12.82 ;
        RECT 14.3 12.7 16.63 12.795 ;
        RECT 14.37 12.66 16.63 12.795 ;
        RECT 14.37 12.645 16.56 12.795 ;
        RECT 14.41 12.625 16.56 12.795 ;
        RECT 14.23 12.77 14.46 12.82 ;
        RECT 14.23 12.77 14.41 12.865 ;
        RECT 14.16 12.84 14.37 12.92 ;
        RECT 14.11 12.9 14.3 12.99 ;
        RECT 13.87 12.925 14.23 13.06 ;
        RECT 13.91 12.925 14.16 13.095 ;
        RECT 13.73 12.9 13.96 12.95 ;
        RECT 13.73 12.855 13.91 12.95 ;
        RECT 13.87 12.925 14.16 13.075 ;
        RECT 13.66 12.8 13.87 12.88 ;
        RECT 13.8 12.925 14.23 13.02 ;
        RECT 13.61 12.73 13.8 12.82 ;
        RECT 11.325 12.66 13.73 12.795 ;
        RECT 11.325 12.625 13.66 12.795 ;
        RECT 11.34 12.625 11.56 12.8 ;
        RECT 11.34 12.625 11.55 12.84 ;
        RECT 10.9 12.925 11.34 13.02 ;
        RECT 11.21 12.9 11.41 12.98 ;
        RECT 11.33 12.8 11.34 13.02 ;
        RECT 10.97 12.925 11.33 13.06 ;
        RECT 11.26 12.84 11.48 12.91 ;
        RECT 11.01 12.925 11.26 13.095 ;
        RECT 10.83 12.9 11.06 12.95 ;
        RECT 10.83 12.855 11.01 12.95 ;
        RECT 10.97 12.925 11.26 13.075 ;
        RECT 10.76 12.8 10.97 12.88 ;
        RECT 10.71 12.73 10.9 12.82 ;
        RECT 8.5 12.7 10.83 12.795 ;
        RECT 8.57 12.66 10.83 12.795 ;
        RECT 8.57 12.645 10.76 12.795 ;
        RECT 8.61 12.625 10.76 12.795 ;
        RECT 8.43 12.77 8.66 12.82 ;
        RECT 8.43 12.77 8.61 12.865 ;
        RECT 8.36 12.84 8.57 12.92 ;
        RECT 8.31 12.9 8.5 12.99 ;
        RECT 8.07 12.925 8.43 13.06 ;
        RECT 8.11 12.925 8.36 13.095 ;
        RECT 7.93 12.9 8.16 12.95 ;
        RECT 7.93 12.855 8.11 12.95 ;
        RECT 8.07 12.925 8.36 13.075 ;
        RECT 7.86 12.8 8.07 12.88 ;
        RECT 8 12.925 8.43 13.02 ;
        RECT 7.81 12.73 8 12.82 ;
        RECT 5.525 12.66 7.93 12.795 ;
        RECT 5.525 12.625 7.86 12.795 ;
        RECT 5.54 12.625 5.76 12.8 ;
        RECT 5.54 12.625 5.75 12.84 ;
        RECT 5.1 12.925 5.54 13.02 ;
        RECT 5.41 12.9 5.61 12.98 ;
        RECT 5.53 12.8 5.54 13.02 ;
        RECT 5.17 12.925 5.53 13.06 ;
        RECT 5.46 12.84 5.68 12.91 ;
        RECT 5.21 12.925 5.46 13.095 ;
        RECT 5.03 12.9 5.26 12.95 ;
        RECT 5.03 12.855 5.21 12.95 ;
        RECT 5.17 12.925 5.46 13.075 ;
        RECT 4.96 12.8 5.17 12.88 ;
        RECT 4.91 12.73 5.1 12.82 ;
        RECT 2.7 12.7 5.03 12.795 ;
        RECT 2.77 12.66 5.03 12.795 ;
        RECT 2.77 12.645 4.96 12.795 ;
        RECT 2.81 12.625 4.96 12.795 ;
        RECT 2.63 12.77 2.86 12.82 ;
        RECT 2.63 12.77 2.81 12.865 ;
        RECT 2.56 12.84 2.77 12.92 ;
        RECT 2.51 12.9 2.7 12.99 ;
        RECT 2.27 12.925 2.63 13.06 ;
        RECT 2.31 12.925 2.56 13.095 ;
        RECT 2.13 12.9 2.36 12.95 ;
        RECT 2.13 12.855 2.31 12.95 ;
        RECT 2.27 12.925 2.56 13.075 ;
        RECT 2.06 12.8 2.27 12.88 ;
        RECT 2.2 12.925 2.63 13.02 ;
        RECT 2.01 12.73 2.2 12.82 ;
        RECT -0.455 12.66 2.13 12.795 ;
        RECT -0.455 12.625 2.06 12.795 ;
    END
  END RWL1_9
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -0.455 1.095 34.625 1.165 ;
        RECT -0.455 2.445 34.625 2.515 ;
        RECT -0.455 3.795 34.625 3.865 ;
        RECT -0.455 5.145 34.625 5.215 ;
        RECT -0.455 6.495 34.625 6.565 ;
        RECT -0.455 7.845 34.625 7.915 ;
        RECT -0.455 9.195 34.625 9.265 ;
        RECT -0.455 10.545 34.625 10.615 ;
        RECT -0.455 11.895 34.625 11.965 ;
        RECT -0.455 13.245 34.625 13.315 ;
        RECT -0.455 14.595 34.625 14.665 ;
        RECT -0.455 15.945 34.625 16.015 ;
        RECT -0.455 17.295 34.625 17.365 ;
        RECT -0.455 18.645 34.625 18.715 ;
        RECT -0.455 19.995 34.625 20.065 ;
        RECT -0.455 21.345 34.625 21.415 ;
    END
  END VDD
  OBS
    LAYER met2 ;
      RECT -0.455 0.475 34.76 0.645 ;
      RECT -0.455 1.825 34.76 1.995 ;
      RECT -0.455 3.175 34.76 3.345 ;
      RECT -0.455 4.525 34.76 4.695 ;
      RECT -0.455 5.875 34.76 6.045 ;
      RECT -0.455 7.225 34.76 7.395 ;
      RECT -0.455 8.575 34.76 8.745 ;
      RECT -0.455 9.925 34.76 10.095 ;
      RECT -0.455 11.275 34.76 11.445 ;
      RECT -0.455 12.625 34.76 12.795 ;
      RECT -0.455 13.975 34.76 14.145 ;
      RECT -0.455 15.325 34.76 15.495 ;
      RECT -0.455 16.675 34.76 16.845 ;
      RECT -0.455 18.025 34.76 18.195 ;
      RECT -0.455 19.375 34.76 19.545 ;
      RECT -0.455 20.725 34.76 20.895 ;
    LAYER met1 ;
      RECT 34.26 0.475 34.41 0.645 ;
      RECT 34.26 1.825 34.41 1.995 ;
      RECT 34.26 3.175 34.41 3.345 ;
      RECT 34.26 4.525 34.41 4.695 ;
      RECT 34.26 5.875 34.41 6.045 ;
      RECT 34.26 7.225 34.41 7.395 ;
      RECT 34.26 8.575 34.41 8.745 ;
      RECT 34.26 9.925 34.41 10.095 ;
      RECT 34.26 11.275 34.41 11.445 ;
      RECT 34.26 12.625 34.41 12.795 ;
      RECT 34.26 13.975 34.41 14.145 ;
      RECT 34.26 15.325 34.41 15.495 ;
      RECT 34.26 16.675 34.41 16.845 ;
      RECT 34.26 18.025 34.41 18.195 ;
      RECT 34.26 19.375 34.41 19.545 ;
      RECT 34.26 20.725 34.41 20.895 ;
      RECT 31.36 0.475 31.51 0.645 ;
      RECT 31.36 1.825 31.51 1.995 ;
      RECT 31.36 3.175 31.51 3.345 ;
      RECT 31.36 4.525 31.51 4.695 ;
      RECT 31.36 5.875 31.51 6.045 ;
      RECT 31.36 7.225 31.51 7.395 ;
      RECT 31.36 8.575 31.51 8.745 ;
      RECT 31.36 9.925 31.51 10.095 ;
      RECT 31.36 11.275 31.51 11.445 ;
      RECT 31.36 12.625 31.51 12.795 ;
      RECT 31.36 13.975 31.51 14.145 ;
      RECT 31.36 15.325 31.51 15.495 ;
      RECT 31.36 16.675 31.51 16.845 ;
      RECT 31.36 18.025 31.51 18.195 ;
      RECT 31.36 19.375 31.51 19.545 ;
      RECT 31.36 20.725 31.51 20.895 ;
      RECT 28.46 0.475 28.61 0.645 ;
      RECT 28.46 1.825 28.61 1.995 ;
      RECT 28.46 3.175 28.61 3.345 ;
      RECT 28.46 4.525 28.61 4.695 ;
      RECT 28.46 5.875 28.61 6.045 ;
      RECT 28.46 7.225 28.61 7.395 ;
      RECT 28.46 8.575 28.61 8.745 ;
      RECT 28.46 9.925 28.61 10.095 ;
      RECT 28.46 11.275 28.61 11.445 ;
      RECT 28.46 12.625 28.61 12.795 ;
      RECT 28.46 13.975 28.61 14.145 ;
      RECT 28.46 15.325 28.61 15.495 ;
      RECT 28.46 16.675 28.61 16.845 ;
      RECT 28.46 18.025 28.61 18.195 ;
      RECT 28.46 19.375 28.61 19.545 ;
      RECT 28.46 20.725 28.61 20.895 ;
      RECT 25.56 0.475 25.71 0.645 ;
      RECT 25.56 1.825 25.71 1.995 ;
      RECT 25.56 3.175 25.71 3.345 ;
      RECT 25.56 4.525 25.71 4.695 ;
      RECT 25.56 5.875 25.71 6.045 ;
      RECT 25.56 7.225 25.71 7.395 ;
      RECT 25.56 8.575 25.71 8.745 ;
      RECT 25.56 9.925 25.71 10.095 ;
      RECT 25.56 11.275 25.71 11.445 ;
      RECT 25.56 12.625 25.71 12.795 ;
      RECT 25.56 13.975 25.71 14.145 ;
      RECT 25.56 15.325 25.71 15.495 ;
      RECT 25.56 16.675 25.71 16.845 ;
      RECT 25.56 18.025 25.71 18.195 ;
      RECT 25.56 19.375 25.71 19.545 ;
      RECT 25.56 20.725 25.71 20.895 ;
      RECT 22.66 0.475 22.81 0.645 ;
      RECT 22.66 1.825 22.81 1.995 ;
      RECT 22.66 3.175 22.81 3.345 ;
      RECT 22.66 4.525 22.81 4.695 ;
      RECT 22.66 5.875 22.81 6.045 ;
      RECT 22.66 7.225 22.81 7.395 ;
      RECT 22.66 8.575 22.81 8.745 ;
      RECT 22.66 9.925 22.81 10.095 ;
      RECT 22.66 11.275 22.81 11.445 ;
      RECT 22.66 12.625 22.81 12.795 ;
      RECT 22.66 13.975 22.81 14.145 ;
      RECT 22.66 15.325 22.81 15.495 ;
      RECT 22.66 16.675 22.81 16.845 ;
      RECT 22.66 18.025 22.81 18.195 ;
      RECT 22.66 19.375 22.81 19.545 ;
      RECT 22.66 20.725 22.81 20.895 ;
      RECT 19.76 0.475 19.91 0.645 ;
      RECT 19.76 1.825 19.91 1.995 ;
      RECT 19.76 3.175 19.91 3.345 ;
      RECT 19.76 4.525 19.91 4.695 ;
      RECT 19.76 5.875 19.91 6.045 ;
      RECT 19.76 7.225 19.91 7.395 ;
      RECT 19.76 8.575 19.91 8.745 ;
      RECT 19.76 9.925 19.91 10.095 ;
      RECT 19.76 11.275 19.91 11.445 ;
      RECT 19.76 12.625 19.91 12.795 ;
      RECT 19.76 13.975 19.91 14.145 ;
      RECT 19.76 15.325 19.91 15.495 ;
      RECT 19.76 16.675 19.91 16.845 ;
      RECT 19.76 18.025 19.91 18.195 ;
      RECT 19.76 19.375 19.91 19.545 ;
      RECT 19.76 20.725 19.91 20.895 ;
      RECT 16.86 0.475 17.01 0.645 ;
      RECT 16.86 1.825 17.01 1.995 ;
      RECT 16.86 3.175 17.01 3.345 ;
      RECT 16.86 4.525 17.01 4.695 ;
      RECT 16.86 5.875 17.01 6.045 ;
      RECT 16.86 7.225 17.01 7.395 ;
      RECT 16.86 8.575 17.01 8.745 ;
      RECT 16.86 9.925 17.01 10.095 ;
      RECT 16.86 11.275 17.01 11.445 ;
      RECT 16.86 12.625 17.01 12.795 ;
      RECT 16.86 13.975 17.01 14.145 ;
      RECT 16.86 15.325 17.01 15.495 ;
      RECT 16.86 16.675 17.01 16.845 ;
      RECT 16.86 18.025 17.01 18.195 ;
      RECT 16.86 19.375 17.01 19.545 ;
      RECT 16.86 20.725 17.01 20.895 ;
      RECT 13.96 0.475 14.11 0.645 ;
      RECT 13.96 1.825 14.11 1.995 ;
      RECT 13.96 3.175 14.11 3.345 ;
      RECT 13.96 4.525 14.11 4.695 ;
      RECT 13.96 5.875 14.11 6.045 ;
      RECT 13.96 7.225 14.11 7.395 ;
      RECT 13.96 8.575 14.11 8.745 ;
      RECT 13.96 9.925 14.11 10.095 ;
      RECT 13.96 11.275 14.11 11.445 ;
      RECT 13.96 12.625 14.11 12.795 ;
      RECT 13.96 13.975 14.11 14.145 ;
      RECT 13.96 15.325 14.11 15.495 ;
      RECT 13.96 16.675 14.11 16.845 ;
      RECT 13.96 18.025 14.11 18.195 ;
      RECT 13.96 19.375 14.11 19.545 ;
      RECT 13.96 20.725 14.11 20.895 ;
      RECT 11.06 0.475 11.21 0.645 ;
      RECT 11.06 1.825 11.21 1.995 ;
      RECT 11.06 3.175 11.21 3.345 ;
      RECT 11.06 4.525 11.21 4.695 ;
      RECT 11.06 5.875 11.21 6.045 ;
      RECT 11.06 7.225 11.21 7.395 ;
      RECT 11.06 8.575 11.21 8.745 ;
      RECT 11.06 9.925 11.21 10.095 ;
      RECT 11.06 11.275 11.21 11.445 ;
      RECT 11.06 12.625 11.21 12.795 ;
      RECT 11.06 13.975 11.21 14.145 ;
      RECT 11.06 15.325 11.21 15.495 ;
      RECT 11.06 16.675 11.21 16.845 ;
      RECT 11.06 18.025 11.21 18.195 ;
      RECT 11.06 19.375 11.21 19.545 ;
      RECT 11.06 20.725 11.21 20.895 ;
      RECT 8.16 0.475 8.31 0.645 ;
      RECT 8.16 1.825 8.31 1.995 ;
      RECT 8.16 3.175 8.31 3.345 ;
      RECT 8.16 4.525 8.31 4.695 ;
      RECT 8.16 5.875 8.31 6.045 ;
      RECT 8.16 7.225 8.31 7.395 ;
      RECT 8.16 8.575 8.31 8.745 ;
      RECT 8.16 9.925 8.31 10.095 ;
      RECT 8.16 11.275 8.31 11.445 ;
      RECT 8.16 12.625 8.31 12.795 ;
      RECT 8.16 13.975 8.31 14.145 ;
      RECT 8.16 15.325 8.31 15.495 ;
      RECT 8.16 16.675 8.31 16.845 ;
      RECT 8.16 18.025 8.31 18.195 ;
      RECT 8.16 19.375 8.31 19.545 ;
      RECT 8.16 20.725 8.31 20.895 ;
      RECT 5.26 0.475 5.41 0.645 ;
      RECT 5.26 1.825 5.41 1.995 ;
      RECT 5.26 3.175 5.41 3.345 ;
      RECT 5.26 4.525 5.41 4.695 ;
      RECT 5.26 5.875 5.41 6.045 ;
      RECT 5.26 7.225 5.41 7.395 ;
      RECT 5.26 8.575 5.41 8.745 ;
      RECT 5.26 9.925 5.41 10.095 ;
      RECT 5.26 11.275 5.41 11.445 ;
      RECT 5.26 12.625 5.41 12.795 ;
      RECT 5.26 13.975 5.41 14.145 ;
      RECT 5.26 15.325 5.41 15.495 ;
      RECT 5.26 16.675 5.41 16.845 ;
      RECT 5.26 18.025 5.41 18.195 ;
      RECT 5.26 19.375 5.41 19.545 ;
      RECT 5.26 20.725 5.41 20.895 ;
      RECT 2.36 0.475 2.51 0.645 ;
      RECT 2.36 1.825 2.51 1.995 ;
      RECT 2.36 3.175 2.51 3.345 ;
      RECT 2.36 4.525 2.51 4.695 ;
      RECT 2.36 5.875 2.51 6.045 ;
      RECT 2.36 7.225 2.51 7.395 ;
      RECT 2.36 8.575 2.51 8.745 ;
      RECT 2.36 9.925 2.51 10.095 ;
      RECT 2.36 11.275 2.51 11.445 ;
      RECT 2.36 12.625 2.51 12.795 ;
      RECT 2.36 13.975 2.51 14.145 ;
      RECT 2.36 15.325 2.51 15.495 ;
      RECT 2.36 16.675 2.51 16.845 ;
      RECT 2.36 18.025 2.51 18.195 ;
      RECT 2.36 19.375 2.51 19.545 ;
      RECT 2.36 20.725 2.51 20.895 ;
  END
END 10T_16x12_2r1w_magic_flattened

END LIBRARY
