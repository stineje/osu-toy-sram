magic
tech sky130A
magscale 1 2
timestamp 1655151742
<< error_s >>
rect -15 258 -2 274
rect 86 272 99 274
rect 52 258 67 272
rect 83 258 113 272
rect 174 270 327 316
rect 156 258 348 270
rect 391 258 421 272
rect 433 258 446 274
rect 534 258 547 274
rect 583 258 596 274
rect 684 272 697 274
rect 650 258 665 272
rect 681 258 711 272
rect 772 270 925 316
rect 754 258 946 270
rect 989 258 1019 272
rect 1031 258 1044 274
rect 1132 258 1145 274
rect -30 244 1145 258
rect -15 140 -2 244
rect 42 222 43 232
rect 58 222 71 232
rect 42 218 71 222
rect 83 218 113 244
rect 131 230 147 232
rect 219 230 285 244
rect 220 228 284 230
rect 327 228 342 244
rect 391 241 421 244
rect 391 238 433 241
rect 357 230 373 232
rect 131 218 146 222
rect 42 216 146 218
rect 174 216 342 228
rect 358 218 373 222
rect 391 219 436 238
rect 455 232 462 233
rect 461 225 462 232
rect 445 222 446 225
rect 461 222 474 225
rect 391 218 421 219
rect 436 218 442 219
rect 445 218 474 222
rect 358 217 474 218
rect 358 216 480 217
rect 33 208 77 216
rect 33 196 51 208
rect 58 196 77 208
rect 115 208 165 216
rect 115 200 131 208
rect 138 206 165 208
rect 174 206 395 216
rect 138 196 395 206
rect 430 208 480 216
rect 430 201 446 208
rect 33 188 77 196
rect 131 188 395 196
rect 445 196 446 201
rect 453 196 480 208
rect 445 188 480 196
rect 42 172 43 188
rect 58 168 71 188
rect 43 156 71 168
rect 13 140 71 156
rect -15 126 61 140
rect 63 132 71 140
rect 83 132 113 188
rect 148 178 356 188
rect 174 148 363 178
rect 189 145 363 148
rect 182 142 363 145
rect 391 164 421 188
rect 427 167 442 179
rect 445 172 446 188
rect 461 168 474 188
rect 446 167 474 168
rect 427 164 461 167
rect 391 151 427 164
rect 433 156 461 164
rect -15 124 59 126
rect -15 122 -2 124
rect 13 122 47 124
rect -15 106 59 122
rect 61 120 67 126
rect 86 118 99 132
rect 114 118 131 134
rect 182 129 193 142
rect -31 84 -30 100
rect -15 84 -2 106
rect 13 84 43 106
rect 86 102 148 118
rect 182 111 193 127
rect 198 122 208 142
rect 218 122 232 142
rect 235 129 244 142
rect 260 129 269 142
rect 198 111 232 122
rect 235 111 244 127
rect 260 111 269 127
rect 276 122 286 142
rect 296 122 310 142
rect 311 129 322 142
rect 276 111 310 122
rect 311 111 322 127
rect 373 126 390 142
rect 391 132 421 151
rect 433 145 491 156
rect 433 140 446 145
rect 461 140 491 145
rect 360 116 406 126
rect 360 108 370 116
rect 389 110 406 116
rect 433 124 507 140
rect 433 122 446 124
rect 461 122 495 124
rect 389 108 394 110
rect 86 100 99 102
rect 114 100 148 102
rect 86 84 151 100
rect 198 96 199 102
rect 198 95 214 96
rect 276 95 306 106
rect 360 92 406 108
rect 433 106 507 122
rect 373 84 390 92
rect 433 84 446 106
rect 461 84 491 106
rect 518 84 519 100
rect 534 84 547 244
rect 583 140 596 244
rect 640 222 641 232
rect 656 222 669 232
rect 640 218 669 222
rect 681 218 711 244
rect 729 230 745 232
rect 817 230 883 244
rect 818 228 882 230
rect 925 228 940 244
rect 989 241 1019 244
rect 989 238 1031 241
rect 955 230 971 232
rect 729 218 744 222
rect 640 216 744 218
rect 772 216 940 228
rect 956 218 971 222
rect 989 219 1034 238
rect 1053 232 1060 233
rect 1059 225 1060 232
rect 1043 222 1044 225
rect 1059 222 1072 225
rect 989 218 1019 219
rect 1034 218 1040 219
rect 1043 218 1072 222
rect 956 217 1072 218
rect 956 216 1078 217
rect 631 208 675 216
rect 631 196 649 208
rect 656 196 675 208
rect 713 208 763 216
rect 713 200 729 208
rect 736 206 763 208
rect 772 206 993 216
rect 736 196 993 206
rect 1028 208 1078 216
rect 1028 201 1044 208
rect 631 188 675 196
rect 729 188 993 196
rect 1043 196 1044 201
rect 1051 196 1078 208
rect 1043 188 1078 196
rect 640 172 641 188
rect 656 168 669 188
rect 641 156 669 168
rect 611 140 669 156
rect 583 126 659 140
rect 661 132 669 140
rect 681 132 711 188
rect 746 178 954 188
rect 772 148 961 178
rect 787 145 961 148
rect 780 142 961 145
rect 989 164 1019 188
rect 1025 167 1040 179
rect 1043 172 1044 188
rect 1059 168 1072 188
rect 1044 167 1072 168
rect 1025 164 1059 167
rect 989 151 1025 164
rect 1031 156 1059 164
rect 583 124 657 126
rect 583 122 596 124
rect 611 122 645 124
rect 583 106 657 122
rect 659 120 665 126
rect 684 118 697 132
rect 712 118 729 134
rect 780 129 791 142
rect 567 84 568 100
rect 583 84 596 106
rect 611 84 641 106
rect 684 102 746 118
rect 780 111 791 127
rect 796 122 806 142
rect 816 122 830 142
rect 833 129 842 142
rect 858 129 867 142
rect 796 111 830 122
rect 833 111 842 127
rect 858 111 867 127
rect 874 122 884 142
rect 894 122 908 142
rect 909 129 920 142
rect 874 111 908 122
rect 909 111 920 127
rect 971 126 988 142
rect 989 132 1019 151
rect 1031 145 1089 156
rect 1031 140 1044 145
rect 1059 140 1089 145
rect 958 116 1004 126
rect 958 108 968 116
rect 987 110 1004 116
rect 1031 124 1105 140
rect 1031 122 1044 124
rect 1059 122 1093 124
rect 987 108 992 110
rect 684 100 697 102
rect 712 100 746 102
rect 684 84 749 100
rect 796 96 797 102
rect 796 95 812 96
rect 874 95 904 106
rect 958 92 1004 108
rect 1031 106 1105 122
rect 971 84 988 92
rect 1031 84 1044 106
rect 1059 84 1089 106
rect 1116 84 1117 100
rect 1132 84 1145 244
rect -37 76 4 84
rect -37 50 -22 76
rect -15 50 4 76
rect 66 72 99 84
rect 105 72 135 84
rect 148 72 223 84
rect 281 72 356 84
rect 369 72 399 84
rect 411 72 446 84
rect 66 70 236 72
rect -37 42 4 50
rect -31 32 -30 42
rect -15 32 -2 42
rect 13 32 43 46
rect 86 32 99 70
rect 114 68 131 70
rect 105 32 135 46
rect 156 42 166 51
rect 169 46 236 70
rect 268 70 446 72
rect 268 46 348 70
rect 169 42 348 46
rect 142 32 172 42
rect 174 32 327 42
rect 335 32 365 42
rect 369 32 399 46
rect 433 32 446 70
rect 518 76 553 84
rect 518 50 519 76
rect 526 50 553 76
rect 461 32 491 46
rect 518 42 553 50
rect 561 76 602 84
rect 561 50 576 76
rect 583 50 602 76
rect 664 72 697 84
rect 703 72 733 84
rect 746 72 821 84
rect 879 72 954 84
rect 967 72 997 84
rect 1009 72 1044 84
rect 664 70 834 72
rect 561 42 602 50
rect 518 32 519 42
rect 534 32 547 42
rect 567 32 568 42
rect 583 32 596 42
rect 611 32 641 46
rect 684 32 697 70
rect 712 68 729 70
rect 703 32 733 46
rect 754 42 764 51
rect 767 46 834 70
rect 866 70 1044 72
rect 866 46 946 70
rect 767 42 946 46
rect 740 32 770 42
rect 772 32 925 42
rect 933 32 963 42
rect 967 32 997 46
rect 1031 32 1044 70
rect 1116 76 1151 84
rect 1116 50 1117 76
rect 1124 50 1151 76
rect 1059 32 1089 46
rect 1116 42 1151 50
rect 1116 32 1117 42
rect 1132 32 1145 42
rect -31 26 1145 32
rect -30 18 1145 26
rect -15 -12 -2 18
rect 13 0 43 18
rect 86 2 99 18
rect 142 4 362 18
rect 52 -12 67 2
rect 83 -12 113 2
rect 174 0 327 4
rect 156 -12 348 0
rect 391 -12 421 2
rect 433 -12 446 18
rect 461 0 491 18
rect 534 -12 547 18
rect 583 -12 596 18
rect 611 0 641 18
rect 684 2 697 18
rect 740 4 960 18
rect 650 -12 665 2
rect 681 -12 711 2
rect 772 0 925 4
rect 754 -12 946 0
rect 989 -12 1019 2
rect 1031 -12 1044 18
rect 1059 0 1089 18
rect 1132 -12 1145 18
rect -30 -26 1145 -12
rect -15 -130 -2 -26
rect 42 -48 43 -38
rect 58 -48 71 -38
rect 42 -52 71 -48
rect 83 -52 113 -26
rect 131 -40 147 -38
rect 219 -40 285 -26
rect 220 -42 284 -40
rect 131 -52 146 -48
rect 42 -54 146 -52
rect 33 -62 77 -54
rect 33 -74 51 -62
rect 58 -74 77 -62
rect 115 -62 165 -54
rect 115 -70 131 -62
rect 138 -64 165 -62
rect 174 -62 189 -58
rect 236 -62 268 -42
rect 327 -54 342 -26
rect 391 -29 421 -26
rect 391 -32 433 -29
rect 357 -40 373 -38
rect 358 -52 373 -48
rect 391 -51 436 -32
rect 455 -38 462 -37
rect 461 -45 462 -38
rect 445 -48 446 -45
rect 461 -48 474 -45
rect 391 -52 421 -51
rect 436 -52 442 -51
rect 445 -52 474 -48
rect 358 -53 474 -52
rect 358 -54 480 -53
rect 327 -62 395 -54
rect 174 -64 395 -62
rect 138 -74 210 -64
rect 228 -65 236 -64
rect 268 -65 276 -64
rect 33 -82 77 -74
rect 131 -78 210 -74
rect 291 -78 395 -64
rect 430 -62 480 -54
rect 430 -69 446 -62
rect 131 -82 395 -78
rect 445 -74 446 -69
rect 453 -74 480 -62
rect 445 -82 480 -74
rect 42 -98 43 -82
rect 58 -102 71 -82
rect 43 -114 71 -102
rect 13 -130 71 -114
rect -15 -144 61 -130
rect 63 -138 71 -130
rect 83 -138 113 -82
rect 148 -92 356 -82
rect 315 -96 363 -92
rect 198 -118 228 -109
rect 291 -116 306 -109
rect 327 -118 363 -96
rect 174 -122 363 -118
rect 189 -125 363 -122
rect 182 -128 363 -125
rect 391 -106 421 -82
rect 427 -103 442 -91
rect 445 -98 446 -82
rect 461 -102 474 -82
rect 446 -103 474 -102
rect 427 -106 461 -103
rect 391 -119 427 -106
rect 433 -114 461 -106
rect -15 -146 59 -144
rect -15 -148 -2 -146
rect 13 -148 47 -146
rect -15 -164 59 -148
rect 61 -150 67 -144
rect 86 -152 99 -138
rect 114 -152 131 -136
rect 182 -141 193 -128
rect -31 -186 -30 -170
rect -15 -186 -2 -164
rect 13 -186 43 -164
rect 86 -168 148 -152
rect 182 -159 193 -143
rect 198 -148 208 -128
rect 218 -148 232 -128
rect 235 -141 244 -128
rect 260 -141 269 -128
rect 198 -159 232 -148
rect 235 -159 244 -143
rect 260 -159 269 -143
rect 276 -148 286 -128
rect 296 -148 310 -128
rect 311 -141 322 -128
rect 276 -159 310 -148
rect 311 -159 322 -143
rect 373 -144 390 -128
rect 391 -138 421 -119
rect 433 -125 491 -114
rect 433 -130 446 -125
rect 461 -130 491 -125
rect 360 -154 406 -144
rect 360 -162 370 -154
rect 389 -160 406 -154
rect 433 -146 507 -130
rect 433 -148 446 -146
rect 461 -148 495 -146
rect 389 -162 394 -160
rect 86 -170 99 -168
rect 114 -170 148 -168
rect 86 -186 151 -170
rect 198 -174 199 -168
rect 198 -175 214 -174
rect 276 -175 306 -164
rect 360 -178 406 -162
rect 433 -164 507 -148
rect 373 -186 390 -178
rect 433 -186 446 -164
rect 461 -186 491 -164
rect 518 -186 519 -170
rect 534 -186 547 -26
rect 583 -130 596 -26
rect 640 -48 641 -38
rect 656 -48 669 -38
rect 640 -52 669 -48
rect 681 -52 711 -26
rect 729 -40 745 -38
rect 817 -40 883 -26
rect 818 -42 882 -40
rect 729 -52 744 -48
rect 640 -54 744 -52
rect 631 -62 675 -54
rect 631 -74 649 -62
rect 656 -74 675 -62
rect 713 -62 763 -54
rect 713 -70 729 -62
rect 736 -64 763 -62
rect 772 -62 787 -58
rect 834 -62 866 -42
rect 925 -54 940 -26
rect 989 -29 1019 -26
rect 989 -32 1031 -29
rect 955 -40 971 -38
rect 956 -52 971 -48
rect 989 -51 1034 -32
rect 1053 -38 1060 -37
rect 1059 -45 1060 -38
rect 1043 -48 1044 -45
rect 1059 -48 1072 -45
rect 989 -52 1019 -51
rect 1034 -52 1040 -51
rect 1043 -52 1072 -48
rect 956 -53 1072 -52
rect 956 -54 1078 -53
rect 925 -62 993 -54
rect 772 -64 993 -62
rect 736 -74 808 -64
rect 826 -65 834 -64
rect 866 -65 874 -64
rect 631 -82 675 -74
rect 729 -78 808 -74
rect 889 -78 993 -64
rect 1028 -62 1078 -54
rect 1028 -69 1044 -62
rect 729 -82 993 -78
rect 1043 -74 1044 -69
rect 1051 -74 1078 -62
rect 1043 -82 1078 -74
rect 640 -98 641 -82
rect 656 -102 669 -82
rect 641 -114 669 -102
rect 611 -130 669 -114
rect 583 -144 659 -130
rect 661 -138 669 -130
rect 681 -138 711 -82
rect 746 -92 954 -82
rect 913 -96 961 -92
rect 796 -118 826 -109
rect 889 -116 904 -109
rect 925 -118 961 -96
rect 772 -122 961 -118
rect 787 -125 961 -122
rect 780 -128 961 -125
rect 989 -106 1019 -82
rect 1025 -103 1040 -91
rect 1043 -98 1044 -82
rect 1059 -102 1072 -82
rect 1044 -103 1072 -102
rect 1025 -106 1059 -103
rect 989 -119 1025 -106
rect 1031 -114 1059 -106
rect 583 -146 657 -144
rect 583 -148 596 -146
rect 611 -148 645 -146
rect 583 -164 657 -148
rect 659 -150 665 -144
rect 684 -152 697 -138
rect 712 -152 729 -136
rect 780 -141 791 -128
rect 567 -186 568 -170
rect 583 -186 596 -164
rect 611 -186 641 -164
rect 684 -168 746 -152
rect 780 -159 791 -143
rect 796 -148 806 -128
rect 816 -148 830 -128
rect 833 -141 842 -128
rect 858 -141 867 -128
rect 796 -159 830 -148
rect 833 -159 842 -143
rect 858 -159 867 -143
rect 874 -148 884 -128
rect 894 -148 908 -128
rect 909 -141 920 -128
rect 874 -159 908 -148
rect 909 -159 920 -143
rect 971 -144 988 -128
rect 989 -138 1019 -119
rect 1031 -125 1089 -114
rect 1031 -130 1044 -125
rect 1059 -130 1089 -125
rect 958 -154 1004 -144
rect 958 -162 968 -154
rect 987 -160 1004 -154
rect 1031 -146 1105 -130
rect 1031 -148 1044 -146
rect 1059 -148 1093 -146
rect 987 -162 992 -160
rect 684 -170 697 -168
rect 712 -170 746 -168
rect 684 -186 749 -170
rect 796 -174 797 -168
rect 796 -175 812 -174
rect 874 -175 904 -164
rect 958 -178 1004 -162
rect 1031 -164 1105 -148
rect 971 -186 988 -178
rect 1031 -186 1044 -164
rect 1059 -186 1089 -164
rect 1116 -186 1117 -170
rect 1132 -186 1145 -26
rect -37 -194 4 -186
rect -37 -220 -22 -194
rect -15 -220 4 -194
rect 66 -198 99 -186
rect 105 -198 135 -186
rect 148 -198 223 -186
rect 281 -198 356 -186
rect 369 -198 399 -186
rect 411 -198 446 -186
rect 66 -200 236 -198
rect -37 -228 4 -220
rect -31 -238 -30 -228
rect -15 -238 -2 -228
rect 13 -238 43 -228
rect 86 -238 99 -200
rect 114 -202 131 -200
rect 105 -238 135 -228
rect 142 -238 150 -228
rect 156 -229 166 -219
rect 169 -227 236 -200
rect 268 -200 446 -198
rect 268 -227 348 -200
rect 169 -228 348 -227
rect 169 -236 172 -228
rect 236 -236 268 -228
rect 169 -238 335 -236
rect 354 -238 365 -228
rect 369 -238 399 -228
rect 433 -238 446 -200
rect 518 -194 553 -186
rect 518 -220 519 -194
rect 526 -220 553 -194
rect 518 -228 553 -220
rect 561 -194 602 -186
rect 561 -220 576 -194
rect 583 -220 602 -194
rect 664 -198 697 -186
rect 703 -198 733 -186
rect 746 -198 821 -186
rect 879 -198 954 -186
rect 967 -198 997 -186
rect 1009 -198 1044 -186
rect 664 -200 834 -198
rect 561 -228 602 -220
rect 461 -238 491 -228
rect 518 -238 519 -228
rect 534 -238 547 -228
rect 567 -238 568 -228
rect 583 -238 596 -228
rect 611 -238 641 -228
rect 684 -238 697 -200
rect 712 -202 729 -200
rect 703 -238 733 -228
rect 740 -238 748 -228
rect 754 -229 764 -219
rect 767 -227 834 -200
rect 866 -200 1044 -198
rect 866 -227 946 -200
rect 767 -228 946 -227
rect 767 -236 770 -228
rect 834 -236 866 -228
rect 767 -238 933 -236
rect 952 -238 963 -228
rect 967 -238 997 -228
rect 1031 -238 1044 -200
rect 1116 -194 1151 -186
rect 1116 -220 1117 -194
rect 1124 -220 1151 -194
rect 1116 -228 1151 -220
rect 1059 -238 1089 -228
rect 1116 -238 1117 -228
rect 1132 -238 1145 -228
rect -31 -244 1145 -238
rect -30 -252 1145 -244
rect -15 -266 -2 -252
rect 13 -270 43 -252
rect 86 -266 99 -252
rect 142 -265 150 -252
rect 183 -261 321 -252
rect 183 -265 276 -261
rect 205 -266 276 -265
rect 285 -265 321 -261
rect 354 -265 362 -252
rect 285 -266 299 -265
rect 433 -266 446 -252
rect 220 -268 284 -266
rect 228 -274 236 -268
rect 268 -274 276 -268
rect 461 -270 491 -252
rect 534 -266 547 -252
rect 583 -266 596 -252
rect 611 -270 641 -252
rect 684 -266 697 -252
rect 740 -265 748 -252
rect 781 -261 919 -252
rect 781 -265 874 -261
rect 803 -266 874 -265
rect 883 -265 919 -261
rect 952 -265 960 -252
rect 883 -266 897 -265
rect 1031 -266 1044 -252
rect 818 -268 882 -266
rect 826 -274 834 -268
rect 866 -274 874 -268
rect 1059 -270 1089 -252
rect 1132 -266 1145 -252
<< poly >>
rect 534 244 568 274
rect 534 -26 568 4
<< metal1 >>
rect 537 230 568 244
rect 537 4 568 18
rect 537 -40 568 -26
rect 537 -266 568 -252
use 10T_toy_magic  10T_toy_magic_1
timestamp 1655151675
transform 1 0 674 0 1 23
box -113 -27 477 293
use 10T_toy_magic  10T_toy_magic_3
timestamp 1655151675
transform 1 0 674 0 1 -247
box -113 -27 477 293
use 10T_toy_magic  10T_toy_magic_0
timestamp 1655151675
transform 1 0 76 0 1 23
box -113 -27 477 293
use 10T_toy_magic  10T_toy_magic_2
timestamp 1655151675
transform 1 0 76 0 1 -247
box -113 -27 477 293
<< end >>
