magic
tech sky130A
magscale 1 2
timestamp 1656030011
<< error_s >>
rect 15 8624 28 8640
rect 117 8638 130 8640
rect 83 8624 98 8638
rect 107 8624 137 8638
rect 198 8636 351 8682
rect 180 8624 372 8636
rect 415 8624 445 8638
rect 451 8624 464 8640
rect 552 8624 565 8640
rect 595 8624 608 8640
rect 697 8638 710 8640
rect 663 8624 678 8638
rect 687 8624 717 8638
rect 778 8636 931 8682
rect 760 8624 952 8636
rect 995 8624 1025 8638
rect 1031 8624 1044 8640
rect 1132 8624 1145 8640
rect 1175 8624 1188 8640
rect 1277 8638 1290 8640
rect 1243 8624 1258 8638
rect 1267 8624 1297 8638
rect 1358 8636 1511 8682
rect 1340 8624 1532 8636
rect 1575 8624 1605 8638
rect 1611 8624 1624 8640
rect 1712 8624 1725 8640
rect 1755 8624 1768 8640
rect 1857 8638 1870 8640
rect 1823 8624 1838 8638
rect 1847 8624 1877 8638
rect 1938 8636 2091 8682
rect 1920 8624 2112 8636
rect 2155 8624 2185 8638
rect 2191 8624 2204 8640
rect 2292 8624 2305 8640
rect 2335 8624 2348 8640
rect 2437 8638 2450 8640
rect 2403 8624 2418 8638
rect 2427 8624 2457 8638
rect 2518 8636 2671 8682
rect 2500 8624 2692 8636
rect 2735 8624 2765 8638
rect 2771 8624 2784 8640
rect 2872 8624 2885 8640
rect 2915 8624 2928 8640
rect 3017 8638 3030 8640
rect 2983 8624 2998 8638
rect 3007 8624 3037 8638
rect 3098 8636 3251 8682
rect 3080 8624 3272 8636
rect 3315 8624 3345 8638
rect 3351 8624 3364 8640
rect 3452 8624 3465 8640
rect 3495 8624 3508 8640
rect 3597 8638 3610 8640
rect 3563 8624 3578 8638
rect 3587 8624 3617 8638
rect 3678 8636 3831 8682
rect 3660 8624 3852 8636
rect 3895 8624 3925 8638
rect 3931 8624 3944 8640
rect 4032 8624 4045 8640
rect 4075 8624 4088 8640
rect 4177 8638 4190 8640
rect 4143 8624 4158 8638
rect 4167 8624 4197 8638
rect 4258 8636 4411 8682
rect 4240 8624 4432 8636
rect 4475 8624 4505 8638
rect 4511 8624 4524 8640
rect 4612 8624 4625 8640
rect 4655 8624 4668 8640
rect 4757 8638 4770 8640
rect 4723 8624 4738 8638
rect 4747 8624 4777 8638
rect 4838 8636 4991 8682
rect 4820 8624 5012 8636
rect 5055 8624 5085 8638
rect 5091 8624 5104 8640
rect 5192 8624 5205 8640
rect 5235 8624 5248 8640
rect 5337 8638 5350 8640
rect 5303 8624 5318 8638
rect 5327 8624 5357 8638
rect 5418 8636 5571 8682
rect 5400 8624 5592 8636
rect 5635 8624 5665 8638
rect 5671 8624 5684 8640
rect 5772 8624 5785 8640
rect 5815 8624 5828 8640
rect 5917 8638 5930 8640
rect 5883 8624 5898 8638
rect 5907 8624 5937 8638
rect 5998 8636 6151 8682
rect 5980 8624 6172 8636
rect 6215 8624 6245 8638
rect 6251 8624 6264 8640
rect 6352 8624 6365 8640
rect 6395 8624 6408 8640
rect 6497 8638 6510 8640
rect 6463 8624 6478 8638
rect 6487 8624 6517 8638
rect 6578 8636 6731 8682
rect 6560 8624 6752 8636
rect 6795 8624 6825 8638
rect 6831 8624 6844 8640
rect 6932 8624 6945 8640
rect 6975 8624 6988 8640
rect 7077 8638 7090 8640
rect 7043 8624 7058 8638
rect 7067 8624 7097 8638
rect 7158 8636 7311 8682
rect 7140 8624 7332 8636
rect 7375 8624 7405 8638
rect 7411 8624 7424 8640
rect 7512 8624 7525 8640
rect 7555 8624 7568 8640
rect 7657 8638 7670 8640
rect 7623 8624 7638 8638
rect 7647 8624 7677 8638
rect 7738 8636 7891 8682
rect 7720 8624 7912 8636
rect 7955 8624 7985 8638
rect 7991 8624 8004 8640
rect 8092 8624 8105 8640
rect 8135 8624 8148 8640
rect 8237 8638 8250 8640
rect 8203 8624 8218 8638
rect 8227 8624 8257 8638
rect 8318 8636 8471 8682
rect 8300 8624 8492 8636
rect 8535 8624 8565 8638
rect 8571 8624 8584 8640
rect 8672 8624 8685 8640
rect 8715 8624 8728 8640
rect 8817 8638 8830 8640
rect 8783 8624 8798 8638
rect 8807 8624 8837 8638
rect 8898 8636 9051 8682
rect 8880 8624 9072 8636
rect 9115 8624 9145 8638
rect 9151 8624 9164 8640
rect 9252 8624 9265 8640
rect 0 8610 9265 8624
rect 15 8506 28 8610
rect 73 8588 74 8598
rect 89 8588 102 8598
rect 73 8584 102 8588
rect 107 8584 137 8610
rect 155 8596 171 8598
rect 243 8596 296 8610
rect 244 8594 308 8596
rect 351 8594 366 8610
rect 415 8607 445 8610
rect 415 8604 451 8607
rect 381 8596 397 8598
rect 155 8584 170 8588
rect 73 8582 170 8584
rect 198 8582 366 8594
rect 382 8584 397 8588
rect 415 8585 454 8604
rect 473 8598 480 8599
rect 479 8591 480 8598
rect 463 8588 464 8591
rect 479 8588 492 8591
rect 415 8584 445 8585
rect 454 8584 460 8585
rect 463 8584 492 8588
rect 382 8583 492 8584
rect 382 8582 498 8583
rect 57 8574 108 8582
rect 57 8562 82 8574
rect 89 8562 108 8574
rect 139 8574 189 8582
rect 139 8566 155 8574
rect 162 8572 189 8574
rect 198 8572 419 8582
rect 162 8562 419 8572
rect 448 8574 498 8582
rect 448 8565 464 8574
rect 57 8554 108 8562
rect 155 8554 419 8562
rect 445 8562 464 8565
rect 471 8562 498 8574
rect 445 8554 498 8562
rect 73 8546 74 8554
rect 89 8546 102 8554
rect 73 8538 89 8546
rect 70 8531 89 8534
rect 70 8522 92 8531
rect 43 8512 92 8522
rect 43 8506 73 8512
rect 92 8507 97 8512
rect 15 8490 89 8506
rect 107 8498 137 8554
rect 172 8544 380 8554
rect 415 8550 460 8554
rect 463 8553 464 8554
rect 479 8553 492 8554
rect 198 8514 387 8544
rect 213 8511 387 8514
rect 206 8508 387 8511
rect 15 8488 28 8490
rect 43 8488 77 8490
rect 15 8472 89 8488
rect 116 8484 129 8498
rect 144 8484 160 8500
rect 206 8495 217 8508
rect -1 8450 0 8466
rect 15 8450 28 8472
rect 43 8450 73 8472
rect 116 8468 178 8484
rect 206 8477 217 8493
rect 222 8488 232 8508
rect 242 8488 256 8508
rect 259 8495 268 8508
rect 284 8495 293 8508
rect 222 8477 256 8488
rect 259 8477 268 8493
rect 284 8477 293 8493
rect 300 8488 310 8508
rect 320 8488 334 8508
rect 335 8495 346 8508
rect 300 8477 334 8488
rect 335 8477 346 8493
rect 392 8484 408 8500
rect 415 8498 445 8550
rect 479 8546 480 8553
rect 464 8538 480 8546
rect 451 8506 464 8525
rect 479 8506 509 8522
rect 451 8490 525 8506
rect 451 8488 464 8490
rect 479 8488 513 8490
rect 116 8466 129 8468
rect 144 8466 178 8468
rect 116 8450 178 8466
rect 222 8461 238 8464
rect 300 8461 330 8472
rect 378 8468 424 8484
rect 451 8472 525 8488
rect 378 8466 412 8468
rect 377 8450 424 8466
rect 451 8450 464 8472
rect 479 8450 509 8472
rect 536 8450 537 8466
rect 552 8450 565 8610
rect 595 8506 608 8610
rect 653 8588 654 8598
rect 669 8588 682 8598
rect 653 8584 682 8588
rect 687 8584 717 8610
rect 735 8596 751 8598
rect 823 8596 876 8610
rect 824 8594 888 8596
rect 931 8594 946 8610
rect 995 8607 1025 8610
rect 995 8604 1031 8607
rect 961 8596 977 8598
rect 735 8584 750 8588
rect 653 8582 750 8584
rect 778 8582 946 8594
rect 962 8584 977 8588
rect 995 8585 1034 8604
rect 1053 8598 1060 8599
rect 1059 8591 1060 8598
rect 1043 8588 1044 8591
rect 1059 8588 1072 8591
rect 995 8584 1025 8585
rect 1034 8584 1040 8585
rect 1043 8584 1072 8588
rect 962 8583 1072 8584
rect 962 8582 1078 8583
rect 637 8574 688 8582
rect 637 8562 662 8574
rect 669 8562 688 8574
rect 719 8574 769 8582
rect 719 8566 735 8574
rect 742 8572 769 8574
rect 778 8572 999 8582
rect 742 8562 999 8572
rect 1028 8574 1078 8582
rect 1028 8565 1044 8574
rect 637 8554 688 8562
rect 735 8554 999 8562
rect 1025 8562 1044 8565
rect 1051 8562 1078 8574
rect 1025 8554 1078 8562
rect 653 8546 654 8554
rect 669 8546 682 8554
rect 653 8538 669 8546
rect 650 8531 669 8534
rect 650 8522 672 8531
rect 623 8512 672 8522
rect 623 8506 653 8512
rect 672 8507 677 8512
rect 595 8490 669 8506
rect 687 8498 717 8554
rect 752 8544 960 8554
rect 995 8550 1040 8554
rect 1043 8553 1044 8554
rect 1059 8553 1072 8554
rect 778 8514 967 8544
rect 793 8511 967 8514
rect 786 8508 967 8511
rect 595 8488 608 8490
rect 623 8488 657 8490
rect 595 8472 669 8488
rect 696 8484 709 8498
rect 724 8484 740 8500
rect 786 8495 797 8508
rect 579 8450 580 8466
rect 595 8450 608 8472
rect 623 8450 653 8472
rect 696 8468 758 8484
rect 786 8477 797 8493
rect 802 8488 812 8508
rect 822 8488 836 8508
rect 839 8495 848 8508
rect 864 8495 873 8508
rect 802 8477 836 8488
rect 839 8477 848 8493
rect 864 8477 873 8493
rect 880 8488 890 8508
rect 900 8488 914 8508
rect 915 8495 926 8508
rect 880 8477 914 8488
rect 915 8477 926 8493
rect 972 8484 988 8500
rect 995 8498 1025 8550
rect 1059 8546 1060 8553
rect 1044 8538 1060 8546
rect 1031 8506 1044 8525
rect 1059 8506 1089 8522
rect 1031 8490 1105 8506
rect 1031 8488 1044 8490
rect 1059 8488 1093 8490
rect 696 8466 709 8468
rect 724 8466 758 8468
rect 696 8450 758 8466
rect 802 8461 818 8464
rect 880 8461 910 8472
rect 958 8468 1004 8484
rect 1031 8472 1105 8488
rect 958 8466 992 8468
rect 957 8450 1004 8466
rect 1031 8450 1044 8472
rect 1059 8450 1089 8472
rect 1116 8450 1117 8466
rect 1132 8450 1145 8610
rect 1175 8506 1188 8610
rect 1233 8588 1234 8598
rect 1249 8588 1262 8598
rect 1233 8584 1262 8588
rect 1267 8584 1297 8610
rect 1315 8596 1331 8598
rect 1403 8596 1456 8610
rect 1404 8594 1468 8596
rect 1511 8594 1526 8610
rect 1575 8607 1605 8610
rect 1575 8604 1611 8607
rect 1541 8596 1557 8598
rect 1315 8584 1330 8588
rect 1233 8582 1330 8584
rect 1358 8582 1526 8594
rect 1542 8584 1557 8588
rect 1575 8585 1614 8604
rect 1633 8598 1640 8599
rect 1639 8591 1640 8598
rect 1623 8588 1624 8591
rect 1639 8588 1652 8591
rect 1575 8584 1605 8585
rect 1614 8584 1620 8585
rect 1623 8584 1652 8588
rect 1542 8583 1652 8584
rect 1542 8582 1658 8583
rect 1217 8574 1268 8582
rect 1217 8562 1242 8574
rect 1249 8562 1268 8574
rect 1299 8574 1349 8582
rect 1299 8566 1315 8574
rect 1322 8572 1349 8574
rect 1358 8572 1579 8582
rect 1322 8562 1579 8572
rect 1608 8574 1658 8582
rect 1608 8565 1624 8574
rect 1217 8554 1268 8562
rect 1315 8554 1579 8562
rect 1605 8562 1624 8565
rect 1631 8562 1658 8574
rect 1605 8554 1658 8562
rect 1233 8546 1234 8554
rect 1249 8546 1262 8554
rect 1233 8538 1249 8546
rect 1230 8531 1249 8534
rect 1230 8522 1252 8531
rect 1203 8512 1252 8522
rect 1203 8506 1233 8512
rect 1252 8507 1257 8512
rect 1175 8490 1249 8506
rect 1267 8498 1297 8554
rect 1332 8544 1540 8554
rect 1575 8550 1620 8554
rect 1623 8553 1624 8554
rect 1639 8553 1652 8554
rect 1358 8514 1547 8544
rect 1373 8511 1547 8514
rect 1366 8508 1547 8511
rect 1175 8488 1188 8490
rect 1203 8488 1237 8490
rect 1175 8472 1249 8488
rect 1276 8484 1289 8498
rect 1304 8484 1320 8500
rect 1366 8495 1377 8508
rect 1159 8450 1160 8466
rect 1175 8450 1188 8472
rect 1203 8450 1233 8472
rect 1276 8468 1338 8484
rect 1366 8477 1377 8493
rect 1382 8488 1392 8508
rect 1402 8488 1416 8508
rect 1419 8495 1428 8508
rect 1444 8495 1453 8508
rect 1382 8477 1416 8488
rect 1419 8477 1428 8493
rect 1444 8477 1453 8493
rect 1460 8488 1470 8508
rect 1480 8488 1494 8508
rect 1495 8495 1506 8508
rect 1460 8477 1494 8488
rect 1495 8477 1506 8493
rect 1552 8484 1568 8500
rect 1575 8498 1605 8550
rect 1639 8546 1640 8553
rect 1624 8538 1640 8546
rect 1611 8506 1624 8525
rect 1639 8506 1669 8522
rect 1611 8490 1685 8506
rect 1611 8488 1624 8490
rect 1639 8488 1673 8490
rect 1276 8466 1289 8468
rect 1304 8466 1338 8468
rect 1276 8450 1338 8466
rect 1382 8461 1398 8464
rect 1460 8461 1490 8472
rect 1538 8468 1584 8484
rect 1611 8472 1685 8488
rect 1538 8466 1572 8468
rect 1537 8450 1584 8466
rect 1611 8450 1624 8472
rect 1639 8450 1669 8472
rect 1696 8450 1697 8466
rect 1712 8450 1725 8610
rect 1755 8506 1768 8610
rect 1813 8588 1814 8598
rect 1829 8588 1842 8598
rect 1813 8584 1842 8588
rect 1847 8584 1877 8610
rect 1895 8596 1911 8598
rect 1983 8596 2036 8610
rect 1984 8594 2048 8596
rect 2091 8594 2106 8610
rect 2155 8607 2185 8610
rect 2155 8604 2191 8607
rect 2121 8596 2137 8598
rect 1895 8584 1910 8588
rect 1813 8582 1910 8584
rect 1938 8582 2106 8594
rect 2122 8584 2137 8588
rect 2155 8585 2194 8604
rect 2213 8598 2220 8599
rect 2219 8591 2220 8598
rect 2203 8588 2204 8591
rect 2219 8588 2232 8591
rect 2155 8584 2185 8585
rect 2194 8584 2200 8585
rect 2203 8584 2232 8588
rect 2122 8583 2232 8584
rect 2122 8582 2238 8583
rect 1797 8574 1848 8582
rect 1797 8562 1822 8574
rect 1829 8562 1848 8574
rect 1879 8574 1929 8582
rect 1879 8566 1895 8574
rect 1902 8572 1929 8574
rect 1938 8572 2159 8582
rect 1902 8562 2159 8572
rect 2188 8574 2238 8582
rect 2188 8565 2204 8574
rect 1797 8554 1848 8562
rect 1895 8554 2159 8562
rect 2185 8562 2204 8565
rect 2211 8562 2238 8574
rect 2185 8554 2238 8562
rect 1813 8546 1814 8554
rect 1829 8546 1842 8554
rect 1813 8538 1829 8546
rect 1810 8531 1829 8534
rect 1810 8522 1832 8531
rect 1783 8512 1832 8522
rect 1783 8506 1813 8512
rect 1832 8507 1837 8512
rect 1755 8490 1829 8506
rect 1847 8498 1877 8554
rect 1912 8544 2120 8554
rect 2155 8550 2200 8554
rect 2203 8553 2204 8554
rect 2219 8553 2232 8554
rect 1938 8514 2127 8544
rect 1953 8511 2127 8514
rect 1946 8508 2127 8511
rect 1755 8488 1768 8490
rect 1783 8488 1817 8490
rect 1755 8472 1829 8488
rect 1856 8484 1869 8498
rect 1884 8484 1900 8500
rect 1946 8495 1957 8508
rect 1739 8450 1740 8466
rect 1755 8450 1768 8472
rect 1783 8450 1813 8472
rect 1856 8468 1918 8484
rect 1946 8477 1957 8493
rect 1962 8488 1972 8508
rect 1982 8488 1996 8508
rect 1999 8495 2008 8508
rect 2024 8495 2033 8508
rect 1962 8477 1996 8488
rect 1999 8477 2008 8493
rect 2024 8477 2033 8493
rect 2040 8488 2050 8508
rect 2060 8488 2074 8508
rect 2075 8495 2086 8508
rect 2040 8477 2074 8488
rect 2075 8477 2086 8493
rect 2132 8484 2148 8500
rect 2155 8498 2185 8550
rect 2219 8546 2220 8553
rect 2204 8538 2220 8546
rect 2191 8506 2204 8525
rect 2219 8506 2249 8522
rect 2191 8490 2265 8506
rect 2191 8488 2204 8490
rect 2219 8488 2253 8490
rect 1856 8466 1869 8468
rect 1884 8466 1918 8468
rect 1856 8450 1918 8466
rect 1962 8461 1976 8464
rect 2040 8461 2070 8472
rect 2118 8468 2164 8484
rect 2191 8472 2265 8488
rect 2118 8466 2152 8468
rect 2117 8450 2164 8466
rect 2191 8450 2204 8472
rect 2219 8450 2249 8472
rect 2276 8450 2277 8466
rect 2292 8450 2305 8610
rect 2335 8506 2348 8610
rect 2393 8588 2394 8598
rect 2409 8588 2422 8598
rect 2393 8584 2422 8588
rect 2427 8584 2457 8610
rect 2475 8596 2491 8598
rect 2563 8596 2616 8610
rect 2564 8594 2628 8596
rect 2671 8594 2686 8610
rect 2735 8607 2765 8610
rect 2735 8604 2771 8607
rect 2701 8596 2717 8598
rect 2475 8584 2490 8588
rect 2393 8582 2490 8584
rect 2518 8582 2686 8594
rect 2702 8584 2717 8588
rect 2735 8585 2774 8604
rect 2793 8598 2800 8599
rect 2799 8591 2800 8598
rect 2783 8588 2784 8591
rect 2799 8588 2812 8591
rect 2735 8584 2765 8585
rect 2774 8584 2780 8585
rect 2783 8584 2812 8588
rect 2702 8583 2812 8584
rect 2702 8582 2818 8583
rect 2377 8574 2428 8582
rect 2377 8562 2402 8574
rect 2409 8562 2428 8574
rect 2459 8574 2509 8582
rect 2459 8566 2475 8574
rect 2482 8572 2509 8574
rect 2518 8572 2739 8582
rect 2482 8562 2739 8572
rect 2768 8574 2818 8582
rect 2768 8565 2784 8574
rect 2377 8554 2428 8562
rect 2475 8554 2739 8562
rect 2765 8562 2784 8565
rect 2791 8562 2818 8574
rect 2765 8554 2818 8562
rect 2393 8546 2394 8554
rect 2409 8546 2422 8554
rect 2393 8538 2409 8546
rect 2390 8531 2409 8534
rect 2390 8522 2412 8531
rect 2363 8512 2412 8522
rect 2363 8506 2393 8512
rect 2412 8507 2417 8512
rect 2335 8490 2409 8506
rect 2427 8498 2457 8554
rect 2492 8544 2700 8554
rect 2735 8550 2780 8554
rect 2783 8553 2784 8554
rect 2799 8553 2812 8554
rect 2518 8514 2707 8544
rect 2533 8511 2707 8514
rect 2526 8508 2707 8511
rect 2335 8488 2348 8490
rect 2363 8488 2397 8490
rect 2335 8472 2409 8488
rect 2436 8484 2449 8498
rect 2464 8484 2480 8500
rect 2526 8495 2537 8508
rect 2319 8450 2320 8466
rect 2335 8450 2348 8472
rect 2363 8450 2393 8472
rect 2436 8468 2498 8484
rect 2526 8477 2537 8493
rect 2542 8488 2552 8508
rect 2562 8488 2576 8508
rect 2579 8495 2588 8508
rect 2604 8495 2613 8508
rect 2542 8477 2576 8488
rect 2579 8477 2588 8493
rect 2604 8477 2613 8493
rect 2620 8488 2630 8508
rect 2640 8488 2654 8508
rect 2655 8495 2666 8508
rect 2620 8477 2654 8488
rect 2655 8477 2666 8493
rect 2712 8484 2728 8500
rect 2735 8498 2765 8550
rect 2799 8546 2800 8553
rect 2784 8538 2800 8546
rect 2771 8506 2784 8525
rect 2799 8506 2829 8522
rect 2771 8490 2845 8506
rect 2771 8488 2784 8490
rect 2799 8488 2833 8490
rect 2436 8466 2449 8468
rect 2464 8466 2498 8468
rect 2436 8450 2498 8466
rect 2542 8461 2558 8464
rect 2620 8461 2650 8472
rect 2698 8468 2744 8484
rect 2771 8472 2845 8488
rect 2698 8466 2732 8468
rect 2697 8450 2744 8466
rect 2771 8450 2784 8472
rect 2799 8450 2829 8472
rect 2856 8450 2857 8466
rect 2872 8450 2885 8610
rect 2915 8506 2928 8610
rect 2973 8588 2974 8598
rect 2989 8588 3002 8598
rect 2973 8584 3002 8588
rect 3007 8584 3037 8610
rect 3055 8596 3071 8598
rect 3143 8596 3196 8610
rect 3144 8594 3208 8596
rect 3251 8594 3266 8610
rect 3315 8607 3345 8610
rect 3315 8604 3351 8607
rect 3281 8596 3297 8598
rect 3055 8584 3070 8588
rect 2973 8582 3070 8584
rect 3098 8582 3266 8594
rect 3282 8584 3297 8588
rect 3315 8585 3354 8604
rect 3373 8598 3380 8599
rect 3379 8591 3380 8598
rect 3363 8588 3364 8591
rect 3379 8588 3392 8591
rect 3315 8584 3345 8585
rect 3354 8584 3360 8585
rect 3363 8584 3392 8588
rect 3282 8583 3392 8584
rect 3282 8582 3398 8583
rect 2957 8574 3008 8582
rect 2957 8562 2982 8574
rect 2989 8562 3008 8574
rect 3039 8574 3089 8582
rect 3039 8566 3055 8574
rect 3062 8572 3089 8574
rect 3098 8572 3319 8582
rect 3062 8562 3319 8572
rect 3348 8574 3398 8582
rect 3348 8565 3364 8574
rect 2957 8554 3008 8562
rect 3055 8554 3319 8562
rect 3345 8562 3364 8565
rect 3371 8562 3398 8574
rect 3345 8554 3398 8562
rect 2973 8546 2974 8554
rect 2989 8546 3002 8554
rect 2973 8538 2989 8546
rect 2970 8531 2989 8534
rect 2970 8522 2992 8531
rect 2943 8512 2992 8522
rect 2943 8506 2973 8512
rect 2992 8507 2997 8512
rect 2915 8490 2989 8506
rect 3007 8498 3037 8554
rect 3072 8544 3280 8554
rect 3315 8550 3360 8554
rect 3363 8553 3364 8554
rect 3379 8553 3392 8554
rect 3098 8514 3287 8544
rect 3113 8511 3287 8514
rect 3106 8508 3287 8511
rect 2915 8488 2928 8490
rect 2943 8488 2977 8490
rect 2915 8472 2989 8488
rect 3016 8484 3029 8498
rect 3044 8484 3060 8500
rect 3106 8495 3117 8508
rect 2899 8450 2900 8466
rect 2915 8450 2928 8472
rect 2943 8450 2973 8472
rect 3016 8468 3078 8484
rect 3106 8477 3117 8493
rect 3122 8488 3132 8508
rect 3142 8488 3156 8508
rect 3159 8495 3168 8508
rect 3184 8495 3193 8508
rect 3122 8477 3156 8488
rect 3159 8477 3168 8493
rect 3184 8477 3193 8493
rect 3200 8488 3210 8508
rect 3220 8488 3234 8508
rect 3235 8495 3246 8508
rect 3200 8477 3234 8488
rect 3235 8477 3246 8493
rect 3292 8484 3308 8500
rect 3315 8498 3345 8550
rect 3379 8546 3380 8553
rect 3364 8538 3380 8546
rect 3351 8506 3364 8525
rect 3379 8506 3409 8522
rect 3351 8490 3425 8506
rect 3351 8488 3364 8490
rect 3379 8488 3413 8490
rect 3016 8466 3029 8468
rect 3044 8466 3078 8468
rect 3016 8450 3078 8466
rect 3122 8461 3138 8464
rect 3200 8461 3230 8472
rect 3278 8468 3324 8484
rect 3351 8472 3425 8488
rect 3278 8466 3312 8468
rect 3277 8450 3324 8466
rect 3351 8450 3364 8472
rect 3379 8450 3409 8472
rect 3436 8450 3437 8466
rect 3452 8450 3465 8610
rect 3495 8506 3508 8610
rect 3553 8588 3554 8598
rect 3569 8588 3582 8598
rect 3553 8584 3582 8588
rect 3587 8584 3617 8610
rect 3635 8596 3651 8598
rect 3723 8596 3776 8610
rect 3724 8594 3788 8596
rect 3831 8594 3846 8610
rect 3895 8607 3925 8610
rect 3895 8604 3931 8607
rect 3861 8596 3877 8598
rect 3635 8584 3650 8588
rect 3553 8582 3650 8584
rect 3678 8582 3846 8594
rect 3862 8584 3877 8588
rect 3895 8585 3934 8604
rect 3953 8598 3960 8599
rect 3959 8591 3960 8598
rect 3943 8588 3944 8591
rect 3959 8588 3972 8591
rect 3895 8584 3925 8585
rect 3934 8584 3940 8585
rect 3943 8584 3972 8588
rect 3862 8583 3972 8584
rect 3862 8582 3978 8583
rect 3537 8574 3588 8582
rect 3537 8562 3562 8574
rect 3569 8562 3588 8574
rect 3619 8574 3669 8582
rect 3619 8566 3635 8574
rect 3642 8572 3669 8574
rect 3678 8572 3899 8582
rect 3642 8562 3899 8572
rect 3928 8574 3978 8582
rect 3928 8565 3944 8574
rect 3537 8554 3588 8562
rect 3635 8554 3899 8562
rect 3925 8562 3944 8565
rect 3951 8562 3978 8574
rect 3925 8554 3978 8562
rect 3553 8546 3554 8554
rect 3569 8546 3582 8554
rect 3553 8538 3569 8546
rect 3550 8531 3569 8534
rect 3550 8522 3572 8531
rect 3523 8512 3572 8522
rect 3523 8506 3553 8512
rect 3572 8507 3577 8512
rect 3495 8490 3569 8506
rect 3587 8498 3617 8554
rect 3652 8544 3860 8554
rect 3895 8550 3940 8554
rect 3943 8553 3944 8554
rect 3959 8553 3972 8554
rect 3678 8514 3867 8544
rect 3693 8511 3867 8514
rect 3686 8508 3867 8511
rect 3495 8488 3508 8490
rect 3523 8488 3557 8490
rect 3495 8472 3569 8488
rect 3596 8484 3609 8498
rect 3624 8484 3640 8500
rect 3686 8495 3697 8508
rect 3479 8450 3480 8466
rect 3495 8450 3508 8472
rect 3523 8450 3553 8472
rect 3596 8468 3658 8484
rect 3686 8477 3697 8493
rect 3702 8488 3712 8508
rect 3722 8488 3736 8508
rect 3739 8495 3748 8508
rect 3764 8495 3773 8508
rect 3702 8477 3736 8488
rect 3739 8477 3748 8493
rect 3764 8477 3773 8493
rect 3780 8488 3790 8508
rect 3800 8488 3814 8508
rect 3815 8495 3826 8508
rect 3780 8477 3814 8488
rect 3815 8477 3826 8493
rect 3872 8484 3888 8500
rect 3895 8498 3925 8550
rect 3959 8546 3960 8553
rect 3944 8538 3960 8546
rect 3931 8506 3944 8525
rect 3959 8506 3989 8522
rect 3931 8490 4005 8506
rect 3931 8488 3944 8490
rect 3959 8488 3993 8490
rect 3596 8466 3609 8468
rect 3624 8466 3658 8468
rect 3596 8450 3658 8466
rect 3702 8461 3718 8464
rect 3780 8461 3810 8472
rect 3858 8468 3904 8484
rect 3931 8472 4005 8488
rect 3858 8466 3892 8468
rect 3857 8450 3904 8466
rect 3931 8450 3944 8472
rect 3959 8450 3989 8472
rect 4016 8450 4017 8466
rect 4032 8450 4045 8610
rect 4075 8506 4088 8610
rect 4133 8588 4134 8598
rect 4149 8588 4162 8598
rect 4133 8584 4162 8588
rect 4167 8584 4197 8610
rect 4215 8596 4231 8598
rect 4303 8596 4356 8610
rect 4304 8594 4368 8596
rect 4411 8594 4426 8610
rect 4475 8607 4505 8610
rect 4475 8604 4511 8607
rect 4441 8596 4457 8598
rect 4215 8584 4230 8588
rect 4133 8582 4230 8584
rect 4258 8582 4426 8594
rect 4442 8584 4457 8588
rect 4475 8585 4514 8604
rect 4533 8598 4540 8599
rect 4539 8591 4540 8598
rect 4523 8588 4524 8591
rect 4539 8588 4552 8591
rect 4475 8584 4505 8585
rect 4514 8584 4520 8585
rect 4523 8584 4552 8588
rect 4442 8583 4552 8584
rect 4442 8582 4558 8583
rect 4117 8574 4168 8582
rect 4117 8562 4142 8574
rect 4149 8562 4168 8574
rect 4199 8574 4249 8582
rect 4199 8566 4215 8574
rect 4222 8572 4249 8574
rect 4258 8572 4479 8582
rect 4222 8562 4479 8572
rect 4508 8574 4558 8582
rect 4508 8565 4524 8574
rect 4117 8554 4168 8562
rect 4215 8554 4479 8562
rect 4505 8562 4524 8565
rect 4531 8562 4558 8574
rect 4505 8554 4558 8562
rect 4133 8546 4134 8554
rect 4149 8546 4162 8554
rect 4133 8538 4149 8546
rect 4130 8531 4149 8534
rect 4130 8522 4152 8531
rect 4103 8512 4152 8522
rect 4103 8506 4133 8512
rect 4152 8507 4157 8512
rect 4075 8490 4149 8506
rect 4167 8498 4197 8554
rect 4232 8544 4440 8554
rect 4475 8550 4520 8554
rect 4523 8553 4524 8554
rect 4539 8553 4552 8554
rect 4258 8514 4447 8544
rect 4273 8511 4447 8514
rect 4266 8508 4447 8511
rect 4075 8488 4088 8490
rect 4103 8488 4137 8490
rect 4075 8472 4149 8488
rect 4176 8484 4189 8498
rect 4204 8484 4220 8500
rect 4266 8495 4277 8508
rect 4059 8450 4060 8466
rect 4075 8450 4088 8472
rect 4103 8450 4133 8472
rect 4176 8468 4238 8484
rect 4266 8477 4277 8493
rect 4282 8488 4292 8508
rect 4302 8488 4316 8508
rect 4319 8495 4328 8508
rect 4344 8495 4353 8508
rect 4282 8477 4316 8488
rect 4319 8477 4328 8493
rect 4344 8477 4353 8493
rect 4360 8488 4370 8508
rect 4380 8488 4394 8508
rect 4395 8495 4406 8508
rect 4360 8477 4394 8488
rect 4395 8477 4406 8493
rect 4452 8484 4468 8500
rect 4475 8498 4505 8550
rect 4539 8546 4540 8553
rect 4524 8538 4540 8546
rect 4511 8506 4524 8525
rect 4539 8506 4569 8522
rect 4511 8490 4585 8506
rect 4511 8488 4524 8490
rect 4539 8488 4573 8490
rect 4176 8466 4189 8468
rect 4204 8466 4238 8468
rect 4176 8450 4238 8466
rect 4282 8461 4298 8464
rect 4360 8461 4390 8472
rect 4438 8468 4484 8484
rect 4511 8472 4585 8488
rect 4438 8466 4472 8468
rect 4437 8450 4484 8466
rect 4511 8450 4524 8472
rect 4539 8450 4569 8472
rect 4596 8450 4597 8466
rect 4612 8450 4625 8610
rect 4655 8506 4668 8610
rect 4713 8588 4714 8598
rect 4729 8588 4742 8598
rect 4713 8584 4742 8588
rect 4747 8584 4777 8610
rect 4795 8596 4811 8598
rect 4883 8596 4936 8610
rect 4884 8594 4948 8596
rect 4991 8594 5006 8610
rect 5055 8607 5085 8610
rect 5055 8604 5091 8607
rect 5021 8596 5037 8598
rect 4795 8584 4810 8588
rect 4713 8582 4810 8584
rect 4838 8582 5006 8594
rect 5022 8584 5037 8588
rect 5055 8585 5094 8604
rect 5113 8598 5120 8599
rect 5119 8591 5120 8598
rect 5103 8588 5104 8591
rect 5119 8588 5132 8591
rect 5055 8584 5085 8585
rect 5094 8584 5100 8585
rect 5103 8584 5132 8588
rect 5022 8583 5132 8584
rect 5022 8582 5138 8583
rect 4697 8574 4748 8582
rect 4697 8562 4722 8574
rect 4729 8562 4748 8574
rect 4779 8574 4829 8582
rect 4779 8566 4795 8574
rect 4802 8572 4829 8574
rect 4838 8572 5059 8582
rect 4802 8562 5059 8572
rect 5088 8574 5138 8582
rect 5088 8565 5104 8574
rect 4697 8554 4748 8562
rect 4795 8554 5059 8562
rect 5085 8562 5104 8565
rect 5111 8562 5138 8574
rect 5085 8554 5138 8562
rect 4713 8546 4714 8554
rect 4729 8546 4742 8554
rect 4713 8538 4729 8546
rect 4710 8531 4729 8534
rect 4710 8522 4732 8531
rect 4683 8512 4732 8522
rect 4683 8506 4713 8512
rect 4732 8507 4737 8512
rect 4655 8490 4729 8506
rect 4747 8498 4777 8554
rect 4812 8544 5020 8554
rect 5055 8550 5100 8554
rect 5103 8553 5104 8554
rect 5119 8553 5132 8554
rect 4838 8514 5027 8544
rect 4853 8511 5027 8514
rect 4846 8508 5027 8511
rect 4655 8488 4668 8490
rect 4683 8488 4717 8490
rect 4655 8472 4729 8488
rect 4756 8484 4769 8498
rect 4784 8484 4800 8500
rect 4846 8495 4857 8508
rect 4639 8450 4640 8466
rect 4655 8450 4668 8472
rect 4683 8450 4713 8472
rect 4756 8468 4818 8484
rect 4846 8477 4857 8493
rect 4862 8488 4872 8508
rect 4882 8488 4896 8508
rect 4899 8495 4908 8508
rect 4924 8495 4933 8508
rect 4862 8477 4896 8488
rect 4899 8477 4908 8493
rect 4924 8477 4933 8493
rect 4940 8488 4950 8508
rect 4960 8488 4974 8508
rect 4975 8495 4986 8508
rect 4940 8477 4974 8488
rect 4975 8477 4986 8493
rect 5032 8484 5048 8500
rect 5055 8498 5085 8550
rect 5119 8546 5120 8553
rect 5104 8538 5120 8546
rect 5091 8506 5104 8525
rect 5119 8506 5149 8522
rect 5091 8490 5165 8506
rect 5091 8488 5104 8490
rect 5119 8488 5153 8490
rect 4756 8466 4769 8468
rect 4784 8466 4818 8468
rect 4756 8450 4818 8466
rect 4862 8461 4878 8464
rect 4940 8461 4970 8472
rect 5018 8468 5064 8484
rect 5091 8472 5165 8488
rect 5018 8466 5052 8468
rect 5017 8450 5064 8466
rect 5091 8450 5104 8472
rect 5119 8450 5149 8472
rect 5176 8450 5177 8466
rect 5192 8450 5205 8610
rect 5235 8506 5248 8610
rect 5293 8588 5294 8598
rect 5309 8588 5322 8598
rect 5293 8584 5322 8588
rect 5327 8584 5357 8610
rect 5375 8596 5391 8598
rect 5463 8596 5516 8610
rect 5464 8594 5528 8596
rect 5571 8594 5586 8610
rect 5635 8607 5665 8610
rect 5635 8604 5671 8607
rect 5601 8596 5617 8598
rect 5375 8584 5390 8588
rect 5293 8582 5390 8584
rect 5418 8582 5586 8594
rect 5602 8584 5617 8588
rect 5635 8585 5674 8604
rect 5693 8598 5700 8599
rect 5699 8591 5700 8598
rect 5683 8588 5684 8591
rect 5699 8588 5712 8591
rect 5635 8584 5665 8585
rect 5674 8584 5680 8585
rect 5683 8584 5712 8588
rect 5602 8583 5712 8584
rect 5602 8582 5718 8583
rect 5277 8574 5328 8582
rect 5277 8562 5302 8574
rect 5309 8562 5328 8574
rect 5359 8574 5409 8582
rect 5359 8566 5375 8574
rect 5382 8572 5409 8574
rect 5418 8572 5639 8582
rect 5382 8562 5639 8572
rect 5668 8574 5718 8582
rect 5668 8565 5684 8574
rect 5277 8554 5328 8562
rect 5375 8554 5639 8562
rect 5665 8562 5684 8565
rect 5691 8562 5718 8574
rect 5665 8554 5718 8562
rect 5293 8546 5294 8554
rect 5309 8546 5322 8554
rect 5293 8538 5309 8546
rect 5290 8531 5309 8534
rect 5290 8522 5312 8531
rect 5263 8512 5312 8522
rect 5263 8506 5293 8512
rect 5312 8507 5317 8512
rect 5235 8490 5309 8506
rect 5327 8498 5357 8554
rect 5392 8544 5600 8554
rect 5635 8550 5680 8554
rect 5683 8553 5684 8554
rect 5699 8553 5712 8554
rect 5418 8514 5607 8544
rect 5433 8511 5607 8514
rect 5426 8508 5607 8511
rect 5235 8488 5248 8490
rect 5263 8488 5297 8490
rect 5235 8472 5309 8488
rect 5336 8484 5349 8498
rect 5364 8484 5380 8500
rect 5426 8495 5437 8508
rect 5219 8450 5220 8466
rect 5235 8450 5248 8472
rect 5263 8450 5293 8472
rect 5336 8468 5398 8484
rect 5426 8477 5437 8493
rect 5442 8488 5452 8508
rect 5462 8488 5476 8508
rect 5479 8495 5488 8508
rect 5504 8495 5513 8508
rect 5442 8477 5476 8488
rect 5479 8477 5488 8493
rect 5504 8477 5513 8493
rect 5520 8488 5530 8508
rect 5540 8488 5554 8508
rect 5555 8495 5566 8508
rect 5520 8477 5554 8488
rect 5555 8477 5566 8493
rect 5612 8484 5628 8500
rect 5635 8498 5665 8550
rect 5699 8546 5700 8553
rect 5684 8538 5700 8546
rect 5671 8506 5684 8525
rect 5699 8506 5729 8522
rect 5671 8490 5745 8506
rect 5671 8488 5684 8490
rect 5699 8488 5733 8490
rect 5336 8466 5349 8468
rect 5364 8466 5398 8468
rect 5336 8450 5398 8466
rect 5442 8461 5458 8464
rect 5520 8461 5550 8472
rect 5598 8468 5644 8484
rect 5671 8472 5745 8488
rect 5598 8466 5632 8468
rect 5597 8450 5644 8466
rect 5671 8450 5684 8472
rect 5699 8450 5729 8472
rect 5756 8450 5757 8466
rect 5772 8450 5785 8610
rect 5815 8506 5828 8610
rect 5873 8588 5874 8598
rect 5889 8588 5902 8598
rect 5873 8584 5902 8588
rect 5907 8584 5937 8610
rect 5955 8596 5971 8598
rect 6043 8596 6096 8610
rect 6044 8594 6108 8596
rect 6151 8594 6166 8610
rect 6215 8607 6245 8610
rect 6215 8604 6251 8607
rect 6181 8596 6197 8598
rect 5955 8584 5970 8588
rect 5873 8582 5970 8584
rect 5998 8582 6166 8594
rect 6182 8584 6197 8588
rect 6215 8585 6254 8604
rect 6273 8598 6280 8599
rect 6279 8591 6280 8598
rect 6263 8588 6264 8591
rect 6279 8588 6292 8591
rect 6215 8584 6245 8585
rect 6254 8584 6260 8585
rect 6263 8584 6292 8588
rect 6182 8583 6292 8584
rect 6182 8582 6298 8583
rect 5857 8574 5908 8582
rect 5857 8562 5882 8574
rect 5889 8562 5908 8574
rect 5939 8574 5989 8582
rect 5939 8566 5955 8574
rect 5962 8572 5989 8574
rect 5998 8572 6219 8582
rect 5962 8562 6219 8572
rect 6248 8574 6298 8582
rect 6248 8565 6264 8574
rect 5857 8554 5908 8562
rect 5955 8554 6219 8562
rect 6245 8562 6264 8565
rect 6271 8562 6298 8574
rect 6245 8554 6298 8562
rect 5873 8546 5874 8554
rect 5889 8546 5902 8554
rect 5873 8538 5889 8546
rect 5870 8531 5889 8534
rect 5870 8522 5892 8531
rect 5843 8512 5892 8522
rect 5843 8506 5873 8512
rect 5892 8507 5897 8512
rect 5815 8490 5889 8506
rect 5907 8498 5937 8554
rect 5972 8544 6180 8554
rect 6215 8550 6260 8554
rect 6263 8553 6264 8554
rect 6279 8553 6292 8554
rect 5998 8514 6187 8544
rect 6013 8511 6187 8514
rect 6006 8508 6187 8511
rect 5815 8488 5828 8490
rect 5843 8488 5877 8490
rect 5815 8472 5889 8488
rect 5916 8484 5929 8498
rect 5944 8484 5960 8500
rect 6006 8495 6017 8508
rect 5799 8450 5800 8466
rect 5815 8450 5828 8472
rect 5843 8450 5873 8472
rect 5916 8468 5978 8484
rect 6006 8477 6017 8493
rect 6022 8488 6032 8508
rect 6042 8488 6056 8508
rect 6059 8495 6068 8508
rect 6084 8495 6093 8508
rect 6022 8477 6056 8488
rect 6059 8477 6068 8493
rect 6084 8477 6093 8493
rect 6100 8488 6110 8508
rect 6120 8488 6134 8508
rect 6135 8495 6146 8508
rect 6100 8477 6134 8488
rect 6135 8477 6146 8493
rect 6192 8484 6208 8500
rect 6215 8498 6245 8550
rect 6279 8546 6280 8553
rect 6264 8538 6280 8546
rect 6251 8506 6264 8525
rect 6279 8506 6309 8522
rect 6251 8490 6325 8506
rect 6251 8488 6264 8490
rect 6279 8488 6313 8490
rect 5916 8466 5929 8468
rect 5944 8466 5978 8468
rect 5916 8450 5978 8466
rect 6022 8461 6038 8464
rect 6100 8461 6130 8472
rect 6178 8468 6224 8484
rect 6251 8472 6325 8488
rect 6178 8466 6212 8468
rect 6177 8450 6224 8466
rect 6251 8450 6264 8472
rect 6279 8450 6309 8472
rect 6336 8450 6337 8466
rect 6352 8450 6365 8610
rect 6395 8506 6408 8610
rect 6453 8588 6454 8598
rect 6469 8588 6482 8598
rect 6453 8584 6482 8588
rect 6487 8584 6517 8610
rect 6535 8596 6551 8598
rect 6623 8596 6676 8610
rect 6624 8594 6688 8596
rect 6731 8594 6746 8610
rect 6795 8607 6825 8610
rect 6795 8604 6831 8607
rect 6761 8596 6777 8598
rect 6535 8584 6550 8588
rect 6453 8582 6550 8584
rect 6578 8582 6746 8594
rect 6762 8584 6777 8588
rect 6795 8585 6834 8604
rect 6853 8598 6860 8599
rect 6859 8591 6860 8598
rect 6843 8588 6844 8591
rect 6859 8588 6872 8591
rect 6795 8584 6825 8585
rect 6834 8584 6840 8585
rect 6843 8584 6872 8588
rect 6762 8583 6872 8584
rect 6762 8582 6878 8583
rect 6437 8574 6488 8582
rect 6437 8562 6462 8574
rect 6469 8562 6488 8574
rect 6519 8574 6569 8582
rect 6519 8566 6535 8574
rect 6542 8572 6569 8574
rect 6578 8572 6799 8582
rect 6542 8562 6799 8572
rect 6828 8574 6878 8582
rect 6828 8565 6844 8574
rect 6437 8554 6488 8562
rect 6535 8554 6799 8562
rect 6825 8562 6844 8565
rect 6851 8562 6878 8574
rect 6825 8554 6878 8562
rect 6453 8546 6454 8554
rect 6469 8546 6482 8554
rect 6453 8538 6469 8546
rect 6450 8531 6469 8534
rect 6450 8522 6472 8531
rect 6423 8512 6472 8522
rect 6423 8506 6453 8512
rect 6472 8507 6477 8512
rect 6395 8490 6469 8506
rect 6487 8498 6517 8554
rect 6552 8544 6760 8554
rect 6795 8550 6840 8554
rect 6843 8553 6844 8554
rect 6859 8553 6872 8554
rect 6578 8514 6767 8544
rect 6593 8511 6767 8514
rect 6586 8508 6767 8511
rect 6395 8488 6408 8490
rect 6423 8488 6457 8490
rect 6395 8472 6469 8488
rect 6496 8484 6509 8498
rect 6524 8484 6540 8500
rect 6586 8495 6597 8508
rect 6379 8450 6380 8466
rect 6395 8450 6408 8472
rect 6423 8450 6453 8472
rect 6496 8468 6558 8484
rect 6586 8477 6597 8493
rect 6602 8488 6612 8508
rect 6622 8488 6636 8508
rect 6639 8495 6648 8508
rect 6664 8495 6673 8508
rect 6602 8477 6636 8488
rect 6639 8477 6648 8493
rect 6664 8477 6673 8493
rect 6680 8488 6690 8508
rect 6700 8488 6714 8508
rect 6715 8495 6726 8508
rect 6680 8477 6714 8488
rect 6715 8477 6726 8493
rect 6772 8484 6788 8500
rect 6795 8498 6825 8550
rect 6859 8546 6860 8553
rect 6844 8538 6860 8546
rect 6831 8506 6844 8525
rect 6859 8506 6889 8522
rect 6831 8490 6905 8506
rect 6831 8488 6844 8490
rect 6859 8488 6893 8490
rect 6496 8466 6509 8468
rect 6524 8466 6558 8468
rect 6496 8450 6558 8466
rect 6602 8461 6618 8464
rect 6680 8461 6710 8472
rect 6758 8468 6804 8484
rect 6831 8472 6905 8488
rect 6758 8466 6792 8468
rect 6757 8450 6804 8466
rect 6831 8450 6844 8472
rect 6859 8450 6889 8472
rect 6916 8450 6917 8466
rect 6932 8450 6945 8610
rect 6975 8506 6988 8610
rect 7033 8588 7034 8598
rect 7049 8588 7062 8598
rect 7033 8584 7062 8588
rect 7067 8584 7097 8610
rect 7115 8596 7131 8598
rect 7203 8596 7256 8610
rect 7204 8594 7268 8596
rect 7311 8594 7326 8610
rect 7375 8607 7405 8610
rect 7375 8604 7411 8607
rect 7341 8596 7357 8598
rect 7115 8584 7130 8588
rect 7033 8582 7130 8584
rect 7158 8582 7326 8594
rect 7342 8584 7357 8588
rect 7375 8585 7414 8604
rect 7433 8598 7440 8599
rect 7439 8591 7440 8598
rect 7423 8588 7424 8591
rect 7439 8588 7452 8591
rect 7375 8584 7405 8585
rect 7414 8584 7420 8585
rect 7423 8584 7452 8588
rect 7342 8583 7452 8584
rect 7342 8582 7458 8583
rect 7017 8574 7068 8582
rect 7017 8562 7042 8574
rect 7049 8562 7068 8574
rect 7099 8574 7149 8582
rect 7099 8566 7115 8574
rect 7122 8572 7149 8574
rect 7158 8572 7379 8582
rect 7122 8562 7379 8572
rect 7408 8574 7458 8582
rect 7408 8565 7424 8574
rect 7017 8554 7068 8562
rect 7115 8554 7379 8562
rect 7405 8562 7424 8565
rect 7431 8562 7458 8574
rect 7405 8554 7458 8562
rect 7033 8546 7034 8554
rect 7049 8546 7062 8554
rect 7033 8538 7049 8546
rect 7030 8531 7049 8534
rect 7030 8522 7052 8531
rect 7003 8512 7052 8522
rect 7003 8506 7033 8512
rect 7052 8507 7057 8512
rect 6975 8490 7049 8506
rect 7067 8498 7097 8554
rect 7132 8544 7340 8554
rect 7375 8550 7420 8554
rect 7423 8553 7424 8554
rect 7439 8553 7452 8554
rect 7158 8514 7347 8544
rect 7173 8511 7347 8514
rect 7166 8508 7347 8511
rect 6975 8488 6988 8490
rect 7003 8488 7037 8490
rect 6975 8472 7049 8488
rect 7076 8484 7089 8498
rect 7104 8484 7120 8500
rect 7166 8495 7177 8508
rect 6959 8450 6960 8466
rect 6975 8450 6988 8472
rect 7003 8450 7033 8472
rect 7076 8468 7138 8484
rect 7166 8477 7177 8493
rect 7182 8488 7192 8508
rect 7202 8488 7216 8508
rect 7219 8495 7228 8508
rect 7244 8495 7253 8508
rect 7182 8477 7216 8488
rect 7219 8477 7228 8493
rect 7244 8477 7253 8493
rect 7260 8488 7270 8508
rect 7280 8488 7294 8508
rect 7295 8495 7306 8508
rect 7260 8477 7294 8488
rect 7295 8477 7306 8493
rect 7352 8484 7368 8500
rect 7375 8498 7405 8550
rect 7439 8546 7440 8553
rect 7424 8538 7440 8546
rect 7411 8506 7424 8525
rect 7439 8506 7469 8522
rect 7411 8490 7485 8506
rect 7411 8488 7424 8490
rect 7439 8488 7473 8490
rect 7076 8466 7089 8468
rect 7104 8466 7138 8468
rect 7076 8450 7138 8466
rect 7182 8461 7198 8464
rect 7260 8461 7290 8472
rect 7338 8468 7384 8484
rect 7411 8472 7485 8488
rect 7338 8466 7372 8468
rect 7337 8450 7384 8466
rect 7411 8450 7424 8472
rect 7439 8450 7469 8472
rect 7496 8450 7497 8466
rect 7512 8450 7525 8610
rect 7555 8506 7568 8610
rect 7613 8588 7614 8598
rect 7629 8588 7642 8598
rect 7613 8584 7642 8588
rect 7647 8584 7677 8610
rect 7695 8596 7711 8598
rect 7783 8596 7836 8610
rect 7784 8594 7848 8596
rect 7891 8594 7906 8610
rect 7955 8607 7985 8610
rect 7955 8604 7991 8607
rect 7921 8596 7937 8598
rect 7695 8584 7710 8588
rect 7613 8582 7710 8584
rect 7738 8582 7906 8594
rect 7922 8584 7937 8588
rect 7955 8585 7994 8604
rect 8013 8598 8020 8599
rect 8019 8591 8020 8598
rect 8003 8588 8004 8591
rect 8019 8588 8032 8591
rect 7955 8584 7985 8585
rect 7994 8584 8000 8585
rect 8003 8584 8032 8588
rect 7922 8583 8032 8584
rect 7922 8582 8038 8583
rect 7597 8574 7648 8582
rect 7597 8562 7622 8574
rect 7629 8562 7648 8574
rect 7679 8574 7729 8582
rect 7679 8566 7695 8574
rect 7702 8572 7729 8574
rect 7738 8572 7959 8582
rect 7702 8562 7959 8572
rect 7988 8574 8038 8582
rect 7988 8565 8004 8574
rect 7597 8554 7648 8562
rect 7695 8554 7959 8562
rect 7985 8562 8004 8565
rect 8011 8562 8038 8574
rect 7985 8554 8038 8562
rect 7613 8546 7614 8554
rect 7629 8546 7642 8554
rect 7613 8538 7629 8546
rect 7610 8531 7629 8534
rect 7610 8522 7632 8531
rect 7583 8512 7632 8522
rect 7583 8506 7613 8512
rect 7632 8507 7637 8512
rect 7555 8490 7629 8506
rect 7647 8498 7677 8554
rect 7712 8544 7920 8554
rect 7955 8550 8000 8554
rect 8003 8553 8004 8554
rect 8019 8553 8032 8554
rect 7738 8514 7927 8544
rect 7753 8511 7927 8514
rect 7746 8508 7927 8511
rect 7555 8488 7568 8490
rect 7583 8488 7617 8490
rect 7555 8472 7629 8488
rect 7656 8484 7669 8498
rect 7684 8484 7700 8500
rect 7746 8495 7757 8508
rect 7539 8450 7540 8466
rect 7555 8450 7568 8472
rect 7583 8450 7613 8472
rect 7656 8468 7718 8484
rect 7746 8477 7757 8493
rect 7762 8488 7772 8508
rect 7782 8488 7796 8508
rect 7799 8495 7808 8508
rect 7824 8495 7833 8508
rect 7762 8477 7796 8488
rect 7799 8477 7808 8493
rect 7824 8477 7833 8493
rect 7840 8488 7850 8508
rect 7860 8488 7874 8508
rect 7875 8495 7886 8508
rect 7840 8477 7874 8488
rect 7875 8477 7886 8493
rect 7932 8484 7948 8500
rect 7955 8498 7985 8550
rect 8019 8546 8020 8553
rect 8004 8538 8020 8546
rect 7991 8506 8004 8525
rect 8019 8506 8049 8522
rect 7991 8490 8065 8506
rect 7991 8488 8004 8490
rect 8019 8488 8053 8490
rect 7656 8466 7669 8468
rect 7684 8466 7718 8468
rect 7656 8450 7718 8466
rect 7762 8461 7778 8464
rect 7840 8461 7870 8472
rect 7918 8468 7964 8484
rect 7991 8472 8065 8488
rect 7918 8466 7952 8468
rect 7917 8450 7964 8466
rect 7991 8450 8004 8472
rect 8019 8450 8049 8472
rect 8076 8450 8077 8466
rect 8092 8450 8105 8610
rect 8135 8506 8148 8610
rect 8193 8588 8194 8598
rect 8209 8588 8222 8598
rect 8193 8584 8222 8588
rect 8227 8584 8257 8610
rect 8275 8596 8291 8598
rect 8363 8596 8416 8610
rect 8364 8594 8428 8596
rect 8471 8594 8486 8610
rect 8535 8607 8565 8610
rect 8535 8604 8571 8607
rect 8501 8596 8517 8598
rect 8275 8584 8290 8588
rect 8193 8582 8290 8584
rect 8318 8582 8486 8594
rect 8502 8584 8517 8588
rect 8535 8585 8574 8604
rect 8593 8598 8600 8599
rect 8599 8591 8600 8598
rect 8583 8588 8584 8591
rect 8599 8588 8612 8591
rect 8535 8584 8565 8585
rect 8574 8584 8580 8585
rect 8583 8584 8612 8588
rect 8502 8583 8612 8584
rect 8502 8582 8618 8583
rect 8177 8574 8228 8582
rect 8177 8562 8202 8574
rect 8209 8562 8228 8574
rect 8259 8574 8309 8582
rect 8259 8566 8275 8574
rect 8282 8572 8309 8574
rect 8318 8572 8539 8582
rect 8282 8562 8539 8572
rect 8568 8574 8618 8582
rect 8568 8565 8584 8574
rect 8177 8554 8228 8562
rect 8275 8554 8539 8562
rect 8565 8562 8584 8565
rect 8591 8562 8618 8574
rect 8565 8554 8618 8562
rect 8193 8546 8194 8554
rect 8209 8546 8222 8554
rect 8193 8538 8209 8546
rect 8190 8531 8209 8534
rect 8190 8522 8212 8531
rect 8163 8512 8212 8522
rect 8163 8506 8193 8512
rect 8212 8507 8217 8512
rect 8135 8490 8209 8506
rect 8227 8498 8257 8554
rect 8292 8544 8500 8554
rect 8535 8550 8580 8554
rect 8583 8553 8584 8554
rect 8599 8553 8612 8554
rect 8318 8514 8507 8544
rect 8333 8511 8507 8514
rect 8326 8508 8507 8511
rect 8135 8488 8148 8490
rect 8163 8488 8197 8490
rect 8135 8472 8209 8488
rect 8236 8484 8249 8498
rect 8264 8484 8280 8500
rect 8326 8495 8337 8508
rect 8119 8450 8120 8466
rect 8135 8450 8148 8472
rect 8163 8450 8193 8472
rect 8236 8468 8298 8484
rect 8326 8477 8337 8493
rect 8342 8488 8352 8508
rect 8362 8488 8376 8508
rect 8379 8495 8388 8508
rect 8404 8495 8413 8508
rect 8342 8477 8376 8488
rect 8379 8477 8388 8493
rect 8404 8477 8413 8493
rect 8420 8488 8430 8508
rect 8440 8488 8454 8508
rect 8455 8495 8466 8508
rect 8420 8477 8454 8488
rect 8455 8477 8466 8493
rect 8512 8484 8528 8500
rect 8535 8498 8565 8550
rect 8599 8546 8600 8553
rect 8584 8538 8600 8546
rect 8571 8506 8584 8525
rect 8599 8506 8629 8522
rect 8571 8490 8645 8506
rect 8571 8488 8584 8490
rect 8599 8488 8633 8490
rect 8236 8466 8249 8468
rect 8264 8466 8298 8468
rect 8236 8450 8298 8466
rect 8342 8461 8358 8464
rect 8420 8461 8450 8472
rect 8498 8468 8544 8484
rect 8571 8472 8645 8488
rect 8498 8466 8532 8468
rect 8497 8450 8544 8466
rect 8571 8450 8584 8472
rect 8599 8450 8629 8472
rect 8656 8450 8657 8466
rect 8672 8450 8685 8610
rect 8715 8506 8728 8610
rect 8773 8588 8774 8598
rect 8789 8588 8802 8598
rect 8773 8584 8802 8588
rect 8807 8584 8837 8610
rect 8855 8596 8871 8598
rect 8943 8596 8996 8610
rect 8944 8594 9008 8596
rect 9051 8594 9066 8610
rect 9115 8607 9145 8610
rect 9115 8604 9151 8607
rect 9081 8596 9097 8598
rect 8855 8584 8870 8588
rect 8773 8582 8870 8584
rect 8898 8582 9066 8594
rect 9082 8584 9097 8588
rect 9115 8585 9154 8604
rect 9173 8598 9180 8599
rect 9179 8591 9180 8598
rect 9163 8588 9164 8591
rect 9179 8588 9192 8591
rect 9115 8584 9145 8585
rect 9154 8584 9160 8585
rect 9163 8584 9192 8588
rect 9082 8583 9192 8584
rect 9082 8582 9198 8583
rect 8757 8574 8808 8582
rect 8757 8562 8782 8574
rect 8789 8562 8808 8574
rect 8839 8574 8889 8582
rect 8839 8566 8855 8574
rect 8862 8572 8889 8574
rect 8898 8572 9119 8582
rect 8862 8562 9119 8572
rect 9148 8574 9198 8582
rect 9148 8565 9164 8574
rect 8757 8554 8808 8562
rect 8855 8554 9119 8562
rect 9145 8562 9164 8565
rect 9171 8562 9198 8574
rect 9145 8554 9198 8562
rect 8773 8546 8774 8554
rect 8789 8546 8802 8554
rect 8773 8538 8789 8546
rect 8770 8531 8789 8534
rect 8770 8522 8792 8531
rect 8743 8512 8792 8522
rect 8743 8506 8773 8512
rect 8792 8507 8797 8512
rect 8715 8490 8789 8506
rect 8807 8498 8837 8554
rect 8872 8544 9080 8554
rect 9115 8550 9160 8554
rect 9163 8553 9164 8554
rect 9179 8553 9192 8554
rect 8898 8514 9087 8544
rect 8913 8511 9087 8514
rect 8906 8508 9087 8511
rect 8715 8488 8728 8490
rect 8743 8488 8777 8490
rect 8715 8472 8789 8488
rect 8816 8484 8829 8498
rect 8844 8484 8860 8500
rect 8906 8495 8917 8508
rect 8699 8450 8700 8466
rect 8715 8450 8728 8472
rect 8743 8450 8773 8472
rect 8816 8468 8878 8484
rect 8906 8477 8917 8493
rect 8922 8488 8932 8508
rect 8942 8488 8956 8508
rect 8959 8495 8968 8508
rect 8984 8495 8993 8508
rect 8922 8477 8956 8488
rect 8959 8477 8968 8493
rect 8984 8477 8993 8493
rect 9000 8488 9010 8508
rect 9020 8488 9034 8508
rect 9035 8495 9046 8508
rect 9000 8477 9034 8488
rect 9035 8477 9046 8493
rect 9092 8484 9108 8500
rect 9115 8498 9145 8550
rect 9179 8546 9180 8553
rect 9164 8538 9180 8546
rect 9151 8506 9164 8525
rect 9179 8506 9209 8522
rect 9151 8490 9225 8506
rect 9151 8488 9164 8490
rect 9179 8488 9213 8490
rect 8816 8466 8829 8468
rect 8844 8466 8878 8468
rect 8816 8450 8878 8466
rect 8922 8461 8938 8464
rect 9000 8461 9030 8472
rect 9078 8468 9124 8484
rect 9151 8472 9225 8488
rect 9078 8466 9112 8468
rect 9077 8450 9124 8466
rect 9151 8450 9164 8472
rect 9179 8450 9209 8472
rect 9236 8450 9237 8466
rect 9252 8450 9265 8610
rect -7 8442 34 8450
rect -7 8416 8 8442
rect 15 8416 34 8442
rect 98 8438 160 8450
rect 172 8438 247 8450
rect 305 8438 380 8450
rect 392 8438 423 8450
rect 429 8438 464 8450
rect 98 8436 260 8438
rect -7 8408 34 8416
rect 116 8412 129 8436
rect 144 8434 159 8436
rect -1 8398 0 8408
rect 15 8398 28 8408
rect 43 8398 73 8412
rect 116 8398 159 8412
rect 183 8409 190 8416
rect 193 8412 260 8436
rect 292 8436 464 8438
rect 262 8414 290 8418
rect 292 8414 372 8436
rect 393 8434 408 8436
rect 262 8412 372 8414
rect 193 8408 372 8412
rect 166 8398 196 8408
rect 198 8398 351 8408
rect 359 8398 389 8408
rect 393 8398 423 8412
rect 451 8398 464 8436
rect 536 8442 571 8450
rect 536 8416 537 8442
rect 544 8416 571 8442
rect 479 8398 509 8412
rect 536 8408 571 8416
rect 573 8442 614 8450
rect 573 8416 588 8442
rect 595 8416 614 8442
rect 678 8438 740 8450
rect 752 8438 827 8450
rect 885 8438 960 8450
rect 972 8438 1003 8450
rect 1009 8438 1044 8450
rect 678 8436 840 8438
rect 573 8408 614 8416
rect 696 8412 709 8436
rect 724 8434 739 8436
rect 536 8398 537 8408
rect 552 8398 565 8408
rect 579 8398 580 8408
rect 595 8398 608 8408
rect 623 8398 653 8412
rect 696 8398 739 8412
rect 763 8409 770 8416
rect 773 8412 840 8436
rect 872 8436 1044 8438
rect 842 8414 870 8418
rect 872 8414 952 8436
rect 973 8434 988 8436
rect 842 8412 952 8414
rect 773 8408 952 8412
rect 746 8398 776 8408
rect 778 8398 931 8408
rect 939 8398 969 8408
rect 973 8398 1003 8412
rect 1031 8398 1044 8436
rect 1116 8442 1151 8450
rect 1116 8416 1117 8442
rect 1124 8416 1151 8442
rect 1059 8398 1089 8412
rect 1116 8408 1151 8416
rect 1153 8442 1194 8450
rect 1153 8416 1168 8442
rect 1175 8416 1194 8442
rect 1258 8438 1320 8450
rect 1332 8438 1407 8450
rect 1465 8438 1540 8450
rect 1552 8438 1583 8450
rect 1589 8438 1624 8450
rect 1258 8436 1420 8438
rect 1153 8408 1194 8416
rect 1276 8412 1289 8436
rect 1304 8434 1319 8436
rect 1116 8398 1117 8408
rect 1132 8398 1145 8408
rect 1159 8398 1160 8408
rect 1175 8398 1188 8408
rect 1203 8398 1233 8412
rect 1276 8398 1319 8412
rect 1343 8409 1350 8416
rect 1353 8412 1420 8436
rect 1452 8436 1624 8438
rect 1422 8414 1450 8418
rect 1452 8414 1532 8436
rect 1553 8434 1568 8436
rect 1422 8412 1532 8414
rect 1353 8408 1532 8412
rect 1326 8398 1356 8408
rect 1358 8398 1511 8408
rect 1519 8398 1549 8408
rect 1553 8398 1583 8412
rect 1611 8398 1624 8436
rect 1696 8442 1731 8450
rect 1696 8416 1697 8442
rect 1704 8416 1731 8442
rect 1639 8398 1669 8412
rect 1696 8408 1731 8416
rect 1733 8442 1774 8450
rect 1733 8416 1748 8442
rect 1755 8416 1774 8442
rect 1838 8438 1900 8450
rect 1912 8438 1987 8450
rect 2045 8438 2120 8450
rect 2132 8438 2163 8450
rect 2169 8438 2204 8450
rect 1838 8436 2000 8438
rect 1733 8408 1774 8416
rect 1856 8412 1869 8436
rect 1884 8434 1899 8436
rect 1696 8398 1697 8408
rect 1712 8398 1725 8408
rect 1739 8398 1740 8408
rect 1755 8398 1768 8408
rect 1783 8398 1813 8412
rect 1856 8398 1899 8412
rect 1923 8409 1930 8416
rect 1933 8412 2000 8436
rect 2032 8436 2204 8438
rect 2002 8414 2030 8418
rect 2032 8414 2112 8436
rect 2133 8434 2148 8436
rect 2002 8412 2112 8414
rect 1933 8408 2112 8412
rect 1906 8398 1936 8408
rect 1938 8398 2091 8408
rect 2099 8398 2129 8408
rect 2133 8398 2163 8412
rect 2191 8398 2204 8436
rect 2276 8442 2311 8450
rect 2276 8416 2277 8442
rect 2284 8416 2311 8442
rect 2219 8398 2249 8412
rect 2276 8408 2311 8416
rect 2313 8442 2354 8450
rect 2313 8416 2328 8442
rect 2335 8416 2354 8442
rect 2418 8438 2480 8450
rect 2492 8438 2567 8450
rect 2625 8438 2700 8450
rect 2712 8438 2743 8450
rect 2749 8438 2784 8450
rect 2418 8436 2580 8438
rect 2313 8408 2354 8416
rect 2436 8412 2449 8436
rect 2464 8434 2479 8436
rect 2276 8398 2277 8408
rect 2292 8398 2305 8408
rect 2319 8398 2320 8408
rect 2335 8398 2348 8408
rect 2363 8398 2393 8412
rect 2436 8398 2479 8412
rect 2503 8409 2510 8416
rect 2513 8412 2580 8436
rect 2612 8436 2784 8438
rect 2582 8414 2610 8418
rect 2612 8414 2692 8436
rect 2713 8434 2728 8436
rect 2582 8412 2692 8414
rect 2513 8408 2692 8412
rect 2486 8398 2516 8408
rect 2518 8398 2671 8408
rect 2679 8398 2709 8408
rect 2713 8398 2743 8412
rect 2771 8398 2784 8436
rect 2856 8442 2891 8450
rect 2856 8416 2857 8442
rect 2864 8416 2891 8442
rect 2799 8398 2829 8412
rect 2856 8408 2891 8416
rect 2893 8442 2934 8450
rect 2893 8416 2908 8442
rect 2915 8416 2934 8442
rect 2998 8438 3060 8450
rect 3072 8438 3147 8450
rect 3205 8438 3280 8450
rect 3292 8438 3323 8450
rect 3329 8438 3364 8450
rect 2998 8436 3160 8438
rect 2893 8408 2934 8416
rect 3016 8412 3029 8436
rect 3044 8434 3059 8436
rect 2856 8398 2857 8408
rect 2872 8398 2885 8408
rect 2899 8398 2900 8408
rect 2915 8398 2928 8408
rect 2943 8398 2973 8412
rect 3016 8398 3059 8412
rect 3083 8409 3090 8416
rect 3093 8412 3160 8436
rect 3192 8436 3364 8438
rect 3162 8414 3190 8418
rect 3192 8414 3272 8436
rect 3293 8434 3308 8436
rect 3162 8412 3272 8414
rect 3093 8408 3272 8412
rect 3066 8398 3096 8408
rect 3098 8398 3251 8408
rect 3259 8398 3289 8408
rect 3293 8398 3323 8412
rect 3351 8398 3364 8436
rect 3436 8442 3471 8450
rect 3436 8416 3437 8442
rect 3444 8416 3471 8442
rect 3379 8398 3409 8412
rect 3436 8408 3471 8416
rect 3473 8442 3514 8450
rect 3473 8416 3488 8442
rect 3495 8416 3514 8442
rect 3578 8438 3640 8450
rect 3652 8438 3727 8450
rect 3785 8438 3860 8450
rect 3872 8438 3903 8450
rect 3909 8438 3944 8450
rect 3578 8436 3740 8438
rect 3473 8408 3514 8416
rect 3596 8412 3609 8436
rect 3624 8434 3639 8436
rect 3436 8398 3437 8408
rect 3452 8398 3465 8408
rect 3479 8398 3480 8408
rect 3495 8398 3508 8408
rect 3523 8398 3553 8412
rect 3596 8398 3639 8412
rect 3663 8409 3670 8416
rect 3673 8412 3740 8436
rect 3772 8436 3944 8438
rect 3742 8414 3770 8418
rect 3772 8414 3852 8436
rect 3873 8434 3888 8436
rect 3742 8412 3852 8414
rect 3673 8408 3852 8412
rect 3646 8398 3676 8408
rect 3678 8398 3831 8408
rect 3839 8398 3869 8408
rect 3873 8398 3903 8412
rect 3931 8398 3944 8436
rect 4016 8442 4051 8450
rect 4016 8416 4017 8442
rect 4024 8416 4051 8442
rect 3959 8398 3989 8412
rect 4016 8408 4051 8416
rect 4053 8442 4094 8450
rect 4053 8416 4068 8442
rect 4075 8416 4094 8442
rect 4158 8438 4220 8450
rect 4232 8438 4307 8450
rect 4365 8438 4440 8450
rect 4452 8438 4483 8450
rect 4489 8438 4524 8450
rect 4158 8436 4320 8438
rect 4053 8408 4094 8416
rect 4176 8412 4189 8436
rect 4204 8434 4219 8436
rect 4016 8398 4017 8408
rect 4032 8398 4045 8408
rect 4059 8398 4060 8408
rect 4075 8398 4088 8408
rect 4103 8398 4133 8412
rect 4176 8398 4219 8412
rect 4243 8409 4250 8416
rect 4253 8412 4320 8436
rect 4352 8436 4524 8438
rect 4322 8414 4350 8418
rect 4352 8414 4432 8436
rect 4453 8434 4468 8436
rect 4322 8412 4432 8414
rect 4253 8408 4432 8412
rect 4226 8398 4256 8408
rect 4258 8398 4411 8408
rect 4419 8398 4449 8408
rect 4453 8398 4483 8412
rect 4511 8398 4524 8436
rect 4596 8442 4631 8450
rect 4596 8416 4597 8442
rect 4604 8416 4631 8442
rect 4539 8398 4569 8412
rect 4596 8408 4631 8416
rect 4633 8442 4674 8450
rect 4633 8416 4648 8442
rect 4655 8416 4674 8442
rect 4738 8438 4800 8450
rect 4812 8438 4887 8450
rect 4945 8438 5020 8450
rect 5032 8438 5063 8450
rect 5069 8438 5104 8450
rect 4738 8436 4900 8438
rect 4633 8408 4674 8416
rect 4756 8412 4769 8436
rect 4784 8434 4799 8436
rect 4596 8398 4597 8408
rect 4612 8398 4625 8408
rect 4639 8398 4640 8408
rect 4655 8398 4668 8408
rect 4683 8398 4713 8412
rect 4756 8398 4799 8412
rect 4823 8409 4830 8416
rect 4833 8412 4900 8436
rect 4932 8436 5104 8438
rect 4902 8414 4930 8418
rect 4932 8414 5012 8436
rect 5033 8434 5048 8436
rect 4902 8412 5012 8414
rect 4833 8408 5012 8412
rect 4806 8398 4836 8408
rect 4838 8398 4991 8408
rect 4999 8398 5029 8408
rect 5033 8398 5063 8412
rect 5091 8398 5104 8436
rect 5176 8442 5211 8450
rect 5176 8416 5177 8442
rect 5184 8416 5211 8442
rect 5119 8398 5149 8412
rect 5176 8408 5211 8416
rect 5213 8442 5254 8450
rect 5213 8416 5228 8442
rect 5235 8416 5254 8442
rect 5318 8438 5380 8450
rect 5392 8438 5467 8450
rect 5525 8438 5600 8450
rect 5612 8438 5643 8450
rect 5649 8438 5684 8450
rect 5318 8436 5480 8438
rect 5213 8408 5254 8416
rect 5336 8412 5349 8436
rect 5364 8434 5379 8436
rect 5176 8398 5177 8408
rect 5192 8398 5205 8408
rect 5219 8398 5220 8408
rect 5235 8398 5248 8408
rect 5263 8398 5293 8412
rect 5336 8398 5379 8412
rect 5403 8409 5410 8416
rect 5413 8412 5480 8436
rect 5512 8436 5684 8438
rect 5482 8414 5510 8418
rect 5512 8414 5592 8436
rect 5613 8434 5628 8436
rect 5482 8412 5592 8414
rect 5413 8408 5592 8412
rect 5386 8398 5416 8408
rect 5418 8398 5571 8408
rect 5579 8398 5609 8408
rect 5613 8398 5643 8412
rect 5671 8398 5684 8436
rect 5756 8442 5791 8450
rect 5756 8416 5757 8442
rect 5764 8416 5791 8442
rect 5699 8398 5729 8412
rect 5756 8408 5791 8416
rect 5793 8442 5834 8450
rect 5793 8416 5808 8442
rect 5815 8416 5834 8442
rect 5898 8438 5960 8450
rect 5972 8438 6047 8450
rect 6105 8438 6180 8450
rect 6192 8438 6223 8450
rect 6229 8438 6264 8450
rect 5898 8436 6060 8438
rect 5793 8408 5834 8416
rect 5916 8412 5929 8436
rect 5944 8434 5959 8436
rect 5756 8398 5757 8408
rect 5772 8398 5785 8408
rect 5799 8398 5800 8408
rect 5815 8398 5828 8408
rect 5843 8398 5873 8412
rect 5916 8398 5959 8412
rect 5983 8409 5990 8416
rect 5993 8412 6060 8436
rect 6092 8436 6264 8438
rect 6062 8414 6090 8418
rect 6092 8414 6172 8436
rect 6193 8434 6208 8436
rect 6062 8412 6172 8414
rect 5993 8408 6172 8412
rect 5966 8398 5996 8408
rect 5998 8398 6151 8408
rect 6159 8398 6189 8408
rect 6193 8398 6223 8412
rect 6251 8398 6264 8436
rect 6336 8442 6371 8450
rect 6336 8416 6337 8442
rect 6344 8416 6371 8442
rect 6279 8398 6309 8412
rect 6336 8408 6371 8416
rect 6373 8442 6414 8450
rect 6373 8416 6388 8442
rect 6395 8416 6414 8442
rect 6478 8438 6540 8450
rect 6552 8438 6627 8450
rect 6685 8438 6760 8450
rect 6772 8438 6803 8450
rect 6809 8438 6844 8450
rect 6478 8436 6640 8438
rect 6373 8408 6414 8416
rect 6496 8412 6509 8436
rect 6524 8434 6539 8436
rect 6336 8398 6337 8408
rect 6352 8398 6365 8408
rect 6379 8398 6380 8408
rect 6395 8398 6408 8408
rect 6423 8398 6453 8412
rect 6496 8398 6539 8412
rect 6563 8409 6570 8416
rect 6573 8412 6640 8436
rect 6672 8436 6844 8438
rect 6642 8414 6670 8418
rect 6672 8414 6752 8436
rect 6773 8434 6788 8436
rect 6642 8412 6752 8414
rect 6573 8408 6752 8412
rect 6546 8398 6576 8408
rect 6578 8398 6731 8408
rect 6739 8398 6769 8408
rect 6773 8398 6803 8412
rect 6831 8398 6844 8436
rect 6916 8442 6951 8450
rect 6916 8416 6917 8442
rect 6924 8416 6951 8442
rect 6859 8398 6889 8412
rect 6916 8408 6951 8416
rect 6953 8442 6994 8450
rect 6953 8416 6968 8442
rect 6975 8416 6994 8442
rect 7058 8438 7120 8450
rect 7132 8438 7207 8450
rect 7265 8438 7340 8450
rect 7352 8438 7383 8450
rect 7389 8438 7424 8450
rect 7058 8436 7220 8438
rect 6953 8408 6994 8416
rect 7076 8412 7089 8436
rect 7104 8434 7119 8436
rect 6916 8398 6917 8408
rect 6932 8398 6945 8408
rect 6959 8398 6960 8408
rect 6975 8398 6988 8408
rect 7003 8398 7033 8412
rect 7076 8398 7119 8412
rect 7143 8409 7150 8416
rect 7153 8412 7220 8436
rect 7252 8436 7424 8438
rect 7222 8414 7250 8418
rect 7252 8414 7332 8436
rect 7353 8434 7368 8436
rect 7222 8412 7332 8414
rect 7153 8408 7332 8412
rect 7126 8398 7156 8408
rect 7158 8398 7311 8408
rect 7319 8398 7349 8408
rect 7353 8398 7383 8412
rect 7411 8398 7424 8436
rect 7496 8442 7531 8450
rect 7496 8416 7497 8442
rect 7504 8416 7531 8442
rect 7439 8398 7469 8412
rect 7496 8408 7531 8416
rect 7533 8442 7574 8450
rect 7533 8416 7548 8442
rect 7555 8416 7574 8442
rect 7638 8438 7700 8450
rect 7712 8438 7787 8450
rect 7845 8438 7920 8450
rect 7932 8438 7963 8450
rect 7969 8438 8004 8450
rect 7638 8436 7800 8438
rect 7533 8408 7574 8416
rect 7656 8412 7669 8436
rect 7684 8434 7699 8436
rect 7496 8398 7497 8408
rect 7512 8398 7525 8408
rect 7539 8398 7540 8408
rect 7555 8398 7568 8408
rect 7583 8398 7613 8412
rect 7656 8398 7699 8412
rect 7723 8409 7730 8416
rect 7733 8412 7800 8436
rect 7832 8436 8004 8438
rect 7802 8414 7830 8418
rect 7832 8414 7912 8436
rect 7933 8434 7948 8436
rect 7802 8412 7912 8414
rect 7733 8408 7912 8412
rect 7706 8398 7736 8408
rect 7738 8398 7891 8408
rect 7899 8398 7929 8408
rect 7933 8398 7963 8412
rect 7991 8398 8004 8436
rect 8076 8442 8111 8450
rect 8076 8416 8077 8442
rect 8084 8416 8111 8442
rect 8019 8398 8049 8412
rect 8076 8408 8111 8416
rect 8113 8442 8154 8450
rect 8113 8416 8128 8442
rect 8135 8416 8154 8442
rect 8218 8438 8280 8450
rect 8292 8438 8367 8450
rect 8425 8438 8500 8450
rect 8512 8438 8543 8450
rect 8549 8438 8584 8450
rect 8218 8436 8380 8438
rect 8113 8408 8154 8416
rect 8236 8412 8249 8436
rect 8264 8434 8279 8436
rect 8076 8398 8077 8408
rect 8092 8398 8105 8408
rect 8119 8398 8120 8408
rect 8135 8398 8148 8408
rect 8163 8398 8193 8412
rect 8236 8398 8279 8412
rect 8303 8409 8310 8416
rect 8313 8412 8380 8436
rect 8412 8436 8584 8438
rect 8382 8414 8410 8418
rect 8412 8414 8492 8436
rect 8513 8434 8528 8436
rect 8382 8412 8492 8414
rect 8313 8408 8492 8412
rect 8286 8398 8316 8408
rect 8318 8398 8471 8408
rect 8479 8398 8509 8408
rect 8513 8398 8543 8412
rect 8571 8398 8584 8436
rect 8656 8442 8691 8450
rect 8656 8416 8657 8442
rect 8664 8416 8691 8442
rect 8599 8398 8629 8412
rect 8656 8408 8691 8416
rect 8693 8442 8734 8450
rect 8693 8416 8708 8442
rect 8715 8416 8734 8442
rect 8798 8438 8860 8450
rect 8872 8438 8947 8450
rect 9005 8438 9080 8450
rect 9092 8438 9123 8450
rect 9129 8438 9164 8450
rect 8798 8436 8960 8438
rect 8693 8408 8734 8416
rect 8816 8412 8829 8436
rect 8844 8434 8859 8436
rect 8656 8398 8657 8408
rect 8672 8398 8685 8408
rect 8699 8398 8700 8408
rect 8715 8398 8728 8408
rect 8743 8398 8773 8412
rect 8816 8398 8859 8412
rect 8883 8409 8890 8416
rect 8893 8412 8960 8436
rect 8992 8436 9164 8438
rect 8962 8414 8990 8418
rect 8992 8414 9072 8436
rect 9093 8434 9108 8436
rect 8962 8412 9072 8414
rect 8893 8408 9072 8412
rect 8866 8398 8896 8408
rect 8898 8398 9051 8408
rect 9059 8398 9089 8408
rect 9093 8398 9123 8412
rect 9151 8398 9164 8436
rect 9236 8442 9271 8450
rect 9236 8416 9237 8442
rect 9244 8416 9271 8442
rect 9179 8398 9209 8412
rect 9236 8408 9271 8416
rect 9236 8398 9237 8408
rect 9252 8398 9265 8408
rect -1 8392 9265 8398
rect 0 8384 9265 8392
rect 15 8354 28 8384
rect 43 8366 73 8384
rect 116 8370 130 8384
rect 166 8370 386 8384
rect 117 8368 130 8370
rect 83 8356 98 8368
rect 80 8354 102 8356
rect 107 8354 137 8368
rect 198 8366 351 8370
rect 180 8354 372 8366
rect 415 8354 445 8368
rect 451 8354 464 8384
rect 479 8366 509 8384
rect 552 8354 565 8384
rect 595 8354 608 8384
rect 623 8366 653 8384
rect 696 8370 710 8384
rect 746 8370 966 8384
rect 697 8368 710 8370
rect 663 8356 678 8368
rect 660 8354 682 8356
rect 687 8354 717 8368
rect 778 8366 931 8370
rect 760 8354 952 8366
rect 995 8354 1025 8368
rect 1031 8354 1044 8384
rect 1059 8366 1089 8384
rect 1132 8354 1145 8384
rect 1175 8354 1188 8384
rect 1203 8366 1233 8384
rect 1276 8370 1290 8384
rect 1326 8370 1546 8384
rect 1277 8368 1290 8370
rect 1243 8356 1258 8368
rect 1240 8354 1262 8356
rect 1267 8354 1297 8368
rect 1358 8366 1511 8370
rect 1340 8354 1532 8366
rect 1575 8354 1605 8368
rect 1611 8354 1624 8384
rect 1639 8366 1669 8384
rect 1712 8354 1725 8384
rect 1755 8354 1768 8384
rect 1783 8366 1813 8384
rect 1856 8370 1870 8384
rect 1906 8370 2126 8384
rect 1857 8368 1870 8370
rect 1823 8356 1838 8368
rect 1820 8354 1842 8356
rect 1847 8354 1877 8368
rect 1938 8366 2091 8370
rect 1920 8354 2112 8366
rect 2155 8354 2185 8368
rect 2191 8354 2204 8384
rect 2219 8366 2249 8384
rect 2292 8354 2305 8384
rect 2335 8354 2348 8384
rect 2363 8366 2393 8384
rect 2436 8370 2450 8384
rect 2486 8370 2706 8384
rect 2437 8368 2450 8370
rect 2403 8356 2418 8368
rect 2400 8354 2422 8356
rect 2427 8354 2457 8368
rect 2518 8366 2671 8370
rect 2500 8354 2692 8366
rect 2735 8354 2765 8368
rect 2771 8354 2784 8384
rect 2799 8366 2829 8384
rect 2872 8354 2885 8384
rect 2915 8354 2928 8384
rect 2943 8366 2973 8384
rect 3016 8370 3030 8384
rect 3066 8370 3286 8384
rect 3017 8368 3030 8370
rect 2983 8356 2998 8368
rect 2980 8354 3002 8356
rect 3007 8354 3037 8368
rect 3098 8366 3251 8370
rect 3080 8354 3272 8366
rect 3315 8354 3345 8368
rect 3351 8354 3364 8384
rect 3379 8366 3409 8384
rect 3452 8354 3465 8384
rect 3495 8354 3508 8384
rect 3523 8366 3553 8384
rect 3596 8370 3610 8384
rect 3646 8370 3866 8384
rect 3597 8368 3610 8370
rect 3563 8356 3578 8368
rect 3560 8354 3582 8356
rect 3587 8354 3617 8368
rect 3678 8366 3831 8370
rect 3660 8354 3852 8366
rect 3895 8354 3925 8368
rect 3931 8354 3944 8384
rect 3959 8366 3989 8384
rect 4032 8354 4045 8384
rect 4075 8354 4088 8384
rect 4103 8366 4133 8384
rect 4176 8370 4190 8384
rect 4226 8370 4446 8384
rect 4177 8368 4190 8370
rect 4143 8356 4158 8368
rect 4140 8354 4162 8356
rect 4167 8354 4197 8368
rect 4258 8366 4411 8370
rect 4240 8354 4432 8366
rect 4475 8354 4505 8368
rect 4511 8354 4524 8384
rect 4539 8366 4569 8384
rect 4612 8354 4625 8384
rect 4655 8354 4668 8384
rect 4683 8366 4713 8384
rect 4756 8370 4770 8384
rect 4806 8370 5026 8384
rect 4757 8368 4770 8370
rect 4723 8356 4738 8368
rect 4720 8354 4742 8356
rect 4747 8354 4777 8368
rect 4838 8366 4991 8370
rect 4820 8354 5012 8366
rect 5055 8354 5085 8368
rect 5091 8354 5104 8384
rect 5119 8366 5149 8384
rect 5192 8354 5205 8384
rect 5235 8354 5248 8384
rect 5263 8366 5293 8384
rect 5336 8370 5350 8384
rect 5386 8370 5606 8384
rect 5337 8368 5350 8370
rect 5303 8356 5318 8368
rect 5300 8354 5322 8356
rect 5327 8354 5357 8368
rect 5418 8366 5571 8370
rect 5400 8354 5592 8366
rect 5635 8354 5665 8368
rect 5671 8354 5684 8384
rect 5699 8366 5729 8384
rect 5772 8354 5785 8384
rect 5815 8354 5828 8384
rect 5843 8366 5873 8384
rect 5916 8370 5930 8384
rect 5966 8370 6186 8384
rect 5917 8368 5930 8370
rect 5883 8356 5898 8368
rect 5880 8354 5902 8356
rect 5907 8354 5937 8368
rect 5998 8366 6151 8370
rect 5980 8354 6172 8366
rect 6215 8354 6245 8368
rect 6251 8354 6264 8384
rect 6279 8366 6309 8384
rect 6352 8354 6365 8384
rect 6395 8354 6408 8384
rect 6423 8366 6453 8384
rect 6496 8370 6510 8384
rect 6546 8370 6766 8384
rect 6497 8368 6510 8370
rect 6463 8356 6478 8368
rect 6460 8354 6482 8356
rect 6487 8354 6517 8368
rect 6578 8366 6731 8370
rect 6560 8354 6752 8366
rect 6795 8354 6825 8368
rect 6831 8354 6844 8384
rect 6859 8366 6889 8384
rect 6932 8354 6945 8384
rect 6975 8354 6988 8384
rect 7003 8366 7033 8384
rect 7076 8370 7090 8384
rect 7126 8370 7346 8384
rect 7077 8368 7090 8370
rect 7043 8356 7058 8368
rect 7040 8354 7062 8356
rect 7067 8354 7097 8368
rect 7158 8366 7311 8370
rect 7140 8354 7332 8366
rect 7375 8354 7405 8368
rect 7411 8354 7424 8384
rect 7439 8366 7469 8384
rect 7512 8354 7525 8384
rect 7555 8354 7568 8384
rect 7583 8366 7613 8384
rect 7656 8370 7670 8384
rect 7706 8370 7926 8384
rect 7657 8368 7670 8370
rect 7623 8356 7638 8368
rect 7620 8354 7642 8356
rect 7647 8354 7677 8368
rect 7738 8366 7891 8370
rect 7720 8354 7912 8366
rect 7955 8354 7985 8368
rect 7991 8354 8004 8384
rect 8019 8366 8049 8384
rect 8092 8354 8105 8384
rect 8135 8354 8148 8384
rect 8163 8366 8193 8384
rect 8236 8370 8250 8384
rect 8286 8370 8506 8384
rect 8237 8368 8250 8370
rect 8203 8356 8218 8368
rect 8200 8354 8222 8356
rect 8227 8354 8257 8368
rect 8318 8366 8471 8370
rect 8300 8354 8492 8366
rect 8535 8354 8565 8368
rect 8571 8354 8584 8384
rect 8599 8366 8629 8384
rect 8672 8354 8685 8384
rect 8715 8354 8728 8384
rect 8743 8366 8773 8384
rect 8816 8370 8830 8384
rect 8866 8370 9086 8384
rect 8817 8368 8830 8370
rect 8783 8356 8798 8368
rect 8780 8354 8802 8356
rect 8807 8354 8837 8368
rect 8898 8366 9051 8370
rect 8880 8354 9072 8366
rect 9115 8354 9145 8368
rect 9151 8354 9164 8384
rect 9179 8366 9209 8384
rect 9252 8354 9265 8384
rect 0 8340 9265 8354
rect 15 8236 28 8340
rect 73 8318 74 8328
rect 89 8318 102 8328
rect 73 8314 102 8318
rect 107 8314 137 8340
rect 155 8326 171 8328
rect 243 8326 296 8340
rect 244 8324 308 8326
rect 351 8324 366 8340
rect 415 8337 445 8340
rect 415 8334 451 8337
rect 381 8326 397 8328
rect 155 8314 170 8318
rect 73 8312 170 8314
rect 198 8312 366 8324
rect 382 8314 397 8318
rect 415 8315 454 8334
rect 473 8328 480 8329
rect 479 8321 480 8328
rect 463 8318 464 8321
rect 479 8318 492 8321
rect 415 8314 445 8315
rect 454 8314 460 8315
rect 463 8314 492 8318
rect 382 8313 492 8314
rect 382 8312 498 8313
rect 57 8304 108 8312
rect 57 8292 82 8304
rect 89 8292 108 8304
rect 139 8304 189 8312
rect 139 8296 155 8304
rect 162 8302 189 8304
rect 198 8302 419 8312
rect 162 8292 419 8302
rect 448 8304 498 8312
rect 448 8295 464 8304
rect 57 8284 108 8292
rect 155 8284 419 8292
rect 445 8292 464 8295
rect 471 8292 498 8304
rect 445 8284 498 8292
rect 73 8276 74 8284
rect 89 8276 102 8284
rect 73 8268 89 8276
rect 70 8261 89 8264
rect 70 8252 92 8261
rect 43 8242 92 8252
rect 43 8236 73 8242
rect 92 8237 97 8242
rect 15 8220 89 8236
rect 107 8228 137 8284
rect 172 8274 380 8284
rect 415 8280 460 8284
rect 463 8283 464 8284
rect 479 8283 492 8284
rect 198 8244 387 8274
rect 213 8241 387 8244
rect 206 8238 387 8241
rect 15 8218 28 8220
rect 43 8218 77 8220
rect 15 8202 89 8218
rect 116 8214 129 8228
rect 144 8214 160 8230
rect 206 8225 217 8238
rect -1 8180 0 8196
rect 15 8180 28 8202
rect 43 8180 73 8202
rect 116 8198 178 8214
rect 206 8207 217 8223
rect 222 8218 232 8238
rect 242 8218 256 8238
rect 259 8225 268 8238
rect 284 8225 293 8238
rect 222 8207 256 8218
rect 259 8207 268 8223
rect 284 8207 293 8223
rect 300 8218 310 8238
rect 320 8218 334 8238
rect 335 8225 346 8238
rect 300 8207 334 8218
rect 335 8207 346 8223
rect 392 8214 408 8230
rect 415 8228 445 8280
rect 479 8276 480 8283
rect 464 8268 480 8276
rect 451 8236 464 8255
rect 479 8236 509 8252
rect 451 8220 525 8236
rect 451 8218 464 8220
rect 479 8218 513 8220
rect 116 8196 129 8198
rect 144 8196 178 8198
rect 116 8180 178 8196
rect 222 8191 238 8194
rect 300 8191 330 8202
rect 378 8198 424 8214
rect 451 8202 525 8218
rect 378 8196 412 8198
rect 377 8180 424 8196
rect 451 8180 464 8202
rect 479 8180 509 8202
rect 536 8180 537 8196
rect 552 8180 565 8340
rect 595 8236 608 8340
rect 653 8318 654 8328
rect 669 8318 682 8328
rect 653 8314 682 8318
rect 687 8314 717 8340
rect 735 8326 751 8328
rect 823 8326 876 8340
rect 824 8324 888 8326
rect 931 8324 946 8340
rect 995 8337 1025 8340
rect 995 8334 1031 8337
rect 961 8326 977 8328
rect 735 8314 750 8318
rect 653 8312 750 8314
rect 778 8312 946 8324
rect 962 8314 977 8318
rect 995 8315 1034 8334
rect 1053 8328 1060 8329
rect 1059 8321 1060 8328
rect 1043 8318 1044 8321
rect 1059 8318 1072 8321
rect 995 8314 1025 8315
rect 1034 8314 1040 8315
rect 1043 8314 1072 8318
rect 962 8313 1072 8314
rect 962 8312 1078 8313
rect 637 8304 688 8312
rect 637 8292 662 8304
rect 669 8292 688 8304
rect 719 8304 769 8312
rect 719 8296 735 8304
rect 742 8302 769 8304
rect 778 8302 999 8312
rect 742 8292 999 8302
rect 1028 8304 1078 8312
rect 1028 8295 1044 8304
rect 637 8284 688 8292
rect 735 8284 999 8292
rect 1025 8292 1044 8295
rect 1051 8292 1078 8304
rect 1025 8284 1078 8292
rect 653 8276 654 8284
rect 669 8276 682 8284
rect 653 8268 669 8276
rect 650 8261 669 8264
rect 650 8252 672 8261
rect 623 8242 672 8252
rect 623 8236 653 8242
rect 672 8237 677 8242
rect 595 8220 669 8236
rect 687 8228 717 8284
rect 752 8274 960 8284
rect 995 8280 1040 8284
rect 1043 8283 1044 8284
rect 1059 8283 1072 8284
rect 778 8244 967 8274
rect 793 8241 967 8244
rect 786 8238 967 8241
rect 595 8218 608 8220
rect 623 8218 657 8220
rect 595 8202 669 8218
rect 696 8214 709 8228
rect 724 8214 740 8230
rect 786 8225 797 8238
rect 579 8180 580 8196
rect 595 8180 608 8202
rect 623 8180 653 8202
rect 696 8198 758 8214
rect 786 8207 797 8223
rect 802 8218 812 8238
rect 822 8218 836 8238
rect 839 8225 848 8238
rect 864 8225 873 8238
rect 802 8207 836 8218
rect 839 8207 848 8223
rect 864 8207 873 8223
rect 880 8218 890 8238
rect 900 8218 914 8238
rect 915 8225 926 8238
rect 880 8207 914 8218
rect 915 8207 926 8223
rect 972 8214 988 8230
rect 995 8228 1025 8280
rect 1059 8276 1060 8283
rect 1044 8268 1060 8276
rect 1031 8236 1044 8255
rect 1059 8236 1089 8252
rect 1031 8220 1105 8236
rect 1031 8218 1044 8220
rect 1059 8218 1093 8220
rect 696 8196 709 8198
rect 724 8196 758 8198
rect 696 8180 758 8196
rect 802 8191 818 8194
rect 880 8191 910 8202
rect 958 8198 1004 8214
rect 1031 8202 1105 8218
rect 958 8196 992 8198
rect 957 8180 1004 8196
rect 1031 8180 1044 8202
rect 1059 8180 1089 8202
rect 1116 8180 1117 8196
rect 1132 8180 1145 8340
rect 1175 8236 1188 8340
rect 1233 8318 1234 8328
rect 1249 8318 1262 8328
rect 1233 8314 1262 8318
rect 1267 8314 1297 8340
rect 1315 8326 1331 8328
rect 1403 8326 1456 8340
rect 1404 8324 1468 8326
rect 1511 8324 1526 8340
rect 1575 8337 1605 8340
rect 1575 8334 1611 8337
rect 1541 8326 1557 8328
rect 1315 8314 1330 8318
rect 1233 8312 1330 8314
rect 1358 8312 1526 8324
rect 1542 8314 1557 8318
rect 1575 8315 1614 8334
rect 1633 8328 1640 8329
rect 1639 8321 1640 8328
rect 1623 8318 1624 8321
rect 1639 8318 1652 8321
rect 1575 8314 1605 8315
rect 1614 8314 1620 8315
rect 1623 8314 1652 8318
rect 1542 8313 1652 8314
rect 1542 8312 1658 8313
rect 1217 8304 1268 8312
rect 1217 8292 1242 8304
rect 1249 8292 1268 8304
rect 1299 8304 1349 8312
rect 1299 8296 1315 8304
rect 1322 8302 1349 8304
rect 1358 8302 1579 8312
rect 1322 8292 1579 8302
rect 1608 8304 1658 8312
rect 1608 8295 1624 8304
rect 1217 8284 1268 8292
rect 1315 8284 1579 8292
rect 1605 8292 1624 8295
rect 1631 8292 1658 8304
rect 1605 8284 1658 8292
rect 1233 8276 1234 8284
rect 1249 8276 1262 8284
rect 1233 8268 1249 8276
rect 1230 8261 1249 8264
rect 1230 8252 1252 8261
rect 1203 8242 1252 8252
rect 1203 8236 1233 8242
rect 1252 8237 1257 8242
rect 1175 8220 1249 8236
rect 1267 8228 1297 8284
rect 1332 8274 1540 8284
rect 1575 8280 1620 8284
rect 1623 8283 1624 8284
rect 1639 8283 1652 8284
rect 1358 8244 1547 8274
rect 1373 8241 1547 8244
rect 1366 8238 1547 8241
rect 1175 8218 1188 8220
rect 1203 8218 1237 8220
rect 1175 8202 1249 8218
rect 1276 8214 1289 8228
rect 1304 8214 1320 8230
rect 1366 8225 1377 8238
rect 1159 8180 1160 8196
rect 1175 8180 1188 8202
rect 1203 8180 1233 8202
rect 1276 8198 1338 8214
rect 1366 8207 1377 8223
rect 1382 8218 1392 8238
rect 1402 8218 1416 8238
rect 1419 8225 1428 8238
rect 1444 8225 1453 8238
rect 1382 8207 1416 8218
rect 1419 8207 1428 8223
rect 1444 8207 1453 8223
rect 1460 8218 1470 8238
rect 1480 8218 1494 8238
rect 1495 8225 1506 8238
rect 1460 8207 1494 8218
rect 1495 8207 1506 8223
rect 1552 8214 1568 8230
rect 1575 8228 1605 8280
rect 1639 8276 1640 8283
rect 1624 8268 1640 8276
rect 1611 8236 1624 8255
rect 1639 8236 1669 8252
rect 1611 8220 1685 8236
rect 1611 8218 1624 8220
rect 1639 8218 1673 8220
rect 1276 8196 1289 8198
rect 1304 8196 1338 8198
rect 1276 8180 1338 8196
rect 1382 8191 1398 8194
rect 1460 8191 1490 8202
rect 1538 8198 1584 8214
rect 1611 8202 1685 8218
rect 1538 8196 1572 8198
rect 1537 8180 1584 8196
rect 1611 8180 1624 8202
rect 1639 8180 1669 8202
rect 1696 8180 1697 8196
rect 1712 8180 1725 8340
rect 1755 8236 1768 8340
rect 1813 8318 1814 8328
rect 1829 8318 1842 8328
rect 1813 8314 1842 8318
rect 1847 8314 1877 8340
rect 1895 8326 1911 8328
rect 1983 8326 2036 8340
rect 1984 8324 2048 8326
rect 2091 8324 2106 8340
rect 2155 8337 2185 8340
rect 2155 8334 2191 8337
rect 2121 8326 2137 8328
rect 1895 8314 1910 8318
rect 1813 8312 1910 8314
rect 1938 8312 2106 8324
rect 2122 8314 2137 8318
rect 2155 8315 2194 8334
rect 2213 8328 2220 8329
rect 2219 8321 2220 8328
rect 2203 8318 2204 8321
rect 2219 8318 2232 8321
rect 2155 8314 2185 8315
rect 2194 8314 2200 8315
rect 2203 8314 2232 8318
rect 2122 8313 2232 8314
rect 2122 8312 2238 8313
rect 1797 8304 1848 8312
rect 1797 8292 1822 8304
rect 1829 8292 1848 8304
rect 1879 8304 1929 8312
rect 1879 8296 1895 8304
rect 1902 8302 1929 8304
rect 1938 8302 2159 8312
rect 1902 8292 2159 8302
rect 2188 8304 2238 8312
rect 2188 8295 2204 8304
rect 1797 8284 1848 8292
rect 1895 8284 2159 8292
rect 2185 8292 2204 8295
rect 2211 8292 2238 8304
rect 2185 8284 2238 8292
rect 1813 8276 1814 8284
rect 1829 8276 1842 8284
rect 1813 8268 1829 8276
rect 1810 8261 1829 8264
rect 1810 8252 1832 8261
rect 1783 8242 1832 8252
rect 1783 8236 1813 8242
rect 1832 8237 1837 8242
rect 1755 8220 1829 8236
rect 1847 8228 1877 8284
rect 1912 8274 2120 8284
rect 2155 8280 2200 8284
rect 2203 8283 2204 8284
rect 2219 8283 2232 8284
rect 1938 8244 2127 8274
rect 1953 8241 2127 8244
rect 1946 8238 2127 8241
rect 1755 8218 1768 8220
rect 1783 8218 1817 8220
rect 1755 8202 1829 8218
rect 1856 8214 1869 8228
rect 1884 8214 1900 8230
rect 1946 8225 1957 8238
rect 1739 8180 1740 8196
rect 1755 8180 1768 8202
rect 1783 8180 1813 8202
rect 1856 8198 1918 8214
rect 1946 8207 1957 8223
rect 1962 8218 1972 8238
rect 1982 8218 1996 8238
rect 1999 8225 2008 8238
rect 2024 8225 2033 8238
rect 1962 8207 1996 8218
rect 1999 8207 2008 8223
rect 2024 8207 2033 8223
rect 2040 8218 2050 8238
rect 2060 8218 2074 8238
rect 2075 8225 2086 8238
rect 2040 8207 2074 8218
rect 2075 8207 2086 8223
rect 2132 8214 2148 8230
rect 2155 8228 2185 8280
rect 2219 8276 2220 8283
rect 2204 8268 2220 8276
rect 2191 8236 2204 8255
rect 2219 8236 2249 8252
rect 2191 8220 2265 8236
rect 2191 8218 2204 8220
rect 2219 8218 2253 8220
rect 1856 8196 1869 8198
rect 1884 8196 1918 8198
rect 1856 8180 1918 8196
rect 1962 8191 1976 8194
rect 2040 8191 2070 8202
rect 2118 8198 2164 8214
rect 2191 8202 2265 8218
rect 2118 8196 2152 8198
rect 2117 8180 2164 8196
rect 2191 8180 2204 8202
rect 2219 8180 2249 8202
rect 2276 8180 2277 8196
rect 2292 8180 2305 8340
rect 2335 8236 2348 8340
rect 2393 8318 2394 8328
rect 2409 8318 2422 8328
rect 2393 8314 2422 8318
rect 2427 8314 2457 8340
rect 2475 8326 2491 8328
rect 2563 8326 2616 8340
rect 2564 8324 2628 8326
rect 2671 8324 2686 8340
rect 2735 8337 2765 8340
rect 2735 8334 2771 8337
rect 2701 8326 2717 8328
rect 2475 8314 2490 8318
rect 2393 8312 2490 8314
rect 2518 8312 2686 8324
rect 2702 8314 2717 8318
rect 2735 8315 2774 8334
rect 2793 8328 2800 8329
rect 2799 8321 2800 8328
rect 2783 8318 2784 8321
rect 2799 8318 2812 8321
rect 2735 8314 2765 8315
rect 2774 8314 2780 8315
rect 2783 8314 2812 8318
rect 2702 8313 2812 8314
rect 2702 8312 2818 8313
rect 2377 8304 2428 8312
rect 2377 8292 2402 8304
rect 2409 8292 2428 8304
rect 2459 8304 2509 8312
rect 2459 8296 2475 8304
rect 2482 8302 2509 8304
rect 2518 8302 2739 8312
rect 2482 8292 2739 8302
rect 2768 8304 2818 8312
rect 2768 8295 2784 8304
rect 2377 8284 2428 8292
rect 2475 8284 2739 8292
rect 2765 8292 2784 8295
rect 2791 8292 2818 8304
rect 2765 8284 2818 8292
rect 2393 8276 2394 8284
rect 2409 8276 2422 8284
rect 2393 8268 2409 8276
rect 2390 8261 2409 8264
rect 2390 8252 2412 8261
rect 2363 8242 2412 8252
rect 2363 8236 2393 8242
rect 2412 8237 2417 8242
rect 2335 8220 2409 8236
rect 2427 8228 2457 8284
rect 2492 8274 2700 8284
rect 2735 8280 2780 8284
rect 2783 8283 2784 8284
rect 2799 8283 2812 8284
rect 2518 8244 2707 8274
rect 2533 8241 2707 8244
rect 2526 8238 2707 8241
rect 2335 8218 2348 8220
rect 2363 8218 2397 8220
rect 2335 8202 2409 8218
rect 2436 8214 2449 8228
rect 2464 8214 2480 8230
rect 2526 8225 2537 8238
rect 2319 8180 2320 8196
rect 2335 8180 2348 8202
rect 2363 8180 2393 8202
rect 2436 8198 2498 8214
rect 2526 8207 2537 8223
rect 2542 8218 2552 8238
rect 2562 8218 2576 8238
rect 2579 8225 2588 8238
rect 2604 8225 2613 8238
rect 2542 8207 2576 8218
rect 2579 8207 2588 8223
rect 2604 8207 2613 8223
rect 2620 8218 2630 8238
rect 2640 8218 2654 8238
rect 2655 8225 2666 8238
rect 2620 8207 2654 8218
rect 2655 8207 2666 8223
rect 2712 8214 2728 8230
rect 2735 8228 2765 8280
rect 2799 8276 2800 8283
rect 2784 8268 2800 8276
rect 2771 8236 2784 8255
rect 2799 8236 2829 8252
rect 2771 8220 2845 8236
rect 2771 8218 2784 8220
rect 2799 8218 2833 8220
rect 2436 8196 2449 8198
rect 2464 8196 2498 8198
rect 2436 8180 2498 8196
rect 2542 8191 2558 8194
rect 2620 8191 2650 8202
rect 2698 8198 2744 8214
rect 2771 8202 2845 8218
rect 2698 8196 2732 8198
rect 2697 8180 2744 8196
rect 2771 8180 2784 8202
rect 2799 8180 2829 8202
rect 2856 8180 2857 8196
rect 2872 8180 2885 8340
rect 2915 8236 2928 8340
rect 2973 8318 2974 8328
rect 2989 8318 3002 8328
rect 2973 8314 3002 8318
rect 3007 8314 3037 8340
rect 3055 8326 3071 8328
rect 3143 8326 3196 8340
rect 3144 8324 3208 8326
rect 3251 8324 3266 8340
rect 3315 8337 3345 8340
rect 3315 8334 3351 8337
rect 3281 8326 3297 8328
rect 3055 8314 3070 8318
rect 2973 8312 3070 8314
rect 3098 8312 3266 8324
rect 3282 8314 3297 8318
rect 3315 8315 3354 8334
rect 3373 8328 3380 8329
rect 3379 8321 3380 8328
rect 3363 8318 3364 8321
rect 3379 8318 3392 8321
rect 3315 8314 3345 8315
rect 3354 8314 3360 8315
rect 3363 8314 3392 8318
rect 3282 8313 3392 8314
rect 3282 8312 3398 8313
rect 2957 8304 3008 8312
rect 2957 8292 2982 8304
rect 2989 8292 3008 8304
rect 3039 8304 3089 8312
rect 3039 8296 3055 8304
rect 3062 8302 3089 8304
rect 3098 8302 3319 8312
rect 3062 8292 3319 8302
rect 3348 8304 3398 8312
rect 3348 8295 3364 8304
rect 2957 8284 3008 8292
rect 3055 8284 3319 8292
rect 3345 8292 3364 8295
rect 3371 8292 3398 8304
rect 3345 8284 3398 8292
rect 2973 8276 2974 8284
rect 2989 8276 3002 8284
rect 2973 8268 2989 8276
rect 2970 8261 2989 8264
rect 2970 8252 2992 8261
rect 2943 8242 2992 8252
rect 2943 8236 2973 8242
rect 2992 8237 2997 8242
rect 2915 8220 2989 8236
rect 3007 8228 3037 8284
rect 3072 8274 3280 8284
rect 3315 8280 3360 8284
rect 3363 8283 3364 8284
rect 3379 8283 3392 8284
rect 3098 8244 3287 8274
rect 3113 8241 3287 8244
rect 3106 8238 3287 8241
rect 2915 8218 2928 8220
rect 2943 8218 2977 8220
rect 2915 8202 2989 8218
rect 3016 8214 3029 8228
rect 3044 8214 3060 8230
rect 3106 8225 3117 8238
rect 2899 8180 2900 8196
rect 2915 8180 2928 8202
rect 2943 8180 2973 8202
rect 3016 8198 3078 8214
rect 3106 8207 3117 8223
rect 3122 8218 3132 8238
rect 3142 8218 3156 8238
rect 3159 8225 3168 8238
rect 3184 8225 3193 8238
rect 3122 8207 3156 8218
rect 3159 8207 3168 8223
rect 3184 8207 3193 8223
rect 3200 8218 3210 8238
rect 3220 8218 3234 8238
rect 3235 8225 3246 8238
rect 3200 8207 3234 8218
rect 3235 8207 3246 8223
rect 3292 8214 3308 8230
rect 3315 8228 3345 8280
rect 3379 8276 3380 8283
rect 3364 8268 3380 8276
rect 3351 8236 3364 8255
rect 3379 8236 3409 8252
rect 3351 8220 3425 8236
rect 3351 8218 3364 8220
rect 3379 8218 3413 8220
rect 3016 8196 3029 8198
rect 3044 8196 3078 8198
rect 3016 8180 3078 8196
rect 3122 8191 3138 8194
rect 3200 8191 3230 8202
rect 3278 8198 3324 8214
rect 3351 8202 3425 8218
rect 3278 8196 3312 8198
rect 3277 8180 3324 8196
rect 3351 8180 3364 8202
rect 3379 8180 3409 8202
rect 3436 8180 3437 8196
rect 3452 8180 3465 8340
rect 3495 8236 3508 8340
rect 3553 8318 3554 8328
rect 3569 8318 3582 8328
rect 3553 8314 3582 8318
rect 3587 8314 3617 8340
rect 3635 8326 3651 8328
rect 3723 8326 3776 8340
rect 3724 8324 3788 8326
rect 3831 8324 3846 8340
rect 3895 8337 3925 8340
rect 3895 8334 3931 8337
rect 3861 8326 3877 8328
rect 3635 8314 3650 8318
rect 3553 8312 3650 8314
rect 3678 8312 3846 8324
rect 3862 8314 3877 8318
rect 3895 8315 3934 8334
rect 3953 8328 3960 8329
rect 3959 8321 3960 8328
rect 3943 8318 3944 8321
rect 3959 8318 3972 8321
rect 3895 8314 3925 8315
rect 3934 8314 3940 8315
rect 3943 8314 3972 8318
rect 3862 8313 3972 8314
rect 3862 8312 3978 8313
rect 3537 8304 3588 8312
rect 3537 8292 3562 8304
rect 3569 8292 3588 8304
rect 3619 8304 3669 8312
rect 3619 8296 3635 8304
rect 3642 8302 3669 8304
rect 3678 8302 3899 8312
rect 3642 8292 3899 8302
rect 3928 8304 3978 8312
rect 3928 8295 3944 8304
rect 3537 8284 3588 8292
rect 3635 8284 3899 8292
rect 3925 8292 3944 8295
rect 3951 8292 3978 8304
rect 3925 8284 3978 8292
rect 3553 8276 3554 8284
rect 3569 8276 3582 8284
rect 3553 8268 3569 8276
rect 3550 8261 3569 8264
rect 3550 8252 3572 8261
rect 3523 8242 3572 8252
rect 3523 8236 3553 8242
rect 3572 8237 3577 8242
rect 3495 8220 3569 8236
rect 3587 8228 3617 8284
rect 3652 8274 3860 8284
rect 3895 8280 3940 8284
rect 3943 8283 3944 8284
rect 3959 8283 3972 8284
rect 3678 8244 3867 8274
rect 3693 8241 3867 8244
rect 3686 8238 3867 8241
rect 3495 8218 3508 8220
rect 3523 8218 3557 8220
rect 3495 8202 3569 8218
rect 3596 8214 3609 8228
rect 3624 8214 3640 8230
rect 3686 8225 3697 8238
rect 3479 8180 3480 8196
rect 3495 8180 3508 8202
rect 3523 8180 3553 8202
rect 3596 8198 3658 8214
rect 3686 8207 3697 8223
rect 3702 8218 3712 8238
rect 3722 8218 3736 8238
rect 3739 8225 3748 8238
rect 3764 8225 3773 8238
rect 3702 8207 3736 8218
rect 3739 8207 3748 8223
rect 3764 8207 3773 8223
rect 3780 8218 3790 8238
rect 3800 8218 3814 8238
rect 3815 8225 3826 8238
rect 3780 8207 3814 8218
rect 3815 8207 3826 8223
rect 3872 8214 3888 8230
rect 3895 8228 3925 8280
rect 3959 8276 3960 8283
rect 3944 8268 3960 8276
rect 3931 8236 3944 8255
rect 3959 8236 3989 8252
rect 3931 8220 4005 8236
rect 3931 8218 3944 8220
rect 3959 8218 3993 8220
rect 3596 8196 3609 8198
rect 3624 8196 3658 8198
rect 3596 8180 3658 8196
rect 3702 8191 3718 8194
rect 3780 8191 3810 8202
rect 3858 8198 3904 8214
rect 3931 8202 4005 8218
rect 3858 8196 3892 8198
rect 3857 8180 3904 8196
rect 3931 8180 3944 8202
rect 3959 8180 3989 8202
rect 4016 8180 4017 8196
rect 4032 8180 4045 8340
rect 4075 8236 4088 8340
rect 4133 8318 4134 8328
rect 4149 8318 4162 8328
rect 4133 8314 4162 8318
rect 4167 8314 4197 8340
rect 4215 8326 4231 8328
rect 4303 8326 4356 8340
rect 4304 8324 4368 8326
rect 4411 8324 4426 8340
rect 4475 8337 4505 8340
rect 4475 8334 4511 8337
rect 4441 8326 4457 8328
rect 4215 8314 4230 8318
rect 4133 8312 4230 8314
rect 4258 8312 4426 8324
rect 4442 8314 4457 8318
rect 4475 8315 4514 8334
rect 4533 8328 4540 8329
rect 4539 8321 4540 8328
rect 4523 8318 4524 8321
rect 4539 8318 4552 8321
rect 4475 8314 4505 8315
rect 4514 8314 4520 8315
rect 4523 8314 4552 8318
rect 4442 8313 4552 8314
rect 4442 8312 4558 8313
rect 4117 8304 4168 8312
rect 4117 8292 4142 8304
rect 4149 8292 4168 8304
rect 4199 8304 4249 8312
rect 4199 8296 4215 8304
rect 4222 8302 4249 8304
rect 4258 8302 4479 8312
rect 4222 8292 4479 8302
rect 4508 8304 4558 8312
rect 4508 8295 4524 8304
rect 4117 8284 4168 8292
rect 4215 8284 4479 8292
rect 4505 8292 4524 8295
rect 4531 8292 4558 8304
rect 4505 8284 4558 8292
rect 4133 8276 4134 8284
rect 4149 8276 4162 8284
rect 4133 8268 4149 8276
rect 4130 8261 4149 8264
rect 4130 8252 4152 8261
rect 4103 8242 4152 8252
rect 4103 8236 4133 8242
rect 4152 8237 4157 8242
rect 4075 8220 4149 8236
rect 4167 8228 4197 8284
rect 4232 8274 4440 8284
rect 4475 8280 4520 8284
rect 4523 8283 4524 8284
rect 4539 8283 4552 8284
rect 4258 8244 4447 8274
rect 4273 8241 4447 8244
rect 4266 8238 4447 8241
rect 4075 8218 4088 8220
rect 4103 8218 4137 8220
rect 4075 8202 4149 8218
rect 4176 8214 4189 8228
rect 4204 8214 4220 8230
rect 4266 8225 4277 8238
rect 4059 8180 4060 8196
rect 4075 8180 4088 8202
rect 4103 8180 4133 8202
rect 4176 8198 4238 8214
rect 4266 8207 4277 8223
rect 4282 8218 4292 8238
rect 4302 8218 4316 8238
rect 4319 8225 4328 8238
rect 4344 8225 4353 8238
rect 4282 8207 4316 8218
rect 4319 8207 4328 8223
rect 4344 8207 4353 8223
rect 4360 8218 4370 8238
rect 4380 8218 4394 8238
rect 4395 8225 4406 8238
rect 4360 8207 4394 8218
rect 4395 8207 4406 8223
rect 4452 8214 4468 8230
rect 4475 8228 4505 8280
rect 4539 8276 4540 8283
rect 4524 8268 4540 8276
rect 4511 8236 4524 8255
rect 4539 8236 4569 8252
rect 4511 8220 4585 8236
rect 4511 8218 4524 8220
rect 4539 8218 4573 8220
rect 4176 8196 4189 8198
rect 4204 8196 4238 8198
rect 4176 8180 4238 8196
rect 4282 8191 4298 8194
rect 4360 8191 4390 8202
rect 4438 8198 4484 8214
rect 4511 8202 4585 8218
rect 4438 8196 4472 8198
rect 4437 8180 4484 8196
rect 4511 8180 4524 8202
rect 4539 8180 4569 8202
rect 4596 8180 4597 8196
rect 4612 8180 4625 8340
rect 4655 8236 4668 8340
rect 4713 8318 4714 8328
rect 4729 8318 4742 8328
rect 4713 8314 4742 8318
rect 4747 8314 4777 8340
rect 4795 8326 4811 8328
rect 4883 8326 4936 8340
rect 4884 8324 4948 8326
rect 4991 8324 5006 8340
rect 5055 8337 5085 8340
rect 5055 8334 5091 8337
rect 5021 8326 5037 8328
rect 4795 8314 4810 8318
rect 4713 8312 4810 8314
rect 4838 8312 5006 8324
rect 5022 8314 5037 8318
rect 5055 8315 5094 8334
rect 5113 8328 5120 8329
rect 5119 8321 5120 8328
rect 5103 8318 5104 8321
rect 5119 8318 5132 8321
rect 5055 8314 5085 8315
rect 5094 8314 5100 8315
rect 5103 8314 5132 8318
rect 5022 8313 5132 8314
rect 5022 8312 5138 8313
rect 4697 8304 4748 8312
rect 4697 8292 4722 8304
rect 4729 8292 4748 8304
rect 4779 8304 4829 8312
rect 4779 8296 4795 8304
rect 4802 8302 4829 8304
rect 4838 8302 5059 8312
rect 4802 8292 5059 8302
rect 5088 8304 5138 8312
rect 5088 8295 5104 8304
rect 4697 8284 4748 8292
rect 4795 8284 5059 8292
rect 5085 8292 5104 8295
rect 5111 8292 5138 8304
rect 5085 8284 5138 8292
rect 4713 8276 4714 8284
rect 4729 8276 4742 8284
rect 4713 8268 4729 8276
rect 4710 8261 4729 8264
rect 4710 8252 4732 8261
rect 4683 8242 4732 8252
rect 4683 8236 4713 8242
rect 4732 8237 4737 8242
rect 4655 8220 4729 8236
rect 4747 8228 4777 8284
rect 4812 8274 5020 8284
rect 5055 8280 5100 8284
rect 5103 8283 5104 8284
rect 5119 8283 5132 8284
rect 4838 8244 5027 8274
rect 4853 8241 5027 8244
rect 4846 8238 5027 8241
rect 4655 8218 4668 8220
rect 4683 8218 4717 8220
rect 4655 8202 4729 8218
rect 4756 8214 4769 8228
rect 4784 8214 4800 8230
rect 4846 8225 4857 8238
rect 4639 8180 4640 8196
rect 4655 8180 4668 8202
rect 4683 8180 4713 8202
rect 4756 8198 4818 8214
rect 4846 8207 4857 8223
rect 4862 8218 4872 8238
rect 4882 8218 4896 8238
rect 4899 8225 4908 8238
rect 4924 8225 4933 8238
rect 4862 8207 4896 8218
rect 4899 8207 4908 8223
rect 4924 8207 4933 8223
rect 4940 8218 4950 8238
rect 4960 8218 4974 8238
rect 4975 8225 4986 8238
rect 4940 8207 4974 8218
rect 4975 8207 4986 8223
rect 5032 8214 5048 8230
rect 5055 8228 5085 8280
rect 5119 8276 5120 8283
rect 5104 8268 5120 8276
rect 5091 8236 5104 8255
rect 5119 8236 5149 8252
rect 5091 8220 5165 8236
rect 5091 8218 5104 8220
rect 5119 8218 5153 8220
rect 4756 8196 4769 8198
rect 4784 8196 4818 8198
rect 4756 8180 4818 8196
rect 4862 8191 4878 8194
rect 4940 8191 4970 8202
rect 5018 8198 5064 8214
rect 5091 8202 5165 8218
rect 5018 8196 5052 8198
rect 5017 8180 5064 8196
rect 5091 8180 5104 8202
rect 5119 8180 5149 8202
rect 5176 8180 5177 8196
rect 5192 8180 5205 8340
rect 5235 8236 5248 8340
rect 5293 8318 5294 8328
rect 5309 8318 5322 8328
rect 5293 8314 5322 8318
rect 5327 8314 5357 8340
rect 5375 8326 5391 8328
rect 5463 8326 5516 8340
rect 5464 8324 5528 8326
rect 5571 8324 5586 8340
rect 5635 8337 5665 8340
rect 5635 8334 5671 8337
rect 5601 8326 5617 8328
rect 5375 8314 5390 8318
rect 5293 8312 5390 8314
rect 5418 8312 5586 8324
rect 5602 8314 5617 8318
rect 5635 8315 5674 8334
rect 5693 8328 5700 8329
rect 5699 8321 5700 8328
rect 5683 8318 5684 8321
rect 5699 8318 5712 8321
rect 5635 8314 5665 8315
rect 5674 8314 5680 8315
rect 5683 8314 5712 8318
rect 5602 8313 5712 8314
rect 5602 8312 5718 8313
rect 5277 8304 5328 8312
rect 5277 8292 5302 8304
rect 5309 8292 5328 8304
rect 5359 8304 5409 8312
rect 5359 8296 5375 8304
rect 5382 8302 5409 8304
rect 5418 8302 5639 8312
rect 5382 8292 5639 8302
rect 5668 8304 5718 8312
rect 5668 8295 5684 8304
rect 5277 8284 5328 8292
rect 5375 8284 5639 8292
rect 5665 8292 5684 8295
rect 5691 8292 5718 8304
rect 5665 8284 5718 8292
rect 5293 8276 5294 8284
rect 5309 8276 5322 8284
rect 5293 8268 5309 8276
rect 5290 8261 5309 8264
rect 5290 8252 5312 8261
rect 5263 8242 5312 8252
rect 5263 8236 5293 8242
rect 5312 8237 5317 8242
rect 5235 8220 5309 8236
rect 5327 8228 5357 8284
rect 5392 8274 5600 8284
rect 5635 8280 5680 8284
rect 5683 8283 5684 8284
rect 5699 8283 5712 8284
rect 5418 8244 5607 8274
rect 5433 8241 5607 8244
rect 5426 8238 5607 8241
rect 5235 8218 5248 8220
rect 5263 8218 5297 8220
rect 5235 8202 5309 8218
rect 5336 8214 5349 8228
rect 5364 8214 5380 8230
rect 5426 8225 5437 8238
rect 5219 8180 5220 8196
rect 5235 8180 5248 8202
rect 5263 8180 5293 8202
rect 5336 8198 5398 8214
rect 5426 8207 5437 8223
rect 5442 8218 5452 8238
rect 5462 8218 5476 8238
rect 5479 8225 5488 8238
rect 5504 8225 5513 8238
rect 5442 8207 5476 8218
rect 5479 8207 5488 8223
rect 5504 8207 5513 8223
rect 5520 8218 5530 8238
rect 5540 8218 5554 8238
rect 5555 8225 5566 8238
rect 5520 8207 5554 8218
rect 5555 8207 5566 8223
rect 5612 8214 5628 8230
rect 5635 8228 5665 8280
rect 5699 8276 5700 8283
rect 5684 8268 5700 8276
rect 5671 8236 5684 8255
rect 5699 8236 5729 8252
rect 5671 8220 5745 8236
rect 5671 8218 5684 8220
rect 5699 8218 5733 8220
rect 5336 8196 5349 8198
rect 5364 8196 5398 8198
rect 5336 8180 5398 8196
rect 5442 8191 5458 8194
rect 5520 8191 5550 8202
rect 5598 8198 5644 8214
rect 5671 8202 5745 8218
rect 5598 8196 5632 8198
rect 5597 8180 5644 8196
rect 5671 8180 5684 8202
rect 5699 8180 5729 8202
rect 5756 8180 5757 8196
rect 5772 8180 5785 8340
rect 5815 8236 5828 8340
rect 5873 8318 5874 8328
rect 5889 8318 5902 8328
rect 5873 8314 5902 8318
rect 5907 8314 5937 8340
rect 5955 8326 5971 8328
rect 6043 8326 6096 8340
rect 6044 8324 6108 8326
rect 6151 8324 6166 8340
rect 6215 8337 6245 8340
rect 6215 8334 6251 8337
rect 6181 8326 6197 8328
rect 5955 8314 5970 8318
rect 5873 8312 5970 8314
rect 5998 8312 6166 8324
rect 6182 8314 6197 8318
rect 6215 8315 6254 8334
rect 6273 8328 6280 8329
rect 6279 8321 6280 8328
rect 6263 8318 6264 8321
rect 6279 8318 6292 8321
rect 6215 8314 6245 8315
rect 6254 8314 6260 8315
rect 6263 8314 6292 8318
rect 6182 8313 6292 8314
rect 6182 8312 6298 8313
rect 5857 8304 5908 8312
rect 5857 8292 5882 8304
rect 5889 8292 5908 8304
rect 5939 8304 5989 8312
rect 5939 8296 5955 8304
rect 5962 8302 5989 8304
rect 5998 8302 6219 8312
rect 5962 8292 6219 8302
rect 6248 8304 6298 8312
rect 6248 8295 6264 8304
rect 5857 8284 5908 8292
rect 5955 8284 6219 8292
rect 6245 8292 6264 8295
rect 6271 8292 6298 8304
rect 6245 8284 6298 8292
rect 5873 8276 5874 8284
rect 5889 8276 5902 8284
rect 5873 8268 5889 8276
rect 5870 8261 5889 8264
rect 5870 8252 5892 8261
rect 5843 8242 5892 8252
rect 5843 8236 5873 8242
rect 5892 8237 5897 8242
rect 5815 8220 5889 8236
rect 5907 8228 5937 8284
rect 5972 8274 6180 8284
rect 6215 8280 6260 8284
rect 6263 8283 6264 8284
rect 6279 8283 6292 8284
rect 5998 8244 6187 8274
rect 6013 8241 6187 8244
rect 6006 8238 6187 8241
rect 5815 8218 5828 8220
rect 5843 8218 5877 8220
rect 5815 8202 5889 8218
rect 5916 8214 5929 8228
rect 5944 8214 5960 8230
rect 6006 8225 6017 8238
rect 5799 8180 5800 8196
rect 5815 8180 5828 8202
rect 5843 8180 5873 8202
rect 5916 8198 5978 8214
rect 6006 8207 6017 8223
rect 6022 8218 6032 8238
rect 6042 8218 6056 8238
rect 6059 8225 6068 8238
rect 6084 8225 6093 8238
rect 6022 8207 6056 8218
rect 6059 8207 6068 8223
rect 6084 8207 6093 8223
rect 6100 8218 6110 8238
rect 6120 8218 6134 8238
rect 6135 8225 6146 8238
rect 6100 8207 6134 8218
rect 6135 8207 6146 8223
rect 6192 8214 6208 8230
rect 6215 8228 6245 8280
rect 6279 8276 6280 8283
rect 6264 8268 6280 8276
rect 6251 8236 6264 8255
rect 6279 8236 6309 8252
rect 6251 8220 6325 8236
rect 6251 8218 6264 8220
rect 6279 8218 6313 8220
rect 5916 8196 5929 8198
rect 5944 8196 5978 8198
rect 5916 8180 5978 8196
rect 6022 8191 6038 8194
rect 6100 8191 6130 8202
rect 6178 8198 6224 8214
rect 6251 8202 6325 8218
rect 6178 8196 6212 8198
rect 6177 8180 6224 8196
rect 6251 8180 6264 8202
rect 6279 8180 6309 8202
rect 6336 8180 6337 8196
rect 6352 8180 6365 8340
rect 6395 8236 6408 8340
rect 6453 8318 6454 8328
rect 6469 8318 6482 8328
rect 6453 8314 6482 8318
rect 6487 8314 6517 8340
rect 6535 8326 6551 8328
rect 6623 8326 6676 8340
rect 6624 8324 6688 8326
rect 6731 8324 6746 8340
rect 6795 8337 6825 8340
rect 6795 8334 6831 8337
rect 6761 8326 6777 8328
rect 6535 8314 6550 8318
rect 6453 8312 6550 8314
rect 6578 8312 6746 8324
rect 6762 8314 6777 8318
rect 6795 8315 6834 8334
rect 6853 8328 6860 8329
rect 6859 8321 6860 8328
rect 6843 8318 6844 8321
rect 6859 8318 6872 8321
rect 6795 8314 6825 8315
rect 6834 8314 6840 8315
rect 6843 8314 6872 8318
rect 6762 8313 6872 8314
rect 6762 8312 6878 8313
rect 6437 8304 6488 8312
rect 6437 8292 6462 8304
rect 6469 8292 6488 8304
rect 6519 8304 6569 8312
rect 6519 8296 6535 8304
rect 6542 8302 6569 8304
rect 6578 8302 6799 8312
rect 6542 8292 6799 8302
rect 6828 8304 6878 8312
rect 6828 8295 6844 8304
rect 6437 8284 6488 8292
rect 6535 8284 6799 8292
rect 6825 8292 6844 8295
rect 6851 8292 6878 8304
rect 6825 8284 6878 8292
rect 6453 8276 6454 8284
rect 6469 8276 6482 8284
rect 6453 8268 6469 8276
rect 6450 8261 6469 8264
rect 6450 8252 6472 8261
rect 6423 8242 6472 8252
rect 6423 8236 6453 8242
rect 6472 8237 6477 8242
rect 6395 8220 6469 8236
rect 6487 8228 6517 8284
rect 6552 8274 6760 8284
rect 6795 8280 6840 8284
rect 6843 8283 6844 8284
rect 6859 8283 6872 8284
rect 6578 8244 6767 8274
rect 6593 8241 6767 8244
rect 6586 8238 6767 8241
rect 6395 8218 6408 8220
rect 6423 8218 6457 8220
rect 6395 8202 6469 8218
rect 6496 8214 6509 8228
rect 6524 8214 6540 8230
rect 6586 8225 6597 8238
rect 6379 8180 6380 8196
rect 6395 8180 6408 8202
rect 6423 8180 6453 8202
rect 6496 8198 6558 8214
rect 6586 8207 6597 8223
rect 6602 8218 6612 8238
rect 6622 8218 6636 8238
rect 6639 8225 6648 8238
rect 6664 8225 6673 8238
rect 6602 8207 6636 8218
rect 6639 8207 6648 8223
rect 6664 8207 6673 8223
rect 6680 8218 6690 8238
rect 6700 8218 6714 8238
rect 6715 8225 6726 8238
rect 6680 8207 6714 8218
rect 6715 8207 6726 8223
rect 6772 8214 6788 8230
rect 6795 8228 6825 8280
rect 6859 8276 6860 8283
rect 6844 8268 6860 8276
rect 6831 8236 6844 8255
rect 6859 8236 6889 8252
rect 6831 8220 6905 8236
rect 6831 8218 6844 8220
rect 6859 8218 6893 8220
rect 6496 8196 6509 8198
rect 6524 8196 6558 8198
rect 6496 8180 6558 8196
rect 6602 8191 6618 8194
rect 6680 8191 6710 8202
rect 6758 8198 6804 8214
rect 6831 8202 6905 8218
rect 6758 8196 6792 8198
rect 6757 8180 6804 8196
rect 6831 8180 6844 8202
rect 6859 8180 6889 8202
rect 6916 8180 6917 8196
rect 6932 8180 6945 8340
rect 6975 8236 6988 8340
rect 7033 8318 7034 8328
rect 7049 8318 7062 8328
rect 7033 8314 7062 8318
rect 7067 8314 7097 8340
rect 7115 8326 7131 8328
rect 7203 8326 7256 8340
rect 7204 8324 7268 8326
rect 7311 8324 7326 8340
rect 7375 8337 7405 8340
rect 7375 8334 7411 8337
rect 7341 8326 7357 8328
rect 7115 8314 7130 8318
rect 7033 8312 7130 8314
rect 7158 8312 7326 8324
rect 7342 8314 7357 8318
rect 7375 8315 7414 8334
rect 7433 8328 7440 8329
rect 7439 8321 7440 8328
rect 7423 8318 7424 8321
rect 7439 8318 7452 8321
rect 7375 8314 7405 8315
rect 7414 8314 7420 8315
rect 7423 8314 7452 8318
rect 7342 8313 7452 8314
rect 7342 8312 7458 8313
rect 7017 8304 7068 8312
rect 7017 8292 7042 8304
rect 7049 8292 7068 8304
rect 7099 8304 7149 8312
rect 7099 8296 7115 8304
rect 7122 8302 7149 8304
rect 7158 8302 7379 8312
rect 7122 8292 7379 8302
rect 7408 8304 7458 8312
rect 7408 8295 7424 8304
rect 7017 8284 7068 8292
rect 7115 8284 7379 8292
rect 7405 8292 7424 8295
rect 7431 8292 7458 8304
rect 7405 8284 7458 8292
rect 7033 8276 7034 8284
rect 7049 8276 7062 8284
rect 7033 8268 7049 8276
rect 7030 8261 7049 8264
rect 7030 8252 7052 8261
rect 7003 8242 7052 8252
rect 7003 8236 7033 8242
rect 7052 8237 7057 8242
rect 6975 8220 7049 8236
rect 7067 8228 7097 8284
rect 7132 8274 7340 8284
rect 7375 8280 7420 8284
rect 7423 8283 7424 8284
rect 7439 8283 7452 8284
rect 7158 8244 7347 8274
rect 7173 8241 7347 8244
rect 7166 8238 7347 8241
rect 6975 8218 6988 8220
rect 7003 8218 7037 8220
rect 6975 8202 7049 8218
rect 7076 8214 7089 8228
rect 7104 8214 7120 8230
rect 7166 8225 7177 8238
rect 6959 8180 6960 8196
rect 6975 8180 6988 8202
rect 7003 8180 7033 8202
rect 7076 8198 7138 8214
rect 7166 8207 7177 8223
rect 7182 8218 7192 8238
rect 7202 8218 7216 8238
rect 7219 8225 7228 8238
rect 7244 8225 7253 8238
rect 7182 8207 7216 8218
rect 7219 8207 7228 8223
rect 7244 8207 7253 8223
rect 7260 8218 7270 8238
rect 7280 8218 7294 8238
rect 7295 8225 7306 8238
rect 7260 8207 7294 8218
rect 7295 8207 7306 8223
rect 7352 8214 7368 8230
rect 7375 8228 7405 8280
rect 7439 8276 7440 8283
rect 7424 8268 7440 8276
rect 7411 8236 7424 8255
rect 7439 8236 7469 8252
rect 7411 8220 7485 8236
rect 7411 8218 7424 8220
rect 7439 8218 7473 8220
rect 7076 8196 7089 8198
rect 7104 8196 7138 8198
rect 7076 8180 7138 8196
rect 7182 8191 7198 8194
rect 7260 8191 7290 8202
rect 7338 8198 7384 8214
rect 7411 8202 7485 8218
rect 7338 8196 7372 8198
rect 7337 8180 7384 8196
rect 7411 8180 7424 8202
rect 7439 8180 7469 8202
rect 7496 8180 7497 8196
rect 7512 8180 7525 8340
rect 7555 8236 7568 8340
rect 7613 8318 7614 8328
rect 7629 8318 7642 8328
rect 7613 8314 7642 8318
rect 7647 8314 7677 8340
rect 7695 8326 7711 8328
rect 7783 8326 7836 8340
rect 7784 8324 7848 8326
rect 7891 8324 7906 8340
rect 7955 8337 7985 8340
rect 7955 8334 7991 8337
rect 7921 8326 7937 8328
rect 7695 8314 7710 8318
rect 7613 8312 7710 8314
rect 7738 8312 7906 8324
rect 7922 8314 7937 8318
rect 7955 8315 7994 8334
rect 8013 8328 8020 8329
rect 8019 8321 8020 8328
rect 8003 8318 8004 8321
rect 8019 8318 8032 8321
rect 7955 8314 7985 8315
rect 7994 8314 8000 8315
rect 8003 8314 8032 8318
rect 7922 8313 8032 8314
rect 7922 8312 8038 8313
rect 7597 8304 7648 8312
rect 7597 8292 7622 8304
rect 7629 8292 7648 8304
rect 7679 8304 7729 8312
rect 7679 8296 7695 8304
rect 7702 8302 7729 8304
rect 7738 8302 7959 8312
rect 7702 8292 7959 8302
rect 7988 8304 8038 8312
rect 7988 8295 8004 8304
rect 7597 8284 7648 8292
rect 7695 8284 7959 8292
rect 7985 8292 8004 8295
rect 8011 8292 8038 8304
rect 7985 8284 8038 8292
rect 7613 8276 7614 8284
rect 7629 8276 7642 8284
rect 7613 8268 7629 8276
rect 7610 8261 7629 8264
rect 7610 8252 7632 8261
rect 7583 8242 7632 8252
rect 7583 8236 7613 8242
rect 7632 8237 7637 8242
rect 7555 8220 7629 8236
rect 7647 8228 7677 8284
rect 7712 8274 7920 8284
rect 7955 8280 8000 8284
rect 8003 8283 8004 8284
rect 8019 8283 8032 8284
rect 7738 8244 7927 8274
rect 7753 8241 7927 8244
rect 7746 8238 7927 8241
rect 7555 8218 7568 8220
rect 7583 8218 7617 8220
rect 7555 8202 7629 8218
rect 7656 8214 7669 8228
rect 7684 8214 7700 8230
rect 7746 8225 7757 8238
rect 7539 8180 7540 8196
rect 7555 8180 7568 8202
rect 7583 8180 7613 8202
rect 7656 8198 7718 8214
rect 7746 8207 7757 8223
rect 7762 8218 7772 8238
rect 7782 8218 7796 8238
rect 7799 8225 7808 8238
rect 7824 8225 7833 8238
rect 7762 8207 7796 8218
rect 7799 8207 7808 8223
rect 7824 8207 7833 8223
rect 7840 8218 7850 8238
rect 7860 8218 7874 8238
rect 7875 8225 7886 8238
rect 7840 8207 7874 8218
rect 7875 8207 7886 8223
rect 7932 8214 7948 8230
rect 7955 8228 7985 8280
rect 8019 8276 8020 8283
rect 8004 8268 8020 8276
rect 7991 8236 8004 8255
rect 8019 8236 8049 8252
rect 7991 8220 8065 8236
rect 7991 8218 8004 8220
rect 8019 8218 8053 8220
rect 7656 8196 7669 8198
rect 7684 8196 7718 8198
rect 7656 8180 7718 8196
rect 7762 8191 7778 8194
rect 7840 8191 7870 8202
rect 7918 8198 7964 8214
rect 7991 8202 8065 8218
rect 7918 8196 7952 8198
rect 7917 8180 7964 8196
rect 7991 8180 8004 8202
rect 8019 8180 8049 8202
rect 8076 8180 8077 8196
rect 8092 8180 8105 8340
rect 8135 8236 8148 8340
rect 8193 8318 8194 8328
rect 8209 8318 8222 8328
rect 8193 8314 8222 8318
rect 8227 8314 8257 8340
rect 8275 8326 8291 8328
rect 8363 8326 8416 8340
rect 8364 8324 8428 8326
rect 8471 8324 8486 8340
rect 8535 8337 8565 8340
rect 8535 8334 8571 8337
rect 8501 8326 8517 8328
rect 8275 8314 8290 8318
rect 8193 8312 8290 8314
rect 8318 8312 8486 8324
rect 8502 8314 8517 8318
rect 8535 8315 8574 8334
rect 8593 8328 8600 8329
rect 8599 8321 8600 8328
rect 8583 8318 8584 8321
rect 8599 8318 8612 8321
rect 8535 8314 8565 8315
rect 8574 8314 8580 8315
rect 8583 8314 8612 8318
rect 8502 8313 8612 8314
rect 8502 8312 8618 8313
rect 8177 8304 8228 8312
rect 8177 8292 8202 8304
rect 8209 8292 8228 8304
rect 8259 8304 8309 8312
rect 8259 8296 8275 8304
rect 8282 8302 8309 8304
rect 8318 8302 8539 8312
rect 8282 8292 8539 8302
rect 8568 8304 8618 8312
rect 8568 8295 8584 8304
rect 8177 8284 8228 8292
rect 8275 8284 8539 8292
rect 8565 8292 8584 8295
rect 8591 8292 8618 8304
rect 8565 8284 8618 8292
rect 8193 8276 8194 8284
rect 8209 8276 8222 8284
rect 8193 8268 8209 8276
rect 8190 8261 8209 8264
rect 8190 8252 8212 8261
rect 8163 8242 8212 8252
rect 8163 8236 8193 8242
rect 8212 8237 8217 8242
rect 8135 8220 8209 8236
rect 8227 8228 8257 8284
rect 8292 8274 8500 8284
rect 8535 8280 8580 8284
rect 8583 8283 8584 8284
rect 8599 8283 8612 8284
rect 8318 8244 8507 8274
rect 8333 8241 8507 8244
rect 8326 8238 8507 8241
rect 8135 8218 8148 8220
rect 8163 8218 8197 8220
rect 8135 8202 8209 8218
rect 8236 8214 8249 8228
rect 8264 8214 8280 8230
rect 8326 8225 8337 8238
rect 8119 8180 8120 8196
rect 8135 8180 8148 8202
rect 8163 8180 8193 8202
rect 8236 8198 8298 8214
rect 8326 8207 8337 8223
rect 8342 8218 8352 8238
rect 8362 8218 8376 8238
rect 8379 8225 8388 8238
rect 8404 8225 8413 8238
rect 8342 8207 8376 8218
rect 8379 8207 8388 8223
rect 8404 8207 8413 8223
rect 8420 8218 8430 8238
rect 8440 8218 8454 8238
rect 8455 8225 8466 8238
rect 8420 8207 8454 8218
rect 8455 8207 8466 8223
rect 8512 8214 8528 8230
rect 8535 8228 8565 8280
rect 8599 8276 8600 8283
rect 8584 8268 8600 8276
rect 8571 8236 8584 8255
rect 8599 8236 8629 8252
rect 8571 8220 8645 8236
rect 8571 8218 8584 8220
rect 8599 8218 8633 8220
rect 8236 8196 8249 8198
rect 8264 8196 8298 8198
rect 8236 8180 8298 8196
rect 8342 8191 8358 8194
rect 8420 8191 8450 8202
rect 8498 8198 8544 8214
rect 8571 8202 8645 8218
rect 8498 8196 8532 8198
rect 8497 8180 8544 8196
rect 8571 8180 8584 8202
rect 8599 8180 8629 8202
rect 8656 8180 8657 8196
rect 8672 8180 8685 8340
rect 8715 8236 8728 8340
rect 8773 8318 8774 8328
rect 8789 8318 8802 8328
rect 8773 8314 8802 8318
rect 8807 8314 8837 8340
rect 8855 8326 8871 8328
rect 8943 8326 8996 8340
rect 8944 8324 9008 8326
rect 9051 8324 9066 8340
rect 9115 8337 9145 8340
rect 9115 8334 9151 8337
rect 9081 8326 9097 8328
rect 8855 8314 8870 8318
rect 8773 8312 8870 8314
rect 8898 8312 9066 8324
rect 9082 8314 9097 8318
rect 9115 8315 9154 8334
rect 9173 8328 9180 8329
rect 9179 8321 9180 8328
rect 9163 8318 9164 8321
rect 9179 8318 9192 8321
rect 9115 8314 9145 8315
rect 9154 8314 9160 8315
rect 9163 8314 9192 8318
rect 9082 8313 9192 8314
rect 9082 8312 9198 8313
rect 8757 8304 8808 8312
rect 8757 8292 8782 8304
rect 8789 8292 8808 8304
rect 8839 8304 8889 8312
rect 8839 8296 8855 8304
rect 8862 8302 8889 8304
rect 8898 8302 9119 8312
rect 8862 8292 9119 8302
rect 9148 8304 9198 8312
rect 9148 8295 9164 8304
rect 8757 8284 8808 8292
rect 8855 8284 9119 8292
rect 9145 8292 9164 8295
rect 9171 8292 9198 8304
rect 9145 8284 9198 8292
rect 8773 8276 8774 8284
rect 8789 8276 8802 8284
rect 8773 8268 8789 8276
rect 8770 8261 8789 8264
rect 8770 8252 8792 8261
rect 8743 8242 8792 8252
rect 8743 8236 8773 8242
rect 8792 8237 8797 8242
rect 8715 8220 8789 8236
rect 8807 8228 8837 8284
rect 8872 8274 9080 8284
rect 9115 8280 9160 8284
rect 9163 8283 9164 8284
rect 9179 8283 9192 8284
rect 8898 8244 9087 8274
rect 8913 8241 9087 8244
rect 8906 8238 9087 8241
rect 8715 8218 8728 8220
rect 8743 8218 8777 8220
rect 8715 8202 8789 8218
rect 8816 8214 8829 8228
rect 8844 8214 8860 8230
rect 8906 8225 8917 8238
rect 8699 8180 8700 8196
rect 8715 8180 8728 8202
rect 8743 8180 8773 8202
rect 8816 8198 8878 8214
rect 8906 8207 8917 8223
rect 8922 8218 8932 8238
rect 8942 8218 8956 8238
rect 8959 8225 8968 8238
rect 8984 8225 8993 8238
rect 8922 8207 8956 8218
rect 8959 8207 8968 8223
rect 8984 8207 8993 8223
rect 9000 8218 9010 8238
rect 9020 8218 9034 8238
rect 9035 8225 9046 8238
rect 9000 8207 9034 8218
rect 9035 8207 9046 8223
rect 9092 8214 9108 8230
rect 9115 8228 9145 8280
rect 9179 8276 9180 8283
rect 9164 8268 9180 8276
rect 9151 8236 9164 8255
rect 9179 8236 9209 8252
rect 9151 8220 9225 8236
rect 9151 8218 9164 8220
rect 9179 8218 9213 8220
rect 8816 8196 8829 8198
rect 8844 8196 8878 8198
rect 8816 8180 8878 8196
rect 8922 8191 8938 8194
rect 9000 8191 9030 8202
rect 9078 8198 9124 8214
rect 9151 8202 9225 8218
rect 9078 8196 9112 8198
rect 9077 8180 9124 8196
rect 9151 8180 9164 8202
rect 9179 8180 9209 8202
rect 9236 8180 9237 8196
rect 9252 8180 9265 8340
rect -7 8172 34 8180
rect -7 8146 8 8172
rect 15 8146 34 8172
rect 98 8168 160 8180
rect 172 8168 247 8180
rect 305 8168 380 8180
rect 392 8168 423 8180
rect 429 8168 464 8180
rect 98 8166 260 8168
rect -7 8138 34 8146
rect 116 8142 129 8166
rect 144 8164 159 8166
rect -1 8128 0 8138
rect 15 8128 28 8138
rect 43 8128 73 8142
rect 116 8128 159 8142
rect 183 8139 190 8146
rect 193 8142 260 8166
rect 292 8166 464 8168
rect 262 8144 290 8148
rect 292 8144 372 8166
rect 393 8164 408 8166
rect 262 8142 372 8144
rect 193 8138 372 8142
rect 166 8128 196 8138
rect 198 8128 351 8138
rect 359 8128 389 8138
rect 393 8128 423 8142
rect 451 8128 464 8166
rect 536 8172 571 8180
rect 536 8146 537 8172
rect 544 8146 571 8172
rect 479 8128 509 8142
rect 536 8138 571 8146
rect 573 8172 614 8180
rect 573 8146 588 8172
rect 595 8146 614 8172
rect 678 8168 740 8180
rect 752 8168 827 8180
rect 885 8168 960 8180
rect 972 8168 1003 8180
rect 1009 8168 1044 8180
rect 678 8166 840 8168
rect 573 8138 614 8146
rect 696 8142 709 8166
rect 724 8164 739 8166
rect 536 8128 537 8138
rect 552 8128 565 8138
rect 579 8128 580 8138
rect 595 8128 608 8138
rect 623 8128 653 8142
rect 696 8128 739 8142
rect 763 8139 770 8146
rect 773 8142 840 8166
rect 872 8166 1044 8168
rect 842 8144 870 8148
rect 872 8144 952 8166
rect 973 8164 988 8166
rect 842 8142 952 8144
rect 773 8138 952 8142
rect 746 8128 776 8138
rect 778 8128 931 8138
rect 939 8128 969 8138
rect 973 8128 1003 8142
rect 1031 8128 1044 8166
rect 1116 8172 1151 8180
rect 1116 8146 1117 8172
rect 1124 8146 1151 8172
rect 1059 8128 1089 8142
rect 1116 8138 1151 8146
rect 1153 8172 1194 8180
rect 1153 8146 1168 8172
rect 1175 8146 1194 8172
rect 1258 8168 1320 8180
rect 1332 8168 1407 8180
rect 1465 8168 1540 8180
rect 1552 8168 1583 8180
rect 1589 8168 1624 8180
rect 1258 8166 1420 8168
rect 1153 8138 1194 8146
rect 1276 8142 1289 8166
rect 1304 8164 1319 8166
rect 1116 8128 1117 8138
rect 1132 8128 1145 8138
rect 1159 8128 1160 8138
rect 1175 8128 1188 8138
rect 1203 8128 1233 8142
rect 1276 8128 1319 8142
rect 1343 8139 1350 8146
rect 1353 8142 1420 8166
rect 1452 8166 1624 8168
rect 1422 8144 1450 8148
rect 1452 8144 1532 8166
rect 1553 8164 1568 8166
rect 1422 8142 1532 8144
rect 1353 8138 1532 8142
rect 1326 8128 1356 8138
rect 1358 8128 1511 8138
rect 1519 8128 1549 8138
rect 1553 8128 1583 8142
rect 1611 8128 1624 8166
rect 1696 8172 1731 8180
rect 1696 8146 1697 8172
rect 1704 8146 1731 8172
rect 1639 8128 1669 8142
rect 1696 8138 1731 8146
rect 1733 8172 1774 8180
rect 1733 8146 1748 8172
rect 1755 8146 1774 8172
rect 1838 8168 1900 8180
rect 1912 8168 1987 8180
rect 2045 8168 2120 8180
rect 2132 8168 2163 8180
rect 2169 8168 2204 8180
rect 1838 8166 2000 8168
rect 1733 8138 1774 8146
rect 1856 8142 1869 8166
rect 1884 8164 1899 8166
rect 1696 8128 1697 8138
rect 1712 8128 1725 8138
rect 1739 8128 1740 8138
rect 1755 8128 1768 8138
rect 1783 8128 1813 8142
rect 1856 8128 1899 8142
rect 1923 8139 1930 8146
rect 1933 8142 2000 8166
rect 2032 8166 2204 8168
rect 2002 8144 2030 8148
rect 2032 8144 2112 8166
rect 2133 8164 2148 8166
rect 2002 8142 2112 8144
rect 1933 8138 2112 8142
rect 1906 8128 1936 8138
rect 1938 8128 2091 8138
rect 2099 8128 2129 8138
rect 2133 8128 2163 8142
rect 2191 8128 2204 8166
rect 2276 8172 2311 8180
rect 2276 8146 2277 8172
rect 2284 8146 2311 8172
rect 2219 8128 2249 8142
rect 2276 8138 2311 8146
rect 2313 8172 2354 8180
rect 2313 8146 2328 8172
rect 2335 8146 2354 8172
rect 2418 8168 2480 8180
rect 2492 8168 2567 8180
rect 2625 8168 2700 8180
rect 2712 8168 2743 8180
rect 2749 8168 2784 8180
rect 2418 8166 2580 8168
rect 2313 8138 2354 8146
rect 2436 8142 2449 8166
rect 2464 8164 2479 8166
rect 2276 8128 2277 8138
rect 2292 8128 2305 8138
rect 2319 8128 2320 8138
rect 2335 8128 2348 8138
rect 2363 8128 2393 8142
rect 2436 8128 2479 8142
rect 2503 8139 2510 8146
rect 2513 8142 2580 8166
rect 2612 8166 2784 8168
rect 2582 8144 2610 8148
rect 2612 8144 2692 8166
rect 2713 8164 2728 8166
rect 2582 8142 2692 8144
rect 2513 8138 2692 8142
rect 2486 8128 2516 8138
rect 2518 8128 2671 8138
rect 2679 8128 2709 8138
rect 2713 8128 2743 8142
rect 2771 8128 2784 8166
rect 2856 8172 2891 8180
rect 2856 8146 2857 8172
rect 2864 8146 2891 8172
rect 2799 8128 2829 8142
rect 2856 8138 2891 8146
rect 2893 8172 2934 8180
rect 2893 8146 2908 8172
rect 2915 8146 2934 8172
rect 2998 8168 3060 8180
rect 3072 8168 3147 8180
rect 3205 8168 3280 8180
rect 3292 8168 3323 8180
rect 3329 8168 3364 8180
rect 2998 8166 3160 8168
rect 2893 8138 2934 8146
rect 3016 8142 3029 8166
rect 3044 8164 3059 8166
rect 2856 8128 2857 8138
rect 2872 8128 2885 8138
rect 2899 8128 2900 8138
rect 2915 8128 2928 8138
rect 2943 8128 2973 8142
rect 3016 8128 3059 8142
rect 3083 8139 3090 8146
rect 3093 8142 3160 8166
rect 3192 8166 3364 8168
rect 3162 8144 3190 8148
rect 3192 8144 3272 8166
rect 3293 8164 3308 8166
rect 3162 8142 3272 8144
rect 3093 8138 3272 8142
rect 3066 8128 3096 8138
rect 3098 8128 3251 8138
rect 3259 8128 3289 8138
rect 3293 8128 3323 8142
rect 3351 8128 3364 8166
rect 3436 8172 3471 8180
rect 3436 8146 3437 8172
rect 3444 8146 3471 8172
rect 3379 8128 3409 8142
rect 3436 8138 3471 8146
rect 3473 8172 3514 8180
rect 3473 8146 3488 8172
rect 3495 8146 3514 8172
rect 3578 8168 3640 8180
rect 3652 8168 3727 8180
rect 3785 8168 3860 8180
rect 3872 8168 3903 8180
rect 3909 8168 3944 8180
rect 3578 8166 3740 8168
rect 3473 8138 3514 8146
rect 3596 8142 3609 8166
rect 3624 8164 3639 8166
rect 3436 8128 3437 8138
rect 3452 8128 3465 8138
rect 3479 8128 3480 8138
rect 3495 8128 3508 8138
rect 3523 8128 3553 8142
rect 3596 8128 3639 8142
rect 3663 8139 3670 8146
rect 3673 8142 3740 8166
rect 3772 8166 3944 8168
rect 3742 8144 3770 8148
rect 3772 8144 3852 8166
rect 3873 8164 3888 8166
rect 3742 8142 3852 8144
rect 3673 8138 3852 8142
rect 3646 8128 3676 8138
rect 3678 8128 3831 8138
rect 3839 8128 3869 8138
rect 3873 8128 3903 8142
rect 3931 8128 3944 8166
rect 4016 8172 4051 8180
rect 4016 8146 4017 8172
rect 4024 8146 4051 8172
rect 3959 8128 3989 8142
rect 4016 8138 4051 8146
rect 4053 8172 4094 8180
rect 4053 8146 4068 8172
rect 4075 8146 4094 8172
rect 4158 8168 4220 8180
rect 4232 8168 4307 8180
rect 4365 8168 4440 8180
rect 4452 8168 4483 8180
rect 4489 8168 4524 8180
rect 4158 8166 4320 8168
rect 4053 8138 4094 8146
rect 4176 8142 4189 8166
rect 4204 8164 4219 8166
rect 4016 8128 4017 8138
rect 4032 8128 4045 8138
rect 4059 8128 4060 8138
rect 4075 8128 4088 8138
rect 4103 8128 4133 8142
rect 4176 8128 4219 8142
rect 4243 8139 4250 8146
rect 4253 8142 4320 8166
rect 4352 8166 4524 8168
rect 4322 8144 4350 8148
rect 4352 8144 4432 8166
rect 4453 8164 4468 8166
rect 4322 8142 4432 8144
rect 4253 8138 4432 8142
rect 4226 8128 4256 8138
rect 4258 8128 4411 8138
rect 4419 8128 4449 8138
rect 4453 8128 4483 8142
rect 4511 8128 4524 8166
rect 4596 8172 4631 8180
rect 4596 8146 4597 8172
rect 4604 8146 4631 8172
rect 4539 8128 4569 8142
rect 4596 8138 4631 8146
rect 4633 8172 4674 8180
rect 4633 8146 4648 8172
rect 4655 8146 4674 8172
rect 4738 8168 4800 8180
rect 4812 8168 4887 8180
rect 4945 8168 5020 8180
rect 5032 8168 5063 8180
rect 5069 8168 5104 8180
rect 4738 8166 4900 8168
rect 4633 8138 4674 8146
rect 4756 8142 4769 8166
rect 4784 8164 4799 8166
rect 4596 8128 4597 8138
rect 4612 8128 4625 8138
rect 4639 8128 4640 8138
rect 4655 8128 4668 8138
rect 4683 8128 4713 8142
rect 4756 8128 4799 8142
rect 4823 8139 4830 8146
rect 4833 8142 4900 8166
rect 4932 8166 5104 8168
rect 4902 8144 4930 8148
rect 4932 8144 5012 8166
rect 5033 8164 5048 8166
rect 4902 8142 5012 8144
rect 4833 8138 5012 8142
rect 4806 8128 4836 8138
rect 4838 8128 4991 8138
rect 4999 8128 5029 8138
rect 5033 8128 5063 8142
rect 5091 8128 5104 8166
rect 5176 8172 5211 8180
rect 5176 8146 5177 8172
rect 5184 8146 5211 8172
rect 5119 8128 5149 8142
rect 5176 8138 5211 8146
rect 5213 8172 5254 8180
rect 5213 8146 5228 8172
rect 5235 8146 5254 8172
rect 5318 8168 5380 8180
rect 5392 8168 5467 8180
rect 5525 8168 5600 8180
rect 5612 8168 5643 8180
rect 5649 8168 5684 8180
rect 5318 8166 5480 8168
rect 5213 8138 5254 8146
rect 5336 8142 5349 8166
rect 5364 8164 5379 8166
rect 5176 8128 5177 8138
rect 5192 8128 5205 8138
rect 5219 8128 5220 8138
rect 5235 8128 5248 8138
rect 5263 8128 5293 8142
rect 5336 8128 5379 8142
rect 5403 8139 5410 8146
rect 5413 8142 5480 8166
rect 5512 8166 5684 8168
rect 5482 8144 5510 8148
rect 5512 8144 5592 8166
rect 5613 8164 5628 8166
rect 5482 8142 5592 8144
rect 5413 8138 5592 8142
rect 5386 8128 5416 8138
rect 5418 8128 5571 8138
rect 5579 8128 5609 8138
rect 5613 8128 5643 8142
rect 5671 8128 5684 8166
rect 5756 8172 5791 8180
rect 5756 8146 5757 8172
rect 5764 8146 5791 8172
rect 5699 8128 5729 8142
rect 5756 8138 5791 8146
rect 5793 8172 5834 8180
rect 5793 8146 5808 8172
rect 5815 8146 5834 8172
rect 5898 8168 5960 8180
rect 5972 8168 6047 8180
rect 6105 8168 6180 8180
rect 6192 8168 6223 8180
rect 6229 8168 6264 8180
rect 5898 8166 6060 8168
rect 5793 8138 5834 8146
rect 5916 8142 5929 8166
rect 5944 8164 5959 8166
rect 5756 8128 5757 8138
rect 5772 8128 5785 8138
rect 5799 8128 5800 8138
rect 5815 8128 5828 8138
rect 5843 8128 5873 8142
rect 5916 8128 5959 8142
rect 5983 8139 5990 8146
rect 5993 8142 6060 8166
rect 6092 8166 6264 8168
rect 6062 8144 6090 8148
rect 6092 8144 6172 8166
rect 6193 8164 6208 8166
rect 6062 8142 6172 8144
rect 5993 8138 6172 8142
rect 5966 8128 5996 8138
rect 5998 8128 6151 8138
rect 6159 8128 6189 8138
rect 6193 8128 6223 8142
rect 6251 8128 6264 8166
rect 6336 8172 6371 8180
rect 6336 8146 6337 8172
rect 6344 8146 6371 8172
rect 6279 8128 6309 8142
rect 6336 8138 6371 8146
rect 6373 8172 6414 8180
rect 6373 8146 6388 8172
rect 6395 8146 6414 8172
rect 6478 8168 6540 8180
rect 6552 8168 6627 8180
rect 6685 8168 6760 8180
rect 6772 8168 6803 8180
rect 6809 8168 6844 8180
rect 6478 8166 6640 8168
rect 6373 8138 6414 8146
rect 6496 8142 6509 8166
rect 6524 8164 6539 8166
rect 6336 8128 6337 8138
rect 6352 8128 6365 8138
rect 6379 8128 6380 8138
rect 6395 8128 6408 8138
rect 6423 8128 6453 8142
rect 6496 8128 6539 8142
rect 6563 8139 6570 8146
rect 6573 8142 6640 8166
rect 6672 8166 6844 8168
rect 6642 8144 6670 8148
rect 6672 8144 6752 8166
rect 6773 8164 6788 8166
rect 6642 8142 6752 8144
rect 6573 8138 6752 8142
rect 6546 8128 6576 8138
rect 6578 8128 6731 8138
rect 6739 8128 6769 8138
rect 6773 8128 6803 8142
rect 6831 8128 6844 8166
rect 6916 8172 6951 8180
rect 6916 8146 6917 8172
rect 6924 8146 6951 8172
rect 6859 8128 6889 8142
rect 6916 8138 6951 8146
rect 6953 8172 6994 8180
rect 6953 8146 6968 8172
rect 6975 8146 6994 8172
rect 7058 8168 7120 8180
rect 7132 8168 7207 8180
rect 7265 8168 7340 8180
rect 7352 8168 7383 8180
rect 7389 8168 7424 8180
rect 7058 8166 7220 8168
rect 6953 8138 6994 8146
rect 7076 8142 7089 8166
rect 7104 8164 7119 8166
rect 6916 8128 6917 8138
rect 6932 8128 6945 8138
rect 6959 8128 6960 8138
rect 6975 8128 6988 8138
rect 7003 8128 7033 8142
rect 7076 8128 7119 8142
rect 7143 8139 7150 8146
rect 7153 8142 7220 8166
rect 7252 8166 7424 8168
rect 7222 8144 7250 8148
rect 7252 8144 7332 8166
rect 7353 8164 7368 8166
rect 7222 8142 7332 8144
rect 7153 8138 7332 8142
rect 7126 8128 7156 8138
rect 7158 8128 7311 8138
rect 7319 8128 7349 8138
rect 7353 8128 7383 8142
rect 7411 8128 7424 8166
rect 7496 8172 7531 8180
rect 7496 8146 7497 8172
rect 7504 8146 7531 8172
rect 7439 8128 7469 8142
rect 7496 8138 7531 8146
rect 7533 8172 7574 8180
rect 7533 8146 7548 8172
rect 7555 8146 7574 8172
rect 7638 8168 7700 8180
rect 7712 8168 7787 8180
rect 7845 8168 7920 8180
rect 7932 8168 7963 8180
rect 7969 8168 8004 8180
rect 7638 8166 7800 8168
rect 7533 8138 7574 8146
rect 7656 8142 7669 8166
rect 7684 8164 7699 8166
rect 7496 8128 7497 8138
rect 7512 8128 7525 8138
rect 7539 8128 7540 8138
rect 7555 8128 7568 8138
rect 7583 8128 7613 8142
rect 7656 8128 7699 8142
rect 7723 8139 7730 8146
rect 7733 8142 7800 8166
rect 7832 8166 8004 8168
rect 7802 8144 7830 8148
rect 7832 8144 7912 8166
rect 7933 8164 7948 8166
rect 7802 8142 7912 8144
rect 7733 8138 7912 8142
rect 7706 8128 7736 8138
rect 7738 8128 7891 8138
rect 7899 8128 7929 8138
rect 7933 8128 7963 8142
rect 7991 8128 8004 8166
rect 8076 8172 8111 8180
rect 8076 8146 8077 8172
rect 8084 8146 8111 8172
rect 8019 8128 8049 8142
rect 8076 8138 8111 8146
rect 8113 8172 8154 8180
rect 8113 8146 8128 8172
rect 8135 8146 8154 8172
rect 8218 8168 8280 8180
rect 8292 8168 8367 8180
rect 8425 8168 8500 8180
rect 8512 8168 8543 8180
rect 8549 8168 8584 8180
rect 8218 8166 8380 8168
rect 8113 8138 8154 8146
rect 8236 8142 8249 8166
rect 8264 8164 8279 8166
rect 8076 8128 8077 8138
rect 8092 8128 8105 8138
rect 8119 8128 8120 8138
rect 8135 8128 8148 8138
rect 8163 8128 8193 8142
rect 8236 8128 8279 8142
rect 8303 8139 8310 8146
rect 8313 8142 8380 8166
rect 8412 8166 8584 8168
rect 8382 8144 8410 8148
rect 8412 8144 8492 8166
rect 8513 8164 8528 8166
rect 8382 8142 8492 8144
rect 8313 8138 8492 8142
rect 8286 8128 8316 8138
rect 8318 8128 8471 8138
rect 8479 8128 8509 8138
rect 8513 8128 8543 8142
rect 8571 8128 8584 8166
rect 8656 8172 8691 8180
rect 8656 8146 8657 8172
rect 8664 8146 8691 8172
rect 8599 8128 8629 8142
rect 8656 8138 8691 8146
rect 8693 8172 8734 8180
rect 8693 8146 8708 8172
rect 8715 8146 8734 8172
rect 8798 8168 8860 8180
rect 8872 8168 8947 8180
rect 9005 8168 9080 8180
rect 9092 8168 9123 8180
rect 9129 8168 9164 8180
rect 8798 8166 8960 8168
rect 8693 8138 8734 8146
rect 8816 8142 8829 8166
rect 8844 8164 8859 8166
rect 8656 8128 8657 8138
rect 8672 8128 8685 8138
rect 8699 8128 8700 8138
rect 8715 8128 8728 8138
rect 8743 8128 8773 8142
rect 8816 8128 8859 8142
rect 8883 8139 8890 8146
rect 8893 8142 8960 8166
rect 8992 8166 9164 8168
rect 8962 8144 8990 8148
rect 8992 8144 9072 8166
rect 9093 8164 9108 8166
rect 8962 8142 9072 8144
rect 8893 8138 9072 8142
rect 8866 8128 8896 8138
rect 8898 8128 9051 8138
rect 9059 8128 9089 8138
rect 9093 8128 9123 8142
rect 9151 8128 9164 8166
rect 9236 8172 9271 8180
rect 9236 8146 9237 8172
rect 9244 8146 9271 8172
rect 9179 8128 9209 8142
rect 9236 8138 9271 8146
rect 9236 8128 9237 8138
rect 9252 8128 9265 8138
rect -1 8122 9265 8128
rect 0 8114 9265 8122
rect 15 8084 28 8114
rect 43 8096 73 8114
rect 116 8100 130 8114
rect 166 8100 386 8114
rect 117 8098 130 8100
rect 83 8086 98 8098
rect 80 8084 102 8086
rect 107 8084 137 8098
rect 198 8096 351 8100
rect 180 8084 372 8096
rect 415 8084 445 8098
rect 451 8084 464 8114
rect 479 8096 509 8114
rect 552 8084 565 8114
rect 595 8084 608 8114
rect 623 8096 653 8114
rect 696 8100 710 8114
rect 746 8100 966 8114
rect 697 8098 710 8100
rect 663 8086 678 8098
rect 660 8084 682 8086
rect 687 8084 717 8098
rect 778 8096 931 8100
rect 760 8084 952 8096
rect 995 8084 1025 8098
rect 1031 8084 1044 8114
rect 1059 8096 1089 8114
rect 1132 8084 1145 8114
rect 1175 8084 1188 8114
rect 1203 8096 1233 8114
rect 1276 8100 1290 8114
rect 1326 8100 1546 8114
rect 1277 8098 1290 8100
rect 1243 8086 1258 8098
rect 1240 8084 1262 8086
rect 1267 8084 1297 8098
rect 1358 8096 1511 8100
rect 1340 8084 1532 8096
rect 1575 8084 1605 8098
rect 1611 8084 1624 8114
rect 1639 8096 1669 8114
rect 1712 8084 1725 8114
rect 1755 8084 1768 8114
rect 1783 8096 1813 8114
rect 1856 8100 1870 8114
rect 1906 8100 2126 8114
rect 1857 8098 1870 8100
rect 1823 8086 1838 8098
rect 1820 8084 1842 8086
rect 1847 8084 1877 8098
rect 1938 8096 2091 8100
rect 1920 8084 2112 8096
rect 2155 8084 2185 8098
rect 2191 8084 2204 8114
rect 2219 8096 2249 8114
rect 2292 8084 2305 8114
rect 2335 8084 2348 8114
rect 2363 8096 2393 8114
rect 2436 8100 2450 8114
rect 2486 8100 2706 8114
rect 2437 8098 2450 8100
rect 2403 8086 2418 8098
rect 2400 8084 2422 8086
rect 2427 8084 2457 8098
rect 2518 8096 2671 8100
rect 2500 8084 2692 8096
rect 2735 8084 2765 8098
rect 2771 8084 2784 8114
rect 2799 8096 2829 8114
rect 2872 8084 2885 8114
rect 2915 8084 2928 8114
rect 2943 8096 2973 8114
rect 3016 8100 3030 8114
rect 3066 8100 3286 8114
rect 3017 8098 3030 8100
rect 2983 8086 2998 8098
rect 2980 8084 3002 8086
rect 3007 8084 3037 8098
rect 3098 8096 3251 8100
rect 3080 8084 3272 8096
rect 3315 8084 3345 8098
rect 3351 8084 3364 8114
rect 3379 8096 3409 8114
rect 3452 8084 3465 8114
rect 3495 8084 3508 8114
rect 3523 8096 3553 8114
rect 3596 8100 3610 8114
rect 3646 8100 3866 8114
rect 3597 8098 3610 8100
rect 3563 8086 3578 8098
rect 3560 8084 3582 8086
rect 3587 8084 3617 8098
rect 3678 8096 3831 8100
rect 3660 8084 3852 8096
rect 3895 8084 3925 8098
rect 3931 8084 3944 8114
rect 3959 8096 3989 8114
rect 4032 8084 4045 8114
rect 4075 8084 4088 8114
rect 4103 8096 4133 8114
rect 4176 8100 4190 8114
rect 4226 8100 4446 8114
rect 4177 8098 4190 8100
rect 4143 8086 4158 8098
rect 4140 8084 4162 8086
rect 4167 8084 4197 8098
rect 4258 8096 4411 8100
rect 4240 8084 4432 8096
rect 4475 8084 4505 8098
rect 4511 8084 4524 8114
rect 4539 8096 4569 8114
rect 4612 8084 4625 8114
rect 4655 8084 4668 8114
rect 4683 8096 4713 8114
rect 4756 8100 4770 8114
rect 4806 8100 5026 8114
rect 4757 8098 4770 8100
rect 4723 8086 4738 8098
rect 4720 8084 4742 8086
rect 4747 8084 4777 8098
rect 4838 8096 4991 8100
rect 4820 8084 5012 8096
rect 5055 8084 5085 8098
rect 5091 8084 5104 8114
rect 5119 8096 5149 8114
rect 5192 8084 5205 8114
rect 5235 8084 5248 8114
rect 5263 8096 5293 8114
rect 5336 8100 5350 8114
rect 5386 8100 5606 8114
rect 5337 8098 5350 8100
rect 5303 8086 5318 8098
rect 5300 8084 5322 8086
rect 5327 8084 5357 8098
rect 5418 8096 5571 8100
rect 5400 8084 5592 8096
rect 5635 8084 5665 8098
rect 5671 8084 5684 8114
rect 5699 8096 5729 8114
rect 5772 8084 5785 8114
rect 5815 8084 5828 8114
rect 5843 8096 5873 8114
rect 5916 8100 5930 8114
rect 5966 8100 6186 8114
rect 5917 8098 5930 8100
rect 5883 8086 5898 8098
rect 5880 8084 5902 8086
rect 5907 8084 5937 8098
rect 5998 8096 6151 8100
rect 5980 8084 6172 8096
rect 6215 8084 6245 8098
rect 6251 8084 6264 8114
rect 6279 8096 6309 8114
rect 6352 8084 6365 8114
rect 6395 8084 6408 8114
rect 6423 8096 6453 8114
rect 6496 8100 6510 8114
rect 6546 8100 6766 8114
rect 6497 8098 6510 8100
rect 6463 8086 6478 8098
rect 6460 8084 6482 8086
rect 6487 8084 6517 8098
rect 6578 8096 6731 8100
rect 6560 8084 6752 8096
rect 6795 8084 6825 8098
rect 6831 8084 6844 8114
rect 6859 8096 6889 8114
rect 6932 8084 6945 8114
rect 6975 8084 6988 8114
rect 7003 8096 7033 8114
rect 7076 8100 7090 8114
rect 7126 8100 7346 8114
rect 7077 8098 7090 8100
rect 7043 8086 7058 8098
rect 7040 8084 7062 8086
rect 7067 8084 7097 8098
rect 7158 8096 7311 8100
rect 7140 8084 7332 8096
rect 7375 8084 7405 8098
rect 7411 8084 7424 8114
rect 7439 8096 7469 8114
rect 7512 8084 7525 8114
rect 7555 8084 7568 8114
rect 7583 8096 7613 8114
rect 7656 8100 7670 8114
rect 7706 8100 7926 8114
rect 7657 8098 7670 8100
rect 7623 8086 7638 8098
rect 7620 8084 7642 8086
rect 7647 8084 7677 8098
rect 7738 8096 7891 8100
rect 7720 8084 7912 8096
rect 7955 8084 7985 8098
rect 7991 8084 8004 8114
rect 8019 8096 8049 8114
rect 8092 8084 8105 8114
rect 8135 8084 8148 8114
rect 8163 8096 8193 8114
rect 8236 8100 8250 8114
rect 8286 8100 8506 8114
rect 8237 8098 8250 8100
rect 8203 8086 8218 8098
rect 8200 8084 8222 8086
rect 8227 8084 8257 8098
rect 8318 8096 8471 8100
rect 8300 8084 8492 8096
rect 8535 8084 8565 8098
rect 8571 8084 8584 8114
rect 8599 8096 8629 8114
rect 8672 8084 8685 8114
rect 8715 8084 8728 8114
rect 8743 8096 8773 8114
rect 8816 8100 8830 8114
rect 8866 8100 9086 8114
rect 8817 8098 8830 8100
rect 8783 8086 8798 8098
rect 8780 8084 8802 8086
rect 8807 8084 8837 8098
rect 8898 8096 9051 8100
rect 8880 8084 9072 8096
rect 9115 8084 9145 8098
rect 9151 8084 9164 8114
rect 9179 8096 9209 8114
rect 9252 8084 9265 8114
rect 0 8070 9265 8084
rect 15 7966 28 8070
rect 73 8048 74 8058
rect 89 8048 102 8058
rect 73 8044 102 8048
rect 107 8044 137 8070
rect 155 8056 171 8058
rect 243 8056 296 8070
rect 244 8054 308 8056
rect 351 8054 366 8070
rect 415 8067 445 8070
rect 415 8064 451 8067
rect 381 8056 397 8058
rect 155 8044 170 8048
rect 73 8042 170 8044
rect 198 8042 366 8054
rect 382 8044 397 8048
rect 415 8045 454 8064
rect 473 8058 480 8059
rect 479 8051 480 8058
rect 463 8048 464 8051
rect 479 8048 492 8051
rect 415 8044 445 8045
rect 454 8044 460 8045
rect 463 8044 492 8048
rect 382 8043 492 8044
rect 382 8042 498 8043
rect 57 8034 108 8042
rect 57 8022 82 8034
rect 89 8022 108 8034
rect 139 8034 189 8042
rect 139 8026 155 8034
rect 162 8032 189 8034
rect 198 8032 419 8042
rect 162 8022 419 8032
rect 448 8034 498 8042
rect 448 8025 464 8034
rect 57 8014 108 8022
rect 155 8014 419 8022
rect 445 8022 464 8025
rect 471 8022 498 8034
rect 445 8014 498 8022
rect 73 8006 74 8014
rect 89 8006 102 8014
rect 73 7998 89 8006
rect 70 7991 89 7994
rect 70 7982 92 7991
rect 43 7972 92 7982
rect 43 7966 73 7972
rect 92 7967 97 7972
rect 15 7950 89 7966
rect 107 7958 137 8014
rect 172 8004 380 8014
rect 415 8010 460 8014
rect 463 8013 464 8014
rect 479 8013 492 8014
rect 198 7974 387 8004
rect 213 7971 387 7974
rect 206 7968 387 7971
rect 15 7948 28 7950
rect 43 7948 77 7950
rect 15 7932 89 7948
rect 116 7944 129 7958
rect 144 7944 160 7960
rect 206 7955 217 7968
rect -1 7910 0 7926
rect 15 7910 28 7932
rect 43 7910 73 7932
rect 116 7928 178 7944
rect 206 7937 217 7953
rect 222 7948 232 7968
rect 242 7948 256 7968
rect 259 7955 268 7968
rect 284 7955 293 7968
rect 222 7937 256 7948
rect 259 7937 268 7953
rect 284 7937 293 7953
rect 300 7948 310 7968
rect 320 7948 334 7968
rect 335 7955 346 7968
rect 300 7937 334 7948
rect 335 7937 346 7953
rect 392 7944 408 7960
rect 415 7958 445 8010
rect 479 8006 480 8013
rect 464 7998 480 8006
rect 451 7966 464 7985
rect 479 7966 509 7982
rect 451 7950 525 7966
rect 451 7948 464 7950
rect 479 7948 513 7950
rect 116 7926 129 7928
rect 144 7926 178 7928
rect 116 7910 178 7926
rect 222 7921 238 7924
rect 300 7921 330 7932
rect 378 7928 424 7944
rect 451 7932 525 7948
rect 378 7926 412 7928
rect 377 7910 424 7926
rect 451 7910 464 7932
rect 479 7910 509 7932
rect 536 7910 537 7926
rect 552 7910 565 8070
rect 595 7966 608 8070
rect 653 8048 654 8058
rect 669 8048 682 8058
rect 653 8044 682 8048
rect 687 8044 717 8070
rect 735 8056 751 8058
rect 823 8056 876 8070
rect 824 8054 888 8056
rect 931 8054 946 8070
rect 995 8067 1025 8070
rect 995 8064 1031 8067
rect 961 8056 977 8058
rect 735 8044 750 8048
rect 653 8042 750 8044
rect 778 8042 946 8054
rect 962 8044 977 8048
rect 995 8045 1034 8064
rect 1053 8058 1060 8059
rect 1059 8051 1060 8058
rect 1043 8048 1044 8051
rect 1059 8048 1072 8051
rect 995 8044 1025 8045
rect 1034 8044 1040 8045
rect 1043 8044 1072 8048
rect 962 8043 1072 8044
rect 962 8042 1078 8043
rect 637 8034 688 8042
rect 637 8022 662 8034
rect 669 8022 688 8034
rect 719 8034 769 8042
rect 719 8026 735 8034
rect 742 8032 769 8034
rect 778 8032 999 8042
rect 742 8022 999 8032
rect 1028 8034 1078 8042
rect 1028 8025 1044 8034
rect 637 8014 688 8022
rect 735 8014 999 8022
rect 1025 8022 1044 8025
rect 1051 8022 1078 8034
rect 1025 8014 1078 8022
rect 653 8006 654 8014
rect 669 8006 682 8014
rect 653 7998 669 8006
rect 650 7991 669 7994
rect 650 7982 672 7991
rect 623 7972 672 7982
rect 623 7966 653 7972
rect 672 7967 677 7972
rect 595 7950 669 7966
rect 687 7958 717 8014
rect 752 8004 960 8014
rect 995 8010 1040 8014
rect 1043 8013 1044 8014
rect 1059 8013 1072 8014
rect 778 7974 967 8004
rect 793 7971 967 7974
rect 786 7968 967 7971
rect 595 7948 608 7950
rect 623 7948 657 7950
rect 595 7932 669 7948
rect 696 7944 709 7958
rect 724 7944 740 7960
rect 786 7955 797 7968
rect 579 7910 580 7926
rect 595 7910 608 7932
rect 623 7910 653 7932
rect 696 7928 758 7944
rect 786 7937 797 7953
rect 802 7948 812 7968
rect 822 7948 836 7968
rect 839 7955 848 7968
rect 864 7955 873 7968
rect 802 7937 836 7948
rect 839 7937 848 7953
rect 864 7937 873 7953
rect 880 7948 890 7968
rect 900 7948 914 7968
rect 915 7955 926 7968
rect 880 7937 914 7948
rect 915 7937 926 7953
rect 972 7944 988 7960
rect 995 7958 1025 8010
rect 1059 8006 1060 8013
rect 1044 7998 1060 8006
rect 1031 7966 1044 7985
rect 1059 7966 1089 7982
rect 1031 7950 1105 7966
rect 1031 7948 1044 7950
rect 1059 7948 1093 7950
rect 696 7926 709 7928
rect 724 7926 758 7928
rect 696 7910 758 7926
rect 802 7921 818 7924
rect 880 7921 910 7932
rect 958 7928 1004 7944
rect 1031 7932 1105 7948
rect 958 7926 992 7928
rect 957 7910 1004 7926
rect 1031 7910 1044 7932
rect 1059 7910 1089 7932
rect 1116 7910 1117 7926
rect 1132 7910 1145 8070
rect 1175 7966 1188 8070
rect 1233 8048 1234 8058
rect 1249 8048 1262 8058
rect 1233 8044 1262 8048
rect 1267 8044 1297 8070
rect 1315 8056 1331 8058
rect 1403 8056 1456 8070
rect 1404 8054 1468 8056
rect 1511 8054 1526 8070
rect 1575 8067 1605 8070
rect 1575 8064 1611 8067
rect 1541 8056 1557 8058
rect 1315 8044 1330 8048
rect 1233 8042 1330 8044
rect 1358 8042 1526 8054
rect 1542 8044 1557 8048
rect 1575 8045 1614 8064
rect 1633 8058 1640 8059
rect 1639 8051 1640 8058
rect 1623 8048 1624 8051
rect 1639 8048 1652 8051
rect 1575 8044 1605 8045
rect 1614 8044 1620 8045
rect 1623 8044 1652 8048
rect 1542 8043 1652 8044
rect 1542 8042 1658 8043
rect 1217 8034 1268 8042
rect 1217 8022 1242 8034
rect 1249 8022 1268 8034
rect 1299 8034 1349 8042
rect 1299 8026 1315 8034
rect 1322 8032 1349 8034
rect 1358 8032 1579 8042
rect 1322 8022 1579 8032
rect 1608 8034 1658 8042
rect 1608 8025 1624 8034
rect 1217 8014 1268 8022
rect 1315 8014 1579 8022
rect 1605 8022 1624 8025
rect 1631 8022 1658 8034
rect 1605 8014 1658 8022
rect 1233 8006 1234 8014
rect 1249 8006 1262 8014
rect 1233 7998 1249 8006
rect 1230 7991 1249 7994
rect 1230 7982 1252 7991
rect 1203 7972 1252 7982
rect 1203 7966 1233 7972
rect 1252 7967 1257 7972
rect 1175 7950 1249 7966
rect 1267 7958 1297 8014
rect 1332 8004 1540 8014
rect 1575 8010 1620 8014
rect 1623 8013 1624 8014
rect 1639 8013 1652 8014
rect 1358 7974 1547 8004
rect 1373 7971 1547 7974
rect 1366 7968 1547 7971
rect 1175 7948 1188 7950
rect 1203 7948 1237 7950
rect 1175 7932 1249 7948
rect 1276 7944 1289 7958
rect 1304 7944 1320 7960
rect 1366 7955 1377 7968
rect 1159 7910 1160 7926
rect 1175 7910 1188 7932
rect 1203 7910 1233 7932
rect 1276 7928 1338 7944
rect 1366 7937 1377 7953
rect 1382 7948 1392 7968
rect 1402 7948 1416 7968
rect 1419 7955 1428 7968
rect 1444 7955 1453 7968
rect 1382 7937 1416 7948
rect 1419 7937 1428 7953
rect 1444 7937 1453 7953
rect 1460 7948 1470 7968
rect 1480 7948 1494 7968
rect 1495 7955 1506 7968
rect 1460 7937 1494 7948
rect 1495 7937 1506 7953
rect 1552 7944 1568 7960
rect 1575 7958 1605 8010
rect 1639 8006 1640 8013
rect 1624 7998 1640 8006
rect 1611 7966 1624 7985
rect 1639 7966 1669 7982
rect 1611 7950 1685 7966
rect 1611 7948 1624 7950
rect 1639 7948 1673 7950
rect 1276 7926 1289 7928
rect 1304 7926 1338 7928
rect 1276 7910 1338 7926
rect 1382 7921 1398 7924
rect 1460 7921 1490 7932
rect 1538 7928 1584 7944
rect 1611 7932 1685 7948
rect 1538 7926 1572 7928
rect 1537 7910 1584 7926
rect 1611 7910 1624 7932
rect 1639 7910 1669 7932
rect 1696 7910 1697 7926
rect 1712 7910 1725 8070
rect 1755 7966 1768 8070
rect 1813 8048 1814 8058
rect 1829 8048 1842 8058
rect 1813 8044 1842 8048
rect 1847 8044 1877 8070
rect 1895 8056 1911 8058
rect 1983 8056 2036 8070
rect 1984 8054 2048 8056
rect 2091 8054 2106 8070
rect 2155 8067 2185 8070
rect 2155 8064 2191 8067
rect 2121 8056 2137 8058
rect 1895 8044 1910 8048
rect 1813 8042 1910 8044
rect 1938 8042 2106 8054
rect 2122 8044 2137 8048
rect 2155 8045 2194 8064
rect 2213 8058 2220 8059
rect 2219 8051 2220 8058
rect 2203 8048 2204 8051
rect 2219 8048 2232 8051
rect 2155 8044 2185 8045
rect 2194 8044 2200 8045
rect 2203 8044 2232 8048
rect 2122 8043 2232 8044
rect 2122 8042 2238 8043
rect 1797 8034 1848 8042
rect 1797 8022 1822 8034
rect 1829 8022 1848 8034
rect 1879 8034 1929 8042
rect 1879 8026 1895 8034
rect 1902 8032 1929 8034
rect 1938 8032 2159 8042
rect 1902 8022 2159 8032
rect 2188 8034 2238 8042
rect 2188 8025 2204 8034
rect 1797 8014 1848 8022
rect 1895 8014 2159 8022
rect 2185 8022 2204 8025
rect 2211 8022 2238 8034
rect 2185 8014 2238 8022
rect 1813 8006 1814 8014
rect 1829 8006 1842 8014
rect 1813 7998 1829 8006
rect 1810 7991 1829 7994
rect 1810 7982 1832 7991
rect 1783 7972 1832 7982
rect 1783 7966 1813 7972
rect 1832 7967 1837 7972
rect 1755 7950 1829 7966
rect 1847 7958 1877 8014
rect 1912 8004 2120 8014
rect 2155 8010 2200 8014
rect 2203 8013 2204 8014
rect 2219 8013 2232 8014
rect 1938 7974 2127 8004
rect 1953 7971 2127 7974
rect 1946 7968 2127 7971
rect 1755 7948 1768 7950
rect 1783 7948 1817 7950
rect 1755 7932 1829 7948
rect 1856 7944 1869 7958
rect 1884 7944 1900 7960
rect 1946 7955 1957 7968
rect 1739 7910 1740 7926
rect 1755 7910 1768 7932
rect 1783 7910 1813 7932
rect 1856 7928 1918 7944
rect 1946 7937 1957 7953
rect 1962 7948 1972 7968
rect 1982 7948 1996 7968
rect 1999 7955 2008 7968
rect 2024 7955 2033 7968
rect 1962 7937 1996 7948
rect 1999 7937 2008 7953
rect 2024 7937 2033 7953
rect 2040 7948 2050 7968
rect 2060 7948 2074 7968
rect 2075 7955 2086 7968
rect 2040 7937 2074 7948
rect 2075 7937 2086 7953
rect 2132 7944 2148 7960
rect 2155 7958 2185 8010
rect 2219 8006 2220 8013
rect 2204 7998 2220 8006
rect 2191 7966 2204 7985
rect 2219 7966 2249 7982
rect 2191 7950 2265 7966
rect 2191 7948 2204 7950
rect 2219 7948 2253 7950
rect 1856 7926 1869 7928
rect 1884 7926 1918 7928
rect 1856 7910 1918 7926
rect 1962 7921 1976 7924
rect 2040 7921 2070 7932
rect 2118 7928 2164 7944
rect 2191 7932 2265 7948
rect 2118 7926 2152 7928
rect 2117 7910 2164 7926
rect 2191 7910 2204 7932
rect 2219 7910 2249 7932
rect 2276 7910 2277 7926
rect 2292 7910 2305 8070
rect 2335 7966 2348 8070
rect 2393 8048 2394 8058
rect 2409 8048 2422 8058
rect 2393 8044 2422 8048
rect 2427 8044 2457 8070
rect 2475 8056 2491 8058
rect 2563 8056 2616 8070
rect 2564 8054 2628 8056
rect 2671 8054 2686 8070
rect 2735 8067 2765 8070
rect 2735 8064 2771 8067
rect 2701 8056 2717 8058
rect 2475 8044 2490 8048
rect 2393 8042 2490 8044
rect 2518 8042 2686 8054
rect 2702 8044 2717 8048
rect 2735 8045 2774 8064
rect 2793 8058 2800 8059
rect 2799 8051 2800 8058
rect 2783 8048 2784 8051
rect 2799 8048 2812 8051
rect 2735 8044 2765 8045
rect 2774 8044 2780 8045
rect 2783 8044 2812 8048
rect 2702 8043 2812 8044
rect 2702 8042 2818 8043
rect 2377 8034 2428 8042
rect 2377 8022 2402 8034
rect 2409 8022 2428 8034
rect 2459 8034 2509 8042
rect 2459 8026 2475 8034
rect 2482 8032 2509 8034
rect 2518 8032 2739 8042
rect 2482 8022 2739 8032
rect 2768 8034 2818 8042
rect 2768 8025 2784 8034
rect 2377 8014 2428 8022
rect 2475 8014 2739 8022
rect 2765 8022 2784 8025
rect 2791 8022 2818 8034
rect 2765 8014 2818 8022
rect 2393 8006 2394 8014
rect 2409 8006 2422 8014
rect 2393 7998 2409 8006
rect 2390 7991 2409 7994
rect 2390 7982 2412 7991
rect 2363 7972 2412 7982
rect 2363 7966 2393 7972
rect 2412 7967 2417 7972
rect 2335 7950 2409 7966
rect 2427 7958 2457 8014
rect 2492 8004 2700 8014
rect 2735 8010 2780 8014
rect 2783 8013 2784 8014
rect 2799 8013 2812 8014
rect 2518 7974 2707 8004
rect 2533 7971 2707 7974
rect 2526 7968 2707 7971
rect 2335 7948 2348 7950
rect 2363 7948 2397 7950
rect 2335 7932 2409 7948
rect 2436 7944 2449 7958
rect 2464 7944 2480 7960
rect 2526 7955 2537 7968
rect 2319 7910 2320 7926
rect 2335 7910 2348 7932
rect 2363 7910 2393 7932
rect 2436 7928 2498 7944
rect 2526 7937 2537 7953
rect 2542 7948 2552 7968
rect 2562 7948 2576 7968
rect 2579 7955 2588 7968
rect 2604 7955 2613 7968
rect 2542 7937 2576 7948
rect 2579 7937 2588 7953
rect 2604 7937 2613 7953
rect 2620 7948 2630 7968
rect 2640 7948 2654 7968
rect 2655 7955 2666 7968
rect 2620 7937 2654 7948
rect 2655 7937 2666 7953
rect 2712 7944 2728 7960
rect 2735 7958 2765 8010
rect 2799 8006 2800 8013
rect 2784 7998 2800 8006
rect 2771 7966 2784 7985
rect 2799 7966 2829 7982
rect 2771 7950 2845 7966
rect 2771 7948 2784 7950
rect 2799 7948 2833 7950
rect 2436 7926 2449 7928
rect 2464 7926 2498 7928
rect 2436 7910 2498 7926
rect 2542 7921 2558 7924
rect 2620 7921 2650 7932
rect 2698 7928 2744 7944
rect 2771 7932 2845 7948
rect 2698 7926 2732 7928
rect 2697 7910 2744 7926
rect 2771 7910 2784 7932
rect 2799 7910 2829 7932
rect 2856 7910 2857 7926
rect 2872 7910 2885 8070
rect 2915 7966 2928 8070
rect 2973 8048 2974 8058
rect 2989 8048 3002 8058
rect 2973 8044 3002 8048
rect 3007 8044 3037 8070
rect 3055 8056 3071 8058
rect 3143 8056 3196 8070
rect 3144 8054 3208 8056
rect 3251 8054 3266 8070
rect 3315 8067 3345 8070
rect 3315 8064 3351 8067
rect 3281 8056 3297 8058
rect 3055 8044 3070 8048
rect 2973 8042 3070 8044
rect 3098 8042 3266 8054
rect 3282 8044 3297 8048
rect 3315 8045 3354 8064
rect 3373 8058 3380 8059
rect 3379 8051 3380 8058
rect 3363 8048 3364 8051
rect 3379 8048 3392 8051
rect 3315 8044 3345 8045
rect 3354 8044 3360 8045
rect 3363 8044 3392 8048
rect 3282 8043 3392 8044
rect 3282 8042 3398 8043
rect 2957 8034 3008 8042
rect 2957 8022 2982 8034
rect 2989 8022 3008 8034
rect 3039 8034 3089 8042
rect 3039 8026 3055 8034
rect 3062 8032 3089 8034
rect 3098 8032 3319 8042
rect 3062 8022 3319 8032
rect 3348 8034 3398 8042
rect 3348 8025 3364 8034
rect 2957 8014 3008 8022
rect 3055 8014 3319 8022
rect 3345 8022 3364 8025
rect 3371 8022 3398 8034
rect 3345 8014 3398 8022
rect 2973 8006 2974 8014
rect 2989 8006 3002 8014
rect 2973 7998 2989 8006
rect 2970 7991 2989 7994
rect 2970 7982 2992 7991
rect 2943 7972 2992 7982
rect 2943 7966 2973 7972
rect 2992 7967 2997 7972
rect 2915 7950 2989 7966
rect 3007 7958 3037 8014
rect 3072 8004 3280 8014
rect 3315 8010 3360 8014
rect 3363 8013 3364 8014
rect 3379 8013 3392 8014
rect 3098 7974 3287 8004
rect 3113 7971 3287 7974
rect 3106 7968 3287 7971
rect 2915 7948 2928 7950
rect 2943 7948 2977 7950
rect 2915 7932 2989 7948
rect 3016 7944 3029 7958
rect 3044 7944 3060 7960
rect 3106 7955 3117 7968
rect 2899 7910 2900 7926
rect 2915 7910 2928 7932
rect 2943 7910 2973 7932
rect 3016 7928 3078 7944
rect 3106 7937 3117 7953
rect 3122 7948 3132 7968
rect 3142 7948 3156 7968
rect 3159 7955 3168 7968
rect 3184 7955 3193 7968
rect 3122 7937 3156 7948
rect 3159 7937 3168 7953
rect 3184 7937 3193 7953
rect 3200 7948 3210 7968
rect 3220 7948 3234 7968
rect 3235 7955 3246 7968
rect 3200 7937 3234 7948
rect 3235 7937 3246 7953
rect 3292 7944 3308 7960
rect 3315 7958 3345 8010
rect 3379 8006 3380 8013
rect 3364 7998 3380 8006
rect 3351 7966 3364 7985
rect 3379 7966 3409 7982
rect 3351 7950 3425 7966
rect 3351 7948 3364 7950
rect 3379 7948 3413 7950
rect 3016 7926 3029 7928
rect 3044 7926 3078 7928
rect 3016 7910 3078 7926
rect 3122 7921 3138 7924
rect 3200 7921 3230 7932
rect 3278 7928 3324 7944
rect 3351 7932 3425 7948
rect 3278 7926 3312 7928
rect 3277 7910 3324 7926
rect 3351 7910 3364 7932
rect 3379 7910 3409 7932
rect 3436 7910 3437 7926
rect 3452 7910 3465 8070
rect 3495 7966 3508 8070
rect 3553 8048 3554 8058
rect 3569 8048 3582 8058
rect 3553 8044 3582 8048
rect 3587 8044 3617 8070
rect 3635 8056 3651 8058
rect 3723 8056 3776 8070
rect 3724 8054 3788 8056
rect 3831 8054 3846 8070
rect 3895 8067 3925 8070
rect 3895 8064 3931 8067
rect 3861 8056 3877 8058
rect 3635 8044 3650 8048
rect 3553 8042 3650 8044
rect 3678 8042 3846 8054
rect 3862 8044 3877 8048
rect 3895 8045 3934 8064
rect 3953 8058 3960 8059
rect 3959 8051 3960 8058
rect 3943 8048 3944 8051
rect 3959 8048 3972 8051
rect 3895 8044 3925 8045
rect 3934 8044 3940 8045
rect 3943 8044 3972 8048
rect 3862 8043 3972 8044
rect 3862 8042 3978 8043
rect 3537 8034 3588 8042
rect 3537 8022 3562 8034
rect 3569 8022 3588 8034
rect 3619 8034 3669 8042
rect 3619 8026 3635 8034
rect 3642 8032 3669 8034
rect 3678 8032 3899 8042
rect 3642 8022 3899 8032
rect 3928 8034 3978 8042
rect 3928 8025 3944 8034
rect 3537 8014 3588 8022
rect 3635 8014 3899 8022
rect 3925 8022 3944 8025
rect 3951 8022 3978 8034
rect 3925 8014 3978 8022
rect 3553 8006 3554 8014
rect 3569 8006 3582 8014
rect 3553 7998 3569 8006
rect 3550 7991 3569 7994
rect 3550 7982 3572 7991
rect 3523 7972 3572 7982
rect 3523 7966 3553 7972
rect 3572 7967 3577 7972
rect 3495 7950 3569 7966
rect 3587 7958 3617 8014
rect 3652 8004 3860 8014
rect 3895 8010 3940 8014
rect 3943 8013 3944 8014
rect 3959 8013 3972 8014
rect 3678 7974 3867 8004
rect 3693 7971 3867 7974
rect 3686 7968 3867 7971
rect 3495 7948 3508 7950
rect 3523 7948 3557 7950
rect 3495 7932 3569 7948
rect 3596 7944 3609 7958
rect 3624 7944 3640 7960
rect 3686 7955 3697 7968
rect 3479 7910 3480 7926
rect 3495 7910 3508 7932
rect 3523 7910 3553 7932
rect 3596 7928 3658 7944
rect 3686 7937 3697 7953
rect 3702 7948 3712 7968
rect 3722 7948 3736 7968
rect 3739 7955 3748 7968
rect 3764 7955 3773 7968
rect 3702 7937 3736 7948
rect 3739 7937 3748 7953
rect 3764 7937 3773 7953
rect 3780 7948 3790 7968
rect 3800 7948 3814 7968
rect 3815 7955 3826 7968
rect 3780 7937 3814 7948
rect 3815 7937 3826 7953
rect 3872 7944 3888 7960
rect 3895 7958 3925 8010
rect 3959 8006 3960 8013
rect 3944 7998 3960 8006
rect 3931 7966 3944 7985
rect 3959 7966 3989 7982
rect 3931 7950 4005 7966
rect 3931 7948 3944 7950
rect 3959 7948 3993 7950
rect 3596 7926 3609 7928
rect 3624 7926 3658 7928
rect 3596 7910 3658 7926
rect 3702 7921 3718 7924
rect 3780 7921 3810 7932
rect 3858 7928 3904 7944
rect 3931 7932 4005 7948
rect 3858 7926 3892 7928
rect 3857 7910 3904 7926
rect 3931 7910 3944 7932
rect 3959 7910 3989 7932
rect 4016 7910 4017 7926
rect 4032 7910 4045 8070
rect 4075 7966 4088 8070
rect 4133 8048 4134 8058
rect 4149 8048 4162 8058
rect 4133 8044 4162 8048
rect 4167 8044 4197 8070
rect 4215 8056 4231 8058
rect 4303 8056 4356 8070
rect 4304 8054 4368 8056
rect 4411 8054 4426 8070
rect 4475 8067 4505 8070
rect 4475 8064 4511 8067
rect 4441 8056 4457 8058
rect 4215 8044 4230 8048
rect 4133 8042 4230 8044
rect 4258 8042 4426 8054
rect 4442 8044 4457 8048
rect 4475 8045 4514 8064
rect 4533 8058 4540 8059
rect 4539 8051 4540 8058
rect 4523 8048 4524 8051
rect 4539 8048 4552 8051
rect 4475 8044 4505 8045
rect 4514 8044 4520 8045
rect 4523 8044 4552 8048
rect 4442 8043 4552 8044
rect 4442 8042 4558 8043
rect 4117 8034 4168 8042
rect 4117 8022 4142 8034
rect 4149 8022 4168 8034
rect 4199 8034 4249 8042
rect 4199 8026 4215 8034
rect 4222 8032 4249 8034
rect 4258 8032 4479 8042
rect 4222 8022 4479 8032
rect 4508 8034 4558 8042
rect 4508 8025 4524 8034
rect 4117 8014 4168 8022
rect 4215 8014 4479 8022
rect 4505 8022 4524 8025
rect 4531 8022 4558 8034
rect 4505 8014 4558 8022
rect 4133 8006 4134 8014
rect 4149 8006 4162 8014
rect 4133 7998 4149 8006
rect 4130 7991 4149 7994
rect 4130 7982 4152 7991
rect 4103 7972 4152 7982
rect 4103 7966 4133 7972
rect 4152 7967 4157 7972
rect 4075 7950 4149 7966
rect 4167 7958 4197 8014
rect 4232 8004 4440 8014
rect 4475 8010 4520 8014
rect 4523 8013 4524 8014
rect 4539 8013 4552 8014
rect 4258 7974 4447 8004
rect 4273 7971 4447 7974
rect 4266 7968 4447 7971
rect 4075 7948 4088 7950
rect 4103 7948 4137 7950
rect 4075 7932 4149 7948
rect 4176 7944 4189 7958
rect 4204 7944 4220 7960
rect 4266 7955 4277 7968
rect 4059 7910 4060 7926
rect 4075 7910 4088 7932
rect 4103 7910 4133 7932
rect 4176 7928 4238 7944
rect 4266 7937 4277 7953
rect 4282 7948 4292 7968
rect 4302 7948 4316 7968
rect 4319 7955 4328 7968
rect 4344 7955 4353 7968
rect 4282 7937 4316 7948
rect 4319 7937 4328 7953
rect 4344 7937 4353 7953
rect 4360 7948 4370 7968
rect 4380 7948 4394 7968
rect 4395 7955 4406 7968
rect 4360 7937 4394 7948
rect 4395 7937 4406 7953
rect 4452 7944 4468 7960
rect 4475 7958 4505 8010
rect 4539 8006 4540 8013
rect 4524 7998 4540 8006
rect 4511 7966 4524 7985
rect 4539 7966 4569 7982
rect 4511 7950 4585 7966
rect 4511 7948 4524 7950
rect 4539 7948 4573 7950
rect 4176 7926 4189 7928
rect 4204 7926 4238 7928
rect 4176 7910 4238 7926
rect 4282 7921 4298 7924
rect 4360 7921 4390 7932
rect 4438 7928 4484 7944
rect 4511 7932 4585 7948
rect 4438 7926 4472 7928
rect 4437 7910 4484 7926
rect 4511 7910 4524 7932
rect 4539 7910 4569 7932
rect 4596 7910 4597 7926
rect 4612 7910 4625 8070
rect 4655 7966 4668 8070
rect 4713 8048 4714 8058
rect 4729 8048 4742 8058
rect 4713 8044 4742 8048
rect 4747 8044 4777 8070
rect 4795 8056 4811 8058
rect 4883 8056 4936 8070
rect 4884 8054 4948 8056
rect 4991 8054 5006 8070
rect 5055 8067 5085 8070
rect 5055 8064 5091 8067
rect 5021 8056 5037 8058
rect 4795 8044 4810 8048
rect 4713 8042 4810 8044
rect 4838 8042 5006 8054
rect 5022 8044 5037 8048
rect 5055 8045 5094 8064
rect 5113 8058 5120 8059
rect 5119 8051 5120 8058
rect 5103 8048 5104 8051
rect 5119 8048 5132 8051
rect 5055 8044 5085 8045
rect 5094 8044 5100 8045
rect 5103 8044 5132 8048
rect 5022 8043 5132 8044
rect 5022 8042 5138 8043
rect 4697 8034 4748 8042
rect 4697 8022 4722 8034
rect 4729 8022 4748 8034
rect 4779 8034 4829 8042
rect 4779 8026 4795 8034
rect 4802 8032 4829 8034
rect 4838 8032 5059 8042
rect 4802 8022 5059 8032
rect 5088 8034 5138 8042
rect 5088 8025 5104 8034
rect 4697 8014 4748 8022
rect 4795 8014 5059 8022
rect 5085 8022 5104 8025
rect 5111 8022 5138 8034
rect 5085 8014 5138 8022
rect 4713 8006 4714 8014
rect 4729 8006 4742 8014
rect 4713 7998 4729 8006
rect 4710 7991 4729 7994
rect 4710 7982 4732 7991
rect 4683 7972 4732 7982
rect 4683 7966 4713 7972
rect 4732 7967 4737 7972
rect 4655 7950 4729 7966
rect 4747 7958 4777 8014
rect 4812 8004 5020 8014
rect 5055 8010 5100 8014
rect 5103 8013 5104 8014
rect 5119 8013 5132 8014
rect 4838 7974 5027 8004
rect 4853 7971 5027 7974
rect 4846 7968 5027 7971
rect 4655 7948 4668 7950
rect 4683 7948 4717 7950
rect 4655 7932 4729 7948
rect 4756 7944 4769 7958
rect 4784 7944 4800 7960
rect 4846 7955 4857 7968
rect 4639 7910 4640 7926
rect 4655 7910 4668 7932
rect 4683 7910 4713 7932
rect 4756 7928 4818 7944
rect 4846 7937 4857 7953
rect 4862 7948 4872 7968
rect 4882 7948 4896 7968
rect 4899 7955 4908 7968
rect 4924 7955 4933 7968
rect 4862 7937 4896 7948
rect 4899 7937 4908 7953
rect 4924 7937 4933 7953
rect 4940 7948 4950 7968
rect 4960 7948 4974 7968
rect 4975 7955 4986 7968
rect 4940 7937 4974 7948
rect 4975 7937 4986 7953
rect 5032 7944 5048 7960
rect 5055 7958 5085 8010
rect 5119 8006 5120 8013
rect 5104 7998 5120 8006
rect 5091 7966 5104 7985
rect 5119 7966 5149 7982
rect 5091 7950 5165 7966
rect 5091 7948 5104 7950
rect 5119 7948 5153 7950
rect 4756 7926 4769 7928
rect 4784 7926 4818 7928
rect 4756 7910 4818 7926
rect 4862 7921 4878 7924
rect 4940 7921 4970 7932
rect 5018 7928 5064 7944
rect 5091 7932 5165 7948
rect 5018 7926 5052 7928
rect 5017 7910 5064 7926
rect 5091 7910 5104 7932
rect 5119 7910 5149 7932
rect 5176 7910 5177 7926
rect 5192 7910 5205 8070
rect 5235 7966 5248 8070
rect 5293 8048 5294 8058
rect 5309 8048 5322 8058
rect 5293 8044 5322 8048
rect 5327 8044 5357 8070
rect 5375 8056 5391 8058
rect 5463 8056 5516 8070
rect 5464 8054 5528 8056
rect 5571 8054 5586 8070
rect 5635 8067 5665 8070
rect 5635 8064 5671 8067
rect 5601 8056 5617 8058
rect 5375 8044 5390 8048
rect 5293 8042 5390 8044
rect 5418 8042 5586 8054
rect 5602 8044 5617 8048
rect 5635 8045 5674 8064
rect 5693 8058 5700 8059
rect 5699 8051 5700 8058
rect 5683 8048 5684 8051
rect 5699 8048 5712 8051
rect 5635 8044 5665 8045
rect 5674 8044 5680 8045
rect 5683 8044 5712 8048
rect 5602 8043 5712 8044
rect 5602 8042 5718 8043
rect 5277 8034 5328 8042
rect 5277 8022 5302 8034
rect 5309 8022 5328 8034
rect 5359 8034 5409 8042
rect 5359 8026 5375 8034
rect 5382 8032 5409 8034
rect 5418 8032 5639 8042
rect 5382 8022 5639 8032
rect 5668 8034 5718 8042
rect 5668 8025 5684 8034
rect 5277 8014 5328 8022
rect 5375 8014 5639 8022
rect 5665 8022 5684 8025
rect 5691 8022 5718 8034
rect 5665 8014 5718 8022
rect 5293 8006 5294 8014
rect 5309 8006 5322 8014
rect 5293 7998 5309 8006
rect 5290 7991 5309 7994
rect 5290 7982 5312 7991
rect 5263 7972 5312 7982
rect 5263 7966 5293 7972
rect 5312 7967 5317 7972
rect 5235 7950 5309 7966
rect 5327 7958 5357 8014
rect 5392 8004 5600 8014
rect 5635 8010 5680 8014
rect 5683 8013 5684 8014
rect 5699 8013 5712 8014
rect 5418 7974 5607 8004
rect 5433 7971 5607 7974
rect 5426 7968 5607 7971
rect 5235 7948 5248 7950
rect 5263 7948 5297 7950
rect 5235 7932 5309 7948
rect 5336 7944 5349 7958
rect 5364 7944 5380 7960
rect 5426 7955 5437 7968
rect 5219 7910 5220 7926
rect 5235 7910 5248 7932
rect 5263 7910 5293 7932
rect 5336 7928 5398 7944
rect 5426 7937 5437 7953
rect 5442 7948 5452 7968
rect 5462 7948 5476 7968
rect 5479 7955 5488 7968
rect 5504 7955 5513 7968
rect 5442 7937 5476 7948
rect 5479 7937 5488 7953
rect 5504 7937 5513 7953
rect 5520 7948 5530 7968
rect 5540 7948 5554 7968
rect 5555 7955 5566 7968
rect 5520 7937 5554 7948
rect 5555 7937 5566 7953
rect 5612 7944 5628 7960
rect 5635 7958 5665 8010
rect 5699 8006 5700 8013
rect 5684 7998 5700 8006
rect 5671 7966 5684 7985
rect 5699 7966 5729 7982
rect 5671 7950 5745 7966
rect 5671 7948 5684 7950
rect 5699 7948 5733 7950
rect 5336 7926 5349 7928
rect 5364 7926 5398 7928
rect 5336 7910 5398 7926
rect 5442 7921 5458 7924
rect 5520 7921 5550 7932
rect 5598 7928 5644 7944
rect 5671 7932 5745 7948
rect 5598 7926 5632 7928
rect 5597 7910 5644 7926
rect 5671 7910 5684 7932
rect 5699 7910 5729 7932
rect 5756 7910 5757 7926
rect 5772 7910 5785 8070
rect 5815 7966 5828 8070
rect 5873 8048 5874 8058
rect 5889 8048 5902 8058
rect 5873 8044 5902 8048
rect 5907 8044 5937 8070
rect 5955 8056 5971 8058
rect 6043 8056 6096 8070
rect 6044 8054 6108 8056
rect 6151 8054 6166 8070
rect 6215 8067 6245 8070
rect 6215 8064 6251 8067
rect 6181 8056 6197 8058
rect 5955 8044 5970 8048
rect 5873 8042 5970 8044
rect 5998 8042 6166 8054
rect 6182 8044 6197 8048
rect 6215 8045 6254 8064
rect 6273 8058 6280 8059
rect 6279 8051 6280 8058
rect 6263 8048 6264 8051
rect 6279 8048 6292 8051
rect 6215 8044 6245 8045
rect 6254 8044 6260 8045
rect 6263 8044 6292 8048
rect 6182 8043 6292 8044
rect 6182 8042 6298 8043
rect 5857 8034 5908 8042
rect 5857 8022 5882 8034
rect 5889 8022 5908 8034
rect 5939 8034 5989 8042
rect 5939 8026 5955 8034
rect 5962 8032 5989 8034
rect 5998 8032 6219 8042
rect 5962 8022 6219 8032
rect 6248 8034 6298 8042
rect 6248 8025 6264 8034
rect 5857 8014 5908 8022
rect 5955 8014 6219 8022
rect 6245 8022 6264 8025
rect 6271 8022 6298 8034
rect 6245 8014 6298 8022
rect 5873 8006 5874 8014
rect 5889 8006 5902 8014
rect 5873 7998 5889 8006
rect 5870 7991 5889 7994
rect 5870 7982 5892 7991
rect 5843 7972 5892 7982
rect 5843 7966 5873 7972
rect 5892 7967 5897 7972
rect 5815 7950 5889 7966
rect 5907 7958 5937 8014
rect 5972 8004 6180 8014
rect 6215 8010 6260 8014
rect 6263 8013 6264 8014
rect 6279 8013 6292 8014
rect 5998 7974 6187 8004
rect 6013 7971 6187 7974
rect 6006 7968 6187 7971
rect 5815 7948 5828 7950
rect 5843 7948 5877 7950
rect 5815 7932 5889 7948
rect 5916 7944 5929 7958
rect 5944 7944 5960 7960
rect 6006 7955 6017 7968
rect 5799 7910 5800 7926
rect 5815 7910 5828 7932
rect 5843 7910 5873 7932
rect 5916 7928 5978 7944
rect 6006 7937 6017 7953
rect 6022 7948 6032 7968
rect 6042 7948 6056 7968
rect 6059 7955 6068 7968
rect 6084 7955 6093 7968
rect 6022 7937 6056 7948
rect 6059 7937 6068 7953
rect 6084 7937 6093 7953
rect 6100 7948 6110 7968
rect 6120 7948 6134 7968
rect 6135 7955 6146 7968
rect 6100 7937 6134 7948
rect 6135 7937 6146 7953
rect 6192 7944 6208 7960
rect 6215 7958 6245 8010
rect 6279 8006 6280 8013
rect 6264 7998 6280 8006
rect 6251 7966 6264 7985
rect 6279 7966 6309 7982
rect 6251 7950 6325 7966
rect 6251 7948 6264 7950
rect 6279 7948 6313 7950
rect 5916 7926 5929 7928
rect 5944 7926 5978 7928
rect 5916 7910 5978 7926
rect 6022 7921 6038 7924
rect 6100 7921 6130 7932
rect 6178 7928 6224 7944
rect 6251 7932 6325 7948
rect 6178 7926 6212 7928
rect 6177 7910 6224 7926
rect 6251 7910 6264 7932
rect 6279 7910 6309 7932
rect 6336 7910 6337 7926
rect 6352 7910 6365 8070
rect 6395 7966 6408 8070
rect 6453 8048 6454 8058
rect 6469 8048 6482 8058
rect 6453 8044 6482 8048
rect 6487 8044 6517 8070
rect 6535 8056 6551 8058
rect 6623 8056 6676 8070
rect 6624 8054 6688 8056
rect 6731 8054 6746 8070
rect 6795 8067 6825 8070
rect 6795 8064 6831 8067
rect 6761 8056 6777 8058
rect 6535 8044 6550 8048
rect 6453 8042 6550 8044
rect 6578 8042 6746 8054
rect 6762 8044 6777 8048
rect 6795 8045 6834 8064
rect 6853 8058 6860 8059
rect 6859 8051 6860 8058
rect 6843 8048 6844 8051
rect 6859 8048 6872 8051
rect 6795 8044 6825 8045
rect 6834 8044 6840 8045
rect 6843 8044 6872 8048
rect 6762 8043 6872 8044
rect 6762 8042 6878 8043
rect 6437 8034 6488 8042
rect 6437 8022 6462 8034
rect 6469 8022 6488 8034
rect 6519 8034 6569 8042
rect 6519 8026 6535 8034
rect 6542 8032 6569 8034
rect 6578 8032 6799 8042
rect 6542 8022 6799 8032
rect 6828 8034 6878 8042
rect 6828 8025 6844 8034
rect 6437 8014 6488 8022
rect 6535 8014 6799 8022
rect 6825 8022 6844 8025
rect 6851 8022 6878 8034
rect 6825 8014 6878 8022
rect 6453 8006 6454 8014
rect 6469 8006 6482 8014
rect 6453 7998 6469 8006
rect 6450 7991 6469 7994
rect 6450 7982 6472 7991
rect 6423 7972 6472 7982
rect 6423 7966 6453 7972
rect 6472 7967 6477 7972
rect 6395 7950 6469 7966
rect 6487 7958 6517 8014
rect 6552 8004 6760 8014
rect 6795 8010 6840 8014
rect 6843 8013 6844 8014
rect 6859 8013 6872 8014
rect 6578 7974 6767 8004
rect 6593 7971 6767 7974
rect 6586 7968 6767 7971
rect 6395 7948 6408 7950
rect 6423 7948 6457 7950
rect 6395 7932 6469 7948
rect 6496 7944 6509 7958
rect 6524 7944 6540 7960
rect 6586 7955 6597 7968
rect 6379 7910 6380 7926
rect 6395 7910 6408 7932
rect 6423 7910 6453 7932
rect 6496 7928 6558 7944
rect 6586 7937 6597 7953
rect 6602 7948 6612 7968
rect 6622 7948 6636 7968
rect 6639 7955 6648 7968
rect 6664 7955 6673 7968
rect 6602 7937 6636 7948
rect 6639 7937 6648 7953
rect 6664 7937 6673 7953
rect 6680 7948 6690 7968
rect 6700 7948 6714 7968
rect 6715 7955 6726 7968
rect 6680 7937 6714 7948
rect 6715 7937 6726 7953
rect 6772 7944 6788 7960
rect 6795 7958 6825 8010
rect 6859 8006 6860 8013
rect 6844 7998 6860 8006
rect 6831 7966 6844 7985
rect 6859 7966 6889 7982
rect 6831 7950 6905 7966
rect 6831 7948 6844 7950
rect 6859 7948 6893 7950
rect 6496 7926 6509 7928
rect 6524 7926 6558 7928
rect 6496 7910 6558 7926
rect 6602 7921 6618 7924
rect 6680 7921 6710 7932
rect 6758 7928 6804 7944
rect 6831 7932 6905 7948
rect 6758 7926 6792 7928
rect 6757 7910 6804 7926
rect 6831 7910 6844 7932
rect 6859 7910 6889 7932
rect 6916 7910 6917 7926
rect 6932 7910 6945 8070
rect 6975 7966 6988 8070
rect 7033 8048 7034 8058
rect 7049 8048 7062 8058
rect 7033 8044 7062 8048
rect 7067 8044 7097 8070
rect 7115 8056 7131 8058
rect 7203 8056 7256 8070
rect 7204 8054 7268 8056
rect 7311 8054 7326 8070
rect 7375 8067 7405 8070
rect 7375 8064 7411 8067
rect 7341 8056 7357 8058
rect 7115 8044 7130 8048
rect 7033 8042 7130 8044
rect 7158 8042 7326 8054
rect 7342 8044 7357 8048
rect 7375 8045 7414 8064
rect 7433 8058 7440 8059
rect 7439 8051 7440 8058
rect 7423 8048 7424 8051
rect 7439 8048 7452 8051
rect 7375 8044 7405 8045
rect 7414 8044 7420 8045
rect 7423 8044 7452 8048
rect 7342 8043 7452 8044
rect 7342 8042 7458 8043
rect 7017 8034 7068 8042
rect 7017 8022 7042 8034
rect 7049 8022 7068 8034
rect 7099 8034 7149 8042
rect 7099 8026 7115 8034
rect 7122 8032 7149 8034
rect 7158 8032 7379 8042
rect 7122 8022 7379 8032
rect 7408 8034 7458 8042
rect 7408 8025 7424 8034
rect 7017 8014 7068 8022
rect 7115 8014 7379 8022
rect 7405 8022 7424 8025
rect 7431 8022 7458 8034
rect 7405 8014 7458 8022
rect 7033 8006 7034 8014
rect 7049 8006 7062 8014
rect 7033 7998 7049 8006
rect 7030 7991 7049 7994
rect 7030 7982 7052 7991
rect 7003 7972 7052 7982
rect 7003 7966 7033 7972
rect 7052 7967 7057 7972
rect 6975 7950 7049 7966
rect 7067 7958 7097 8014
rect 7132 8004 7340 8014
rect 7375 8010 7420 8014
rect 7423 8013 7424 8014
rect 7439 8013 7452 8014
rect 7158 7974 7347 8004
rect 7173 7971 7347 7974
rect 7166 7968 7347 7971
rect 6975 7948 6988 7950
rect 7003 7948 7037 7950
rect 6975 7932 7049 7948
rect 7076 7944 7089 7958
rect 7104 7944 7120 7960
rect 7166 7955 7177 7968
rect 6959 7910 6960 7926
rect 6975 7910 6988 7932
rect 7003 7910 7033 7932
rect 7076 7928 7138 7944
rect 7166 7937 7177 7953
rect 7182 7948 7192 7968
rect 7202 7948 7216 7968
rect 7219 7955 7228 7968
rect 7244 7955 7253 7968
rect 7182 7937 7216 7948
rect 7219 7937 7228 7953
rect 7244 7937 7253 7953
rect 7260 7948 7270 7968
rect 7280 7948 7294 7968
rect 7295 7955 7306 7968
rect 7260 7937 7294 7948
rect 7295 7937 7306 7953
rect 7352 7944 7368 7960
rect 7375 7958 7405 8010
rect 7439 8006 7440 8013
rect 7424 7998 7440 8006
rect 7411 7966 7424 7985
rect 7439 7966 7469 7982
rect 7411 7950 7485 7966
rect 7411 7948 7424 7950
rect 7439 7948 7473 7950
rect 7076 7926 7089 7928
rect 7104 7926 7138 7928
rect 7076 7910 7138 7926
rect 7182 7921 7198 7924
rect 7260 7921 7290 7932
rect 7338 7928 7384 7944
rect 7411 7932 7485 7948
rect 7338 7926 7372 7928
rect 7337 7910 7384 7926
rect 7411 7910 7424 7932
rect 7439 7910 7469 7932
rect 7496 7910 7497 7926
rect 7512 7910 7525 8070
rect 7555 7966 7568 8070
rect 7613 8048 7614 8058
rect 7629 8048 7642 8058
rect 7613 8044 7642 8048
rect 7647 8044 7677 8070
rect 7695 8056 7711 8058
rect 7783 8056 7836 8070
rect 7784 8054 7848 8056
rect 7891 8054 7906 8070
rect 7955 8067 7985 8070
rect 7955 8064 7991 8067
rect 7921 8056 7937 8058
rect 7695 8044 7710 8048
rect 7613 8042 7710 8044
rect 7738 8042 7906 8054
rect 7922 8044 7937 8048
rect 7955 8045 7994 8064
rect 8013 8058 8020 8059
rect 8019 8051 8020 8058
rect 8003 8048 8004 8051
rect 8019 8048 8032 8051
rect 7955 8044 7985 8045
rect 7994 8044 8000 8045
rect 8003 8044 8032 8048
rect 7922 8043 8032 8044
rect 7922 8042 8038 8043
rect 7597 8034 7648 8042
rect 7597 8022 7622 8034
rect 7629 8022 7648 8034
rect 7679 8034 7729 8042
rect 7679 8026 7695 8034
rect 7702 8032 7729 8034
rect 7738 8032 7959 8042
rect 7702 8022 7959 8032
rect 7988 8034 8038 8042
rect 7988 8025 8004 8034
rect 7597 8014 7648 8022
rect 7695 8014 7959 8022
rect 7985 8022 8004 8025
rect 8011 8022 8038 8034
rect 7985 8014 8038 8022
rect 7613 8006 7614 8014
rect 7629 8006 7642 8014
rect 7613 7998 7629 8006
rect 7610 7991 7629 7994
rect 7610 7982 7632 7991
rect 7583 7972 7632 7982
rect 7583 7966 7613 7972
rect 7632 7967 7637 7972
rect 7555 7950 7629 7966
rect 7647 7958 7677 8014
rect 7712 8004 7920 8014
rect 7955 8010 8000 8014
rect 8003 8013 8004 8014
rect 8019 8013 8032 8014
rect 7738 7974 7927 8004
rect 7753 7971 7927 7974
rect 7746 7968 7927 7971
rect 7555 7948 7568 7950
rect 7583 7948 7617 7950
rect 7555 7932 7629 7948
rect 7656 7944 7669 7958
rect 7684 7944 7700 7960
rect 7746 7955 7757 7968
rect 7539 7910 7540 7926
rect 7555 7910 7568 7932
rect 7583 7910 7613 7932
rect 7656 7928 7718 7944
rect 7746 7937 7757 7953
rect 7762 7948 7772 7968
rect 7782 7948 7796 7968
rect 7799 7955 7808 7968
rect 7824 7955 7833 7968
rect 7762 7937 7796 7948
rect 7799 7937 7808 7953
rect 7824 7937 7833 7953
rect 7840 7948 7850 7968
rect 7860 7948 7874 7968
rect 7875 7955 7886 7968
rect 7840 7937 7874 7948
rect 7875 7937 7886 7953
rect 7932 7944 7948 7960
rect 7955 7958 7985 8010
rect 8019 8006 8020 8013
rect 8004 7998 8020 8006
rect 7991 7966 8004 7985
rect 8019 7966 8049 7982
rect 7991 7950 8065 7966
rect 7991 7948 8004 7950
rect 8019 7948 8053 7950
rect 7656 7926 7669 7928
rect 7684 7926 7718 7928
rect 7656 7910 7718 7926
rect 7762 7921 7778 7924
rect 7840 7921 7870 7932
rect 7918 7928 7964 7944
rect 7991 7932 8065 7948
rect 7918 7926 7952 7928
rect 7917 7910 7964 7926
rect 7991 7910 8004 7932
rect 8019 7910 8049 7932
rect 8076 7910 8077 7926
rect 8092 7910 8105 8070
rect 8135 7966 8148 8070
rect 8193 8048 8194 8058
rect 8209 8048 8222 8058
rect 8193 8044 8222 8048
rect 8227 8044 8257 8070
rect 8275 8056 8291 8058
rect 8363 8056 8416 8070
rect 8364 8054 8428 8056
rect 8471 8054 8486 8070
rect 8535 8067 8565 8070
rect 8535 8064 8571 8067
rect 8501 8056 8517 8058
rect 8275 8044 8290 8048
rect 8193 8042 8290 8044
rect 8318 8042 8486 8054
rect 8502 8044 8517 8048
rect 8535 8045 8574 8064
rect 8593 8058 8600 8059
rect 8599 8051 8600 8058
rect 8583 8048 8584 8051
rect 8599 8048 8612 8051
rect 8535 8044 8565 8045
rect 8574 8044 8580 8045
rect 8583 8044 8612 8048
rect 8502 8043 8612 8044
rect 8502 8042 8618 8043
rect 8177 8034 8228 8042
rect 8177 8022 8202 8034
rect 8209 8022 8228 8034
rect 8259 8034 8309 8042
rect 8259 8026 8275 8034
rect 8282 8032 8309 8034
rect 8318 8032 8539 8042
rect 8282 8022 8539 8032
rect 8568 8034 8618 8042
rect 8568 8025 8584 8034
rect 8177 8014 8228 8022
rect 8275 8014 8539 8022
rect 8565 8022 8584 8025
rect 8591 8022 8618 8034
rect 8565 8014 8618 8022
rect 8193 8006 8194 8014
rect 8209 8006 8222 8014
rect 8193 7998 8209 8006
rect 8190 7991 8209 7994
rect 8190 7982 8212 7991
rect 8163 7972 8212 7982
rect 8163 7966 8193 7972
rect 8212 7967 8217 7972
rect 8135 7950 8209 7966
rect 8227 7958 8257 8014
rect 8292 8004 8500 8014
rect 8535 8010 8580 8014
rect 8583 8013 8584 8014
rect 8599 8013 8612 8014
rect 8318 7974 8507 8004
rect 8333 7971 8507 7974
rect 8326 7968 8507 7971
rect 8135 7948 8148 7950
rect 8163 7948 8197 7950
rect 8135 7932 8209 7948
rect 8236 7944 8249 7958
rect 8264 7944 8280 7960
rect 8326 7955 8337 7968
rect 8119 7910 8120 7926
rect 8135 7910 8148 7932
rect 8163 7910 8193 7932
rect 8236 7928 8298 7944
rect 8326 7937 8337 7953
rect 8342 7948 8352 7968
rect 8362 7948 8376 7968
rect 8379 7955 8388 7968
rect 8404 7955 8413 7968
rect 8342 7937 8376 7948
rect 8379 7937 8388 7953
rect 8404 7937 8413 7953
rect 8420 7948 8430 7968
rect 8440 7948 8454 7968
rect 8455 7955 8466 7968
rect 8420 7937 8454 7948
rect 8455 7937 8466 7953
rect 8512 7944 8528 7960
rect 8535 7958 8565 8010
rect 8599 8006 8600 8013
rect 8584 7998 8600 8006
rect 8571 7966 8584 7985
rect 8599 7966 8629 7982
rect 8571 7950 8645 7966
rect 8571 7948 8584 7950
rect 8599 7948 8633 7950
rect 8236 7926 8249 7928
rect 8264 7926 8298 7928
rect 8236 7910 8298 7926
rect 8342 7921 8358 7924
rect 8420 7921 8450 7932
rect 8498 7928 8544 7944
rect 8571 7932 8645 7948
rect 8498 7926 8532 7928
rect 8497 7910 8544 7926
rect 8571 7910 8584 7932
rect 8599 7910 8629 7932
rect 8656 7910 8657 7926
rect 8672 7910 8685 8070
rect 8715 7966 8728 8070
rect 8773 8048 8774 8058
rect 8789 8048 8802 8058
rect 8773 8044 8802 8048
rect 8807 8044 8837 8070
rect 8855 8056 8871 8058
rect 8943 8056 8996 8070
rect 8944 8054 9008 8056
rect 9051 8054 9066 8070
rect 9115 8067 9145 8070
rect 9115 8064 9151 8067
rect 9081 8056 9097 8058
rect 8855 8044 8870 8048
rect 8773 8042 8870 8044
rect 8898 8042 9066 8054
rect 9082 8044 9097 8048
rect 9115 8045 9154 8064
rect 9173 8058 9180 8059
rect 9179 8051 9180 8058
rect 9163 8048 9164 8051
rect 9179 8048 9192 8051
rect 9115 8044 9145 8045
rect 9154 8044 9160 8045
rect 9163 8044 9192 8048
rect 9082 8043 9192 8044
rect 9082 8042 9198 8043
rect 8757 8034 8808 8042
rect 8757 8022 8782 8034
rect 8789 8022 8808 8034
rect 8839 8034 8889 8042
rect 8839 8026 8855 8034
rect 8862 8032 8889 8034
rect 8898 8032 9119 8042
rect 8862 8022 9119 8032
rect 9148 8034 9198 8042
rect 9148 8025 9164 8034
rect 8757 8014 8808 8022
rect 8855 8014 9119 8022
rect 9145 8022 9164 8025
rect 9171 8022 9198 8034
rect 9145 8014 9198 8022
rect 8773 8006 8774 8014
rect 8789 8006 8802 8014
rect 8773 7998 8789 8006
rect 8770 7991 8789 7994
rect 8770 7982 8792 7991
rect 8743 7972 8792 7982
rect 8743 7966 8773 7972
rect 8792 7967 8797 7972
rect 8715 7950 8789 7966
rect 8807 7958 8837 8014
rect 8872 8004 9080 8014
rect 9115 8010 9160 8014
rect 9163 8013 9164 8014
rect 9179 8013 9192 8014
rect 8898 7974 9087 8004
rect 8913 7971 9087 7974
rect 8906 7968 9087 7971
rect 8715 7948 8728 7950
rect 8743 7948 8777 7950
rect 8715 7932 8789 7948
rect 8816 7944 8829 7958
rect 8844 7944 8860 7960
rect 8906 7955 8917 7968
rect 8699 7910 8700 7926
rect 8715 7910 8728 7932
rect 8743 7910 8773 7932
rect 8816 7928 8878 7944
rect 8906 7937 8917 7953
rect 8922 7948 8932 7968
rect 8942 7948 8956 7968
rect 8959 7955 8968 7968
rect 8984 7955 8993 7968
rect 8922 7937 8956 7948
rect 8959 7937 8968 7953
rect 8984 7937 8993 7953
rect 9000 7948 9010 7968
rect 9020 7948 9034 7968
rect 9035 7955 9046 7968
rect 9000 7937 9034 7948
rect 9035 7937 9046 7953
rect 9092 7944 9108 7960
rect 9115 7958 9145 8010
rect 9179 8006 9180 8013
rect 9164 7998 9180 8006
rect 9151 7966 9164 7985
rect 9179 7966 9209 7982
rect 9151 7950 9225 7966
rect 9151 7948 9164 7950
rect 9179 7948 9213 7950
rect 8816 7926 8829 7928
rect 8844 7926 8878 7928
rect 8816 7910 8878 7926
rect 8922 7921 8938 7924
rect 9000 7921 9030 7932
rect 9078 7928 9124 7944
rect 9151 7932 9225 7948
rect 9078 7926 9112 7928
rect 9077 7910 9124 7926
rect 9151 7910 9164 7932
rect 9179 7910 9209 7932
rect 9236 7910 9237 7926
rect 9252 7910 9265 8070
rect -7 7902 34 7910
rect -7 7876 8 7902
rect 15 7876 34 7902
rect 98 7898 160 7910
rect 172 7898 247 7910
rect 305 7898 380 7910
rect 392 7898 423 7910
rect 429 7898 464 7910
rect 98 7896 260 7898
rect -7 7868 34 7876
rect 116 7872 129 7896
rect 144 7894 159 7896
rect -1 7858 0 7868
rect 15 7858 28 7868
rect 43 7858 73 7872
rect 116 7858 159 7872
rect 183 7869 190 7876
rect 193 7872 260 7896
rect 292 7896 464 7898
rect 262 7874 290 7878
rect 292 7874 372 7896
rect 393 7894 408 7896
rect 262 7872 372 7874
rect 193 7868 372 7872
rect 166 7858 196 7868
rect 198 7858 351 7868
rect 359 7858 389 7868
rect 393 7858 423 7872
rect 451 7858 464 7896
rect 536 7902 571 7910
rect 536 7876 537 7902
rect 544 7876 571 7902
rect 479 7858 509 7872
rect 536 7868 571 7876
rect 573 7902 614 7910
rect 573 7876 588 7902
rect 595 7876 614 7902
rect 678 7898 740 7910
rect 752 7898 827 7910
rect 885 7898 960 7910
rect 972 7898 1003 7910
rect 1009 7898 1044 7910
rect 678 7896 840 7898
rect 573 7868 614 7876
rect 696 7872 709 7896
rect 724 7894 739 7896
rect 536 7858 537 7868
rect 552 7858 565 7868
rect 579 7858 580 7868
rect 595 7858 608 7868
rect 623 7858 653 7872
rect 696 7858 739 7872
rect 763 7869 770 7876
rect 773 7872 840 7896
rect 872 7896 1044 7898
rect 842 7874 870 7878
rect 872 7874 952 7896
rect 973 7894 988 7896
rect 842 7872 952 7874
rect 773 7868 952 7872
rect 746 7858 776 7868
rect 778 7858 931 7868
rect 939 7858 969 7868
rect 973 7858 1003 7872
rect 1031 7858 1044 7896
rect 1116 7902 1151 7910
rect 1116 7876 1117 7902
rect 1124 7876 1151 7902
rect 1059 7858 1089 7872
rect 1116 7868 1151 7876
rect 1153 7902 1194 7910
rect 1153 7876 1168 7902
rect 1175 7876 1194 7902
rect 1258 7898 1320 7910
rect 1332 7898 1407 7910
rect 1465 7898 1540 7910
rect 1552 7898 1583 7910
rect 1589 7898 1624 7910
rect 1258 7896 1420 7898
rect 1153 7868 1194 7876
rect 1276 7872 1289 7896
rect 1304 7894 1319 7896
rect 1116 7858 1117 7868
rect 1132 7858 1145 7868
rect 1159 7858 1160 7868
rect 1175 7858 1188 7868
rect 1203 7858 1233 7872
rect 1276 7858 1319 7872
rect 1343 7869 1350 7876
rect 1353 7872 1420 7896
rect 1452 7896 1624 7898
rect 1422 7874 1450 7878
rect 1452 7874 1532 7896
rect 1553 7894 1568 7896
rect 1422 7872 1532 7874
rect 1353 7868 1532 7872
rect 1326 7858 1356 7868
rect 1358 7858 1511 7868
rect 1519 7858 1549 7868
rect 1553 7858 1583 7872
rect 1611 7858 1624 7896
rect 1696 7902 1731 7910
rect 1696 7876 1697 7902
rect 1704 7876 1731 7902
rect 1639 7858 1669 7872
rect 1696 7868 1731 7876
rect 1733 7902 1774 7910
rect 1733 7876 1748 7902
rect 1755 7876 1774 7902
rect 1838 7898 1900 7910
rect 1912 7898 1987 7910
rect 2045 7898 2120 7910
rect 2132 7898 2163 7910
rect 2169 7898 2204 7910
rect 1838 7896 2000 7898
rect 1733 7868 1774 7876
rect 1856 7872 1869 7896
rect 1884 7894 1899 7896
rect 1696 7858 1697 7868
rect 1712 7858 1725 7868
rect 1739 7858 1740 7868
rect 1755 7858 1768 7868
rect 1783 7858 1813 7872
rect 1856 7858 1899 7872
rect 1923 7869 1930 7876
rect 1933 7872 2000 7896
rect 2032 7896 2204 7898
rect 2002 7874 2030 7878
rect 2032 7874 2112 7896
rect 2133 7894 2148 7896
rect 2002 7872 2112 7874
rect 1933 7868 2112 7872
rect 1906 7858 1936 7868
rect 1938 7858 2091 7868
rect 2099 7858 2129 7868
rect 2133 7858 2163 7872
rect 2191 7858 2204 7896
rect 2276 7902 2311 7910
rect 2276 7876 2277 7902
rect 2284 7876 2311 7902
rect 2219 7858 2249 7872
rect 2276 7868 2311 7876
rect 2313 7902 2354 7910
rect 2313 7876 2328 7902
rect 2335 7876 2354 7902
rect 2418 7898 2480 7910
rect 2492 7898 2567 7910
rect 2625 7898 2700 7910
rect 2712 7898 2743 7910
rect 2749 7898 2784 7910
rect 2418 7896 2580 7898
rect 2313 7868 2354 7876
rect 2436 7872 2449 7896
rect 2464 7894 2479 7896
rect 2276 7858 2277 7868
rect 2292 7858 2305 7868
rect 2319 7858 2320 7868
rect 2335 7858 2348 7868
rect 2363 7858 2393 7872
rect 2436 7858 2479 7872
rect 2503 7869 2510 7876
rect 2513 7872 2580 7896
rect 2612 7896 2784 7898
rect 2582 7874 2610 7878
rect 2612 7874 2692 7896
rect 2713 7894 2728 7896
rect 2582 7872 2692 7874
rect 2513 7868 2692 7872
rect 2486 7858 2516 7868
rect 2518 7858 2671 7868
rect 2679 7858 2709 7868
rect 2713 7858 2743 7872
rect 2771 7858 2784 7896
rect 2856 7902 2891 7910
rect 2856 7876 2857 7902
rect 2864 7876 2891 7902
rect 2799 7858 2829 7872
rect 2856 7868 2891 7876
rect 2893 7902 2934 7910
rect 2893 7876 2908 7902
rect 2915 7876 2934 7902
rect 2998 7898 3060 7910
rect 3072 7898 3147 7910
rect 3205 7898 3280 7910
rect 3292 7898 3323 7910
rect 3329 7898 3364 7910
rect 2998 7896 3160 7898
rect 2893 7868 2934 7876
rect 3016 7872 3029 7896
rect 3044 7894 3059 7896
rect 2856 7858 2857 7868
rect 2872 7858 2885 7868
rect 2899 7858 2900 7868
rect 2915 7858 2928 7868
rect 2943 7858 2973 7872
rect 3016 7858 3059 7872
rect 3083 7869 3090 7876
rect 3093 7872 3160 7896
rect 3192 7896 3364 7898
rect 3162 7874 3190 7878
rect 3192 7874 3272 7896
rect 3293 7894 3308 7896
rect 3162 7872 3272 7874
rect 3093 7868 3272 7872
rect 3066 7858 3096 7868
rect 3098 7858 3251 7868
rect 3259 7858 3289 7868
rect 3293 7858 3323 7872
rect 3351 7858 3364 7896
rect 3436 7902 3471 7910
rect 3436 7876 3437 7902
rect 3444 7876 3471 7902
rect 3379 7858 3409 7872
rect 3436 7868 3471 7876
rect 3473 7902 3514 7910
rect 3473 7876 3488 7902
rect 3495 7876 3514 7902
rect 3578 7898 3640 7910
rect 3652 7898 3727 7910
rect 3785 7898 3860 7910
rect 3872 7898 3903 7910
rect 3909 7898 3944 7910
rect 3578 7896 3740 7898
rect 3473 7868 3514 7876
rect 3596 7872 3609 7896
rect 3624 7894 3639 7896
rect 3436 7858 3437 7868
rect 3452 7858 3465 7868
rect 3479 7858 3480 7868
rect 3495 7858 3508 7868
rect 3523 7858 3553 7872
rect 3596 7858 3639 7872
rect 3663 7869 3670 7876
rect 3673 7872 3740 7896
rect 3772 7896 3944 7898
rect 3742 7874 3770 7878
rect 3772 7874 3852 7896
rect 3873 7894 3888 7896
rect 3742 7872 3852 7874
rect 3673 7868 3852 7872
rect 3646 7858 3676 7868
rect 3678 7858 3831 7868
rect 3839 7858 3869 7868
rect 3873 7858 3903 7872
rect 3931 7858 3944 7896
rect 4016 7902 4051 7910
rect 4016 7876 4017 7902
rect 4024 7876 4051 7902
rect 3959 7858 3989 7872
rect 4016 7868 4051 7876
rect 4053 7902 4094 7910
rect 4053 7876 4068 7902
rect 4075 7876 4094 7902
rect 4158 7898 4220 7910
rect 4232 7898 4307 7910
rect 4365 7898 4440 7910
rect 4452 7898 4483 7910
rect 4489 7898 4524 7910
rect 4158 7896 4320 7898
rect 4053 7868 4094 7876
rect 4176 7872 4189 7896
rect 4204 7894 4219 7896
rect 4016 7858 4017 7868
rect 4032 7858 4045 7868
rect 4059 7858 4060 7868
rect 4075 7858 4088 7868
rect 4103 7858 4133 7872
rect 4176 7858 4219 7872
rect 4243 7869 4250 7876
rect 4253 7872 4320 7896
rect 4352 7896 4524 7898
rect 4322 7874 4350 7878
rect 4352 7874 4432 7896
rect 4453 7894 4468 7896
rect 4322 7872 4432 7874
rect 4253 7868 4432 7872
rect 4226 7858 4256 7868
rect 4258 7858 4411 7868
rect 4419 7858 4449 7868
rect 4453 7858 4483 7872
rect 4511 7858 4524 7896
rect 4596 7902 4631 7910
rect 4596 7876 4597 7902
rect 4604 7876 4631 7902
rect 4539 7858 4569 7872
rect 4596 7868 4631 7876
rect 4633 7902 4674 7910
rect 4633 7876 4648 7902
rect 4655 7876 4674 7902
rect 4738 7898 4800 7910
rect 4812 7898 4887 7910
rect 4945 7898 5020 7910
rect 5032 7898 5063 7910
rect 5069 7898 5104 7910
rect 4738 7896 4900 7898
rect 4633 7868 4674 7876
rect 4756 7872 4769 7896
rect 4784 7894 4799 7896
rect 4596 7858 4597 7868
rect 4612 7858 4625 7868
rect 4639 7858 4640 7868
rect 4655 7858 4668 7868
rect 4683 7858 4713 7872
rect 4756 7858 4799 7872
rect 4823 7869 4830 7876
rect 4833 7872 4900 7896
rect 4932 7896 5104 7898
rect 4902 7874 4930 7878
rect 4932 7874 5012 7896
rect 5033 7894 5048 7896
rect 4902 7872 5012 7874
rect 4833 7868 5012 7872
rect 4806 7858 4836 7868
rect 4838 7858 4991 7868
rect 4999 7858 5029 7868
rect 5033 7858 5063 7872
rect 5091 7858 5104 7896
rect 5176 7902 5211 7910
rect 5176 7876 5177 7902
rect 5184 7876 5211 7902
rect 5119 7858 5149 7872
rect 5176 7868 5211 7876
rect 5213 7902 5254 7910
rect 5213 7876 5228 7902
rect 5235 7876 5254 7902
rect 5318 7898 5380 7910
rect 5392 7898 5467 7910
rect 5525 7898 5600 7910
rect 5612 7898 5643 7910
rect 5649 7898 5684 7910
rect 5318 7896 5480 7898
rect 5213 7868 5254 7876
rect 5336 7872 5349 7896
rect 5364 7894 5379 7896
rect 5176 7858 5177 7868
rect 5192 7858 5205 7868
rect 5219 7858 5220 7868
rect 5235 7858 5248 7868
rect 5263 7858 5293 7872
rect 5336 7858 5379 7872
rect 5403 7869 5410 7876
rect 5413 7872 5480 7896
rect 5512 7896 5684 7898
rect 5482 7874 5510 7878
rect 5512 7874 5592 7896
rect 5613 7894 5628 7896
rect 5482 7872 5592 7874
rect 5413 7868 5592 7872
rect 5386 7858 5416 7868
rect 5418 7858 5571 7868
rect 5579 7858 5609 7868
rect 5613 7858 5643 7872
rect 5671 7858 5684 7896
rect 5756 7902 5791 7910
rect 5756 7876 5757 7902
rect 5764 7876 5791 7902
rect 5699 7858 5729 7872
rect 5756 7868 5791 7876
rect 5793 7902 5834 7910
rect 5793 7876 5808 7902
rect 5815 7876 5834 7902
rect 5898 7898 5960 7910
rect 5972 7898 6047 7910
rect 6105 7898 6180 7910
rect 6192 7898 6223 7910
rect 6229 7898 6264 7910
rect 5898 7896 6060 7898
rect 5793 7868 5834 7876
rect 5916 7872 5929 7896
rect 5944 7894 5959 7896
rect 5756 7858 5757 7868
rect 5772 7858 5785 7868
rect 5799 7858 5800 7868
rect 5815 7858 5828 7868
rect 5843 7858 5873 7872
rect 5916 7858 5959 7872
rect 5983 7869 5990 7876
rect 5993 7872 6060 7896
rect 6092 7896 6264 7898
rect 6062 7874 6090 7878
rect 6092 7874 6172 7896
rect 6193 7894 6208 7896
rect 6062 7872 6172 7874
rect 5993 7868 6172 7872
rect 5966 7858 5996 7868
rect 5998 7858 6151 7868
rect 6159 7858 6189 7868
rect 6193 7858 6223 7872
rect 6251 7858 6264 7896
rect 6336 7902 6371 7910
rect 6336 7876 6337 7902
rect 6344 7876 6371 7902
rect 6279 7858 6309 7872
rect 6336 7868 6371 7876
rect 6373 7902 6414 7910
rect 6373 7876 6388 7902
rect 6395 7876 6414 7902
rect 6478 7898 6540 7910
rect 6552 7898 6627 7910
rect 6685 7898 6760 7910
rect 6772 7898 6803 7910
rect 6809 7898 6844 7910
rect 6478 7896 6640 7898
rect 6373 7868 6414 7876
rect 6496 7872 6509 7896
rect 6524 7894 6539 7896
rect 6336 7858 6337 7868
rect 6352 7858 6365 7868
rect 6379 7858 6380 7868
rect 6395 7858 6408 7868
rect 6423 7858 6453 7872
rect 6496 7858 6539 7872
rect 6563 7869 6570 7876
rect 6573 7872 6640 7896
rect 6672 7896 6844 7898
rect 6642 7874 6670 7878
rect 6672 7874 6752 7896
rect 6773 7894 6788 7896
rect 6642 7872 6752 7874
rect 6573 7868 6752 7872
rect 6546 7858 6576 7868
rect 6578 7858 6731 7868
rect 6739 7858 6769 7868
rect 6773 7858 6803 7872
rect 6831 7858 6844 7896
rect 6916 7902 6951 7910
rect 6916 7876 6917 7902
rect 6924 7876 6951 7902
rect 6859 7858 6889 7872
rect 6916 7868 6951 7876
rect 6953 7902 6994 7910
rect 6953 7876 6968 7902
rect 6975 7876 6994 7902
rect 7058 7898 7120 7910
rect 7132 7898 7207 7910
rect 7265 7898 7340 7910
rect 7352 7898 7383 7910
rect 7389 7898 7424 7910
rect 7058 7896 7220 7898
rect 6953 7868 6994 7876
rect 7076 7872 7089 7896
rect 7104 7894 7119 7896
rect 6916 7858 6917 7868
rect 6932 7858 6945 7868
rect 6959 7858 6960 7868
rect 6975 7858 6988 7868
rect 7003 7858 7033 7872
rect 7076 7858 7119 7872
rect 7143 7869 7150 7876
rect 7153 7872 7220 7896
rect 7252 7896 7424 7898
rect 7222 7874 7250 7878
rect 7252 7874 7332 7896
rect 7353 7894 7368 7896
rect 7222 7872 7332 7874
rect 7153 7868 7332 7872
rect 7126 7858 7156 7868
rect 7158 7858 7311 7868
rect 7319 7858 7349 7868
rect 7353 7858 7383 7872
rect 7411 7858 7424 7896
rect 7496 7902 7531 7910
rect 7496 7876 7497 7902
rect 7504 7876 7531 7902
rect 7439 7858 7469 7872
rect 7496 7868 7531 7876
rect 7533 7902 7574 7910
rect 7533 7876 7548 7902
rect 7555 7876 7574 7902
rect 7638 7898 7700 7910
rect 7712 7898 7787 7910
rect 7845 7898 7920 7910
rect 7932 7898 7963 7910
rect 7969 7898 8004 7910
rect 7638 7896 7800 7898
rect 7533 7868 7574 7876
rect 7656 7872 7669 7896
rect 7684 7894 7699 7896
rect 7496 7858 7497 7868
rect 7512 7858 7525 7868
rect 7539 7858 7540 7868
rect 7555 7858 7568 7868
rect 7583 7858 7613 7872
rect 7656 7858 7699 7872
rect 7723 7869 7730 7876
rect 7733 7872 7800 7896
rect 7832 7896 8004 7898
rect 7802 7874 7830 7878
rect 7832 7874 7912 7896
rect 7933 7894 7948 7896
rect 7802 7872 7912 7874
rect 7733 7868 7912 7872
rect 7706 7858 7736 7868
rect 7738 7858 7891 7868
rect 7899 7858 7929 7868
rect 7933 7858 7963 7872
rect 7991 7858 8004 7896
rect 8076 7902 8111 7910
rect 8076 7876 8077 7902
rect 8084 7876 8111 7902
rect 8019 7858 8049 7872
rect 8076 7868 8111 7876
rect 8113 7902 8154 7910
rect 8113 7876 8128 7902
rect 8135 7876 8154 7902
rect 8218 7898 8280 7910
rect 8292 7898 8367 7910
rect 8425 7898 8500 7910
rect 8512 7898 8543 7910
rect 8549 7898 8584 7910
rect 8218 7896 8380 7898
rect 8113 7868 8154 7876
rect 8236 7872 8249 7896
rect 8264 7894 8279 7896
rect 8076 7858 8077 7868
rect 8092 7858 8105 7868
rect 8119 7858 8120 7868
rect 8135 7858 8148 7868
rect 8163 7858 8193 7872
rect 8236 7858 8279 7872
rect 8303 7869 8310 7876
rect 8313 7872 8380 7896
rect 8412 7896 8584 7898
rect 8382 7874 8410 7878
rect 8412 7874 8492 7896
rect 8513 7894 8528 7896
rect 8382 7872 8492 7874
rect 8313 7868 8492 7872
rect 8286 7858 8316 7868
rect 8318 7858 8471 7868
rect 8479 7858 8509 7868
rect 8513 7858 8543 7872
rect 8571 7858 8584 7896
rect 8656 7902 8691 7910
rect 8656 7876 8657 7902
rect 8664 7876 8691 7902
rect 8599 7858 8629 7872
rect 8656 7868 8691 7876
rect 8693 7902 8734 7910
rect 8693 7876 8708 7902
rect 8715 7876 8734 7902
rect 8798 7898 8860 7910
rect 8872 7898 8947 7910
rect 9005 7898 9080 7910
rect 9092 7898 9123 7910
rect 9129 7898 9164 7910
rect 8798 7896 8960 7898
rect 8693 7868 8734 7876
rect 8816 7872 8829 7896
rect 8844 7894 8859 7896
rect 8656 7858 8657 7868
rect 8672 7858 8685 7868
rect 8699 7858 8700 7868
rect 8715 7858 8728 7868
rect 8743 7858 8773 7872
rect 8816 7858 8859 7872
rect 8883 7869 8890 7876
rect 8893 7872 8960 7896
rect 8992 7896 9164 7898
rect 8962 7874 8990 7878
rect 8992 7874 9072 7896
rect 9093 7894 9108 7896
rect 8962 7872 9072 7874
rect 8893 7868 9072 7872
rect 8866 7858 8896 7868
rect 8898 7858 9051 7868
rect 9059 7858 9089 7868
rect 9093 7858 9123 7872
rect 9151 7858 9164 7896
rect 9236 7902 9271 7910
rect 9236 7876 9237 7902
rect 9244 7876 9271 7902
rect 9179 7858 9209 7872
rect 9236 7868 9271 7876
rect 9236 7858 9237 7868
rect 9252 7858 9265 7868
rect -1 7852 9265 7858
rect 0 7844 9265 7852
rect 15 7814 28 7844
rect 43 7826 73 7844
rect 116 7830 130 7844
rect 166 7830 386 7844
rect 117 7828 130 7830
rect 83 7816 98 7828
rect 80 7814 102 7816
rect 107 7814 137 7828
rect 198 7826 351 7830
rect 180 7814 372 7826
rect 415 7814 445 7828
rect 451 7814 464 7844
rect 479 7826 509 7844
rect 552 7814 565 7844
rect 595 7814 608 7844
rect 623 7826 653 7844
rect 696 7830 710 7844
rect 746 7830 966 7844
rect 697 7828 710 7830
rect 663 7816 678 7828
rect 660 7814 682 7816
rect 687 7814 717 7828
rect 778 7826 931 7830
rect 760 7814 952 7826
rect 995 7814 1025 7828
rect 1031 7814 1044 7844
rect 1059 7826 1089 7844
rect 1132 7814 1145 7844
rect 1175 7814 1188 7844
rect 1203 7826 1233 7844
rect 1276 7830 1290 7844
rect 1326 7830 1546 7844
rect 1277 7828 1290 7830
rect 1243 7816 1258 7828
rect 1240 7814 1262 7816
rect 1267 7814 1297 7828
rect 1358 7826 1511 7830
rect 1340 7814 1532 7826
rect 1575 7814 1605 7828
rect 1611 7814 1624 7844
rect 1639 7826 1669 7844
rect 1712 7814 1725 7844
rect 1755 7814 1768 7844
rect 1783 7826 1813 7844
rect 1856 7830 1870 7844
rect 1906 7830 2126 7844
rect 1857 7828 1870 7830
rect 1823 7816 1838 7828
rect 1820 7814 1842 7816
rect 1847 7814 1877 7828
rect 1938 7826 2091 7830
rect 1920 7814 2112 7826
rect 2155 7814 2185 7828
rect 2191 7814 2204 7844
rect 2219 7826 2249 7844
rect 2292 7814 2305 7844
rect 2335 7814 2348 7844
rect 2363 7826 2393 7844
rect 2436 7830 2450 7844
rect 2486 7830 2706 7844
rect 2437 7828 2450 7830
rect 2403 7816 2418 7828
rect 2400 7814 2422 7816
rect 2427 7814 2457 7828
rect 2518 7826 2671 7830
rect 2500 7814 2692 7826
rect 2735 7814 2765 7828
rect 2771 7814 2784 7844
rect 2799 7826 2829 7844
rect 2872 7814 2885 7844
rect 2915 7814 2928 7844
rect 2943 7826 2973 7844
rect 3016 7830 3030 7844
rect 3066 7830 3286 7844
rect 3017 7828 3030 7830
rect 2983 7816 2998 7828
rect 2980 7814 3002 7816
rect 3007 7814 3037 7828
rect 3098 7826 3251 7830
rect 3080 7814 3272 7826
rect 3315 7814 3345 7828
rect 3351 7814 3364 7844
rect 3379 7826 3409 7844
rect 3452 7814 3465 7844
rect 3495 7814 3508 7844
rect 3523 7826 3553 7844
rect 3596 7830 3610 7844
rect 3646 7830 3866 7844
rect 3597 7828 3610 7830
rect 3563 7816 3578 7828
rect 3560 7814 3582 7816
rect 3587 7814 3617 7828
rect 3678 7826 3831 7830
rect 3660 7814 3852 7826
rect 3895 7814 3925 7828
rect 3931 7814 3944 7844
rect 3959 7826 3989 7844
rect 4032 7814 4045 7844
rect 4075 7814 4088 7844
rect 4103 7826 4133 7844
rect 4176 7830 4190 7844
rect 4226 7830 4446 7844
rect 4177 7828 4190 7830
rect 4143 7816 4158 7828
rect 4140 7814 4162 7816
rect 4167 7814 4197 7828
rect 4258 7826 4411 7830
rect 4240 7814 4432 7826
rect 4475 7814 4505 7828
rect 4511 7814 4524 7844
rect 4539 7826 4569 7844
rect 4612 7814 4625 7844
rect 4655 7814 4668 7844
rect 4683 7826 4713 7844
rect 4756 7830 4770 7844
rect 4806 7830 5026 7844
rect 4757 7828 4770 7830
rect 4723 7816 4738 7828
rect 4720 7814 4742 7816
rect 4747 7814 4777 7828
rect 4838 7826 4991 7830
rect 4820 7814 5012 7826
rect 5055 7814 5085 7828
rect 5091 7814 5104 7844
rect 5119 7826 5149 7844
rect 5192 7814 5205 7844
rect 5235 7814 5248 7844
rect 5263 7826 5293 7844
rect 5336 7830 5350 7844
rect 5386 7830 5606 7844
rect 5337 7828 5350 7830
rect 5303 7816 5318 7828
rect 5300 7814 5322 7816
rect 5327 7814 5357 7828
rect 5418 7826 5571 7830
rect 5400 7814 5592 7826
rect 5635 7814 5665 7828
rect 5671 7814 5684 7844
rect 5699 7826 5729 7844
rect 5772 7814 5785 7844
rect 5815 7814 5828 7844
rect 5843 7826 5873 7844
rect 5916 7830 5930 7844
rect 5966 7830 6186 7844
rect 5917 7828 5930 7830
rect 5883 7816 5898 7828
rect 5880 7814 5902 7816
rect 5907 7814 5937 7828
rect 5998 7826 6151 7830
rect 5980 7814 6172 7826
rect 6215 7814 6245 7828
rect 6251 7814 6264 7844
rect 6279 7826 6309 7844
rect 6352 7814 6365 7844
rect 6395 7814 6408 7844
rect 6423 7826 6453 7844
rect 6496 7830 6510 7844
rect 6546 7830 6766 7844
rect 6497 7828 6510 7830
rect 6463 7816 6478 7828
rect 6460 7814 6482 7816
rect 6487 7814 6517 7828
rect 6578 7826 6731 7830
rect 6560 7814 6752 7826
rect 6795 7814 6825 7828
rect 6831 7814 6844 7844
rect 6859 7826 6889 7844
rect 6932 7814 6945 7844
rect 6975 7814 6988 7844
rect 7003 7826 7033 7844
rect 7076 7830 7090 7844
rect 7126 7830 7346 7844
rect 7077 7828 7090 7830
rect 7043 7816 7058 7828
rect 7040 7814 7062 7816
rect 7067 7814 7097 7828
rect 7158 7826 7311 7830
rect 7140 7814 7332 7826
rect 7375 7814 7405 7828
rect 7411 7814 7424 7844
rect 7439 7826 7469 7844
rect 7512 7814 7525 7844
rect 7555 7814 7568 7844
rect 7583 7826 7613 7844
rect 7656 7830 7670 7844
rect 7706 7830 7926 7844
rect 7657 7828 7670 7830
rect 7623 7816 7638 7828
rect 7620 7814 7642 7816
rect 7647 7814 7677 7828
rect 7738 7826 7891 7830
rect 7720 7814 7912 7826
rect 7955 7814 7985 7828
rect 7991 7814 8004 7844
rect 8019 7826 8049 7844
rect 8092 7814 8105 7844
rect 8135 7814 8148 7844
rect 8163 7826 8193 7844
rect 8236 7830 8250 7844
rect 8286 7830 8506 7844
rect 8237 7828 8250 7830
rect 8203 7816 8218 7828
rect 8200 7814 8222 7816
rect 8227 7814 8257 7828
rect 8318 7826 8471 7830
rect 8300 7814 8492 7826
rect 8535 7814 8565 7828
rect 8571 7814 8584 7844
rect 8599 7826 8629 7844
rect 8672 7814 8685 7844
rect 8715 7814 8728 7844
rect 8743 7826 8773 7844
rect 8816 7830 8830 7844
rect 8866 7830 9086 7844
rect 8817 7828 8830 7830
rect 8783 7816 8798 7828
rect 8780 7814 8802 7816
rect 8807 7814 8837 7828
rect 8898 7826 9051 7830
rect 8880 7814 9072 7826
rect 9115 7814 9145 7828
rect 9151 7814 9164 7844
rect 9179 7826 9209 7844
rect 9252 7814 9265 7844
rect 0 7800 9265 7814
rect 15 7696 28 7800
rect 73 7778 74 7788
rect 89 7778 102 7788
rect 73 7774 102 7778
rect 107 7774 137 7800
rect 155 7786 171 7788
rect 243 7786 296 7800
rect 244 7784 308 7786
rect 351 7784 366 7800
rect 415 7797 445 7800
rect 415 7794 451 7797
rect 381 7786 397 7788
rect 155 7774 170 7778
rect 73 7772 170 7774
rect 198 7772 366 7784
rect 382 7774 397 7778
rect 415 7775 454 7794
rect 473 7788 480 7789
rect 479 7781 480 7788
rect 463 7778 464 7781
rect 479 7778 492 7781
rect 415 7774 445 7775
rect 454 7774 460 7775
rect 463 7774 492 7778
rect 382 7773 492 7774
rect 382 7772 498 7773
rect 57 7764 108 7772
rect 57 7752 82 7764
rect 89 7752 108 7764
rect 139 7764 189 7772
rect 139 7756 155 7764
rect 162 7762 189 7764
rect 198 7762 419 7772
rect 162 7752 419 7762
rect 448 7764 498 7772
rect 448 7755 464 7764
rect 57 7744 108 7752
rect 155 7744 419 7752
rect 445 7752 464 7755
rect 471 7752 498 7764
rect 445 7744 498 7752
rect 73 7736 74 7744
rect 89 7736 102 7744
rect 73 7728 89 7736
rect 70 7721 89 7724
rect 70 7712 92 7721
rect 43 7702 92 7712
rect 43 7696 73 7702
rect 92 7697 97 7702
rect 15 7680 89 7696
rect 107 7688 137 7744
rect 172 7734 380 7744
rect 415 7740 460 7744
rect 463 7743 464 7744
rect 479 7743 492 7744
rect 198 7704 387 7734
rect 213 7701 387 7704
rect 206 7698 387 7701
rect 15 7678 28 7680
rect 43 7678 77 7680
rect 15 7662 89 7678
rect 116 7674 129 7688
rect 144 7674 160 7690
rect 206 7685 217 7698
rect -1 7640 0 7656
rect 15 7640 28 7662
rect 43 7640 73 7662
rect 116 7658 178 7674
rect 206 7667 217 7683
rect 222 7678 232 7698
rect 242 7678 256 7698
rect 259 7685 268 7698
rect 284 7685 293 7698
rect 222 7667 256 7678
rect 259 7667 268 7683
rect 284 7667 293 7683
rect 300 7678 310 7698
rect 320 7678 334 7698
rect 335 7685 346 7698
rect 300 7667 334 7678
rect 335 7667 346 7683
rect 392 7674 408 7690
rect 415 7688 445 7740
rect 479 7736 480 7743
rect 464 7728 480 7736
rect 451 7696 464 7715
rect 479 7696 509 7712
rect 451 7680 525 7696
rect 451 7678 464 7680
rect 479 7678 513 7680
rect 116 7656 129 7658
rect 144 7656 178 7658
rect 116 7640 178 7656
rect 222 7651 238 7654
rect 300 7651 330 7662
rect 378 7658 424 7674
rect 451 7662 525 7678
rect 378 7656 412 7658
rect 377 7640 424 7656
rect 451 7640 464 7662
rect 479 7640 509 7662
rect 536 7640 537 7656
rect 552 7640 565 7800
rect 595 7696 608 7800
rect 653 7778 654 7788
rect 669 7778 682 7788
rect 653 7774 682 7778
rect 687 7774 717 7800
rect 735 7786 751 7788
rect 823 7786 876 7800
rect 824 7784 888 7786
rect 931 7784 946 7800
rect 995 7797 1025 7800
rect 995 7794 1031 7797
rect 961 7786 977 7788
rect 735 7774 750 7778
rect 653 7772 750 7774
rect 778 7772 946 7784
rect 962 7774 977 7778
rect 995 7775 1034 7794
rect 1053 7788 1060 7789
rect 1059 7781 1060 7788
rect 1043 7778 1044 7781
rect 1059 7778 1072 7781
rect 995 7774 1025 7775
rect 1034 7774 1040 7775
rect 1043 7774 1072 7778
rect 962 7773 1072 7774
rect 962 7772 1078 7773
rect 637 7764 688 7772
rect 637 7752 662 7764
rect 669 7752 688 7764
rect 719 7764 769 7772
rect 719 7756 735 7764
rect 742 7762 769 7764
rect 778 7762 999 7772
rect 742 7752 999 7762
rect 1028 7764 1078 7772
rect 1028 7755 1044 7764
rect 637 7744 688 7752
rect 735 7744 999 7752
rect 1025 7752 1044 7755
rect 1051 7752 1078 7764
rect 1025 7744 1078 7752
rect 653 7736 654 7744
rect 669 7736 682 7744
rect 653 7728 669 7736
rect 650 7721 669 7724
rect 650 7712 672 7721
rect 623 7702 672 7712
rect 623 7696 653 7702
rect 672 7697 677 7702
rect 595 7680 669 7696
rect 687 7688 717 7744
rect 752 7734 960 7744
rect 995 7740 1040 7744
rect 1043 7743 1044 7744
rect 1059 7743 1072 7744
rect 778 7704 967 7734
rect 793 7701 967 7704
rect 786 7698 967 7701
rect 595 7678 608 7680
rect 623 7678 657 7680
rect 595 7662 669 7678
rect 696 7674 709 7688
rect 724 7674 740 7690
rect 786 7685 797 7698
rect 579 7640 580 7656
rect 595 7640 608 7662
rect 623 7640 653 7662
rect 696 7658 758 7674
rect 786 7667 797 7683
rect 802 7678 812 7698
rect 822 7678 836 7698
rect 839 7685 848 7698
rect 864 7685 873 7698
rect 802 7667 836 7678
rect 839 7667 848 7683
rect 864 7667 873 7683
rect 880 7678 890 7698
rect 900 7678 914 7698
rect 915 7685 926 7698
rect 880 7667 914 7678
rect 915 7667 926 7683
rect 972 7674 988 7690
rect 995 7688 1025 7740
rect 1059 7736 1060 7743
rect 1044 7728 1060 7736
rect 1031 7696 1044 7715
rect 1059 7696 1089 7712
rect 1031 7680 1105 7696
rect 1031 7678 1044 7680
rect 1059 7678 1093 7680
rect 696 7656 709 7658
rect 724 7656 758 7658
rect 696 7640 758 7656
rect 802 7651 818 7654
rect 880 7651 910 7662
rect 958 7658 1004 7674
rect 1031 7662 1105 7678
rect 958 7656 992 7658
rect 957 7640 1004 7656
rect 1031 7640 1044 7662
rect 1059 7640 1089 7662
rect 1116 7640 1117 7656
rect 1132 7640 1145 7800
rect 1175 7696 1188 7800
rect 1233 7778 1234 7788
rect 1249 7778 1262 7788
rect 1233 7774 1262 7778
rect 1267 7774 1297 7800
rect 1315 7786 1331 7788
rect 1403 7786 1456 7800
rect 1404 7784 1468 7786
rect 1511 7784 1526 7800
rect 1575 7797 1605 7800
rect 1575 7794 1611 7797
rect 1541 7786 1557 7788
rect 1315 7774 1330 7778
rect 1233 7772 1330 7774
rect 1358 7772 1526 7784
rect 1542 7774 1557 7778
rect 1575 7775 1614 7794
rect 1633 7788 1640 7789
rect 1639 7781 1640 7788
rect 1623 7778 1624 7781
rect 1639 7778 1652 7781
rect 1575 7774 1605 7775
rect 1614 7774 1620 7775
rect 1623 7774 1652 7778
rect 1542 7773 1652 7774
rect 1542 7772 1658 7773
rect 1217 7764 1268 7772
rect 1217 7752 1242 7764
rect 1249 7752 1268 7764
rect 1299 7764 1349 7772
rect 1299 7756 1315 7764
rect 1322 7762 1349 7764
rect 1358 7762 1579 7772
rect 1322 7752 1579 7762
rect 1608 7764 1658 7772
rect 1608 7755 1624 7764
rect 1217 7744 1268 7752
rect 1315 7744 1579 7752
rect 1605 7752 1624 7755
rect 1631 7752 1658 7764
rect 1605 7744 1658 7752
rect 1233 7736 1234 7744
rect 1249 7736 1262 7744
rect 1233 7728 1249 7736
rect 1230 7721 1249 7724
rect 1230 7712 1252 7721
rect 1203 7702 1252 7712
rect 1203 7696 1233 7702
rect 1252 7697 1257 7702
rect 1175 7680 1249 7696
rect 1267 7688 1297 7744
rect 1332 7734 1540 7744
rect 1575 7740 1620 7744
rect 1623 7743 1624 7744
rect 1639 7743 1652 7744
rect 1358 7704 1547 7734
rect 1373 7701 1547 7704
rect 1366 7698 1547 7701
rect 1175 7678 1188 7680
rect 1203 7678 1237 7680
rect 1175 7662 1249 7678
rect 1276 7674 1289 7688
rect 1304 7674 1320 7690
rect 1366 7685 1377 7698
rect 1159 7640 1160 7656
rect 1175 7640 1188 7662
rect 1203 7640 1233 7662
rect 1276 7658 1338 7674
rect 1366 7667 1377 7683
rect 1382 7678 1392 7698
rect 1402 7678 1416 7698
rect 1419 7685 1428 7698
rect 1444 7685 1453 7698
rect 1382 7667 1416 7678
rect 1419 7667 1428 7683
rect 1444 7667 1453 7683
rect 1460 7678 1470 7698
rect 1480 7678 1494 7698
rect 1495 7685 1506 7698
rect 1460 7667 1494 7678
rect 1495 7667 1506 7683
rect 1552 7674 1568 7690
rect 1575 7688 1605 7740
rect 1639 7736 1640 7743
rect 1624 7728 1640 7736
rect 1611 7696 1624 7715
rect 1639 7696 1669 7712
rect 1611 7680 1685 7696
rect 1611 7678 1624 7680
rect 1639 7678 1673 7680
rect 1276 7656 1289 7658
rect 1304 7656 1338 7658
rect 1276 7640 1338 7656
rect 1382 7651 1398 7654
rect 1460 7651 1490 7662
rect 1538 7658 1584 7674
rect 1611 7662 1685 7678
rect 1538 7656 1572 7658
rect 1537 7640 1584 7656
rect 1611 7640 1624 7662
rect 1639 7640 1669 7662
rect 1696 7640 1697 7656
rect 1712 7640 1725 7800
rect 1755 7696 1768 7800
rect 1813 7778 1814 7788
rect 1829 7778 1842 7788
rect 1813 7774 1842 7778
rect 1847 7774 1877 7800
rect 1895 7786 1911 7788
rect 1983 7786 2036 7800
rect 1984 7784 2048 7786
rect 2091 7784 2106 7800
rect 2155 7797 2185 7800
rect 2155 7794 2191 7797
rect 2121 7786 2137 7788
rect 1895 7774 1910 7778
rect 1813 7772 1910 7774
rect 1938 7772 2106 7784
rect 2122 7774 2137 7778
rect 2155 7775 2194 7794
rect 2213 7788 2220 7789
rect 2219 7781 2220 7788
rect 2203 7778 2204 7781
rect 2219 7778 2232 7781
rect 2155 7774 2185 7775
rect 2194 7774 2200 7775
rect 2203 7774 2232 7778
rect 2122 7773 2232 7774
rect 2122 7772 2238 7773
rect 1797 7764 1848 7772
rect 1797 7752 1822 7764
rect 1829 7752 1848 7764
rect 1879 7764 1929 7772
rect 1879 7756 1895 7764
rect 1902 7762 1929 7764
rect 1938 7762 2159 7772
rect 1902 7752 2159 7762
rect 2188 7764 2238 7772
rect 2188 7755 2204 7764
rect 1797 7744 1848 7752
rect 1895 7744 2159 7752
rect 2185 7752 2204 7755
rect 2211 7752 2238 7764
rect 2185 7744 2238 7752
rect 1813 7736 1814 7744
rect 1829 7736 1842 7744
rect 1813 7728 1829 7736
rect 1810 7721 1829 7724
rect 1810 7712 1832 7721
rect 1783 7702 1832 7712
rect 1783 7696 1813 7702
rect 1832 7697 1837 7702
rect 1755 7680 1829 7696
rect 1847 7688 1877 7744
rect 1912 7734 2120 7744
rect 2155 7740 2200 7744
rect 2203 7743 2204 7744
rect 2219 7743 2232 7744
rect 1938 7704 2127 7734
rect 1953 7701 2127 7704
rect 1946 7698 2127 7701
rect 1755 7678 1768 7680
rect 1783 7678 1817 7680
rect 1755 7662 1829 7678
rect 1856 7674 1869 7688
rect 1884 7674 1900 7690
rect 1946 7685 1957 7698
rect 1739 7640 1740 7656
rect 1755 7640 1768 7662
rect 1783 7640 1813 7662
rect 1856 7658 1918 7674
rect 1946 7667 1957 7683
rect 1962 7678 1972 7698
rect 1982 7678 1996 7698
rect 1999 7685 2008 7698
rect 2024 7685 2033 7698
rect 1962 7667 1996 7678
rect 1999 7667 2008 7683
rect 2024 7667 2033 7683
rect 2040 7678 2050 7698
rect 2060 7678 2074 7698
rect 2075 7685 2086 7698
rect 2040 7667 2074 7678
rect 2075 7667 2086 7683
rect 2132 7674 2148 7690
rect 2155 7688 2185 7740
rect 2219 7736 2220 7743
rect 2204 7728 2220 7736
rect 2191 7696 2204 7715
rect 2219 7696 2249 7712
rect 2191 7680 2265 7696
rect 2191 7678 2204 7680
rect 2219 7678 2253 7680
rect 1856 7656 1869 7658
rect 1884 7656 1918 7658
rect 1856 7640 1918 7656
rect 1962 7651 1976 7654
rect 2040 7651 2070 7662
rect 2118 7658 2164 7674
rect 2191 7662 2265 7678
rect 2118 7656 2152 7658
rect 2117 7640 2164 7656
rect 2191 7640 2204 7662
rect 2219 7640 2249 7662
rect 2276 7640 2277 7656
rect 2292 7640 2305 7800
rect 2335 7696 2348 7800
rect 2393 7778 2394 7788
rect 2409 7778 2422 7788
rect 2393 7774 2422 7778
rect 2427 7774 2457 7800
rect 2475 7786 2491 7788
rect 2563 7786 2616 7800
rect 2564 7784 2628 7786
rect 2671 7784 2686 7800
rect 2735 7797 2765 7800
rect 2735 7794 2771 7797
rect 2701 7786 2717 7788
rect 2475 7774 2490 7778
rect 2393 7772 2490 7774
rect 2518 7772 2686 7784
rect 2702 7774 2717 7778
rect 2735 7775 2774 7794
rect 2793 7788 2800 7789
rect 2799 7781 2800 7788
rect 2783 7778 2784 7781
rect 2799 7778 2812 7781
rect 2735 7774 2765 7775
rect 2774 7774 2780 7775
rect 2783 7774 2812 7778
rect 2702 7773 2812 7774
rect 2702 7772 2818 7773
rect 2377 7764 2428 7772
rect 2377 7752 2402 7764
rect 2409 7752 2428 7764
rect 2459 7764 2509 7772
rect 2459 7756 2475 7764
rect 2482 7762 2509 7764
rect 2518 7762 2739 7772
rect 2482 7752 2739 7762
rect 2768 7764 2818 7772
rect 2768 7755 2784 7764
rect 2377 7744 2428 7752
rect 2475 7744 2739 7752
rect 2765 7752 2784 7755
rect 2791 7752 2818 7764
rect 2765 7744 2818 7752
rect 2393 7736 2394 7744
rect 2409 7736 2422 7744
rect 2393 7728 2409 7736
rect 2390 7721 2409 7724
rect 2390 7712 2412 7721
rect 2363 7702 2412 7712
rect 2363 7696 2393 7702
rect 2412 7697 2417 7702
rect 2335 7680 2409 7696
rect 2427 7688 2457 7744
rect 2492 7734 2700 7744
rect 2735 7740 2780 7744
rect 2783 7743 2784 7744
rect 2799 7743 2812 7744
rect 2518 7704 2707 7734
rect 2533 7701 2707 7704
rect 2526 7698 2707 7701
rect 2335 7678 2348 7680
rect 2363 7678 2397 7680
rect 2335 7662 2409 7678
rect 2436 7674 2449 7688
rect 2464 7674 2480 7690
rect 2526 7685 2537 7698
rect 2319 7640 2320 7656
rect 2335 7640 2348 7662
rect 2363 7640 2393 7662
rect 2436 7658 2498 7674
rect 2526 7667 2537 7683
rect 2542 7678 2552 7698
rect 2562 7678 2576 7698
rect 2579 7685 2588 7698
rect 2604 7685 2613 7698
rect 2542 7667 2576 7678
rect 2579 7667 2588 7683
rect 2604 7667 2613 7683
rect 2620 7678 2630 7698
rect 2640 7678 2654 7698
rect 2655 7685 2666 7698
rect 2620 7667 2654 7678
rect 2655 7667 2666 7683
rect 2712 7674 2728 7690
rect 2735 7688 2765 7740
rect 2799 7736 2800 7743
rect 2784 7728 2800 7736
rect 2771 7696 2784 7715
rect 2799 7696 2829 7712
rect 2771 7680 2845 7696
rect 2771 7678 2784 7680
rect 2799 7678 2833 7680
rect 2436 7656 2449 7658
rect 2464 7656 2498 7658
rect 2436 7640 2498 7656
rect 2542 7651 2558 7654
rect 2620 7651 2650 7662
rect 2698 7658 2744 7674
rect 2771 7662 2845 7678
rect 2698 7656 2732 7658
rect 2697 7640 2744 7656
rect 2771 7640 2784 7662
rect 2799 7640 2829 7662
rect 2856 7640 2857 7656
rect 2872 7640 2885 7800
rect 2915 7696 2928 7800
rect 2973 7778 2974 7788
rect 2989 7778 3002 7788
rect 2973 7774 3002 7778
rect 3007 7774 3037 7800
rect 3055 7786 3071 7788
rect 3143 7786 3196 7800
rect 3144 7784 3208 7786
rect 3251 7784 3266 7800
rect 3315 7797 3345 7800
rect 3315 7794 3351 7797
rect 3281 7786 3297 7788
rect 3055 7774 3070 7778
rect 2973 7772 3070 7774
rect 3098 7772 3266 7784
rect 3282 7774 3297 7778
rect 3315 7775 3354 7794
rect 3373 7788 3380 7789
rect 3379 7781 3380 7788
rect 3363 7778 3364 7781
rect 3379 7778 3392 7781
rect 3315 7774 3345 7775
rect 3354 7774 3360 7775
rect 3363 7774 3392 7778
rect 3282 7773 3392 7774
rect 3282 7772 3398 7773
rect 2957 7764 3008 7772
rect 2957 7752 2982 7764
rect 2989 7752 3008 7764
rect 3039 7764 3089 7772
rect 3039 7756 3055 7764
rect 3062 7762 3089 7764
rect 3098 7762 3319 7772
rect 3062 7752 3319 7762
rect 3348 7764 3398 7772
rect 3348 7755 3364 7764
rect 2957 7744 3008 7752
rect 3055 7744 3319 7752
rect 3345 7752 3364 7755
rect 3371 7752 3398 7764
rect 3345 7744 3398 7752
rect 2973 7736 2974 7744
rect 2989 7736 3002 7744
rect 2973 7728 2989 7736
rect 2970 7721 2989 7724
rect 2970 7712 2992 7721
rect 2943 7702 2992 7712
rect 2943 7696 2973 7702
rect 2992 7697 2997 7702
rect 2915 7680 2989 7696
rect 3007 7688 3037 7744
rect 3072 7734 3280 7744
rect 3315 7740 3360 7744
rect 3363 7743 3364 7744
rect 3379 7743 3392 7744
rect 3098 7704 3287 7734
rect 3113 7701 3287 7704
rect 3106 7698 3287 7701
rect 2915 7678 2928 7680
rect 2943 7678 2977 7680
rect 2915 7662 2989 7678
rect 3016 7674 3029 7688
rect 3044 7674 3060 7690
rect 3106 7685 3117 7698
rect 2899 7640 2900 7656
rect 2915 7640 2928 7662
rect 2943 7640 2973 7662
rect 3016 7658 3078 7674
rect 3106 7667 3117 7683
rect 3122 7678 3132 7698
rect 3142 7678 3156 7698
rect 3159 7685 3168 7698
rect 3184 7685 3193 7698
rect 3122 7667 3156 7678
rect 3159 7667 3168 7683
rect 3184 7667 3193 7683
rect 3200 7678 3210 7698
rect 3220 7678 3234 7698
rect 3235 7685 3246 7698
rect 3200 7667 3234 7678
rect 3235 7667 3246 7683
rect 3292 7674 3308 7690
rect 3315 7688 3345 7740
rect 3379 7736 3380 7743
rect 3364 7728 3380 7736
rect 3351 7696 3364 7715
rect 3379 7696 3409 7712
rect 3351 7680 3425 7696
rect 3351 7678 3364 7680
rect 3379 7678 3413 7680
rect 3016 7656 3029 7658
rect 3044 7656 3078 7658
rect 3016 7640 3078 7656
rect 3122 7651 3138 7654
rect 3200 7651 3230 7662
rect 3278 7658 3324 7674
rect 3351 7662 3425 7678
rect 3278 7656 3312 7658
rect 3277 7640 3324 7656
rect 3351 7640 3364 7662
rect 3379 7640 3409 7662
rect 3436 7640 3437 7656
rect 3452 7640 3465 7800
rect 3495 7696 3508 7800
rect 3553 7778 3554 7788
rect 3569 7778 3582 7788
rect 3553 7774 3582 7778
rect 3587 7774 3617 7800
rect 3635 7786 3651 7788
rect 3723 7786 3776 7800
rect 3724 7784 3788 7786
rect 3831 7784 3846 7800
rect 3895 7797 3925 7800
rect 3895 7794 3931 7797
rect 3861 7786 3877 7788
rect 3635 7774 3650 7778
rect 3553 7772 3650 7774
rect 3678 7772 3846 7784
rect 3862 7774 3877 7778
rect 3895 7775 3934 7794
rect 3953 7788 3960 7789
rect 3959 7781 3960 7788
rect 3943 7778 3944 7781
rect 3959 7778 3972 7781
rect 3895 7774 3925 7775
rect 3934 7774 3940 7775
rect 3943 7774 3972 7778
rect 3862 7773 3972 7774
rect 3862 7772 3978 7773
rect 3537 7764 3588 7772
rect 3537 7752 3562 7764
rect 3569 7752 3588 7764
rect 3619 7764 3669 7772
rect 3619 7756 3635 7764
rect 3642 7762 3669 7764
rect 3678 7762 3899 7772
rect 3642 7752 3899 7762
rect 3928 7764 3978 7772
rect 3928 7755 3944 7764
rect 3537 7744 3588 7752
rect 3635 7744 3899 7752
rect 3925 7752 3944 7755
rect 3951 7752 3978 7764
rect 3925 7744 3978 7752
rect 3553 7736 3554 7744
rect 3569 7736 3582 7744
rect 3553 7728 3569 7736
rect 3550 7721 3569 7724
rect 3550 7712 3572 7721
rect 3523 7702 3572 7712
rect 3523 7696 3553 7702
rect 3572 7697 3577 7702
rect 3495 7680 3569 7696
rect 3587 7688 3617 7744
rect 3652 7734 3860 7744
rect 3895 7740 3940 7744
rect 3943 7743 3944 7744
rect 3959 7743 3972 7744
rect 3678 7704 3867 7734
rect 3693 7701 3867 7704
rect 3686 7698 3867 7701
rect 3495 7678 3508 7680
rect 3523 7678 3557 7680
rect 3495 7662 3569 7678
rect 3596 7674 3609 7688
rect 3624 7674 3640 7690
rect 3686 7685 3697 7698
rect 3479 7640 3480 7656
rect 3495 7640 3508 7662
rect 3523 7640 3553 7662
rect 3596 7658 3658 7674
rect 3686 7667 3697 7683
rect 3702 7678 3712 7698
rect 3722 7678 3736 7698
rect 3739 7685 3748 7698
rect 3764 7685 3773 7698
rect 3702 7667 3736 7678
rect 3739 7667 3748 7683
rect 3764 7667 3773 7683
rect 3780 7678 3790 7698
rect 3800 7678 3814 7698
rect 3815 7685 3826 7698
rect 3780 7667 3814 7678
rect 3815 7667 3826 7683
rect 3872 7674 3888 7690
rect 3895 7688 3925 7740
rect 3959 7736 3960 7743
rect 3944 7728 3960 7736
rect 3931 7696 3944 7715
rect 3959 7696 3989 7712
rect 3931 7680 4005 7696
rect 3931 7678 3944 7680
rect 3959 7678 3993 7680
rect 3596 7656 3609 7658
rect 3624 7656 3658 7658
rect 3596 7640 3658 7656
rect 3702 7651 3718 7654
rect 3780 7651 3810 7662
rect 3858 7658 3904 7674
rect 3931 7662 4005 7678
rect 3858 7656 3892 7658
rect 3857 7640 3904 7656
rect 3931 7640 3944 7662
rect 3959 7640 3989 7662
rect 4016 7640 4017 7656
rect 4032 7640 4045 7800
rect 4075 7696 4088 7800
rect 4133 7778 4134 7788
rect 4149 7778 4162 7788
rect 4133 7774 4162 7778
rect 4167 7774 4197 7800
rect 4215 7786 4231 7788
rect 4303 7786 4356 7800
rect 4304 7784 4368 7786
rect 4411 7784 4426 7800
rect 4475 7797 4505 7800
rect 4475 7794 4511 7797
rect 4441 7786 4457 7788
rect 4215 7774 4230 7778
rect 4133 7772 4230 7774
rect 4258 7772 4426 7784
rect 4442 7774 4457 7778
rect 4475 7775 4514 7794
rect 4533 7788 4540 7789
rect 4539 7781 4540 7788
rect 4523 7778 4524 7781
rect 4539 7778 4552 7781
rect 4475 7774 4505 7775
rect 4514 7774 4520 7775
rect 4523 7774 4552 7778
rect 4442 7773 4552 7774
rect 4442 7772 4558 7773
rect 4117 7764 4168 7772
rect 4117 7752 4142 7764
rect 4149 7752 4168 7764
rect 4199 7764 4249 7772
rect 4199 7756 4215 7764
rect 4222 7762 4249 7764
rect 4258 7762 4479 7772
rect 4222 7752 4479 7762
rect 4508 7764 4558 7772
rect 4508 7755 4524 7764
rect 4117 7744 4168 7752
rect 4215 7744 4479 7752
rect 4505 7752 4524 7755
rect 4531 7752 4558 7764
rect 4505 7744 4558 7752
rect 4133 7736 4134 7744
rect 4149 7736 4162 7744
rect 4133 7728 4149 7736
rect 4130 7721 4149 7724
rect 4130 7712 4152 7721
rect 4103 7702 4152 7712
rect 4103 7696 4133 7702
rect 4152 7697 4157 7702
rect 4075 7680 4149 7696
rect 4167 7688 4197 7744
rect 4232 7734 4440 7744
rect 4475 7740 4520 7744
rect 4523 7743 4524 7744
rect 4539 7743 4552 7744
rect 4258 7704 4447 7734
rect 4273 7701 4447 7704
rect 4266 7698 4447 7701
rect 4075 7678 4088 7680
rect 4103 7678 4137 7680
rect 4075 7662 4149 7678
rect 4176 7674 4189 7688
rect 4204 7674 4220 7690
rect 4266 7685 4277 7698
rect 4059 7640 4060 7656
rect 4075 7640 4088 7662
rect 4103 7640 4133 7662
rect 4176 7658 4238 7674
rect 4266 7667 4277 7683
rect 4282 7678 4292 7698
rect 4302 7678 4316 7698
rect 4319 7685 4328 7698
rect 4344 7685 4353 7698
rect 4282 7667 4316 7678
rect 4319 7667 4328 7683
rect 4344 7667 4353 7683
rect 4360 7678 4370 7698
rect 4380 7678 4394 7698
rect 4395 7685 4406 7698
rect 4360 7667 4394 7678
rect 4395 7667 4406 7683
rect 4452 7674 4468 7690
rect 4475 7688 4505 7740
rect 4539 7736 4540 7743
rect 4524 7728 4540 7736
rect 4511 7696 4524 7715
rect 4539 7696 4569 7712
rect 4511 7680 4585 7696
rect 4511 7678 4524 7680
rect 4539 7678 4573 7680
rect 4176 7656 4189 7658
rect 4204 7656 4238 7658
rect 4176 7640 4238 7656
rect 4282 7651 4298 7654
rect 4360 7651 4390 7662
rect 4438 7658 4484 7674
rect 4511 7662 4585 7678
rect 4438 7656 4472 7658
rect 4437 7640 4484 7656
rect 4511 7640 4524 7662
rect 4539 7640 4569 7662
rect 4596 7640 4597 7656
rect 4612 7640 4625 7800
rect 4655 7696 4668 7800
rect 4713 7778 4714 7788
rect 4729 7778 4742 7788
rect 4713 7774 4742 7778
rect 4747 7774 4777 7800
rect 4795 7786 4811 7788
rect 4883 7786 4936 7800
rect 4884 7784 4948 7786
rect 4991 7784 5006 7800
rect 5055 7797 5085 7800
rect 5055 7794 5091 7797
rect 5021 7786 5037 7788
rect 4795 7774 4810 7778
rect 4713 7772 4810 7774
rect 4838 7772 5006 7784
rect 5022 7774 5037 7778
rect 5055 7775 5094 7794
rect 5113 7788 5120 7789
rect 5119 7781 5120 7788
rect 5103 7778 5104 7781
rect 5119 7778 5132 7781
rect 5055 7774 5085 7775
rect 5094 7774 5100 7775
rect 5103 7774 5132 7778
rect 5022 7773 5132 7774
rect 5022 7772 5138 7773
rect 4697 7764 4748 7772
rect 4697 7752 4722 7764
rect 4729 7752 4748 7764
rect 4779 7764 4829 7772
rect 4779 7756 4795 7764
rect 4802 7762 4829 7764
rect 4838 7762 5059 7772
rect 4802 7752 5059 7762
rect 5088 7764 5138 7772
rect 5088 7755 5104 7764
rect 4697 7744 4748 7752
rect 4795 7744 5059 7752
rect 5085 7752 5104 7755
rect 5111 7752 5138 7764
rect 5085 7744 5138 7752
rect 4713 7736 4714 7744
rect 4729 7736 4742 7744
rect 4713 7728 4729 7736
rect 4710 7721 4729 7724
rect 4710 7712 4732 7721
rect 4683 7702 4732 7712
rect 4683 7696 4713 7702
rect 4732 7697 4737 7702
rect 4655 7680 4729 7696
rect 4747 7688 4777 7744
rect 4812 7734 5020 7744
rect 5055 7740 5100 7744
rect 5103 7743 5104 7744
rect 5119 7743 5132 7744
rect 4838 7704 5027 7734
rect 4853 7701 5027 7704
rect 4846 7698 5027 7701
rect 4655 7678 4668 7680
rect 4683 7678 4717 7680
rect 4655 7662 4729 7678
rect 4756 7674 4769 7688
rect 4784 7674 4800 7690
rect 4846 7685 4857 7698
rect 4639 7640 4640 7656
rect 4655 7640 4668 7662
rect 4683 7640 4713 7662
rect 4756 7658 4818 7674
rect 4846 7667 4857 7683
rect 4862 7678 4872 7698
rect 4882 7678 4896 7698
rect 4899 7685 4908 7698
rect 4924 7685 4933 7698
rect 4862 7667 4896 7678
rect 4899 7667 4908 7683
rect 4924 7667 4933 7683
rect 4940 7678 4950 7698
rect 4960 7678 4974 7698
rect 4975 7685 4986 7698
rect 4940 7667 4974 7678
rect 4975 7667 4986 7683
rect 5032 7674 5048 7690
rect 5055 7688 5085 7740
rect 5119 7736 5120 7743
rect 5104 7728 5120 7736
rect 5091 7696 5104 7715
rect 5119 7696 5149 7712
rect 5091 7680 5165 7696
rect 5091 7678 5104 7680
rect 5119 7678 5153 7680
rect 4756 7656 4769 7658
rect 4784 7656 4818 7658
rect 4756 7640 4818 7656
rect 4862 7651 4878 7654
rect 4940 7651 4970 7662
rect 5018 7658 5064 7674
rect 5091 7662 5165 7678
rect 5018 7656 5052 7658
rect 5017 7640 5064 7656
rect 5091 7640 5104 7662
rect 5119 7640 5149 7662
rect 5176 7640 5177 7656
rect 5192 7640 5205 7800
rect 5235 7696 5248 7800
rect 5293 7778 5294 7788
rect 5309 7778 5322 7788
rect 5293 7774 5322 7778
rect 5327 7774 5357 7800
rect 5375 7786 5391 7788
rect 5463 7786 5516 7800
rect 5464 7784 5528 7786
rect 5571 7784 5586 7800
rect 5635 7797 5665 7800
rect 5635 7794 5671 7797
rect 5601 7786 5617 7788
rect 5375 7774 5390 7778
rect 5293 7772 5390 7774
rect 5418 7772 5586 7784
rect 5602 7774 5617 7778
rect 5635 7775 5674 7794
rect 5693 7788 5700 7789
rect 5699 7781 5700 7788
rect 5683 7778 5684 7781
rect 5699 7778 5712 7781
rect 5635 7774 5665 7775
rect 5674 7774 5680 7775
rect 5683 7774 5712 7778
rect 5602 7773 5712 7774
rect 5602 7772 5718 7773
rect 5277 7764 5328 7772
rect 5277 7752 5302 7764
rect 5309 7752 5328 7764
rect 5359 7764 5409 7772
rect 5359 7756 5375 7764
rect 5382 7762 5409 7764
rect 5418 7762 5639 7772
rect 5382 7752 5639 7762
rect 5668 7764 5718 7772
rect 5668 7755 5684 7764
rect 5277 7744 5328 7752
rect 5375 7744 5639 7752
rect 5665 7752 5684 7755
rect 5691 7752 5718 7764
rect 5665 7744 5718 7752
rect 5293 7736 5294 7744
rect 5309 7736 5322 7744
rect 5293 7728 5309 7736
rect 5290 7721 5309 7724
rect 5290 7712 5312 7721
rect 5263 7702 5312 7712
rect 5263 7696 5293 7702
rect 5312 7697 5317 7702
rect 5235 7680 5309 7696
rect 5327 7688 5357 7744
rect 5392 7734 5600 7744
rect 5635 7740 5680 7744
rect 5683 7743 5684 7744
rect 5699 7743 5712 7744
rect 5418 7704 5607 7734
rect 5433 7701 5607 7704
rect 5426 7698 5607 7701
rect 5235 7678 5248 7680
rect 5263 7678 5297 7680
rect 5235 7662 5309 7678
rect 5336 7674 5349 7688
rect 5364 7674 5380 7690
rect 5426 7685 5437 7698
rect 5219 7640 5220 7656
rect 5235 7640 5248 7662
rect 5263 7640 5293 7662
rect 5336 7658 5398 7674
rect 5426 7667 5437 7683
rect 5442 7678 5452 7698
rect 5462 7678 5476 7698
rect 5479 7685 5488 7698
rect 5504 7685 5513 7698
rect 5442 7667 5476 7678
rect 5479 7667 5488 7683
rect 5504 7667 5513 7683
rect 5520 7678 5530 7698
rect 5540 7678 5554 7698
rect 5555 7685 5566 7698
rect 5520 7667 5554 7678
rect 5555 7667 5566 7683
rect 5612 7674 5628 7690
rect 5635 7688 5665 7740
rect 5699 7736 5700 7743
rect 5684 7728 5700 7736
rect 5671 7696 5684 7715
rect 5699 7696 5729 7712
rect 5671 7680 5745 7696
rect 5671 7678 5684 7680
rect 5699 7678 5733 7680
rect 5336 7656 5349 7658
rect 5364 7656 5398 7658
rect 5336 7640 5398 7656
rect 5442 7651 5458 7654
rect 5520 7651 5550 7662
rect 5598 7658 5644 7674
rect 5671 7662 5745 7678
rect 5598 7656 5632 7658
rect 5597 7640 5644 7656
rect 5671 7640 5684 7662
rect 5699 7640 5729 7662
rect 5756 7640 5757 7656
rect 5772 7640 5785 7800
rect 5815 7696 5828 7800
rect 5873 7778 5874 7788
rect 5889 7778 5902 7788
rect 5873 7774 5902 7778
rect 5907 7774 5937 7800
rect 5955 7786 5971 7788
rect 6043 7786 6096 7800
rect 6044 7784 6108 7786
rect 6151 7784 6166 7800
rect 6215 7797 6245 7800
rect 6215 7794 6251 7797
rect 6181 7786 6197 7788
rect 5955 7774 5970 7778
rect 5873 7772 5970 7774
rect 5998 7772 6166 7784
rect 6182 7774 6197 7778
rect 6215 7775 6254 7794
rect 6273 7788 6280 7789
rect 6279 7781 6280 7788
rect 6263 7778 6264 7781
rect 6279 7778 6292 7781
rect 6215 7774 6245 7775
rect 6254 7774 6260 7775
rect 6263 7774 6292 7778
rect 6182 7773 6292 7774
rect 6182 7772 6298 7773
rect 5857 7764 5908 7772
rect 5857 7752 5882 7764
rect 5889 7752 5908 7764
rect 5939 7764 5989 7772
rect 5939 7756 5955 7764
rect 5962 7762 5989 7764
rect 5998 7762 6219 7772
rect 5962 7752 6219 7762
rect 6248 7764 6298 7772
rect 6248 7755 6264 7764
rect 5857 7744 5908 7752
rect 5955 7744 6219 7752
rect 6245 7752 6264 7755
rect 6271 7752 6298 7764
rect 6245 7744 6298 7752
rect 5873 7736 5874 7744
rect 5889 7736 5902 7744
rect 5873 7728 5889 7736
rect 5870 7721 5889 7724
rect 5870 7712 5892 7721
rect 5843 7702 5892 7712
rect 5843 7696 5873 7702
rect 5892 7697 5897 7702
rect 5815 7680 5889 7696
rect 5907 7688 5937 7744
rect 5972 7734 6180 7744
rect 6215 7740 6260 7744
rect 6263 7743 6264 7744
rect 6279 7743 6292 7744
rect 5998 7704 6187 7734
rect 6013 7701 6187 7704
rect 6006 7698 6187 7701
rect 5815 7678 5828 7680
rect 5843 7678 5877 7680
rect 5815 7662 5889 7678
rect 5916 7674 5929 7688
rect 5944 7674 5960 7690
rect 6006 7685 6017 7698
rect 5799 7640 5800 7656
rect 5815 7640 5828 7662
rect 5843 7640 5873 7662
rect 5916 7658 5978 7674
rect 6006 7667 6017 7683
rect 6022 7678 6032 7698
rect 6042 7678 6056 7698
rect 6059 7685 6068 7698
rect 6084 7685 6093 7698
rect 6022 7667 6056 7678
rect 6059 7667 6068 7683
rect 6084 7667 6093 7683
rect 6100 7678 6110 7698
rect 6120 7678 6134 7698
rect 6135 7685 6146 7698
rect 6100 7667 6134 7678
rect 6135 7667 6146 7683
rect 6192 7674 6208 7690
rect 6215 7688 6245 7740
rect 6279 7736 6280 7743
rect 6264 7728 6280 7736
rect 6251 7696 6264 7715
rect 6279 7696 6309 7712
rect 6251 7680 6325 7696
rect 6251 7678 6264 7680
rect 6279 7678 6313 7680
rect 5916 7656 5929 7658
rect 5944 7656 5978 7658
rect 5916 7640 5978 7656
rect 6022 7651 6038 7654
rect 6100 7651 6130 7662
rect 6178 7658 6224 7674
rect 6251 7662 6325 7678
rect 6178 7656 6212 7658
rect 6177 7640 6224 7656
rect 6251 7640 6264 7662
rect 6279 7640 6309 7662
rect 6336 7640 6337 7656
rect 6352 7640 6365 7800
rect 6395 7696 6408 7800
rect 6453 7778 6454 7788
rect 6469 7778 6482 7788
rect 6453 7774 6482 7778
rect 6487 7774 6517 7800
rect 6535 7786 6551 7788
rect 6623 7786 6676 7800
rect 6624 7784 6688 7786
rect 6731 7784 6746 7800
rect 6795 7797 6825 7800
rect 6795 7794 6831 7797
rect 6761 7786 6777 7788
rect 6535 7774 6550 7778
rect 6453 7772 6550 7774
rect 6578 7772 6746 7784
rect 6762 7774 6777 7778
rect 6795 7775 6834 7794
rect 6853 7788 6860 7789
rect 6859 7781 6860 7788
rect 6843 7778 6844 7781
rect 6859 7778 6872 7781
rect 6795 7774 6825 7775
rect 6834 7774 6840 7775
rect 6843 7774 6872 7778
rect 6762 7773 6872 7774
rect 6762 7772 6878 7773
rect 6437 7764 6488 7772
rect 6437 7752 6462 7764
rect 6469 7752 6488 7764
rect 6519 7764 6569 7772
rect 6519 7756 6535 7764
rect 6542 7762 6569 7764
rect 6578 7762 6799 7772
rect 6542 7752 6799 7762
rect 6828 7764 6878 7772
rect 6828 7755 6844 7764
rect 6437 7744 6488 7752
rect 6535 7744 6799 7752
rect 6825 7752 6844 7755
rect 6851 7752 6878 7764
rect 6825 7744 6878 7752
rect 6453 7736 6454 7744
rect 6469 7736 6482 7744
rect 6453 7728 6469 7736
rect 6450 7721 6469 7724
rect 6450 7712 6472 7721
rect 6423 7702 6472 7712
rect 6423 7696 6453 7702
rect 6472 7697 6477 7702
rect 6395 7680 6469 7696
rect 6487 7688 6517 7744
rect 6552 7734 6760 7744
rect 6795 7740 6840 7744
rect 6843 7743 6844 7744
rect 6859 7743 6872 7744
rect 6578 7704 6767 7734
rect 6593 7701 6767 7704
rect 6586 7698 6767 7701
rect 6395 7678 6408 7680
rect 6423 7678 6457 7680
rect 6395 7662 6469 7678
rect 6496 7674 6509 7688
rect 6524 7674 6540 7690
rect 6586 7685 6597 7698
rect 6379 7640 6380 7656
rect 6395 7640 6408 7662
rect 6423 7640 6453 7662
rect 6496 7658 6558 7674
rect 6586 7667 6597 7683
rect 6602 7678 6612 7698
rect 6622 7678 6636 7698
rect 6639 7685 6648 7698
rect 6664 7685 6673 7698
rect 6602 7667 6636 7678
rect 6639 7667 6648 7683
rect 6664 7667 6673 7683
rect 6680 7678 6690 7698
rect 6700 7678 6714 7698
rect 6715 7685 6726 7698
rect 6680 7667 6714 7678
rect 6715 7667 6726 7683
rect 6772 7674 6788 7690
rect 6795 7688 6825 7740
rect 6859 7736 6860 7743
rect 6844 7728 6860 7736
rect 6831 7696 6844 7715
rect 6859 7696 6889 7712
rect 6831 7680 6905 7696
rect 6831 7678 6844 7680
rect 6859 7678 6893 7680
rect 6496 7656 6509 7658
rect 6524 7656 6558 7658
rect 6496 7640 6558 7656
rect 6602 7651 6618 7654
rect 6680 7651 6710 7662
rect 6758 7658 6804 7674
rect 6831 7662 6905 7678
rect 6758 7656 6792 7658
rect 6757 7640 6804 7656
rect 6831 7640 6844 7662
rect 6859 7640 6889 7662
rect 6916 7640 6917 7656
rect 6932 7640 6945 7800
rect 6975 7696 6988 7800
rect 7033 7778 7034 7788
rect 7049 7778 7062 7788
rect 7033 7774 7062 7778
rect 7067 7774 7097 7800
rect 7115 7786 7131 7788
rect 7203 7786 7256 7800
rect 7204 7784 7268 7786
rect 7311 7784 7326 7800
rect 7375 7797 7405 7800
rect 7375 7794 7411 7797
rect 7341 7786 7357 7788
rect 7115 7774 7130 7778
rect 7033 7772 7130 7774
rect 7158 7772 7326 7784
rect 7342 7774 7357 7778
rect 7375 7775 7414 7794
rect 7433 7788 7440 7789
rect 7439 7781 7440 7788
rect 7423 7778 7424 7781
rect 7439 7778 7452 7781
rect 7375 7774 7405 7775
rect 7414 7774 7420 7775
rect 7423 7774 7452 7778
rect 7342 7773 7452 7774
rect 7342 7772 7458 7773
rect 7017 7764 7068 7772
rect 7017 7752 7042 7764
rect 7049 7752 7068 7764
rect 7099 7764 7149 7772
rect 7099 7756 7115 7764
rect 7122 7762 7149 7764
rect 7158 7762 7379 7772
rect 7122 7752 7379 7762
rect 7408 7764 7458 7772
rect 7408 7755 7424 7764
rect 7017 7744 7068 7752
rect 7115 7744 7379 7752
rect 7405 7752 7424 7755
rect 7431 7752 7458 7764
rect 7405 7744 7458 7752
rect 7033 7736 7034 7744
rect 7049 7736 7062 7744
rect 7033 7728 7049 7736
rect 7030 7721 7049 7724
rect 7030 7712 7052 7721
rect 7003 7702 7052 7712
rect 7003 7696 7033 7702
rect 7052 7697 7057 7702
rect 6975 7680 7049 7696
rect 7067 7688 7097 7744
rect 7132 7734 7340 7744
rect 7375 7740 7420 7744
rect 7423 7743 7424 7744
rect 7439 7743 7452 7744
rect 7158 7704 7347 7734
rect 7173 7701 7347 7704
rect 7166 7698 7347 7701
rect 6975 7678 6988 7680
rect 7003 7678 7037 7680
rect 6975 7662 7049 7678
rect 7076 7674 7089 7688
rect 7104 7674 7120 7690
rect 7166 7685 7177 7698
rect 6959 7640 6960 7656
rect 6975 7640 6988 7662
rect 7003 7640 7033 7662
rect 7076 7658 7138 7674
rect 7166 7667 7177 7683
rect 7182 7678 7192 7698
rect 7202 7678 7216 7698
rect 7219 7685 7228 7698
rect 7244 7685 7253 7698
rect 7182 7667 7216 7678
rect 7219 7667 7228 7683
rect 7244 7667 7253 7683
rect 7260 7678 7270 7698
rect 7280 7678 7294 7698
rect 7295 7685 7306 7698
rect 7260 7667 7294 7678
rect 7295 7667 7306 7683
rect 7352 7674 7368 7690
rect 7375 7688 7405 7740
rect 7439 7736 7440 7743
rect 7424 7728 7440 7736
rect 7411 7696 7424 7715
rect 7439 7696 7469 7712
rect 7411 7680 7485 7696
rect 7411 7678 7424 7680
rect 7439 7678 7473 7680
rect 7076 7656 7089 7658
rect 7104 7656 7138 7658
rect 7076 7640 7138 7656
rect 7182 7651 7198 7654
rect 7260 7651 7290 7662
rect 7338 7658 7384 7674
rect 7411 7662 7485 7678
rect 7338 7656 7372 7658
rect 7337 7640 7384 7656
rect 7411 7640 7424 7662
rect 7439 7640 7469 7662
rect 7496 7640 7497 7656
rect 7512 7640 7525 7800
rect 7555 7696 7568 7800
rect 7613 7778 7614 7788
rect 7629 7778 7642 7788
rect 7613 7774 7642 7778
rect 7647 7774 7677 7800
rect 7695 7786 7711 7788
rect 7783 7786 7836 7800
rect 7784 7784 7848 7786
rect 7891 7784 7906 7800
rect 7955 7797 7985 7800
rect 7955 7794 7991 7797
rect 7921 7786 7937 7788
rect 7695 7774 7710 7778
rect 7613 7772 7710 7774
rect 7738 7772 7906 7784
rect 7922 7774 7937 7778
rect 7955 7775 7994 7794
rect 8013 7788 8020 7789
rect 8019 7781 8020 7788
rect 8003 7778 8004 7781
rect 8019 7778 8032 7781
rect 7955 7774 7985 7775
rect 7994 7774 8000 7775
rect 8003 7774 8032 7778
rect 7922 7773 8032 7774
rect 7922 7772 8038 7773
rect 7597 7764 7648 7772
rect 7597 7752 7622 7764
rect 7629 7752 7648 7764
rect 7679 7764 7729 7772
rect 7679 7756 7695 7764
rect 7702 7762 7729 7764
rect 7738 7762 7959 7772
rect 7702 7752 7959 7762
rect 7988 7764 8038 7772
rect 7988 7755 8004 7764
rect 7597 7744 7648 7752
rect 7695 7744 7959 7752
rect 7985 7752 8004 7755
rect 8011 7752 8038 7764
rect 7985 7744 8038 7752
rect 7613 7736 7614 7744
rect 7629 7736 7642 7744
rect 7613 7728 7629 7736
rect 7610 7721 7629 7724
rect 7610 7712 7632 7721
rect 7583 7702 7632 7712
rect 7583 7696 7613 7702
rect 7632 7697 7637 7702
rect 7555 7680 7629 7696
rect 7647 7688 7677 7744
rect 7712 7734 7920 7744
rect 7955 7740 8000 7744
rect 8003 7743 8004 7744
rect 8019 7743 8032 7744
rect 7738 7704 7927 7734
rect 7753 7701 7927 7704
rect 7746 7698 7927 7701
rect 7555 7678 7568 7680
rect 7583 7678 7617 7680
rect 7555 7662 7629 7678
rect 7656 7674 7669 7688
rect 7684 7674 7700 7690
rect 7746 7685 7757 7698
rect 7539 7640 7540 7656
rect 7555 7640 7568 7662
rect 7583 7640 7613 7662
rect 7656 7658 7718 7674
rect 7746 7667 7757 7683
rect 7762 7678 7772 7698
rect 7782 7678 7796 7698
rect 7799 7685 7808 7698
rect 7824 7685 7833 7698
rect 7762 7667 7796 7678
rect 7799 7667 7808 7683
rect 7824 7667 7833 7683
rect 7840 7678 7850 7698
rect 7860 7678 7874 7698
rect 7875 7685 7886 7698
rect 7840 7667 7874 7678
rect 7875 7667 7886 7683
rect 7932 7674 7948 7690
rect 7955 7688 7985 7740
rect 8019 7736 8020 7743
rect 8004 7728 8020 7736
rect 7991 7696 8004 7715
rect 8019 7696 8049 7712
rect 7991 7680 8065 7696
rect 7991 7678 8004 7680
rect 8019 7678 8053 7680
rect 7656 7656 7669 7658
rect 7684 7656 7718 7658
rect 7656 7640 7718 7656
rect 7762 7651 7778 7654
rect 7840 7651 7870 7662
rect 7918 7658 7964 7674
rect 7991 7662 8065 7678
rect 7918 7656 7952 7658
rect 7917 7640 7964 7656
rect 7991 7640 8004 7662
rect 8019 7640 8049 7662
rect 8076 7640 8077 7656
rect 8092 7640 8105 7800
rect 8135 7696 8148 7800
rect 8193 7778 8194 7788
rect 8209 7778 8222 7788
rect 8193 7774 8222 7778
rect 8227 7774 8257 7800
rect 8275 7786 8291 7788
rect 8363 7786 8416 7800
rect 8364 7784 8428 7786
rect 8471 7784 8486 7800
rect 8535 7797 8565 7800
rect 8535 7794 8571 7797
rect 8501 7786 8517 7788
rect 8275 7774 8290 7778
rect 8193 7772 8290 7774
rect 8318 7772 8486 7784
rect 8502 7774 8517 7778
rect 8535 7775 8574 7794
rect 8593 7788 8600 7789
rect 8599 7781 8600 7788
rect 8583 7778 8584 7781
rect 8599 7778 8612 7781
rect 8535 7774 8565 7775
rect 8574 7774 8580 7775
rect 8583 7774 8612 7778
rect 8502 7773 8612 7774
rect 8502 7772 8618 7773
rect 8177 7764 8228 7772
rect 8177 7752 8202 7764
rect 8209 7752 8228 7764
rect 8259 7764 8309 7772
rect 8259 7756 8275 7764
rect 8282 7762 8309 7764
rect 8318 7762 8539 7772
rect 8282 7752 8539 7762
rect 8568 7764 8618 7772
rect 8568 7755 8584 7764
rect 8177 7744 8228 7752
rect 8275 7744 8539 7752
rect 8565 7752 8584 7755
rect 8591 7752 8618 7764
rect 8565 7744 8618 7752
rect 8193 7736 8194 7744
rect 8209 7736 8222 7744
rect 8193 7728 8209 7736
rect 8190 7721 8209 7724
rect 8190 7712 8212 7721
rect 8163 7702 8212 7712
rect 8163 7696 8193 7702
rect 8212 7697 8217 7702
rect 8135 7680 8209 7696
rect 8227 7688 8257 7744
rect 8292 7734 8500 7744
rect 8535 7740 8580 7744
rect 8583 7743 8584 7744
rect 8599 7743 8612 7744
rect 8318 7704 8507 7734
rect 8333 7701 8507 7704
rect 8326 7698 8507 7701
rect 8135 7678 8148 7680
rect 8163 7678 8197 7680
rect 8135 7662 8209 7678
rect 8236 7674 8249 7688
rect 8264 7674 8280 7690
rect 8326 7685 8337 7698
rect 8119 7640 8120 7656
rect 8135 7640 8148 7662
rect 8163 7640 8193 7662
rect 8236 7658 8298 7674
rect 8326 7667 8337 7683
rect 8342 7678 8352 7698
rect 8362 7678 8376 7698
rect 8379 7685 8388 7698
rect 8404 7685 8413 7698
rect 8342 7667 8376 7678
rect 8379 7667 8388 7683
rect 8404 7667 8413 7683
rect 8420 7678 8430 7698
rect 8440 7678 8454 7698
rect 8455 7685 8466 7698
rect 8420 7667 8454 7678
rect 8455 7667 8466 7683
rect 8512 7674 8528 7690
rect 8535 7688 8565 7740
rect 8599 7736 8600 7743
rect 8584 7728 8600 7736
rect 8571 7696 8584 7715
rect 8599 7696 8629 7712
rect 8571 7680 8645 7696
rect 8571 7678 8584 7680
rect 8599 7678 8633 7680
rect 8236 7656 8249 7658
rect 8264 7656 8298 7658
rect 8236 7640 8298 7656
rect 8342 7651 8358 7654
rect 8420 7651 8450 7662
rect 8498 7658 8544 7674
rect 8571 7662 8645 7678
rect 8498 7656 8532 7658
rect 8497 7640 8544 7656
rect 8571 7640 8584 7662
rect 8599 7640 8629 7662
rect 8656 7640 8657 7656
rect 8672 7640 8685 7800
rect 8715 7696 8728 7800
rect 8773 7778 8774 7788
rect 8789 7778 8802 7788
rect 8773 7774 8802 7778
rect 8807 7774 8837 7800
rect 8855 7786 8871 7788
rect 8943 7786 8996 7800
rect 8944 7784 9008 7786
rect 9051 7784 9066 7800
rect 9115 7797 9145 7800
rect 9115 7794 9151 7797
rect 9081 7786 9097 7788
rect 8855 7774 8870 7778
rect 8773 7772 8870 7774
rect 8898 7772 9066 7784
rect 9082 7774 9097 7778
rect 9115 7775 9154 7794
rect 9173 7788 9180 7789
rect 9179 7781 9180 7788
rect 9163 7778 9164 7781
rect 9179 7778 9192 7781
rect 9115 7774 9145 7775
rect 9154 7774 9160 7775
rect 9163 7774 9192 7778
rect 9082 7773 9192 7774
rect 9082 7772 9198 7773
rect 8757 7764 8808 7772
rect 8757 7752 8782 7764
rect 8789 7752 8808 7764
rect 8839 7764 8889 7772
rect 8839 7756 8855 7764
rect 8862 7762 8889 7764
rect 8898 7762 9119 7772
rect 8862 7752 9119 7762
rect 9148 7764 9198 7772
rect 9148 7755 9164 7764
rect 8757 7744 8808 7752
rect 8855 7744 9119 7752
rect 9145 7752 9164 7755
rect 9171 7752 9198 7764
rect 9145 7744 9198 7752
rect 8773 7736 8774 7744
rect 8789 7736 8802 7744
rect 8773 7728 8789 7736
rect 8770 7721 8789 7724
rect 8770 7712 8792 7721
rect 8743 7702 8792 7712
rect 8743 7696 8773 7702
rect 8792 7697 8797 7702
rect 8715 7680 8789 7696
rect 8807 7688 8837 7744
rect 8872 7734 9080 7744
rect 9115 7740 9160 7744
rect 9163 7743 9164 7744
rect 9179 7743 9192 7744
rect 8898 7704 9087 7734
rect 8913 7701 9087 7704
rect 8906 7698 9087 7701
rect 8715 7678 8728 7680
rect 8743 7678 8777 7680
rect 8715 7662 8789 7678
rect 8816 7674 8829 7688
rect 8844 7674 8860 7690
rect 8906 7685 8917 7698
rect 8699 7640 8700 7656
rect 8715 7640 8728 7662
rect 8743 7640 8773 7662
rect 8816 7658 8878 7674
rect 8906 7667 8917 7683
rect 8922 7678 8932 7698
rect 8942 7678 8956 7698
rect 8959 7685 8968 7698
rect 8984 7685 8993 7698
rect 8922 7667 8956 7678
rect 8959 7667 8968 7683
rect 8984 7667 8993 7683
rect 9000 7678 9010 7698
rect 9020 7678 9034 7698
rect 9035 7685 9046 7698
rect 9000 7667 9034 7678
rect 9035 7667 9046 7683
rect 9092 7674 9108 7690
rect 9115 7688 9145 7740
rect 9179 7736 9180 7743
rect 9164 7728 9180 7736
rect 9151 7696 9164 7715
rect 9179 7696 9209 7712
rect 9151 7680 9225 7696
rect 9151 7678 9164 7680
rect 9179 7678 9213 7680
rect 8816 7656 8829 7658
rect 8844 7656 8878 7658
rect 8816 7640 8878 7656
rect 8922 7651 8938 7654
rect 9000 7651 9030 7662
rect 9078 7658 9124 7674
rect 9151 7662 9225 7678
rect 9078 7656 9112 7658
rect 9077 7640 9124 7656
rect 9151 7640 9164 7662
rect 9179 7640 9209 7662
rect 9236 7640 9237 7656
rect 9252 7640 9265 7800
rect -7 7632 34 7640
rect -7 7606 8 7632
rect 15 7606 34 7632
rect 98 7628 160 7640
rect 172 7628 247 7640
rect 305 7628 380 7640
rect 392 7628 423 7640
rect 429 7628 464 7640
rect 98 7626 260 7628
rect -7 7598 34 7606
rect 116 7602 129 7626
rect 144 7624 159 7626
rect -1 7588 0 7598
rect 15 7588 28 7598
rect 43 7588 73 7602
rect 116 7588 159 7602
rect 183 7599 190 7606
rect 193 7602 260 7626
rect 292 7626 464 7628
rect 262 7604 290 7608
rect 292 7604 372 7626
rect 393 7624 408 7626
rect 262 7602 372 7604
rect 193 7598 372 7602
rect 166 7588 196 7598
rect 198 7588 351 7598
rect 359 7588 389 7598
rect 393 7588 423 7602
rect 451 7588 464 7626
rect 536 7632 571 7640
rect 536 7606 537 7632
rect 544 7606 571 7632
rect 479 7588 509 7602
rect 536 7598 571 7606
rect 573 7632 614 7640
rect 573 7606 588 7632
rect 595 7606 614 7632
rect 678 7628 740 7640
rect 752 7628 827 7640
rect 885 7628 960 7640
rect 972 7628 1003 7640
rect 1009 7628 1044 7640
rect 678 7626 840 7628
rect 573 7598 614 7606
rect 696 7602 709 7626
rect 724 7624 739 7626
rect 536 7588 537 7598
rect 552 7588 565 7598
rect 579 7588 580 7598
rect 595 7588 608 7598
rect 623 7588 653 7602
rect 696 7588 739 7602
rect 763 7599 770 7606
rect 773 7602 840 7626
rect 872 7626 1044 7628
rect 842 7604 870 7608
rect 872 7604 952 7626
rect 973 7624 988 7626
rect 842 7602 952 7604
rect 773 7598 952 7602
rect 746 7588 776 7598
rect 778 7588 931 7598
rect 939 7588 969 7598
rect 973 7588 1003 7602
rect 1031 7588 1044 7626
rect 1116 7632 1151 7640
rect 1116 7606 1117 7632
rect 1124 7606 1151 7632
rect 1059 7588 1089 7602
rect 1116 7598 1151 7606
rect 1153 7632 1194 7640
rect 1153 7606 1168 7632
rect 1175 7606 1194 7632
rect 1258 7628 1320 7640
rect 1332 7628 1407 7640
rect 1465 7628 1540 7640
rect 1552 7628 1583 7640
rect 1589 7628 1624 7640
rect 1258 7626 1420 7628
rect 1153 7598 1194 7606
rect 1276 7602 1289 7626
rect 1304 7624 1319 7626
rect 1116 7588 1117 7598
rect 1132 7588 1145 7598
rect 1159 7588 1160 7598
rect 1175 7588 1188 7598
rect 1203 7588 1233 7602
rect 1276 7588 1319 7602
rect 1343 7599 1350 7606
rect 1353 7602 1420 7626
rect 1452 7626 1624 7628
rect 1422 7604 1450 7608
rect 1452 7604 1532 7626
rect 1553 7624 1568 7626
rect 1422 7602 1532 7604
rect 1353 7598 1532 7602
rect 1326 7588 1356 7598
rect 1358 7588 1511 7598
rect 1519 7588 1549 7598
rect 1553 7588 1583 7602
rect 1611 7588 1624 7626
rect 1696 7632 1731 7640
rect 1696 7606 1697 7632
rect 1704 7606 1731 7632
rect 1639 7588 1669 7602
rect 1696 7598 1731 7606
rect 1733 7632 1774 7640
rect 1733 7606 1748 7632
rect 1755 7606 1774 7632
rect 1838 7628 1900 7640
rect 1912 7628 1987 7640
rect 2045 7628 2120 7640
rect 2132 7628 2163 7640
rect 2169 7628 2204 7640
rect 1838 7626 2000 7628
rect 1733 7598 1774 7606
rect 1856 7602 1869 7626
rect 1884 7624 1899 7626
rect 1696 7588 1697 7598
rect 1712 7588 1725 7598
rect 1739 7588 1740 7598
rect 1755 7588 1768 7598
rect 1783 7588 1813 7602
rect 1856 7588 1899 7602
rect 1923 7599 1930 7606
rect 1933 7602 2000 7626
rect 2032 7626 2204 7628
rect 2002 7604 2030 7608
rect 2032 7604 2112 7626
rect 2133 7624 2148 7626
rect 2002 7602 2112 7604
rect 1933 7598 2112 7602
rect 1906 7588 1936 7598
rect 1938 7588 2091 7598
rect 2099 7588 2129 7598
rect 2133 7588 2163 7602
rect 2191 7588 2204 7626
rect 2276 7632 2311 7640
rect 2276 7606 2277 7632
rect 2284 7606 2311 7632
rect 2219 7588 2249 7602
rect 2276 7598 2311 7606
rect 2313 7632 2354 7640
rect 2313 7606 2328 7632
rect 2335 7606 2354 7632
rect 2418 7628 2480 7640
rect 2492 7628 2567 7640
rect 2625 7628 2700 7640
rect 2712 7628 2743 7640
rect 2749 7628 2784 7640
rect 2418 7626 2580 7628
rect 2313 7598 2354 7606
rect 2436 7602 2449 7626
rect 2464 7624 2479 7626
rect 2276 7588 2277 7598
rect 2292 7588 2305 7598
rect 2319 7588 2320 7598
rect 2335 7588 2348 7598
rect 2363 7588 2393 7602
rect 2436 7588 2479 7602
rect 2503 7599 2510 7606
rect 2513 7602 2580 7626
rect 2612 7626 2784 7628
rect 2582 7604 2610 7608
rect 2612 7604 2692 7626
rect 2713 7624 2728 7626
rect 2582 7602 2692 7604
rect 2513 7598 2692 7602
rect 2486 7588 2516 7598
rect 2518 7588 2671 7598
rect 2679 7588 2709 7598
rect 2713 7588 2743 7602
rect 2771 7588 2784 7626
rect 2856 7632 2891 7640
rect 2856 7606 2857 7632
rect 2864 7606 2891 7632
rect 2799 7588 2829 7602
rect 2856 7598 2891 7606
rect 2893 7632 2934 7640
rect 2893 7606 2908 7632
rect 2915 7606 2934 7632
rect 2998 7628 3060 7640
rect 3072 7628 3147 7640
rect 3205 7628 3280 7640
rect 3292 7628 3323 7640
rect 3329 7628 3364 7640
rect 2998 7626 3160 7628
rect 2893 7598 2934 7606
rect 3016 7602 3029 7626
rect 3044 7624 3059 7626
rect 2856 7588 2857 7598
rect 2872 7588 2885 7598
rect 2899 7588 2900 7598
rect 2915 7588 2928 7598
rect 2943 7588 2973 7602
rect 3016 7588 3059 7602
rect 3083 7599 3090 7606
rect 3093 7602 3160 7626
rect 3192 7626 3364 7628
rect 3162 7604 3190 7608
rect 3192 7604 3272 7626
rect 3293 7624 3308 7626
rect 3162 7602 3272 7604
rect 3093 7598 3272 7602
rect 3066 7588 3096 7598
rect 3098 7588 3251 7598
rect 3259 7588 3289 7598
rect 3293 7588 3323 7602
rect 3351 7588 3364 7626
rect 3436 7632 3471 7640
rect 3436 7606 3437 7632
rect 3444 7606 3471 7632
rect 3379 7588 3409 7602
rect 3436 7598 3471 7606
rect 3473 7632 3514 7640
rect 3473 7606 3488 7632
rect 3495 7606 3514 7632
rect 3578 7628 3640 7640
rect 3652 7628 3727 7640
rect 3785 7628 3860 7640
rect 3872 7628 3903 7640
rect 3909 7628 3944 7640
rect 3578 7626 3740 7628
rect 3473 7598 3514 7606
rect 3596 7602 3609 7626
rect 3624 7624 3639 7626
rect 3436 7588 3437 7598
rect 3452 7588 3465 7598
rect 3479 7588 3480 7598
rect 3495 7588 3508 7598
rect 3523 7588 3553 7602
rect 3596 7588 3639 7602
rect 3663 7599 3670 7606
rect 3673 7602 3740 7626
rect 3772 7626 3944 7628
rect 3742 7604 3770 7608
rect 3772 7604 3852 7626
rect 3873 7624 3888 7626
rect 3742 7602 3852 7604
rect 3673 7598 3852 7602
rect 3646 7588 3676 7598
rect 3678 7588 3831 7598
rect 3839 7588 3869 7598
rect 3873 7588 3903 7602
rect 3931 7588 3944 7626
rect 4016 7632 4051 7640
rect 4016 7606 4017 7632
rect 4024 7606 4051 7632
rect 3959 7588 3989 7602
rect 4016 7598 4051 7606
rect 4053 7632 4094 7640
rect 4053 7606 4068 7632
rect 4075 7606 4094 7632
rect 4158 7628 4220 7640
rect 4232 7628 4307 7640
rect 4365 7628 4440 7640
rect 4452 7628 4483 7640
rect 4489 7628 4524 7640
rect 4158 7626 4320 7628
rect 4053 7598 4094 7606
rect 4176 7602 4189 7626
rect 4204 7624 4219 7626
rect 4016 7588 4017 7598
rect 4032 7588 4045 7598
rect 4059 7588 4060 7598
rect 4075 7588 4088 7598
rect 4103 7588 4133 7602
rect 4176 7588 4219 7602
rect 4243 7599 4250 7606
rect 4253 7602 4320 7626
rect 4352 7626 4524 7628
rect 4322 7604 4350 7608
rect 4352 7604 4432 7626
rect 4453 7624 4468 7626
rect 4322 7602 4432 7604
rect 4253 7598 4432 7602
rect 4226 7588 4256 7598
rect 4258 7588 4411 7598
rect 4419 7588 4449 7598
rect 4453 7588 4483 7602
rect 4511 7588 4524 7626
rect 4596 7632 4631 7640
rect 4596 7606 4597 7632
rect 4604 7606 4631 7632
rect 4539 7588 4569 7602
rect 4596 7598 4631 7606
rect 4633 7632 4674 7640
rect 4633 7606 4648 7632
rect 4655 7606 4674 7632
rect 4738 7628 4800 7640
rect 4812 7628 4887 7640
rect 4945 7628 5020 7640
rect 5032 7628 5063 7640
rect 5069 7628 5104 7640
rect 4738 7626 4900 7628
rect 4633 7598 4674 7606
rect 4756 7602 4769 7626
rect 4784 7624 4799 7626
rect 4596 7588 4597 7598
rect 4612 7588 4625 7598
rect 4639 7588 4640 7598
rect 4655 7588 4668 7598
rect 4683 7588 4713 7602
rect 4756 7588 4799 7602
rect 4823 7599 4830 7606
rect 4833 7602 4900 7626
rect 4932 7626 5104 7628
rect 4902 7604 4930 7608
rect 4932 7604 5012 7626
rect 5033 7624 5048 7626
rect 4902 7602 5012 7604
rect 4833 7598 5012 7602
rect 4806 7588 4836 7598
rect 4838 7588 4991 7598
rect 4999 7588 5029 7598
rect 5033 7588 5063 7602
rect 5091 7588 5104 7626
rect 5176 7632 5211 7640
rect 5176 7606 5177 7632
rect 5184 7606 5211 7632
rect 5119 7588 5149 7602
rect 5176 7598 5211 7606
rect 5213 7632 5254 7640
rect 5213 7606 5228 7632
rect 5235 7606 5254 7632
rect 5318 7628 5380 7640
rect 5392 7628 5467 7640
rect 5525 7628 5600 7640
rect 5612 7628 5643 7640
rect 5649 7628 5684 7640
rect 5318 7626 5480 7628
rect 5213 7598 5254 7606
rect 5336 7602 5349 7626
rect 5364 7624 5379 7626
rect 5176 7588 5177 7598
rect 5192 7588 5205 7598
rect 5219 7588 5220 7598
rect 5235 7588 5248 7598
rect 5263 7588 5293 7602
rect 5336 7588 5379 7602
rect 5403 7599 5410 7606
rect 5413 7602 5480 7626
rect 5512 7626 5684 7628
rect 5482 7604 5510 7608
rect 5512 7604 5592 7626
rect 5613 7624 5628 7626
rect 5482 7602 5592 7604
rect 5413 7598 5592 7602
rect 5386 7588 5416 7598
rect 5418 7588 5571 7598
rect 5579 7588 5609 7598
rect 5613 7588 5643 7602
rect 5671 7588 5684 7626
rect 5756 7632 5791 7640
rect 5756 7606 5757 7632
rect 5764 7606 5791 7632
rect 5699 7588 5729 7602
rect 5756 7598 5791 7606
rect 5793 7632 5834 7640
rect 5793 7606 5808 7632
rect 5815 7606 5834 7632
rect 5898 7628 5960 7640
rect 5972 7628 6047 7640
rect 6105 7628 6180 7640
rect 6192 7628 6223 7640
rect 6229 7628 6264 7640
rect 5898 7626 6060 7628
rect 5793 7598 5834 7606
rect 5916 7602 5929 7626
rect 5944 7624 5959 7626
rect 5756 7588 5757 7598
rect 5772 7588 5785 7598
rect 5799 7588 5800 7598
rect 5815 7588 5828 7598
rect 5843 7588 5873 7602
rect 5916 7588 5959 7602
rect 5983 7599 5990 7606
rect 5993 7602 6060 7626
rect 6092 7626 6264 7628
rect 6062 7604 6090 7608
rect 6092 7604 6172 7626
rect 6193 7624 6208 7626
rect 6062 7602 6172 7604
rect 5993 7598 6172 7602
rect 5966 7588 5996 7598
rect 5998 7588 6151 7598
rect 6159 7588 6189 7598
rect 6193 7588 6223 7602
rect 6251 7588 6264 7626
rect 6336 7632 6371 7640
rect 6336 7606 6337 7632
rect 6344 7606 6371 7632
rect 6279 7588 6309 7602
rect 6336 7598 6371 7606
rect 6373 7632 6414 7640
rect 6373 7606 6388 7632
rect 6395 7606 6414 7632
rect 6478 7628 6540 7640
rect 6552 7628 6627 7640
rect 6685 7628 6760 7640
rect 6772 7628 6803 7640
rect 6809 7628 6844 7640
rect 6478 7626 6640 7628
rect 6373 7598 6414 7606
rect 6496 7602 6509 7626
rect 6524 7624 6539 7626
rect 6336 7588 6337 7598
rect 6352 7588 6365 7598
rect 6379 7588 6380 7598
rect 6395 7588 6408 7598
rect 6423 7588 6453 7602
rect 6496 7588 6539 7602
rect 6563 7599 6570 7606
rect 6573 7602 6640 7626
rect 6672 7626 6844 7628
rect 6642 7604 6670 7608
rect 6672 7604 6752 7626
rect 6773 7624 6788 7626
rect 6642 7602 6752 7604
rect 6573 7598 6752 7602
rect 6546 7588 6576 7598
rect 6578 7588 6731 7598
rect 6739 7588 6769 7598
rect 6773 7588 6803 7602
rect 6831 7588 6844 7626
rect 6916 7632 6951 7640
rect 6916 7606 6917 7632
rect 6924 7606 6951 7632
rect 6859 7588 6889 7602
rect 6916 7598 6951 7606
rect 6953 7632 6994 7640
rect 6953 7606 6968 7632
rect 6975 7606 6994 7632
rect 7058 7628 7120 7640
rect 7132 7628 7207 7640
rect 7265 7628 7340 7640
rect 7352 7628 7383 7640
rect 7389 7628 7424 7640
rect 7058 7626 7220 7628
rect 6953 7598 6994 7606
rect 7076 7602 7089 7626
rect 7104 7624 7119 7626
rect 6916 7588 6917 7598
rect 6932 7588 6945 7598
rect 6959 7588 6960 7598
rect 6975 7588 6988 7598
rect 7003 7588 7033 7602
rect 7076 7588 7119 7602
rect 7143 7599 7150 7606
rect 7153 7602 7220 7626
rect 7252 7626 7424 7628
rect 7222 7604 7250 7608
rect 7252 7604 7332 7626
rect 7353 7624 7368 7626
rect 7222 7602 7332 7604
rect 7153 7598 7332 7602
rect 7126 7588 7156 7598
rect 7158 7588 7311 7598
rect 7319 7588 7349 7598
rect 7353 7588 7383 7602
rect 7411 7588 7424 7626
rect 7496 7632 7531 7640
rect 7496 7606 7497 7632
rect 7504 7606 7531 7632
rect 7439 7588 7469 7602
rect 7496 7598 7531 7606
rect 7533 7632 7574 7640
rect 7533 7606 7548 7632
rect 7555 7606 7574 7632
rect 7638 7628 7700 7640
rect 7712 7628 7787 7640
rect 7845 7628 7920 7640
rect 7932 7628 7963 7640
rect 7969 7628 8004 7640
rect 7638 7626 7800 7628
rect 7533 7598 7574 7606
rect 7656 7602 7669 7626
rect 7684 7624 7699 7626
rect 7496 7588 7497 7598
rect 7512 7588 7525 7598
rect 7539 7588 7540 7598
rect 7555 7588 7568 7598
rect 7583 7588 7613 7602
rect 7656 7588 7699 7602
rect 7723 7599 7730 7606
rect 7733 7602 7800 7626
rect 7832 7626 8004 7628
rect 7802 7604 7830 7608
rect 7832 7604 7912 7626
rect 7933 7624 7948 7626
rect 7802 7602 7912 7604
rect 7733 7598 7912 7602
rect 7706 7588 7736 7598
rect 7738 7588 7891 7598
rect 7899 7588 7929 7598
rect 7933 7588 7963 7602
rect 7991 7588 8004 7626
rect 8076 7632 8111 7640
rect 8076 7606 8077 7632
rect 8084 7606 8111 7632
rect 8019 7588 8049 7602
rect 8076 7598 8111 7606
rect 8113 7632 8154 7640
rect 8113 7606 8128 7632
rect 8135 7606 8154 7632
rect 8218 7628 8280 7640
rect 8292 7628 8367 7640
rect 8425 7628 8500 7640
rect 8512 7628 8543 7640
rect 8549 7628 8584 7640
rect 8218 7626 8380 7628
rect 8113 7598 8154 7606
rect 8236 7602 8249 7626
rect 8264 7624 8279 7626
rect 8076 7588 8077 7598
rect 8092 7588 8105 7598
rect 8119 7588 8120 7598
rect 8135 7588 8148 7598
rect 8163 7588 8193 7602
rect 8236 7588 8279 7602
rect 8303 7599 8310 7606
rect 8313 7602 8380 7626
rect 8412 7626 8584 7628
rect 8382 7604 8410 7608
rect 8412 7604 8492 7626
rect 8513 7624 8528 7626
rect 8382 7602 8492 7604
rect 8313 7598 8492 7602
rect 8286 7588 8316 7598
rect 8318 7588 8471 7598
rect 8479 7588 8509 7598
rect 8513 7588 8543 7602
rect 8571 7588 8584 7626
rect 8656 7632 8691 7640
rect 8656 7606 8657 7632
rect 8664 7606 8691 7632
rect 8599 7588 8629 7602
rect 8656 7598 8691 7606
rect 8693 7632 8734 7640
rect 8693 7606 8708 7632
rect 8715 7606 8734 7632
rect 8798 7628 8860 7640
rect 8872 7628 8947 7640
rect 9005 7628 9080 7640
rect 9092 7628 9123 7640
rect 9129 7628 9164 7640
rect 8798 7626 8960 7628
rect 8693 7598 8734 7606
rect 8816 7602 8829 7626
rect 8844 7624 8859 7626
rect 8656 7588 8657 7598
rect 8672 7588 8685 7598
rect 8699 7588 8700 7598
rect 8715 7588 8728 7598
rect 8743 7588 8773 7602
rect 8816 7588 8859 7602
rect 8883 7599 8890 7606
rect 8893 7602 8960 7626
rect 8992 7626 9164 7628
rect 8962 7604 8990 7608
rect 8992 7604 9072 7626
rect 9093 7624 9108 7626
rect 8962 7602 9072 7604
rect 8893 7598 9072 7602
rect 8866 7588 8896 7598
rect 8898 7588 9051 7598
rect 9059 7588 9089 7598
rect 9093 7588 9123 7602
rect 9151 7588 9164 7626
rect 9236 7632 9271 7640
rect 9236 7606 9237 7632
rect 9244 7606 9271 7632
rect 9179 7588 9209 7602
rect 9236 7598 9271 7606
rect 9236 7588 9237 7598
rect 9252 7588 9265 7598
rect -1 7582 9265 7588
rect 0 7574 9265 7582
rect 15 7544 28 7574
rect 43 7556 73 7574
rect 116 7560 130 7574
rect 166 7560 386 7574
rect 117 7558 130 7560
rect 83 7546 98 7558
rect 80 7544 102 7546
rect 107 7544 137 7558
rect 198 7556 351 7560
rect 180 7544 372 7556
rect 415 7544 445 7558
rect 451 7544 464 7574
rect 479 7556 509 7574
rect 552 7544 565 7574
rect 595 7544 608 7574
rect 623 7556 653 7574
rect 696 7560 710 7574
rect 746 7560 966 7574
rect 697 7558 710 7560
rect 663 7546 678 7558
rect 660 7544 682 7546
rect 687 7544 717 7558
rect 778 7556 931 7560
rect 760 7544 952 7556
rect 995 7544 1025 7558
rect 1031 7544 1044 7574
rect 1059 7556 1089 7574
rect 1132 7544 1145 7574
rect 1175 7544 1188 7574
rect 1203 7556 1233 7574
rect 1276 7560 1290 7574
rect 1326 7560 1546 7574
rect 1277 7558 1290 7560
rect 1243 7546 1258 7558
rect 1240 7544 1262 7546
rect 1267 7544 1297 7558
rect 1358 7556 1511 7560
rect 1340 7544 1532 7556
rect 1575 7544 1605 7558
rect 1611 7544 1624 7574
rect 1639 7556 1669 7574
rect 1712 7544 1725 7574
rect 1755 7544 1768 7574
rect 1783 7556 1813 7574
rect 1856 7560 1870 7574
rect 1906 7560 2126 7574
rect 1857 7558 1870 7560
rect 1823 7546 1838 7558
rect 1820 7544 1842 7546
rect 1847 7544 1877 7558
rect 1938 7556 2091 7560
rect 1920 7544 2112 7556
rect 2155 7544 2185 7558
rect 2191 7544 2204 7574
rect 2219 7556 2249 7574
rect 2292 7544 2305 7574
rect 2335 7544 2348 7574
rect 2363 7556 2393 7574
rect 2436 7560 2450 7574
rect 2486 7560 2706 7574
rect 2437 7558 2450 7560
rect 2403 7546 2418 7558
rect 2400 7544 2422 7546
rect 2427 7544 2457 7558
rect 2518 7556 2671 7560
rect 2500 7544 2692 7556
rect 2735 7544 2765 7558
rect 2771 7544 2784 7574
rect 2799 7556 2829 7574
rect 2872 7544 2885 7574
rect 2915 7544 2928 7574
rect 2943 7556 2973 7574
rect 3016 7560 3030 7574
rect 3066 7560 3286 7574
rect 3017 7558 3030 7560
rect 2983 7546 2998 7558
rect 2980 7544 3002 7546
rect 3007 7544 3037 7558
rect 3098 7556 3251 7560
rect 3080 7544 3272 7556
rect 3315 7544 3345 7558
rect 3351 7544 3364 7574
rect 3379 7556 3409 7574
rect 3452 7544 3465 7574
rect 3495 7544 3508 7574
rect 3523 7556 3553 7574
rect 3596 7560 3610 7574
rect 3646 7560 3866 7574
rect 3597 7558 3610 7560
rect 3563 7546 3578 7558
rect 3560 7544 3582 7546
rect 3587 7544 3617 7558
rect 3678 7556 3831 7560
rect 3660 7544 3852 7556
rect 3895 7544 3925 7558
rect 3931 7544 3944 7574
rect 3959 7556 3989 7574
rect 4032 7544 4045 7574
rect 4075 7544 4088 7574
rect 4103 7556 4133 7574
rect 4176 7560 4190 7574
rect 4226 7560 4446 7574
rect 4177 7558 4190 7560
rect 4143 7546 4158 7558
rect 4140 7544 4162 7546
rect 4167 7544 4197 7558
rect 4258 7556 4411 7560
rect 4240 7544 4432 7556
rect 4475 7544 4505 7558
rect 4511 7544 4524 7574
rect 4539 7556 4569 7574
rect 4612 7544 4625 7574
rect 4655 7544 4668 7574
rect 4683 7556 4713 7574
rect 4756 7560 4770 7574
rect 4806 7560 5026 7574
rect 4757 7558 4770 7560
rect 4723 7546 4738 7558
rect 4720 7544 4742 7546
rect 4747 7544 4777 7558
rect 4838 7556 4991 7560
rect 4820 7544 5012 7556
rect 5055 7544 5085 7558
rect 5091 7544 5104 7574
rect 5119 7556 5149 7574
rect 5192 7544 5205 7574
rect 5235 7544 5248 7574
rect 5263 7556 5293 7574
rect 5336 7560 5350 7574
rect 5386 7560 5606 7574
rect 5337 7558 5350 7560
rect 5303 7546 5318 7558
rect 5300 7544 5322 7546
rect 5327 7544 5357 7558
rect 5418 7556 5571 7560
rect 5400 7544 5592 7556
rect 5635 7544 5665 7558
rect 5671 7544 5684 7574
rect 5699 7556 5729 7574
rect 5772 7544 5785 7574
rect 5815 7544 5828 7574
rect 5843 7556 5873 7574
rect 5916 7560 5930 7574
rect 5966 7560 6186 7574
rect 5917 7558 5930 7560
rect 5883 7546 5898 7558
rect 5880 7544 5902 7546
rect 5907 7544 5937 7558
rect 5998 7556 6151 7560
rect 5980 7544 6172 7556
rect 6215 7544 6245 7558
rect 6251 7544 6264 7574
rect 6279 7556 6309 7574
rect 6352 7544 6365 7574
rect 6395 7544 6408 7574
rect 6423 7556 6453 7574
rect 6496 7560 6510 7574
rect 6546 7560 6766 7574
rect 6497 7558 6510 7560
rect 6463 7546 6478 7558
rect 6460 7544 6482 7546
rect 6487 7544 6517 7558
rect 6578 7556 6731 7560
rect 6560 7544 6752 7556
rect 6795 7544 6825 7558
rect 6831 7544 6844 7574
rect 6859 7556 6889 7574
rect 6932 7544 6945 7574
rect 6975 7544 6988 7574
rect 7003 7556 7033 7574
rect 7076 7560 7090 7574
rect 7126 7560 7346 7574
rect 7077 7558 7090 7560
rect 7043 7546 7058 7558
rect 7040 7544 7062 7546
rect 7067 7544 7097 7558
rect 7158 7556 7311 7560
rect 7140 7544 7332 7556
rect 7375 7544 7405 7558
rect 7411 7544 7424 7574
rect 7439 7556 7469 7574
rect 7512 7544 7525 7574
rect 7555 7544 7568 7574
rect 7583 7556 7613 7574
rect 7656 7560 7670 7574
rect 7706 7560 7926 7574
rect 7657 7558 7670 7560
rect 7623 7546 7638 7558
rect 7620 7544 7642 7546
rect 7647 7544 7677 7558
rect 7738 7556 7891 7560
rect 7720 7544 7912 7556
rect 7955 7544 7985 7558
rect 7991 7544 8004 7574
rect 8019 7556 8049 7574
rect 8092 7544 8105 7574
rect 8135 7544 8148 7574
rect 8163 7556 8193 7574
rect 8236 7560 8250 7574
rect 8286 7560 8506 7574
rect 8237 7558 8250 7560
rect 8203 7546 8218 7558
rect 8200 7544 8222 7546
rect 8227 7544 8257 7558
rect 8318 7556 8471 7560
rect 8300 7544 8492 7556
rect 8535 7544 8565 7558
rect 8571 7544 8584 7574
rect 8599 7556 8629 7574
rect 8672 7544 8685 7574
rect 8715 7544 8728 7574
rect 8743 7556 8773 7574
rect 8816 7560 8830 7574
rect 8866 7560 9086 7574
rect 8817 7558 8830 7560
rect 8783 7546 8798 7558
rect 8780 7544 8802 7546
rect 8807 7544 8837 7558
rect 8898 7556 9051 7560
rect 8880 7544 9072 7556
rect 9115 7544 9145 7558
rect 9151 7544 9164 7574
rect 9179 7556 9209 7574
rect 9252 7544 9265 7574
rect 0 7530 9265 7544
rect 15 7426 28 7530
rect 73 7508 74 7518
rect 89 7508 102 7518
rect 73 7504 102 7508
rect 107 7504 137 7530
rect 155 7516 171 7518
rect 243 7516 296 7530
rect 244 7514 308 7516
rect 351 7514 366 7530
rect 415 7527 445 7530
rect 415 7524 451 7527
rect 381 7516 397 7518
rect 155 7504 170 7508
rect 73 7502 170 7504
rect 198 7502 366 7514
rect 382 7504 397 7508
rect 415 7505 454 7524
rect 473 7518 480 7519
rect 479 7511 480 7518
rect 463 7508 464 7511
rect 479 7508 492 7511
rect 415 7504 445 7505
rect 454 7504 460 7505
rect 463 7504 492 7508
rect 382 7503 492 7504
rect 382 7502 498 7503
rect 57 7494 108 7502
rect 57 7482 82 7494
rect 89 7482 108 7494
rect 139 7494 189 7502
rect 139 7486 155 7494
rect 162 7492 189 7494
rect 198 7492 419 7502
rect 162 7482 419 7492
rect 448 7494 498 7502
rect 448 7485 464 7494
rect 57 7474 108 7482
rect 155 7474 419 7482
rect 445 7482 464 7485
rect 471 7482 498 7494
rect 445 7474 498 7482
rect 73 7466 74 7474
rect 89 7466 102 7474
rect 73 7458 89 7466
rect 70 7451 89 7454
rect 70 7442 92 7451
rect 43 7432 92 7442
rect 43 7426 73 7432
rect 92 7427 97 7432
rect 15 7410 89 7426
rect 107 7418 137 7474
rect 172 7464 380 7474
rect 415 7470 460 7474
rect 463 7473 464 7474
rect 479 7473 492 7474
rect 198 7434 387 7464
rect 213 7431 387 7434
rect 206 7428 387 7431
rect 15 7408 28 7410
rect 43 7408 77 7410
rect 15 7392 89 7408
rect 116 7404 129 7418
rect 144 7404 160 7420
rect 206 7415 217 7428
rect -1 7370 0 7386
rect 15 7370 28 7392
rect 43 7370 73 7392
rect 116 7388 178 7404
rect 206 7397 217 7413
rect 222 7408 232 7428
rect 242 7408 256 7428
rect 259 7415 268 7428
rect 284 7415 293 7428
rect 222 7397 256 7408
rect 259 7397 268 7413
rect 284 7397 293 7413
rect 300 7408 310 7428
rect 320 7408 334 7428
rect 335 7415 346 7428
rect 300 7397 334 7408
rect 335 7397 346 7413
rect 392 7404 408 7420
rect 415 7418 445 7470
rect 479 7466 480 7473
rect 464 7458 480 7466
rect 451 7426 464 7445
rect 479 7426 509 7442
rect 451 7410 525 7426
rect 451 7408 464 7410
rect 479 7408 513 7410
rect 116 7386 129 7388
rect 144 7386 178 7388
rect 116 7370 178 7386
rect 222 7381 238 7384
rect 300 7381 330 7392
rect 378 7388 424 7404
rect 451 7392 525 7408
rect 378 7386 412 7388
rect 377 7370 424 7386
rect 451 7370 464 7392
rect 479 7370 509 7392
rect 536 7370 537 7386
rect 552 7370 565 7530
rect 595 7426 608 7530
rect 653 7508 654 7518
rect 669 7508 682 7518
rect 653 7504 682 7508
rect 687 7504 717 7530
rect 735 7516 751 7518
rect 823 7516 876 7530
rect 824 7514 888 7516
rect 931 7514 946 7530
rect 995 7527 1025 7530
rect 995 7524 1031 7527
rect 961 7516 977 7518
rect 735 7504 750 7508
rect 653 7502 750 7504
rect 778 7502 946 7514
rect 962 7504 977 7508
rect 995 7505 1034 7524
rect 1053 7518 1060 7519
rect 1059 7511 1060 7518
rect 1043 7508 1044 7511
rect 1059 7508 1072 7511
rect 995 7504 1025 7505
rect 1034 7504 1040 7505
rect 1043 7504 1072 7508
rect 962 7503 1072 7504
rect 962 7502 1078 7503
rect 637 7494 688 7502
rect 637 7482 662 7494
rect 669 7482 688 7494
rect 719 7494 769 7502
rect 719 7486 735 7494
rect 742 7492 769 7494
rect 778 7492 999 7502
rect 742 7482 999 7492
rect 1028 7494 1078 7502
rect 1028 7485 1044 7494
rect 637 7474 688 7482
rect 735 7474 999 7482
rect 1025 7482 1044 7485
rect 1051 7482 1078 7494
rect 1025 7474 1078 7482
rect 653 7466 654 7474
rect 669 7466 682 7474
rect 653 7458 669 7466
rect 650 7451 669 7454
rect 650 7442 672 7451
rect 623 7432 672 7442
rect 623 7426 653 7432
rect 672 7427 677 7432
rect 595 7410 669 7426
rect 687 7418 717 7474
rect 752 7464 960 7474
rect 995 7470 1040 7474
rect 1043 7473 1044 7474
rect 1059 7473 1072 7474
rect 778 7434 967 7464
rect 793 7431 967 7434
rect 786 7428 967 7431
rect 595 7408 608 7410
rect 623 7408 657 7410
rect 595 7392 669 7408
rect 696 7404 709 7418
rect 724 7404 740 7420
rect 786 7415 797 7428
rect 579 7370 580 7386
rect 595 7370 608 7392
rect 623 7370 653 7392
rect 696 7388 758 7404
rect 786 7397 797 7413
rect 802 7408 812 7428
rect 822 7408 836 7428
rect 839 7415 848 7428
rect 864 7415 873 7428
rect 802 7397 836 7408
rect 839 7397 848 7413
rect 864 7397 873 7413
rect 880 7408 890 7428
rect 900 7408 914 7428
rect 915 7415 926 7428
rect 880 7397 914 7408
rect 915 7397 926 7413
rect 972 7404 988 7420
rect 995 7418 1025 7470
rect 1059 7466 1060 7473
rect 1044 7458 1060 7466
rect 1031 7426 1044 7445
rect 1059 7426 1089 7442
rect 1031 7410 1105 7426
rect 1031 7408 1044 7410
rect 1059 7408 1093 7410
rect 696 7386 709 7388
rect 724 7386 758 7388
rect 696 7370 758 7386
rect 802 7381 818 7384
rect 880 7381 910 7392
rect 958 7388 1004 7404
rect 1031 7392 1105 7408
rect 958 7386 992 7388
rect 957 7370 1004 7386
rect 1031 7370 1044 7392
rect 1059 7370 1089 7392
rect 1116 7370 1117 7386
rect 1132 7370 1145 7530
rect 1175 7426 1188 7530
rect 1233 7508 1234 7518
rect 1249 7508 1262 7518
rect 1233 7504 1262 7508
rect 1267 7504 1297 7530
rect 1315 7516 1331 7518
rect 1403 7516 1456 7530
rect 1404 7514 1468 7516
rect 1511 7514 1526 7530
rect 1575 7527 1605 7530
rect 1575 7524 1611 7527
rect 1541 7516 1557 7518
rect 1315 7504 1330 7508
rect 1233 7502 1330 7504
rect 1358 7502 1526 7514
rect 1542 7504 1557 7508
rect 1575 7505 1614 7524
rect 1633 7518 1640 7519
rect 1639 7511 1640 7518
rect 1623 7508 1624 7511
rect 1639 7508 1652 7511
rect 1575 7504 1605 7505
rect 1614 7504 1620 7505
rect 1623 7504 1652 7508
rect 1542 7503 1652 7504
rect 1542 7502 1658 7503
rect 1217 7494 1268 7502
rect 1217 7482 1242 7494
rect 1249 7482 1268 7494
rect 1299 7494 1349 7502
rect 1299 7486 1315 7494
rect 1322 7492 1349 7494
rect 1358 7492 1579 7502
rect 1322 7482 1579 7492
rect 1608 7494 1658 7502
rect 1608 7485 1624 7494
rect 1217 7474 1268 7482
rect 1315 7474 1579 7482
rect 1605 7482 1624 7485
rect 1631 7482 1658 7494
rect 1605 7474 1658 7482
rect 1233 7466 1234 7474
rect 1249 7466 1262 7474
rect 1233 7458 1249 7466
rect 1230 7451 1249 7454
rect 1230 7442 1252 7451
rect 1203 7432 1252 7442
rect 1203 7426 1233 7432
rect 1252 7427 1257 7432
rect 1175 7410 1249 7426
rect 1267 7418 1297 7474
rect 1332 7464 1540 7474
rect 1575 7470 1620 7474
rect 1623 7473 1624 7474
rect 1639 7473 1652 7474
rect 1358 7434 1547 7464
rect 1373 7431 1547 7434
rect 1366 7428 1547 7431
rect 1175 7408 1188 7410
rect 1203 7408 1237 7410
rect 1175 7392 1249 7408
rect 1276 7404 1289 7418
rect 1304 7404 1320 7420
rect 1366 7415 1377 7428
rect 1159 7370 1160 7386
rect 1175 7370 1188 7392
rect 1203 7370 1233 7392
rect 1276 7388 1338 7404
rect 1366 7397 1377 7413
rect 1382 7408 1392 7428
rect 1402 7408 1416 7428
rect 1419 7415 1428 7428
rect 1444 7415 1453 7428
rect 1382 7397 1416 7408
rect 1419 7397 1428 7413
rect 1444 7397 1453 7413
rect 1460 7408 1470 7428
rect 1480 7408 1494 7428
rect 1495 7415 1506 7428
rect 1460 7397 1494 7408
rect 1495 7397 1506 7413
rect 1552 7404 1568 7420
rect 1575 7418 1605 7470
rect 1639 7466 1640 7473
rect 1624 7458 1640 7466
rect 1611 7426 1624 7445
rect 1639 7426 1669 7442
rect 1611 7410 1685 7426
rect 1611 7408 1624 7410
rect 1639 7408 1673 7410
rect 1276 7386 1289 7388
rect 1304 7386 1338 7388
rect 1276 7370 1338 7386
rect 1382 7381 1398 7384
rect 1460 7381 1490 7392
rect 1538 7388 1584 7404
rect 1611 7392 1685 7408
rect 1538 7386 1572 7388
rect 1537 7370 1584 7386
rect 1611 7370 1624 7392
rect 1639 7370 1669 7392
rect 1696 7370 1697 7386
rect 1712 7370 1725 7530
rect 1755 7426 1768 7530
rect 1813 7508 1814 7518
rect 1829 7508 1842 7518
rect 1813 7504 1842 7508
rect 1847 7504 1877 7530
rect 1895 7516 1911 7518
rect 1983 7516 2036 7530
rect 1984 7514 2048 7516
rect 2091 7514 2106 7530
rect 2155 7527 2185 7530
rect 2155 7524 2191 7527
rect 2121 7516 2137 7518
rect 1895 7504 1910 7508
rect 1813 7502 1910 7504
rect 1938 7502 2106 7514
rect 2122 7504 2137 7508
rect 2155 7505 2194 7524
rect 2213 7518 2220 7519
rect 2219 7511 2220 7518
rect 2203 7508 2204 7511
rect 2219 7508 2232 7511
rect 2155 7504 2185 7505
rect 2194 7504 2200 7505
rect 2203 7504 2232 7508
rect 2122 7503 2232 7504
rect 2122 7502 2238 7503
rect 1797 7494 1848 7502
rect 1797 7482 1822 7494
rect 1829 7482 1848 7494
rect 1879 7494 1929 7502
rect 1879 7486 1895 7494
rect 1902 7492 1929 7494
rect 1938 7492 2159 7502
rect 1902 7482 2159 7492
rect 2188 7494 2238 7502
rect 2188 7485 2204 7494
rect 1797 7474 1848 7482
rect 1895 7474 2159 7482
rect 2185 7482 2204 7485
rect 2211 7482 2238 7494
rect 2185 7474 2238 7482
rect 1813 7466 1814 7474
rect 1829 7466 1842 7474
rect 1813 7458 1829 7466
rect 1810 7451 1829 7454
rect 1810 7442 1832 7451
rect 1783 7432 1832 7442
rect 1783 7426 1813 7432
rect 1832 7427 1837 7432
rect 1755 7410 1829 7426
rect 1847 7418 1877 7474
rect 1912 7464 2120 7474
rect 2155 7470 2200 7474
rect 2203 7473 2204 7474
rect 2219 7473 2232 7474
rect 1938 7434 2127 7464
rect 1953 7431 2127 7434
rect 1946 7428 2127 7431
rect 1755 7408 1768 7410
rect 1783 7408 1817 7410
rect 1755 7392 1829 7408
rect 1856 7404 1869 7418
rect 1884 7404 1900 7420
rect 1946 7415 1957 7428
rect 1739 7370 1740 7386
rect 1755 7370 1768 7392
rect 1783 7370 1813 7392
rect 1856 7388 1918 7404
rect 1946 7397 1957 7413
rect 1962 7408 1972 7428
rect 1982 7408 1996 7428
rect 1999 7415 2008 7428
rect 2024 7415 2033 7428
rect 1962 7397 1996 7408
rect 1999 7397 2008 7413
rect 2024 7397 2033 7413
rect 2040 7408 2050 7428
rect 2060 7408 2074 7428
rect 2075 7415 2086 7428
rect 2040 7397 2074 7408
rect 2075 7397 2086 7413
rect 2132 7404 2148 7420
rect 2155 7418 2185 7470
rect 2219 7466 2220 7473
rect 2204 7458 2220 7466
rect 2191 7426 2204 7445
rect 2219 7426 2249 7442
rect 2191 7410 2265 7426
rect 2191 7408 2204 7410
rect 2219 7408 2253 7410
rect 1856 7386 1869 7388
rect 1884 7386 1918 7388
rect 1856 7370 1918 7386
rect 1962 7381 1976 7384
rect 2040 7381 2070 7392
rect 2118 7388 2164 7404
rect 2191 7392 2265 7408
rect 2118 7386 2152 7388
rect 2117 7370 2164 7386
rect 2191 7370 2204 7392
rect 2219 7370 2249 7392
rect 2276 7370 2277 7386
rect 2292 7370 2305 7530
rect 2335 7426 2348 7530
rect 2393 7508 2394 7518
rect 2409 7508 2422 7518
rect 2393 7504 2422 7508
rect 2427 7504 2457 7530
rect 2475 7516 2491 7518
rect 2563 7516 2616 7530
rect 2564 7514 2628 7516
rect 2671 7514 2686 7530
rect 2735 7527 2765 7530
rect 2735 7524 2771 7527
rect 2701 7516 2717 7518
rect 2475 7504 2490 7508
rect 2393 7502 2490 7504
rect 2518 7502 2686 7514
rect 2702 7504 2717 7508
rect 2735 7505 2774 7524
rect 2793 7518 2800 7519
rect 2799 7511 2800 7518
rect 2783 7508 2784 7511
rect 2799 7508 2812 7511
rect 2735 7504 2765 7505
rect 2774 7504 2780 7505
rect 2783 7504 2812 7508
rect 2702 7503 2812 7504
rect 2702 7502 2818 7503
rect 2377 7494 2428 7502
rect 2377 7482 2402 7494
rect 2409 7482 2428 7494
rect 2459 7494 2509 7502
rect 2459 7486 2475 7494
rect 2482 7492 2509 7494
rect 2518 7492 2739 7502
rect 2482 7482 2739 7492
rect 2768 7494 2818 7502
rect 2768 7485 2784 7494
rect 2377 7474 2428 7482
rect 2475 7474 2739 7482
rect 2765 7482 2784 7485
rect 2791 7482 2818 7494
rect 2765 7474 2818 7482
rect 2393 7466 2394 7474
rect 2409 7466 2422 7474
rect 2393 7458 2409 7466
rect 2390 7451 2409 7454
rect 2390 7442 2412 7451
rect 2363 7432 2412 7442
rect 2363 7426 2393 7432
rect 2412 7427 2417 7432
rect 2335 7410 2409 7426
rect 2427 7418 2457 7474
rect 2492 7464 2700 7474
rect 2735 7470 2780 7474
rect 2783 7473 2784 7474
rect 2799 7473 2812 7474
rect 2518 7434 2707 7464
rect 2533 7431 2707 7434
rect 2526 7428 2707 7431
rect 2335 7408 2348 7410
rect 2363 7408 2397 7410
rect 2335 7392 2409 7408
rect 2436 7404 2449 7418
rect 2464 7404 2480 7420
rect 2526 7415 2537 7428
rect 2319 7370 2320 7386
rect 2335 7370 2348 7392
rect 2363 7370 2393 7392
rect 2436 7388 2498 7404
rect 2526 7397 2537 7413
rect 2542 7408 2552 7428
rect 2562 7408 2576 7428
rect 2579 7415 2588 7428
rect 2604 7415 2613 7428
rect 2542 7397 2576 7408
rect 2579 7397 2588 7413
rect 2604 7397 2613 7413
rect 2620 7408 2630 7428
rect 2640 7408 2654 7428
rect 2655 7415 2666 7428
rect 2620 7397 2654 7408
rect 2655 7397 2666 7413
rect 2712 7404 2728 7420
rect 2735 7418 2765 7470
rect 2799 7466 2800 7473
rect 2784 7458 2800 7466
rect 2771 7426 2784 7445
rect 2799 7426 2829 7442
rect 2771 7410 2845 7426
rect 2771 7408 2784 7410
rect 2799 7408 2833 7410
rect 2436 7386 2449 7388
rect 2464 7386 2498 7388
rect 2436 7370 2498 7386
rect 2542 7381 2558 7384
rect 2620 7381 2650 7392
rect 2698 7388 2744 7404
rect 2771 7392 2845 7408
rect 2698 7386 2732 7388
rect 2697 7370 2744 7386
rect 2771 7370 2784 7392
rect 2799 7370 2829 7392
rect 2856 7370 2857 7386
rect 2872 7370 2885 7530
rect 2915 7426 2928 7530
rect 2973 7508 2974 7518
rect 2989 7508 3002 7518
rect 2973 7504 3002 7508
rect 3007 7504 3037 7530
rect 3055 7516 3071 7518
rect 3143 7516 3196 7530
rect 3144 7514 3208 7516
rect 3251 7514 3266 7530
rect 3315 7527 3345 7530
rect 3315 7524 3351 7527
rect 3281 7516 3297 7518
rect 3055 7504 3070 7508
rect 2973 7502 3070 7504
rect 3098 7502 3266 7514
rect 3282 7504 3297 7508
rect 3315 7505 3354 7524
rect 3373 7518 3380 7519
rect 3379 7511 3380 7518
rect 3363 7508 3364 7511
rect 3379 7508 3392 7511
rect 3315 7504 3345 7505
rect 3354 7504 3360 7505
rect 3363 7504 3392 7508
rect 3282 7503 3392 7504
rect 3282 7502 3398 7503
rect 2957 7494 3008 7502
rect 2957 7482 2982 7494
rect 2989 7482 3008 7494
rect 3039 7494 3089 7502
rect 3039 7486 3055 7494
rect 3062 7492 3089 7494
rect 3098 7492 3319 7502
rect 3062 7482 3319 7492
rect 3348 7494 3398 7502
rect 3348 7485 3364 7494
rect 2957 7474 3008 7482
rect 3055 7474 3319 7482
rect 3345 7482 3364 7485
rect 3371 7482 3398 7494
rect 3345 7474 3398 7482
rect 2973 7466 2974 7474
rect 2989 7466 3002 7474
rect 2973 7458 2989 7466
rect 2970 7451 2989 7454
rect 2970 7442 2992 7451
rect 2943 7432 2992 7442
rect 2943 7426 2973 7432
rect 2992 7427 2997 7432
rect 2915 7410 2989 7426
rect 3007 7418 3037 7474
rect 3072 7464 3280 7474
rect 3315 7470 3360 7474
rect 3363 7473 3364 7474
rect 3379 7473 3392 7474
rect 3098 7434 3287 7464
rect 3113 7431 3287 7434
rect 3106 7428 3287 7431
rect 2915 7408 2928 7410
rect 2943 7408 2977 7410
rect 2915 7392 2989 7408
rect 3016 7404 3029 7418
rect 3044 7404 3060 7420
rect 3106 7415 3117 7428
rect 2899 7370 2900 7386
rect 2915 7370 2928 7392
rect 2943 7370 2973 7392
rect 3016 7388 3078 7404
rect 3106 7397 3117 7413
rect 3122 7408 3132 7428
rect 3142 7408 3156 7428
rect 3159 7415 3168 7428
rect 3184 7415 3193 7428
rect 3122 7397 3156 7408
rect 3159 7397 3168 7413
rect 3184 7397 3193 7413
rect 3200 7408 3210 7428
rect 3220 7408 3234 7428
rect 3235 7415 3246 7428
rect 3200 7397 3234 7408
rect 3235 7397 3246 7413
rect 3292 7404 3308 7420
rect 3315 7418 3345 7470
rect 3379 7466 3380 7473
rect 3364 7458 3380 7466
rect 3351 7426 3364 7445
rect 3379 7426 3409 7442
rect 3351 7410 3425 7426
rect 3351 7408 3364 7410
rect 3379 7408 3413 7410
rect 3016 7386 3029 7388
rect 3044 7386 3078 7388
rect 3016 7370 3078 7386
rect 3122 7381 3138 7384
rect 3200 7381 3230 7392
rect 3278 7388 3324 7404
rect 3351 7392 3425 7408
rect 3278 7386 3312 7388
rect 3277 7370 3324 7386
rect 3351 7370 3364 7392
rect 3379 7370 3409 7392
rect 3436 7370 3437 7386
rect 3452 7370 3465 7530
rect 3495 7426 3508 7530
rect 3553 7508 3554 7518
rect 3569 7508 3582 7518
rect 3553 7504 3582 7508
rect 3587 7504 3617 7530
rect 3635 7516 3651 7518
rect 3723 7516 3776 7530
rect 3724 7514 3788 7516
rect 3831 7514 3846 7530
rect 3895 7527 3925 7530
rect 3895 7524 3931 7527
rect 3861 7516 3877 7518
rect 3635 7504 3650 7508
rect 3553 7502 3650 7504
rect 3678 7502 3846 7514
rect 3862 7504 3877 7508
rect 3895 7505 3934 7524
rect 3953 7518 3960 7519
rect 3959 7511 3960 7518
rect 3943 7508 3944 7511
rect 3959 7508 3972 7511
rect 3895 7504 3925 7505
rect 3934 7504 3940 7505
rect 3943 7504 3972 7508
rect 3862 7503 3972 7504
rect 3862 7502 3978 7503
rect 3537 7494 3588 7502
rect 3537 7482 3562 7494
rect 3569 7482 3588 7494
rect 3619 7494 3669 7502
rect 3619 7486 3635 7494
rect 3642 7492 3669 7494
rect 3678 7492 3899 7502
rect 3642 7482 3899 7492
rect 3928 7494 3978 7502
rect 3928 7485 3944 7494
rect 3537 7474 3588 7482
rect 3635 7474 3899 7482
rect 3925 7482 3944 7485
rect 3951 7482 3978 7494
rect 3925 7474 3978 7482
rect 3553 7466 3554 7474
rect 3569 7466 3582 7474
rect 3553 7458 3569 7466
rect 3550 7451 3569 7454
rect 3550 7442 3572 7451
rect 3523 7432 3572 7442
rect 3523 7426 3553 7432
rect 3572 7427 3577 7432
rect 3495 7410 3569 7426
rect 3587 7418 3617 7474
rect 3652 7464 3860 7474
rect 3895 7470 3940 7474
rect 3943 7473 3944 7474
rect 3959 7473 3972 7474
rect 3678 7434 3867 7464
rect 3693 7431 3867 7434
rect 3686 7428 3867 7431
rect 3495 7408 3508 7410
rect 3523 7408 3557 7410
rect 3495 7392 3569 7408
rect 3596 7404 3609 7418
rect 3624 7404 3640 7420
rect 3686 7415 3697 7428
rect 3479 7370 3480 7386
rect 3495 7370 3508 7392
rect 3523 7370 3553 7392
rect 3596 7388 3658 7404
rect 3686 7397 3697 7413
rect 3702 7408 3712 7428
rect 3722 7408 3736 7428
rect 3739 7415 3748 7428
rect 3764 7415 3773 7428
rect 3702 7397 3736 7408
rect 3739 7397 3748 7413
rect 3764 7397 3773 7413
rect 3780 7408 3790 7428
rect 3800 7408 3814 7428
rect 3815 7415 3826 7428
rect 3780 7397 3814 7408
rect 3815 7397 3826 7413
rect 3872 7404 3888 7420
rect 3895 7418 3925 7470
rect 3959 7466 3960 7473
rect 3944 7458 3960 7466
rect 3931 7426 3944 7445
rect 3959 7426 3989 7442
rect 3931 7410 4005 7426
rect 3931 7408 3944 7410
rect 3959 7408 3993 7410
rect 3596 7386 3609 7388
rect 3624 7386 3658 7388
rect 3596 7370 3658 7386
rect 3702 7381 3718 7384
rect 3780 7381 3810 7392
rect 3858 7388 3904 7404
rect 3931 7392 4005 7408
rect 3858 7386 3892 7388
rect 3857 7370 3904 7386
rect 3931 7370 3944 7392
rect 3959 7370 3989 7392
rect 4016 7370 4017 7386
rect 4032 7370 4045 7530
rect 4075 7426 4088 7530
rect 4133 7508 4134 7518
rect 4149 7508 4162 7518
rect 4133 7504 4162 7508
rect 4167 7504 4197 7530
rect 4215 7516 4231 7518
rect 4303 7516 4356 7530
rect 4304 7514 4368 7516
rect 4411 7514 4426 7530
rect 4475 7527 4505 7530
rect 4475 7524 4511 7527
rect 4441 7516 4457 7518
rect 4215 7504 4230 7508
rect 4133 7502 4230 7504
rect 4258 7502 4426 7514
rect 4442 7504 4457 7508
rect 4475 7505 4514 7524
rect 4533 7518 4540 7519
rect 4539 7511 4540 7518
rect 4523 7508 4524 7511
rect 4539 7508 4552 7511
rect 4475 7504 4505 7505
rect 4514 7504 4520 7505
rect 4523 7504 4552 7508
rect 4442 7503 4552 7504
rect 4442 7502 4558 7503
rect 4117 7494 4168 7502
rect 4117 7482 4142 7494
rect 4149 7482 4168 7494
rect 4199 7494 4249 7502
rect 4199 7486 4215 7494
rect 4222 7492 4249 7494
rect 4258 7492 4479 7502
rect 4222 7482 4479 7492
rect 4508 7494 4558 7502
rect 4508 7485 4524 7494
rect 4117 7474 4168 7482
rect 4215 7474 4479 7482
rect 4505 7482 4524 7485
rect 4531 7482 4558 7494
rect 4505 7474 4558 7482
rect 4133 7466 4134 7474
rect 4149 7466 4162 7474
rect 4133 7458 4149 7466
rect 4130 7451 4149 7454
rect 4130 7442 4152 7451
rect 4103 7432 4152 7442
rect 4103 7426 4133 7432
rect 4152 7427 4157 7432
rect 4075 7410 4149 7426
rect 4167 7418 4197 7474
rect 4232 7464 4440 7474
rect 4475 7470 4520 7474
rect 4523 7473 4524 7474
rect 4539 7473 4552 7474
rect 4258 7434 4447 7464
rect 4273 7431 4447 7434
rect 4266 7428 4447 7431
rect 4075 7408 4088 7410
rect 4103 7408 4137 7410
rect 4075 7392 4149 7408
rect 4176 7404 4189 7418
rect 4204 7404 4220 7420
rect 4266 7415 4277 7428
rect 4059 7370 4060 7386
rect 4075 7370 4088 7392
rect 4103 7370 4133 7392
rect 4176 7388 4238 7404
rect 4266 7397 4277 7413
rect 4282 7408 4292 7428
rect 4302 7408 4316 7428
rect 4319 7415 4328 7428
rect 4344 7415 4353 7428
rect 4282 7397 4316 7408
rect 4319 7397 4328 7413
rect 4344 7397 4353 7413
rect 4360 7408 4370 7428
rect 4380 7408 4394 7428
rect 4395 7415 4406 7428
rect 4360 7397 4394 7408
rect 4395 7397 4406 7413
rect 4452 7404 4468 7420
rect 4475 7418 4505 7470
rect 4539 7466 4540 7473
rect 4524 7458 4540 7466
rect 4511 7426 4524 7445
rect 4539 7426 4569 7442
rect 4511 7410 4585 7426
rect 4511 7408 4524 7410
rect 4539 7408 4573 7410
rect 4176 7386 4189 7388
rect 4204 7386 4238 7388
rect 4176 7370 4238 7386
rect 4282 7381 4298 7384
rect 4360 7381 4390 7392
rect 4438 7388 4484 7404
rect 4511 7392 4585 7408
rect 4438 7386 4472 7388
rect 4437 7370 4484 7386
rect 4511 7370 4524 7392
rect 4539 7370 4569 7392
rect 4596 7370 4597 7386
rect 4612 7370 4625 7530
rect 4655 7426 4668 7530
rect 4713 7508 4714 7518
rect 4729 7508 4742 7518
rect 4713 7504 4742 7508
rect 4747 7504 4777 7530
rect 4795 7516 4811 7518
rect 4883 7516 4936 7530
rect 4884 7514 4948 7516
rect 4991 7514 5006 7530
rect 5055 7527 5085 7530
rect 5055 7524 5091 7527
rect 5021 7516 5037 7518
rect 4795 7504 4810 7508
rect 4713 7502 4810 7504
rect 4838 7502 5006 7514
rect 5022 7504 5037 7508
rect 5055 7505 5094 7524
rect 5113 7518 5120 7519
rect 5119 7511 5120 7518
rect 5103 7508 5104 7511
rect 5119 7508 5132 7511
rect 5055 7504 5085 7505
rect 5094 7504 5100 7505
rect 5103 7504 5132 7508
rect 5022 7503 5132 7504
rect 5022 7502 5138 7503
rect 4697 7494 4748 7502
rect 4697 7482 4722 7494
rect 4729 7482 4748 7494
rect 4779 7494 4829 7502
rect 4779 7486 4795 7494
rect 4802 7492 4829 7494
rect 4838 7492 5059 7502
rect 4802 7482 5059 7492
rect 5088 7494 5138 7502
rect 5088 7485 5104 7494
rect 4697 7474 4748 7482
rect 4795 7474 5059 7482
rect 5085 7482 5104 7485
rect 5111 7482 5138 7494
rect 5085 7474 5138 7482
rect 4713 7466 4714 7474
rect 4729 7466 4742 7474
rect 4713 7458 4729 7466
rect 4710 7451 4729 7454
rect 4710 7442 4732 7451
rect 4683 7432 4732 7442
rect 4683 7426 4713 7432
rect 4732 7427 4737 7432
rect 4655 7410 4729 7426
rect 4747 7418 4777 7474
rect 4812 7464 5020 7474
rect 5055 7470 5100 7474
rect 5103 7473 5104 7474
rect 5119 7473 5132 7474
rect 4838 7434 5027 7464
rect 4853 7431 5027 7434
rect 4846 7428 5027 7431
rect 4655 7408 4668 7410
rect 4683 7408 4717 7410
rect 4655 7392 4729 7408
rect 4756 7404 4769 7418
rect 4784 7404 4800 7420
rect 4846 7415 4857 7428
rect 4639 7370 4640 7386
rect 4655 7370 4668 7392
rect 4683 7370 4713 7392
rect 4756 7388 4818 7404
rect 4846 7397 4857 7413
rect 4862 7408 4872 7428
rect 4882 7408 4896 7428
rect 4899 7415 4908 7428
rect 4924 7415 4933 7428
rect 4862 7397 4896 7408
rect 4899 7397 4908 7413
rect 4924 7397 4933 7413
rect 4940 7408 4950 7428
rect 4960 7408 4974 7428
rect 4975 7415 4986 7428
rect 4940 7397 4974 7408
rect 4975 7397 4986 7413
rect 5032 7404 5048 7420
rect 5055 7418 5085 7470
rect 5119 7466 5120 7473
rect 5104 7458 5120 7466
rect 5091 7426 5104 7445
rect 5119 7426 5149 7442
rect 5091 7410 5165 7426
rect 5091 7408 5104 7410
rect 5119 7408 5153 7410
rect 4756 7386 4769 7388
rect 4784 7386 4818 7388
rect 4756 7370 4818 7386
rect 4862 7381 4878 7384
rect 4940 7381 4970 7392
rect 5018 7388 5064 7404
rect 5091 7392 5165 7408
rect 5018 7386 5052 7388
rect 5017 7370 5064 7386
rect 5091 7370 5104 7392
rect 5119 7370 5149 7392
rect 5176 7370 5177 7386
rect 5192 7370 5205 7530
rect 5235 7426 5248 7530
rect 5293 7508 5294 7518
rect 5309 7508 5322 7518
rect 5293 7504 5322 7508
rect 5327 7504 5357 7530
rect 5375 7516 5391 7518
rect 5463 7516 5516 7530
rect 5464 7514 5528 7516
rect 5571 7514 5586 7530
rect 5635 7527 5665 7530
rect 5635 7524 5671 7527
rect 5601 7516 5617 7518
rect 5375 7504 5390 7508
rect 5293 7502 5390 7504
rect 5418 7502 5586 7514
rect 5602 7504 5617 7508
rect 5635 7505 5674 7524
rect 5693 7518 5700 7519
rect 5699 7511 5700 7518
rect 5683 7508 5684 7511
rect 5699 7508 5712 7511
rect 5635 7504 5665 7505
rect 5674 7504 5680 7505
rect 5683 7504 5712 7508
rect 5602 7503 5712 7504
rect 5602 7502 5718 7503
rect 5277 7494 5328 7502
rect 5277 7482 5302 7494
rect 5309 7482 5328 7494
rect 5359 7494 5409 7502
rect 5359 7486 5375 7494
rect 5382 7492 5409 7494
rect 5418 7492 5639 7502
rect 5382 7482 5639 7492
rect 5668 7494 5718 7502
rect 5668 7485 5684 7494
rect 5277 7474 5328 7482
rect 5375 7474 5639 7482
rect 5665 7482 5684 7485
rect 5691 7482 5718 7494
rect 5665 7474 5718 7482
rect 5293 7466 5294 7474
rect 5309 7466 5322 7474
rect 5293 7458 5309 7466
rect 5290 7451 5309 7454
rect 5290 7442 5312 7451
rect 5263 7432 5312 7442
rect 5263 7426 5293 7432
rect 5312 7427 5317 7432
rect 5235 7410 5309 7426
rect 5327 7418 5357 7474
rect 5392 7464 5600 7474
rect 5635 7470 5680 7474
rect 5683 7473 5684 7474
rect 5699 7473 5712 7474
rect 5418 7434 5607 7464
rect 5433 7431 5607 7434
rect 5426 7428 5607 7431
rect 5235 7408 5248 7410
rect 5263 7408 5297 7410
rect 5235 7392 5309 7408
rect 5336 7404 5349 7418
rect 5364 7404 5380 7420
rect 5426 7415 5437 7428
rect 5219 7370 5220 7386
rect 5235 7370 5248 7392
rect 5263 7370 5293 7392
rect 5336 7388 5398 7404
rect 5426 7397 5437 7413
rect 5442 7408 5452 7428
rect 5462 7408 5476 7428
rect 5479 7415 5488 7428
rect 5504 7415 5513 7428
rect 5442 7397 5476 7408
rect 5479 7397 5488 7413
rect 5504 7397 5513 7413
rect 5520 7408 5530 7428
rect 5540 7408 5554 7428
rect 5555 7415 5566 7428
rect 5520 7397 5554 7408
rect 5555 7397 5566 7413
rect 5612 7404 5628 7420
rect 5635 7418 5665 7470
rect 5699 7466 5700 7473
rect 5684 7458 5700 7466
rect 5671 7426 5684 7445
rect 5699 7426 5729 7442
rect 5671 7410 5745 7426
rect 5671 7408 5684 7410
rect 5699 7408 5733 7410
rect 5336 7386 5349 7388
rect 5364 7386 5398 7388
rect 5336 7370 5398 7386
rect 5442 7381 5458 7384
rect 5520 7381 5550 7392
rect 5598 7388 5644 7404
rect 5671 7392 5745 7408
rect 5598 7386 5632 7388
rect 5597 7370 5644 7386
rect 5671 7370 5684 7392
rect 5699 7370 5729 7392
rect 5756 7370 5757 7386
rect 5772 7370 5785 7530
rect 5815 7426 5828 7530
rect 5873 7508 5874 7518
rect 5889 7508 5902 7518
rect 5873 7504 5902 7508
rect 5907 7504 5937 7530
rect 5955 7516 5971 7518
rect 6043 7516 6096 7530
rect 6044 7514 6108 7516
rect 6151 7514 6166 7530
rect 6215 7527 6245 7530
rect 6215 7524 6251 7527
rect 6181 7516 6197 7518
rect 5955 7504 5970 7508
rect 5873 7502 5970 7504
rect 5998 7502 6166 7514
rect 6182 7504 6197 7508
rect 6215 7505 6254 7524
rect 6273 7518 6280 7519
rect 6279 7511 6280 7518
rect 6263 7508 6264 7511
rect 6279 7508 6292 7511
rect 6215 7504 6245 7505
rect 6254 7504 6260 7505
rect 6263 7504 6292 7508
rect 6182 7503 6292 7504
rect 6182 7502 6298 7503
rect 5857 7494 5908 7502
rect 5857 7482 5882 7494
rect 5889 7482 5908 7494
rect 5939 7494 5989 7502
rect 5939 7486 5955 7494
rect 5962 7492 5989 7494
rect 5998 7492 6219 7502
rect 5962 7482 6219 7492
rect 6248 7494 6298 7502
rect 6248 7485 6264 7494
rect 5857 7474 5908 7482
rect 5955 7474 6219 7482
rect 6245 7482 6264 7485
rect 6271 7482 6298 7494
rect 6245 7474 6298 7482
rect 5873 7466 5874 7474
rect 5889 7466 5902 7474
rect 5873 7458 5889 7466
rect 5870 7451 5889 7454
rect 5870 7442 5892 7451
rect 5843 7432 5892 7442
rect 5843 7426 5873 7432
rect 5892 7427 5897 7432
rect 5815 7410 5889 7426
rect 5907 7418 5937 7474
rect 5972 7464 6180 7474
rect 6215 7470 6260 7474
rect 6263 7473 6264 7474
rect 6279 7473 6292 7474
rect 5998 7434 6187 7464
rect 6013 7431 6187 7434
rect 6006 7428 6187 7431
rect 5815 7408 5828 7410
rect 5843 7408 5877 7410
rect 5815 7392 5889 7408
rect 5916 7404 5929 7418
rect 5944 7404 5960 7420
rect 6006 7415 6017 7428
rect 5799 7370 5800 7386
rect 5815 7370 5828 7392
rect 5843 7370 5873 7392
rect 5916 7388 5978 7404
rect 6006 7397 6017 7413
rect 6022 7408 6032 7428
rect 6042 7408 6056 7428
rect 6059 7415 6068 7428
rect 6084 7415 6093 7428
rect 6022 7397 6056 7408
rect 6059 7397 6068 7413
rect 6084 7397 6093 7413
rect 6100 7408 6110 7428
rect 6120 7408 6134 7428
rect 6135 7415 6146 7428
rect 6100 7397 6134 7408
rect 6135 7397 6146 7413
rect 6192 7404 6208 7420
rect 6215 7418 6245 7470
rect 6279 7466 6280 7473
rect 6264 7458 6280 7466
rect 6251 7426 6264 7445
rect 6279 7426 6309 7442
rect 6251 7410 6325 7426
rect 6251 7408 6264 7410
rect 6279 7408 6313 7410
rect 5916 7386 5929 7388
rect 5944 7386 5978 7388
rect 5916 7370 5978 7386
rect 6022 7381 6038 7384
rect 6100 7381 6130 7392
rect 6178 7388 6224 7404
rect 6251 7392 6325 7408
rect 6178 7386 6212 7388
rect 6177 7370 6224 7386
rect 6251 7370 6264 7392
rect 6279 7370 6309 7392
rect 6336 7370 6337 7386
rect 6352 7370 6365 7530
rect 6395 7426 6408 7530
rect 6453 7508 6454 7518
rect 6469 7508 6482 7518
rect 6453 7504 6482 7508
rect 6487 7504 6517 7530
rect 6535 7516 6551 7518
rect 6623 7516 6676 7530
rect 6624 7514 6688 7516
rect 6731 7514 6746 7530
rect 6795 7527 6825 7530
rect 6795 7524 6831 7527
rect 6761 7516 6777 7518
rect 6535 7504 6550 7508
rect 6453 7502 6550 7504
rect 6578 7502 6746 7514
rect 6762 7504 6777 7508
rect 6795 7505 6834 7524
rect 6853 7518 6860 7519
rect 6859 7511 6860 7518
rect 6843 7508 6844 7511
rect 6859 7508 6872 7511
rect 6795 7504 6825 7505
rect 6834 7504 6840 7505
rect 6843 7504 6872 7508
rect 6762 7503 6872 7504
rect 6762 7502 6878 7503
rect 6437 7494 6488 7502
rect 6437 7482 6462 7494
rect 6469 7482 6488 7494
rect 6519 7494 6569 7502
rect 6519 7486 6535 7494
rect 6542 7492 6569 7494
rect 6578 7492 6799 7502
rect 6542 7482 6799 7492
rect 6828 7494 6878 7502
rect 6828 7485 6844 7494
rect 6437 7474 6488 7482
rect 6535 7474 6799 7482
rect 6825 7482 6844 7485
rect 6851 7482 6878 7494
rect 6825 7474 6878 7482
rect 6453 7466 6454 7474
rect 6469 7466 6482 7474
rect 6453 7458 6469 7466
rect 6450 7451 6469 7454
rect 6450 7442 6472 7451
rect 6423 7432 6472 7442
rect 6423 7426 6453 7432
rect 6472 7427 6477 7432
rect 6395 7410 6469 7426
rect 6487 7418 6517 7474
rect 6552 7464 6760 7474
rect 6795 7470 6840 7474
rect 6843 7473 6844 7474
rect 6859 7473 6872 7474
rect 6578 7434 6767 7464
rect 6593 7431 6767 7434
rect 6586 7428 6767 7431
rect 6395 7408 6408 7410
rect 6423 7408 6457 7410
rect 6395 7392 6469 7408
rect 6496 7404 6509 7418
rect 6524 7404 6540 7420
rect 6586 7415 6597 7428
rect 6379 7370 6380 7386
rect 6395 7370 6408 7392
rect 6423 7370 6453 7392
rect 6496 7388 6558 7404
rect 6586 7397 6597 7413
rect 6602 7408 6612 7428
rect 6622 7408 6636 7428
rect 6639 7415 6648 7428
rect 6664 7415 6673 7428
rect 6602 7397 6636 7408
rect 6639 7397 6648 7413
rect 6664 7397 6673 7413
rect 6680 7408 6690 7428
rect 6700 7408 6714 7428
rect 6715 7415 6726 7428
rect 6680 7397 6714 7408
rect 6715 7397 6726 7413
rect 6772 7404 6788 7420
rect 6795 7418 6825 7470
rect 6859 7466 6860 7473
rect 6844 7458 6860 7466
rect 6831 7426 6844 7445
rect 6859 7426 6889 7442
rect 6831 7410 6905 7426
rect 6831 7408 6844 7410
rect 6859 7408 6893 7410
rect 6496 7386 6509 7388
rect 6524 7386 6558 7388
rect 6496 7370 6558 7386
rect 6602 7381 6618 7384
rect 6680 7381 6710 7392
rect 6758 7388 6804 7404
rect 6831 7392 6905 7408
rect 6758 7386 6792 7388
rect 6757 7370 6804 7386
rect 6831 7370 6844 7392
rect 6859 7370 6889 7392
rect 6916 7370 6917 7386
rect 6932 7370 6945 7530
rect 6975 7426 6988 7530
rect 7033 7508 7034 7518
rect 7049 7508 7062 7518
rect 7033 7504 7062 7508
rect 7067 7504 7097 7530
rect 7115 7516 7131 7518
rect 7203 7516 7256 7530
rect 7204 7514 7268 7516
rect 7311 7514 7326 7530
rect 7375 7527 7405 7530
rect 7375 7524 7411 7527
rect 7341 7516 7357 7518
rect 7115 7504 7130 7508
rect 7033 7502 7130 7504
rect 7158 7502 7326 7514
rect 7342 7504 7357 7508
rect 7375 7505 7414 7524
rect 7433 7518 7440 7519
rect 7439 7511 7440 7518
rect 7423 7508 7424 7511
rect 7439 7508 7452 7511
rect 7375 7504 7405 7505
rect 7414 7504 7420 7505
rect 7423 7504 7452 7508
rect 7342 7503 7452 7504
rect 7342 7502 7458 7503
rect 7017 7494 7068 7502
rect 7017 7482 7042 7494
rect 7049 7482 7068 7494
rect 7099 7494 7149 7502
rect 7099 7486 7115 7494
rect 7122 7492 7149 7494
rect 7158 7492 7379 7502
rect 7122 7482 7379 7492
rect 7408 7494 7458 7502
rect 7408 7485 7424 7494
rect 7017 7474 7068 7482
rect 7115 7474 7379 7482
rect 7405 7482 7424 7485
rect 7431 7482 7458 7494
rect 7405 7474 7458 7482
rect 7033 7466 7034 7474
rect 7049 7466 7062 7474
rect 7033 7458 7049 7466
rect 7030 7451 7049 7454
rect 7030 7442 7052 7451
rect 7003 7432 7052 7442
rect 7003 7426 7033 7432
rect 7052 7427 7057 7432
rect 6975 7410 7049 7426
rect 7067 7418 7097 7474
rect 7132 7464 7340 7474
rect 7375 7470 7420 7474
rect 7423 7473 7424 7474
rect 7439 7473 7452 7474
rect 7158 7434 7347 7464
rect 7173 7431 7347 7434
rect 7166 7428 7347 7431
rect 6975 7408 6988 7410
rect 7003 7408 7037 7410
rect 6975 7392 7049 7408
rect 7076 7404 7089 7418
rect 7104 7404 7120 7420
rect 7166 7415 7177 7428
rect 6959 7370 6960 7386
rect 6975 7370 6988 7392
rect 7003 7370 7033 7392
rect 7076 7388 7138 7404
rect 7166 7397 7177 7413
rect 7182 7408 7192 7428
rect 7202 7408 7216 7428
rect 7219 7415 7228 7428
rect 7244 7415 7253 7428
rect 7182 7397 7216 7408
rect 7219 7397 7228 7413
rect 7244 7397 7253 7413
rect 7260 7408 7270 7428
rect 7280 7408 7294 7428
rect 7295 7415 7306 7428
rect 7260 7397 7294 7408
rect 7295 7397 7306 7413
rect 7352 7404 7368 7420
rect 7375 7418 7405 7470
rect 7439 7466 7440 7473
rect 7424 7458 7440 7466
rect 7411 7426 7424 7445
rect 7439 7426 7469 7442
rect 7411 7410 7485 7426
rect 7411 7408 7424 7410
rect 7439 7408 7473 7410
rect 7076 7386 7089 7388
rect 7104 7386 7138 7388
rect 7076 7370 7138 7386
rect 7182 7381 7198 7384
rect 7260 7381 7290 7392
rect 7338 7388 7384 7404
rect 7411 7392 7485 7408
rect 7338 7386 7372 7388
rect 7337 7370 7384 7386
rect 7411 7370 7424 7392
rect 7439 7370 7469 7392
rect 7496 7370 7497 7386
rect 7512 7370 7525 7530
rect 7555 7426 7568 7530
rect 7613 7508 7614 7518
rect 7629 7508 7642 7518
rect 7613 7504 7642 7508
rect 7647 7504 7677 7530
rect 7695 7516 7711 7518
rect 7783 7516 7836 7530
rect 7784 7514 7848 7516
rect 7891 7514 7906 7530
rect 7955 7527 7985 7530
rect 7955 7524 7991 7527
rect 7921 7516 7937 7518
rect 7695 7504 7710 7508
rect 7613 7502 7710 7504
rect 7738 7502 7906 7514
rect 7922 7504 7937 7508
rect 7955 7505 7994 7524
rect 8013 7518 8020 7519
rect 8019 7511 8020 7518
rect 8003 7508 8004 7511
rect 8019 7508 8032 7511
rect 7955 7504 7985 7505
rect 7994 7504 8000 7505
rect 8003 7504 8032 7508
rect 7922 7503 8032 7504
rect 7922 7502 8038 7503
rect 7597 7494 7648 7502
rect 7597 7482 7622 7494
rect 7629 7482 7648 7494
rect 7679 7494 7729 7502
rect 7679 7486 7695 7494
rect 7702 7492 7729 7494
rect 7738 7492 7959 7502
rect 7702 7482 7959 7492
rect 7988 7494 8038 7502
rect 7988 7485 8004 7494
rect 7597 7474 7648 7482
rect 7695 7474 7959 7482
rect 7985 7482 8004 7485
rect 8011 7482 8038 7494
rect 7985 7474 8038 7482
rect 7613 7466 7614 7474
rect 7629 7466 7642 7474
rect 7613 7458 7629 7466
rect 7610 7451 7629 7454
rect 7610 7442 7632 7451
rect 7583 7432 7632 7442
rect 7583 7426 7613 7432
rect 7632 7427 7637 7432
rect 7555 7410 7629 7426
rect 7647 7418 7677 7474
rect 7712 7464 7920 7474
rect 7955 7470 8000 7474
rect 8003 7473 8004 7474
rect 8019 7473 8032 7474
rect 7738 7434 7927 7464
rect 7753 7431 7927 7434
rect 7746 7428 7927 7431
rect 7555 7408 7568 7410
rect 7583 7408 7617 7410
rect 7555 7392 7629 7408
rect 7656 7404 7669 7418
rect 7684 7404 7700 7420
rect 7746 7415 7757 7428
rect 7539 7370 7540 7386
rect 7555 7370 7568 7392
rect 7583 7370 7613 7392
rect 7656 7388 7718 7404
rect 7746 7397 7757 7413
rect 7762 7408 7772 7428
rect 7782 7408 7796 7428
rect 7799 7415 7808 7428
rect 7824 7415 7833 7428
rect 7762 7397 7796 7408
rect 7799 7397 7808 7413
rect 7824 7397 7833 7413
rect 7840 7408 7850 7428
rect 7860 7408 7874 7428
rect 7875 7415 7886 7428
rect 7840 7397 7874 7408
rect 7875 7397 7886 7413
rect 7932 7404 7948 7420
rect 7955 7418 7985 7470
rect 8019 7466 8020 7473
rect 8004 7458 8020 7466
rect 7991 7426 8004 7445
rect 8019 7426 8049 7442
rect 7991 7410 8065 7426
rect 7991 7408 8004 7410
rect 8019 7408 8053 7410
rect 7656 7386 7669 7388
rect 7684 7386 7718 7388
rect 7656 7370 7718 7386
rect 7762 7381 7778 7384
rect 7840 7381 7870 7392
rect 7918 7388 7964 7404
rect 7991 7392 8065 7408
rect 7918 7386 7952 7388
rect 7917 7370 7964 7386
rect 7991 7370 8004 7392
rect 8019 7370 8049 7392
rect 8076 7370 8077 7386
rect 8092 7370 8105 7530
rect 8135 7426 8148 7530
rect 8193 7508 8194 7518
rect 8209 7508 8222 7518
rect 8193 7504 8222 7508
rect 8227 7504 8257 7530
rect 8275 7516 8291 7518
rect 8363 7516 8416 7530
rect 8364 7514 8428 7516
rect 8471 7514 8486 7530
rect 8535 7527 8565 7530
rect 8535 7524 8571 7527
rect 8501 7516 8517 7518
rect 8275 7504 8290 7508
rect 8193 7502 8290 7504
rect 8318 7502 8486 7514
rect 8502 7504 8517 7508
rect 8535 7505 8574 7524
rect 8593 7518 8600 7519
rect 8599 7511 8600 7518
rect 8583 7508 8584 7511
rect 8599 7508 8612 7511
rect 8535 7504 8565 7505
rect 8574 7504 8580 7505
rect 8583 7504 8612 7508
rect 8502 7503 8612 7504
rect 8502 7502 8618 7503
rect 8177 7494 8228 7502
rect 8177 7482 8202 7494
rect 8209 7482 8228 7494
rect 8259 7494 8309 7502
rect 8259 7486 8275 7494
rect 8282 7492 8309 7494
rect 8318 7492 8539 7502
rect 8282 7482 8539 7492
rect 8568 7494 8618 7502
rect 8568 7485 8584 7494
rect 8177 7474 8228 7482
rect 8275 7474 8539 7482
rect 8565 7482 8584 7485
rect 8591 7482 8618 7494
rect 8565 7474 8618 7482
rect 8193 7466 8194 7474
rect 8209 7466 8222 7474
rect 8193 7458 8209 7466
rect 8190 7451 8209 7454
rect 8190 7442 8212 7451
rect 8163 7432 8212 7442
rect 8163 7426 8193 7432
rect 8212 7427 8217 7432
rect 8135 7410 8209 7426
rect 8227 7418 8257 7474
rect 8292 7464 8500 7474
rect 8535 7470 8580 7474
rect 8583 7473 8584 7474
rect 8599 7473 8612 7474
rect 8318 7434 8507 7464
rect 8333 7431 8507 7434
rect 8326 7428 8507 7431
rect 8135 7408 8148 7410
rect 8163 7408 8197 7410
rect 8135 7392 8209 7408
rect 8236 7404 8249 7418
rect 8264 7404 8280 7420
rect 8326 7415 8337 7428
rect 8119 7370 8120 7386
rect 8135 7370 8148 7392
rect 8163 7370 8193 7392
rect 8236 7388 8298 7404
rect 8326 7397 8337 7413
rect 8342 7408 8352 7428
rect 8362 7408 8376 7428
rect 8379 7415 8388 7428
rect 8404 7415 8413 7428
rect 8342 7397 8376 7408
rect 8379 7397 8388 7413
rect 8404 7397 8413 7413
rect 8420 7408 8430 7428
rect 8440 7408 8454 7428
rect 8455 7415 8466 7428
rect 8420 7397 8454 7408
rect 8455 7397 8466 7413
rect 8512 7404 8528 7420
rect 8535 7418 8565 7470
rect 8599 7466 8600 7473
rect 8584 7458 8600 7466
rect 8571 7426 8584 7445
rect 8599 7426 8629 7442
rect 8571 7410 8645 7426
rect 8571 7408 8584 7410
rect 8599 7408 8633 7410
rect 8236 7386 8249 7388
rect 8264 7386 8298 7388
rect 8236 7370 8298 7386
rect 8342 7381 8358 7384
rect 8420 7381 8450 7392
rect 8498 7388 8544 7404
rect 8571 7392 8645 7408
rect 8498 7386 8532 7388
rect 8497 7370 8544 7386
rect 8571 7370 8584 7392
rect 8599 7370 8629 7392
rect 8656 7370 8657 7386
rect 8672 7370 8685 7530
rect 8715 7426 8728 7530
rect 8773 7508 8774 7518
rect 8789 7508 8802 7518
rect 8773 7504 8802 7508
rect 8807 7504 8837 7530
rect 8855 7516 8871 7518
rect 8943 7516 8996 7530
rect 8944 7514 9008 7516
rect 9051 7514 9066 7530
rect 9115 7527 9145 7530
rect 9115 7524 9151 7527
rect 9081 7516 9097 7518
rect 8855 7504 8870 7508
rect 8773 7502 8870 7504
rect 8898 7502 9066 7514
rect 9082 7504 9097 7508
rect 9115 7505 9154 7524
rect 9173 7518 9180 7519
rect 9179 7511 9180 7518
rect 9163 7508 9164 7511
rect 9179 7508 9192 7511
rect 9115 7504 9145 7505
rect 9154 7504 9160 7505
rect 9163 7504 9192 7508
rect 9082 7503 9192 7504
rect 9082 7502 9198 7503
rect 8757 7494 8808 7502
rect 8757 7482 8782 7494
rect 8789 7482 8808 7494
rect 8839 7494 8889 7502
rect 8839 7486 8855 7494
rect 8862 7492 8889 7494
rect 8898 7492 9119 7502
rect 8862 7482 9119 7492
rect 9148 7494 9198 7502
rect 9148 7485 9164 7494
rect 8757 7474 8808 7482
rect 8855 7474 9119 7482
rect 9145 7482 9164 7485
rect 9171 7482 9198 7494
rect 9145 7474 9198 7482
rect 8773 7466 8774 7474
rect 8789 7466 8802 7474
rect 8773 7458 8789 7466
rect 8770 7451 8789 7454
rect 8770 7442 8792 7451
rect 8743 7432 8792 7442
rect 8743 7426 8773 7432
rect 8792 7427 8797 7432
rect 8715 7410 8789 7426
rect 8807 7418 8837 7474
rect 8872 7464 9080 7474
rect 9115 7470 9160 7474
rect 9163 7473 9164 7474
rect 9179 7473 9192 7474
rect 8898 7434 9087 7464
rect 8913 7431 9087 7434
rect 8906 7428 9087 7431
rect 8715 7408 8728 7410
rect 8743 7408 8777 7410
rect 8715 7392 8789 7408
rect 8816 7404 8829 7418
rect 8844 7404 8860 7420
rect 8906 7415 8917 7428
rect 8699 7370 8700 7386
rect 8715 7370 8728 7392
rect 8743 7370 8773 7392
rect 8816 7388 8878 7404
rect 8906 7397 8917 7413
rect 8922 7408 8932 7428
rect 8942 7408 8956 7428
rect 8959 7415 8968 7428
rect 8984 7415 8993 7428
rect 8922 7397 8956 7408
rect 8959 7397 8968 7413
rect 8984 7397 8993 7413
rect 9000 7408 9010 7428
rect 9020 7408 9034 7428
rect 9035 7415 9046 7428
rect 9000 7397 9034 7408
rect 9035 7397 9046 7413
rect 9092 7404 9108 7420
rect 9115 7418 9145 7470
rect 9179 7466 9180 7473
rect 9164 7458 9180 7466
rect 9151 7426 9164 7445
rect 9179 7426 9209 7442
rect 9151 7410 9225 7426
rect 9151 7408 9164 7410
rect 9179 7408 9213 7410
rect 8816 7386 8829 7388
rect 8844 7386 8878 7388
rect 8816 7370 8878 7386
rect 8922 7381 8938 7384
rect 9000 7381 9030 7392
rect 9078 7388 9124 7404
rect 9151 7392 9225 7408
rect 9078 7386 9112 7388
rect 9077 7370 9124 7386
rect 9151 7370 9164 7392
rect 9179 7370 9209 7392
rect 9236 7370 9237 7386
rect 9252 7370 9265 7530
rect -7 7362 34 7370
rect -7 7336 8 7362
rect 15 7336 34 7362
rect 98 7358 160 7370
rect 172 7358 247 7370
rect 305 7358 380 7370
rect 392 7358 423 7370
rect 429 7358 464 7370
rect 98 7356 260 7358
rect -7 7328 34 7336
rect 116 7332 129 7356
rect 144 7354 159 7356
rect -1 7318 0 7328
rect 15 7318 28 7328
rect 43 7318 73 7332
rect 116 7318 159 7332
rect 183 7329 190 7336
rect 193 7332 260 7356
rect 292 7356 464 7358
rect 262 7334 290 7338
rect 292 7334 372 7356
rect 393 7354 408 7356
rect 262 7332 372 7334
rect 193 7328 372 7332
rect 166 7318 196 7328
rect 198 7318 351 7328
rect 359 7318 389 7328
rect 393 7318 423 7332
rect 451 7318 464 7356
rect 536 7362 571 7370
rect 536 7336 537 7362
rect 544 7336 571 7362
rect 479 7318 509 7332
rect 536 7328 571 7336
rect 573 7362 614 7370
rect 573 7336 588 7362
rect 595 7336 614 7362
rect 678 7358 740 7370
rect 752 7358 827 7370
rect 885 7358 960 7370
rect 972 7358 1003 7370
rect 1009 7358 1044 7370
rect 678 7356 840 7358
rect 573 7328 614 7336
rect 696 7332 709 7356
rect 724 7354 739 7356
rect 536 7318 537 7328
rect 552 7318 565 7328
rect 579 7318 580 7328
rect 595 7318 608 7328
rect 623 7318 653 7332
rect 696 7318 739 7332
rect 763 7329 770 7336
rect 773 7332 840 7356
rect 872 7356 1044 7358
rect 842 7334 870 7338
rect 872 7334 952 7356
rect 973 7354 988 7356
rect 842 7332 952 7334
rect 773 7328 952 7332
rect 746 7318 776 7328
rect 778 7318 931 7328
rect 939 7318 969 7328
rect 973 7318 1003 7332
rect 1031 7318 1044 7356
rect 1116 7362 1151 7370
rect 1116 7336 1117 7362
rect 1124 7336 1151 7362
rect 1059 7318 1089 7332
rect 1116 7328 1151 7336
rect 1153 7362 1194 7370
rect 1153 7336 1168 7362
rect 1175 7336 1194 7362
rect 1258 7358 1320 7370
rect 1332 7358 1407 7370
rect 1465 7358 1540 7370
rect 1552 7358 1583 7370
rect 1589 7358 1624 7370
rect 1258 7356 1420 7358
rect 1153 7328 1194 7336
rect 1276 7332 1289 7356
rect 1304 7354 1319 7356
rect 1116 7318 1117 7328
rect 1132 7318 1145 7328
rect 1159 7318 1160 7328
rect 1175 7318 1188 7328
rect 1203 7318 1233 7332
rect 1276 7318 1319 7332
rect 1343 7329 1350 7336
rect 1353 7332 1420 7356
rect 1452 7356 1624 7358
rect 1422 7334 1450 7338
rect 1452 7334 1532 7356
rect 1553 7354 1568 7356
rect 1422 7332 1532 7334
rect 1353 7328 1532 7332
rect 1326 7318 1356 7328
rect 1358 7318 1511 7328
rect 1519 7318 1549 7328
rect 1553 7318 1583 7332
rect 1611 7318 1624 7356
rect 1696 7362 1731 7370
rect 1696 7336 1697 7362
rect 1704 7336 1731 7362
rect 1639 7318 1669 7332
rect 1696 7328 1731 7336
rect 1733 7362 1774 7370
rect 1733 7336 1748 7362
rect 1755 7336 1774 7362
rect 1838 7358 1900 7370
rect 1912 7358 1987 7370
rect 2045 7358 2120 7370
rect 2132 7358 2163 7370
rect 2169 7358 2204 7370
rect 1838 7356 2000 7358
rect 1733 7328 1774 7336
rect 1856 7332 1869 7356
rect 1884 7354 1899 7356
rect 1696 7318 1697 7328
rect 1712 7318 1725 7328
rect 1739 7318 1740 7328
rect 1755 7318 1768 7328
rect 1783 7318 1813 7332
rect 1856 7318 1899 7332
rect 1923 7329 1930 7336
rect 1933 7332 2000 7356
rect 2032 7356 2204 7358
rect 2002 7334 2030 7338
rect 2032 7334 2112 7356
rect 2133 7354 2148 7356
rect 2002 7332 2112 7334
rect 1933 7328 2112 7332
rect 1906 7318 1936 7328
rect 1938 7318 2091 7328
rect 2099 7318 2129 7328
rect 2133 7318 2163 7332
rect 2191 7318 2204 7356
rect 2276 7362 2311 7370
rect 2276 7336 2277 7362
rect 2284 7336 2311 7362
rect 2219 7318 2249 7332
rect 2276 7328 2311 7336
rect 2313 7362 2354 7370
rect 2313 7336 2328 7362
rect 2335 7336 2354 7362
rect 2418 7358 2480 7370
rect 2492 7358 2567 7370
rect 2625 7358 2700 7370
rect 2712 7358 2743 7370
rect 2749 7358 2784 7370
rect 2418 7356 2580 7358
rect 2313 7328 2354 7336
rect 2436 7332 2449 7356
rect 2464 7354 2479 7356
rect 2276 7318 2277 7328
rect 2292 7318 2305 7328
rect 2319 7318 2320 7328
rect 2335 7318 2348 7328
rect 2363 7318 2393 7332
rect 2436 7318 2479 7332
rect 2503 7329 2510 7336
rect 2513 7332 2580 7356
rect 2612 7356 2784 7358
rect 2582 7334 2610 7338
rect 2612 7334 2692 7356
rect 2713 7354 2728 7356
rect 2582 7332 2692 7334
rect 2513 7328 2692 7332
rect 2486 7318 2516 7328
rect 2518 7318 2671 7328
rect 2679 7318 2709 7328
rect 2713 7318 2743 7332
rect 2771 7318 2784 7356
rect 2856 7362 2891 7370
rect 2856 7336 2857 7362
rect 2864 7336 2891 7362
rect 2799 7318 2829 7332
rect 2856 7328 2891 7336
rect 2893 7362 2934 7370
rect 2893 7336 2908 7362
rect 2915 7336 2934 7362
rect 2998 7358 3060 7370
rect 3072 7358 3147 7370
rect 3205 7358 3280 7370
rect 3292 7358 3323 7370
rect 3329 7358 3364 7370
rect 2998 7356 3160 7358
rect 2893 7328 2934 7336
rect 3016 7332 3029 7356
rect 3044 7354 3059 7356
rect 2856 7318 2857 7328
rect 2872 7318 2885 7328
rect 2899 7318 2900 7328
rect 2915 7318 2928 7328
rect 2943 7318 2973 7332
rect 3016 7318 3059 7332
rect 3083 7329 3090 7336
rect 3093 7332 3160 7356
rect 3192 7356 3364 7358
rect 3162 7334 3190 7338
rect 3192 7334 3272 7356
rect 3293 7354 3308 7356
rect 3162 7332 3272 7334
rect 3093 7328 3272 7332
rect 3066 7318 3096 7328
rect 3098 7318 3251 7328
rect 3259 7318 3289 7328
rect 3293 7318 3323 7332
rect 3351 7318 3364 7356
rect 3436 7362 3471 7370
rect 3436 7336 3437 7362
rect 3444 7336 3471 7362
rect 3379 7318 3409 7332
rect 3436 7328 3471 7336
rect 3473 7362 3514 7370
rect 3473 7336 3488 7362
rect 3495 7336 3514 7362
rect 3578 7358 3640 7370
rect 3652 7358 3727 7370
rect 3785 7358 3860 7370
rect 3872 7358 3903 7370
rect 3909 7358 3944 7370
rect 3578 7356 3740 7358
rect 3473 7328 3514 7336
rect 3596 7332 3609 7356
rect 3624 7354 3639 7356
rect 3436 7318 3437 7328
rect 3452 7318 3465 7328
rect 3479 7318 3480 7328
rect 3495 7318 3508 7328
rect 3523 7318 3553 7332
rect 3596 7318 3639 7332
rect 3663 7329 3670 7336
rect 3673 7332 3740 7356
rect 3772 7356 3944 7358
rect 3742 7334 3770 7338
rect 3772 7334 3852 7356
rect 3873 7354 3888 7356
rect 3742 7332 3852 7334
rect 3673 7328 3852 7332
rect 3646 7318 3676 7328
rect 3678 7318 3831 7328
rect 3839 7318 3869 7328
rect 3873 7318 3903 7332
rect 3931 7318 3944 7356
rect 4016 7362 4051 7370
rect 4016 7336 4017 7362
rect 4024 7336 4051 7362
rect 3959 7318 3989 7332
rect 4016 7328 4051 7336
rect 4053 7362 4094 7370
rect 4053 7336 4068 7362
rect 4075 7336 4094 7362
rect 4158 7358 4220 7370
rect 4232 7358 4307 7370
rect 4365 7358 4440 7370
rect 4452 7358 4483 7370
rect 4489 7358 4524 7370
rect 4158 7356 4320 7358
rect 4053 7328 4094 7336
rect 4176 7332 4189 7356
rect 4204 7354 4219 7356
rect 4016 7318 4017 7328
rect 4032 7318 4045 7328
rect 4059 7318 4060 7328
rect 4075 7318 4088 7328
rect 4103 7318 4133 7332
rect 4176 7318 4219 7332
rect 4243 7329 4250 7336
rect 4253 7332 4320 7356
rect 4352 7356 4524 7358
rect 4322 7334 4350 7338
rect 4352 7334 4432 7356
rect 4453 7354 4468 7356
rect 4322 7332 4432 7334
rect 4253 7328 4432 7332
rect 4226 7318 4256 7328
rect 4258 7318 4411 7328
rect 4419 7318 4449 7328
rect 4453 7318 4483 7332
rect 4511 7318 4524 7356
rect 4596 7362 4631 7370
rect 4596 7336 4597 7362
rect 4604 7336 4631 7362
rect 4539 7318 4569 7332
rect 4596 7328 4631 7336
rect 4633 7362 4674 7370
rect 4633 7336 4648 7362
rect 4655 7336 4674 7362
rect 4738 7358 4800 7370
rect 4812 7358 4887 7370
rect 4945 7358 5020 7370
rect 5032 7358 5063 7370
rect 5069 7358 5104 7370
rect 4738 7356 4900 7358
rect 4633 7328 4674 7336
rect 4756 7332 4769 7356
rect 4784 7354 4799 7356
rect 4596 7318 4597 7328
rect 4612 7318 4625 7328
rect 4639 7318 4640 7328
rect 4655 7318 4668 7328
rect 4683 7318 4713 7332
rect 4756 7318 4799 7332
rect 4823 7329 4830 7336
rect 4833 7332 4900 7356
rect 4932 7356 5104 7358
rect 4902 7334 4930 7338
rect 4932 7334 5012 7356
rect 5033 7354 5048 7356
rect 4902 7332 5012 7334
rect 4833 7328 5012 7332
rect 4806 7318 4836 7328
rect 4838 7318 4991 7328
rect 4999 7318 5029 7328
rect 5033 7318 5063 7332
rect 5091 7318 5104 7356
rect 5176 7362 5211 7370
rect 5176 7336 5177 7362
rect 5184 7336 5211 7362
rect 5119 7318 5149 7332
rect 5176 7328 5211 7336
rect 5213 7362 5254 7370
rect 5213 7336 5228 7362
rect 5235 7336 5254 7362
rect 5318 7358 5380 7370
rect 5392 7358 5467 7370
rect 5525 7358 5600 7370
rect 5612 7358 5643 7370
rect 5649 7358 5684 7370
rect 5318 7356 5480 7358
rect 5213 7328 5254 7336
rect 5336 7332 5349 7356
rect 5364 7354 5379 7356
rect 5176 7318 5177 7328
rect 5192 7318 5205 7328
rect 5219 7318 5220 7328
rect 5235 7318 5248 7328
rect 5263 7318 5293 7332
rect 5336 7318 5379 7332
rect 5403 7329 5410 7336
rect 5413 7332 5480 7356
rect 5512 7356 5684 7358
rect 5482 7334 5510 7338
rect 5512 7334 5592 7356
rect 5613 7354 5628 7356
rect 5482 7332 5592 7334
rect 5413 7328 5592 7332
rect 5386 7318 5416 7328
rect 5418 7318 5571 7328
rect 5579 7318 5609 7328
rect 5613 7318 5643 7332
rect 5671 7318 5684 7356
rect 5756 7362 5791 7370
rect 5756 7336 5757 7362
rect 5764 7336 5791 7362
rect 5699 7318 5729 7332
rect 5756 7328 5791 7336
rect 5793 7362 5834 7370
rect 5793 7336 5808 7362
rect 5815 7336 5834 7362
rect 5898 7358 5960 7370
rect 5972 7358 6047 7370
rect 6105 7358 6180 7370
rect 6192 7358 6223 7370
rect 6229 7358 6264 7370
rect 5898 7356 6060 7358
rect 5793 7328 5834 7336
rect 5916 7332 5929 7356
rect 5944 7354 5959 7356
rect 5756 7318 5757 7328
rect 5772 7318 5785 7328
rect 5799 7318 5800 7328
rect 5815 7318 5828 7328
rect 5843 7318 5873 7332
rect 5916 7318 5959 7332
rect 5983 7329 5990 7336
rect 5993 7332 6060 7356
rect 6092 7356 6264 7358
rect 6062 7334 6090 7338
rect 6092 7334 6172 7356
rect 6193 7354 6208 7356
rect 6062 7332 6172 7334
rect 5993 7328 6172 7332
rect 5966 7318 5996 7328
rect 5998 7318 6151 7328
rect 6159 7318 6189 7328
rect 6193 7318 6223 7332
rect 6251 7318 6264 7356
rect 6336 7362 6371 7370
rect 6336 7336 6337 7362
rect 6344 7336 6371 7362
rect 6279 7318 6309 7332
rect 6336 7328 6371 7336
rect 6373 7362 6414 7370
rect 6373 7336 6388 7362
rect 6395 7336 6414 7362
rect 6478 7358 6540 7370
rect 6552 7358 6627 7370
rect 6685 7358 6760 7370
rect 6772 7358 6803 7370
rect 6809 7358 6844 7370
rect 6478 7356 6640 7358
rect 6373 7328 6414 7336
rect 6496 7332 6509 7356
rect 6524 7354 6539 7356
rect 6336 7318 6337 7328
rect 6352 7318 6365 7328
rect 6379 7318 6380 7328
rect 6395 7318 6408 7328
rect 6423 7318 6453 7332
rect 6496 7318 6539 7332
rect 6563 7329 6570 7336
rect 6573 7332 6640 7356
rect 6672 7356 6844 7358
rect 6642 7334 6670 7338
rect 6672 7334 6752 7356
rect 6773 7354 6788 7356
rect 6642 7332 6752 7334
rect 6573 7328 6752 7332
rect 6546 7318 6576 7328
rect 6578 7318 6731 7328
rect 6739 7318 6769 7328
rect 6773 7318 6803 7332
rect 6831 7318 6844 7356
rect 6916 7362 6951 7370
rect 6916 7336 6917 7362
rect 6924 7336 6951 7362
rect 6859 7318 6889 7332
rect 6916 7328 6951 7336
rect 6953 7362 6994 7370
rect 6953 7336 6968 7362
rect 6975 7336 6994 7362
rect 7058 7358 7120 7370
rect 7132 7358 7207 7370
rect 7265 7358 7340 7370
rect 7352 7358 7383 7370
rect 7389 7358 7424 7370
rect 7058 7356 7220 7358
rect 6953 7328 6994 7336
rect 7076 7332 7089 7356
rect 7104 7354 7119 7356
rect 6916 7318 6917 7328
rect 6932 7318 6945 7328
rect 6959 7318 6960 7328
rect 6975 7318 6988 7328
rect 7003 7318 7033 7332
rect 7076 7318 7119 7332
rect 7143 7329 7150 7336
rect 7153 7332 7220 7356
rect 7252 7356 7424 7358
rect 7222 7334 7250 7338
rect 7252 7334 7332 7356
rect 7353 7354 7368 7356
rect 7222 7332 7332 7334
rect 7153 7328 7332 7332
rect 7126 7318 7156 7328
rect 7158 7318 7311 7328
rect 7319 7318 7349 7328
rect 7353 7318 7383 7332
rect 7411 7318 7424 7356
rect 7496 7362 7531 7370
rect 7496 7336 7497 7362
rect 7504 7336 7531 7362
rect 7439 7318 7469 7332
rect 7496 7328 7531 7336
rect 7533 7362 7574 7370
rect 7533 7336 7548 7362
rect 7555 7336 7574 7362
rect 7638 7358 7700 7370
rect 7712 7358 7787 7370
rect 7845 7358 7920 7370
rect 7932 7358 7963 7370
rect 7969 7358 8004 7370
rect 7638 7356 7800 7358
rect 7533 7328 7574 7336
rect 7656 7332 7669 7356
rect 7684 7354 7699 7356
rect 7496 7318 7497 7328
rect 7512 7318 7525 7328
rect 7539 7318 7540 7328
rect 7555 7318 7568 7328
rect 7583 7318 7613 7332
rect 7656 7318 7699 7332
rect 7723 7329 7730 7336
rect 7733 7332 7800 7356
rect 7832 7356 8004 7358
rect 7802 7334 7830 7338
rect 7832 7334 7912 7356
rect 7933 7354 7948 7356
rect 7802 7332 7912 7334
rect 7733 7328 7912 7332
rect 7706 7318 7736 7328
rect 7738 7318 7891 7328
rect 7899 7318 7929 7328
rect 7933 7318 7963 7332
rect 7991 7318 8004 7356
rect 8076 7362 8111 7370
rect 8076 7336 8077 7362
rect 8084 7336 8111 7362
rect 8019 7318 8049 7332
rect 8076 7328 8111 7336
rect 8113 7362 8154 7370
rect 8113 7336 8128 7362
rect 8135 7336 8154 7362
rect 8218 7358 8280 7370
rect 8292 7358 8367 7370
rect 8425 7358 8500 7370
rect 8512 7358 8543 7370
rect 8549 7358 8584 7370
rect 8218 7356 8380 7358
rect 8113 7328 8154 7336
rect 8236 7332 8249 7356
rect 8264 7354 8279 7356
rect 8076 7318 8077 7328
rect 8092 7318 8105 7328
rect 8119 7318 8120 7328
rect 8135 7318 8148 7328
rect 8163 7318 8193 7332
rect 8236 7318 8279 7332
rect 8303 7329 8310 7336
rect 8313 7332 8380 7356
rect 8412 7356 8584 7358
rect 8382 7334 8410 7338
rect 8412 7334 8492 7356
rect 8513 7354 8528 7356
rect 8382 7332 8492 7334
rect 8313 7328 8492 7332
rect 8286 7318 8316 7328
rect 8318 7318 8471 7328
rect 8479 7318 8509 7328
rect 8513 7318 8543 7332
rect 8571 7318 8584 7356
rect 8656 7362 8691 7370
rect 8656 7336 8657 7362
rect 8664 7336 8691 7362
rect 8599 7318 8629 7332
rect 8656 7328 8691 7336
rect 8693 7362 8734 7370
rect 8693 7336 8708 7362
rect 8715 7336 8734 7362
rect 8798 7358 8860 7370
rect 8872 7358 8947 7370
rect 9005 7358 9080 7370
rect 9092 7358 9123 7370
rect 9129 7358 9164 7370
rect 8798 7356 8960 7358
rect 8693 7328 8734 7336
rect 8816 7332 8829 7356
rect 8844 7354 8859 7356
rect 8656 7318 8657 7328
rect 8672 7318 8685 7328
rect 8699 7318 8700 7328
rect 8715 7318 8728 7328
rect 8743 7318 8773 7332
rect 8816 7318 8859 7332
rect 8883 7329 8890 7336
rect 8893 7332 8960 7356
rect 8992 7356 9164 7358
rect 8962 7334 8990 7338
rect 8992 7334 9072 7356
rect 9093 7354 9108 7356
rect 8962 7332 9072 7334
rect 8893 7328 9072 7332
rect 8866 7318 8896 7328
rect 8898 7318 9051 7328
rect 9059 7318 9089 7328
rect 9093 7318 9123 7332
rect 9151 7318 9164 7356
rect 9236 7362 9271 7370
rect 9236 7336 9237 7362
rect 9244 7336 9271 7362
rect 9179 7318 9209 7332
rect 9236 7328 9271 7336
rect 9236 7318 9237 7328
rect 9252 7318 9265 7328
rect -1 7312 9265 7318
rect 0 7304 9265 7312
rect 15 7274 28 7304
rect 43 7286 73 7304
rect 116 7290 130 7304
rect 166 7290 386 7304
rect 117 7288 130 7290
rect 83 7276 98 7288
rect 80 7274 102 7276
rect 107 7274 137 7288
rect 198 7286 351 7290
rect 180 7274 372 7286
rect 415 7274 445 7288
rect 451 7274 464 7304
rect 479 7286 509 7304
rect 552 7274 565 7304
rect 595 7274 608 7304
rect 623 7286 653 7304
rect 696 7290 710 7304
rect 746 7290 966 7304
rect 697 7288 710 7290
rect 663 7276 678 7288
rect 660 7274 682 7276
rect 687 7274 717 7288
rect 778 7286 931 7290
rect 760 7274 952 7286
rect 995 7274 1025 7288
rect 1031 7274 1044 7304
rect 1059 7286 1089 7304
rect 1132 7274 1145 7304
rect 1175 7274 1188 7304
rect 1203 7286 1233 7304
rect 1276 7290 1290 7304
rect 1326 7290 1546 7304
rect 1277 7288 1290 7290
rect 1243 7276 1258 7288
rect 1240 7274 1262 7276
rect 1267 7274 1297 7288
rect 1358 7286 1511 7290
rect 1340 7274 1532 7286
rect 1575 7274 1605 7288
rect 1611 7274 1624 7304
rect 1639 7286 1669 7304
rect 1712 7274 1725 7304
rect 1755 7274 1768 7304
rect 1783 7286 1813 7304
rect 1856 7290 1870 7304
rect 1906 7290 2126 7304
rect 1857 7288 1870 7290
rect 1823 7276 1838 7288
rect 1820 7274 1842 7276
rect 1847 7274 1877 7288
rect 1938 7286 2091 7290
rect 1920 7274 2112 7286
rect 2155 7274 2185 7288
rect 2191 7274 2204 7304
rect 2219 7286 2249 7304
rect 2292 7274 2305 7304
rect 2335 7274 2348 7304
rect 2363 7286 2393 7304
rect 2436 7290 2450 7304
rect 2486 7290 2706 7304
rect 2437 7288 2450 7290
rect 2403 7276 2418 7288
rect 2400 7274 2422 7276
rect 2427 7274 2457 7288
rect 2518 7286 2671 7290
rect 2500 7274 2692 7286
rect 2735 7274 2765 7288
rect 2771 7274 2784 7304
rect 2799 7286 2829 7304
rect 2872 7274 2885 7304
rect 2915 7274 2928 7304
rect 2943 7286 2973 7304
rect 3016 7290 3030 7304
rect 3066 7290 3286 7304
rect 3017 7288 3030 7290
rect 2983 7276 2998 7288
rect 2980 7274 3002 7276
rect 3007 7274 3037 7288
rect 3098 7286 3251 7290
rect 3080 7274 3272 7286
rect 3315 7274 3345 7288
rect 3351 7274 3364 7304
rect 3379 7286 3409 7304
rect 3452 7274 3465 7304
rect 3495 7274 3508 7304
rect 3523 7286 3553 7304
rect 3596 7290 3610 7304
rect 3646 7290 3866 7304
rect 3597 7288 3610 7290
rect 3563 7276 3578 7288
rect 3560 7274 3582 7276
rect 3587 7274 3617 7288
rect 3678 7286 3831 7290
rect 3660 7274 3852 7286
rect 3895 7274 3925 7288
rect 3931 7274 3944 7304
rect 3959 7286 3989 7304
rect 4032 7274 4045 7304
rect 4075 7274 4088 7304
rect 4103 7286 4133 7304
rect 4176 7290 4190 7304
rect 4226 7290 4446 7304
rect 4177 7288 4190 7290
rect 4143 7276 4158 7288
rect 4140 7274 4162 7276
rect 4167 7274 4197 7288
rect 4258 7286 4411 7290
rect 4240 7274 4432 7286
rect 4475 7274 4505 7288
rect 4511 7274 4524 7304
rect 4539 7286 4569 7304
rect 4612 7274 4625 7304
rect 4655 7274 4668 7304
rect 4683 7286 4713 7304
rect 4756 7290 4770 7304
rect 4806 7290 5026 7304
rect 4757 7288 4770 7290
rect 4723 7276 4738 7288
rect 4720 7274 4742 7276
rect 4747 7274 4777 7288
rect 4838 7286 4991 7290
rect 4820 7274 5012 7286
rect 5055 7274 5085 7288
rect 5091 7274 5104 7304
rect 5119 7286 5149 7304
rect 5192 7274 5205 7304
rect 5235 7274 5248 7304
rect 5263 7286 5293 7304
rect 5336 7290 5350 7304
rect 5386 7290 5606 7304
rect 5337 7288 5350 7290
rect 5303 7276 5318 7288
rect 5300 7274 5322 7276
rect 5327 7274 5357 7288
rect 5418 7286 5571 7290
rect 5400 7274 5592 7286
rect 5635 7274 5665 7288
rect 5671 7274 5684 7304
rect 5699 7286 5729 7304
rect 5772 7274 5785 7304
rect 5815 7274 5828 7304
rect 5843 7286 5873 7304
rect 5916 7290 5930 7304
rect 5966 7290 6186 7304
rect 5917 7288 5930 7290
rect 5883 7276 5898 7288
rect 5880 7274 5902 7276
rect 5907 7274 5937 7288
rect 5998 7286 6151 7290
rect 5980 7274 6172 7286
rect 6215 7274 6245 7288
rect 6251 7274 6264 7304
rect 6279 7286 6309 7304
rect 6352 7274 6365 7304
rect 6395 7274 6408 7304
rect 6423 7286 6453 7304
rect 6496 7290 6510 7304
rect 6546 7290 6766 7304
rect 6497 7288 6510 7290
rect 6463 7276 6478 7288
rect 6460 7274 6482 7276
rect 6487 7274 6517 7288
rect 6578 7286 6731 7290
rect 6560 7274 6752 7286
rect 6795 7274 6825 7288
rect 6831 7274 6844 7304
rect 6859 7286 6889 7304
rect 6932 7274 6945 7304
rect 6975 7274 6988 7304
rect 7003 7286 7033 7304
rect 7076 7290 7090 7304
rect 7126 7290 7346 7304
rect 7077 7288 7090 7290
rect 7043 7276 7058 7288
rect 7040 7274 7062 7276
rect 7067 7274 7097 7288
rect 7158 7286 7311 7290
rect 7140 7274 7332 7286
rect 7375 7274 7405 7288
rect 7411 7274 7424 7304
rect 7439 7286 7469 7304
rect 7512 7274 7525 7304
rect 7555 7274 7568 7304
rect 7583 7286 7613 7304
rect 7656 7290 7670 7304
rect 7706 7290 7926 7304
rect 7657 7288 7670 7290
rect 7623 7276 7638 7288
rect 7620 7274 7642 7276
rect 7647 7274 7677 7288
rect 7738 7286 7891 7290
rect 7720 7274 7912 7286
rect 7955 7274 7985 7288
rect 7991 7274 8004 7304
rect 8019 7286 8049 7304
rect 8092 7274 8105 7304
rect 8135 7274 8148 7304
rect 8163 7286 8193 7304
rect 8236 7290 8250 7304
rect 8286 7290 8506 7304
rect 8237 7288 8250 7290
rect 8203 7276 8218 7288
rect 8200 7274 8222 7276
rect 8227 7274 8257 7288
rect 8318 7286 8471 7290
rect 8300 7274 8492 7286
rect 8535 7274 8565 7288
rect 8571 7274 8584 7304
rect 8599 7286 8629 7304
rect 8672 7274 8685 7304
rect 8715 7274 8728 7304
rect 8743 7286 8773 7304
rect 8816 7290 8830 7304
rect 8866 7290 9086 7304
rect 8817 7288 8830 7290
rect 8783 7276 8798 7288
rect 8780 7274 8802 7276
rect 8807 7274 8837 7288
rect 8898 7286 9051 7290
rect 8880 7274 9072 7286
rect 9115 7274 9145 7288
rect 9151 7274 9164 7304
rect 9179 7286 9209 7304
rect 9252 7274 9265 7304
rect 0 7260 9265 7274
rect 15 7156 28 7260
rect 73 7238 74 7248
rect 89 7238 102 7248
rect 73 7234 102 7238
rect 107 7234 137 7260
rect 155 7246 171 7248
rect 243 7246 296 7260
rect 244 7244 308 7246
rect 351 7244 366 7260
rect 415 7257 445 7260
rect 415 7254 451 7257
rect 381 7246 397 7248
rect 155 7234 170 7238
rect 73 7232 170 7234
rect 198 7232 366 7244
rect 382 7234 397 7238
rect 415 7235 454 7254
rect 473 7248 480 7249
rect 479 7241 480 7248
rect 463 7238 464 7241
rect 479 7238 492 7241
rect 415 7234 445 7235
rect 454 7234 460 7235
rect 463 7234 492 7238
rect 382 7233 492 7234
rect 382 7232 498 7233
rect 57 7224 108 7232
rect 57 7212 82 7224
rect 89 7212 108 7224
rect 139 7224 189 7232
rect 139 7216 155 7224
rect 162 7222 189 7224
rect 198 7222 419 7232
rect 162 7212 419 7222
rect 448 7224 498 7232
rect 448 7215 464 7224
rect 57 7204 108 7212
rect 155 7204 419 7212
rect 445 7212 464 7215
rect 471 7212 498 7224
rect 445 7204 498 7212
rect 73 7196 74 7204
rect 89 7196 102 7204
rect 73 7188 89 7196
rect 70 7181 89 7184
rect 70 7172 92 7181
rect 43 7162 92 7172
rect 43 7156 73 7162
rect 92 7157 97 7162
rect 15 7140 89 7156
rect 107 7148 137 7204
rect 172 7194 380 7204
rect 415 7200 460 7204
rect 463 7203 464 7204
rect 479 7203 492 7204
rect 198 7164 387 7194
rect 213 7161 387 7164
rect 206 7158 387 7161
rect 15 7138 28 7140
rect 43 7138 77 7140
rect 15 7122 89 7138
rect 116 7134 129 7148
rect 144 7134 160 7150
rect 206 7145 217 7158
rect -1 7100 0 7116
rect 15 7100 28 7122
rect 43 7100 73 7122
rect 116 7118 178 7134
rect 206 7127 217 7143
rect 222 7138 232 7158
rect 242 7138 256 7158
rect 259 7145 268 7158
rect 284 7145 293 7158
rect 222 7127 256 7138
rect 259 7127 268 7143
rect 284 7127 293 7143
rect 300 7138 310 7158
rect 320 7138 334 7158
rect 335 7145 346 7158
rect 300 7127 334 7138
rect 335 7127 346 7143
rect 392 7134 408 7150
rect 415 7148 445 7200
rect 479 7196 480 7203
rect 464 7188 480 7196
rect 451 7156 464 7175
rect 479 7156 509 7172
rect 451 7140 525 7156
rect 451 7138 464 7140
rect 479 7138 513 7140
rect 116 7116 129 7118
rect 144 7116 178 7118
rect 116 7100 178 7116
rect 222 7111 238 7114
rect 300 7111 330 7122
rect 378 7118 424 7134
rect 451 7122 525 7138
rect 378 7116 412 7118
rect 377 7100 424 7116
rect 451 7100 464 7122
rect 479 7100 509 7122
rect 536 7100 537 7116
rect 552 7100 565 7260
rect 595 7156 608 7260
rect 653 7238 654 7248
rect 669 7238 682 7248
rect 653 7234 682 7238
rect 687 7234 717 7260
rect 735 7246 751 7248
rect 823 7246 876 7260
rect 824 7244 888 7246
rect 931 7244 946 7260
rect 995 7257 1025 7260
rect 995 7254 1031 7257
rect 961 7246 977 7248
rect 735 7234 750 7238
rect 653 7232 750 7234
rect 778 7232 946 7244
rect 962 7234 977 7238
rect 995 7235 1034 7254
rect 1053 7248 1060 7249
rect 1059 7241 1060 7248
rect 1043 7238 1044 7241
rect 1059 7238 1072 7241
rect 995 7234 1025 7235
rect 1034 7234 1040 7235
rect 1043 7234 1072 7238
rect 962 7233 1072 7234
rect 962 7232 1078 7233
rect 637 7224 688 7232
rect 637 7212 662 7224
rect 669 7212 688 7224
rect 719 7224 769 7232
rect 719 7216 735 7224
rect 742 7222 769 7224
rect 778 7222 999 7232
rect 742 7212 999 7222
rect 1028 7224 1078 7232
rect 1028 7215 1044 7224
rect 637 7204 688 7212
rect 735 7204 999 7212
rect 1025 7212 1044 7215
rect 1051 7212 1078 7224
rect 1025 7204 1078 7212
rect 653 7196 654 7204
rect 669 7196 682 7204
rect 653 7188 669 7196
rect 650 7181 669 7184
rect 650 7172 672 7181
rect 623 7162 672 7172
rect 623 7156 653 7162
rect 672 7157 677 7162
rect 595 7140 669 7156
rect 687 7148 717 7204
rect 752 7194 960 7204
rect 995 7200 1040 7204
rect 1043 7203 1044 7204
rect 1059 7203 1072 7204
rect 778 7164 967 7194
rect 793 7161 967 7164
rect 786 7158 967 7161
rect 595 7138 608 7140
rect 623 7138 657 7140
rect 595 7122 669 7138
rect 696 7134 709 7148
rect 724 7134 740 7150
rect 786 7145 797 7158
rect 579 7100 580 7116
rect 595 7100 608 7122
rect 623 7100 653 7122
rect 696 7118 758 7134
rect 786 7127 797 7143
rect 802 7138 812 7158
rect 822 7138 836 7158
rect 839 7145 848 7158
rect 864 7145 873 7158
rect 802 7127 836 7138
rect 839 7127 848 7143
rect 864 7127 873 7143
rect 880 7138 890 7158
rect 900 7138 914 7158
rect 915 7145 926 7158
rect 880 7127 914 7138
rect 915 7127 926 7143
rect 972 7134 988 7150
rect 995 7148 1025 7200
rect 1059 7196 1060 7203
rect 1044 7188 1060 7196
rect 1031 7156 1044 7175
rect 1059 7156 1089 7172
rect 1031 7140 1105 7156
rect 1031 7138 1044 7140
rect 1059 7138 1093 7140
rect 696 7116 709 7118
rect 724 7116 758 7118
rect 696 7100 758 7116
rect 802 7111 818 7114
rect 880 7111 910 7122
rect 958 7118 1004 7134
rect 1031 7122 1105 7138
rect 958 7116 992 7118
rect 957 7100 1004 7116
rect 1031 7100 1044 7122
rect 1059 7100 1089 7122
rect 1116 7100 1117 7116
rect 1132 7100 1145 7260
rect 1175 7156 1188 7260
rect 1233 7238 1234 7248
rect 1249 7238 1262 7248
rect 1233 7234 1262 7238
rect 1267 7234 1297 7260
rect 1315 7246 1331 7248
rect 1403 7246 1456 7260
rect 1404 7244 1468 7246
rect 1511 7244 1526 7260
rect 1575 7257 1605 7260
rect 1575 7254 1611 7257
rect 1541 7246 1557 7248
rect 1315 7234 1330 7238
rect 1233 7232 1330 7234
rect 1358 7232 1526 7244
rect 1542 7234 1557 7238
rect 1575 7235 1614 7254
rect 1633 7248 1640 7249
rect 1639 7241 1640 7248
rect 1623 7238 1624 7241
rect 1639 7238 1652 7241
rect 1575 7234 1605 7235
rect 1614 7234 1620 7235
rect 1623 7234 1652 7238
rect 1542 7233 1652 7234
rect 1542 7232 1658 7233
rect 1217 7224 1268 7232
rect 1217 7212 1242 7224
rect 1249 7212 1268 7224
rect 1299 7224 1349 7232
rect 1299 7216 1315 7224
rect 1322 7222 1349 7224
rect 1358 7222 1579 7232
rect 1322 7212 1579 7222
rect 1608 7224 1658 7232
rect 1608 7215 1624 7224
rect 1217 7204 1268 7212
rect 1315 7204 1579 7212
rect 1605 7212 1624 7215
rect 1631 7212 1658 7224
rect 1605 7204 1658 7212
rect 1233 7196 1234 7204
rect 1249 7196 1262 7204
rect 1233 7188 1249 7196
rect 1230 7181 1249 7184
rect 1230 7172 1252 7181
rect 1203 7162 1252 7172
rect 1203 7156 1233 7162
rect 1252 7157 1257 7162
rect 1175 7140 1249 7156
rect 1267 7148 1297 7204
rect 1332 7194 1540 7204
rect 1575 7200 1620 7204
rect 1623 7203 1624 7204
rect 1639 7203 1652 7204
rect 1358 7164 1547 7194
rect 1373 7161 1547 7164
rect 1366 7158 1547 7161
rect 1175 7138 1188 7140
rect 1203 7138 1237 7140
rect 1175 7122 1249 7138
rect 1276 7134 1289 7148
rect 1304 7134 1320 7150
rect 1366 7145 1377 7158
rect 1159 7100 1160 7116
rect 1175 7100 1188 7122
rect 1203 7100 1233 7122
rect 1276 7118 1338 7134
rect 1366 7127 1377 7143
rect 1382 7138 1392 7158
rect 1402 7138 1416 7158
rect 1419 7145 1428 7158
rect 1444 7145 1453 7158
rect 1382 7127 1416 7138
rect 1419 7127 1428 7143
rect 1444 7127 1453 7143
rect 1460 7138 1470 7158
rect 1480 7138 1494 7158
rect 1495 7145 1506 7158
rect 1460 7127 1494 7138
rect 1495 7127 1506 7143
rect 1552 7134 1568 7150
rect 1575 7148 1605 7200
rect 1639 7196 1640 7203
rect 1624 7188 1640 7196
rect 1611 7156 1624 7175
rect 1639 7156 1669 7172
rect 1611 7140 1685 7156
rect 1611 7138 1624 7140
rect 1639 7138 1673 7140
rect 1276 7116 1289 7118
rect 1304 7116 1338 7118
rect 1276 7100 1338 7116
rect 1382 7111 1398 7114
rect 1460 7111 1490 7122
rect 1538 7118 1584 7134
rect 1611 7122 1685 7138
rect 1538 7116 1572 7118
rect 1537 7100 1584 7116
rect 1611 7100 1624 7122
rect 1639 7100 1669 7122
rect 1696 7100 1697 7116
rect 1712 7100 1725 7260
rect 1755 7156 1768 7260
rect 1813 7238 1814 7248
rect 1829 7238 1842 7248
rect 1813 7234 1842 7238
rect 1847 7234 1877 7260
rect 1895 7246 1911 7248
rect 1983 7246 2036 7260
rect 1984 7244 2048 7246
rect 2091 7244 2106 7260
rect 2155 7257 2185 7260
rect 2155 7254 2191 7257
rect 2121 7246 2137 7248
rect 1895 7234 1910 7238
rect 1813 7232 1910 7234
rect 1938 7232 2106 7244
rect 2122 7234 2137 7238
rect 2155 7235 2194 7254
rect 2213 7248 2220 7249
rect 2219 7241 2220 7248
rect 2203 7238 2204 7241
rect 2219 7238 2232 7241
rect 2155 7234 2185 7235
rect 2194 7234 2200 7235
rect 2203 7234 2232 7238
rect 2122 7233 2232 7234
rect 2122 7232 2238 7233
rect 1797 7224 1848 7232
rect 1797 7212 1822 7224
rect 1829 7212 1848 7224
rect 1879 7224 1929 7232
rect 1879 7216 1895 7224
rect 1902 7222 1929 7224
rect 1938 7222 2159 7232
rect 1902 7212 2159 7222
rect 2188 7224 2238 7232
rect 2188 7215 2204 7224
rect 1797 7204 1848 7212
rect 1895 7204 2159 7212
rect 2185 7212 2204 7215
rect 2211 7212 2238 7224
rect 2185 7204 2238 7212
rect 1813 7196 1814 7204
rect 1829 7196 1842 7204
rect 1813 7188 1829 7196
rect 1810 7181 1829 7184
rect 1810 7172 1832 7181
rect 1783 7162 1832 7172
rect 1783 7156 1813 7162
rect 1832 7157 1837 7162
rect 1755 7140 1829 7156
rect 1847 7148 1877 7204
rect 1912 7194 2120 7204
rect 2155 7200 2200 7204
rect 2203 7203 2204 7204
rect 2219 7203 2232 7204
rect 1938 7164 2127 7194
rect 1953 7161 2127 7164
rect 1946 7158 2127 7161
rect 1755 7138 1768 7140
rect 1783 7138 1817 7140
rect 1755 7122 1829 7138
rect 1856 7134 1869 7148
rect 1884 7134 1900 7150
rect 1946 7145 1957 7158
rect 1739 7100 1740 7116
rect 1755 7100 1768 7122
rect 1783 7100 1813 7122
rect 1856 7118 1918 7134
rect 1946 7127 1957 7143
rect 1962 7138 1972 7158
rect 1982 7138 1996 7158
rect 1999 7145 2008 7158
rect 2024 7145 2033 7158
rect 1962 7127 1996 7138
rect 1999 7127 2008 7143
rect 2024 7127 2033 7143
rect 2040 7138 2050 7158
rect 2060 7138 2074 7158
rect 2075 7145 2086 7158
rect 2040 7127 2074 7138
rect 2075 7127 2086 7143
rect 2132 7134 2148 7150
rect 2155 7148 2185 7200
rect 2219 7196 2220 7203
rect 2204 7188 2220 7196
rect 2191 7156 2204 7175
rect 2219 7156 2249 7172
rect 2191 7140 2265 7156
rect 2191 7138 2204 7140
rect 2219 7138 2253 7140
rect 1856 7116 1869 7118
rect 1884 7116 1918 7118
rect 1856 7100 1918 7116
rect 1962 7111 1976 7114
rect 2040 7111 2070 7122
rect 2118 7118 2164 7134
rect 2191 7122 2265 7138
rect 2118 7116 2152 7118
rect 2117 7100 2164 7116
rect 2191 7100 2204 7122
rect 2219 7100 2249 7122
rect 2276 7100 2277 7116
rect 2292 7100 2305 7260
rect 2335 7156 2348 7260
rect 2393 7238 2394 7248
rect 2409 7238 2422 7248
rect 2393 7234 2422 7238
rect 2427 7234 2457 7260
rect 2475 7246 2491 7248
rect 2563 7246 2616 7260
rect 2564 7244 2628 7246
rect 2671 7244 2686 7260
rect 2735 7257 2765 7260
rect 2735 7254 2771 7257
rect 2701 7246 2717 7248
rect 2475 7234 2490 7238
rect 2393 7232 2490 7234
rect 2518 7232 2686 7244
rect 2702 7234 2717 7238
rect 2735 7235 2774 7254
rect 2793 7248 2800 7249
rect 2799 7241 2800 7248
rect 2783 7238 2784 7241
rect 2799 7238 2812 7241
rect 2735 7234 2765 7235
rect 2774 7234 2780 7235
rect 2783 7234 2812 7238
rect 2702 7233 2812 7234
rect 2702 7232 2818 7233
rect 2377 7224 2428 7232
rect 2377 7212 2402 7224
rect 2409 7212 2428 7224
rect 2459 7224 2509 7232
rect 2459 7216 2475 7224
rect 2482 7222 2509 7224
rect 2518 7222 2739 7232
rect 2482 7212 2739 7222
rect 2768 7224 2818 7232
rect 2768 7215 2784 7224
rect 2377 7204 2428 7212
rect 2475 7204 2739 7212
rect 2765 7212 2784 7215
rect 2791 7212 2818 7224
rect 2765 7204 2818 7212
rect 2393 7196 2394 7204
rect 2409 7196 2422 7204
rect 2393 7188 2409 7196
rect 2390 7181 2409 7184
rect 2390 7172 2412 7181
rect 2363 7162 2412 7172
rect 2363 7156 2393 7162
rect 2412 7157 2417 7162
rect 2335 7140 2409 7156
rect 2427 7148 2457 7204
rect 2492 7194 2700 7204
rect 2735 7200 2780 7204
rect 2783 7203 2784 7204
rect 2799 7203 2812 7204
rect 2518 7164 2707 7194
rect 2533 7161 2707 7164
rect 2526 7158 2707 7161
rect 2335 7138 2348 7140
rect 2363 7138 2397 7140
rect 2335 7122 2409 7138
rect 2436 7134 2449 7148
rect 2464 7134 2480 7150
rect 2526 7145 2537 7158
rect 2319 7100 2320 7116
rect 2335 7100 2348 7122
rect 2363 7100 2393 7122
rect 2436 7118 2498 7134
rect 2526 7127 2537 7143
rect 2542 7138 2552 7158
rect 2562 7138 2576 7158
rect 2579 7145 2588 7158
rect 2604 7145 2613 7158
rect 2542 7127 2576 7138
rect 2579 7127 2588 7143
rect 2604 7127 2613 7143
rect 2620 7138 2630 7158
rect 2640 7138 2654 7158
rect 2655 7145 2666 7158
rect 2620 7127 2654 7138
rect 2655 7127 2666 7143
rect 2712 7134 2728 7150
rect 2735 7148 2765 7200
rect 2799 7196 2800 7203
rect 2784 7188 2800 7196
rect 2771 7156 2784 7175
rect 2799 7156 2829 7172
rect 2771 7140 2845 7156
rect 2771 7138 2784 7140
rect 2799 7138 2833 7140
rect 2436 7116 2449 7118
rect 2464 7116 2498 7118
rect 2436 7100 2498 7116
rect 2542 7111 2558 7114
rect 2620 7111 2650 7122
rect 2698 7118 2744 7134
rect 2771 7122 2845 7138
rect 2698 7116 2732 7118
rect 2697 7100 2744 7116
rect 2771 7100 2784 7122
rect 2799 7100 2829 7122
rect 2856 7100 2857 7116
rect 2872 7100 2885 7260
rect 2915 7156 2928 7260
rect 2973 7238 2974 7248
rect 2989 7238 3002 7248
rect 2973 7234 3002 7238
rect 3007 7234 3037 7260
rect 3055 7246 3071 7248
rect 3143 7246 3196 7260
rect 3144 7244 3208 7246
rect 3251 7244 3266 7260
rect 3315 7257 3345 7260
rect 3315 7254 3351 7257
rect 3281 7246 3297 7248
rect 3055 7234 3070 7238
rect 2973 7232 3070 7234
rect 3098 7232 3266 7244
rect 3282 7234 3297 7238
rect 3315 7235 3354 7254
rect 3373 7248 3380 7249
rect 3379 7241 3380 7248
rect 3363 7238 3364 7241
rect 3379 7238 3392 7241
rect 3315 7234 3345 7235
rect 3354 7234 3360 7235
rect 3363 7234 3392 7238
rect 3282 7233 3392 7234
rect 3282 7232 3398 7233
rect 2957 7224 3008 7232
rect 2957 7212 2982 7224
rect 2989 7212 3008 7224
rect 3039 7224 3089 7232
rect 3039 7216 3055 7224
rect 3062 7222 3089 7224
rect 3098 7222 3319 7232
rect 3062 7212 3319 7222
rect 3348 7224 3398 7232
rect 3348 7215 3364 7224
rect 2957 7204 3008 7212
rect 3055 7204 3319 7212
rect 3345 7212 3364 7215
rect 3371 7212 3398 7224
rect 3345 7204 3398 7212
rect 2973 7196 2974 7204
rect 2989 7196 3002 7204
rect 2973 7188 2989 7196
rect 2970 7181 2989 7184
rect 2970 7172 2992 7181
rect 2943 7162 2992 7172
rect 2943 7156 2973 7162
rect 2992 7157 2997 7162
rect 2915 7140 2989 7156
rect 3007 7148 3037 7204
rect 3072 7194 3280 7204
rect 3315 7200 3360 7204
rect 3363 7203 3364 7204
rect 3379 7203 3392 7204
rect 3098 7164 3287 7194
rect 3113 7161 3287 7164
rect 3106 7158 3287 7161
rect 2915 7138 2928 7140
rect 2943 7138 2977 7140
rect 2915 7122 2989 7138
rect 3016 7134 3029 7148
rect 3044 7134 3060 7150
rect 3106 7145 3117 7158
rect 2899 7100 2900 7116
rect 2915 7100 2928 7122
rect 2943 7100 2973 7122
rect 3016 7118 3078 7134
rect 3106 7127 3117 7143
rect 3122 7138 3132 7158
rect 3142 7138 3156 7158
rect 3159 7145 3168 7158
rect 3184 7145 3193 7158
rect 3122 7127 3156 7138
rect 3159 7127 3168 7143
rect 3184 7127 3193 7143
rect 3200 7138 3210 7158
rect 3220 7138 3234 7158
rect 3235 7145 3246 7158
rect 3200 7127 3234 7138
rect 3235 7127 3246 7143
rect 3292 7134 3308 7150
rect 3315 7148 3345 7200
rect 3379 7196 3380 7203
rect 3364 7188 3380 7196
rect 3351 7156 3364 7175
rect 3379 7156 3409 7172
rect 3351 7140 3425 7156
rect 3351 7138 3364 7140
rect 3379 7138 3413 7140
rect 3016 7116 3029 7118
rect 3044 7116 3078 7118
rect 3016 7100 3078 7116
rect 3122 7111 3138 7114
rect 3200 7111 3230 7122
rect 3278 7118 3324 7134
rect 3351 7122 3425 7138
rect 3278 7116 3312 7118
rect 3277 7100 3324 7116
rect 3351 7100 3364 7122
rect 3379 7100 3409 7122
rect 3436 7100 3437 7116
rect 3452 7100 3465 7260
rect 3495 7156 3508 7260
rect 3553 7238 3554 7248
rect 3569 7238 3582 7248
rect 3553 7234 3582 7238
rect 3587 7234 3617 7260
rect 3635 7246 3651 7248
rect 3723 7246 3776 7260
rect 3724 7244 3788 7246
rect 3831 7244 3846 7260
rect 3895 7257 3925 7260
rect 3895 7254 3931 7257
rect 3861 7246 3877 7248
rect 3635 7234 3650 7238
rect 3553 7232 3650 7234
rect 3678 7232 3846 7244
rect 3862 7234 3877 7238
rect 3895 7235 3934 7254
rect 3953 7248 3960 7249
rect 3959 7241 3960 7248
rect 3943 7238 3944 7241
rect 3959 7238 3972 7241
rect 3895 7234 3925 7235
rect 3934 7234 3940 7235
rect 3943 7234 3972 7238
rect 3862 7233 3972 7234
rect 3862 7232 3978 7233
rect 3537 7224 3588 7232
rect 3537 7212 3562 7224
rect 3569 7212 3588 7224
rect 3619 7224 3669 7232
rect 3619 7216 3635 7224
rect 3642 7222 3669 7224
rect 3678 7222 3899 7232
rect 3642 7212 3899 7222
rect 3928 7224 3978 7232
rect 3928 7215 3944 7224
rect 3537 7204 3588 7212
rect 3635 7204 3899 7212
rect 3925 7212 3944 7215
rect 3951 7212 3978 7224
rect 3925 7204 3978 7212
rect 3553 7196 3554 7204
rect 3569 7196 3582 7204
rect 3553 7188 3569 7196
rect 3550 7181 3569 7184
rect 3550 7172 3572 7181
rect 3523 7162 3572 7172
rect 3523 7156 3553 7162
rect 3572 7157 3577 7162
rect 3495 7140 3569 7156
rect 3587 7148 3617 7204
rect 3652 7194 3860 7204
rect 3895 7200 3940 7204
rect 3943 7203 3944 7204
rect 3959 7203 3972 7204
rect 3678 7164 3867 7194
rect 3693 7161 3867 7164
rect 3686 7158 3867 7161
rect 3495 7138 3508 7140
rect 3523 7138 3557 7140
rect 3495 7122 3569 7138
rect 3596 7134 3609 7148
rect 3624 7134 3640 7150
rect 3686 7145 3697 7158
rect 3479 7100 3480 7116
rect 3495 7100 3508 7122
rect 3523 7100 3553 7122
rect 3596 7118 3658 7134
rect 3686 7127 3697 7143
rect 3702 7138 3712 7158
rect 3722 7138 3736 7158
rect 3739 7145 3748 7158
rect 3764 7145 3773 7158
rect 3702 7127 3736 7138
rect 3739 7127 3748 7143
rect 3764 7127 3773 7143
rect 3780 7138 3790 7158
rect 3800 7138 3814 7158
rect 3815 7145 3826 7158
rect 3780 7127 3814 7138
rect 3815 7127 3826 7143
rect 3872 7134 3888 7150
rect 3895 7148 3925 7200
rect 3959 7196 3960 7203
rect 3944 7188 3960 7196
rect 3931 7156 3944 7175
rect 3959 7156 3989 7172
rect 3931 7140 4005 7156
rect 3931 7138 3944 7140
rect 3959 7138 3993 7140
rect 3596 7116 3609 7118
rect 3624 7116 3658 7118
rect 3596 7100 3658 7116
rect 3702 7111 3718 7114
rect 3780 7111 3810 7122
rect 3858 7118 3904 7134
rect 3931 7122 4005 7138
rect 3858 7116 3892 7118
rect 3857 7100 3904 7116
rect 3931 7100 3944 7122
rect 3959 7100 3989 7122
rect 4016 7100 4017 7116
rect 4032 7100 4045 7260
rect 4075 7156 4088 7260
rect 4133 7238 4134 7248
rect 4149 7238 4162 7248
rect 4133 7234 4162 7238
rect 4167 7234 4197 7260
rect 4215 7246 4231 7248
rect 4303 7246 4356 7260
rect 4304 7244 4368 7246
rect 4411 7244 4426 7260
rect 4475 7257 4505 7260
rect 4475 7254 4511 7257
rect 4441 7246 4457 7248
rect 4215 7234 4230 7238
rect 4133 7232 4230 7234
rect 4258 7232 4426 7244
rect 4442 7234 4457 7238
rect 4475 7235 4514 7254
rect 4533 7248 4540 7249
rect 4539 7241 4540 7248
rect 4523 7238 4524 7241
rect 4539 7238 4552 7241
rect 4475 7234 4505 7235
rect 4514 7234 4520 7235
rect 4523 7234 4552 7238
rect 4442 7233 4552 7234
rect 4442 7232 4558 7233
rect 4117 7224 4168 7232
rect 4117 7212 4142 7224
rect 4149 7212 4168 7224
rect 4199 7224 4249 7232
rect 4199 7216 4215 7224
rect 4222 7222 4249 7224
rect 4258 7222 4479 7232
rect 4222 7212 4479 7222
rect 4508 7224 4558 7232
rect 4508 7215 4524 7224
rect 4117 7204 4168 7212
rect 4215 7204 4479 7212
rect 4505 7212 4524 7215
rect 4531 7212 4558 7224
rect 4505 7204 4558 7212
rect 4133 7196 4134 7204
rect 4149 7196 4162 7204
rect 4133 7188 4149 7196
rect 4130 7181 4149 7184
rect 4130 7172 4152 7181
rect 4103 7162 4152 7172
rect 4103 7156 4133 7162
rect 4152 7157 4157 7162
rect 4075 7140 4149 7156
rect 4167 7148 4197 7204
rect 4232 7194 4440 7204
rect 4475 7200 4520 7204
rect 4523 7203 4524 7204
rect 4539 7203 4552 7204
rect 4258 7164 4447 7194
rect 4273 7161 4447 7164
rect 4266 7158 4447 7161
rect 4075 7138 4088 7140
rect 4103 7138 4137 7140
rect 4075 7122 4149 7138
rect 4176 7134 4189 7148
rect 4204 7134 4220 7150
rect 4266 7145 4277 7158
rect 4059 7100 4060 7116
rect 4075 7100 4088 7122
rect 4103 7100 4133 7122
rect 4176 7118 4238 7134
rect 4266 7127 4277 7143
rect 4282 7138 4292 7158
rect 4302 7138 4316 7158
rect 4319 7145 4328 7158
rect 4344 7145 4353 7158
rect 4282 7127 4316 7138
rect 4319 7127 4328 7143
rect 4344 7127 4353 7143
rect 4360 7138 4370 7158
rect 4380 7138 4394 7158
rect 4395 7145 4406 7158
rect 4360 7127 4394 7138
rect 4395 7127 4406 7143
rect 4452 7134 4468 7150
rect 4475 7148 4505 7200
rect 4539 7196 4540 7203
rect 4524 7188 4540 7196
rect 4511 7156 4524 7175
rect 4539 7156 4569 7172
rect 4511 7140 4585 7156
rect 4511 7138 4524 7140
rect 4539 7138 4573 7140
rect 4176 7116 4189 7118
rect 4204 7116 4238 7118
rect 4176 7100 4238 7116
rect 4282 7111 4298 7114
rect 4360 7111 4390 7122
rect 4438 7118 4484 7134
rect 4511 7122 4585 7138
rect 4438 7116 4472 7118
rect 4437 7100 4484 7116
rect 4511 7100 4524 7122
rect 4539 7100 4569 7122
rect 4596 7100 4597 7116
rect 4612 7100 4625 7260
rect 4655 7156 4668 7260
rect 4713 7238 4714 7248
rect 4729 7238 4742 7248
rect 4713 7234 4742 7238
rect 4747 7234 4777 7260
rect 4795 7246 4811 7248
rect 4883 7246 4936 7260
rect 4884 7244 4948 7246
rect 4991 7244 5006 7260
rect 5055 7257 5085 7260
rect 5055 7254 5091 7257
rect 5021 7246 5037 7248
rect 4795 7234 4810 7238
rect 4713 7232 4810 7234
rect 4838 7232 5006 7244
rect 5022 7234 5037 7238
rect 5055 7235 5094 7254
rect 5113 7248 5120 7249
rect 5119 7241 5120 7248
rect 5103 7238 5104 7241
rect 5119 7238 5132 7241
rect 5055 7234 5085 7235
rect 5094 7234 5100 7235
rect 5103 7234 5132 7238
rect 5022 7233 5132 7234
rect 5022 7232 5138 7233
rect 4697 7224 4748 7232
rect 4697 7212 4722 7224
rect 4729 7212 4748 7224
rect 4779 7224 4829 7232
rect 4779 7216 4795 7224
rect 4802 7222 4829 7224
rect 4838 7222 5059 7232
rect 4802 7212 5059 7222
rect 5088 7224 5138 7232
rect 5088 7215 5104 7224
rect 4697 7204 4748 7212
rect 4795 7204 5059 7212
rect 5085 7212 5104 7215
rect 5111 7212 5138 7224
rect 5085 7204 5138 7212
rect 4713 7196 4714 7204
rect 4729 7196 4742 7204
rect 4713 7188 4729 7196
rect 4710 7181 4729 7184
rect 4710 7172 4732 7181
rect 4683 7162 4732 7172
rect 4683 7156 4713 7162
rect 4732 7157 4737 7162
rect 4655 7140 4729 7156
rect 4747 7148 4777 7204
rect 4812 7194 5020 7204
rect 5055 7200 5100 7204
rect 5103 7203 5104 7204
rect 5119 7203 5132 7204
rect 4838 7164 5027 7194
rect 4853 7161 5027 7164
rect 4846 7158 5027 7161
rect 4655 7138 4668 7140
rect 4683 7138 4717 7140
rect 4655 7122 4729 7138
rect 4756 7134 4769 7148
rect 4784 7134 4800 7150
rect 4846 7145 4857 7158
rect 4639 7100 4640 7116
rect 4655 7100 4668 7122
rect 4683 7100 4713 7122
rect 4756 7118 4818 7134
rect 4846 7127 4857 7143
rect 4862 7138 4872 7158
rect 4882 7138 4896 7158
rect 4899 7145 4908 7158
rect 4924 7145 4933 7158
rect 4862 7127 4896 7138
rect 4899 7127 4908 7143
rect 4924 7127 4933 7143
rect 4940 7138 4950 7158
rect 4960 7138 4974 7158
rect 4975 7145 4986 7158
rect 4940 7127 4974 7138
rect 4975 7127 4986 7143
rect 5032 7134 5048 7150
rect 5055 7148 5085 7200
rect 5119 7196 5120 7203
rect 5104 7188 5120 7196
rect 5091 7156 5104 7175
rect 5119 7156 5149 7172
rect 5091 7140 5165 7156
rect 5091 7138 5104 7140
rect 5119 7138 5153 7140
rect 4756 7116 4769 7118
rect 4784 7116 4818 7118
rect 4756 7100 4818 7116
rect 4862 7111 4878 7114
rect 4940 7111 4970 7122
rect 5018 7118 5064 7134
rect 5091 7122 5165 7138
rect 5018 7116 5052 7118
rect 5017 7100 5064 7116
rect 5091 7100 5104 7122
rect 5119 7100 5149 7122
rect 5176 7100 5177 7116
rect 5192 7100 5205 7260
rect 5235 7156 5248 7260
rect 5293 7238 5294 7248
rect 5309 7238 5322 7248
rect 5293 7234 5322 7238
rect 5327 7234 5357 7260
rect 5375 7246 5391 7248
rect 5463 7246 5516 7260
rect 5464 7244 5528 7246
rect 5571 7244 5586 7260
rect 5635 7257 5665 7260
rect 5635 7254 5671 7257
rect 5601 7246 5617 7248
rect 5375 7234 5390 7238
rect 5293 7232 5390 7234
rect 5418 7232 5586 7244
rect 5602 7234 5617 7238
rect 5635 7235 5674 7254
rect 5693 7248 5700 7249
rect 5699 7241 5700 7248
rect 5683 7238 5684 7241
rect 5699 7238 5712 7241
rect 5635 7234 5665 7235
rect 5674 7234 5680 7235
rect 5683 7234 5712 7238
rect 5602 7233 5712 7234
rect 5602 7232 5718 7233
rect 5277 7224 5328 7232
rect 5277 7212 5302 7224
rect 5309 7212 5328 7224
rect 5359 7224 5409 7232
rect 5359 7216 5375 7224
rect 5382 7222 5409 7224
rect 5418 7222 5639 7232
rect 5382 7212 5639 7222
rect 5668 7224 5718 7232
rect 5668 7215 5684 7224
rect 5277 7204 5328 7212
rect 5375 7204 5639 7212
rect 5665 7212 5684 7215
rect 5691 7212 5718 7224
rect 5665 7204 5718 7212
rect 5293 7196 5294 7204
rect 5309 7196 5322 7204
rect 5293 7188 5309 7196
rect 5290 7181 5309 7184
rect 5290 7172 5312 7181
rect 5263 7162 5312 7172
rect 5263 7156 5293 7162
rect 5312 7157 5317 7162
rect 5235 7140 5309 7156
rect 5327 7148 5357 7204
rect 5392 7194 5600 7204
rect 5635 7200 5680 7204
rect 5683 7203 5684 7204
rect 5699 7203 5712 7204
rect 5418 7164 5607 7194
rect 5433 7161 5607 7164
rect 5426 7158 5607 7161
rect 5235 7138 5248 7140
rect 5263 7138 5297 7140
rect 5235 7122 5309 7138
rect 5336 7134 5349 7148
rect 5364 7134 5380 7150
rect 5426 7145 5437 7158
rect 5219 7100 5220 7116
rect 5235 7100 5248 7122
rect 5263 7100 5293 7122
rect 5336 7118 5398 7134
rect 5426 7127 5437 7143
rect 5442 7138 5452 7158
rect 5462 7138 5476 7158
rect 5479 7145 5488 7158
rect 5504 7145 5513 7158
rect 5442 7127 5476 7138
rect 5479 7127 5488 7143
rect 5504 7127 5513 7143
rect 5520 7138 5530 7158
rect 5540 7138 5554 7158
rect 5555 7145 5566 7158
rect 5520 7127 5554 7138
rect 5555 7127 5566 7143
rect 5612 7134 5628 7150
rect 5635 7148 5665 7200
rect 5699 7196 5700 7203
rect 5684 7188 5700 7196
rect 5671 7156 5684 7175
rect 5699 7156 5729 7172
rect 5671 7140 5745 7156
rect 5671 7138 5684 7140
rect 5699 7138 5733 7140
rect 5336 7116 5349 7118
rect 5364 7116 5398 7118
rect 5336 7100 5398 7116
rect 5442 7111 5458 7114
rect 5520 7111 5550 7122
rect 5598 7118 5644 7134
rect 5671 7122 5745 7138
rect 5598 7116 5632 7118
rect 5597 7100 5644 7116
rect 5671 7100 5684 7122
rect 5699 7100 5729 7122
rect 5756 7100 5757 7116
rect 5772 7100 5785 7260
rect 5815 7156 5828 7260
rect 5873 7238 5874 7248
rect 5889 7238 5902 7248
rect 5873 7234 5902 7238
rect 5907 7234 5937 7260
rect 5955 7246 5971 7248
rect 6043 7246 6096 7260
rect 6044 7244 6108 7246
rect 6151 7244 6166 7260
rect 6215 7257 6245 7260
rect 6215 7254 6251 7257
rect 6181 7246 6197 7248
rect 5955 7234 5970 7238
rect 5873 7232 5970 7234
rect 5998 7232 6166 7244
rect 6182 7234 6197 7238
rect 6215 7235 6254 7254
rect 6273 7248 6280 7249
rect 6279 7241 6280 7248
rect 6263 7238 6264 7241
rect 6279 7238 6292 7241
rect 6215 7234 6245 7235
rect 6254 7234 6260 7235
rect 6263 7234 6292 7238
rect 6182 7233 6292 7234
rect 6182 7232 6298 7233
rect 5857 7224 5908 7232
rect 5857 7212 5882 7224
rect 5889 7212 5908 7224
rect 5939 7224 5989 7232
rect 5939 7216 5955 7224
rect 5962 7222 5989 7224
rect 5998 7222 6219 7232
rect 5962 7212 6219 7222
rect 6248 7224 6298 7232
rect 6248 7215 6264 7224
rect 5857 7204 5908 7212
rect 5955 7204 6219 7212
rect 6245 7212 6264 7215
rect 6271 7212 6298 7224
rect 6245 7204 6298 7212
rect 5873 7196 5874 7204
rect 5889 7196 5902 7204
rect 5873 7188 5889 7196
rect 5870 7181 5889 7184
rect 5870 7172 5892 7181
rect 5843 7162 5892 7172
rect 5843 7156 5873 7162
rect 5892 7157 5897 7162
rect 5815 7140 5889 7156
rect 5907 7148 5937 7204
rect 5972 7194 6180 7204
rect 6215 7200 6260 7204
rect 6263 7203 6264 7204
rect 6279 7203 6292 7204
rect 5998 7164 6187 7194
rect 6013 7161 6187 7164
rect 6006 7158 6187 7161
rect 5815 7138 5828 7140
rect 5843 7138 5877 7140
rect 5815 7122 5889 7138
rect 5916 7134 5929 7148
rect 5944 7134 5960 7150
rect 6006 7145 6017 7158
rect 5799 7100 5800 7116
rect 5815 7100 5828 7122
rect 5843 7100 5873 7122
rect 5916 7118 5978 7134
rect 6006 7127 6017 7143
rect 6022 7138 6032 7158
rect 6042 7138 6056 7158
rect 6059 7145 6068 7158
rect 6084 7145 6093 7158
rect 6022 7127 6056 7138
rect 6059 7127 6068 7143
rect 6084 7127 6093 7143
rect 6100 7138 6110 7158
rect 6120 7138 6134 7158
rect 6135 7145 6146 7158
rect 6100 7127 6134 7138
rect 6135 7127 6146 7143
rect 6192 7134 6208 7150
rect 6215 7148 6245 7200
rect 6279 7196 6280 7203
rect 6264 7188 6280 7196
rect 6251 7156 6264 7175
rect 6279 7156 6309 7172
rect 6251 7140 6325 7156
rect 6251 7138 6264 7140
rect 6279 7138 6313 7140
rect 5916 7116 5929 7118
rect 5944 7116 5978 7118
rect 5916 7100 5978 7116
rect 6022 7111 6038 7114
rect 6100 7111 6130 7122
rect 6178 7118 6224 7134
rect 6251 7122 6325 7138
rect 6178 7116 6212 7118
rect 6177 7100 6224 7116
rect 6251 7100 6264 7122
rect 6279 7100 6309 7122
rect 6336 7100 6337 7116
rect 6352 7100 6365 7260
rect 6395 7156 6408 7260
rect 6453 7238 6454 7248
rect 6469 7238 6482 7248
rect 6453 7234 6482 7238
rect 6487 7234 6517 7260
rect 6535 7246 6551 7248
rect 6623 7246 6676 7260
rect 6624 7244 6688 7246
rect 6731 7244 6746 7260
rect 6795 7257 6825 7260
rect 6795 7254 6831 7257
rect 6761 7246 6777 7248
rect 6535 7234 6550 7238
rect 6453 7232 6550 7234
rect 6578 7232 6746 7244
rect 6762 7234 6777 7238
rect 6795 7235 6834 7254
rect 6853 7248 6860 7249
rect 6859 7241 6860 7248
rect 6843 7238 6844 7241
rect 6859 7238 6872 7241
rect 6795 7234 6825 7235
rect 6834 7234 6840 7235
rect 6843 7234 6872 7238
rect 6762 7233 6872 7234
rect 6762 7232 6878 7233
rect 6437 7224 6488 7232
rect 6437 7212 6462 7224
rect 6469 7212 6488 7224
rect 6519 7224 6569 7232
rect 6519 7216 6535 7224
rect 6542 7222 6569 7224
rect 6578 7222 6799 7232
rect 6542 7212 6799 7222
rect 6828 7224 6878 7232
rect 6828 7215 6844 7224
rect 6437 7204 6488 7212
rect 6535 7204 6799 7212
rect 6825 7212 6844 7215
rect 6851 7212 6878 7224
rect 6825 7204 6878 7212
rect 6453 7196 6454 7204
rect 6469 7196 6482 7204
rect 6453 7188 6469 7196
rect 6450 7181 6469 7184
rect 6450 7172 6472 7181
rect 6423 7162 6472 7172
rect 6423 7156 6453 7162
rect 6472 7157 6477 7162
rect 6395 7140 6469 7156
rect 6487 7148 6517 7204
rect 6552 7194 6760 7204
rect 6795 7200 6840 7204
rect 6843 7203 6844 7204
rect 6859 7203 6872 7204
rect 6578 7164 6767 7194
rect 6593 7161 6767 7164
rect 6586 7158 6767 7161
rect 6395 7138 6408 7140
rect 6423 7138 6457 7140
rect 6395 7122 6469 7138
rect 6496 7134 6509 7148
rect 6524 7134 6540 7150
rect 6586 7145 6597 7158
rect 6379 7100 6380 7116
rect 6395 7100 6408 7122
rect 6423 7100 6453 7122
rect 6496 7118 6558 7134
rect 6586 7127 6597 7143
rect 6602 7138 6612 7158
rect 6622 7138 6636 7158
rect 6639 7145 6648 7158
rect 6664 7145 6673 7158
rect 6602 7127 6636 7138
rect 6639 7127 6648 7143
rect 6664 7127 6673 7143
rect 6680 7138 6690 7158
rect 6700 7138 6714 7158
rect 6715 7145 6726 7158
rect 6680 7127 6714 7138
rect 6715 7127 6726 7143
rect 6772 7134 6788 7150
rect 6795 7148 6825 7200
rect 6859 7196 6860 7203
rect 6844 7188 6860 7196
rect 6831 7156 6844 7175
rect 6859 7156 6889 7172
rect 6831 7140 6905 7156
rect 6831 7138 6844 7140
rect 6859 7138 6893 7140
rect 6496 7116 6509 7118
rect 6524 7116 6558 7118
rect 6496 7100 6558 7116
rect 6602 7111 6618 7114
rect 6680 7111 6710 7122
rect 6758 7118 6804 7134
rect 6831 7122 6905 7138
rect 6758 7116 6792 7118
rect 6757 7100 6804 7116
rect 6831 7100 6844 7122
rect 6859 7100 6889 7122
rect 6916 7100 6917 7116
rect 6932 7100 6945 7260
rect 6975 7156 6988 7260
rect 7033 7238 7034 7248
rect 7049 7238 7062 7248
rect 7033 7234 7062 7238
rect 7067 7234 7097 7260
rect 7115 7246 7131 7248
rect 7203 7246 7256 7260
rect 7204 7244 7268 7246
rect 7311 7244 7326 7260
rect 7375 7257 7405 7260
rect 7375 7254 7411 7257
rect 7341 7246 7357 7248
rect 7115 7234 7130 7238
rect 7033 7232 7130 7234
rect 7158 7232 7326 7244
rect 7342 7234 7357 7238
rect 7375 7235 7414 7254
rect 7433 7248 7440 7249
rect 7439 7241 7440 7248
rect 7423 7238 7424 7241
rect 7439 7238 7452 7241
rect 7375 7234 7405 7235
rect 7414 7234 7420 7235
rect 7423 7234 7452 7238
rect 7342 7233 7452 7234
rect 7342 7232 7458 7233
rect 7017 7224 7068 7232
rect 7017 7212 7042 7224
rect 7049 7212 7068 7224
rect 7099 7224 7149 7232
rect 7099 7216 7115 7224
rect 7122 7222 7149 7224
rect 7158 7222 7379 7232
rect 7122 7212 7379 7222
rect 7408 7224 7458 7232
rect 7408 7215 7424 7224
rect 7017 7204 7068 7212
rect 7115 7204 7379 7212
rect 7405 7212 7424 7215
rect 7431 7212 7458 7224
rect 7405 7204 7458 7212
rect 7033 7196 7034 7204
rect 7049 7196 7062 7204
rect 7033 7188 7049 7196
rect 7030 7181 7049 7184
rect 7030 7172 7052 7181
rect 7003 7162 7052 7172
rect 7003 7156 7033 7162
rect 7052 7157 7057 7162
rect 6975 7140 7049 7156
rect 7067 7148 7097 7204
rect 7132 7194 7340 7204
rect 7375 7200 7420 7204
rect 7423 7203 7424 7204
rect 7439 7203 7452 7204
rect 7158 7164 7347 7194
rect 7173 7161 7347 7164
rect 7166 7158 7347 7161
rect 6975 7138 6988 7140
rect 7003 7138 7037 7140
rect 6975 7122 7049 7138
rect 7076 7134 7089 7148
rect 7104 7134 7120 7150
rect 7166 7145 7177 7158
rect 6959 7100 6960 7116
rect 6975 7100 6988 7122
rect 7003 7100 7033 7122
rect 7076 7118 7138 7134
rect 7166 7127 7177 7143
rect 7182 7138 7192 7158
rect 7202 7138 7216 7158
rect 7219 7145 7228 7158
rect 7244 7145 7253 7158
rect 7182 7127 7216 7138
rect 7219 7127 7228 7143
rect 7244 7127 7253 7143
rect 7260 7138 7270 7158
rect 7280 7138 7294 7158
rect 7295 7145 7306 7158
rect 7260 7127 7294 7138
rect 7295 7127 7306 7143
rect 7352 7134 7368 7150
rect 7375 7148 7405 7200
rect 7439 7196 7440 7203
rect 7424 7188 7440 7196
rect 7411 7156 7424 7175
rect 7439 7156 7469 7172
rect 7411 7140 7485 7156
rect 7411 7138 7424 7140
rect 7439 7138 7473 7140
rect 7076 7116 7089 7118
rect 7104 7116 7138 7118
rect 7076 7100 7138 7116
rect 7182 7111 7198 7114
rect 7260 7111 7290 7122
rect 7338 7118 7384 7134
rect 7411 7122 7485 7138
rect 7338 7116 7372 7118
rect 7337 7100 7384 7116
rect 7411 7100 7424 7122
rect 7439 7100 7469 7122
rect 7496 7100 7497 7116
rect 7512 7100 7525 7260
rect 7555 7156 7568 7260
rect 7613 7238 7614 7248
rect 7629 7238 7642 7248
rect 7613 7234 7642 7238
rect 7647 7234 7677 7260
rect 7695 7246 7711 7248
rect 7783 7246 7836 7260
rect 7784 7244 7848 7246
rect 7891 7244 7906 7260
rect 7955 7257 7985 7260
rect 7955 7254 7991 7257
rect 7921 7246 7937 7248
rect 7695 7234 7710 7238
rect 7613 7232 7710 7234
rect 7738 7232 7906 7244
rect 7922 7234 7937 7238
rect 7955 7235 7994 7254
rect 8013 7248 8020 7249
rect 8019 7241 8020 7248
rect 8003 7238 8004 7241
rect 8019 7238 8032 7241
rect 7955 7234 7985 7235
rect 7994 7234 8000 7235
rect 8003 7234 8032 7238
rect 7922 7233 8032 7234
rect 7922 7232 8038 7233
rect 7597 7224 7648 7232
rect 7597 7212 7622 7224
rect 7629 7212 7648 7224
rect 7679 7224 7729 7232
rect 7679 7216 7695 7224
rect 7702 7222 7729 7224
rect 7738 7222 7959 7232
rect 7702 7212 7959 7222
rect 7988 7224 8038 7232
rect 7988 7215 8004 7224
rect 7597 7204 7648 7212
rect 7695 7204 7959 7212
rect 7985 7212 8004 7215
rect 8011 7212 8038 7224
rect 7985 7204 8038 7212
rect 7613 7196 7614 7204
rect 7629 7196 7642 7204
rect 7613 7188 7629 7196
rect 7610 7181 7629 7184
rect 7610 7172 7632 7181
rect 7583 7162 7632 7172
rect 7583 7156 7613 7162
rect 7632 7157 7637 7162
rect 7555 7140 7629 7156
rect 7647 7148 7677 7204
rect 7712 7194 7920 7204
rect 7955 7200 8000 7204
rect 8003 7203 8004 7204
rect 8019 7203 8032 7204
rect 7738 7164 7927 7194
rect 7753 7161 7927 7164
rect 7746 7158 7927 7161
rect 7555 7138 7568 7140
rect 7583 7138 7617 7140
rect 7555 7122 7629 7138
rect 7656 7134 7669 7148
rect 7684 7134 7700 7150
rect 7746 7145 7757 7158
rect 7539 7100 7540 7116
rect 7555 7100 7568 7122
rect 7583 7100 7613 7122
rect 7656 7118 7718 7134
rect 7746 7127 7757 7143
rect 7762 7138 7772 7158
rect 7782 7138 7796 7158
rect 7799 7145 7808 7158
rect 7824 7145 7833 7158
rect 7762 7127 7796 7138
rect 7799 7127 7808 7143
rect 7824 7127 7833 7143
rect 7840 7138 7850 7158
rect 7860 7138 7874 7158
rect 7875 7145 7886 7158
rect 7840 7127 7874 7138
rect 7875 7127 7886 7143
rect 7932 7134 7948 7150
rect 7955 7148 7985 7200
rect 8019 7196 8020 7203
rect 8004 7188 8020 7196
rect 7991 7156 8004 7175
rect 8019 7156 8049 7172
rect 7991 7140 8065 7156
rect 7991 7138 8004 7140
rect 8019 7138 8053 7140
rect 7656 7116 7669 7118
rect 7684 7116 7718 7118
rect 7656 7100 7718 7116
rect 7762 7111 7778 7114
rect 7840 7111 7870 7122
rect 7918 7118 7964 7134
rect 7991 7122 8065 7138
rect 7918 7116 7952 7118
rect 7917 7100 7964 7116
rect 7991 7100 8004 7122
rect 8019 7100 8049 7122
rect 8076 7100 8077 7116
rect 8092 7100 8105 7260
rect 8135 7156 8148 7260
rect 8193 7238 8194 7248
rect 8209 7238 8222 7248
rect 8193 7234 8222 7238
rect 8227 7234 8257 7260
rect 8275 7246 8291 7248
rect 8363 7246 8416 7260
rect 8364 7244 8428 7246
rect 8471 7244 8486 7260
rect 8535 7257 8565 7260
rect 8535 7254 8571 7257
rect 8501 7246 8517 7248
rect 8275 7234 8290 7238
rect 8193 7232 8290 7234
rect 8318 7232 8486 7244
rect 8502 7234 8517 7238
rect 8535 7235 8574 7254
rect 8593 7248 8600 7249
rect 8599 7241 8600 7248
rect 8583 7238 8584 7241
rect 8599 7238 8612 7241
rect 8535 7234 8565 7235
rect 8574 7234 8580 7235
rect 8583 7234 8612 7238
rect 8502 7233 8612 7234
rect 8502 7232 8618 7233
rect 8177 7224 8228 7232
rect 8177 7212 8202 7224
rect 8209 7212 8228 7224
rect 8259 7224 8309 7232
rect 8259 7216 8275 7224
rect 8282 7222 8309 7224
rect 8318 7222 8539 7232
rect 8282 7212 8539 7222
rect 8568 7224 8618 7232
rect 8568 7215 8584 7224
rect 8177 7204 8228 7212
rect 8275 7204 8539 7212
rect 8565 7212 8584 7215
rect 8591 7212 8618 7224
rect 8565 7204 8618 7212
rect 8193 7196 8194 7204
rect 8209 7196 8222 7204
rect 8193 7188 8209 7196
rect 8190 7181 8209 7184
rect 8190 7172 8212 7181
rect 8163 7162 8212 7172
rect 8163 7156 8193 7162
rect 8212 7157 8217 7162
rect 8135 7140 8209 7156
rect 8227 7148 8257 7204
rect 8292 7194 8500 7204
rect 8535 7200 8580 7204
rect 8583 7203 8584 7204
rect 8599 7203 8612 7204
rect 8318 7164 8507 7194
rect 8333 7161 8507 7164
rect 8326 7158 8507 7161
rect 8135 7138 8148 7140
rect 8163 7138 8197 7140
rect 8135 7122 8209 7138
rect 8236 7134 8249 7148
rect 8264 7134 8280 7150
rect 8326 7145 8337 7158
rect 8119 7100 8120 7116
rect 8135 7100 8148 7122
rect 8163 7100 8193 7122
rect 8236 7118 8298 7134
rect 8326 7127 8337 7143
rect 8342 7138 8352 7158
rect 8362 7138 8376 7158
rect 8379 7145 8388 7158
rect 8404 7145 8413 7158
rect 8342 7127 8376 7138
rect 8379 7127 8388 7143
rect 8404 7127 8413 7143
rect 8420 7138 8430 7158
rect 8440 7138 8454 7158
rect 8455 7145 8466 7158
rect 8420 7127 8454 7138
rect 8455 7127 8466 7143
rect 8512 7134 8528 7150
rect 8535 7148 8565 7200
rect 8599 7196 8600 7203
rect 8584 7188 8600 7196
rect 8571 7156 8584 7175
rect 8599 7156 8629 7172
rect 8571 7140 8645 7156
rect 8571 7138 8584 7140
rect 8599 7138 8633 7140
rect 8236 7116 8249 7118
rect 8264 7116 8298 7118
rect 8236 7100 8298 7116
rect 8342 7111 8358 7114
rect 8420 7111 8450 7122
rect 8498 7118 8544 7134
rect 8571 7122 8645 7138
rect 8498 7116 8532 7118
rect 8497 7100 8544 7116
rect 8571 7100 8584 7122
rect 8599 7100 8629 7122
rect 8656 7100 8657 7116
rect 8672 7100 8685 7260
rect 8715 7156 8728 7260
rect 8773 7238 8774 7248
rect 8789 7238 8802 7248
rect 8773 7234 8802 7238
rect 8807 7234 8837 7260
rect 8855 7246 8871 7248
rect 8943 7246 8996 7260
rect 8944 7244 9008 7246
rect 9051 7244 9066 7260
rect 9115 7257 9145 7260
rect 9115 7254 9151 7257
rect 9081 7246 9097 7248
rect 8855 7234 8870 7238
rect 8773 7232 8870 7234
rect 8898 7232 9066 7244
rect 9082 7234 9097 7238
rect 9115 7235 9154 7254
rect 9173 7248 9180 7249
rect 9179 7241 9180 7248
rect 9163 7238 9164 7241
rect 9179 7238 9192 7241
rect 9115 7234 9145 7235
rect 9154 7234 9160 7235
rect 9163 7234 9192 7238
rect 9082 7233 9192 7234
rect 9082 7232 9198 7233
rect 8757 7224 8808 7232
rect 8757 7212 8782 7224
rect 8789 7212 8808 7224
rect 8839 7224 8889 7232
rect 8839 7216 8855 7224
rect 8862 7222 8889 7224
rect 8898 7222 9119 7232
rect 8862 7212 9119 7222
rect 9148 7224 9198 7232
rect 9148 7215 9164 7224
rect 8757 7204 8808 7212
rect 8855 7204 9119 7212
rect 9145 7212 9164 7215
rect 9171 7212 9198 7224
rect 9145 7204 9198 7212
rect 8773 7196 8774 7204
rect 8789 7196 8802 7204
rect 8773 7188 8789 7196
rect 8770 7181 8789 7184
rect 8770 7172 8792 7181
rect 8743 7162 8792 7172
rect 8743 7156 8773 7162
rect 8792 7157 8797 7162
rect 8715 7140 8789 7156
rect 8807 7148 8837 7204
rect 8872 7194 9080 7204
rect 9115 7200 9160 7204
rect 9163 7203 9164 7204
rect 9179 7203 9192 7204
rect 8898 7164 9087 7194
rect 8913 7161 9087 7164
rect 8906 7158 9087 7161
rect 8715 7138 8728 7140
rect 8743 7138 8777 7140
rect 8715 7122 8789 7138
rect 8816 7134 8829 7148
rect 8844 7134 8860 7150
rect 8906 7145 8917 7158
rect 8699 7100 8700 7116
rect 8715 7100 8728 7122
rect 8743 7100 8773 7122
rect 8816 7118 8878 7134
rect 8906 7127 8917 7143
rect 8922 7138 8932 7158
rect 8942 7138 8956 7158
rect 8959 7145 8968 7158
rect 8984 7145 8993 7158
rect 8922 7127 8956 7138
rect 8959 7127 8968 7143
rect 8984 7127 8993 7143
rect 9000 7138 9010 7158
rect 9020 7138 9034 7158
rect 9035 7145 9046 7158
rect 9000 7127 9034 7138
rect 9035 7127 9046 7143
rect 9092 7134 9108 7150
rect 9115 7148 9145 7200
rect 9179 7196 9180 7203
rect 9164 7188 9180 7196
rect 9151 7156 9164 7175
rect 9179 7156 9209 7172
rect 9151 7140 9225 7156
rect 9151 7138 9164 7140
rect 9179 7138 9213 7140
rect 8816 7116 8829 7118
rect 8844 7116 8878 7118
rect 8816 7100 8878 7116
rect 8922 7111 8938 7114
rect 9000 7111 9030 7122
rect 9078 7118 9124 7134
rect 9151 7122 9225 7138
rect 9078 7116 9112 7118
rect 9077 7100 9124 7116
rect 9151 7100 9164 7122
rect 9179 7100 9209 7122
rect 9236 7100 9237 7116
rect 9252 7100 9265 7260
rect -7 7092 34 7100
rect -7 7066 8 7092
rect 15 7066 34 7092
rect 98 7088 160 7100
rect 172 7088 247 7100
rect 305 7088 380 7100
rect 392 7088 423 7100
rect 429 7088 464 7100
rect 98 7086 260 7088
rect -7 7058 34 7066
rect 116 7062 129 7086
rect 144 7084 159 7086
rect -1 7048 0 7058
rect 15 7048 28 7058
rect 43 7048 73 7062
rect 116 7048 159 7062
rect 183 7059 190 7066
rect 193 7062 260 7086
rect 292 7086 464 7088
rect 262 7064 290 7068
rect 292 7064 372 7086
rect 393 7084 408 7086
rect 262 7062 372 7064
rect 193 7058 372 7062
rect 166 7048 196 7058
rect 198 7048 351 7058
rect 359 7048 389 7058
rect 393 7048 423 7062
rect 451 7048 464 7086
rect 536 7092 571 7100
rect 536 7066 537 7092
rect 544 7066 571 7092
rect 479 7048 509 7062
rect 536 7058 571 7066
rect 573 7092 614 7100
rect 573 7066 588 7092
rect 595 7066 614 7092
rect 678 7088 740 7100
rect 752 7088 827 7100
rect 885 7088 960 7100
rect 972 7088 1003 7100
rect 1009 7088 1044 7100
rect 678 7086 840 7088
rect 573 7058 614 7066
rect 696 7062 709 7086
rect 724 7084 739 7086
rect 536 7048 537 7058
rect 552 7048 565 7058
rect 579 7048 580 7058
rect 595 7048 608 7058
rect 623 7048 653 7062
rect 696 7048 739 7062
rect 763 7059 770 7066
rect 773 7062 840 7086
rect 872 7086 1044 7088
rect 842 7064 870 7068
rect 872 7064 952 7086
rect 973 7084 988 7086
rect 842 7062 952 7064
rect 773 7058 952 7062
rect 746 7048 776 7058
rect 778 7048 931 7058
rect 939 7048 969 7058
rect 973 7048 1003 7062
rect 1031 7048 1044 7086
rect 1116 7092 1151 7100
rect 1116 7066 1117 7092
rect 1124 7066 1151 7092
rect 1059 7048 1089 7062
rect 1116 7058 1151 7066
rect 1153 7092 1194 7100
rect 1153 7066 1168 7092
rect 1175 7066 1194 7092
rect 1258 7088 1320 7100
rect 1332 7088 1407 7100
rect 1465 7088 1540 7100
rect 1552 7088 1583 7100
rect 1589 7088 1624 7100
rect 1258 7086 1420 7088
rect 1153 7058 1194 7066
rect 1276 7062 1289 7086
rect 1304 7084 1319 7086
rect 1116 7048 1117 7058
rect 1132 7048 1145 7058
rect 1159 7048 1160 7058
rect 1175 7048 1188 7058
rect 1203 7048 1233 7062
rect 1276 7048 1319 7062
rect 1343 7059 1350 7066
rect 1353 7062 1420 7086
rect 1452 7086 1624 7088
rect 1422 7064 1450 7068
rect 1452 7064 1532 7086
rect 1553 7084 1568 7086
rect 1422 7062 1532 7064
rect 1353 7058 1532 7062
rect 1326 7048 1356 7058
rect 1358 7048 1511 7058
rect 1519 7048 1549 7058
rect 1553 7048 1583 7062
rect 1611 7048 1624 7086
rect 1696 7092 1731 7100
rect 1696 7066 1697 7092
rect 1704 7066 1731 7092
rect 1639 7048 1669 7062
rect 1696 7058 1731 7066
rect 1733 7092 1774 7100
rect 1733 7066 1748 7092
rect 1755 7066 1774 7092
rect 1838 7088 1900 7100
rect 1912 7088 1987 7100
rect 2045 7088 2120 7100
rect 2132 7088 2163 7100
rect 2169 7088 2204 7100
rect 1838 7086 2000 7088
rect 1733 7058 1774 7066
rect 1856 7062 1869 7086
rect 1884 7084 1899 7086
rect 1696 7048 1697 7058
rect 1712 7048 1725 7058
rect 1739 7048 1740 7058
rect 1755 7048 1768 7058
rect 1783 7048 1813 7062
rect 1856 7048 1899 7062
rect 1923 7059 1930 7066
rect 1933 7062 2000 7086
rect 2032 7086 2204 7088
rect 2002 7064 2030 7068
rect 2032 7064 2112 7086
rect 2133 7084 2148 7086
rect 2002 7062 2112 7064
rect 1933 7058 2112 7062
rect 1906 7048 1936 7058
rect 1938 7048 2091 7058
rect 2099 7048 2129 7058
rect 2133 7048 2163 7062
rect 2191 7048 2204 7086
rect 2276 7092 2311 7100
rect 2276 7066 2277 7092
rect 2284 7066 2311 7092
rect 2219 7048 2249 7062
rect 2276 7058 2311 7066
rect 2313 7092 2354 7100
rect 2313 7066 2328 7092
rect 2335 7066 2354 7092
rect 2418 7088 2480 7100
rect 2492 7088 2567 7100
rect 2625 7088 2700 7100
rect 2712 7088 2743 7100
rect 2749 7088 2784 7100
rect 2418 7086 2580 7088
rect 2313 7058 2354 7066
rect 2436 7062 2449 7086
rect 2464 7084 2479 7086
rect 2276 7048 2277 7058
rect 2292 7048 2305 7058
rect 2319 7048 2320 7058
rect 2335 7048 2348 7058
rect 2363 7048 2393 7062
rect 2436 7048 2479 7062
rect 2503 7059 2510 7066
rect 2513 7062 2580 7086
rect 2612 7086 2784 7088
rect 2582 7064 2610 7068
rect 2612 7064 2692 7086
rect 2713 7084 2728 7086
rect 2582 7062 2692 7064
rect 2513 7058 2692 7062
rect 2486 7048 2516 7058
rect 2518 7048 2671 7058
rect 2679 7048 2709 7058
rect 2713 7048 2743 7062
rect 2771 7048 2784 7086
rect 2856 7092 2891 7100
rect 2856 7066 2857 7092
rect 2864 7066 2891 7092
rect 2799 7048 2829 7062
rect 2856 7058 2891 7066
rect 2893 7092 2934 7100
rect 2893 7066 2908 7092
rect 2915 7066 2934 7092
rect 2998 7088 3060 7100
rect 3072 7088 3147 7100
rect 3205 7088 3280 7100
rect 3292 7088 3323 7100
rect 3329 7088 3364 7100
rect 2998 7086 3160 7088
rect 2893 7058 2934 7066
rect 3016 7062 3029 7086
rect 3044 7084 3059 7086
rect 2856 7048 2857 7058
rect 2872 7048 2885 7058
rect 2899 7048 2900 7058
rect 2915 7048 2928 7058
rect 2943 7048 2973 7062
rect 3016 7048 3059 7062
rect 3083 7059 3090 7066
rect 3093 7062 3160 7086
rect 3192 7086 3364 7088
rect 3162 7064 3190 7068
rect 3192 7064 3272 7086
rect 3293 7084 3308 7086
rect 3162 7062 3272 7064
rect 3093 7058 3272 7062
rect 3066 7048 3096 7058
rect 3098 7048 3251 7058
rect 3259 7048 3289 7058
rect 3293 7048 3323 7062
rect 3351 7048 3364 7086
rect 3436 7092 3471 7100
rect 3436 7066 3437 7092
rect 3444 7066 3471 7092
rect 3379 7048 3409 7062
rect 3436 7058 3471 7066
rect 3473 7092 3514 7100
rect 3473 7066 3488 7092
rect 3495 7066 3514 7092
rect 3578 7088 3640 7100
rect 3652 7088 3727 7100
rect 3785 7088 3860 7100
rect 3872 7088 3903 7100
rect 3909 7088 3944 7100
rect 3578 7086 3740 7088
rect 3473 7058 3514 7066
rect 3596 7062 3609 7086
rect 3624 7084 3639 7086
rect 3436 7048 3437 7058
rect 3452 7048 3465 7058
rect 3479 7048 3480 7058
rect 3495 7048 3508 7058
rect 3523 7048 3553 7062
rect 3596 7048 3639 7062
rect 3663 7059 3670 7066
rect 3673 7062 3740 7086
rect 3772 7086 3944 7088
rect 3742 7064 3770 7068
rect 3772 7064 3852 7086
rect 3873 7084 3888 7086
rect 3742 7062 3852 7064
rect 3673 7058 3852 7062
rect 3646 7048 3676 7058
rect 3678 7048 3831 7058
rect 3839 7048 3869 7058
rect 3873 7048 3903 7062
rect 3931 7048 3944 7086
rect 4016 7092 4051 7100
rect 4016 7066 4017 7092
rect 4024 7066 4051 7092
rect 3959 7048 3989 7062
rect 4016 7058 4051 7066
rect 4053 7092 4094 7100
rect 4053 7066 4068 7092
rect 4075 7066 4094 7092
rect 4158 7088 4220 7100
rect 4232 7088 4307 7100
rect 4365 7088 4440 7100
rect 4452 7088 4483 7100
rect 4489 7088 4524 7100
rect 4158 7086 4320 7088
rect 4053 7058 4094 7066
rect 4176 7062 4189 7086
rect 4204 7084 4219 7086
rect 4016 7048 4017 7058
rect 4032 7048 4045 7058
rect 4059 7048 4060 7058
rect 4075 7048 4088 7058
rect 4103 7048 4133 7062
rect 4176 7048 4219 7062
rect 4243 7059 4250 7066
rect 4253 7062 4320 7086
rect 4352 7086 4524 7088
rect 4322 7064 4350 7068
rect 4352 7064 4432 7086
rect 4453 7084 4468 7086
rect 4322 7062 4432 7064
rect 4253 7058 4432 7062
rect 4226 7048 4256 7058
rect 4258 7048 4411 7058
rect 4419 7048 4449 7058
rect 4453 7048 4483 7062
rect 4511 7048 4524 7086
rect 4596 7092 4631 7100
rect 4596 7066 4597 7092
rect 4604 7066 4631 7092
rect 4539 7048 4569 7062
rect 4596 7058 4631 7066
rect 4633 7092 4674 7100
rect 4633 7066 4648 7092
rect 4655 7066 4674 7092
rect 4738 7088 4800 7100
rect 4812 7088 4887 7100
rect 4945 7088 5020 7100
rect 5032 7088 5063 7100
rect 5069 7088 5104 7100
rect 4738 7086 4900 7088
rect 4633 7058 4674 7066
rect 4756 7062 4769 7086
rect 4784 7084 4799 7086
rect 4596 7048 4597 7058
rect 4612 7048 4625 7058
rect 4639 7048 4640 7058
rect 4655 7048 4668 7058
rect 4683 7048 4713 7062
rect 4756 7048 4799 7062
rect 4823 7059 4830 7066
rect 4833 7062 4900 7086
rect 4932 7086 5104 7088
rect 4902 7064 4930 7068
rect 4932 7064 5012 7086
rect 5033 7084 5048 7086
rect 4902 7062 5012 7064
rect 4833 7058 5012 7062
rect 4806 7048 4836 7058
rect 4838 7048 4991 7058
rect 4999 7048 5029 7058
rect 5033 7048 5063 7062
rect 5091 7048 5104 7086
rect 5176 7092 5211 7100
rect 5176 7066 5177 7092
rect 5184 7066 5211 7092
rect 5119 7048 5149 7062
rect 5176 7058 5211 7066
rect 5213 7092 5254 7100
rect 5213 7066 5228 7092
rect 5235 7066 5254 7092
rect 5318 7088 5380 7100
rect 5392 7088 5467 7100
rect 5525 7088 5600 7100
rect 5612 7088 5643 7100
rect 5649 7088 5684 7100
rect 5318 7086 5480 7088
rect 5213 7058 5254 7066
rect 5336 7062 5349 7086
rect 5364 7084 5379 7086
rect 5176 7048 5177 7058
rect 5192 7048 5205 7058
rect 5219 7048 5220 7058
rect 5235 7048 5248 7058
rect 5263 7048 5293 7062
rect 5336 7048 5379 7062
rect 5403 7059 5410 7066
rect 5413 7062 5480 7086
rect 5512 7086 5684 7088
rect 5482 7064 5510 7068
rect 5512 7064 5592 7086
rect 5613 7084 5628 7086
rect 5482 7062 5592 7064
rect 5413 7058 5592 7062
rect 5386 7048 5416 7058
rect 5418 7048 5571 7058
rect 5579 7048 5609 7058
rect 5613 7048 5643 7062
rect 5671 7048 5684 7086
rect 5756 7092 5791 7100
rect 5756 7066 5757 7092
rect 5764 7066 5791 7092
rect 5699 7048 5729 7062
rect 5756 7058 5791 7066
rect 5793 7092 5834 7100
rect 5793 7066 5808 7092
rect 5815 7066 5834 7092
rect 5898 7088 5960 7100
rect 5972 7088 6047 7100
rect 6105 7088 6180 7100
rect 6192 7088 6223 7100
rect 6229 7088 6264 7100
rect 5898 7086 6060 7088
rect 5793 7058 5834 7066
rect 5916 7062 5929 7086
rect 5944 7084 5959 7086
rect 5756 7048 5757 7058
rect 5772 7048 5785 7058
rect 5799 7048 5800 7058
rect 5815 7048 5828 7058
rect 5843 7048 5873 7062
rect 5916 7048 5959 7062
rect 5983 7059 5990 7066
rect 5993 7062 6060 7086
rect 6092 7086 6264 7088
rect 6062 7064 6090 7068
rect 6092 7064 6172 7086
rect 6193 7084 6208 7086
rect 6062 7062 6172 7064
rect 5993 7058 6172 7062
rect 5966 7048 5996 7058
rect 5998 7048 6151 7058
rect 6159 7048 6189 7058
rect 6193 7048 6223 7062
rect 6251 7048 6264 7086
rect 6336 7092 6371 7100
rect 6336 7066 6337 7092
rect 6344 7066 6371 7092
rect 6279 7048 6309 7062
rect 6336 7058 6371 7066
rect 6373 7092 6414 7100
rect 6373 7066 6388 7092
rect 6395 7066 6414 7092
rect 6478 7088 6540 7100
rect 6552 7088 6627 7100
rect 6685 7088 6760 7100
rect 6772 7088 6803 7100
rect 6809 7088 6844 7100
rect 6478 7086 6640 7088
rect 6373 7058 6414 7066
rect 6496 7062 6509 7086
rect 6524 7084 6539 7086
rect 6336 7048 6337 7058
rect 6352 7048 6365 7058
rect 6379 7048 6380 7058
rect 6395 7048 6408 7058
rect 6423 7048 6453 7062
rect 6496 7048 6539 7062
rect 6563 7059 6570 7066
rect 6573 7062 6640 7086
rect 6672 7086 6844 7088
rect 6642 7064 6670 7068
rect 6672 7064 6752 7086
rect 6773 7084 6788 7086
rect 6642 7062 6752 7064
rect 6573 7058 6752 7062
rect 6546 7048 6576 7058
rect 6578 7048 6731 7058
rect 6739 7048 6769 7058
rect 6773 7048 6803 7062
rect 6831 7048 6844 7086
rect 6916 7092 6951 7100
rect 6916 7066 6917 7092
rect 6924 7066 6951 7092
rect 6859 7048 6889 7062
rect 6916 7058 6951 7066
rect 6953 7092 6994 7100
rect 6953 7066 6968 7092
rect 6975 7066 6994 7092
rect 7058 7088 7120 7100
rect 7132 7088 7207 7100
rect 7265 7088 7340 7100
rect 7352 7088 7383 7100
rect 7389 7088 7424 7100
rect 7058 7086 7220 7088
rect 6953 7058 6994 7066
rect 7076 7062 7089 7086
rect 7104 7084 7119 7086
rect 6916 7048 6917 7058
rect 6932 7048 6945 7058
rect 6959 7048 6960 7058
rect 6975 7048 6988 7058
rect 7003 7048 7033 7062
rect 7076 7048 7119 7062
rect 7143 7059 7150 7066
rect 7153 7062 7220 7086
rect 7252 7086 7424 7088
rect 7222 7064 7250 7068
rect 7252 7064 7332 7086
rect 7353 7084 7368 7086
rect 7222 7062 7332 7064
rect 7153 7058 7332 7062
rect 7126 7048 7156 7058
rect 7158 7048 7311 7058
rect 7319 7048 7349 7058
rect 7353 7048 7383 7062
rect 7411 7048 7424 7086
rect 7496 7092 7531 7100
rect 7496 7066 7497 7092
rect 7504 7066 7531 7092
rect 7439 7048 7469 7062
rect 7496 7058 7531 7066
rect 7533 7092 7574 7100
rect 7533 7066 7548 7092
rect 7555 7066 7574 7092
rect 7638 7088 7700 7100
rect 7712 7088 7787 7100
rect 7845 7088 7920 7100
rect 7932 7088 7963 7100
rect 7969 7088 8004 7100
rect 7638 7086 7800 7088
rect 7533 7058 7574 7066
rect 7656 7062 7669 7086
rect 7684 7084 7699 7086
rect 7496 7048 7497 7058
rect 7512 7048 7525 7058
rect 7539 7048 7540 7058
rect 7555 7048 7568 7058
rect 7583 7048 7613 7062
rect 7656 7048 7699 7062
rect 7723 7059 7730 7066
rect 7733 7062 7800 7086
rect 7832 7086 8004 7088
rect 7802 7064 7830 7068
rect 7832 7064 7912 7086
rect 7933 7084 7948 7086
rect 7802 7062 7912 7064
rect 7733 7058 7912 7062
rect 7706 7048 7736 7058
rect 7738 7048 7891 7058
rect 7899 7048 7929 7058
rect 7933 7048 7963 7062
rect 7991 7048 8004 7086
rect 8076 7092 8111 7100
rect 8076 7066 8077 7092
rect 8084 7066 8111 7092
rect 8019 7048 8049 7062
rect 8076 7058 8111 7066
rect 8113 7092 8154 7100
rect 8113 7066 8128 7092
rect 8135 7066 8154 7092
rect 8218 7088 8280 7100
rect 8292 7088 8367 7100
rect 8425 7088 8500 7100
rect 8512 7088 8543 7100
rect 8549 7088 8584 7100
rect 8218 7086 8380 7088
rect 8113 7058 8154 7066
rect 8236 7062 8249 7086
rect 8264 7084 8279 7086
rect 8076 7048 8077 7058
rect 8092 7048 8105 7058
rect 8119 7048 8120 7058
rect 8135 7048 8148 7058
rect 8163 7048 8193 7062
rect 8236 7048 8279 7062
rect 8303 7059 8310 7066
rect 8313 7062 8380 7086
rect 8412 7086 8584 7088
rect 8382 7064 8410 7068
rect 8412 7064 8492 7086
rect 8513 7084 8528 7086
rect 8382 7062 8492 7064
rect 8313 7058 8492 7062
rect 8286 7048 8316 7058
rect 8318 7048 8471 7058
rect 8479 7048 8509 7058
rect 8513 7048 8543 7062
rect 8571 7048 8584 7086
rect 8656 7092 8691 7100
rect 8656 7066 8657 7092
rect 8664 7066 8691 7092
rect 8599 7048 8629 7062
rect 8656 7058 8691 7066
rect 8693 7092 8734 7100
rect 8693 7066 8708 7092
rect 8715 7066 8734 7092
rect 8798 7088 8860 7100
rect 8872 7088 8947 7100
rect 9005 7088 9080 7100
rect 9092 7088 9123 7100
rect 9129 7088 9164 7100
rect 8798 7086 8960 7088
rect 8693 7058 8734 7066
rect 8816 7062 8829 7086
rect 8844 7084 8859 7086
rect 8656 7048 8657 7058
rect 8672 7048 8685 7058
rect 8699 7048 8700 7058
rect 8715 7048 8728 7058
rect 8743 7048 8773 7062
rect 8816 7048 8859 7062
rect 8883 7059 8890 7066
rect 8893 7062 8960 7086
rect 8992 7086 9164 7088
rect 8962 7064 8990 7068
rect 8992 7064 9072 7086
rect 9093 7084 9108 7086
rect 8962 7062 9072 7064
rect 8893 7058 9072 7062
rect 8866 7048 8896 7058
rect 8898 7048 9051 7058
rect 9059 7048 9089 7058
rect 9093 7048 9123 7062
rect 9151 7048 9164 7086
rect 9236 7092 9271 7100
rect 9236 7066 9237 7092
rect 9244 7066 9271 7092
rect 9179 7048 9209 7062
rect 9236 7058 9271 7066
rect 9236 7048 9237 7058
rect 9252 7048 9265 7058
rect -1 7042 9265 7048
rect 0 7034 9265 7042
rect 15 7004 28 7034
rect 43 7016 73 7034
rect 116 7020 130 7034
rect 166 7020 386 7034
rect 117 7018 130 7020
rect 83 7006 98 7018
rect 80 7004 102 7006
rect 107 7004 137 7018
rect 198 7016 351 7020
rect 180 7004 372 7016
rect 415 7004 445 7018
rect 451 7004 464 7034
rect 479 7016 509 7034
rect 552 7004 565 7034
rect 595 7004 608 7034
rect 623 7016 653 7034
rect 696 7020 710 7034
rect 746 7020 966 7034
rect 697 7018 710 7020
rect 663 7006 678 7018
rect 660 7004 682 7006
rect 687 7004 717 7018
rect 778 7016 931 7020
rect 760 7004 952 7016
rect 995 7004 1025 7018
rect 1031 7004 1044 7034
rect 1059 7016 1089 7034
rect 1132 7004 1145 7034
rect 1175 7004 1188 7034
rect 1203 7016 1233 7034
rect 1276 7020 1290 7034
rect 1326 7020 1546 7034
rect 1277 7018 1290 7020
rect 1243 7006 1258 7018
rect 1240 7004 1262 7006
rect 1267 7004 1297 7018
rect 1358 7016 1511 7020
rect 1340 7004 1532 7016
rect 1575 7004 1605 7018
rect 1611 7004 1624 7034
rect 1639 7016 1669 7034
rect 1712 7004 1725 7034
rect 1755 7004 1768 7034
rect 1783 7016 1813 7034
rect 1856 7020 1870 7034
rect 1906 7020 2126 7034
rect 1857 7018 1870 7020
rect 1823 7006 1838 7018
rect 1820 7004 1842 7006
rect 1847 7004 1877 7018
rect 1938 7016 2091 7020
rect 1920 7004 2112 7016
rect 2155 7004 2185 7018
rect 2191 7004 2204 7034
rect 2219 7016 2249 7034
rect 2292 7004 2305 7034
rect 2335 7004 2348 7034
rect 2363 7016 2393 7034
rect 2436 7020 2450 7034
rect 2486 7020 2706 7034
rect 2437 7018 2450 7020
rect 2403 7006 2418 7018
rect 2400 7004 2422 7006
rect 2427 7004 2457 7018
rect 2518 7016 2671 7020
rect 2500 7004 2692 7016
rect 2735 7004 2765 7018
rect 2771 7004 2784 7034
rect 2799 7016 2829 7034
rect 2872 7004 2885 7034
rect 2915 7004 2928 7034
rect 2943 7016 2973 7034
rect 3016 7020 3030 7034
rect 3066 7020 3286 7034
rect 3017 7018 3030 7020
rect 2983 7006 2998 7018
rect 2980 7004 3002 7006
rect 3007 7004 3037 7018
rect 3098 7016 3251 7020
rect 3080 7004 3272 7016
rect 3315 7004 3345 7018
rect 3351 7004 3364 7034
rect 3379 7016 3409 7034
rect 3452 7004 3465 7034
rect 3495 7004 3508 7034
rect 3523 7016 3553 7034
rect 3596 7020 3610 7034
rect 3646 7020 3866 7034
rect 3597 7018 3610 7020
rect 3563 7006 3578 7018
rect 3560 7004 3582 7006
rect 3587 7004 3617 7018
rect 3678 7016 3831 7020
rect 3660 7004 3852 7016
rect 3895 7004 3925 7018
rect 3931 7004 3944 7034
rect 3959 7016 3989 7034
rect 4032 7004 4045 7034
rect 4075 7004 4088 7034
rect 4103 7016 4133 7034
rect 4176 7020 4190 7034
rect 4226 7020 4446 7034
rect 4177 7018 4190 7020
rect 4143 7006 4158 7018
rect 4140 7004 4162 7006
rect 4167 7004 4197 7018
rect 4258 7016 4411 7020
rect 4240 7004 4432 7016
rect 4475 7004 4505 7018
rect 4511 7004 4524 7034
rect 4539 7016 4569 7034
rect 4612 7004 4625 7034
rect 4655 7004 4668 7034
rect 4683 7016 4713 7034
rect 4756 7020 4770 7034
rect 4806 7020 5026 7034
rect 4757 7018 4770 7020
rect 4723 7006 4738 7018
rect 4720 7004 4742 7006
rect 4747 7004 4777 7018
rect 4838 7016 4991 7020
rect 4820 7004 5012 7016
rect 5055 7004 5085 7018
rect 5091 7004 5104 7034
rect 5119 7016 5149 7034
rect 5192 7004 5205 7034
rect 5235 7004 5248 7034
rect 5263 7016 5293 7034
rect 5336 7020 5350 7034
rect 5386 7020 5606 7034
rect 5337 7018 5350 7020
rect 5303 7006 5318 7018
rect 5300 7004 5322 7006
rect 5327 7004 5357 7018
rect 5418 7016 5571 7020
rect 5400 7004 5592 7016
rect 5635 7004 5665 7018
rect 5671 7004 5684 7034
rect 5699 7016 5729 7034
rect 5772 7004 5785 7034
rect 5815 7004 5828 7034
rect 5843 7016 5873 7034
rect 5916 7020 5930 7034
rect 5966 7020 6186 7034
rect 5917 7018 5930 7020
rect 5883 7006 5898 7018
rect 5880 7004 5902 7006
rect 5907 7004 5937 7018
rect 5998 7016 6151 7020
rect 5980 7004 6172 7016
rect 6215 7004 6245 7018
rect 6251 7004 6264 7034
rect 6279 7016 6309 7034
rect 6352 7004 6365 7034
rect 6395 7004 6408 7034
rect 6423 7016 6453 7034
rect 6496 7020 6510 7034
rect 6546 7020 6766 7034
rect 6497 7018 6510 7020
rect 6463 7006 6478 7018
rect 6460 7004 6482 7006
rect 6487 7004 6517 7018
rect 6578 7016 6731 7020
rect 6560 7004 6752 7016
rect 6795 7004 6825 7018
rect 6831 7004 6844 7034
rect 6859 7016 6889 7034
rect 6932 7004 6945 7034
rect 6975 7004 6988 7034
rect 7003 7016 7033 7034
rect 7076 7020 7090 7034
rect 7126 7020 7346 7034
rect 7077 7018 7090 7020
rect 7043 7006 7058 7018
rect 7040 7004 7062 7006
rect 7067 7004 7097 7018
rect 7158 7016 7311 7020
rect 7140 7004 7332 7016
rect 7375 7004 7405 7018
rect 7411 7004 7424 7034
rect 7439 7016 7469 7034
rect 7512 7004 7525 7034
rect 7555 7004 7568 7034
rect 7583 7016 7613 7034
rect 7656 7020 7670 7034
rect 7706 7020 7926 7034
rect 7657 7018 7670 7020
rect 7623 7006 7638 7018
rect 7620 7004 7642 7006
rect 7647 7004 7677 7018
rect 7738 7016 7891 7020
rect 7720 7004 7912 7016
rect 7955 7004 7985 7018
rect 7991 7004 8004 7034
rect 8019 7016 8049 7034
rect 8092 7004 8105 7034
rect 8135 7004 8148 7034
rect 8163 7016 8193 7034
rect 8236 7020 8250 7034
rect 8286 7020 8506 7034
rect 8237 7018 8250 7020
rect 8203 7006 8218 7018
rect 8200 7004 8222 7006
rect 8227 7004 8257 7018
rect 8318 7016 8471 7020
rect 8300 7004 8492 7016
rect 8535 7004 8565 7018
rect 8571 7004 8584 7034
rect 8599 7016 8629 7034
rect 8672 7004 8685 7034
rect 8715 7004 8728 7034
rect 8743 7016 8773 7034
rect 8816 7020 8830 7034
rect 8866 7020 9086 7034
rect 8817 7018 8830 7020
rect 8783 7006 8798 7018
rect 8780 7004 8802 7006
rect 8807 7004 8837 7018
rect 8898 7016 9051 7020
rect 8880 7004 9072 7016
rect 9115 7004 9145 7018
rect 9151 7004 9164 7034
rect 9179 7016 9209 7034
rect 9252 7004 9265 7034
rect 0 6990 9265 7004
rect 15 6886 28 6990
rect 73 6968 74 6978
rect 89 6968 102 6978
rect 73 6964 102 6968
rect 107 6964 137 6990
rect 155 6976 171 6978
rect 243 6976 296 6990
rect 244 6974 308 6976
rect 351 6974 366 6990
rect 415 6987 445 6990
rect 415 6984 451 6987
rect 381 6976 397 6978
rect 155 6964 170 6968
rect 73 6962 170 6964
rect 198 6962 366 6974
rect 382 6964 397 6968
rect 415 6965 454 6984
rect 473 6978 480 6979
rect 479 6971 480 6978
rect 463 6968 464 6971
rect 479 6968 492 6971
rect 415 6964 445 6965
rect 454 6964 460 6965
rect 463 6964 492 6968
rect 382 6963 492 6964
rect 382 6962 498 6963
rect 57 6954 108 6962
rect 57 6942 82 6954
rect 89 6942 108 6954
rect 139 6954 189 6962
rect 139 6946 155 6954
rect 162 6952 189 6954
rect 198 6952 419 6962
rect 162 6942 419 6952
rect 448 6954 498 6962
rect 448 6945 464 6954
rect 57 6934 108 6942
rect 155 6934 419 6942
rect 445 6942 464 6945
rect 471 6942 498 6954
rect 445 6934 498 6942
rect 73 6926 74 6934
rect 89 6926 102 6934
rect 73 6918 89 6926
rect 70 6911 89 6914
rect 70 6902 92 6911
rect 43 6892 92 6902
rect 43 6886 73 6892
rect 92 6887 97 6892
rect 15 6870 89 6886
rect 107 6878 137 6934
rect 172 6924 380 6934
rect 415 6930 460 6934
rect 463 6933 464 6934
rect 479 6933 492 6934
rect 198 6894 387 6924
rect 213 6891 387 6894
rect 206 6888 387 6891
rect 15 6868 28 6870
rect 43 6868 77 6870
rect 15 6852 89 6868
rect 116 6864 129 6878
rect 144 6864 160 6880
rect 206 6875 217 6888
rect -1 6830 0 6846
rect 15 6830 28 6852
rect 43 6830 73 6852
rect 116 6848 178 6864
rect 206 6857 217 6873
rect 222 6868 232 6888
rect 242 6868 256 6888
rect 259 6875 268 6888
rect 284 6875 293 6888
rect 222 6857 256 6868
rect 259 6857 268 6873
rect 284 6857 293 6873
rect 300 6868 310 6888
rect 320 6868 334 6888
rect 335 6875 346 6888
rect 300 6857 334 6868
rect 335 6857 346 6873
rect 392 6864 408 6880
rect 415 6878 445 6930
rect 479 6926 480 6933
rect 464 6918 480 6926
rect 451 6886 464 6905
rect 479 6886 509 6902
rect 451 6870 525 6886
rect 451 6868 464 6870
rect 479 6868 513 6870
rect 116 6846 129 6848
rect 144 6846 178 6848
rect 116 6830 178 6846
rect 222 6841 238 6844
rect 300 6841 330 6852
rect 378 6848 424 6864
rect 451 6852 525 6868
rect 378 6846 412 6848
rect 377 6830 424 6846
rect 451 6830 464 6852
rect 479 6830 509 6852
rect 536 6830 537 6846
rect 552 6830 565 6990
rect 595 6886 608 6990
rect 653 6968 654 6978
rect 669 6968 682 6978
rect 653 6964 682 6968
rect 687 6964 717 6990
rect 735 6976 751 6978
rect 823 6976 876 6990
rect 824 6974 888 6976
rect 931 6974 946 6990
rect 995 6987 1025 6990
rect 995 6984 1031 6987
rect 961 6976 977 6978
rect 735 6964 750 6968
rect 653 6962 750 6964
rect 778 6962 946 6974
rect 962 6964 977 6968
rect 995 6965 1034 6984
rect 1053 6978 1060 6979
rect 1059 6971 1060 6978
rect 1043 6968 1044 6971
rect 1059 6968 1072 6971
rect 995 6964 1025 6965
rect 1034 6964 1040 6965
rect 1043 6964 1072 6968
rect 962 6963 1072 6964
rect 962 6962 1078 6963
rect 637 6954 688 6962
rect 637 6942 662 6954
rect 669 6942 688 6954
rect 719 6954 769 6962
rect 719 6946 735 6954
rect 742 6952 769 6954
rect 778 6952 999 6962
rect 742 6942 999 6952
rect 1028 6954 1078 6962
rect 1028 6945 1044 6954
rect 637 6934 688 6942
rect 735 6934 999 6942
rect 1025 6942 1044 6945
rect 1051 6942 1078 6954
rect 1025 6934 1078 6942
rect 653 6926 654 6934
rect 669 6926 682 6934
rect 653 6918 669 6926
rect 650 6911 669 6914
rect 650 6902 672 6911
rect 623 6892 672 6902
rect 623 6886 653 6892
rect 672 6887 677 6892
rect 595 6870 669 6886
rect 687 6878 717 6934
rect 752 6924 960 6934
rect 995 6930 1040 6934
rect 1043 6933 1044 6934
rect 1059 6933 1072 6934
rect 778 6894 967 6924
rect 793 6891 967 6894
rect 786 6888 967 6891
rect 595 6868 608 6870
rect 623 6868 657 6870
rect 595 6852 669 6868
rect 696 6864 709 6878
rect 724 6864 740 6880
rect 786 6875 797 6888
rect 579 6830 580 6846
rect 595 6830 608 6852
rect 623 6830 653 6852
rect 696 6848 758 6864
rect 786 6857 797 6873
rect 802 6868 812 6888
rect 822 6868 836 6888
rect 839 6875 848 6888
rect 864 6875 873 6888
rect 802 6857 836 6868
rect 839 6857 848 6873
rect 864 6857 873 6873
rect 880 6868 890 6888
rect 900 6868 914 6888
rect 915 6875 926 6888
rect 880 6857 914 6868
rect 915 6857 926 6873
rect 972 6864 988 6880
rect 995 6878 1025 6930
rect 1059 6926 1060 6933
rect 1044 6918 1060 6926
rect 1031 6886 1044 6905
rect 1059 6886 1089 6902
rect 1031 6870 1105 6886
rect 1031 6868 1044 6870
rect 1059 6868 1093 6870
rect 696 6846 709 6848
rect 724 6846 758 6848
rect 696 6830 758 6846
rect 802 6841 818 6844
rect 880 6841 910 6852
rect 958 6848 1004 6864
rect 1031 6852 1105 6868
rect 958 6846 992 6848
rect 957 6830 1004 6846
rect 1031 6830 1044 6852
rect 1059 6830 1089 6852
rect 1116 6830 1117 6846
rect 1132 6830 1145 6990
rect 1175 6886 1188 6990
rect 1233 6968 1234 6978
rect 1249 6968 1262 6978
rect 1233 6964 1262 6968
rect 1267 6964 1297 6990
rect 1315 6976 1331 6978
rect 1403 6976 1456 6990
rect 1404 6974 1468 6976
rect 1511 6974 1526 6990
rect 1575 6987 1605 6990
rect 1575 6984 1611 6987
rect 1541 6976 1557 6978
rect 1315 6964 1330 6968
rect 1233 6962 1330 6964
rect 1358 6962 1526 6974
rect 1542 6964 1557 6968
rect 1575 6965 1614 6984
rect 1633 6978 1640 6979
rect 1639 6971 1640 6978
rect 1623 6968 1624 6971
rect 1639 6968 1652 6971
rect 1575 6964 1605 6965
rect 1614 6964 1620 6965
rect 1623 6964 1652 6968
rect 1542 6963 1652 6964
rect 1542 6962 1658 6963
rect 1217 6954 1268 6962
rect 1217 6942 1242 6954
rect 1249 6942 1268 6954
rect 1299 6954 1349 6962
rect 1299 6946 1315 6954
rect 1322 6952 1349 6954
rect 1358 6952 1579 6962
rect 1322 6942 1579 6952
rect 1608 6954 1658 6962
rect 1608 6945 1624 6954
rect 1217 6934 1268 6942
rect 1315 6934 1579 6942
rect 1605 6942 1624 6945
rect 1631 6942 1658 6954
rect 1605 6934 1658 6942
rect 1233 6926 1234 6934
rect 1249 6926 1262 6934
rect 1233 6918 1249 6926
rect 1230 6911 1249 6914
rect 1230 6902 1252 6911
rect 1203 6892 1252 6902
rect 1203 6886 1233 6892
rect 1252 6887 1257 6892
rect 1175 6870 1249 6886
rect 1267 6878 1297 6934
rect 1332 6924 1540 6934
rect 1575 6930 1620 6934
rect 1623 6933 1624 6934
rect 1639 6933 1652 6934
rect 1358 6894 1547 6924
rect 1373 6891 1547 6894
rect 1366 6888 1547 6891
rect 1175 6868 1188 6870
rect 1203 6868 1237 6870
rect 1175 6852 1249 6868
rect 1276 6864 1289 6878
rect 1304 6864 1320 6880
rect 1366 6875 1377 6888
rect 1159 6830 1160 6846
rect 1175 6830 1188 6852
rect 1203 6830 1233 6852
rect 1276 6848 1338 6864
rect 1366 6857 1377 6873
rect 1382 6868 1392 6888
rect 1402 6868 1416 6888
rect 1419 6875 1428 6888
rect 1444 6875 1453 6888
rect 1382 6857 1416 6868
rect 1419 6857 1428 6873
rect 1444 6857 1453 6873
rect 1460 6868 1470 6888
rect 1480 6868 1494 6888
rect 1495 6875 1506 6888
rect 1460 6857 1494 6868
rect 1495 6857 1506 6873
rect 1552 6864 1568 6880
rect 1575 6878 1605 6930
rect 1639 6926 1640 6933
rect 1624 6918 1640 6926
rect 1611 6886 1624 6905
rect 1639 6886 1669 6902
rect 1611 6870 1685 6886
rect 1611 6868 1624 6870
rect 1639 6868 1673 6870
rect 1276 6846 1289 6848
rect 1304 6846 1338 6848
rect 1276 6830 1338 6846
rect 1382 6841 1398 6844
rect 1460 6841 1490 6852
rect 1538 6848 1584 6864
rect 1611 6852 1685 6868
rect 1538 6846 1572 6848
rect 1537 6830 1584 6846
rect 1611 6830 1624 6852
rect 1639 6830 1669 6852
rect 1696 6830 1697 6846
rect 1712 6830 1725 6990
rect 1755 6886 1768 6990
rect 1813 6968 1814 6978
rect 1829 6968 1842 6978
rect 1813 6964 1842 6968
rect 1847 6964 1877 6990
rect 1895 6976 1911 6978
rect 1983 6976 2036 6990
rect 1984 6974 2048 6976
rect 2091 6974 2106 6990
rect 2155 6987 2185 6990
rect 2155 6984 2191 6987
rect 2121 6976 2137 6978
rect 1895 6964 1910 6968
rect 1813 6962 1910 6964
rect 1938 6962 2106 6974
rect 2122 6964 2137 6968
rect 2155 6965 2194 6984
rect 2213 6978 2220 6979
rect 2219 6971 2220 6978
rect 2203 6968 2204 6971
rect 2219 6968 2232 6971
rect 2155 6964 2185 6965
rect 2194 6964 2200 6965
rect 2203 6964 2232 6968
rect 2122 6963 2232 6964
rect 2122 6962 2238 6963
rect 1797 6954 1848 6962
rect 1797 6942 1822 6954
rect 1829 6942 1848 6954
rect 1879 6954 1929 6962
rect 1879 6946 1895 6954
rect 1902 6952 1929 6954
rect 1938 6952 2159 6962
rect 1902 6942 2159 6952
rect 2188 6954 2238 6962
rect 2188 6945 2204 6954
rect 1797 6934 1848 6942
rect 1895 6934 2159 6942
rect 2185 6942 2204 6945
rect 2211 6942 2238 6954
rect 2185 6934 2238 6942
rect 1813 6926 1814 6934
rect 1829 6926 1842 6934
rect 1813 6918 1829 6926
rect 1810 6911 1829 6914
rect 1810 6902 1832 6911
rect 1783 6892 1832 6902
rect 1783 6886 1813 6892
rect 1832 6887 1837 6892
rect 1755 6870 1829 6886
rect 1847 6878 1877 6934
rect 1912 6924 2120 6934
rect 2155 6930 2200 6934
rect 2203 6933 2204 6934
rect 2219 6933 2232 6934
rect 1938 6894 2127 6924
rect 1953 6891 2127 6894
rect 1946 6888 2127 6891
rect 1755 6868 1768 6870
rect 1783 6868 1817 6870
rect 1755 6852 1829 6868
rect 1856 6864 1869 6878
rect 1884 6864 1900 6880
rect 1946 6875 1957 6888
rect 1739 6830 1740 6846
rect 1755 6830 1768 6852
rect 1783 6830 1813 6852
rect 1856 6848 1918 6864
rect 1946 6857 1957 6873
rect 1962 6868 1972 6888
rect 1982 6868 1996 6888
rect 1999 6875 2008 6888
rect 2024 6875 2033 6888
rect 1962 6857 1996 6868
rect 1999 6857 2008 6873
rect 2024 6857 2033 6873
rect 2040 6868 2050 6888
rect 2060 6868 2074 6888
rect 2075 6875 2086 6888
rect 2040 6857 2074 6868
rect 2075 6857 2086 6873
rect 2132 6864 2148 6880
rect 2155 6878 2185 6930
rect 2219 6926 2220 6933
rect 2204 6918 2220 6926
rect 2191 6886 2204 6905
rect 2219 6886 2249 6902
rect 2191 6870 2265 6886
rect 2191 6868 2204 6870
rect 2219 6868 2253 6870
rect 1856 6846 1869 6848
rect 1884 6846 1918 6848
rect 1856 6830 1918 6846
rect 1962 6841 1976 6844
rect 2040 6841 2070 6852
rect 2118 6848 2164 6864
rect 2191 6852 2265 6868
rect 2118 6846 2152 6848
rect 2117 6830 2164 6846
rect 2191 6830 2204 6852
rect 2219 6830 2249 6852
rect 2276 6830 2277 6846
rect 2292 6830 2305 6990
rect 2335 6886 2348 6990
rect 2393 6968 2394 6978
rect 2409 6968 2422 6978
rect 2393 6964 2422 6968
rect 2427 6964 2457 6990
rect 2475 6976 2491 6978
rect 2563 6976 2616 6990
rect 2564 6974 2628 6976
rect 2671 6974 2686 6990
rect 2735 6987 2765 6990
rect 2735 6984 2771 6987
rect 2701 6976 2717 6978
rect 2475 6964 2490 6968
rect 2393 6962 2490 6964
rect 2518 6962 2686 6974
rect 2702 6964 2717 6968
rect 2735 6965 2774 6984
rect 2793 6978 2800 6979
rect 2799 6971 2800 6978
rect 2783 6968 2784 6971
rect 2799 6968 2812 6971
rect 2735 6964 2765 6965
rect 2774 6964 2780 6965
rect 2783 6964 2812 6968
rect 2702 6963 2812 6964
rect 2702 6962 2818 6963
rect 2377 6954 2428 6962
rect 2377 6942 2402 6954
rect 2409 6942 2428 6954
rect 2459 6954 2509 6962
rect 2459 6946 2475 6954
rect 2482 6952 2509 6954
rect 2518 6952 2739 6962
rect 2482 6942 2739 6952
rect 2768 6954 2818 6962
rect 2768 6945 2784 6954
rect 2377 6934 2428 6942
rect 2475 6934 2739 6942
rect 2765 6942 2784 6945
rect 2791 6942 2818 6954
rect 2765 6934 2818 6942
rect 2393 6926 2394 6934
rect 2409 6926 2422 6934
rect 2393 6918 2409 6926
rect 2390 6911 2409 6914
rect 2390 6902 2412 6911
rect 2363 6892 2412 6902
rect 2363 6886 2393 6892
rect 2412 6887 2417 6892
rect 2335 6870 2409 6886
rect 2427 6878 2457 6934
rect 2492 6924 2700 6934
rect 2735 6930 2780 6934
rect 2783 6933 2784 6934
rect 2799 6933 2812 6934
rect 2518 6894 2707 6924
rect 2533 6891 2707 6894
rect 2526 6888 2707 6891
rect 2335 6868 2348 6870
rect 2363 6868 2397 6870
rect 2335 6852 2409 6868
rect 2436 6864 2449 6878
rect 2464 6864 2480 6880
rect 2526 6875 2537 6888
rect 2319 6830 2320 6846
rect 2335 6830 2348 6852
rect 2363 6830 2393 6852
rect 2436 6848 2498 6864
rect 2526 6857 2537 6873
rect 2542 6868 2552 6888
rect 2562 6868 2576 6888
rect 2579 6875 2588 6888
rect 2604 6875 2613 6888
rect 2542 6857 2576 6868
rect 2579 6857 2588 6873
rect 2604 6857 2613 6873
rect 2620 6868 2630 6888
rect 2640 6868 2654 6888
rect 2655 6875 2666 6888
rect 2620 6857 2654 6868
rect 2655 6857 2666 6873
rect 2712 6864 2728 6880
rect 2735 6878 2765 6930
rect 2799 6926 2800 6933
rect 2784 6918 2800 6926
rect 2771 6886 2784 6905
rect 2799 6886 2829 6902
rect 2771 6870 2845 6886
rect 2771 6868 2784 6870
rect 2799 6868 2833 6870
rect 2436 6846 2449 6848
rect 2464 6846 2498 6848
rect 2436 6830 2498 6846
rect 2542 6841 2558 6844
rect 2620 6841 2650 6852
rect 2698 6848 2744 6864
rect 2771 6852 2845 6868
rect 2698 6846 2732 6848
rect 2697 6830 2744 6846
rect 2771 6830 2784 6852
rect 2799 6830 2829 6852
rect 2856 6830 2857 6846
rect 2872 6830 2885 6990
rect 2915 6886 2928 6990
rect 2973 6968 2974 6978
rect 2989 6968 3002 6978
rect 2973 6964 3002 6968
rect 3007 6964 3037 6990
rect 3055 6976 3071 6978
rect 3143 6976 3196 6990
rect 3144 6974 3208 6976
rect 3251 6974 3266 6990
rect 3315 6987 3345 6990
rect 3315 6984 3351 6987
rect 3281 6976 3297 6978
rect 3055 6964 3070 6968
rect 2973 6962 3070 6964
rect 3098 6962 3266 6974
rect 3282 6964 3297 6968
rect 3315 6965 3354 6984
rect 3373 6978 3380 6979
rect 3379 6971 3380 6978
rect 3363 6968 3364 6971
rect 3379 6968 3392 6971
rect 3315 6964 3345 6965
rect 3354 6964 3360 6965
rect 3363 6964 3392 6968
rect 3282 6963 3392 6964
rect 3282 6962 3398 6963
rect 2957 6954 3008 6962
rect 2957 6942 2982 6954
rect 2989 6942 3008 6954
rect 3039 6954 3089 6962
rect 3039 6946 3055 6954
rect 3062 6952 3089 6954
rect 3098 6952 3319 6962
rect 3062 6942 3319 6952
rect 3348 6954 3398 6962
rect 3348 6945 3364 6954
rect 2957 6934 3008 6942
rect 3055 6934 3319 6942
rect 3345 6942 3364 6945
rect 3371 6942 3398 6954
rect 3345 6934 3398 6942
rect 2973 6926 2974 6934
rect 2989 6926 3002 6934
rect 2973 6918 2989 6926
rect 2970 6911 2989 6914
rect 2970 6902 2992 6911
rect 2943 6892 2992 6902
rect 2943 6886 2973 6892
rect 2992 6887 2997 6892
rect 2915 6870 2989 6886
rect 3007 6878 3037 6934
rect 3072 6924 3280 6934
rect 3315 6930 3360 6934
rect 3363 6933 3364 6934
rect 3379 6933 3392 6934
rect 3098 6894 3287 6924
rect 3113 6891 3287 6894
rect 3106 6888 3287 6891
rect 2915 6868 2928 6870
rect 2943 6868 2977 6870
rect 2915 6852 2989 6868
rect 3016 6864 3029 6878
rect 3044 6864 3060 6880
rect 3106 6875 3117 6888
rect 2899 6830 2900 6846
rect 2915 6830 2928 6852
rect 2943 6830 2973 6852
rect 3016 6848 3078 6864
rect 3106 6857 3117 6873
rect 3122 6868 3132 6888
rect 3142 6868 3156 6888
rect 3159 6875 3168 6888
rect 3184 6875 3193 6888
rect 3122 6857 3156 6868
rect 3159 6857 3168 6873
rect 3184 6857 3193 6873
rect 3200 6868 3210 6888
rect 3220 6868 3234 6888
rect 3235 6875 3246 6888
rect 3200 6857 3234 6868
rect 3235 6857 3246 6873
rect 3292 6864 3308 6880
rect 3315 6878 3345 6930
rect 3379 6926 3380 6933
rect 3364 6918 3380 6926
rect 3351 6886 3364 6905
rect 3379 6886 3409 6902
rect 3351 6870 3425 6886
rect 3351 6868 3364 6870
rect 3379 6868 3413 6870
rect 3016 6846 3029 6848
rect 3044 6846 3078 6848
rect 3016 6830 3078 6846
rect 3122 6841 3138 6844
rect 3200 6841 3230 6852
rect 3278 6848 3324 6864
rect 3351 6852 3425 6868
rect 3278 6846 3312 6848
rect 3277 6830 3324 6846
rect 3351 6830 3364 6852
rect 3379 6830 3409 6852
rect 3436 6830 3437 6846
rect 3452 6830 3465 6990
rect 3495 6886 3508 6990
rect 3553 6968 3554 6978
rect 3569 6968 3582 6978
rect 3553 6964 3582 6968
rect 3587 6964 3617 6990
rect 3635 6976 3651 6978
rect 3723 6976 3776 6990
rect 3724 6974 3788 6976
rect 3831 6974 3846 6990
rect 3895 6987 3925 6990
rect 3895 6984 3931 6987
rect 3861 6976 3877 6978
rect 3635 6964 3650 6968
rect 3553 6962 3650 6964
rect 3678 6962 3846 6974
rect 3862 6964 3877 6968
rect 3895 6965 3934 6984
rect 3953 6978 3960 6979
rect 3959 6971 3960 6978
rect 3943 6968 3944 6971
rect 3959 6968 3972 6971
rect 3895 6964 3925 6965
rect 3934 6964 3940 6965
rect 3943 6964 3972 6968
rect 3862 6963 3972 6964
rect 3862 6962 3978 6963
rect 3537 6954 3588 6962
rect 3537 6942 3562 6954
rect 3569 6942 3588 6954
rect 3619 6954 3669 6962
rect 3619 6946 3635 6954
rect 3642 6952 3669 6954
rect 3678 6952 3899 6962
rect 3642 6942 3899 6952
rect 3928 6954 3978 6962
rect 3928 6945 3944 6954
rect 3537 6934 3588 6942
rect 3635 6934 3899 6942
rect 3925 6942 3944 6945
rect 3951 6942 3978 6954
rect 3925 6934 3978 6942
rect 3553 6926 3554 6934
rect 3569 6926 3582 6934
rect 3553 6918 3569 6926
rect 3550 6911 3569 6914
rect 3550 6902 3572 6911
rect 3523 6892 3572 6902
rect 3523 6886 3553 6892
rect 3572 6887 3577 6892
rect 3495 6870 3569 6886
rect 3587 6878 3617 6934
rect 3652 6924 3860 6934
rect 3895 6930 3940 6934
rect 3943 6933 3944 6934
rect 3959 6933 3972 6934
rect 3678 6894 3867 6924
rect 3693 6891 3867 6894
rect 3686 6888 3867 6891
rect 3495 6868 3508 6870
rect 3523 6868 3557 6870
rect 3495 6852 3569 6868
rect 3596 6864 3609 6878
rect 3624 6864 3640 6880
rect 3686 6875 3697 6888
rect 3479 6830 3480 6846
rect 3495 6830 3508 6852
rect 3523 6830 3553 6852
rect 3596 6848 3658 6864
rect 3686 6857 3697 6873
rect 3702 6868 3712 6888
rect 3722 6868 3736 6888
rect 3739 6875 3748 6888
rect 3764 6875 3773 6888
rect 3702 6857 3736 6868
rect 3739 6857 3748 6873
rect 3764 6857 3773 6873
rect 3780 6868 3790 6888
rect 3800 6868 3814 6888
rect 3815 6875 3826 6888
rect 3780 6857 3814 6868
rect 3815 6857 3826 6873
rect 3872 6864 3888 6880
rect 3895 6878 3925 6930
rect 3959 6926 3960 6933
rect 3944 6918 3960 6926
rect 3931 6886 3944 6905
rect 3959 6886 3989 6902
rect 3931 6870 4005 6886
rect 3931 6868 3944 6870
rect 3959 6868 3993 6870
rect 3596 6846 3609 6848
rect 3624 6846 3658 6848
rect 3596 6830 3658 6846
rect 3702 6841 3718 6844
rect 3780 6841 3810 6852
rect 3858 6848 3904 6864
rect 3931 6852 4005 6868
rect 3858 6846 3892 6848
rect 3857 6830 3904 6846
rect 3931 6830 3944 6852
rect 3959 6830 3989 6852
rect 4016 6830 4017 6846
rect 4032 6830 4045 6990
rect 4075 6886 4088 6990
rect 4133 6968 4134 6978
rect 4149 6968 4162 6978
rect 4133 6964 4162 6968
rect 4167 6964 4197 6990
rect 4215 6976 4231 6978
rect 4303 6976 4356 6990
rect 4304 6974 4368 6976
rect 4411 6974 4426 6990
rect 4475 6987 4505 6990
rect 4475 6984 4511 6987
rect 4441 6976 4457 6978
rect 4215 6964 4230 6968
rect 4133 6962 4230 6964
rect 4258 6962 4426 6974
rect 4442 6964 4457 6968
rect 4475 6965 4514 6984
rect 4533 6978 4540 6979
rect 4539 6971 4540 6978
rect 4523 6968 4524 6971
rect 4539 6968 4552 6971
rect 4475 6964 4505 6965
rect 4514 6964 4520 6965
rect 4523 6964 4552 6968
rect 4442 6963 4552 6964
rect 4442 6962 4558 6963
rect 4117 6954 4168 6962
rect 4117 6942 4142 6954
rect 4149 6942 4168 6954
rect 4199 6954 4249 6962
rect 4199 6946 4215 6954
rect 4222 6952 4249 6954
rect 4258 6952 4479 6962
rect 4222 6942 4479 6952
rect 4508 6954 4558 6962
rect 4508 6945 4524 6954
rect 4117 6934 4168 6942
rect 4215 6934 4479 6942
rect 4505 6942 4524 6945
rect 4531 6942 4558 6954
rect 4505 6934 4558 6942
rect 4133 6926 4134 6934
rect 4149 6926 4162 6934
rect 4133 6918 4149 6926
rect 4130 6911 4149 6914
rect 4130 6902 4152 6911
rect 4103 6892 4152 6902
rect 4103 6886 4133 6892
rect 4152 6887 4157 6892
rect 4075 6870 4149 6886
rect 4167 6878 4197 6934
rect 4232 6924 4440 6934
rect 4475 6930 4520 6934
rect 4523 6933 4524 6934
rect 4539 6933 4552 6934
rect 4258 6894 4447 6924
rect 4273 6891 4447 6894
rect 4266 6888 4447 6891
rect 4075 6868 4088 6870
rect 4103 6868 4137 6870
rect 4075 6852 4149 6868
rect 4176 6864 4189 6878
rect 4204 6864 4220 6880
rect 4266 6875 4277 6888
rect 4059 6830 4060 6846
rect 4075 6830 4088 6852
rect 4103 6830 4133 6852
rect 4176 6848 4238 6864
rect 4266 6857 4277 6873
rect 4282 6868 4292 6888
rect 4302 6868 4316 6888
rect 4319 6875 4328 6888
rect 4344 6875 4353 6888
rect 4282 6857 4316 6868
rect 4319 6857 4328 6873
rect 4344 6857 4353 6873
rect 4360 6868 4370 6888
rect 4380 6868 4394 6888
rect 4395 6875 4406 6888
rect 4360 6857 4394 6868
rect 4395 6857 4406 6873
rect 4452 6864 4468 6880
rect 4475 6878 4505 6930
rect 4539 6926 4540 6933
rect 4524 6918 4540 6926
rect 4511 6886 4524 6905
rect 4539 6886 4569 6902
rect 4511 6870 4585 6886
rect 4511 6868 4524 6870
rect 4539 6868 4573 6870
rect 4176 6846 4189 6848
rect 4204 6846 4238 6848
rect 4176 6830 4238 6846
rect 4282 6841 4298 6844
rect 4360 6841 4390 6852
rect 4438 6848 4484 6864
rect 4511 6852 4585 6868
rect 4438 6846 4472 6848
rect 4437 6830 4484 6846
rect 4511 6830 4524 6852
rect 4539 6830 4569 6852
rect 4596 6830 4597 6846
rect 4612 6830 4625 6990
rect 4655 6886 4668 6990
rect 4713 6968 4714 6978
rect 4729 6968 4742 6978
rect 4713 6964 4742 6968
rect 4747 6964 4777 6990
rect 4795 6976 4811 6978
rect 4883 6976 4936 6990
rect 4884 6974 4948 6976
rect 4991 6974 5006 6990
rect 5055 6987 5085 6990
rect 5055 6984 5091 6987
rect 5021 6976 5037 6978
rect 4795 6964 4810 6968
rect 4713 6962 4810 6964
rect 4838 6962 5006 6974
rect 5022 6964 5037 6968
rect 5055 6965 5094 6984
rect 5113 6978 5120 6979
rect 5119 6971 5120 6978
rect 5103 6968 5104 6971
rect 5119 6968 5132 6971
rect 5055 6964 5085 6965
rect 5094 6964 5100 6965
rect 5103 6964 5132 6968
rect 5022 6963 5132 6964
rect 5022 6962 5138 6963
rect 4697 6954 4748 6962
rect 4697 6942 4722 6954
rect 4729 6942 4748 6954
rect 4779 6954 4829 6962
rect 4779 6946 4795 6954
rect 4802 6952 4829 6954
rect 4838 6952 5059 6962
rect 4802 6942 5059 6952
rect 5088 6954 5138 6962
rect 5088 6945 5104 6954
rect 4697 6934 4748 6942
rect 4795 6934 5059 6942
rect 5085 6942 5104 6945
rect 5111 6942 5138 6954
rect 5085 6934 5138 6942
rect 4713 6926 4714 6934
rect 4729 6926 4742 6934
rect 4713 6918 4729 6926
rect 4710 6911 4729 6914
rect 4710 6902 4732 6911
rect 4683 6892 4732 6902
rect 4683 6886 4713 6892
rect 4732 6887 4737 6892
rect 4655 6870 4729 6886
rect 4747 6878 4777 6934
rect 4812 6924 5020 6934
rect 5055 6930 5100 6934
rect 5103 6933 5104 6934
rect 5119 6933 5132 6934
rect 4838 6894 5027 6924
rect 4853 6891 5027 6894
rect 4846 6888 5027 6891
rect 4655 6868 4668 6870
rect 4683 6868 4717 6870
rect 4655 6852 4729 6868
rect 4756 6864 4769 6878
rect 4784 6864 4800 6880
rect 4846 6875 4857 6888
rect 4639 6830 4640 6846
rect 4655 6830 4668 6852
rect 4683 6830 4713 6852
rect 4756 6848 4818 6864
rect 4846 6857 4857 6873
rect 4862 6868 4872 6888
rect 4882 6868 4896 6888
rect 4899 6875 4908 6888
rect 4924 6875 4933 6888
rect 4862 6857 4896 6868
rect 4899 6857 4908 6873
rect 4924 6857 4933 6873
rect 4940 6868 4950 6888
rect 4960 6868 4974 6888
rect 4975 6875 4986 6888
rect 4940 6857 4974 6868
rect 4975 6857 4986 6873
rect 5032 6864 5048 6880
rect 5055 6878 5085 6930
rect 5119 6926 5120 6933
rect 5104 6918 5120 6926
rect 5091 6886 5104 6905
rect 5119 6886 5149 6902
rect 5091 6870 5165 6886
rect 5091 6868 5104 6870
rect 5119 6868 5153 6870
rect 4756 6846 4769 6848
rect 4784 6846 4818 6848
rect 4756 6830 4818 6846
rect 4862 6841 4878 6844
rect 4940 6841 4970 6852
rect 5018 6848 5064 6864
rect 5091 6852 5165 6868
rect 5018 6846 5052 6848
rect 5017 6830 5064 6846
rect 5091 6830 5104 6852
rect 5119 6830 5149 6852
rect 5176 6830 5177 6846
rect 5192 6830 5205 6990
rect 5235 6886 5248 6990
rect 5293 6968 5294 6978
rect 5309 6968 5322 6978
rect 5293 6964 5322 6968
rect 5327 6964 5357 6990
rect 5375 6976 5391 6978
rect 5463 6976 5516 6990
rect 5464 6974 5528 6976
rect 5571 6974 5586 6990
rect 5635 6987 5665 6990
rect 5635 6984 5671 6987
rect 5601 6976 5617 6978
rect 5375 6964 5390 6968
rect 5293 6962 5390 6964
rect 5418 6962 5586 6974
rect 5602 6964 5617 6968
rect 5635 6965 5674 6984
rect 5693 6978 5700 6979
rect 5699 6971 5700 6978
rect 5683 6968 5684 6971
rect 5699 6968 5712 6971
rect 5635 6964 5665 6965
rect 5674 6964 5680 6965
rect 5683 6964 5712 6968
rect 5602 6963 5712 6964
rect 5602 6962 5718 6963
rect 5277 6954 5328 6962
rect 5277 6942 5302 6954
rect 5309 6942 5328 6954
rect 5359 6954 5409 6962
rect 5359 6946 5375 6954
rect 5382 6952 5409 6954
rect 5418 6952 5639 6962
rect 5382 6942 5639 6952
rect 5668 6954 5718 6962
rect 5668 6945 5684 6954
rect 5277 6934 5328 6942
rect 5375 6934 5639 6942
rect 5665 6942 5684 6945
rect 5691 6942 5718 6954
rect 5665 6934 5718 6942
rect 5293 6926 5294 6934
rect 5309 6926 5322 6934
rect 5293 6918 5309 6926
rect 5290 6911 5309 6914
rect 5290 6902 5312 6911
rect 5263 6892 5312 6902
rect 5263 6886 5293 6892
rect 5312 6887 5317 6892
rect 5235 6870 5309 6886
rect 5327 6878 5357 6934
rect 5392 6924 5600 6934
rect 5635 6930 5680 6934
rect 5683 6933 5684 6934
rect 5699 6933 5712 6934
rect 5418 6894 5607 6924
rect 5433 6891 5607 6894
rect 5426 6888 5607 6891
rect 5235 6868 5248 6870
rect 5263 6868 5297 6870
rect 5235 6852 5309 6868
rect 5336 6864 5349 6878
rect 5364 6864 5380 6880
rect 5426 6875 5437 6888
rect 5219 6830 5220 6846
rect 5235 6830 5248 6852
rect 5263 6830 5293 6852
rect 5336 6848 5398 6864
rect 5426 6857 5437 6873
rect 5442 6868 5452 6888
rect 5462 6868 5476 6888
rect 5479 6875 5488 6888
rect 5504 6875 5513 6888
rect 5442 6857 5476 6868
rect 5479 6857 5488 6873
rect 5504 6857 5513 6873
rect 5520 6868 5530 6888
rect 5540 6868 5554 6888
rect 5555 6875 5566 6888
rect 5520 6857 5554 6868
rect 5555 6857 5566 6873
rect 5612 6864 5628 6880
rect 5635 6878 5665 6930
rect 5699 6926 5700 6933
rect 5684 6918 5700 6926
rect 5671 6886 5684 6905
rect 5699 6886 5729 6902
rect 5671 6870 5745 6886
rect 5671 6868 5684 6870
rect 5699 6868 5733 6870
rect 5336 6846 5349 6848
rect 5364 6846 5398 6848
rect 5336 6830 5398 6846
rect 5442 6841 5458 6844
rect 5520 6841 5550 6852
rect 5598 6848 5644 6864
rect 5671 6852 5745 6868
rect 5598 6846 5632 6848
rect 5597 6830 5644 6846
rect 5671 6830 5684 6852
rect 5699 6830 5729 6852
rect 5756 6830 5757 6846
rect 5772 6830 5785 6990
rect 5815 6886 5828 6990
rect 5873 6968 5874 6978
rect 5889 6968 5902 6978
rect 5873 6964 5902 6968
rect 5907 6964 5937 6990
rect 5955 6976 5971 6978
rect 6043 6976 6096 6990
rect 6044 6974 6108 6976
rect 6151 6974 6166 6990
rect 6215 6987 6245 6990
rect 6215 6984 6251 6987
rect 6181 6976 6197 6978
rect 5955 6964 5970 6968
rect 5873 6962 5970 6964
rect 5998 6962 6166 6974
rect 6182 6964 6197 6968
rect 6215 6965 6254 6984
rect 6273 6978 6280 6979
rect 6279 6971 6280 6978
rect 6263 6968 6264 6971
rect 6279 6968 6292 6971
rect 6215 6964 6245 6965
rect 6254 6964 6260 6965
rect 6263 6964 6292 6968
rect 6182 6963 6292 6964
rect 6182 6962 6298 6963
rect 5857 6954 5908 6962
rect 5857 6942 5882 6954
rect 5889 6942 5908 6954
rect 5939 6954 5989 6962
rect 5939 6946 5955 6954
rect 5962 6952 5989 6954
rect 5998 6952 6219 6962
rect 5962 6942 6219 6952
rect 6248 6954 6298 6962
rect 6248 6945 6264 6954
rect 5857 6934 5908 6942
rect 5955 6934 6219 6942
rect 6245 6942 6264 6945
rect 6271 6942 6298 6954
rect 6245 6934 6298 6942
rect 5873 6926 5874 6934
rect 5889 6926 5902 6934
rect 5873 6918 5889 6926
rect 5870 6911 5889 6914
rect 5870 6902 5892 6911
rect 5843 6892 5892 6902
rect 5843 6886 5873 6892
rect 5892 6887 5897 6892
rect 5815 6870 5889 6886
rect 5907 6878 5937 6934
rect 5972 6924 6180 6934
rect 6215 6930 6260 6934
rect 6263 6933 6264 6934
rect 6279 6933 6292 6934
rect 5998 6894 6187 6924
rect 6013 6891 6187 6894
rect 6006 6888 6187 6891
rect 5815 6868 5828 6870
rect 5843 6868 5877 6870
rect 5815 6852 5889 6868
rect 5916 6864 5929 6878
rect 5944 6864 5960 6880
rect 6006 6875 6017 6888
rect 5799 6830 5800 6846
rect 5815 6830 5828 6852
rect 5843 6830 5873 6852
rect 5916 6848 5978 6864
rect 6006 6857 6017 6873
rect 6022 6868 6032 6888
rect 6042 6868 6056 6888
rect 6059 6875 6068 6888
rect 6084 6875 6093 6888
rect 6022 6857 6056 6868
rect 6059 6857 6068 6873
rect 6084 6857 6093 6873
rect 6100 6868 6110 6888
rect 6120 6868 6134 6888
rect 6135 6875 6146 6888
rect 6100 6857 6134 6868
rect 6135 6857 6146 6873
rect 6192 6864 6208 6880
rect 6215 6878 6245 6930
rect 6279 6926 6280 6933
rect 6264 6918 6280 6926
rect 6251 6886 6264 6905
rect 6279 6886 6309 6902
rect 6251 6870 6325 6886
rect 6251 6868 6264 6870
rect 6279 6868 6313 6870
rect 5916 6846 5929 6848
rect 5944 6846 5978 6848
rect 5916 6830 5978 6846
rect 6022 6841 6038 6844
rect 6100 6841 6130 6852
rect 6178 6848 6224 6864
rect 6251 6852 6325 6868
rect 6178 6846 6212 6848
rect 6177 6830 6224 6846
rect 6251 6830 6264 6852
rect 6279 6830 6309 6852
rect 6336 6830 6337 6846
rect 6352 6830 6365 6990
rect 6395 6886 6408 6990
rect 6453 6968 6454 6978
rect 6469 6968 6482 6978
rect 6453 6964 6482 6968
rect 6487 6964 6517 6990
rect 6535 6976 6551 6978
rect 6623 6976 6676 6990
rect 6624 6974 6688 6976
rect 6731 6974 6746 6990
rect 6795 6987 6825 6990
rect 6795 6984 6831 6987
rect 6761 6976 6777 6978
rect 6535 6964 6550 6968
rect 6453 6962 6550 6964
rect 6578 6962 6746 6974
rect 6762 6964 6777 6968
rect 6795 6965 6834 6984
rect 6853 6978 6860 6979
rect 6859 6971 6860 6978
rect 6843 6968 6844 6971
rect 6859 6968 6872 6971
rect 6795 6964 6825 6965
rect 6834 6964 6840 6965
rect 6843 6964 6872 6968
rect 6762 6963 6872 6964
rect 6762 6962 6878 6963
rect 6437 6954 6488 6962
rect 6437 6942 6462 6954
rect 6469 6942 6488 6954
rect 6519 6954 6569 6962
rect 6519 6946 6535 6954
rect 6542 6952 6569 6954
rect 6578 6952 6799 6962
rect 6542 6942 6799 6952
rect 6828 6954 6878 6962
rect 6828 6945 6844 6954
rect 6437 6934 6488 6942
rect 6535 6934 6799 6942
rect 6825 6942 6844 6945
rect 6851 6942 6878 6954
rect 6825 6934 6878 6942
rect 6453 6926 6454 6934
rect 6469 6926 6482 6934
rect 6453 6918 6469 6926
rect 6450 6911 6469 6914
rect 6450 6902 6472 6911
rect 6423 6892 6472 6902
rect 6423 6886 6453 6892
rect 6472 6887 6477 6892
rect 6395 6870 6469 6886
rect 6487 6878 6517 6934
rect 6552 6924 6760 6934
rect 6795 6930 6840 6934
rect 6843 6933 6844 6934
rect 6859 6933 6872 6934
rect 6578 6894 6767 6924
rect 6593 6891 6767 6894
rect 6586 6888 6767 6891
rect 6395 6868 6408 6870
rect 6423 6868 6457 6870
rect 6395 6852 6469 6868
rect 6496 6864 6509 6878
rect 6524 6864 6540 6880
rect 6586 6875 6597 6888
rect 6379 6830 6380 6846
rect 6395 6830 6408 6852
rect 6423 6830 6453 6852
rect 6496 6848 6558 6864
rect 6586 6857 6597 6873
rect 6602 6868 6612 6888
rect 6622 6868 6636 6888
rect 6639 6875 6648 6888
rect 6664 6875 6673 6888
rect 6602 6857 6636 6868
rect 6639 6857 6648 6873
rect 6664 6857 6673 6873
rect 6680 6868 6690 6888
rect 6700 6868 6714 6888
rect 6715 6875 6726 6888
rect 6680 6857 6714 6868
rect 6715 6857 6726 6873
rect 6772 6864 6788 6880
rect 6795 6878 6825 6930
rect 6859 6926 6860 6933
rect 6844 6918 6860 6926
rect 6831 6886 6844 6905
rect 6859 6886 6889 6902
rect 6831 6870 6905 6886
rect 6831 6868 6844 6870
rect 6859 6868 6893 6870
rect 6496 6846 6509 6848
rect 6524 6846 6558 6848
rect 6496 6830 6558 6846
rect 6602 6841 6618 6844
rect 6680 6841 6710 6852
rect 6758 6848 6804 6864
rect 6831 6852 6905 6868
rect 6758 6846 6792 6848
rect 6757 6830 6804 6846
rect 6831 6830 6844 6852
rect 6859 6830 6889 6852
rect 6916 6830 6917 6846
rect 6932 6830 6945 6990
rect 6975 6886 6988 6990
rect 7033 6968 7034 6978
rect 7049 6968 7062 6978
rect 7033 6964 7062 6968
rect 7067 6964 7097 6990
rect 7115 6976 7131 6978
rect 7203 6976 7256 6990
rect 7204 6974 7268 6976
rect 7311 6974 7326 6990
rect 7375 6987 7405 6990
rect 7375 6984 7411 6987
rect 7341 6976 7357 6978
rect 7115 6964 7130 6968
rect 7033 6962 7130 6964
rect 7158 6962 7326 6974
rect 7342 6964 7357 6968
rect 7375 6965 7414 6984
rect 7433 6978 7440 6979
rect 7439 6971 7440 6978
rect 7423 6968 7424 6971
rect 7439 6968 7452 6971
rect 7375 6964 7405 6965
rect 7414 6964 7420 6965
rect 7423 6964 7452 6968
rect 7342 6963 7452 6964
rect 7342 6962 7458 6963
rect 7017 6954 7068 6962
rect 7017 6942 7042 6954
rect 7049 6942 7068 6954
rect 7099 6954 7149 6962
rect 7099 6946 7115 6954
rect 7122 6952 7149 6954
rect 7158 6952 7379 6962
rect 7122 6942 7379 6952
rect 7408 6954 7458 6962
rect 7408 6945 7424 6954
rect 7017 6934 7068 6942
rect 7115 6934 7379 6942
rect 7405 6942 7424 6945
rect 7431 6942 7458 6954
rect 7405 6934 7458 6942
rect 7033 6926 7034 6934
rect 7049 6926 7062 6934
rect 7033 6918 7049 6926
rect 7030 6911 7049 6914
rect 7030 6902 7052 6911
rect 7003 6892 7052 6902
rect 7003 6886 7033 6892
rect 7052 6887 7057 6892
rect 6975 6870 7049 6886
rect 7067 6878 7097 6934
rect 7132 6924 7340 6934
rect 7375 6930 7420 6934
rect 7423 6933 7424 6934
rect 7439 6933 7452 6934
rect 7158 6894 7347 6924
rect 7173 6891 7347 6894
rect 7166 6888 7347 6891
rect 6975 6868 6988 6870
rect 7003 6868 7037 6870
rect 6975 6852 7049 6868
rect 7076 6864 7089 6878
rect 7104 6864 7120 6880
rect 7166 6875 7177 6888
rect 6959 6830 6960 6846
rect 6975 6830 6988 6852
rect 7003 6830 7033 6852
rect 7076 6848 7138 6864
rect 7166 6857 7177 6873
rect 7182 6868 7192 6888
rect 7202 6868 7216 6888
rect 7219 6875 7228 6888
rect 7244 6875 7253 6888
rect 7182 6857 7216 6868
rect 7219 6857 7228 6873
rect 7244 6857 7253 6873
rect 7260 6868 7270 6888
rect 7280 6868 7294 6888
rect 7295 6875 7306 6888
rect 7260 6857 7294 6868
rect 7295 6857 7306 6873
rect 7352 6864 7368 6880
rect 7375 6878 7405 6930
rect 7439 6926 7440 6933
rect 7424 6918 7440 6926
rect 7411 6886 7424 6905
rect 7439 6886 7469 6902
rect 7411 6870 7485 6886
rect 7411 6868 7424 6870
rect 7439 6868 7473 6870
rect 7076 6846 7089 6848
rect 7104 6846 7138 6848
rect 7076 6830 7138 6846
rect 7182 6841 7198 6844
rect 7260 6841 7290 6852
rect 7338 6848 7384 6864
rect 7411 6852 7485 6868
rect 7338 6846 7372 6848
rect 7337 6830 7384 6846
rect 7411 6830 7424 6852
rect 7439 6830 7469 6852
rect 7496 6830 7497 6846
rect 7512 6830 7525 6990
rect 7555 6886 7568 6990
rect 7613 6968 7614 6978
rect 7629 6968 7642 6978
rect 7613 6964 7642 6968
rect 7647 6964 7677 6990
rect 7695 6976 7711 6978
rect 7783 6976 7836 6990
rect 7784 6974 7848 6976
rect 7891 6974 7906 6990
rect 7955 6987 7985 6990
rect 7955 6984 7991 6987
rect 7921 6976 7937 6978
rect 7695 6964 7710 6968
rect 7613 6962 7710 6964
rect 7738 6962 7906 6974
rect 7922 6964 7937 6968
rect 7955 6965 7994 6984
rect 8013 6978 8020 6979
rect 8019 6971 8020 6978
rect 8003 6968 8004 6971
rect 8019 6968 8032 6971
rect 7955 6964 7985 6965
rect 7994 6964 8000 6965
rect 8003 6964 8032 6968
rect 7922 6963 8032 6964
rect 7922 6962 8038 6963
rect 7597 6954 7648 6962
rect 7597 6942 7622 6954
rect 7629 6942 7648 6954
rect 7679 6954 7729 6962
rect 7679 6946 7695 6954
rect 7702 6952 7729 6954
rect 7738 6952 7959 6962
rect 7702 6942 7959 6952
rect 7988 6954 8038 6962
rect 7988 6945 8004 6954
rect 7597 6934 7648 6942
rect 7695 6934 7959 6942
rect 7985 6942 8004 6945
rect 8011 6942 8038 6954
rect 7985 6934 8038 6942
rect 7613 6926 7614 6934
rect 7629 6926 7642 6934
rect 7613 6918 7629 6926
rect 7610 6911 7629 6914
rect 7610 6902 7632 6911
rect 7583 6892 7632 6902
rect 7583 6886 7613 6892
rect 7632 6887 7637 6892
rect 7555 6870 7629 6886
rect 7647 6878 7677 6934
rect 7712 6924 7920 6934
rect 7955 6930 8000 6934
rect 8003 6933 8004 6934
rect 8019 6933 8032 6934
rect 7738 6894 7927 6924
rect 7753 6891 7927 6894
rect 7746 6888 7927 6891
rect 7555 6868 7568 6870
rect 7583 6868 7617 6870
rect 7555 6852 7629 6868
rect 7656 6864 7669 6878
rect 7684 6864 7700 6880
rect 7746 6875 7757 6888
rect 7539 6830 7540 6846
rect 7555 6830 7568 6852
rect 7583 6830 7613 6852
rect 7656 6848 7718 6864
rect 7746 6857 7757 6873
rect 7762 6868 7772 6888
rect 7782 6868 7796 6888
rect 7799 6875 7808 6888
rect 7824 6875 7833 6888
rect 7762 6857 7796 6868
rect 7799 6857 7808 6873
rect 7824 6857 7833 6873
rect 7840 6868 7850 6888
rect 7860 6868 7874 6888
rect 7875 6875 7886 6888
rect 7840 6857 7874 6868
rect 7875 6857 7886 6873
rect 7932 6864 7948 6880
rect 7955 6878 7985 6930
rect 8019 6926 8020 6933
rect 8004 6918 8020 6926
rect 7991 6886 8004 6905
rect 8019 6886 8049 6902
rect 7991 6870 8065 6886
rect 7991 6868 8004 6870
rect 8019 6868 8053 6870
rect 7656 6846 7669 6848
rect 7684 6846 7718 6848
rect 7656 6830 7718 6846
rect 7762 6841 7778 6844
rect 7840 6841 7870 6852
rect 7918 6848 7964 6864
rect 7991 6852 8065 6868
rect 7918 6846 7952 6848
rect 7917 6830 7964 6846
rect 7991 6830 8004 6852
rect 8019 6830 8049 6852
rect 8076 6830 8077 6846
rect 8092 6830 8105 6990
rect 8135 6886 8148 6990
rect 8193 6968 8194 6978
rect 8209 6968 8222 6978
rect 8193 6964 8222 6968
rect 8227 6964 8257 6990
rect 8275 6976 8291 6978
rect 8363 6976 8416 6990
rect 8364 6974 8428 6976
rect 8471 6974 8486 6990
rect 8535 6987 8565 6990
rect 8535 6984 8571 6987
rect 8501 6976 8517 6978
rect 8275 6964 8290 6968
rect 8193 6962 8290 6964
rect 8318 6962 8486 6974
rect 8502 6964 8517 6968
rect 8535 6965 8574 6984
rect 8593 6978 8600 6979
rect 8599 6971 8600 6978
rect 8583 6968 8584 6971
rect 8599 6968 8612 6971
rect 8535 6964 8565 6965
rect 8574 6964 8580 6965
rect 8583 6964 8612 6968
rect 8502 6963 8612 6964
rect 8502 6962 8618 6963
rect 8177 6954 8228 6962
rect 8177 6942 8202 6954
rect 8209 6942 8228 6954
rect 8259 6954 8309 6962
rect 8259 6946 8275 6954
rect 8282 6952 8309 6954
rect 8318 6952 8539 6962
rect 8282 6942 8539 6952
rect 8568 6954 8618 6962
rect 8568 6945 8584 6954
rect 8177 6934 8228 6942
rect 8275 6934 8539 6942
rect 8565 6942 8584 6945
rect 8591 6942 8618 6954
rect 8565 6934 8618 6942
rect 8193 6926 8194 6934
rect 8209 6926 8222 6934
rect 8193 6918 8209 6926
rect 8190 6911 8209 6914
rect 8190 6902 8212 6911
rect 8163 6892 8212 6902
rect 8163 6886 8193 6892
rect 8212 6887 8217 6892
rect 8135 6870 8209 6886
rect 8227 6878 8257 6934
rect 8292 6924 8500 6934
rect 8535 6930 8580 6934
rect 8583 6933 8584 6934
rect 8599 6933 8612 6934
rect 8318 6894 8507 6924
rect 8333 6891 8507 6894
rect 8326 6888 8507 6891
rect 8135 6868 8148 6870
rect 8163 6868 8197 6870
rect 8135 6852 8209 6868
rect 8236 6864 8249 6878
rect 8264 6864 8280 6880
rect 8326 6875 8337 6888
rect 8119 6830 8120 6846
rect 8135 6830 8148 6852
rect 8163 6830 8193 6852
rect 8236 6848 8298 6864
rect 8326 6857 8337 6873
rect 8342 6868 8352 6888
rect 8362 6868 8376 6888
rect 8379 6875 8388 6888
rect 8404 6875 8413 6888
rect 8342 6857 8376 6868
rect 8379 6857 8388 6873
rect 8404 6857 8413 6873
rect 8420 6868 8430 6888
rect 8440 6868 8454 6888
rect 8455 6875 8466 6888
rect 8420 6857 8454 6868
rect 8455 6857 8466 6873
rect 8512 6864 8528 6880
rect 8535 6878 8565 6930
rect 8599 6926 8600 6933
rect 8584 6918 8600 6926
rect 8571 6886 8584 6905
rect 8599 6886 8629 6902
rect 8571 6870 8645 6886
rect 8571 6868 8584 6870
rect 8599 6868 8633 6870
rect 8236 6846 8249 6848
rect 8264 6846 8298 6848
rect 8236 6830 8298 6846
rect 8342 6841 8358 6844
rect 8420 6841 8450 6852
rect 8498 6848 8544 6864
rect 8571 6852 8645 6868
rect 8498 6846 8532 6848
rect 8497 6830 8544 6846
rect 8571 6830 8584 6852
rect 8599 6830 8629 6852
rect 8656 6830 8657 6846
rect 8672 6830 8685 6990
rect 8715 6886 8728 6990
rect 8773 6968 8774 6978
rect 8789 6968 8802 6978
rect 8773 6964 8802 6968
rect 8807 6964 8837 6990
rect 8855 6976 8871 6978
rect 8943 6976 8996 6990
rect 8944 6974 9008 6976
rect 9051 6974 9066 6990
rect 9115 6987 9145 6990
rect 9115 6984 9151 6987
rect 9081 6976 9097 6978
rect 8855 6964 8870 6968
rect 8773 6962 8870 6964
rect 8898 6962 9066 6974
rect 9082 6964 9097 6968
rect 9115 6965 9154 6984
rect 9173 6978 9180 6979
rect 9179 6971 9180 6978
rect 9163 6968 9164 6971
rect 9179 6968 9192 6971
rect 9115 6964 9145 6965
rect 9154 6964 9160 6965
rect 9163 6964 9192 6968
rect 9082 6963 9192 6964
rect 9082 6962 9198 6963
rect 8757 6954 8808 6962
rect 8757 6942 8782 6954
rect 8789 6942 8808 6954
rect 8839 6954 8889 6962
rect 8839 6946 8855 6954
rect 8862 6952 8889 6954
rect 8898 6952 9119 6962
rect 8862 6942 9119 6952
rect 9148 6954 9198 6962
rect 9148 6945 9164 6954
rect 8757 6934 8808 6942
rect 8855 6934 9119 6942
rect 9145 6942 9164 6945
rect 9171 6942 9198 6954
rect 9145 6934 9198 6942
rect 8773 6926 8774 6934
rect 8789 6926 8802 6934
rect 8773 6918 8789 6926
rect 8770 6911 8789 6914
rect 8770 6902 8792 6911
rect 8743 6892 8792 6902
rect 8743 6886 8773 6892
rect 8792 6887 8797 6892
rect 8715 6870 8789 6886
rect 8807 6878 8837 6934
rect 8872 6924 9080 6934
rect 9115 6930 9160 6934
rect 9163 6933 9164 6934
rect 9179 6933 9192 6934
rect 8898 6894 9087 6924
rect 8913 6891 9087 6894
rect 8906 6888 9087 6891
rect 8715 6868 8728 6870
rect 8743 6868 8777 6870
rect 8715 6852 8789 6868
rect 8816 6864 8829 6878
rect 8844 6864 8860 6880
rect 8906 6875 8917 6888
rect 8699 6830 8700 6846
rect 8715 6830 8728 6852
rect 8743 6830 8773 6852
rect 8816 6848 8878 6864
rect 8906 6857 8917 6873
rect 8922 6868 8932 6888
rect 8942 6868 8956 6888
rect 8959 6875 8968 6888
rect 8984 6875 8993 6888
rect 8922 6857 8956 6868
rect 8959 6857 8968 6873
rect 8984 6857 8993 6873
rect 9000 6868 9010 6888
rect 9020 6868 9034 6888
rect 9035 6875 9046 6888
rect 9000 6857 9034 6868
rect 9035 6857 9046 6873
rect 9092 6864 9108 6880
rect 9115 6878 9145 6930
rect 9179 6926 9180 6933
rect 9164 6918 9180 6926
rect 9151 6886 9164 6905
rect 9179 6886 9209 6902
rect 9151 6870 9225 6886
rect 9151 6868 9164 6870
rect 9179 6868 9213 6870
rect 8816 6846 8829 6848
rect 8844 6846 8878 6848
rect 8816 6830 8878 6846
rect 8922 6841 8938 6844
rect 9000 6841 9030 6852
rect 9078 6848 9124 6864
rect 9151 6852 9225 6868
rect 9078 6846 9112 6848
rect 9077 6830 9124 6846
rect 9151 6830 9164 6852
rect 9179 6830 9209 6852
rect 9236 6830 9237 6846
rect 9252 6830 9265 6990
rect -7 6822 34 6830
rect -7 6796 8 6822
rect 15 6796 34 6822
rect 98 6818 160 6830
rect 172 6818 247 6830
rect 305 6818 380 6830
rect 392 6818 423 6830
rect 429 6818 464 6830
rect 98 6816 260 6818
rect -7 6788 34 6796
rect 116 6792 129 6816
rect 144 6814 159 6816
rect -1 6778 0 6788
rect 15 6778 28 6788
rect 43 6778 73 6792
rect 116 6778 159 6792
rect 183 6789 190 6796
rect 193 6792 260 6816
rect 292 6816 464 6818
rect 262 6794 290 6798
rect 292 6794 372 6816
rect 393 6814 408 6816
rect 262 6792 372 6794
rect 193 6788 372 6792
rect 166 6778 196 6788
rect 198 6778 351 6788
rect 359 6778 389 6788
rect 393 6778 423 6792
rect 451 6778 464 6816
rect 536 6822 571 6830
rect 536 6796 537 6822
rect 544 6796 571 6822
rect 479 6778 509 6792
rect 536 6788 571 6796
rect 573 6822 614 6830
rect 573 6796 588 6822
rect 595 6796 614 6822
rect 678 6818 740 6830
rect 752 6818 827 6830
rect 885 6818 960 6830
rect 972 6818 1003 6830
rect 1009 6818 1044 6830
rect 678 6816 840 6818
rect 573 6788 614 6796
rect 696 6792 709 6816
rect 724 6814 739 6816
rect 536 6778 537 6788
rect 552 6778 565 6788
rect 579 6778 580 6788
rect 595 6778 608 6788
rect 623 6778 653 6792
rect 696 6778 739 6792
rect 763 6789 770 6796
rect 773 6792 840 6816
rect 872 6816 1044 6818
rect 842 6794 870 6798
rect 872 6794 952 6816
rect 973 6814 988 6816
rect 842 6792 952 6794
rect 773 6788 952 6792
rect 746 6778 776 6788
rect 778 6778 931 6788
rect 939 6778 969 6788
rect 973 6778 1003 6792
rect 1031 6778 1044 6816
rect 1116 6822 1151 6830
rect 1116 6796 1117 6822
rect 1124 6796 1151 6822
rect 1059 6778 1089 6792
rect 1116 6788 1151 6796
rect 1153 6822 1194 6830
rect 1153 6796 1168 6822
rect 1175 6796 1194 6822
rect 1258 6818 1320 6830
rect 1332 6818 1407 6830
rect 1465 6818 1540 6830
rect 1552 6818 1583 6830
rect 1589 6818 1624 6830
rect 1258 6816 1420 6818
rect 1153 6788 1194 6796
rect 1276 6792 1289 6816
rect 1304 6814 1319 6816
rect 1116 6778 1117 6788
rect 1132 6778 1145 6788
rect 1159 6778 1160 6788
rect 1175 6778 1188 6788
rect 1203 6778 1233 6792
rect 1276 6778 1319 6792
rect 1343 6789 1350 6796
rect 1353 6792 1420 6816
rect 1452 6816 1624 6818
rect 1422 6794 1450 6798
rect 1452 6794 1532 6816
rect 1553 6814 1568 6816
rect 1422 6792 1532 6794
rect 1353 6788 1532 6792
rect 1326 6778 1356 6788
rect 1358 6778 1511 6788
rect 1519 6778 1549 6788
rect 1553 6778 1583 6792
rect 1611 6778 1624 6816
rect 1696 6822 1731 6830
rect 1696 6796 1697 6822
rect 1704 6796 1731 6822
rect 1639 6778 1669 6792
rect 1696 6788 1731 6796
rect 1733 6822 1774 6830
rect 1733 6796 1748 6822
rect 1755 6796 1774 6822
rect 1838 6818 1900 6830
rect 1912 6818 1987 6830
rect 2045 6818 2120 6830
rect 2132 6818 2163 6830
rect 2169 6818 2204 6830
rect 1838 6816 2000 6818
rect 1733 6788 1774 6796
rect 1856 6792 1869 6816
rect 1884 6814 1899 6816
rect 1696 6778 1697 6788
rect 1712 6778 1725 6788
rect 1739 6778 1740 6788
rect 1755 6778 1768 6788
rect 1783 6778 1813 6792
rect 1856 6778 1899 6792
rect 1923 6789 1930 6796
rect 1933 6792 2000 6816
rect 2032 6816 2204 6818
rect 2002 6794 2030 6798
rect 2032 6794 2112 6816
rect 2133 6814 2148 6816
rect 2002 6792 2112 6794
rect 1933 6788 2112 6792
rect 1906 6778 1936 6788
rect 1938 6778 2091 6788
rect 2099 6778 2129 6788
rect 2133 6778 2163 6792
rect 2191 6778 2204 6816
rect 2276 6822 2311 6830
rect 2276 6796 2277 6822
rect 2284 6796 2311 6822
rect 2219 6778 2249 6792
rect 2276 6788 2311 6796
rect 2313 6822 2354 6830
rect 2313 6796 2328 6822
rect 2335 6796 2354 6822
rect 2418 6818 2480 6830
rect 2492 6818 2567 6830
rect 2625 6818 2700 6830
rect 2712 6818 2743 6830
rect 2749 6818 2784 6830
rect 2418 6816 2580 6818
rect 2313 6788 2354 6796
rect 2436 6792 2449 6816
rect 2464 6814 2479 6816
rect 2276 6778 2277 6788
rect 2292 6778 2305 6788
rect 2319 6778 2320 6788
rect 2335 6778 2348 6788
rect 2363 6778 2393 6792
rect 2436 6778 2479 6792
rect 2503 6789 2510 6796
rect 2513 6792 2580 6816
rect 2612 6816 2784 6818
rect 2582 6794 2610 6798
rect 2612 6794 2692 6816
rect 2713 6814 2728 6816
rect 2582 6792 2692 6794
rect 2513 6788 2692 6792
rect 2486 6778 2516 6788
rect 2518 6778 2671 6788
rect 2679 6778 2709 6788
rect 2713 6778 2743 6792
rect 2771 6778 2784 6816
rect 2856 6822 2891 6830
rect 2856 6796 2857 6822
rect 2864 6796 2891 6822
rect 2799 6778 2829 6792
rect 2856 6788 2891 6796
rect 2893 6822 2934 6830
rect 2893 6796 2908 6822
rect 2915 6796 2934 6822
rect 2998 6818 3060 6830
rect 3072 6818 3147 6830
rect 3205 6818 3280 6830
rect 3292 6818 3323 6830
rect 3329 6818 3364 6830
rect 2998 6816 3160 6818
rect 2893 6788 2934 6796
rect 3016 6792 3029 6816
rect 3044 6814 3059 6816
rect 2856 6778 2857 6788
rect 2872 6778 2885 6788
rect 2899 6778 2900 6788
rect 2915 6778 2928 6788
rect 2943 6778 2973 6792
rect 3016 6778 3059 6792
rect 3083 6789 3090 6796
rect 3093 6792 3160 6816
rect 3192 6816 3364 6818
rect 3162 6794 3190 6798
rect 3192 6794 3272 6816
rect 3293 6814 3308 6816
rect 3162 6792 3272 6794
rect 3093 6788 3272 6792
rect 3066 6778 3096 6788
rect 3098 6778 3251 6788
rect 3259 6778 3289 6788
rect 3293 6778 3323 6792
rect 3351 6778 3364 6816
rect 3436 6822 3471 6830
rect 3436 6796 3437 6822
rect 3444 6796 3471 6822
rect 3379 6778 3409 6792
rect 3436 6788 3471 6796
rect 3473 6822 3514 6830
rect 3473 6796 3488 6822
rect 3495 6796 3514 6822
rect 3578 6818 3640 6830
rect 3652 6818 3727 6830
rect 3785 6818 3860 6830
rect 3872 6818 3903 6830
rect 3909 6818 3944 6830
rect 3578 6816 3740 6818
rect 3473 6788 3514 6796
rect 3596 6792 3609 6816
rect 3624 6814 3639 6816
rect 3436 6778 3437 6788
rect 3452 6778 3465 6788
rect 3479 6778 3480 6788
rect 3495 6778 3508 6788
rect 3523 6778 3553 6792
rect 3596 6778 3639 6792
rect 3663 6789 3670 6796
rect 3673 6792 3740 6816
rect 3772 6816 3944 6818
rect 3742 6794 3770 6798
rect 3772 6794 3852 6816
rect 3873 6814 3888 6816
rect 3742 6792 3852 6794
rect 3673 6788 3852 6792
rect 3646 6778 3676 6788
rect 3678 6778 3831 6788
rect 3839 6778 3869 6788
rect 3873 6778 3903 6792
rect 3931 6778 3944 6816
rect 4016 6822 4051 6830
rect 4016 6796 4017 6822
rect 4024 6796 4051 6822
rect 3959 6778 3989 6792
rect 4016 6788 4051 6796
rect 4053 6822 4094 6830
rect 4053 6796 4068 6822
rect 4075 6796 4094 6822
rect 4158 6818 4220 6830
rect 4232 6818 4307 6830
rect 4365 6818 4440 6830
rect 4452 6818 4483 6830
rect 4489 6818 4524 6830
rect 4158 6816 4320 6818
rect 4053 6788 4094 6796
rect 4176 6792 4189 6816
rect 4204 6814 4219 6816
rect 4016 6778 4017 6788
rect 4032 6778 4045 6788
rect 4059 6778 4060 6788
rect 4075 6778 4088 6788
rect 4103 6778 4133 6792
rect 4176 6778 4219 6792
rect 4243 6789 4250 6796
rect 4253 6792 4320 6816
rect 4352 6816 4524 6818
rect 4322 6794 4350 6798
rect 4352 6794 4432 6816
rect 4453 6814 4468 6816
rect 4322 6792 4432 6794
rect 4253 6788 4432 6792
rect 4226 6778 4256 6788
rect 4258 6778 4411 6788
rect 4419 6778 4449 6788
rect 4453 6778 4483 6792
rect 4511 6778 4524 6816
rect 4596 6822 4631 6830
rect 4596 6796 4597 6822
rect 4604 6796 4631 6822
rect 4539 6778 4569 6792
rect 4596 6788 4631 6796
rect 4633 6822 4674 6830
rect 4633 6796 4648 6822
rect 4655 6796 4674 6822
rect 4738 6818 4800 6830
rect 4812 6818 4887 6830
rect 4945 6818 5020 6830
rect 5032 6818 5063 6830
rect 5069 6818 5104 6830
rect 4738 6816 4900 6818
rect 4633 6788 4674 6796
rect 4756 6792 4769 6816
rect 4784 6814 4799 6816
rect 4596 6778 4597 6788
rect 4612 6778 4625 6788
rect 4639 6778 4640 6788
rect 4655 6778 4668 6788
rect 4683 6778 4713 6792
rect 4756 6778 4799 6792
rect 4823 6789 4830 6796
rect 4833 6792 4900 6816
rect 4932 6816 5104 6818
rect 4902 6794 4930 6798
rect 4932 6794 5012 6816
rect 5033 6814 5048 6816
rect 4902 6792 5012 6794
rect 4833 6788 5012 6792
rect 4806 6778 4836 6788
rect 4838 6778 4991 6788
rect 4999 6778 5029 6788
rect 5033 6778 5063 6792
rect 5091 6778 5104 6816
rect 5176 6822 5211 6830
rect 5176 6796 5177 6822
rect 5184 6796 5211 6822
rect 5119 6778 5149 6792
rect 5176 6788 5211 6796
rect 5213 6822 5254 6830
rect 5213 6796 5228 6822
rect 5235 6796 5254 6822
rect 5318 6818 5380 6830
rect 5392 6818 5467 6830
rect 5525 6818 5600 6830
rect 5612 6818 5643 6830
rect 5649 6818 5684 6830
rect 5318 6816 5480 6818
rect 5213 6788 5254 6796
rect 5336 6792 5349 6816
rect 5364 6814 5379 6816
rect 5176 6778 5177 6788
rect 5192 6778 5205 6788
rect 5219 6778 5220 6788
rect 5235 6778 5248 6788
rect 5263 6778 5293 6792
rect 5336 6778 5379 6792
rect 5403 6789 5410 6796
rect 5413 6792 5480 6816
rect 5512 6816 5684 6818
rect 5482 6794 5510 6798
rect 5512 6794 5592 6816
rect 5613 6814 5628 6816
rect 5482 6792 5592 6794
rect 5413 6788 5592 6792
rect 5386 6778 5416 6788
rect 5418 6778 5571 6788
rect 5579 6778 5609 6788
rect 5613 6778 5643 6792
rect 5671 6778 5684 6816
rect 5756 6822 5791 6830
rect 5756 6796 5757 6822
rect 5764 6796 5791 6822
rect 5699 6778 5729 6792
rect 5756 6788 5791 6796
rect 5793 6822 5834 6830
rect 5793 6796 5808 6822
rect 5815 6796 5834 6822
rect 5898 6818 5960 6830
rect 5972 6818 6047 6830
rect 6105 6818 6180 6830
rect 6192 6818 6223 6830
rect 6229 6818 6264 6830
rect 5898 6816 6060 6818
rect 5793 6788 5834 6796
rect 5916 6792 5929 6816
rect 5944 6814 5959 6816
rect 5756 6778 5757 6788
rect 5772 6778 5785 6788
rect 5799 6778 5800 6788
rect 5815 6778 5828 6788
rect 5843 6778 5873 6792
rect 5916 6778 5959 6792
rect 5983 6789 5990 6796
rect 5993 6792 6060 6816
rect 6092 6816 6264 6818
rect 6062 6794 6090 6798
rect 6092 6794 6172 6816
rect 6193 6814 6208 6816
rect 6062 6792 6172 6794
rect 5993 6788 6172 6792
rect 5966 6778 5996 6788
rect 5998 6778 6151 6788
rect 6159 6778 6189 6788
rect 6193 6778 6223 6792
rect 6251 6778 6264 6816
rect 6336 6822 6371 6830
rect 6336 6796 6337 6822
rect 6344 6796 6371 6822
rect 6279 6778 6309 6792
rect 6336 6788 6371 6796
rect 6373 6822 6414 6830
rect 6373 6796 6388 6822
rect 6395 6796 6414 6822
rect 6478 6818 6540 6830
rect 6552 6818 6627 6830
rect 6685 6818 6760 6830
rect 6772 6818 6803 6830
rect 6809 6818 6844 6830
rect 6478 6816 6640 6818
rect 6373 6788 6414 6796
rect 6496 6792 6509 6816
rect 6524 6814 6539 6816
rect 6336 6778 6337 6788
rect 6352 6778 6365 6788
rect 6379 6778 6380 6788
rect 6395 6778 6408 6788
rect 6423 6778 6453 6792
rect 6496 6778 6539 6792
rect 6563 6789 6570 6796
rect 6573 6792 6640 6816
rect 6672 6816 6844 6818
rect 6642 6794 6670 6798
rect 6672 6794 6752 6816
rect 6773 6814 6788 6816
rect 6642 6792 6752 6794
rect 6573 6788 6752 6792
rect 6546 6778 6576 6788
rect 6578 6778 6731 6788
rect 6739 6778 6769 6788
rect 6773 6778 6803 6792
rect 6831 6778 6844 6816
rect 6916 6822 6951 6830
rect 6916 6796 6917 6822
rect 6924 6796 6951 6822
rect 6859 6778 6889 6792
rect 6916 6788 6951 6796
rect 6953 6822 6994 6830
rect 6953 6796 6968 6822
rect 6975 6796 6994 6822
rect 7058 6818 7120 6830
rect 7132 6818 7207 6830
rect 7265 6818 7340 6830
rect 7352 6818 7383 6830
rect 7389 6818 7424 6830
rect 7058 6816 7220 6818
rect 6953 6788 6994 6796
rect 7076 6792 7089 6816
rect 7104 6814 7119 6816
rect 6916 6778 6917 6788
rect 6932 6778 6945 6788
rect 6959 6778 6960 6788
rect 6975 6778 6988 6788
rect 7003 6778 7033 6792
rect 7076 6778 7119 6792
rect 7143 6789 7150 6796
rect 7153 6792 7220 6816
rect 7252 6816 7424 6818
rect 7222 6794 7250 6798
rect 7252 6794 7332 6816
rect 7353 6814 7368 6816
rect 7222 6792 7332 6794
rect 7153 6788 7332 6792
rect 7126 6778 7156 6788
rect 7158 6778 7311 6788
rect 7319 6778 7349 6788
rect 7353 6778 7383 6792
rect 7411 6778 7424 6816
rect 7496 6822 7531 6830
rect 7496 6796 7497 6822
rect 7504 6796 7531 6822
rect 7439 6778 7469 6792
rect 7496 6788 7531 6796
rect 7533 6822 7574 6830
rect 7533 6796 7548 6822
rect 7555 6796 7574 6822
rect 7638 6818 7700 6830
rect 7712 6818 7787 6830
rect 7845 6818 7920 6830
rect 7932 6818 7963 6830
rect 7969 6818 8004 6830
rect 7638 6816 7800 6818
rect 7533 6788 7574 6796
rect 7656 6792 7669 6816
rect 7684 6814 7699 6816
rect 7496 6778 7497 6788
rect 7512 6778 7525 6788
rect 7539 6778 7540 6788
rect 7555 6778 7568 6788
rect 7583 6778 7613 6792
rect 7656 6778 7699 6792
rect 7723 6789 7730 6796
rect 7733 6792 7800 6816
rect 7832 6816 8004 6818
rect 7802 6794 7830 6798
rect 7832 6794 7912 6816
rect 7933 6814 7948 6816
rect 7802 6792 7912 6794
rect 7733 6788 7912 6792
rect 7706 6778 7736 6788
rect 7738 6778 7891 6788
rect 7899 6778 7929 6788
rect 7933 6778 7963 6792
rect 7991 6778 8004 6816
rect 8076 6822 8111 6830
rect 8076 6796 8077 6822
rect 8084 6796 8111 6822
rect 8019 6778 8049 6792
rect 8076 6788 8111 6796
rect 8113 6822 8154 6830
rect 8113 6796 8128 6822
rect 8135 6796 8154 6822
rect 8218 6818 8280 6830
rect 8292 6818 8367 6830
rect 8425 6818 8500 6830
rect 8512 6818 8543 6830
rect 8549 6818 8584 6830
rect 8218 6816 8380 6818
rect 8113 6788 8154 6796
rect 8236 6792 8249 6816
rect 8264 6814 8279 6816
rect 8076 6778 8077 6788
rect 8092 6778 8105 6788
rect 8119 6778 8120 6788
rect 8135 6778 8148 6788
rect 8163 6778 8193 6792
rect 8236 6778 8279 6792
rect 8303 6789 8310 6796
rect 8313 6792 8380 6816
rect 8412 6816 8584 6818
rect 8382 6794 8410 6798
rect 8412 6794 8492 6816
rect 8513 6814 8528 6816
rect 8382 6792 8492 6794
rect 8313 6788 8492 6792
rect 8286 6778 8316 6788
rect 8318 6778 8471 6788
rect 8479 6778 8509 6788
rect 8513 6778 8543 6792
rect 8571 6778 8584 6816
rect 8656 6822 8691 6830
rect 8656 6796 8657 6822
rect 8664 6796 8691 6822
rect 8599 6778 8629 6792
rect 8656 6788 8691 6796
rect 8693 6822 8734 6830
rect 8693 6796 8708 6822
rect 8715 6796 8734 6822
rect 8798 6818 8860 6830
rect 8872 6818 8947 6830
rect 9005 6818 9080 6830
rect 9092 6818 9123 6830
rect 9129 6818 9164 6830
rect 8798 6816 8960 6818
rect 8693 6788 8734 6796
rect 8816 6792 8829 6816
rect 8844 6814 8859 6816
rect 8656 6778 8657 6788
rect 8672 6778 8685 6788
rect 8699 6778 8700 6788
rect 8715 6778 8728 6788
rect 8743 6778 8773 6792
rect 8816 6778 8859 6792
rect 8883 6789 8890 6796
rect 8893 6792 8960 6816
rect 8992 6816 9164 6818
rect 8962 6794 8990 6798
rect 8992 6794 9072 6816
rect 9093 6814 9108 6816
rect 8962 6792 9072 6794
rect 8893 6788 9072 6792
rect 8866 6778 8896 6788
rect 8898 6778 9051 6788
rect 9059 6778 9089 6788
rect 9093 6778 9123 6792
rect 9151 6778 9164 6816
rect 9236 6822 9271 6830
rect 9236 6796 9237 6822
rect 9244 6796 9271 6822
rect 9179 6778 9209 6792
rect 9236 6788 9271 6796
rect 9236 6778 9237 6788
rect 9252 6778 9265 6788
rect -1 6772 9265 6778
rect 0 6764 9265 6772
rect 15 6734 28 6764
rect 43 6746 73 6764
rect 116 6750 130 6764
rect 166 6750 386 6764
rect 117 6748 130 6750
rect 83 6736 98 6748
rect 80 6734 102 6736
rect 107 6734 137 6748
rect 198 6746 351 6750
rect 180 6734 372 6746
rect 415 6734 445 6748
rect 451 6734 464 6764
rect 479 6746 509 6764
rect 552 6734 565 6764
rect 595 6734 608 6764
rect 623 6746 653 6764
rect 696 6750 710 6764
rect 746 6750 966 6764
rect 697 6748 710 6750
rect 663 6736 678 6748
rect 660 6734 682 6736
rect 687 6734 717 6748
rect 778 6746 931 6750
rect 760 6734 952 6746
rect 995 6734 1025 6748
rect 1031 6734 1044 6764
rect 1059 6746 1089 6764
rect 1132 6734 1145 6764
rect 1175 6734 1188 6764
rect 1203 6746 1233 6764
rect 1276 6750 1290 6764
rect 1326 6750 1546 6764
rect 1277 6748 1290 6750
rect 1243 6736 1258 6748
rect 1240 6734 1262 6736
rect 1267 6734 1297 6748
rect 1358 6746 1511 6750
rect 1340 6734 1532 6746
rect 1575 6734 1605 6748
rect 1611 6734 1624 6764
rect 1639 6746 1669 6764
rect 1712 6734 1725 6764
rect 1755 6734 1768 6764
rect 1783 6746 1813 6764
rect 1856 6750 1870 6764
rect 1906 6750 2126 6764
rect 1857 6748 1870 6750
rect 1823 6736 1838 6748
rect 1820 6734 1842 6736
rect 1847 6734 1877 6748
rect 1938 6746 2091 6750
rect 1920 6734 2112 6746
rect 2155 6734 2185 6748
rect 2191 6734 2204 6764
rect 2219 6746 2249 6764
rect 2292 6734 2305 6764
rect 2335 6734 2348 6764
rect 2363 6746 2393 6764
rect 2436 6750 2450 6764
rect 2486 6750 2706 6764
rect 2437 6748 2450 6750
rect 2403 6736 2418 6748
rect 2400 6734 2422 6736
rect 2427 6734 2457 6748
rect 2518 6746 2671 6750
rect 2500 6734 2692 6746
rect 2735 6734 2765 6748
rect 2771 6734 2784 6764
rect 2799 6746 2829 6764
rect 2872 6734 2885 6764
rect 2915 6734 2928 6764
rect 2943 6746 2973 6764
rect 3016 6750 3030 6764
rect 3066 6750 3286 6764
rect 3017 6748 3030 6750
rect 2983 6736 2998 6748
rect 2980 6734 3002 6736
rect 3007 6734 3037 6748
rect 3098 6746 3251 6750
rect 3080 6734 3272 6746
rect 3315 6734 3345 6748
rect 3351 6734 3364 6764
rect 3379 6746 3409 6764
rect 3452 6734 3465 6764
rect 3495 6734 3508 6764
rect 3523 6746 3553 6764
rect 3596 6750 3610 6764
rect 3646 6750 3866 6764
rect 3597 6748 3610 6750
rect 3563 6736 3578 6748
rect 3560 6734 3582 6736
rect 3587 6734 3617 6748
rect 3678 6746 3831 6750
rect 3660 6734 3852 6746
rect 3895 6734 3925 6748
rect 3931 6734 3944 6764
rect 3959 6746 3989 6764
rect 4032 6734 4045 6764
rect 4075 6734 4088 6764
rect 4103 6746 4133 6764
rect 4176 6750 4190 6764
rect 4226 6750 4446 6764
rect 4177 6748 4190 6750
rect 4143 6736 4158 6748
rect 4140 6734 4162 6736
rect 4167 6734 4197 6748
rect 4258 6746 4411 6750
rect 4240 6734 4432 6746
rect 4475 6734 4505 6748
rect 4511 6734 4524 6764
rect 4539 6746 4569 6764
rect 4612 6734 4625 6764
rect 4655 6734 4668 6764
rect 4683 6746 4713 6764
rect 4756 6750 4770 6764
rect 4806 6750 5026 6764
rect 4757 6748 4770 6750
rect 4723 6736 4738 6748
rect 4720 6734 4742 6736
rect 4747 6734 4777 6748
rect 4838 6746 4991 6750
rect 4820 6734 5012 6746
rect 5055 6734 5085 6748
rect 5091 6734 5104 6764
rect 5119 6746 5149 6764
rect 5192 6734 5205 6764
rect 5235 6734 5248 6764
rect 5263 6746 5293 6764
rect 5336 6750 5350 6764
rect 5386 6750 5606 6764
rect 5337 6748 5350 6750
rect 5303 6736 5318 6748
rect 5300 6734 5322 6736
rect 5327 6734 5357 6748
rect 5418 6746 5571 6750
rect 5400 6734 5592 6746
rect 5635 6734 5665 6748
rect 5671 6734 5684 6764
rect 5699 6746 5729 6764
rect 5772 6734 5785 6764
rect 5815 6734 5828 6764
rect 5843 6746 5873 6764
rect 5916 6750 5930 6764
rect 5966 6750 6186 6764
rect 5917 6748 5930 6750
rect 5883 6736 5898 6748
rect 5880 6734 5902 6736
rect 5907 6734 5937 6748
rect 5998 6746 6151 6750
rect 5980 6734 6172 6746
rect 6215 6734 6245 6748
rect 6251 6734 6264 6764
rect 6279 6746 6309 6764
rect 6352 6734 6365 6764
rect 6395 6734 6408 6764
rect 6423 6746 6453 6764
rect 6496 6750 6510 6764
rect 6546 6750 6766 6764
rect 6497 6748 6510 6750
rect 6463 6736 6478 6748
rect 6460 6734 6482 6736
rect 6487 6734 6517 6748
rect 6578 6746 6731 6750
rect 6560 6734 6752 6746
rect 6795 6734 6825 6748
rect 6831 6734 6844 6764
rect 6859 6746 6889 6764
rect 6932 6734 6945 6764
rect 6975 6734 6988 6764
rect 7003 6746 7033 6764
rect 7076 6750 7090 6764
rect 7126 6750 7346 6764
rect 7077 6748 7090 6750
rect 7043 6736 7058 6748
rect 7040 6734 7062 6736
rect 7067 6734 7097 6748
rect 7158 6746 7311 6750
rect 7140 6734 7332 6746
rect 7375 6734 7405 6748
rect 7411 6734 7424 6764
rect 7439 6746 7469 6764
rect 7512 6734 7525 6764
rect 7555 6734 7568 6764
rect 7583 6746 7613 6764
rect 7656 6750 7670 6764
rect 7706 6750 7926 6764
rect 7657 6748 7670 6750
rect 7623 6736 7638 6748
rect 7620 6734 7642 6736
rect 7647 6734 7677 6748
rect 7738 6746 7891 6750
rect 7720 6734 7912 6746
rect 7955 6734 7985 6748
rect 7991 6734 8004 6764
rect 8019 6746 8049 6764
rect 8092 6734 8105 6764
rect 8135 6734 8148 6764
rect 8163 6746 8193 6764
rect 8236 6750 8250 6764
rect 8286 6750 8506 6764
rect 8237 6748 8250 6750
rect 8203 6736 8218 6748
rect 8200 6734 8222 6736
rect 8227 6734 8257 6748
rect 8318 6746 8471 6750
rect 8300 6734 8492 6746
rect 8535 6734 8565 6748
rect 8571 6734 8584 6764
rect 8599 6746 8629 6764
rect 8672 6734 8685 6764
rect 8715 6734 8728 6764
rect 8743 6746 8773 6764
rect 8816 6750 8830 6764
rect 8866 6750 9086 6764
rect 8817 6748 8830 6750
rect 8783 6736 8798 6748
rect 8780 6734 8802 6736
rect 8807 6734 8837 6748
rect 8898 6746 9051 6750
rect 8880 6734 9072 6746
rect 9115 6734 9145 6748
rect 9151 6734 9164 6764
rect 9179 6746 9209 6764
rect 9252 6734 9265 6764
rect 0 6720 9265 6734
rect 15 6616 28 6720
rect 73 6698 74 6708
rect 89 6698 102 6708
rect 73 6694 102 6698
rect 107 6694 137 6720
rect 155 6706 171 6708
rect 243 6706 296 6720
rect 244 6704 308 6706
rect 351 6704 366 6720
rect 415 6717 445 6720
rect 415 6714 451 6717
rect 381 6706 397 6708
rect 155 6694 170 6698
rect 73 6692 170 6694
rect 198 6692 366 6704
rect 382 6694 397 6698
rect 415 6695 454 6714
rect 473 6708 480 6709
rect 479 6701 480 6708
rect 463 6698 464 6701
rect 479 6698 492 6701
rect 415 6694 445 6695
rect 454 6694 460 6695
rect 463 6694 492 6698
rect 382 6693 492 6694
rect 382 6692 498 6693
rect 57 6684 108 6692
rect 57 6672 82 6684
rect 89 6672 108 6684
rect 139 6684 189 6692
rect 139 6676 155 6684
rect 162 6682 189 6684
rect 198 6682 419 6692
rect 162 6672 419 6682
rect 448 6684 498 6692
rect 448 6675 464 6684
rect 57 6664 108 6672
rect 155 6664 419 6672
rect 445 6672 464 6675
rect 471 6672 498 6684
rect 445 6664 498 6672
rect 73 6656 74 6664
rect 89 6656 102 6664
rect 73 6648 89 6656
rect 70 6641 89 6644
rect 70 6632 92 6641
rect 43 6622 92 6632
rect 43 6616 73 6622
rect 92 6617 97 6622
rect 15 6600 89 6616
rect 107 6608 137 6664
rect 172 6654 380 6664
rect 415 6660 460 6664
rect 463 6663 464 6664
rect 479 6663 492 6664
rect 198 6624 387 6654
rect 213 6621 387 6624
rect 206 6618 387 6621
rect 15 6598 28 6600
rect 43 6598 77 6600
rect 15 6582 89 6598
rect 116 6594 129 6608
rect 144 6594 160 6610
rect 206 6605 217 6618
rect -1 6560 0 6576
rect 15 6560 28 6582
rect 43 6560 73 6582
rect 116 6578 178 6594
rect 206 6587 217 6603
rect 222 6598 232 6618
rect 242 6598 256 6618
rect 259 6605 268 6618
rect 284 6605 293 6618
rect 222 6587 256 6598
rect 259 6587 268 6603
rect 284 6587 293 6603
rect 300 6598 310 6618
rect 320 6598 334 6618
rect 335 6605 346 6618
rect 300 6587 334 6598
rect 335 6587 346 6603
rect 392 6594 408 6610
rect 415 6608 445 6660
rect 479 6656 480 6663
rect 464 6648 480 6656
rect 451 6616 464 6635
rect 479 6616 509 6632
rect 451 6600 525 6616
rect 451 6598 464 6600
rect 479 6598 513 6600
rect 116 6576 129 6578
rect 144 6576 178 6578
rect 116 6560 178 6576
rect 222 6571 238 6574
rect 300 6571 330 6582
rect 378 6578 424 6594
rect 451 6582 525 6598
rect 378 6576 412 6578
rect 377 6560 424 6576
rect 451 6560 464 6582
rect 479 6560 509 6582
rect 536 6560 537 6576
rect 552 6560 565 6720
rect 595 6616 608 6720
rect 653 6698 654 6708
rect 669 6698 682 6708
rect 653 6694 682 6698
rect 687 6694 717 6720
rect 735 6706 751 6708
rect 823 6706 876 6720
rect 824 6704 888 6706
rect 931 6704 946 6720
rect 995 6717 1025 6720
rect 995 6714 1031 6717
rect 961 6706 977 6708
rect 735 6694 750 6698
rect 653 6692 750 6694
rect 778 6692 946 6704
rect 962 6694 977 6698
rect 995 6695 1034 6714
rect 1053 6708 1060 6709
rect 1059 6701 1060 6708
rect 1043 6698 1044 6701
rect 1059 6698 1072 6701
rect 995 6694 1025 6695
rect 1034 6694 1040 6695
rect 1043 6694 1072 6698
rect 962 6693 1072 6694
rect 962 6692 1078 6693
rect 637 6684 688 6692
rect 637 6672 662 6684
rect 669 6672 688 6684
rect 719 6684 769 6692
rect 719 6676 735 6684
rect 742 6682 769 6684
rect 778 6682 999 6692
rect 742 6672 999 6682
rect 1028 6684 1078 6692
rect 1028 6675 1044 6684
rect 637 6664 688 6672
rect 735 6664 999 6672
rect 1025 6672 1044 6675
rect 1051 6672 1078 6684
rect 1025 6664 1078 6672
rect 653 6656 654 6664
rect 669 6656 682 6664
rect 653 6648 669 6656
rect 650 6641 669 6644
rect 650 6632 672 6641
rect 623 6622 672 6632
rect 623 6616 653 6622
rect 672 6617 677 6622
rect 595 6600 669 6616
rect 687 6608 717 6664
rect 752 6654 960 6664
rect 995 6660 1040 6664
rect 1043 6663 1044 6664
rect 1059 6663 1072 6664
rect 778 6624 967 6654
rect 793 6621 967 6624
rect 786 6618 967 6621
rect 595 6598 608 6600
rect 623 6598 657 6600
rect 595 6582 669 6598
rect 696 6594 709 6608
rect 724 6594 740 6610
rect 786 6605 797 6618
rect 579 6560 580 6576
rect 595 6560 608 6582
rect 623 6560 653 6582
rect 696 6578 758 6594
rect 786 6587 797 6603
rect 802 6598 812 6618
rect 822 6598 836 6618
rect 839 6605 848 6618
rect 864 6605 873 6618
rect 802 6587 836 6598
rect 839 6587 848 6603
rect 864 6587 873 6603
rect 880 6598 890 6618
rect 900 6598 914 6618
rect 915 6605 926 6618
rect 880 6587 914 6598
rect 915 6587 926 6603
rect 972 6594 988 6610
rect 995 6608 1025 6660
rect 1059 6656 1060 6663
rect 1044 6648 1060 6656
rect 1031 6616 1044 6635
rect 1059 6616 1089 6632
rect 1031 6600 1105 6616
rect 1031 6598 1044 6600
rect 1059 6598 1093 6600
rect 696 6576 709 6578
rect 724 6576 758 6578
rect 696 6560 758 6576
rect 802 6571 818 6574
rect 880 6571 910 6582
rect 958 6578 1004 6594
rect 1031 6582 1105 6598
rect 958 6576 992 6578
rect 957 6560 1004 6576
rect 1031 6560 1044 6582
rect 1059 6560 1089 6582
rect 1116 6560 1117 6576
rect 1132 6560 1145 6720
rect 1175 6616 1188 6720
rect 1233 6698 1234 6708
rect 1249 6698 1262 6708
rect 1233 6694 1262 6698
rect 1267 6694 1297 6720
rect 1315 6706 1331 6708
rect 1403 6706 1456 6720
rect 1404 6704 1468 6706
rect 1511 6704 1526 6720
rect 1575 6717 1605 6720
rect 1575 6714 1611 6717
rect 1541 6706 1557 6708
rect 1315 6694 1330 6698
rect 1233 6692 1330 6694
rect 1358 6692 1526 6704
rect 1542 6694 1557 6698
rect 1575 6695 1614 6714
rect 1633 6708 1640 6709
rect 1639 6701 1640 6708
rect 1623 6698 1624 6701
rect 1639 6698 1652 6701
rect 1575 6694 1605 6695
rect 1614 6694 1620 6695
rect 1623 6694 1652 6698
rect 1542 6693 1652 6694
rect 1542 6692 1658 6693
rect 1217 6684 1268 6692
rect 1217 6672 1242 6684
rect 1249 6672 1268 6684
rect 1299 6684 1349 6692
rect 1299 6676 1315 6684
rect 1322 6682 1349 6684
rect 1358 6682 1579 6692
rect 1322 6672 1579 6682
rect 1608 6684 1658 6692
rect 1608 6675 1624 6684
rect 1217 6664 1268 6672
rect 1315 6664 1579 6672
rect 1605 6672 1624 6675
rect 1631 6672 1658 6684
rect 1605 6664 1658 6672
rect 1233 6656 1234 6664
rect 1249 6656 1262 6664
rect 1233 6648 1249 6656
rect 1230 6641 1249 6644
rect 1230 6632 1252 6641
rect 1203 6622 1252 6632
rect 1203 6616 1233 6622
rect 1252 6617 1257 6622
rect 1175 6600 1249 6616
rect 1267 6608 1297 6664
rect 1332 6654 1540 6664
rect 1575 6660 1620 6664
rect 1623 6663 1624 6664
rect 1639 6663 1652 6664
rect 1358 6624 1547 6654
rect 1373 6621 1547 6624
rect 1366 6618 1547 6621
rect 1175 6598 1188 6600
rect 1203 6598 1237 6600
rect 1175 6582 1249 6598
rect 1276 6594 1289 6608
rect 1304 6594 1320 6610
rect 1366 6605 1377 6618
rect 1159 6560 1160 6576
rect 1175 6560 1188 6582
rect 1203 6560 1233 6582
rect 1276 6578 1338 6594
rect 1366 6587 1377 6603
rect 1382 6598 1392 6618
rect 1402 6598 1416 6618
rect 1419 6605 1428 6618
rect 1444 6605 1453 6618
rect 1382 6587 1416 6598
rect 1419 6587 1428 6603
rect 1444 6587 1453 6603
rect 1460 6598 1470 6618
rect 1480 6598 1494 6618
rect 1495 6605 1506 6618
rect 1460 6587 1494 6598
rect 1495 6587 1506 6603
rect 1552 6594 1568 6610
rect 1575 6608 1605 6660
rect 1639 6656 1640 6663
rect 1624 6648 1640 6656
rect 1611 6616 1624 6635
rect 1639 6616 1669 6632
rect 1611 6600 1685 6616
rect 1611 6598 1624 6600
rect 1639 6598 1673 6600
rect 1276 6576 1289 6578
rect 1304 6576 1338 6578
rect 1276 6560 1338 6576
rect 1382 6571 1398 6574
rect 1460 6571 1490 6582
rect 1538 6578 1584 6594
rect 1611 6582 1685 6598
rect 1538 6576 1572 6578
rect 1537 6560 1584 6576
rect 1611 6560 1624 6582
rect 1639 6560 1669 6582
rect 1696 6560 1697 6576
rect 1712 6560 1725 6720
rect 1755 6616 1768 6720
rect 1813 6698 1814 6708
rect 1829 6698 1842 6708
rect 1813 6694 1842 6698
rect 1847 6694 1877 6720
rect 1895 6706 1911 6708
rect 1983 6706 2036 6720
rect 1984 6704 2048 6706
rect 2091 6704 2106 6720
rect 2155 6717 2185 6720
rect 2155 6714 2191 6717
rect 2121 6706 2137 6708
rect 1895 6694 1910 6698
rect 1813 6692 1910 6694
rect 1938 6692 2106 6704
rect 2122 6694 2137 6698
rect 2155 6695 2194 6714
rect 2213 6708 2220 6709
rect 2219 6701 2220 6708
rect 2203 6698 2204 6701
rect 2219 6698 2232 6701
rect 2155 6694 2185 6695
rect 2194 6694 2200 6695
rect 2203 6694 2232 6698
rect 2122 6693 2232 6694
rect 2122 6692 2238 6693
rect 1797 6684 1848 6692
rect 1797 6672 1822 6684
rect 1829 6672 1848 6684
rect 1879 6684 1929 6692
rect 1879 6676 1895 6684
rect 1902 6682 1929 6684
rect 1938 6682 2159 6692
rect 1902 6672 2159 6682
rect 2188 6684 2238 6692
rect 2188 6675 2204 6684
rect 1797 6664 1848 6672
rect 1895 6664 2159 6672
rect 2185 6672 2204 6675
rect 2211 6672 2238 6684
rect 2185 6664 2238 6672
rect 1813 6656 1814 6664
rect 1829 6656 1842 6664
rect 1813 6648 1829 6656
rect 1810 6641 1829 6644
rect 1810 6632 1832 6641
rect 1783 6622 1832 6632
rect 1783 6616 1813 6622
rect 1832 6617 1837 6622
rect 1755 6600 1829 6616
rect 1847 6608 1877 6664
rect 1912 6654 2120 6664
rect 2155 6660 2200 6664
rect 2203 6663 2204 6664
rect 2219 6663 2232 6664
rect 1938 6624 2127 6654
rect 1953 6621 2127 6624
rect 1946 6618 2127 6621
rect 1755 6598 1768 6600
rect 1783 6598 1817 6600
rect 1755 6582 1829 6598
rect 1856 6594 1869 6608
rect 1884 6594 1900 6610
rect 1946 6605 1957 6618
rect 1739 6560 1740 6576
rect 1755 6560 1768 6582
rect 1783 6560 1813 6582
rect 1856 6578 1918 6594
rect 1946 6587 1957 6603
rect 1962 6598 1972 6618
rect 1982 6598 1996 6618
rect 1999 6605 2008 6618
rect 2024 6605 2033 6618
rect 1962 6587 1996 6598
rect 1999 6587 2008 6603
rect 2024 6587 2033 6603
rect 2040 6598 2050 6618
rect 2060 6598 2074 6618
rect 2075 6605 2086 6618
rect 2040 6587 2074 6598
rect 2075 6587 2086 6603
rect 2132 6594 2148 6610
rect 2155 6608 2185 6660
rect 2219 6656 2220 6663
rect 2204 6648 2220 6656
rect 2191 6616 2204 6635
rect 2219 6616 2249 6632
rect 2191 6600 2265 6616
rect 2191 6598 2204 6600
rect 2219 6598 2253 6600
rect 1856 6576 1869 6578
rect 1884 6576 1918 6578
rect 1856 6560 1918 6576
rect 1962 6571 1976 6574
rect 2040 6571 2070 6582
rect 2118 6578 2164 6594
rect 2191 6582 2265 6598
rect 2118 6576 2152 6578
rect 2117 6560 2164 6576
rect 2191 6560 2204 6582
rect 2219 6560 2249 6582
rect 2276 6560 2277 6576
rect 2292 6560 2305 6720
rect 2335 6616 2348 6720
rect 2393 6698 2394 6708
rect 2409 6698 2422 6708
rect 2393 6694 2422 6698
rect 2427 6694 2457 6720
rect 2475 6706 2491 6708
rect 2563 6706 2616 6720
rect 2564 6704 2628 6706
rect 2671 6704 2686 6720
rect 2735 6717 2765 6720
rect 2735 6714 2771 6717
rect 2701 6706 2717 6708
rect 2475 6694 2490 6698
rect 2393 6692 2490 6694
rect 2518 6692 2686 6704
rect 2702 6694 2717 6698
rect 2735 6695 2774 6714
rect 2793 6708 2800 6709
rect 2799 6701 2800 6708
rect 2783 6698 2784 6701
rect 2799 6698 2812 6701
rect 2735 6694 2765 6695
rect 2774 6694 2780 6695
rect 2783 6694 2812 6698
rect 2702 6693 2812 6694
rect 2702 6692 2818 6693
rect 2377 6684 2428 6692
rect 2377 6672 2402 6684
rect 2409 6672 2428 6684
rect 2459 6684 2509 6692
rect 2459 6676 2475 6684
rect 2482 6682 2509 6684
rect 2518 6682 2739 6692
rect 2482 6672 2739 6682
rect 2768 6684 2818 6692
rect 2768 6675 2784 6684
rect 2377 6664 2428 6672
rect 2475 6664 2739 6672
rect 2765 6672 2784 6675
rect 2791 6672 2818 6684
rect 2765 6664 2818 6672
rect 2393 6656 2394 6664
rect 2409 6656 2422 6664
rect 2393 6648 2409 6656
rect 2390 6641 2409 6644
rect 2390 6632 2412 6641
rect 2363 6622 2412 6632
rect 2363 6616 2393 6622
rect 2412 6617 2417 6622
rect 2335 6600 2409 6616
rect 2427 6608 2457 6664
rect 2492 6654 2700 6664
rect 2735 6660 2780 6664
rect 2783 6663 2784 6664
rect 2799 6663 2812 6664
rect 2518 6624 2707 6654
rect 2533 6621 2707 6624
rect 2526 6618 2707 6621
rect 2335 6598 2348 6600
rect 2363 6598 2397 6600
rect 2335 6582 2409 6598
rect 2436 6594 2449 6608
rect 2464 6594 2480 6610
rect 2526 6605 2537 6618
rect 2319 6560 2320 6576
rect 2335 6560 2348 6582
rect 2363 6560 2393 6582
rect 2436 6578 2498 6594
rect 2526 6587 2537 6603
rect 2542 6598 2552 6618
rect 2562 6598 2576 6618
rect 2579 6605 2588 6618
rect 2604 6605 2613 6618
rect 2542 6587 2576 6598
rect 2579 6587 2588 6603
rect 2604 6587 2613 6603
rect 2620 6598 2630 6618
rect 2640 6598 2654 6618
rect 2655 6605 2666 6618
rect 2620 6587 2654 6598
rect 2655 6587 2666 6603
rect 2712 6594 2728 6610
rect 2735 6608 2765 6660
rect 2799 6656 2800 6663
rect 2784 6648 2800 6656
rect 2771 6616 2784 6635
rect 2799 6616 2829 6632
rect 2771 6600 2845 6616
rect 2771 6598 2784 6600
rect 2799 6598 2833 6600
rect 2436 6576 2449 6578
rect 2464 6576 2498 6578
rect 2436 6560 2498 6576
rect 2542 6571 2558 6574
rect 2620 6571 2650 6582
rect 2698 6578 2744 6594
rect 2771 6582 2845 6598
rect 2698 6576 2732 6578
rect 2697 6560 2744 6576
rect 2771 6560 2784 6582
rect 2799 6560 2829 6582
rect 2856 6560 2857 6576
rect 2872 6560 2885 6720
rect 2915 6616 2928 6720
rect 2973 6698 2974 6708
rect 2989 6698 3002 6708
rect 2973 6694 3002 6698
rect 3007 6694 3037 6720
rect 3055 6706 3071 6708
rect 3143 6706 3196 6720
rect 3144 6704 3208 6706
rect 3251 6704 3266 6720
rect 3315 6717 3345 6720
rect 3315 6714 3351 6717
rect 3281 6706 3297 6708
rect 3055 6694 3070 6698
rect 2973 6692 3070 6694
rect 3098 6692 3266 6704
rect 3282 6694 3297 6698
rect 3315 6695 3354 6714
rect 3373 6708 3380 6709
rect 3379 6701 3380 6708
rect 3363 6698 3364 6701
rect 3379 6698 3392 6701
rect 3315 6694 3345 6695
rect 3354 6694 3360 6695
rect 3363 6694 3392 6698
rect 3282 6693 3392 6694
rect 3282 6692 3398 6693
rect 2957 6684 3008 6692
rect 2957 6672 2982 6684
rect 2989 6672 3008 6684
rect 3039 6684 3089 6692
rect 3039 6676 3055 6684
rect 3062 6682 3089 6684
rect 3098 6682 3319 6692
rect 3062 6672 3319 6682
rect 3348 6684 3398 6692
rect 3348 6675 3364 6684
rect 2957 6664 3008 6672
rect 3055 6664 3319 6672
rect 3345 6672 3364 6675
rect 3371 6672 3398 6684
rect 3345 6664 3398 6672
rect 2973 6656 2974 6664
rect 2989 6656 3002 6664
rect 2973 6648 2989 6656
rect 2970 6641 2989 6644
rect 2970 6632 2992 6641
rect 2943 6622 2992 6632
rect 2943 6616 2973 6622
rect 2992 6617 2997 6622
rect 2915 6600 2989 6616
rect 3007 6608 3037 6664
rect 3072 6654 3280 6664
rect 3315 6660 3360 6664
rect 3363 6663 3364 6664
rect 3379 6663 3392 6664
rect 3098 6624 3287 6654
rect 3113 6621 3287 6624
rect 3106 6618 3287 6621
rect 2915 6598 2928 6600
rect 2943 6598 2977 6600
rect 2915 6582 2989 6598
rect 3016 6594 3029 6608
rect 3044 6594 3060 6610
rect 3106 6605 3117 6618
rect 2899 6560 2900 6576
rect 2915 6560 2928 6582
rect 2943 6560 2973 6582
rect 3016 6578 3078 6594
rect 3106 6587 3117 6603
rect 3122 6598 3132 6618
rect 3142 6598 3156 6618
rect 3159 6605 3168 6618
rect 3184 6605 3193 6618
rect 3122 6587 3156 6598
rect 3159 6587 3168 6603
rect 3184 6587 3193 6603
rect 3200 6598 3210 6618
rect 3220 6598 3234 6618
rect 3235 6605 3246 6618
rect 3200 6587 3234 6598
rect 3235 6587 3246 6603
rect 3292 6594 3308 6610
rect 3315 6608 3345 6660
rect 3379 6656 3380 6663
rect 3364 6648 3380 6656
rect 3351 6616 3364 6635
rect 3379 6616 3409 6632
rect 3351 6600 3425 6616
rect 3351 6598 3364 6600
rect 3379 6598 3413 6600
rect 3016 6576 3029 6578
rect 3044 6576 3078 6578
rect 3016 6560 3078 6576
rect 3122 6571 3138 6574
rect 3200 6571 3230 6582
rect 3278 6578 3324 6594
rect 3351 6582 3425 6598
rect 3278 6576 3312 6578
rect 3277 6560 3324 6576
rect 3351 6560 3364 6582
rect 3379 6560 3409 6582
rect 3436 6560 3437 6576
rect 3452 6560 3465 6720
rect 3495 6616 3508 6720
rect 3553 6698 3554 6708
rect 3569 6698 3582 6708
rect 3553 6694 3582 6698
rect 3587 6694 3617 6720
rect 3635 6706 3651 6708
rect 3723 6706 3776 6720
rect 3724 6704 3788 6706
rect 3831 6704 3846 6720
rect 3895 6717 3925 6720
rect 3895 6714 3931 6717
rect 3861 6706 3877 6708
rect 3635 6694 3650 6698
rect 3553 6692 3650 6694
rect 3678 6692 3846 6704
rect 3862 6694 3877 6698
rect 3895 6695 3934 6714
rect 3953 6708 3960 6709
rect 3959 6701 3960 6708
rect 3943 6698 3944 6701
rect 3959 6698 3972 6701
rect 3895 6694 3925 6695
rect 3934 6694 3940 6695
rect 3943 6694 3972 6698
rect 3862 6693 3972 6694
rect 3862 6692 3978 6693
rect 3537 6684 3588 6692
rect 3537 6672 3562 6684
rect 3569 6672 3588 6684
rect 3619 6684 3669 6692
rect 3619 6676 3635 6684
rect 3642 6682 3669 6684
rect 3678 6682 3899 6692
rect 3642 6672 3899 6682
rect 3928 6684 3978 6692
rect 3928 6675 3944 6684
rect 3537 6664 3588 6672
rect 3635 6664 3899 6672
rect 3925 6672 3944 6675
rect 3951 6672 3978 6684
rect 3925 6664 3978 6672
rect 3553 6656 3554 6664
rect 3569 6656 3582 6664
rect 3553 6648 3569 6656
rect 3550 6641 3569 6644
rect 3550 6632 3572 6641
rect 3523 6622 3572 6632
rect 3523 6616 3553 6622
rect 3572 6617 3577 6622
rect 3495 6600 3569 6616
rect 3587 6608 3617 6664
rect 3652 6654 3860 6664
rect 3895 6660 3940 6664
rect 3943 6663 3944 6664
rect 3959 6663 3972 6664
rect 3678 6624 3867 6654
rect 3693 6621 3867 6624
rect 3686 6618 3867 6621
rect 3495 6598 3508 6600
rect 3523 6598 3557 6600
rect 3495 6582 3569 6598
rect 3596 6594 3609 6608
rect 3624 6594 3640 6610
rect 3686 6605 3697 6618
rect 3479 6560 3480 6576
rect 3495 6560 3508 6582
rect 3523 6560 3553 6582
rect 3596 6578 3658 6594
rect 3686 6587 3697 6603
rect 3702 6598 3712 6618
rect 3722 6598 3736 6618
rect 3739 6605 3748 6618
rect 3764 6605 3773 6618
rect 3702 6587 3736 6598
rect 3739 6587 3748 6603
rect 3764 6587 3773 6603
rect 3780 6598 3790 6618
rect 3800 6598 3814 6618
rect 3815 6605 3826 6618
rect 3780 6587 3814 6598
rect 3815 6587 3826 6603
rect 3872 6594 3888 6610
rect 3895 6608 3925 6660
rect 3959 6656 3960 6663
rect 3944 6648 3960 6656
rect 3931 6616 3944 6635
rect 3959 6616 3989 6632
rect 3931 6600 4005 6616
rect 3931 6598 3944 6600
rect 3959 6598 3993 6600
rect 3596 6576 3609 6578
rect 3624 6576 3658 6578
rect 3596 6560 3658 6576
rect 3702 6571 3718 6574
rect 3780 6571 3810 6582
rect 3858 6578 3904 6594
rect 3931 6582 4005 6598
rect 3858 6576 3892 6578
rect 3857 6560 3904 6576
rect 3931 6560 3944 6582
rect 3959 6560 3989 6582
rect 4016 6560 4017 6576
rect 4032 6560 4045 6720
rect 4075 6616 4088 6720
rect 4133 6698 4134 6708
rect 4149 6698 4162 6708
rect 4133 6694 4162 6698
rect 4167 6694 4197 6720
rect 4215 6706 4231 6708
rect 4303 6706 4356 6720
rect 4304 6704 4368 6706
rect 4411 6704 4426 6720
rect 4475 6717 4505 6720
rect 4475 6714 4511 6717
rect 4441 6706 4457 6708
rect 4215 6694 4230 6698
rect 4133 6692 4230 6694
rect 4258 6692 4426 6704
rect 4442 6694 4457 6698
rect 4475 6695 4514 6714
rect 4533 6708 4540 6709
rect 4539 6701 4540 6708
rect 4523 6698 4524 6701
rect 4539 6698 4552 6701
rect 4475 6694 4505 6695
rect 4514 6694 4520 6695
rect 4523 6694 4552 6698
rect 4442 6693 4552 6694
rect 4442 6692 4558 6693
rect 4117 6684 4168 6692
rect 4117 6672 4142 6684
rect 4149 6672 4168 6684
rect 4199 6684 4249 6692
rect 4199 6676 4215 6684
rect 4222 6682 4249 6684
rect 4258 6682 4479 6692
rect 4222 6672 4479 6682
rect 4508 6684 4558 6692
rect 4508 6675 4524 6684
rect 4117 6664 4168 6672
rect 4215 6664 4479 6672
rect 4505 6672 4524 6675
rect 4531 6672 4558 6684
rect 4505 6664 4558 6672
rect 4133 6656 4134 6664
rect 4149 6656 4162 6664
rect 4133 6648 4149 6656
rect 4130 6641 4149 6644
rect 4130 6632 4152 6641
rect 4103 6622 4152 6632
rect 4103 6616 4133 6622
rect 4152 6617 4157 6622
rect 4075 6600 4149 6616
rect 4167 6608 4197 6664
rect 4232 6654 4440 6664
rect 4475 6660 4520 6664
rect 4523 6663 4524 6664
rect 4539 6663 4552 6664
rect 4258 6624 4447 6654
rect 4273 6621 4447 6624
rect 4266 6618 4447 6621
rect 4075 6598 4088 6600
rect 4103 6598 4137 6600
rect 4075 6582 4149 6598
rect 4176 6594 4189 6608
rect 4204 6594 4220 6610
rect 4266 6605 4277 6618
rect 4059 6560 4060 6576
rect 4075 6560 4088 6582
rect 4103 6560 4133 6582
rect 4176 6578 4238 6594
rect 4266 6587 4277 6603
rect 4282 6598 4292 6618
rect 4302 6598 4316 6618
rect 4319 6605 4328 6618
rect 4344 6605 4353 6618
rect 4282 6587 4316 6598
rect 4319 6587 4328 6603
rect 4344 6587 4353 6603
rect 4360 6598 4370 6618
rect 4380 6598 4394 6618
rect 4395 6605 4406 6618
rect 4360 6587 4394 6598
rect 4395 6587 4406 6603
rect 4452 6594 4468 6610
rect 4475 6608 4505 6660
rect 4539 6656 4540 6663
rect 4524 6648 4540 6656
rect 4511 6616 4524 6635
rect 4539 6616 4569 6632
rect 4511 6600 4585 6616
rect 4511 6598 4524 6600
rect 4539 6598 4573 6600
rect 4176 6576 4189 6578
rect 4204 6576 4238 6578
rect 4176 6560 4238 6576
rect 4282 6571 4298 6574
rect 4360 6571 4390 6582
rect 4438 6578 4484 6594
rect 4511 6582 4585 6598
rect 4438 6576 4472 6578
rect 4437 6560 4484 6576
rect 4511 6560 4524 6582
rect 4539 6560 4569 6582
rect 4596 6560 4597 6576
rect 4612 6560 4625 6720
rect 4655 6616 4668 6720
rect 4713 6698 4714 6708
rect 4729 6698 4742 6708
rect 4713 6694 4742 6698
rect 4747 6694 4777 6720
rect 4795 6706 4811 6708
rect 4883 6706 4936 6720
rect 4884 6704 4948 6706
rect 4991 6704 5006 6720
rect 5055 6717 5085 6720
rect 5055 6714 5091 6717
rect 5021 6706 5037 6708
rect 4795 6694 4810 6698
rect 4713 6692 4810 6694
rect 4838 6692 5006 6704
rect 5022 6694 5037 6698
rect 5055 6695 5094 6714
rect 5113 6708 5120 6709
rect 5119 6701 5120 6708
rect 5103 6698 5104 6701
rect 5119 6698 5132 6701
rect 5055 6694 5085 6695
rect 5094 6694 5100 6695
rect 5103 6694 5132 6698
rect 5022 6693 5132 6694
rect 5022 6692 5138 6693
rect 4697 6684 4748 6692
rect 4697 6672 4722 6684
rect 4729 6672 4748 6684
rect 4779 6684 4829 6692
rect 4779 6676 4795 6684
rect 4802 6682 4829 6684
rect 4838 6682 5059 6692
rect 4802 6672 5059 6682
rect 5088 6684 5138 6692
rect 5088 6675 5104 6684
rect 4697 6664 4748 6672
rect 4795 6664 5059 6672
rect 5085 6672 5104 6675
rect 5111 6672 5138 6684
rect 5085 6664 5138 6672
rect 4713 6656 4714 6664
rect 4729 6656 4742 6664
rect 4713 6648 4729 6656
rect 4710 6641 4729 6644
rect 4710 6632 4732 6641
rect 4683 6622 4732 6632
rect 4683 6616 4713 6622
rect 4732 6617 4737 6622
rect 4655 6600 4729 6616
rect 4747 6608 4777 6664
rect 4812 6654 5020 6664
rect 5055 6660 5100 6664
rect 5103 6663 5104 6664
rect 5119 6663 5132 6664
rect 4838 6624 5027 6654
rect 4853 6621 5027 6624
rect 4846 6618 5027 6621
rect 4655 6598 4668 6600
rect 4683 6598 4717 6600
rect 4655 6582 4729 6598
rect 4756 6594 4769 6608
rect 4784 6594 4800 6610
rect 4846 6605 4857 6618
rect 4639 6560 4640 6576
rect 4655 6560 4668 6582
rect 4683 6560 4713 6582
rect 4756 6578 4818 6594
rect 4846 6587 4857 6603
rect 4862 6598 4872 6618
rect 4882 6598 4896 6618
rect 4899 6605 4908 6618
rect 4924 6605 4933 6618
rect 4862 6587 4896 6598
rect 4899 6587 4908 6603
rect 4924 6587 4933 6603
rect 4940 6598 4950 6618
rect 4960 6598 4974 6618
rect 4975 6605 4986 6618
rect 4940 6587 4974 6598
rect 4975 6587 4986 6603
rect 5032 6594 5048 6610
rect 5055 6608 5085 6660
rect 5119 6656 5120 6663
rect 5104 6648 5120 6656
rect 5091 6616 5104 6635
rect 5119 6616 5149 6632
rect 5091 6600 5165 6616
rect 5091 6598 5104 6600
rect 5119 6598 5153 6600
rect 4756 6576 4769 6578
rect 4784 6576 4818 6578
rect 4756 6560 4818 6576
rect 4862 6571 4878 6574
rect 4940 6571 4970 6582
rect 5018 6578 5064 6594
rect 5091 6582 5165 6598
rect 5018 6576 5052 6578
rect 5017 6560 5064 6576
rect 5091 6560 5104 6582
rect 5119 6560 5149 6582
rect 5176 6560 5177 6576
rect 5192 6560 5205 6720
rect 5235 6616 5248 6720
rect 5293 6698 5294 6708
rect 5309 6698 5322 6708
rect 5293 6694 5322 6698
rect 5327 6694 5357 6720
rect 5375 6706 5391 6708
rect 5463 6706 5516 6720
rect 5464 6704 5528 6706
rect 5571 6704 5586 6720
rect 5635 6717 5665 6720
rect 5635 6714 5671 6717
rect 5601 6706 5617 6708
rect 5375 6694 5390 6698
rect 5293 6692 5390 6694
rect 5418 6692 5586 6704
rect 5602 6694 5617 6698
rect 5635 6695 5674 6714
rect 5693 6708 5700 6709
rect 5699 6701 5700 6708
rect 5683 6698 5684 6701
rect 5699 6698 5712 6701
rect 5635 6694 5665 6695
rect 5674 6694 5680 6695
rect 5683 6694 5712 6698
rect 5602 6693 5712 6694
rect 5602 6692 5718 6693
rect 5277 6684 5328 6692
rect 5277 6672 5302 6684
rect 5309 6672 5328 6684
rect 5359 6684 5409 6692
rect 5359 6676 5375 6684
rect 5382 6682 5409 6684
rect 5418 6682 5639 6692
rect 5382 6672 5639 6682
rect 5668 6684 5718 6692
rect 5668 6675 5684 6684
rect 5277 6664 5328 6672
rect 5375 6664 5639 6672
rect 5665 6672 5684 6675
rect 5691 6672 5718 6684
rect 5665 6664 5718 6672
rect 5293 6656 5294 6664
rect 5309 6656 5322 6664
rect 5293 6648 5309 6656
rect 5290 6641 5309 6644
rect 5290 6632 5312 6641
rect 5263 6622 5312 6632
rect 5263 6616 5293 6622
rect 5312 6617 5317 6622
rect 5235 6600 5309 6616
rect 5327 6608 5357 6664
rect 5392 6654 5600 6664
rect 5635 6660 5680 6664
rect 5683 6663 5684 6664
rect 5699 6663 5712 6664
rect 5418 6624 5607 6654
rect 5433 6621 5607 6624
rect 5426 6618 5607 6621
rect 5235 6598 5248 6600
rect 5263 6598 5297 6600
rect 5235 6582 5309 6598
rect 5336 6594 5349 6608
rect 5364 6594 5380 6610
rect 5426 6605 5437 6618
rect 5219 6560 5220 6576
rect 5235 6560 5248 6582
rect 5263 6560 5293 6582
rect 5336 6578 5398 6594
rect 5426 6587 5437 6603
rect 5442 6598 5452 6618
rect 5462 6598 5476 6618
rect 5479 6605 5488 6618
rect 5504 6605 5513 6618
rect 5442 6587 5476 6598
rect 5479 6587 5488 6603
rect 5504 6587 5513 6603
rect 5520 6598 5530 6618
rect 5540 6598 5554 6618
rect 5555 6605 5566 6618
rect 5520 6587 5554 6598
rect 5555 6587 5566 6603
rect 5612 6594 5628 6610
rect 5635 6608 5665 6660
rect 5699 6656 5700 6663
rect 5684 6648 5700 6656
rect 5671 6616 5684 6635
rect 5699 6616 5729 6632
rect 5671 6600 5745 6616
rect 5671 6598 5684 6600
rect 5699 6598 5733 6600
rect 5336 6576 5349 6578
rect 5364 6576 5398 6578
rect 5336 6560 5398 6576
rect 5442 6571 5458 6574
rect 5520 6571 5550 6582
rect 5598 6578 5644 6594
rect 5671 6582 5745 6598
rect 5598 6576 5632 6578
rect 5597 6560 5644 6576
rect 5671 6560 5684 6582
rect 5699 6560 5729 6582
rect 5756 6560 5757 6576
rect 5772 6560 5785 6720
rect 5815 6616 5828 6720
rect 5873 6698 5874 6708
rect 5889 6698 5902 6708
rect 5873 6694 5902 6698
rect 5907 6694 5937 6720
rect 5955 6706 5971 6708
rect 6043 6706 6096 6720
rect 6044 6704 6108 6706
rect 6151 6704 6166 6720
rect 6215 6717 6245 6720
rect 6215 6714 6251 6717
rect 6181 6706 6197 6708
rect 5955 6694 5970 6698
rect 5873 6692 5970 6694
rect 5998 6692 6166 6704
rect 6182 6694 6197 6698
rect 6215 6695 6254 6714
rect 6273 6708 6280 6709
rect 6279 6701 6280 6708
rect 6263 6698 6264 6701
rect 6279 6698 6292 6701
rect 6215 6694 6245 6695
rect 6254 6694 6260 6695
rect 6263 6694 6292 6698
rect 6182 6693 6292 6694
rect 6182 6692 6298 6693
rect 5857 6684 5908 6692
rect 5857 6672 5882 6684
rect 5889 6672 5908 6684
rect 5939 6684 5989 6692
rect 5939 6676 5955 6684
rect 5962 6682 5989 6684
rect 5998 6682 6219 6692
rect 5962 6672 6219 6682
rect 6248 6684 6298 6692
rect 6248 6675 6264 6684
rect 5857 6664 5908 6672
rect 5955 6664 6219 6672
rect 6245 6672 6264 6675
rect 6271 6672 6298 6684
rect 6245 6664 6298 6672
rect 5873 6656 5874 6664
rect 5889 6656 5902 6664
rect 5873 6648 5889 6656
rect 5870 6641 5889 6644
rect 5870 6632 5892 6641
rect 5843 6622 5892 6632
rect 5843 6616 5873 6622
rect 5892 6617 5897 6622
rect 5815 6600 5889 6616
rect 5907 6608 5937 6664
rect 5972 6654 6180 6664
rect 6215 6660 6260 6664
rect 6263 6663 6264 6664
rect 6279 6663 6292 6664
rect 5998 6624 6187 6654
rect 6013 6621 6187 6624
rect 6006 6618 6187 6621
rect 5815 6598 5828 6600
rect 5843 6598 5877 6600
rect 5815 6582 5889 6598
rect 5916 6594 5929 6608
rect 5944 6594 5960 6610
rect 6006 6605 6017 6618
rect 5799 6560 5800 6576
rect 5815 6560 5828 6582
rect 5843 6560 5873 6582
rect 5916 6578 5978 6594
rect 6006 6587 6017 6603
rect 6022 6598 6032 6618
rect 6042 6598 6056 6618
rect 6059 6605 6068 6618
rect 6084 6605 6093 6618
rect 6022 6587 6056 6598
rect 6059 6587 6068 6603
rect 6084 6587 6093 6603
rect 6100 6598 6110 6618
rect 6120 6598 6134 6618
rect 6135 6605 6146 6618
rect 6100 6587 6134 6598
rect 6135 6587 6146 6603
rect 6192 6594 6208 6610
rect 6215 6608 6245 6660
rect 6279 6656 6280 6663
rect 6264 6648 6280 6656
rect 6251 6616 6264 6635
rect 6279 6616 6309 6632
rect 6251 6600 6325 6616
rect 6251 6598 6264 6600
rect 6279 6598 6313 6600
rect 5916 6576 5929 6578
rect 5944 6576 5978 6578
rect 5916 6560 5978 6576
rect 6022 6571 6038 6574
rect 6100 6571 6130 6582
rect 6178 6578 6224 6594
rect 6251 6582 6325 6598
rect 6178 6576 6212 6578
rect 6177 6560 6224 6576
rect 6251 6560 6264 6582
rect 6279 6560 6309 6582
rect 6336 6560 6337 6576
rect 6352 6560 6365 6720
rect 6395 6616 6408 6720
rect 6453 6698 6454 6708
rect 6469 6698 6482 6708
rect 6453 6694 6482 6698
rect 6487 6694 6517 6720
rect 6535 6706 6551 6708
rect 6623 6706 6676 6720
rect 6624 6704 6688 6706
rect 6731 6704 6746 6720
rect 6795 6717 6825 6720
rect 6795 6714 6831 6717
rect 6761 6706 6777 6708
rect 6535 6694 6550 6698
rect 6453 6692 6550 6694
rect 6578 6692 6746 6704
rect 6762 6694 6777 6698
rect 6795 6695 6834 6714
rect 6853 6708 6860 6709
rect 6859 6701 6860 6708
rect 6843 6698 6844 6701
rect 6859 6698 6872 6701
rect 6795 6694 6825 6695
rect 6834 6694 6840 6695
rect 6843 6694 6872 6698
rect 6762 6693 6872 6694
rect 6762 6692 6878 6693
rect 6437 6684 6488 6692
rect 6437 6672 6462 6684
rect 6469 6672 6488 6684
rect 6519 6684 6569 6692
rect 6519 6676 6535 6684
rect 6542 6682 6569 6684
rect 6578 6682 6799 6692
rect 6542 6672 6799 6682
rect 6828 6684 6878 6692
rect 6828 6675 6844 6684
rect 6437 6664 6488 6672
rect 6535 6664 6799 6672
rect 6825 6672 6844 6675
rect 6851 6672 6878 6684
rect 6825 6664 6878 6672
rect 6453 6656 6454 6664
rect 6469 6656 6482 6664
rect 6453 6648 6469 6656
rect 6450 6641 6469 6644
rect 6450 6632 6472 6641
rect 6423 6622 6472 6632
rect 6423 6616 6453 6622
rect 6472 6617 6477 6622
rect 6395 6600 6469 6616
rect 6487 6608 6517 6664
rect 6552 6654 6760 6664
rect 6795 6660 6840 6664
rect 6843 6663 6844 6664
rect 6859 6663 6872 6664
rect 6578 6624 6767 6654
rect 6593 6621 6767 6624
rect 6586 6618 6767 6621
rect 6395 6598 6408 6600
rect 6423 6598 6457 6600
rect 6395 6582 6469 6598
rect 6496 6594 6509 6608
rect 6524 6594 6540 6610
rect 6586 6605 6597 6618
rect 6379 6560 6380 6576
rect 6395 6560 6408 6582
rect 6423 6560 6453 6582
rect 6496 6578 6558 6594
rect 6586 6587 6597 6603
rect 6602 6598 6612 6618
rect 6622 6598 6636 6618
rect 6639 6605 6648 6618
rect 6664 6605 6673 6618
rect 6602 6587 6636 6598
rect 6639 6587 6648 6603
rect 6664 6587 6673 6603
rect 6680 6598 6690 6618
rect 6700 6598 6714 6618
rect 6715 6605 6726 6618
rect 6680 6587 6714 6598
rect 6715 6587 6726 6603
rect 6772 6594 6788 6610
rect 6795 6608 6825 6660
rect 6859 6656 6860 6663
rect 6844 6648 6860 6656
rect 6831 6616 6844 6635
rect 6859 6616 6889 6632
rect 6831 6600 6905 6616
rect 6831 6598 6844 6600
rect 6859 6598 6893 6600
rect 6496 6576 6509 6578
rect 6524 6576 6558 6578
rect 6496 6560 6558 6576
rect 6602 6571 6618 6574
rect 6680 6571 6710 6582
rect 6758 6578 6804 6594
rect 6831 6582 6905 6598
rect 6758 6576 6792 6578
rect 6757 6560 6804 6576
rect 6831 6560 6844 6582
rect 6859 6560 6889 6582
rect 6916 6560 6917 6576
rect 6932 6560 6945 6720
rect 6975 6616 6988 6720
rect 7033 6698 7034 6708
rect 7049 6698 7062 6708
rect 7033 6694 7062 6698
rect 7067 6694 7097 6720
rect 7115 6706 7131 6708
rect 7203 6706 7256 6720
rect 7204 6704 7268 6706
rect 7311 6704 7326 6720
rect 7375 6717 7405 6720
rect 7375 6714 7411 6717
rect 7341 6706 7357 6708
rect 7115 6694 7130 6698
rect 7033 6692 7130 6694
rect 7158 6692 7326 6704
rect 7342 6694 7357 6698
rect 7375 6695 7414 6714
rect 7433 6708 7440 6709
rect 7439 6701 7440 6708
rect 7423 6698 7424 6701
rect 7439 6698 7452 6701
rect 7375 6694 7405 6695
rect 7414 6694 7420 6695
rect 7423 6694 7452 6698
rect 7342 6693 7452 6694
rect 7342 6692 7458 6693
rect 7017 6684 7068 6692
rect 7017 6672 7042 6684
rect 7049 6672 7068 6684
rect 7099 6684 7149 6692
rect 7099 6676 7115 6684
rect 7122 6682 7149 6684
rect 7158 6682 7379 6692
rect 7122 6672 7379 6682
rect 7408 6684 7458 6692
rect 7408 6675 7424 6684
rect 7017 6664 7068 6672
rect 7115 6664 7379 6672
rect 7405 6672 7424 6675
rect 7431 6672 7458 6684
rect 7405 6664 7458 6672
rect 7033 6656 7034 6664
rect 7049 6656 7062 6664
rect 7033 6648 7049 6656
rect 7030 6641 7049 6644
rect 7030 6632 7052 6641
rect 7003 6622 7052 6632
rect 7003 6616 7033 6622
rect 7052 6617 7057 6622
rect 6975 6600 7049 6616
rect 7067 6608 7097 6664
rect 7132 6654 7340 6664
rect 7375 6660 7420 6664
rect 7423 6663 7424 6664
rect 7439 6663 7452 6664
rect 7158 6624 7347 6654
rect 7173 6621 7347 6624
rect 7166 6618 7347 6621
rect 6975 6598 6988 6600
rect 7003 6598 7037 6600
rect 6975 6582 7049 6598
rect 7076 6594 7089 6608
rect 7104 6594 7120 6610
rect 7166 6605 7177 6618
rect 6959 6560 6960 6576
rect 6975 6560 6988 6582
rect 7003 6560 7033 6582
rect 7076 6578 7138 6594
rect 7166 6587 7177 6603
rect 7182 6598 7192 6618
rect 7202 6598 7216 6618
rect 7219 6605 7228 6618
rect 7244 6605 7253 6618
rect 7182 6587 7216 6598
rect 7219 6587 7228 6603
rect 7244 6587 7253 6603
rect 7260 6598 7270 6618
rect 7280 6598 7294 6618
rect 7295 6605 7306 6618
rect 7260 6587 7294 6598
rect 7295 6587 7306 6603
rect 7352 6594 7368 6610
rect 7375 6608 7405 6660
rect 7439 6656 7440 6663
rect 7424 6648 7440 6656
rect 7411 6616 7424 6635
rect 7439 6616 7469 6632
rect 7411 6600 7485 6616
rect 7411 6598 7424 6600
rect 7439 6598 7473 6600
rect 7076 6576 7089 6578
rect 7104 6576 7138 6578
rect 7076 6560 7138 6576
rect 7182 6571 7198 6574
rect 7260 6571 7290 6582
rect 7338 6578 7384 6594
rect 7411 6582 7485 6598
rect 7338 6576 7372 6578
rect 7337 6560 7384 6576
rect 7411 6560 7424 6582
rect 7439 6560 7469 6582
rect 7496 6560 7497 6576
rect 7512 6560 7525 6720
rect 7555 6616 7568 6720
rect 7613 6698 7614 6708
rect 7629 6698 7642 6708
rect 7613 6694 7642 6698
rect 7647 6694 7677 6720
rect 7695 6706 7711 6708
rect 7783 6706 7836 6720
rect 7784 6704 7848 6706
rect 7891 6704 7906 6720
rect 7955 6717 7985 6720
rect 7955 6714 7991 6717
rect 7921 6706 7937 6708
rect 7695 6694 7710 6698
rect 7613 6692 7710 6694
rect 7738 6692 7906 6704
rect 7922 6694 7937 6698
rect 7955 6695 7994 6714
rect 8013 6708 8020 6709
rect 8019 6701 8020 6708
rect 8003 6698 8004 6701
rect 8019 6698 8032 6701
rect 7955 6694 7985 6695
rect 7994 6694 8000 6695
rect 8003 6694 8032 6698
rect 7922 6693 8032 6694
rect 7922 6692 8038 6693
rect 7597 6684 7648 6692
rect 7597 6672 7622 6684
rect 7629 6672 7648 6684
rect 7679 6684 7729 6692
rect 7679 6676 7695 6684
rect 7702 6682 7729 6684
rect 7738 6682 7959 6692
rect 7702 6672 7959 6682
rect 7988 6684 8038 6692
rect 7988 6675 8004 6684
rect 7597 6664 7648 6672
rect 7695 6664 7959 6672
rect 7985 6672 8004 6675
rect 8011 6672 8038 6684
rect 7985 6664 8038 6672
rect 7613 6656 7614 6664
rect 7629 6656 7642 6664
rect 7613 6648 7629 6656
rect 7610 6641 7629 6644
rect 7610 6632 7632 6641
rect 7583 6622 7632 6632
rect 7583 6616 7613 6622
rect 7632 6617 7637 6622
rect 7555 6600 7629 6616
rect 7647 6608 7677 6664
rect 7712 6654 7920 6664
rect 7955 6660 8000 6664
rect 8003 6663 8004 6664
rect 8019 6663 8032 6664
rect 7738 6624 7927 6654
rect 7753 6621 7927 6624
rect 7746 6618 7927 6621
rect 7555 6598 7568 6600
rect 7583 6598 7617 6600
rect 7555 6582 7629 6598
rect 7656 6594 7669 6608
rect 7684 6594 7700 6610
rect 7746 6605 7757 6618
rect 7539 6560 7540 6576
rect 7555 6560 7568 6582
rect 7583 6560 7613 6582
rect 7656 6578 7718 6594
rect 7746 6587 7757 6603
rect 7762 6598 7772 6618
rect 7782 6598 7796 6618
rect 7799 6605 7808 6618
rect 7824 6605 7833 6618
rect 7762 6587 7796 6598
rect 7799 6587 7808 6603
rect 7824 6587 7833 6603
rect 7840 6598 7850 6618
rect 7860 6598 7874 6618
rect 7875 6605 7886 6618
rect 7840 6587 7874 6598
rect 7875 6587 7886 6603
rect 7932 6594 7948 6610
rect 7955 6608 7985 6660
rect 8019 6656 8020 6663
rect 8004 6648 8020 6656
rect 7991 6616 8004 6635
rect 8019 6616 8049 6632
rect 7991 6600 8065 6616
rect 7991 6598 8004 6600
rect 8019 6598 8053 6600
rect 7656 6576 7669 6578
rect 7684 6576 7718 6578
rect 7656 6560 7718 6576
rect 7762 6571 7778 6574
rect 7840 6571 7870 6582
rect 7918 6578 7964 6594
rect 7991 6582 8065 6598
rect 7918 6576 7952 6578
rect 7917 6560 7964 6576
rect 7991 6560 8004 6582
rect 8019 6560 8049 6582
rect 8076 6560 8077 6576
rect 8092 6560 8105 6720
rect 8135 6616 8148 6720
rect 8193 6698 8194 6708
rect 8209 6698 8222 6708
rect 8193 6694 8222 6698
rect 8227 6694 8257 6720
rect 8275 6706 8291 6708
rect 8363 6706 8416 6720
rect 8364 6704 8428 6706
rect 8471 6704 8486 6720
rect 8535 6717 8565 6720
rect 8535 6714 8571 6717
rect 8501 6706 8517 6708
rect 8275 6694 8290 6698
rect 8193 6692 8290 6694
rect 8318 6692 8486 6704
rect 8502 6694 8517 6698
rect 8535 6695 8574 6714
rect 8593 6708 8600 6709
rect 8599 6701 8600 6708
rect 8583 6698 8584 6701
rect 8599 6698 8612 6701
rect 8535 6694 8565 6695
rect 8574 6694 8580 6695
rect 8583 6694 8612 6698
rect 8502 6693 8612 6694
rect 8502 6692 8618 6693
rect 8177 6684 8228 6692
rect 8177 6672 8202 6684
rect 8209 6672 8228 6684
rect 8259 6684 8309 6692
rect 8259 6676 8275 6684
rect 8282 6682 8309 6684
rect 8318 6682 8539 6692
rect 8282 6672 8539 6682
rect 8568 6684 8618 6692
rect 8568 6675 8584 6684
rect 8177 6664 8228 6672
rect 8275 6664 8539 6672
rect 8565 6672 8584 6675
rect 8591 6672 8618 6684
rect 8565 6664 8618 6672
rect 8193 6656 8194 6664
rect 8209 6656 8222 6664
rect 8193 6648 8209 6656
rect 8190 6641 8209 6644
rect 8190 6632 8212 6641
rect 8163 6622 8212 6632
rect 8163 6616 8193 6622
rect 8212 6617 8217 6622
rect 8135 6600 8209 6616
rect 8227 6608 8257 6664
rect 8292 6654 8500 6664
rect 8535 6660 8580 6664
rect 8583 6663 8584 6664
rect 8599 6663 8612 6664
rect 8318 6624 8507 6654
rect 8333 6621 8507 6624
rect 8326 6618 8507 6621
rect 8135 6598 8148 6600
rect 8163 6598 8197 6600
rect 8135 6582 8209 6598
rect 8236 6594 8249 6608
rect 8264 6594 8280 6610
rect 8326 6605 8337 6618
rect 8119 6560 8120 6576
rect 8135 6560 8148 6582
rect 8163 6560 8193 6582
rect 8236 6578 8298 6594
rect 8326 6587 8337 6603
rect 8342 6598 8352 6618
rect 8362 6598 8376 6618
rect 8379 6605 8388 6618
rect 8404 6605 8413 6618
rect 8342 6587 8376 6598
rect 8379 6587 8388 6603
rect 8404 6587 8413 6603
rect 8420 6598 8430 6618
rect 8440 6598 8454 6618
rect 8455 6605 8466 6618
rect 8420 6587 8454 6598
rect 8455 6587 8466 6603
rect 8512 6594 8528 6610
rect 8535 6608 8565 6660
rect 8599 6656 8600 6663
rect 8584 6648 8600 6656
rect 8571 6616 8584 6635
rect 8599 6616 8629 6632
rect 8571 6600 8645 6616
rect 8571 6598 8584 6600
rect 8599 6598 8633 6600
rect 8236 6576 8249 6578
rect 8264 6576 8298 6578
rect 8236 6560 8298 6576
rect 8342 6571 8358 6574
rect 8420 6571 8450 6582
rect 8498 6578 8544 6594
rect 8571 6582 8645 6598
rect 8498 6576 8532 6578
rect 8497 6560 8544 6576
rect 8571 6560 8584 6582
rect 8599 6560 8629 6582
rect 8656 6560 8657 6576
rect 8672 6560 8685 6720
rect 8715 6616 8728 6720
rect 8773 6698 8774 6708
rect 8789 6698 8802 6708
rect 8773 6694 8802 6698
rect 8807 6694 8837 6720
rect 8855 6706 8871 6708
rect 8943 6706 8996 6720
rect 8944 6704 9008 6706
rect 9051 6704 9066 6720
rect 9115 6717 9145 6720
rect 9115 6714 9151 6717
rect 9081 6706 9097 6708
rect 8855 6694 8870 6698
rect 8773 6692 8870 6694
rect 8898 6692 9066 6704
rect 9082 6694 9097 6698
rect 9115 6695 9154 6714
rect 9173 6708 9180 6709
rect 9179 6701 9180 6708
rect 9163 6698 9164 6701
rect 9179 6698 9192 6701
rect 9115 6694 9145 6695
rect 9154 6694 9160 6695
rect 9163 6694 9192 6698
rect 9082 6693 9192 6694
rect 9082 6692 9198 6693
rect 8757 6684 8808 6692
rect 8757 6672 8782 6684
rect 8789 6672 8808 6684
rect 8839 6684 8889 6692
rect 8839 6676 8855 6684
rect 8862 6682 8889 6684
rect 8898 6682 9119 6692
rect 8862 6672 9119 6682
rect 9148 6684 9198 6692
rect 9148 6675 9164 6684
rect 8757 6664 8808 6672
rect 8855 6664 9119 6672
rect 9145 6672 9164 6675
rect 9171 6672 9198 6684
rect 9145 6664 9198 6672
rect 8773 6656 8774 6664
rect 8789 6656 8802 6664
rect 8773 6648 8789 6656
rect 8770 6641 8789 6644
rect 8770 6632 8792 6641
rect 8743 6622 8792 6632
rect 8743 6616 8773 6622
rect 8792 6617 8797 6622
rect 8715 6600 8789 6616
rect 8807 6608 8837 6664
rect 8872 6654 9080 6664
rect 9115 6660 9160 6664
rect 9163 6663 9164 6664
rect 9179 6663 9192 6664
rect 8898 6624 9087 6654
rect 8913 6621 9087 6624
rect 8906 6618 9087 6621
rect 8715 6598 8728 6600
rect 8743 6598 8777 6600
rect 8715 6582 8789 6598
rect 8816 6594 8829 6608
rect 8844 6594 8860 6610
rect 8906 6605 8917 6618
rect 8699 6560 8700 6576
rect 8715 6560 8728 6582
rect 8743 6560 8773 6582
rect 8816 6578 8878 6594
rect 8906 6587 8917 6603
rect 8922 6598 8932 6618
rect 8942 6598 8956 6618
rect 8959 6605 8968 6618
rect 8984 6605 8993 6618
rect 8922 6587 8956 6598
rect 8959 6587 8968 6603
rect 8984 6587 8993 6603
rect 9000 6598 9010 6618
rect 9020 6598 9034 6618
rect 9035 6605 9046 6618
rect 9000 6587 9034 6598
rect 9035 6587 9046 6603
rect 9092 6594 9108 6610
rect 9115 6608 9145 6660
rect 9179 6656 9180 6663
rect 9164 6648 9180 6656
rect 9151 6616 9164 6635
rect 9179 6616 9209 6632
rect 9151 6600 9225 6616
rect 9151 6598 9164 6600
rect 9179 6598 9213 6600
rect 8816 6576 8829 6578
rect 8844 6576 8878 6578
rect 8816 6560 8878 6576
rect 8922 6571 8938 6574
rect 9000 6571 9030 6582
rect 9078 6578 9124 6594
rect 9151 6582 9225 6598
rect 9078 6576 9112 6578
rect 9077 6560 9124 6576
rect 9151 6560 9164 6582
rect 9179 6560 9209 6582
rect 9236 6560 9237 6576
rect 9252 6560 9265 6720
rect -7 6552 34 6560
rect -7 6526 8 6552
rect 15 6526 34 6552
rect 98 6548 160 6560
rect 172 6548 247 6560
rect 305 6548 380 6560
rect 392 6548 423 6560
rect 429 6548 464 6560
rect 98 6546 260 6548
rect -7 6518 34 6526
rect 116 6522 129 6546
rect 144 6544 159 6546
rect -1 6508 0 6518
rect 15 6508 28 6518
rect 43 6508 73 6522
rect 116 6508 159 6522
rect 183 6519 190 6526
rect 193 6522 260 6546
rect 292 6546 464 6548
rect 262 6524 290 6528
rect 292 6524 372 6546
rect 393 6544 408 6546
rect 262 6522 372 6524
rect 193 6518 372 6522
rect 166 6508 196 6518
rect 198 6508 351 6518
rect 359 6508 389 6518
rect 393 6508 423 6522
rect 451 6508 464 6546
rect 536 6552 571 6560
rect 536 6526 537 6552
rect 544 6526 571 6552
rect 479 6508 509 6522
rect 536 6518 571 6526
rect 573 6552 614 6560
rect 573 6526 588 6552
rect 595 6526 614 6552
rect 678 6548 740 6560
rect 752 6548 827 6560
rect 885 6548 960 6560
rect 972 6548 1003 6560
rect 1009 6548 1044 6560
rect 678 6546 840 6548
rect 573 6518 614 6526
rect 696 6522 709 6546
rect 724 6544 739 6546
rect 536 6508 537 6518
rect 552 6508 565 6518
rect 579 6508 580 6518
rect 595 6508 608 6518
rect 623 6508 653 6522
rect 696 6508 739 6522
rect 763 6519 770 6526
rect 773 6522 840 6546
rect 872 6546 1044 6548
rect 842 6524 870 6528
rect 872 6524 952 6546
rect 973 6544 988 6546
rect 842 6522 952 6524
rect 773 6518 952 6522
rect 746 6508 776 6518
rect 778 6508 931 6518
rect 939 6508 969 6518
rect 973 6508 1003 6522
rect 1031 6508 1044 6546
rect 1116 6552 1151 6560
rect 1116 6526 1117 6552
rect 1124 6526 1151 6552
rect 1059 6508 1089 6522
rect 1116 6518 1151 6526
rect 1153 6552 1194 6560
rect 1153 6526 1168 6552
rect 1175 6526 1194 6552
rect 1258 6548 1320 6560
rect 1332 6548 1407 6560
rect 1465 6548 1540 6560
rect 1552 6548 1583 6560
rect 1589 6548 1624 6560
rect 1258 6546 1420 6548
rect 1153 6518 1194 6526
rect 1276 6522 1289 6546
rect 1304 6544 1319 6546
rect 1116 6508 1117 6518
rect 1132 6508 1145 6518
rect 1159 6508 1160 6518
rect 1175 6508 1188 6518
rect 1203 6508 1233 6522
rect 1276 6508 1319 6522
rect 1343 6519 1350 6526
rect 1353 6522 1420 6546
rect 1452 6546 1624 6548
rect 1422 6524 1450 6528
rect 1452 6524 1532 6546
rect 1553 6544 1568 6546
rect 1422 6522 1532 6524
rect 1353 6518 1532 6522
rect 1326 6508 1356 6518
rect 1358 6508 1511 6518
rect 1519 6508 1549 6518
rect 1553 6508 1583 6522
rect 1611 6508 1624 6546
rect 1696 6552 1731 6560
rect 1696 6526 1697 6552
rect 1704 6526 1731 6552
rect 1639 6508 1669 6522
rect 1696 6518 1731 6526
rect 1733 6552 1774 6560
rect 1733 6526 1748 6552
rect 1755 6526 1774 6552
rect 1838 6548 1900 6560
rect 1912 6548 1987 6560
rect 2045 6548 2120 6560
rect 2132 6548 2163 6560
rect 2169 6548 2204 6560
rect 1838 6546 2000 6548
rect 1733 6518 1774 6526
rect 1856 6522 1869 6546
rect 1884 6544 1899 6546
rect 1696 6508 1697 6518
rect 1712 6508 1725 6518
rect 1739 6508 1740 6518
rect 1755 6508 1768 6518
rect 1783 6508 1813 6522
rect 1856 6508 1899 6522
rect 1923 6519 1930 6526
rect 1933 6522 2000 6546
rect 2032 6546 2204 6548
rect 2002 6524 2030 6528
rect 2032 6524 2112 6546
rect 2133 6544 2148 6546
rect 2002 6522 2112 6524
rect 1933 6518 2112 6522
rect 1906 6508 1936 6518
rect 1938 6508 2091 6518
rect 2099 6508 2129 6518
rect 2133 6508 2163 6522
rect 2191 6508 2204 6546
rect 2276 6552 2311 6560
rect 2276 6526 2277 6552
rect 2284 6526 2311 6552
rect 2219 6508 2249 6522
rect 2276 6518 2311 6526
rect 2313 6552 2354 6560
rect 2313 6526 2328 6552
rect 2335 6526 2354 6552
rect 2418 6548 2480 6560
rect 2492 6548 2567 6560
rect 2625 6548 2700 6560
rect 2712 6548 2743 6560
rect 2749 6548 2784 6560
rect 2418 6546 2580 6548
rect 2313 6518 2354 6526
rect 2436 6522 2449 6546
rect 2464 6544 2479 6546
rect 2276 6508 2277 6518
rect 2292 6508 2305 6518
rect 2319 6508 2320 6518
rect 2335 6508 2348 6518
rect 2363 6508 2393 6522
rect 2436 6508 2479 6522
rect 2503 6519 2510 6526
rect 2513 6522 2580 6546
rect 2612 6546 2784 6548
rect 2582 6524 2610 6528
rect 2612 6524 2692 6546
rect 2713 6544 2728 6546
rect 2582 6522 2692 6524
rect 2513 6518 2692 6522
rect 2486 6508 2516 6518
rect 2518 6508 2671 6518
rect 2679 6508 2709 6518
rect 2713 6508 2743 6522
rect 2771 6508 2784 6546
rect 2856 6552 2891 6560
rect 2856 6526 2857 6552
rect 2864 6526 2891 6552
rect 2799 6508 2829 6522
rect 2856 6518 2891 6526
rect 2893 6552 2934 6560
rect 2893 6526 2908 6552
rect 2915 6526 2934 6552
rect 2998 6548 3060 6560
rect 3072 6548 3147 6560
rect 3205 6548 3280 6560
rect 3292 6548 3323 6560
rect 3329 6548 3364 6560
rect 2998 6546 3160 6548
rect 2893 6518 2934 6526
rect 3016 6522 3029 6546
rect 3044 6544 3059 6546
rect 2856 6508 2857 6518
rect 2872 6508 2885 6518
rect 2899 6508 2900 6518
rect 2915 6508 2928 6518
rect 2943 6508 2973 6522
rect 3016 6508 3059 6522
rect 3083 6519 3090 6526
rect 3093 6522 3160 6546
rect 3192 6546 3364 6548
rect 3162 6524 3190 6528
rect 3192 6524 3272 6546
rect 3293 6544 3308 6546
rect 3162 6522 3272 6524
rect 3093 6518 3272 6522
rect 3066 6508 3096 6518
rect 3098 6508 3251 6518
rect 3259 6508 3289 6518
rect 3293 6508 3323 6522
rect 3351 6508 3364 6546
rect 3436 6552 3471 6560
rect 3436 6526 3437 6552
rect 3444 6526 3471 6552
rect 3379 6508 3409 6522
rect 3436 6518 3471 6526
rect 3473 6552 3514 6560
rect 3473 6526 3488 6552
rect 3495 6526 3514 6552
rect 3578 6548 3640 6560
rect 3652 6548 3727 6560
rect 3785 6548 3860 6560
rect 3872 6548 3903 6560
rect 3909 6548 3944 6560
rect 3578 6546 3740 6548
rect 3473 6518 3514 6526
rect 3596 6522 3609 6546
rect 3624 6544 3639 6546
rect 3436 6508 3437 6518
rect 3452 6508 3465 6518
rect 3479 6508 3480 6518
rect 3495 6508 3508 6518
rect 3523 6508 3553 6522
rect 3596 6508 3639 6522
rect 3663 6519 3670 6526
rect 3673 6522 3740 6546
rect 3772 6546 3944 6548
rect 3742 6524 3770 6528
rect 3772 6524 3852 6546
rect 3873 6544 3888 6546
rect 3742 6522 3852 6524
rect 3673 6518 3852 6522
rect 3646 6508 3676 6518
rect 3678 6508 3831 6518
rect 3839 6508 3869 6518
rect 3873 6508 3903 6522
rect 3931 6508 3944 6546
rect 4016 6552 4051 6560
rect 4016 6526 4017 6552
rect 4024 6526 4051 6552
rect 3959 6508 3989 6522
rect 4016 6518 4051 6526
rect 4053 6552 4094 6560
rect 4053 6526 4068 6552
rect 4075 6526 4094 6552
rect 4158 6548 4220 6560
rect 4232 6548 4307 6560
rect 4365 6548 4440 6560
rect 4452 6548 4483 6560
rect 4489 6548 4524 6560
rect 4158 6546 4320 6548
rect 4053 6518 4094 6526
rect 4176 6522 4189 6546
rect 4204 6544 4219 6546
rect 4016 6508 4017 6518
rect 4032 6508 4045 6518
rect 4059 6508 4060 6518
rect 4075 6508 4088 6518
rect 4103 6508 4133 6522
rect 4176 6508 4219 6522
rect 4243 6519 4250 6526
rect 4253 6522 4320 6546
rect 4352 6546 4524 6548
rect 4322 6524 4350 6528
rect 4352 6524 4432 6546
rect 4453 6544 4468 6546
rect 4322 6522 4432 6524
rect 4253 6518 4432 6522
rect 4226 6508 4256 6518
rect 4258 6508 4411 6518
rect 4419 6508 4449 6518
rect 4453 6508 4483 6522
rect 4511 6508 4524 6546
rect 4596 6552 4631 6560
rect 4596 6526 4597 6552
rect 4604 6526 4631 6552
rect 4539 6508 4569 6522
rect 4596 6518 4631 6526
rect 4633 6552 4674 6560
rect 4633 6526 4648 6552
rect 4655 6526 4674 6552
rect 4738 6548 4800 6560
rect 4812 6548 4887 6560
rect 4945 6548 5020 6560
rect 5032 6548 5063 6560
rect 5069 6548 5104 6560
rect 4738 6546 4900 6548
rect 4633 6518 4674 6526
rect 4756 6522 4769 6546
rect 4784 6544 4799 6546
rect 4596 6508 4597 6518
rect 4612 6508 4625 6518
rect 4639 6508 4640 6518
rect 4655 6508 4668 6518
rect 4683 6508 4713 6522
rect 4756 6508 4799 6522
rect 4823 6519 4830 6526
rect 4833 6522 4900 6546
rect 4932 6546 5104 6548
rect 4902 6524 4930 6528
rect 4932 6524 5012 6546
rect 5033 6544 5048 6546
rect 4902 6522 5012 6524
rect 4833 6518 5012 6522
rect 4806 6508 4836 6518
rect 4838 6508 4991 6518
rect 4999 6508 5029 6518
rect 5033 6508 5063 6522
rect 5091 6508 5104 6546
rect 5176 6552 5211 6560
rect 5176 6526 5177 6552
rect 5184 6526 5211 6552
rect 5119 6508 5149 6522
rect 5176 6518 5211 6526
rect 5213 6552 5254 6560
rect 5213 6526 5228 6552
rect 5235 6526 5254 6552
rect 5318 6548 5380 6560
rect 5392 6548 5467 6560
rect 5525 6548 5600 6560
rect 5612 6548 5643 6560
rect 5649 6548 5684 6560
rect 5318 6546 5480 6548
rect 5213 6518 5254 6526
rect 5336 6522 5349 6546
rect 5364 6544 5379 6546
rect 5176 6508 5177 6518
rect 5192 6508 5205 6518
rect 5219 6508 5220 6518
rect 5235 6508 5248 6518
rect 5263 6508 5293 6522
rect 5336 6508 5379 6522
rect 5403 6519 5410 6526
rect 5413 6522 5480 6546
rect 5512 6546 5684 6548
rect 5482 6524 5510 6528
rect 5512 6524 5592 6546
rect 5613 6544 5628 6546
rect 5482 6522 5592 6524
rect 5413 6518 5592 6522
rect 5386 6508 5416 6518
rect 5418 6508 5571 6518
rect 5579 6508 5609 6518
rect 5613 6508 5643 6522
rect 5671 6508 5684 6546
rect 5756 6552 5791 6560
rect 5756 6526 5757 6552
rect 5764 6526 5791 6552
rect 5699 6508 5729 6522
rect 5756 6518 5791 6526
rect 5793 6552 5834 6560
rect 5793 6526 5808 6552
rect 5815 6526 5834 6552
rect 5898 6548 5960 6560
rect 5972 6548 6047 6560
rect 6105 6548 6180 6560
rect 6192 6548 6223 6560
rect 6229 6548 6264 6560
rect 5898 6546 6060 6548
rect 5793 6518 5834 6526
rect 5916 6522 5929 6546
rect 5944 6544 5959 6546
rect 5756 6508 5757 6518
rect 5772 6508 5785 6518
rect 5799 6508 5800 6518
rect 5815 6508 5828 6518
rect 5843 6508 5873 6522
rect 5916 6508 5959 6522
rect 5983 6519 5990 6526
rect 5993 6522 6060 6546
rect 6092 6546 6264 6548
rect 6062 6524 6090 6528
rect 6092 6524 6172 6546
rect 6193 6544 6208 6546
rect 6062 6522 6172 6524
rect 5993 6518 6172 6522
rect 5966 6508 5996 6518
rect 5998 6508 6151 6518
rect 6159 6508 6189 6518
rect 6193 6508 6223 6522
rect 6251 6508 6264 6546
rect 6336 6552 6371 6560
rect 6336 6526 6337 6552
rect 6344 6526 6371 6552
rect 6279 6508 6309 6522
rect 6336 6518 6371 6526
rect 6373 6552 6414 6560
rect 6373 6526 6388 6552
rect 6395 6526 6414 6552
rect 6478 6548 6540 6560
rect 6552 6548 6627 6560
rect 6685 6548 6760 6560
rect 6772 6548 6803 6560
rect 6809 6548 6844 6560
rect 6478 6546 6640 6548
rect 6373 6518 6414 6526
rect 6496 6522 6509 6546
rect 6524 6544 6539 6546
rect 6336 6508 6337 6518
rect 6352 6508 6365 6518
rect 6379 6508 6380 6518
rect 6395 6508 6408 6518
rect 6423 6508 6453 6522
rect 6496 6508 6539 6522
rect 6563 6519 6570 6526
rect 6573 6522 6640 6546
rect 6672 6546 6844 6548
rect 6642 6524 6670 6528
rect 6672 6524 6752 6546
rect 6773 6544 6788 6546
rect 6642 6522 6752 6524
rect 6573 6518 6752 6522
rect 6546 6508 6576 6518
rect 6578 6508 6731 6518
rect 6739 6508 6769 6518
rect 6773 6508 6803 6522
rect 6831 6508 6844 6546
rect 6916 6552 6951 6560
rect 6916 6526 6917 6552
rect 6924 6526 6951 6552
rect 6859 6508 6889 6522
rect 6916 6518 6951 6526
rect 6953 6552 6994 6560
rect 6953 6526 6968 6552
rect 6975 6526 6994 6552
rect 7058 6548 7120 6560
rect 7132 6548 7207 6560
rect 7265 6548 7340 6560
rect 7352 6548 7383 6560
rect 7389 6548 7424 6560
rect 7058 6546 7220 6548
rect 6953 6518 6994 6526
rect 7076 6522 7089 6546
rect 7104 6544 7119 6546
rect 6916 6508 6917 6518
rect 6932 6508 6945 6518
rect 6959 6508 6960 6518
rect 6975 6508 6988 6518
rect 7003 6508 7033 6522
rect 7076 6508 7119 6522
rect 7143 6519 7150 6526
rect 7153 6522 7220 6546
rect 7252 6546 7424 6548
rect 7222 6524 7250 6528
rect 7252 6524 7332 6546
rect 7353 6544 7368 6546
rect 7222 6522 7332 6524
rect 7153 6518 7332 6522
rect 7126 6508 7156 6518
rect 7158 6508 7311 6518
rect 7319 6508 7349 6518
rect 7353 6508 7383 6522
rect 7411 6508 7424 6546
rect 7496 6552 7531 6560
rect 7496 6526 7497 6552
rect 7504 6526 7531 6552
rect 7439 6508 7469 6522
rect 7496 6518 7531 6526
rect 7533 6552 7574 6560
rect 7533 6526 7548 6552
rect 7555 6526 7574 6552
rect 7638 6548 7700 6560
rect 7712 6548 7787 6560
rect 7845 6548 7920 6560
rect 7932 6548 7963 6560
rect 7969 6548 8004 6560
rect 7638 6546 7800 6548
rect 7533 6518 7574 6526
rect 7656 6522 7669 6546
rect 7684 6544 7699 6546
rect 7496 6508 7497 6518
rect 7512 6508 7525 6518
rect 7539 6508 7540 6518
rect 7555 6508 7568 6518
rect 7583 6508 7613 6522
rect 7656 6508 7699 6522
rect 7723 6519 7730 6526
rect 7733 6522 7800 6546
rect 7832 6546 8004 6548
rect 7802 6524 7830 6528
rect 7832 6524 7912 6546
rect 7933 6544 7948 6546
rect 7802 6522 7912 6524
rect 7733 6518 7912 6522
rect 7706 6508 7736 6518
rect 7738 6508 7891 6518
rect 7899 6508 7929 6518
rect 7933 6508 7963 6522
rect 7991 6508 8004 6546
rect 8076 6552 8111 6560
rect 8076 6526 8077 6552
rect 8084 6526 8111 6552
rect 8019 6508 8049 6522
rect 8076 6518 8111 6526
rect 8113 6552 8154 6560
rect 8113 6526 8128 6552
rect 8135 6526 8154 6552
rect 8218 6548 8280 6560
rect 8292 6548 8367 6560
rect 8425 6548 8500 6560
rect 8512 6548 8543 6560
rect 8549 6548 8584 6560
rect 8218 6546 8380 6548
rect 8113 6518 8154 6526
rect 8236 6522 8249 6546
rect 8264 6544 8279 6546
rect 8076 6508 8077 6518
rect 8092 6508 8105 6518
rect 8119 6508 8120 6518
rect 8135 6508 8148 6518
rect 8163 6508 8193 6522
rect 8236 6508 8279 6522
rect 8303 6519 8310 6526
rect 8313 6522 8380 6546
rect 8412 6546 8584 6548
rect 8382 6524 8410 6528
rect 8412 6524 8492 6546
rect 8513 6544 8528 6546
rect 8382 6522 8492 6524
rect 8313 6518 8492 6522
rect 8286 6508 8316 6518
rect 8318 6508 8471 6518
rect 8479 6508 8509 6518
rect 8513 6508 8543 6522
rect 8571 6508 8584 6546
rect 8656 6552 8691 6560
rect 8656 6526 8657 6552
rect 8664 6526 8691 6552
rect 8599 6508 8629 6522
rect 8656 6518 8691 6526
rect 8693 6552 8734 6560
rect 8693 6526 8708 6552
rect 8715 6526 8734 6552
rect 8798 6548 8860 6560
rect 8872 6548 8947 6560
rect 9005 6548 9080 6560
rect 9092 6548 9123 6560
rect 9129 6548 9164 6560
rect 8798 6546 8960 6548
rect 8693 6518 8734 6526
rect 8816 6522 8829 6546
rect 8844 6544 8859 6546
rect 8656 6508 8657 6518
rect 8672 6508 8685 6518
rect 8699 6508 8700 6518
rect 8715 6508 8728 6518
rect 8743 6508 8773 6522
rect 8816 6508 8859 6522
rect 8883 6519 8890 6526
rect 8893 6522 8960 6546
rect 8992 6546 9164 6548
rect 8962 6524 8990 6528
rect 8992 6524 9072 6546
rect 9093 6544 9108 6546
rect 8962 6522 9072 6524
rect 8893 6518 9072 6522
rect 8866 6508 8896 6518
rect 8898 6508 9051 6518
rect 9059 6508 9089 6518
rect 9093 6508 9123 6522
rect 9151 6508 9164 6546
rect 9236 6552 9271 6560
rect 9236 6526 9237 6552
rect 9244 6526 9271 6552
rect 9179 6508 9209 6522
rect 9236 6518 9271 6526
rect 9236 6508 9237 6518
rect 9252 6508 9265 6518
rect -1 6502 9265 6508
rect 0 6494 9265 6502
rect 15 6464 28 6494
rect 43 6476 73 6494
rect 116 6480 130 6494
rect 166 6480 386 6494
rect 117 6478 130 6480
rect 83 6466 98 6478
rect 80 6464 102 6466
rect 107 6464 137 6478
rect 198 6476 351 6480
rect 180 6464 372 6476
rect 415 6464 445 6478
rect 451 6464 464 6494
rect 479 6476 509 6494
rect 552 6464 565 6494
rect 595 6464 608 6494
rect 623 6476 653 6494
rect 696 6480 710 6494
rect 746 6480 966 6494
rect 697 6478 710 6480
rect 663 6466 678 6478
rect 660 6464 682 6466
rect 687 6464 717 6478
rect 778 6476 931 6480
rect 760 6464 952 6476
rect 995 6464 1025 6478
rect 1031 6464 1044 6494
rect 1059 6476 1089 6494
rect 1132 6464 1145 6494
rect 1175 6464 1188 6494
rect 1203 6476 1233 6494
rect 1276 6480 1290 6494
rect 1326 6480 1546 6494
rect 1277 6478 1290 6480
rect 1243 6466 1258 6478
rect 1240 6464 1262 6466
rect 1267 6464 1297 6478
rect 1358 6476 1511 6480
rect 1340 6464 1532 6476
rect 1575 6464 1605 6478
rect 1611 6464 1624 6494
rect 1639 6476 1669 6494
rect 1712 6464 1725 6494
rect 1755 6464 1768 6494
rect 1783 6476 1813 6494
rect 1856 6480 1870 6494
rect 1906 6480 2126 6494
rect 1857 6478 1870 6480
rect 1823 6466 1838 6478
rect 1820 6464 1842 6466
rect 1847 6464 1877 6478
rect 1938 6476 2091 6480
rect 1920 6464 2112 6476
rect 2155 6464 2185 6478
rect 2191 6464 2204 6494
rect 2219 6476 2249 6494
rect 2292 6464 2305 6494
rect 2335 6464 2348 6494
rect 2363 6476 2393 6494
rect 2436 6480 2450 6494
rect 2486 6480 2706 6494
rect 2437 6478 2450 6480
rect 2403 6466 2418 6478
rect 2400 6464 2422 6466
rect 2427 6464 2457 6478
rect 2518 6476 2671 6480
rect 2500 6464 2692 6476
rect 2735 6464 2765 6478
rect 2771 6464 2784 6494
rect 2799 6476 2829 6494
rect 2872 6464 2885 6494
rect 2915 6464 2928 6494
rect 2943 6476 2973 6494
rect 3016 6480 3030 6494
rect 3066 6480 3286 6494
rect 3017 6478 3030 6480
rect 2983 6466 2998 6478
rect 2980 6464 3002 6466
rect 3007 6464 3037 6478
rect 3098 6476 3251 6480
rect 3080 6464 3272 6476
rect 3315 6464 3345 6478
rect 3351 6464 3364 6494
rect 3379 6476 3409 6494
rect 3452 6464 3465 6494
rect 3495 6464 3508 6494
rect 3523 6476 3553 6494
rect 3596 6480 3610 6494
rect 3646 6480 3866 6494
rect 3597 6478 3610 6480
rect 3563 6466 3578 6478
rect 3560 6464 3582 6466
rect 3587 6464 3617 6478
rect 3678 6476 3831 6480
rect 3660 6464 3852 6476
rect 3895 6464 3925 6478
rect 3931 6464 3944 6494
rect 3959 6476 3989 6494
rect 4032 6464 4045 6494
rect 4075 6464 4088 6494
rect 4103 6476 4133 6494
rect 4176 6480 4190 6494
rect 4226 6480 4446 6494
rect 4177 6478 4190 6480
rect 4143 6466 4158 6478
rect 4140 6464 4162 6466
rect 4167 6464 4197 6478
rect 4258 6476 4411 6480
rect 4240 6464 4432 6476
rect 4475 6464 4505 6478
rect 4511 6464 4524 6494
rect 4539 6476 4569 6494
rect 4612 6464 4625 6494
rect 4655 6464 4668 6494
rect 4683 6476 4713 6494
rect 4756 6480 4770 6494
rect 4806 6480 5026 6494
rect 4757 6478 4770 6480
rect 4723 6466 4738 6478
rect 4720 6464 4742 6466
rect 4747 6464 4777 6478
rect 4838 6476 4991 6480
rect 4820 6464 5012 6476
rect 5055 6464 5085 6478
rect 5091 6464 5104 6494
rect 5119 6476 5149 6494
rect 5192 6464 5205 6494
rect 5235 6464 5248 6494
rect 5263 6476 5293 6494
rect 5336 6480 5350 6494
rect 5386 6480 5606 6494
rect 5337 6478 5350 6480
rect 5303 6466 5318 6478
rect 5300 6464 5322 6466
rect 5327 6464 5357 6478
rect 5418 6476 5571 6480
rect 5400 6464 5592 6476
rect 5635 6464 5665 6478
rect 5671 6464 5684 6494
rect 5699 6476 5729 6494
rect 5772 6464 5785 6494
rect 5815 6464 5828 6494
rect 5843 6476 5873 6494
rect 5916 6480 5930 6494
rect 5966 6480 6186 6494
rect 5917 6478 5930 6480
rect 5883 6466 5898 6478
rect 5880 6464 5902 6466
rect 5907 6464 5937 6478
rect 5998 6476 6151 6480
rect 5980 6464 6172 6476
rect 6215 6464 6245 6478
rect 6251 6464 6264 6494
rect 6279 6476 6309 6494
rect 6352 6464 6365 6494
rect 6395 6464 6408 6494
rect 6423 6476 6453 6494
rect 6496 6480 6510 6494
rect 6546 6480 6766 6494
rect 6497 6478 6510 6480
rect 6463 6466 6478 6478
rect 6460 6464 6482 6466
rect 6487 6464 6517 6478
rect 6578 6476 6731 6480
rect 6560 6464 6752 6476
rect 6795 6464 6825 6478
rect 6831 6464 6844 6494
rect 6859 6476 6889 6494
rect 6932 6464 6945 6494
rect 6975 6464 6988 6494
rect 7003 6476 7033 6494
rect 7076 6480 7090 6494
rect 7126 6480 7346 6494
rect 7077 6478 7090 6480
rect 7043 6466 7058 6478
rect 7040 6464 7062 6466
rect 7067 6464 7097 6478
rect 7158 6476 7311 6480
rect 7140 6464 7332 6476
rect 7375 6464 7405 6478
rect 7411 6464 7424 6494
rect 7439 6476 7469 6494
rect 7512 6464 7525 6494
rect 7555 6464 7568 6494
rect 7583 6476 7613 6494
rect 7656 6480 7670 6494
rect 7706 6480 7926 6494
rect 7657 6478 7670 6480
rect 7623 6466 7638 6478
rect 7620 6464 7642 6466
rect 7647 6464 7677 6478
rect 7738 6476 7891 6480
rect 7720 6464 7912 6476
rect 7955 6464 7985 6478
rect 7991 6464 8004 6494
rect 8019 6476 8049 6494
rect 8092 6464 8105 6494
rect 8135 6464 8148 6494
rect 8163 6476 8193 6494
rect 8236 6480 8250 6494
rect 8286 6480 8506 6494
rect 8237 6478 8250 6480
rect 8203 6466 8218 6478
rect 8200 6464 8222 6466
rect 8227 6464 8257 6478
rect 8318 6476 8471 6480
rect 8300 6464 8492 6476
rect 8535 6464 8565 6478
rect 8571 6464 8584 6494
rect 8599 6476 8629 6494
rect 8672 6464 8685 6494
rect 8715 6464 8728 6494
rect 8743 6476 8773 6494
rect 8816 6480 8830 6494
rect 8866 6480 9086 6494
rect 8817 6478 8830 6480
rect 8783 6466 8798 6478
rect 8780 6464 8802 6466
rect 8807 6464 8837 6478
rect 8898 6476 9051 6480
rect 8880 6464 9072 6476
rect 9115 6464 9145 6478
rect 9151 6464 9164 6494
rect 9179 6476 9209 6494
rect 9252 6464 9265 6494
rect 0 6450 9265 6464
rect 15 6346 28 6450
rect 73 6428 74 6438
rect 89 6428 102 6438
rect 73 6424 102 6428
rect 107 6424 137 6450
rect 155 6436 171 6438
rect 243 6436 296 6450
rect 244 6434 308 6436
rect 351 6434 366 6450
rect 415 6447 445 6450
rect 415 6444 451 6447
rect 381 6436 397 6438
rect 155 6424 170 6428
rect 73 6422 170 6424
rect 198 6422 366 6434
rect 382 6424 397 6428
rect 415 6425 454 6444
rect 473 6438 480 6439
rect 479 6431 480 6438
rect 463 6428 464 6431
rect 479 6428 492 6431
rect 415 6424 445 6425
rect 454 6424 460 6425
rect 463 6424 492 6428
rect 382 6423 492 6424
rect 382 6422 498 6423
rect 57 6414 108 6422
rect 57 6402 82 6414
rect 89 6402 108 6414
rect 139 6414 189 6422
rect 139 6406 155 6414
rect 162 6412 189 6414
rect 198 6412 419 6422
rect 162 6402 419 6412
rect 448 6414 498 6422
rect 448 6405 464 6414
rect 57 6394 108 6402
rect 155 6394 419 6402
rect 445 6402 464 6405
rect 471 6402 498 6414
rect 445 6394 498 6402
rect 73 6386 74 6394
rect 89 6386 102 6394
rect 73 6378 89 6386
rect 70 6371 89 6374
rect 70 6362 92 6371
rect 43 6352 92 6362
rect 43 6346 73 6352
rect 92 6347 97 6352
rect 15 6330 89 6346
rect 107 6338 137 6394
rect 172 6384 380 6394
rect 415 6390 460 6394
rect 463 6393 464 6394
rect 479 6393 492 6394
rect 198 6354 387 6384
rect 213 6351 387 6354
rect 206 6348 387 6351
rect 15 6328 28 6330
rect 43 6328 77 6330
rect 15 6312 89 6328
rect 116 6324 129 6338
rect 144 6324 160 6340
rect 206 6335 217 6348
rect -1 6290 0 6306
rect 15 6290 28 6312
rect 43 6290 73 6312
rect 116 6308 178 6324
rect 206 6317 217 6333
rect 222 6328 232 6348
rect 242 6328 256 6348
rect 259 6335 268 6348
rect 284 6335 293 6348
rect 222 6317 256 6328
rect 259 6317 268 6333
rect 284 6317 293 6333
rect 300 6328 310 6348
rect 320 6328 334 6348
rect 335 6335 346 6348
rect 300 6317 334 6328
rect 335 6317 346 6333
rect 392 6324 408 6340
rect 415 6338 445 6390
rect 479 6386 480 6393
rect 464 6378 480 6386
rect 451 6346 464 6365
rect 479 6346 509 6362
rect 451 6330 525 6346
rect 451 6328 464 6330
rect 479 6328 513 6330
rect 116 6306 129 6308
rect 144 6306 178 6308
rect 116 6290 178 6306
rect 222 6301 238 6304
rect 300 6301 330 6312
rect 378 6308 424 6324
rect 451 6312 525 6328
rect 378 6306 412 6308
rect 377 6290 424 6306
rect 451 6290 464 6312
rect 479 6290 509 6312
rect 536 6290 537 6306
rect 552 6290 565 6450
rect 595 6346 608 6450
rect 653 6428 654 6438
rect 669 6428 682 6438
rect 653 6424 682 6428
rect 687 6424 717 6450
rect 735 6436 751 6438
rect 823 6436 876 6450
rect 824 6434 888 6436
rect 931 6434 946 6450
rect 995 6447 1025 6450
rect 995 6444 1031 6447
rect 961 6436 977 6438
rect 735 6424 750 6428
rect 653 6422 750 6424
rect 778 6422 946 6434
rect 962 6424 977 6428
rect 995 6425 1034 6444
rect 1053 6438 1060 6439
rect 1059 6431 1060 6438
rect 1043 6428 1044 6431
rect 1059 6428 1072 6431
rect 995 6424 1025 6425
rect 1034 6424 1040 6425
rect 1043 6424 1072 6428
rect 962 6423 1072 6424
rect 962 6422 1078 6423
rect 637 6414 688 6422
rect 637 6402 662 6414
rect 669 6402 688 6414
rect 719 6414 769 6422
rect 719 6406 735 6414
rect 742 6412 769 6414
rect 778 6412 999 6422
rect 742 6402 999 6412
rect 1028 6414 1078 6422
rect 1028 6405 1044 6414
rect 637 6394 688 6402
rect 735 6394 999 6402
rect 1025 6402 1044 6405
rect 1051 6402 1078 6414
rect 1025 6394 1078 6402
rect 653 6386 654 6394
rect 669 6386 682 6394
rect 653 6378 669 6386
rect 650 6371 669 6374
rect 650 6362 672 6371
rect 623 6352 672 6362
rect 623 6346 653 6352
rect 672 6347 677 6352
rect 595 6330 669 6346
rect 687 6338 717 6394
rect 752 6384 960 6394
rect 995 6390 1040 6394
rect 1043 6393 1044 6394
rect 1059 6393 1072 6394
rect 778 6354 967 6384
rect 793 6351 967 6354
rect 786 6348 967 6351
rect 595 6328 608 6330
rect 623 6328 657 6330
rect 595 6312 669 6328
rect 696 6324 709 6338
rect 724 6324 740 6340
rect 786 6335 797 6348
rect 579 6290 580 6306
rect 595 6290 608 6312
rect 623 6290 653 6312
rect 696 6308 758 6324
rect 786 6317 797 6333
rect 802 6328 812 6348
rect 822 6328 836 6348
rect 839 6335 848 6348
rect 864 6335 873 6348
rect 802 6317 836 6328
rect 839 6317 848 6333
rect 864 6317 873 6333
rect 880 6328 890 6348
rect 900 6328 914 6348
rect 915 6335 926 6348
rect 880 6317 914 6328
rect 915 6317 926 6333
rect 972 6324 988 6340
rect 995 6338 1025 6390
rect 1059 6386 1060 6393
rect 1044 6378 1060 6386
rect 1031 6346 1044 6365
rect 1059 6346 1089 6362
rect 1031 6330 1105 6346
rect 1031 6328 1044 6330
rect 1059 6328 1093 6330
rect 696 6306 709 6308
rect 724 6306 758 6308
rect 696 6290 758 6306
rect 802 6301 818 6304
rect 880 6301 910 6312
rect 958 6308 1004 6324
rect 1031 6312 1105 6328
rect 958 6306 992 6308
rect 957 6290 1004 6306
rect 1031 6290 1044 6312
rect 1059 6290 1089 6312
rect 1116 6290 1117 6306
rect 1132 6290 1145 6450
rect 1175 6346 1188 6450
rect 1233 6428 1234 6438
rect 1249 6428 1262 6438
rect 1233 6424 1262 6428
rect 1267 6424 1297 6450
rect 1315 6436 1331 6438
rect 1403 6436 1456 6450
rect 1404 6434 1468 6436
rect 1511 6434 1526 6450
rect 1575 6447 1605 6450
rect 1575 6444 1611 6447
rect 1541 6436 1557 6438
rect 1315 6424 1330 6428
rect 1233 6422 1330 6424
rect 1358 6422 1526 6434
rect 1542 6424 1557 6428
rect 1575 6425 1614 6444
rect 1633 6438 1640 6439
rect 1639 6431 1640 6438
rect 1623 6428 1624 6431
rect 1639 6428 1652 6431
rect 1575 6424 1605 6425
rect 1614 6424 1620 6425
rect 1623 6424 1652 6428
rect 1542 6423 1652 6424
rect 1542 6422 1658 6423
rect 1217 6414 1268 6422
rect 1217 6402 1242 6414
rect 1249 6402 1268 6414
rect 1299 6414 1349 6422
rect 1299 6406 1315 6414
rect 1322 6412 1349 6414
rect 1358 6412 1579 6422
rect 1322 6402 1579 6412
rect 1608 6414 1658 6422
rect 1608 6405 1624 6414
rect 1217 6394 1268 6402
rect 1315 6394 1579 6402
rect 1605 6402 1624 6405
rect 1631 6402 1658 6414
rect 1605 6394 1658 6402
rect 1233 6386 1234 6394
rect 1249 6386 1262 6394
rect 1233 6378 1249 6386
rect 1230 6371 1249 6374
rect 1230 6362 1252 6371
rect 1203 6352 1252 6362
rect 1203 6346 1233 6352
rect 1252 6347 1257 6352
rect 1175 6330 1249 6346
rect 1267 6338 1297 6394
rect 1332 6384 1540 6394
rect 1575 6390 1620 6394
rect 1623 6393 1624 6394
rect 1639 6393 1652 6394
rect 1358 6354 1547 6384
rect 1373 6351 1547 6354
rect 1366 6348 1547 6351
rect 1175 6328 1188 6330
rect 1203 6328 1237 6330
rect 1175 6312 1249 6328
rect 1276 6324 1289 6338
rect 1304 6324 1320 6340
rect 1366 6335 1377 6348
rect 1159 6290 1160 6306
rect 1175 6290 1188 6312
rect 1203 6290 1233 6312
rect 1276 6308 1338 6324
rect 1366 6317 1377 6333
rect 1382 6328 1392 6348
rect 1402 6328 1416 6348
rect 1419 6335 1428 6348
rect 1444 6335 1453 6348
rect 1382 6317 1416 6328
rect 1419 6317 1428 6333
rect 1444 6317 1453 6333
rect 1460 6328 1470 6348
rect 1480 6328 1494 6348
rect 1495 6335 1506 6348
rect 1460 6317 1494 6328
rect 1495 6317 1506 6333
rect 1552 6324 1568 6340
rect 1575 6338 1605 6390
rect 1639 6386 1640 6393
rect 1624 6378 1640 6386
rect 1611 6346 1624 6365
rect 1639 6346 1669 6362
rect 1611 6330 1685 6346
rect 1611 6328 1624 6330
rect 1639 6328 1673 6330
rect 1276 6306 1289 6308
rect 1304 6306 1338 6308
rect 1276 6290 1338 6306
rect 1382 6301 1398 6304
rect 1460 6301 1490 6312
rect 1538 6308 1584 6324
rect 1611 6312 1685 6328
rect 1538 6306 1572 6308
rect 1537 6290 1584 6306
rect 1611 6290 1624 6312
rect 1639 6290 1669 6312
rect 1696 6290 1697 6306
rect 1712 6290 1725 6450
rect 1755 6346 1768 6450
rect 1813 6428 1814 6438
rect 1829 6428 1842 6438
rect 1813 6424 1842 6428
rect 1847 6424 1877 6450
rect 1895 6436 1911 6438
rect 1983 6436 2036 6450
rect 1984 6434 2048 6436
rect 2091 6434 2106 6450
rect 2155 6447 2185 6450
rect 2155 6444 2191 6447
rect 2121 6436 2137 6438
rect 1895 6424 1910 6428
rect 1813 6422 1910 6424
rect 1938 6422 2106 6434
rect 2122 6424 2137 6428
rect 2155 6425 2194 6444
rect 2213 6438 2220 6439
rect 2219 6431 2220 6438
rect 2203 6428 2204 6431
rect 2219 6428 2232 6431
rect 2155 6424 2185 6425
rect 2194 6424 2200 6425
rect 2203 6424 2232 6428
rect 2122 6423 2232 6424
rect 2122 6422 2238 6423
rect 1797 6414 1848 6422
rect 1797 6402 1822 6414
rect 1829 6402 1848 6414
rect 1879 6414 1929 6422
rect 1879 6406 1895 6414
rect 1902 6412 1929 6414
rect 1938 6412 2159 6422
rect 1902 6402 2159 6412
rect 2188 6414 2238 6422
rect 2188 6405 2204 6414
rect 1797 6394 1848 6402
rect 1895 6394 2159 6402
rect 2185 6402 2204 6405
rect 2211 6402 2238 6414
rect 2185 6394 2238 6402
rect 1813 6386 1814 6394
rect 1829 6386 1842 6394
rect 1813 6378 1829 6386
rect 1810 6371 1829 6374
rect 1810 6362 1832 6371
rect 1783 6352 1832 6362
rect 1783 6346 1813 6352
rect 1832 6347 1837 6352
rect 1755 6330 1829 6346
rect 1847 6338 1877 6394
rect 1912 6384 2120 6394
rect 2155 6390 2200 6394
rect 2203 6393 2204 6394
rect 2219 6393 2232 6394
rect 1938 6354 2127 6384
rect 1953 6351 2127 6354
rect 1946 6348 2127 6351
rect 1755 6328 1768 6330
rect 1783 6328 1817 6330
rect 1755 6312 1829 6328
rect 1856 6324 1869 6338
rect 1884 6324 1900 6340
rect 1946 6335 1957 6348
rect 1739 6290 1740 6306
rect 1755 6290 1768 6312
rect 1783 6290 1813 6312
rect 1856 6308 1918 6324
rect 1946 6317 1957 6333
rect 1962 6328 1972 6348
rect 1982 6328 1996 6348
rect 1999 6335 2008 6348
rect 2024 6335 2033 6348
rect 1962 6317 1996 6328
rect 1999 6317 2008 6333
rect 2024 6317 2033 6333
rect 2040 6328 2050 6348
rect 2060 6328 2074 6348
rect 2075 6335 2086 6348
rect 2040 6317 2074 6328
rect 2075 6317 2086 6333
rect 2132 6324 2148 6340
rect 2155 6338 2185 6390
rect 2219 6386 2220 6393
rect 2204 6378 2220 6386
rect 2191 6346 2204 6365
rect 2219 6346 2249 6362
rect 2191 6330 2265 6346
rect 2191 6328 2204 6330
rect 2219 6328 2253 6330
rect 1856 6306 1869 6308
rect 1884 6306 1918 6308
rect 1856 6290 1918 6306
rect 1962 6301 1976 6304
rect 2040 6301 2070 6312
rect 2118 6308 2164 6324
rect 2191 6312 2265 6328
rect 2118 6306 2152 6308
rect 2117 6290 2164 6306
rect 2191 6290 2204 6312
rect 2219 6290 2249 6312
rect 2276 6290 2277 6306
rect 2292 6290 2305 6450
rect 2335 6346 2348 6450
rect 2393 6428 2394 6438
rect 2409 6428 2422 6438
rect 2393 6424 2422 6428
rect 2427 6424 2457 6450
rect 2475 6436 2491 6438
rect 2563 6436 2616 6450
rect 2564 6434 2628 6436
rect 2671 6434 2686 6450
rect 2735 6447 2765 6450
rect 2735 6444 2771 6447
rect 2701 6436 2717 6438
rect 2475 6424 2490 6428
rect 2393 6422 2490 6424
rect 2518 6422 2686 6434
rect 2702 6424 2717 6428
rect 2735 6425 2774 6444
rect 2793 6438 2800 6439
rect 2799 6431 2800 6438
rect 2783 6428 2784 6431
rect 2799 6428 2812 6431
rect 2735 6424 2765 6425
rect 2774 6424 2780 6425
rect 2783 6424 2812 6428
rect 2702 6423 2812 6424
rect 2702 6422 2818 6423
rect 2377 6414 2428 6422
rect 2377 6402 2402 6414
rect 2409 6402 2428 6414
rect 2459 6414 2509 6422
rect 2459 6406 2475 6414
rect 2482 6412 2509 6414
rect 2518 6412 2739 6422
rect 2482 6402 2739 6412
rect 2768 6414 2818 6422
rect 2768 6405 2784 6414
rect 2377 6394 2428 6402
rect 2475 6394 2739 6402
rect 2765 6402 2784 6405
rect 2791 6402 2818 6414
rect 2765 6394 2818 6402
rect 2393 6386 2394 6394
rect 2409 6386 2422 6394
rect 2393 6378 2409 6386
rect 2390 6371 2409 6374
rect 2390 6362 2412 6371
rect 2363 6352 2412 6362
rect 2363 6346 2393 6352
rect 2412 6347 2417 6352
rect 2335 6330 2409 6346
rect 2427 6338 2457 6394
rect 2492 6384 2700 6394
rect 2735 6390 2780 6394
rect 2783 6393 2784 6394
rect 2799 6393 2812 6394
rect 2518 6354 2707 6384
rect 2533 6351 2707 6354
rect 2526 6348 2707 6351
rect 2335 6328 2348 6330
rect 2363 6328 2397 6330
rect 2335 6312 2409 6328
rect 2436 6324 2449 6338
rect 2464 6324 2480 6340
rect 2526 6335 2537 6348
rect 2319 6290 2320 6306
rect 2335 6290 2348 6312
rect 2363 6290 2393 6312
rect 2436 6308 2498 6324
rect 2526 6317 2537 6333
rect 2542 6328 2552 6348
rect 2562 6328 2576 6348
rect 2579 6335 2588 6348
rect 2604 6335 2613 6348
rect 2542 6317 2576 6328
rect 2579 6317 2588 6333
rect 2604 6317 2613 6333
rect 2620 6328 2630 6348
rect 2640 6328 2654 6348
rect 2655 6335 2666 6348
rect 2620 6317 2654 6328
rect 2655 6317 2666 6333
rect 2712 6324 2728 6340
rect 2735 6338 2765 6390
rect 2799 6386 2800 6393
rect 2784 6378 2800 6386
rect 2771 6346 2784 6365
rect 2799 6346 2829 6362
rect 2771 6330 2845 6346
rect 2771 6328 2784 6330
rect 2799 6328 2833 6330
rect 2436 6306 2449 6308
rect 2464 6306 2498 6308
rect 2436 6290 2498 6306
rect 2542 6301 2558 6304
rect 2620 6301 2650 6312
rect 2698 6308 2744 6324
rect 2771 6312 2845 6328
rect 2698 6306 2732 6308
rect 2697 6290 2744 6306
rect 2771 6290 2784 6312
rect 2799 6290 2829 6312
rect 2856 6290 2857 6306
rect 2872 6290 2885 6450
rect 2915 6346 2928 6450
rect 2973 6428 2974 6438
rect 2989 6428 3002 6438
rect 2973 6424 3002 6428
rect 3007 6424 3037 6450
rect 3055 6436 3071 6438
rect 3143 6436 3196 6450
rect 3144 6434 3208 6436
rect 3251 6434 3266 6450
rect 3315 6447 3345 6450
rect 3315 6444 3351 6447
rect 3281 6436 3297 6438
rect 3055 6424 3070 6428
rect 2973 6422 3070 6424
rect 3098 6422 3266 6434
rect 3282 6424 3297 6428
rect 3315 6425 3354 6444
rect 3373 6438 3380 6439
rect 3379 6431 3380 6438
rect 3363 6428 3364 6431
rect 3379 6428 3392 6431
rect 3315 6424 3345 6425
rect 3354 6424 3360 6425
rect 3363 6424 3392 6428
rect 3282 6423 3392 6424
rect 3282 6422 3398 6423
rect 2957 6414 3008 6422
rect 2957 6402 2982 6414
rect 2989 6402 3008 6414
rect 3039 6414 3089 6422
rect 3039 6406 3055 6414
rect 3062 6412 3089 6414
rect 3098 6412 3319 6422
rect 3062 6402 3319 6412
rect 3348 6414 3398 6422
rect 3348 6405 3364 6414
rect 2957 6394 3008 6402
rect 3055 6394 3319 6402
rect 3345 6402 3364 6405
rect 3371 6402 3398 6414
rect 3345 6394 3398 6402
rect 2973 6386 2974 6394
rect 2989 6386 3002 6394
rect 2973 6378 2989 6386
rect 2970 6371 2989 6374
rect 2970 6362 2992 6371
rect 2943 6352 2992 6362
rect 2943 6346 2973 6352
rect 2992 6347 2997 6352
rect 2915 6330 2989 6346
rect 3007 6338 3037 6394
rect 3072 6384 3280 6394
rect 3315 6390 3360 6394
rect 3363 6393 3364 6394
rect 3379 6393 3392 6394
rect 3098 6354 3287 6384
rect 3113 6351 3287 6354
rect 3106 6348 3287 6351
rect 2915 6328 2928 6330
rect 2943 6328 2977 6330
rect 2915 6312 2989 6328
rect 3016 6324 3029 6338
rect 3044 6324 3060 6340
rect 3106 6335 3117 6348
rect 2899 6290 2900 6306
rect 2915 6290 2928 6312
rect 2943 6290 2973 6312
rect 3016 6308 3078 6324
rect 3106 6317 3117 6333
rect 3122 6328 3132 6348
rect 3142 6328 3156 6348
rect 3159 6335 3168 6348
rect 3184 6335 3193 6348
rect 3122 6317 3156 6328
rect 3159 6317 3168 6333
rect 3184 6317 3193 6333
rect 3200 6328 3210 6348
rect 3220 6328 3234 6348
rect 3235 6335 3246 6348
rect 3200 6317 3234 6328
rect 3235 6317 3246 6333
rect 3292 6324 3308 6340
rect 3315 6338 3345 6390
rect 3379 6386 3380 6393
rect 3364 6378 3380 6386
rect 3351 6346 3364 6365
rect 3379 6346 3409 6362
rect 3351 6330 3425 6346
rect 3351 6328 3364 6330
rect 3379 6328 3413 6330
rect 3016 6306 3029 6308
rect 3044 6306 3078 6308
rect 3016 6290 3078 6306
rect 3122 6301 3138 6304
rect 3200 6301 3230 6312
rect 3278 6308 3324 6324
rect 3351 6312 3425 6328
rect 3278 6306 3312 6308
rect 3277 6290 3324 6306
rect 3351 6290 3364 6312
rect 3379 6290 3409 6312
rect 3436 6290 3437 6306
rect 3452 6290 3465 6450
rect 3495 6346 3508 6450
rect 3553 6428 3554 6438
rect 3569 6428 3582 6438
rect 3553 6424 3582 6428
rect 3587 6424 3617 6450
rect 3635 6436 3651 6438
rect 3723 6436 3776 6450
rect 3724 6434 3788 6436
rect 3831 6434 3846 6450
rect 3895 6447 3925 6450
rect 3895 6444 3931 6447
rect 3861 6436 3877 6438
rect 3635 6424 3650 6428
rect 3553 6422 3650 6424
rect 3678 6422 3846 6434
rect 3862 6424 3877 6428
rect 3895 6425 3934 6444
rect 3953 6438 3960 6439
rect 3959 6431 3960 6438
rect 3943 6428 3944 6431
rect 3959 6428 3972 6431
rect 3895 6424 3925 6425
rect 3934 6424 3940 6425
rect 3943 6424 3972 6428
rect 3862 6423 3972 6424
rect 3862 6422 3978 6423
rect 3537 6414 3588 6422
rect 3537 6402 3562 6414
rect 3569 6402 3588 6414
rect 3619 6414 3669 6422
rect 3619 6406 3635 6414
rect 3642 6412 3669 6414
rect 3678 6412 3899 6422
rect 3642 6402 3899 6412
rect 3928 6414 3978 6422
rect 3928 6405 3944 6414
rect 3537 6394 3588 6402
rect 3635 6394 3899 6402
rect 3925 6402 3944 6405
rect 3951 6402 3978 6414
rect 3925 6394 3978 6402
rect 3553 6386 3554 6394
rect 3569 6386 3582 6394
rect 3553 6378 3569 6386
rect 3550 6371 3569 6374
rect 3550 6362 3572 6371
rect 3523 6352 3572 6362
rect 3523 6346 3553 6352
rect 3572 6347 3577 6352
rect 3495 6330 3569 6346
rect 3587 6338 3617 6394
rect 3652 6384 3860 6394
rect 3895 6390 3940 6394
rect 3943 6393 3944 6394
rect 3959 6393 3972 6394
rect 3678 6354 3867 6384
rect 3693 6351 3867 6354
rect 3686 6348 3867 6351
rect 3495 6328 3508 6330
rect 3523 6328 3557 6330
rect 3495 6312 3569 6328
rect 3596 6324 3609 6338
rect 3624 6324 3640 6340
rect 3686 6335 3697 6348
rect 3479 6290 3480 6306
rect 3495 6290 3508 6312
rect 3523 6290 3553 6312
rect 3596 6308 3658 6324
rect 3686 6317 3697 6333
rect 3702 6328 3712 6348
rect 3722 6328 3736 6348
rect 3739 6335 3748 6348
rect 3764 6335 3773 6348
rect 3702 6317 3736 6328
rect 3739 6317 3748 6333
rect 3764 6317 3773 6333
rect 3780 6328 3790 6348
rect 3800 6328 3814 6348
rect 3815 6335 3826 6348
rect 3780 6317 3814 6328
rect 3815 6317 3826 6333
rect 3872 6324 3888 6340
rect 3895 6338 3925 6390
rect 3959 6386 3960 6393
rect 3944 6378 3960 6386
rect 3931 6346 3944 6365
rect 3959 6346 3989 6362
rect 3931 6330 4005 6346
rect 3931 6328 3944 6330
rect 3959 6328 3993 6330
rect 3596 6306 3609 6308
rect 3624 6306 3658 6308
rect 3596 6290 3658 6306
rect 3702 6301 3718 6304
rect 3780 6301 3810 6312
rect 3858 6308 3904 6324
rect 3931 6312 4005 6328
rect 3858 6306 3892 6308
rect 3857 6290 3904 6306
rect 3931 6290 3944 6312
rect 3959 6290 3989 6312
rect 4016 6290 4017 6306
rect 4032 6290 4045 6450
rect 4075 6346 4088 6450
rect 4133 6428 4134 6438
rect 4149 6428 4162 6438
rect 4133 6424 4162 6428
rect 4167 6424 4197 6450
rect 4215 6436 4231 6438
rect 4303 6436 4356 6450
rect 4304 6434 4368 6436
rect 4411 6434 4426 6450
rect 4475 6447 4505 6450
rect 4475 6444 4511 6447
rect 4441 6436 4457 6438
rect 4215 6424 4230 6428
rect 4133 6422 4230 6424
rect 4258 6422 4426 6434
rect 4442 6424 4457 6428
rect 4475 6425 4514 6444
rect 4533 6438 4540 6439
rect 4539 6431 4540 6438
rect 4523 6428 4524 6431
rect 4539 6428 4552 6431
rect 4475 6424 4505 6425
rect 4514 6424 4520 6425
rect 4523 6424 4552 6428
rect 4442 6423 4552 6424
rect 4442 6422 4558 6423
rect 4117 6414 4168 6422
rect 4117 6402 4142 6414
rect 4149 6402 4168 6414
rect 4199 6414 4249 6422
rect 4199 6406 4215 6414
rect 4222 6412 4249 6414
rect 4258 6412 4479 6422
rect 4222 6402 4479 6412
rect 4508 6414 4558 6422
rect 4508 6405 4524 6414
rect 4117 6394 4168 6402
rect 4215 6394 4479 6402
rect 4505 6402 4524 6405
rect 4531 6402 4558 6414
rect 4505 6394 4558 6402
rect 4133 6386 4134 6394
rect 4149 6386 4162 6394
rect 4133 6378 4149 6386
rect 4130 6371 4149 6374
rect 4130 6362 4152 6371
rect 4103 6352 4152 6362
rect 4103 6346 4133 6352
rect 4152 6347 4157 6352
rect 4075 6330 4149 6346
rect 4167 6338 4197 6394
rect 4232 6384 4440 6394
rect 4475 6390 4520 6394
rect 4523 6393 4524 6394
rect 4539 6393 4552 6394
rect 4258 6354 4447 6384
rect 4273 6351 4447 6354
rect 4266 6348 4447 6351
rect 4075 6328 4088 6330
rect 4103 6328 4137 6330
rect 4075 6312 4149 6328
rect 4176 6324 4189 6338
rect 4204 6324 4220 6340
rect 4266 6335 4277 6348
rect 4059 6290 4060 6306
rect 4075 6290 4088 6312
rect 4103 6290 4133 6312
rect 4176 6308 4238 6324
rect 4266 6317 4277 6333
rect 4282 6328 4292 6348
rect 4302 6328 4316 6348
rect 4319 6335 4328 6348
rect 4344 6335 4353 6348
rect 4282 6317 4316 6328
rect 4319 6317 4328 6333
rect 4344 6317 4353 6333
rect 4360 6328 4370 6348
rect 4380 6328 4394 6348
rect 4395 6335 4406 6348
rect 4360 6317 4394 6328
rect 4395 6317 4406 6333
rect 4452 6324 4468 6340
rect 4475 6338 4505 6390
rect 4539 6386 4540 6393
rect 4524 6378 4540 6386
rect 4511 6346 4524 6365
rect 4539 6346 4569 6362
rect 4511 6330 4585 6346
rect 4511 6328 4524 6330
rect 4539 6328 4573 6330
rect 4176 6306 4189 6308
rect 4204 6306 4238 6308
rect 4176 6290 4238 6306
rect 4282 6301 4298 6304
rect 4360 6301 4390 6312
rect 4438 6308 4484 6324
rect 4511 6312 4585 6328
rect 4438 6306 4472 6308
rect 4437 6290 4484 6306
rect 4511 6290 4524 6312
rect 4539 6290 4569 6312
rect 4596 6290 4597 6306
rect 4612 6290 4625 6450
rect 4655 6346 4668 6450
rect 4713 6428 4714 6438
rect 4729 6428 4742 6438
rect 4713 6424 4742 6428
rect 4747 6424 4777 6450
rect 4795 6436 4811 6438
rect 4883 6436 4936 6450
rect 4884 6434 4948 6436
rect 4991 6434 5006 6450
rect 5055 6447 5085 6450
rect 5055 6444 5091 6447
rect 5021 6436 5037 6438
rect 4795 6424 4810 6428
rect 4713 6422 4810 6424
rect 4838 6422 5006 6434
rect 5022 6424 5037 6428
rect 5055 6425 5094 6444
rect 5113 6438 5120 6439
rect 5119 6431 5120 6438
rect 5103 6428 5104 6431
rect 5119 6428 5132 6431
rect 5055 6424 5085 6425
rect 5094 6424 5100 6425
rect 5103 6424 5132 6428
rect 5022 6423 5132 6424
rect 5022 6422 5138 6423
rect 4697 6414 4748 6422
rect 4697 6402 4722 6414
rect 4729 6402 4748 6414
rect 4779 6414 4829 6422
rect 4779 6406 4795 6414
rect 4802 6412 4829 6414
rect 4838 6412 5059 6422
rect 4802 6402 5059 6412
rect 5088 6414 5138 6422
rect 5088 6405 5104 6414
rect 4697 6394 4748 6402
rect 4795 6394 5059 6402
rect 5085 6402 5104 6405
rect 5111 6402 5138 6414
rect 5085 6394 5138 6402
rect 4713 6386 4714 6394
rect 4729 6386 4742 6394
rect 4713 6378 4729 6386
rect 4710 6371 4729 6374
rect 4710 6362 4732 6371
rect 4683 6352 4732 6362
rect 4683 6346 4713 6352
rect 4732 6347 4737 6352
rect 4655 6330 4729 6346
rect 4747 6338 4777 6394
rect 4812 6384 5020 6394
rect 5055 6390 5100 6394
rect 5103 6393 5104 6394
rect 5119 6393 5132 6394
rect 4838 6354 5027 6384
rect 4853 6351 5027 6354
rect 4846 6348 5027 6351
rect 4655 6328 4668 6330
rect 4683 6328 4717 6330
rect 4655 6312 4729 6328
rect 4756 6324 4769 6338
rect 4784 6324 4800 6340
rect 4846 6335 4857 6348
rect 4639 6290 4640 6306
rect 4655 6290 4668 6312
rect 4683 6290 4713 6312
rect 4756 6308 4818 6324
rect 4846 6317 4857 6333
rect 4862 6328 4872 6348
rect 4882 6328 4896 6348
rect 4899 6335 4908 6348
rect 4924 6335 4933 6348
rect 4862 6317 4896 6328
rect 4899 6317 4908 6333
rect 4924 6317 4933 6333
rect 4940 6328 4950 6348
rect 4960 6328 4974 6348
rect 4975 6335 4986 6348
rect 4940 6317 4974 6328
rect 4975 6317 4986 6333
rect 5032 6324 5048 6340
rect 5055 6338 5085 6390
rect 5119 6386 5120 6393
rect 5104 6378 5120 6386
rect 5091 6346 5104 6365
rect 5119 6346 5149 6362
rect 5091 6330 5165 6346
rect 5091 6328 5104 6330
rect 5119 6328 5153 6330
rect 4756 6306 4769 6308
rect 4784 6306 4818 6308
rect 4756 6290 4818 6306
rect 4862 6301 4878 6304
rect 4940 6301 4970 6312
rect 5018 6308 5064 6324
rect 5091 6312 5165 6328
rect 5018 6306 5052 6308
rect 5017 6290 5064 6306
rect 5091 6290 5104 6312
rect 5119 6290 5149 6312
rect 5176 6290 5177 6306
rect 5192 6290 5205 6450
rect 5235 6346 5248 6450
rect 5293 6428 5294 6438
rect 5309 6428 5322 6438
rect 5293 6424 5322 6428
rect 5327 6424 5357 6450
rect 5375 6436 5391 6438
rect 5463 6436 5516 6450
rect 5464 6434 5528 6436
rect 5571 6434 5586 6450
rect 5635 6447 5665 6450
rect 5635 6444 5671 6447
rect 5601 6436 5617 6438
rect 5375 6424 5390 6428
rect 5293 6422 5390 6424
rect 5418 6422 5586 6434
rect 5602 6424 5617 6428
rect 5635 6425 5674 6444
rect 5693 6438 5700 6439
rect 5699 6431 5700 6438
rect 5683 6428 5684 6431
rect 5699 6428 5712 6431
rect 5635 6424 5665 6425
rect 5674 6424 5680 6425
rect 5683 6424 5712 6428
rect 5602 6423 5712 6424
rect 5602 6422 5718 6423
rect 5277 6414 5328 6422
rect 5277 6402 5302 6414
rect 5309 6402 5328 6414
rect 5359 6414 5409 6422
rect 5359 6406 5375 6414
rect 5382 6412 5409 6414
rect 5418 6412 5639 6422
rect 5382 6402 5639 6412
rect 5668 6414 5718 6422
rect 5668 6405 5684 6414
rect 5277 6394 5328 6402
rect 5375 6394 5639 6402
rect 5665 6402 5684 6405
rect 5691 6402 5718 6414
rect 5665 6394 5718 6402
rect 5293 6386 5294 6394
rect 5309 6386 5322 6394
rect 5293 6378 5309 6386
rect 5290 6371 5309 6374
rect 5290 6362 5312 6371
rect 5263 6352 5312 6362
rect 5263 6346 5293 6352
rect 5312 6347 5317 6352
rect 5235 6330 5309 6346
rect 5327 6338 5357 6394
rect 5392 6384 5600 6394
rect 5635 6390 5680 6394
rect 5683 6393 5684 6394
rect 5699 6393 5712 6394
rect 5418 6354 5607 6384
rect 5433 6351 5607 6354
rect 5426 6348 5607 6351
rect 5235 6328 5248 6330
rect 5263 6328 5297 6330
rect 5235 6312 5309 6328
rect 5336 6324 5349 6338
rect 5364 6324 5380 6340
rect 5426 6335 5437 6348
rect 5219 6290 5220 6306
rect 5235 6290 5248 6312
rect 5263 6290 5293 6312
rect 5336 6308 5398 6324
rect 5426 6317 5437 6333
rect 5442 6328 5452 6348
rect 5462 6328 5476 6348
rect 5479 6335 5488 6348
rect 5504 6335 5513 6348
rect 5442 6317 5476 6328
rect 5479 6317 5488 6333
rect 5504 6317 5513 6333
rect 5520 6328 5530 6348
rect 5540 6328 5554 6348
rect 5555 6335 5566 6348
rect 5520 6317 5554 6328
rect 5555 6317 5566 6333
rect 5612 6324 5628 6340
rect 5635 6338 5665 6390
rect 5699 6386 5700 6393
rect 5684 6378 5700 6386
rect 5671 6346 5684 6365
rect 5699 6346 5729 6362
rect 5671 6330 5745 6346
rect 5671 6328 5684 6330
rect 5699 6328 5733 6330
rect 5336 6306 5349 6308
rect 5364 6306 5398 6308
rect 5336 6290 5398 6306
rect 5442 6301 5458 6304
rect 5520 6301 5550 6312
rect 5598 6308 5644 6324
rect 5671 6312 5745 6328
rect 5598 6306 5632 6308
rect 5597 6290 5644 6306
rect 5671 6290 5684 6312
rect 5699 6290 5729 6312
rect 5756 6290 5757 6306
rect 5772 6290 5785 6450
rect 5815 6346 5828 6450
rect 5873 6428 5874 6438
rect 5889 6428 5902 6438
rect 5873 6424 5902 6428
rect 5907 6424 5937 6450
rect 5955 6436 5971 6438
rect 6043 6436 6096 6450
rect 6044 6434 6108 6436
rect 6151 6434 6166 6450
rect 6215 6447 6245 6450
rect 6215 6444 6251 6447
rect 6181 6436 6197 6438
rect 5955 6424 5970 6428
rect 5873 6422 5970 6424
rect 5998 6422 6166 6434
rect 6182 6424 6197 6428
rect 6215 6425 6254 6444
rect 6273 6438 6280 6439
rect 6279 6431 6280 6438
rect 6263 6428 6264 6431
rect 6279 6428 6292 6431
rect 6215 6424 6245 6425
rect 6254 6424 6260 6425
rect 6263 6424 6292 6428
rect 6182 6423 6292 6424
rect 6182 6422 6298 6423
rect 5857 6414 5908 6422
rect 5857 6402 5882 6414
rect 5889 6402 5908 6414
rect 5939 6414 5989 6422
rect 5939 6406 5955 6414
rect 5962 6412 5989 6414
rect 5998 6412 6219 6422
rect 5962 6402 6219 6412
rect 6248 6414 6298 6422
rect 6248 6405 6264 6414
rect 5857 6394 5908 6402
rect 5955 6394 6219 6402
rect 6245 6402 6264 6405
rect 6271 6402 6298 6414
rect 6245 6394 6298 6402
rect 5873 6386 5874 6394
rect 5889 6386 5902 6394
rect 5873 6378 5889 6386
rect 5870 6371 5889 6374
rect 5870 6362 5892 6371
rect 5843 6352 5892 6362
rect 5843 6346 5873 6352
rect 5892 6347 5897 6352
rect 5815 6330 5889 6346
rect 5907 6338 5937 6394
rect 5972 6384 6180 6394
rect 6215 6390 6260 6394
rect 6263 6393 6264 6394
rect 6279 6393 6292 6394
rect 5998 6354 6187 6384
rect 6013 6351 6187 6354
rect 6006 6348 6187 6351
rect 5815 6328 5828 6330
rect 5843 6328 5877 6330
rect 5815 6312 5889 6328
rect 5916 6324 5929 6338
rect 5944 6324 5960 6340
rect 6006 6335 6017 6348
rect 5799 6290 5800 6306
rect 5815 6290 5828 6312
rect 5843 6290 5873 6312
rect 5916 6308 5978 6324
rect 6006 6317 6017 6333
rect 6022 6328 6032 6348
rect 6042 6328 6056 6348
rect 6059 6335 6068 6348
rect 6084 6335 6093 6348
rect 6022 6317 6056 6328
rect 6059 6317 6068 6333
rect 6084 6317 6093 6333
rect 6100 6328 6110 6348
rect 6120 6328 6134 6348
rect 6135 6335 6146 6348
rect 6100 6317 6134 6328
rect 6135 6317 6146 6333
rect 6192 6324 6208 6340
rect 6215 6338 6245 6390
rect 6279 6386 6280 6393
rect 6264 6378 6280 6386
rect 6251 6346 6264 6365
rect 6279 6346 6309 6362
rect 6251 6330 6325 6346
rect 6251 6328 6264 6330
rect 6279 6328 6313 6330
rect 5916 6306 5929 6308
rect 5944 6306 5978 6308
rect 5916 6290 5978 6306
rect 6022 6301 6038 6304
rect 6100 6301 6130 6312
rect 6178 6308 6224 6324
rect 6251 6312 6325 6328
rect 6178 6306 6212 6308
rect 6177 6290 6224 6306
rect 6251 6290 6264 6312
rect 6279 6290 6309 6312
rect 6336 6290 6337 6306
rect 6352 6290 6365 6450
rect 6395 6346 6408 6450
rect 6453 6428 6454 6438
rect 6469 6428 6482 6438
rect 6453 6424 6482 6428
rect 6487 6424 6517 6450
rect 6535 6436 6551 6438
rect 6623 6436 6676 6450
rect 6624 6434 6688 6436
rect 6731 6434 6746 6450
rect 6795 6447 6825 6450
rect 6795 6444 6831 6447
rect 6761 6436 6777 6438
rect 6535 6424 6550 6428
rect 6453 6422 6550 6424
rect 6578 6422 6746 6434
rect 6762 6424 6777 6428
rect 6795 6425 6834 6444
rect 6853 6438 6860 6439
rect 6859 6431 6860 6438
rect 6843 6428 6844 6431
rect 6859 6428 6872 6431
rect 6795 6424 6825 6425
rect 6834 6424 6840 6425
rect 6843 6424 6872 6428
rect 6762 6423 6872 6424
rect 6762 6422 6878 6423
rect 6437 6414 6488 6422
rect 6437 6402 6462 6414
rect 6469 6402 6488 6414
rect 6519 6414 6569 6422
rect 6519 6406 6535 6414
rect 6542 6412 6569 6414
rect 6578 6412 6799 6422
rect 6542 6402 6799 6412
rect 6828 6414 6878 6422
rect 6828 6405 6844 6414
rect 6437 6394 6488 6402
rect 6535 6394 6799 6402
rect 6825 6402 6844 6405
rect 6851 6402 6878 6414
rect 6825 6394 6878 6402
rect 6453 6386 6454 6394
rect 6469 6386 6482 6394
rect 6453 6378 6469 6386
rect 6450 6371 6469 6374
rect 6450 6362 6472 6371
rect 6423 6352 6472 6362
rect 6423 6346 6453 6352
rect 6472 6347 6477 6352
rect 6395 6330 6469 6346
rect 6487 6338 6517 6394
rect 6552 6384 6760 6394
rect 6795 6390 6840 6394
rect 6843 6393 6844 6394
rect 6859 6393 6872 6394
rect 6578 6354 6767 6384
rect 6593 6351 6767 6354
rect 6586 6348 6767 6351
rect 6395 6328 6408 6330
rect 6423 6328 6457 6330
rect 6395 6312 6469 6328
rect 6496 6324 6509 6338
rect 6524 6324 6540 6340
rect 6586 6335 6597 6348
rect 6379 6290 6380 6306
rect 6395 6290 6408 6312
rect 6423 6290 6453 6312
rect 6496 6308 6558 6324
rect 6586 6317 6597 6333
rect 6602 6328 6612 6348
rect 6622 6328 6636 6348
rect 6639 6335 6648 6348
rect 6664 6335 6673 6348
rect 6602 6317 6636 6328
rect 6639 6317 6648 6333
rect 6664 6317 6673 6333
rect 6680 6328 6690 6348
rect 6700 6328 6714 6348
rect 6715 6335 6726 6348
rect 6680 6317 6714 6328
rect 6715 6317 6726 6333
rect 6772 6324 6788 6340
rect 6795 6338 6825 6390
rect 6859 6386 6860 6393
rect 6844 6378 6860 6386
rect 6831 6346 6844 6365
rect 6859 6346 6889 6362
rect 6831 6330 6905 6346
rect 6831 6328 6844 6330
rect 6859 6328 6893 6330
rect 6496 6306 6509 6308
rect 6524 6306 6558 6308
rect 6496 6290 6558 6306
rect 6602 6301 6618 6304
rect 6680 6301 6710 6312
rect 6758 6308 6804 6324
rect 6831 6312 6905 6328
rect 6758 6306 6792 6308
rect 6757 6290 6804 6306
rect 6831 6290 6844 6312
rect 6859 6290 6889 6312
rect 6916 6290 6917 6306
rect 6932 6290 6945 6450
rect 6975 6346 6988 6450
rect 7033 6428 7034 6438
rect 7049 6428 7062 6438
rect 7033 6424 7062 6428
rect 7067 6424 7097 6450
rect 7115 6436 7131 6438
rect 7203 6436 7256 6450
rect 7204 6434 7268 6436
rect 7311 6434 7326 6450
rect 7375 6447 7405 6450
rect 7375 6444 7411 6447
rect 7341 6436 7357 6438
rect 7115 6424 7130 6428
rect 7033 6422 7130 6424
rect 7158 6422 7326 6434
rect 7342 6424 7357 6428
rect 7375 6425 7414 6444
rect 7433 6438 7440 6439
rect 7439 6431 7440 6438
rect 7423 6428 7424 6431
rect 7439 6428 7452 6431
rect 7375 6424 7405 6425
rect 7414 6424 7420 6425
rect 7423 6424 7452 6428
rect 7342 6423 7452 6424
rect 7342 6422 7458 6423
rect 7017 6414 7068 6422
rect 7017 6402 7042 6414
rect 7049 6402 7068 6414
rect 7099 6414 7149 6422
rect 7099 6406 7115 6414
rect 7122 6412 7149 6414
rect 7158 6412 7379 6422
rect 7122 6402 7379 6412
rect 7408 6414 7458 6422
rect 7408 6405 7424 6414
rect 7017 6394 7068 6402
rect 7115 6394 7379 6402
rect 7405 6402 7424 6405
rect 7431 6402 7458 6414
rect 7405 6394 7458 6402
rect 7033 6386 7034 6394
rect 7049 6386 7062 6394
rect 7033 6378 7049 6386
rect 7030 6371 7049 6374
rect 7030 6362 7052 6371
rect 7003 6352 7052 6362
rect 7003 6346 7033 6352
rect 7052 6347 7057 6352
rect 6975 6330 7049 6346
rect 7067 6338 7097 6394
rect 7132 6384 7340 6394
rect 7375 6390 7420 6394
rect 7423 6393 7424 6394
rect 7439 6393 7452 6394
rect 7158 6354 7347 6384
rect 7173 6351 7347 6354
rect 7166 6348 7347 6351
rect 6975 6328 6988 6330
rect 7003 6328 7037 6330
rect 6975 6312 7049 6328
rect 7076 6324 7089 6338
rect 7104 6324 7120 6340
rect 7166 6335 7177 6348
rect 6959 6290 6960 6306
rect 6975 6290 6988 6312
rect 7003 6290 7033 6312
rect 7076 6308 7138 6324
rect 7166 6317 7177 6333
rect 7182 6328 7192 6348
rect 7202 6328 7216 6348
rect 7219 6335 7228 6348
rect 7244 6335 7253 6348
rect 7182 6317 7216 6328
rect 7219 6317 7228 6333
rect 7244 6317 7253 6333
rect 7260 6328 7270 6348
rect 7280 6328 7294 6348
rect 7295 6335 7306 6348
rect 7260 6317 7294 6328
rect 7295 6317 7306 6333
rect 7352 6324 7368 6340
rect 7375 6338 7405 6390
rect 7439 6386 7440 6393
rect 7424 6378 7440 6386
rect 7411 6346 7424 6365
rect 7439 6346 7469 6362
rect 7411 6330 7485 6346
rect 7411 6328 7424 6330
rect 7439 6328 7473 6330
rect 7076 6306 7089 6308
rect 7104 6306 7138 6308
rect 7076 6290 7138 6306
rect 7182 6301 7198 6304
rect 7260 6301 7290 6312
rect 7338 6308 7384 6324
rect 7411 6312 7485 6328
rect 7338 6306 7372 6308
rect 7337 6290 7384 6306
rect 7411 6290 7424 6312
rect 7439 6290 7469 6312
rect 7496 6290 7497 6306
rect 7512 6290 7525 6450
rect 7555 6346 7568 6450
rect 7613 6428 7614 6438
rect 7629 6428 7642 6438
rect 7613 6424 7642 6428
rect 7647 6424 7677 6450
rect 7695 6436 7711 6438
rect 7783 6436 7836 6450
rect 7784 6434 7848 6436
rect 7891 6434 7906 6450
rect 7955 6447 7985 6450
rect 7955 6444 7991 6447
rect 7921 6436 7937 6438
rect 7695 6424 7710 6428
rect 7613 6422 7710 6424
rect 7738 6422 7906 6434
rect 7922 6424 7937 6428
rect 7955 6425 7994 6444
rect 8013 6438 8020 6439
rect 8019 6431 8020 6438
rect 8003 6428 8004 6431
rect 8019 6428 8032 6431
rect 7955 6424 7985 6425
rect 7994 6424 8000 6425
rect 8003 6424 8032 6428
rect 7922 6423 8032 6424
rect 7922 6422 8038 6423
rect 7597 6414 7648 6422
rect 7597 6402 7622 6414
rect 7629 6402 7648 6414
rect 7679 6414 7729 6422
rect 7679 6406 7695 6414
rect 7702 6412 7729 6414
rect 7738 6412 7959 6422
rect 7702 6402 7959 6412
rect 7988 6414 8038 6422
rect 7988 6405 8004 6414
rect 7597 6394 7648 6402
rect 7695 6394 7959 6402
rect 7985 6402 8004 6405
rect 8011 6402 8038 6414
rect 7985 6394 8038 6402
rect 7613 6386 7614 6394
rect 7629 6386 7642 6394
rect 7613 6378 7629 6386
rect 7610 6371 7629 6374
rect 7610 6362 7632 6371
rect 7583 6352 7632 6362
rect 7583 6346 7613 6352
rect 7632 6347 7637 6352
rect 7555 6330 7629 6346
rect 7647 6338 7677 6394
rect 7712 6384 7920 6394
rect 7955 6390 8000 6394
rect 8003 6393 8004 6394
rect 8019 6393 8032 6394
rect 7738 6354 7927 6384
rect 7753 6351 7927 6354
rect 7746 6348 7927 6351
rect 7555 6328 7568 6330
rect 7583 6328 7617 6330
rect 7555 6312 7629 6328
rect 7656 6324 7669 6338
rect 7684 6324 7700 6340
rect 7746 6335 7757 6348
rect 7539 6290 7540 6306
rect 7555 6290 7568 6312
rect 7583 6290 7613 6312
rect 7656 6308 7718 6324
rect 7746 6317 7757 6333
rect 7762 6328 7772 6348
rect 7782 6328 7796 6348
rect 7799 6335 7808 6348
rect 7824 6335 7833 6348
rect 7762 6317 7796 6328
rect 7799 6317 7808 6333
rect 7824 6317 7833 6333
rect 7840 6328 7850 6348
rect 7860 6328 7874 6348
rect 7875 6335 7886 6348
rect 7840 6317 7874 6328
rect 7875 6317 7886 6333
rect 7932 6324 7948 6340
rect 7955 6338 7985 6390
rect 8019 6386 8020 6393
rect 8004 6378 8020 6386
rect 7991 6346 8004 6365
rect 8019 6346 8049 6362
rect 7991 6330 8065 6346
rect 7991 6328 8004 6330
rect 8019 6328 8053 6330
rect 7656 6306 7669 6308
rect 7684 6306 7718 6308
rect 7656 6290 7718 6306
rect 7762 6301 7778 6304
rect 7840 6301 7870 6312
rect 7918 6308 7964 6324
rect 7991 6312 8065 6328
rect 7918 6306 7952 6308
rect 7917 6290 7964 6306
rect 7991 6290 8004 6312
rect 8019 6290 8049 6312
rect 8076 6290 8077 6306
rect 8092 6290 8105 6450
rect 8135 6346 8148 6450
rect 8193 6428 8194 6438
rect 8209 6428 8222 6438
rect 8193 6424 8222 6428
rect 8227 6424 8257 6450
rect 8275 6436 8291 6438
rect 8363 6436 8416 6450
rect 8364 6434 8428 6436
rect 8471 6434 8486 6450
rect 8535 6447 8565 6450
rect 8535 6444 8571 6447
rect 8501 6436 8517 6438
rect 8275 6424 8290 6428
rect 8193 6422 8290 6424
rect 8318 6422 8486 6434
rect 8502 6424 8517 6428
rect 8535 6425 8574 6444
rect 8593 6438 8600 6439
rect 8599 6431 8600 6438
rect 8583 6428 8584 6431
rect 8599 6428 8612 6431
rect 8535 6424 8565 6425
rect 8574 6424 8580 6425
rect 8583 6424 8612 6428
rect 8502 6423 8612 6424
rect 8502 6422 8618 6423
rect 8177 6414 8228 6422
rect 8177 6402 8202 6414
rect 8209 6402 8228 6414
rect 8259 6414 8309 6422
rect 8259 6406 8275 6414
rect 8282 6412 8309 6414
rect 8318 6412 8539 6422
rect 8282 6402 8539 6412
rect 8568 6414 8618 6422
rect 8568 6405 8584 6414
rect 8177 6394 8228 6402
rect 8275 6394 8539 6402
rect 8565 6402 8584 6405
rect 8591 6402 8618 6414
rect 8565 6394 8618 6402
rect 8193 6386 8194 6394
rect 8209 6386 8222 6394
rect 8193 6378 8209 6386
rect 8190 6371 8209 6374
rect 8190 6362 8212 6371
rect 8163 6352 8212 6362
rect 8163 6346 8193 6352
rect 8212 6347 8217 6352
rect 8135 6330 8209 6346
rect 8227 6338 8257 6394
rect 8292 6384 8500 6394
rect 8535 6390 8580 6394
rect 8583 6393 8584 6394
rect 8599 6393 8612 6394
rect 8318 6354 8507 6384
rect 8333 6351 8507 6354
rect 8326 6348 8507 6351
rect 8135 6328 8148 6330
rect 8163 6328 8197 6330
rect 8135 6312 8209 6328
rect 8236 6324 8249 6338
rect 8264 6324 8280 6340
rect 8326 6335 8337 6348
rect 8119 6290 8120 6306
rect 8135 6290 8148 6312
rect 8163 6290 8193 6312
rect 8236 6308 8298 6324
rect 8326 6317 8337 6333
rect 8342 6328 8352 6348
rect 8362 6328 8376 6348
rect 8379 6335 8388 6348
rect 8404 6335 8413 6348
rect 8342 6317 8376 6328
rect 8379 6317 8388 6333
rect 8404 6317 8413 6333
rect 8420 6328 8430 6348
rect 8440 6328 8454 6348
rect 8455 6335 8466 6348
rect 8420 6317 8454 6328
rect 8455 6317 8466 6333
rect 8512 6324 8528 6340
rect 8535 6338 8565 6390
rect 8599 6386 8600 6393
rect 8584 6378 8600 6386
rect 8571 6346 8584 6365
rect 8599 6346 8629 6362
rect 8571 6330 8645 6346
rect 8571 6328 8584 6330
rect 8599 6328 8633 6330
rect 8236 6306 8249 6308
rect 8264 6306 8298 6308
rect 8236 6290 8298 6306
rect 8342 6301 8358 6304
rect 8420 6301 8450 6312
rect 8498 6308 8544 6324
rect 8571 6312 8645 6328
rect 8498 6306 8532 6308
rect 8497 6290 8544 6306
rect 8571 6290 8584 6312
rect 8599 6290 8629 6312
rect 8656 6290 8657 6306
rect 8672 6290 8685 6450
rect 8715 6346 8728 6450
rect 8773 6428 8774 6438
rect 8789 6428 8802 6438
rect 8773 6424 8802 6428
rect 8807 6424 8837 6450
rect 8855 6436 8871 6438
rect 8943 6436 8996 6450
rect 8944 6434 9008 6436
rect 9051 6434 9066 6450
rect 9115 6447 9145 6450
rect 9115 6444 9151 6447
rect 9081 6436 9097 6438
rect 8855 6424 8870 6428
rect 8773 6422 8870 6424
rect 8898 6422 9066 6434
rect 9082 6424 9097 6428
rect 9115 6425 9154 6444
rect 9173 6438 9180 6439
rect 9179 6431 9180 6438
rect 9163 6428 9164 6431
rect 9179 6428 9192 6431
rect 9115 6424 9145 6425
rect 9154 6424 9160 6425
rect 9163 6424 9192 6428
rect 9082 6423 9192 6424
rect 9082 6422 9198 6423
rect 8757 6414 8808 6422
rect 8757 6402 8782 6414
rect 8789 6402 8808 6414
rect 8839 6414 8889 6422
rect 8839 6406 8855 6414
rect 8862 6412 8889 6414
rect 8898 6412 9119 6422
rect 8862 6402 9119 6412
rect 9148 6414 9198 6422
rect 9148 6405 9164 6414
rect 8757 6394 8808 6402
rect 8855 6394 9119 6402
rect 9145 6402 9164 6405
rect 9171 6402 9198 6414
rect 9145 6394 9198 6402
rect 8773 6386 8774 6394
rect 8789 6386 8802 6394
rect 8773 6378 8789 6386
rect 8770 6371 8789 6374
rect 8770 6362 8792 6371
rect 8743 6352 8792 6362
rect 8743 6346 8773 6352
rect 8792 6347 8797 6352
rect 8715 6330 8789 6346
rect 8807 6338 8837 6394
rect 8872 6384 9080 6394
rect 9115 6390 9160 6394
rect 9163 6393 9164 6394
rect 9179 6393 9192 6394
rect 8898 6354 9087 6384
rect 8913 6351 9087 6354
rect 8906 6348 9087 6351
rect 8715 6328 8728 6330
rect 8743 6328 8777 6330
rect 8715 6312 8789 6328
rect 8816 6324 8829 6338
rect 8844 6324 8860 6340
rect 8906 6335 8917 6348
rect 8699 6290 8700 6306
rect 8715 6290 8728 6312
rect 8743 6290 8773 6312
rect 8816 6308 8878 6324
rect 8906 6317 8917 6333
rect 8922 6328 8932 6348
rect 8942 6328 8956 6348
rect 8959 6335 8968 6348
rect 8984 6335 8993 6348
rect 8922 6317 8956 6328
rect 8959 6317 8968 6333
rect 8984 6317 8993 6333
rect 9000 6328 9010 6348
rect 9020 6328 9034 6348
rect 9035 6335 9046 6348
rect 9000 6317 9034 6328
rect 9035 6317 9046 6333
rect 9092 6324 9108 6340
rect 9115 6338 9145 6390
rect 9179 6386 9180 6393
rect 9164 6378 9180 6386
rect 9151 6346 9164 6365
rect 9179 6346 9209 6362
rect 9151 6330 9225 6346
rect 9151 6328 9164 6330
rect 9179 6328 9213 6330
rect 8816 6306 8829 6308
rect 8844 6306 8878 6308
rect 8816 6290 8878 6306
rect 8922 6301 8938 6304
rect 9000 6301 9030 6312
rect 9078 6308 9124 6324
rect 9151 6312 9225 6328
rect 9078 6306 9112 6308
rect 9077 6290 9124 6306
rect 9151 6290 9164 6312
rect 9179 6290 9209 6312
rect 9236 6290 9237 6306
rect 9252 6290 9265 6450
rect -7 6282 34 6290
rect -7 6256 8 6282
rect 15 6256 34 6282
rect 98 6278 160 6290
rect 172 6278 247 6290
rect 305 6278 380 6290
rect 392 6278 423 6290
rect 429 6278 464 6290
rect 98 6276 260 6278
rect -7 6248 34 6256
rect 116 6252 129 6276
rect 144 6274 159 6276
rect -1 6238 0 6248
rect 15 6238 28 6248
rect 43 6238 73 6252
rect 116 6238 159 6252
rect 183 6249 190 6256
rect 193 6252 260 6276
rect 292 6276 464 6278
rect 262 6254 290 6258
rect 292 6254 372 6276
rect 393 6274 408 6276
rect 262 6252 372 6254
rect 193 6248 372 6252
rect 166 6238 196 6248
rect 198 6238 351 6248
rect 359 6238 389 6248
rect 393 6238 423 6252
rect 451 6238 464 6276
rect 536 6282 571 6290
rect 536 6256 537 6282
rect 544 6256 571 6282
rect 479 6238 509 6252
rect 536 6248 571 6256
rect 573 6282 614 6290
rect 573 6256 588 6282
rect 595 6256 614 6282
rect 678 6278 740 6290
rect 752 6278 827 6290
rect 885 6278 960 6290
rect 972 6278 1003 6290
rect 1009 6278 1044 6290
rect 678 6276 840 6278
rect 573 6248 614 6256
rect 696 6252 709 6276
rect 724 6274 739 6276
rect 536 6238 537 6248
rect 552 6238 565 6248
rect 579 6238 580 6248
rect 595 6238 608 6248
rect 623 6238 653 6252
rect 696 6238 739 6252
rect 763 6249 770 6256
rect 773 6252 840 6276
rect 872 6276 1044 6278
rect 842 6254 870 6258
rect 872 6254 952 6276
rect 973 6274 988 6276
rect 842 6252 952 6254
rect 773 6248 952 6252
rect 746 6238 776 6248
rect 778 6238 931 6248
rect 939 6238 969 6248
rect 973 6238 1003 6252
rect 1031 6238 1044 6276
rect 1116 6282 1151 6290
rect 1116 6256 1117 6282
rect 1124 6256 1151 6282
rect 1059 6238 1089 6252
rect 1116 6248 1151 6256
rect 1153 6282 1194 6290
rect 1153 6256 1168 6282
rect 1175 6256 1194 6282
rect 1258 6278 1320 6290
rect 1332 6278 1407 6290
rect 1465 6278 1540 6290
rect 1552 6278 1583 6290
rect 1589 6278 1624 6290
rect 1258 6276 1420 6278
rect 1153 6248 1194 6256
rect 1276 6252 1289 6276
rect 1304 6274 1319 6276
rect 1116 6238 1117 6248
rect 1132 6238 1145 6248
rect 1159 6238 1160 6248
rect 1175 6238 1188 6248
rect 1203 6238 1233 6252
rect 1276 6238 1319 6252
rect 1343 6249 1350 6256
rect 1353 6252 1420 6276
rect 1452 6276 1624 6278
rect 1422 6254 1450 6258
rect 1452 6254 1532 6276
rect 1553 6274 1568 6276
rect 1422 6252 1532 6254
rect 1353 6248 1532 6252
rect 1326 6238 1356 6248
rect 1358 6238 1511 6248
rect 1519 6238 1549 6248
rect 1553 6238 1583 6252
rect 1611 6238 1624 6276
rect 1696 6282 1731 6290
rect 1696 6256 1697 6282
rect 1704 6256 1731 6282
rect 1639 6238 1669 6252
rect 1696 6248 1731 6256
rect 1733 6282 1774 6290
rect 1733 6256 1748 6282
rect 1755 6256 1774 6282
rect 1838 6278 1900 6290
rect 1912 6278 1987 6290
rect 2045 6278 2120 6290
rect 2132 6278 2163 6290
rect 2169 6278 2204 6290
rect 1838 6276 2000 6278
rect 1733 6248 1774 6256
rect 1856 6252 1869 6276
rect 1884 6274 1899 6276
rect 1696 6238 1697 6248
rect 1712 6238 1725 6248
rect 1739 6238 1740 6248
rect 1755 6238 1768 6248
rect 1783 6238 1813 6252
rect 1856 6238 1899 6252
rect 1923 6249 1930 6256
rect 1933 6252 2000 6276
rect 2032 6276 2204 6278
rect 2002 6254 2030 6258
rect 2032 6254 2112 6276
rect 2133 6274 2148 6276
rect 2002 6252 2112 6254
rect 1933 6248 2112 6252
rect 1906 6238 1936 6248
rect 1938 6238 2091 6248
rect 2099 6238 2129 6248
rect 2133 6238 2163 6252
rect 2191 6238 2204 6276
rect 2276 6282 2311 6290
rect 2276 6256 2277 6282
rect 2284 6256 2311 6282
rect 2219 6238 2249 6252
rect 2276 6248 2311 6256
rect 2313 6282 2354 6290
rect 2313 6256 2328 6282
rect 2335 6256 2354 6282
rect 2418 6278 2480 6290
rect 2492 6278 2567 6290
rect 2625 6278 2700 6290
rect 2712 6278 2743 6290
rect 2749 6278 2784 6290
rect 2418 6276 2580 6278
rect 2313 6248 2354 6256
rect 2436 6252 2449 6276
rect 2464 6274 2479 6276
rect 2276 6238 2277 6248
rect 2292 6238 2305 6248
rect 2319 6238 2320 6248
rect 2335 6238 2348 6248
rect 2363 6238 2393 6252
rect 2436 6238 2479 6252
rect 2503 6249 2510 6256
rect 2513 6252 2580 6276
rect 2612 6276 2784 6278
rect 2582 6254 2610 6258
rect 2612 6254 2692 6276
rect 2713 6274 2728 6276
rect 2582 6252 2692 6254
rect 2513 6248 2692 6252
rect 2486 6238 2516 6248
rect 2518 6238 2671 6248
rect 2679 6238 2709 6248
rect 2713 6238 2743 6252
rect 2771 6238 2784 6276
rect 2856 6282 2891 6290
rect 2856 6256 2857 6282
rect 2864 6256 2891 6282
rect 2799 6238 2829 6252
rect 2856 6248 2891 6256
rect 2893 6282 2934 6290
rect 2893 6256 2908 6282
rect 2915 6256 2934 6282
rect 2998 6278 3060 6290
rect 3072 6278 3147 6290
rect 3205 6278 3280 6290
rect 3292 6278 3323 6290
rect 3329 6278 3364 6290
rect 2998 6276 3160 6278
rect 2893 6248 2934 6256
rect 3016 6252 3029 6276
rect 3044 6274 3059 6276
rect 2856 6238 2857 6248
rect 2872 6238 2885 6248
rect 2899 6238 2900 6248
rect 2915 6238 2928 6248
rect 2943 6238 2973 6252
rect 3016 6238 3059 6252
rect 3083 6249 3090 6256
rect 3093 6252 3160 6276
rect 3192 6276 3364 6278
rect 3162 6254 3190 6258
rect 3192 6254 3272 6276
rect 3293 6274 3308 6276
rect 3162 6252 3272 6254
rect 3093 6248 3272 6252
rect 3066 6238 3096 6248
rect 3098 6238 3251 6248
rect 3259 6238 3289 6248
rect 3293 6238 3323 6252
rect 3351 6238 3364 6276
rect 3436 6282 3471 6290
rect 3436 6256 3437 6282
rect 3444 6256 3471 6282
rect 3379 6238 3409 6252
rect 3436 6248 3471 6256
rect 3473 6282 3514 6290
rect 3473 6256 3488 6282
rect 3495 6256 3514 6282
rect 3578 6278 3640 6290
rect 3652 6278 3727 6290
rect 3785 6278 3860 6290
rect 3872 6278 3903 6290
rect 3909 6278 3944 6290
rect 3578 6276 3740 6278
rect 3473 6248 3514 6256
rect 3596 6252 3609 6276
rect 3624 6274 3639 6276
rect 3436 6238 3437 6248
rect 3452 6238 3465 6248
rect 3479 6238 3480 6248
rect 3495 6238 3508 6248
rect 3523 6238 3553 6252
rect 3596 6238 3639 6252
rect 3663 6249 3670 6256
rect 3673 6252 3740 6276
rect 3772 6276 3944 6278
rect 3742 6254 3770 6258
rect 3772 6254 3852 6276
rect 3873 6274 3888 6276
rect 3742 6252 3852 6254
rect 3673 6248 3852 6252
rect 3646 6238 3676 6248
rect 3678 6238 3831 6248
rect 3839 6238 3869 6248
rect 3873 6238 3903 6252
rect 3931 6238 3944 6276
rect 4016 6282 4051 6290
rect 4016 6256 4017 6282
rect 4024 6256 4051 6282
rect 3959 6238 3989 6252
rect 4016 6248 4051 6256
rect 4053 6282 4094 6290
rect 4053 6256 4068 6282
rect 4075 6256 4094 6282
rect 4158 6278 4220 6290
rect 4232 6278 4307 6290
rect 4365 6278 4440 6290
rect 4452 6278 4483 6290
rect 4489 6278 4524 6290
rect 4158 6276 4320 6278
rect 4053 6248 4094 6256
rect 4176 6252 4189 6276
rect 4204 6274 4219 6276
rect 4016 6238 4017 6248
rect 4032 6238 4045 6248
rect 4059 6238 4060 6248
rect 4075 6238 4088 6248
rect 4103 6238 4133 6252
rect 4176 6238 4219 6252
rect 4243 6249 4250 6256
rect 4253 6252 4320 6276
rect 4352 6276 4524 6278
rect 4322 6254 4350 6258
rect 4352 6254 4432 6276
rect 4453 6274 4468 6276
rect 4322 6252 4432 6254
rect 4253 6248 4432 6252
rect 4226 6238 4256 6248
rect 4258 6238 4411 6248
rect 4419 6238 4449 6248
rect 4453 6238 4483 6252
rect 4511 6238 4524 6276
rect 4596 6282 4631 6290
rect 4596 6256 4597 6282
rect 4604 6256 4631 6282
rect 4539 6238 4569 6252
rect 4596 6248 4631 6256
rect 4633 6282 4674 6290
rect 4633 6256 4648 6282
rect 4655 6256 4674 6282
rect 4738 6278 4800 6290
rect 4812 6278 4887 6290
rect 4945 6278 5020 6290
rect 5032 6278 5063 6290
rect 5069 6278 5104 6290
rect 4738 6276 4900 6278
rect 4633 6248 4674 6256
rect 4756 6252 4769 6276
rect 4784 6274 4799 6276
rect 4596 6238 4597 6248
rect 4612 6238 4625 6248
rect 4639 6238 4640 6248
rect 4655 6238 4668 6248
rect 4683 6238 4713 6252
rect 4756 6238 4799 6252
rect 4823 6249 4830 6256
rect 4833 6252 4900 6276
rect 4932 6276 5104 6278
rect 4902 6254 4930 6258
rect 4932 6254 5012 6276
rect 5033 6274 5048 6276
rect 4902 6252 5012 6254
rect 4833 6248 5012 6252
rect 4806 6238 4836 6248
rect 4838 6238 4991 6248
rect 4999 6238 5029 6248
rect 5033 6238 5063 6252
rect 5091 6238 5104 6276
rect 5176 6282 5211 6290
rect 5176 6256 5177 6282
rect 5184 6256 5211 6282
rect 5119 6238 5149 6252
rect 5176 6248 5211 6256
rect 5213 6282 5254 6290
rect 5213 6256 5228 6282
rect 5235 6256 5254 6282
rect 5318 6278 5380 6290
rect 5392 6278 5467 6290
rect 5525 6278 5600 6290
rect 5612 6278 5643 6290
rect 5649 6278 5684 6290
rect 5318 6276 5480 6278
rect 5213 6248 5254 6256
rect 5336 6252 5349 6276
rect 5364 6274 5379 6276
rect 5176 6238 5177 6248
rect 5192 6238 5205 6248
rect 5219 6238 5220 6248
rect 5235 6238 5248 6248
rect 5263 6238 5293 6252
rect 5336 6238 5379 6252
rect 5403 6249 5410 6256
rect 5413 6252 5480 6276
rect 5512 6276 5684 6278
rect 5482 6254 5510 6258
rect 5512 6254 5592 6276
rect 5613 6274 5628 6276
rect 5482 6252 5592 6254
rect 5413 6248 5592 6252
rect 5386 6238 5416 6248
rect 5418 6238 5571 6248
rect 5579 6238 5609 6248
rect 5613 6238 5643 6252
rect 5671 6238 5684 6276
rect 5756 6282 5791 6290
rect 5756 6256 5757 6282
rect 5764 6256 5791 6282
rect 5699 6238 5729 6252
rect 5756 6248 5791 6256
rect 5793 6282 5834 6290
rect 5793 6256 5808 6282
rect 5815 6256 5834 6282
rect 5898 6278 5960 6290
rect 5972 6278 6047 6290
rect 6105 6278 6180 6290
rect 6192 6278 6223 6290
rect 6229 6278 6264 6290
rect 5898 6276 6060 6278
rect 5793 6248 5834 6256
rect 5916 6252 5929 6276
rect 5944 6274 5959 6276
rect 5756 6238 5757 6248
rect 5772 6238 5785 6248
rect 5799 6238 5800 6248
rect 5815 6238 5828 6248
rect 5843 6238 5873 6252
rect 5916 6238 5959 6252
rect 5983 6249 5990 6256
rect 5993 6252 6060 6276
rect 6092 6276 6264 6278
rect 6062 6254 6090 6258
rect 6092 6254 6172 6276
rect 6193 6274 6208 6276
rect 6062 6252 6172 6254
rect 5993 6248 6172 6252
rect 5966 6238 5996 6248
rect 5998 6238 6151 6248
rect 6159 6238 6189 6248
rect 6193 6238 6223 6252
rect 6251 6238 6264 6276
rect 6336 6282 6371 6290
rect 6336 6256 6337 6282
rect 6344 6256 6371 6282
rect 6279 6238 6309 6252
rect 6336 6248 6371 6256
rect 6373 6282 6414 6290
rect 6373 6256 6388 6282
rect 6395 6256 6414 6282
rect 6478 6278 6540 6290
rect 6552 6278 6627 6290
rect 6685 6278 6760 6290
rect 6772 6278 6803 6290
rect 6809 6278 6844 6290
rect 6478 6276 6640 6278
rect 6373 6248 6414 6256
rect 6496 6252 6509 6276
rect 6524 6274 6539 6276
rect 6336 6238 6337 6248
rect 6352 6238 6365 6248
rect 6379 6238 6380 6248
rect 6395 6238 6408 6248
rect 6423 6238 6453 6252
rect 6496 6238 6539 6252
rect 6563 6249 6570 6256
rect 6573 6252 6640 6276
rect 6672 6276 6844 6278
rect 6642 6254 6670 6258
rect 6672 6254 6752 6276
rect 6773 6274 6788 6276
rect 6642 6252 6752 6254
rect 6573 6248 6752 6252
rect 6546 6238 6576 6248
rect 6578 6238 6731 6248
rect 6739 6238 6769 6248
rect 6773 6238 6803 6252
rect 6831 6238 6844 6276
rect 6916 6282 6951 6290
rect 6916 6256 6917 6282
rect 6924 6256 6951 6282
rect 6859 6238 6889 6252
rect 6916 6248 6951 6256
rect 6953 6282 6994 6290
rect 6953 6256 6968 6282
rect 6975 6256 6994 6282
rect 7058 6278 7120 6290
rect 7132 6278 7207 6290
rect 7265 6278 7340 6290
rect 7352 6278 7383 6290
rect 7389 6278 7424 6290
rect 7058 6276 7220 6278
rect 6953 6248 6994 6256
rect 7076 6252 7089 6276
rect 7104 6274 7119 6276
rect 6916 6238 6917 6248
rect 6932 6238 6945 6248
rect 6959 6238 6960 6248
rect 6975 6238 6988 6248
rect 7003 6238 7033 6252
rect 7076 6238 7119 6252
rect 7143 6249 7150 6256
rect 7153 6252 7220 6276
rect 7252 6276 7424 6278
rect 7222 6254 7250 6258
rect 7252 6254 7332 6276
rect 7353 6274 7368 6276
rect 7222 6252 7332 6254
rect 7153 6248 7332 6252
rect 7126 6238 7156 6248
rect 7158 6238 7311 6248
rect 7319 6238 7349 6248
rect 7353 6238 7383 6252
rect 7411 6238 7424 6276
rect 7496 6282 7531 6290
rect 7496 6256 7497 6282
rect 7504 6256 7531 6282
rect 7439 6238 7469 6252
rect 7496 6248 7531 6256
rect 7533 6282 7574 6290
rect 7533 6256 7548 6282
rect 7555 6256 7574 6282
rect 7638 6278 7700 6290
rect 7712 6278 7787 6290
rect 7845 6278 7920 6290
rect 7932 6278 7963 6290
rect 7969 6278 8004 6290
rect 7638 6276 7800 6278
rect 7533 6248 7574 6256
rect 7656 6252 7669 6276
rect 7684 6274 7699 6276
rect 7496 6238 7497 6248
rect 7512 6238 7525 6248
rect 7539 6238 7540 6248
rect 7555 6238 7568 6248
rect 7583 6238 7613 6252
rect 7656 6238 7699 6252
rect 7723 6249 7730 6256
rect 7733 6252 7800 6276
rect 7832 6276 8004 6278
rect 7802 6254 7830 6258
rect 7832 6254 7912 6276
rect 7933 6274 7948 6276
rect 7802 6252 7912 6254
rect 7733 6248 7912 6252
rect 7706 6238 7736 6248
rect 7738 6238 7891 6248
rect 7899 6238 7929 6248
rect 7933 6238 7963 6252
rect 7991 6238 8004 6276
rect 8076 6282 8111 6290
rect 8076 6256 8077 6282
rect 8084 6256 8111 6282
rect 8019 6238 8049 6252
rect 8076 6248 8111 6256
rect 8113 6282 8154 6290
rect 8113 6256 8128 6282
rect 8135 6256 8154 6282
rect 8218 6278 8280 6290
rect 8292 6278 8367 6290
rect 8425 6278 8500 6290
rect 8512 6278 8543 6290
rect 8549 6278 8584 6290
rect 8218 6276 8380 6278
rect 8113 6248 8154 6256
rect 8236 6252 8249 6276
rect 8264 6274 8279 6276
rect 8076 6238 8077 6248
rect 8092 6238 8105 6248
rect 8119 6238 8120 6248
rect 8135 6238 8148 6248
rect 8163 6238 8193 6252
rect 8236 6238 8279 6252
rect 8303 6249 8310 6256
rect 8313 6252 8380 6276
rect 8412 6276 8584 6278
rect 8382 6254 8410 6258
rect 8412 6254 8492 6276
rect 8513 6274 8528 6276
rect 8382 6252 8492 6254
rect 8313 6248 8492 6252
rect 8286 6238 8316 6248
rect 8318 6238 8471 6248
rect 8479 6238 8509 6248
rect 8513 6238 8543 6252
rect 8571 6238 8584 6276
rect 8656 6282 8691 6290
rect 8656 6256 8657 6282
rect 8664 6256 8691 6282
rect 8599 6238 8629 6252
rect 8656 6248 8691 6256
rect 8693 6282 8734 6290
rect 8693 6256 8708 6282
rect 8715 6256 8734 6282
rect 8798 6278 8860 6290
rect 8872 6278 8947 6290
rect 9005 6278 9080 6290
rect 9092 6278 9123 6290
rect 9129 6278 9164 6290
rect 8798 6276 8960 6278
rect 8693 6248 8734 6256
rect 8816 6252 8829 6276
rect 8844 6274 8859 6276
rect 8656 6238 8657 6248
rect 8672 6238 8685 6248
rect 8699 6238 8700 6248
rect 8715 6238 8728 6248
rect 8743 6238 8773 6252
rect 8816 6238 8859 6252
rect 8883 6249 8890 6256
rect 8893 6252 8960 6276
rect 8992 6276 9164 6278
rect 8962 6254 8990 6258
rect 8992 6254 9072 6276
rect 9093 6274 9108 6276
rect 8962 6252 9072 6254
rect 8893 6248 9072 6252
rect 8866 6238 8896 6248
rect 8898 6238 9051 6248
rect 9059 6238 9089 6248
rect 9093 6238 9123 6252
rect 9151 6238 9164 6276
rect 9236 6282 9271 6290
rect 9236 6256 9237 6282
rect 9244 6256 9271 6282
rect 9179 6238 9209 6252
rect 9236 6248 9271 6256
rect 9236 6238 9237 6248
rect 9252 6238 9265 6248
rect -1 6232 9265 6238
rect 0 6224 9265 6232
rect 15 6194 28 6224
rect 43 6206 73 6224
rect 116 6210 130 6224
rect 166 6210 386 6224
rect 117 6208 130 6210
rect 83 6196 98 6208
rect 80 6194 102 6196
rect 107 6194 137 6208
rect 198 6206 351 6210
rect 180 6194 372 6206
rect 415 6194 445 6208
rect 451 6194 464 6224
rect 479 6206 509 6224
rect 552 6194 565 6224
rect 595 6194 608 6224
rect 623 6206 653 6224
rect 696 6210 710 6224
rect 746 6210 966 6224
rect 697 6208 710 6210
rect 663 6196 678 6208
rect 660 6194 682 6196
rect 687 6194 717 6208
rect 778 6206 931 6210
rect 760 6194 952 6206
rect 995 6194 1025 6208
rect 1031 6194 1044 6224
rect 1059 6206 1089 6224
rect 1132 6194 1145 6224
rect 1175 6194 1188 6224
rect 1203 6206 1233 6224
rect 1276 6210 1290 6224
rect 1326 6210 1546 6224
rect 1277 6208 1290 6210
rect 1243 6196 1258 6208
rect 1240 6194 1262 6196
rect 1267 6194 1297 6208
rect 1358 6206 1511 6210
rect 1340 6194 1532 6206
rect 1575 6194 1605 6208
rect 1611 6194 1624 6224
rect 1639 6206 1669 6224
rect 1712 6194 1725 6224
rect 1755 6194 1768 6224
rect 1783 6206 1813 6224
rect 1856 6210 1870 6224
rect 1906 6210 2126 6224
rect 1857 6208 1870 6210
rect 1823 6196 1838 6208
rect 1820 6194 1842 6196
rect 1847 6194 1877 6208
rect 1938 6206 2091 6210
rect 1920 6194 2112 6206
rect 2155 6194 2185 6208
rect 2191 6194 2204 6224
rect 2219 6206 2249 6224
rect 2292 6194 2305 6224
rect 2335 6194 2348 6224
rect 2363 6206 2393 6224
rect 2436 6210 2450 6224
rect 2486 6210 2706 6224
rect 2437 6208 2450 6210
rect 2403 6196 2418 6208
rect 2400 6194 2422 6196
rect 2427 6194 2457 6208
rect 2518 6206 2671 6210
rect 2500 6194 2692 6206
rect 2735 6194 2765 6208
rect 2771 6194 2784 6224
rect 2799 6206 2829 6224
rect 2872 6194 2885 6224
rect 2915 6194 2928 6224
rect 2943 6206 2973 6224
rect 3016 6210 3030 6224
rect 3066 6210 3286 6224
rect 3017 6208 3030 6210
rect 2983 6196 2998 6208
rect 2980 6194 3002 6196
rect 3007 6194 3037 6208
rect 3098 6206 3251 6210
rect 3080 6194 3272 6206
rect 3315 6194 3345 6208
rect 3351 6194 3364 6224
rect 3379 6206 3409 6224
rect 3452 6194 3465 6224
rect 3495 6194 3508 6224
rect 3523 6206 3553 6224
rect 3596 6210 3610 6224
rect 3646 6210 3866 6224
rect 3597 6208 3610 6210
rect 3563 6196 3578 6208
rect 3560 6194 3582 6196
rect 3587 6194 3617 6208
rect 3678 6206 3831 6210
rect 3660 6194 3852 6206
rect 3895 6194 3925 6208
rect 3931 6194 3944 6224
rect 3959 6206 3989 6224
rect 4032 6194 4045 6224
rect 4075 6194 4088 6224
rect 4103 6206 4133 6224
rect 4176 6210 4190 6224
rect 4226 6210 4446 6224
rect 4177 6208 4190 6210
rect 4143 6196 4158 6208
rect 4140 6194 4162 6196
rect 4167 6194 4197 6208
rect 4258 6206 4411 6210
rect 4240 6194 4432 6206
rect 4475 6194 4505 6208
rect 4511 6194 4524 6224
rect 4539 6206 4569 6224
rect 4612 6194 4625 6224
rect 4655 6194 4668 6224
rect 4683 6206 4713 6224
rect 4756 6210 4770 6224
rect 4806 6210 5026 6224
rect 4757 6208 4770 6210
rect 4723 6196 4738 6208
rect 4720 6194 4742 6196
rect 4747 6194 4777 6208
rect 4838 6206 4991 6210
rect 4820 6194 5012 6206
rect 5055 6194 5085 6208
rect 5091 6194 5104 6224
rect 5119 6206 5149 6224
rect 5192 6194 5205 6224
rect 5235 6194 5248 6224
rect 5263 6206 5293 6224
rect 5336 6210 5350 6224
rect 5386 6210 5606 6224
rect 5337 6208 5350 6210
rect 5303 6196 5318 6208
rect 5300 6194 5322 6196
rect 5327 6194 5357 6208
rect 5418 6206 5571 6210
rect 5400 6194 5592 6206
rect 5635 6194 5665 6208
rect 5671 6194 5684 6224
rect 5699 6206 5729 6224
rect 5772 6194 5785 6224
rect 5815 6194 5828 6224
rect 5843 6206 5873 6224
rect 5916 6210 5930 6224
rect 5966 6210 6186 6224
rect 5917 6208 5930 6210
rect 5883 6196 5898 6208
rect 5880 6194 5902 6196
rect 5907 6194 5937 6208
rect 5998 6206 6151 6210
rect 5980 6194 6172 6206
rect 6215 6194 6245 6208
rect 6251 6194 6264 6224
rect 6279 6206 6309 6224
rect 6352 6194 6365 6224
rect 6395 6194 6408 6224
rect 6423 6206 6453 6224
rect 6496 6210 6510 6224
rect 6546 6210 6766 6224
rect 6497 6208 6510 6210
rect 6463 6196 6478 6208
rect 6460 6194 6482 6196
rect 6487 6194 6517 6208
rect 6578 6206 6731 6210
rect 6560 6194 6752 6206
rect 6795 6194 6825 6208
rect 6831 6194 6844 6224
rect 6859 6206 6889 6224
rect 6932 6194 6945 6224
rect 6975 6194 6988 6224
rect 7003 6206 7033 6224
rect 7076 6210 7090 6224
rect 7126 6210 7346 6224
rect 7077 6208 7090 6210
rect 7043 6196 7058 6208
rect 7040 6194 7062 6196
rect 7067 6194 7097 6208
rect 7158 6206 7311 6210
rect 7140 6194 7332 6206
rect 7375 6194 7405 6208
rect 7411 6194 7424 6224
rect 7439 6206 7469 6224
rect 7512 6194 7525 6224
rect 7555 6194 7568 6224
rect 7583 6206 7613 6224
rect 7656 6210 7670 6224
rect 7706 6210 7926 6224
rect 7657 6208 7670 6210
rect 7623 6196 7638 6208
rect 7620 6194 7642 6196
rect 7647 6194 7677 6208
rect 7738 6206 7891 6210
rect 7720 6194 7912 6206
rect 7955 6194 7985 6208
rect 7991 6194 8004 6224
rect 8019 6206 8049 6224
rect 8092 6194 8105 6224
rect 8135 6194 8148 6224
rect 8163 6206 8193 6224
rect 8236 6210 8250 6224
rect 8286 6210 8506 6224
rect 8237 6208 8250 6210
rect 8203 6196 8218 6208
rect 8200 6194 8222 6196
rect 8227 6194 8257 6208
rect 8318 6206 8471 6210
rect 8300 6194 8492 6206
rect 8535 6194 8565 6208
rect 8571 6194 8584 6224
rect 8599 6206 8629 6224
rect 8672 6194 8685 6224
rect 8715 6194 8728 6224
rect 8743 6206 8773 6224
rect 8816 6210 8830 6224
rect 8866 6210 9086 6224
rect 8817 6208 8830 6210
rect 8783 6196 8798 6208
rect 8780 6194 8802 6196
rect 8807 6194 8837 6208
rect 8898 6206 9051 6210
rect 8880 6194 9072 6206
rect 9115 6194 9145 6208
rect 9151 6194 9164 6224
rect 9179 6206 9209 6224
rect 9252 6194 9265 6224
rect 0 6180 9265 6194
rect 15 6076 28 6180
rect 73 6158 74 6168
rect 89 6158 102 6168
rect 73 6154 102 6158
rect 107 6154 137 6180
rect 155 6166 171 6168
rect 243 6166 296 6180
rect 244 6164 308 6166
rect 351 6164 366 6180
rect 415 6177 445 6180
rect 415 6174 451 6177
rect 381 6166 397 6168
rect 155 6154 170 6158
rect 73 6152 170 6154
rect 198 6152 366 6164
rect 382 6154 397 6158
rect 415 6155 454 6174
rect 473 6168 480 6169
rect 479 6161 480 6168
rect 463 6158 464 6161
rect 479 6158 492 6161
rect 415 6154 445 6155
rect 454 6154 460 6155
rect 463 6154 492 6158
rect 382 6153 492 6154
rect 382 6152 498 6153
rect 57 6144 108 6152
rect 57 6132 82 6144
rect 89 6132 108 6144
rect 139 6144 189 6152
rect 139 6136 155 6144
rect 162 6142 189 6144
rect 198 6142 419 6152
rect 162 6132 419 6142
rect 448 6144 498 6152
rect 448 6135 464 6144
rect 57 6124 108 6132
rect 155 6124 419 6132
rect 445 6132 464 6135
rect 471 6132 498 6144
rect 445 6124 498 6132
rect 73 6116 74 6124
rect 89 6116 102 6124
rect 73 6108 89 6116
rect 70 6101 89 6104
rect 70 6092 92 6101
rect 43 6082 92 6092
rect 43 6076 73 6082
rect 92 6077 97 6082
rect 15 6060 89 6076
rect 107 6068 137 6124
rect 172 6114 380 6124
rect 415 6120 460 6124
rect 463 6123 464 6124
rect 479 6123 492 6124
rect 198 6084 387 6114
rect 213 6081 387 6084
rect 206 6078 387 6081
rect 15 6058 28 6060
rect 43 6058 77 6060
rect 15 6042 89 6058
rect 116 6054 129 6068
rect 144 6054 160 6070
rect 206 6065 217 6078
rect -1 6020 0 6036
rect 15 6020 28 6042
rect 43 6020 73 6042
rect 116 6038 178 6054
rect 206 6047 217 6063
rect 222 6058 232 6078
rect 242 6058 256 6078
rect 259 6065 268 6078
rect 284 6065 293 6078
rect 222 6047 256 6058
rect 259 6047 268 6063
rect 284 6047 293 6063
rect 300 6058 310 6078
rect 320 6058 334 6078
rect 335 6065 346 6078
rect 300 6047 334 6058
rect 335 6047 346 6063
rect 392 6054 408 6070
rect 415 6068 445 6120
rect 479 6116 480 6123
rect 464 6108 480 6116
rect 451 6076 464 6095
rect 479 6076 509 6092
rect 451 6060 525 6076
rect 451 6058 464 6060
rect 479 6058 513 6060
rect 116 6036 129 6038
rect 144 6036 178 6038
rect 116 6020 178 6036
rect 222 6031 238 6034
rect 300 6031 330 6042
rect 378 6038 424 6054
rect 451 6042 525 6058
rect 378 6036 412 6038
rect 377 6020 424 6036
rect 451 6020 464 6042
rect 479 6020 509 6042
rect 536 6020 537 6036
rect 552 6020 565 6180
rect 595 6076 608 6180
rect 653 6158 654 6168
rect 669 6158 682 6168
rect 653 6154 682 6158
rect 687 6154 717 6180
rect 735 6166 751 6168
rect 823 6166 876 6180
rect 824 6164 888 6166
rect 931 6164 946 6180
rect 995 6177 1025 6180
rect 995 6174 1031 6177
rect 961 6166 977 6168
rect 735 6154 750 6158
rect 653 6152 750 6154
rect 778 6152 946 6164
rect 962 6154 977 6158
rect 995 6155 1034 6174
rect 1053 6168 1060 6169
rect 1059 6161 1060 6168
rect 1043 6158 1044 6161
rect 1059 6158 1072 6161
rect 995 6154 1025 6155
rect 1034 6154 1040 6155
rect 1043 6154 1072 6158
rect 962 6153 1072 6154
rect 962 6152 1078 6153
rect 637 6144 688 6152
rect 637 6132 662 6144
rect 669 6132 688 6144
rect 719 6144 769 6152
rect 719 6136 735 6144
rect 742 6142 769 6144
rect 778 6142 999 6152
rect 742 6132 999 6142
rect 1028 6144 1078 6152
rect 1028 6135 1044 6144
rect 637 6124 688 6132
rect 735 6124 999 6132
rect 1025 6132 1044 6135
rect 1051 6132 1078 6144
rect 1025 6124 1078 6132
rect 653 6116 654 6124
rect 669 6116 682 6124
rect 653 6108 669 6116
rect 650 6101 669 6104
rect 650 6092 672 6101
rect 623 6082 672 6092
rect 623 6076 653 6082
rect 672 6077 677 6082
rect 595 6060 669 6076
rect 687 6068 717 6124
rect 752 6114 960 6124
rect 995 6120 1040 6124
rect 1043 6123 1044 6124
rect 1059 6123 1072 6124
rect 778 6084 967 6114
rect 793 6081 967 6084
rect 786 6078 967 6081
rect 595 6058 608 6060
rect 623 6058 657 6060
rect 595 6042 669 6058
rect 696 6054 709 6068
rect 724 6054 740 6070
rect 786 6065 797 6078
rect 579 6020 580 6036
rect 595 6020 608 6042
rect 623 6020 653 6042
rect 696 6038 758 6054
rect 786 6047 797 6063
rect 802 6058 812 6078
rect 822 6058 836 6078
rect 839 6065 848 6078
rect 864 6065 873 6078
rect 802 6047 836 6058
rect 839 6047 848 6063
rect 864 6047 873 6063
rect 880 6058 890 6078
rect 900 6058 914 6078
rect 915 6065 926 6078
rect 880 6047 914 6058
rect 915 6047 926 6063
rect 972 6054 988 6070
rect 995 6068 1025 6120
rect 1059 6116 1060 6123
rect 1044 6108 1060 6116
rect 1031 6076 1044 6095
rect 1059 6076 1089 6092
rect 1031 6060 1105 6076
rect 1031 6058 1044 6060
rect 1059 6058 1093 6060
rect 696 6036 709 6038
rect 724 6036 758 6038
rect 696 6020 758 6036
rect 802 6031 818 6034
rect 880 6031 910 6042
rect 958 6038 1004 6054
rect 1031 6042 1105 6058
rect 958 6036 992 6038
rect 957 6020 1004 6036
rect 1031 6020 1044 6042
rect 1059 6020 1089 6042
rect 1116 6020 1117 6036
rect 1132 6020 1145 6180
rect 1175 6076 1188 6180
rect 1233 6158 1234 6168
rect 1249 6158 1262 6168
rect 1233 6154 1262 6158
rect 1267 6154 1297 6180
rect 1315 6166 1331 6168
rect 1403 6166 1456 6180
rect 1404 6164 1468 6166
rect 1511 6164 1526 6180
rect 1575 6177 1605 6180
rect 1575 6174 1611 6177
rect 1541 6166 1557 6168
rect 1315 6154 1330 6158
rect 1233 6152 1330 6154
rect 1358 6152 1526 6164
rect 1542 6154 1557 6158
rect 1575 6155 1614 6174
rect 1633 6168 1640 6169
rect 1639 6161 1640 6168
rect 1623 6158 1624 6161
rect 1639 6158 1652 6161
rect 1575 6154 1605 6155
rect 1614 6154 1620 6155
rect 1623 6154 1652 6158
rect 1542 6153 1652 6154
rect 1542 6152 1658 6153
rect 1217 6144 1268 6152
rect 1217 6132 1242 6144
rect 1249 6132 1268 6144
rect 1299 6144 1349 6152
rect 1299 6136 1315 6144
rect 1322 6142 1349 6144
rect 1358 6142 1579 6152
rect 1322 6132 1579 6142
rect 1608 6144 1658 6152
rect 1608 6135 1624 6144
rect 1217 6124 1268 6132
rect 1315 6124 1579 6132
rect 1605 6132 1624 6135
rect 1631 6132 1658 6144
rect 1605 6124 1658 6132
rect 1233 6116 1234 6124
rect 1249 6116 1262 6124
rect 1233 6108 1249 6116
rect 1230 6101 1249 6104
rect 1230 6092 1252 6101
rect 1203 6082 1252 6092
rect 1203 6076 1233 6082
rect 1252 6077 1257 6082
rect 1175 6060 1249 6076
rect 1267 6068 1297 6124
rect 1332 6114 1540 6124
rect 1575 6120 1620 6124
rect 1623 6123 1624 6124
rect 1639 6123 1652 6124
rect 1358 6084 1547 6114
rect 1373 6081 1547 6084
rect 1366 6078 1547 6081
rect 1175 6058 1188 6060
rect 1203 6058 1237 6060
rect 1175 6042 1249 6058
rect 1276 6054 1289 6068
rect 1304 6054 1320 6070
rect 1366 6065 1377 6078
rect 1159 6020 1160 6036
rect 1175 6020 1188 6042
rect 1203 6020 1233 6042
rect 1276 6038 1338 6054
rect 1366 6047 1377 6063
rect 1382 6058 1392 6078
rect 1402 6058 1416 6078
rect 1419 6065 1428 6078
rect 1444 6065 1453 6078
rect 1382 6047 1416 6058
rect 1419 6047 1428 6063
rect 1444 6047 1453 6063
rect 1460 6058 1470 6078
rect 1480 6058 1494 6078
rect 1495 6065 1506 6078
rect 1460 6047 1494 6058
rect 1495 6047 1506 6063
rect 1552 6054 1568 6070
rect 1575 6068 1605 6120
rect 1639 6116 1640 6123
rect 1624 6108 1640 6116
rect 1611 6076 1624 6095
rect 1639 6076 1669 6092
rect 1611 6060 1685 6076
rect 1611 6058 1624 6060
rect 1639 6058 1673 6060
rect 1276 6036 1289 6038
rect 1304 6036 1338 6038
rect 1276 6020 1338 6036
rect 1382 6031 1398 6034
rect 1460 6031 1490 6042
rect 1538 6038 1584 6054
rect 1611 6042 1685 6058
rect 1538 6036 1572 6038
rect 1537 6020 1584 6036
rect 1611 6020 1624 6042
rect 1639 6020 1669 6042
rect 1696 6020 1697 6036
rect 1712 6020 1725 6180
rect 1755 6076 1768 6180
rect 1813 6158 1814 6168
rect 1829 6158 1842 6168
rect 1813 6154 1842 6158
rect 1847 6154 1877 6180
rect 1895 6166 1911 6168
rect 1983 6166 2036 6180
rect 1984 6164 2048 6166
rect 2091 6164 2106 6180
rect 2155 6177 2185 6180
rect 2155 6174 2191 6177
rect 2121 6166 2137 6168
rect 1895 6154 1910 6158
rect 1813 6152 1910 6154
rect 1938 6152 2106 6164
rect 2122 6154 2137 6158
rect 2155 6155 2194 6174
rect 2213 6168 2220 6169
rect 2219 6161 2220 6168
rect 2203 6158 2204 6161
rect 2219 6158 2232 6161
rect 2155 6154 2185 6155
rect 2194 6154 2200 6155
rect 2203 6154 2232 6158
rect 2122 6153 2232 6154
rect 2122 6152 2238 6153
rect 1797 6144 1848 6152
rect 1797 6132 1822 6144
rect 1829 6132 1848 6144
rect 1879 6144 1929 6152
rect 1879 6136 1895 6144
rect 1902 6142 1929 6144
rect 1938 6142 2159 6152
rect 1902 6132 2159 6142
rect 2188 6144 2238 6152
rect 2188 6135 2204 6144
rect 1797 6124 1848 6132
rect 1895 6124 2159 6132
rect 2185 6132 2204 6135
rect 2211 6132 2238 6144
rect 2185 6124 2238 6132
rect 1813 6116 1814 6124
rect 1829 6116 1842 6124
rect 1813 6108 1829 6116
rect 1810 6101 1829 6104
rect 1810 6092 1832 6101
rect 1783 6082 1832 6092
rect 1783 6076 1813 6082
rect 1832 6077 1837 6082
rect 1755 6060 1829 6076
rect 1847 6068 1877 6124
rect 1912 6114 2120 6124
rect 2155 6120 2200 6124
rect 2203 6123 2204 6124
rect 2219 6123 2232 6124
rect 1938 6084 2127 6114
rect 1953 6081 2127 6084
rect 1946 6078 2127 6081
rect 1755 6058 1768 6060
rect 1783 6058 1817 6060
rect 1755 6042 1829 6058
rect 1856 6054 1869 6068
rect 1884 6054 1900 6070
rect 1946 6065 1957 6078
rect 1739 6020 1740 6036
rect 1755 6020 1768 6042
rect 1783 6020 1813 6042
rect 1856 6038 1918 6054
rect 1946 6047 1957 6063
rect 1962 6058 1972 6078
rect 1982 6058 1996 6078
rect 1999 6065 2008 6078
rect 2024 6065 2033 6078
rect 1962 6047 1996 6058
rect 1999 6047 2008 6063
rect 2024 6047 2033 6063
rect 2040 6058 2050 6078
rect 2060 6058 2074 6078
rect 2075 6065 2086 6078
rect 2040 6047 2074 6058
rect 2075 6047 2086 6063
rect 2132 6054 2148 6070
rect 2155 6068 2185 6120
rect 2219 6116 2220 6123
rect 2204 6108 2220 6116
rect 2191 6076 2204 6095
rect 2219 6076 2249 6092
rect 2191 6060 2265 6076
rect 2191 6058 2204 6060
rect 2219 6058 2253 6060
rect 1856 6036 1869 6038
rect 1884 6036 1918 6038
rect 1856 6020 1918 6036
rect 1962 6031 1976 6034
rect 2040 6031 2070 6042
rect 2118 6038 2164 6054
rect 2191 6042 2265 6058
rect 2118 6036 2152 6038
rect 2117 6020 2164 6036
rect 2191 6020 2204 6042
rect 2219 6020 2249 6042
rect 2276 6020 2277 6036
rect 2292 6020 2305 6180
rect 2335 6076 2348 6180
rect 2393 6158 2394 6168
rect 2409 6158 2422 6168
rect 2393 6154 2422 6158
rect 2427 6154 2457 6180
rect 2475 6166 2491 6168
rect 2563 6166 2616 6180
rect 2564 6164 2628 6166
rect 2671 6164 2686 6180
rect 2735 6177 2765 6180
rect 2735 6174 2771 6177
rect 2701 6166 2717 6168
rect 2475 6154 2490 6158
rect 2393 6152 2490 6154
rect 2518 6152 2686 6164
rect 2702 6154 2717 6158
rect 2735 6155 2774 6174
rect 2793 6168 2800 6169
rect 2799 6161 2800 6168
rect 2783 6158 2784 6161
rect 2799 6158 2812 6161
rect 2735 6154 2765 6155
rect 2774 6154 2780 6155
rect 2783 6154 2812 6158
rect 2702 6153 2812 6154
rect 2702 6152 2818 6153
rect 2377 6144 2428 6152
rect 2377 6132 2402 6144
rect 2409 6132 2428 6144
rect 2459 6144 2509 6152
rect 2459 6136 2475 6144
rect 2482 6142 2509 6144
rect 2518 6142 2739 6152
rect 2482 6132 2739 6142
rect 2768 6144 2818 6152
rect 2768 6135 2784 6144
rect 2377 6124 2428 6132
rect 2475 6124 2739 6132
rect 2765 6132 2784 6135
rect 2791 6132 2818 6144
rect 2765 6124 2818 6132
rect 2393 6116 2394 6124
rect 2409 6116 2422 6124
rect 2393 6108 2409 6116
rect 2390 6101 2409 6104
rect 2390 6092 2412 6101
rect 2363 6082 2412 6092
rect 2363 6076 2393 6082
rect 2412 6077 2417 6082
rect 2335 6060 2409 6076
rect 2427 6068 2457 6124
rect 2492 6114 2700 6124
rect 2735 6120 2780 6124
rect 2783 6123 2784 6124
rect 2799 6123 2812 6124
rect 2518 6084 2707 6114
rect 2533 6081 2707 6084
rect 2526 6078 2707 6081
rect 2335 6058 2348 6060
rect 2363 6058 2397 6060
rect 2335 6042 2409 6058
rect 2436 6054 2449 6068
rect 2464 6054 2480 6070
rect 2526 6065 2537 6078
rect 2319 6020 2320 6036
rect 2335 6020 2348 6042
rect 2363 6020 2393 6042
rect 2436 6038 2498 6054
rect 2526 6047 2537 6063
rect 2542 6058 2552 6078
rect 2562 6058 2576 6078
rect 2579 6065 2588 6078
rect 2604 6065 2613 6078
rect 2542 6047 2576 6058
rect 2579 6047 2588 6063
rect 2604 6047 2613 6063
rect 2620 6058 2630 6078
rect 2640 6058 2654 6078
rect 2655 6065 2666 6078
rect 2620 6047 2654 6058
rect 2655 6047 2666 6063
rect 2712 6054 2728 6070
rect 2735 6068 2765 6120
rect 2799 6116 2800 6123
rect 2784 6108 2800 6116
rect 2771 6076 2784 6095
rect 2799 6076 2829 6092
rect 2771 6060 2845 6076
rect 2771 6058 2784 6060
rect 2799 6058 2833 6060
rect 2436 6036 2449 6038
rect 2464 6036 2498 6038
rect 2436 6020 2498 6036
rect 2542 6031 2558 6034
rect 2620 6031 2650 6042
rect 2698 6038 2744 6054
rect 2771 6042 2845 6058
rect 2698 6036 2732 6038
rect 2697 6020 2744 6036
rect 2771 6020 2784 6042
rect 2799 6020 2829 6042
rect 2856 6020 2857 6036
rect 2872 6020 2885 6180
rect 2915 6076 2928 6180
rect 2973 6158 2974 6168
rect 2989 6158 3002 6168
rect 2973 6154 3002 6158
rect 3007 6154 3037 6180
rect 3055 6166 3071 6168
rect 3143 6166 3196 6180
rect 3144 6164 3208 6166
rect 3251 6164 3266 6180
rect 3315 6177 3345 6180
rect 3315 6174 3351 6177
rect 3281 6166 3297 6168
rect 3055 6154 3070 6158
rect 2973 6152 3070 6154
rect 3098 6152 3266 6164
rect 3282 6154 3297 6158
rect 3315 6155 3354 6174
rect 3373 6168 3380 6169
rect 3379 6161 3380 6168
rect 3363 6158 3364 6161
rect 3379 6158 3392 6161
rect 3315 6154 3345 6155
rect 3354 6154 3360 6155
rect 3363 6154 3392 6158
rect 3282 6153 3392 6154
rect 3282 6152 3398 6153
rect 2957 6144 3008 6152
rect 2957 6132 2982 6144
rect 2989 6132 3008 6144
rect 3039 6144 3089 6152
rect 3039 6136 3055 6144
rect 3062 6142 3089 6144
rect 3098 6142 3319 6152
rect 3062 6132 3319 6142
rect 3348 6144 3398 6152
rect 3348 6135 3364 6144
rect 2957 6124 3008 6132
rect 3055 6124 3319 6132
rect 3345 6132 3364 6135
rect 3371 6132 3398 6144
rect 3345 6124 3398 6132
rect 2973 6116 2974 6124
rect 2989 6116 3002 6124
rect 2973 6108 2989 6116
rect 2970 6101 2989 6104
rect 2970 6092 2992 6101
rect 2943 6082 2992 6092
rect 2943 6076 2973 6082
rect 2992 6077 2997 6082
rect 2915 6060 2989 6076
rect 3007 6068 3037 6124
rect 3072 6114 3280 6124
rect 3315 6120 3360 6124
rect 3363 6123 3364 6124
rect 3379 6123 3392 6124
rect 3098 6084 3287 6114
rect 3113 6081 3287 6084
rect 3106 6078 3287 6081
rect 2915 6058 2928 6060
rect 2943 6058 2977 6060
rect 2915 6042 2989 6058
rect 3016 6054 3029 6068
rect 3044 6054 3060 6070
rect 3106 6065 3117 6078
rect 2899 6020 2900 6036
rect 2915 6020 2928 6042
rect 2943 6020 2973 6042
rect 3016 6038 3078 6054
rect 3106 6047 3117 6063
rect 3122 6058 3132 6078
rect 3142 6058 3156 6078
rect 3159 6065 3168 6078
rect 3184 6065 3193 6078
rect 3122 6047 3156 6058
rect 3159 6047 3168 6063
rect 3184 6047 3193 6063
rect 3200 6058 3210 6078
rect 3220 6058 3234 6078
rect 3235 6065 3246 6078
rect 3200 6047 3234 6058
rect 3235 6047 3246 6063
rect 3292 6054 3308 6070
rect 3315 6068 3345 6120
rect 3379 6116 3380 6123
rect 3364 6108 3380 6116
rect 3351 6076 3364 6095
rect 3379 6076 3409 6092
rect 3351 6060 3425 6076
rect 3351 6058 3364 6060
rect 3379 6058 3413 6060
rect 3016 6036 3029 6038
rect 3044 6036 3078 6038
rect 3016 6020 3078 6036
rect 3122 6031 3138 6034
rect 3200 6031 3230 6042
rect 3278 6038 3324 6054
rect 3351 6042 3425 6058
rect 3278 6036 3312 6038
rect 3277 6020 3324 6036
rect 3351 6020 3364 6042
rect 3379 6020 3409 6042
rect 3436 6020 3437 6036
rect 3452 6020 3465 6180
rect 3495 6076 3508 6180
rect 3553 6158 3554 6168
rect 3569 6158 3582 6168
rect 3553 6154 3582 6158
rect 3587 6154 3617 6180
rect 3635 6166 3651 6168
rect 3723 6166 3776 6180
rect 3724 6164 3788 6166
rect 3831 6164 3846 6180
rect 3895 6177 3925 6180
rect 3895 6174 3931 6177
rect 3861 6166 3877 6168
rect 3635 6154 3650 6158
rect 3553 6152 3650 6154
rect 3678 6152 3846 6164
rect 3862 6154 3877 6158
rect 3895 6155 3934 6174
rect 3953 6168 3960 6169
rect 3959 6161 3960 6168
rect 3943 6158 3944 6161
rect 3959 6158 3972 6161
rect 3895 6154 3925 6155
rect 3934 6154 3940 6155
rect 3943 6154 3972 6158
rect 3862 6153 3972 6154
rect 3862 6152 3978 6153
rect 3537 6144 3588 6152
rect 3537 6132 3562 6144
rect 3569 6132 3588 6144
rect 3619 6144 3669 6152
rect 3619 6136 3635 6144
rect 3642 6142 3669 6144
rect 3678 6142 3899 6152
rect 3642 6132 3899 6142
rect 3928 6144 3978 6152
rect 3928 6135 3944 6144
rect 3537 6124 3588 6132
rect 3635 6124 3899 6132
rect 3925 6132 3944 6135
rect 3951 6132 3978 6144
rect 3925 6124 3978 6132
rect 3553 6116 3554 6124
rect 3569 6116 3582 6124
rect 3553 6108 3569 6116
rect 3550 6101 3569 6104
rect 3550 6092 3572 6101
rect 3523 6082 3572 6092
rect 3523 6076 3553 6082
rect 3572 6077 3577 6082
rect 3495 6060 3569 6076
rect 3587 6068 3617 6124
rect 3652 6114 3860 6124
rect 3895 6120 3940 6124
rect 3943 6123 3944 6124
rect 3959 6123 3972 6124
rect 3678 6084 3867 6114
rect 3693 6081 3867 6084
rect 3686 6078 3867 6081
rect 3495 6058 3508 6060
rect 3523 6058 3557 6060
rect 3495 6042 3569 6058
rect 3596 6054 3609 6068
rect 3624 6054 3640 6070
rect 3686 6065 3697 6078
rect 3479 6020 3480 6036
rect 3495 6020 3508 6042
rect 3523 6020 3553 6042
rect 3596 6038 3658 6054
rect 3686 6047 3697 6063
rect 3702 6058 3712 6078
rect 3722 6058 3736 6078
rect 3739 6065 3748 6078
rect 3764 6065 3773 6078
rect 3702 6047 3736 6058
rect 3739 6047 3748 6063
rect 3764 6047 3773 6063
rect 3780 6058 3790 6078
rect 3800 6058 3814 6078
rect 3815 6065 3826 6078
rect 3780 6047 3814 6058
rect 3815 6047 3826 6063
rect 3872 6054 3888 6070
rect 3895 6068 3925 6120
rect 3959 6116 3960 6123
rect 3944 6108 3960 6116
rect 3931 6076 3944 6095
rect 3959 6076 3989 6092
rect 3931 6060 4005 6076
rect 3931 6058 3944 6060
rect 3959 6058 3993 6060
rect 3596 6036 3609 6038
rect 3624 6036 3658 6038
rect 3596 6020 3658 6036
rect 3702 6031 3718 6034
rect 3780 6031 3810 6042
rect 3858 6038 3904 6054
rect 3931 6042 4005 6058
rect 3858 6036 3892 6038
rect 3857 6020 3904 6036
rect 3931 6020 3944 6042
rect 3959 6020 3989 6042
rect 4016 6020 4017 6036
rect 4032 6020 4045 6180
rect 4075 6076 4088 6180
rect 4133 6158 4134 6168
rect 4149 6158 4162 6168
rect 4133 6154 4162 6158
rect 4167 6154 4197 6180
rect 4215 6166 4231 6168
rect 4303 6166 4356 6180
rect 4304 6164 4368 6166
rect 4411 6164 4426 6180
rect 4475 6177 4505 6180
rect 4475 6174 4511 6177
rect 4441 6166 4457 6168
rect 4215 6154 4230 6158
rect 4133 6152 4230 6154
rect 4258 6152 4426 6164
rect 4442 6154 4457 6158
rect 4475 6155 4514 6174
rect 4533 6168 4540 6169
rect 4539 6161 4540 6168
rect 4523 6158 4524 6161
rect 4539 6158 4552 6161
rect 4475 6154 4505 6155
rect 4514 6154 4520 6155
rect 4523 6154 4552 6158
rect 4442 6153 4552 6154
rect 4442 6152 4558 6153
rect 4117 6144 4168 6152
rect 4117 6132 4142 6144
rect 4149 6132 4168 6144
rect 4199 6144 4249 6152
rect 4199 6136 4215 6144
rect 4222 6142 4249 6144
rect 4258 6142 4479 6152
rect 4222 6132 4479 6142
rect 4508 6144 4558 6152
rect 4508 6135 4524 6144
rect 4117 6124 4168 6132
rect 4215 6124 4479 6132
rect 4505 6132 4524 6135
rect 4531 6132 4558 6144
rect 4505 6124 4558 6132
rect 4133 6116 4134 6124
rect 4149 6116 4162 6124
rect 4133 6108 4149 6116
rect 4130 6101 4149 6104
rect 4130 6092 4152 6101
rect 4103 6082 4152 6092
rect 4103 6076 4133 6082
rect 4152 6077 4157 6082
rect 4075 6060 4149 6076
rect 4167 6068 4197 6124
rect 4232 6114 4440 6124
rect 4475 6120 4520 6124
rect 4523 6123 4524 6124
rect 4539 6123 4552 6124
rect 4258 6084 4447 6114
rect 4273 6081 4447 6084
rect 4266 6078 4447 6081
rect 4075 6058 4088 6060
rect 4103 6058 4137 6060
rect 4075 6042 4149 6058
rect 4176 6054 4189 6068
rect 4204 6054 4220 6070
rect 4266 6065 4277 6078
rect 4059 6020 4060 6036
rect 4075 6020 4088 6042
rect 4103 6020 4133 6042
rect 4176 6038 4238 6054
rect 4266 6047 4277 6063
rect 4282 6058 4292 6078
rect 4302 6058 4316 6078
rect 4319 6065 4328 6078
rect 4344 6065 4353 6078
rect 4282 6047 4316 6058
rect 4319 6047 4328 6063
rect 4344 6047 4353 6063
rect 4360 6058 4370 6078
rect 4380 6058 4394 6078
rect 4395 6065 4406 6078
rect 4360 6047 4394 6058
rect 4395 6047 4406 6063
rect 4452 6054 4468 6070
rect 4475 6068 4505 6120
rect 4539 6116 4540 6123
rect 4524 6108 4540 6116
rect 4511 6076 4524 6095
rect 4539 6076 4569 6092
rect 4511 6060 4585 6076
rect 4511 6058 4524 6060
rect 4539 6058 4573 6060
rect 4176 6036 4189 6038
rect 4204 6036 4238 6038
rect 4176 6020 4238 6036
rect 4282 6031 4298 6034
rect 4360 6031 4390 6042
rect 4438 6038 4484 6054
rect 4511 6042 4585 6058
rect 4438 6036 4472 6038
rect 4437 6020 4484 6036
rect 4511 6020 4524 6042
rect 4539 6020 4569 6042
rect 4596 6020 4597 6036
rect 4612 6020 4625 6180
rect 4655 6076 4668 6180
rect 4713 6158 4714 6168
rect 4729 6158 4742 6168
rect 4713 6154 4742 6158
rect 4747 6154 4777 6180
rect 4795 6166 4811 6168
rect 4883 6166 4936 6180
rect 4884 6164 4948 6166
rect 4991 6164 5006 6180
rect 5055 6177 5085 6180
rect 5055 6174 5091 6177
rect 5021 6166 5037 6168
rect 4795 6154 4810 6158
rect 4713 6152 4810 6154
rect 4838 6152 5006 6164
rect 5022 6154 5037 6158
rect 5055 6155 5094 6174
rect 5113 6168 5120 6169
rect 5119 6161 5120 6168
rect 5103 6158 5104 6161
rect 5119 6158 5132 6161
rect 5055 6154 5085 6155
rect 5094 6154 5100 6155
rect 5103 6154 5132 6158
rect 5022 6153 5132 6154
rect 5022 6152 5138 6153
rect 4697 6144 4748 6152
rect 4697 6132 4722 6144
rect 4729 6132 4748 6144
rect 4779 6144 4829 6152
rect 4779 6136 4795 6144
rect 4802 6142 4829 6144
rect 4838 6142 5059 6152
rect 4802 6132 5059 6142
rect 5088 6144 5138 6152
rect 5088 6135 5104 6144
rect 4697 6124 4748 6132
rect 4795 6124 5059 6132
rect 5085 6132 5104 6135
rect 5111 6132 5138 6144
rect 5085 6124 5138 6132
rect 4713 6116 4714 6124
rect 4729 6116 4742 6124
rect 4713 6108 4729 6116
rect 4710 6101 4729 6104
rect 4710 6092 4732 6101
rect 4683 6082 4732 6092
rect 4683 6076 4713 6082
rect 4732 6077 4737 6082
rect 4655 6060 4729 6076
rect 4747 6068 4777 6124
rect 4812 6114 5020 6124
rect 5055 6120 5100 6124
rect 5103 6123 5104 6124
rect 5119 6123 5132 6124
rect 4838 6084 5027 6114
rect 4853 6081 5027 6084
rect 4846 6078 5027 6081
rect 4655 6058 4668 6060
rect 4683 6058 4717 6060
rect 4655 6042 4729 6058
rect 4756 6054 4769 6068
rect 4784 6054 4800 6070
rect 4846 6065 4857 6078
rect 4639 6020 4640 6036
rect 4655 6020 4668 6042
rect 4683 6020 4713 6042
rect 4756 6038 4818 6054
rect 4846 6047 4857 6063
rect 4862 6058 4872 6078
rect 4882 6058 4896 6078
rect 4899 6065 4908 6078
rect 4924 6065 4933 6078
rect 4862 6047 4896 6058
rect 4899 6047 4908 6063
rect 4924 6047 4933 6063
rect 4940 6058 4950 6078
rect 4960 6058 4974 6078
rect 4975 6065 4986 6078
rect 4940 6047 4974 6058
rect 4975 6047 4986 6063
rect 5032 6054 5048 6070
rect 5055 6068 5085 6120
rect 5119 6116 5120 6123
rect 5104 6108 5120 6116
rect 5091 6076 5104 6095
rect 5119 6076 5149 6092
rect 5091 6060 5165 6076
rect 5091 6058 5104 6060
rect 5119 6058 5153 6060
rect 4756 6036 4769 6038
rect 4784 6036 4818 6038
rect 4756 6020 4818 6036
rect 4862 6031 4878 6034
rect 4940 6031 4970 6042
rect 5018 6038 5064 6054
rect 5091 6042 5165 6058
rect 5018 6036 5052 6038
rect 5017 6020 5064 6036
rect 5091 6020 5104 6042
rect 5119 6020 5149 6042
rect 5176 6020 5177 6036
rect 5192 6020 5205 6180
rect 5235 6076 5248 6180
rect 5293 6158 5294 6168
rect 5309 6158 5322 6168
rect 5293 6154 5322 6158
rect 5327 6154 5357 6180
rect 5375 6166 5391 6168
rect 5463 6166 5516 6180
rect 5464 6164 5528 6166
rect 5571 6164 5586 6180
rect 5635 6177 5665 6180
rect 5635 6174 5671 6177
rect 5601 6166 5617 6168
rect 5375 6154 5390 6158
rect 5293 6152 5390 6154
rect 5418 6152 5586 6164
rect 5602 6154 5617 6158
rect 5635 6155 5674 6174
rect 5693 6168 5700 6169
rect 5699 6161 5700 6168
rect 5683 6158 5684 6161
rect 5699 6158 5712 6161
rect 5635 6154 5665 6155
rect 5674 6154 5680 6155
rect 5683 6154 5712 6158
rect 5602 6153 5712 6154
rect 5602 6152 5718 6153
rect 5277 6144 5328 6152
rect 5277 6132 5302 6144
rect 5309 6132 5328 6144
rect 5359 6144 5409 6152
rect 5359 6136 5375 6144
rect 5382 6142 5409 6144
rect 5418 6142 5639 6152
rect 5382 6132 5639 6142
rect 5668 6144 5718 6152
rect 5668 6135 5684 6144
rect 5277 6124 5328 6132
rect 5375 6124 5639 6132
rect 5665 6132 5684 6135
rect 5691 6132 5718 6144
rect 5665 6124 5718 6132
rect 5293 6116 5294 6124
rect 5309 6116 5322 6124
rect 5293 6108 5309 6116
rect 5290 6101 5309 6104
rect 5290 6092 5312 6101
rect 5263 6082 5312 6092
rect 5263 6076 5293 6082
rect 5312 6077 5317 6082
rect 5235 6060 5309 6076
rect 5327 6068 5357 6124
rect 5392 6114 5600 6124
rect 5635 6120 5680 6124
rect 5683 6123 5684 6124
rect 5699 6123 5712 6124
rect 5418 6084 5607 6114
rect 5433 6081 5607 6084
rect 5426 6078 5607 6081
rect 5235 6058 5248 6060
rect 5263 6058 5297 6060
rect 5235 6042 5309 6058
rect 5336 6054 5349 6068
rect 5364 6054 5380 6070
rect 5426 6065 5437 6078
rect 5219 6020 5220 6036
rect 5235 6020 5248 6042
rect 5263 6020 5293 6042
rect 5336 6038 5398 6054
rect 5426 6047 5437 6063
rect 5442 6058 5452 6078
rect 5462 6058 5476 6078
rect 5479 6065 5488 6078
rect 5504 6065 5513 6078
rect 5442 6047 5476 6058
rect 5479 6047 5488 6063
rect 5504 6047 5513 6063
rect 5520 6058 5530 6078
rect 5540 6058 5554 6078
rect 5555 6065 5566 6078
rect 5520 6047 5554 6058
rect 5555 6047 5566 6063
rect 5612 6054 5628 6070
rect 5635 6068 5665 6120
rect 5699 6116 5700 6123
rect 5684 6108 5700 6116
rect 5671 6076 5684 6095
rect 5699 6076 5729 6092
rect 5671 6060 5745 6076
rect 5671 6058 5684 6060
rect 5699 6058 5733 6060
rect 5336 6036 5349 6038
rect 5364 6036 5398 6038
rect 5336 6020 5398 6036
rect 5442 6031 5458 6034
rect 5520 6031 5550 6042
rect 5598 6038 5644 6054
rect 5671 6042 5745 6058
rect 5598 6036 5632 6038
rect 5597 6020 5644 6036
rect 5671 6020 5684 6042
rect 5699 6020 5729 6042
rect 5756 6020 5757 6036
rect 5772 6020 5785 6180
rect 5815 6076 5828 6180
rect 5873 6158 5874 6168
rect 5889 6158 5902 6168
rect 5873 6154 5902 6158
rect 5907 6154 5937 6180
rect 5955 6166 5971 6168
rect 6043 6166 6096 6180
rect 6044 6164 6108 6166
rect 6151 6164 6166 6180
rect 6215 6177 6245 6180
rect 6215 6174 6251 6177
rect 6181 6166 6197 6168
rect 5955 6154 5970 6158
rect 5873 6152 5970 6154
rect 5998 6152 6166 6164
rect 6182 6154 6197 6158
rect 6215 6155 6254 6174
rect 6273 6168 6280 6169
rect 6279 6161 6280 6168
rect 6263 6158 6264 6161
rect 6279 6158 6292 6161
rect 6215 6154 6245 6155
rect 6254 6154 6260 6155
rect 6263 6154 6292 6158
rect 6182 6153 6292 6154
rect 6182 6152 6298 6153
rect 5857 6144 5908 6152
rect 5857 6132 5882 6144
rect 5889 6132 5908 6144
rect 5939 6144 5989 6152
rect 5939 6136 5955 6144
rect 5962 6142 5989 6144
rect 5998 6142 6219 6152
rect 5962 6132 6219 6142
rect 6248 6144 6298 6152
rect 6248 6135 6264 6144
rect 5857 6124 5908 6132
rect 5955 6124 6219 6132
rect 6245 6132 6264 6135
rect 6271 6132 6298 6144
rect 6245 6124 6298 6132
rect 5873 6116 5874 6124
rect 5889 6116 5902 6124
rect 5873 6108 5889 6116
rect 5870 6101 5889 6104
rect 5870 6092 5892 6101
rect 5843 6082 5892 6092
rect 5843 6076 5873 6082
rect 5892 6077 5897 6082
rect 5815 6060 5889 6076
rect 5907 6068 5937 6124
rect 5972 6114 6180 6124
rect 6215 6120 6260 6124
rect 6263 6123 6264 6124
rect 6279 6123 6292 6124
rect 5998 6084 6187 6114
rect 6013 6081 6187 6084
rect 6006 6078 6187 6081
rect 5815 6058 5828 6060
rect 5843 6058 5877 6060
rect 5815 6042 5889 6058
rect 5916 6054 5929 6068
rect 5944 6054 5960 6070
rect 6006 6065 6017 6078
rect 5799 6020 5800 6036
rect 5815 6020 5828 6042
rect 5843 6020 5873 6042
rect 5916 6038 5978 6054
rect 6006 6047 6017 6063
rect 6022 6058 6032 6078
rect 6042 6058 6056 6078
rect 6059 6065 6068 6078
rect 6084 6065 6093 6078
rect 6022 6047 6056 6058
rect 6059 6047 6068 6063
rect 6084 6047 6093 6063
rect 6100 6058 6110 6078
rect 6120 6058 6134 6078
rect 6135 6065 6146 6078
rect 6100 6047 6134 6058
rect 6135 6047 6146 6063
rect 6192 6054 6208 6070
rect 6215 6068 6245 6120
rect 6279 6116 6280 6123
rect 6264 6108 6280 6116
rect 6251 6076 6264 6095
rect 6279 6076 6309 6092
rect 6251 6060 6325 6076
rect 6251 6058 6264 6060
rect 6279 6058 6313 6060
rect 5916 6036 5929 6038
rect 5944 6036 5978 6038
rect 5916 6020 5978 6036
rect 6022 6031 6038 6034
rect 6100 6031 6130 6042
rect 6178 6038 6224 6054
rect 6251 6042 6325 6058
rect 6178 6036 6212 6038
rect 6177 6020 6224 6036
rect 6251 6020 6264 6042
rect 6279 6020 6309 6042
rect 6336 6020 6337 6036
rect 6352 6020 6365 6180
rect 6395 6076 6408 6180
rect 6453 6158 6454 6168
rect 6469 6158 6482 6168
rect 6453 6154 6482 6158
rect 6487 6154 6517 6180
rect 6535 6166 6551 6168
rect 6623 6166 6676 6180
rect 6624 6164 6688 6166
rect 6731 6164 6746 6180
rect 6795 6177 6825 6180
rect 6795 6174 6831 6177
rect 6761 6166 6777 6168
rect 6535 6154 6550 6158
rect 6453 6152 6550 6154
rect 6578 6152 6746 6164
rect 6762 6154 6777 6158
rect 6795 6155 6834 6174
rect 6853 6168 6860 6169
rect 6859 6161 6860 6168
rect 6843 6158 6844 6161
rect 6859 6158 6872 6161
rect 6795 6154 6825 6155
rect 6834 6154 6840 6155
rect 6843 6154 6872 6158
rect 6762 6153 6872 6154
rect 6762 6152 6878 6153
rect 6437 6144 6488 6152
rect 6437 6132 6462 6144
rect 6469 6132 6488 6144
rect 6519 6144 6569 6152
rect 6519 6136 6535 6144
rect 6542 6142 6569 6144
rect 6578 6142 6799 6152
rect 6542 6132 6799 6142
rect 6828 6144 6878 6152
rect 6828 6135 6844 6144
rect 6437 6124 6488 6132
rect 6535 6124 6799 6132
rect 6825 6132 6844 6135
rect 6851 6132 6878 6144
rect 6825 6124 6878 6132
rect 6453 6116 6454 6124
rect 6469 6116 6482 6124
rect 6453 6108 6469 6116
rect 6450 6101 6469 6104
rect 6450 6092 6472 6101
rect 6423 6082 6472 6092
rect 6423 6076 6453 6082
rect 6472 6077 6477 6082
rect 6395 6060 6469 6076
rect 6487 6068 6517 6124
rect 6552 6114 6760 6124
rect 6795 6120 6840 6124
rect 6843 6123 6844 6124
rect 6859 6123 6872 6124
rect 6578 6084 6767 6114
rect 6593 6081 6767 6084
rect 6586 6078 6767 6081
rect 6395 6058 6408 6060
rect 6423 6058 6457 6060
rect 6395 6042 6469 6058
rect 6496 6054 6509 6068
rect 6524 6054 6540 6070
rect 6586 6065 6597 6078
rect 6379 6020 6380 6036
rect 6395 6020 6408 6042
rect 6423 6020 6453 6042
rect 6496 6038 6558 6054
rect 6586 6047 6597 6063
rect 6602 6058 6612 6078
rect 6622 6058 6636 6078
rect 6639 6065 6648 6078
rect 6664 6065 6673 6078
rect 6602 6047 6636 6058
rect 6639 6047 6648 6063
rect 6664 6047 6673 6063
rect 6680 6058 6690 6078
rect 6700 6058 6714 6078
rect 6715 6065 6726 6078
rect 6680 6047 6714 6058
rect 6715 6047 6726 6063
rect 6772 6054 6788 6070
rect 6795 6068 6825 6120
rect 6859 6116 6860 6123
rect 6844 6108 6860 6116
rect 6831 6076 6844 6095
rect 6859 6076 6889 6092
rect 6831 6060 6905 6076
rect 6831 6058 6844 6060
rect 6859 6058 6893 6060
rect 6496 6036 6509 6038
rect 6524 6036 6558 6038
rect 6496 6020 6558 6036
rect 6602 6031 6618 6034
rect 6680 6031 6710 6042
rect 6758 6038 6804 6054
rect 6831 6042 6905 6058
rect 6758 6036 6792 6038
rect 6757 6020 6804 6036
rect 6831 6020 6844 6042
rect 6859 6020 6889 6042
rect 6916 6020 6917 6036
rect 6932 6020 6945 6180
rect 6975 6076 6988 6180
rect 7033 6158 7034 6168
rect 7049 6158 7062 6168
rect 7033 6154 7062 6158
rect 7067 6154 7097 6180
rect 7115 6166 7131 6168
rect 7203 6166 7256 6180
rect 7204 6164 7268 6166
rect 7311 6164 7326 6180
rect 7375 6177 7405 6180
rect 7375 6174 7411 6177
rect 7341 6166 7357 6168
rect 7115 6154 7130 6158
rect 7033 6152 7130 6154
rect 7158 6152 7326 6164
rect 7342 6154 7357 6158
rect 7375 6155 7414 6174
rect 7433 6168 7440 6169
rect 7439 6161 7440 6168
rect 7423 6158 7424 6161
rect 7439 6158 7452 6161
rect 7375 6154 7405 6155
rect 7414 6154 7420 6155
rect 7423 6154 7452 6158
rect 7342 6153 7452 6154
rect 7342 6152 7458 6153
rect 7017 6144 7068 6152
rect 7017 6132 7042 6144
rect 7049 6132 7068 6144
rect 7099 6144 7149 6152
rect 7099 6136 7115 6144
rect 7122 6142 7149 6144
rect 7158 6142 7379 6152
rect 7122 6132 7379 6142
rect 7408 6144 7458 6152
rect 7408 6135 7424 6144
rect 7017 6124 7068 6132
rect 7115 6124 7379 6132
rect 7405 6132 7424 6135
rect 7431 6132 7458 6144
rect 7405 6124 7458 6132
rect 7033 6116 7034 6124
rect 7049 6116 7062 6124
rect 7033 6108 7049 6116
rect 7030 6101 7049 6104
rect 7030 6092 7052 6101
rect 7003 6082 7052 6092
rect 7003 6076 7033 6082
rect 7052 6077 7057 6082
rect 6975 6060 7049 6076
rect 7067 6068 7097 6124
rect 7132 6114 7340 6124
rect 7375 6120 7420 6124
rect 7423 6123 7424 6124
rect 7439 6123 7452 6124
rect 7158 6084 7347 6114
rect 7173 6081 7347 6084
rect 7166 6078 7347 6081
rect 6975 6058 6988 6060
rect 7003 6058 7037 6060
rect 6975 6042 7049 6058
rect 7076 6054 7089 6068
rect 7104 6054 7120 6070
rect 7166 6065 7177 6078
rect 6959 6020 6960 6036
rect 6975 6020 6988 6042
rect 7003 6020 7033 6042
rect 7076 6038 7138 6054
rect 7166 6047 7177 6063
rect 7182 6058 7192 6078
rect 7202 6058 7216 6078
rect 7219 6065 7228 6078
rect 7244 6065 7253 6078
rect 7182 6047 7216 6058
rect 7219 6047 7228 6063
rect 7244 6047 7253 6063
rect 7260 6058 7270 6078
rect 7280 6058 7294 6078
rect 7295 6065 7306 6078
rect 7260 6047 7294 6058
rect 7295 6047 7306 6063
rect 7352 6054 7368 6070
rect 7375 6068 7405 6120
rect 7439 6116 7440 6123
rect 7424 6108 7440 6116
rect 7411 6076 7424 6095
rect 7439 6076 7469 6092
rect 7411 6060 7485 6076
rect 7411 6058 7424 6060
rect 7439 6058 7473 6060
rect 7076 6036 7089 6038
rect 7104 6036 7138 6038
rect 7076 6020 7138 6036
rect 7182 6031 7198 6034
rect 7260 6031 7290 6042
rect 7338 6038 7384 6054
rect 7411 6042 7485 6058
rect 7338 6036 7372 6038
rect 7337 6020 7384 6036
rect 7411 6020 7424 6042
rect 7439 6020 7469 6042
rect 7496 6020 7497 6036
rect 7512 6020 7525 6180
rect 7555 6076 7568 6180
rect 7613 6158 7614 6168
rect 7629 6158 7642 6168
rect 7613 6154 7642 6158
rect 7647 6154 7677 6180
rect 7695 6166 7711 6168
rect 7783 6166 7836 6180
rect 7784 6164 7848 6166
rect 7891 6164 7906 6180
rect 7955 6177 7985 6180
rect 7955 6174 7991 6177
rect 7921 6166 7937 6168
rect 7695 6154 7710 6158
rect 7613 6152 7710 6154
rect 7738 6152 7906 6164
rect 7922 6154 7937 6158
rect 7955 6155 7994 6174
rect 8013 6168 8020 6169
rect 8019 6161 8020 6168
rect 8003 6158 8004 6161
rect 8019 6158 8032 6161
rect 7955 6154 7985 6155
rect 7994 6154 8000 6155
rect 8003 6154 8032 6158
rect 7922 6153 8032 6154
rect 7922 6152 8038 6153
rect 7597 6144 7648 6152
rect 7597 6132 7622 6144
rect 7629 6132 7648 6144
rect 7679 6144 7729 6152
rect 7679 6136 7695 6144
rect 7702 6142 7729 6144
rect 7738 6142 7959 6152
rect 7702 6132 7959 6142
rect 7988 6144 8038 6152
rect 7988 6135 8004 6144
rect 7597 6124 7648 6132
rect 7695 6124 7959 6132
rect 7985 6132 8004 6135
rect 8011 6132 8038 6144
rect 7985 6124 8038 6132
rect 7613 6116 7614 6124
rect 7629 6116 7642 6124
rect 7613 6108 7629 6116
rect 7610 6101 7629 6104
rect 7610 6092 7632 6101
rect 7583 6082 7632 6092
rect 7583 6076 7613 6082
rect 7632 6077 7637 6082
rect 7555 6060 7629 6076
rect 7647 6068 7677 6124
rect 7712 6114 7920 6124
rect 7955 6120 8000 6124
rect 8003 6123 8004 6124
rect 8019 6123 8032 6124
rect 7738 6084 7927 6114
rect 7753 6081 7927 6084
rect 7746 6078 7927 6081
rect 7555 6058 7568 6060
rect 7583 6058 7617 6060
rect 7555 6042 7629 6058
rect 7656 6054 7669 6068
rect 7684 6054 7700 6070
rect 7746 6065 7757 6078
rect 7539 6020 7540 6036
rect 7555 6020 7568 6042
rect 7583 6020 7613 6042
rect 7656 6038 7718 6054
rect 7746 6047 7757 6063
rect 7762 6058 7772 6078
rect 7782 6058 7796 6078
rect 7799 6065 7808 6078
rect 7824 6065 7833 6078
rect 7762 6047 7796 6058
rect 7799 6047 7808 6063
rect 7824 6047 7833 6063
rect 7840 6058 7850 6078
rect 7860 6058 7874 6078
rect 7875 6065 7886 6078
rect 7840 6047 7874 6058
rect 7875 6047 7886 6063
rect 7932 6054 7948 6070
rect 7955 6068 7985 6120
rect 8019 6116 8020 6123
rect 8004 6108 8020 6116
rect 7991 6076 8004 6095
rect 8019 6076 8049 6092
rect 7991 6060 8065 6076
rect 7991 6058 8004 6060
rect 8019 6058 8053 6060
rect 7656 6036 7669 6038
rect 7684 6036 7718 6038
rect 7656 6020 7718 6036
rect 7762 6031 7778 6034
rect 7840 6031 7870 6042
rect 7918 6038 7964 6054
rect 7991 6042 8065 6058
rect 7918 6036 7952 6038
rect 7917 6020 7964 6036
rect 7991 6020 8004 6042
rect 8019 6020 8049 6042
rect 8076 6020 8077 6036
rect 8092 6020 8105 6180
rect 8135 6076 8148 6180
rect 8193 6158 8194 6168
rect 8209 6158 8222 6168
rect 8193 6154 8222 6158
rect 8227 6154 8257 6180
rect 8275 6166 8291 6168
rect 8363 6166 8416 6180
rect 8364 6164 8428 6166
rect 8471 6164 8486 6180
rect 8535 6177 8565 6180
rect 8535 6174 8571 6177
rect 8501 6166 8517 6168
rect 8275 6154 8290 6158
rect 8193 6152 8290 6154
rect 8318 6152 8486 6164
rect 8502 6154 8517 6158
rect 8535 6155 8574 6174
rect 8593 6168 8600 6169
rect 8599 6161 8600 6168
rect 8583 6158 8584 6161
rect 8599 6158 8612 6161
rect 8535 6154 8565 6155
rect 8574 6154 8580 6155
rect 8583 6154 8612 6158
rect 8502 6153 8612 6154
rect 8502 6152 8618 6153
rect 8177 6144 8228 6152
rect 8177 6132 8202 6144
rect 8209 6132 8228 6144
rect 8259 6144 8309 6152
rect 8259 6136 8275 6144
rect 8282 6142 8309 6144
rect 8318 6142 8539 6152
rect 8282 6132 8539 6142
rect 8568 6144 8618 6152
rect 8568 6135 8584 6144
rect 8177 6124 8228 6132
rect 8275 6124 8539 6132
rect 8565 6132 8584 6135
rect 8591 6132 8618 6144
rect 8565 6124 8618 6132
rect 8193 6116 8194 6124
rect 8209 6116 8222 6124
rect 8193 6108 8209 6116
rect 8190 6101 8209 6104
rect 8190 6092 8212 6101
rect 8163 6082 8212 6092
rect 8163 6076 8193 6082
rect 8212 6077 8217 6082
rect 8135 6060 8209 6076
rect 8227 6068 8257 6124
rect 8292 6114 8500 6124
rect 8535 6120 8580 6124
rect 8583 6123 8584 6124
rect 8599 6123 8612 6124
rect 8318 6084 8507 6114
rect 8333 6081 8507 6084
rect 8326 6078 8507 6081
rect 8135 6058 8148 6060
rect 8163 6058 8197 6060
rect 8135 6042 8209 6058
rect 8236 6054 8249 6068
rect 8264 6054 8280 6070
rect 8326 6065 8337 6078
rect 8119 6020 8120 6036
rect 8135 6020 8148 6042
rect 8163 6020 8193 6042
rect 8236 6038 8298 6054
rect 8326 6047 8337 6063
rect 8342 6058 8352 6078
rect 8362 6058 8376 6078
rect 8379 6065 8388 6078
rect 8404 6065 8413 6078
rect 8342 6047 8376 6058
rect 8379 6047 8388 6063
rect 8404 6047 8413 6063
rect 8420 6058 8430 6078
rect 8440 6058 8454 6078
rect 8455 6065 8466 6078
rect 8420 6047 8454 6058
rect 8455 6047 8466 6063
rect 8512 6054 8528 6070
rect 8535 6068 8565 6120
rect 8599 6116 8600 6123
rect 8584 6108 8600 6116
rect 8571 6076 8584 6095
rect 8599 6076 8629 6092
rect 8571 6060 8645 6076
rect 8571 6058 8584 6060
rect 8599 6058 8633 6060
rect 8236 6036 8249 6038
rect 8264 6036 8298 6038
rect 8236 6020 8298 6036
rect 8342 6031 8358 6034
rect 8420 6031 8450 6042
rect 8498 6038 8544 6054
rect 8571 6042 8645 6058
rect 8498 6036 8532 6038
rect 8497 6020 8544 6036
rect 8571 6020 8584 6042
rect 8599 6020 8629 6042
rect 8656 6020 8657 6036
rect 8672 6020 8685 6180
rect 8715 6076 8728 6180
rect 8773 6158 8774 6168
rect 8789 6158 8802 6168
rect 8773 6154 8802 6158
rect 8807 6154 8837 6180
rect 8855 6166 8871 6168
rect 8943 6166 8996 6180
rect 8944 6164 9008 6166
rect 9051 6164 9066 6180
rect 9115 6177 9145 6180
rect 9115 6174 9151 6177
rect 9081 6166 9097 6168
rect 8855 6154 8870 6158
rect 8773 6152 8870 6154
rect 8898 6152 9066 6164
rect 9082 6154 9097 6158
rect 9115 6155 9154 6174
rect 9173 6168 9180 6169
rect 9179 6161 9180 6168
rect 9163 6158 9164 6161
rect 9179 6158 9192 6161
rect 9115 6154 9145 6155
rect 9154 6154 9160 6155
rect 9163 6154 9192 6158
rect 9082 6153 9192 6154
rect 9082 6152 9198 6153
rect 8757 6144 8808 6152
rect 8757 6132 8782 6144
rect 8789 6132 8808 6144
rect 8839 6144 8889 6152
rect 8839 6136 8855 6144
rect 8862 6142 8889 6144
rect 8898 6142 9119 6152
rect 8862 6132 9119 6142
rect 9148 6144 9198 6152
rect 9148 6135 9164 6144
rect 8757 6124 8808 6132
rect 8855 6124 9119 6132
rect 9145 6132 9164 6135
rect 9171 6132 9198 6144
rect 9145 6124 9198 6132
rect 8773 6116 8774 6124
rect 8789 6116 8802 6124
rect 8773 6108 8789 6116
rect 8770 6101 8789 6104
rect 8770 6092 8792 6101
rect 8743 6082 8792 6092
rect 8743 6076 8773 6082
rect 8792 6077 8797 6082
rect 8715 6060 8789 6076
rect 8807 6068 8837 6124
rect 8872 6114 9080 6124
rect 9115 6120 9160 6124
rect 9163 6123 9164 6124
rect 9179 6123 9192 6124
rect 8898 6084 9087 6114
rect 8913 6081 9087 6084
rect 8906 6078 9087 6081
rect 8715 6058 8728 6060
rect 8743 6058 8777 6060
rect 8715 6042 8789 6058
rect 8816 6054 8829 6068
rect 8844 6054 8860 6070
rect 8906 6065 8917 6078
rect 8699 6020 8700 6036
rect 8715 6020 8728 6042
rect 8743 6020 8773 6042
rect 8816 6038 8878 6054
rect 8906 6047 8917 6063
rect 8922 6058 8932 6078
rect 8942 6058 8956 6078
rect 8959 6065 8968 6078
rect 8984 6065 8993 6078
rect 8922 6047 8956 6058
rect 8959 6047 8968 6063
rect 8984 6047 8993 6063
rect 9000 6058 9010 6078
rect 9020 6058 9034 6078
rect 9035 6065 9046 6078
rect 9000 6047 9034 6058
rect 9035 6047 9046 6063
rect 9092 6054 9108 6070
rect 9115 6068 9145 6120
rect 9179 6116 9180 6123
rect 9164 6108 9180 6116
rect 9151 6076 9164 6095
rect 9179 6076 9209 6092
rect 9151 6060 9225 6076
rect 9151 6058 9164 6060
rect 9179 6058 9213 6060
rect 8816 6036 8829 6038
rect 8844 6036 8878 6038
rect 8816 6020 8878 6036
rect 8922 6031 8938 6034
rect 9000 6031 9030 6042
rect 9078 6038 9124 6054
rect 9151 6042 9225 6058
rect 9078 6036 9112 6038
rect 9077 6020 9124 6036
rect 9151 6020 9164 6042
rect 9179 6020 9209 6042
rect 9236 6020 9237 6036
rect 9252 6020 9265 6180
rect -7 6012 34 6020
rect -7 5986 8 6012
rect 15 5986 34 6012
rect 98 6008 160 6020
rect 172 6008 247 6020
rect 305 6008 380 6020
rect 392 6008 423 6020
rect 429 6008 464 6020
rect 98 6006 260 6008
rect -7 5978 34 5986
rect 116 5982 129 6006
rect 144 6004 159 6006
rect -1 5968 0 5978
rect 15 5968 28 5978
rect 43 5968 73 5982
rect 116 5968 159 5982
rect 183 5979 190 5986
rect 193 5982 260 6006
rect 292 6006 464 6008
rect 262 5984 290 5988
rect 292 5984 372 6006
rect 393 6004 408 6006
rect 262 5982 372 5984
rect 193 5978 372 5982
rect 166 5968 196 5978
rect 198 5968 351 5978
rect 359 5968 389 5978
rect 393 5968 423 5982
rect 451 5968 464 6006
rect 536 6012 571 6020
rect 536 5986 537 6012
rect 544 5986 571 6012
rect 479 5968 509 5982
rect 536 5978 571 5986
rect 573 6012 614 6020
rect 573 5986 588 6012
rect 595 5986 614 6012
rect 678 6008 740 6020
rect 752 6008 827 6020
rect 885 6008 960 6020
rect 972 6008 1003 6020
rect 1009 6008 1044 6020
rect 678 6006 840 6008
rect 573 5978 614 5986
rect 696 5982 709 6006
rect 724 6004 739 6006
rect 536 5968 537 5978
rect 552 5968 565 5978
rect 579 5968 580 5978
rect 595 5968 608 5978
rect 623 5968 653 5982
rect 696 5968 739 5982
rect 763 5979 770 5986
rect 773 5982 840 6006
rect 872 6006 1044 6008
rect 842 5984 870 5988
rect 872 5984 952 6006
rect 973 6004 988 6006
rect 842 5982 952 5984
rect 773 5978 952 5982
rect 746 5968 776 5978
rect 778 5968 931 5978
rect 939 5968 969 5978
rect 973 5968 1003 5982
rect 1031 5968 1044 6006
rect 1116 6012 1151 6020
rect 1116 5986 1117 6012
rect 1124 5986 1151 6012
rect 1059 5968 1089 5982
rect 1116 5978 1151 5986
rect 1153 6012 1194 6020
rect 1153 5986 1168 6012
rect 1175 5986 1194 6012
rect 1258 6008 1320 6020
rect 1332 6008 1407 6020
rect 1465 6008 1540 6020
rect 1552 6008 1583 6020
rect 1589 6008 1624 6020
rect 1258 6006 1420 6008
rect 1153 5978 1194 5986
rect 1276 5982 1289 6006
rect 1304 6004 1319 6006
rect 1116 5968 1117 5978
rect 1132 5968 1145 5978
rect 1159 5968 1160 5978
rect 1175 5968 1188 5978
rect 1203 5968 1233 5982
rect 1276 5968 1319 5982
rect 1343 5979 1350 5986
rect 1353 5982 1420 6006
rect 1452 6006 1624 6008
rect 1422 5984 1450 5988
rect 1452 5984 1532 6006
rect 1553 6004 1568 6006
rect 1422 5982 1532 5984
rect 1353 5978 1532 5982
rect 1326 5968 1356 5978
rect 1358 5968 1511 5978
rect 1519 5968 1549 5978
rect 1553 5968 1583 5982
rect 1611 5968 1624 6006
rect 1696 6012 1731 6020
rect 1696 5986 1697 6012
rect 1704 5986 1731 6012
rect 1639 5968 1669 5982
rect 1696 5978 1731 5986
rect 1733 6012 1774 6020
rect 1733 5986 1748 6012
rect 1755 5986 1774 6012
rect 1838 6008 1900 6020
rect 1912 6008 1987 6020
rect 2045 6008 2120 6020
rect 2132 6008 2163 6020
rect 2169 6008 2204 6020
rect 1838 6006 2000 6008
rect 1733 5978 1774 5986
rect 1856 5982 1869 6006
rect 1884 6004 1899 6006
rect 1696 5968 1697 5978
rect 1712 5968 1725 5978
rect 1739 5968 1740 5978
rect 1755 5968 1768 5978
rect 1783 5968 1813 5982
rect 1856 5968 1899 5982
rect 1923 5979 1930 5986
rect 1933 5982 2000 6006
rect 2032 6006 2204 6008
rect 2002 5984 2030 5988
rect 2032 5984 2112 6006
rect 2133 6004 2148 6006
rect 2002 5982 2112 5984
rect 1933 5978 2112 5982
rect 1906 5968 1936 5978
rect 1938 5968 2091 5978
rect 2099 5968 2129 5978
rect 2133 5968 2163 5982
rect 2191 5968 2204 6006
rect 2276 6012 2311 6020
rect 2276 5986 2277 6012
rect 2284 5986 2311 6012
rect 2219 5968 2249 5982
rect 2276 5978 2311 5986
rect 2313 6012 2354 6020
rect 2313 5986 2328 6012
rect 2335 5986 2354 6012
rect 2418 6008 2480 6020
rect 2492 6008 2567 6020
rect 2625 6008 2700 6020
rect 2712 6008 2743 6020
rect 2749 6008 2784 6020
rect 2418 6006 2580 6008
rect 2313 5978 2354 5986
rect 2436 5982 2449 6006
rect 2464 6004 2479 6006
rect 2276 5968 2277 5978
rect 2292 5968 2305 5978
rect 2319 5968 2320 5978
rect 2335 5968 2348 5978
rect 2363 5968 2393 5982
rect 2436 5968 2479 5982
rect 2503 5979 2510 5986
rect 2513 5982 2580 6006
rect 2612 6006 2784 6008
rect 2582 5984 2610 5988
rect 2612 5984 2692 6006
rect 2713 6004 2728 6006
rect 2582 5982 2692 5984
rect 2513 5978 2692 5982
rect 2486 5968 2516 5978
rect 2518 5968 2671 5978
rect 2679 5968 2709 5978
rect 2713 5968 2743 5982
rect 2771 5968 2784 6006
rect 2856 6012 2891 6020
rect 2856 5986 2857 6012
rect 2864 5986 2891 6012
rect 2799 5968 2829 5982
rect 2856 5978 2891 5986
rect 2893 6012 2934 6020
rect 2893 5986 2908 6012
rect 2915 5986 2934 6012
rect 2998 6008 3060 6020
rect 3072 6008 3147 6020
rect 3205 6008 3280 6020
rect 3292 6008 3323 6020
rect 3329 6008 3364 6020
rect 2998 6006 3160 6008
rect 2893 5978 2934 5986
rect 3016 5982 3029 6006
rect 3044 6004 3059 6006
rect 2856 5968 2857 5978
rect 2872 5968 2885 5978
rect 2899 5968 2900 5978
rect 2915 5968 2928 5978
rect 2943 5968 2973 5982
rect 3016 5968 3059 5982
rect 3083 5979 3090 5986
rect 3093 5982 3160 6006
rect 3192 6006 3364 6008
rect 3162 5984 3190 5988
rect 3192 5984 3272 6006
rect 3293 6004 3308 6006
rect 3162 5982 3272 5984
rect 3093 5978 3272 5982
rect 3066 5968 3096 5978
rect 3098 5968 3251 5978
rect 3259 5968 3289 5978
rect 3293 5968 3323 5982
rect 3351 5968 3364 6006
rect 3436 6012 3471 6020
rect 3436 5986 3437 6012
rect 3444 5986 3471 6012
rect 3379 5968 3409 5982
rect 3436 5978 3471 5986
rect 3473 6012 3514 6020
rect 3473 5986 3488 6012
rect 3495 5986 3514 6012
rect 3578 6008 3640 6020
rect 3652 6008 3727 6020
rect 3785 6008 3860 6020
rect 3872 6008 3903 6020
rect 3909 6008 3944 6020
rect 3578 6006 3740 6008
rect 3473 5978 3514 5986
rect 3596 5982 3609 6006
rect 3624 6004 3639 6006
rect 3436 5968 3437 5978
rect 3452 5968 3465 5978
rect 3479 5968 3480 5978
rect 3495 5968 3508 5978
rect 3523 5968 3553 5982
rect 3596 5968 3639 5982
rect 3663 5979 3670 5986
rect 3673 5982 3740 6006
rect 3772 6006 3944 6008
rect 3742 5984 3770 5988
rect 3772 5984 3852 6006
rect 3873 6004 3888 6006
rect 3742 5982 3852 5984
rect 3673 5978 3852 5982
rect 3646 5968 3676 5978
rect 3678 5968 3831 5978
rect 3839 5968 3869 5978
rect 3873 5968 3903 5982
rect 3931 5968 3944 6006
rect 4016 6012 4051 6020
rect 4016 5986 4017 6012
rect 4024 5986 4051 6012
rect 3959 5968 3989 5982
rect 4016 5978 4051 5986
rect 4053 6012 4094 6020
rect 4053 5986 4068 6012
rect 4075 5986 4094 6012
rect 4158 6008 4220 6020
rect 4232 6008 4307 6020
rect 4365 6008 4440 6020
rect 4452 6008 4483 6020
rect 4489 6008 4524 6020
rect 4158 6006 4320 6008
rect 4053 5978 4094 5986
rect 4176 5982 4189 6006
rect 4204 6004 4219 6006
rect 4016 5968 4017 5978
rect 4032 5968 4045 5978
rect 4059 5968 4060 5978
rect 4075 5968 4088 5978
rect 4103 5968 4133 5982
rect 4176 5968 4219 5982
rect 4243 5979 4250 5986
rect 4253 5982 4320 6006
rect 4352 6006 4524 6008
rect 4322 5984 4350 5988
rect 4352 5984 4432 6006
rect 4453 6004 4468 6006
rect 4322 5982 4432 5984
rect 4253 5978 4432 5982
rect 4226 5968 4256 5978
rect 4258 5968 4411 5978
rect 4419 5968 4449 5978
rect 4453 5968 4483 5982
rect 4511 5968 4524 6006
rect 4596 6012 4631 6020
rect 4596 5986 4597 6012
rect 4604 5986 4631 6012
rect 4539 5968 4569 5982
rect 4596 5978 4631 5986
rect 4633 6012 4674 6020
rect 4633 5986 4648 6012
rect 4655 5986 4674 6012
rect 4738 6008 4800 6020
rect 4812 6008 4887 6020
rect 4945 6008 5020 6020
rect 5032 6008 5063 6020
rect 5069 6008 5104 6020
rect 4738 6006 4900 6008
rect 4633 5978 4674 5986
rect 4756 5982 4769 6006
rect 4784 6004 4799 6006
rect 4596 5968 4597 5978
rect 4612 5968 4625 5978
rect 4639 5968 4640 5978
rect 4655 5968 4668 5978
rect 4683 5968 4713 5982
rect 4756 5968 4799 5982
rect 4823 5979 4830 5986
rect 4833 5982 4900 6006
rect 4932 6006 5104 6008
rect 4902 5984 4930 5988
rect 4932 5984 5012 6006
rect 5033 6004 5048 6006
rect 4902 5982 5012 5984
rect 4833 5978 5012 5982
rect 4806 5968 4836 5978
rect 4838 5968 4991 5978
rect 4999 5968 5029 5978
rect 5033 5968 5063 5982
rect 5091 5968 5104 6006
rect 5176 6012 5211 6020
rect 5176 5986 5177 6012
rect 5184 5986 5211 6012
rect 5119 5968 5149 5982
rect 5176 5978 5211 5986
rect 5213 6012 5254 6020
rect 5213 5986 5228 6012
rect 5235 5986 5254 6012
rect 5318 6008 5380 6020
rect 5392 6008 5467 6020
rect 5525 6008 5600 6020
rect 5612 6008 5643 6020
rect 5649 6008 5684 6020
rect 5318 6006 5480 6008
rect 5213 5978 5254 5986
rect 5336 5982 5349 6006
rect 5364 6004 5379 6006
rect 5176 5968 5177 5978
rect 5192 5968 5205 5978
rect 5219 5968 5220 5978
rect 5235 5968 5248 5978
rect 5263 5968 5293 5982
rect 5336 5968 5379 5982
rect 5403 5979 5410 5986
rect 5413 5982 5480 6006
rect 5512 6006 5684 6008
rect 5482 5984 5510 5988
rect 5512 5984 5592 6006
rect 5613 6004 5628 6006
rect 5482 5982 5592 5984
rect 5413 5978 5592 5982
rect 5386 5968 5416 5978
rect 5418 5968 5571 5978
rect 5579 5968 5609 5978
rect 5613 5968 5643 5982
rect 5671 5968 5684 6006
rect 5756 6012 5791 6020
rect 5756 5986 5757 6012
rect 5764 5986 5791 6012
rect 5699 5968 5729 5982
rect 5756 5978 5791 5986
rect 5793 6012 5834 6020
rect 5793 5986 5808 6012
rect 5815 5986 5834 6012
rect 5898 6008 5960 6020
rect 5972 6008 6047 6020
rect 6105 6008 6180 6020
rect 6192 6008 6223 6020
rect 6229 6008 6264 6020
rect 5898 6006 6060 6008
rect 5793 5978 5834 5986
rect 5916 5982 5929 6006
rect 5944 6004 5959 6006
rect 5756 5968 5757 5978
rect 5772 5968 5785 5978
rect 5799 5968 5800 5978
rect 5815 5968 5828 5978
rect 5843 5968 5873 5982
rect 5916 5968 5959 5982
rect 5983 5979 5990 5986
rect 5993 5982 6060 6006
rect 6092 6006 6264 6008
rect 6062 5984 6090 5988
rect 6092 5984 6172 6006
rect 6193 6004 6208 6006
rect 6062 5982 6172 5984
rect 5993 5978 6172 5982
rect 5966 5968 5996 5978
rect 5998 5968 6151 5978
rect 6159 5968 6189 5978
rect 6193 5968 6223 5982
rect 6251 5968 6264 6006
rect 6336 6012 6371 6020
rect 6336 5986 6337 6012
rect 6344 5986 6371 6012
rect 6279 5968 6309 5982
rect 6336 5978 6371 5986
rect 6373 6012 6414 6020
rect 6373 5986 6388 6012
rect 6395 5986 6414 6012
rect 6478 6008 6540 6020
rect 6552 6008 6627 6020
rect 6685 6008 6760 6020
rect 6772 6008 6803 6020
rect 6809 6008 6844 6020
rect 6478 6006 6640 6008
rect 6373 5978 6414 5986
rect 6496 5982 6509 6006
rect 6524 6004 6539 6006
rect 6336 5968 6337 5978
rect 6352 5968 6365 5978
rect 6379 5968 6380 5978
rect 6395 5968 6408 5978
rect 6423 5968 6453 5982
rect 6496 5968 6539 5982
rect 6563 5979 6570 5986
rect 6573 5982 6640 6006
rect 6672 6006 6844 6008
rect 6642 5984 6670 5988
rect 6672 5984 6752 6006
rect 6773 6004 6788 6006
rect 6642 5982 6752 5984
rect 6573 5978 6752 5982
rect 6546 5968 6576 5978
rect 6578 5968 6731 5978
rect 6739 5968 6769 5978
rect 6773 5968 6803 5982
rect 6831 5968 6844 6006
rect 6916 6012 6951 6020
rect 6916 5986 6917 6012
rect 6924 5986 6951 6012
rect 6859 5968 6889 5982
rect 6916 5978 6951 5986
rect 6953 6012 6994 6020
rect 6953 5986 6968 6012
rect 6975 5986 6994 6012
rect 7058 6008 7120 6020
rect 7132 6008 7207 6020
rect 7265 6008 7340 6020
rect 7352 6008 7383 6020
rect 7389 6008 7424 6020
rect 7058 6006 7220 6008
rect 6953 5978 6994 5986
rect 7076 5982 7089 6006
rect 7104 6004 7119 6006
rect 6916 5968 6917 5978
rect 6932 5968 6945 5978
rect 6959 5968 6960 5978
rect 6975 5968 6988 5978
rect 7003 5968 7033 5982
rect 7076 5968 7119 5982
rect 7143 5979 7150 5986
rect 7153 5982 7220 6006
rect 7252 6006 7424 6008
rect 7222 5984 7250 5988
rect 7252 5984 7332 6006
rect 7353 6004 7368 6006
rect 7222 5982 7332 5984
rect 7153 5978 7332 5982
rect 7126 5968 7156 5978
rect 7158 5968 7311 5978
rect 7319 5968 7349 5978
rect 7353 5968 7383 5982
rect 7411 5968 7424 6006
rect 7496 6012 7531 6020
rect 7496 5986 7497 6012
rect 7504 5986 7531 6012
rect 7439 5968 7469 5982
rect 7496 5978 7531 5986
rect 7533 6012 7574 6020
rect 7533 5986 7548 6012
rect 7555 5986 7574 6012
rect 7638 6008 7700 6020
rect 7712 6008 7787 6020
rect 7845 6008 7920 6020
rect 7932 6008 7963 6020
rect 7969 6008 8004 6020
rect 7638 6006 7800 6008
rect 7533 5978 7574 5986
rect 7656 5982 7669 6006
rect 7684 6004 7699 6006
rect 7496 5968 7497 5978
rect 7512 5968 7525 5978
rect 7539 5968 7540 5978
rect 7555 5968 7568 5978
rect 7583 5968 7613 5982
rect 7656 5968 7699 5982
rect 7723 5979 7730 5986
rect 7733 5982 7800 6006
rect 7832 6006 8004 6008
rect 7802 5984 7830 5988
rect 7832 5984 7912 6006
rect 7933 6004 7948 6006
rect 7802 5982 7912 5984
rect 7733 5978 7912 5982
rect 7706 5968 7736 5978
rect 7738 5968 7891 5978
rect 7899 5968 7929 5978
rect 7933 5968 7963 5982
rect 7991 5968 8004 6006
rect 8076 6012 8111 6020
rect 8076 5986 8077 6012
rect 8084 5986 8111 6012
rect 8019 5968 8049 5982
rect 8076 5978 8111 5986
rect 8113 6012 8154 6020
rect 8113 5986 8128 6012
rect 8135 5986 8154 6012
rect 8218 6008 8280 6020
rect 8292 6008 8367 6020
rect 8425 6008 8500 6020
rect 8512 6008 8543 6020
rect 8549 6008 8584 6020
rect 8218 6006 8380 6008
rect 8113 5978 8154 5986
rect 8236 5982 8249 6006
rect 8264 6004 8279 6006
rect 8076 5968 8077 5978
rect 8092 5968 8105 5978
rect 8119 5968 8120 5978
rect 8135 5968 8148 5978
rect 8163 5968 8193 5982
rect 8236 5968 8279 5982
rect 8303 5979 8310 5986
rect 8313 5982 8380 6006
rect 8412 6006 8584 6008
rect 8382 5984 8410 5988
rect 8412 5984 8492 6006
rect 8513 6004 8528 6006
rect 8382 5982 8492 5984
rect 8313 5978 8492 5982
rect 8286 5968 8316 5978
rect 8318 5968 8471 5978
rect 8479 5968 8509 5978
rect 8513 5968 8543 5982
rect 8571 5968 8584 6006
rect 8656 6012 8691 6020
rect 8656 5986 8657 6012
rect 8664 5986 8691 6012
rect 8599 5968 8629 5982
rect 8656 5978 8691 5986
rect 8693 6012 8734 6020
rect 8693 5986 8708 6012
rect 8715 5986 8734 6012
rect 8798 6008 8860 6020
rect 8872 6008 8947 6020
rect 9005 6008 9080 6020
rect 9092 6008 9123 6020
rect 9129 6008 9164 6020
rect 8798 6006 8960 6008
rect 8693 5978 8734 5986
rect 8816 5982 8829 6006
rect 8844 6004 8859 6006
rect 8656 5968 8657 5978
rect 8672 5968 8685 5978
rect 8699 5968 8700 5978
rect 8715 5968 8728 5978
rect 8743 5968 8773 5982
rect 8816 5968 8859 5982
rect 8883 5979 8890 5986
rect 8893 5982 8960 6006
rect 8992 6006 9164 6008
rect 8962 5984 8990 5988
rect 8992 5984 9072 6006
rect 9093 6004 9108 6006
rect 8962 5982 9072 5984
rect 8893 5978 9072 5982
rect 8866 5968 8896 5978
rect 8898 5968 9051 5978
rect 9059 5968 9089 5978
rect 9093 5968 9123 5982
rect 9151 5968 9164 6006
rect 9236 6012 9271 6020
rect 9236 5986 9237 6012
rect 9244 5986 9271 6012
rect 9179 5968 9209 5982
rect 9236 5978 9271 5986
rect 9236 5968 9237 5978
rect 9252 5968 9265 5978
rect -1 5962 9265 5968
rect 0 5954 9265 5962
rect 15 5924 28 5954
rect 43 5936 73 5954
rect 116 5940 130 5954
rect 166 5940 386 5954
rect 117 5938 130 5940
rect 83 5926 98 5938
rect 80 5924 102 5926
rect 107 5924 137 5938
rect 198 5936 351 5940
rect 180 5924 372 5936
rect 415 5924 445 5938
rect 451 5924 464 5954
rect 479 5936 509 5954
rect 552 5924 565 5954
rect 595 5924 608 5954
rect 623 5936 653 5954
rect 696 5940 710 5954
rect 746 5940 966 5954
rect 697 5938 710 5940
rect 663 5926 678 5938
rect 660 5924 682 5926
rect 687 5924 717 5938
rect 778 5936 931 5940
rect 760 5924 952 5936
rect 995 5924 1025 5938
rect 1031 5924 1044 5954
rect 1059 5936 1089 5954
rect 1132 5924 1145 5954
rect 1175 5924 1188 5954
rect 1203 5936 1233 5954
rect 1276 5940 1290 5954
rect 1326 5940 1546 5954
rect 1277 5938 1290 5940
rect 1243 5926 1258 5938
rect 1240 5924 1262 5926
rect 1267 5924 1297 5938
rect 1358 5936 1511 5940
rect 1340 5924 1532 5936
rect 1575 5924 1605 5938
rect 1611 5924 1624 5954
rect 1639 5936 1669 5954
rect 1712 5924 1725 5954
rect 1755 5924 1768 5954
rect 1783 5936 1813 5954
rect 1856 5940 1870 5954
rect 1906 5940 2126 5954
rect 1857 5938 1870 5940
rect 1823 5926 1838 5938
rect 1820 5924 1842 5926
rect 1847 5924 1877 5938
rect 1938 5936 2091 5940
rect 1920 5924 2112 5936
rect 2155 5924 2185 5938
rect 2191 5924 2204 5954
rect 2219 5936 2249 5954
rect 2292 5924 2305 5954
rect 2335 5924 2348 5954
rect 2363 5936 2393 5954
rect 2436 5940 2450 5954
rect 2486 5940 2706 5954
rect 2437 5938 2450 5940
rect 2403 5926 2418 5938
rect 2400 5924 2422 5926
rect 2427 5924 2457 5938
rect 2518 5936 2671 5940
rect 2500 5924 2692 5936
rect 2735 5924 2765 5938
rect 2771 5924 2784 5954
rect 2799 5936 2829 5954
rect 2872 5924 2885 5954
rect 2915 5924 2928 5954
rect 2943 5936 2973 5954
rect 3016 5940 3030 5954
rect 3066 5940 3286 5954
rect 3017 5938 3030 5940
rect 2983 5926 2998 5938
rect 2980 5924 3002 5926
rect 3007 5924 3037 5938
rect 3098 5936 3251 5940
rect 3080 5924 3272 5936
rect 3315 5924 3345 5938
rect 3351 5924 3364 5954
rect 3379 5936 3409 5954
rect 3452 5924 3465 5954
rect 3495 5924 3508 5954
rect 3523 5936 3553 5954
rect 3596 5940 3610 5954
rect 3646 5940 3866 5954
rect 3597 5938 3610 5940
rect 3563 5926 3578 5938
rect 3560 5924 3582 5926
rect 3587 5924 3617 5938
rect 3678 5936 3831 5940
rect 3660 5924 3852 5936
rect 3895 5924 3925 5938
rect 3931 5924 3944 5954
rect 3959 5936 3989 5954
rect 4032 5924 4045 5954
rect 4075 5924 4088 5954
rect 4103 5936 4133 5954
rect 4176 5940 4190 5954
rect 4226 5940 4446 5954
rect 4177 5938 4190 5940
rect 4143 5926 4158 5938
rect 4140 5924 4162 5926
rect 4167 5924 4197 5938
rect 4258 5936 4411 5940
rect 4240 5924 4432 5936
rect 4475 5924 4505 5938
rect 4511 5924 4524 5954
rect 4539 5936 4569 5954
rect 4612 5924 4625 5954
rect 4655 5924 4668 5954
rect 4683 5936 4713 5954
rect 4756 5940 4770 5954
rect 4806 5940 5026 5954
rect 4757 5938 4770 5940
rect 4723 5926 4738 5938
rect 4720 5924 4742 5926
rect 4747 5924 4777 5938
rect 4838 5936 4991 5940
rect 4820 5924 5012 5936
rect 5055 5924 5085 5938
rect 5091 5924 5104 5954
rect 5119 5936 5149 5954
rect 5192 5924 5205 5954
rect 5235 5924 5248 5954
rect 5263 5936 5293 5954
rect 5336 5940 5350 5954
rect 5386 5940 5606 5954
rect 5337 5938 5350 5940
rect 5303 5926 5318 5938
rect 5300 5924 5322 5926
rect 5327 5924 5357 5938
rect 5418 5936 5571 5940
rect 5400 5924 5592 5936
rect 5635 5924 5665 5938
rect 5671 5924 5684 5954
rect 5699 5936 5729 5954
rect 5772 5924 5785 5954
rect 5815 5924 5828 5954
rect 5843 5936 5873 5954
rect 5916 5940 5930 5954
rect 5966 5940 6186 5954
rect 5917 5938 5930 5940
rect 5883 5926 5898 5938
rect 5880 5924 5902 5926
rect 5907 5924 5937 5938
rect 5998 5936 6151 5940
rect 5980 5924 6172 5936
rect 6215 5924 6245 5938
rect 6251 5924 6264 5954
rect 6279 5936 6309 5954
rect 6352 5924 6365 5954
rect 6395 5924 6408 5954
rect 6423 5936 6453 5954
rect 6496 5940 6510 5954
rect 6546 5940 6766 5954
rect 6497 5938 6510 5940
rect 6463 5926 6478 5938
rect 6460 5924 6482 5926
rect 6487 5924 6517 5938
rect 6578 5936 6731 5940
rect 6560 5924 6752 5936
rect 6795 5924 6825 5938
rect 6831 5924 6844 5954
rect 6859 5936 6889 5954
rect 6932 5924 6945 5954
rect 6975 5924 6988 5954
rect 7003 5936 7033 5954
rect 7076 5940 7090 5954
rect 7126 5940 7346 5954
rect 7077 5938 7090 5940
rect 7043 5926 7058 5938
rect 7040 5924 7062 5926
rect 7067 5924 7097 5938
rect 7158 5936 7311 5940
rect 7140 5924 7332 5936
rect 7375 5924 7405 5938
rect 7411 5924 7424 5954
rect 7439 5936 7469 5954
rect 7512 5924 7525 5954
rect 7555 5924 7568 5954
rect 7583 5936 7613 5954
rect 7656 5940 7670 5954
rect 7706 5940 7926 5954
rect 7657 5938 7670 5940
rect 7623 5926 7638 5938
rect 7620 5924 7642 5926
rect 7647 5924 7677 5938
rect 7738 5936 7891 5940
rect 7720 5924 7912 5936
rect 7955 5924 7985 5938
rect 7991 5924 8004 5954
rect 8019 5936 8049 5954
rect 8092 5924 8105 5954
rect 8135 5924 8148 5954
rect 8163 5936 8193 5954
rect 8236 5940 8250 5954
rect 8286 5940 8506 5954
rect 8237 5938 8250 5940
rect 8203 5926 8218 5938
rect 8200 5924 8222 5926
rect 8227 5924 8257 5938
rect 8318 5936 8471 5940
rect 8300 5924 8492 5936
rect 8535 5924 8565 5938
rect 8571 5924 8584 5954
rect 8599 5936 8629 5954
rect 8672 5924 8685 5954
rect 8715 5924 8728 5954
rect 8743 5936 8773 5954
rect 8816 5940 8830 5954
rect 8866 5940 9086 5954
rect 8817 5938 8830 5940
rect 8783 5926 8798 5938
rect 8780 5924 8802 5926
rect 8807 5924 8837 5938
rect 8898 5936 9051 5940
rect 8880 5924 9072 5936
rect 9115 5924 9145 5938
rect 9151 5924 9164 5954
rect 9179 5936 9209 5954
rect 9252 5924 9265 5954
rect 0 5910 9265 5924
rect 15 5806 28 5910
rect 73 5888 74 5898
rect 89 5888 102 5898
rect 73 5884 102 5888
rect 107 5884 137 5910
rect 155 5896 171 5898
rect 243 5896 296 5910
rect 244 5894 308 5896
rect 351 5894 366 5910
rect 415 5907 445 5910
rect 415 5904 451 5907
rect 381 5896 397 5898
rect 155 5884 170 5888
rect 73 5882 170 5884
rect 198 5882 366 5894
rect 382 5884 397 5888
rect 415 5885 454 5904
rect 473 5898 480 5899
rect 479 5891 480 5898
rect 463 5888 464 5891
rect 479 5888 492 5891
rect 415 5884 445 5885
rect 454 5884 460 5885
rect 463 5884 492 5888
rect 382 5883 492 5884
rect 382 5882 498 5883
rect 57 5874 108 5882
rect 57 5862 82 5874
rect 89 5862 108 5874
rect 139 5874 189 5882
rect 139 5866 155 5874
rect 162 5872 189 5874
rect 198 5872 419 5882
rect 162 5862 419 5872
rect 448 5874 498 5882
rect 448 5865 464 5874
rect 57 5854 108 5862
rect 155 5854 419 5862
rect 445 5862 464 5865
rect 471 5862 498 5874
rect 445 5854 498 5862
rect 73 5846 74 5854
rect 89 5846 102 5854
rect 73 5838 89 5846
rect 70 5831 89 5834
rect 70 5822 92 5831
rect 43 5812 92 5822
rect 43 5806 73 5812
rect 92 5807 97 5812
rect 15 5790 89 5806
rect 107 5798 137 5854
rect 172 5844 380 5854
rect 415 5850 460 5854
rect 463 5853 464 5854
rect 479 5853 492 5854
rect 198 5814 387 5844
rect 213 5811 387 5814
rect 206 5808 387 5811
rect 15 5788 28 5790
rect 43 5788 77 5790
rect 15 5772 89 5788
rect 116 5784 129 5798
rect 144 5784 160 5800
rect 206 5795 217 5808
rect -1 5750 0 5766
rect 15 5750 28 5772
rect 43 5750 73 5772
rect 116 5768 178 5784
rect 206 5777 217 5793
rect 222 5788 232 5808
rect 242 5788 256 5808
rect 259 5795 268 5808
rect 284 5795 293 5808
rect 222 5777 256 5788
rect 259 5777 268 5793
rect 284 5777 293 5793
rect 300 5788 310 5808
rect 320 5788 334 5808
rect 335 5795 346 5808
rect 300 5777 334 5788
rect 335 5777 346 5793
rect 392 5784 408 5800
rect 415 5798 445 5850
rect 479 5846 480 5853
rect 464 5838 480 5846
rect 451 5806 464 5825
rect 479 5806 509 5822
rect 451 5790 525 5806
rect 451 5788 464 5790
rect 479 5788 513 5790
rect 116 5766 129 5768
rect 144 5766 178 5768
rect 116 5750 178 5766
rect 222 5761 238 5764
rect 300 5761 330 5772
rect 378 5768 424 5784
rect 451 5772 525 5788
rect 378 5766 412 5768
rect 377 5750 424 5766
rect 451 5750 464 5772
rect 479 5750 509 5772
rect 536 5750 537 5766
rect 552 5750 565 5910
rect 595 5806 608 5910
rect 653 5888 654 5898
rect 669 5888 682 5898
rect 653 5884 682 5888
rect 687 5884 717 5910
rect 735 5896 751 5898
rect 823 5896 876 5910
rect 824 5894 888 5896
rect 931 5894 946 5910
rect 995 5907 1025 5910
rect 995 5904 1031 5907
rect 961 5896 977 5898
rect 735 5884 750 5888
rect 653 5882 750 5884
rect 778 5882 946 5894
rect 962 5884 977 5888
rect 995 5885 1034 5904
rect 1053 5898 1060 5899
rect 1059 5891 1060 5898
rect 1043 5888 1044 5891
rect 1059 5888 1072 5891
rect 995 5884 1025 5885
rect 1034 5884 1040 5885
rect 1043 5884 1072 5888
rect 962 5883 1072 5884
rect 962 5882 1078 5883
rect 637 5874 688 5882
rect 637 5862 662 5874
rect 669 5862 688 5874
rect 719 5874 769 5882
rect 719 5866 735 5874
rect 742 5872 769 5874
rect 778 5872 999 5882
rect 742 5862 999 5872
rect 1028 5874 1078 5882
rect 1028 5865 1044 5874
rect 637 5854 688 5862
rect 735 5854 999 5862
rect 1025 5862 1044 5865
rect 1051 5862 1078 5874
rect 1025 5854 1078 5862
rect 653 5846 654 5854
rect 669 5846 682 5854
rect 653 5838 669 5846
rect 650 5831 669 5834
rect 650 5822 672 5831
rect 623 5812 672 5822
rect 623 5806 653 5812
rect 672 5807 677 5812
rect 595 5790 669 5806
rect 687 5798 717 5854
rect 752 5844 960 5854
rect 995 5850 1040 5854
rect 1043 5853 1044 5854
rect 1059 5853 1072 5854
rect 778 5814 967 5844
rect 793 5811 967 5814
rect 786 5808 967 5811
rect 595 5788 608 5790
rect 623 5788 657 5790
rect 595 5772 669 5788
rect 696 5784 709 5798
rect 724 5784 740 5800
rect 786 5795 797 5808
rect 579 5750 580 5766
rect 595 5750 608 5772
rect 623 5750 653 5772
rect 696 5768 758 5784
rect 786 5777 797 5793
rect 802 5788 812 5808
rect 822 5788 836 5808
rect 839 5795 848 5808
rect 864 5795 873 5808
rect 802 5777 836 5788
rect 839 5777 848 5793
rect 864 5777 873 5793
rect 880 5788 890 5808
rect 900 5788 914 5808
rect 915 5795 926 5808
rect 880 5777 914 5788
rect 915 5777 926 5793
rect 972 5784 988 5800
rect 995 5798 1025 5850
rect 1059 5846 1060 5853
rect 1044 5838 1060 5846
rect 1031 5806 1044 5825
rect 1059 5806 1089 5822
rect 1031 5790 1105 5806
rect 1031 5788 1044 5790
rect 1059 5788 1093 5790
rect 696 5766 709 5768
rect 724 5766 758 5768
rect 696 5750 758 5766
rect 802 5761 818 5764
rect 880 5761 910 5772
rect 958 5768 1004 5784
rect 1031 5772 1105 5788
rect 958 5766 992 5768
rect 957 5750 1004 5766
rect 1031 5750 1044 5772
rect 1059 5750 1089 5772
rect 1116 5750 1117 5766
rect 1132 5750 1145 5910
rect 1175 5806 1188 5910
rect 1233 5888 1234 5898
rect 1249 5888 1262 5898
rect 1233 5884 1262 5888
rect 1267 5884 1297 5910
rect 1315 5896 1331 5898
rect 1403 5896 1456 5910
rect 1404 5894 1468 5896
rect 1511 5894 1526 5910
rect 1575 5907 1605 5910
rect 1575 5904 1611 5907
rect 1541 5896 1557 5898
rect 1315 5884 1330 5888
rect 1233 5882 1330 5884
rect 1358 5882 1526 5894
rect 1542 5884 1557 5888
rect 1575 5885 1614 5904
rect 1633 5898 1640 5899
rect 1639 5891 1640 5898
rect 1623 5888 1624 5891
rect 1639 5888 1652 5891
rect 1575 5884 1605 5885
rect 1614 5884 1620 5885
rect 1623 5884 1652 5888
rect 1542 5883 1652 5884
rect 1542 5882 1658 5883
rect 1217 5874 1268 5882
rect 1217 5862 1242 5874
rect 1249 5862 1268 5874
rect 1299 5874 1349 5882
rect 1299 5866 1315 5874
rect 1322 5872 1349 5874
rect 1358 5872 1579 5882
rect 1322 5862 1579 5872
rect 1608 5874 1658 5882
rect 1608 5865 1624 5874
rect 1217 5854 1268 5862
rect 1315 5854 1579 5862
rect 1605 5862 1624 5865
rect 1631 5862 1658 5874
rect 1605 5854 1658 5862
rect 1233 5846 1234 5854
rect 1249 5846 1262 5854
rect 1233 5838 1249 5846
rect 1230 5831 1249 5834
rect 1230 5822 1252 5831
rect 1203 5812 1252 5822
rect 1203 5806 1233 5812
rect 1252 5807 1257 5812
rect 1175 5790 1249 5806
rect 1267 5798 1297 5854
rect 1332 5844 1540 5854
rect 1575 5850 1620 5854
rect 1623 5853 1624 5854
rect 1639 5853 1652 5854
rect 1358 5814 1547 5844
rect 1373 5811 1547 5814
rect 1366 5808 1547 5811
rect 1175 5788 1188 5790
rect 1203 5788 1237 5790
rect 1175 5772 1249 5788
rect 1276 5784 1289 5798
rect 1304 5784 1320 5800
rect 1366 5795 1377 5808
rect 1159 5750 1160 5766
rect 1175 5750 1188 5772
rect 1203 5750 1233 5772
rect 1276 5768 1338 5784
rect 1366 5777 1377 5793
rect 1382 5788 1392 5808
rect 1402 5788 1416 5808
rect 1419 5795 1428 5808
rect 1444 5795 1453 5808
rect 1382 5777 1416 5788
rect 1419 5777 1428 5793
rect 1444 5777 1453 5793
rect 1460 5788 1470 5808
rect 1480 5788 1494 5808
rect 1495 5795 1506 5808
rect 1460 5777 1494 5788
rect 1495 5777 1506 5793
rect 1552 5784 1568 5800
rect 1575 5798 1605 5850
rect 1639 5846 1640 5853
rect 1624 5838 1640 5846
rect 1611 5806 1624 5825
rect 1639 5806 1669 5822
rect 1611 5790 1685 5806
rect 1611 5788 1624 5790
rect 1639 5788 1673 5790
rect 1276 5766 1289 5768
rect 1304 5766 1338 5768
rect 1276 5750 1338 5766
rect 1382 5761 1398 5764
rect 1460 5761 1490 5772
rect 1538 5768 1584 5784
rect 1611 5772 1685 5788
rect 1538 5766 1572 5768
rect 1537 5750 1584 5766
rect 1611 5750 1624 5772
rect 1639 5750 1669 5772
rect 1696 5750 1697 5766
rect 1712 5750 1725 5910
rect 1755 5806 1768 5910
rect 1813 5888 1814 5898
rect 1829 5888 1842 5898
rect 1813 5884 1842 5888
rect 1847 5884 1877 5910
rect 1895 5896 1911 5898
rect 1983 5896 2036 5910
rect 1984 5894 2048 5896
rect 2091 5894 2106 5910
rect 2155 5907 2185 5910
rect 2155 5904 2191 5907
rect 2121 5896 2137 5898
rect 1895 5884 1910 5888
rect 1813 5882 1910 5884
rect 1938 5882 2106 5894
rect 2122 5884 2137 5888
rect 2155 5885 2194 5904
rect 2213 5898 2220 5899
rect 2219 5891 2220 5898
rect 2203 5888 2204 5891
rect 2219 5888 2232 5891
rect 2155 5884 2185 5885
rect 2194 5884 2200 5885
rect 2203 5884 2232 5888
rect 2122 5883 2232 5884
rect 2122 5882 2238 5883
rect 1797 5874 1848 5882
rect 1797 5862 1822 5874
rect 1829 5862 1848 5874
rect 1879 5874 1929 5882
rect 1879 5866 1895 5874
rect 1902 5872 1929 5874
rect 1938 5872 2159 5882
rect 1902 5862 2159 5872
rect 2188 5874 2238 5882
rect 2188 5865 2204 5874
rect 1797 5854 1848 5862
rect 1895 5854 2159 5862
rect 2185 5862 2204 5865
rect 2211 5862 2238 5874
rect 2185 5854 2238 5862
rect 1813 5846 1814 5854
rect 1829 5846 1842 5854
rect 1813 5838 1829 5846
rect 1810 5831 1829 5834
rect 1810 5822 1832 5831
rect 1783 5812 1832 5822
rect 1783 5806 1813 5812
rect 1832 5807 1837 5812
rect 1755 5790 1829 5806
rect 1847 5798 1877 5854
rect 1912 5844 2120 5854
rect 2155 5850 2200 5854
rect 2203 5853 2204 5854
rect 2219 5853 2232 5854
rect 1938 5814 2127 5844
rect 1953 5811 2127 5814
rect 1946 5808 2127 5811
rect 1755 5788 1768 5790
rect 1783 5788 1817 5790
rect 1755 5772 1829 5788
rect 1856 5784 1869 5798
rect 1884 5784 1900 5800
rect 1946 5795 1957 5808
rect 1739 5750 1740 5766
rect 1755 5750 1768 5772
rect 1783 5750 1813 5772
rect 1856 5768 1918 5784
rect 1946 5777 1957 5793
rect 1962 5788 1972 5808
rect 1982 5788 1996 5808
rect 1999 5795 2008 5808
rect 2024 5795 2033 5808
rect 1962 5777 1996 5788
rect 1999 5777 2008 5793
rect 2024 5777 2033 5793
rect 2040 5788 2050 5808
rect 2060 5788 2074 5808
rect 2075 5795 2086 5808
rect 2040 5777 2074 5788
rect 2075 5777 2086 5793
rect 2132 5784 2148 5800
rect 2155 5798 2185 5850
rect 2219 5846 2220 5853
rect 2204 5838 2220 5846
rect 2191 5806 2204 5825
rect 2219 5806 2249 5822
rect 2191 5790 2265 5806
rect 2191 5788 2204 5790
rect 2219 5788 2253 5790
rect 1856 5766 1869 5768
rect 1884 5766 1918 5768
rect 1856 5750 1918 5766
rect 1962 5761 1976 5764
rect 2040 5761 2070 5772
rect 2118 5768 2164 5784
rect 2191 5772 2265 5788
rect 2118 5766 2152 5768
rect 2117 5750 2164 5766
rect 2191 5750 2204 5772
rect 2219 5750 2249 5772
rect 2276 5750 2277 5766
rect 2292 5750 2305 5910
rect 2335 5806 2348 5910
rect 2393 5888 2394 5898
rect 2409 5888 2422 5898
rect 2393 5884 2422 5888
rect 2427 5884 2457 5910
rect 2475 5896 2491 5898
rect 2563 5896 2616 5910
rect 2564 5894 2628 5896
rect 2671 5894 2686 5910
rect 2735 5907 2765 5910
rect 2735 5904 2771 5907
rect 2701 5896 2717 5898
rect 2475 5884 2490 5888
rect 2393 5882 2490 5884
rect 2518 5882 2686 5894
rect 2702 5884 2717 5888
rect 2735 5885 2774 5904
rect 2793 5898 2800 5899
rect 2799 5891 2800 5898
rect 2783 5888 2784 5891
rect 2799 5888 2812 5891
rect 2735 5884 2765 5885
rect 2774 5884 2780 5885
rect 2783 5884 2812 5888
rect 2702 5883 2812 5884
rect 2702 5882 2818 5883
rect 2377 5874 2428 5882
rect 2377 5862 2402 5874
rect 2409 5862 2428 5874
rect 2459 5874 2509 5882
rect 2459 5866 2475 5874
rect 2482 5872 2509 5874
rect 2518 5872 2739 5882
rect 2482 5862 2739 5872
rect 2768 5874 2818 5882
rect 2768 5865 2784 5874
rect 2377 5854 2428 5862
rect 2475 5854 2739 5862
rect 2765 5862 2784 5865
rect 2791 5862 2818 5874
rect 2765 5854 2818 5862
rect 2393 5846 2394 5854
rect 2409 5846 2422 5854
rect 2393 5838 2409 5846
rect 2390 5831 2409 5834
rect 2390 5822 2412 5831
rect 2363 5812 2412 5822
rect 2363 5806 2393 5812
rect 2412 5807 2417 5812
rect 2335 5790 2409 5806
rect 2427 5798 2457 5854
rect 2492 5844 2700 5854
rect 2735 5850 2780 5854
rect 2783 5853 2784 5854
rect 2799 5853 2812 5854
rect 2518 5814 2707 5844
rect 2533 5811 2707 5814
rect 2526 5808 2707 5811
rect 2335 5788 2348 5790
rect 2363 5788 2397 5790
rect 2335 5772 2409 5788
rect 2436 5784 2449 5798
rect 2464 5784 2480 5800
rect 2526 5795 2537 5808
rect 2319 5750 2320 5766
rect 2335 5750 2348 5772
rect 2363 5750 2393 5772
rect 2436 5768 2498 5784
rect 2526 5777 2537 5793
rect 2542 5788 2552 5808
rect 2562 5788 2576 5808
rect 2579 5795 2588 5808
rect 2604 5795 2613 5808
rect 2542 5777 2576 5788
rect 2579 5777 2588 5793
rect 2604 5777 2613 5793
rect 2620 5788 2630 5808
rect 2640 5788 2654 5808
rect 2655 5795 2666 5808
rect 2620 5777 2654 5788
rect 2655 5777 2666 5793
rect 2712 5784 2728 5800
rect 2735 5798 2765 5850
rect 2799 5846 2800 5853
rect 2784 5838 2800 5846
rect 2771 5806 2784 5825
rect 2799 5806 2829 5822
rect 2771 5790 2845 5806
rect 2771 5788 2784 5790
rect 2799 5788 2833 5790
rect 2436 5766 2449 5768
rect 2464 5766 2498 5768
rect 2436 5750 2498 5766
rect 2542 5761 2558 5764
rect 2620 5761 2650 5772
rect 2698 5768 2744 5784
rect 2771 5772 2845 5788
rect 2698 5766 2732 5768
rect 2697 5750 2744 5766
rect 2771 5750 2784 5772
rect 2799 5750 2829 5772
rect 2856 5750 2857 5766
rect 2872 5750 2885 5910
rect 2915 5806 2928 5910
rect 2973 5888 2974 5898
rect 2989 5888 3002 5898
rect 2973 5884 3002 5888
rect 3007 5884 3037 5910
rect 3055 5896 3071 5898
rect 3143 5896 3196 5910
rect 3144 5894 3208 5896
rect 3251 5894 3266 5910
rect 3315 5907 3345 5910
rect 3315 5904 3351 5907
rect 3281 5896 3297 5898
rect 3055 5884 3070 5888
rect 2973 5882 3070 5884
rect 3098 5882 3266 5894
rect 3282 5884 3297 5888
rect 3315 5885 3354 5904
rect 3373 5898 3380 5899
rect 3379 5891 3380 5898
rect 3363 5888 3364 5891
rect 3379 5888 3392 5891
rect 3315 5884 3345 5885
rect 3354 5884 3360 5885
rect 3363 5884 3392 5888
rect 3282 5883 3392 5884
rect 3282 5882 3398 5883
rect 2957 5874 3008 5882
rect 2957 5862 2982 5874
rect 2989 5862 3008 5874
rect 3039 5874 3089 5882
rect 3039 5866 3055 5874
rect 3062 5872 3089 5874
rect 3098 5872 3319 5882
rect 3062 5862 3319 5872
rect 3348 5874 3398 5882
rect 3348 5865 3364 5874
rect 2957 5854 3008 5862
rect 3055 5854 3319 5862
rect 3345 5862 3364 5865
rect 3371 5862 3398 5874
rect 3345 5854 3398 5862
rect 2973 5846 2974 5854
rect 2989 5846 3002 5854
rect 2973 5838 2989 5846
rect 2970 5831 2989 5834
rect 2970 5822 2992 5831
rect 2943 5812 2992 5822
rect 2943 5806 2973 5812
rect 2992 5807 2997 5812
rect 2915 5790 2989 5806
rect 3007 5798 3037 5854
rect 3072 5844 3280 5854
rect 3315 5850 3360 5854
rect 3363 5853 3364 5854
rect 3379 5853 3392 5854
rect 3098 5814 3287 5844
rect 3113 5811 3287 5814
rect 3106 5808 3287 5811
rect 2915 5788 2928 5790
rect 2943 5788 2977 5790
rect 2915 5772 2989 5788
rect 3016 5784 3029 5798
rect 3044 5784 3060 5800
rect 3106 5795 3117 5808
rect 2899 5750 2900 5766
rect 2915 5750 2928 5772
rect 2943 5750 2973 5772
rect 3016 5768 3078 5784
rect 3106 5777 3117 5793
rect 3122 5788 3132 5808
rect 3142 5788 3156 5808
rect 3159 5795 3168 5808
rect 3184 5795 3193 5808
rect 3122 5777 3156 5788
rect 3159 5777 3168 5793
rect 3184 5777 3193 5793
rect 3200 5788 3210 5808
rect 3220 5788 3234 5808
rect 3235 5795 3246 5808
rect 3200 5777 3234 5788
rect 3235 5777 3246 5793
rect 3292 5784 3308 5800
rect 3315 5798 3345 5850
rect 3379 5846 3380 5853
rect 3364 5838 3380 5846
rect 3351 5806 3364 5825
rect 3379 5806 3409 5822
rect 3351 5790 3425 5806
rect 3351 5788 3364 5790
rect 3379 5788 3413 5790
rect 3016 5766 3029 5768
rect 3044 5766 3078 5768
rect 3016 5750 3078 5766
rect 3122 5761 3138 5764
rect 3200 5761 3230 5772
rect 3278 5768 3324 5784
rect 3351 5772 3425 5788
rect 3278 5766 3312 5768
rect 3277 5750 3324 5766
rect 3351 5750 3364 5772
rect 3379 5750 3409 5772
rect 3436 5750 3437 5766
rect 3452 5750 3465 5910
rect 3495 5806 3508 5910
rect 3553 5888 3554 5898
rect 3569 5888 3582 5898
rect 3553 5884 3582 5888
rect 3587 5884 3617 5910
rect 3635 5896 3651 5898
rect 3723 5896 3776 5910
rect 3724 5894 3788 5896
rect 3831 5894 3846 5910
rect 3895 5907 3925 5910
rect 3895 5904 3931 5907
rect 3861 5896 3877 5898
rect 3635 5884 3650 5888
rect 3553 5882 3650 5884
rect 3678 5882 3846 5894
rect 3862 5884 3877 5888
rect 3895 5885 3934 5904
rect 3953 5898 3960 5899
rect 3959 5891 3960 5898
rect 3943 5888 3944 5891
rect 3959 5888 3972 5891
rect 3895 5884 3925 5885
rect 3934 5884 3940 5885
rect 3943 5884 3972 5888
rect 3862 5883 3972 5884
rect 3862 5882 3978 5883
rect 3537 5874 3588 5882
rect 3537 5862 3562 5874
rect 3569 5862 3588 5874
rect 3619 5874 3669 5882
rect 3619 5866 3635 5874
rect 3642 5872 3669 5874
rect 3678 5872 3899 5882
rect 3642 5862 3899 5872
rect 3928 5874 3978 5882
rect 3928 5865 3944 5874
rect 3537 5854 3588 5862
rect 3635 5854 3899 5862
rect 3925 5862 3944 5865
rect 3951 5862 3978 5874
rect 3925 5854 3978 5862
rect 3553 5846 3554 5854
rect 3569 5846 3582 5854
rect 3553 5838 3569 5846
rect 3550 5831 3569 5834
rect 3550 5822 3572 5831
rect 3523 5812 3572 5822
rect 3523 5806 3553 5812
rect 3572 5807 3577 5812
rect 3495 5790 3569 5806
rect 3587 5798 3617 5854
rect 3652 5844 3860 5854
rect 3895 5850 3940 5854
rect 3943 5853 3944 5854
rect 3959 5853 3972 5854
rect 3678 5814 3867 5844
rect 3693 5811 3867 5814
rect 3686 5808 3867 5811
rect 3495 5788 3508 5790
rect 3523 5788 3557 5790
rect 3495 5772 3569 5788
rect 3596 5784 3609 5798
rect 3624 5784 3640 5800
rect 3686 5795 3697 5808
rect 3479 5750 3480 5766
rect 3495 5750 3508 5772
rect 3523 5750 3553 5772
rect 3596 5768 3658 5784
rect 3686 5777 3697 5793
rect 3702 5788 3712 5808
rect 3722 5788 3736 5808
rect 3739 5795 3748 5808
rect 3764 5795 3773 5808
rect 3702 5777 3736 5788
rect 3739 5777 3748 5793
rect 3764 5777 3773 5793
rect 3780 5788 3790 5808
rect 3800 5788 3814 5808
rect 3815 5795 3826 5808
rect 3780 5777 3814 5788
rect 3815 5777 3826 5793
rect 3872 5784 3888 5800
rect 3895 5798 3925 5850
rect 3959 5846 3960 5853
rect 3944 5838 3960 5846
rect 3931 5806 3944 5825
rect 3959 5806 3989 5822
rect 3931 5790 4005 5806
rect 3931 5788 3944 5790
rect 3959 5788 3993 5790
rect 3596 5766 3609 5768
rect 3624 5766 3658 5768
rect 3596 5750 3658 5766
rect 3702 5761 3718 5764
rect 3780 5761 3810 5772
rect 3858 5768 3904 5784
rect 3931 5772 4005 5788
rect 3858 5766 3892 5768
rect 3857 5750 3904 5766
rect 3931 5750 3944 5772
rect 3959 5750 3989 5772
rect 4016 5750 4017 5766
rect 4032 5750 4045 5910
rect 4075 5806 4088 5910
rect 4133 5888 4134 5898
rect 4149 5888 4162 5898
rect 4133 5884 4162 5888
rect 4167 5884 4197 5910
rect 4215 5896 4231 5898
rect 4303 5896 4356 5910
rect 4304 5894 4368 5896
rect 4411 5894 4426 5910
rect 4475 5907 4505 5910
rect 4475 5904 4511 5907
rect 4441 5896 4457 5898
rect 4215 5884 4230 5888
rect 4133 5882 4230 5884
rect 4258 5882 4426 5894
rect 4442 5884 4457 5888
rect 4475 5885 4514 5904
rect 4533 5898 4540 5899
rect 4539 5891 4540 5898
rect 4523 5888 4524 5891
rect 4539 5888 4552 5891
rect 4475 5884 4505 5885
rect 4514 5884 4520 5885
rect 4523 5884 4552 5888
rect 4442 5883 4552 5884
rect 4442 5882 4558 5883
rect 4117 5874 4168 5882
rect 4117 5862 4142 5874
rect 4149 5862 4168 5874
rect 4199 5874 4249 5882
rect 4199 5866 4215 5874
rect 4222 5872 4249 5874
rect 4258 5872 4479 5882
rect 4222 5862 4479 5872
rect 4508 5874 4558 5882
rect 4508 5865 4524 5874
rect 4117 5854 4168 5862
rect 4215 5854 4479 5862
rect 4505 5862 4524 5865
rect 4531 5862 4558 5874
rect 4505 5854 4558 5862
rect 4133 5846 4134 5854
rect 4149 5846 4162 5854
rect 4133 5838 4149 5846
rect 4130 5831 4149 5834
rect 4130 5822 4152 5831
rect 4103 5812 4152 5822
rect 4103 5806 4133 5812
rect 4152 5807 4157 5812
rect 4075 5790 4149 5806
rect 4167 5798 4197 5854
rect 4232 5844 4440 5854
rect 4475 5850 4520 5854
rect 4523 5853 4524 5854
rect 4539 5853 4552 5854
rect 4258 5814 4447 5844
rect 4273 5811 4447 5814
rect 4266 5808 4447 5811
rect 4075 5788 4088 5790
rect 4103 5788 4137 5790
rect 4075 5772 4149 5788
rect 4176 5784 4189 5798
rect 4204 5784 4220 5800
rect 4266 5795 4277 5808
rect 4059 5750 4060 5766
rect 4075 5750 4088 5772
rect 4103 5750 4133 5772
rect 4176 5768 4238 5784
rect 4266 5777 4277 5793
rect 4282 5788 4292 5808
rect 4302 5788 4316 5808
rect 4319 5795 4328 5808
rect 4344 5795 4353 5808
rect 4282 5777 4316 5788
rect 4319 5777 4328 5793
rect 4344 5777 4353 5793
rect 4360 5788 4370 5808
rect 4380 5788 4394 5808
rect 4395 5795 4406 5808
rect 4360 5777 4394 5788
rect 4395 5777 4406 5793
rect 4452 5784 4468 5800
rect 4475 5798 4505 5850
rect 4539 5846 4540 5853
rect 4524 5838 4540 5846
rect 4511 5806 4524 5825
rect 4539 5806 4569 5822
rect 4511 5790 4585 5806
rect 4511 5788 4524 5790
rect 4539 5788 4573 5790
rect 4176 5766 4189 5768
rect 4204 5766 4238 5768
rect 4176 5750 4238 5766
rect 4282 5761 4298 5764
rect 4360 5761 4390 5772
rect 4438 5768 4484 5784
rect 4511 5772 4585 5788
rect 4438 5766 4472 5768
rect 4437 5750 4484 5766
rect 4511 5750 4524 5772
rect 4539 5750 4569 5772
rect 4596 5750 4597 5766
rect 4612 5750 4625 5910
rect 4655 5806 4668 5910
rect 4713 5888 4714 5898
rect 4729 5888 4742 5898
rect 4713 5884 4742 5888
rect 4747 5884 4777 5910
rect 4795 5896 4811 5898
rect 4883 5896 4936 5910
rect 4884 5894 4948 5896
rect 4991 5894 5006 5910
rect 5055 5907 5085 5910
rect 5055 5904 5091 5907
rect 5021 5896 5037 5898
rect 4795 5884 4810 5888
rect 4713 5882 4810 5884
rect 4838 5882 5006 5894
rect 5022 5884 5037 5888
rect 5055 5885 5094 5904
rect 5113 5898 5120 5899
rect 5119 5891 5120 5898
rect 5103 5888 5104 5891
rect 5119 5888 5132 5891
rect 5055 5884 5085 5885
rect 5094 5884 5100 5885
rect 5103 5884 5132 5888
rect 5022 5883 5132 5884
rect 5022 5882 5138 5883
rect 4697 5874 4748 5882
rect 4697 5862 4722 5874
rect 4729 5862 4748 5874
rect 4779 5874 4829 5882
rect 4779 5866 4795 5874
rect 4802 5872 4829 5874
rect 4838 5872 5059 5882
rect 4802 5862 5059 5872
rect 5088 5874 5138 5882
rect 5088 5865 5104 5874
rect 4697 5854 4748 5862
rect 4795 5854 5059 5862
rect 5085 5862 5104 5865
rect 5111 5862 5138 5874
rect 5085 5854 5138 5862
rect 4713 5846 4714 5854
rect 4729 5846 4742 5854
rect 4713 5838 4729 5846
rect 4710 5831 4729 5834
rect 4710 5822 4732 5831
rect 4683 5812 4732 5822
rect 4683 5806 4713 5812
rect 4732 5807 4737 5812
rect 4655 5790 4729 5806
rect 4747 5798 4777 5854
rect 4812 5844 5020 5854
rect 5055 5850 5100 5854
rect 5103 5853 5104 5854
rect 5119 5853 5132 5854
rect 4838 5814 5027 5844
rect 4853 5811 5027 5814
rect 4846 5808 5027 5811
rect 4655 5788 4668 5790
rect 4683 5788 4717 5790
rect 4655 5772 4729 5788
rect 4756 5784 4769 5798
rect 4784 5784 4800 5800
rect 4846 5795 4857 5808
rect 4639 5750 4640 5766
rect 4655 5750 4668 5772
rect 4683 5750 4713 5772
rect 4756 5768 4818 5784
rect 4846 5777 4857 5793
rect 4862 5788 4872 5808
rect 4882 5788 4896 5808
rect 4899 5795 4908 5808
rect 4924 5795 4933 5808
rect 4862 5777 4896 5788
rect 4899 5777 4908 5793
rect 4924 5777 4933 5793
rect 4940 5788 4950 5808
rect 4960 5788 4974 5808
rect 4975 5795 4986 5808
rect 4940 5777 4974 5788
rect 4975 5777 4986 5793
rect 5032 5784 5048 5800
rect 5055 5798 5085 5850
rect 5119 5846 5120 5853
rect 5104 5838 5120 5846
rect 5091 5806 5104 5825
rect 5119 5806 5149 5822
rect 5091 5790 5165 5806
rect 5091 5788 5104 5790
rect 5119 5788 5153 5790
rect 4756 5766 4769 5768
rect 4784 5766 4818 5768
rect 4756 5750 4818 5766
rect 4862 5761 4878 5764
rect 4940 5761 4970 5772
rect 5018 5768 5064 5784
rect 5091 5772 5165 5788
rect 5018 5766 5052 5768
rect 5017 5750 5064 5766
rect 5091 5750 5104 5772
rect 5119 5750 5149 5772
rect 5176 5750 5177 5766
rect 5192 5750 5205 5910
rect 5235 5806 5248 5910
rect 5293 5888 5294 5898
rect 5309 5888 5322 5898
rect 5293 5884 5322 5888
rect 5327 5884 5357 5910
rect 5375 5896 5391 5898
rect 5463 5896 5516 5910
rect 5464 5894 5528 5896
rect 5571 5894 5586 5910
rect 5635 5907 5665 5910
rect 5635 5904 5671 5907
rect 5601 5896 5617 5898
rect 5375 5884 5390 5888
rect 5293 5882 5390 5884
rect 5418 5882 5586 5894
rect 5602 5884 5617 5888
rect 5635 5885 5674 5904
rect 5693 5898 5700 5899
rect 5699 5891 5700 5898
rect 5683 5888 5684 5891
rect 5699 5888 5712 5891
rect 5635 5884 5665 5885
rect 5674 5884 5680 5885
rect 5683 5884 5712 5888
rect 5602 5883 5712 5884
rect 5602 5882 5718 5883
rect 5277 5874 5328 5882
rect 5277 5862 5302 5874
rect 5309 5862 5328 5874
rect 5359 5874 5409 5882
rect 5359 5866 5375 5874
rect 5382 5872 5409 5874
rect 5418 5872 5639 5882
rect 5382 5862 5639 5872
rect 5668 5874 5718 5882
rect 5668 5865 5684 5874
rect 5277 5854 5328 5862
rect 5375 5854 5639 5862
rect 5665 5862 5684 5865
rect 5691 5862 5718 5874
rect 5665 5854 5718 5862
rect 5293 5846 5294 5854
rect 5309 5846 5322 5854
rect 5293 5838 5309 5846
rect 5290 5831 5309 5834
rect 5290 5822 5312 5831
rect 5263 5812 5312 5822
rect 5263 5806 5293 5812
rect 5312 5807 5317 5812
rect 5235 5790 5309 5806
rect 5327 5798 5357 5854
rect 5392 5844 5600 5854
rect 5635 5850 5680 5854
rect 5683 5853 5684 5854
rect 5699 5853 5712 5854
rect 5418 5814 5607 5844
rect 5433 5811 5607 5814
rect 5426 5808 5607 5811
rect 5235 5788 5248 5790
rect 5263 5788 5297 5790
rect 5235 5772 5309 5788
rect 5336 5784 5349 5798
rect 5364 5784 5380 5800
rect 5426 5795 5437 5808
rect 5219 5750 5220 5766
rect 5235 5750 5248 5772
rect 5263 5750 5293 5772
rect 5336 5768 5398 5784
rect 5426 5777 5437 5793
rect 5442 5788 5452 5808
rect 5462 5788 5476 5808
rect 5479 5795 5488 5808
rect 5504 5795 5513 5808
rect 5442 5777 5476 5788
rect 5479 5777 5488 5793
rect 5504 5777 5513 5793
rect 5520 5788 5530 5808
rect 5540 5788 5554 5808
rect 5555 5795 5566 5808
rect 5520 5777 5554 5788
rect 5555 5777 5566 5793
rect 5612 5784 5628 5800
rect 5635 5798 5665 5850
rect 5699 5846 5700 5853
rect 5684 5838 5700 5846
rect 5671 5806 5684 5825
rect 5699 5806 5729 5822
rect 5671 5790 5745 5806
rect 5671 5788 5684 5790
rect 5699 5788 5733 5790
rect 5336 5766 5349 5768
rect 5364 5766 5398 5768
rect 5336 5750 5398 5766
rect 5442 5761 5458 5764
rect 5520 5761 5550 5772
rect 5598 5768 5644 5784
rect 5671 5772 5745 5788
rect 5598 5766 5632 5768
rect 5597 5750 5644 5766
rect 5671 5750 5684 5772
rect 5699 5750 5729 5772
rect 5756 5750 5757 5766
rect 5772 5750 5785 5910
rect 5815 5806 5828 5910
rect 5873 5888 5874 5898
rect 5889 5888 5902 5898
rect 5873 5884 5902 5888
rect 5907 5884 5937 5910
rect 5955 5896 5971 5898
rect 6043 5896 6096 5910
rect 6044 5894 6108 5896
rect 6151 5894 6166 5910
rect 6215 5907 6245 5910
rect 6215 5904 6251 5907
rect 6181 5896 6197 5898
rect 5955 5884 5970 5888
rect 5873 5882 5970 5884
rect 5998 5882 6166 5894
rect 6182 5884 6197 5888
rect 6215 5885 6254 5904
rect 6273 5898 6280 5899
rect 6279 5891 6280 5898
rect 6263 5888 6264 5891
rect 6279 5888 6292 5891
rect 6215 5884 6245 5885
rect 6254 5884 6260 5885
rect 6263 5884 6292 5888
rect 6182 5883 6292 5884
rect 6182 5882 6298 5883
rect 5857 5874 5908 5882
rect 5857 5862 5882 5874
rect 5889 5862 5908 5874
rect 5939 5874 5989 5882
rect 5939 5866 5955 5874
rect 5962 5872 5989 5874
rect 5998 5872 6219 5882
rect 5962 5862 6219 5872
rect 6248 5874 6298 5882
rect 6248 5865 6264 5874
rect 5857 5854 5908 5862
rect 5955 5854 6219 5862
rect 6245 5862 6264 5865
rect 6271 5862 6298 5874
rect 6245 5854 6298 5862
rect 5873 5846 5874 5854
rect 5889 5846 5902 5854
rect 5873 5838 5889 5846
rect 5870 5831 5889 5834
rect 5870 5822 5892 5831
rect 5843 5812 5892 5822
rect 5843 5806 5873 5812
rect 5892 5807 5897 5812
rect 5815 5790 5889 5806
rect 5907 5798 5937 5854
rect 5972 5844 6180 5854
rect 6215 5850 6260 5854
rect 6263 5853 6264 5854
rect 6279 5853 6292 5854
rect 5998 5814 6187 5844
rect 6013 5811 6187 5814
rect 6006 5808 6187 5811
rect 5815 5788 5828 5790
rect 5843 5788 5877 5790
rect 5815 5772 5889 5788
rect 5916 5784 5929 5798
rect 5944 5784 5960 5800
rect 6006 5795 6017 5808
rect 5799 5750 5800 5766
rect 5815 5750 5828 5772
rect 5843 5750 5873 5772
rect 5916 5768 5978 5784
rect 6006 5777 6017 5793
rect 6022 5788 6032 5808
rect 6042 5788 6056 5808
rect 6059 5795 6068 5808
rect 6084 5795 6093 5808
rect 6022 5777 6056 5788
rect 6059 5777 6068 5793
rect 6084 5777 6093 5793
rect 6100 5788 6110 5808
rect 6120 5788 6134 5808
rect 6135 5795 6146 5808
rect 6100 5777 6134 5788
rect 6135 5777 6146 5793
rect 6192 5784 6208 5800
rect 6215 5798 6245 5850
rect 6279 5846 6280 5853
rect 6264 5838 6280 5846
rect 6251 5806 6264 5825
rect 6279 5806 6309 5822
rect 6251 5790 6325 5806
rect 6251 5788 6264 5790
rect 6279 5788 6313 5790
rect 5916 5766 5929 5768
rect 5944 5766 5978 5768
rect 5916 5750 5978 5766
rect 6022 5761 6038 5764
rect 6100 5761 6130 5772
rect 6178 5768 6224 5784
rect 6251 5772 6325 5788
rect 6178 5766 6212 5768
rect 6177 5750 6224 5766
rect 6251 5750 6264 5772
rect 6279 5750 6309 5772
rect 6336 5750 6337 5766
rect 6352 5750 6365 5910
rect 6395 5806 6408 5910
rect 6453 5888 6454 5898
rect 6469 5888 6482 5898
rect 6453 5884 6482 5888
rect 6487 5884 6517 5910
rect 6535 5896 6551 5898
rect 6623 5896 6676 5910
rect 6624 5894 6688 5896
rect 6731 5894 6746 5910
rect 6795 5907 6825 5910
rect 6795 5904 6831 5907
rect 6761 5896 6777 5898
rect 6535 5884 6550 5888
rect 6453 5882 6550 5884
rect 6578 5882 6746 5894
rect 6762 5884 6777 5888
rect 6795 5885 6834 5904
rect 6853 5898 6860 5899
rect 6859 5891 6860 5898
rect 6843 5888 6844 5891
rect 6859 5888 6872 5891
rect 6795 5884 6825 5885
rect 6834 5884 6840 5885
rect 6843 5884 6872 5888
rect 6762 5883 6872 5884
rect 6762 5882 6878 5883
rect 6437 5874 6488 5882
rect 6437 5862 6462 5874
rect 6469 5862 6488 5874
rect 6519 5874 6569 5882
rect 6519 5866 6535 5874
rect 6542 5872 6569 5874
rect 6578 5872 6799 5882
rect 6542 5862 6799 5872
rect 6828 5874 6878 5882
rect 6828 5865 6844 5874
rect 6437 5854 6488 5862
rect 6535 5854 6799 5862
rect 6825 5862 6844 5865
rect 6851 5862 6878 5874
rect 6825 5854 6878 5862
rect 6453 5846 6454 5854
rect 6469 5846 6482 5854
rect 6453 5838 6469 5846
rect 6450 5831 6469 5834
rect 6450 5822 6472 5831
rect 6423 5812 6472 5822
rect 6423 5806 6453 5812
rect 6472 5807 6477 5812
rect 6395 5790 6469 5806
rect 6487 5798 6517 5854
rect 6552 5844 6760 5854
rect 6795 5850 6840 5854
rect 6843 5853 6844 5854
rect 6859 5853 6872 5854
rect 6578 5814 6767 5844
rect 6593 5811 6767 5814
rect 6586 5808 6767 5811
rect 6395 5788 6408 5790
rect 6423 5788 6457 5790
rect 6395 5772 6469 5788
rect 6496 5784 6509 5798
rect 6524 5784 6540 5800
rect 6586 5795 6597 5808
rect 6379 5750 6380 5766
rect 6395 5750 6408 5772
rect 6423 5750 6453 5772
rect 6496 5768 6558 5784
rect 6586 5777 6597 5793
rect 6602 5788 6612 5808
rect 6622 5788 6636 5808
rect 6639 5795 6648 5808
rect 6664 5795 6673 5808
rect 6602 5777 6636 5788
rect 6639 5777 6648 5793
rect 6664 5777 6673 5793
rect 6680 5788 6690 5808
rect 6700 5788 6714 5808
rect 6715 5795 6726 5808
rect 6680 5777 6714 5788
rect 6715 5777 6726 5793
rect 6772 5784 6788 5800
rect 6795 5798 6825 5850
rect 6859 5846 6860 5853
rect 6844 5838 6860 5846
rect 6831 5806 6844 5825
rect 6859 5806 6889 5822
rect 6831 5790 6905 5806
rect 6831 5788 6844 5790
rect 6859 5788 6893 5790
rect 6496 5766 6509 5768
rect 6524 5766 6558 5768
rect 6496 5750 6558 5766
rect 6602 5761 6618 5764
rect 6680 5761 6710 5772
rect 6758 5768 6804 5784
rect 6831 5772 6905 5788
rect 6758 5766 6792 5768
rect 6757 5750 6804 5766
rect 6831 5750 6844 5772
rect 6859 5750 6889 5772
rect 6916 5750 6917 5766
rect 6932 5750 6945 5910
rect 6975 5806 6988 5910
rect 7033 5888 7034 5898
rect 7049 5888 7062 5898
rect 7033 5884 7062 5888
rect 7067 5884 7097 5910
rect 7115 5896 7131 5898
rect 7203 5896 7256 5910
rect 7204 5894 7268 5896
rect 7311 5894 7326 5910
rect 7375 5907 7405 5910
rect 7375 5904 7411 5907
rect 7341 5896 7357 5898
rect 7115 5884 7130 5888
rect 7033 5882 7130 5884
rect 7158 5882 7326 5894
rect 7342 5884 7357 5888
rect 7375 5885 7414 5904
rect 7433 5898 7440 5899
rect 7439 5891 7440 5898
rect 7423 5888 7424 5891
rect 7439 5888 7452 5891
rect 7375 5884 7405 5885
rect 7414 5884 7420 5885
rect 7423 5884 7452 5888
rect 7342 5883 7452 5884
rect 7342 5882 7458 5883
rect 7017 5874 7068 5882
rect 7017 5862 7042 5874
rect 7049 5862 7068 5874
rect 7099 5874 7149 5882
rect 7099 5866 7115 5874
rect 7122 5872 7149 5874
rect 7158 5872 7379 5882
rect 7122 5862 7379 5872
rect 7408 5874 7458 5882
rect 7408 5865 7424 5874
rect 7017 5854 7068 5862
rect 7115 5854 7379 5862
rect 7405 5862 7424 5865
rect 7431 5862 7458 5874
rect 7405 5854 7458 5862
rect 7033 5846 7034 5854
rect 7049 5846 7062 5854
rect 7033 5838 7049 5846
rect 7030 5831 7049 5834
rect 7030 5822 7052 5831
rect 7003 5812 7052 5822
rect 7003 5806 7033 5812
rect 7052 5807 7057 5812
rect 6975 5790 7049 5806
rect 7067 5798 7097 5854
rect 7132 5844 7340 5854
rect 7375 5850 7420 5854
rect 7423 5853 7424 5854
rect 7439 5853 7452 5854
rect 7158 5814 7347 5844
rect 7173 5811 7347 5814
rect 7166 5808 7347 5811
rect 6975 5788 6988 5790
rect 7003 5788 7037 5790
rect 6975 5772 7049 5788
rect 7076 5784 7089 5798
rect 7104 5784 7120 5800
rect 7166 5795 7177 5808
rect 6959 5750 6960 5766
rect 6975 5750 6988 5772
rect 7003 5750 7033 5772
rect 7076 5768 7138 5784
rect 7166 5777 7177 5793
rect 7182 5788 7192 5808
rect 7202 5788 7216 5808
rect 7219 5795 7228 5808
rect 7244 5795 7253 5808
rect 7182 5777 7216 5788
rect 7219 5777 7228 5793
rect 7244 5777 7253 5793
rect 7260 5788 7270 5808
rect 7280 5788 7294 5808
rect 7295 5795 7306 5808
rect 7260 5777 7294 5788
rect 7295 5777 7306 5793
rect 7352 5784 7368 5800
rect 7375 5798 7405 5850
rect 7439 5846 7440 5853
rect 7424 5838 7440 5846
rect 7411 5806 7424 5825
rect 7439 5806 7469 5822
rect 7411 5790 7485 5806
rect 7411 5788 7424 5790
rect 7439 5788 7473 5790
rect 7076 5766 7089 5768
rect 7104 5766 7138 5768
rect 7076 5750 7138 5766
rect 7182 5761 7198 5764
rect 7260 5761 7290 5772
rect 7338 5768 7384 5784
rect 7411 5772 7485 5788
rect 7338 5766 7372 5768
rect 7337 5750 7384 5766
rect 7411 5750 7424 5772
rect 7439 5750 7469 5772
rect 7496 5750 7497 5766
rect 7512 5750 7525 5910
rect 7555 5806 7568 5910
rect 7613 5888 7614 5898
rect 7629 5888 7642 5898
rect 7613 5884 7642 5888
rect 7647 5884 7677 5910
rect 7695 5896 7711 5898
rect 7783 5896 7836 5910
rect 7784 5894 7848 5896
rect 7891 5894 7906 5910
rect 7955 5907 7985 5910
rect 7955 5904 7991 5907
rect 7921 5896 7937 5898
rect 7695 5884 7710 5888
rect 7613 5882 7710 5884
rect 7738 5882 7906 5894
rect 7922 5884 7937 5888
rect 7955 5885 7994 5904
rect 8013 5898 8020 5899
rect 8019 5891 8020 5898
rect 8003 5888 8004 5891
rect 8019 5888 8032 5891
rect 7955 5884 7985 5885
rect 7994 5884 8000 5885
rect 8003 5884 8032 5888
rect 7922 5883 8032 5884
rect 7922 5882 8038 5883
rect 7597 5874 7648 5882
rect 7597 5862 7622 5874
rect 7629 5862 7648 5874
rect 7679 5874 7729 5882
rect 7679 5866 7695 5874
rect 7702 5872 7729 5874
rect 7738 5872 7959 5882
rect 7702 5862 7959 5872
rect 7988 5874 8038 5882
rect 7988 5865 8004 5874
rect 7597 5854 7648 5862
rect 7695 5854 7959 5862
rect 7985 5862 8004 5865
rect 8011 5862 8038 5874
rect 7985 5854 8038 5862
rect 7613 5846 7614 5854
rect 7629 5846 7642 5854
rect 7613 5838 7629 5846
rect 7610 5831 7629 5834
rect 7610 5822 7632 5831
rect 7583 5812 7632 5822
rect 7583 5806 7613 5812
rect 7632 5807 7637 5812
rect 7555 5790 7629 5806
rect 7647 5798 7677 5854
rect 7712 5844 7920 5854
rect 7955 5850 8000 5854
rect 8003 5853 8004 5854
rect 8019 5853 8032 5854
rect 7738 5814 7927 5844
rect 7753 5811 7927 5814
rect 7746 5808 7927 5811
rect 7555 5788 7568 5790
rect 7583 5788 7617 5790
rect 7555 5772 7629 5788
rect 7656 5784 7669 5798
rect 7684 5784 7700 5800
rect 7746 5795 7757 5808
rect 7539 5750 7540 5766
rect 7555 5750 7568 5772
rect 7583 5750 7613 5772
rect 7656 5768 7718 5784
rect 7746 5777 7757 5793
rect 7762 5788 7772 5808
rect 7782 5788 7796 5808
rect 7799 5795 7808 5808
rect 7824 5795 7833 5808
rect 7762 5777 7796 5788
rect 7799 5777 7808 5793
rect 7824 5777 7833 5793
rect 7840 5788 7850 5808
rect 7860 5788 7874 5808
rect 7875 5795 7886 5808
rect 7840 5777 7874 5788
rect 7875 5777 7886 5793
rect 7932 5784 7948 5800
rect 7955 5798 7985 5850
rect 8019 5846 8020 5853
rect 8004 5838 8020 5846
rect 7991 5806 8004 5825
rect 8019 5806 8049 5822
rect 7991 5790 8065 5806
rect 7991 5788 8004 5790
rect 8019 5788 8053 5790
rect 7656 5766 7669 5768
rect 7684 5766 7718 5768
rect 7656 5750 7718 5766
rect 7762 5761 7778 5764
rect 7840 5761 7870 5772
rect 7918 5768 7964 5784
rect 7991 5772 8065 5788
rect 7918 5766 7952 5768
rect 7917 5750 7964 5766
rect 7991 5750 8004 5772
rect 8019 5750 8049 5772
rect 8076 5750 8077 5766
rect 8092 5750 8105 5910
rect 8135 5806 8148 5910
rect 8193 5888 8194 5898
rect 8209 5888 8222 5898
rect 8193 5884 8222 5888
rect 8227 5884 8257 5910
rect 8275 5896 8291 5898
rect 8363 5896 8416 5910
rect 8364 5894 8428 5896
rect 8471 5894 8486 5910
rect 8535 5907 8565 5910
rect 8535 5904 8571 5907
rect 8501 5896 8517 5898
rect 8275 5884 8290 5888
rect 8193 5882 8290 5884
rect 8318 5882 8486 5894
rect 8502 5884 8517 5888
rect 8535 5885 8574 5904
rect 8593 5898 8600 5899
rect 8599 5891 8600 5898
rect 8583 5888 8584 5891
rect 8599 5888 8612 5891
rect 8535 5884 8565 5885
rect 8574 5884 8580 5885
rect 8583 5884 8612 5888
rect 8502 5883 8612 5884
rect 8502 5882 8618 5883
rect 8177 5874 8228 5882
rect 8177 5862 8202 5874
rect 8209 5862 8228 5874
rect 8259 5874 8309 5882
rect 8259 5866 8275 5874
rect 8282 5872 8309 5874
rect 8318 5872 8539 5882
rect 8282 5862 8539 5872
rect 8568 5874 8618 5882
rect 8568 5865 8584 5874
rect 8177 5854 8228 5862
rect 8275 5854 8539 5862
rect 8565 5862 8584 5865
rect 8591 5862 8618 5874
rect 8565 5854 8618 5862
rect 8193 5846 8194 5854
rect 8209 5846 8222 5854
rect 8193 5838 8209 5846
rect 8190 5831 8209 5834
rect 8190 5822 8212 5831
rect 8163 5812 8212 5822
rect 8163 5806 8193 5812
rect 8212 5807 8217 5812
rect 8135 5790 8209 5806
rect 8227 5798 8257 5854
rect 8292 5844 8500 5854
rect 8535 5850 8580 5854
rect 8583 5853 8584 5854
rect 8599 5853 8612 5854
rect 8318 5814 8507 5844
rect 8333 5811 8507 5814
rect 8326 5808 8507 5811
rect 8135 5788 8148 5790
rect 8163 5788 8197 5790
rect 8135 5772 8209 5788
rect 8236 5784 8249 5798
rect 8264 5784 8280 5800
rect 8326 5795 8337 5808
rect 8119 5750 8120 5766
rect 8135 5750 8148 5772
rect 8163 5750 8193 5772
rect 8236 5768 8298 5784
rect 8326 5777 8337 5793
rect 8342 5788 8352 5808
rect 8362 5788 8376 5808
rect 8379 5795 8388 5808
rect 8404 5795 8413 5808
rect 8342 5777 8376 5788
rect 8379 5777 8388 5793
rect 8404 5777 8413 5793
rect 8420 5788 8430 5808
rect 8440 5788 8454 5808
rect 8455 5795 8466 5808
rect 8420 5777 8454 5788
rect 8455 5777 8466 5793
rect 8512 5784 8528 5800
rect 8535 5798 8565 5850
rect 8599 5846 8600 5853
rect 8584 5838 8600 5846
rect 8571 5806 8584 5825
rect 8599 5806 8629 5822
rect 8571 5790 8645 5806
rect 8571 5788 8584 5790
rect 8599 5788 8633 5790
rect 8236 5766 8249 5768
rect 8264 5766 8298 5768
rect 8236 5750 8298 5766
rect 8342 5761 8358 5764
rect 8420 5761 8450 5772
rect 8498 5768 8544 5784
rect 8571 5772 8645 5788
rect 8498 5766 8532 5768
rect 8497 5750 8544 5766
rect 8571 5750 8584 5772
rect 8599 5750 8629 5772
rect 8656 5750 8657 5766
rect 8672 5750 8685 5910
rect 8715 5806 8728 5910
rect 8773 5888 8774 5898
rect 8789 5888 8802 5898
rect 8773 5884 8802 5888
rect 8807 5884 8837 5910
rect 8855 5896 8871 5898
rect 8943 5896 8996 5910
rect 8944 5894 9008 5896
rect 9051 5894 9066 5910
rect 9115 5907 9145 5910
rect 9115 5904 9151 5907
rect 9081 5896 9097 5898
rect 8855 5884 8870 5888
rect 8773 5882 8870 5884
rect 8898 5882 9066 5894
rect 9082 5884 9097 5888
rect 9115 5885 9154 5904
rect 9173 5898 9180 5899
rect 9179 5891 9180 5898
rect 9163 5888 9164 5891
rect 9179 5888 9192 5891
rect 9115 5884 9145 5885
rect 9154 5884 9160 5885
rect 9163 5884 9192 5888
rect 9082 5883 9192 5884
rect 9082 5882 9198 5883
rect 8757 5874 8808 5882
rect 8757 5862 8782 5874
rect 8789 5862 8808 5874
rect 8839 5874 8889 5882
rect 8839 5866 8855 5874
rect 8862 5872 8889 5874
rect 8898 5872 9119 5882
rect 8862 5862 9119 5872
rect 9148 5874 9198 5882
rect 9148 5865 9164 5874
rect 8757 5854 8808 5862
rect 8855 5854 9119 5862
rect 9145 5862 9164 5865
rect 9171 5862 9198 5874
rect 9145 5854 9198 5862
rect 8773 5846 8774 5854
rect 8789 5846 8802 5854
rect 8773 5838 8789 5846
rect 8770 5831 8789 5834
rect 8770 5822 8792 5831
rect 8743 5812 8792 5822
rect 8743 5806 8773 5812
rect 8792 5807 8797 5812
rect 8715 5790 8789 5806
rect 8807 5798 8837 5854
rect 8872 5844 9080 5854
rect 9115 5850 9160 5854
rect 9163 5853 9164 5854
rect 9179 5853 9192 5854
rect 8898 5814 9087 5844
rect 8913 5811 9087 5814
rect 8906 5808 9087 5811
rect 8715 5788 8728 5790
rect 8743 5788 8777 5790
rect 8715 5772 8789 5788
rect 8816 5784 8829 5798
rect 8844 5784 8860 5800
rect 8906 5795 8917 5808
rect 8699 5750 8700 5766
rect 8715 5750 8728 5772
rect 8743 5750 8773 5772
rect 8816 5768 8878 5784
rect 8906 5777 8917 5793
rect 8922 5788 8932 5808
rect 8942 5788 8956 5808
rect 8959 5795 8968 5808
rect 8984 5795 8993 5808
rect 8922 5777 8956 5788
rect 8959 5777 8968 5793
rect 8984 5777 8993 5793
rect 9000 5788 9010 5808
rect 9020 5788 9034 5808
rect 9035 5795 9046 5808
rect 9000 5777 9034 5788
rect 9035 5777 9046 5793
rect 9092 5784 9108 5800
rect 9115 5798 9145 5850
rect 9179 5846 9180 5853
rect 9164 5838 9180 5846
rect 9151 5806 9164 5825
rect 9179 5806 9209 5822
rect 9151 5790 9225 5806
rect 9151 5788 9164 5790
rect 9179 5788 9213 5790
rect 8816 5766 8829 5768
rect 8844 5766 8878 5768
rect 8816 5750 8878 5766
rect 8922 5761 8938 5764
rect 9000 5761 9030 5772
rect 9078 5768 9124 5784
rect 9151 5772 9225 5788
rect 9078 5766 9112 5768
rect 9077 5750 9124 5766
rect 9151 5750 9164 5772
rect 9179 5750 9209 5772
rect 9236 5750 9237 5766
rect 9252 5750 9265 5910
rect -7 5742 34 5750
rect -7 5716 8 5742
rect 15 5716 34 5742
rect 98 5738 160 5750
rect 172 5738 247 5750
rect 305 5738 380 5750
rect 392 5738 423 5750
rect 429 5738 464 5750
rect 98 5736 260 5738
rect -7 5708 34 5716
rect 116 5712 129 5736
rect 144 5734 159 5736
rect -1 5698 0 5708
rect 15 5698 28 5708
rect 43 5698 73 5712
rect 116 5698 159 5712
rect 183 5709 190 5716
rect 193 5712 260 5736
rect 292 5736 464 5738
rect 262 5714 290 5718
rect 292 5714 372 5736
rect 393 5734 408 5736
rect 262 5712 372 5714
rect 193 5708 372 5712
rect 166 5698 196 5708
rect 198 5698 351 5708
rect 359 5698 389 5708
rect 393 5698 423 5712
rect 451 5698 464 5736
rect 536 5742 571 5750
rect 536 5716 537 5742
rect 544 5716 571 5742
rect 479 5698 509 5712
rect 536 5708 571 5716
rect 573 5742 614 5750
rect 573 5716 588 5742
rect 595 5716 614 5742
rect 678 5738 740 5750
rect 752 5738 827 5750
rect 885 5738 960 5750
rect 972 5738 1003 5750
rect 1009 5738 1044 5750
rect 678 5736 840 5738
rect 573 5708 614 5716
rect 696 5712 709 5736
rect 724 5734 739 5736
rect 536 5698 537 5708
rect 552 5698 565 5708
rect 579 5698 580 5708
rect 595 5698 608 5708
rect 623 5698 653 5712
rect 696 5698 739 5712
rect 763 5709 770 5716
rect 773 5712 840 5736
rect 872 5736 1044 5738
rect 842 5714 870 5718
rect 872 5714 952 5736
rect 973 5734 988 5736
rect 842 5712 952 5714
rect 773 5708 952 5712
rect 746 5698 776 5708
rect 778 5698 931 5708
rect 939 5698 969 5708
rect 973 5698 1003 5712
rect 1031 5698 1044 5736
rect 1116 5742 1151 5750
rect 1116 5716 1117 5742
rect 1124 5716 1151 5742
rect 1059 5698 1089 5712
rect 1116 5708 1151 5716
rect 1153 5742 1194 5750
rect 1153 5716 1168 5742
rect 1175 5716 1194 5742
rect 1258 5738 1320 5750
rect 1332 5738 1407 5750
rect 1465 5738 1540 5750
rect 1552 5738 1583 5750
rect 1589 5738 1624 5750
rect 1258 5736 1420 5738
rect 1153 5708 1194 5716
rect 1276 5712 1289 5736
rect 1304 5734 1319 5736
rect 1116 5698 1117 5708
rect 1132 5698 1145 5708
rect 1159 5698 1160 5708
rect 1175 5698 1188 5708
rect 1203 5698 1233 5712
rect 1276 5698 1319 5712
rect 1343 5709 1350 5716
rect 1353 5712 1420 5736
rect 1452 5736 1624 5738
rect 1422 5714 1450 5718
rect 1452 5714 1532 5736
rect 1553 5734 1568 5736
rect 1422 5712 1532 5714
rect 1353 5708 1532 5712
rect 1326 5698 1356 5708
rect 1358 5698 1511 5708
rect 1519 5698 1549 5708
rect 1553 5698 1583 5712
rect 1611 5698 1624 5736
rect 1696 5742 1731 5750
rect 1696 5716 1697 5742
rect 1704 5716 1731 5742
rect 1639 5698 1669 5712
rect 1696 5708 1731 5716
rect 1733 5742 1774 5750
rect 1733 5716 1748 5742
rect 1755 5716 1774 5742
rect 1838 5738 1900 5750
rect 1912 5738 1987 5750
rect 2045 5738 2120 5750
rect 2132 5738 2163 5750
rect 2169 5738 2204 5750
rect 1838 5736 2000 5738
rect 1733 5708 1774 5716
rect 1856 5712 1869 5736
rect 1884 5734 1899 5736
rect 1696 5698 1697 5708
rect 1712 5698 1725 5708
rect 1739 5698 1740 5708
rect 1755 5698 1768 5708
rect 1783 5698 1813 5712
rect 1856 5698 1899 5712
rect 1923 5709 1930 5716
rect 1933 5712 2000 5736
rect 2032 5736 2204 5738
rect 2002 5714 2030 5718
rect 2032 5714 2112 5736
rect 2133 5734 2148 5736
rect 2002 5712 2112 5714
rect 1933 5708 2112 5712
rect 1906 5698 1936 5708
rect 1938 5698 2091 5708
rect 2099 5698 2129 5708
rect 2133 5698 2163 5712
rect 2191 5698 2204 5736
rect 2276 5742 2311 5750
rect 2276 5716 2277 5742
rect 2284 5716 2311 5742
rect 2219 5698 2249 5712
rect 2276 5708 2311 5716
rect 2313 5742 2354 5750
rect 2313 5716 2328 5742
rect 2335 5716 2354 5742
rect 2418 5738 2480 5750
rect 2492 5738 2567 5750
rect 2625 5738 2700 5750
rect 2712 5738 2743 5750
rect 2749 5738 2784 5750
rect 2418 5736 2580 5738
rect 2313 5708 2354 5716
rect 2436 5712 2449 5736
rect 2464 5734 2479 5736
rect 2276 5698 2277 5708
rect 2292 5698 2305 5708
rect 2319 5698 2320 5708
rect 2335 5698 2348 5708
rect 2363 5698 2393 5712
rect 2436 5698 2479 5712
rect 2503 5709 2510 5716
rect 2513 5712 2580 5736
rect 2612 5736 2784 5738
rect 2582 5714 2610 5718
rect 2612 5714 2692 5736
rect 2713 5734 2728 5736
rect 2582 5712 2692 5714
rect 2513 5708 2692 5712
rect 2486 5698 2516 5708
rect 2518 5698 2671 5708
rect 2679 5698 2709 5708
rect 2713 5698 2743 5712
rect 2771 5698 2784 5736
rect 2856 5742 2891 5750
rect 2856 5716 2857 5742
rect 2864 5716 2891 5742
rect 2799 5698 2829 5712
rect 2856 5708 2891 5716
rect 2893 5742 2934 5750
rect 2893 5716 2908 5742
rect 2915 5716 2934 5742
rect 2998 5738 3060 5750
rect 3072 5738 3147 5750
rect 3205 5738 3280 5750
rect 3292 5738 3323 5750
rect 3329 5738 3364 5750
rect 2998 5736 3160 5738
rect 2893 5708 2934 5716
rect 3016 5712 3029 5736
rect 3044 5734 3059 5736
rect 2856 5698 2857 5708
rect 2872 5698 2885 5708
rect 2899 5698 2900 5708
rect 2915 5698 2928 5708
rect 2943 5698 2973 5712
rect 3016 5698 3059 5712
rect 3083 5709 3090 5716
rect 3093 5712 3160 5736
rect 3192 5736 3364 5738
rect 3162 5714 3190 5718
rect 3192 5714 3272 5736
rect 3293 5734 3308 5736
rect 3162 5712 3272 5714
rect 3093 5708 3272 5712
rect 3066 5698 3096 5708
rect 3098 5698 3251 5708
rect 3259 5698 3289 5708
rect 3293 5698 3323 5712
rect 3351 5698 3364 5736
rect 3436 5742 3471 5750
rect 3436 5716 3437 5742
rect 3444 5716 3471 5742
rect 3379 5698 3409 5712
rect 3436 5708 3471 5716
rect 3473 5742 3514 5750
rect 3473 5716 3488 5742
rect 3495 5716 3514 5742
rect 3578 5738 3640 5750
rect 3652 5738 3727 5750
rect 3785 5738 3860 5750
rect 3872 5738 3903 5750
rect 3909 5738 3944 5750
rect 3578 5736 3740 5738
rect 3473 5708 3514 5716
rect 3596 5712 3609 5736
rect 3624 5734 3639 5736
rect 3436 5698 3437 5708
rect 3452 5698 3465 5708
rect 3479 5698 3480 5708
rect 3495 5698 3508 5708
rect 3523 5698 3553 5712
rect 3596 5698 3639 5712
rect 3663 5709 3670 5716
rect 3673 5712 3740 5736
rect 3772 5736 3944 5738
rect 3742 5714 3770 5718
rect 3772 5714 3852 5736
rect 3873 5734 3888 5736
rect 3742 5712 3852 5714
rect 3673 5708 3852 5712
rect 3646 5698 3676 5708
rect 3678 5698 3831 5708
rect 3839 5698 3869 5708
rect 3873 5698 3903 5712
rect 3931 5698 3944 5736
rect 4016 5742 4051 5750
rect 4016 5716 4017 5742
rect 4024 5716 4051 5742
rect 3959 5698 3989 5712
rect 4016 5708 4051 5716
rect 4053 5742 4094 5750
rect 4053 5716 4068 5742
rect 4075 5716 4094 5742
rect 4158 5738 4220 5750
rect 4232 5738 4307 5750
rect 4365 5738 4440 5750
rect 4452 5738 4483 5750
rect 4489 5738 4524 5750
rect 4158 5736 4320 5738
rect 4053 5708 4094 5716
rect 4176 5712 4189 5736
rect 4204 5734 4219 5736
rect 4016 5698 4017 5708
rect 4032 5698 4045 5708
rect 4059 5698 4060 5708
rect 4075 5698 4088 5708
rect 4103 5698 4133 5712
rect 4176 5698 4219 5712
rect 4243 5709 4250 5716
rect 4253 5712 4320 5736
rect 4352 5736 4524 5738
rect 4322 5714 4350 5718
rect 4352 5714 4432 5736
rect 4453 5734 4468 5736
rect 4322 5712 4432 5714
rect 4253 5708 4432 5712
rect 4226 5698 4256 5708
rect 4258 5698 4411 5708
rect 4419 5698 4449 5708
rect 4453 5698 4483 5712
rect 4511 5698 4524 5736
rect 4596 5742 4631 5750
rect 4596 5716 4597 5742
rect 4604 5716 4631 5742
rect 4539 5698 4569 5712
rect 4596 5708 4631 5716
rect 4633 5742 4674 5750
rect 4633 5716 4648 5742
rect 4655 5716 4674 5742
rect 4738 5738 4800 5750
rect 4812 5738 4887 5750
rect 4945 5738 5020 5750
rect 5032 5738 5063 5750
rect 5069 5738 5104 5750
rect 4738 5736 4900 5738
rect 4633 5708 4674 5716
rect 4756 5712 4769 5736
rect 4784 5734 4799 5736
rect 4596 5698 4597 5708
rect 4612 5698 4625 5708
rect 4639 5698 4640 5708
rect 4655 5698 4668 5708
rect 4683 5698 4713 5712
rect 4756 5698 4799 5712
rect 4823 5709 4830 5716
rect 4833 5712 4900 5736
rect 4932 5736 5104 5738
rect 4902 5714 4930 5718
rect 4932 5714 5012 5736
rect 5033 5734 5048 5736
rect 4902 5712 5012 5714
rect 4833 5708 5012 5712
rect 4806 5698 4836 5708
rect 4838 5698 4991 5708
rect 4999 5698 5029 5708
rect 5033 5698 5063 5712
rect 5091 5698 5104 5736
rect 5176 5742 5211 5750
rect 5176 5716 5177 5742
rect 5184 5716 5211 5742
rect 5119 5698 5149 5712
rect 5176 5708 5211 5716
rect 5213 5742 5254 5750
rect 5213 5716 5228 5742
rect 5235 5716 5254 5742
rect 5318 5738 5380 5750
rect 5392 5738 5467 5750
rect 5525 5738 5600 5750
rect 5612 5738 5643 5750
rect 5649 5738 5684 5750
rect 5318 5736 5480 5738
rect 5213 5708 5254 5716
rect 5336 5712 5349 5736
rect 5364 5734 5379 5736
rect 5176 5698 5177 5708
rect 5192 5698 5205 5708
rect 5219 5698 5220 5708
rect 5235 5698 5248 5708
rect 5263 5698 5293 5712
rect 5336 5698 5379 5712
rect 5403 5709 5410 5716
rect 5413 5712 5480 5736
rect 5512 5736 5684 5738
rect 5482 5714 5510 5718
rect 5512 5714 5592 5736
rect 5613 5734 5628 5736
rect 5482 5712 5592 5714
rect 5413 5708 5592 5712
rect 5386 5698 5416 5708
rect 5418 5698 5571 5708
rect 5579 5698 5609 5708
rect 5613 5698 5643 5712
rect 5671 5698 5684 5736
rect 5756 5742 5791 5750
rect 5756 5716 5757 5742
rect 5764 5716 5791 5742
rect 5699 5698 5729 5712
rect 5756 5708 5791 5716
rect 5793 5742 5834 5750
rect 5793 5716 5808 5742
rect 5815 5716 5834 5742
rect 5898 5738 5960 5750
rect 5972 5738 6047 5750
rect 6105 5738 6180 5750
rect 6192 5738 6223 5750
rect 6229 5738 6264 5750
rect 5898 5736 6060 5738
rect 5793 5708 5834 5716
rect 5916 5712 5929 5736
rect 5944 5734 5959 5736
rect 5756 5698 5757 5708
rect 5772 5698 5785 5708
rect 5799 5698 5800 5708
rect 5815 5698 5828 5708
rect 5843 5698 5873 5712
rect 5916 5698 5959 5712
rect 5983 5709 5990 5716
rect 5993 5712 6060 5736
rect 6092 5736 6264 5738
rect 6062 5714 6090 5718
rect 6092 5714 6172 5736
rect 6193 5734 6208 5736
rect 6062 5712 6172 5714
rect 5993 5708 6172 5712
rect 5966 5698 5996 5708
rect 5998 5698 6151 5708
rect 6159 5698 6189 5708
rect 6193 5698 6223 5712
rect 6251 5698 6264 5736
rect 6336 5742 6371 5750
rect 6336 5716 6337 5742
rect 6344 5716 6371 5742
rect 6279 5698 6309 5712
rect 6336 5708 6371 5716
rect 6373 5742 6414 5750
rect 6373 5716 6388 5742
rect 6395 5716 6414 5742
rect 6478 5738 6540 5750
rect 6552 5738 6627 5750
rect 6685 5738 6760 5750
rect 6772 5738 6803 5750
rect 6809 5738 6844 5750
rect 6478 5736 6640 5738
rect 6373 5708 6414 5716
rect 6496 5712 6509 5736
rect 6524 5734 6539 5736
rect 6336 5698 6337 5708
rect 6352 5698 6365 5708
rect 6379 5698 6380 5708
rect 6395 5698 6408 5708
rect 6423 5698 6453 5712
rect 6496 5698 6539 5712
rect 6563 5709 6570 5716
rect 6573 5712 6640 5736
rect 6672 5736 6844 5738
rect 6642 5714 6670 5718
rect 6672 5714 6752 5736
rect 6773 5734 6788 5736
rect 6642 5712 6752 5714
rect 6573 5708 6752 5712
rect 6546 5698 6576 5708
rect 6578 5698 6731 5708
rect 6739 5698 6769 5708
rect 6773 5698 6803 5712
rect 6831 5698 6844 5736
rect 6916 5742 6951 5750
rect 6916 5716 6917 5742
rect 6924 5716 6951 5742
rect 6859 5698 6889 5712
rect 6916 5708 6951 5716
rect 6953 5742 6994 5750
rect 6953 5716 6968 5742
rect 6975 5716 6994 5742
rect 7058 5738 7120 5750
rect 7132 5738 7207 5750
rect 7265 5738 7340 5750
rect 7352 5738 7383 5750
rect 7389 5738 7424 5750
rect 7058 5736 7220 5738
rect 6953 5708 6994 5716
rect 7076 5712 7089 5736
rect 7104 5734 7119 5736
rect 6916 5698 6917 5708
rect 6932 5698 6945 5708
rect 6959 5698 6960 5708
rect 6975 5698 6988 5708
rect 7003 5698 7033 5712
rect 7076 5698 7119 5712
rect 7143 5709 7150 5716
rect 7153 5712 7220 5736
rect 7252 5736 7424 5738
rect 7222 5714 7250 5718
rect 7252 5714 7332 5736
rect 7353 5734 7368 5736
rect 7222 5712 7332 5714
rect 7153 5708 7332 5712
rect 7126 5698 7156 5708
rect 7158 5698 7311 5708
rect 7319 5698 7349 5708
rect 7353 5698 7383 5712
rect 7411 5698 7424 5736
rect 7496 5742 7531 5750
rect 7496 5716 7497 5742
rect 7504 5716 7531 5742
rect 7439 5698 7469 5712
rect 7496 5708 7531 5716
rect 7533 5742 7574 5750
rect 7533 5716 7548 5742
rect 7555 5716 7574 5742
rect 7638 5738 7700 5750
rect 7712 5738 7787 5750
rect 7845 5738 7920 5750
rect 7932 5738 7963 5750
rect 7969 5738 8004 5750
rect 7638 5736 7800 5738
rect 7533 5708 7574 5716
rect 7656 5712 7669 5736
rect 7684 5734 7699 5736
rect 7496 5698 7497 5708
rect 7512 5698 7525 5708
rect 7539 5698 7540 5708
rect 7555 5698 7568 5708
rect 7583 5698 7613 5712
rect 7656 5698 7699 5712
rect 7723 5709 7730 5716
rect 7733 5712 7800 5736
rect 7832 5736 8004 5738
rect 7802 5714 7830 5718
rect 7832 5714 7912 5736
rect 7933 5734 7948 5736
rect 7802 5712 7912 5714
rect 7733 5708 7912 5712
rect 7706 5698 7736 5708
rect 7738 5698 7891 5708
rect 7899 5698 7929 5708
rect 7933 5698 7963 5712
rect 7991 5698 8004 5736
rect 8076 5742 8111 5750
rect 8076 5716 8077 5742
rect 8084 5716 8111 5742
rect 8019 5698 8049 5712
rect 8076 5708 8111 5716
rect 8113 5742 8154 5750
rect 8113 5716 8128 5742
rect 8135 5716 8154 5742
rect 8218 5738 8280 5750
rect 8292 5738 8367 5750
rect 8425 5738 8500 5750
rect 8512 5738 8543 5750
rect 8549 5738 8584 5750
rect 8218 5736 8380 5738
rect 8113 5708 8154 5716
rect 8236 5712 8249 5736
rect 8264 5734 8279 5736
rect 8076 5698 8077 5708
rect 8092 5698 8105 5708
rect 8119 5698 8120 5708
rect 8135 5698 8148 5708
rect 8163 5698 8193 5712
rect 8236 5698 8279 5712
rect 8303 5709 8310 5716
rect 8313 5712 8380 5736
rect 8412 5736 8584 5738
rect 8382 5714 8410 5718
rect 8412 5714 8492 5736
rect 8513 5734 8528 5736
rect 8382 5712 8492 5714
rect 8313 5708 8492 5712
rect 8286 5698 8316 5708
rect 8318 5698 8471 5708
rect 8479 5698 8509 5708
rect 8513 5698 8543 5712
rect 8571 5698 8584 5736
rect 8656 5742 8691 5750
rect 8656 5716 8657 5742
rect 8664 5716 8691 5742
rect 8599 5698 8629 5712
rect 8656 5708 8691 5716
rect 8693 5742 8734 5750
rect 8693 5716 8708 5742
rect 8715 5716 8734 5742
rect 8798 5738 8860 5750
rect 8872 5738 8947 5750
rect 9005 5738 9080 5750
rect 9092 5738 9123 5750
rect 9129 5738 9164 5750
rect 8798 5736 8960 5738
rect 8693 5708 8734 5716
rect 8816 5712 8829 5736
rect 8844 5734 8859 5736
rect 8656 5698 8657 5708
rect 8672 5698 8685 5708
rect 8699 5698 8700 5708
rect 8715 5698 8728 5708
rect 8743 5698 8773 5712
rect 8816 5698 8859 5712
rect 8883 5709 8890 5716
rect 8893 5712 8960 5736
rect 8992 5736 9164 5738
rect 8962 5714 8990 5718
rect 8992 5714 9072 5736
rect 9093 5734 9108 5736
rect 8962 5712 9072 5714
rect 8893 5708 9072 5712
rect 8866 5698 8896 5708
rect 8898 5698 9051 5708
rect 9059 5698 9089 5708
rect 9093 5698 9123 5712
rect 9151 5698 9164 5736
rect 9236 5742 9271 5750
rect 9236 5716 9237 5742
rect 9244 5716 9271 5742
rect 9179 5698 9209 5712
rect 9236 5708 9271 5716
rect 9236 5698 9237 5708
rect 9252 5698 9265 5708
rect -1 5692 9265 5698
rect 0 5684 9265 5692
rect 15 5654 28 5684
rect 43 5666 73 5684
rect 116 5670 130 5684
rect 166 5670 386 5684
rect 117 5668 130 5670
rect 83 5656 98 5668
rect 80 5654 102 5656
rect 107 5654 137 5668
rect 198 5666 351 5670
rect 180 5654 372 5666
rect 415 5654 445 5668
rect 451 5654 464 5684
rect 479 5666 509 5684
rect 552 5654 565 5684
rect 595 5654 608 5684
rect 623 5666 653 5684
rect 696 5670 710 5684
rect 746 5670 966 5684
rect 697 5668 710 5670
rect 663 5656 678 5668
rect 660 5654 682 5656
rect 687 5654 717 5668
rect 778 5666 931 5670
rect 760 5654 952 5666
rect 995 5654 1025 5668
rect 1031 5654 1044 5684
rect 1059 5666 1089 5684
rect 1132 5654 1145 5684
rect 1175 5654 1188 5684
rect 1203 5666 1233 5684
rect 1276 5670 1290 5684
rect 1326 5670 1546 5684
rect 1277 5668 1290 5670
rect 1243 5656 1258 5668
rect 1240 5654 1262 5656
rect 1267 5654 1297 5668
rect 1358 5666 1511 5670
rect 1340 5654 1532 5666
rect 1575 5654 1605 5668
rect 1611 5654 1624 5684
rect 1639 5666 1669 5684
rect 1712 5654 1725 5684
rect 1755 5654 1768 5684
rect 1783 5666 1813 5684
rect 1856 5670 1870 5684
rect 1906 5670 2126 5684
rect 1857 5668 1870 5670
rect 1823 5656 1838 5668
rect 1820 5654 1842 5656
rect 1847 5654 1877 5668
rect 1938 5666 2091 5670
rect 1920 5654 2112 5666
rect 2155 5654 2185 5668
rect 2191 5654 2204 5684
rect 2219 5666 2249 5684
rect 2292 5654 2305 5684
rect 2335 5654 2348 5684
rect 2363 5666 2393 5684
rect 2436 5670 2450 5684
rect 2486 5670 2706 5684
rect 2437 5668 2450 5670
rect 2403 5656 2418 5668
rect 2400 5654 2422 5656
rect 2427 5654 2457 5668
rect 2518 5666 2671 5670
rect 2500 5654 2692 5666
rect 2735 5654 2765 5668
rect 2771 5654 2784 5684
rect 2799 5666 2829 5684
rect 2872 5654 2885 5684
rect 2915 5654 2928 5684
rect 2943 5666 2973 5684
rect 3016 5670 3030 5684
rect 3066 5670 3286 5684
rect 3017 5668 3030 5670
rect 2983 5656 2998 5668
rect 2980 5654 3002 5656
rect 3007 5654 3037 5668
rect 3098 5666 3251 5670
rect 3080 5654 3272 5666
rect 3315 5654 3345 5668
rect 3351 5654 3364 5684
rect 3379 5666 3409 5684
rect 3452 5654 3465 5684
rect 3495 5654 3508 5684
rect 3523 5666 3553 5684
rect 3596 5670 3610 5684
rect 3646 5670 3866 5684
rect 3597 5668 3610 5670
rect 3563 5656 3578 5668
rect 3560 5654 3582 5656
rect 3587 5654 3617 5668
rect 3678 5666 3831 5670
rect 3660 5654 3852 5666
rect 3895 5654 3925 5668
rect 3931 5654 3944 5684
rect 3959 5666 3989 5684
rect 4032 5654 4045 5684
rect 4075 5654 4088 5684
rect 4103 5666 4133 5684
rect 4176 5670 4190 5684
rect 4226 5670 4446 5684
rect 4177 5668 4190 5670
rect 4143 5656 4158 5668
rect 4140 5654 4162 5656
rect 4167 5654 4197 5668
rect 4258 5666 4411 5670
rect 4240 5654 4432 5666
rect 4475 5654 4505 5668
rect 4511 5654 4524 5684
rect 4539 5666 4569 5684
rect 4612 5654 4625 5684
rect 4655 5654 4668 5684
rect 4683 5666 4713 5684
rect 4756 5670 4770 5684
rect 4806 5670 5026 5684
rect 4757 5668 4770 5670
rect 4723 5656 4738 5668
rect 4720 5654 4742 5656
rect 4747 5654 4777 5668
rect 4838 5666 4991 5670
rect 4820 5654 5012 5666
rect 5055 5654 5085 5668
rect 5091 5654 5104 5684
rect 5119 5666 5149 5684
rect 5192 5654 5205 5684
rect 5235 5654 5248 5684
rect 5263 5666 5293 5684
rect 5336 5670 5350 5684
rect 5386 5670 5606 5684
rect 5337 5668 5350 5670
rect 5303 5656 5318 5668
rect 5300 5654 5322 5656
rect 5327 5654 5357 5668
rect 5418 5666 5571 5670
rect 5400 5654 5592 5666
rect 5635 5654 5665 5668
rect 5671 5654 5684 5684
rect 5699 5666 5729 5684
rect 5772 5654 5785 5684
rect 5815 5654 5828 5684
rect 5843 5666 5873 5684
rect 5916 5670 5930 5684
rect 5966 5670 6186 5684
rect 5917 5668 5930 5670
rect 5883 5656 5898 5668
rect 5880 5654 5902 5656
rect 5907 5654 5937 5668
rect 5998 5666 6151 5670
rect 5980 5654 6172 5666
rect 6215 5654 6245 5668
rect 6251 5654 6264 5684
rect 6279 5666 6309 5684
rect 6352 5654 6365 5684
rect 6395 5654 6408 5684
rect 6423 5666 6453 5684
rect 6496 5670 6510 5684
rect 6546 5670 6766 5684
rect 6497 5668 6510 5670
rect 6463 5656 6478 5668
rect 6460 5654 6482 5656
rect 6487 5654 6517 5668
rect 6578 5666 6731 5670
rect 6560 5654 6752 5666
rect 6795 5654 6825 5668
rect 6831 5654 6844 5684
rect 6859 5666 6889 5684
rect 6932 5654 6945 5684
rect 6975 5654 6988 5684
rect 7003 5666 7033 5684
rect 7076 5670 7090 5684
rect 7126 5670 7346 5684
rect 7077 5668 7090 5670
rect 7043 5656 7058 5668
rect 7040 5654 7062 5656
rect 7067 5654 7097 5668
rect 7158 5666 7311 5670
rect 7140 5654 7332 5666
rect 7375 5654 7405 5668
rect 7411 5654 7424 5684
rect 7439 5666 7469 5684
rect 7512 5654 7525 5684
rect 7555 5654 7568 5684
rect 7583 5666 7613 5684
rect 7656 5670 7670 5684
rect 7706 5670 7926 5684
rect 7657 5668 7670 5670
rect 7623 5656 7638 5668
rect 7620 5654 7642 5656
rect 7647 5654 7677 5668
rect 7738 5666 7891 5670
rect 7720 5654 7912 5666
rect 7955 5654 7985 5668
rect 7991 5654 8004 5684
rect 8019 5666 8049 5684
rect 8092 5654 8105 5684
rect 8135 5654 8148 5684
rect 8163 5666 8193 5684
rect 8236 5670 8250 5684
rect 8286 5670 8506 5684
rect 8237 5668 8250 5670
rect 8203 5656 8218 5668
rect 8200 5654 8222 5656
rect 8227 5654 8257 5668
rect 8318 5666 8471 5670
rect 8300 5654 8492 5666
rect 8535 5654 8565 5668
rect 8571 5654 8584 5684
rect 8599 5666 8629 5684
rect 8672 5654 8685 5684
rect 8715 5654 8728 5684
rect 8743 5666 8773 5684
rect 8816 5670 8830 5684
rect 8866 5670 9086 5684
rect 8817 5668 8830 5670
rect 8783 5656 8798 5668
rect 8780 5654 8802 5656
rect 8807 5654 8837 5668
rect 8898 5666 9051 5670
rect 8880 5654 9072 5666
rect 9115 5654 9145 5668
rect 9151 5654 9164 5684
rect 9179 5666 9209 5684
rect 9252 5654 9265 5684
rect 0 5640 9265 5654
rect 15 5536 28 5640
rect 73 5618 74 5628
rect 89 5618 102 5628
rect 73 5614 102 5618
rect 107 5614 137 5640
rect 155 5626 171 5628
rect 243 5626 296 5640
rect 244 5624 308 5626
rect 351 5624 366 5640
rect 415 5637 445 5640
rect 415 5634 451 5637
rect 381 5626 397 5628
rect 155 5614 170 5618
rect 73 5612 170 5614
rect 198 5612 366 5624
rect 382 5614 397 5618
rect 415 5615 454 5634
rect 473 5628 480 5629
rect 479 5621 480 5628
rect 463 5618 464 5621
rect 479 5618 492 5621
rect 415 5614 445 5615
rect 454 5614 460 5615
rect 463 5614 492 5618
rect 382 5613 492 5614
rect 382 5612 498 5613
rect 57 5604 108 5612
rect 57 5592 82 5604
rect 89 5592 108 5604
rect 139 5604 189 5612
rect 139 5596 155 5604
rect 162 5602 189 5604
rect 198 5602 419 5612
rect 162 5592 419 5602
rect 448 5604 498 5612
rect 448 5595 464 5604
rect 57 5584 108 5592
rect 155 5584 419 5592
rect 445 5592 464 5595
rect 471 5592 498 5604
rect 445 5584 498 5592
rect 73 5576 74 5584
rect 89 5576 102 5584
rect 73 5568 89 5576
rect 70 5561 89 5564
rect 70 5552 92 5561
rect 43 5542 92 5552
rect 43 5536 73 5542
rect 92 5537 97 5542
rect 15 5520 89 5536
rect 107 5528 137 5584
rect 172 5574 380 5584
rect 415 5580 460 5584
rect 463 5583 464 5584
rect 479 5583 492 5584
rect 198 5544 387 5574
rect 213 5541 387 5544
rect 206 5538 387 5541
rect 15 5518 28 5520
rect 43 5518 77 5520
rect 15 5502 89 5518
rect 116 5514 129 5528
rect 144 5514 160 5530
rect 206 5525 217 5538
rect -1 5480 0 5496
rect 15 5480 28 5502
rect 43 5480 73 5502
rect 116 5498 178 5514
rect 206 5507 217 5523
rect 222 5518 232 5538
rect 242 5518 256 5538
rect 259 5525 268 5538
rect 284 5525 293 5538
rect 222 5507 256 5518
rect 259 5507 268 5523
rect 284 5507 293 5523
rect 300 5518 310 5538
rect 320 5518 334 5538
rect 335 5525 346 5538
rect 300 5507 334 5518
rect 335 5507 346 5523
rect 392 5514 408 5530
rect 415 5528 445 5580
rect 479 5576 480 5583
rect 464 5568 480 5576
rect 451 5536 464 5555
rect 479 5536 509 5552
rect 451 5520 525 5536
rect 451 5518 464 5520
rect 479 5518 513 5520
rect 116 5496 129 5498
rect 144 5496 178 5498
rect 116 5480 178 5496
rect 222 5491 238 5494
rect 300 5491 330 5502
rect 378 5498 424 5514
rect 451 5502 525 5518
rect 378 5496 412 5498
rect 377 5480 424 5496
rect 451 5480 464 5502
rect 479 5480 509 5502
rect 536 5480 537 5496
rect 552 5480 565 5640
rect 595 5536 608 5640
rect 653 5618 654 5628
rect 669 5618 682 5628
rect 653 5614 682 5618
rect 687 5614 717 5640
rect 735 5626 751 5628
rect 823 5626 876 5640
rect 824 5624 888 5626
rect 931 5624 946 5640
rect 995 5637 1025 5640
rect 995 5634 1031 5637
rect 961 5626 977 5628
rect 735 5614 750 5618
rect 653 5612 750 5614
rect 778 5612 946 5624
rect 962 5614 977 5618
rect 995 5615 1034 5634
rect 1053 5628 1060 5629
rect 1059 5621 1060 5628
rect 1043 5618 1044 5621
rect 1059 5618 1072 5621
rect 995 5614 1025 5615
rect 1034 5614 1040 5615
rect 1043 5614 1072 5618
rect 962 5613 1072 5614
rect 962 5612 1078 5613
rect 637 5604 688 5612
rect 637 5592 662 5604
rect 669 5592 688 5604
rect 719 5604 769 5612
rect 719 5596 735 5604
rect 742 5602 769 5604
rect 778 5602 999 5612
rect 742 5592 999 5602
rect 1028 5604 1078 5612
rect 1028 5595 1044 5604
rect 637 5584 688 5592
rect 735 5584 999 5592
rect 1025 5592 1044 5595
rect 1051 5592 1078 5604
rect 1025 5584 1078 5592
rect 653 5576 654 5584
rect 669 5576 682 5584
rect 653 5568 669 5576
rect 650 5561 669 5564
rect 650 5552 672 5561
rect 623 5542 672 5552
rect 623 5536 653 5542
rect 672 5537 677 5542
rect 595 5520 669 5536
rect 687 5528 717 5584
rect 752 5574 960 5584
rect 995 5580 1040 5584
rect 1043 5583 1044 5584
rect 1059 5583 1072 5584
rect 778 5544 967 5574
rect 793 5541 967 5544
rect 786 5538 967 5541
rect 595 5518 608 5520
rect 623 5518 657 5520
rect 595 5502 669 5518
rect 696 5514 709 5528
rect 724 5514 740 5530
rect 786 5525 797 5538
rect 579 5480 580 5496
rect 595 5480 608 5502
rect 623 5480 653 5502
rect 696 5498 758 5514
rect 786 5507 797 5523
rect 802 5518 812 5538
rect 822 5518 836 5538
rect 839 5525 848 5538
rect 864 5525 873 5538
rect 802 5507 836 5518
rect 839 5507 848 5523
rect 864 5507 873 5523
rect 880 5518 890 5538
rect 900 5518 914 5538
rect 915 5525 926 5538
rect 880 5507 914 5518
rect 915 5507 926 5523
rect 972 5514 988 5530
rect 995 5528 1025 5580
rect 1059 5576 1060 5583
rect 1044 5568 1060 5576
rect 1031 5536 1044 5555
rect 1059 5536 1089 5552
rect 1031 5520 1105 5536
rect 1031 5518 1044 5520
rect 1059 5518 1093 5520
rect 696 5496 709 5498
rect 724 5496 758 5498
rect 696 5480 758 5496
rect 802 5491 818 5494
rect 880 5491 910 5502
rect 958 5498 1004 5514
rect 1031 5502 1105 5518
rect 958 5496 992 5498
rect 957 5480 1004 5496
rect 1031 5480 1044 5502
rect 1059 5480 1089 5502
rect 1116 5480 1117 5496
rect 1132 5480 1145 5640
rect 1175 5536 1188 5640
rect 1233 5618 1234 5628
rect 1249 5618 1262 5628
rect 1233 5614 1262 5618
rect 1267 5614 1297 5640
rect 1315 5626 1331 5628
rect 1403 5626 1456 5640
rect 1404 5624 1468 5626
rect 1511 5624 1526 5640
rect 1575 5637 1605 5640
rect 1575 5634 1611 5637
rect 1541 5626 1557 5628
rect 1315 5614 1330 5618
rect 1233 5612 1330 5614
rect 1358 5612 1526 5624
rect 1542 5614 1557 5618
rect 1575 5615 1614 5634
rect 1633 5628 1640 5629
rect 1639 5621 1640 5628
rect 1623 5618 1624 5621
rect 1639 5618 1652 5621
rect 1575 5614 1605 5615
rect 1614 5614 1620 5615
rect 1623 5614 1652 5618
rect 1542 5613 1652 5614
rect 1542 5612 1658 5613
rect 1217 5604 1268 5612
rect 1217 5592 1242 5604
rect 1249 5592 1268 5604
rect 1299 5604 1349 5612
rect 1299 5596 1315 5604
rect 1322 5602 1349 5604
rect 1358 5602 1579 5612
rect 1322 5592 1579 5602
rect 1608 5604 1658 5612
rect 1608 5595 1624 5604
rect 1217 5584 1268 5592
rect 1315 5584 1579 5592
rect 1605 5592 1624 5595
rect 1631 5592 1658 5604
rect 1605 5584 1658 5592
rect 1233 5576 1234 5584
rect 1249 5576 1262 5584
rect 1233 5568 1249 5576
rect 1230 5561 1249 5564
rect 1230 5552 1252 5561
rect 1203 5542 1252 5552
rect 1203 5536 1233 5542
rect 1252 5537 1257 5542
rect 1175 5520 1249 5536
rect 1267 5528 1297 5584
rect 1332 5574 1540 5584
rect 1575 5580 1620 5584
rect 1623 5583 1624 5584
rect 1639 5583 1652 5584
rect 1358 5544 1547 5574
rect 1373 5541 1547 5544
rect 1366 5538 1547 5541
rect 1175 5518 1188 5520
rect 1203 5518 1237 5520
rect 1175 5502 1249 5518
rect 1276 5514 1289 5528
rect 1304 5514 1320 5530
rect 1366 5525 1377 5538
rect 1159 5480 1160 5496
rect 1175 5480 1188 5502
rect 1203 5480 1233 5502
rect 1276 5498 1338 5514
rect 1366 5507 1377 5523
rect 1382 5518 1392 5538
rect 1402 5518 1416 5538
rect 1419 5525 1428 5538
rect 1444 5525 1453 5538
rect 1382 5507 1416 5518
rect 1419 5507 1428 5523
rect 1444 5507 1453 5523
rect 1460 5518 1470 5538
rect 1480 5518 1494 5538
rect 1495 5525 1506 5538
rect 1460 5507 1494 5518
rect 1495 5507 1506 5523
rect 1552 5514 1568 5530
rect 1575 5528 1605 5580
rect 1639 5576 1640 5583
rect 1624 5568 1640 5576
rect 1611 5536 1624 5555
rect 1639 5536 1669 5552
rect 1611 5520 1685 5536
rect 1611 5518 1624 5520
rect 1639 5518 1673 5520
rect 1276 5496 1289 5498
rect 1304 5496 1338 5498
rect 1276 5480 1338 5496
rect 1382 5491 1398 5494
rect 1460 5491 1490 5502
rect 1538 5498 1584 5514
rect 1611 5502 1685 5518
rect 1538 5496 1572 5498
rect 1537 5480 1584 5496
rect 1611 5480 1624 5502
rect 1639 5480 1669 5502
rect 1696 5480 1697 5496
rect 1712 5480 1725 5640
rect 1755 5536 1768 5640
rect 1813 5618 1814 5628
rect 1829 5618 1842 5628
rect 1813 5614 1842 5618
rect 1847 5614 1877 5640
rect 1895 5626 1911 5628
rect 1983 5626 2036 5640
rect 1984 5624 2048 5626
rect 2091 5624 2106 5640
rect 2155 5637 2185 5640
rect 2155 5634 2191 5637
rect 2121 5626 2137 5628
rect 1895 5614 1910 5618
rect 1813 5612 1910 5614
rect 1938 5612 2106 5624
rect 2122 5614 2137 5618
rect 2155 5615 2194 5634
rect 2213 5628 2220 5629
rect 2219 5621 2220 5628
rect 2203 5618 2204 5621
rect 2219 5618 2232 5621
rect 2155 5614 2185 5615
rect 2194 5614 2200 5615
rect 2203 5614 2232 5618
rect 2122 5613 2232 5614
rect 2122 5612 2238 5613
rect 1797 5604 1848 5612
rect 1797 5592 1822 5604
rect 1829 5592 1848 5604
rect 1879 5604 1929 5612
rect 1879 5596 1895 5604
rect 1902 5602 1929 5604
rect 1938 5602 2159 5612
rect 1902 5592 2159 5602
rect 2188 5604 2238 5612
rect 2188 5595 2204 5604
rect 1797 5584 1848 5592
rect 1895 5584 2159 5592
rect 2185 5592 2204 5595
rect 2211 5592 2238 5604
rect 2185 5584 2238 5592
rect 1813 5576 1814 5584
rect 1829 5576 1842 5584
rect 1813 5568 1829 5576
rect 1810 5561 1829 5564
rect 1810 5552 1832 5561
rect 1783 5542 1832 5552
rect 1783 5536 1813 5542
rect 1832 5537 1837 5542
rect 1755 5520 1829 5536
rect 1847 5528 1877 5584
rect 1912 5574 2120 5584
rect 2155 5580 2200 5584
rect 2203 5583 2204 5584
rect 2219 5583 2232 5584
rect 1938 5544 2127 5574
rect 1953 5541 2127 5544
rect 1946 5538 2127 5541
rect 1755 5518 1768 5520
rect 1783 5518 1817 5520
rect 1755 5502 1829 5518
rect 1856 5514 1869 5528
rect 1884 5514 1900 5530
rect 1946 5525 1957 5538
rect 1739 5480 1740 5496
rect 1755 5480 1768 5502
rect 1783 5480 1813 5502
rect 1856 5498 1918 5514
rect 1946 5507 1957 5523
rect 1962 5518 1972 5538
rect 1982 5518 1996 5538
rect 1999 5525 2008 5538
rect 2024 5525 2033 5538
rect 1962 5507 1996 5518
rect 1999 5507 2008 5523
rect 2024 5507 2033 5523
rect 2040 5518 2050 5538
rect 2060 5518 2074 5538
rect 2075 5525 2086 5538
rect 2040 5507 2074 5518
rect 2075 5507 2086 5523
rect 2132 5514 2148 5530
rect 2155 5528 2185 5580
rect 2219 5576 2220 5583
rect 2204 5568 2220 5576
rect 2191 5536 2204 5555
rect 2219 5536 2249 5552
rect 2191 5520 2265 5536
rect 2191 5518 2204 5520
rect 2219 5518 2253 5520
rect 1856 5496 1869 5498
rect 1884 5496 1918 5498
rect 1856 5480 1918 5496
rect 1962 5491 1976 5494
rect 2040 5491 2070 5502
rect 2118 5498 2164 5514
rect 2191 5502 2265 5518
rect 2118 5496 2152 5498
rect 2117 5480 2164 5496
rect 2191 5480 2204 5502
rect 2219 5480 2249 5502
rect 2276 5480 2277 5496
rect 2292 5480 2305 5640
rect 2335 5536 2348 5640
rect 2393 5618 2394 5628
rect 2409 5618 2422 5628
rect 2393 5614 2422 5618
rect 2427 5614 2457 5640
rect 2475 5626 2491 5628
rect 2563 5626 2616 5640
rect 2564 5624 2628 5626
rect 2671 5624 2686 5640
rect 2735 5637 2765 5640
rect 2735 5634 2771 5637
rect 2701 5626 2717 5628
rect 2475 5614 2490 5618
rect 2393 5612 2490 5614
rect 2518 5612 2686 5624
rect 2702 5614 2717 5618
rect 2735 5615 2774 5634
rect 2793 5628 2800 5629
rect 2799 5621 2800 5628
rect 2783 5618 2784 5621
rect 2799 5618 2812 5621
rect 2735 5614 2765 5615
rect 2774 5614 2780 5615
rect 2783 5614 2812 5618
rect 2702 5613 2812 5614
rect 2702 5612 2818 5613
rect 2377 5604 2428 5612
rect 2377 5592 2402 5604
rect 2409 5592 2428 5604
rect 2459 5604 2509 5612
rect 2459 5596 2475 5604
rect 2482 5602 2509 5604
rect 2518 5602 2739 5612
rect 2482 5592 2739 5602
rect 2768 5604 2818 5612
rect 2768 5595 2784 5604
rect 2377 5584 2428 5592
rect 2475 5584 2739 5592
rect 2765 5592 2784 5595
rect 2791 5592 2818 5604
rect 2765 5584 2818 5592
rect 2393 5576 2394 5584
rect 2409 5576 2422 5584
rect 2393 5568 2409 5576
rect 2390 5561 2409 5564
rect 2390 5552 2412 5561
rect 2363 5542 2412 5552
rect 2363 5536 2393 5542
rect 2412 5537 2417 5542
rect 2335 5520 2409 5536
rect 2427 5528 2457 5584
rect 2492 5574 2700 5584
rect 2735 5580 2780 5584
rect 2783 5583 2784 5584
rect 2799 5583 2812 5584
rect 2518 5544 2707 5574
rect 2533 5541 2707 5544
rect 2526 5538 2707 5541
rect 2335 5518 2348 5520
rect 2363 5518 2397 5520
rect 2335 5502 2409 5518
rect 2436 5514 2449 5528
rect 2464 5514 2480 5530
rect 2526 5525 2537 5538
rect 2319 5480 2320 5496
rect 2335 5480 2348 5502
rect 2363 5480 2393 5502
rect 2436 5498 2498 5514
rect 2526 5507 2537 5523
rect 2542 5518 2552 5538
rect 2562 5518 2576 5538
rect 2579 5525 2588 5538
rect 2604 5525 2613 5538
rect 2542 5507 2576 5518
rect 2579 5507 2588 5523
rect 2604 5507 2613 5523
rect 2620 5518 2630 5538
rect 2640 5518 2654 5538
rect 2655 5525 2666 5538
rect 2620 5507 2654 5518
rect 2655 5507 2666 5523
rect 2712 5514 2728 5530
rect 2735 5528 2765 5580
rect 2799 5576 2800 5583
rect 2784 5568 2800 5576
rect 2771 5536 2784 5555
rect 2799 5536 2829 5552
rect 2771 5520 2845 5536
rect 2771 5518 2784 5520
rect 2799 5518 2833 5520
rect 2436 5496 2449 5498
rect 2464 5496 2498 5498
rect 2436 5480 2498 5496
rect 2542 5491 2558 5494
rect 2620 5491 2650 5502
rect 2698 5498 2744 5514
rect 2771 5502 2845 5518
rect 2698 5496 2732 5498
rect 2697 5480 2744 5496
rect 2771 5480 2784 5502
rect 2799 5480 2829 5502
rect 2856 5480 2857 5496
rect 2872 5480 2885 5640
rect 2915 5536 2928 5640
rect 2973 5618 2974 5628
rect 2989 5618 3002 5628
rect 2973 5614 3002 5618
rect 3007 5614 3037 5640
rect 3055 5626 3071 5628
rect 3143 5626 3196 5640
rect 3144 5624 3208 5626
rect 3251 5624 3266 5640
rect 3315 5637 3345 5640
rect 3315 5634 3351 5637
rect 3281 5626 3297 5628
rect 3055 5614 3070 5618
rect 2973 5612 3070 5614
rect 3098 5612 3266 5624
rect 3282 5614 3297 5618
rect 3315 5615 3354 5634
rect 3373 5628 3380 5629
rect 3379 5621 3380 5628
rect 3363 5618 3364 5621
rect 3379 5618 3392 5621
rect 3315 5614 3345 5615
rect 3354 5614 3360 5615
rect 3363 5614 3392 5618
rect 3282 5613 3392 5614
rect 3282 5612 3398 5613
rect 2957 5604 3008 5612
rect 2957 5592 2982 5604
rect 2989 5592 3008 5604
rect 3039 5604 3089 5612
rect 3039 5596 3055 5604
rect 3062 5602 3089 5604
rect 3098 5602 3319 5612
rect 3062 5592 3319 5602
rect 3348 5604 3398 5612
rect 3348 5595 3364 5604
rect 2957 5584 3008 5592
rect 3055 5584 3319 5592
rect 3345 5592 3364 5595
rect 3371 5592 3398 5604
rect 3345 5584 3398 5592
rect 2973 5576 2974 5584
rect 2989 5576 3002 5584
rect 2973 5568 2989 5576
rect 2970 5561 2989 5564
rect 2970 5552 2992 5561
rect 2943 5542 2992 5552
rect 2943 5536 2973 5542
rect 2992 5537 2997 5542
rect 2915 5520 2989 5536
rect 3007 5528 3037 5584
rect 3072 5574 3280 5584
rect 3315 5580 3360 5584
rect 3363 5583 3364 5584
rect 3379 5583 3392 5584
rect 3098 5544 3287 5574
rect 3113 5541 3287 5544
rect 3106 5538 3287 5541
rect 2915 5518 2928 5520
rect 2943 5518 2977 5520
rect 2915 5502 2989 5518
rect 3016 5514 3029 5528
rect 3044 5514 3060 5530
rect 3106 5525 3117 5538
rect 2899 5480 2900 5496
rect 2915 5480 2928 5502
rect 2943 5480 2973 5502
rect 3016 5498 3078 5514
rect 3106 5507 3117 5523
rect 3122 5518 3132 5538
rect 3142 5518 3156 5538
rect 3159 5525 3168 5538
rect 3184 5525 3193 5538
rect 3122 5507 3156 5518
rect 3159 5507 3168 5523
rect 3184 5507 3193 5523
rect 3200 5518 3210 5538
rect 3220 5518 3234 5538
rect 3235 5525 3246 5538
rect 3200 5507 3234 5518
rect 3235 5507 3246 5523
rect 3292 5514 3308 5530
rect 3315 5528 3345 5580
rect 3379 5576 3380 5583
rect 3364 5568 3380 5576
rect 3351 5536 3364 5555
rect 3379 5536 3409 5552
rect 3351 5520 3425 5536
rect 3351 5518 3364 5520
rect 3379 5518 3413 5520
rect 3016 5496 3029 5498
rect 3044 5496 3078 5498
rect 3016 5480 3078 5496
rect 3122 5491 3138 5494
rect 3200 5491 3230 5502
rect 3278 5498 3324 5514
rect 3351 5502 3425 5518
rect 3278 5496 3312 5498
rect 3277 5480 3324 5496
rect 3351 5480 3364 5502
rect 3379 5480 3409 5502
rect 3436 5480 3437 5496
rect 3452 5480 3465 5640
rect 3495 5536 3508 5640
rect 3553 5618 3554 5628
rect 3569 5618 3582 5628
rect 3553 5614 3582 5618
rect 3587 5614 3617 5640
rect 3635 5626 3651 5628
rect 3723 5626 3776 5640
rect 3724 5624 3788 5626
rect 3831 5624 3846 5640
rect 3895 5637 3925 5640
rect 3895 5634 3931 5637
rect 3861 5626 3877 5628
rect 3635 5614 3650 5618
rect 3553 5612 3650 5614
rect 3678 5612 3846 5624
rect 3862 5614 3877 5618
rect 3895 5615 3934 5634
rect 3953 5628 3960 5629
rect 3959 5621 3960 5628
rect 3943 5618 3944 5621
rect 3959 5618 3972 5621
rect 3895 5614 3925 5615
rect 3934 5614 3940 5615
rect 3943 5614 3972 5618
rect 3862 5613 3972 5614
rect 3862 5612 3978 5613
rect 3537 5604 3588 5612
rect 3537 5592 3562 5604
rect 3569 5592 3588 5604
rect 3619 5604 3669 5612
rect 3619 5596 3635 5604
rect 3642 5602 3669 5604
rect 3678 5602 3899 5612
rect 3642 5592 3899 5602
rect 3928 5604 3978 5612
rect 3928 5595 3944 5604
rect 3537 5584 3588 5592
rect 3635 5584 3899 5592
rect 3925 5592 3944 5595
rect 3951 5592 3978 5604
rect 3925 5584 3978 5592
rect 3553 5576 3554 5584
rect 3569 5576 3582 5584
rect 3553 5568 3569 5576
rect 3550 5561 3569 5564
rect 3550 5552 3572 5561
rect 3523 5542 3572 5552
rect 3523 5536 3553 5542
rect 3572 5537 3577 5542
rect 3495 5520 3569 5536
rect 3587 5528 3617 5584
rect 3652 5574 3860 5584
rect 3895 5580 3940 5584
rect 3943 5583 3944 5584
rect 3959 5583 3972 5584
rect 3678 5544 3867 5574
rect 3693 5541 3867 5544
rect 3686 5538 3867 5541
rect 3495 5518 3508 5520
rect 3523 5518 3557 5520
rect 3495 5502 3569 5518
rect 3596 5514 3609 5528
rect 3624 5514 3640 5530
rect 3686 5525 3697 5538
rect 3479 5480 3480 5496
rect 3495 5480 3508 5502
rect 3523 5480 3553 5502
rect 3596 5498 3658 5514
rect 3686 5507 3697 5523
rect 3702 5518 3712 5538
rect 3722 5518 3736 5538
rect 3739 5525 3748 5538
rect 3764 5525 3773 5538
rect 3702 5507 3736 5518
rect 3739 5507 3748 5523
rect 3764 5507 3773 5523
rect 3780 5518 3790 5538
rect 3800 5518 3814 5538
rect 3815 5525 3826 5538
rect 3780 5507 3814 5518
rect 3815 5507 3826 5523
rect 3872 5514 3888 5530
rect 3895 5528 3925 5580
rect 3959 5576 3960 5583
rect 3944 5568 3960 5576
rect 3931 5536 3944 5555
rect 3959 5536 3989 5552
rect 3931 5520 4005 5536
rect 3931 5518 3944 5520
rect 3959 5518 3993 5520
rect 3596 5496 3609 5498
rect 3624 5496 3658 5498
rect 3596 5480 3658 5496
rect 3702 5491 3718 5494
rect 3780 5491 3810 5502
rect 3858 5498 3904 5514
rect 3931 5502 4005 5518
rect 3858 5496 3892 5498
rect 3857 5480 3904 5496
rect 3931 5480 3944 5502
rect 3959 5480 3989 5502
rect 4016 5480 4017 5496
rect 4032 5480 4045 5640
rect 4075 5536 4088 5640
rect 4133 5618 4134 5628
rect 4149 5618 4162 5628
rect 4133 5614 4162 5618
rect 4167 5614 4197 5640
rect 4215 5626 4231 5628
rect 4303 5626 4356 5640
rect 4304 5624 4368 5626
rect 4411 5624 4426 5640
rect 4475 5637 4505 5640
rect 4475 5634 4511 5637
rect 4441 5626 4457 5628
rect 4215 5614 4230 5618
rect 4133 5612 4230 5614
rect 4258 5612 4426 5624
rect 4442 5614 4457 5618
rect 4475 5615 4514 5634
rect 4533 5628 4540 5629
rect 4539 5621 4540 5628
rect 4523 5618 4524 5621
rect 4539 5618 4552 5621
rect 4475 5614 4505 5615
rect 4514 5614 4520 5615
rect 4523 5614 4552 5618
rect 4442 5613 4552 5614
rect 4442 5612 4558 5613
rect 4117 5604 4168 5612
rect 4117 5592 4142 5604
rect 4149 5592 4168 5604
rect 4199 5604 4249 5612
rect 4199 5596 4215 5604
rect 4222 5602 4249 5604
rect 4258 5602 4479 5612
rect 4222 5592 4479 5602
rect 4508 5604 4558 5612
rect 4508 5595 4524 5604
rect 4117 5584 4168 5592
rect 4215 5584 4479 5592
rect 4505 5592 4524 5595
rect 4531 5592 4558 5604
rect 4505 5584 4558 5592
rect 4133 5576 4134 5584
rect 4149 5576 4162 5584
rect 4133 5568 4149 5576
rect 4130 5561 4149 5564
rect 4130 5552 4152 5561
rect 4103 5542 4152 5552
rect 4103 5536 4133 5542
rect 4152 5537 4157 5542
rect 4075 5520 4149 5536
rect 4167 5528 4197 5584
rect 4232 5574 4440 5584
rect 4475 5580 4520 5584
rect 4523 5583 4524 5584
rect 4539 5583 4552 5584
rect 4258 5544 4447 5574
rect 4273 5541 4447 5544
rect 4266 5538 4447 5541
rect 4075 5518 4088 5520
rect 4103 5518 4137 5520
rect 4075 5502 4149 5518
rect 4176 5514 4189 5528
rect 4204 5514 4220 5530
rect 4266 5525 4277 5538
rect 4059 5480 4060 5496
rect 4075 5480 4088 5502
rect 4103 5480 4133 5502
rect 4176 5498 4238 5514
rect 4266 5507 4277 5523
rect 4282 5518 4292 5538
rect 4302 5518 4316 5538
rect 4319 5525 4328 5538
rect 4344 5525 4353 5538
rect 4282 5507 4316 5518
rect 4319 5507 4328 5523
rect 4344 5507 4353 5523
rect 4360 5518 4370 5538
rect 4380 5518 4394 5538
rect 4395 5525 4406 5538
rect 4360 5507 4394 5518
rect 4395 5507 4406 5523
rect 4452 5514 4468 5530
rect 4475 5528 4505 5580
rect 4539 5576 4540 5583
rect 4524 5568 4540 5576
rect 4511 5536 4524 5555
rect 4539 5536 4569 5552
rect 4511 5520 4585 5536
rect 4511 5518 4524 5520
rect 4539 5518 4573 5520
rect 4176 5496 4189 5498
rect 4204 5496 4238 5498
rect 4176 5480 4238 5496
rect 4282 5491 4298 5494
rect 4360 5491 4390 5502
rect 4438 5498 4484 5514
rect 4511 5502 4585 5518
rect 4438 5496 4472 5498
rect 4437 5480 4484 5496
rect 4511 5480 4524 5502
rect 4539 5480 4569 5502
rect 4596 5480 4597 5496
rect 4612 5480 4625 5640
rect 4655 5536 4668 5640
rect 4713 5618 4714 5628
rect 4729 5618 4742 5628
rect 4713 5614 4742 5618
rect 4747 5614 4777 5640
rect 4795 5626 4811 5628
rect 4883 5626 4936 5640
rect 4884 5624 4948 5626
rect 4991 5624 5006 5640
rect 5055 5637 5085 5640
rect 5055 5634 5091 5637
rect 5021 5626 5037 5628
rect 4795 5614 4810 5618
rect 4713 5612 4810 5614
rect 4838 5612 5006 5624
rect 5022 5614 5037 5618
rect 5055 5615 5094 5634
rect 5113 5628 5120 5629
rect 5119 5621 5120 5628
rect 5103 5618 5104 5621
rect 5119 5618 5132 5621
rect 5055 5614 5085 5615
rect 5094 5614 5100 5615
rect 5103 5614 5132 5618
rect 5022 5613 5132 5614
rect 5022 5612 5138 5613
rect 4697 5604 4748 5612
rect 4697 5592 4722 5604
rect 4729 5592 4748 5604
rect 4779 5604 4829 5612
rect 4779 5596 4795 5604
rect 4802 5602 4829 5604
rect 4838 5602 5059 5612
rect 4802 5592 5059 5602
rect 5088 5604 5138 5612
rect 5088 5595 5104 5604
rect 4697 5584 4748 5592
rect 4795 5584 5059 5592
rect 5085 5592 5104 5595
rect 5111 5592 5138 5604
rect 5085 5584 5138 5592
rect 4713 5576 4714 5584
rect 4729 5576 4742 5584
rect 4713 5568 4729 5576
rect 4710 5561 4729 5564
rect 4710 5552 4732 5561
rect 4683 5542 4732 5552
rect 4683 5536 4713 5542
rect 4732 5537 4737 5542
rect 4655 5520 4729 5536
rect 4747 5528 4777 5584
rect 4812 5574 5020 5584
rect 5055 5580 5100 5584
rect 5103 5583 5104 5584
rect 5119 5583 5132 5584
rect 4838 5544 5027 5574
rect 4853 5541 5027 5544
rect 4846 5538 5027 5541
rect 4655 5518 4668 5520
rect 4683 5518 4717 5520
rect 4655 5502 4729 5518
rect 4756 5514 4769 5528
rect 4784 5514 4800 5530
rect 4846 5525 4857 5538
rect 4639 5480 4640 5496
rect 4655 5480 4668 5502
rect 4683 5480 4713 5502
rect 4756 5498 4818 5514
rect 4846 5507 4857 5523
rect 4862 5518 4872 5538
rect 4882 5518 4896 5538
rect 4899 5525 4908 5538
rect 4924 5525 4933 5538
rect 4862 5507 4896 5518
rect 4899 5507 4908 5523
rect 4924 5507 4933 5523
rect 4940 5518 4950 5538
rect 4960 5518 4974 5538
rect 4975 5525 4986 5538
rect 4940 5507 4974 5518
rect 4975 5507 4986 5523
rect 5032 5514 5048 5530
rect 5055 5528 5085 5580
rect 5119 5576 5120 5583
rect 5104 5568 5120 5576
rect 5091 5536 5104 5555
rect 5119 5536 5149 5552
rect 5091 5520 5165 5536
rect 5091 5518 5104 5520
rect 5119 5518 5153 5520
rect 4756 5496 4769 5498
rect 4784 5496 4818 5498
rect 4756 5480 4818 5496
rect 4862 5491 4878 5494
rect 4940 5491 4970 5502
rect 5018 5498 5064 5514
rect 5091 5502 5165 5518
rect 5018 5496 5052 5498
rect 5017 5480 5064 5496
rect 5091 5480 5104 5502
rect 5119 5480 5149 5502
rect 5176 5480 5177 5496
rect 5192 5480 5205 5640
rect 5235 5536 5248 5640
rect 5293 5618 5294 5628
rect 5309 5618 5322 5628
rect 5293 5614 5322 5618
rect 5327 5614 5357 5640
rect 5375 5626 5391 5628
rect 5463 5626 5516 5640
rect 5464 5624 5528 5626
rect 5571 5624 5586 5640
rect 5635 5637 5665 5640
rect 5635 5634 5671 5637
rect 5601 5626 5617 5628
rect 5375 5614 5390 5618
rect 5293 5612 5390 5614
rect 5418 5612 5586 5624
rect 5602 5614 5617 5618
rect 5635 5615 5674 5634
rect 5693 5628 5700 5629
rect 5699 5621 5700 5628
rect 5683 5618 5684 5621
rect 5699 5618 5712 5621
rect 5635 5614 5665 5615
rect 5674 5614 5680 5615
rect 5683 5614 5712 5618
rect 5602 5613 5712 5614
rect 5602 5612 5718 5613
rect 5277 5604 5328 5612
rect 5277 5592 5302 5604
rect 5309 5592 5328 5604
rect 5359 5604 5409 5612
rect 5359 5596 5375 5604
rect 5382 5602 5409 5604
rect 5418 5602 5639 5612
rect 5382 5592 5639 5602
rect 5668 5604 5718 5612
rect 5668 5595 5684 5604
rect 5277 5584 5328 5592
rect 5375 5584 5639 5592
rect 5665 5592 5684 5595
rect 5691 5592 5718 5604
rect 5665 5584 5718 5592
rect 5293 5576 5294 5584
rect 5309 5576 5322 5584
rect 5293 5568 5309 5576
rect 5290 5561 5309 5564
rect 5290 5552 5312 5561
rect 5263 5542 5312 5552
rect 5263 5536 5293 5542
rect 5312 5537 5317 5542
rect 5235 5520 5309 5536
rect 5327 5528 5357 5584
rect 5392 5574 5600 5584
rect 5635 5580 5680 5584
rect 5683 5583 5684 5584
rect 5699 5583 5712 5584
rect 5418 5544 5607 5574
rect 5433 5541 5607 5544
rect 5426 5538 5607 5541
rect 5235 5518 5248 5520
rect 5263 5518 5297 5520
rect 5235 5502 5309 5518
rect 5336 5514 5349 5528
rect 5364 5514 5380 5530
rect 5426 5525 5437 5538
rect 5219 5480 5220 5496
rect 5235 5480 5248 5502
rect 5263 5480 5293 5502
rect 5336 5498 5398 5514
rect 5426 5507 5437 5523
rect 5442 5518 5452 5538
rect 5462 5518 5476 5538
rect 5479 5525 5488 5538
rect 5504 5525 5513 5538
rect 5442 5507 5476 5518
rect 5479 5507 5488 5523
rect 5504 5507 5513 5523
rect 5520 5518 5530 5538
rect 5540 5518 5554 5538
rect 5555 5525 5566 5538
rect 5520 5507 5554 5518
rect 5555 5507 5566 5523
rect 5612 5514 5628 5530
rect 5635 5528 5665 5580
rect 5699 5576 5700 5583
rect 5684 5568 5700 5576
rect 5671 5536 5684 5555
rect 5699 5536 5729 5552
rect 5671 5520 5745 5536
rect 5671 5518 5684 5520
rect 5699 5518 5733 5520
rect 5336 5496 5349 5498
rect 5364 5496 5398 5498
rect 5336 5480 5398 5496
rect 5442 5491 5458 5494
rect 5520 5491 5550 5502
rect 5598 5498 5644 5514
rect 5671 5502 5745 5518
rect 5598 5496 5632 5498
rect 5597 5480 5644 5496
rect 5671 5480 5684 5502
rect 5699 5480 5729 5502
rect 5756 5480 5757 5496
rect 5772 5480 5785 5640
rect 5815 5536 5828 5640
rect 5873 5618 5874 5628
rect 5889 5618 5902 5628
rect 5873 5614 5902 5618
rect 5907 5614 5937 5640
rect 5955 5626 5971 5628
rect 6043 5626 6096 5640
rect 6044 5624 6108 5626
rect 6151 5624 6166 5640
rect 6215 5637 6245 5640
rect 6215 5634 6251 5637
rect 6181 5626 6197 5628
rect 5955 5614 5970 5618
rect 5873 5612 5970 5614
rect 5998 5612 6166 5624
rect 6182 5614 6197 5618
rect 6215 5615 6254 5634
rect 6273 5628 6280 5629
rect 6279 5621 6280 5628
rect 6263 5618 6264 5621
rect 6279 5618 6292 5621
rect 6215 5614 6245 5615
rect 6254 5614 6260 5615
rect 6263 5614 6292 5618
rect 6182 5613 6292 5614
rect 6182 5612 6298 5613
rect 5857 5604 5908 5612
rect 5857 5592 5882 5604
rect 5889 5592 5908 5604
rect 5939 5604 5989 5612
rect 5939 5596 5955 5604
rect 5962 5602 5989 5604
rect 5998 5602 6219 5612
rect 5962 5592 6219 5602
rect 6248 5604 6298 5612
rect 6248 5595 6264 5604
rect 5857 5584 5908 5592
rect 5955 5584 6219 5592
rect 6245 5592 6264 5595
rect 6271 5592 6298 5604
rect 6245 5584 6298 5592
rect 5873 5576 5874 5584
rect 5889 5576 5902 5584
rect 5873 5568 5889 5576
rect 5870 5561 5889 5564
rect 5870 5552 5892 5561
rect 5843 5542 5892 5552
rect 5843 5536 5873 5542
rect 5892 5537 5897 5542
rect 5815 5520 5889 5536
rect 5907 5528 5937 5584
rect 5972 5574 6180 5584
rect 6215 5580 6260 5584
rect 6263 5583 6264 5584
rect 6279 5583 6292 5584
rect 5998 5544 6187 5574
rect 6013 5541 6187 5544
rect 6006 5538 6187 5541
rect 5815 5518 5828 5520
rect 5843 5518 5877 5520
rect 5815 5502 5889 5518
rect 5916 5514 5929 5528
rect 5944 5514 5960 5530
rect 6006 5525 6017 5538
rect 5799 5480 5800 5496
rect 5815 5480 5828 5502
rect 5843 5480 5873 5502
rect 5916 5498 5978 5514
rect 6006 5507 6017 5523
rect 6022 5518 6032 5538
rect 6042 5518 6056 5538
rect 6059 5525 6068 5538
rect 6084 5525 6093 5538
rect 6022 5507 6056 5518
rect 6059 5507 6068 5523
rect 6084 5507 6093 5523
rect 6100 5518 6110 5538
rect 6120 5518 6134 5538
rect 6135 5525 6146 5538
rect 6100 5507 6134 5518
rect 6135 5507 6146 5523
rect 6192 5514 6208 5530
rect 6215 5528 6245 5580
rect 6279 5576 6280 5583
rect 6264 5568 6280 5576
rect 6251 5536 6264 5555
rect 6279 5536 6309 5552
rect 6251 5520 6325 5536
rect 6251 5518 6264 5520
rect 6279 5518 6313 5520
rect 5916 5496 5929 5498
rect 5944 5496 5978 5498
rect 5916 5480 5978 5496
rect 6022 5491 6038 5494
rect 6100 5491 6130 5502
rect 6178 5498 6224 5514
rect 6251 5502 6325 5518
rect 6178 5496 6212 5498
rect 6177 5480 6224 5496
rect 6251 5480 6264 5502
rect 6279 5480 6309 5502
rect 6336 5480 6337 5496
rect 6352 5480 6365 5640
rect 6395 5536 6408 5640
rect 6453 5618 6454 5628
rect 6469 5618 6482 5628
rect 6453 5614 6482 5618
rect 6487 5614 6517 5640
rect 6535 5626 6551 5628
rect 6623 5626 6676 5640
rect 6624 5624 6688 5626
rect 6731 5624 6746 5640
rect 6795 5637 6825 5640
rect 6795 5634 6831 5637
rect 6761 5626 6777 5628
rect 6535 5614 6550 5618
rect 6453 5612 6550 5614
rect 6578 5612 6746 5624
rect 6762 5614 6777 5618
rect 6795 5615 6834 5634
rect 6853 5628 6860 5629
rect 6859 5621 6860 5628
rect 6843 5618 6844 5621
rect 6859 5618 6872 5621
rect 6795 5614 6825 5615
rect 6834 5614 6840 5615
rect 6843 5614 6872 5618
rect 6762 5613 6872 5614
rect 6762 5612 6878 5613
rect 6437 5604 6488 5612
rect 6437 5592 6462 5604
rect 6469 5592 6488 5604
rect 6519 5604 6569 5612
rect 6519 5596 6535 5604
rect 6542 5602 6569 5604
rect 6578 5602 6799 5612
rect 6542 5592 6799 5602
rect 6828 5604 6878 5612
rect 6828 5595 6844 5604
rect 6437 5584 6488 5592
rect 6535 5584 6799 5592
rect 6825 5592 6844 5595
rect 6851 5592 6878 5604
rect 6825 5584 6878 5592
rect 6453 5576 6454 5584
rect 6469 5576 6482 5584
rect 6453 5568 6469 5576
rect 6450 5561 6469 5564
rect 6450 5552 6472 5561
rect 6423 5542 6472 5552
rect 6423 5536 6453 5542
rect 6472 5537 6477 5542
rect 6395 5520 6469 5536
rect 6487 5528 6517 5584
rect 6552 5574 6760 5584
rect 6795 5580 6840 5584
rect 6843 5583 6844 5584
rect 6859 5583 6872 5584
rect 6578 5544 6767 5574
rect 6593 5541 6767 5544
rect 6586 5538 6767 5541
rect 6395 5518 6408 5520
rect 6423 5518 6457 5520
rect 6395 5502 6469 5518
rect 6496 5514 6509 5528
rect 6524 5514 6540 5530
rect 6586 5525 6597 5538
rect 6379 5480 6380 5496
rect 6395 5480 6408 5502
rect 6423 5480 6453 5502
rect 6496 5498 6558 5514
rect 6586 5507 6597 5523
rect 6602 5518 6612 5538
rect 6622 5518 6636 5538
rect 6639 5525 6648 5538
rect 6664 5525 6673 5538
rect 6602 5507 6636 5518
rect 6639 5507 6648 5523
rect 6664 5507 6673 5523
rect 6680 5518 6690 5538
rect 6700 5518 6714 5538
rect 6715 5525 6726 5538
rect 6680 5507 6714 5518
rect 6715 5507 6726 5523
rect 6772 5514 6788 5530
rect 6795 5528 6825 5580
rect 6859 5576 6860 5583
rect 6844 5568 6860 5576
rect 6831 5536 6844 5555
rect 6859 5536 6889 5552
rect 6831 5520 6905 5536
rect 6831 5518 6844 5520
rect 6859 5518 6893 5520
rect 6496 5496 6509 5498
rect 6524 5496 6558 5498
rect 6496 5480 6558 5496
rect 6602 5491 6618 5494
rect 6680 5491 6710 5502
rect 6758 5498 6804 5514
rect 6831 5502 6905 5518
rect 6758 5496 6792 5498
rect 6757 5480 6804 5496
rect 6831 5480 6844 5502
rect 6859 5480 6889 5502
rect 6916 5480 6917 5496
rect 6932 5480 6945 5640
rect 6975 5536 6988 5640
rect 7033 5618 7034 5628
rect 7049 5618 7062 5628
rect 7033 5614 7062 5618
rect 7067 5614 7097 5640
rect 7115 5626 7131 5628
rect 7203 5626 7256 5640
rect 7204 5624 7268 5626
rect 7311 5624 7326 5640
rect 7375 5637 7405 5640
rect 7375 5634 7411 5637
rect 7341 5626 7357 5628
rect 7115 5614 7130 5618
rect 7033 5612 7130 5614
rect 7158 5612 7326 5624
rect 7342 5614 7357 5618
rect 7375 5615 7414 5634
rect 7433 5628 7440 5629
rect 7439 5621 7440 5628
rect 7423 5618 7424 5621
rect 7439 5618 7452 5621
rect 7375 5614 7405 5615
rect 7414 5614 7420 5615
rect 7423 5614 7452 5618
rect 7342 5613 7452 5614
rect 7342 5612 7458 5613
rect 7017 5604 7068 5612
rect 7017 5592 7042 5604
rect 7049 5592 7068 5604
rect 7099 5604 7149 5612
rect 7099 5596 7115 5604
rect 7122 5602 7149 5604
rect 7158 5602 7379 5612
rect 7122 5592 7379 5602
rect 7408 5604 7458 5612
rect 7408 5595 7424 5604
rect 7017 5584 7068 5592
rect 7115 5584 7379 5592
rect 7405 5592 7424 5595
rect 7431 5592 7458 5604
rect 7405 5584 7458 5592
rect 7033 5576 7034 5584
rect 7049 5576 7062 5584
rect 7033 5568 7049 5576
rect 7030 5561 7049 5564
rect 7030 5552 7052 5561
rect 7003 5542 7052 5552
rect 7003 5536 7033 5542
rect 7052 5537 7057 5542
rect 6975 5520 7049 5536
rect 7067 5528 7097 5584
rect 7132 5574 7340 5584
rect 7375 5580 7420 5584
rect 7423 5583 7424 5584
rect 7439 5583 7452 5584
rect 7158 5544 7347 5574
rect 7173 5541 7347 5544
rect 7166 5538 7347 5541
rect 6975 5518 6988 5520
rect 7003 5518 7037 5520
rect 6975 5502 7049 5518
rect 7076 5514 7089 5528
rect 7104 5514 7120 5530
rect 7166 5525 7177 5538
rect 6959 5480 6960 5496
rect 6975 5480 6988 5502
rect 7003 5480 7033 5502
rect 7076 5498 7138 5514
rect 7166 5507 7177 5523
rect 7182 5518 7192 5538
rect 7202 5518 7216 5538
rect 7219 5525 7228 5538
rect 7244 5525 7253 5538
rect 7182 5507 7216 5518
rect 7219 5507 7228 5523
rect 7244 5507 7253 5523
rect 7260 5518 7270 5538
rect 7280 5518 7294 5538
rect 7295 5525 7306 5538
rect 7260 5507 7294 5518
rect 7295 5507 7306 5523
rect 7352 5514 7368 5530
rect 7375 5528 7405 5580
rect 7439 5576 7440 5583
rect 7424 5568 7440 5576
rect 7411 5536 7424 5555
rect 7439 5536 7469 5552
rect 7411 5520 7485 5536
rect 7411 5518 7424 5520
rect 7439 5518 7473 5520
rect 7076 5496 7089 5498
rect 7104 5496 7138 5498
rect 7076 5480 7138 5496
rect 7182 5491 7198 5494
rect 7260 5491 7290 5502
rect 7338 5498 7384 5514
rect 7411 5502 7485 5518
rect 7338 5496 7372 5498
rect 7337 5480 7384 5496
rect 7411 5480 7424 5502
rect 7439 5480 7469 5502
rect 7496 5480 7497 5496
rect 7512 5480 7525 5640
rect 7555 5536 7568 5640
rect 7613 5618 7614 5628
rect 7629 5618 7642 5628
rect 7613 5614 7642 5618
rect 7647 5614 7677 5640
rect 7695 5626 7711 5628
rect 7783 5626 7836 5640
rect 7784 5624 7848 5626
rect 7891 5624 7906 5640
rect 7955 5637 7985 5640
rect 7955 5634 7991 5637
rect 7921 5626 7937 5628
rect 7695 5614 7710 5618
rect 7613 5612 7710 5614
rect 7738 5612 7906 5624
rect 7922 5614 7937 5618
rect 7955 5615 7994 5634
rect 8013 5628 8020 5629
rect 8019 5621 8020 5628
rect 8003 5618 8004 5621
rect 8019 5618 8032 5621
rect 7955 5614 7985 5615
rect 7994 5614 8000 5615
rect 8003 5614 8032 5618
rect 7922 5613 8032 5614
rect 7922 5612 8038 5613
rect 7597 5604 7648 5612
rect 7597 5592 7622 5604
rect 7629 5592 7648 5604
rect 7679 5604 7729 5612
rect 7679 5596 7695 5604
rect 7702 5602 7729 5604
rect 7738 5602 7959 5612
rect 7702 5592 7959 5602
rect 7988 5604 8038 5612
rect 7988 5595 8004 5604
rect 7597 5584 7648 5592
rect 7695 5584 7959 5592
rect 7985 5592 8004 5595
rect 8011 5592 8038 5604
rect 7985 5584 8038 5592
rect 7613 5576 7614 5584
rect 7629 5576 7642 5584
rect 7613 5568 7629 5576
rect 7610 5561 7629 5564
rect 7610 5552 7632 5561
rect 7583 5542 7632 5552
rect 7583 5536 7613 5542
rect 7632 5537 7637 5542
rect 7555 5520 7629 5536
rect 7647 5528 7677 5584
rect 7712 5574 7920 5584
rect 7955 5580 8000 5584
rect 8003 5583 8004 5584
rect 8019 5583 8032 5584
rect 7738 5544 7927 5574
rect 7753 5541 7927 5544
rect 7746 5538 7927 5541
rect 7555 5518 7568 5520
rect 7583 5518 7617 5520
rect 7555 5502 7629 5518
rect 7656 5514 7669 5528
rect 7684 5514 7700 5530
rect 7746 5525 7757 5538
rect 7539 5480 7540 5496
rect 7555 5480 7568 5502
rect 7583 5480 7613 5502
rect 7656 5498 7718 5514
rect 7746 5507 7757 5523
rect 7762 5518 7772 5538
rect 7782 5518 7796 5538
rect 7799 5525 7808 5538
rect 7824 5525 7833 5538
rect 7762 5507 7796 5518
rect 7799 5507 7808 5523
rect 7824 5507 7833 5523
rect 7840 5518 7850 5538
rect 7860 5518 7874 5538
rect 7875 5525 7886 5538
rect 7840 5507 7874 5518
rect 7875 5507 7886 5523
rect 7932 5514 7948 5530
rect 7955 5528 7985 5580
rect 8019 5576 8020 5583
rect 8004 5568 8020 5576
rect 7991 5536 8004 5555
rect 8019 5536 8049 5552
rect 7991 5520 8065 5536
rect 7991 5518 8004 5520
rect 8019 5518 8053 5520
rect 7656 5496 7669 5498
rect 7684 5496 7718 5498
rect 7656 5480 7718 5496
rect 7762 5491 7778 5494
rect 7840 5491 7870 5502
rect 7918 5498 7964 5514
rect 7991 5502 8065 5518
rect 7918 5496 7952 5498
rect 7917 5480 7964 5496
rect 7991 5480 8004 5502
rect 8019 5480 8049 5502
rect 8076 5480 8077 5496
rect 8092 5480 8105 5640
rect 8135 5536 8148 5640
rect 8193 5618 8194 5628
rect 8209 5618 8222 5628
rect 8193 5614 8222 5618
rect 8227 5614 8257 5640
rect 8275 5626 8291 5628
rect 8363 5626 8416 5640
rect 8364 5624 8428 5626
rect 8471 5624 8486 5640
rect 8535 5637 8565 5640
rect 8535 5634 8571 5637
rect 8501 5626 8517 5628
rect 8275 5614 8290 5618
rect 8193 5612 8290 5614
rect 8318 5612 8486 5624
rect 8502 5614 8517 5618
rect 8535 5615 8574 5634
rect 8593 5628 8600 5629
rect 8599 5621 8600 5628
rect 8583 5618 8584 5621
rect 8599 5618 8612 5621
rect 8535 5614 8565 5615
rect 8574 5614 8580 5615
rect 8583 5614 8612 5618
rect 8502 5613 8612 5614
rect 8502 5612 8618 5613
rect 8177 5604 8228 5612
rect 8177 5592 8202 5604
rect 8209 5592 8228 5604
rect 8259 5604 8309 5612
rect 8259 5596 8275 5604
rect 8282 5602 8309 5604
rect 8318 5602 8539 5612
rect 8282 5592 8539 5602
rect 8568 5604 8618 5612
rect 8568 5595 8584 5604
rect 8177 5584 8228 5592
rect 8275 5584 8539 5592
rect 8565 5592 8584 5595
rect 8591 5592 8618 5604
rect 8565 5584 8618 5592
rect 8193 5576 8194 5584
rect 8209 5576 8222 5584
rect 8193 5568 8209 5576
rect 8190 5561 8209 5564
rect 8190 5552 8212 5561
rect 8163 5542 8212 5552
rect 8163 5536 8193 5542
rect 8212 5537 8217 5542
rect 8135 5520 8209 5536
rect 8227 5528 8257 5584
rect 8292 5574 8500 5584
rect 8535 5580 8580 5584
rect 8583 5583 8584 5584
rect 8599 5583 8612 5584
rect 8318 5544 8507 5574
rect 8333 5541 8507 5544
rect 8326 5538 8507 5541
rect 8135 5518 8148 5520
rect 8163 5518 8197 5520
rect 8135 5502 8209 5518
rect 8236 5514 8249 5528
rect 8264 5514 8280 5530
rect 8326 5525 8337 5538
rect 8119 5480 8120 5496
rect 8135 5480 8148 5502
rect 8163 5480 8193 5502
rect 8236 5498 8298 5514
rect 8326 5507 8337 5523
rect 8342 5518 8352 5538
rect 8362 5518 8376 5538
rect 8379 5525 8388 5538
rect 8404 5525 8413 5538
rect 8342 5507 8376 5518
rect 8379 5507 8388 5523
rect 8404 5507 8413 5523
rect 8420 5518 8430 5538
rect 8440 5518 8454 5538
rect 8455 5525 8466 5538
rect 8420 5507 8454 5518
rect 8455 5507 8466 5523
rect 8512 5514 8528 5530
rect 8535 5528 8565 5580
rect 8599 5576 8600 5583
rect 8584 5568 8600 5576
rect 8571 5536 8584 5555
rect 8599 5536 8629 5552
rect 8571 5520 8645 5536
rect 8571 5518 8584 5520
rect 8599 5518 8633 5520
rect 8236 5496 8249 5498
rect 8264 5496 8298 5498
rect 8236 5480 8298 5496
rect 8342 5491 8358 5494
rect 8420 5491 8450 5502
rect 8498 5498 8544 5514
rect 8571 5502 8645 5518
rect 8498 5496 8532 5498
rect 8497 5480 8544 5496
rect 8571 5480 8584 5502
rect 8599 5480 8629 5502
rect 8656 5480 8657 5496
rect 8672 5480 8685 5640
rect 8715 5536 8728 5640
rect 8773 5618 8774 5628
rect 8789 5618 8802 5628
rect 8773 5614 8802 5618
rect 8807 5614 8837 5640
rect 8855 5626 8871 5628
rect 8943 5626 8996 5640
rect 8944 5624 9008 5626
rect 9051 5624 9066 5640
rect 9115 5637 9145 5640
rect 9115 5634 9151 5637
rect 9081 5626 9097 5628
rect 8855 5614 8870 5618
rect 8773 5612 8870 5614
rect 8898 5612 9066 5624
rect 9082 5614 9097 5618
rect 9115 5615 9154 5634
rect 9173 5628 9180 5629
rect 9179 5621 9180 5628
rect 9163 5618 9164 5621
rect 9179 5618 9192 5621
rect 9115 5614 9145 5615
rect 9154 5614 9160 5615
rect 9163 5614 9192 5618
rect 9082 5613 9192 5614
rect 9082 5612 9198 5613
rect 8757 5604 8808 5612
rect 8757 5592 8782 5604
rect 8789 5592 8808 5604
rect 8839 5604 8889 5612
rect 8839 5596 8855 5604
rect 8862 5602 8889 5604
rect 8898 5602 9119 5612
rect 8862 5592 9119 5602
rect 9148 5604 9198 5612
rect 9148 5595 9164 5604
rect 8757 5584 8808 5592
rect 8855 5584 9119 5592
rect 9145 5592 9164 5595
rect 9171 5592 9198 5604
rect 9145 5584 9198 5592
rect 8773 5576 8774 5584
rect 8789 5576 8802 5584
rect 8773 5568 8789 5576
rect 8770 5561 8789 5564
rect 8770 5552 8792 5561
rect 8743 5542 8792 5552
rect 8743 5536 8773 5542
rect 8792 5537 8797 5542
rect 8715 5520 8789 5536
rect 8807 5528 8837 5584
rect 8872 5574 9080 5584
rect 9115 5580 9160 5584
rect 9163 5583 9164 5584
rect 9179 5583 9192 5584
rect 8898 5544 9087 5574
rect 8913 5541 9087 5544
rect 8906 5538 9087 5541
rect 8715 5518 8728 5520
rect 8743 5518 8777 5520
rect 8715 5502 8789 5518
rect 8816 5514 8829 5528
rect 8844 5514 8860 5530
rect 8906 5525 8917 5538
rect 8699 5480 8700 5496
rect 8715 5480 8728 5502
rect 8743 5480 8773 5502
rect 8816 5498 8878 5514
rect 8906 5507 8917 5523
rect 8922 5518 8932 5538
rect 8942 5518 8956 5538
rect 8959 5525 8968 5538
rect 8984 5525 8993 5538
rect 8922 5507 8956 5518
rect 8959 5507 8968 5523
rect 8984 5507 8993 5523
rect 9000 5518 9010 5538
rect 9020 5518 9034 5538
rect 9035 5525 9046 5538
rect 9000 5507 9034 5518
rect 9035 5507 9046 5523
rect 9092 5514 9108 5530
rect 9115 5528 9145 5580
rect 9179 5576 9180 5583
rect 9164 5568 9180 5576
rect 9151 5536 9164 5555
rect 9179 5536 9209 5552
rect 9151 5520 9225 5536
rect 9151 5518 9164 5520
rect 9179 5518 9213 5520
rect 8816 5496 8829 5498
rect 8844 5496 8878 5498
rect 8816 5480 8878 5496
rect 8922 5491 8938 5494
rect 9000 5491 9030 5502
rect 9078 5498 9124 5514
rect 9151 5502 9225 5518
rect 9078 5496 9112 5498
rect 9077 5480 9124 5496
rect 9151 5480 9164 5502
rect 9179 5480 9209 5502
rect 9236 5480 9237 5496
rect 9252 5480 9265 5640
rect -7 5472 34 5480
rect -7 5446 8 5472
rect 15 5446 34 5472
rect 98 5468 160 5480
rect 172 5468 247 5480
rect 305 5468 380 5480
rect 392 5468 423 5480
rect 429 5468 464 5480
rect 98 5466 260 5468
rect -7 5438 34 5446
rect 116 5442 129 5466
rect 144 5464 159 5466
rect -1 5428 0 5438
rect 15 5428 28 5438
rect 43 5428 73 5442
rect 116 5428 159 5442
rect 183 5439 190 5446
rect 193 5442 260 5466
rect 292 5466 464 5468
rect 262 5444 290 5448
rect 292 5444 372 5466
rect 393 5464 408 5466
rect 262 5442 372 5444
rect 193 5438 372 5442
rect 166 5428 196 5438
rect 198 5428 351 5438
rect 359 5428 389 5438
rect 393 5428 423 5442
rect 451 5428 464 5466
rect 536 5472 571 5480
rect 536 5446 537 5472
rect 544 5446 571 5472
rect 479 5428 509 5442
rect 536 5438 571 5446
rect 573 5472 614 5480
rect 573 5446 588 5472
rect 595 5446 614 5472
rect 678 5468 740 5480
rect 752 5468 827 5480
rect 885 5468 960 5480
rect 972 5468 1003 5480
rect 1009 5468 1044 5480
rect 678 5466 840 5468
rect 573 5438 614 5446
rect 696 5442 709 5466
rect 724 5464 739 5466
rect 536 5428 537 5438
rect 552 5428 565 5438
rect 579 5428 580 5438
rect 595 5428 608 5438
rect 623 5428 653 5442
rect 696 5428 739 5442
rect 763 5439 770 5446
rect 773 5442 840 5466
rect 872 5466 1044 5468
rect 842 5444 870 5448
rect 872 5444 952 5466
rect 973 5464 988 5466
rect 842 5442 952 5444
rect 773 5438 952 5442
rect 746 5428 776 5438
rect 778 5428 931 5438
rect 939 5428 969 5438
rect 973 5428 1003 5442
rect 1031 5428 1044 5466
rect 1116 5472 1151 5480
rect 1116 5446 1117 5472
rect 1124 5446 1151 5472
rect 1059 5428 1089 5442
rect 1116 5438 1151 5446
rect 1153 5472 1194 5480
rect 1153 5446 1168 5472
rect 1175 5446 1194 5472
rect 1258 5468 1320 5480
rect 1332 5468 1407 5480
rect 1465 5468 1540 5480
rect 1552 5468 1583 5480
rect 1589 5468 1624 5480
rect 1258 5466 1420 5468
rect 1153 5438 1194 5446
rect 1276 5442 1289 5466
rect 1304 5464 1319 5466
rect 1116 5428 1117 5438
rect 1132 5428 1145 5438
rect 1159 5428 1160 5438
rect 1175 5428 1188 5438
rect 1203 5428 1233 5442
rect 1276 5428 1319 5442
rect 1343 5439 1350 5446
rect 1353 5442 1420 5466
rect 1452 5466 1624 5468
rect 1422 5444 1450 5448
rect 1452 5444 1532 5466
rect 1553 5464 1568 5466
rect 1422 5442 1532 5444
rect 1353 5438 1532 5442
rect 1326 5428 1356 5438
rect 1358 5428 1511 5438
rect 1519 5428 1549 5438
rect 1553 5428 1583 5442
rect 1611 5428 1624 5466
rect 1696 5472 1731 5480
rect 1696 5446 1697 5472
rect 1704 5446 1731 5472
rect 1639 5428 1669 5442
rect 1696 5438 1731 5446
rect 1733 5472 1774 5480
rect 1733 5446 1748 5472
rect 1755 5446 1774 5472
rect 1838 5468 1900 5480
rect 1912 5468 1987 5480
rect 2045 5468 2120 5480
rect 2132 5468 2163 5480
rect 2169 5468 2204 5480
rect 1838 5466 2000 5468
rect 1733 5438 1774 5446
rect 1856 5442 1869 5466
rect 1884 5464 1899 5466
rect 1696 5428 1697 5438
rect 1712 5428 1725 5438
rect 1739 5428 1740 5438
rect 1755 5428 1768 5438
rect 1783 5428 1813 5442
rect 1856 5428 1899 5442
rect 1923 5439 1930 5446
rect 1933 5442 2000 5466
rect 2032 5466 2204 5468
rect 2002 5444 2030 5448
rect 2032 5444 2112 5466
rect 2133 5464 2148 5466
rect 2002 5442 2112 5444
rect 1933 5438 2112 5442
rect 1906 5428 1936 5438
rect 1938 5428 2091 5438
rect 2099 5428 2129 5438
rect 2133 5428 2163 5442
rect 2191 5428 2204 5466
rect 2276 5472 2311 5480
rect 2276 5446 2277 5472
rect 2284 5446 2311 5472
rect 2219 5428 2249 5442
rect 2276 5438 2311 5446
rect 2313 5472 2354 5480
rect 2313 5446 2328 5472
rect 2335 5446 2354 5472
rect 2418 5468 2480 5480
rect 2492 5468 2567 5480
rect 2625 5468 2700 5480
rect 2712 5468 2743 5480
rect 2749 5468 2784 5480
rect 2418 5466 2580 5468
rect 2313 5438 2354 5446
rect 2436 5442 2449 5466
rect 2464 5464 2479 5466
rect 2276 5428 2277 5438
rect 2292 5428 2305 5438
rect 2319 5428 2320 5438
rect 2335 5428 2348 5438
rect 2363 5428 2393 5442
rect 2436 5428 2479 5442
rect 2503 5439 2510 5446
rect 2513 5442 2580 5466
rect 2612 5466 2784 5468
rect 2582 5444 2610 5448
rect 2612 5444 2692 5466
rect 2713 5464 2728 5466
rect 2582 5442 2692 5444
rect 2513 5438 2692 5442
rect 2486 5428 2516 5438
rect 2518 5428 2671 5438
rect 2679 5428 2709 5438
rect 2713 5428 2743 5442
rect 2771 5428 2784 5466
rect 2856 5472 2891 5480
rect 2856 5446 2857 5472
rect 2864 5446 2891 5472
rect 2799 5428 2829 5442
rect 2856 5438 2891 5446
rect 2893 5472 2934 5480
rect 2893 5446 2908 5472
rect 2915 5446 2934 5472
rect 2998 5468 3060 5480
rect 3072 5468 3147 5480
rect 3205 5468 3280 5480
rect 3292 5468 3323 5480
rect 3329 5468 3364 5480
rect 2998 5466 3160 5468
rect 2893 5438 2934 5446
rect 3016 5442 3029 5466
rect 3044 5464 3059 5466
rect 2856 5428 2857 5438
rect 2872 5428 2885 5438
rect 2899 5428 2900 5438
rect 2915 5428 2928 5438
rect 2943 5428 2973 5442
rect 3016 5428 3059 5442
rect 3083 5439 3090 5446
rect 3093 5442 3160 5466
rect 3192 5466 3364 5468
rect 3162 5444 3190 5448
rect 3192 5444 3272 5466
rect 3293 5464 3308 5466
rect 3162 5442 3272 5444
rect 3093 5438 3272 5442
rect 3066 5428 3096 5438
rect 3098 5428 3251 5438
rect 3259 5428 3289 5438
rect 3293 5428 3323 5442
rect 3351 5428 3364 5466
rect 3436 5472 3471 5480
rect 3436 5446 3437 5472
rect 3444 5446 3471 5472
rect 3379 5428 3409 5442
rect 3436 5438 3471 5446
rect 3473 5472 3514 5480
rect 3473 5446 3488 5472
rect 3495 5446 3514 5472
rect 3578 5468 3640 5480
rect 3652 5468 3727 5480
rect 3785 5468 3860 5480
rect 3872 5468 3903 5480
rect 3909 5468 3944 5480
rect 3578 5466 3740 5468
rect 3473 5438 3514 5446
rect 3596 5442 3609 5466
rect 3624 5464 3639 5466
rect 3436 5428 3437 5438
rect 3452 5428 3465 5438
rect 3479 5428 3480 5438
rect 3495 5428 3508 5438
rect 3523 5428 3553 5442
rect 3596 5428 3639 5442
rect 3663 5439 3670 5446
rect 3673 5442 3740 5466
rect 3772 5466 3944 5468
rect 3742 5444 3770 5448
rect 3772 5444 3852 5466
rect 3873 5464 3888 5466
rect 3742 5442 3852 5444
rect 3673 5438 3852 5442
rect 3646 5428 3676 5438
rect 3678 5428 3831 5438
rect 3839 5428 3869 5438
rect 3873 5428 3903 5442
rect 3931 5428 3944 5466
rect 4016 5472 4051 5480
rect 4016 5446 4017 5472
rect 4024 5446 4051 5472
rect 3959 5428 3989 5442
rect 4016 5438 4051 5446
rect 4053 5472 4094 5480
rect 4053 5446 4068 5472
rect 4075 5446 4094 5472
rect 4158 5468 4220 5480
rect 4232 5468 4307 5480
rect 4365 5468 4440 5480
rect 4452 5468 4483 5480
rect 4489 5468 4524 5480
rect 4158 5466 4320 5468
rect 4053 5438 4094 5446
rect 4176 5442 4189 5466
rect 4204 5464 4219 5466
rect 4016 5428 4017 5438
rect 4032 5428 4045 5438
rect 4059 5428 4060 5438
rect 4075 5428 4088 5438
rect 4103 5428 4133 5442
rect 4176 5428 4219 5442
rect 4243 5439 4250 5446
rect 4253 5442 4320 5466
rect 4352 5466 4524 5468
rect 4322 5444 4350 5448
rect 4352 5444 4432 5466
rect 4453 5464 4468 5466
rect 4322 5442 4432 5444
rect 4253 5438 4432 5442
rect 4226 5428 4256 5438
rect 4258 5428 4411 5438
rect 4419 5428 4449 5438
rect 4453 5428 4483 5442
rect 4511 5428 4524 5466
rect 4596 5472 4631 5480
rect 4596 5446 4597 5472
rect 4604 5446 4631 5472
rect 4539 5428 4569 5442
rect 4596 5438 4631 5446
rect 4633 5472 4674 5480
rect 4633 5446 4648 5472
rect 4655 5446 4674 5472
rect 4738 5468 4800 5480
rect 4812 5468 4887 5480
rect 4945 5468 5020 5480
rect 5032 5468 5063 5480
rect 5069 5468 5104 5480
rect 4738 5466 4900 5468
rect 4633 5438 4674 5446
rect 4756 5442 4769 5466
rect 4784 5464 4799 5466
rect 4596 5428 4597 5438
rect 4612 5428 4625 5438
rect 4639 5428 4640 5438
rect 4655 5428 4668 5438
rect 4683 5428 4713 5442
rect 4756 5428 4799 5442
rect 4823 5439 4830 5446
rect 4833 5442 4900 5466
rect 4932 5466 5104 5468
rect 4902 5444 4930 5448
rect 4932 5444 5012 5466
rect 5033 5464 5048 5466
rect 4902 5442 5012 5444
rect 4833 5438 5012 5442
rect 4806 5428 4836 5438
rect 4838 5428 4991 5438
rect 4999 5428 5029 5438
rect 5033 5428 5063 5442
rect 5091 5428 5104 5466
rect 5176 5472 5211 5480
rect 5176 5446 5177 5472
rect 5184 5446 5211 5472
rect 5119 5428 5149 5442
rect 5176 5438 5211 5446
rect 5213 5472 5254 5480
rect 5213 5446 5228 5472
rect 5235 5446 5254 5472
rect 5318 5468 5380 5480
rect 5392 5468 5467 5480
rect 5525 5468 5600 5480
rect 5612 5468 5643 5480
rect 5649 5468 5684 5480
rect 5318 5466 5480 5468
rect 5213 5438 5254 5446
rect 5336 5442 5349 5466
rect 5364 5464 5379 5466
rect 5176 5428 5177 5438
rect 5192 5428 5205 5438
rect 5219 5428 5220 5438
rect 5235 5428 5248 5438
rect 5263 5428 5293 5442
rect 5336 5428 5379 5442
rect 5403 5439 5410 5446
rect 5413 5442 5480 5466
rect 5512 5466 5684 5468
rect 5482 5444 5510 5448
rect 5512 5444 5592 5466
rect 5613 5464 5628 5466
rect 5482 5442 5592 5444
rect 5413 5438 5592 5442
rect 5386 5428 5416 5438
rect 5418 5428 5571 5438
rect 5579 5428 5609 5438
rect 5613 5428 5643 5442
rect 5671 5428 5684 5466
rect 5756 5472 5791 5480
rect 5756 5446 5757 5472
rect 5764 5446 5791 5472
rect 5699 5428 5729 5442
rect 5756 5438 5791 5446
rect 5793 5472 5834 5480
rect 5793 5446 5808 5472
rect 5815 5446 5834 5472
rect 5898 5468 5960 5480
rect 5972 5468 6047 5480
rect 6105 5468 6180 5480
rect 6192 5468 6223 5480
rect 6229 5468 6264 5480
rect 5898 5466 6060 5468
rect 5793 5438 5834 5446
rect 5916 5442 5929 5466
rect 5944 5464 5959 5466
rect 5756 5428 5757 5438
rect 5772 5428 5785 5438
rect 5799 5428 5800 5438
rect 5815 5428 5828 5438
rect 5843 5428 5873 5442
rect 5916 5428 5959 5442
rect 5983 5439 5990 5446
rect 5993 5442 6060 5466
rect 6092 5466 6264 5468
rect 6062 5444 6090 5448
rect 6092 5444 6172 5466
rect 6193 5464 6208 5466
rect 6062 5442 6172 5444
rect 5993 5438 6172 5442
rect 5966 5428 5996 5438
rect 5998 5428 6151 5438
rect 6159 5428 6189 5438
rect 6193 5428 6223 5442
rect 6251 5428 6264 5466
rect 6336 5472 6371 5480
rect 6336 5446 6337 5472
rect 6344 5446 6371 5472
rect 6279 5428 6309 5442
rect 6336 5438 6371 5446
rect 6373 5472 6414 5480
rect 6373 5446 6388 5472
rect 6395 5446 6414 5472
rect 6478 5468 6540 5480
rect 6552 5468 6627 5480
rect 6685 5468 6760 5480
rect 6772 5468 6803 5480
rect 6809 5468 6844 5480
rect 6478 5466 6640 5468
rect 6373 5438 6414 5446
rect 6496 5442 6509 5466
rect 6524 5464 6539 5466
rect 6336 5428 6337 5438
rect 6352 5428 6365 5438
rect 6379 5428 6380 5438
rect 6395 5428 6408 5438
rect 6423 5428 6453 5442
rect 6496 5428 6539 5442
rect 6563 5439 6570 5446
rect 6573 5442 6640 5466
rect 6672 5466 6844 5468
rect 6642 5444 6670 5448
rect 6672 5444 6752 5466
rect 6773 5464 6788 5466
rect 6642 5442 6752 5444
rect 6573 5438 6752 5442
rect 6546 5428 6576 5438
rect 6578 5428 6731 5438
rect 6739 5428 6769 5438
rect 6773 5428 6803 5442
rect 6831 5428 6844 5466
rect 6916 5472 6951 5480
rect 6916 5446 6917 5472
rect 6924 5446 6951 5472
rect 6859 5428 6889 5442
rect 6916 5438 6951 5446
rect 6953 5472 6994 5480
rect 6953 5446 6968 5472
rect 6975 5446 6994 5472
rect 7058 5468 7120 5480
rect 7132 5468 7207 5480
rect 7265 5468 7340 5480
rect 7352 5468 7383 5480
rect 7389 5468 7424 5480
rect 7058 5466 7220 5468
rect 6953 5438 6994 5446
rect 7076 5442 7089 5466
rect 7104 5464 7119 5466
rect 6916 5428 6917 5438
rect 6932 5428 6945 5438
rect 6959 5428 6960 5438
rect 6975 5428 6988 5438
rect 7003 5428 7033 5442
rect 7076 5428 7119 5442
rect 7143 5439 7150 5446
rect 7153 5442 7220 5466
rect 7252 5466 7424 5468
rect 7222 5444 7250 5448
rect 7252 5444 7332 5466
rect 7353 5464 7368 5466
rect 7222 5442 7332 5444
rect 7153 5438 7332 5442
rect 7126 5428 7156 5438
rect 7158 5428 7311 5438
rect 7319 5428 7349 5438
rect 7353 5428 7383 5442
rect 7411 5428 7424 5466
rect 7496 5472 7531 5480
rect 7496 5446 7497 5472
rect 7504 5446 7531 5472
rect 7439 5428 7469 5442
rect 7496 5438 7531 5446
rect 7533 5472 7574 5480
rect 7533 5446 7548 5472
rect 7555 5446 7574 5472
rect 7638 5468 7700 5480
rect 7712 5468 7787 5480
rect 7845 5468 7920 5480
rect 7932 5468 7963 5480
rect 7969 5468 8004 5480
rect 7638 5466 7800 5468
rect 7533 5438 7574 5446
rect 7656 5442 7669 5466
rect 7684 5464 7699 5466
rect 7496 5428 7497 5438
rect 7512 5428 7525 5438
rect 7539 5428 7540 5438
rect 7555 5428 7568 5438
rect 7583 5428 7613 5442
rect 7656 5428 7699 5442
rect 7723 5439 7730 5446
rect 7733 5442 7800 5466
rect 7832 5466 8004 5468
rect 7802 5444 7830 5448
rect 7832 5444 7912 5466
rect 7933 5464 7948 5466
rect 7802 5442 7912 5444
rect 7733 5438 7912 5442
rect 7706 5428 7736 5438
rect 7738 5428 7891 5438
rect 7899 5428 7929 5438
rect 7933 5428 7963 5442
rect 7991 5428 8004 5466
rect 8076 5472 8111 5480
rect 8076 5446 8077 5472
rect 8084 5446 8111 5472
rect 8019 5428 8049 5442
rect 8076 5438 8111 5446
rect 8113 5472 8154 5480
rect 8113 5446 8128 5472
rect 8135 5446 8154 5472
rect 8218 5468 8280 5480
rect 8292 5468 8367 5480
rect 8425 5468 8500 5480
rect 8512 5468 8543 5480
rect 8549 5468 8584 5480
rect 8218 5466 8380 5468
rect 8113 5438 8154 5446
rect 8236 5442 8249 5466
rect 8264 5464 8279 5466
rect 8076 5428 8077 5438
rect 8092 5428 8105 5438
rect 8119 5428 8120 5438
rect 8135 5428 8148 5438
rect 8163 5428 8193 5442
rect 8236 5428 8279 5442
rect 8303 5439 8310 5446
rect 8313 5442 8380 5466
rect 8412 5466 8584 5468
rect 8382 5444 8410 5448
rect 8412 5444 8492 5466
rect 8513 5464 8528 5466
rect 8382 5442 8492 5444
rect 8313 5438 8492 5442
rect 8286 5428 8316 5438
rect 8318 5428 8471 5438
rect 8479 5428 8509 5438
rect 8513 5428 8543 5442
rect 8571 5428 8584 5466
rect 8656 5472 8691 5480
rect 8656 5446 8657 5472
rect 8664 5446 8691 5472
rect 8599 5428 8629 5442
rect 8656 5438 8691 5446
rect 8693 5472 8734 5480
rect 8693 5446 8708 5472
rect 8715 5446 8734 5472
rect 8798 5468 8860 5480
rect 8872 5468 8947 5480
rect 9005 5468 9080 5480
rect 9092 5468 9123 5480
rect 9129 5468 9164 5480
rect 8798 5466 8960 5468
rect 8693 5438 8734 5446
rect 8816 5442 8829 5466
rect 8844 5464 8859 5466
rect 8656 5428 8657 5438
rect 8672 5428 8685 5438
rect 8699 5428 8700 5438
rect 8715 5428 8728 5438
rect 8743 5428 8773 5442
rect 8816 5428 8859 5442
rect 8883 5439 8890 5446
rect 8893 5442 8960 5466
rect 8992 5466 9164 5468
rect 8962 5444 8990 5448
rect 8992 5444 9072 5466
rect 9093 5464 9108 5466
rect 8962 5442 9072 5444
rect 8893 5438 9072 5442
rect 8866 5428 8896 5438
rect 8898 5428 9051 5438
rect 9059 5428 9089 5438
rect 9093 5428 9123 5442
rect 9151 5428 9164 5466
rect 9236 5472 9271 5480
rect 9236 5446 9237 5472
rect 9244 5446 9271 5472
rect 9179 5428 9209 5442
rect 9236 5438 9271 5446
rect 9236 5428 9237 5438
rect 9252 5428 9265 5438
rect -1 5422 9265 5428
rect 0 5414 9265 5422
rect 15 5384 28 5414
rect 43 5396 73 5414
rect 116 5400 130 5414
rect 166 5400 386 5414
rect 117 5398 130 5400
rect 83 5386 98 5398
rect 80 5384 102 5386
rect 107 5384 137 5398
rect 198 5396 351 5400
rect 180 5384 372 5396
rect 415 5384 445 5398
rect 451 5384 464 5414
rect 479 5396 509 5414
rect 552 5384 565 5414
rect 595 5384 608 5414
rect 623 5396 653 5414
rect 696 5400 710 5414
rect 746 5400 966 5414
rect 697 5398 710 5400
rect 663 5386 678 5398
rect 660 5384 682 5386
rect 687 5384 717 5398
rect 778 5396 931 5400
rect 760 5384 952 5396
rect 995 5384 1025 5398
rect 1031 5384 1044 5414
rect 1059 5396 1089 5414
rect 1132 5384 1145 5414
rect 1175 5384 1188 5414
rect 1203 5396 1233 5414
rect 1276 5400 1290 5414
rect 1326 5400 1546 5414
rect 1277 5398 1290 5400
rect 1243 5386 1258 5398
rect 1240 5384 1262 5386
rect 1267 5384 1297 5398
rect 1358 5396 1511 5400
rect 1340 5384 1532 5396
rect 1575 5384 1605 5398
rect 1611 5384 1624 5414
rect 1639 5396 1669 5414
rect 1712 5384 1725 5414
rect 1755 5384 1768 5414
rect 1783 5396 1813 5414
rect 1856 5400 1870 5414
rect 1906 5400 2126 5414
rect 1857 5398 1870 5400
rect 1823 5386 1838 5398
rect 1820 5384 1842 5386
rect 1847 5384 1877 5398
rect 1938 5396 2091 5400
rect 1920 5384 2112 5396
rect 2155 5384 2185 5398
rect 2191 5384 2204 5414
rect 2219 5396 2249 5414
rect 2292 5384 2305 5414
rect 2335 5384 2348 5414
rect 2363 5396 2393 5414
rect 2436 5400 2450 5414
rect 2486 5400 2706 5414
rect 2437 5398 2450 5400
rect 2403 5386 2418 5398
rect 2400 5384 2422 5386
rect 2427 5384 2457 5398
rect 2518 5396 2671 5400
rect 2500 5384 2692 5396
rect 2735 5384 2765 5398
rect 2771 5384 2784 5414
rect 2799 5396 2829 5414
rect 2872 5384 2885 5414
rect 2915 5384 2928 5414
rect 2943 5396 2973 5414
rect 3016 5400 3030 5414
rect 3066 5400 3286 5414
rect 3017 5398 3030 5400
rect 2983 5386 2998 5398
rect 2980 5384 3002 5386
rect 3007 5384 3037 5398
rect 3098 5396 3251 5400
rect 3080 5384 3272 5396
rect 3315 5384 3345 5398
rect 3351 5384 3364 5414
rect 3379 5396 3409 5414
rect 3452 5384 3465 5414
rect 3495 5384 3508 5414
rect 3523 5396 3553 5414
rect 3596 5400 3610 5414
rect 3646 5400 3866 5414
rect 3597 5398 3610 5400
rect 3563 5386 3578 5398
rect 3560 5384 3582 5386
rect 3587 5384 3617 5398
rect 3678 5396 3831 5400
rect 3660 5384 3852 5396
rect 3895 5384 3925 5398
rect 3931 5384 3944 5414
rect 3959 5396 3989 5414
rect 4032 5384 4045 5414
rect 4075 5384 4088 5414
rect 4103 5396 4133 5414
rect 4176 5400 4190 5414
rect 4226 5400 4446 5414
rect 4177 5398 4190 5400
rect 4143 5386 4158 5398
rect 4140 5384 4162 5386
rect 4167 5384 4197 5398
rect 4258 5396 4411 5400
rect 4240 5384 4432 5396
rect 4475 5384 4505 5398
rect 4511 5384 4524 5414
rect 4539 5396 4569 5414
rect 4612 5384 4625 5414
rect 4655 5384 4668 5414
rect 4683 5396 4713 5414
rect 4756 5400 4770 5414
rect 4806 5400 5026 5414
rect 4757 5398 4770 5400
rect 4723 5386 4738 5398
rect 4720 5384 4742 5386
rect 4747 5384 4777 5398
rect 4838 5396 4991 5400
rect 4820 5384 5012 5396
rect 5055 5384 5085 5398
rect 5091 5384 5104 5414
rect 5119 5396 5149 5414
rect 5192 5384 5205 5414
rect 5235 5384 5248 5414
rect 5263 5396 5293 5414
rect 5336 5400 5350 5414
rect 5386 5400 5606 5414
rect 5337 5398 5350 5400
rect 5303 5386 5318 5398
rect 5300 5384 5322 5386
rect 5327 5384 5357 5398
rect 5418 5396 5571 5400
rect 5400 5384 5592 5396
rect 5635 5384 5665 5398
rect 5671 5384 5684 5414
rect 5699 5396 5729 5414
rect 5772 5384 5785 5414
rect 5815 5384 5828 5414
rect 5843 5396 5873 5414
rect 5916 5400 5930 5414
rect 5966 5400 6186 5414
rect 5917 5398 5930 5400
rect 5883 5386 5898 5398
rect 5880 5384 5902 5386
rect 5907 5384 5937 5398
rect 5998 5396 6151 5400
rect 5980 5384 6172 5396
rect 6215 5384 6245 5398
rect 6251 5384 6264 5414
rect 6279 5396 6309 5414
rect 6352 5384 6365 5414
rect 6395 5384 6408 5414
rect 6423 5396 6453 5414
rect 6496 5400 6510 5414
rect 6546 5400 6766 5414
rect 6497 5398 6510 5400
rect 6463 5386 6478 5398
rect 6460 5384 6482 5386
rect 6487 5384 6517 5398
rect 6578 5396 6731 5400
rect 6560 5384 6752 5396
rect 6795 5384 6825 5398
rect 6831 5384 6844 5414
rect 6859 5396 6889 5414
rect 6932 5384 6945 5414
rect 6975 5384 6988 5414
rect 7003 5396 7033 5414
rect 7076 5400 7090 5414
rect 7126 5400 7346 5414
rect 7077 5398 7090 5400
rect 7043 5386 7058 5398
rect 7040 5384 7062 5386
rect 7067 5384 7097 5398
rect 7158 5396 7311 5400
rect 7140 5384 7332 5396
rect 7375 5384 7405 5398
rect 7411 5384 7424 5414
rect 7439 5396 7469 5414
rect 7512 5384 7525 5414
rect 7555 5384 7568 5414
rect 7583 5396 7613 5414
rect 7656 5400 7670 5414
rect 7706 5400 7926 5414
rect 7657 5398 7670 5400
rect 7623 5386 7638 5398
rect 7620 5384 7642 5386
rect 7647 5384 7677 5398
rect 7738 5396 7891 5400
rect 7720 5384 7912 5396
rect 7955 5384 7985 5398
rect 7991 5384 8004 5414
rect 8019 5396 8049 5414
rect 8092 5384 8105 5414
rect 8135 5384 8148 5414
rect 8163 5396 8193 5414
rect 8236 5400 8250 5414
rect 8286 5400 8506 5414
rect 8237 5398 8250 5400
rect 8203 5386 8218 5398
rect 8200 5384 8222 5386
rect 8227 5384 8257 5398
rect 8318 5396 8471 5400
rect 8300 5384 8492 5396
rect 8535 5384 8565 5398
rect 8571 5384 8584 5414
rect 8599 5396 8629 5414
rect 8672 5384 8685 5414
rect 8715 5384 8728 5414
rect 8743 5396 8773 5414
rect 8816 5400 8830 5414
rect 8866 5400 9086 5414
rect 8817 5398 8830 5400
rect 8783 5386 8798 5398
rect 8780 5384 8802 5386
rect 8807 5384 8837 5398
rect 8898 5396 9051 5400
rect 8880 5384 9072 5396
rect 9115 5384 9145 5398
rect 9151 5384 9164 5414
rect 9179 5396 9209 5414
rect 9252 5384 9265 5414
rect 0 5370 9265 5384
rect 15 5266 28 5370
rect 73 5348 74 5358
rect 89 5348 102 5358
rect 73 5344 102 5348
rect 107 5344 137 5370
rect 155 5356 171 5358
rect 243 5356 296 5370
rect 244 5354 308 5356
rect 351 5354 366 5370
rect 415 5367 445 5370
rect 415 5364 451 5367
rect 381 5356 397 5358
rect 155 5344 170 5348
rect 73 5342 170 5344
rect 198 5342 366 5354
rect 382 5344 397 5348
rect 415 5345 454 5364
rect 473 5358 480 5359
rect 479 5351 480 5358
rect 463 5348 464 5351
rect 479 5348 492 5351
rect 415 5344 445 5345
rect 454 5344 460 5345
rect 463 5344 492 5348
rect 382 5343 492 5344
rect 382 5342 498 5343
rect 57 5334 108 5342
rect 57 5322 82 5334
rect 89 5322 108 5334
rect 139 5334 189 5342
rect 139 5326 155 5334
rect 162 5332 189 5334
rect 198 5332 419 5342
rect 162 5322 419 5332
rect 448 5334 498 5342
rect 448 5325 464 5334
rect 57 5314 108 5322
rect 155 5314 419 5322
rect 445 5322 464 5325
rect 471 5322 498 5334
rect 445 5314 498 5322
rect 73 5306 74 5314
rect 89 5306 102 5314
rect 73 5298 89 5306
rect 70 5291 89 5294
rect 70 5282 92 5291
rect 43 5272 92 5282
rect 43 5266 73 5272
rect 92 5267 97 5272
rect 15 5250 89 5266
rect 107 5258 137 5314
rect 172 5304 380 5314
rect 415 5310 460 5314
rect 463 5313 464 5314
rect 479 5313 492 5314
rect 198 5274 387 5304
rect 213 5271 387 5274
rect 206 5268 387 5271
rect 15 5248 28 5250
rect 43 5248 77 5250
rect 15 5232 89 5248
rect 116 5244 129 5258
rect 144 5244 160 5260
rect 206 5255 217 5268
rect -1 5210 0 5226
rect 15 5210 28 5232
rect 43 5210 73 5232
rect 116 5228 178 5244
rect 206 5237 217 5253
rect 222 5248 232 5268
rect 242 5248 256 5268
rect 259 5255 268 5268
rect 284 5255 293 5268
rect 222 5237 256 5248
rect 259 5237 268 5253
rect 284 5237 293 5253
rect 300 5248 310 5268
rect 320 5248 334 5268
rect 335 5255 346 5268
rect 300 5237 334 5248
rect 335 5237 346 5253
rect 392 5244 408 5260
rect 415 5258 445 5310
rect 479 5306 480 5313
rect 464 5298 480 5306
rect 451 5266 464 5285
rect 479 5266 509 5282
rect 451 5250 525 5266
rect 451 5248 464 5250
rect 479 5248 513 5250
rect 116 5226 129 5228
rect 144 5226 178 5228
rect 116 5210 178 5226
rect 222 5221 238 5224
rect 300 5221 330 5232
rect 378 5228 424 5244
rect 451 5232 525 5248
rect 378 5226 412 5228
rect 377 5210 424 5226
rect 451 5210 464 5232
rect 479 5210 509 5232
rect 536 5210 537 5226
rect 552 5210 565 5370
rect 595 5266 608 5370
rect 653 5348 654 5358
rect 669 5348 682 5358
rect 653 5344 682 5348
rect 687 5344 717 5370
rect 735 5356 751 5358
rect 823 5356 876 5370
rect 824 5354 888 5356
rect 931 5354 946 5370
rect 995 5367 1025 5370
rect 995 5364 1031 5367
rect 961 5356 977 5358
rect 735 5344 750 5348
rect 653 5342 750 5344
rect 778 5342 946 5354
rect 962 5344 977 5348
rect 995 5345 1034 5364
rect 1053 5358 1060 5359
rect 1059 5351 1060 5358
rect 1043 5348 1044 5351
rect 1059 5348 1072 5351
rect 995 5344 1025 5345
rect 1034 5344 1040 5345
rect 1043 5344 1072 5348
rect 962 5343 1072 5344
rect 962 5342 1078 5343
rect 637 5334 688 5342
rect 637 5322 662 5334
rect 669 5322 688 5334
rect 719 5334 769 5342
rect 719 5326 735 5334
rect 742 5332 769 5334
rect 778 5332 999 5342
rect 742 5322 999 5332
rect 1028 5334 1078 5342
rect 1028 5325 1044 5334
rect 637 5314 688 5322
rect 735 5314 999 5322
rect 1025 5322 1044 5325
rect 1051 5322 1078 5334
rect 1025 5314 1078 5322
rect 653 5306 654 5314
rect 669 5306 682 5314
rect 653 5298 669 5306
rect 650 5291 669 5294
rect 650 5282 672 5291
rect 623 5272 672 5282
rect 623 5266 653 5272
rect 672 5267 677 5272
rect 595 5250 669 5266
rect 687 5258 717 5314
rect 752 5304 960 5314
rect 995 5310 1040 5314
rect 1043 5313 1044 5314
rect 1059 5313 1072 5314
rect 778 5274 967 5304
rect 793 5271 967 5274
rect 786 5268 967 5271
rect 595 5248 608 5250
rect 623 5248 657 5250
rect 595 5232 669 5248
rect 696 5244 709 5258
rect 724 5244 740 5260
rect 786 5255 797 5268
rect 579 5210 580 5226
rect 595 5210 608 5232
rect 623 5210 653 5232
rect 696 5228 758 5244
rect 786 5237 797 5253
rect 802 5248 812 5268
rect 822 5248 836 5268
rect 839 5255 848 5268
rect 864 5255 873 5268
rect 802 5237 836 5248
rect 839 5237 848 5253
rect 864 5237 873 5253
rect 880 5248 890 5268
rect 900 5248 914 5268
rect 915 5255 926 5268
rect 880 5237 914 5248
rect 915 5237 926 5253
rect 972 5244 988 5260
rect 995 5258 1025 5310
rect 1059 5306 1060 5313
rect 1044 5298 1060 5306
rect 1031 5266 1044 5285
rect 1059 5266 1089 5282
rect 1031 5250 1105 5266
rect 1031 5248 1044 5250
rect 1059 5248 1093 5250
rect 696 5226 709 5228
rect 724 5226 758 5228
rect 696 5210 758 5226
rect 802 5221 818 5224
rect 880 5221 910 5232
rect 958 5228 1004 5244
rect 1031 5232 1105 5248
rect 958 5226 992 5228
rect 957 5210 1004 5226
rect 1031 5210 1044 5232
rect 1059 5210 1089 5232
rect 1116 5210 1117 5226
rect 1132 5210 1145 5370
rect 1175 5266 1188 5370
rect 1233 5348 1234 5358
rect 1249 5348 1262 5358
rect 1233 5344 1262 5348
rect 1267 5344 1297 5370
rect 1315 5356 1331 5358
rect 1403 5356 1456 5370
rect 1404 5354 1468 5356
rect 1511 5354 1526 5370
rect 1575 5367 1605 5370
rect 1575 5364 1611 5367
rect 1541 5356 1557 5358
rect 1315 5344 1330 5348
rect 1233 5342 1330 5344
rect 1358 5342 1526 5354
rect 1542 5344 1557 5348
rect 1575 5345 1614 5364
rect 1633 5358 1640 5359
rect 1639 5351 1640 5358
rect 1623 5348 1624 5351
rect 1639 5348 1652 5351
rect 1575 5344 1605 5345
rect 1614 5344 1620 5345
rect 1623 5344 1652 5348
rect 1542 5343 1652 5344
rect 1542 5342 1658 5343
rect 1217 5334 1268 5342
rect 1217 5322 1242 5334
rect 1249 5322 1268 5334
rect 1299 5334 1349 5342
rect 1299 5326 1315 5334
rect 1322 5332 1349 5334
rect 1358 5332 1579 5342
rect 1322 5322 1579 5332
rect 1608 5334 1658 5342
rect 1608 5325 1624 5334
rect 1217 5314 1268 5322
rect 1315 5314 1579 5322
rect 1605 5322 1624 5325
rect 1631 5322 1658 5334
rect 1605 5314 1658 5322
rect 1233 5306 1234 5314
rect 1249 5306 1262 5314
rect 1233 5298 1249 5306
rect 1230 5291 1249 5294
rect 1230 5282 1252 5291
rect 1203 5272 1252 5282
rect 1203 5266 1233 5272
rect 1252 5267 1257 5272
rect 1175 5250 1249 5266
rect 1267 5258 1297 5314
rect 1332 5304 1540 5314
rect 1575 5310 1620 5314
rect 1623 5313 1624 5314
rect 1639 5313 1652 5314
rect 1358 5274 1547 5304
rect 1373 5271 1547 5274
rect 1366 5268 1547 5271
rect 1175 5248 1188 5250
rect 1203 5248 1237 5250
rect 1175 5232 1249 5248
rect 1276 5244 1289 5258
rect 1304 5244 1320 5260
rect 1366 5255 1377 5268
rect 1159 5210 1160 5226
rect 1175 5210 1188 5232
rect 1203 5210 1233 5232
rect 1276 5228 1338 5244
rect 1366 5237 1377 5253
rect 1382 5248 1392 5268
rect 1402 5248 1416 5268
rect 1419 5255 1428 5268
rect 1444 5255 1453 5268
rect 1382 5237 1416 5248
rect 1419 5237 1428 5253
rect 1444 5237 1453 5253
rect 1460 5248 1470 5268
rect 1480 5248 1494 5268
rect 1495 5255 1506 5268
rect 1460 5237 1494 5248
rect 1495 5237 1506 5253
rect 1552 5244 1568 5260
rect 1575 5258 1605 5310
rect 1639 5306 1640 5313
rect 1624 5298 1640 5306
rect 1611 5266 1624 5285
rect 1639 5266 1669 5282
rect 1611 5250 1685 5266
rect 1611 5248 1624 5250
rect 1639 5248 1673 5250
rect 1276 5226 1289 5228
rect 1304 5226 1338 5228
rect 1276 5210 1338 5226
rect 1382 5221 1398 5224
rect 1460 5221 1490 5232
rect 1538 5228 1584 5244
rect 1611 5232 1685 5248
rect 1538 5226 1572 5228
rect 1537 5210 1584 5226
rect 1611 5210 1624 5232
rect 1639 5210 1669 5232
rect 1696 5210 1697 5226
rect 1712 5210 1725 5370
rect 1755 5266 1768 5370
rect 1813 5348 1814 5358
rect 1829 5348 1842 5358
rect 1813 5344 1842 5348
rect 1847 5344 1877 5370
rect 1895 5356 1911 5358
rect 1983 5356 2036 5370
rect 1984 5354 2048 5356
rect 2091 5354 2106 5370
rect 2155 5367 2185 5370
rect 2155 5364 2191 5367
rect 2121 5356 2137 5358
rect 1895 5344 1910 5348
rect 1813 5342 1910 5344
rect 1938 5342 2106 5354
rect 2122 5344 2137 5348
rect 2155 5345 2194 5364
rect 2213 5358 2220 5359
rect 2219 5351 2220 5358
rect 2203 5348 2204 5351
rect 2219 5348 2232 5351
rect 2155 5344 2185 5345
rect 2194 5344 2200 5345
rect 2203 5344 2232 5348
rect 2122 5343 2232 5344
rect 2122 5342 2238 5343
rect 1797 5334 1848 5342
rect 1797 5322 1822 5334
rect 1829 5322 1848 5334
rect 1879 5334 1929 5342
rect 1879 5326 1895 5334
rect 1902 5332 1929 5334
rect 1938 5332 2159 5342
rect 1902 5322 2159 5332
rect 2188 5334 2238 5342
rect 2188 5325 2204 5334
rect 1797 5314 1848 5322
rect 1895 5314 2159 5322
rect 2185 5322 2204 5325
rect 2211 5322 2238 5334
rect 2185 5314 2238 5322
rect 1813 5306 1814 5314
rect 1829 5306 1842 5314
rect 1813 5298 1829 5306
rect 1810 5291 1829 5294
rect 1810 5282 1832 5291
rect 1783 5272 1832 5282
rect 1783 5266 1813 5272
rect 1832 5267 1837 5272
rect 1755 5250 1829 5266
rect 1847 5258 1877 5314
rect 1912 5304 2120 5314
rect 2155 5310 2200 5314
rect 2203 5313 2204 5314
rect 2219 5313 2232 5314
rect 1938 5274 2127 5304
rect 1953 5271 2127 5274
rect 1946 5268 2127 5271
rect 1755 5248 1768 5250
rect 1783 5248 1817 5250
rect 1755 5232 1829 5248
rect 1856 5244 1869 5258
rect 1884 5244 1900 5260
rect 1946 5255 1957 5268
rect 1739 5210 1740 5226
rect 1755 5210 1768 5232
rect 1783 5210 1813 5232
rect 1856 5228 1918 5244
rect 1946 5237 1957 5253
rect 1962 5248 1972 5268
rect 1982 5248 1996 5268
rect 1999 5255 2008 5268
rect 2024 5255 2033 5268
rect 1962 5237 1996 5248
rect 1999 5237 2008 5253
rect 2024 5237 2033 5253
rect 2040 5248 2050 5268
rect 2060 5248 2074 5268
rect 2075 5255 2086 5268
rect 2040 5237 2074 5248
rect 2075 5237 2086 5253
rect 2132 5244 2148 5260
rect 2155 5258 2185 5310
rect 2219 5306 2220 5313
rect 2204 5298 2220 5306
rect 2191 5266 2204 5285
rect 2219 5266 2249 5282
rect 2191 5250 2265 5266
rect 2191 5248 2204 5250
rect 2219 5248 2253 5250
rect 1856 5226 1869 5228
rect 1884 5226 1918 5228
rect 1856 5210 1918 5226
rect 1962 5221 1976 5224
rect 2040 5221 2070 5232
rect 2118 5228 2164 5244
rect 2191 5232 2265 5248
rect 2118 5226 2152 5228
rect 2117 5210 2164 5226
rect 2191 5210 2204 5232
rect 2219 5210 2249 5232
rect 2276 5210 2277 5226
rect 2292 5210 2305 5370
rect 2335 5266 2348 5370
rect 2393 5348 2394 5358
rect 2409 5348 2422 5358
rect 2393 5344 2422 5348
rect 2427 5344 2457 5370
rect 2475 5356 2491 5358
rect 2563 5356 2616 5370
rect 2564 5354 2628 5356
rect 2671 5354 2686 5370
rect 2735 5367 2765 5370
rect 2735 5364 2771 5367
rect 2701 5356 2717 5358
rect 2475 5344 2490 5348
rect 2393 5342 2490 5344
rect 2518 5342 2686 5354
rect 2702 5344 2717 5348
rect 2735 5345 2774 5364
rect 2793 5358 2800 5359
rect 2799 5351 2800 5358
rect 2783 5348 2784 5351
rect 2799 5348 2812 5351
rect 2735 5344 2765 5345
rect 2774 5344 2780 5345
rect 2783 5344 2812 5348
rect 2702 5343 2812 5344
rect 2702 5342 2818 5343
rect 2377 5334 2428 5342
rect 2377 5322 2402 5334
rect 2409 5322 2428 5334
rect 2459 5334 2509 5342
rect 2459 5326 2475 5334
rect 2482 5332 2509 5334
rect 2518 5332 2739 5342
rect 2482 5322 2739 5332
rect 2768 5334 2818 5342
rect 2768 5325 2784 5334
rect 2377 5314 2428 5322
rect 2475 5314 2739 5322
rect 2765 5322 2784 5325
rect 2791 5322 2818 5334
rect 2765 5314 2818 5322
rect 2393 5306 2394 5314
rect 2409 5306 2422 5314
rect 2393 5298 2409 5306
rect 2390 5291 2409 5294
rect 2390 5282 2412 5291
rect 2363 5272 2412 5282
rect 2363 5266 2393 5272
rect 2412 5267 2417 5272
rect 2335 5250 2409 5266
rect 2427 5258 2457 5314
rect 2492 5304 2700 5314
rect 2735 5310 2780 5314
rect 2783 5313 2784 5314
rect 2799 5313 2812 5314
rect 2518 5274 2707 5304
rect 2533 5271 2707 5274
rect 2526 5268 2707 5271
rect 2335 5248 2348 5250
rect 2363 5248 2397 5250
rect 2335 5232 2409 5248
rect 2436 5244 2449 5258
rect 2464 5244 2480 5260
rect 2526 5255 2537 5268
rect 2319 5210 2320 5226
rect 2335 5210 2348 5232
rect 2363 5210 2393 5232
rect 2436 5228 2498 5244
rect 2526 5237 2537 5253
rect 2542 5248 2552 5268
rect 2562 5248 2576 5268
rect 2579 5255 2588 5268
rect 2604 5255 2613 5268
rect 2542 5237 2576 5248
rect 2579 5237 2588 5253
rect 2604 5237 2613 5253
rect 2620 5248 2630 5268
rect 2640 5248 2654 5268
rect 2655 5255 2666 5268
rect 2620 5237 2654 5248
rect 2655 5237 2666 5253
rect 2712 5244 2728 5260
rect 2735 5258 2765 5310
rect 2799 5306 2800 5313
rect 2784 5298 2800 5306
rect 2771 5266 2784 5285
rect 2799 5266 2829 5282
rect 2771 5250 2845 5266
rect 2771 5248 2784 5250
rect 2799 5248 2833 5250
rect 2436 5226 2449 5228
rect 2464 5226 2498 5228
rect 2436 5210 2498 5226
rect 2542 5221 2558 5224
rect 2620 5221 2650 5232
rect 2698 5228 2744 5244
rect 2771 5232 2845 5248
rect 2698 5226 2732 5228
rect 2697 5210 2744 5226
rect 2771 5210 2784 5232
rect 2799 5210 2829 5232
rect 2856 5210 2857 5226
rect 2872 5210 2885 5370
rect 2915 5266 2928 5370
rect 2973 5348 2974 5358
rect 2989 5348 3002 5358
rect 2973 5344 3002 5348
rect 3007 5344 3037 5370
rect 3055 5356 3071 5358
rect 3143 5356 3196 5370
rect 3144 5354 3208 5356
rect 3251 5354 3266 5370
rect 3315 5367 3345 5370
rect 3315 5364 3351 5367
rect 3281 5356 3297 5358
rect 3055 5344 3070 5348
rect 2973 5342 3070 5344
rect 3098 5342 3266 5354
rect 3282 5344 3297 5348
rect 3315 5345 3354 5364
rect 3373 5358 3380 5359
rect 3379 5351 3380 5358
rect 3363 5348 3364 5351
rect 3379 5348 3392 5351
rect 3315 5344 3345 5345
rect 3354 5344 3360 5345
rect 3363 5344 3392 5348
rect 3282 5343 3392 5344
rect 3282 5342 3398 5343
rect 2957 5334 3008 5342
rect 2957 5322 2982 5334
rect 2989 5322 3008 5334
rect 3039 5334 3089 5342
rect 3039 5326 3055 5334
rect 3062 5332 3089 5334
rect 3098 5332 3319 5342
rect 3062 5322 3319 5332
rect 3348 5334 3398 5342
rect 3348 5325 3364 5334
rect 2957 5314 3008 5322
rect 3055 5314 3319 5322
rect 3345 5322 3364 5325
rect 3371 5322 3398 5334
rect 3345 5314 3398 5322
rect 2973 5306 2974 5314
rect 2989 5306 3002 5314
rect 2973 5298 2989 5306
rect 2970 5291 2989 5294
rect 2970 5282 2992 5291
rect 2943 5272 2992 5282
rect 2943 5266 2973 5272
rect 2992 5267 2997 5272
rect 2915 5250 2989 5266
rect 3007 5258 3037 5314
rect 3072 5304 3280 5314
rect 3315 5310 3360 5314
rect 3363 5313 3364 5314
rect 3379 5313 3392 5314
rect 3098 5274 3287 5304
rect 3113 5271 3287 5274
rect 3106 5268 3287 5271
rect 2915 5248 2928 5250
rect 2943 5248 2977 5250
rect 2915 5232 2989 5248
rect 3016 5244 3029 5258
rect 3044 5244 3060 5260
rect 3106 5255 3117 5268
rect 2899 5210 2900 5226
rect 2915 5210 2928 5232
rect 2943 5210 2973 5232
rect 3016 5228 3078 5244
rect 3106 5237 3117 5253
rect 3122 5248 3132 5268
rect 3142 5248 3156 5268
rect 3159 5255 3168 5268
rect 3184 5255 3193 5268
rect 3122 5237 3156 5248
rect 3159 5237 3168 5253
rect 3184 5237 3193 5253
rect 3200 5248 3210 5268
rect 3220 5248 3234 5268
rect 3235 5255 3246 5268
rect 3200 5237 3234 5248
rect 3235 5237 3246 5253
rect 3292 5244 3308 5260
rect 3315 5258 3345 5310
rect 3379 5306 3380 5313
rect 3364 5298 3380 5306
rect 3351 5266 3364 5285
rect 3379 5266 3409 5282
rect 3351 5250 3425 5266
rect 3351 5248 3364 5250
rect 3379 5248 3413 5250
rect 3016 5226 3029 5228
rect 3044 5226 3078 5228
rect 3016 5210 3078 5226
rect 3122 5221 3138 5224
rect 3200 5221 3230 5232
rect 3278 5228 3324 5244
rect 3351 5232 3425 5248
rect 3278 5226 3312 5228
rect 3277 5210 3324 5226
rect 3351 5210 3364 5232
rect 3379 5210 3409 5232
rect 3436 5210 3437 5226
rect 3452 5210 3465 5370
rect 3495 5266 3508 5370
rect 3553 5348 3554 5358
rect 3569 5348 3582 5358
rect 3553 5344 3582 5348
rect 3587 5344 3617 5370
rect 3635 5356 3651 5358
rect 3723 5356 3776 5370
rect 3724 5354 3788 5356
rect 3831 5354 3846 5370
rect 3895 5367 3925 5370
rect 3895 5364 3931 5367
rect 3861 5356 3877 5358
rect 3635 5344 3650 5348
rect 3553 5342 3650 5344
rect 3678 5342 3846 5354
rect 3862 5344 3877 5348
rect 3895 5345 3934 5364
rect 3953 5358 3960 5359
rect 3959 5351 3960 5358
rect 3943 5348 3944 5351
rect 3959 5348 3972 5351
rect 3895 5344 3925 5345
rect 3934 5344 3940 5345
rect 3943 5344 3972 5348
rect 3862 5343 3972 5344
rect 3862 5342 3978 5343
rect 3537 5334 3588 5342
rect 3537 5322 3562 5334
rect 3569 5322 3588 5334
rect 3619 5334 3669 5342
rect 3619 5326 3635 5334
rect 3642 5332 3669 5334
rect 3678 5332 3899 5342
rect 3642 5322 3899 5332
rect 3928 5334 3978 5342
rect 3928 5325 3944 5334
rect 3537 5314 3588 5322
rect 3635 5314 3899 5322
rect 3925 5322 3944 5325
rect 3951 5322 3978 5334
rect 3925 5314 3978 5322
rect 3553 5306 3554 5314
rect 3569 5306 3582 5314
rect 3553 5298 3569 5306
rect 3550 5291 3569 5294
rect 3550 5282 3572 5291
rect 3523 5272 3572 5282
rect 3523 5266 3553 5272
rect 3572 5267 3577 5272
rect 3495 5250 3569 5266
rect 3587 5258 3617 5314
rect 3652 5304 3860 5314
rect 3895 5310 3940 5314
rect 3943 5313 3944 5314
rect 3959 5313 3972 5314
rect 3678 5274 3867 5304
rect 3693 5271 3867 5274
rect 3686 5268 3867 5271
rect 3495 5248 3508 5250
rect 3523 5248 3557 5250
rect 3495 5232 3569 5248
rect 3596 5244 3609 5258
rect 3624 5244 3640 5260
rect 3686 5255 3697 5268
rect 3479 5210 3480 5226
rect 3495 5210 3508 5232
rect 3523 5210 3553 5232
rect 3596 5228 3658 5244
rect 3686 5237 3697 5253
rect 3702 5248 3712 5268
rect 3722 5248 3736 5268
rect 3739 5255 3748 5268
rect 3764 5255 3773 5268
rect 3702 5237 3736 5248
rect 3739 5237 3748 5253
rect 3764 5237 3773 5253
rect 3780 5248 3790 5268
rect 3800 5248 3814 5268
rect 3815 5255 3826 5268
rect 3780 5237 3814 5248
rect 3815 5237 3826 5253
rect 3872 5244 3888 5260
rect 3895 5258 3925 5310
rect 3959 5306 3960 5313
rect 3944 5298 3960 5306
rect 3931 5266 3944 5285
rect 3959 5266 3989 5282
rect 3931 5250 4005 5266
rect 3931 5248 3944 5250
rect 3959 5248 3993 5250
rect 3596 5226 3609 5228
rect 3624 5226 3658 5228
rect 3596 5210 3658 5226
rect 3702 5221 3718 5224
rect 3780 5221 3810 5232
rect 3858 5228 3904 5244
rect 3931 5232 4005 5248
rect 3858 5226 3892 5228
rect 3857 5210 3904 5226
rect 3931 5210 3944 5232
rect 3959 5210 3989 5232
rect 4016 5210 4017 5226
rect 4032 5210 4045 5370
rect 4075 5266 4088 5370
rect 4133 5348 4134 5358
rect 4149 5348 4162 5358
rect 4133 5344 4162 5348
rect 4167 5344 4197 5370
rect 4215 5356 4231 5358
rect 4303 5356 4356 5370
rect 4304 5354 4368 5356
rect 4411 5354 4426 5370
rect 4475 5367 4505 5370
rect 4475 5364 4511 5367
rect 4441 5356 4457 5358
rect 4215 5344 4230 5348
rect 4133 5342 4230 5344
rect 4258 5342 4426 5354
rect 4442 5344 4457 5348
rect 4475 5345 4514 5364
rect 4533 5358 4540 5359
rect 4539 5351 4540 5358
rect 4523 5348 4524 5351
rect 4539 5348 4552 5351
rect 4475 5344 4505 5345
rect 4514 5344 4520 5345
rect 4523 5344 4552 5348
rect 4442 5343 4552 5344
rect 4442 5342 4558 5343
rect 4117 5334 4168 5342
rect 4117 5322 4142 5334
rect 4149 5322 4168 5334
rect 4199 5334 4249 5342
rect 4199 5326 4215 5334
rect 4222 5332 4249 5334
rect 4258 5332 4479 5342
rect 4222 5322 4479 5332
rect 4508 5334 4558 5342
rect 4508 5325 4524 5334
rect 4117 5314 4168 5322
rect 4215 5314 4479 5322
rect 4505 5322 4524 5325
rect 4531 5322 4558 5334
rect 4505 5314 4558 5322
rect 4133 5306 4134 5314
rect 4149 5306 4162 5314
rect 4133 5298 4149 5306
rect 4130 5291 4149 5294
rect 4130 5282 4152 5291
rect 4103 5272 4152 5282
rect 4103 5266 4133 5272
rect 4152 5267 4157 5272
rect 4075 5250 4149 5266
rect 4167 5258 4197 5314
rect 4232 5304 4440 5314
rect 4475 5310 4520 5314
rect 4523 5313 4524 5314
rect 4539 5313 4552 5314
rect 4258 5274 4447 5304
rect 4273 5271 4447 5274
rect 4266 5268 4447 5271
rect 4075 5248 4088 5250
rect 4103 5248 4137 5250
rect 4075 5232 4149 5248
rect 4176 5244 4189 5258
rect 4204 5244 4220 5260
rect 4266 5255 4277 5268
rect 4059 5210 4060 5226
rect 4075 5210 4088 5232
rect 4103 5210 4133 5232
rect 4176 5228 4238 5244
rect 4266 5237 4277 5253
rect 4282 5248 4292 5268
rect 4302 5248 4316 5268
rect 4319 5255 4328 5268
rect 4344 5255 4353 5268
rect 4282 5237 4316 5248
rect 4319 5237 4328 5253
rect 4344 5237 4353 5253
rect 4360 5248 4370 5268
rect 4380 5248 4394 5268
rect 4395 5255 4406 5268
rect 4360 5237 4394 5248
rect 4395 5237 4406 5253
rect 4452 5244 4468 5260
rect 4475 5258 4505 5310
rect 4539 5306 4540 5313
rect 4524 5298 4540 5306
rect 4511 5266 4524 5285
rect 4539 5266 4569 5282
rect 4511 5250 4585 5266
rect 4511 5248 4524 5250
rect 4539 5248 4573 5250
rect 4176 5226 4189 5228
rect 4204 5226 4238 5228
rect 4176 5210 4238 5226
rect 4282 5221 4298 5224
rect 4360 5221 4390 5232
rect 4438 5228 4484 5244
rect 4511 5232 4585 5248
rect 4438 5226 4472 5228
rect 4437 5210 4484 5226
rect 4511 5210 4524 5232
rect 4539 5210 4569 5232
rect 4596 5210 4597 5226
rect 4612 5210 4625 5370
rect 4655 5266 4668 5370
rect 4713 5348 4714 5358
rect 4729 5348 4742 5358
rect 4713 5344 4742 5348
rect 4747 5344 4777 5370
rect 4795 5356 4811 5358
rect 4883 5356 4936 5370
rect 4884 5354 4948 5356
rect 4991 5354 5006 5370
rect 5055 5367 5085 5370
rect 5055 5364 5091 5367
rect 5021 5356 5037 5358
rect 4795 5344 4810 5348
rect 4713 5342 4810 5344
rect 4838 5342 5006 5354
rect 5022 5344 5037 5348
rect 5055 5345 5094 5364
rect 5113 5358 5120 5359
rect 5119 5351 5120 5358
rect 5103 5348 5104 5351
rect 5119 5348 5132 5351
rect 5055 5344 5085 5345
rect 5094 5344 5100 5345
rect 5103 5344 5132 5348
rect 5022 5343 5132 5344
rect 5022 5342 5138 5343
rect 4697 5334 4748 5342
rect 4697 5322 4722 5334
rect 4729 5322 4748 5334
rect 4779 5334 4829 5342
rect 4779 5326 4795 5334
rect 4802 5332 4829 5334
rect 4838 5332 5059 5342
rect 4802 5322 5059 5332
rect 5088 5334 5138 5342
rect 5088 5325 5104 5334
rect 4697 5314 4748 5322
rect 4795 5314 5059 5322
rect 5085 5322 5104 5325
rect 5111 5322 5138 5334
rect 5085 5314 5138 5322
rect 4713 5306 4714 5314
rect 4729 5306 4742 5314
rect 4713 5298 4729 5306
rect 4710 5291 4729 5294
rect 4710 5282 4732 5291
rect 4683 5272 4732 5282
rect 4683 5266 4713 5272
rect 4732 5267 4737 5272
rect 4655 5250 4729 5266
rect 4747 5258 4777 5314
rect 4812 5304 5020 5314
rect 5055 5310 5100 5314
rect 5103 5313 5104 5314
rect 5119 5313 5132 5314
rect 4838 5274 5027 5304
rect 4853 5271 5027 5274
rect 4846 5268 5027 5271
rect 4655 5248 4668 5250
rect 4683 5248 4717 5250
rect 4655 5232 4729 5248
rect 4756 5244 4769 5258
rect 4784 5244 4800 5260
rect 4846 5255 4857 5268
rect 4639 5210 4640 5226
rect 4655 5210 4668 5232
rect 4683 5210 4713 5232
rect 4756 5228 4818 5244
rect 4846 5237 4857 5253
rect 4862 5248 4872 5268
rect 4882 5248 4896 5268
rect 4899 5255 4908 5268
rect 4924 5255 4933 5268
rect 4862 5237 4896 5248
rect 4899 5237 4908 5253
rect 4924 5237 4933 5253
rect 4940 5248 4950 5268
rect 4960 5248 4974 5268
rect 4975 5255 4986 5268
rect 4940 5237 4974 5248
rect 4975 5237 4986 5253
rect 5032 5244 5048 5260
rect 5055 5258 5085 5310
rect 5119 5306 5120 5313
rect 5104 5298 5120 5306
rect 5091 5266 5104 5285
rect 5119 5266 5149 5282
rect 5091 5250 5165 5266
rect 5091 5248 5104 5250
rect 5119 5248 5153 5250
rect 4756 5226 4769 5228
rect 4784 5226 4818 5228
rect 4756 5210 4818 5226
rect 4862 5221 4878 5224
rect 4940 5221 4970 5232
rect 5018 5228 5064 5244
rect 5091 5232 5165 5248
rect 5018 5226 5052 5228
rect 5017 5210 5064 5226
rect 5091 5210 5104 5232
rect 5119 5210 5149 5232
rect 5176 5210 5177 5226
rect 5192 5210 5205 5370
rect 5235 5266 5248 5370
rect 5293 5348 5294 5358
rect 5309 5348 5322 5358
rect 5293 5344 5322 5348
rect 5327 5344 5357 5370
rect 5375 5356 5391 5358
rect 5463 5356 5516 5370
rect 5464 5354 5528 5356
rect 5571 5354 5586 5370
rect 5635 5367 5665 5370
rect 5635 5364 5671 5367
rect 5601 5356 5617 5358
rect 5375 5344 5390 5348
rect 5293 5342 5390 5344
rect 5418 5342 5586 5354
rect 5602 5344 5617 5348
rect 5635 5345 5674 5364
rect 5693 5358 5700 5359
rect 5699 5351 5700 5358
rect 5683 5348 5684 5351
rect 5699 5348 5712 5351
rect 5635 5344 5665 5345
rect 5674 5344 5680 5345
rect 5683 5344 5712 5348
rect 5602 5343 5712 5344
rect 5602 5342 5718 5343
rect 5277 5334 5328 5342
rect 5277 5322 5302 5334
rect 5309 5322 5328 5334
rect 5359 5334 5409 5342
rect 5359 5326 5375 5334
rect 5382 5332 5409 5334
rect 5418 5332 5639 5342
rect 5382 5322 5639 5332
rect 5668 5334 5718 5342
rect 5668 5325 5684 5334
rect 5277 5314 5328 5322
rect 5375 5314 5639 5322
rect 5665 5322 5684 5325
rect 5691 5322 5718 5334
rect 5665 5314 5718 5322
rect 5293 5306 5294 5314
rect 5309 5306 5322 5314
rect 5293 5298 5309 5306
rect 5290 5291 5309 5294
rect 5290 5282 5312 5291
rect 5263 5272 5312 5282
rect 5263 5266 5293 5272
rect 5312 5267 5317 5272
rect 5235 5250 5309 5266
rect 5327 5258 5357 5314
rect 5392 5304 5600 5314
rect 5635 5310 5680 5314
rect 5683 5313 5684 5314
rect 5699 5313 5712 5314
rect 5418 5274 5607 5304
rect 5433 5271 5607 5274
rect 5426 5268 5607 5271
rect 5235 5248 5248 5250
rect 5263 5248 5297 5250
rect 5235 5232 5309 5248
rect 5336 5244 5349 5258
rect 5364 5244 5380 5260
rect 5426 5255 5437 5268
rect 5219 5210 5220 5226
rect 5235 5210 5248 5232
rect 5263 5210 5293 5232
rect 5336 5228 5398 5244
rect 5426 5237 5437 5253
rect 5442 5248 5452 5268
rect 5462 5248 5476 5268
rect 5479 5255 5488 5268
rect 5504 5255 5513 5268
rect 5442 5237 5476 5248
rect 5479 5237 5488 5253
rect 5504 5237 5513 5253
rect 5520 5248 5530 5268
rect 5540 5248 5554 5268
rect 5555 5255 5566 5268
rect 5520 5237 5554 5248
rect 5555 5237 5566 5253
rect 5612 5244 5628 5260
rect 5635 5258 5665 5310
rect 5699 5306 5700 5313
rect 5684 5298 5700 5306
rect 5671 5266 5684 5285
rect 5699 5266 5729 5282
rect 5671 5250 5745 5266
rect 5671 5248 5684 5250
rect 5699 5248 5733 5250
rect 5336 5226 5349 5228
rect 5364 5226 5398 5228
rect 5336 5210 5398 5226
rect 5442 5221 5458 5224
rect 5520 5221 5550 5232
rect 5598 5228 5644 5244
rect 5671 5232 5745 5248
rect 5598 5226 5632 5228
rect 5597 5210 5644 5226
rect 5671 5210 5684 5232
rect 5699 5210 5729 5232
rect 5756 5210 5757 5226
rect 5772 5210 5785 5370
rect 5815 5266 5828 5370
rect 5873 5348 5874 5358
rect 5889 5348 5902 5358
rect 5873 5344 5902 5348
rect 5907 5344 5937 5370
rect 5955 5356 5971 5358
rect 6043 5356 6096 5370
rect 6044 5354 6108 5356
rect 6151 5354 6166 5370
rect 6215 5367 6245 5370
rect 6215 5364 6251 5367
rect 6181 5356 6197 5358
rect 5955 5344 5970 5348
rect 5873 5342 5970 5344
rect 5998 5342 6166 5354
rect 6182 5344 6197 5348
rect 6215 5345 6254 5364
rect 6273 5358 6280 5359
rect 6279 5351 6280 5358
rect 6263 5348 6264 5351
rect 6279 5348 6292 5351
rect 6215 5344 6245 5345
rect 6254 5344 6260 5345
rect 6263 5344 6292 5348
rect 6182 5343 6292 5344
rect 6182 5342 6298 5343
rect 5857 5334 5908 5342
rect 5857 5322 5882 5334
rect 5889 5322 5908 5334
rect 5939 5334 5989 5342
rect 5939 5326 5955 5334
rect 5962 5332 5989 5334
rect 5998 5332 6219 5342
rect 5962 5322 6219 5332
rect 6248 5334 6298 5342
rect 6248 5325 6264 5334
rect 5857 5314 5908 5322
rect 5955 5314 6219 5322
rect 6245 5322 6264 5325
rect 6271 5322 6298 5334
rect 6245 5314 6298 5322
rect 5873 5306 5874 5314
rect 5889 5306 5902 5314
rect 5873 5298 5889 5306
rect 5870 5291 5889 5294
rect 5870 5282 5892 5291
rect 5843 5272 5892 5282
rect 5843 5266 5873 5272
rect 5892 5267 5897 5272
rect 5815 5250 5889 5266
rect 5907 5258 5937 5314
rect 5972 5304 6180 5314
rect 6215 5310 6260 5314
rect 6263 5313 6264 5314
rect 6279 5313 6292 5314
rect 5998 5274 6187 5304
rect 6013 5271 6187 5274
rect 6006 5268 6187 5271
rect 5815 5248 5828 5250
rect 5843 5248 5877 5250
rect 5815 5232 5889 5248
rect 5916 5244 5929 5258
rect 5944 5244 5960 5260
rect 6006 5255 6017 5268
rect 5799 5210 5800 5226
rect 5815 5210 5828 5232
rect 5843 5210 5873 5232
rect 5916 5228 5978 5244
rect 6006 5237 6017 5253
rect 6022 5248 6032 5268
rect 6042 5248 6056 5268
rect 6059 5255 6068 5268
rect 6084 5255 6093 5268
rect 6022 5237 6056 5248
rect 6059 5237 6068 5253
rect 6084 5237 6093 5253
rect 6100 5248 6110 5268
rect 6120 5248 6134 5268
rect 6135 5255 6146 5268
rect 6100 5237 6134 5248
rect 6135 5237 6146 5253
rect 6192 5244 6208 5260
rect 6215 5258 6245 5310
rect 6279 5306 6280 5313
rect 6264 5298 6280 5306
rect 6251 5266 6264 5285
rect 6279 5266 6309 5282
rect 6251 5250 6325 5266
rect 6251 5248 6264 5250
rect 6279 5248 6313 5250
rect 5916 5226 5929 5228
rect 5944 5226 5978 5228
rect 5916 5210 5978 5226
rect 6022 5221 6038 5224
rect 6100 5221 6130 5232
rect 6178 5228 6224 5244
rect 6251 5232 6325 5248
rect 6178 5226 6212 5228
rect 6177 5210 6224 5226
rect 6251 5210 6264 5232
rect 6279 5210 6309 5232
rect 6336 5210 6337 5226
rect 6352 5210 6365 5370
rect 6395 5266 6408 5370
rect 6453 5348 6454 5358
rect 6469 5348 6482 5358
rect 6453 5344 6482 5348
rect 6487 5344 6517 5370
rect 6535 5356 6551 5358
rect 6623 5356 6676 5370
rect 6624 5354 6688 5356
rect 6731 5354 6746 5370
rect 6795 5367 6825 5370
rect 6795 5364 6831 5367
rect 6761 5356 6777 5358
rect 6535 5344 6550 5348
rect 6453 5342 6550 5344
rect 6578 5342 6746 5354
rect 6762 5344 6777 5348
rect 6795 5345 6834 5364
rect 6853 5358 6860 5359
rect 6859 5351 6860 5358
rect 6843 5348 6844 5351
rect 6859 5348 6872 5351
rect 6795 5344 6825 5345
rect 6834 5344 6840 5345
rect 6843 5344 6872 5348
rect 6762 5343 6872 5344
rect 6762 5342 6878 5343
rect 6437 5334 6488 5342
rect 6437 5322 6462 5334
rect 6469 5322 6488 5334
rect 6519 5334 6569 5342
rect 6519 5326 6535 5334
rect 6542 5332 6569 5334
rect 6578 5332 6799 5342
rect 6542 5322 6799 5332
rect 6828 5334 6878 5342
rect 6828 5325 6844 5334
rect 6437 5314 6488 5322
rect 6535 5314 6799 5322
rect 6825 5322 6844 5325
rect 6851 5322 6878 5334
rect 6825 5314 6878 5322
rect 6453 5306 6454 5314
rect 6469 5306 6482 5314
rect 6453 5298 6469 5306
rect 6450 5291 6469 5294
rect 6450 5282 6472 5291
rect 6423 5272 6472 5282
rect 6423 5266 6453 5272
rect 6472 5267 6477 5272
rect 6395 5250 6469 5266
rect 6487 5258 6517 5314
rect 6552 5304 6760 5314
rect 6795 5310 6840 5314
rect 6843 5313 6844 5314
rect 6859 5313 6872 5314
rect 6578 5274 6767 5304
rect 6593 5271 6767 5274
rect 6586 5268 6767 5271
rect 6395 5248 6408 5250
rect 6423 5248 6457 5250
rect 6395 5232 6469 5248
rect 6496 5244 6509 5258
rect 6524 5244 6540 5260
rect 6586 5255 6597 5268
rect 6379 5210 6380 5226
rect 6395 5210 6408 5232
rect 6423 5210 6453 5232
rect 6496 5228 6558 5244
rect 6586 5237 6597 5253
rect 6602 5248 6612 5268
rect 6622 5248 6636 5268
rect 6639 5255 6648 5268
rect 6664 5255 6673 5268
rect 6602 5237 6636 5248
rect 6639 5237 6648 5253
rect 6664 5237 6673 5253
rect 6680 5248 6690 5268
rect 6700 5248 6714 5268
rect 6715 5255 6726 5268
rect 6680 5237 6714 5248
rect 6715 5237 6726 5253
rect 6772 5244 6788 5260
rect 6795 5258 6825 5310
rect 6859 5306 6860 5313
rect 6844 5298 6860 5306
rect 6831 5266 6844 5285
rect 6859 5266 6889 5282
rect 6831 5250 6905 5266
rect 6831 5248 6844 5250
rect 6859 5248 6893 5250
rect 6496 5226 6509 5228
rect 6524 5226 6558 5228
rect 6496 5210 6558 5226
rect 6602 5221 6618 5224
rect 6680 5221 6710 5232
rect 6758 5228 6804 5244
rect 6831 5232 6905 5248
rect 6758 5226 6792 5228
rect 6757 5210 6804 5226
rect 6831 5210 6844 5232
rect 6859 5210 6889 5232
rect 6916 5210 6917 5226
rect 6932 5210 6945 5370
rect 6975 5266 6988 5370
rect 7033 5348 7034 5358
rect 7049 5348 7062 5358
rect 7033 5344 7062 5348
rect 7067 5344 7097 5370
rect 7115 5356 7131 5358
rect 7203 5356 7256 5370
rect 7204 5354 7268 5356
rect 7311 5354 7326 5370
rect 7375 5367 7405 5370
rect 7375 5364 7411 5367
rect 7341 5356 7357 5358
rect 7115 5344 7130 5348
rect 7033 5342 7130 5344
rect 7158 5342 7326 5354
rect 7342 5344 7357 5348
rect 7375 5345 7414 5364
rect 7433 5358 7440 5359
rect 7439 5351 7440 5358
rect 7423 5348 7424 5351
rect 7439 5348 7452 5351
rect 7375 5344 7405 5345
rect 7414 5344 7420 5345
rect 7423 5344 7452 5348
rect 7342 5343 7452 5344
rect 7342 5342 7458 5343
rect 7017 5334 7068 5342
rect 7017 5322 7042 5334
rect 7049 5322 7068 5334
rect 7099 5334 7149 5342
rect 7099 5326 7115 5334
rect 7122 5332 7149 5334
rect 7158 5332 7379 5342
rect 7122 5322 7379 5332
rect 7408 5334 7458 5342
rect 7408 5325 7424 5334
rect 7017 5314 7068 5322
rect 7115 5314 7379 5322
rect 7405 5322 7424 5325
rect 7431 5322 7458 5334
rect 7405 5314 7458 5322
rect 7033 5306 7034 5314
rect 7049 5306 7062 5314
rect 7033 5298 7049 5306
rect 7030 5291 7049 5294
rect 7030 5282 7052 5291
rect 7003 5272 7052 5282
rect 7003 5266 7033 5272
rect 7052 5267 7057 5272
rect 6975 5250 7049 5266
rect 7067 5258 7097 5314
rect 7132 5304 7340 5314
rect 7375 5310 7420 5314
rect 7423 5313 7424 5314
rect 7439 5313 7452 5314
rect 7158 5274 7347 5304
rect 7173 5271 7347 5274
rect 7166 5268 7347 5271
rect 6975 5248 6988 5250
rect 7003 5248 7037 5250
rect 6975 5232 7049 5248
rect 7076 5244 7089 5258
rect 7104 5244 7120 5260
rect 7166 5255 7177 5268
rect 6959 5210 6960 5226
rect 6975 5210 6988 5232
rect 7003 5210 7033 5232
rect 7076 5228 7138 5244
rect 7166 5237 7177 5253
rect 7182 5248 7192 5268
rect 7202 5248 7216 5268
rect 7219 5255 7228 5268
rect 7244 5255 7253 5268
rect 7182 5237 7216 5248
rect 7219 5237 7228 5253
rect 7244 5237 7253 5253
rect 7260 5248 7270 5268
rect 7280 5248 7294 5268
rect 7295 5255 7306 5268
rect 7260 5237 7294 5248
rect 7295 5237 7306 5253
rect 7352 5244 7368 5260
rect 7375 5258 7405 5310
rect 7439 5306 7440 5313
rect 7424 5298 7440 5306
rect 7411 5266 7424 5285
rect 7439 5266 7469 5282
rect 7411 5250 7485 5266
rect 7411 5248 7424 5250
rect 7439 5248 7473 5250
rect 7076 5226 7089 5228
rect 7104 5226 7138 5228
rect 7076 5210 7138 5226
rect 7182 5221 7198 5224
rect 7260 5221 7290 5232
rect 7338 5228 7384 5244
rect 7411 5232 7485 5248
rect 7338 5226 7372 5228
rect 7337 5210 7384 5226
rect 7411 5210 7424 5232
rect 7439 5210 7469 5232
rect 7496 5210 7497 5226
rect 7512 5210 7525 5370
rect 7555 5266 7568 5370
rect 7613 5348 7614 5358
rect 7629 5348 7642 5358
rect 7613 5344 7642 5348
rect 7647 5344 7677 5370
rect 7695 5356 7711 5358
rect 7783 5356 7836 5370
rect 7784 5354 7848 5356
rect 7891 5354 7906 5370
rect 7955 5367 7985 5370
rect 7955 5364 7991 5367
rect 7921 5356 7937 5358
rect 7695 5344 7710 5348
rect 7613 5342 7710 5344
rect 7738 5342 7906 5354
rect 7922 5344 7937 5348
rect 7955 5345 7994 5364
rect 8013 5358 8020 5359
rect 8019 5351 8020 5358
rect 8003 5348 8004 5351
rect 8019 5348 8032 5351
rect 7955 5344 7985 5345
rect 7994 5344 8000 5345
rect 8003 5344 8032 5348
rect 7922 5343 8032 5344
rect 7922 5342 8038 5343
rect 7597 5334 7648 5342
rect 7597 5322 7622 5334
rect 7629 5322 7648 5334
rect 7679 5334 7729 5342
rect 7679 5326 7695 5334
rect 7702 5332 7729 5334
rect 7738 5332 7959 5342
rect 7702 5322 7959 5332
rect 7988 5334 8038 5342
rect 7988 5325 8004 5334
rect 7597 5314 7648 5322
rect 7695 5314 7959 5322
rect 7985 5322 8004 5325
rect 8011 5322 8038 5334
rect 7985 5314 8038 5322
rect 7613 5306 7614 5314
rect 7629 5306 7642 5314
rect 7613 5298 7629 5306
rect 7610 5291 7629 5294
rect 7610 5282 7632 5291
rect 7583 5272 7632 5282
rect 7583 5266 7613 5272
rect 7632 5267 7637 5272
rect 7555 5250 7629 5266
rect 7647 5258 7677 5314
rect 7712 5304 7920 5314
rect 7955 5310 8000 5314
rect 8003 5313 8004 5314
rect 8019 5313 8032 5314
rect 7738 5274 7927 5304
rect 7753 5271 7927 5274
rect 7746 5268 7927 5271
rect 7555 5248 7568 5250
rect 7583 5248 7617 5250
rect 7555 5232 7629 5248
rect 7656 5244 7669 5258
rect 7684 5244 7700 5260
rect 7746 5255 7757 5268
rect 7539 5210 7540 5226
rect 7555 5210 7568 5232
rect 7583 5210 7613 5232
rect 7656 5228 7718 5244
rect 7746 5237 7757 5253
rect 7762 5248 7772 5268
rect 7782 5248 7796 5268
rect 7799 5255 7808 5268
rect 7824 5255 7833 5268
rect 7762 5237 7796 5248
rect 7799 5237 7808 5253
rect 7824 5237 7833 5253
rect 7840 5248 7850 5268
rect 7860 5248 7874 5268
rect 7875 5255 7886 5268
rect 7840 5237 7874 5248
rect 7875 5237 7886 5253
rect 7932 5244 7948 5260
rect 7955 5258 7985 5310
rect 8019 5306 8020 5313
rect 8004 5298 8020 5306
rect 7991 5266 8004 5285
rect 8019 5266 8049 5282
rect 7991 5250 8065 5266
rect 7991 5248 8004 5250
rect 8019 5248 8053 5250
rect 7656 5226 7669 5228
rect 7684 5226 7718 5228
rect 7656 5210 7718 5226
rect 7762 5221 7778 5224
rect 7840 5221 7870 5232
rect 7918 5228 7964 5244
rect 7991 5232 8065 5248
rect 7918 5226 7952 5228
rect 7917 5210 7964 5226
rect 7991 5210 8004 5232
rect 8019 5210 8049 5232
rect 8076 5210 8077 5226
rect 8092 5210 8105 5370
rect 8135 5266 8148 5370
rect 8193 5348 8194 5358
rect 8209 5348 8222 5358
rect 8193 5344 8222 5348
rect 8227 5344 8257 5370
rect 8275 5356 8291 5358
rect 8363 5356 8416 5370
rect 8364 5354 8428 5356
rect 8471 5354 8486 5370
rect 8535 5367 8565 5370
rect 8535 5364 8571 5367
rect 8501 5356 8517 5358
rect 8275 5344 8290 5348
rect 8193 5342 8290 5344
rect 8318 5342 8486 5354
rect 8502 5344 8517 5348
rect 8535 5345 8574 5364
rect 8593 5358 8600 5359
rect 8599 5351 8600 5358
rect 8583 5348 8584 5351
rect 8599 5348 8612 5351
rect 8535 5344 8565 5345
rect 8574 5344 8580 5345
rect 8583 5344 8612 5348
rect 8502 5343 8612 5344
rect 8502 5342 8618 5343
rect 8177 5334 8228 5342
rect 8177 5322 8202 5334
rect 8209 5322 8228 5334
rect 8259 5334 8309 5342
rect 8259 5326 8275 5334
rect 8282 5332 8309 5334
rect 8318 5332 8539 5342
rect 8282 5322 8539 5332
rect 8568 5334 8618 5342
rect 8568 5325 8584 5334
rect 8177 5314 8228 5322
rect 8275 5314 8539 5322
rect 8565 5322 8584 5325
rect 8591 5322 8618 5334
rect 8565 5314 8618 5322
rect 8193 5306 8194 5314
rect 8209 5306 8222 5314
rect 8193 5298 8209 5306
rect 8190 5291 8209 5294
rect 8190 5282 8212 5291
rect 8163 5272 8212 5282
rect 8163 5266 8193 5272
rect 8212 5267 8217 5272
rect 8135 5250 8209 5266
rect 8227 5258 8257 5314
rect 8292 5304 8500 5314
rect 8535 5310 8580 5314
rect 8583 5313 8584 5314
rect 8599 5313 8612 5314
rect 8318 5274 8507 5304
rect 8333 5271 8507 5274
rect 8326 5268 8507 5271
rect 8135 5248 8148 5250
rect 8163 5248 8197 5250
rect 8135 5232 8209 5248
rect 8236 5244 8249 5258
rect 8264 5244 8280 5260
rect 8326 5255 8337 5268
rect 8119 5210 8120 5226
rect 8135 5210 8148 5232
rect 8163 5210 8193 5232
rect 8236 5228 8298 5244
rect 8326 5237 8337 5253
rect 8342 5248 8352 5268
rect 8362 5248 8376 5268
rect 8379 5255 8388 5268
rect 8404 5255 8413 5268
rect 8342 5237 8376 5248
rect 8379 5237 8388 5253
rect 8404 5237 8413 5253
rect 8420 5248 8430 5268
rect 8440 5248 8454 5268
rect 8455 5255 8466 5268
rect 8420 5237 8454 5248
rect 8455 5237 8466 5253
rect 8512 5244 8528 5260
rect 8535 5258 8565 5310
rect 8599 5306 8600 5313
rect 8584 5298 8600 5306
rect 8571 5266 8584 5285
rect 8599 5266 8629 5282
rect 8571 5250 8645 5266
rect 8571 5248 8584 5250
rect 8599 5248 8633 5250
rect 8236 5226 8249 5228
rect 8264 5226 8298 5228
rect 8236 5210 8298 5226
rect 8342 5221 8358 5224
rect 8420 5221 8450 5232
rect 8498 5228 8544 5244
rect 8571 5232 8645 5248
rect 8498 5226 8532 5228
rect 8497 5210 8544 5226
rect 8571 5210 8584 5232
rect 8599 5210 8629 5232
rect 8656 5210 8657 5226
rect 8672 5210 8685 5370
rect 8715 5266 8728 5370
rect 8773 5348 8774 5358
rect 8789 5348 8802 5358
rect 8773 5344 8802 5348
rect 8807 5344 8837 5370
rect 8855 5356 8871 5358
rect 8943 5356 8996 5370
rect 8944 5354 9008 5356
rect 9051 5354 9066 5370
rect 9115 5367 9145 5370
rect 9115 5364 9151 5367
rect 9081 5356 9097 5358
rect 8855 5344 8870 5348
rect 8773 5342 8870 5344
rect 8898 5342 9066 5354
rect 9082 5344 9097 5348
rect 9115 5345 9154 5364
rect 9173 5358 9180 5359
rect 9179 5351 9180 5358
rect 9163 5348 9164 5351
rect 9179 5348 9192 5351
rect 9115 5344 9145 5345
rect 9154 5344 9160 5345
rect 9163 5344 9192 5348
rect 9082 5343 9192 5344
rect 9082 5342 9198 5343
rect 8757 5334 8808 5342
rect 8757 5322 8782 5334
rect 8789 5322 8808 5334
rect 8839 5334 8889 5342
rect 8839 5326 8855 5334
rect 8862 5332 8889 5334
rect 8898 5332 9119 5342
rect 8862 5322 9119 5332
rect 9148 5334 9198 5342
rect 9148 5325 9164 5334
rect 8757 5314 8808 5322
rect 8855 5314 9119 5322
rect 9145 5322 9164 5325
rect 9171 5322 9198 5334
rect 9145 5314 9198 5322
rect 8773 5306 8774 5314
rect 8789 5306 8802 5314
rect 8773 5298 8789 5306
rect 8770 5291 8789 5294
rect 8770 5282 8792 5291
rect 8743 5272 8792 5282
rect 8743 5266 8773 5272
rect 8792 5267 8797 5272
rect 8715 5250 8789 5266
rect 8807 5258 8837 5314
rect 8872 5304 9080 5314
rect 9115 5310 9160 5314
rect 9163 5313 9164 5314
rect 9179 5313 9192 5314
rect 8898 5274 9087 5304
rect 8913 5271 9087 5274
rect 8906 5268 9087 5271
rect 8715 5248 8728 5250
rect 8743 5248 8777 5250
rect 8715 5232 8789 5248
rect 8816 5244 8829 5258
rect 8844 5244 8860 5260
rect 8906 5255 8917 5268
rect 8699 5210 8700 5226
rect 8715 5210 8728 5232
rect 8743 5210 8773 5232
rect 8816 5228 8878 5244
rect 8906 5237 8917 5253
rect 8922 5248 8932 5268
rect 8942 5248 8956 5268
rect 8959 5255 8968 5268
rect 8984 5255 8993 5268
rect 8922 5237 8956 5248
rect 8959 5237 8968 5253
rect 8984 5237 8993 5253
rect 9000 5248 9010 5268
rect 9020 5248 9034 5268
rect 9035 5255 9046 5268
rect 9000 5237 9034 5248
rect 9035 5237 9046 5253
rect 9092 5244 9108 5260
rect 9115 5258 9145 5310
rect 9179 5306 9180 5313
rect 9164 5298 9180 5306
rect 9151 5266 9164 5285
rect 9179 5266 9209 5282
rect 9151 5250 9225 5266
rect 9151 5248 9164 5250
rect 9179 5248 9213 5250
rect 8816 5226 8829 5228
rect 8844 5226 8878 5228
rect 8816 5210 8878 5226
rect 8922 5221 8938 5224
rect 9000 5221 9030 5232
rect 9078 5228 9124 5244
rect 9151 5232 9225 5248
rect 9078 5226 9112 5228
rect 9077 5210 9124 5226
rect 9151 5210 9164 5232
rect 9179 5210 9209 5232
rect 9236 5210 9237 5226
rect 9252 5210 9265 5370
rect -7 5202 34 5210
rect -7 5176 8 5202
rect 15 5176 34 5202
rect 98 5198 160 5210
rect 172 5198 247 5210
rect 305 5198 380 5210
rect 392 5198 423 5210
rect 429 5198 464 5210
rect 98 5196 260 5198
rect -7 5168 34 5176
rect 116 5172 129 5196
rect 144 5194 159 5196
rect -1 5158 0 5168
rect 15 5158 28 5168
rect 43 5158 73 5172
rect 116 5158 159 5172
rect 183 5169 190 5176
rect 193 5172 260 5196
rect 292 5196 464 5198
rect 262 5174 290 5178
rect 292 5174 372 5196
rect 393 5194 408 5196
rect 262 5172 372 5174
rect 193 5168 372 5172
rect 166 5158 196 5168
rect 198 5158 351 5168
rect 359 5158 389 5168
rect 393 5158 423 5172
rect 451 5158 464 5196
rect 536 5202 571 5210
rect 536 5176 537 5202
rect 544 5176 571 5202
rect 479 5158 509 5172
rect 536 5168 571 5176
rect 573 5202 614 5210
rect 573 5176 588 5202
rect 595 5176 614 5202
rect 678 5198 740 5210
rect 752 5198 827 5210
rect 885 5198 960 5210
rect 972 5198 1003 5210
rect 1009 5198 1044 5210
rect 678 5196 840 5198
rect 573 5168 614 5176
rect 696 5172 709 5196
rect 724 5194 739 5196
rect 536 5158 537 5168
rect 552 5158 565 5168
rect 579 5158 580 5168
rect 595 5158 608 5168
rect 623 5158 653 5172
rect 696 5158 739 5172
rect 763 5169 770 5176
rect 773 5172 840 5196
rect 872 5196 1044 5198
rect 842 5174 870 5178
rect 872 5174 952 5196
rect 973 5194 988 5196
rect 842 5172 952 5174
rect 773 5168 952 5172
rect 746 5158 776 5168
rect 778 5158 931 5168
rect 939 5158 969 5168
rect 973 5158 1003 5172
rect 1031 5158 1044 5196
rect 1116 5202 1151 5210
rect 1116 5176 1117 5202
rect 1124 5176 1151 5202
rect 1059 5158 1089 5172
rect 1116 5168 1151 5176
rect 1153 5202 1194 5210
rect 1153 5176 1168 5202
rect 1175 5176 1194 5202
rect 1258 5198 1320 5210
rect 1332 5198 1407 5210
rect 1465 5198 1540 5210
rect 1552 5198 1583 5210
rect 1589 5198 1624 5210
rect 1258 5196 1420 5198
rect 1153 5168 1194 5176
rect 1276 5172 1289 5196
rect 1304 5194 1319 5196
rect 1116 5158 1117 5168
rect 1132 5158 1145 5168
rect 1159 5158 1160 5168
rect 1175 5158 1188 5168
rect 1203 5158 1233 5172
rect 1276 5158 1319 5172
rect 1343 5169 1350 5176
rect 1353 5172 1420 5196
rect 1452 5196 1624 5198
rect 1422 5174 1450 5178
rect 1452 5174 1532 5196
rect 1553 5194 1568 5196
rect 1422 5172 1532 5174
rect 1353 5168 1532 5172
rect 1326 5158 1356 5168
rect 1358 5158 1511 5168
rect 1519 5158 1549 5168
rect 1553 5158 1583 5172
rect 1611 5158 1624 5196
rect 1696 5202 1731 5210
rect 1696 5176 1697 5202
rect 1704 5176 1731 5202
rect 1639 5158 1669 5172
rect 1696 5168 1731 5176
rect 1733 5202 1774 5210
rect 1733 5176 1748 5202
rect 1755 5176 1774 5202
rect 1838 5198 1900 5210
rect 1912 5198 1987 5210
rect 2045 5198 2120 5210
rect 2132 5198 2163 5210
rect 2169 5198 2204 5210
rect 1838 5196 2000 5198
rect 1733 5168 1774 5176
rect 1856 5172 1869 5196
rect 1884 5194 1899 5196
rect 1696 5158 1697 5168
rect 1712 5158 1725 5168
rect 1739 5158 1740 5168
rect 1755 5158 1768 5168
rect 1783 5158 1813 5172
rect 1856 5158 1899 5172
rect 1923 5169 1930 5176
rect 1933 5172 2000 5196
rect 2032 5196 2204 5198
rect 2002 5174 2030 5178
rect 2032 5174 2112 5196
rect 2133 5194 2148 5196
rect 2002 5172 2112 5174
rect 1933 5168 2112 5172
rect 1906 5158 1936 5168
rect 1938 5158 2091 5168
rect 2099 5158 2129 5168
rect 2133 5158 2163 5172
rect 2191 5158 2204 5196
rect 2276 5202 2311 5210
rect 2276 5176 2277 5202
rect 2284 5176 2311 5202
rect 2219 5158 2249 5172
rect 2276 5168 2311 5176
rect 2313 5202 2354 5210
rect 2313 5176 2328 5202
rect 2335 5176 2354 5202
rect 2418 5198 2480 5210
rect 2492 5198 2567 5210
rect 2625 5198 2700 5210
rect 2712 5198 2743 5210
rect 2749 5198 2784 5210
rect 2418 5196 2580 5198
rect 2313 5168 2354 5176
rect 2436 5172 2449 5196
rect 2464 5194 2479 5196
rect 2276 5158 2277 5168
rect 2292 5158 2305 5168
rect 2319 5158 2320 5168
rect 2335 5158 2348 5168
rect 2363 5158 2393 5172
rect 2436 5158 2479 5172
rect 2503 5169 2510 5176
rect 2513 5172 2580 5196
rect 2612 5196 2784 5198
rect 2582 5174 2610 5178
rect 2612 5174 2692 5196
rect 2713 5194 2728 5196
rect 2582 5172 2692 5174
rect 2513 5168 2692 5172
rect 2486 5158 2516 5168
rect 2518 5158 2671 5168
rect 2679 5158 2709 5168
rect 2713 5158 2743 5172
rect 2771 5158 2784 5196
rect 2856 5202 2891 5210
rect 2856 5176 2857 5202
rect 2864 5176 2891 5202
rect 2799 5158 2829 5172
rect 2856 5168 2891 5176
rect 2893 5202 2934 5210
rect 2893 5176 2908 5202
rect 2915 5176 2934 5202
rect 2998 5198 3060 5210
rect 3072 5198 3147 5210
rect 3205 5198 3280 5210
rect 3292 5198 3323 5210
rect 3329 5198 3364 5210
rect 2998 5196 3160 5198
rect 2893 5168 2934 5176
rect 3016 5172 3029 5196
rect 3044 5194 3059 5196
rect 2856 5158 2857 5168
rect 2872 5158 2885 5168
rect 2899 5158 2900 5168
rect 2915 5158 2928 5168
rect 2943 5158 2973 5172
rect 3016 5158 3059 5172
rect 3083 5169 3090 5176
rect 3093 5172 3160 5196
rect 3192 5196 3364 5198
rect 3162 5174 3190 5178
rect 3192 5174 3272 5196
rect 3293 5194 3308 5196
rect 3162 5172 3272 5174
rect 3093 5168 3272 5172
rect 3066 5158 3096 5168
rect 3098 5158 3251 5168
rect 3259 5158 3289 5168
rect 3293 5158 3323 5172
rect 3351 5158 3364 5196
rect 3436 5202 3471 5210
rect 3436 5176 3437 5202
rect 3444 5176 3471 5202
rect 3379 5158 3409 5172
rect 3436 5168 3471 5176
rect 3473 5202 3514 5210
rect 3473 5176 3488 5202
rect 3495 5176 3514 5202
rect 3578 5198 3640 5210
rect 3652 5198 3727 5210
rect 3785 5198 3860 5210
rect 3872 5198 3903 5210
rect 3909 5198 3944 5210
rect 3578 5196 3740 5198
rect 3473 5168 3514 5176
rect 3596 5172 3609 5196
rect 3624 5194 3639 5196
rect 3436 5158 3437 5168
rect 3452 5158 3465 5168
rect 3479 5158 3480 5168
rect 3495 5158 3508 5168
rect 3523 5158 3553 5172
rect 3596 5158 3639 5172
rect 3663 5169 3670 5176
rect 3673 5172 3740 5196
rect 3772 5196 3944 5198
rect 3742 5174 3770 5178
rect 3772 5174 3852 5196
rect 3873 5194 3888 5196
rect 3742 5172 3852 5174
rect 3673 5168 3852 5172
rect 3646 5158 3676 5168
rect 3678 5158 3831 5168
rect 3839 5158 3869 5168
rect 3873 5158 3903 5172
rect 3931 5158 3944 5196
rect 4016 5202 4051 5210
rect 4016 5176 4017 5202
rect 4024 5176 4051 5202
rect 3959 5158 3989 5172
rect 4016 5168 4051 5176
rect 4053 5202 4094 5210
rect 4053 5176 4068 5202
rect 4075 5176 4094 5202
rect 4158 5198 4220 5210
rect 4232 5198 4307 5210
rect 4365 5198 4440 5210
rect 4452 5198 4483 5210
rect 4489 5198 4524 5210
rect 4158 5196 4320 5198
rect 4053 5168 4094 5176
rect 4176 5172 4189 5196
rect 4204 5194 4219 5196
rect 4016 5158 4017 5168
rect 4032 5158 4045 5168
rect 4059 5158 4060 5168
rect 4075 5158 4088 5168
rect 4103 5158 4133 5172
rect 4176 5158 4219 5172
rect 4243 5169 4250 5176
rect 4253 5172 4320 5196
rect 4352 5196 4524 5198
rect 4322 5174 4350 5178
rect 4352 5174 4432 5196
rect 4453 5194 4468 5196
rect 4322 5172 4432 5174
rect 4253 5168 4432 5172
rect 4226 5158 4256 5168
rect 4258 5158 4411 5168
rect 4419 5158 4449 5168
rect 4453 5158 4483 5172
rect 4511 5158 4524 5196
rect 4596 5202 4631 5210
rect 4596 5176 4597 5202
rect 4604 5176 4631 5202
rect 4539 5158 4569 5172
rect 4596 5168 4631 5176
rect 4633 5202 4674 5210
rect 4633 5176 4648 5202
rect 4655 5176 4674 5202
rect 4738 5198 4800 5210
rect 4812 5198 4887 5210
rect 4945 5198 5020 5210
rect 5032 5198 5063 5210
rect 5069 5198 5104 5210
rect 4738 5196 4900 5198
rect 4633 5168 4674 5176
rect 4756 5172 4769 5196
rect 4784 5194 4799 5196
rect 4596 5158 4597 5168
rect 4612 5158 4625 5168
rect 4639 5158 4640 5168
rect 4655 5158 4668 5168
rect 4683 5158 4713 5172
rect 4756 5158 4799 5172
rect 4823 5169 4830 5176
rect 4833 5172 4900 5196
rect 4932 5196 5104 5198
rect 4902 5174 4930 5178
rect 4932 5174 5012 5196
rect 5033 5194 5048 5196
rect 4902 5172 5012 5174
rect 4833 5168 5012 5172
rect 4806 5158 4836 5168
rect 4838 5158 4991 5168
rect 4999 5158 5029 5168
rect 5033 5158 5063 5172
rect 5091 5158 5104 5196
rect 5176 5202 5211 5210
rect 5176 5176 5177 5202
rect 5184 5176 5211 5202
rect 5119 5158 5149 5172
rect 5176 5168 5211 5176
rect 5213 5202 5254 5210
rect 5213 5176 5228 5202
rect 5235 5176 5254 5202
rect 5318 5198 5380 5210
rect 5392 5198 5467 5210
rect 5525 5198 5600 5210
rect 5612 5198 5643 5210
rect 5649 5198 5684 5210
rect 5318 5196 5480 5198
rect 5213 5168 5254 5176
rect 5336 5172 5349 5196
rect 5364 5194 5379 5196
rect 5176 5158 5177 5168
rect 5192 5158 5205 5168
rect 5219 5158 5220 5168
rect 5235 5158 5248 5168
rect 5263 5158 5293 5172
rect 5336 5158 5379 5172
rect 5403 5169 5410 5176
rect 5413 5172 5480 5196
rect 5512 5196 5684 5198
rect 5482 5174 5510 5178
rect 5512 5174 5592 5196
rect 5613 5194 5628 5196
rect 5482 5172 5592 5174
rect 5413 5168 5592 5172
rect 5386 5158 5416 5168
rect 5418 5158 5571 5168
rect 5579 5158 5609 5168
rect 5613 5158 5643 5172
rect 5671 5158 5684 5196
rect 5756 5202 5791 5210
rect 5756 5176 5757 5202
rect 5764 5176 5791 5202
rect 5699 5158 5729 5172
rect 5756 5168 5791 5176
rect 5793 5202 5834 5210
rect 5793 5176 5808 5202
rect 5815 5176 5834 5202
rect 5898 5198 5960 5210
rect 5972 5198 6047 5210
rect 6105 5198 6180 5210
rect 6192 5198 6223 5210
rect 6229 5198 6264 5210
rect 5898 5196 6060 5198
rect 5793 5168 5834 5176
rect 5916 5172 5929 5196
rect 5944 5194 5959 5196
rect 5756 5158 5757 5168
rect 5772 5158 5785 5168
rect 5799 5158 5800 5168
rect 5815 5158 5828 5168
rect 5843 5158 5873 5172
rect 5916 5158 5959 5172
rect 5983 5169 5990 5176
rect 5993 5172 6060 5196
rect 6092 5196 6264 5198
rect 6062 5174 6090 5178
rect 6092 5174 6172 5196
rect 6193 5194 6208 5196
rect 6062 5172 6172 5174
rect 5993 5168 6172 5172
rect 5966 5158 5996 5168
rect 5998 5158 6151 5168
rect 6159 5158 6189 5168
rect 6193 5158 6223 5172
rect 6251 5158 6264 5196
rect 6336 5202 6371 5210
rect 6336 5176 6337 5202
rect 6344 5176 6371 5202
rect 6279 5158 6309 5172
rect 6336 5168 6371 5176
rect 6373 5202 6414 5210
rect 6373 5176 6388 5202
rect 6395 5176 6414 5202
rect 6478 5198 6540 5210
rect 6552 5198 6627 5210
rect 6685 5198 6760 5210
rect 6772 5198 6803 5210
rect 6809 5198 6844 5210
rect 6478 5196 6640 5198
rect 6373 5168 6414 5176
rect 6496 5172 6509 5196
rect 6524 5194 6539 5196
rect 6336 5158 6337 5168
rect 6352 5158 6365 5168
rect 6379 5158 6380 5168
rect 6395 5158 6408 5168
rect 6423 5158 6453 5172
rect 6496 5158 6539 5172
rect 6563 5169 6570 5176
rect 6573 5172 6640 5196
rect 6672 5196 6844 5198
rect 6642 5174 6670 5178
rect 6672 5174 6752 5196
rect 6773 5194 6788 5196
rect 6642 5172 6752 5174
rect 6573 5168 6752 5172
rect 6546 5158 6576 5168
rect 6578 5158 6731 5168
rect 6739 5158 6769 5168
rect 6773 5158 6803 5172
rect 6831 5158 6844 5196
rect 6916 5202 6951 5210
rect 6916 5176 6917 5202
rect 6924 5176 6951 5202
rect 6859 5158 6889 5172
rect 6916 5168 6951 5176
rect 6953 5202 6994 5210
rect 6953 5176 6968 5202
rect 6975 5176 6994 5202
rect 7058 5198 7120 5210
rect 7132 5198 7207 5210
rect 7265 5198 7340 5210
rect 7352 5198 7383 5210
rect 7389 5198 7424 5210
rect 7058 5196 7220 5198
rect 6953 5168 6994 5176
rect 7076 5172 7089 5196
rect 7104 5194 7119 5196
rect 6916 5158 6917 5168
rect 6932 5158 6945 5168
rect 6959 5158 6960 5168
rect 6975 5158 6988 5168
rect 7003 5158 7033 5172
rect 7076 5158 7119 5172
rect 7143 5169 7150 5176
rect 7153 5172 7220 5196
rect 7252 5196 7424 5198
rect 7222 5174 7250 5178
rect 7252 5174 7332 5196
rect 7353 5194 7368 5196
rect 7222 5172 7332 5174
rect 7153 5168 7332 5172
rect 7126 5158 7156 5168
rect 7158 5158 7311 5168
rect 7319 5158 7349 5168
rect 7353 5158 7383 5172
rect 7411 5158 7424 5196
rect 7496 5202 7531 5210
rect 7496 5176 7497 5202
rect 7504 5176 7531 5202
rect 7439 5158 7469 5172
rect 7496 5168 7531 5176
rect 7533 5202 7574 5210
rect 7533 5176 7548 5202
rect 7555 5176 7574 5202
rect 7638 5198 7700 5210
rect 7712 5198 7787 5210
rect 7845 5198 7920 5210
rect 7932 5198 7963 5210
rect 7969 5198 8004 5210
rect 7638 5196 7800 5198
rect 7533 5168 7574 5176
rect 7656 5172 7669 5196
rect 7684 5194 7699 5196
rect 7496 5158 7497 5168
rect 7512 5158 7525 5168
rect 7539 5158 7540 5168
rect 7555 5158 7568 5168
rect 7583 5158 7613 5172
rect 7656 5158 7699 5172
rect 7723 5169 7730 5176
rect 7733 5172 7800 5196
rect 7832 5196 8004 5198
rect 7802 5174 7830 5178
rect 7832 5174 7912 5196
rect 7933 5194 7948 5196
rect 7802 5172 7912 5174
rect 7733 5168 7912 5172
rect 7706 5158 7736 5168
rect 7738 5158 7891 5168
rect 7899 5158 7929 5168
rect 7933 5158 7963 5172
rect 7991 5158 8004 5196
rect 8076 5202 8111 5210
rect 8076 5176 8077 5202
rect 8084 5176 8111 5202
rect 8019 5158 8049 5172
rect 8076 5168 8111 5176
rect 8113 5202 8154 5210
rect 8113 5176 8128 5202
rect 8135 5176 8154 5202
rect 8218 5198 8280 5210
rect 8292 5198 8367 5210
rect 8425 5198 8500 5210
rect 8512 5198 8543 5210
rect 8549 5198 8584 5210
rect 8218 5196 8380 5198
rect 8113 5168 8154 5176
rect 8236 5172 8249 5196
rect 8264 5194 8279 5196
rect 8076 5158 8077 5168
rect 8092 5158 8105 5168
rect 8119 5158 8120 5168
rect 8135 5158 8148 5168
rect 8163 5158 8193 5172
rect 8236 5158 8279 5172
rect 8303 5169 8310 5176
rect 8313 5172 8380 5196
rect 8412 5196 8584 5198
rect 8382 5174 8410 5178
rect 8412 5174 8492 5196
rect 8513 5194 8528 5196
rect 8382 5172 8492 5174
rect 8313 5168 8492 5172
rect 8286 5158 8316 5168
rect 8318 5158 8471 5168
rect 8479 5158 8509 5168
rect 8513 5158 8543 5172
rect 8571 5158 8584 5196
rect 8656 5202 8691 5210
rect 8656 5176 8657 5202
rect 8664 5176 8691 5202
rect 8599 5158 8629 5172
rect 8656 5168 8691 5176
rect 8693 5202 8734 5210
rect 8693 5176 8708 5202
rect 8715 5176 8734 5202
rect 8798 5198 8860 5210
rect 8872 5198 8947 5210
rect 9005 5198 9080 5210
rect 9092 5198 9123 5210
rect 9129 5198 9164 5210
rect 8798 5196 8960 5198
rect 8693 5168 8734 5176
rect 8816 5172 8829 5196
rect 8844 5194 8859 5196
rect 8656 5158 8657 5168
rect 8672 5158 8685 5168
rect 8699 5158 8700 5168
rect 8715 5158 8728 5168
rect 8743 5158 8773 5172
rect 8816 5158 8859 5172
rect 8883 5169 8890 5176
rect 8893 5172 8960 5196
rect 8992 5196 9164 5198
rect 8962 5174 8990 5178
rect 8992 5174 9072 5196
rect 9093 5194 9108 5196
rect 8962 5172 9072 5174
rect 8893 5168 9072 5172
rect 8866 5158 8896 5168
rect 8898 5158 9051 5168
rect 9059 5158 9089 5168
rect 9093 5158 9123 5172
rect 9151 5158 9164 5196
rect 9236 5202 9271 5210
rect 9236 5176 9237 5202
rect 9244 5176 9271 5202
rect 9179 5158 9209 5172
rect 9236 5168 9271 5176
rect 9236 5158 9237 5168
rect 9252 5158 9265 5168
rect -1 5152 9265 5158
rect 0 5144 9265 5152
rect 15 5114 28 5144
rect 43 5126 73 5144
rect 116 5130 130 5144
rect 166 5130 386 5144
rect 117 5128 130 5130
rect 83 5116 98 5128
rect 80 5114 102 5116
rect 107 5114 137 5128
rect 198 5126 351 5130
rect 180 5114 372 5126
rect 415 5114 445 5128
rect 451 5114 464 5144
rect 479 5126 509 5144
rect 552 5114 565 5144
rect 595 5114 608 5144
rect 623 5126 653 5144
rect 696 5130 710 5144
rect 746 5130 966 5144
rect 697 5128 710 5130
rect 663 5116 678 5128
rect 660 5114 682 5116
rect 687 5114 717 5128
rect 778 5126 931 5130
rect 760 5114 952 5126
rect 995 5114 1025 5128
rect 1031 5114 1044 5144
rect 1059 5126 1089 5144
rect 1132 5114 1145 5144
rect 1175 5114 1188 5144
rect 1203 5126 1233 5144
rect 1276 5130 1290 5144
rect 1326 5130 1546 5144
rect 1277 5128 1290 5130
rect 1243 5116 1258 5128
rect 1240 5114 1262 5116
rect 1267 5114 1297 5128
rect 1358 5126 1511 5130
rect 1340 5114 1532 5126
rect 1575 5114 1605 5128
rect 1611 5114 1624 5144
rect 1639 5126 1669 5144
rect 1712 5114 1725 5144
rect 1755 5114 1768 5144
rect 1783 5126 1813 5144
rect 1856 5130 1870 5144
rect 1906 5130 2126 5144
rect 1857 5128 1870 5130
rect 1823 5116 1838 5128
rect 1820 5114 1842 5116
rect 1847 5114 1877 5128
rect 1938 5126 2091 5130
rect 1920 5114 2112 5126
rect 2155 5114 2185 5128
rect 2191 5114 2204 5144
rect 2219 5126 2249 5144
rect 2292 5114 2305 5144
rect 2335 5114 2348 5144
rect 2363 5126 2393 5144
rect 2436 5130 2450 5144
rect 2486 5130 2706 5144
rect 2437 5128 2450 5130
rect 2403 5116 2418 5128
rect 2400 5114 2422 5116
rect 2427 5114 2457 5128
rect 2518 5126 2671 5130
rect 2500 5114 2692 5126
rect 2735 5114 2765 5128
rect 2771 5114 2784 5144
rect 2799 5126 2829 5144
rect 2872 5114 2885 5144
rect 2915 5114 2928 5144
rect 2943 5126 2973 5144
rect 3016 5130 3030 5144
rect 3066 5130 3286 5144
rect 3017 5128 3030 5130
rect 2983 5116 2998 5128
rect 2980 5114 3002 5116
rect 3007 5114 3037 5128
rect 3098 5126 3251 5130
rect 3080 5114 3272 5126
rect 3315 5114 3345 5128
rect 3351 5114 3364 5144
rect 3379 5126 3409 5144
rect 3452 5114 3465 5144
rect 3495 5114 3508 5144
rect 3523 5126 3553 5144
rect 3596 5130 3610 5144
rect 3646 5130 3866 5144
rect 3597 5128 3610 5130
rect 3563 5116 3578 5128
rect 3560 5114 3582 5116
rect 3587 5114 3617 5128
rect 3678 5126 3831 5130
rect 3660 5114 3852 5126
rect 3895 5114 3925 5128
rect 3931 5114 3944 5144
rect 3959 5126 3989 5144
rect 4032 5114 4045 5144
rect 4075 5114 4088 5144
rect 4103 5126 4133 5144
rect 4176 5130 4190 5144
rect 4226 5130 4446 5144
rect 4177 5128 4190 5130
rect 4143 5116 4158 5128
rect 4140 5114 4162 5116
rect 4167 5114 4197 5128
rect 4258 5126 4411 5130
rect 4240 5114 4432 5126
rect 4475 5114 4505 5128
rect 4511 5114 4524 5144
rect 4539 5126 4569 5144
rect 4612 5114 4625 5144
rect 4655 5114 4668 5144
rect 4683 5126 4713 5144
rect 4756 5130 4770 5144
rect 4806 5130 5026 5144
rect 4757 5128 4770 5130
rect 4723 5116 4738 5128
rect 4720 5114 4742 5116
rect 4747 5114 4777 5128
rect 4838 5126 4991 5130
rect 4820 5114 5012 5126
rect 5055 5114 5085 5128
rect 5091 5114 5104 5144
rect 5119 5126 5149 5144
rect 5192 5114 5205 5144
rect 5235 5114 5248 5144
rect 5263 5126 5293 5144
rect 5336 5130 5350 5144
rect 5386 5130 5606 5144
rect 5337 5128 5350 5130
rect 5303 5116 5318 5128
rect 5300 5114 5322 5116
rect 5327 5114 5357 5128
rect 5418 5126 5571 5130
rect 5400 5114 5592 5126
rect 5635 5114 5665 5128
rect 5671 5114 5684 5144
rect 5699 5126 5729 5144
rect 5772 5114 5785 5144
rect 5815 5114 5828 5144
rect 5843 5126 5873 5144
rect 5916 5130 5930 5144
rect 5966 5130 6186 5144
rect 5917 5128 5930 5130
rect 5883 5116 5898 5128
rect 5880 5114 5902 5116
rect 5907 5114 5937 5128
rect 5998 5126 6151 5130
rect 5980 5114 6172 5126
rect 6215 5114 6245 5128
rect 6251 5114 6264 5144
rect 6279 5126 6309 5144
rect 6352 5114 6365 5144
rect 6395 5114 6408 5144
rect 6423 5126 6453 5144
rect 6496 5130 6510 5144
rect 6546 5130 6766 5144
rect 6497 5128 6510 5130
rect 6463 5116 6478 5128
rect 6460 5114 6482 5116
rect 6487 5114 6517 5128
rect 6578 5126 6731 5130
rect 6560 5114 6752 5126
rect 6795 5114 6825 5128
rect 6831 5114 6844 5144
rect 6859 5126 6889 5144
rect 6932 5114 6945 5144
rect 6975 5114 6988 5144
rect 7003 5126 7033 5144
rect 7076 5130 7090 5144
rect 7126 5130 7346 5144
rect 7077 5128 7090 5130
rect 7043 5116 7058 5128
rect 7040 5114 7062 5116
rect 7067 5114 7097 5128
rect 7158 5126 7311 5130
rect 7140 5114 7332 5126
rect 7375 5114 7405 5128
rect 7411 5114 7424 5144
rect 7439 5126 7469 5144
rect 7512 5114 7525 5144
rect 7555 5114 7568 5144
rect 7583 5126 7613 5144
rect 7656 5130 7670 5144
rect 7706 5130 7926 5144
rect 7657 5128 7670 5130
rect 7623 5116 7638 5128
rect 7620 5114 7642 5116
rect 7647 5114 7677 5128
rect 7738 5126 7891 5130
rect 7720 5114 7912 5126
rect 7955 5114 7985 5128
rect 7991 5114 8004 5144
rect 8019 5126 8049 5144
rect 8092 5114 8105 5144
rect 8135 5114 8148 5144
rect 8163 5126 8193 5144
rect 8236 5130 8250 5144
rect 8286 5130 8506 5144
rect 8237 5128 8250 5130
rect 8203 5116 8218 5128
rect 8200 5114 8222 5116
rect 8227 5114 8257 5128
rect 8318 5126 8471 5130
rect 8300 5114 8492 5126
rect 8535 5114 8565 5128
rect 8571 5114 8584 5144
rect 8599 5126 8629 5144
rect 8672 5114 8685 5144
rect 8715 5114 8728 5144
rect 8743 5126 8773 5144
rect 8816 5130 8830 5144
rect 8866 5130 9086 5144
rect 8817 5128 8830 5130
rect 8783 5116 8798 5128
rect 8780 5114 8802 5116
rect 8807 5114 8837 5128
rect 8898 5126 9051 5130
rect 8880 5114 9072 5126
rect 9115 5114 9145 5128
rect 9151 5114 9164 5144
rect 9179 5126 9209 5144
rect 9252 5114 9265 5144
rect 0 5100 9265 5114
rect 15 4996 28 5100
rect 73 5078 74 5088
rect 89 5078 102 5088
rect 73 5074 102 5078
rect 107 5074 137 5100
rect 155 5086 171 5088
rect 243 5086 296 5100
rect 244 5084 308 5086
rect 351 5084 366 5100
rect 415 5097 445 5100
rect 415 5094 451 5097
rect 381 5086 397 5088
rect 155 5074 170 5078
rect 73 5072 170 5074
rect 198 5072 366 5084
rect 382 5074 397 5078
rect 415 5075 454 5094
rect 473 5088 480 5089
rect 479 5081 480 5088
rect 463 5078 464 5081
rect 479 5078 492 5081
rect 415 5074 445 5075
rect 454 5074 460 5075
rect 463 5074 492 5078
rect 382 5073 492 5074
rect 382 5072 498 5073
rect 57 5064 108 5072
rect 57 5052 82 5064
rect 89 5052 108 5064
rect 139 5064 189 5072
rect 139 5056 155 5064
rect 162 5062 189 5064
rect 198 5062 419 5072
rect 162 5052 419 5062
rect 448 5064 498 5072
rect 448 5055 464 5064
rect 57 5044 108 5052
rect 155 5044 419 5052
rect 445 5052 464 5055
rect 471 5052 498 5064
rect 445 5044 498 5052
rect 73 5036 74 5044
rect 89 5036 102 5044
rect 73 5028 89 5036
rect 70 5021 89 5024
rect 70 5012 92 5021
rect 43 5002 92 5012
rect 43 4996 73 5002
rect 92 4997 97 5002
rect 15 4980 89 4996
rect 107 4988 137 5044
rect 172 5034 380 5044
rect 415 5040 460 5044
rect 463 5043 464 5044
rect 479 5043 492 5044
rect 198 5004 387 5034
rect 213 5001 387 5004
rect 206 4998 387 5001
rect 15 4978 28 4980
rect 43 4978 77 4980
rect 15 4962 89 4978
rect 116 4974 129 4988
rect 144 4974 160 4990
rect 206 4985 217 4998
rect -1 4940 0 4956
rect 15 4940 28 4962
rect 43 4940 73 4962
rect 116 4958 178 4974
rect 206 4967 217 4983
rect 222 4978 232 4998
rect 242 4978 256 4998
rect 259 4985 268 4998
rect 284 4985 293 4998
rect 222 4967 256 4978
rect 259 4967 268 4983
rect 284 4967 293 4983
rect 300 4978 310 4998
rect 320 4978 334 4998
rect 335 4985 346 4998
rect 300 4967 334 4978
rect 335 4967 346 4983
rect 392 4974 408 4990
rect 415 4988 445 5040
rect 479 5036 480 5043
rect 464 5028 480 5036
rect 451 4996 464 5015
rect 479 4996 509 5012
rect 451 4980 525 4996
rect 451 4978 464 4980
rect 479 4978 513 4980
rect 116 4956 129 4958
rect 144 4956 178 4958
rect 116 4940 178 4956
rect 222 4951 238 4954
rect 300 4951 330 4962
rect 378 4958 424 4974
rect 451 4962 525 4978
rect 378 4956 412 4958
rect 377 4940 424 4956
rect 451 4940 464 4962
rect 479 4940 509 4962
rect 536 4940 537 4956
rect 552 4940 565 5100
rect 595 4996 608 5100
rect 653 5078 654 5088
rect 669 5078 682 5088
rect 653 5074 682 5078
rect 687 5074 717 5100
rect 735 5086 751 5088
rect 823 5086 876 5100
rect 824 5084 888 5086
rect 931 5084 946 5100
rect 995 5097 1025 5100
rect 995 5094 1031 5097
rect 961 5086 977 5088
rect 735 5074 750 5078
rect 653 5072 750 5074
rect 778 5072 946 5084
rect 962 5074 977 5078
rect 995 5075 1034 5094
rect 1053 5088 1060 5089
rect 1059 5081 1060 5088
rect 1043 5078 1044 5081
rect 1059 5078 1072 5081
rect 995 5074 1025 5075
rect 1034 5074 1040 5075
rect 1043 5074 1072 5078
rect 962 5073 1072 5074
rect 962 5072 1078 5073
rect 637 5064 688 5072
rect 637 5052 662 5064
rect 669 5052 688 5064
rect 719 5064 769 5072
rect 719 5056 735 5064
rect 742 5062 769 5064
rect 778 5062 999 5072
rect 742 5052 999 5062
rect 1028 5064 1078 5072
rect 1028 5055 1044 5064
rect 637 5044 688 5052
rect 735 5044 999 5052
rect 1025 5052 1044 5055
rect 1051 5052 1078 5064
rect 1025 5044 1078 5052
rect 653 5036 654 5044
rect 669 5036 682 5044
rect 653 5028 669 5036
rect 650 5021 669 5024
rect 650 5012 672 5021
rect 623 5002 672 5012
rect 623 4996 653 5002
rect 672 4997 677 5002
rect 595 4980 669 4996
rect 687 4988 717 5044
rect 752 5034 960 5044
rect 995 5040 1040 5044
rect 1043 5043 1044 5044
rect 1059 5043 1072 5044
rect 778 5004 967 5034
rect 793 5001 967 5004
rect 786 4998 967 5001
rect 595 4978 608 4980
rect 623 4978 657 4980
rect 595 4962 669 4978
rect 696 4974 709 4988
rect 724 4974 740 4990
rect 786 4985 797 4998
rect 579 4940 580 4956
rect 595 4940 608 4962
rect 623 4940 653 4962
rect 696 4958 758 4974
rect 786 4967 797 4983
rect 802 4978 812 4998
rect 822 4978 836 4998
rect 839 4985 848 4998
rect 864 4985 873 4998
rect 802 4967 836 4978
rect 839 4967 848 4983
rect 864 4967 873 4983
rect 880 4978 890 4998
rect 900 4978 914 4998
rect 915 4985 926 4998
rect 880 4967 914 4978
rect 915 4967 926 4983
rect 972 4974 988 4990
rect 995 4988 1025 5040
rect 1059 5036 1060 5043
rect 1044 5028 1060 5036
rect 1031 4996 1044 5015
rect 1059 4996 1089 5012
rect 1031 4980 1105 4996
rect 1031 4978 1044 4980
rect 1059 4978 1093 4980
rect 696 4956 709 4958
rect 724 4956 758 4958
rect 696 4940 758 4956
rect 802 4951 818 4954
rect 880 4951 910 4962
rect 958 4958 1004 4974
rect 1031 4962 1105 4978
rect 958 4956 992 4958
rect 957 4940 1004 4956
rect 1031 4940 1044 4962
rect 1059 4940 1089 4962
rect 1116 4940 1117 4956
rect 1132 4940 1145 5100
rect 1175 4996 1188 5100
rect 1233 5078 1234 5088
rect 1249 5078 1262 5088
rect 1233 5074 1262 5078
rect 1267 5074 1297 5100
rect 1315 5086 1331 5088
rect 1403 5086 1456 5100
rect 1404 5084 1468 5086
rect 1511 5084 1526 5100
rect 1575 5097 1605 5100
rect 1575 5094 1611 5097
rect 1541 5086 1557 5088
rect 1315 5074 1330 5078
rect 1233 5072 1330 5074
rect 1358 5072 1526 5084
rect 1542 5074 1557 5078
rect 1575 5075 1614 5094
rect 1633 5088 1640 5089
rect 1639 5081 1640 5088
rect 1623 5078 1624 5081
rect 1639 5078 1652 5081
rect 1575 5074 1605 5075
rect 1614 5074 1620 5075
rect 1623 5074 1652 5078
rect 1542 5073 1652 5074
rect 1542 5072 1658 5073
rect 1217 5064 1268 5072
rect 1217 5052 1242 5064
rect 1249 5052 1268 5064
rect 1299 5064 1349 5072
rect 1299 5056 1315 5064
rect 1322 5062 1349 5064
rect 1358 5062 1579 5072
rect 1322 5052 1579 5062
rect 1608 5064 1658 5072
rect 1608 5055 1624 5064
rect 1217 5044 1268 5052
rect 1315 5044 1579 5052
rect 1605 5052 1624 5055
rect 1631 5052 1658 5064
rect 1605 5044 1658 5052
rect 1233 5036 1234 5044
rect 1249 5036 1262 5044
rect 1233 5028 1249 5036
rect 1230 5021 1249 5024
rect 1230 5012 1252 5021
rect 1203 5002 1252 5012
rect 1203 4996 1233 5002
rect 1252 4997 1257 5002
rect 1175 4980 1249 4996
rect 1267 4988 1297 5044
rect 1332 5034 1540 5044
rect 1575 5040 1620 5044
rect 1623 5043 1624 5044
rect 1639 5043 1652 5044
rect 1358 5004 1547 5034
rect 1373 5001 1547 5004
rect 1366 4998 1547 5001
rect 1175 4978 1188 4980
rect 1203 4978 1237 4980
rect 1175 4962 1249 4978
rect 1276 4974 1289 4988
rect 1304 4974 1320 4990
rect 1366 4985 1377 4998
rect 1159 4940 1160 4956
rect 1175 4940 1188 4962
rect 1203 4940 1233 4962
rect 1276 4958 1338 4974
rect 1366 4967 1377 4983
rect 1382 4978 1392 4998
rect 1402 4978 1416 4998
rect 1419 4985 1428 4998
rect 1444 4985 1453 4998
rect 1382 4967 1416 4978
rect 1419 4967 1428 4983
rect 1444 4967 1453 4983
rect 1460 4978 1470 4998
rect 1480 4978 1494 4998
rect 1495 4985 1506 4998
rect 1460 4967 1494 4978
rect 1495 4967 1506 4983
rect 1552 4974 1568 4990
rect 1575 4988 1605 5040
rect 1639 5036 1640 5043
rect 1624 5028 1640 5036
rect 1611 4996 1624 5015
rect 1639 4996 1669 5012
rect 1611 4980 1685 4996
rect 1611 4978 1624 4980
rect 1639 4978 1673 4980
rect 1276 4956 1289 4958
rect 1304 4956 1338 4958
rect 1276 4940 1338 4956
rect 1382 4951 1398 4954
rect 1460 4951 1490 4962
rect 1538 4958 1584 4974
rect 1611 4962 1685 4978
rect 1538 4956 1572 4958
rect 1537 4940 1584 4956
rect 1611 4940 1624 4962
rect 1639 4940 1669 4962
rect 1696 4940 1697 4956
rect 1712 4940 1725 5100
rect 1755 4996 1768 5100
rect 1813 5078 1814 5088
rect 1829 5078 1842 5088
rect 1813 5074 1842 5078
rect 1847 5074 1877 5100
rect 1895 5086 1911 5088
rect 1983 5086 2036 5100
rect 1984 5084 2048 5086
rect 2091 5084 2106 5100
rect 2155 5097 2185 5100
rect 2155 5094 2191 5097
rect 2121 5086 2137 5088
rect 1895 5074 1910 5078
rect 1813 5072 1910 5074
rect 1938 5072 2106 5084
rect 2122 5074 2137 5078
rect 2155 5075 2194 5094
rect 2213 5088 2220 5089
rect 2219 5081 2220 5088
rect 2203 5078 2204 5081
rect 2219 5078 2232 5081
rect 2155 5074 2185 5075
rect 2194 5074 2200 5075
rect 2203 5074 2232 5078
rect 2122 5073 2232 5074
rect 2122 5072 2238 5073
rect 1797 5064 1848 5072
rect 1797 5052 1822 5064
rect 1829 5052 1848 5064
rect 1879 5064 1929 5072
rect 1879 5056 1895 5064
rect 1902 5062 1929 5064
rect 1938 5062 2159 5072
rect 1902 5052 2159 5062
rect 2188 5064 2238 5072
rect 2188 5055 2204 5064
rect 1797 5044 1848 5052
rect 1895 5044 2159 5052
rect 2185 5052 2204 5055
rect 2211 5052 2238 5064
rect 2185 5044 2238 5052
rect 1813 5036 1814 5044
rect 1829 5036 1842 5044
rect 1813 5028 1829 5036
rect 1810 5021 1829 5024
rect 1810 5012 1832 5021
rect 1783 5002 1832 5012
rect 1783 4996 1813 5002
rect 1832 4997 1837 5002
rect 1755 4980 1829 4996
rect 1847 4988 1877 5044
rect 1912 5034 2120 5044
rect 2155 5040 2200 5044
rect 2203 5043 2204 5044
rect 2219 5043 2232 5044
rect 1938 5004 2127 5034
rect 1953 5001 2127 5004
rect 1946 4998 2127 5001
rect 1755 4978 1768 4980
rect 1783 4978 1817 4980
rect 1755 4962 1829 4978
rect 1856 4974 1869 4988
rect 1884 4974 1900 4990
rect 1946 4985 1957 4998
rect 1739 4940 1740 4956
rect 1755 4940 1768 4962
rect 1783 4940 1813 4962
rect 1856 4958 1918 4974
rect 1946 4967 1957 4983
rect 1962 4978 1972 4998
rect 1982 4978 1996 4998
rect 1999 4985 2008 4998
rect 2024 4985 2033 4998
rect 1962 4967 1996 4978
rect 1999 4967 2008 4983
rect 2024 4967 2033 4983
rect 2040 4978 2050 4998
rect 2060 4978 2074 4998
rect 2075 4985 2086 4998
rect 2040 4967 2074 4978
rect 2075 4967 2086 4983
rect 2132 4974 2148 4990
rect 2155 4988 2185 5040
rect 2219 5036 2220 5043
rect 2204 5028 2220 5036
rect 2191 4996 2204 5015
rect 2219 4996 2249 5012
rect 2191 4980 2265 4996
rect 2191 4978 2204 4980
rect 2219 4978 2253 4980
rect 1856 4956 1869 4958
rect 1884 4956 1918 4958
rect 1856 4940 1918 4956
rect 1962 4951 1976 4954
rect 2040 4951 2070 4962
rect 2118 4958 2164 4974
rect 2191 4962 2265 4978
rect 2118 4956 2152 4958
rect 2117 4940 2164 4956
rect 2191 4940 2204 4962
rect 2219 4940 2249 4962
rect 2276 4940 2277 4956
rect 2292 4940 2305 5100
rect 2335 4996 2348 5100
rect 2393 5078 2394 5088
rect 2409 5078 2422 5088
rect 2393 5074 2422 5078
rect 2427 5074 2457 5100
rect 2475 5086 2491 5088
rect 2563 5086 2616 5100
rect 2564 5084 2628 5086
rect 2671 5084 2686 5100
rect 2735 5097 2765 5100
rect 2735 5094 2771 5097
rect 2701 5086 2717 5088
rect 2475 5074 2490 5078
rect 2393 5072 2490 5074
rect 2518 5072 2686 5084
rect 2702 5074 2717 5078
rect 2735 5075 2774 5094
rect 2793 5088 2800 5089
rect 2799 5081 2800 5088
rect 2783 5078 2784 5081
rect 2799 5078 2812 5081
rect 2735 5074 2765 5075
rect 2774 5074 2780 5075
rect 2783 5074 2812 5078
rect 2702 5073 2812 5074
rect 2702 5072 2818 5073
rect 2377 5064 2428 5072
rect 2377 5052 2402 5064
rect 2409 5052 2428 5064
rect 2459 5064 2509 5072
rect 2459 5056 2475 5064
rect 2482 5062 2509 5064
rect 2518 5062 2739 5072
rect 2482 5052 2739 5062
rect 2768 5064 2818 5072
rect 2768 5055 2784 5064
rect 2377 5044 2428 5052
rect 2475 5044 2739 5052
rect 2765 5052 2784 5055
rect 2791 5052 2818 5064
rect 2765 5044 2818 5052
rect 2393 5036 2394 5044
rect 2409 5036 2422 5044
rect 2393 5028 2409 5036
rect 2390 5021 2409 5024
rect 2390 5012 2412 5021
rect 2363 5002 2412 5012
rect 2363 4996 2393 5002
rect 2412 4997 2417 5002
rect 2335 4980 2409 4996
rect 2427 4988 2457 5044
rect 2492 5034 2700 5044
rect 2735 5040 2780 5044
rect 2783 5043 2784 5044
rect 2799 5043 2812 5044
rect 2518 5004 2707 5034
rect 2533 5001 2707 5004
rect 2526 4998 2707 5001
rect 2335 4978 2348 4980
rect 2363 4978 2397 4980
rect 2335 4962 2409 4978
rect 2436 4974 2449 4988
rect 2464 4974 2480 4990
rect 2526 4985 2537 4998
rect 2319 4940 2320 4956
rect 2335 4940 2348 4962
rect 2363 4940 2393 4962
rect 2436 4958 2498 4974
rect 2526 4967 2537 4983
rect 2542 4978 2552 4998
rect 2562 4978 2576 4998
rect 2579 4985 2588 4998
rect 2604 4985 2613 4998
rect 2542 4967 2576 4978
rect 2579 4967 2588 4983
rect 2604 4967 2613 4983
rect 2620 4978 2630 4998
rect 2640 4978 2654 4998
rect 2655 4985 2666 4998
rect 2620 4967 2654 4978
rect 2655 4967 2666 4983
rect 2712 4974 2728 4990
rect 2735 4988 2765 5040
rect 2799 5036 2800 5043
rect 2784 5028 2800 5036
rect 2771 4996 2784 5015
rect 2799 4996 2829 5012
rect 2771 4980 2845 4996
rect 2771 4978 2784 4980
rect 2799 4978 2833 4980
rect 2436 4956 2449 4958
rect 2464 4956 2498 4958
rect 2436 4940 2498 4956
rect 2542 4951 2558 4954
rect 2620 4951 2650 4962
rect 2698 4958 2744 4974
rect 2771 4962 2845 4978
rect 2698 4956 2732 4958
rect 2697 4940 2744 4956
rect 2771 4940 2784 4962
rect 2799 4940 2829 4962
rect 2856 4940 2857 4956
rect 2872 4940 2885 5100
rect 2915 4996 2928 5100
rect 2973 5078 2974 5088
rect 2989 5078 3002 5088
rect 2973 5074 3002 5078
rect 3007 5074 3037 5100
rect 3055 5086 3071 5088
rect 3143 5086 3196 5100
rect 3144 5084 3208 5086
rect 3251 5084 3266 5100
rect 3315 5097 3345 5100
rect 3315 5094 3351 5097
rect 3281 5086 3297 5088
rect 3055 5074 3070 5078
rect 2973 5072 3070 5074
rect 3098 5072 3266 5084
rect 3282 5074 3297 5078
rect 3315 5075 3354 5094
rect 3373 5088 3380 5089
rect 3379 5081 3380 5088
rect 3363 5078 3364 5081
rect 3379 5078 3392 5081
rect 3315 5074 3345 5075
rect 3354 5074 3360 5075
rect 3363 5074 3392 5078
rect 3282 5073 3392 5074
rect 3282 5072 3398 5073
rect 2957 5064 3008 5072
rect 2957 5052 2982 5064
rect 2989 5052 3008 5064
rect 3039 5064 3089 5072
rect 3039 5056 3055 5064
rect 3062 5062 3089 5064
rect 3098 5062 3319 5072
rect 3062 5052 3319 5062
rect 3348 5064 3398 5072
rect 3348 5055 3364 5064
rect 2957 5044 3008 5052
rect 3055 5044 3319 5052
rect 3345 5052 3364 5055
rect 3371 5052 3398 5064
rect 3345 5044 3398 5052
rect 2973 5036 2974 5044
rect 2989 5036 3002 5044
rect 2973 5028 2989 5036
rect 2970 5021 2989 5024
rect 2970 5012 2992 5021
rect 2943 5002 2992 5012
rect 2943 4996 2973 5002
rect 2992 4997 2997 5002
rect 2915 4980 2989 4996
rect 3007 4988 3037 5044
rect 3072 5034 3280 5044
rect 3315 5040 3360 5044
rect 3363 5043 3364 5044
rect 3379 5043 3392 5044
rect 3098 5004 3287 5034
rect 3113 5001 3287 5004
rect 3106 4998 3287 5001
rect 2915 4978 2928 4980
rect 2943 4978 2977 4980
rect 2915 4962 2989 4978
rect 3016 4974 3029 4988
rect 3044 4974 3060 4990
rect 3106 4985 3117 4998
rect 2899 4940 2900 4956
rect 2915 4940 2928 4962
rect 2943 4940 2973 4962
rect 3016 4958 3078 4974
rect 3106 4967 3117 4983
rect 3122 4978 3132 4998
rect 3142 4978 3156 4998
rect 3159 4985 3168 4998
rect 3184 4985 3193 4998
rect 3122 4967 3156 4978
rect 3159 4967 3168 4983
rect 3184 4967 3193 4983
rect 3200 4978 3210 4998
rect 3220 4978 3234 4998
rect 3235 4985 3246 4998
rect 3200 4967 3234 4978
rect 3235 4967 3246 4983
rect 3292 4974 3308 4990
rect 3315 4988 3345 5040
rect 3379 5036 3380 5043
rect 3364 5028 3380 5036
rect 3351 4996 3364 5015
rect 3379 4996 3409 5012
rect 3351 4980 3425 4996
rect 3351 4978 3364 4980
rect 3379 4978 3413 4980
rect 3016 4956 3029 4958
rect 3044 4956 3078 4958
rect 3016 4940 3078 4956
rect 3122 4951 3138 4954
rect 3200 4951 3230 4962
rect 3278 4958 3324 4974
rect 3351 4962 3425 4978
rect 3278 4956 3312 4958
rect 3277 4940 3324 4956
rect 3351 4940 3364 4962
rect 3379 4940 3409 4962
rect 3436 4940 3437 4956
rect 3452 4940 3465 5100
rect 3495 4996 3508 5100
rect 3553 5078 3554 5088
rect 3569 5078 3582 5088
rect 3553 5074 3582 5078
rect 3587 5074 3617 5100
rect 3635 5086 3651 5088
rect 3723 5086 3776 5100
rect 3724 5084 3788 5086
rect 3831 5084 3846 5100
rect 3895 5097 3925 5100
rect 3895 5094 3931 5097
rect 3861 5086 3877 5088
rect 3635 5074 3650 5078
rect 3553 5072 3650 5074
rect 3678 5072 3846 5084
rect 3862 5074 3877 5078
rect 3895 5075 3934 5094
rect 3953 5088 3960 5089
rect 3959 5081 3960 5088
rect 3943 5078 3944 5081
rect 3959 5078 3972 5081
rect 3895 5074 3925 5075
rect 3934 5074 3940 5075
rect 3943 5074 3972 5078
rect 3862 5073 3972 5074
rect 3862 5072 3978 5073
rect 3537 5064 3588 5072
rect 3537 5052 3562 5064
rect 3569 5052 3588 5064
rect 3619 5064 3669 5072
rect 3619 5056 3635 5064
rect 3642 5062 3669 5064
rect 3678 5062 3899 5072
rect 3642 5052 3899 5062
rect 3928 5064 3978 5072
rect 3928 5055 3944 5064
rect 3537 5044 3588 5052
rect 3635 5044 3899 5052
rect 3925 5052 3944 5055
rect 3951 5052 3978 5064
rect 3925 5044 3978 5052
rect 3553 5036 3554 5044
rect 3569 5036 3582 5044
rect 3553 5028 3569 5036
rect 3550 5021 3569 5024
rect 3550 5012 3572 5021
rect 3523 5002 3572 5012
rect 3523 4996 3553 5002
rect 3572 4997 3577 5002
rect 3495 4980 3569 4996
rect 3587 4988 3617 5044
rect 3652 5034 3860 5044
rect 3895 5040 3940 5044
rect 3943 5043 3944 5044
rect 3959 5043 3972 5044
rect 3678 5004 3867 5034
rect 3693 5001 3867 5004
rect 3686 4998 3867 5001
rect 3495 4978 3508 4980
rect 3523 4978 3557 4980
rect 3495 4962 3569 4978
rect 3596 4974 3609 4988
rect 3624 4974 3640 4990
rect 3686 4985 3697 4998
rect 3479 4940 3480 4956
rect 3495 4940 3508 4962
rect 3523 4940 3553 4962
rect 3596 4958 3658 4974
rect 3686 4967 3697 4983
rect 3702 4978 3712 4998
rect 3722 4978 3736 4998
rect 3739 4985 3748 4998
rect 3764 4985 3773 4998
rect 3702 4967 3736 4978
rect 3739 4967 3748 4983
rect 3764 4967 3773 4983
rect 3780 4978 3790 4998
rect 3800 4978 3814 4998
rect 3815 4985 3826 4998
rect 3780 4967 3814 4978
rect 3815 4967 3826 4983
rect 3872 4974 3888 4990
rect 3895 4988 3925 5040
rect 3959 5036 3960 5043
rect 3944 5028 3960 5036
rect 3931 4996 3944 5015
rect 3959 4996 3989 5012
rect 3931 4980 4005 4996
rect 3931 4978 3944 4980
rect 3959 4978 3993 4980
rect 3596 4956 3609 4958
rect 3624 4956 3658 4958
rect 3596 4940 3658 4956
rect 3702 4951 3718 4954
rect 3780 4951 3810 4962
rect 3858 4958 3904 4974
rect 3931 4962 4005 4978
rect 3858 4956 3892 4958
rect 3857 4940 3904 4956
rect 3931 4940 3944 4962
rect 3959 4940 3989 4962
rect 4016 4940 4017 4956
rect 4032 4940 4045 5100
rect 4075 4996 4088 5100
rect 4133 5078 4134 5088
rect 4149 5078 4162 5088
rect 4133 5074 4162 5078
rect 4167 5074 4197 5100
rect 4215 5086 4231 5088
rect 4303 5086 4356 5100
rect 4304 5084 4368 5086
rect 4411 5084 4426 5100
rect 4475 5097 4505 5100
rect 4475 5094 4511 5097
rect 4441 5086 4457 5088
rect 4215 5074 4230 5078
rect 4133 5072 4230 5074
rect 4258 5072 4426 5084
rect 4442 5074 4457 5078
rect 4475 5075 4514 5094
rect 4533 5088 4540 5089
rect 4539 5081 4540 5088
rect 4523 5078 4524 5081
rect 4539 5078 4552 5081
rect 4475 5074 4505 5075
rect 4514 5074 4520 5075
rect 4523 5074 4552 5078
rect 4442 5073 4552 5074
rect 4442 5072 4558 5073
rect 4117 5064 4168 5072
rect 4117 5052 4142 5064
rect 4149 5052 4168 5064
rect 4199 5064 4249 5072
rect 4199 5056 4215 5064
rect 4222 5062 4249 5064
rect 4258 5062 4479 5072
rect 4222 5052 4479 5062
rect 4508 5064 4558 5072
rect 4508 5055 4524 5064
rect 4117 5044 4168 5052
rect 4215 5044 4479 5052
rect 4505 5052 4524 5055
rect 4531 5052 4558 5064
rect 4505 5044 4558 5052
rect 4133 5036 4134 5044
rect 4149 5036 4162 5044
rect 4133 5028 4149 5036
rect 4130 5021 4149 5024
rect 4130 5012 4152 5021
rect 4103 5002 4152 5012
rect 4103 4996 4133 5002
rect 4152 4997 4157 5002
rect 4075 4980 4149 4996
rect 4167 4988 4197 5044
rect 4232 5034 4440 5044
rect 4475 5040 4520 5044
rect 4523 5043 4524 5044
rect 4539 5043 4552 5044
rect 4258 5004 4447 5034
rect 4273 5001 4447 5004
rect 4266 4998 4447 5001
rect 4075 4978 4088 4980
rect 4103 4978 4137 4980
rect 4075 4962 4149 4978
rect 4176 4974 4189 4988
rect 4204 4974 4220 4990
rect 4266 4985 4277 4998
rect 4059 4940 4060 4956
rect 4075 4940 4088 4962
rect 4103 4940 4133 4962
rect 4176 4958 4238 4974
rect 4266 4967 4277 4983
rect 4282 4978 4292 4998
rect 4302 4978 4316 4998
rect 4319 4985 4328 4998
rect 4344 4985 4353 4998
rect 4282 4967 4316 4978
rect 4319 4967 4328 4983
rect 4344 4967 4353 4983
rect 4360 4978 4370 4998
rect 4380 4978 4394 4998
rect 4395 4985 4406 4998
rect 4360 4967 4394 4978
rect 4395 4967 4406 4983
rect 4452 4974 4468 4990
rect 4475 4988 4505 5040
rect 4539 5036 4540 5043
rect 4524 5028 4540 5036
rect 4511 4996 4524 5015
rect 4539 4996 4569 5012
rect 4511 4980 4585 4996
rect 4511 4978 4524 4980
rect 4539 4978 4573 4980
rect 4176 4956 4189 4958
rect 4204 4956 4238 4958
rect 4176 4940 4238 4956
rect 4282 4951 4298 4954
rect 4360 4951 4390 4962
rect 4438 4958 4484 4974
rect 4511 4962 4585 4978
rect 4438 4956 4472 4958
rect 4437 4940 4484 4956
rect 4511 4940 4524 4962
rect 4539 4940 4569 4962
rect 4596 4940 4597 4956
rect 4612 4940 4625 5100
rect 4655 4996 4668 5100
rect 4713 5078 4714 5088
rect 4729 5078 4742 5088
rect 4713 5074 4742 5078
rect 4747 5074 4777 5100
rect 4795 5086 4811 5088
rect 4883 5086 4936 5100
rect 4884 5084 4948 5086
rect 4991 5084 5006 5100
rect 5055 5097 5085 5100
rect 5055 5094 5091 5097
rect 5021 5086 5037 5088
rect 4795 5074 4810 5078
rect 4713 5072 4810 5074
rect 4838 5072 5006 5084
rect 5022 5074 5037 5078
rect 5055 5075 5094 5094
rect 5113 5088 5120 5089
rect 5119 5081 5120 5088
rect 5103 5078 5104 5081
rect 5119 5078 5132 5081
rect 5055 5074 5085 5075
rect 5094 5074 5100 5075
rect 5103 5074 5132 5078
rect 5022 5073 5132 5074
rect 5022 5072 5138 5073
rect 4697 5064 4748 5072
rect 4697 5052 4722 5064
rect 4729 5052 4748 5064
rect 4779 5064 4829 5072
rect 4779 5056 4795 5064
rect 4802 5062 4829 5064
rect 4838 5062 5059 5072
rect 4802 5052 5059 5062
rect 5088 5064 5138 5072
rect 5088 5055 5104 5064
rect 4697 5044 4748 5052
rect 4795 5044 5059 5052
rect 5085 5052 5104 5055
rect 5111 5052 5138 5064
rect 5085 5044 5138 5052
rect 4713 5036 4714 5044
rect 4729 5036 4742 5044
rect 4713 5028 4729 5036
rect 4710 5021 4729 5024
rect 4710 5012 4732 5021
rect 4683 5002 4732 5012
rect 4683 4996 4713 5002
rect 4732 4997 4737 5002
rect 4655 4980 4729 4996
rect 4747 4988 4777 5044
rect 4812 5034 5020 5044
rect 5055 5040 5100 5044
rect 5103 5043 5104 5044
rect 5119 5043 5132 5044
rect 4838 5004 5027 5034
rect 4853 5001 5027 5004
rect 4846 4998 5027 5001
rect 4655 4978 4668 4980
rect 4683 4978 4717 4980
rect 4655 4962 4729 4978
rect 4756 4974 4769 4988
rect 4784 4974 4800 4990
rect 4846 4985 4857 4998
rect 4639 4940 4640 4956
rect 4655 4940 4668 4962
rect 4683 4940 4713 4962
rect 4756 4958 4818 4974
rect 4846 4967 4857 4983
rect 4862 4978 4872 4998
rect 4882 4978 4896 4998
rect 4899 4985 4908 4998
rect 4924 4985 4933 4998
rect 4862 4967 4896 4978
rect 4899 4967 4908 4983
rect 4924 4967 4933 4983
rect 4940 4978 4950 4998
rect 4960 4978 4974 4998
rect 4975 4985 4986 4998
rect 4940 4967 4974 4978
rect 4975 4967 4986 4983
rect 5032 4974 5048 4990
rect 5055 4988 5085 5040
rect 5119 5036 5120 5043
rect 5104 5028 5120 5036
rect 5091 4996 5104 5015
rect 5119 4996 5149 5012
rect 5091 4980 5165 4996
rect 5091 4978 5104 4980
rect 5119 4978 5153 4980
rect 4756 4956 4769 4958
rect 4784 4956 4818 4958
rect 4756 4940 4818 4956
rect 4862 4951 4878 4954
rect 4940 4951 4970 4962
rect 5018 4958 5064 4974
rect 5091 4962 5165 4978
rect 5018 4956 5052 4958
rect 5017 4940 5064 4956
rect 5091 4940 5104 4962
rect 5119 4940 5149 4962
rect 5176 4940 5177 4956
rect 5192 4940 5205 5100
rect 5235 4996 5248 5100
rect 5293 5078 5294 5088
rect 5309 5078 5322 5088
rect 5293 5074 5322 5078
rect 5327 5074 5357 5100
rect 5375 5086 5391 5088
rect 5463 5086 5516 5100
rect 5464 5084 5528 5086
rect 5571 5084 5586 5100
rect 5635 5097 5665 5100
rect 5635 5094 5671 5097
rect 5601 5086 5617 5088
rect 5375 5074 5390 5078
rect 5293 5072 5390 5074
rect 5418 5072 5586 5084
rect 5602 5074 5617 5078
rect 5635 5075 5674 5094
rect 5693 5088 5700 5089
rect 5699 5081 5700 5088
rect 5683 5078 5684 5081
rect 5699 5078 5712 5081
rect 5635 5074 5665 5075
rect 5674 5074 5680 5075
rect 5683 5074 5712 5078
rect 5602 5073 5712 5074
rect 5602 5072 5718 5073
rect 5277 5064 5328 5072
rect 5277 5052 5302 5064
rect 5309 5052 5328 5064
rect 5359 5064 5409 5072
rect 5359 5056 5375 5064
rect 5382 5062 5409 5064
rect 5418 5062 5639 5072
rect 5382 5052 5639 5062
rect 5668 5064 5718 5072
rect 5668 5055 5684 5064
rect 5277 5044 5328 5052
rect 5375 5044 5639 5052
rect 5665 5052 5684 5055
rect 5691 5052 5718 5064
rect 5665 5044 5718 5052
rect 5293 5036 5294 5044
rect 5309 5036 5322 5044
rect 5293 5028 5309 5036
rect 5290 5021 5309 5024
rect 5290 5012 5312 5021
rect 5263 5002 5312 5012
rect 5263 4996 5293 5002
rect 5312 4997 5317 5002
rect 5235 4980 5309 4996
rect 5327 4988 5357 5044
rect 5392 5034 5600 5044
rect 5635 5040 5680 5044
rect 5683 5043 5684 5044
rect 5699 5043 5712 5044
rect 5418 5004 5607 5034
rect 5433 5001 5607 5004
rect 5426 4998 5607 5001
rect 5235 4978 5248 4980
rect 5263 4978 5297 4980
rect 5235 4962 5309 4978
rect 5336 4974 5349 4988
rect 5364 4974 5380 4990
rect 5426 4985 5437 4998
rect 5219 4940 5220 4956
rect 5235 4940 5248 4962
rect 5263 4940 5293 4962
rect 5336 4958 5398 4974
rect 5426 4967 5437 4983
rect 5442 4978 5452 4998
rect 5462 4978 5476 4998
rect 5479 4985 5488 4998
rect 5504 4985 5513 4998
rect 5442 4967 5476 4978
rect 5479 4967 5488 4983
rect 5504 4967 5513 4983
rect 5520 4978 5530 4998
rect 5540 4978 5554 4998
rect 5555 4985 5566 4998
rect 5520 4967 5554 4978
rect 5555 4967 5566 4983
rect 5612 4974 5628 4990
rect 5635 4988 5665 5040
rect 5699 5036 5700 5043
rect 5684 5028 5700 5036
rect 5671 4996 5684 5015
rect 5699 4996 5729 5012
rect 5671 4980 5745 4996
rect 5671 4978 5684 4980
rect 5699 4978 5733 4980
rect 5336 4956 5349 4958
rect 5364 4956 5398 4958
rect 5336 4940 5398 4956
rect 5442 4951 5458 4954
rect 5520 4951 5550 4962
rect 5598 4958 5644 4974
rect 5671 4962 5745 4978
rect 5598 4956 5632 4958
rect 5597 4940 5644 4956
rect 5671 4940 5684 4962
rect 5699 4940 5729 4962
rect 5756 4940 5757 4956
rect 5772 4940 5785 5100
rect 5815 4996 5828 5100
rect 5873 5078 5874 5088
rect 5889 5078 5902 5088
rect 5873 5074 5902 5078
rect 5907 5074 5937 5100
rect 5955 5086 5971 5088
rect 6043 5086 6096 5100
rect 6044 5084 6108 5086
rect 6151 5084 6166 5100
rect 6215 5097 6245 5100
rect 6215 5094 6251 5097
rect 6181 5086 6197 5088
rect 5955 5074 5970 5078
rect 5873 5072 5970 5074
rect 5998 5072 6166 5084
rect 6182 5074 6197 5078
rect 6215 5075 6254 5094
rect 6273 5088 6280 5089
rect 6279 5081 6280 5088
rect 6263 5078 6264 5081
rect 6279 5078 6292 5081
rect 6215 5074 6245 5075
rect 6254 5074 6260 5075
rect 6263 5074 6292 5078
rect 6182 5073 6292 5074
rect 6182 5072 6298 5073
rect 5857 5064 5908 5072
rect 5857 5052 5882 5064
rect 5889 5052 5908 5064
rect 5939 5064 5989 5072
rect 5939 5056 5955 5064
rect 5962 5062 5989 5064
rect 5998 5062 6219 5072
rect 5962 5052 6219 5062
rect 6248 5064 6298 5072
rect 6248 5055 6264 5064
rect 5857 5044 5908 5052
rect 5955 5044 6219 5052
rect 6245 5052 6264 5055
rect 6271 5052 6298 5064
rect 6245 5044 6298 5052
rect 5873 5036 5874 5044
rect 5889 5036 5902 5044
rect 5873 5028 5889 5036
rect 5870 5021 5889 5024
rect 5870 5012 5892 5021
rect 5843 5002 5892 5012
rect 5843 4996 5873 5002
rect 5892 4997 5897 5002
rect 5815 4980 5889 4996
rect 5907 4988 5937 5044
rect 5972 5034 6180 5044
rect 6215 5040 6260 5044
rect 6263 5043 6264 5044
rect 6279 5043 6292 5044
rect 5998 5004 6187 5034
rect 6013 5001 6187 5004
rect 6006 4998 6187 5001
rect 5815 4978 5828 4980
rect 5843 4978 5877 4980
rect 5815 4962 5889 4978
rect 5916 4974 5929 4988
rect 5944 4974 5960 4990
rect 6006 4985 6017 4998
rect 5799 4940 5800 4956
rect 5815 4940 5828 4962
rect 5843 4940 5873 4962
rect 5916 4958 5978 4974
rect 6006 4967 6017 4983
rect 6022 4978 6032 4998
rect 6042 4978 6056 4998
rect 6059 4985 6068 4998
rect 6084 4985 6093 4998
rect 6022 4967 6056 4978
rect 6059 4967 6068 4983
rect 6084 4967 6093 4983
rect 6100 4978 6110 4998
rect 6120 4978 6134 4998
rect 6135 4985 6146 4998
rect 6100 4967 6134 4978
rect 6135 4967 6146 4983
rect 6192 4974 6208 4990
rect 6215 4988 6245 5040
rect 6279 5036 6280 5043
rect 6264 5028 6280 5036
rect 6251 4996 6264 5015
rect 6279 4996 6309 5012
rect 6251 4980 6325 4996
rect 6251 4978 6264 4980
rect 6279 4978 6313 4980
rect 5916 4956 5929 4958
rect 5944 4956 5978 4958
rect 5916 4940 5978 4956
rect 6022 4951 6038 4954
rect 6100 4951 6130 4962
rect 6178 4958 6224 4974
rect 6251 4962 6325 4978
rect 6178 4956 6212 4958
rect 6177 4940 6224 4956
rect 6251 4940 6264 4962
rect 6279 4940 6309 4962
rect 6336 4940 6337 4956
rect 6352 4940 6365 5100
rect 6395 4996 6408 5100
rect 6453 5078 6454 5088
rect 6469 5078 6482 5088
rect 6453 5074 6482 5078
rect 6487 5074 6517 5100
rect 6535 5086 6551 5088
rect 6623 5086 6676 5100
rect 6624 5084 6688 5086
rect 6731 5084 6746 5100
rect 6795 5097 6825 5100
rect 6795 5094 6831 5097
rect 6761 5086 6777 5088
rect 6535 5074 6550 5078
rect 6453 5072 6550 5074
rect 6578 5072 6746 5084
rect 6762 5074 6777 5078
rect 6795 5075 6834 5094
rect 6853 5088 6860 5089
rect 6859 5081 6860 5088
rect 6843 5078 6844 5081
rect 6859 5078 6872 5081
rect 6795 5074 6825 5075
rect 6834 5074 6840 5075
rect 6843 5074 6872 5078
rect 6762 5073 6872 5074
rect 6762 5072 6878 5073
rect 6437 5064 6488 5072
rect 6437 5052 6462 5064
rect 6469 5052 6488 5064
rect 6519 5064 6569 5072
rect 6519 5056 6535 5064
rect 6542 5062 6569 5064
rect 6578 5062 6799 5072
rect 6542 5052 6799 5062
rect 6828 5064 6878 5072
rect 6828 5055 6844 5064
rect 6437 5044 6488 5052
rect 6535 5044 6799 5052
rect 6825 5052 6844 5055
rect 6851 5052 6878 5064
rect 6825 5044 6878 5052
rect 6453 5036 6454 5044
rect 6469 5036 6482 5044
rect 6453 5028 6469 5036
rect 6450 5021 6469 5024
rect 6450 5012 6472 5021
rect 6423 5002 6472 5012
rect 6423 4996 6453 5002
rect 6472 4997 6477 5002
rect 6395 4980 6469 4996
rect 6487 4988 6517 5044
rect 6552 5034 6760 5044
rect 6795 5040 6840 5044
rect 6843 5043 6844 5044
rect 6859 5043 6872 5044
rect 6578 5004 6767 5034
rect 6593 5001 6767 5004
rect 6586 4998 6767 5001
rect 6395 4978 6408 4980
rect 6423 4978 6457 4980
rect 6395 4962 6469 4978
rect 6496 4974 6509 4988
rect 6524 4974 6540 4990
rect 6586 4985 6597 4998
rect 6379 4940 6380 4956
rect 6395 4940 6408 4962
rect 6423 4940 6453 4962
rect 6496 4958 6558 4974
rect 6586 4967 6597 4983
rect 6602 4978 6612 4998
rect 6622 4978 6636 4998
rect 6639 4985 6648 4998
rect 6664 4985 6673 4998
rect 6602 4967 6636 4978
rect 6639 4967 6648 4983
rect 6664 4967 6673 4983
rect 6680 4978 6690 4998
rect 6700 4978 6714 4998
rect 6715 4985 6726 4998
rect 6680 4967 6714 4978
rect 6715 4967 6726 4983
rect 6772 4974 6788 4990
rect 6795 4988 6825 5040
rect 6859 5036 6860 5043
rect 6844 5028 6860 5036
rect 6831 4996 6844 5015
rect 6859 4996 6889 5012
rect 6831 4980 6905 4996
rect 6831 4978 6844 4980
rect 6859 4978 6893 4980
rect 6496 4956 6509 4958
rect 6524 4956 6558 4958
rect 6496 4940 6558 4956
rect 6602 4951 6618 4954
rect 6680 4951 6710 4962
rect 6758 4958 6804 4974
rect 6831 4962 6905 4978
rect 6758 4956 6792 4958
rect 6757 4940 6804 4956
rect 6831 4940 6844 4962
rect 6859 4940 6889 4962
rect 6916 4940 6917 4956
rect 6932 4940 6945 5100
rect 6975 4996 6988 5100
rect 7033 5078 7034 5088
rect 7049 5078 7062 5088
rect 7033 5074 7062 5078
rect 7067 5074 7097 5100
rect 7115 5086 7131 5088
rect 7203 5086 7256 5100
rect 7204 5084 7268 5086
rect 7311 5084 7326 5100
rect 7375 5097 7405 5100
rect 7375 5094 7411 5097
rect 7341 5086 7357 5088
rect 7115 5074 7130 5078
rect 7033 5072 7130 5074
rect 7158 5072 7326 5084
rect 7342 5074 7357 5078
rect 7375 5075 7414 5094
rect 7433 5088 7440 5089
rect 7439 5081 7440 5088
rect 7423 5078 7424 5081
rect 7439 5078 7452 5081
rect 7375 5074 7405 5075
rect 7414 5074 7420 5075
rect 7423 5074 7452 5078
rect 7342 5073 7452 5074
rect 7342 5072 7458 5073
rect 7017 5064 7068 5072
rect 7017 5052 7042 5064
rect 7049 5052 7068 5064
rect 7099 5064 7149 5072
rect 7099 5056 7115 5064
rect 7122 5062 7149 5064
rect 7158 5062 7379 5072
rect 7122 5052 7379 5062
rect 7408 5064 7458 5072
rect 7408 5055 7424 5064
rect 7017 5044 7068 5052
rect 7115 5044 7379 5052
rect 7405 5052 7424 5055
rect 7431 5052 7458 5064
rect 7405 5044 7458 5052
rect 7033 5036 7034 5044
rect 7049 5036 7062 5044
rect 7033 5028 7049 5036
rect 7030 5021 7049 5024
rect 7030 5012 7052 5021
rect 7003 5002 7052 5012
rect 7003 4996 7033 5002
rect 7052 4997 7057 5002
rect 6975 4980 7049 4996
rect 7067 4988 7097 5044
rect 7132 5034 7340 5044
rect 7375 5040 7420 5044
rect 7423 5043 7424 5044
rect 7439 5043 7452 5044
rect 7158 5004 7347 5034
rect 7173 5001 7347 5004
rect 7166 4998 7347 5001
rect 6975 4978 6988 4980
rect 7003 4978 7037 4980
rect 6975 4962 7049 4978
rect 7076 4974 7089 4988
rect 7104 4974 7120 4990
rect 7166 4985 7177 4998
rect 6959 4940 6960 4956
rect 6975 4940 6988 4962
rect 7003 4940 7033 4962
rect 7076 4958 7138 4974
rect 7166 4967 7177 4983
rect 7182 4978 7192 4998
rect 7202 4978 7216 4998
rect 7219 4985 7228 4998
rect 7244 4985 7253 4998
rect 7182 4967 7216 4978
rect 7219 4967 7228 4983
rect 7244 4967 7253 4983
rect 7260 4978 7270 4998
rect 7280 4978 7294 4998
rect 7295 4985 7306 4998
rect 7260 4967 7294 4978
rect 7295 4967 7306 4983
rect 7352 4974 7368 4990
rect 7375 4988 7405 5040
rect 7439 5036 7440 5043
rect 7424 5028 7440 5036
rect 7411 4996 7424 5015
rect 7439 4996 7469 5012
rect 7411 4980 7485 4996
rect 7411 4978 7424 4980
rect 7439 4978 7473 4980
rect 7076 4956 7089 4958
rect 7104 4956 7138 4958
rect 7076 4940 7138 4956
rect 7182 4951 7198 4954
rect 7260 4951 7290 4962
rect 7338 4958 7384 4974
rect 7411 4962 7485 4978
rect 7338 4956 7372 4958
rect 7337 4940 7384 4956
rect 7411 4940 7424 4962
rect 7439 4940 7469 4962
rect 7496 4940 7497 4956
rect 7512 4940 7525 5100
rect 7555 4996 7568 5100
rect 7613 5078 7614 5088
rect 7629 5078 7642 5088
rect 7613 5074 7642 5078
rect 7647 5074 7677 5100
rect 7695 5086 7711 5088
rect 7783 5086 7836 5100
rect 7784 5084 7848 5086
rect 7891 5084 7906 5100
rect 7955 5097 7985 5100
rect 7955 5094 7991 5097
rect 7921 5086 7937 5088
rect 7695 5074 7710 5078
rect 7613 5072 7710 5074
rect 7738 5072 7906 5084
rect 7922 5074 7937 5078
rect 7955 5075 7994 5094
rect 8013 5088 8020 5089
rect 8019 5081 8020 5088
rect 8003 5078 8004 5081
rect 8019 5078 8032 5081
rect 7955 5074 7985 5075
rect 7994 5074 8000 5075
rect 8003 5074 8032 5078
rect 7922 5073 8032 5074
rect 7922 5072 8038 5073
rect 7597 5064 7648 5072
rect 7597 5052 7622 5064
rect 7629 5052 7648 5064
rect 7679 5064 7729 5072
rect 7679 5056 7695 5064
rect 7702 5062 7729 5064
rect 7738 5062 7959 5072
rect 7702 5052 7959 5062
rect 7988 5064 8038 5072
rect 7988 5055 8004 5064
rect 7597 5044 7648 5052
rect 7695 5044 7959 5052
rect 7985 5052 8004 5055
rect 8011 5052 8038 5064
rect 7985 5044 8038 5052
rect 7613 5036 7614 5044
rect 7629 5036 7642 5044
rect 7613 5028 7629 5036
rect 7610 5021 7629 5024
rect 7610 5012 7632 5021
rect 7583 5002 7632 5012
rect 7583 4996 7613 5002
rect 7632 4997 7637 5002
rect 7555 4980 7629 4996
rect 7647 4988 7677 5044
rect 7712 5034 7920 5044
rect 7955 5040 8000 5044
rect 8003 5043 8004 5044
rect 8019 5043 8032 5044
rect 7738 5004 7927 5034
rect 7753 5001 7927 5004
rect 7746 4998 7927 5001
rect 7555 4978 7568 4980
rect 7583 4978 7617 4980
rect 7555 4962 7629 4978
rect 7656 4974 7669 4988
rect 7684 4974 7700 4990
rect 7746 4985 7757 4998
rect 7539 4940 7540 4956
rect 7555 4940 7568 4962
rect 7583 4940 7613 4962
rect 7656 4958 7718 4974
rect 7746 4967 7757 4983
rect 7762 4978 7772 4998
rect 7782 4978 7796 4998
rect 7799 4985 7808 4998
rect 7824 4985 7833 4998
rect 7762 4967 7796 4978
rect 7799 4967 7808 4983
rect 7824 4967 7833 4983
rect 7840 4978 7850 4998
rect 7860 4978 7874 4998
rect 7875 4985 7886 4998
rect 7840 4967 7874 4978
rect 7875 4967 7886 4983
rect 7932 4974 7948 4990
rect 7955 4988 7985 5040
rect 8019 5036 8020 5043
rect 8004 5028 8020 5036
rect 7991 4996 8004 5015
rect 8019 4996 8049 5012
rect 7991 4980 8065 4996
rect 7991 4978 8004 4980
rect 8019 4978 8053 4980
rect 7656 4956 7669 4958
rect 7684 4956 7718 4958
rect 7656 4940 7718 4956
rect 7762 4951 7778 4954
rect 7840 4951 7870 4962
rect 7918 4958 7964 4974
rect 7991 4962 8065 4978
rect 7918 4956 7952 4958
rect 7917 4940 7964 4956
rect 7991 4940 8004 4962
rect 8019 4940 8049 4962
rect 8076 4940 8077 4956
rect 8092 4940 8105 5100
rect 8135 4996 8148 5100
rect 8193 5078 8194 5088
rect 8209 5078 8222 5088
rect 8193 5074 8222 5078
rect 8227 5074 8257 5100
rect 8275 5086 8291 5088
rect 8363 5086 8416 5100
rect 8364 5084 8428 5086
rect 8471 5084 8486 5100
rect 8535 5097 8565 5100
rect 8535 5094 8571 5097
rect 8501 5086 8517 5088
rect 8275 5074 8290 5078
rect 8193 5072 8290 5074
rect 8318 5072 8486 5084
rect 8502 5074 8517 5078
rect 8535 5075 8574 5094
rect 8593 5088 8600 5089
rect 8599 5081 8600 5088
rect 8583 5078 8584 5081
rect 8599 5078 8612 5081
rect 8535 5074 8565 5075
rect 8574 5074 8580 5075
rect 8583 5074 8612 5078
rect 8502 5073 8612 5074
rect 8502 5072 8618 5073
rect 8177 5064 8228 5072
rect 8177 5052 8202 5064
rect 8209 5052 8228 5064
rect 8259 5064 8309 5072
rect 8259 5056 8275 5064
rect 8282 5062 8309 5064
rect 8318 5062 8539 5072
rect 8282 5052 8539 5062
rect 8568 5064 8618 5072
rect 8568 5055 8584 5064
rect 8177 5044 8228 5052
rect 8275 5044 8539 5052
rect 8565 5052 8584 5055
rect 8591 5052 8618 5064
rect 8565 5044 8618 5052
rect 8193 5036 8194 5044
rect 8209 5036 8222 5044
rect 8193 5028 8209 5036
rect 8190 5021 8209 5024
rect 8190 5012 8212 5021
rect 8163 5002 8212 5012
rect 8163 4996 8193 5002
rect 8212 4997 8217 5002
rect 8135 4980 8209 4996
rect 8227 4988 8257 5044
rect 8292 5034 8500 5044
rect 8535 5040 8580 5044
rect 8583 5043 8584 5044
rect 8599 5043 8612 5044
rect 8318 5004 8507 5034
rect 8333 5001 8507 5004
rect 8326 4998 8507 5001
rect 8135 4978 8148 4980
rect 8163 4978 8197 4980
rect 8135 4962 8209 4978
rect 8236 4974 8249 4988
rect 8264 4974 8280 4990
rect 8326 4985 8337 4998
rect 8119 4940 8120 4956
rect 8135 4940 8148 4962
rect 8163 4940 8193 4962
rect 8236 4958 8298 4974
rect 8326 4967 8337 4983
rect 8342 4978 8352 4998
rect 8362 4978 8376 4998
rect 8379 4985 8388 4998
rect 8404 4985 8413 4998
rect 8342 4967 8376 4978
rect 8379 4967 8388 4983
rect 8404 4967 8413 4983
rect 8420 4978 8430 4998
rect 8440 4978 8454 4998
rect 8455 4985 8466 4998
rect 8420 4967 8454 4978
rect 8455 4967 8466 4983
rect 8512 4974 8528 4990
rect 8535 4988 8565 5040
rect 8599 5036 8600 5043
rect 8584 5028 8600 5036
rect 8571 4996 8584 5015
rect 8599 4996 8629 5012
rect 8571 4980 8645 4996
rect 8571 4978 8584 4980
rect 8599 4978 8633 4980
rect 8236 4956 8249 4958
rect 8264 4956 8298 4958
rect 8236 4940 8298 4956
rect 8342 4951 8358 4954
rect 8420 4951 8450 4962
rect 8498 4958 8544 4974
rect 8571 4962 8645 4978
rect 8498 4956 8532 4958
rect 8497 4940 8544 4956
rect 8571 4940 8584 4962
rect 8599 4940 8629 4962
rect 8656 4940 8657 4956
rect 8672 4940 8685 5100
rect 8715 4996 8728 5100
rect 8773 5078 8774 5088
rect 8789 5078 8802 5088
rect 8773 5074 8802 5078
rect 8807 5074 8837 5100
rect 8855 5086 8871 5088
rect 8943 5086 8996 5100
rect 8944 5084 9008 5086
rect 9051 5084 9066 5100
rect 9115 5097 9145 5100
rect 9115 5094 9151 5097
rect 9081 5086 9097 5088
rect 8855 5074 8870 5078
rect 8773 5072 8870 5074
rect 8898 5072 9066 5084
rect 9082 5074 9097 5078
rect 9115 5075 9154 5094
rect 9173 5088 9180 5089
rect 9179 5081 9180 5088
rect 9163 5078 9164 5081
rect 9179 5078 9192 5081
rect 9115 5074 9145 5075
rect 9154 5074 9160 5075
rect 9163 5074 9192 5078
rect 9082 5073 9192 5074
rect 9082 5072 9198 5073
rect 8757 5064 8808 5072
rect 8757 5052 8782 5064
rect 8789 5052 8808 5064
rect 8839 5064 8889 5072
rect 8839 5056 8855 5064
rect 8862 5062 8889 5064
rect 8898 5062 9119 5072
rect 8862 5052 9119 5062
rect 9148 5064 9198 5072
rect 9148 5055 9164 5064
rect 8757 5044 8808 5052
rect 8855 5044 9119 5052
rect 9145 5052 9164 5055
rect 9171 5052 9198 5064
rect 9145 5044 9198 5052
rect 8773 5036 8774 5044
rect 8789 5036 8802 5044
rect 8773 5028 8789 5036
rect 8770 5021 8789 5024
rect 8770 5012 8792 5021
rect 8743 5002 8792 5012
rect 8743 4996 8773 5002
rect 8792 4997 8797 5002
rect 8715 4980 8789 4996
rect 8807 4988 8837 5044
rect 8872 5034 9080 5044
rect 9115 5040 9160 5044
rect 9163 5043 9164 5044
rect 9179 5043 9192 5044
rect 8898 5004 9087 5034
rect 8913 5001 9087 5004
rect 8906 4998 9087 5001
rect 8715 4978 8728 4980
rect 8743 4978 8777 4980
rect 8715 4962 8789 4978
rect 8816 4974 8829 4988
rect 8844 4974 8860 4990
rect 8906 4985 8917 4998
rect 8699 4940 8700 4956
rect 8715 4940 8728 4962
rect 8743 4940 8773 4962
rect 8816 4958 8878 4974
rect 8906 4967 8917 4983
rect 8922 4978 8932 4998
rect 8942 4978 8956 4998
rect 8959 4985 8968 4998
rect 8984 4985 8993 4998
rect 8922 4967 8956 4978
rect 8959 4967 8968 4983
rect 8984 4967 8993 4983
rect 9000 4978 9010 4998
rect 9020 4978 9034 4998
rect 9035 4985 9046 4998
rect 9000 4967 9034 4978
rect 9035 4967 9046 4983
rect 9092 4974 9108 4990
rect 9115 4988 9145 5040
rect 9179 5036 9180 5043
rect 9164 5028 9180 5036
rect 9151 4996 9164 5015
rect 9179 4996 9209 5012
rect 9151 4980 9225 4996
rect 9151 4978 9164 4980
rect 9179 4978 9213 4980
rect 8816 4956 8829 4958
rect 8844 4956 8878 4958
rect 8816 4940 8878 4956
rect 8922 4951 8938 4954
rect 9000 4951 9030 4962
rect 9078 4958 9124 4974
rect 9151 4962 9225 4978
rect 9078 4956 9112 4958
rect 9077 4940 9124 4956
rect 9151 4940 9164 4962
rect 9179 4940 9209 4962
rect 9236 4940 9237 4956
rect 9252 4940 9265 5100
rect -7 4932 34 4940
rect -7 4906 8 4932
rect 15 4906 34 4932
rect 98 4928 160 4940
rect 172 4928 247 4940
rect 305 4928 380 4940
rect 392 4928 423 4940
rect 429 4928 464 4940
rect 98 4926 260 4928
rect -7 4898 34 4906
rect 116 4902 129 4926
rect 144 4924 159 4926
rect -1 4888 0 4898
rect 15 4888 28 4898
rect 43 4888 73 4902
rect 116 4888 159 4902
rect 183 4899 190 4906
rect 193 4902 260 4926
rect 292 4926 464 4928
rect 262 4904 290 4908
rect 292 4904 372 4926
rect 393 4924 408 4926
rect 262 4902 372 4904
rect 193 4898 372 4902
rect 166 4888 196 4898
rect 198 4888 351 4898
rect 359 4888 389 4898
rect 393 4888 423 4902
rect 451 4888 464 4926
rect 536 4932 571 4940
rect 536 4906 537 4932
rect 544 4906 571 4932
rect 479 4888 509 4902
rect 536 4898 571 4906
rect 573 4932 614 4940
rect 573 4906 588 4932
rect 595 4906 614 4932
rect 678 4928 740 4940
rect 752 4928 827 4940
rect 885 4928 960 4940
rect 972 4928 1003 4940
rect 1009 4928 1044 4940
rect 678 4926 840 4928
rect 573 4898 614 4906
rect 696 4902 709 4926
rect 724 4924 739 4926
rect 536 4888 537 4898
rect 552 4888 565 4898
rect 579 4888 580 4898
rect 595 4888 608 4898
rect 623 4888 653 4902
rect 696 4888 739 4902
rect 763 4899 770 4906
rect 773 4902 840 4926
rect 872 4926 1044 4928
rect 842 4904 870 4908
rect 872 4904 952 4926
rect 973 4924 988 4926
rect 842 4902 952 4904
rect 773 4898 952 4902
rect 746 4888 776 4898
rect 778 4888 931 4898
rect 939 4888 969 4898
rect 973 4888 1003 4902
rect 1031 4888 1044 4926
rect 1116 4932 1151 4940
rect 1116 4906 1117 4932
rect 1124 4906 1151 4932
rect 1059 4888 1089 4902
rect 1116 4898 1151 4906
rect 1153 4932 1194 4940
rect 1153 4906 1168 4932
rect 1175 4906 1194 4932
rect 1258 4928 1320 4940
rect 1332 4928 1407 4940
rect 1465 4928 1540 4940
rect 1552 4928 1583 4940
rect 1589 4928 1624 4940
rect 1258 4926 1420 4928
rect 1153 4898 1194 4906
rect 1276 4902 1289 4926
rect 1304 4924 1319 4926
rect 1116 4888 1117 4898
rect 1132 4888 1145 4898
rect 1159 4888 1160 4898
rect 1175 4888 1188 4898
rect 1203 4888 1233 4902
rect 1276 4888 1319 4902
rect 1343 4899 1350 4906
rect 1353 4902 1420 4926
rect 1452 4926 1624 4928
rect 1422 4904 1450 4908
rect 1452 4904 1532 4926
rect 1553 4924 1568 4926
rect 1422 4902 1532 4904
rect 1353 4898 1532 4902
rect 1326 4888 1356 4898
rect 1358 4888 1511 4898
rect 1519 4888 1549 4898
rect 1553 4888 1583 4902
rect 1611 4888 1624 4926
rect 1696 4932 1731 4940
rect 1696 4906 1697 4932
rect 1704 4906 1731 4932
rect 1639 4888 1669 4902
rect 1696 4898 1731 4906
rect 1733 4932 1774 4940
rect 1733 4906 1748 4932
rect 1755 4906 1774 4932
rect 1838 4928 1900 4940
rect 1912 4928 1987 4940
rect 2045 4928 2120 4940
rect 2132 4928 2163 4940
rect 2169 4928 2204 4940
rect 1838 4926 2000 4928
rect 1733 4898 1774 4906
rect 1856 4902 1869 4926
rect 1884 4924 1899 4926
rect 1696 4888 1697 4898
rect 1712 4888 1725 4898
rect 1739 4888 1740 4898
rect 1755 4888 1768 4898
rect 1783 4888 1813 4902
rect 1856 4888 1899 4902
rect 1923 4899 1930 4906
rect 1933 4902 2000 4926
rect 2032 4926 2204 4928
rect 2002 4904 2030 4908
rect 2032 4904 2112 4926
rect 2133 4924 2148 4926
rect 2002 4902 2112 4904
rect 1933 4898 2112 4902
rect 1906 4888 1936 4898
rect 1938 4888 2091 4898
rect 2099 4888 2129 4898
rect 2133 4888 2163 4902
rect 2191 4888 2204 4926
rect 2276 4932 2311 4940
rect 2276 4906 2277 4932
rect 2284 4906 2311 4932
rect 2219 4888 2249 4902
rect 2276 4898 2311 4906
rect 2313 4932 2354 4940
rect 2313 4906 2328 4932
rect 2335 4906 2354 4932
rect 2418 4928 2480 4940
rect 2492 4928 2567 4940
rect 2625 4928 2700 4940
rect 2712 4928 2743 4940
rect 2749 4928 2784 4940
rect 2418 4926 2580 4928
rect 2313 4898 2354 4906
rect 2436 4902 2449 4926
rect 2464 4924 2479 4926
rect 2276 4888 2277 4898
rect 2292 4888 2305 4898
rect 2319 4888 2320 4898
rect 2335 4888 2348 4898
rect 2363 4888 2393 4902
rect 2436 4888 2479 4902
rect 2503 4899 2510 4906
rect 2513 4902 2580 4926
rect 2612 4926 2784 4928
rect 2582 4904 2610 4908
rect 2612 4904 2692 4926
rect 2713 4924 2728 4926
rect 2582 4902 2692 4904
rect 2513 4898 2692 4902
rect 2486 4888 2516 4898
rect 2518 4888 2671 4898
rect 2679 4888 2709 4898
rect 2713 4888 2743 4902
rect 2771 4888 2784 4926
rect 2856 4932 2891 4940
rect 2856 4906 2857 4932
rect 2864 4906 2891 4932
rect 2799 4888 2829 4902
rect 2856 4898 2891 4906
rect 2893 4932 2934 4940
rect 2893 4906 2908 4932
rect 2915 4906 2934 4932
rect 2998 4928 3060 4940
rect 3072 4928 3147 4940
rect 3205 4928 3280 4940
rect 3292 4928 3323 4940
rect 3329 4928 3364 4940
rect 2998 4926 3160 4928
rect 2893 4898 2934 4906
rect 3016 4902 3029 4926
rect 3044 4924 3059 4926
rect 2856 4888 2857 4898
rect 2872 4888 2885 4898
rect 2899 4888 2900 4898
rect 2915 4888 2928 4898
rect 2943 4888 2973 4902
rect 3016 4888 3059 4902
rect 3083 4899 3090 4906
rect 3093 4902 3160 4926
rect 3192 4926 3364 4928
rect 3162 4904 3190 4908
rect 3192 4904 3272 4926
rect 3293 4924 3308 4926
rect 3162 4902 3272 4904
rect 3093 4898 3272 4902
rect 3066 4888 3096 4898
rect 3098 4888 3251 4898
rect 3259 4888 3289 4898
rect 3293 4888 3323 4902
rect 3351 4888 3364 4926
rect 3436 4932 3471 4940
rect 3436 4906 3437 4932
rect 3444 4906 3471 4932
rect 3379 4888 3409 4902
rect 3436 4898 3471 4906
rect 3473 4932 3514 4940
rect 3473 4906 3488 4932
rect 3495 4906 3514 4932
rect 3578 4928 3640 4940
rect 3652 4928 3727 4940
rect 3785 4928 3860 4940
rect 3872 4928 3903 4940
rect 3909 4928 3944 4940
rect 3578 4926 3740 4928
rect 3473 4898 3514 4906
rect 3596 4902 3609 4926
rect 3624 4924 3639 4926
rect 3436 4888 3437 4898
rect 3452 4888 3465 4898
rect 3479 4888 3480 4898
rect 3495 4888 3508 4898
rect 3523 4888 3553 4902
rect 3596 4888 3639 4902
rect 3663 4899 3670 4906
rect 3673 4902 3740 4926
rect 3772 4926 3944 4928
rect 3742 4904 3770 4908
rect 3772 4904 3852 4926
rect 3873 4924 3888 4926
rect 3742 4902 3852 4904
rect 3673 4898 3852 4902
rect 3646 4888 3676 4898
rect 3678 4888 3831 4898
rect 3839 4888 3869 4898
rect 3873 4888 3903 4902
rect 3931 4888 3944 4926
rect 4016 4932 4051 4940
rect 4016 4906 4017 4932
rect 4024 4906 4051 4932
rect 3959 4888 3989 4902
rect 4016 4898 4051 4906
rect 4053 4932 4094 4940
rect 4053 4906 4068 4932
rect 4075 4906 4094 4932
rect 4158 4928 4220 4940
rect 4232 4928 4307 4940
rect 4365 4928 4440 4940
rect 4452 4928 4483 4940
rect 4489 4928 4524 4940
rect 4158 4926 4320 4928
rect 4053 4898 4094 4906
rect 4176 4902 4189 4926
rect 4204 4924 4219 4926
rect 4016 4888 4017 4898
rect 4032 4888 4045 4898
rect 4059 4888 4060 4898
rect 4075 4888 4088 4898
rect 4103 4888 4133 4902
rect 4176 4888 4219 4902
rect 4243 4899 4250 4906
rect 4253 4902 4320 4926
rect 4352 4926 4524 4928
rect 4322 4904 4350 4908
rect 4352 4904 4432 4926
rect 4453 4924 4468 4926
rect 4322 4902 4432 4904
rect 4253 4898 4432 4902
rect 4226 4888 4256 4898
rect 4258 4888 4411 4898
rect 4419 4888 4449 4898
rect 4453 4888 4483 4902
rect 4511 4888 4524 4926
rect 4596 4932 4631 4940
rect 4596 4906 4597 4932
rect 4604 4906 4631 4932
rect 4539 4888 4569 4902
rect 4596 4898 4631 4906
rect 4633 4932 4674 4940
rect 4633 4906 4648 4932
rect 4655 4906 4674 4932
rect 4738 4928 4800 4940
rect 4812 4928 4887 4940
rect 4945 4928 5020 4940
rect 5032 4928 5063 4940
rect 5069 4928 5104 4940
rect 4738 4926 4900 4928
rect 4633 4898 4674 4906
rect 4756 4902 4769 4926
rect 4784 4924 4799 4926
rect 4596 4888 4597 4898
rect 4612 4888 4625 4898
rect 4639 4888 4640 4898
rect 4655 4888 4668 4898
rect 4683 4888 4713 4902
rect 4756 4888 4799 4902
rect 4823 4899 4830 4906
rect 4833 4902 4900 4926
rect 4932 4926 5104 4928
rect 4902 4904 4930 4908
rect 4932 4904 5012 4926
rect 5033 4924 5048 4926
rect 4902 4902 5012 4904
rect 4833 4898 5012 4902
rect 4806 4888 4836 4898
rect 4838 4888 4991 4898
rect 4999 4888 5029 4898
rect 5033 4888 5063 4902
rect 5091 4888 5104 4926
rect 5176 4932 5211 4940
rect 5176 4906 5177 4932
rect 5184 4906 5211 4932
rect 5119 4888 5149 4902
rect 5176 4898 5211 4906
rect 5213 4932 5254 4940
rect 5213 4906 5228 4932
rect 5235 4906 5254 4932
rect 5318 4928 5380 4940
rect 5392 4928 5467 4940
rect 5525 4928 5600 4940
rect 5612 4928 5643 4940
rect 5649 4928 5684 4940
rect 5318 4926 5480 4928
rect 5213 4898 5254 4906
rect 5336 4902 5349 4926
rect 5364 4924 5379 4926
rect 5176 4888 5177 4898
rect 5192 4888 5205 4898
rect 5219 4888 5220 4898
rect 5235 4888 5248 4898
rect 5263 4888 5293 4902
rect 5336 4888 5379 4902
rect 5403 4899 5410 4906
rect 5413 4902 5480 4926
rect 5512 4926 5684 4928
rect 5482 4904 5510 4908
rect 5512 4904 5592 4926
rect 5613 4924 5628 4926
rect 5482 4902 5592 4904
rect 5413 4898 5592 4902
rect 5386 4888 5416 4898
rect 5418 4888 5571 4898
rect 5579 4888 5609 4898
rect 5613 4888 5643 4902
rect 5671 4888 5684 4926
rect 5756 4932 5791 4940
rect 5756 4906 5757 4932
rect 5764 4906 5791 4932
rect 5699 4888 5729 4902
rect 5756 4898 5791 4906
rect 5793 4932 5834 4940
rect 5793 4906 5808 4932
rect 5815 4906 5834 4932
rect 5898 4928 5960 4940
rect 5972 4928 6047 4940
rect 6105 4928 6180 4940
rect 6192 4928 6223 4940
rect 6229 4928 6264 4940
rect 5898 4926 6060 4928
rect 5793 4898 5834 4906
rect 5916 4902 5929 4926
rect 5944 4924 5959 4926
rect 5756 4888 5757 4898
rect 5772 4888 5785 4898
rect 5799 4888 5800 4898
rect 5815 4888 5828 4898
rect 5843 4888 5873 4902
rect 5916 4888 5959 4902
rect 5983 4899 5990 4906
rect 5993 4902 6060 4926
rect 6092 4926 6264 4928
rect 6062 4904 6090 4908
rect 6092 4904 6172 4926
rect 6193 4924 6208 4926
rect 6062 4902 6172 4904
rect 5993 4898 6172 4902
rect 5966 4888 5996 4898
rect 5998 4888 6151 4898
rect 6159 4888 6189 4898
rect 6193 4888 6223 4902
rect 6251 4888 6264 4926
rect 6336 4932 6371 4940
rect 6336 4906 6337 4932
rect 6344 4906 6371 4932
rect 6279 4888 6309 4902
rect 6336 4898 6371 4906
rect 6373 4932 6414 4940
rect 6373 4906 6388 4932
rect 6395 4906 6414 4932
rect 6478 4928 6540 4940
rect 6552 4928 6627 4940
rect 6685 4928 6760 4940
rect 6772 4928 6803 4940
rect 6809 4928 6844 4940
rect 6478 4926 6640 4928
rect 6373 4898 6414 4906
rect 6496 4902 6509 4926
rect 6524 4924 6539 4926
rect 6336 4888 6337 4898
rect 6352 4888 6365 4898
rect 6379 4888 6380 4898
rect 6395 4888 6408 4898
rect 6423 4888 6453 4902
rect 6496 4888 6539 4902
rect 6563 4899 6570 4906
rect 6573 4902 6640 4926
rect 6672 4926 6844 4928
rect 6642 4904 6670 4908
rect 6672 4904 6752 4926
rect 6773 4924 6788 4926
rect 6642 4902 6752 4904
rect 6573 4898 6752 4902
rect 6546 4888 6576 4898
rect 6578 4888 6731 4898
rect 6739 4888 6769 4898
rect 6773 4888 6803 4902
rect 6831 4888 6844 4926
rect 6916 4932 6951 4940
rect 6916 4906 6917 4932
rect 6924 4906 6951 4932
rect 6859 4888 6889 4902
rect 6916 4898 6951 4906
rect 6953 4932 6994 4940
rect 6953 4906 6968 4932
rect 6975 4906 6994 4932
rect 7058 4928 7120 4940
rect 7132 4928 7207 4940
rect 7265 4928 7340 4940
rect 7352 4928 7383 4940
rect 7389 4928 7424 4940
rect 7058 4926 7220 4928
rect 6953 4898 6994 4906
rect 7076 4902 7089 4926
rect 7104 4924 7119 4926
rect 6916 4888 6917 4898
rect 6932 4888 6945 4898
rect 6959 4888 6960 4898
rect 6975 4888 6988 4898
rect 7003 4888 7033 4902
rect 7076 4888 7119 4902
rect 7143 4899 7150 4906
rect 7153 4902 7220 4926
rect 7252 4926 7424 4928
rect 7222 4904 7250 4908
rect 7252 4904 7332 4926
rect 7353 4924 7368 4926
rect 7222 4902 7332 4904
rect 7153 4898 7332 4902
rect 7126 4888 7156 4898
rect 7158 4888 7311 4898
rect 7319 4888 7349 4898
rect 7353 4888 7383 4902
rect 7411 4888 7424 4926
rect 7496 4932 7531 4940
rect 7496 4906 7497 4932
rect 7504 4906 7531 4932
rect 7439 4888 7469 4902
rect 7496 4898 7531 4906
rect 7533 4932 7574 4940
rect 7533 4906 7548 4932
rect 7555 4906 7574 4932
rect 7638 4928 7700 4940
rect 7712 4928 7787 4940
rect 7845 4928 7920 4940
rect 7932 4928 7963 4940
rect 7969 4928 8004 4940
rect 7638 4926 7800 4928
rect 7533 4898 7574 4906
rect 7656 4902 7669 4926
rect 7684 4924 7699 4926
rect 7496 4888 7497 4898
rect 7512 4888 7525 4898
rect 7539 4888 7540 4898
rect 7555 4888 7568 4898
rect 7583 4888 7613 4902
rect 7656 4888 7699 4902
rect 7723 4899 7730 4906
rect 7733 4902 7800 4926
rect 7832 4926 8004 4928
rect 7802 4904 7830 4908
rect 7832 4904 7912 4926
rect 7933 4924 7948 4926
rect 7802 4902 7912 4904
rect 7733 4898 7912 4902
rect 7706 4888 7736 4898
rect 7738 4888 7891 4898
rect 7899 4888 7929 4898
rect 7933 4888 7963 4902
rect 7991 4888 8004 4926
rect 8076 4932 8111 4940
rect 8076 4906 8077 4932
rect 8084 4906 8111 4932
rect 8019 4888 8049 4902
rect 8076 4898 8111 4906
rect 8113 4932 8154 4940
rect 8113 4906 8128 4932
rect 8135 4906 8154 4932
rect 8218 4928 8280 4940
rect 8292 4928 8367 4940
rect 8425 4928 8500 4940
rect 8512 4928 8543 4940
rect 8549 4928 8584 4940
rect 8218 4926 8380 4928
rect 8113 4898 8154 4906
rect 8236 4902 8249 4926
rect 8264 4924 8279 4926
rect 8076 4888 8077 4898
rect 8092 4888 8105 4898
rect 8119 4888 8120 4898
rect 8135 4888 8148 4898
rect 8163 4888 8193 4902
rect 8236 4888 8279 4902
rect 8303 4899 8310 4906
rect 8313 4902 8380 4926
rect 8412 4926 8584 4928
rect 8382 4904 8410 4908
rect 8412 4904 8492 4926
rect 8513 4924 8528 4926
rect 8382 4902 8492 4904
rect 8313 4898 8492 4902
rect 8286 4888 8316 4898
rect 8318 4888 8471 4898
rect 8479 4888 8509 4898
rect 8513 4888 8543 4902
rect 8571 4888 8584 4926
rect 8656 4932 8691 4940
rect 8656 4906 8657 4932
rect 8664 4906 8691 4932
rect 8599 4888 8629 4902
rect 8656 4898 8691 4906
rect 8693 4932 8734 4940
rect 8693 4906 8708 4932
rect 8715 4906 8734 4932
rect 8798 4928 8860 4940
rect 8872 4928 8947 4940
rect 9005 4928 9080 4940
rect 9092 4928 9123 4940
rect 9129 4928 9164 4940
rect 8798 4926 8960 4928
rect 8693 4898 8734 4906
rect 8816 4902 8829 4926
rect 8844 4924 8859 4926
rect 8656 4888 8657 4898
rect 8672 4888 8685 4898
rect 8699 4888 8700 4898
rect 8715 4888 8728 4898
rect 8743 4888 8773 4902
rect 8816 4888 8859 4902
rect 8883 4899 8890 4906
rect 8893 4902 8960 4926
rect 8992 4926 9164 4928
rect 8962 4904 8990 4908
rect 8992 4904 9072 4926
rect 9093 4924 9108 4926
rect 8962 4902 9072 4904
rect 8893 4898 9072 4902
rect 8866 4888 8896 4898
rect 8898 4888 9051 4898
rect 9059 4888 9089 4898
rect 9093 4888 9123 4902
rect 9151 4888 9164 4926
rect 9236 4932 9271 4940
rect 9236 4906 9237 4932
rect 9244 4906 9271 4932
rect 9179 4888 9209 4902
rect 9236 4898 9271 4906
rect 9236 4888 9237 4898
rect 9252 4888 9265 4898
rect -1 4882 9265 4888
rect 0 4874 9265 4882
rect 15 4844 28 4874
rect 43 4856 73 4874
rect 116 4860 130 4874
rect 166 4860 386 4874
rect 117 4858 130 4860
rect 83 4846 98 4858
rect 80 4844 102 4846
rect 107 4844 137 4858
rect 198 4856 351 4860
rect 180 4844 372 4856
rect 415 4844 445 4858
rect 451 4844 464 4874
rect 479 4856 509 4874
rect 552 4844 565 4874
rect 595 4844 608 4874
rect 623 4856 653 4874
rect 696 4860 710 4874
rect 746 4860 966 4874
rect 697 4858 710 4860
rect 663 4846 678 4858
rect 660 4844 682 4846
rect 687 4844 717 4858
rect 778 4856 931 4860
rect 760 4844 952 4856
rect 995 4844 1025 4858
rect 1031 4844 1044 4874
rect 1059 4856 1089 4874
rect 1132 4844 1145 4874
rect 1175 4844 1188 4874
rect 1203 4856 1233 4874
rect 1276 4860 1290 4874
rect 1326 4860 1546 4874
rect 1277 4858 1290 4860
rect 1243 4846 1258 4858
rect 1240 4844 1262 4846
rect 1267 4844 1297 4858
rect 1358 4856 1511 4860
rect 1340 4844 1532 4856
rect 1575 4844 1605 4858
rect 1611 4844 1624 4874
rect 1639 4856 1669 4874
rect 1712 4844 1725 4874
rect 1755 4844 1768 4874
rect 1783 4856 1813 4874
rect 1856 4860 1870 4874
rect 1906 4860 2126 4874
rect 1857 4858 1870 4860
rect 1823 4846 1838 4858
rect 1820 4844 1842 4846
rect 1847 4844 1877 4858
rect 1938 4856 2091 4860
rect 1920 4844 2112 4856
rect 2155 4844 2185 4858
rect 2191 4844 2204 4874
rect 2219 4856 2249 4874
rect 2292 4844 2305 4874
rect 2335 4844 2348 4874
rect 2363 4856 2393 4874
rect 2436 4860 2450 4874
rect 2486 4860 2706 4874
rect 2437 4858 2450 4860
rect 2403 4846 2418 4858
rect 2400 4844 2422 4846
rect 2427 4844 2457 4858
rect 2518 4856 2671 4860
rect 2500 4844 2692 4856
rect 2735 4844 2765 4858
rect 2771 4844 2784 4874
rect 2799 4856 2829 4874
rect 2872 4844 2885 4874
rect 2915 4844 2928 4874
rect 2943 4856 2973 4874
rect 3016 4860 3030 4874
rect 3066 4860 3286 4874
rect 3017 4858 3030 4860
rect 2983 4846 2998 4858
rect 2980 4844 3002 4846
rect 3007 4844 3037 4858
rect 3098 4856 3251 4860
rect 3080 4844 3272 4856
rect 3315 4844 3345 4858
rect 3351 4844 3364 4874
rect 3379 4856 3409 4874
rect 3452 4844 3465 4874
rect 3495 4844 3508 4874
rect 3523 4856 3553 4874
rect 3596 4860 3610 4874
rect 3646 4860 3866 4874
rect 3597 4858 3610 4860
rect 3563 4846 3578 4858
rect 3560 4844 3582 4846
rect 3587 4844 3617 4858
rect 3678 4856 3831 4860
rect 3660 4844 3852 4856
rect 3895 4844 3925 4858
rect 3931 4844 3944 4874
rect 3959 4856 3989 4874
rect 4032 4844 4045 4874
rect 4075 4844 4088 4874
rect 4103 4856 4133 4874
rect 4176 4860 4190 4874
rect 4226 4860 4446 4874
rect 4177 4858 4190 4860
rect 4143 4846 4158 4858
rect 4140 4844 4162 4846
rect 4167 4844 4197 4858
rect 4258 4856 4411 4860
rect 4240 4844 4432 4856
rect 4475 4844 4505 4858
rect 4511 4844 4524 4874
rect 4539 4856 4569 4874
rect 4612 4844 4625 4874
rect 4655 4844 4668 4874
rect 4683 4856 4713 4874
rect 4756 4860 4770 4874
rect 4806 4860 5026 4874
rect 4757 4858 4770 4860
rect 4723 4846 4738 4858
rect 4720 4844 4742 4846
rect 4747 4844 4777 4858
rect 4838 4856 4991 4860
rect 4820 4844 5012 4856
rect 5055 4844 5085 4858
rect 5091 4844 5104 4874
rect 5119 4856 5149 4874
rect 5192 4844 5205 4874
rect 5235 4844 5248 4874
rect 5263 4856 5293 4874
rect 5336 4860 5350 4874
rect 5386 4860 5606 4874
rect 5337 4858 5350 4860
rect 5303 4846 5318 4858
rect 5300 4844 5322 4846
rect 5327 4844 5357 4858
rect 5418 4856 5571 4860
rect 5400 4844 5592 4856
rect 5635 4844 5665 4858
rect 5671 4844 5684 4874
rect 5699 4856 5729 4874
rect 5772 4844 5785 4874
rect 5815 4844 5828 4874
rect 5843 4856 5873 4874
rect 5916 4860 5930 4874
rect 5966 4860 6186 4874
rect 5917 4858 5930 4860
rect 5883 4846 5898 4858
rect 5880 4844 5902 4846
rect 5907 4844 5937 4858
rect 5998 4856 6151 4860
rect 5980 4844 6172 4856
rect 6215 4844 6245 4858
rect 6251 4844 6264 4874
rect 6279 4856 6309 4874
rect 6352 4844 6365 4874
rect 6395 4844 6408 4874
rect 6423 4856 6453 4874
rect 6496 4860 6510 4874
rect 6546 4860 6766 4874
rect 6497 4858 6510 4860
rect 6463 4846 6478 4858
rect 6460 4844 6482 4846
rect 6487 4844 6517 4858
rect 6578 4856 6731 4860
rect 6560 4844 6752 4856
rect 6795 4844 6825 4858
rect 6831 4844 6844 4874
rect 6859 4856 6889 4874
rect 6932 4844 6945 4874
rect 6975 4844 6988 4874
rect 7003 4856 7033 4874
rect 7076 4860 7090 4874
rect 7126 4860 7346 4874
rect 7077 4858 7090 4860
rect 7043 4846 7058 4858
rect 7040 4844 7062 4846
rect 7067 4844 7097 4858
rect 7158 4856 7311 4860
rect 7140 4844 7332 4856
rect 7375 4844 7405 4858
rect 7411 4844 7424 4874
rect 7439 4856 7469 4874
rect 7512 4844 7525 4874
rect 7555 4844 7568 4874
rect 7583 4856 7613 4874
rect 7656 4860 7670 4874
rect 7706 4860 7926 4874
rect 7657 4858 7670 4860
rect 7623 4846 7638 4858
rect 7620 4844 7642 4846
rect 7647 4844 7677 4858
rect 7738 4856 7891 4860
rect 7720 4844 7912 4856
rect 7955 4844 7985 4858
rect 7991 4844 8004 4874
rect 8019 4856 8049 4874
rect 8092 4844 8105 4874
rect 8135 4844 8148 4874
rect 8163 4856 8193 4874
rect 8236 4860 8250 4874
rect 8286 4860 8506 4874
rect 8237 4858 8250 4860
rect 8203 4846 8218 4858
rect 8200 4844 8222 4846
rect 8227 4844 8257 4858
rect 8318 4856 8471 4860
rect 8300 4844 8492 4856
rect 8535 4844 8565 4858
rect 8571 4844 8584 4874
rect 8599 4856 8629 4874
rect 8672 4844 8685 4874
rect 8715 4844 8728 4874
rect 8743 4856 8773 4874
rect 8816 4860 8830 4874
rect 8866 4860 9086 4874
rect 8817 4858 8830 4860
rect 8783 4846 8798 4858
rect 8780 4844 8802 4846
rect 8807 4844 8837 4858
rect 8898 4856 9051 4860
rect 8880 4844 9072 4856
rect 9115 4844 9145 4858
rect 9151 4844 9164 4874
rect 9179 4856 9209 4874
rect 9252 4844 9265 4874
rect 0 4830 9265 4844
rect 15 4726 28 4830
rect 73 4808 74 4818
rect 89 4808 102 4818
rect 73 4804 102 4808
rect 107 4804 137 4830
rect 155 4816 171 4818
rect 243 4816 296 4830
rect 244 4814 308 4816
rect 351 4814 366 4830
rect 415 4827 445 4830
rect 415 4824 451 4827
rect 381 4816 397 4818
rect 155 4804 170 4808
rect 73 4802 170 4804
rect 198 4802 366 4814
rect 382 4804 397 4808
rect 415 4805 454 4824
rect 473 4818 480 4819
rect 479 4811 480 4818
rect 463 4808 464 4811
rect 479 4808 492 4811
rect 415 4804 445 4805
rect 454 4804 460 4805
rect 463 4804 492 4808
rect 382 4803 492 4804
rect 382 4802 498 4803
rect 57 4794 108 4802
rect 57 4782 82 4794
rect 89 4782 108 4794
rect 139 4794 189 4802
rect 139 4786 155 4794
rect 162 4792 189 4794
rect 198 4792 419 4802
rect 162 4782 419 4792
rect 448 4794 498 4802
rect 448 4785 464 4794
rect 57 4774 108 4782
rect 155 4774 419 4782
rect 445 4782 464 4785
rect 471 4782 498 4794
rect 445 4774 498 4782
rect 73 4766 74 4774
rect 89 4766 102 4774
rect 73 4758 89 4766
rect 70 4751 89 4754
rect 70 4742 92 4751
rect 43 4732 92 4742
rect 43 4726 73 4732
rect 92 4727 97 4732
rect 15 4710 89 4726
rect 107 4718 137 4774
rect 172 4764 380 4774
rect 415 4770 460 4774
rect 463 4773 464 4774
rect 479 4773 492 4774
rect 198 4734 387 4764
rect 213 4731 387 4734
rect 206 4728 387 4731
rect 15 4708 28 4710
rect 43 4708 77 4710
rect 15 4692 89 4708
rect 116 4704 129 4718
rect 144 4704 160 4720
rect 206 4715 217 4728
rect -1 4670 0 4686
rect 15 4670 28 4692
rect 43 4670 73 4692
rect 116 4688 178 4704
rect 206 4697 217 4713
rect 222 4708 232 4728
rect 242 4708 256 4728
rect 259 4715 268 4728
rect 284 4715 293 4728
rect 222 4697 256 4708
rect 259 4697 268 4713
rect 284 4697 293 4713
rect 300 4708 310 4728
rect 320 4708 334 4728
rect 335 4715 346 4728
rect 300 4697 334 4708
rect 335 4697 346 4713
rect 392 4704 408 4720
rect 415 4718 445 4770
rect 479 4766 480 4773
rect 464 4758 480 4766
rect 451 4726 464 4745
rect 479 4726 509 4742
rect 451 4710 525 4726
rect 451 4708 464 4710
rect 479 4708 513 4710
rect 116 4686 129 4688
rect 144 4686 178 4688
rect 116 4670 178 4686
rect 222 4681 238 4684
rect 300 4681 330 4692
rect 378 4688 424 4704
rect 451 4692 525 4708
rect 378 4686 412 4688
rect 377 4670 424 4686
rect 451 4670 464 4692
rect 479 4670 509 4692
rect 536 4670 537 4686
rect 552 4670 565 4830
rect 595 4726 608 4830
rect 653 4808 654 4818
rect 669 4808 682 4818
rect 653 4804 682 4808
rect 687 4804 717 4830
rect 735 4816 751 4818
rect 823 4816 876 4830
rect 824 4814 888 4816
rect 931 4814 946 4830
rect 995 4827 1025 4830
rect 995 4824 1031 4827
rect 961 4816 977 4818
rect 735 4804 750 4808
rect 653 4802 750 4804
rect 778 4802 946 4814
rect 962 4804 977 4808
rect 995 4805 1034 4824
rect 1053 4818 1060 4819
rect 1059 4811 1060 4818
rect 1043 4808 1044 4811
rect 1059 4808 1072 4811
rect 995 4804 1025 4805
rect 1034 4804 1040 4805
rect 1043 4804 1072 4808
rect 962 4803 1072 4804
rect 962 4802 1078 4803
rect 637 4794 688 4802
rect 637 4782 662 4794
rect 669 4782 688 4794
rect 719 4794 769 4802
rect 719 4786 735 4794
rect 742 4792 769 4794
rect 778 4792 999 4802
rect 742 4782 999 4792
rect 1028 4794 1078 4802
rect 1028 4785 1044 4794
rect 637 4774 688 4782
rect 735 4774 999 4782
rect 1025 4782 1044 4785
rect 1051 4782 1078 4794
rect 1025 4774 1078 4782
rect 653 4766 654 4774
rect 669 4766 682 4774
rect 653 4758 669 4766
rect 650 4751 669 4754
rect 650 4742 672 4751
rect 623 4732 672 4742
rect 623 4726 653 4732
rect 672 4727 677 4732
rect 595 4710 669 4726
rect 687 4718 717 4774
rect 752 4764 960 4774
rect 995 4770 1040 4774
rect 1043 4773 1044 4774
rect 1059 4773 1072 4774
rect 778 4734 967 4764
rect 793 4731 967 4734
rect 786 4728 967 4731
rect 595 4708 608 4710
rect 623 4708 657 4710
rect 595 4692 669 4708
rect 696 4704 709 4718
rect 724 4704 740 4720
rect 786 4715 797 4728
rect 579 4670 580 4686
rect 595 4670 608 4692
rect 623 4670 653 4692
rect 696 4688 758 4704
rect 786 4697 797 4713
rect 802 4708 812 4728
rect 822 4708 836 4728
rect 839 4715 848 4728
rect 864 4715 873 4728
rect 802 4697 836 4708
rect 839 4697 848 4713
rect 864 4697 873 4713
rect 880 4708 890 4728
rect 900 4708 914 4728
rect 915 4715 926 4728
rect 880 4697 914 4708
rect 915 4697 926 4713
rect 972 4704 988 4720
rect 995 4718 1025 4770
rect 1059 4766 1060 4773
rect 1044 4758 1060 4766
rect 1031 4726 1044 4745
rect 1059 4726 1089 4742
rect 1031 4710 1105 4726
rect 1031 4708 1044 4710
rect 1059 4708 1093 4710
rect 696 4686 709 4688
rect 724 4686 758 4688
rect 696 4670 758 4686
rect 802 4681 818 4684
rect 880 4681 910 4692
rect 958 4688 1004 4704
rect 1031 4692 1105 4708
rect 958 4686 992 4688
rect 957 4670 1004 4686
rect 1031 4670 1044 4692
rect 1059 4670 1089 4692
rect 1116 4670 1117 4686
rect 1132 4670 1145 4830
rect 1175 4726 1188 4830
rect 1233 4808 1234 4818
rect 1249 4808 1262 4818
rect 1233 4804 1262 4808
rect 1267 4804 1297 4830
rect 1315 4816 1331 4818
rect 1403 4816 1456 4830
rect 1404 4814 1468 4816
rect 1511 4814 1526 4830
rect 1575 4827 1605 4830
rect 1575 4824 1611 4827
rect 1541 4816 1557 4818
rect 1315 4804 1330 4808
rect 1233 4802 1330 4804
rect 1358 4802 1526 4814
rect 1542 4804 1557 4808
rect 1575 4805 1614 4824
rect 1633 4818 1640 4819
rect 1639 4811 1640 4818
rect 1623 4808 1624 4811
rect 1639 4808 1652 4811
rect 1575 4804 1605 4805
rect 1614 4804 1620 4805
rect 1623 4804 1652 4808
rect 1542 4803 1652 4804
rect 1542 4802 1658 4803
rect 1217 4794 1268 4802
rect 1217 4782 1242 4794
rect 1249 4782 1268 4794
rect 1299 4794 1349 4802
rect 1299 4786 1315 4794
rect 1322 4792 1349 4794
rect 1358 4792 1579 4802
rect 1322 4782 1579 4792
rect 1608 4794 1658 4802
rect 1608 4785 1624 4794
rect 1217 4774 1268 4782
rect 1315 4774 1579 4782
rect 1605 4782 1624 4785
rect 1631 4782 1658 4794
rect 1605 4774 1658 4782
rect 1233 4766 1234 4774
rect 1249 4766 1262 4774
rect 1233 4758 1249 4766
rect 1230 4751 1249 4754
rect 1230 4742 1252 4751
rect 1203 4732 1252 4742
rect 1203 4726 1233 4732
rect 1252 4727 1257 4732
rect 1175 4710 1249 4726
rect 1267 4718 1297 4774
rect 1332 4764 1540 4774
rect 1575 4770 1620 4774
rect 1623 4773 1624 4774
rect 1639 4773 1652 4774
rect 1358 4734 1547 4764
rect 1373 4731 1547 4734
rect 1366 4728 1547 4731
rect 1175 4708 1188 4710
rect 1203 4708 1237 4710
rect 1175 4692 1249 4708
rect 1276 4704 1289 4718
rect 1304 4704 1320 4720
rect 1366 4715 1377 4728
rect 1159 4670 1160 4686
rect 1175 4670 1188 4692
rect 1203 4670 1233 4692
rect 1276 4688 1338 4704
rect 1366 4697 1377 4713
rect 1382 4708 1392 4728
rect 1402 4708 1416 4728
rect 1419 4715 1428 4728
rect 1444 4715 1453 4728
rect 1382 4697 1416 4708
rect 1419 4697 1428 4713
rect 1444 4697 1453 4713
rect 1460 4708 1470 4728
rect 1480 4708 1494 4728
rect 1495 4715 1506 4728
rect 1460 4697 1494 4708
rect 1495 4697 1506 4713
rect 1552 4704 1568 4720
rect 1575 4718 1605 4770
rect 1639 4766 1640 4773
rect 1624 4758 1640 4766
rect 1611 4726 1624 4745
rect 1639 4726 1669 4742
rect 1611 4710 1685 4726
rect 1611 4708 1624 4710
rect 1639 4708 1673 4710
rect 1276 4686 1289 4688
rect 1304 4686 1338 4688
rect 1276 4670 1338 4686
rect 1382 4681 1398 4684
rect 1460 4681 1490 4692
rect 1538 4688 1584 4704
rect 1611 4692 1685 4708
rect 1538 4686 1572 4688
rect 1537 4670 1584 4686
rect 1611 4670 1624 4692
rect 1639 4670 1669 4692
rect 1696 4670 1697 4686
rect 1712 4670 1725 4830
rect 1755 4726 1768 4830
rect 1813 4808 1814 4818
rect 1829 4808 1842 4818
rect 1813 4804 1842 4808
rect 1847 4804 1877 4830
rect 1895 4816 1911 4818
rect 1983 4816 2036 4830
rect 1984 4814 2048 4816
rect 2091 4814 2106 4830
rect 2155 4827 2185 4830
rect 2155 4824 2191 4827
rect 2121 4816 2137 4818
rect 1895 4804 1910 4808
rect 1813 4802 1910 4804
rect 1938 4802 2106 4814
rect 2122 4804 2137 4808
rect 2155 4805 2194 4824
rect 2213 4818 2220 4819
rect 2219 4811 2220 4818
rect 2203 4808 2204 4811
rect 2219 4808 2232 4811
rect 2155 4804 2185 4805
rect 2194 4804 2200 4805
rect 2203 4804 2232 4808
rect 2122 4803 2232 4804
rect 2122 4802 2238 4803
rect 1797 4794 1848 4802
rect 1797 4782 1822 4794
rect 1829 4782 1848 4794
rect 1879 4794 1929 4802
rect 1879 4786 1895 4794
rect 1902 4792 1929 4794
rect 1938 4792 2159 4802
rect 1902 4782 2159 4792
rect 2188 4794 2238 4802
rect 2188 4785 2204 4794
rect 1797 4774 1848 4782
rect 1895 4774 2159 4782
rect 2185 4782 2204 4785
rect 2211 4782 2238 4794
rect 2185 4774 2238 4782
rect 1813 4766 1814 4774
rect 1829 4766 1842 4774
rect 1813 4758 1829 4766
rect 1810 4751 1829 4754
rect 1810 4742 1832 4751
rect 1783 4732 1832 4742
rect 1783 4726 1813 4732
rect 1832 4727 1837 4732
rect 1755 4710 1829 4726
rect 1847 4718 1877 4774
rect 1912 4764 2120 4774
rect 2155 4770 2200 4774
rect 2203 4773 2204 4774
rect 2219 4773 2232 4774
rect 1938 4734 2127 4764
rect 1953 4731 2127 4734
rect 1946 4728 2127 4731
rect 1755 4708 1768 4710
rect 1783 4708 1817 4710
rect 1755 4692 1829 4708
rect 1856 4704 1869 4718
rect 1884 4704 1900 4720
rect 1946 4715 1957 4728
rect 1739 4670 1740 4686
rect 1755 4670 1768 4692
rect 1783 4670 1813 4692
rect 1856 4688 1918 4704
rect 1946 4697 1957 4713
rect 1962 4708 1972 4728
rect 1982 4708 1996 4728
rect 1999 4715 2008 4728
rect 2024 4715 2033 4728
rect 1962 4697 1996 4708
rect 1999 4697 2008 4713
rect 2024 4697 2033 4713
rect 2040 4708 2050 4728
rect 2060 4708 2074 4728
rect 2075 4715 2086 4728
rect 2040 4697 2074 4708
rect 2075 4697 2086 4713
rect 2132 4704 2148 4720
rect 2155 4718 2185 4770
rect 2219 4766 2220 4773
rect 2204 4758 2220 4766
rect 2191 4726 2204 4745
rect 2219 4726 2249 4742
rect 2191 4710 2265 4726
rect 2191 4708 2204 4710
rect 2219 4708 2253 4710
rect 1856 4686 1869 4688
rect 1884 4686 1918 4688
rect 1856 4670 1918 4686
rect 1962 4681 1976 4684
rect 2040 4681 2070 4692
rect 2118 4688 2164 4704
rect 2191 4692 2265 4708
rect 2118 4686 2152 4688
rect 2117 4670 2164 4686
rect 2191 4670 2204 4692
rect 2219 4670 2249 4692
rect 2276 4670 2277 4686
rect 2292 4670 2305 4830
rect 2335 4726 2348 4830
rect 2393 4808 2394 4818
rect 2409 4808 2422 4818
rect 2393 4804 2422 4808
rect 2427 4804 2457 4830
rect 2475 4816 2491 4818
rect 2563 4816 2616 4830
rect 2564 4814 2628 4816
rect 2671 4814 2686 4830
rect 2735 4827 2765 4830
rect 2735 4824 2771 4827
rect 2701 4816 2717 4818
rect 2475 4804 2490 4808
rect 2393 4802 2490 4804
rect 2518 4802 2686 4814
rect 2702 4804 2717 4808
rect 2735 4805 2774 4824
rect 2793 4818 2800 4819
rect 2799 4811 2800 4818
rect 2783 4808 2784 4811
rect 2799 4808 2812 4811
rect 2735 4804 2765 4805
rect 2774 4804 2780 4805
rect 2783 4804 2812 4808
rect 2702 4803 2812 4804
rect 2702 4802 2818 4803
rect 2377 4794 2428 4802
rect 2377 4782 2402 4794
rect 2409 4782 2428 4794
rect 2459 4794 2509 4802
rect 2459 4786 2475 4794
rect 2482 4792 2509 4794
rect 2518 4792 2739 4802
rect 2482 4782 2739 4792
rect 2768 4794 2818 4802
rect 2768 4785 2784 4794
rect 2377 4774 2428 4782
rect 2475 4774 2739 4782
rect 2765 4782 2784 4785
rect 2791 4782 2818 4794
rect 2765 4774 2818 4782
rect 2393 4766 2394 4774
rect 2409 4766 2422 4774
rect 2393 4758 2409 4766
rect 2390 4751 2409 4754
rect 2390 4742 2412 4751
rect 2363 4732 2412 4742
rect 2363 4726 2393 4732
rect 2412 4727 2417 4732
rect 2335 4710 2409 4726
rect 2427 4718 2457 4774
rect 2492 4764 2700 4774
rect 2735 4770 2780 4774
rect 2783 4773 2784 4774
rect 2799 4773 2812 4774
rect 2518 4734 2707 4764
rect 2533 4731 2707 4734
rect 2526 4728 2707 4731
rect 2335 4708 2348 4710
rect 2363 4708 2397 4710
rect 2335 4692 2409 4708
rect 2436 4704 2449 4718
rect 2464 4704 2480 4720
rect 2526 4715 2537 4728
rect 2319 4670 2320 4686
rect 2335 4670 2348 4692
rect 2363 4670 2393 4692
rect 2436 4688 2498 4704
rect 2526 4697 2537 4713
rect 2542 4708 2552 4728
rect 2562 4708 2576 4728
rect 2579 4715 2588 4728
rect 2604 4715 2613 4728
rect 2542 4697 2576 4708
rect 2579 4697 2588 4713
rect 2604 4697 2613 4713
rect 2620 4708 2630 4728
rect 2640 4708 2654 4728
rect 2655 4715 2666 4728
rect 2620 4697 2654 4708
rect 2655 4697 2666 4713
rect 2712 4704 2728 4720
rect 2735 4718 2765 4770
rect 2799 4766 2800 4773
rect 2784 4758 2800 4766
rect 2771 4726 2784 4745
rect 2799 4726 2829 4742
rect 2771 4710 2845 4726
rect 2771 4708 2784 4710
rect 2799 4708 2833 4710
rect 2436 4686 2449 4688
rect 2464 4686 2498 4688
rect 2436 4670 2498 4686
rect 2542 4681 2558 4684
rect 2620 4681 2650 4692
rect 2698 4688 2744 4704
rect 2771 4692 2845 4708
rect 2698 4686 2732 4688
rect 2697 4670 2744 4686
rect 2771 4670 2784 4692
rect 2799 4670 2829 4692
rect 2856 4670 2857 4686
rect 2872 4670 2885 4830
rect 2915 4726 2928 4830
rect 2973 4808 2974 4818
rect 2989 4808 3002 4818
rect 2973 4804 3002 4808
rect 3007 4804 3037 4830
rect 3055 4816 3071 4818
rect 3143 4816 3196 4830
rect 3144 4814 3208 4816
rect 3251 4814 3266 4830
rect 3315 4827 3345 4830
rect 3315 4824 3351 4827
rect 3281 4816 3297 4818
rect 3055 4804 3070 4808
rect 2973 4802 3070 4804
rect 3098 4802 3266 4814
rect 3282 4804 3297 4808
rect 3315 4805 3354 4824
rect 3373 4818 3380 4819
rect 3379 4811 3380 4818
rect 3363 4808 3364 4811
rect 3379 4808 3392 4811
rect 3315 4804 3345 4805
rect 3354 4804 3360 4805
rect 3363 4804 3392 4808
rect 3282 4803 3392 4804
rect 3282 4802 3398 4803
rect 2957 4794 3008 4802
rect 2957 4782 2982 4794
rect 2989 4782 3008 4794
rect 3039 4794 3089 4802
rect 3039 4786 3055 4794
rect 3062 4792 3089 4794
rect 3098 4792 3319 4802
rect 3062 4782 3319 4792
rect 3348 4794 3398 4802
rect 3348 4785 3364 4794
rect 2957 4774 3008 4782
rect 3055 4774 3319 4782
rect 3345 4782 3364 4785
rect 3371 4782 3398 4794
rect 3345 4774 3398 4782
rect 2973 4766 2974 4774
rect 2989 4766 3002 4774
rect 2973 4758 2989 4766
rect 2970 4751 2989 4754
rect 2970 4742 2992 4751
rect 2943 4732 2992 4742
rect 2943 4726 2973 4732
rect 2992 4727 2997 4732
rect 2915 4710 2989 4726
rect 3007 4718 3037 4774
rect 3072 4764 3280 4774
rect 3315 4770 3360 4774
rect 3363 4773 3364 4774
rect 3379 4773 3392 4774
rect 3098 4734 3287 4764
rect 3113 4731 3287 4734
rect 3106 4728 3287 4731
rect 2915 4708 2928 4710
rect 2943 4708 2977 4710
rect 2915 4692 2989 4708
rect 3016 4704 3029 4718
rect 3044 4704 3060 4720
rect 3106 4715 3117 4728
rect 2899 4670 2900 4686
rect 2915 4670 2928 4692
rect 2943 4670 2973 4692
rect 3016 4688 3078 4704
rect 3106 4697 3117 4713
rect 3122 4708 3132 4728
rect 3142 4708 3156 4728
rect 3159 4715 3168 4728
rect 3184 4715 3193 4728
rect 3122 4697 3156 4708
rect 3159 4697 3168 4713
rect 3184 4697 3193 4713
rect 3200 4708 3210 4728
rect 3220 4708 3234 4728
rect 3235 4715 3246 4728
rect 3200 4697 3234 4708
rect 3235 4697 3246 4713
rect 3292 4704 3308 4720
rect 3315 4718 3345 4770
rect 3379 4766 3380 4773
rect 3364 4758 3380 4766
rect 3351 4726 3364 4745
rect 3379 4726 3409 4742
rect 3351 4710 3425 4726
rect 3351 4708 3364 4710
rect 3379 4708 3413 4710
rect 3016 4686 3029 4688
rect 3044 4686 3078 4688
rect 3016 4670 3078 4686
rect 3122 4681 3138 4684
rect 3200 4681 3230 4692
rect 3278 4688 3324 4704
rect 3351 4692 3425 4708
rect 3278 4686 3312 4688
rect 3277 4670 3324 4686
rect 3351 4670 3364 4692
rect 3379 4670 3409 4692
rect 3436 4670 3437 4686
rect 3452 4670 3465 4830
rect 3495 4726 3508 4830
rect 3553 4808 3554 4818
rect 3569 4808 3582 4818
rect 3553 4804 3582 4808
rect 3587 4804 3617 4830
rect 3635 4816 3651 4818
rect 3723 4816 3776 4830
rect 3724 4814 3788 4816
rect 3831 4814 3846 4830
rect 3895 4827 3925 4830
rect 3895 4824 3931 4827
rect 3861 4816 3877 4818
rect 3635 4804 3650 4808
rect 3553 4802 3650 4804
rect 3678 4802 3846 4814
rect 3862 4804 3877 4808
rect 3895 4805 3934 4824
rect 3953 4818 3960 4819
rect 3959 4811 3960 4818
rect 3943 4808 3944 4811
rect 3959 4808 3972 4811
rect 3895 4804 3925 4805
rect 3934 4804 3940 4805
rect 3943 4804 3972 4808
rect 3862 4803 3972 4804
rect 3862 4802 3978 4803
rect 3537 4794 3588 4802
rect 3537 4782 3562 4794
rect 3569 4782 3588 4794
rect 3619 4794 3669 4802
rect 3619 4786 3635 4794
rect 3642 4792 3669 4794
rect 3678 4792 3899 4802
rect 3642 4782 3899 4792
rect 3928 4794 3978 4802
rect 3928 4785 3944 4794
rect 3537 4774 3588 4782
rect 3635 4774 3899 4782
rect 3925 4782 3944 4785
rect 3951 4782 3978 4794
rect 3925 4774 3978 4782
rect 3553 4766 3554 4774
rect 3569 4766 3582 4774
rect 3553 4758 3569 4766
rect 3550 4751 3569 4754
rect 3550 4742 3572 4751
rect 3523 4732 3572 4742
rect 3523 4726 3553 4732
rect 3572 4727 3577 4732
rect 3495 4710 3569 4726
rect 3587 4718 3617 4774
rect 3652 4764 3860 4774
rect 3895 4770 3940 4774
rect 3943 4773 3944 4774
rect 3959 4773 3972 4774
rect 3678 4734 3867 4764
rect 3693 4731 3867 4734
rect 3686 4728 3867 4731
rect 3495 4708 3508 4710
rect 3523 4708 3557 4710
rect 3495 4692 3569 4708
rect 3596 4704 3609 4718
rect 3624 4704 3640 4720
rect 3686 4715 3697 4728
rect 3479 4670 3480 4686
rect 3495 4670 3508 4692
rect 3523 4670 3553 4692
rect 3596 4688 3658 4704
rect 3686 4697 3697 4713
rect 3702 4708 3712 4728
rect 3722 4708 3736 4728
rect 3739 4715 3748 4728
rect 3764 4715 3773 4728
rect 3702 4697 3736 4708
rect 3739 4697 3748 4713
rect 3764 4697 3773 4713
rect 3780 4708 3790 4728
rect 3800 4708 3814 4728
rect 3815 4715 3826 4728
rect 3780 4697 3814 4708
rect 3815 4697 3826 4713
rect 3872 4704 3888 4720
rect 3895 4718 3925 4770
rect 3959 4766 3960 4773
rect 3944 4758 3960 4766
rect 3931 4726 3944 4745
rect 3959 4726 3989 4742
rect 3931 4710 4005 4726
rect 3931 4708 3944 4710
rect 3959 4708 3993 4710
rect 3596 4686 3609 4688
rect 3624 4686 3658 4688
rect 3596 4670 3658 4686
rect 3702 4681 3718 4684
rect 3780 4681 3810 4692
rect 3858 4688 3904 4704
rect 3931 4692 4005 4708
rect 3858 4686 3892 4688
rect 3857 4670 3904 4686
rect 3931 4670 3944 4692
rect 3959 4670 3989 4692
rect 4016 4670 4017 4686
rect 4032 4670 4045 4830
rect 4075 4726 4088 4830
rect 4133 4808 4134 4818
rect 4149 4808 4162 4818
rect 4133 4804 4162 4808
rect 4167 4804 4197 4830
rect 4215 4816 4231 4818
rect 4303 4816 4356 4830
rect 4304 4814 4368 4816
rect 4411 4814 4426 4830
rect 4475 4827 4505 4830
rect 4475 4824 4511 4827
rect 4441 4816 4457 4818
rect 4215 4804 4230 4808
rect 4133 4802 4230 4804
rect 4258 4802 4426 4814
rect 4442 4804 4457 4808
rect 4475 4805 4514 4824
rect 4533 4818 4540 4819
rect 4539 4811 4540 4818
rect 4523 4808 4524 4811
rect 4539 4808 4552 4811
rect 4475 4804 4505 4805
rect 4514 4804 4520 4805
rect 4523 4804 4552 4808
rect 4442 4803 4552 4804
rect 4442 4802 4558 4803
rect 4117 4794 4168 4802
rect 4117 4782 4142 4794
rect 4149 4782 4168 4794
rect 4199 4794 4249 4802
rect 4199 4786 4215 4794
rect 4222 4792 4249 4794
rect 4258 4792 4479 4802
rect 4222 4782 4479 4792
rect 4508 4794 4558 4802
rect 4508 4785 4524 4794
rect 4117 4774 4168 4782
rect 4215 4774 4479 4782
rect 4505 4782 4524 4785
rect 4531 4782 4558 4794
rect 4505 4774 4558 4782
rect 4133 4766 4134 4774
rect 4149 4766 4162 4774
rect 4133 4758 4149 4766
rect 4130 4751 4149 4754
rect 4130 4742 4152 4751
rect 4103 4732 4152 4742
rect 4103 4726 4133 4732
rect 4152 4727 4157 4732
rect 4075 4710 4149 4726
rect 4167 4718 4197 4774
rect 4232 4764 4440 4774
rect 4475 4770 4520 4774
rect 4523 4773 4524 4774
rect 4539 4773 4552 4774
rect 4258 4734 4447 4764
rect 4273 4731 4447 4734
rect 4266 4728 4447 4731
rect 4075 4708 4088 4710
rect 4103 4708 4137 4710
rect 4075 4692 4149 4708
rect 4176 4704 4189 4718
rect 4204 4704 4220 4720
rect 4266 4715 4277 4728
rect 4059 4670 4060 4686
rect 4075 4670 4088 4692
rect 4103 4670 4133 4692
rect 4176 4688 4238 4704
rect 4266 4697 4277 4713
rect 4282 4708 4292 4728
rect 4302 4708 4316 4728
rect 4319 4715 4328 4728
rect 4344 4715 4353 4728
rect 4282 4697 4316 4708
rect 4319 4697 4328 4713
rect 4344 4697 4353 4713
rect 4360 4708 4370 4728
rect 4380 4708 4394 4728
rect 4395 4715 4406 4728
rect 4360 4697 4394 4708
rect 4395 4697 4406 4713
rect 4452 4704 4468 4720
rect 4475 4718 4505 4770
rect 4539 4766 4540 4773
rect 4524 4758 4540 4766
rect 4511 4726 4524 4745
rect 4539 4726 4569 4742
rect 4511 4710 4585 4726
rect 4511 4708 4524 4710
rect 4539 4708 4573 4710
rect 4176 4686 4189 4688
rect 4204 4686 4238 4688
rect 4176 4670 4238 4686
rect 4282 4681 4298 4684
rect 4360 4681 4390 4692
rect 4438 4688 4484 4704
rect 4511 4692 4585 4708
rect 4438 4686 4472 4688
rect 4437 4670 4484 4686
rect 4511 4670 4524 4692
rect 4539 4670 4569 4692
rect 4596 4670 4597 4686
rect 4612 4670 4625 4830
rect 4655 4726 4668 4830
rect 4713 4808 4714 4818
rect 4729 4808 4742 4818
rect 4713 4804 4742 4808
rect 4747 4804 4777 4830
rect 4795 4816 4811 4818
rect 4883 4816 4936 4830
rect 4884 4814 4948 4816
rect 4991 4814 5006 4830
rect 5055 4827 5085 4830
rect 5055 4824 5091 4827
rect 5021 4816 5037 4818
rect 4795 4804 4810 4808
rect 4713 4802 4810 4804
rect 4838 4802 5006 4814
rect 5022 4804 5037 4808
rect 5055 4805 5094 4824
rect 5113 4818 5120 4819
rect 5119 4811 5120 4818
rect 5103 4808 5104 4811
rect 5119 4808 5132 4811
rect 5055 4804 5085 4805
rect 5094 4804 5100 4805
rect 5103 4804 5132 4808
rect 5022 4803 5132 4804
rect 5022 4802 5138 4803
rect 4697 4794 4748 4802
rect 4697 4782 4722 4794
rect 4729 4782 4748 4794
rect 4779 4794 4829 4802
rect 4779 4786 4795 4794
rect 4802 4792 4829 4794
rect 4838 4792 5059 4802
rect 4802 4782 5059 4792
rect 5088 4794 5138 4802
rect 5088 4785 5104 4794
rect 4697 4774 4748 4782
rect 4795 4774 5059 4782
rect 5085 4782 5104 4785
rect 5111 4782 5138 4794
rect 5085 4774 5138 4782
rect 4713 4766 4714 4774
rect 4729 4766 4742 4774
rect 4713 4758 4729 4766
rect 4710 4751 4729 4754
rect 4710 4742 4732 4751
rect 4683 4732 4732 4742
rect 4683 4726 4713 4732
rect 4732 4727 4737 4732
rect 4655 4710 4729 4726
rect 4747 4718 4777 4774
rect 4812 4764 5020 4774
rect 5055 4770 5100 4774
rect 5103 4773 5104 4774
rect 5119 4773 5132 4774
rect 4838 4734 5027 4764
rect 4853 4731 5027 4734
rect 4846 4728 5027 4731
rect 4655 4708 4668 4710
rect 4683 4708 4717 4710
rect 4655 4692 4729 4708
rect 4756 4704 4769 4718
rect 4784 4704 4800 4720
rect 4846 4715 4857 4728
rect 4639 4670 4640 4686
rect 4655 4670 4668 4692
rect 4683 4670 4713 4692
rect 4756 4688 4818 4704
rect 4846 4697 4857 4713
rect 4862 4708 4872 4728
rect 4882 4708 4896 4728
rect 4899 4715 4908 4728
rect 4924 4715 4933 4728
rect 4862 4697 4896 4708
rect 4899 4697 4908 4713
rect 4924 4697 4933 4713
rect 4940 4708 4950 4728
rect 4960 4708 4974 4728
rect 4975 4715 4986 4728
rect 4940 4697 4974 4708
rect 4975 4697 4986 4713
rect 5032 4704 5048 4720
rect 5055 4718 5085 4770
rect 5119 4766 5120 4773
rect 5104 4758 5120 4766
rect 5091 4726 5104 4745
rect 5119 4726 5149 4742
rect 5091 4710 5165 4726
rect 5091 4708 5104 4710
rect 5119 4708 5153 4710
rect 4756 4686 4769 4688
rect 4784 4686 4818 4688
rect 4756 4670 4818 4686
rect 4862 4681 4878 4684
rect 4940 4681 4970 4692
rect 5018 4688 5064 4704
rect 5091 4692 5165 4708
rect 5018 4686 5052 4688
rect 5017 4670 5064 4686
rect 5091 4670 5104 4692
rect 5119 4670 5149 4692
rect 5176 4670 5177 4686
rect 5192 4670 5205 4830
rect 5235 4726 5248 4830
rect 5293 4808 5294 4818
rect 5309 4808 5322 4818
rect 5293 4804 5322 4808
rect 5327 4804 5357 4830
rect 5375 4816 5391 4818
rect 5463 4816 5516 4830
rect 5464 4814 5528 4816
rect 5571 4814 5586 4830
rect 5635 4827 5665 4830
rect 5635 4824 5671 4827
rect 5601 4816 5617 4818
rect 5375 4804 5390 4808
rect 5293 4802 5390 4804
rect 5418 4802 5586 4814
rect 5602 4804 5617 4808
rect 5635 4805 5674 4824
rect 5693 4818 5700 4819
rect 5699 4811 5700 4818
rect 5683 4808 5684 4811
rect 5699 4808 5712 4811
rect 5635 4804 5665 4805
rect 5674 4804 5680 4805
rect 5683 4804 5712 4808
rect 5602 4803 5712 4804
rect 5602 4802 5718 4803
rect 5277 4794 5328 4802
rect 5277 4782 5302 4794
rect 5309 4782 5328 4794
rect 5359 4794 5409 4802
rect 5359 4786 5375 4794
rect 5382 4792 5409 4794
rect 5418 4792 5639 4802
rect 5382 4782 5639 4792
rect 5668 4794 5718 4802
rect 5668 4785 5684 4794
rect 5277 4774 5328 4782
rect 5375 4774 5639 4782
rect 5665 4782 5684 4785
rect 5691 4782 5718 4794
rect 5665 4774 5718 4782
rect 5293 4766 5294 4774
rect 5309 4766 5322 4774
rect 5293 4758 5309 4766
rect 5290 4751 5309 4754
rect 5290 4742 5312 4751
rect 5263 4732 5312 4742
rect 5263 4726 5293 4732
rect 5312 4727 5317 4732
rect 5235 4710 5309 4726
rect 5327 4718 5357 4774
rect 5392 4764 5600 4774
rect 5635 4770 5680 4774
rect 5683 4773 5684 4774
rect 5699 4773 5712 4774
rect 5418 4734 5607 4764
rect 5433 4731 5607 4734
rect 5426 4728 5607 4731
rect 5235 4708 5248 4710
rect 5263 4708 5297 4710
rect 5235 4692 5309 4708
rect 5336 4704 5349 4718
rect 5364 4704 5380 4720
rect 5426 4715 5437 4728
rect 5219 4670 5220 4686
rect 5235 4670 5248 4692
rect 5263 4670 5293 4692
rect 5336 4688 5398 4704
rect 5426 4697 5437 4713
rect 5442 4708 5452 4728
rect 5462 4708 5476 4728
rect 5479 4715 5488 4728
rect 5504 4715 5513 4728
rect 5442 4697 5476 4708
rect 5479 4697 5488 4713
rect 5504 4697 5513 4713
rect 5520 4708 5530 4728
rect 5540 4708 5554 4728
rect 5555 4715 5566 4728
rect 5520 4697 5554 4708
rect 5555 4697 5566 4713
rect 5612 4704 5628 4720
rect 5635 4718 5665 4770
rect 5699 4766 5700 4773
rect 5684 4758 5700 4766
rect 5671 4726 5684 4745
rect 5699 4726 5729 4742
rect 5671 4710 5745 4726
rect 5671 4708 5684 4710
rect 5699 4708 5733 4710
rect 5336 4686 5349 4688
rect 5364 4686 5398 4688
rect 5336 4670 5398 4686
rect 5442 4681 5458 4684
rect 5520 4681 5550 4692
rect 5598 4688 5644 4704
rect 5671 4692 5745 4708
rect 5598 4686 5632 4688
rect 5597 4670 5644 4686
rect 5671 4670 5684 4692
rect 5699 4670 5729 4692
rect 5756 4670 5757 4686
rect 5772 4670 5785 4830
rect 5815 4726 5828 4830
rect 5873 4808 5874 4818
rect 5889 4808 5902 4818
rect 5873 4804 5902 4808
rect 5907 4804 5937 4830
rect 5955 4816 5971 4818
rect 6043 4816 6096 4830
rect 6044 4814 6108 4816
rect 6151 4814 6166 4830
rect 6215 4827 6245 4830
rect 6215 4824 6251 4827
rect 6181 4816 6197 4818
rect 5955 4804 5970 4808
rect 5873 4802 5970 4804
rect 5998 4802 6166 4814
rect 6182 4804 6197 4808
rect 6215 4805 6254 4824
rect 6273 4818 6280 4819
rect 6279 4811 6280 4818
rect 6263 4808 6264 4811
rect 6279 4808 6292 4811
rect 6215 4804 6245 4805
rect 6254 4804 6260 4805
rect 6263 4804 6292 4808
rect 6182 4803 6292 4804
rect 6182 4802 6298 4803
rect 5857 4794 5908 4802
rect 5857 4782 5882 4794
rect 5889 4782 5908 4794
rect 5939 4794 5989 4802
rect 5939 4786 5955 4794
rect 5962 4792 5989 4794
rect 5998 4792 6219 4802
rect 5962 4782 6219 4792
rect 6248 4794 6298 4802
rect 6248 4785 6264 4794
rect 5857 4774 5908 4782
rect 5955 4774 6219 4782
rect 6245 4782 6264 4785
rect 6271 4782 6298 4794
rect 6245 4774 6298 4782
rect 5873 4766 5874 4774
rect 5889 4766 5902 4774
rect 5873 4758 5889 4766
rect 5870 4751 5889 4754
rect 5870 4742 5892 4751
rect 5843 4732 5892 4742
rect 5843 4726 5873 4732
rect 5892 4727 5897 4732
rect 5815 4710 5889 4726
rect 5907 4718 5937 4774
rect 5972 4764 6180 4774
rect 6215 4770 6260 4774
rect 6263 4773 6264 4774
rect 6279 4773 6292 4774
rect 5998 4734 6187 4764
rect 6013 4731 6187 4734
rect 6006 4728 6187 4731
rect 5815 4708 5828 4710
rect 5843 4708 5877 4710
rect 5815 4692 5889 4708
rect 5916 4704 5929 4718
rect 5944 4704 5960 4720
rect 6006 4715 6017 4728
rect 5799 4670 5800 4686
rect 5815 4670 5828 4692
rect 5843 4670 5873 4692
rect 5916 4688 5978 4704
rect 6006 4697 6017 4713
rect 6022 4708 6032 4728
rect 6042 4708 6056 4728
rect 6059 4715 6068 4728
rect 6084 4715 6093 4728
rect 6022 4697 6056 4708
rect 6059 4697 6068 4713
rect 6084 4697 6093 4713
rect 6100 4708 6110 4728
rect 6120 4708 6134 4728
rect 6135 4715 6146 4728
rect 6100 4697 6134 4708
rect 6135 4697 6146 4713
rect 6192 4704 6208 4720
rect 6215 4718 6245 4770
rect 6279 4766 6280 4773
rect 6264 4758 6280 4766
rect 6251 4726 6264 4745
rect 6279 4726 6309 4742
rect 6251 4710 6325 4726
rect 6251 4708 6264 4710
rect 6279 4708 6313 4710
rect 5916 4686 5929 4688
rect 5944 4686 5978 4688
rect 5916 4670 5978 4686
rect 6022 4681 6038 4684
rect 6100 4681 6130 4692
rect 6178 4688 6224 4704
rect 6251 4692 6325 4708
rect 6178 4686 6212 4688
rect 6177 4670 6224 4686
rect 6251 4670 6264 4692
rect 6279 4670 6309 4692
rect 6336 4670 6337 4686
rect 6352 4670 6365 4830
rect 6395 4726 6408 4830
rect 6453 4808 6454 4818
rect 6469 4808 6482 4818
rect 6453 4804 6482 4808
rect 6487 4804 6517 4830
rect 6535 4816 6551 4818
rect 6623 4816 6676 4830
rect 6624 4814 6688 4816
rect 6731 4814 6746 4830
rect 6795 4827 6825 4830
rect 6795 4824 6831 4827
rect 6761 4816 6777 4818
rect 6535 4804 6550 4808
rect 6453 4802 6550 4804
rect 6578 4802 6746 4814
rect 6762 4804 6777 4808
rect 6795 4805 6834 4824
rect 6853 4818 6860 4819
rect 6859 4811 6860 4818
rect 6843 4808 6844 4811
rect 6859 4808 6872 4811
rect 6795 4804 6825 4805
rect 6834 4804 6840 4805
rect 6843 4804 6872 4808
rect 6762 4803 6872 4804
rect 6762 4802 6878 4803
rect 6437 4794 6488 4802
rect 6437 4782 6462 4794
rect 6469 4782 6488 4794
rect 6519 4794 6569 4802
rect 6519 4786 6535 4794
rect 6542 4792 6569 4794
rect 6578 4792 6799 4802
rect 6542 4782 6799 4792
rect 6828 4794 6878 4802
rect 6828 4785 6844 4794
rect 6437 4774 6488 4782
rect 6535 4774 6799 4782
rect 6825 4782 6844 4785
rect 6851 4782 6878 4794
rect 6825 4774 6878 4782
rect 6453 4766 6454 4774
rect 6469 4766 6482 4774
rect 6453 4758 6469 4766
rect 6450 4751 6469 4754
rect 6450 4742 6472 4751
rect 6423 4732 6472 4742
rect 6423 4726 6453 4732
rect 6472 4727 6477 4732
rect 6395 4710 6469 4726
rect 6487 4718 6517 4774
rect 6552 4764 6760 4774
rect 6795 4770 6840 4774
rect 6843 4773 6844 4774
rect 6859 4773 6872 4774
rect 6578 4734 6767 4764
rect 6593 4731 6767 4734
rect 6586 4728 6767 4731
rect 6395 4708 6408 4710
rect 6423 4708 6457 4710
rect 6395 4692 6469 4708
rect 6496 4704 6509 4718
rect 6524 4704 6540 4720
rect 6586 4715 6597 4728
rect 6379 4670 6380 4686
rect 6395 4670 6408 4692
rect 6423 4670 6453 4692
rect 6496 4688 6558 4704
rect 6586 4697 6597 4713
rect 6602 4708 6612 4728
rect 6622 4708 6636 4728
rect 6639 4715 6648 4728
rect 6664 4715 6673 4728
rect 6602 4697 6636 4708
rect 6639 4697 6648 4713
rect 6664 4697 6673 4713
rect 6680 4708 6690 4728
rect 6700 4708 6714 4728
rect 6715 4715 6726 4728
rect 6680 4697 6714 4708
rect 6715 4697 6726 4713
rect 6772 4704 6788 4720
rect 6795 4718 6825 4770
rect 6859 4766 6860 4773
rect 6844 4758 6860 4766
rect 6831 4726 6844 4745
rect 6859 4726 6889 4742
rect 6831 4710 6905 4726
rect 6831 4708 6844 4710
rect 6859 4708 6893 4710
rect 6496 4686 6509 4688
rect 6524 4686 6558 4688
rect 6496 4670 6558 4686
rect 6602 4681 6618 4684
rect 6680 4681 6710 4692
rect 6758 4688 6804 4704
rect 6831 4692 6905 4708
rect 6758 4686 6792 4688
rect 6757 4670 6804 4686
rect 6831 4670 6844 4692
rect 6859 4670 6889 4692
rect 6916 4670 6917 4686
rect 6932 4670 6945 4830
rect 6975 4726 6988 4830
rect 7033 4808 7034 4818
rect 7049 4808 7062 4818
rect 7033 4804 7062 4808
rect 7067 4804 7097 4830
rect 7115 4816 7131 4818
rect 7203 4816 7256 4830
rect 7204 4814 7268 4816
rect 7311 4814 7326 4830
rect 7375 4827 7405 4830
rect 7375 4824 7411 4827
rect 7341 4816 7357 4818
rect 7115 4804 7130 4808
rect 7033 4802 7130 4804
rect 7158 4802 7326 4814
rect 7342 4804 7357 4808
rect 7375 4805 7414 4824
rect 7433 4818 7440 4819
rect 7439 4811 7440 4818
rect 7423 4808 7424 4811
rect 7439 4808 7452 4811
rect 7375 4804 7405 4805
rect 7414 4804 7420 4805
rect 7423 4804 7452 4808
rect 7342 4803 7452 4804
rect 7342 4802 7458 4803
rect 7017 4794 7068 4802
rect 7017 4782 7042 4794
rect 7049 4782 7068 4794
rect 7099 4794 7149 4802
rect 7099 4786 7115 4794
rect 7122 4792 7149 4794
rect 7158 4792 7379 4802
rect 7122 4782 7379 4792
rect 7408 4794 7458 4802
rect 7408 4785 7424 4794
rect 7017 4774 7068 4782
rect 7115 4774 7379 4782
rect 7405 4782 7424 4785
rect 7431 4782 7458 4794
rect 7405 4774 7458 4782
rect 7033 4766 7034 4774
rect 7049 4766 7062 4774
rect 7033 4758 7049 4766
rect 7030 4751 7049 4754
rect 7030 4742 7052 4751
rect 7003 4732 7052 4742
rect 7003 4726 7033 4732
rect 7052 4727 7057 4732
rect 6975 4710 7049 4726
rect 7067 4718 7097 4774
rect 7132 4764 7340 4774
rect 7375 4770 7420 4774
rect 7423 4773 7424 4774
rect 7439 4773 7452 4774
rect 7158 4734 7347 4764
rect 7173 4731 7347 4734
rect 7166 4728 7347 4731
rect 6975 4708 6988 4710
rect 7003 4708 7037 4710
rect 6975 4692 7049 4708
rect 7076 4704 7089 4718
rect 7104 4704 7120 4720
rect 7166 4715 7177 4728
rect 6959 4670 6960 4686
rect 6975 4670 6988 4692
rect 7003 4670 7033 4692
rect 7076 4688 7138 4704
rect 7166 4697 7177 4713
rect 7182 4708 7192 4728
rect 7202 4708 7216 4728
rect 7219 4715 7228 4728
rect 7244 4715 7253 4728
rect 7182 4697 7216 4708
rect 7219 4697 7228 4713
rect 7244 4697 7253 4713
rect 7260 4708 7270 4728
rect 7280 4708 7294 4728
rect 7295 4715 7306 4728
rect 7260 4697 7294 4708
rect 7295 4697 7306 4713
rect 7352 4704 7368 4720
rect 7375 4718 7405 4770
rect 7439 4766 7440 4773
rect 7424 4758 7440 4766
rect 7411 4726 7424 4745
rect 7439 4726 7469 4742
rect 7411 4710 7485 4726
rect 7411 4708 7424 4710
rect 7439 4708 7473 4710
rect 7076 4686 7089 4688
rect 7104 4686 7138 4688
rect 7076 4670 7138 4686
rect 7182 4681 7198 4684
rect 7260 4681 7290 4692
rect 7338 4688 7384 4704
rect 7411 4692 7485 4708
rect 7338 4686 7372 4688
rect 7337 4670 7384 4686
rect 7411 4670 7424 4692
rect 7439 4670 7469 4692
rect 7496 4670 7497 4686
rect 7512 4670 7525 4830
rect 7555 4726 7568 4830
rect 7613 4808 7614 4818
rect 7629 4808 7642 4818
rect 7613 4804 7642 4808
rect 7647 4804 7677 4830
rect 7695 4816 7711 4818
rect 7783 4816 7836 4830
rect 7784 4814 7848 4816
rect 7891 4814 7906 4830
rect 7955 4827 7985 4830
rect 7955 4824 7991 4827
rect 7921 4816 7937 4818
rect 7695 4804 7710 4808
rect 7613 4802 7710 4804
rect 7738 4802 7906 4814
rect 7922 4804 7937 4808
rect 7955 4805 7994 4824
rect 8013 4818 8020 4819
rect 8019 4811 8020 4818
rect 8003 4808 8004 4811
rect 8019 4808 8032 4811
rect 7955 4804 7985 4805
rect 7994 4804 8000 4805
rect 8003 4804 8032 4808
rect 7922 4803 8032 4804
rect 7922 4802 8038 4803
rect 7597 4794 7648 4802
rect 7597 4782 7622 4794
rect 7629 4782 7648 4794
rect 7679 4794 7729 4802
rect 7679 4786 7695 4794
rect 7702 4792 7729 4794
rect 7738 4792 7959 4802
rect 7702 4782 7959 4792
rect 7988 4794 8038 4802
rect 7988 4785 8004 4794
rect 7597 4774 7648 4782
rect 7695 4774 7959 4782
rect 7985 4782 8004 4785
rect 8011 4782 8038 4794
rect 7985 4774 8038 4782
rect 7613 4766 7614 4774
rect 7629 4766 7642 4774
rect 7613 4758 7629 4766
rect 7610 4751 7629 4754
rect 7610 4742 7632 4751
rect 7583 4732 7632 4742
rect 7583 4726 7613 4732
rect 7632 4727 7637 4732
rect 7555 4710 7629 4726
rect 7647 4718 7677 4774
rect 7712 4764 7920 4774
rect 7955 4770 8000 4774
rect 8003 4773 8004 4774
rect 8019 4773 8032 4774
rect 7738 4734 7927 4764
rect 7753 4731 7927 4734
rect 7746 4728 7927 4731
rect 7555 4708 7568 4710
rect 7583 4708 7617 4710
rect 7555 4692 7629 4708
rect 7656 4704 7669 4718
rect 7684 4704 7700 4720
rect 7746 4715 7757 4728
rect 7539 4670 7540 4686
rect 7555 4670 7568 4692
rect 7583 4670 7613 4692
rect 7656 4688 7718 4704
rect 7746 4697 7757 4713
rect 7762 4708 7772 4728
rect 7782 4708 7796 4728
rect 7799 4715 7808 4728
rect 7824 4715 7833 4728
rect 7762 4697 7796 4708
rect 7799 4697 7808 4713
rect 7824 4697 7833 4713
rect 7840 4708 7850 4728
rect 7860 4708 7874 4728
rect 7875 4715 7886 4728
rect 7840 4697 7874 4708
rect 7875 4697 7886 4713
rect 7932 4704 7948 4720
rect 7955 4718 7985 4770
rect 8019 4766 8020 4773
rect 8004 4758 8020 4766
rect 7991 4726 8004 4745
rect 8019 4726 8049 4742
rect 7991 4710 8065 4726
rect 7991 4708 8004 4710
rect 8019 4708 8053 4710
rect 7656 4686 7669 4688
rect 7684 4686 7718 4688
rect 7656 4670 7718 4686
rect 7762 4681 7778 4684
rect 7840 4681 7870 4692
rect 7918 4688 7964 4704
rect 7991 4692 8065 4708
rect 7918 4686 7952 4688
rect 7917 4670 7964 4686
rect 7991 4670 8004 4692
rect 8019 4670 8049 4692
rect 8076 4670 8077 4686
rect 8092 4670 8105 4830
rect 8135 4726 8148 4830
rect 8193 4808 8194 4818
rect 8209 4808 8222 4818
rect 8193 4804 8222 4808
rect 8227 4804 8257 4830
rect 8275 4816 8291 4818
rect 8363 4816 8416 4830
rect 8364 4814 8428 4816
rect 8471 4814 8486 4830
rect 8535 4827 8565 4830
rect 8535 4824 8571 4827
rect 8501 4816 8517 4818
rect 8275 4804 8290 4808
rect 8193 4802 8290 4804
rect 8318 4802 8486 4814
rect 8502 4804 8517 4808
rect 8535 4805 8574 4824
rect 8593 4818 8600 4819
rect 8599 4811 8600 4818
rect 8583 4808 8584 4811
rect 8599 4808 8612 4811
rect 8535 4804 8565 4805
rect 8574 4804 8580 4805
rect 8583 4804 8612 4808
rect 8502 4803 8612 4804
rect 8502 4802 8618 4803
rect 8177 4794 8228 4802
rect 8177 4782 8202 4794
rect 8209 4782 8228 4794
rect 8259 4794 8309 4802
rect 8259 4786 8275 4794
rect 8282 4792 8309 4794
rect 8318 4792 8539 4802
rect 8282 4782 8539 4792
rect 8568 4794 8618 4802
rect 8568 4785 8584 4794
rect 8177 4774 8228 4782
rect 8275 4774 8539 4782
rect 8565 4782 8584 4785
rect 8591 4782 8618 4794
rect 8565 4774 8618 4782
rect 8193 4766 8194 4774
rect 8209 4766 8222 4774
rect 8193 4758 8209 4766
rect 8190 4751 8209 4754
rect 8190 4742 8212 4751
rect 8163 4732 8212 4742
rect 8163 4726 8193 4732
rect 8212 4727 8217 4732
rect 8135 4710 8209 4726
rect 8227 4718 8257 4774
rect 8292 4764 8500 4774
rect 8535 4770 8580 4774
rect 8583 4773 8584 4774
rect 8599 4773 8612 4774
rect 8318 4734 8507 4764
rect 8333 4731 8507 4734
rect 8326 4728 8507 4731
rect 8135 4708 8148 4710
rect 8163 4708 8197 4710
rect 8135 4692 8209 4708
rect 8236 4704 8249 4718
rect 8264 4704 8280 4720
rect 8326 4715 8337 4728
rect 8119 4670 8120 4686
rect 8135 4670 8148 4692
rect 8163 4670 8193 4692
rect 8236 4688 8298 4704
rect 8326 4697 8337 4713
rect 8342 4708 8352 4728
rect 8362 4708 8376 4728
rect 8379 4715 8388 4728
rect 8404 4715 8413 4728
rect 8342 4697 8376 4708
rect 8379 4697 8388 4713
rect 8404 4697 8413 4713
rect 8420 4708 8430 4728
rect 8440 4708 8454 4728
rect 8455 4715 8466 4728
rect 8420 4697 8454 4708
rect 8455 4697 8466 4713
rect 8512 4704 8528 4720
rect 8535 4718 8565 4770
rect 8599 4766 8600 4773
rect 8584 4758 8600 4766
rect 8571 4726 8584 4745
rect 8599 4726 8629 4742
rect 8571 4710 8645 4726
rect 8571 4708 8584 4710
rect 8599 4708 8633 4710
rect 8236 4686 8249 4688
rect 8264 4686 8298 4688
rect 8236 4670 8298 4686
rect 8342 4681 8358 4684
rect 8420 4681 8450 4692
rect 8498 4688 8544 4704
rect 8571 4692 8645 4708
rect 8498 4686 8532 4688
rect 8497 4670 8544 4686
rect 8571 4670 8584 4692
rect 8599 4670 8629 4692
rect 8656 4670 8657 4686
rect 8672 4670 8685 4830
rect 8715 4726 8728 4830
rect 8773 4808 8774 4818
rect 8789 4808 8802 4818
rect 8773 4804 8802 4808
rect 8807 4804 8837 4830
rect 8855 4816 8871 4818
rect 8943 4816 8996 4830
rect 8944 4814 9008 4816
rect 9051 4814 9066 4830
rect 9115 4827 9145 4830
rect 9115 4824 9151 4827
rect 9081 4816 9097 4818
rect 8855 4804 8870 4808
rect 8773 4802 8870 4804
rect 8898 4802 9066 4814
rect 9082 4804 9097 4808
rect 9115 4805 9154 4824
rect 9173 4818 9180 4819
rect 9179 4811 9180 4818
rect 9163 4808 9164 4811
rect 9179 4808 9192 4811
rect 9115 4804 9145 4805
rect 9154 4804 9160 4805
rect 9163 4804 9192 4808
rect 9082 4803 9192 4804
rect 9082 4802 9198 4803
rect 8757 4794 8808 4802
rect 8757 4782 8782 4794
rect 8789 4782 8808 4794
rect 8839 4794 8889 4802
rect 8839 4786 8855 4794
rect 8862 4792 8889 4794
rect 8898 4792 9119 4802
rect 8862 4782 9119 4792
rect 9148 4794 9198 4802
rect 9148 4785 9164 4794
rect 8757 4774 8808 4782
rect 8855 4774 9119 4782
rect 9145 4782 9164 4785
rect 9171 4782 9198 4794
rect 9145 4774 9198 4782
rect 8773 4766 8774 4774
rect 8789 4766 8802 4774
rect 8773 4758 8789 4766
rect 8770 4751 8789 4754
rect 8770 4742 8792 4751
rect 8743 4732 8792 4742
rect 8743 4726 8773 4732
rect 8792 4727 8797 4732
rect 8715 4710 8789 4726
rect 8807 4718 8837 4774
rect 8872 4764 9080 4774
rect 9115 4770 9160 4774
rect 9163 4773 9164 4774
rect 9179 4773 9192 4774
rect 8898 4734 9087 4764
rect 8913 4731 9087 4734
rect 8906 4728 9087 4731
rect 8715 4708 8728 4710
rect 8743 4708 8777 4710
rect 8715 4692 8789 4708
rect 8816 4704 8829 4718
rect 8844 4704 8860 4720
rect 8906 4715 8917 4728
rect 8699 4670 8700 4686
rect 8715 4670 8728 4692
rect 8743 4670 8773 4692
rect 8816 4688 8878 4704
rect 8906 4697 8917 4713
rect 8922 4708 8932 4728
rect 8942 4708 8956 4728
rect 8959 4715 8968 4728
rect 8984 4715 8993 4728
rect 8922 4697 8956 4708
rect 8959 4697 8968 4713
rect 8984 4697 8993 4713
rect 9000 4708 9010 4728
rect 9020 4708 9034 4728
rect 9035 4715 9046 4728
rect 9000 4697 9034 4708
rect 9035 4697 9046 4713
rect 9092 4704 9108 4720
rect 9115 4718 9145 4770
rect 9179 4766 9180 4773
rect 9164 4758 9180 4766
rect 9151 4726 9164 4745
rect 9179 4726 9209 4742
rect 9151 4710 9225 4726
rect 9151 4708 9164 4710
rect 9179 4708 9213 4710
rect 8816 4686 8829 4688
rect 8844 4686 8878 4688
rect 8816 4670 8878 4686
rect 8922 4681 8938 4684
rect 9000 4681 9030 4692
rect 9078 4688 9124 4704
rect 9151 4692 9225 4708
rect 9078 4686 9112 4688
rect 9077 4670 9124 4686
rect 9151 4670 9164 4692
rect 9179 4670 9209 4692
rect 9236 4670 9237 4686
rect 9252 4670 9265 4830
rect -7 4662 34 4670
rect -7 4636 8 4662
rect 15 4636 34 4662
rect 98 4658 160 4670
rect 172 4658 247 4670
rect 305 4658 380 4670
rect 392 4658 423 4670
rect 429 4658 464 4670
rect 98 4656 260 4658
rect -7 4628 34 4636
rect 116 4632 129 4656
rect 144 4654 159 4656
rect -1 4618 0 4628
rect 15 4618 28 4628
rect 43 4618 73 4632
rect 116 4618 159 4632
rect 183 4629 190 4636
rect 193 4632 260 4656
rect 292 4656 464 4658
rect 262 4634 290 4638
rect 292 4634 372 4656
rect 393 4654 408 4656
rect 262 4632 372 4634
rect 193 4628 372 4632
rect 166 4618 196 4628
rect 198 4618 351 4628
rect 359 4618 389 4628
rect 393 4618 423 4632
rect 451 4618 464 4656
rect 536 4662 571 4670
rect 536 4636 537 4662
rect 544 4636 571 4662
rect 479 4618 509 4632
rect 536 4628 571 4636
rect 573 4662 614 4670
rect 573 4636 588 4662
rect 595 4636 614 4662
rect 678 4658 740 4670
rect 752 4658 827 4670
rect 885 4658 960 4670
rect 972 4658 1003 4670
rect 1009 4658 1044 4670
rect 678 4656 840 4658
rect 573 4628 614 4636
rect 696 4632 709 4656
rect 724 4654 739 4656
rect 536 4618 537 4628
rect 552 4618 565 4628
rect 579 4618 580 4628
rect 595 4618 608 4628
rect 623 4618 653 4632
rect 696 4618 739 4632
rect 763 4629 770 4636
rect 773 4632 840 4656
rect 872 4656 1044 4658
rect 842 4634 870 4638
rect 872 4634 952 4656
rect 973 4654 988 4656
rect 842 4632 952 4634
rect 773 4628 952 4632
rect 746 4618 776 4628
rect 778 4618 931 4628
rect 939 4618 969 4628
rect 973 4618 1003 4632
rect 1031 4618 1044 4656
rect 1116 4662 1151 4670
rect 1116 4636 1117 4662
rect 1124 4636 1151 4662
rect 1059 4618 1089 4632
rect 1116 4628 1151 4636
rect 1153 4662 1194 4670
rect 1153 4636 1168 4662
rect 1175 4636 1194 4662
rect 1258 4658 1320 4670
rect 1332 4658 1407 4670
rect 1465 4658 1540 4670
rect 1552 4658 1583 4670
rect 1589 4658 1624 4670
rect 1258 4656 1420 4658
rect 1153 4628 1194 4636
rect 1276 4632 1289 4656
rect 1304 4654 1319 4656
rect 1116 4618 1117 4628
rect 1132 4618 1145 4628
rect 1159 4618 1160 4628
rect 1175 4618 1188 4628
rect 1203 4618 1233 4632
rect 1276 4618 1319 4632
rect 1343 4629 1350 4636
rect 1353 4632 1420 4656
rect 1452 4656 1624 4658
rect 1422 4634 1450 4638
rect 1452 4634 1532 4656
rect 1553 4654 1568 4656
rect 1422 4632 1532 4634
rect 1353 4628 1532 4632
rect 1326 4618 1356 4628
rect 1358 4618 1511 4628
rect 1519 4618 1549 4628
rect 1553 4618 1583 4632
rect 1611 4618 1624 4656
rect 1696 4662 1731 4670
rect 1696 4636 1697 4662
rect 1704 4636 1731 4662
rect 1639 4618 1669 4632
rect 1696 4628 1731 4636
rect 1733 4662 1774 4670
rect 1733 4636 1748 4662
rect 1755 4636 1774 4662
rect 1838 4658 1900 4670
rect 1912 4658 1987 4670
rect 2045 4658 2120 4670
rect 2132 4658 2163 4670
rect 2169 4658 2204 4670
rect 1838 4656 2000 4658
rect 1733 4628 1774 4636
rect 1856 4632 1869 4656
rect 1884 4654 1899 4656
rect 1696 4618 1697 4628
rect 1712 4618 1725 4628
rect 1739 4618 1740 4628
rect 1755 4618 1768 4628
rect 1783 4618 1813 4632
rect 1856 4618 1899 4632
rect 1923 4629 1930 4636
rect 1933 4632 2000 4656
rect 2032 4656 2204 4658
rect 2002 4634 2030 4638
rect 2032 4634 2112 4656
rect 2133 4654 2148 4656
rect 2002 4632 2112 4634
rect 1933 4628 2112 4632
rect 1906 4618 1936 4628
rect 1938 4618 2091 4628
rect 2099 4618 2129 4628
rect 2133 4618 2163 4632
rect 2191 4618 2204 4656
rect 2276 4662 2311 4670
rect 2276 4636 2277 4662
rect 2284 4636 2311 4662
rect 2219 4618 2249 4632
rect 2276 4628 2311 4636
rect 2313 4662 2354 4670
rect 2313 4636 2328 4662
rect 2335 4636 2354 4662
rect 2418 4658 2480 4670
rect 2492 4658 2567 4670
rect 2625 4658 2700 4670
rect 2712 4658 2743 4670
rect 2749 4658 2784 4670
rect 2418 4656 2580 4658
rect 2313 4628 2354 4636
rect 2436 4632 2449 4656
rect 2464 4654 2479 4656
rect 2276 4618 2277 4628
rect 2292 4618 2305 4628
rect 2319 4618 2320 4628
rect 2335 4618 2348 4628
rect 2363 4618 2393 4632
rect 2436 4618 2479 4632
rect 2503 4629 2510 4636
rect 2513 4632 2580 4656
rect 2612 4656 2784 4658
rect 2582 4634 2610 4638
rect 2612 4634 2692 4656
rect 2713 4654 2728 4656
rect 2582 4632 2692 4634
rect 2513 4628 2692 4632
rect 2486 4618 2516 4628
rect 2518 4618 2671 4628
rect 2679 4618 2709 4628
rect 2713 4618 2743 4632
rect 2771 4618 2784 4656
rect 2856 4662 2891 4670
rect 2856 4636 2857 4662
rect 2864 4636 2891 4662
rect 2799 4618 2829 4632
rect 2856 4628 2891 4636
rect 2893 4662 2934 4670
rect 2893 4636 2908 4662
rect 2915 4636 2934 4662
rect 2998 4658 3060 4670
rect 3072 4658 3147 4670
rect 3205 4658 3280 4670
rect 3292 4658 3323 4670
rect 3329 4658 3364 4670
rect 2998 4656 3160 4658
rect 2893 4628 2934 4636
rect 3016 4632 3029 4656
rect 3044 4654 3059 4656
rect 2856 4618 2857 4628
rect 2872 4618 2885 4628
rect 2899 4618 2900 4628
rect 2915 4618 2928 4628
rect 2943 4618 2973 4632
rect 3016 4618 3059 4632
rect 3083 4629 3090 4636
rect 3093 4632 3160 4656
rect 3192 4656 3364 4658
rect 3162 4634 3190 4638
rect 3192 4634 3272 4656
rect 3293 4654 3308 4656
rect 3162 4632 3272 4634
rect 3093 4628 3272 4632
rect 3066 4618 3096 4628
rect 3098 4618 3251 4628
rect 3259 4618 3289 4628
rect 3293 4618 3323 4632
rect 3351 4618 3364 4656
rect 3436 4662 3471 4670
rect 3436 4636 3437 4662
rect 3444 4636 3471 4662
rect 3379 4618 3409 4632
rect 3436 4628 3471 4636
rect 3473 4662 3514 4670
rect 3473 4636 3488 4662
rect 3495 4636 3514 4662
rect 3578 4658 3640 4670
rect 3652 4658 3727 4670
rect 3785 4658 3860 4670
rect 3872 4658 3903 4670
rect 3909 4658 3944 4670
rect 3578 4656 3740 4658
rect 3473 4628 3514 4636
rect 3596 4632 3609 4656
rect 3624 4654 3639 4656
rect 3436 4618 3437 4628
rect 3452 4618 3465 4628
rect 3479 4618 3480 4628
rect 3495 4618 3508 4628
rect 3523 4618 3553 4632
rect 3596 4618 3639 4632
rect 3663 4629 3670 4636
rect 3673 4632 3740 4656
rect 3772 4656 3944 4658
rect 3742 4634 3770 4638
rect 3772 4634 3852 4656
rect 3873 4654 3888 4656
rect 3742 4632 3852 4634
rect 3673 4628 3852 4632
rect 3646 4618 3676 4628
rect 3678 4618 3831 4628
rect 3839 4618 3869 4628
rect 3873 4618 3903 4632
rect 3931 4618 3944 4656
rect 4016 4662 4051 4670
rect 4016 4636 4017 4662
rect 4024 4636 4051 4662
rect 3959 4618 3989 4632
rect 4016 4628 4051 4636
rect 4053 4662 4094 4670
rect 4053 4636 4068 4662
rect 4075 4636 4094 4662
rect 4158 4658 4220 4670
rect 4232 4658 4307 4670
rect 4365 4658 4440 4670
rect 4452 4658 4483 4670
rect 4489 4658 4524 4670
rect 4158 4656 4320 4658
rect 4053 4628 4094 4636
rect 4176 4632 4189 4656
rect 4204 4654 4219 4656
rect 4016 4618 4017 4628
rect 4032 4618 4045 4628
rect 4059 4618 4060 4628
rect 4075 4618 4088 4628
rect 4103 4618 4133 4632
rect 4176 4618 4219 4632
rect 4243 4629 4250 4636
rect 4253 4632 4320 4656
rect 4352 4656 4524 4658
rect 4322 4634 4350 4638
rect 4352 4634 4432 4656
rect 4453 4654 4468 4656
rect 4322 4632 4432 4634
rect 4253 4628 4432 4632
rect 4226 4618 4256 4628
rect 4258 4618 4411 4628
rect 4419 4618 4449 4628
rect 4453 4618 4483 4632
rect 4511 4618 4524 4656
rect 4596 4662 4631 4670
rect 4596 4636 4597 4662
rect 4604 4636 4631 4662
rect 4539 4618 4569 4632
rect 4596 4628 4631 4636
rect 4633 4662 4674 4670
rect 4633 4636 4648 4662
rect 4655 4636 4674 4662
rect 4738 4658 4800 4670
rect 4812 4658 4887 4670
rect 4945 4658 5020 4670
rect 5032 4658 5063 4670
rect 5069 4658 5104 4670
rect 4738 4656 4900 4658
rect 4633 4628 4674 4636
rect 4756 4632 4769 4656
rect 4784 4654 4799 4656
rect 4596 4618 4597 4628
rect 4612 4618 4625 4628
rect 4639 4618 4640 4628
rect 4655 4618 4668 4628
rect 4683 4618 4713 4632
rect 4756 4618 4799 4632
rect 4823 4629 4830 4636
rect 4833 4632 4900 4656
rect 4932 4656 5104 4658
rect 4902 4634 4930 4638
rect 4932 4634 5012 4656
rect 5033 4654 5048 4656
rect 4902 4632 5012 4634
rect 4833 4628 5012 4632
rect 4806 4618 4836 4628
rect 4838 4618 4991 4628
rect 4999 4618 5029 4628
rect 5033 4618 5063 4632
rect 5091 4618 5104 4656
rect 5176 4662 5211 4670
rect 5176 4636 5177 4662
rect 5184 4636 5211 4662
rect 5119 4618 5149 4632
rect 5176 4628 5211 4636
rect 5213 4662 5254 4670
rect 5213 4636 5228 4662
rect 5235 4636 5254 4662
rect 5318 4658 5380 4670
rect 5392 4658 5467 4670
rect 5525 4658 5600 4670
rect 5612 4658 5643 4670
rect 5649 4658 5684 4670
rect 5318 4656 5480 4658
rect 5213 4628 5254 4636
rect 5336 4632 5349 4656
rect 5364 4654 5379 4656
rect 5176 4618 5177 4628
rect 5192 4618 5205 4628
rect 5219 4618 5220 4628
rect 5235 4618 5248 4628
rect 5263 4618 5293 4632
rect 5336 4618 5379 4632
rect 5403 4629 5410 4636
rect 5413 4632 5480 4656
rect 5512 4656 5684 4658
rect 5482 4634 5510 4638
rect 5512 4634 5592 4656
rect 5613 4654 5628 4656
rect 5482 4632 5592 4634
rect 5413 4628 5592 4632
rect 5386 4618 5416 4628
rect 5418 4618 5571 4628
rect 5579 4618 5609 4628
rect 5613 4618 5643 4632
rect 5671 4618 5684 4656
rect 5756 4662 5791 4670
rect 5756 4636 5757 4662
rect 5764 4636 5791 4662
rect 5699 4618 5729 4632
rect 5756 4628 5791 4636
rect 5793 4662 5834 4670
rect 5793 4636 5808 4662
rect 5815 4636 5834 4662
rect 5898 4658 5960 4670
rect 5972 4658 6047 4670
rect 6105 4658 6180 4670
rect 6192 4658 6223 4670
rect 6229 4658 6264 4670
rect 5898 4656 6060 4658
rect 5793 4628 5834 4636
rect 5916 4632 5929 4656
rect 5944 4654 5959 4656
rect 5756 4618 5757 4628
rect 5772 4618 5785 4628
rect 5799 4618 5800 4628
rect 5815 4618 5828 4628
rect 5843 4618 5873 4632
rect 5916 4618 5959 4632
rect 5983 4629 5990 4636
rect 5993 4632 6060 4656
rect 6092 4656 6264 4658
rect 6062 4634 6090 4638
rect 6092 4634 6172 4656
rect 6193 4654 6208 4656
rect 6062 4632 6172 4634
rect 5993 4628 6172 4632
rect 5966 4618 5996 4628
rect 5998 4618 6151 4628
rect 6159 4618 6189 4628
rect 6193 4618 6223 4632
rect 6251 4618 6264 4656
rect 6336 4662 6371 4670
rect 6336 4636 6337 4662
rect 6344 4636 6371 4662
rect 6279 4618 6309 4632
rect 6336 4628 6371 4636
rect 6373 4662 6414 4670
rect 6373 4636 6388 4662
rect 6395 4636 6414 4662
rect 6478 4658 6540 4670
rect 6552 4658 6627 4670
rect 6685 4658 6760 4670
rect 6772 4658 6803 4670
rect 6809 4658 6844 4670
rect 6478 4656 6640 4658
rect 6373 4628 6414 4636
rect 6496 4632 6509 4656
rect 6524 4654 6539 4656
rect 6336 4618 6337 4628
rect 6352 4618 6365 4628
rect 6379 4618 6380 4628
rect 6395 4618 6408 4628
rect 6423 4618 6453 4632
rect 6496 4618 6539 4632
rect 6563 4629 6570 4636
rect 6573 4632 6640 4656
rect 6672 4656 6844 4658
rect 6642 4634 6670 4638
rect 6672 4634 6752 4656
rect 6773 4654 6788 4656
rect 6642 4632 6752 4634
rect 6573 4628 6752 4632
rect 6546 4618 6576 4628
rect 6578 4618 6731 4628
rect 6739 4618 6769 4628
rect 6773 4618 6803 4632
rect 6831 4618 6844 4656
rect 6916 4662 6951 4670
rect 6916 4636 6917 4662
rect 6924 4636 6951 4662
rect 6859 4618 6889 4632
rect 6916 4628 6951 4636
rect 6953 4662 6994 4670
rect 6953 4636 6968 4662
rect 6975 4636 6994 4662
rect 7058 4658 7120 4670
rect 7132 4658 7207 4670
rect 7265 4658 7340 4670
rect 7352 4658 7383 4670
rect 7389 4658 7424 4670
rect 7058 4656 7220 4658
rect 6953 4628 6994 4636
rect 7076 4632 7089 4656
rect 7104 4654 7119 4656
rect 6916 4618 6917 4628
rect 6932 4618 6945 4628
rect 6959 4618 6960 4628
rect 6975 4618 6988 4628
rect 7003 4618 7033 4632
rect 7076 4618 7119 4632
rect 7143 4629 7150 4636
rect 7153 4632 7220 4656
rect 7252 4656 7424 4658
rect 7222 4634 7250 4638
rect 7252 4634 7332 4656
rect 7353 4654 7368 4656
rect 7222 4632 7332 4634
rect 7153 4628 7332 4632
rect 7126 4618 7156 4628
rect 7158 4618 7311 4628
rect 7319 4618 7349 4628
rect 7353 4618 7383 4632
rect 7411 4618 7424 4656
rect 7496 4662 7531 4670
rect 7496 4636 7497 4662
rect 7504 4636 7531 4662
rect 7439 4618 7469 4632
rect 7496 4628 7531 4636
rect 7533 4662 7574 4670
rect 7533 4636 7548 4662
rect 7555 4636 7574 4662
rect 7638 4658 7700 4670
rect 7712 4658 7787 4670
rect 7845 4658 7920 4670
rect 7932 4658 7963 4670
rect 7969 4658 8004 4670
rect 7638 4656 7800 4658
rect 7533 4628 7574 4636
rect 7656 4632 7669 4656
rect 7684 4654 7699 4656
rect 7496 4618 7497 4628
rect 7512 4618 7525 4628
rect 7539 4618 7540 4628
rect 7555 4618 7568 4628
rect 7583 4618 7613 4632
rect 7656 4618 7699 4632
rect 7723 4629 7730 4636
rect 7733 4632 7800 4656
rect 7832 4656 8004 4658
rect 7802 4634 7830 4638
rect 7832 4634 7912 4656
rect 7933 4654 7948 4656
rect 7802 4632 7912 4634
rect 7733 4628 7912 4632
rect 7706 4618 7736 4628
rect 7738 4618 7891 4628
rect 7899 4618 7929 4628
rect 7933 4618 7963 4632
rect 7991 4618 8004 4656
rect 8076 4662 8111 4670
rect 8076 4636 8077 4662
rect 8084 4636 8111 4662
rect 8019 4618 8049 4632
rect 8076 4628 8111 4636
rect 8113 4662 8154 4670
rect 8113 4636 8128 4662
rect 8135 4636 8154 4662
rect 8218 4658 8280 4670
rect 8292 4658 8367 4670
rect 8425 4658 8500 4670
rect 8512 4658 8543 4670
rect 8549 4658 8584 4670
rect 8218 4656 8380 4658
rect 8113 4628 8154 4636
rect 8236 4632 8249 4656
rect 8264 4654 8279 4656
rect 8076 4618 8077 4628
rect 8092 4618 8105 4628
rect 8119 4618 8120 4628
rect 8135 4618 8148 4628
rect 8163 4618 8193 4632
rect 8236 4618 8279 4632
rect 8303 4629 8310 4636
rect 8313 4632 8380 4656
rect 8412 4656 8584 4658
rect 8382 4634 8410 4638
rect 8412 4634 8492 4656
rect 8513 4654 8528 4656
rect 8382 4632 8492 4634
rect 8313 4628 8492 4632
rect 8286 4618 8316 4628
rect 8318 4618 8471 4628
rect 8479 4618 8509 4628
rect 8513 4618 8543 4632
rect 8571 4618 8584 4656
rect 8656 4662 8691 4670
rect 8656 4636 8657 4662
rect 8664 4636 8691 4662
rect 8599 4618 8629 4632
rect 8656 4628 8691 4636
rect 8693 4662 8734 4670
rect 8693 4636 8708 4662
rect 8715 4636 8734 4662
rect 8798 4658 8860 4670
rect 8872 4658 8947 4670
rect 9005 4658 9080 4670
rect 9092 4658 9123 4670
rect 9129 4658 9164 4670
rect 8798 4656 8960 4658
rect 8693 4628 8734 4636
rect 8816 4632 8829 4656
rect 8844 4654 8859 4656
rect 8656 4618 8657 4628
rect 8672 4618 8685 4628
rect 8699 4618 8700 4628
rect 8715 4618 8728 4628
rect 8743 4618 8773 4632
rect 8816 4618 8859 4632
rect 8883 4629 8890 4636
rect 8893 4632 8960 4656
rect 8992 4656 9164 4658
rect 8962 4634 8990 4638
rect 8992 4634 9072 4656
rect 9093 4654 9108 4656
rect 8962 4632 9072 4634
rect 8893 4628 9072 4632
rect 8866 4618 8896 4628
rect 8898 4618 9051 4628
rect 9059 4618 9089 4628
rect 9093 4618 9123 4632
rect 9151 4618 9164 4656
rect 9236 4662 9271 4670
rect 9236 4636 9237 4662
rect 9244 4636 9271 4662
rect 9179 4618 9209 4632
rect 9236 4628 9271 4636
rect 9236 4618 9237 4628
rect 9252 4618 9265 4628
rect -1 4612 9265 4618
rect 0 4604 9265 4612
rect 15 4574 28 4604
rect 43 4586 73 4604
rect 116 4590 130 4604
rect 166 4590 386 4604
rect 117 4588 130 4590
rect 83 4576 98 4588
rect 80 4574 102 4576
rect 107 4574 137 4588
rect 198 4586 351 4590
rect 180 4574 372 4586
rect 415 4574 445 4588
rect 451 4574 464 4604
rect 479 4586 509 4604
rect 552 4574 565 4604
rect 595 4574 608 4604
rect 623 4586 653 4604
rect 696 4590 710 4604
rect 746 4590 966 4604
rect 697 4588 710 4590
rect 663 4576 678 4588
rect 660 4574 682 4576
rect 687 4574 717 4588
rect 778 4586 931 4590
rect 760 4574 952 4586
rect 995 4574 1025 4588
rect 1031 4574 1044 4604
rect 1059 4586 1089 4604
rect 1132 4574 1145 4604
rect 1175 4574 1188 4604
rect 1203 4586 1233 4604
rect 1276 4590 1290 4604
rect 1326 4590 1546 4604
rect 1277 4588 1290 4590
rect 1243 4576 1258 4588
rect 1240 4574 1262 4576
rect 1267 4574 1297 4588
rect 1358 4586 1511 4590
rect 1340 4574 1532 4586
rect 1575 4574 1605 4588
rect 1611 4574 1624 4604
rect 1639 4586 1669 4604
rect 1712 4574 1725 4604
rect 1755 4574 1768 4604
rect 1783 4586 1813 4604
rect 1856 4590 1870 4604
rect 1906 4590 2126 4604
rect 1857 4588 1870 4590
rect 1823 4576 1838 4588
rect 1820 4574 1842 4576
rect 1847 4574 1877 4588
rect 1938 4586 2091 4590
rect 1920 4574 2112 4586
rect 2155 4574 2185 4588
rect 2191 4574 2204 4604
rect 2219 4586 2249 4604
rect 2292 4574 2305 4604
rect 2335 4574 2348 4604
rect 2363 4586 2393 4604
rect 2436 4590 2450 4604
rect 2486 4590 2706 4604
rect 2437 4588 2450 4590
rect 2403 4576 2418 4588
rect 2400 4574 2422 4576
rect 2427 4574 2457 4588
rect 2518 4586 2671 4590
rect 2500 4574 2692 4586
rect 2735 4574 2765 4588
rect 2771 4574 2784 4604
rect 2799 4586 2829 4604
rect 2872 4574 2885 4604
rect 2915 4574 2928 4604
rect 2943 4586 2973 4604
rect 3016 4590 3030 4604
rect 3066 4590 3286 4604
rect 3017 4588 3030 4590
rect 2983 4576 2998 4588
rect 2980 4574 3002 4576
rect 3007 4574 3037 4588
rect 3098 4586 3251 4590
rect 3080 4574 3272 4586
rect 3315 4574 3345 4588
rect 3351 4574 3364 4604
rect 3379 4586 3409 4604
rect 3452 4574 3465 4604
rect 3495 4574 3508 4604
rect 3523 4586 3553 4604
rect 3596 4590 3610 4604
rect 3646 4590 3866 4604
rect 3597 4588 3610 4590
rect 3563 4576 3578 4588
rect 3560 4574 3582 4576
rect 3587 4574 3617 4588
rect 3678 4586 3831 4590
rect 3660 4574 3852 4586
rect 3895 4574 3925 4588
rect 3931 4574 3944 4604
rect 3959 4586 3989 4604
rect 4032 4574 4045 4604
rect 4075 4574 4088 4604
rect 4103 4586 4133 4604
rect 4176 4590 4190 4604
rect 4226 4590 4446 4604
rect 4177 4588 4190 4590
rect 4143 4576 4158 4588
rect 4140 4574 4162 4576
rect 4167 4574 4197 4588
rect 4258 4586 4411 4590
rect 4240 4574 4432 4586
rect 4475 4574 4505 4588
rect 4511 4574 4524 4604
rect 4539 4586 4569 4604
rect 4612 4574 4625 4604
rect 4655 4574 4668 4604
rect 4683 4586 4713 4604
rect 4756 4590 4770 4604
rect 4806 4590 5026 4604
rect 4757 4588 4770 4590
rect 4723 4576 4738 4588
rect 4720 4574 4742 4576
rect 4747 4574 4777 4588
rect 4838 4586 4991 4590
rect 4820 4574 5012 4586
rect 5055 4574 5085 4588
rect 5091 4574 5104 4604
rect 5119 4586 5149 4604
rect 5192 4574 5205 4604
rect 5235 4574 5248 4604
rect 5263 4586 5293 4604
rect 5336 4590 5350 4604
rect 5386 4590 5606 4604
rect 5337 4588 5350 4590
rect 5303 4576 5318 4588
rect 5300 4574 5322 4576
rect 5327 4574 5357 4588
rect 5418 4586 5571 4590
rect 5400 4574 5592 4586
rect 5635 4574 5665 4588
rect 5671 4574 5684 4604
rect 5699 4586 5729 4604
rect 5772 4574 5785 4604
rect 5815 4574 5828 4604
rect 5843 4586 5873 4604
rect 5916 4590 5930 4604
rect 5966 4590 6186 4604
rect 5917 4588 5930 4590
rect 5883 4576 5898 4588
rect 5880 4574 5902 4576
rect 5907 4574 5937 4588
rect 5998 4586 6151 4590
rect 5980 4574 6172 4586
rect 6215 4574 6245 4588
rect 6251 4574 6264 4604
rect 6279 4586 6309 4604
rect 6352 4574 6365 4604
rect 6395 4574 6408 4604
rect 6423 4586 6453 4604
rect 6496 4590 6510 4604
rect 6546 4590 6766 4604
rect 6497 4588 6510 4590
rect 6463 4576 6478 4588
rect 6460 4574 6482 4576
rect 6487 4574 6517 4588
rect 6578 4586 6731 4590
rect 6560 4574 6752 4586
rect 6795 4574 6825 4588
rect 6831 4574 6844 4604
rect 6859 4586 6889 4604
rect 6932 4574 6945 4604
rect 6975 4574 6988 4604
rect 7003 4586 7033 4604
rect 7076 4590 7090 4604
rect 7126 4590 7346 4604
rect 7077 4588 7090 4590
rect 7043 4576 7058 4588
rect 7040 4574 7062 4576
rect 7067 4574 7097 4588
rect 7158 4586 7311 4590
rect 7140 4574 7332 4586
rect 7375 4574 7405 4588
rect 7411 4574 7424 4604
rect 7439 4586 7469 4604
rect 7512 4574 7525 4604
rect 7555 4574 7568 4604
rect 7583 4586 7613 4604
rect 7656 4590 7670 4604
rect 7706 4590 7926 4604
rect 7657 4588 7670 4590
rect 7623 4576 7638 4588
rect 7620 4574 7642 4576
rect 7647 4574 7677 4588
rect 7738 4586 7891 4590
rect 7720 4574 7912 4586
rect 7955 4574 7985 4588
rect 7991 4574 8004 4604
rect 8019 4586 8049 4604
rect 8092 4574 8105 4604
rect 8135 4574 8148 4604
rect 8163 4586 8193 4604
rect 8236 4590 8250 4604
rect 8286 4590 8506 4604
rect 8237 4588 8250 4590
rect 8203 4576 8218 4588
rect 8200 4574 8222 4576
rect 8227 4574 8257 4588
rect 8318 4586 8471 4590
rect 8300 4574 8492 4586
rect 8535 4574 8565 4588
rect 8571 4574 8584 4604
rect 8599 4586 8629 4604
rect 8672 4574 8685 4604
rect 8715 4574 8728 4604
rect 8743 4586 8773 4604
rect 8816 4590 8830 4604
rect 8866 4590 9086 4604
rect 8817 4588 8830 4590
rect 8783 4576 8798 4588
rect 8780 4574 8802 4576
rect 8807 4574 8837 4588
rect 8898 4586 9051 4590
rect 8880 4574 9072 4586
rect 9115 4574 9145 4588
rect 9151 4574 9164 4604
rect 9179 4586 9209 4604
rect 9252 4574 9265 4604
rect 0 4560 9265 4574
rect 15 4456 28 4560
rect 73 4538 74 4548
rect 89 4538 102 4548
rect 73 4534 102 4538
rect 107 4534 137 4560
rect 155 4546 171 4548
rect 243 4546 296 4560
rect 244 4544 308 4546
rect 351 4544 366 4560
rect 415 4557 445 4560
rect 415 4554 451 4557
rect 381 4546 397 4548
rect 155 4534 170 4538
rect 73 4532 170 4534
rect 198 4532 366 4544
rect 382 4534 397 4538
rect 415 4535 454 4554
rect 473 4548 480 4549
rect 479 4541 480 4548
rect 463 4538 464 4541
rect 479 4538 492 4541
rect 415 4534 445 4535
rect 454 4534 460 4535
rect 463 4534 492 4538
rect 382 4533 492 4534
rect 382 4532 498 4533
rect 57 4524 108 4532
rect 57 4512 82 4524
rect 89 4512 108 4524
rect 139 4524 189 4532
rect 139 4516 155 4524
rect 162 4522 189 4524
rect 198 4522 419 4532
rect 162 4512 419 4522
rect 448 4524 498 4532
rect 448 4515 464 4524
rect 57 4504 108 4512
rect 155 4504 419 4512
rect 445 4512 464 4515
rect 471 4512 498 4524
rect 445 4504 498 4512
rect 73 4496 74 4504
rect 89 4496 102 4504
rect 73 4488 89 4496
rect 70 4481 89 4484
rect 70 4472 92 4481
rect 43 4462 92 4472
rect 43 4456 73 4462
rect 92 4457 97 4462
rect 15 4440 89 4456
rect 107 4448 137 4504
rect 172 4494 380 4504
rect 415 4500 460 4504
rect 463 4503 464 4504
rect 479 4503 492 4504
rect 198 4464 387 4494
rect 213 4461 387 4464
rect 206 4458 387 4461
rect 15 4438 28 4440
rect 43 4438 77 4440
rect 15 4422 89 4438
rect 116 4434 129 4448
rect 144 4434 160 4450
rect 206 4445 217 4458
rect -1 4400 0 4416
rect 15 4400 28 4422
rect 43 4400 73 4422
rect 116 4418 178 4434
rect 206 4427 217 4443
rect 222 4438 232 4458
rect 242 4438 256 4458
rect 259 4445 268 4458
rect 284 4445 293 4458
rect 222 4427 256 4438
rect 259 4427 268 4443
rect 284 4427 293 4443
rect 300 4438 310 4458
rect 320 4438 334 4458
rect 335 4445 346 4458
rect 300 4427 334 4438
rect 335 4427 346 4443
rect 392 4434 408 4450
rect 415 4448 445 4500
rect 479 4496 480 4503
rect 464 4488 480 4496
rect 451 4456 464 4475
rect 479 4456 509 4472
rect 451 4440 525 4456
rect 451 4438 464 4440
rect 479 4438 513 4440
rect 116 4416 129 4418
rect 144 4416 178 4418
rect 116 4400 178 4416
rect 222 4411 238 4414
rect 300 4411 330 4422
rect 378 4418 424 4434
rect 451 4422 525 4438
rect 378 4416 412 4418
rect 377 4400 424 4416
rect 451 4400 464 4422
rect 479 4400 509 4422
rect 536 4400 537 4416
rect 552 4400 565 4560
rect 595 4456 608 4560
rect 653 4538 654 4548
rect 669 4538 682 4548
rect 653 4534 682 4538
rect 687 4534 717 4560
rect 735 4546 751 4548
rect 823 4546 876 4560
rect 824 4544 888 4546
rect 931 4544 946 4560
rect 995 4557 1025 4560
rect 995 4554 1031 4557
rect 961 4546 977 4548
rect 735 4534 750 4538
rect 653 4532 750 4534
rect 778 4532 946 4544
rect 962 4534 977 4538
rect 995 4535 1034 4554
rect 1053 4548 1060 4549
rect 1059 4541 1060 4548
rect 1043 4538 1044 4541
rect 1059 4538 1072 4541
rect 995 4534 1025 4535
rect 1034 4534 1040 4535
rect 1043 4534 1072 4538
rect 962 4533 1072 4534
rect 962 4532 1078 4533
rect 637 4524 688 4532
rect 637 4512 662 4524
rect 669 4512 688 4524
rect 719 4524 769 4532
rect 719 4516 735 4524
rect 742 4522 769 4524
rect 778 4522 999 4532
rect 742 4512 999 4522
rect 1028 4524 1078 4532
rect 1028 4515 1044 4524
rect 637 4504 688 4512
rect 735 4504 999 4512
rect 1025 4512 1044 4515
rect 1051 4512 1078 4524
rect 1025 4504 1078 4512
rect 653 4496 654 4504
rect 669 4496 682 4504
rect 653 4488 669 4496
rect 650 4481 669 4484
rect 650 4472 672 4481
rect 623 4462 672 4472
rect 623 4456 653 4462
rect 672 4457 677 4462
rect 595 4440 669 4456
rect 687 4448 717 4504
rect 752 4494 960 4504
rect 995 4500 1040 4504
rect 1043 4503 1044 4504
rect 1059 4503 1072 4504
rect 778 4464 967 4494
rect 793 4461 967 4464
rect 786 4458 967 4461
rect 595 4438 608 4440
rect 623 4438 657 4440
rect 595 4422 669 4438
rect 696 4434 709 4448
rect 724 4434 740 4450
rect 786 4445 797 4458
rect 579 4400 580 4416
rect 595 4400 608 4422
rect 623 4400 653 4422
rect 696 4418 758 4434
rect 786 4427 797 4443
rect 802 4438 812 4458
rect 822 4438 836 4458
rect 839 4445 848 4458
rect 864 4445 873 4458
rect 802 4427 836 4438
rect 839 4427 848 4443
rect 864 4427 873 4443
rect 880 4438 890 4458
rect 900 4438 914 4458
rect 915 4445 926 4458
rect 880 4427 914 4438
rect 915 4427 926 4443
rect 972 4434 988 4450
rect 995 4448 1025 4500
rect 1059 4496 1060 4503
rect 1044 4488 1060 4496
rect 1031 4456 1044 4475
rect 1059 4456 1089 4472
rect 1031 4440 1105 4456
rect 1031 4438 1044 4440
rect 1059 4438 1093 4440
rect 696 4416 709 4418
rect 724 4416 758 4418
rect 696 4400 758 4416
rect 802 4411 818 4414
rect 880 4411 910 4422
rect 958 4418 1004 4434
rect 1031 4422 1105 4438
rect 958 4416 992 4418
rect 957 4400 1004 4416
rect 1031 4400 1044 4422
rect 1059 4400 1089 4422
rect 1116 4400 1117 4416
rect 1132 4400 1145 4560
rect 1175 4456 1188 4560
rect 1233 4538 1234 4548
rect 1249 4538 1262 4548
rect 1233 4534 1262 4538
rect 1267 4534 1297 4560
rect 1315 4546 1331 4548
rect 1403 4546 1456 4560
rect 1404 4544 1468 4546
rect 1511 4544 1526 4560
rect 1575 4557 1605 4560
rect 1575 4554 1611 4557
rect 1541 4546 1557 4548
rect 1315 4534 1330 4538
rect 1233 4532 1330 4534
rect 1358 4532 1526 4544
rect 1542 4534 1557 4538
rect 1575 4535 1614 4554
rect 1633 4548 1640 4549
rect 1639 4541 1640 4548
rect 1623 4538 1624 4541
rect 1639 4538 1652 4541
rect 1575 4534 1605 4535
rect 1614 4534 1620 4535
rect 1623 4534 1652 4538
rect 1542 4533 1652 4534
rect 1542 4532 1658 4533
rect 1217 4524 1268 4532
rect 1217 4512 1242 4524
rect 1249 4512 1268 4524
rect 1299 4524 1349 4532
rect 1299 4516 1315 4524
rect 1322 4522 1349 4524
rect 1358 4522 1579 4532
rect 1322 4512 1579 4522
rect 1608 4524 1658 4532
rect 1608 4515 1624 4524
rect 1217 4504 1268 4512
rect 1315 4504 1579 4512
rect 1605 4512 1624 4515
rect 1631 4512 1658 4524
rect 1605 4504 1658 4512
rect 1233 4496 1234 4504
rect 1249 4496 1262 4504
rect 1233 4488 1249 4496
rect 1230 4481 1249 4484
rect 1230 4472 1252 4481
rect 1203 4462 1252 4472
rect 1203 4456 1233 4462
rect 1252 4457 1257 4462
rect 1175 4440 1249 4456
rect 1267 4448 1297 4504
rect 1332 4494 1540 4504
rect 1575 4500 1620 4504
rect 1623 4503 1624 4504
rect 1639 4503 1652 4504
rect 1358 4464 1547 4494
rect 1373 4461 1547 4464
rect 1366 4458 1547 4461
rect 1175 4438 1188 4440
rect 1203 4438 1237 4440
rect 1175 4422 1249 4438
rect 1276 4434 1289 4448
rect 1304 4434 1320 4450
rect 1366 4445 1377 4458
rect 1159 4400 1160 4416
rect 1175 4400 1188 4422
rect 1203 4400 1233 4422
rect 1276 4418 1338 4434
rect 1366 4427 1377 4443
rect 1382 4438 1392 4458
rect 1402 4438 1416 4458
rect 1419 4445 1428 4458
rect 1444 4445 1453 4458
rect 1382 4427 1416 4438
rect 1419 4427 1428 4443
rect 1444 4427 1453 4443
rect 1460 4438 1470 4458
rect 1480 4438 1494 4458
rect 1495 4445 1506 4458
rect 1460 4427 1494 4438
rect 1495 4427 1506 4443
rect 1552 4434 1568 4450
rect 1575 4448 1605 4500
rect 1639 4496 1640 4503
rect 1624 4488 1640 4496
rect 1611 4456 1624 4475
rect 1639 4456 1669 4472
rect 1611 4440 1685 4456
rect 1611 4438 1624 4440
rect 1639 4438 1673 4440
rect 1276 4416 1289 4418
rect 1304 4416 1338 4418
rect 1276 4400 1338 4416
rect 1382 4411 1398 4414
rect 1460 4411 1490 4422
rect 1538 4418 1584 4434
rect 1611 4422 1685 4438
rect 1538 4416 1572 4418
rect 1537 4400 1584 4416
rect 1611 4400 1624 4422
rect 1639 4400 1669 4422
rect 1696 4400 1697 4416
rect 1712 4400 1725 4560
rect 1755 4456 1768 4560
rect 1813 4538 1814 4548
rect 1829 4538 1842 4548
rect 1813 4534 1842 4538
rect 1847 4534 1877 4560
rect 1895 4546 1911 4548
rect 1983 4546 2036 4560
rect 1984 4544 2048 4546
rect 2091 4544 2106 4560
rect 2155 4557 2185 4560
rect 2155 4554 2191 4557
rect 2121 4546 2137 4548
rect 1895 4534 1910 4538
rect 1813 4532 1910 4534
rect 1938 4532 2106 4544
rect 2122 4534 2137 4538
rect 2155 4535 2194 4554
rect 2213 4548 2220 4549
rect 2219 4541 2220 4548
rect 2203 4538 2204 4541
rect 2219 4538 2232 4541
rect 2155 4534 2185 4535
rect 2194 4534 2200 4535
rect 2203 4534 2232 4538
rect 2122 4533 2232 4534
rect 2122 4532 2238 4533
rect 1797 4524 1848 4532
rect 1797 4512 1822 4524
rect 1829 4512 1848 4524
rect 1879 4524 1929 4532
rect 1879 4516 1895 4524
rect 1902 4522 1929 4524
rect 1938 4522 2159 4532
rect 1902 4512 2159 4522
rect 2188 4524 2238 4532
rect 2188 4515 2204 4524
rect 1797 4504 1848 4512
rect 1895 4504 2159 4512
rect 2185 4512 2204 4515
rect 2211 4512 2238 4524
rect 2185 4504 2238 4512
rect 1813 4496 1814 4504
rect 1829 4496 1842 4504
rect 1813 4488 1829 4496
rect 1810 4481 1829 4484
rect 1810 4472 1832 4481
rect 1783 4462 1832 4472
rect 1783 4456 1813 4462
rect 1832 4457 1837 4462
rect 1755 4440 1829 4456
rect 1847 4448 1877 4504
rect 1912 4494 2120 4504
rect 2155 4500 2200 4504
rect 2203 4503 2204 4504
rect 2219 4503 2232 4504
rect 1938 4464 2127 4494
rect 1953 4461 2127 4464
rect 1946 4458 2127 4461
rect 1755 4438 1768 4440
rect 1783 4438 1817 4440
rect 1755 4422 1829 4438
rect 1856 4434 1869 4448
rect 1884 4434 1900 4450
rect 1946 4445 1957 4458
rect 1739 4400 1740 4416
rect 1755 4400 1768 4422
rect 1783 4400 1813 4422
rect 1856 4418 1918 4434
rect 1946 4427 1957 4443
rect 1962 4438 1972 4458
rect 1982 4438 1996 4458
rect 1999 4445 2008 4458
rect 2024 4445 2033 4458
rect 1962 4427 1996 4438
rect 1999 4427 2008 4443
rect 2024 4427 2033 4443
rect 2040 4438 2050 4458
rect 2060 4438 2074 4458
rect 2075 4445 2086 4458
rect 2040 4427 2074 4438
rect 2075 4427 2086 4443
rect 2132 4434 2148 4450
rect 2155 4448 2185 4500
rect 2219 4496 2220 4503
rect 2204 4488 2220 4496
rect 2191 4456 2204 4475
rect 2219 4456 2249 4472
rect 2191 4440 2265 4456
rect 2191 4438 2204 4440
rect 2219 4438 2253 4440
rect 1856 4416 1869 4418
rect 1884 4416 1918 4418
rect 1856 4400 1918 4416
rect 1962 4411 1976 4414
rect 2040 4411 2070 4422
rect 2118 4418 2164 4434
rect 2191 4422 2265 4438
rect 2118 4416 2152 4418
rect 2117 4400 2164 4416
rect 2191 4400 2204 4422
rect 2219 4400 2249 4422
rect 2276 4400 2277 4416
rect 2292 4400 2305 4560
rect 2335 4456 2348 4560
rect 2393 4538 2394 4548
rect 2409 4538 2422 4548
rect 2393 4534 2422 4538
rect 2427 4534 2457 4560
rect 2475 4546 2491 4548
rect 2563 4546 2616 4560
rect 2564 4544 2628 4546
rect 2671 4544 2686 4560
rect 2735 4557 2765 4560
rect 2735 4554 2771 4557
rect 2701 4546 2717 4548
rect 2475 4534 2490 4538
rect 2393 4532 2490 4534
rect 2518 4532 2686 4544
rect 2702 4534 2717 4538
rect 2735 4535 2774 4554
rect 2793 4548 2800 4549
rect 2799 4541 2800 4548
rect 2783 4538 2784 4541
rect 2799 4538 2812 4541
rect 2735 4534 2765 4535
rect 2774 4534 2780 4535
rect 2783 4534 2812 4538
rect 2702 4533 2812 4534
rect 2702 4532 2818 4533
rect 2377 4524 2428 4532
rect 2377 4512 2402 4524
rect 2409 4512 2428 4524
rect 2459 4524 2509 4532
rect 2459 4516 2475 4524
rect 2482 4522 2509 4524
rect 2518 4522 2739 4532
rect 2482 4512 2739 4522
rect 2768 4524 2818 4532
rect 2768 4515 2784 4524
rect 2377 4504 2428 4512
rect 2475 4504 2739 4512
rect 2765 4512 2784 4515
rect 2791 4512 2818 4524
rect 2765 4504 2818 4512
rect 2393 4496 2394 4504
rect 2409 4496 2422 4504
rect 2393 4488 2409 4496
rect 2390 4481 2409 4484
rect 2390 4472 2412 4481
rect 2363 4462 2412 4472
rect 2363 4456 2393 4462
rect 2412 4457 2417 4462
rect 2335 4440 2409 4456
rect 2427 4448 2457 4504
rect 2492 4494 2700 4504
rect 2735 4500 2780 4504
rect 2783 4503 2784 4504
rect 2799 4503 2812 4504
rect 2518 4464 2707 4494
rect 2533 4461 2707 4464
rect 2526 4458 2707 4461
rect 2335 4438 2348 4440
rect 2363 4438 2397 4440
rect 2335 4422 2409 4438
rect 2436 4434 2449 4448
rect 2464 4434 2480 4450
rect 2526 4445 2537 4458
rect 2319 4400 2320 4416
rect 2335 4400 2348 4422
rect 2363 4400 2393 4422
rect 2436 4418 2498 4434
rect 2526 4427 2537 4443
rect 2542 4438 2552 4458
rect 2562 4438 2576 4458
rect 2579 4445 2588 4458
rect 2604 4445 2613 4458
rect 2542 4427 2576 4438
rect 2579 4427 2588 4443
rect 2604 4427 2613 4443
rect 2620 4438 2630 4458
rect 2640 4438 2654 4458
rect 2655 4445 2666 4458
rect 2620 4427 2654 4438
rect 2655 4427 2666 4443
rect 2712 4434 2728 4450
rect 2735 4448 2765 4500
rect 2799 4496 2800 4503
rect 2784 4488 2800 4496
rect 2771 4456 2784 4475
rect 2799 4456 2829 4472
rect 2771 4440 2845 4456
rect 2771 4438 2784 4440
rect 2799 4438 2833 4440
rect 2436 4416 2449 4418
rect 2464 4416 2498 4418
rect 2436 4400 2498 4416
rect 2542 4411 2558 4414
rect 2620 4411 2650 4422
rect 2698 4418 2744 4434
rect 2771 4422 2845 4438
rect 2698 4416 2732 4418
rect 2697 4400 2744 4416
rect 2771 4400 2784 4422
rect 2799 4400 2829 4422
rect 2856 4400 2857 4416
rect 2872 4400 2885 4560
rect 2915 4456 2928 4560
rect 2973 4538 2974 4548
rect 2989 4538 3002 4548
rect 2973 4534 3002 4538
rect 3007 4534 3037 4560
rect 3055 4546 3071 4548
rect 3143 4546 3196 4560
rect 3144 4544 3208 4546
rect 3251 4544 3266 4560
rect 3315 4557 3345 4560
rect 3315 4554 3351 4557
rect 3281 4546 3297 4548
rect 3055 4534 3070 4538
rect 2973 4532 3070 4534
rect 3098 4532 3266 4544
rect 3282 4534 3297 4538
rect 3315 4535 3354 4554
rect 3373 4548 3380 4549
rect 3379 4541 3380 4548
rect 3363 4538 3364 4541
rect 3379 4538 3392 4541
rect 3315 4534 3345 4535
rect 3354 4534 3360 4535
rect 3363 4534 3392 4538
rect 3282 4533 3392 4534
rect 3282 4532 3398 4533
rect 2957 4524 3008 4532
rect 2957 4512 2982 4524
rect 2989 4512 3008 4524
rect 3039 4524 3089 4532
rect 3039 4516 3055 4524
rect 3062 4522 3089 4524
rect 3098 4522 3319 4532
rect 3062 4512 3319 4522
rect 3348 4524 3398 4532
rect 3348 4515 3364 4524
rect 2957 4504 3008 4512
rect 3055 4504 3319 4512
rect 3345 4512 3364 4515
rect 3371 4512 3398 4524
rect 3345 4504 3398 4512
rect 2973 4496 2974 4504
rect 2989 4496 3002 4504
rect 2973 4488 2989 4496
rect 2970 4481 2989 4484
rect 2970 4472 2992 4481
rect 2943 4462 2992 4472
rect 2943 4456 2973 4462
rect 2992 4457 2997 4462
rect 2915 4440 2989 4456
rect 3007 4448 3037 4504
rect 3072 4494 3280 4504
rect 3315 4500 3360 4504
rect 3363 4503 3364 4504
rect 3379 4503 3392 4504
rect 3098 4464 3287 4494
rect 3113 4461 3287 4464
rect 3106 4458 3287 4461
rect 2915 4438 2928 4440
rect 2943 4438 2977 4440
rect 2915 4422 2989 4438
rect 3016 4434 3029 4448
rect 3044 4434 3060 4450
rect 3106 4445 3117 4458
rect 2899 4400 2900 4416
rect 2915 4400 2928 4422
rect 2943 4400 2973 4422
rect 3016 4418 3078 4434
rect 3106 4427 3117 4443
rect 3122 4438 3132 4458
rect 3142 4438 3156 4458
rect 3159 4445 3168 4458
rect 3184 4445 3193 4458
rect 3122 4427 3156 4438
rect 3159 4427 3168 4443
rect 3184 4427 3193 4443
rect 3200 4438 3210 4458
rect 3220 4438 3234 4458
rect 3235 4445 3246 4458
rect 3200 4427 3234 4438
rect 3235 4427 3246 4443
rect 3292 4434 3308 4450
rect 3315 4448 3345 4500
rect 3379 4496 3380 4503
rect 3364 4488 3380 4496
rect 3351 4456 3364 4475
rect 3379 4456 3409 4472
rect 3351 4440 3425 4456
rect 3351 4438 3364 4440
rect 3379 4438 3413 4440
rect 3016 4416 3029 4418
rect 3044 4416 3078 4418
rect 3016 4400 3078 4416
rect 3122 4411 3138 4414
rect 3200 4411 3230 4422
rect 3278 4418 3324 4434
rect 3351 4422 3425 4438
rect 3278 4416 3312 4418
rect 3277 4400 3324 4416
rect 3351 4400 3364 4422
rect 3379 4400 3409 4422
rect 3436 4400 3437 4416
rect 3452 4400 3465 4560
rect 3495 4456 3508 4560
rect 3553 4538 3554 4548
rect 3569 4538 3582 4548
rect 3553 4534 3582 4538
rect 3587 4534 3617 4560
rect 3635 4546 3651 4548
rect 3723 4546 3776 4560
rect 3724 4544 3788 4546
rect 3831 4544 3846 4560
rect 3895 4557 3925 4560
rect 3895 4554 3931 4557
rect 3861 4546 3877 4548
rect 3635 4534 3650 4538
rect 3553 4532 3650 4534
rect 3678 4532 3846 4544
rect 3862 4534 3877 4538
rect 3895 4535 3934 4554
rect 3953 4548 3960 4549
rect 3959 4541 3960 4548
rect 3943 4538 3944 4541
rect 3959 4538 3972 4541
rect 3895 4534 3925 4535
rect 3934 4534 3940 4535
rect 3943 4534 3972 4538
rect 3862 4533 3972 4534
rect 3862 4532 3978 4533
rect 3537 4524 3588 4532
rect 3537 4512 3562 4524
rect 3569 4512 3588 4524
rect 3619 4524 3669 4532
rect 3619 4516 3635 4524
rect 3642 4522 3669 4524
rect 3678 4522 3899 4532
rect 3642 4512 3899 4522
rect 3928 4524 3978 4532
rect 3928 4515 3944 4524
rect 3537 4504 3588 4512
rect 3635 4504 3899 4512
rect 3925 4512 3944 4515
rect 3951 4512 3978 4524
rect 3925 4504 3978 4512
rect 3553 4496 3554 4504
rect 3569 4496 3582 4504
rect 3553 4488 3569 4496
rect 3550 4481 3569 4484
rect 3550 4472 3572 4481
rect 3523 4462 3572 4472
rect 3523 4456 3553 4462
rect 3572 4457 3577 4462
rect 3495 4440 3569 4456
rect 3587 4448 3617 4504
rect 3652 4494 3860 4504
rect 3895 4500 3940 4504
rect 3943 4503 3944 4504
rect 3959 4503 3972 4504
rect 3678 4464 3867 4494
rect 3693 4461 3867 4464
rect 3686 4458 3867 4461
rect 3495 4438 3508 4440
rect 3523 4438 3557 4440
rect 3495 4422 3569 4438
rect 3596 4434 3609 4448
rect 3624 4434 3640 4450
rect 3686 4445 3697 4458
rect 3479 4400 3480 4416
rect 3495 4400 3508 4422
rect 3523 4400 3553 4422
rect 3596 4418 3658 4434
rect 3686 4427 3697 4443
rect 3702 4438 3712 4458
rect 3722 4438 3736 4458
rect 3739 4445 3748 4458
rect 3764 4445 3773 4458
rect 3702 4427 3736 4438
rect 3739 4427 3748 4443
rect 3764 4427 3773 4443
rect 3780 4438 3790 4458
rect 3800 4438 3814 4458
rect 3815 4445 3826 4458
rect 3780 4427 3814 4438
rect 3815 4427 3826 4443
rect 3872 4434 3888 4450
rect 3895 4448 3925 4500
rect 3959 4496 3960 4503
rect 3944 4488 3960 4496
rect 3931 4456 3944 4475
rect 3959 4456 3989 4472
rect 3931 4440 4005 4456
rect 3931 4438 3944 4440
rect 3959 4438 3993 4440
rect 3596 4416 3609 4418
rect 3624 4416 3658 4418
rect 3596 4400 3658 4416
rect 3702 4411 3718 4414
rect 3780 4411 3810 4422
rect 3858 4418 3904 4434
rect 3931 4422 4005 4438
rect 3858 4416 3892 4418
rect 3857 4400 3904 4416
rect 3931 4400 3944 4422
rect 3959 4400 3989 4422
rect 4016 4400 4017 4416
rect 4032 4400 4045 4560
rect 4075 4456 4088 4560
rect 4133 4538 4134 4548
rect 4149 4538 4162 4548
rect 4133 4534 4162 4538
rect 4167 4534 4197 4560
rect 4215 4546 4231 4548
rect 4303 4546 4356 4560
rect 4304 4544 4368 4546
rect 4411 4544 4426 4560
rect 4475 4557 4505 4560
rect 4475 4554 4511 4557
rect 4441 4546 4457 4548
rect 4215 4534 4230 4538
rect 4133 4532 4230 4534
rect 4258 4532 4426 4544
rect 4442 4534 4457 4538
rect 4475 4535 4514 4554
rect 4533 4548 4540 4549
rect 4539 4541 4540 4548
rect 4523 4538 4524 4541
rect 4539 4538 4552 4541
rect 4475 4534 4505 4535
rect 4514 4534 4520 4535
rect 4523 4534 4552 4538
rect 4442 4533 4552 4534
rect 4442 4532 4558 4533
rect 4117 4524 4168 4532
rect 4117 4512 4142 4524
rect 4149 4512 4168 4524
rect 4199 4524 4249 4532
rect 4199 4516 4215 4524
rect 4222 4522 4249 4524
rect 4258 4522 4479 4532
rect 4222 4512 4479 4522
rect 4508 4524 4558 4532
rect 4508 4515 4524 4524
rect 4117 4504 4168 4512
rect 4215 4504 4479 4512
rect 4505 4512 4524 4515
rect 4531 4512 4558 4524
rect 4505 4504 4558 4512
rect 4133 4496 4134 4504
rect 4149 4496 4162 4504
rect 4133 4488 4149 4496
rect 4130 4481 4149 4484
rect 4130 4472 4152 4481
rect 4103 4462 4152 4472
rect 4103 4456 4133 4462
rect 4152 4457 4157 4462
rect 4075 4440 4149 4456
rect 4167 4448 4197 4504
rect 4232 4494 4440 4504
rect 4475 4500 4520 4504
rect 4523 4503 4524 4504
rect 4539 4503 4552 4504
rect 4258 4464 4447 4494
rect 4273 4461 4447 4464
rect 4266 4458 4447 4461
rect 4075 4438 4088 4440
rect 4103 4438 4137 4440
rect 4075 4422 4149 4438
rect 4176 4434 4189 4448
rect 4204 4434 4220 4450
rect 4266 4445 4277 4458
rect 4059 4400 4060 4416
rect 4075 4400 4088 4422
rect 4103 4400 4133 4422
rect 4176 4418 4238 4434
rect 4266 4427 4277 4443
rect 4282 4438 4292 4458
rect 4302 4438 4316 4458
rect 4319 4445 4328 4458
rect 4344 4445 4353 4458
rect 4282 4427 4316 4438
rect 4319 4427 4328 4443
rect 4344 4427 4353 4443
rect 4360 4438 4370 4458
rect 4380 4438 4394 4458
rect 4395 4445 4406 4458
rect 4360 4427 4394 4438
rect 4395 4427 4406 4443
rect 4452 4434 4468 4450
rect 4475 4448 4505 4500
rect 4539 4496 4540 4503
rect 4524 4488 4540 4496
rect 4511 4456 4524 4475
rect 4539 4456 4569 4472
rect 4511 4440 4585 4456
rect 4511 4438 4524 4440
rect 4539 4438 4573 4440
rect 4176 4416 4189 4418
rect 4204 4416 4238 4418
rect 4176 4400 4238 4416
rect 4282 4411 4298 4414
rect 4360 4411 4390 4422
rect 4438 4418 4484 4434
rect 4511 4422 4585 4438
rect 4438 4416 4472 4418
rect 4437 4400 4484 4416
rect 4511 4400 4524 4422
rect 4539 4400 4569 4422
rect 4596 4400 4597 4416
rect 4612 4400 4625 4560
rect 4655 4456 4668 4560
rect 4713 4538 4714 4548
rect 4729 4538 4742 4548
rect 4713 4534 4742 4538
rect 4747 4534 4777 4560
rect 4795 4546 4811 4548
rect 4883 4546 4936 4560
rect 4884 4544 4948 4546
rect 4991 4544 5006 4560
rect 5055 4557 5085 4560
rect 5055 4554 5091 4557
rect 5021 4546 5037 4548
rect 4795 4534 4810 4538
rect 4713 4532 4810 4534
rect 4838 4532 5006 4544
rect 5022 4534 5037 4538
rect 5055 4535 5094 4554
rect 5113 4548 5120 4549
rect 5119 4541 5120 4548
rect 5103 4538 5104 4541
rect 5119 4538 5132 4541
rect 5055 4534 5085 4535
rect 5094 4534 5100 4535
rect 5103 4534 5132 4538
rect 5022 4533 5132 4534
rect 5022 4532 5138 4533
rect 4697 4524 4748 4532
rect 4697 4512 4722 4524
rect 4729 4512 4748 4524
rect 4779 4524 4829 4532
rect 4779 4516 4795 4524
rect 4802 4522 4829 4524
rect 4838 4522 5059 4532
rect 4802 4512 5059 4522
rect 5088 4524 5138 4532
rect 5088 4515 5104 4524
rect 4697 4504 4748 4512
rect 4795 4504 5059 4512
rect 5085 4512 5104 4515
rect 5111 4512 5138 4524
rect 5085 4504 5138 4512
rect 4713 4496 4714 4504
rect 4729 4496 4742 4504
rect 4713 4488 4729 4496
rect 4710 4481 4729 4484
rect 4710 4472 4732 4481
rect 4683 4462 4732 4472
rect 4683 4456 4713 4462
rect 4732 4457 4737 4462
rect 4655 4440 4729 4456
rect 4747 4448 4777 4504
rect 4812 4494 5020 4504
rect 5055 4500 5100 4504
rect 5103 4503 5104 4504
rect 5119 4503 5132 4504
rect 4838 4464 5027 4494
rect 4853 4461 5027 4464
rect 4846 4458 5027 4461
rect 4655 4438 4668 4440
rect 4683 4438 4717 4440
rect 4655 4422 4729 4438
rect 4756 4434 4769 4448
rect 4784 4434 4800 4450
rect 4846 4445 4857 4458
rect 4639 4400 4640 4416
rect 4655 4400 4668 4422
rect 4683 4400 4713 4422
rect 4756 4418 4818 4434
rect 4846 4427 4857 4443
rect 4862 4438 4872 4458
rect 4882 4438 4896 4458
rect 4899 4445 4908 4458
rect 4924 4445 4933 4458
rect 4862 4427 4896 4438
rect 4899 4427 4908 4443
rect 4924 4427 4933 4443
rect 4940 4438 4950 4458
rect 4960 4438 4974 4458
rect 4975 4445 4986 4458
rect 4940 4427 4974 4438
rect 4975 4427 4986 4443
rect 5032 4434 5048 4450
rect 5055 4448 5085 4500
rect 5119 4496 5120 4503
rect 5104 4488 5120 4496
rect 5091 4456 5104 4475
rect 5119 4456 5149 4472
rect 5091 4440 5165 4456
rect 5091 4438 5104 4440
rect 5119 4438 5153 4440
rect 4756 4416 4769 4418
rect 4784 4416 4818 4418
rect 4756 4400 4818 4416
rect 4862 4411 4878 4414
rect 4940 4411 4970 4422
rect 5018 4418 5064 4434
rect 5091 4422 5165 4438
rect 5018 4416 5052 4418
rect 5017 4400 5064 4416
rect 5091 4400 5104 4422
rect 5119 4400 5149 4422
rect 5176 4400 5177 4416
rect 5192 4400 5205 4560
rect 5235 4456 5248 4560
rect 5293 4538 5294 4548
rect 5309 4538 5322 4548
rect 5293 4534 5322 4538
rect 5327 4534 5357 4560
rect 5375 4546 5391 4548
rect 5463 4546 5516 4560
rect 5464 4544 5528 4546
rect 5571 4544 5586 4560
rect 5635 4557 5665 4560
rect 5635 4554 5671 4557
rect 5601 4546 5617 4548
rect 5375 4534 5390 4538
rect 5293 4532 5390 4534
rect 5418 4532 5586 4544
rect 5602 4534 5617 4538
rect 5635 4535 5674 4554
rect 5693 4548 5700 4549
rect 5699 4541 5700 4548
rect 5683 4538 5684 4541
rect 5699 4538 5712 4541
rect 5635 4534 5665 4535
rect 5674 4534 5680 4535
rect 5683 4534 5712 4538
rect 5602 4533 5712 4534
rect 5602 4532 5718 4533
rect 5277 4524 5328 4532
rect 5277 4512 5302 4524
rect 5309 4512 5328 4524
rect 5359 4524 5409 4532
rect 5359 4516 5375 4524
rect 5382 4522 5409 4524
rect 5418 4522 5639 4532
rect 5382 4512 5639 4522
rect 5668 4524 5718 4532
rect 5668 4515 5684 4524
rect 5277 4504 5328 4512
rect 5375 4504 5639 4512
rect 5665 4512 5684 4515
rect 5691 4512 5718 4524
rect 5665 4504 5718 4512
rect 5293 4496 5294 4504
rect 5309 4496 5322 4504
rect 5293 4488 5309 4496
rect 5290 4481 5309 4484
rect 5290 4472 5312 4481
rect 5263 4462 5312 4472
rect 5263 4456 5293 4462
rect 5312 4457 5317 4462
rect 5235 4440 5309 4456
rect 5327 4448 5357 4504
rect 5392 4494 5600 4504
rect 5635 4500 5680 4504
rect 5683 4503 5684 4504
rect 5699 4503 5712 4504
rect 5418 4464 5607 4494
rect 5433 4461 5607 4464
rect 5426 4458 5607 4461
rect 5235 4438 5248 4440
rect 5263 4438 5297 4440
rect 5235 4422 5309 4438
rect 5336 4434 5349 4448
rect 5364 4434 5380 4450
rect 5426 4445 5437 4458
rect 5219 4400 5220 4416
rect 5235 4400 5248 4422
rect 5263 4400 5293 4422
rect 5336 4418 5398 4434
rect 5426 4427 5437 4443
rect 5442 4438 5452 4458
rect 5462 4438 5476 4458
rect 5479 4445 5488 4458
rect 5504 4445 5513 4458
rect 5442 4427 5476 4438
rect 5479 4427 5488 4443
rect 5504 4427 5513 4443
rect 5520 4438 5530 4458
rect 5540 4438 5554 4458
rect 5555 4445 5566 4458
rect 5520 4427 5554 4438
rect 5555 4427 5566 4443
rect 5612 4434 5628 4450
rect 5635 4448 5665 4500
rect 5699 4496 5700 4503
rect 5684 4488 5700 4496
rect 5671 4456 5684 4475
rect 5699 4456 5729 4472
rect 5671 4440 5745 4456
rect 5671 4438 5684 4440
rect 5699 4438 5733 4440
rect 5336 4416 5349 4418
rect 5364 4416 5398 4418
rect 5336 4400 5398 4416
rect 5442 4411 5458 4414
rect 5520 4411 5550 4422
rect 5598 4418 5644 4434
rect 5671 4422 5745 4438
rect 5598 4416 5632 4418
rect 5597 4400 5644 4416
rect 5671 4400 5684 4422
rect 5699 4400 5729 4422
rect 5756 4400 5757 4416
rect 5772 4400 5785 4560
rect 5815 4456 5828 4560
rect 5873 4538 5874 4548
rect 5889 4538 5902 4548
rect 5873 4534 5902 4538
rect 5907 4534 5937 4560
rect 5955 4546 5971 4548
rect 6043 4546 6096 4560
rect 6044 4544 6108 4546
rect 6151 4544 6166 4560
rect 6215 4557 6245 4560
rect 6215 4554 6251 4557
rect 6181 4546 6197 4548
rect 5955 4534 5970 4538
rect 5873 4532 5970 4534
rect 5998 4532 6166 4544
rect 6182 4534 6197 4538
rect 6215 4535 6254 4554
rect 6273 4548 6280 4549
rect 6279 4541 6280 4548
rect 6263 4538 6264 4541
rect 6279 4538 6292 4541
rect 6215 4534 6245 4535
rect 6254 4534 6260 4535
rect 6263 4534 6292 4538
rect 6182 4533 6292 4534
rect 6182 4532 6298 4533
rect 5857 4524 5908 4532
rect 5857 4512 5882 4524
rect 5889 4512 5908 4524
rect 5939 4524 5989 4532
rect 5939 4516 5955 4524
rect 5962 4522 5989 4524
rect 5998 4522 6219 4532
rect 5962 4512 6219 4522
rect 6248 4524 6298 4532
rect 6248 4515 6264 4524
rect 5857 4504 5908 4512
rect 5955 4504 6219 4512
rect 6245 4512 6264 4515
rect 6271 4512 6298 4524
rect 6245 4504 6298 4512
rect 5873 4496 5874 4504
rect 5889 4496 5902 4504
rect 5873 4488 5889 4496
rect 5870 4481 5889 4484
rect 5870 4472 5892 4481
rect 5843 4462 5892 4472
rect 5843 4456 5873 4462
rect 5892 4457 5897 4462
rect 5815 4440 5889 4456
rect 5907 4448 5937 4504
rect 5972 4494 6180 4504
rect 6215 4500 6260 4504
rect 6263 4503 6264 4504
rect 6279 4503 6292 4504
rect 5998 4464 6187 4494
rect 6013 4461 6187 4464
rect 6006 4458 6187 4461
rect 5815 4438 5828 4440
rect 5843 4438 5877 4440
rect 5815 4422 5889 4438
rect 5916 4434 5929 4448
rect 5944 4434 5960 4450
rect 6006 4445 6017 4458
rect 5799 4400 5800 4416
rect 5815 4400 5828 4422
rect 5843 4400 5873 4422
rect 5916 4418 5978 4434
rect 6006 4427 6017 4443
rect 6022 4438 6032 4458
rect 6042 4438 6056 4458
rect 6059 4445 6068 4458
rect 6084 4445 6093 4458
rect 6022 4427 6056 4438
rect 6059 4427 6068 4443
rect 6084 4427 6093 4443
rect 6100 4438 6110 4458
rect 6120 4438 6134 4458
rect 6135 4445 6146 4458
rect 6100 4427 6134 4438
rect 6135 4427 6146 4443
rect 6192 4434 6208 4450
rect 6215 4448 6245 4500
rect 6279 4496 6280 4503
rect 6264 4488 6280 4496
rect 6251 4456 6264 4475
rect 6279 4456 6309 4472
rect 6251 4440 6325 4456
rect 6251 4438 6264 4440
rect 6279 4438 6313 4440
rect 5916 4416 5929 4418
rect 5944 4416 5978 4418
rect 5916 4400 5978 4416
rect 6022 4411 6038 4414
rect 6100 4411 6130 4422
rect 6178 4418 6224 4434
rect 6251 4422 6325 4438
rect 6178 4416 6212 4418
rect 6177 4400 6224 4416
rect 6251 4400 6264 4422
rect 6279 4400 6309 4422
rect 6336 4400 6337 4416
rect 6352 4400 6365 4560
rect 6395 4456 6408 4560
rect 6453 4538 6454 4548
rect 6469 4538 6482 4548
rect 6453 4534 6482 4538
rect 6487 4534 6517 4560
rect 6535 4546 6551 4548
rect 6623 4546 6676 4560
rect 6624 4544 6688 4546
rect 6731 4544 6746 4560
rect 6795 4557 6825 4560
rect 6795 4554 6831 4557
rect 6761 4546 6777 4548
rect 6535 4534 6550 4538
rect 6453 4532 6550 4534
rect 6578 4532 6746 4544
rect 6762 4534 6777 4538
rect 6795 4535 6834 4554
rect 6853 4548 6860 4549
rect 6859 4541 6860 4548
rect 6843 4538 6844 4541
rect 6859 4538 6872 4541
rect 6795 4534 6825 4535
rect 6834 4534 6840 4535
rect 6843 4534 6872 4538
rect 6762 4533 6872 4534
rect 6762 4532 6878 4533
rect 6437 4524 6488 4532
rect 6437 4512 6462 4524
rect 6469 4512 6488 4524
rect 6519 4524 6569 4532
rect 6519 4516 6535 4524
rect 6542 4522 6569 4524
rect 6578 4522 6799 4532
rect 6542 4512 6799 4522
rect 6828 4524 6878 4532
rect 6828 4515 6844 4524
rect 6437 4504 6488 4512
rect 6535 4504 6799 4512
rect 6825 4512 6844 4515
rect 6851 4512 6878 4524
rect 6825 4504 6878 4512
rect 6453 4496 6454 4504
rect 6469 4496 6482 4504
rect 6453 4488 6469 4496
rect 6450 4481 6469 4484
rect 6450 4472 6472 4481
rect 6423 4462 6472 4472
rect 6423 4456 6453 4462
rect 6472 4457 6477 4462
rect 6395 4440 6469 4456
rect 6487 4448 6517 4504
rect 6552 4494 6760 4504
rect 6795 4500 6840 4504
rect 6843 4503 6844 4504
rect 6859 4503 6872 4504
rect 6578 4464 6767 4494
rect 6593 4461 6767 4464
rect 6586 4458 6767 4461
rect 6395 4438 6408 4440
rect 6423 4438 6457 4440
rect 6395 4422 6469 4438
rect 6496 4434 6509 4448
rect 6524 4434 6540 4450
rect 6586 4445 6597 4458
rect 6379 4400 6380 4416
rect 6395 4400 6408 4422
rect 6423 4400 6453 4422
rect 6496 4418 6558 4434
rect 6586 4427 6597 4443
rect 6602 4438 6612 4458
rect 6622 4438 6636 4458
rect 6639 4445 6648 4458
rect 6664 4445 6673 4458
rect 6602 4427 6636 4438
rect 6639 4427 6648 4443
rect 6664 4427 6673 4443
rect 6680 4438 6690 4458
rect 6700 4438 6714 4458
rect 6715 4445 6726 4458
rect 6680 4427 6714 4438
rect 6715 4427 6726 4443
rect 6772 4434 6788 4450
rect 6795 4448 6825 4500
rect 6859 4496 6860 4503
rect 6844 4488 6860 4496
rect 6831 4456 6844 4475
rect 6859 4456 6889 4472
rect 6831 4440 6905 4456
rect 6831 4438 6844 4440
rect 6859 4438 6893 4440
rect 6496 4416 6509 4418
rect 6524 4416 6558 4418
rect 6496 4400 6558 4416
rect 6602 4411 6618 4414
rect 6680 4411 6710 4422
rect 6758 4418 6804 4434
rect 6831 4422 6905 4438
rect 6758 4416 6792 4418
rect 6757 4400 6804 4416
rect 6831 4400 6844 4422
rect 6859 4400 6889 4422
rect 6916 4400 6917 4416
rect 6932 4400 6945 4560
rect 6975 4456 6988 4560
rect 7033 4538 7034 4548
rect 7049 4538 7062 4548
rect 7033 4534 7062 4538
rect 7067 4534 7097 4560
rect 7115 4546 7131 4548
rect 7203 4546 7256 4560
rect 7204 4544 7268 4546
rect 7311 4544 7326 4560
rect 7375 4557 7405 4560
rect 7375 4554 7411 4557
rect 7341 4546 7357 4548
rect 7115 4534 7130 4538
rect 7033 4532 7130 4534
rect 7158 4532 7326 4544
rect 7342 4534 7357 4538
rect 7375 4535 7414 4554
rect 7433 4548 7440 4549
rect 7439 4541 7440 4548
rect 7423 4538 7424 4541
rect 7439 4538 7452 4541
rect 7375 4534 7405 4535
rect 7414 4534 7420 4535
rect 7423 4534 7452 4538
rect 7342 4533 7452 4534
rect 7342 4532 7458 4533
rect 7017 4524 7068 4532
rect 7017 4512 7042 4524
rect 7049 4512 7068 4524
rect 7099 4524 7149 4532
rect 7099 4516 7115 4524
rect 7122 4522 7149 4524
rect 7158 4522 7379 4532
rect 7122 4512 7379 4522
rect 7408 4524 7458 4532
rect 7408 4515 7424 4524
rect 7017 4504 7068 4512
rect 7115 4504 7379 4512
rect 7405 4512 7424 4515
rect 7431 4512 7458 4524
rect 7405 4504 7458 4512
rect 7033 4496 7034 4504
rect 7049 4496 7062 4504
rect 7033 4488 7049 4496
rect 7030 4481 7049 4484
rect 7030 4472 7052 4481
rect 7003 4462 7052 4472
rect 7003 4456 7033 4462
rect 7052 4457 7057 4462
rect 6975 4440 7049 4456
rect 7067 4448 7097 4504
rect 7132 4494 7340 4504
rect 7375 4500 7420 4504
rect 7423 4503 7424 4504
rect 7439 4503 7452 4504
rect 7158 4464 7347 4494
rect 7173 4461 7347 4464
rect 7166 4458 7347 4461
rect 6975 4438 6988 4440
rect 7003 4438 7037 4440
rect 6975 4422 7049 4438
rect 7076 4434 7089 4448
rect 7104 4434 7120 4450
rect 7166 4445 7177 4458
rect 6959 4400 6960 4416
rect 6975 4400 6988 4422
rect 7003 4400 7033 4422
rect 7076 4418 7138 4434
rect 7166 4427 7177 4443
rect 7182 4438 7192 4458
rect 7202 4438 7216 4458
rect 7219 4445 7228 4458
rect 7244 4445 7253 4458
rect 7182 4427 7216 4438
rect 7219 4427 7228 4443
rect 7244 4427 7253 4443
rect 7260 4438 7270 4458
rect 7280 4438 7294 4458
rect 7295 4445 7306 4458
rect 7260 4427 7294 4438
rect 7295 4427 7306 4443
rect 7352 4434 7368 4450
rect 7375 4448 7405 4500
rect 7439 4496 7440 4503
rect 7424 4488 7440 4496
rect 7411 4456 7424 4475
rect 7439 4456 7469 4472
rect 7411 4440 7485 4456
rect 7411 4438 7424 4440
rect 7439 4438 7473 4440
rect 7076 4416 7089 4418
rect 7104 4416 7138 4418
rect 7076 4400 7138 4416
rect 7182 4411 7198 4414
rect 7260 4411 7290 4422
rect 7338 4418 7384 4434
rect 7411 4422 7485 4438
rect 7338 4416 7372 4418
rect 7337 4400 7384 4416
rect 7411 4400 7424 4422
rect 7439 4400 7469 4422
rect 7496 4400 7497 4416
rect 7512 4400 7525 4560
rect 7555 4456 7568 4560
rect 7613 4538 7614 4548
rect 7629 4538 7642 4548
rect 7613 4534 7642 4538
rect 7647 4534 7677 4560
rect 7695 4546 7711 4548
rect 7783 4546 7836 4560
rect 7784 4544 7848 4546
rect 7891 4544 7906 4560
rect 7955 4557 7985 4560
rect 7955 4554 7991 4557
rect 7921 4546 7937 4548
rect 7695 4534 7710 4538
rect 7613 4532 7710 4534
rect 7738 4532 7906 4544
rect 7922 4534 7937 4538
rect 7955 4535 7994 4554
rect 8013 4548 8020 4549
rect 8019 4541 8020 4548
rect 8003 4538 8004 4541
rect 8019 4538 8032 4541
rect 7955 4534 7985 4535
rect 7994 4534 8000 4535
rect 8003 4534 8032 4538
rect 7922 4533 8032 4534
rect 7922 4532 8038 4533
rect 7597 4524 7648 4532
rect 7597 4512 7622 4524
rect 7629 4512 7648 4524
rect 7679 4524 7729 4532
rect 7679 4516 7695 4524
rect 7702 4522 7729 4524
rect 7738 4522 7959 4532
rect 7702 4512 7959 4522
rect 7988 4524 8038 4532
rect 7988 4515 8004 4524
rect 7597 4504 7648 4512
rect 7695 4504 7959 4512
rect 7985 4512 8004 4515
rect 8011 4512 8038 4524
rect 7985 4504 8038 4512
rect 7613 4496 7614 4504
rect 7629 4496 7642 4504
rect 7613 4488 7629 4496
rect 7610 4481 7629 4484
rect 7610 4472 7632 4481
rect 7583 4462 7632 4472
rect 7583 4456 7613 4462
rect 7632 4457 7637 4462
rect 7555 4440 7629 4456
rect 7647 4448 7677 4504
rect 7712 4494 7920 4504
rect 7955 4500 8000 4504
rect 8003 4503 8004 4504
rect 8019 4503 8032 4504
rect 7738 4464 7927 4494
rect 7753 4461 7927 4464
rect 7746 4458 7927 4461
rect 7555 4438 7568 4440
rect 7583 4438 7617 4440
rect 7555 4422 7629 4438
rect 7656 4434 7669 4448
rect 7684 4434 7700 4450
rect 7746 4445 7757 4458
rect 7539 4400 7540 4416
rect 7555 4400 7568 4422
rect 7583 4400 7613 4422
rect 7656 4418 7718 4434
rect 7746 4427 7757 4443
rect 7762 4438 7772 4458
rect 7782 4438 7796 4458
rect 7799 4445 7808 4458
rect 7824 4445 7833 4458
rect 7762 4427 7796 4438
rect 7799 4427 7808 4443
rect 7824 4427 7833 4443
rect 7840 4438 7850 4458
rect 7860 4438 7874 4458
rect 7875 4445 7886 4458
rect 7840 4427 7874 4438
rect 7875 4427 7886 4443
rect 7932 4434 7948 4450
rect 7955 4448 7985 4500
rect 8019 4496 8020 4503
rect 8004 4488 8020 4496
rect 7991 4456 8004 4475
rect 8019 4456 8049 4472
rect 7991 4440 8065 4456
rect 7991 4438 8004 4440
rect 8019 4438 8053 4440
rect 7656 4416 7669 4418
rect 7684 4416 7718 4418
rect 7656 4400 7718 4416
rect 7762 4411 7778 4414
rect 7840 4411 7870 4422
rect 7918 4418 7964 4434
rect 7991 4422 8065 4438
rect 7918 4416 7952 4418
rect 7917 4400 7964 4416
rect 7991 4400 8004 4422
rect 8019 4400 8049 4422
rect 8076 4400 8077 4416
rect 8092 4400 8105 4560
rect 8135 4456 8148 4560
rect 8193 4538 8194 4548
rect 8209 4538 8222 4548
rect 8193 4534 8222 4538
rect 8227 4534 8257 4560
rect 8275 4546 8291 4548
rect 8363 4546 8416 4560
rect 8364 4544 8428 4546
rect 8471 4544 8486 4560
rect 8535 4557 8565 4560
rect 8535 4554 8571 4557
rect 8501 4546 8517 4548
rect 8275 4534 8290 4538
rect 8193 4532 8290 4534
rect 8318 4532 8486 4544
rect 8502 4534 8517 4538
rect 8535 4535 8574 4554
rect 8593 4548 8600 4549
rect 8599 4541 8600 4548
rect 8583 4538 8584 4541
rect 8599 4538 8612 4541
rect 8535 4534 8565 4535
rect 8574 4534 8580 4535
rect 8583 4534 8612 4538
rect 8502 4533 8612 4534
rect 8502 4532 8618 4533
rect 8177 4524 8228 4532
rect 8177 4512 8202 4524
rect 8209 4512 8228 4524
rect 8259 4524 8309 4532
rect 8259 4516 8275 4524
rect 8282 4522 8309 4524
rect 8318 4522 8539 4532
rect 8282 4512 8539 4522
rect 8568 4524 8618 4532
rect 8568 4515 8584 4524
rect 8177 4504 8228 4512
rect 8275 4504 8539 4512
rect 8565 4512 8584 4515
rect 8591 4512 8618 4524
rect 8565 4504 8618 4512
rect 8193 4496 8194 4504
rect 8209 4496 8222 4504
rect 8193 4488 8209 4496
rect 8190 4481 8209 4484
rect 8190 4472 8212 4481
rect 8163 4462 8212 4472
rect 8163 4456 8193 4462
rect 8212 4457 8217 4462
rect 8135 4440 8209 4456
rect 8227 4448 8257 4504
rect 8292 4494 8500 4504
rect 8535 4500 8580 4504
rect 8583 4503 8584 4504
rect 8599 4503 8612 4504
rect 8318 4464 8507 4494
rect 8333 4461 8507 4464
rect 8326 4458 8507 4461
rect 8135 4438 8148 4440
rect 8163 4438 8197 4440
rect 8135 4422 8209 4438
rect 8236 4434 8249 4448
rect 8264 4434 8280 4450
rect 8326 4445 8337 4458
rect 8119 4400 8120 4416
rect 8135 4400 8148 4422
rect 8163 4400 8193 4422
rect 8236 4418 8298 4434
rect 8326 4427 8337 4443
rect 8342 4438 8352 4458
rect 8362 4438 8376 4458
rect 8379 4445 8388 4458
rect 8404 4445 8413 4458
rect 8342 4427 8376 4438
rect 8379 4427 8388 4443
rect 8404 4427 8413 4443
rect 8420 4438 8430 4458
rect 8440 4438 8454 4458
rect 8455 4445 8466 4458
rect 8420 4427 8454 4438
rect 8455 4427 8466 4443
rect 8512 4434 8528 4450
rect 8535 4448 8565 4500
rect 8599 4496 8600 4503
rect 8584 4488 8600 4496
rect 8571 4456 8584 4475
rect 8599 4456 8629 4472
rect 8571 4440 8645 4456
rect 8571 4438 8584 4440
rect 8599 4438 8633 4440
rect 8236 4416 8249 4418
rect 8264 4416 8298 4418
rect 8236 4400 8298 4416
rect 8342 4411 8358 4414
rect 8420 4411 8450 4422
rect 8498 4418 8544 4434
rect 8571 4422 8645 4438
rect 8498 4416 8532 4418
rect 8497 4400 8544 4416
rect 8571 4400 8584 4422
rect 8599 4400 8629 4422
rect 8656 4400 8657 4416
rect 8672 4400 8685 4560
rect 8715 4456 8728 4560
rect 8773 4538 8774 4548
rect 8789 4538 8802 4548
rect 8773 4534 8802 4538
rect 8807 4534 8837 4560
rect 8855 4546 8871 4548
rect 8943 4546 8996 4560
rect 8944 4544 9008 4546
rect 9051 4544 9066 4560
rect 9115 4557 9145 4560
rect 9115 4554 9151 4557
rect 9081 4546 9097 4548
rect 8855 4534 8870 4538
rect 8773 4532 8870 4534
rect 8898 4532 9066 4544
rect 9082 4534 9097 4538
rect 9115 4535 9154 4554
rect 9173 4548 9180 4549
rect 9179 4541 9180 4548
rect 9163 4538 9164 4541
rect 9179 4538 9192 4541
rect 9115 4534 9145 4535
rect 9154 4534 9160 4535
rect 9163 4534 9192 4538
rect 9082 4533 9192 4534
rect 9082 4532 9198 4533
rect 8757 4524 8808 4532
rect 8757 4512 8782 4524
rect 8789 4512 8808 4524
rect 8839 4524 8889 4532
rect 8839 4516 8855 4524
rect 8862 4522 8889 4524
rect 8898 4522 9119 4532
rect 8862 4512 9119 4522
rect 9148 4524 9198 4532
rect 9148 4515 9164 4524
rect 8757 4504 8808 4512
rect 8855 4504 9119 4512
rect 9145 4512 9164 4515
rect 9171 4512 9198 4524
rect 9145 4504 9198 4512
rect 8773 4496 8774 4504
rect 8789 4496 8802 4504
rect 8773 4488 8789 4496
rect 8770 4481 8789 4484
rect 8770 4472 8792 4481
rect 8743 4462 8792 4472
rect 8743 4456 8773 4462
rect 8792 4457 8797 4462
rect 8715 4440 8789 4456
rect 8807 4448 8837 4504
rect 8872 4494 9080 4504
rect 9115 4500 9160 4504
rect 9163 4503 9164 4504
rect 9179 4503 9192 4504
rect 8898 4464 9087 4494
rect 8913 4461 9087 4464
rect 8906 4458 9087 4461
rect 8715 4438 8728 4440
rect 8743 4438 8777 4440
rect 8715 4422 8789 4438
rect 8816 4434 8829 4448
rect 8844 4434 8860 4450
rect 8906 4445 8917 4458
rect 8699 4400 8700 4416
rect 8715 4400 8728 4422
rect 8743 4400 8773 4422
rect 8816 4418 8878 4434
rect 8906 4427 8917 4443
rect 8922 4438 8932 4458
rect 8942 4438 8956 4458
rect 8959 4445 8968 4458
rect 8984 4445 8993 4458
rect 8922 4427 8956 4438
rect 8959 4427 8968 4443
rect 8984 4427 8993 4443
rect 9000 4438 9010 4458
rect 9020 4438 9034 4458
rect 9035 4445 9046 4458
rect 9000 4427 9034 4438
rect 9035 4427 9046 4443
rect 9092 4434 9108 4450
rect 9115 4448 9145 4500
rect 9179 4496 9180 4503
rect 9164 4488 9180 4496
rect 9151 4456 9164 4475
rect 9179 4456 9209 4472
rect 9151 4440 9225 4456
rect 9151 4438 9164 4440
rect 9179 4438 9213 4440
rect 8816 4416 8829 4418
rect 8844 4416 8878 4418
rect 8816 4400 8878 4416
rect 8922 4411 8938 4414
rect 9000 4411 9030 4422
rect 9078 4418 9124 4434
rect 9151 4422 9225 4438
rect 9078 4416 9112 4418
rect 9077 4400 9124 4416
rect 9151 4400 9164 4422
rect 9179 4400 9209 4422
rect 9236 4400 9237 4416
rect 9252 4400 9265 4560
rect -7 4392 34 4400
rect -7 4366 8 4392
rect 15 4366 34 4392
rect 98 4388 160 4400
rect 172 4388 247 4400
rect 305 4388 380 4400
rect 392 4388 423 4400
rect 429 4388 464 4400
rect 98 4386 260 4388
rect -7 4358 34 4366
rect 116 4362 129 4386
rect 144 4384 159 4386
rect -1 4348 0 4358
rect 15 4348 28 4358
rect 43 4348 73 4362
rect 116 4348 159 4362
rect 183 4359 190 4366
rect 193 4362 260 4386
rect 292 4386 464 4388
rect 262 4364 290 4368
rect 292 4364 372 4386
rect 393 4384 408 4386
rect 262 4362 372 4364
rect 193 4358 372 4362
rect 166 4348 196 4358
rect 198 4348 351 4358
rect 359 4348 389 4358
rect 393 4348 423 4362
rect 451 4348 464 4386
rect 536 4392 571 4400
rect 536 4366 537 4392
rect 544 4366 571 4392
rect 479 4348 509 4362
rect 536 4358 571 4366
rect 573 4392 614 4400
rect 573 4366 588 4392
rect 595 4366 614 4392
rect 678 4388 740 4400
rect 752 4388 827 4400
rect 885 4388 960 4400
rect 972 4388 1003 4400
rect 1009 4388 1044 4400
rect 678 4386 840 4388
rect 573 4358 614 4366
rect 696 4362 709 4386
rect 724 4384 739 4386
rect 536 4348 537 4358
rect 552 4348 565 4358
rect 579 4348 580 4358
rect 595 4348 608 4358
rect 623 4348 653 4362
rect 696 4348 739 4362
rect 763 4359 770 4366
rect 773 4362 840 4386
rect 872 4386 1044 4388
rect 842 4364 870 4368
rect 872 4364 952 4386
rect 973 4384 988 4386
rect 842 4362 952 4364
rect 773 4358 952 4362
rect 746 4348 776 4358
rect 778 4348 931 4358
rect 939 4348 969 4358
rect 973 4348 1003 4362
rect 1031 4348 1044 4386
rect 1116 4392 1151 4400
rect 1116 4366 1117 4392
rect 1124 4366 1151 4392
rect 1059 4348 1089 4362
rect 1116 4358 1151 4366
rect 1153 4392 1194 4400
rect 1153 4366 1168 4392
rect 1175 4366 1194 4392
rect 1258 4388 1320 4400
rect 1332 4388 1407 4400
rect 1465 4388 1540 4400
rect 1552 4388 1583 4400
rect 1589 4388 1624 4400
rect 1258 4386 1420 4388
rect 1153 4358 1194 4366
rect 1276 4362 1289 4386
rect 1304 4384 1319 4386
rect 1116 4348 1117 4358
rect 1132 4348 1145 4358
rect 1159 4348 1160 4358
rect 1175 4348 1188 4358
rect 1203 4348 1233 4362
rect 1276 4348 1319 4362
rect 1343 4359 1350 4366
rect 1353 4362 1420 4386
rect 1452 4386 1624 4388
rect 1422 4364 1450 4368
rect 1452 4364 1532 4386
rect 1553 4384 1568 4386
rect 1422 4362 1532 4364
rect 1353 4358 1532 4362
rect 1326 4348 1356 4358
rect 1358 4348 1511 4358
rect 1519 4348 1549 4358
rect 1553 4348 1583 4362
rect 1611 4348 1624 4386
rect 1696 4392 1731 4400
rect 1696 4366 1697 4392
rect 1704 4366 1731 4392
rect 1639 4348 1669 4362
rect 1696 4358 1731 4366
rect 1733 4392 1774 4400
rect 1733 4366 1748 4392
rect 1755 4366 1774 4392
rect 1838 4388 1900 4400
rect 1912 4388 1987 4400
rect 2045 4388 2120 4400
rect 2132 4388 2163 4400
rect 2169 4388 2204 4400
rect 1838 4386 2000 4388
rect 1733 4358 1774 4366
rect 1856 4362 1869 4386
rect 1884 4384 1899 4386
rect 1696 4348 1697 4358
rect 1712 4348 1725 4358
rect 1739 4348 1740 4358
rect 1755 4348 1768 4358
rect 1783 4348 1813 4362
rect 1856 4348 1899 4362
rect 1923 4359 1930 4366
rect 1933 4362 2000 4386
rect 2032 4386 2204 4388
rect 2002 4364 2030 4368
rect 2032 4364 2112 4386
rect 2133 4384 2148 4386
rect 2002 4362 2112 4364
rect 1933 4358 2112 4362
rect 1906 4348 1936 4358
rect 1938 4348 2091 4358
rect 2099 4348 2129 4358
rect 2133 4348 2163 4362
rect 2191 4348 2204 4386
rect 2276 4392 2311 4400
rect 2276 4366 2277 4392
rect 2284 4366 2311 4392
rect 2219 4348 2249 4362
rect 2276 4358 2311 4366
rect 2313 4392 2354 4400
rect 2313 4366 2328 4392
rect 2335 4366 2354 4392
rect 2418 4388 2480 4400
rect 2492 4388 2567 4400
rect 2625 4388 2700 4400
rect 2712 4388 2743 4400
rect 2749 4388 2784 4400
rect 2418 4386 2580 4388
rect 2313 4358 2354 4366
rect 2436 4362 2449 4386
rect 2464 4384 2479 4386
rect 2276 4348 2277 4358
rect 2292 4348 2305 4358
rect 2319 4348 2320 4358
rect 2335 4348 2348 4358
rect 2363 4348 2393 4362
rect 2436 4348 2479 4362
rect 2503 4359 2510 4366
rect 2513 4362 2580 4386
rect 2612 4386 2784 4388
rect 2582 4364 2610 4368
rect 2612 4364 2692 4386
rect 2713 4384 2728 4386
rect 2582 4362 2692 4364
rect 2513 4358 2692 4362
rect 2486 4348 2516 4358
rect 2518 4348 2671 4358
rect 2679 4348 2709 4358
rect 2713 4348 2743 4362
rect 2771 4348 2784 4386
rect 2856 4392 2891 4400
rect 2856 4366 2857 4392
rect 2864 4366 2891 4392
rect 2799 4348 2829 4362
rect 2856 4358 2891 4366
rect 2893 4392 2934 4400
rect 2893 4366 2908 4392
rect 2915 4366 2934 4392
rect 2998 4388 3060 4400
rect 3072 4388 3147 4400
rect 3205 4388 3280 4400
rect 3292 4388 3323 4400
rect 3329 4388 3364 4400
rect 2998 4386 3160 4388
rect 2893 4358 2934 4366
rect 3016 4362 3029 4386
rect 3044 4384 3059 4386
rect 2856 4348 2857 4358
rect 2872 4348 2885 4358
rect 2899 4348 2900 4358
rect 2915 4348 2928 4358
rect 2943 4348 2973 4362
rect 3016 4348 3059 4362
rect 3083 4359 3090 4366
rect 3093 4362 3160 4386
rect 3192 4386 3364 4388
rect 3162 4364 3190 4368
rect 3192 4364 3272 4386
rect 3293 4384 3308 4386
rect 3162 4362 3272 4364
rect 3093 4358 3272 4362
rect 3066 4348 3096 4358
rect 3098 4348 3251 4358
rect 3259 4348 3289 4358
rect 3293 4348 3323 4362
rect 3351 4348 3364 4386
rect 3436 4392 3471 4400
rect 3436 4366 3437 4392
rect 3444 4366 3471 4392
rect 3379 4348 3409 4362
rect 3436 4358 3471 4366
rect 3473 4392 3514 4400
rect 3473 4366 3488 4392
rect 3495 4366 3514 4392
rect 3578 4388 3640 4400
rect 3652 4388 3727 4400
rect 3785 4388 3860 4400
rect 3872 4388 3903 4400
rect 3909 4388 3944 4400
rect 3578 4386 3740 4388
rect 3473 4358 3514 4366
rect 3596 4362 3609 4386
rect 3624 4384 3639 4386
rect 3436 4348 3437 4358
rect 3452 4348 3465 4358
rect 3479 4348 3480 4358
rect 3495 4348 3508 4358
rect 3523 4348 3553 4362
rect 3596 4348 3639 4362
rect 3663 4359 3670 4366
rect 3673 4362 3740 4386
rect 3772 4386 3944 4388
rect 3742 4364 3770 4368
rect 3772 4364 3852 4386
rect 3873 4384 3888 4386
rect 3742 4362 3852 4364
rect 3673 4358 3852 4362
rect 3646 4348 3676 4358
rect 3678 4348 3831 4358
rect 3839 4348 3869 4358
rect 3873 4348 3903 4362
rect 3931 4348 3944 4386
rect 4016 4392 4051 4400
rect 4016 4366 4017 4392
rect 4024 4366 4051 4392
rect 3959 4348 3989 4362
rect 4016 4358 4051 4366
rect 4053 4392 4094 4400
rect 4053 4366 4068 4392
rect 4075 4366 4094 4392
rect 4158 4388 4220 4400
rect 4232 4388 4307 4400
rect 4365 4388 4440 4400
rect 4452 4388 4483 4400
rect 4489 4388 4524 4400
rect 4158 4386 4320 4388
rect 4053 4358 4094 4366
rect 4176 4362 4189 4386
rect 4204 4384 4219 4386
rect 4016 4348 4017 4358
rect 4032 4348 4045 4358
rect 4059 4348 4060 4358
rect 4075 4348 4088 4358
rect 4103 4348 4133 4362
rect 4176 4348 4219 4362
rect 4243 4359 4250 4366
rect 4253 4362 4320 4386
rect 4352 4386 4524 4388
rect 4322 4364 4350 4368
rect 4352 4364 4432 4386
rect 4453 4384 4468 4386
rect 4322 4362 4432 4364
rect 4253 4358 4432 4362
rect 4226 4348 4256 4358
rect 4258 4348 4411 4358
rect 4419 4348 4449 4358
rect 4453 4348 4483 4362
rect 4511 4348 4524 4386
rect 4596 4392 4631 4400
rect 4596 4366 4597 4392
rect 4604 4366 4631 4392
rect 4539 4348 4569 4362
rect 4596 4358 4631 4366
rect 4633 4392 4674 4400
rect 4633 4366 4648 4392
rect 4655 4366 4674 4392
rect 4738 4388 4800 4400
rect 4812 4388 4887 4400
rect 4945 4388 5020 4400
rect 5032 4388 5063 4400
rect 5069 4388 5104 4400
rect 4738 4386 4900 4388
rect 4633 4358 4674 4366
rect 4756 4362 4769 4386
rect 4784 4384 4799 4386
rect 4596 4348 4597 4358
rect 4612 4348 4625 4358
rect 4639 4348 4640 4358
rect 4655 4348 4668 4358
rect 4683 4348 4713 4362
rect 4756 4348 4799 4362
rect 4823 4359 4830 4366
rect 4833 4362 4900 4386
rect 4932 4386 5104 4388
rect 4902 4364 4930 4368
rect 4932 4364 5012 4386
rect 5033 4384 5048 4386
rect 4902 4362 5012 4364
rect 4833 4358 5012 4362
rect 4806 4348 4836 4358
rect 4838 4348 4991 4358
rect 4999 4348 5029 4358
rect 5033 4348 5063 4362
rect 5091 4348 5104 4386
rect 5176 4392 5211 4400
rect 5176 4366 5177 4392
rect 5184 4366 5211 4392
rect 5119 4348 5149 4362
rect 5176 4358 5211 4366
rect 5213 4392 5254 4400
rect 5213 4366 5228 4392
rect 5235 4366 5254 4392
rect 5318 4388 5380 4400
rect 5392 4388 5467 4400
rect 5525 4388 5600 4400
rect 5612 4388 5643 4400
rect 5649 4388 5684 4400
rect 5318 4386 5480 4388
rect 5213 4358 5254 4366
rect 5336 4362 5349 4386
rect 5364 4384 5379 4386
rect 5176 4348 5177 4358
rect 5192 4348 5205 4358
rect 5219 4348 5220 4358
rect 5235 4348 5248 4358
rect 5263 4348 5293 4362
rect 5336 4348 5379 4362
rect 5403 4359 5410 4366
rect 5413 4362 5480 4386
rect 5512 4386 5684 4388
rect 5482 4364 5510 4368
rect 5512 4364 5592 4386
rect 5613 4384 5628 4386
rect 5482 4362 5592 4364
rect 5413 4358 5592 4362
rect 5386 4348 5416 4358
rect 5418 4348 5571 4358
rect 5579 4348 5609 4358
rect 5613 4348 5643 4362
rect 5671 4348 5684 4386
rect 5756 4392 5791 4400
rect 5756 4366 5757 4392
rect 5764 4366 5791 4392
rect 5699 4348 5729 4362
rect 5756 4358 5791 4366
rect 5793 4392 5834 4400
rect 5793 4366 5808 4392
rect 5815 4366 5834 4392
rect 5898 4388 5960 4400
rect 5972 4388 6047 4400
rect 6105 4388 6180 4400
rect 6192 4388 6223 4400
rect 6229 4388 6264 4400
rect 5898 4386 6060 4388
rect 5793 4358 5834 4366
rect 5916 4362 5929 4386
rect 5944 4384 5959 4386
rect 5756 4348 5757 4358
rect 5772 4348 5785 4358
rect 5799 4348 5800 4358
rect 5815 4348 5828 4358
rect 5843 4348 5873 4362
rect 5916 4348 5959 4362
rect 5983 4359 5990 4366
rect 5993 4362 6060 4386
rect 6092 4386 6264 4388
rect 6062 4364 6090 4368
rect 6092 4364 6172 4386
rect 6193 4384 6208 4386
rect 6062 4362 6172 4364
rect 5993 4358 6172 4362
rect 5966 4348 5996 4358
rect 5998 4348 6151 4358
rect 6159 4348 6189 4358
rect 6193 4348 6223 4362
rect 6251 4348 6264 4386
rect 6336 4392 6371 4400
rect 6336 4366 6337 4392
rect 6344 4366 6371 4392
rect 6279 4348 6309 4362
rect 6336 4358 6371 4366
rect 6373 4392 6414 4400
rect 6373 4366 6388 4392
rect 6395 4366 6414 4392
rect 6478 4388 6540 4400
rect 6552 4388 6627 4400
rect 6685 4388 6760 4400
rect 6772 4388 6803 4400
rect 6809 4388 6844 4400
rect 6478 4386 6640 4388
rect 6373 4358 6414 4366
rect 6496 4362 6509 4386
rect 6524 4384 6539 4386
rect 6336 4348 6337 4358
rect 6352 4348 6365 4358
rect 6379 4348 6380 4358
rect 6395 4348 6408 4358
rect 6423 4348 6453 4362
rect 6496 4348 6539 4362
rect 6563 4359 6570 4366
rect 6573 4362 6640 4386
rect 6672 4386 6844 4388
rect 6642 4364 6670 4368
rect 6672 4364 6752 4386
rect 6773 4384 6788 4386
rect 6642 4362 6752 4364
rect 6573 4358 6752 4362
rect 6546 4348 6576 4358
rect 6578 4348 6731 4358
rect 6739 4348 6769 4358
rect 6773 4348 6803 4362
rect 6831 4348 6844 4386
rect 6916 4392 6951 4400
rect 6916 4366 6917 4392
rect 6924 4366 6951 4392
rect 6859 4348 6889 4362
rect 6916 4358 6951 4366
rect 6953 4392 6994 4400
rect 6953 4366 6968 4392
rect 6975 4366 6994 4392
rect 7058 4388 7120 4400
rect 7132 4388 7207 4400
rect 7265 4388 7340 4400
rect 7352 4388 7383 4400
rect 7389 4388 7424 4400
rect 7058 4386 7220 4388
rect 6953 4358 6994 4366
rect 7076 4362 7089 4386
rect 7104 4384 7119 4386
rect 6916 4348 6917 4358
rect 6932 4348 6945 4358
rect 6959 4348 6960 4358
rect 6975 4348 6988 4358
rect 7003 4348 7033 4362
rect 7076 4348 7119 4362
rect 7143 4359 7150 4366
rect 7153 4362 7220 4386
rect 7252 4386 7424 4388
rect 7222 4364 7250 4368
rect 7252 4364 7332 4386
rect 7353 4384 7368 4386
rect 7222 4362 7332 4364
rect 7153 4358 7332 4362
rect 7126 4348 7156 4358
rect 7158 4348 7311 4358
rect 7319 4348 7349 4358
rect 7353 4348 7383 4362
rect 7411 4348 7424 4386
rect 7496 4392 7531 4400
rect 7496 4366 7497 4392
rect 7504 4366 7531 4392
rect 7439 4348 7469 4362
rect 7496 4358 7531 4366
rect 7533 4392 7574 4400
rect 7533 4366 7548 4392
rect 7555 4366 7574 4392
rect 7638 4388 7700 4400
rect 7712 4388 7787 4400
rect 7845 4388 7920 4400
rect 7932 4388 7963 4400
rect 7969 4388 8004 4400
rect 7638 4386 7800 4388
rect 7533 4358 7574 4366
rect 7656 4362 7669 4386
rect 7684 4384 7699 4386
rect 7496 4348 7497 4358
rect 7512 4348 7525 4358
rect 7539 4348 7540 4358
rect 7555 4348 7568 4358
rect 7583 4348 7613 4362
rect 7656 4348 7699 4362
rect 7723 4359 7730 4366
rect 7733 4362 7800 4386
rect 7832 4386 8004 4388
rect 7802 4364 7830 4368
rect 7832 4364 7912 4386
rect 7933 4384 7948 4386
rect 7802 4362 7912 4364
rect 7733 4358 7912 4362
rect 7706 4348 7736 4358
rect 7738 4348 7891 4358
rect 7899 4348 7929 4358
rect 7933 4348 7963 4362
rect 7991 4348 8004 4386
rect 8076 4392 8111 4400
rect 8076 4366 8077 4392
rect 8084 4366 8111 4392
rect 8019 4348 8049 4362
rect 8076 4358 8111 4366
rect 8113 4392 8154 4400
rect 8113 4366 8128 4392
rect 8135 4366 8154 4392
rect 8218 4388 8280 4400
rect 8292 4388 8367 4400
rect 8425 4388 8500 4400
rect 8512 4388 8543 4400
rect 8549 4388 8584 4400
rect 8218 4386 8380 4388
rect 8113 4358 8154 4366
rect 8236 4362 8249 4386
rect 8264 4384 8279 4386
rect 8076 4348 8077 4358
rect 8092 4348 8105 4358
rect 8119 4348 8120 4358
rect 8135 4348 8148 4358
rect 8163 4348 8193 4362
rect 8236 4348 8279 4362
rect 8303 4359 8310 4366
rect 8313 4362 8380 4386
rect 8412 4386 8584 4388
rect 8382 4364 8410 4368
rect 8412 4364 8492 4386
rect 8513 4384 8528 4386
rect 8382 4362 8492 4364
rect 8313 4358 8492 4362
rect 8286 4348 8316 4358
rect 8318 4348 8471 4358
rect 8479 4348 8509 4358
rect 8513 4348 8543 4362
rect 8571 4348 8584 4386
rect 8656 4392 8691 4400
rect 8656 4366 8657 4392
rect 8664 4366 8691 4392
rect 8599 4348 8629 4362
rect 8656 4358 8691 4366
rect 8693 4392 8734 4400
rect 8693 4366 8708 4392
rect 8715 4366 8734 4392
rect 8798 4388 8860 4400
rect 8872 4388 8947 4400
rect 9005 4388 9080 4400
rect 9092 4388 9123 4400
rect 9129 4388 9164 4400
rect 8798 4386 8960 4388
rect 8693 4358 8734 4366
rect 8816 4362 8829 4386
rect 8844 4384 8859 4386
rect 8656 4348 8657 4358
rect 8672 4348 8685 4358
rect 8699 4348 8700 4358
rect 8715 4348 8728 4358
rect 8743 4348 8773 4362
rect 8816 4348 8859 4362
rect 8883 4359 8890 4366
rect 8893 4362 8960 4386
rect 8992 4386 9164 4388
rect 8962 4364 8990 4368
rect 8992 4364 9072 4386
rect 9093 4384 9108 4386
rect 8962 4362 9072 4364
rect 8893 4358 9072 4362
rect 8866 4348 8896 4358
rect 8898 4348 9051 4358
rect 9059 4348 9089 4358
rect 9093 4348 9123 4362
rect 9151 4348 9164 4386
rect 9236 4392 9271 4400
rect 9236 4366 9237 4392
rect 9244 4366 9271 4392
rect 9179 4348 9209 4362
rect 9236 4358 9271 4366
rect 9236 4348 9237 4358
rect 9252 4348 9265 4358
rect -1 4342 9265 4348
rect 0 4334 9265 4342
rect 15 4304 28 4334
rect 43 4316 73 4334
rect 116 4320 130 4334
rect 166 4320 386 4334
rect 117 4318 130 4320
rect 83 4306 98 4318
rect 80 4304 102 4306
rect 107 4304 137 4318
rect 198 4316 351 4320
rect 180 4304 372 4316
rect 415 4304 445 4318
rect 451 4304 464 4334
rect 479 4316 509 4334
rect 552 4304 565 4334
rect 595 4304 608 4334
rect 623 4316 653 4334
rect 696 4320 710 4334
rect 746 4320 966 4334
rect 697 4318 710 4320
rect 663 4306 678 4318
rect 660 4304 682 4306
rect 687 4304 717 4318
rect 778 4316 931 4320
rect 760 4304 952 4316
rect 995 4304 1025 4318
rect 1031 4304 1044 4334
rect 1059 4316 1089 4334
rect 1132 4304 1145 4334
rect 1175 4304 1188 4334
rect 1203 4316 1233 4334
rect 1276 4320 1290 4334
rect 1326 4320 1546 4334
rect 1277 4318 1290 4320
rect 1243 4306 1258 4318
rect 1240 4304 1262 4306
rect 1267 4304 1297 4318
rect 1358 4316 1511 4320
rect 1340 4304 1532 4316
rect 1575 4304 1605 4318
rect 1611 4304 1624 4334
rect 1639 4316 1669 4334
rect 1712 4304 1725 4334
rect 1755 4304 1768 4334
rect 1783 4316 1813 4334
rect 1856 4320 1870 4334
rect 1906 4320 2126 4334
rect 1857 4318 1870 4320
rect 1823 4306 1838 4318
rect 1820 4304 1842 4306
rect 1847 4304 1877 4318
rect 1938 4316 2091 4320
rect 1920 4304 2112 4316
rect 2155 4304 2185 4318
rect 2191 4304 2204 4334
rect 2219 4316 2249 4334
rect 2292 4304 2305 4334
rect 2335 4304 2348 4334
rect 2363 4316 2393 4334
rect 2436 4320 2450 4334
rect 2486 4320 2706 4334
rect 2437 4318 2450 4320
rect 2403 4306 2418 4318
rect 2400 4304 2422 4306
rect 2427 4304 2457 4318
rect 2518 4316 2671 4320
rect 2500 4304 2692 4316
rect 2735 4304 2765 4318
rect 2771 4304 2784 4334
rect 2799 4316 2829 4334
rect 2872 4304 2885 4334
rect 2915 4304 2928 4334
rect 2943 4316 2973 4334
rect 3016 4320 3030 4334
rect 3066 4320 3286 4334
rect 3017 4318 3030 4320
rect 2983 4306 2998 4318
rect 2980 4304 3002 4306
rect 3007 4304 3037 4318
rect 3098 4316 3251 4320
rect 3080 4304 3272 4316
rect 3315 4304 3345 4318
rect 3351 4304 3364 4334
rect 3379 4316 3409 4334
rect 3452 4304 3465 4334
rect 3495 4304 3508 4334
rect 3523 4316 3553 4334
rect 3596 4320 3610 4334
rect 3646 4320 3866 4334
rect 3597 4318 3610 4320
rect 3563 4306 3578 4318
rect 3560 4304 3582 4306
rect 3587 4304 3617 4318
rect 3678 4316 3831 4320
rect 3660 4304 3852 4316
rect 3895 4304 3925 4318
rect 3931 4304 3944 4334
rect 3959 4316 3989 4334
rect 4032 4304 4045 4334
rect 4075 4304 4088 4334
rect 4103 4316 4133 4334
rect 4176 4320 4190 4334
rect 4226 4320 4446 4334
rect 4177 4318 4190 4320
rect 4143 4306 4158 4318
rect 4140 4304 4162 4306
rect 4167 4304 4197 4318
rect 4258 4316 4411 4320
rect 4240 4304 4432 4316
rect 4475 4304 4505 4318
rect 4511 4304 4524 4334
rect 4539 4316 4569 4334
rect 4612 4304 4625 4334
rect 4655 4304 4668 4334
rect 4683 4316 4713 4334
rect 4756 4320 4770 4334
rect 4806 4320 5026 4334
rect 4757 4318 4770 4320
rect 4723 4306 4738 4318
rect 4720 4304 4742 4306
rect 4747 4304 4777 4318
rect 4838 4316 4991 4320
rect 4820 4304 5012 4316
rect 5055 4304 5085 4318
rect 5091 4304 5104 4334
rect 5119 4316 5149 4334
rect 5192 4304 5205 4334
rect 5235 4304 5248 4334
rect 5263 4316 5293 4334
rect 5336 4320 5350 4334
rect 5386 4320 5606 4334
rect 5337 4318 5350 4320
rect 5303 4306 5318 4318
rect 5300 4304 5322 4306
rect 5327 4304 5357 4318
rect 5418 4316 5571 4320
rect 5400 4304 5592 4316
rect 5635 4304 5665 4318
rect 5671 4304 5684 4334
rect 5699 4316 5729 4334
rect 5772 4304 5785 4334
rect 5815 4304 5828 4334
rect 5843 4316 5873 4334
rect 5916 4320 5930 4334
rect 5966 4320 6186 4334
rect 5917 4318 5930 4320
rect 5883 4306 5898 4318
rect 5880 4304 5902 4306
rect 5907 4304 5937 4318
rect 5998 4316 6151 4320
rect 5980 4304 6172 4316
rect 6215 4304 6245 4318
rect 6251 4304 6264 4334
rect 6279 4316 6309 4334
rect 6352 4304 6365 4334
rect 6395 4304 6408 4334
rect 6423 4316 6453 4334
rect 6496 4320 6510 4334
rect 6546 4320 6766 4334
rect 6497 4318 6510 4320
rect 6463 4306 6478 4318
rect 6460 4304 6482 4306
rect 6487 4304 6517 4318
rect 6578 4316 6731 4320
rect 6560 4304 6752 4316
rect 6795 4304 6825 4318
rect 6831 4304 6844 4334
rect 6859 4316 6889 4334
rect 6932 4304 6945 4334
rect 6975 4304 6988 4334
rect 7003 4316 7033 4334
rect 7076 4320 7090 4334
rect 7126 4320 7346 4334
rect 7077 4318 7090 4320
rect 7043 4306 7058 4318
rect 7040 4304 7062 4306
rect 7067 4304 7097 4318
rect 7158 4316 7311 4320
rect 7140 4304 7332 4316
rect 7375 4304 7405 4318
rect 7411 4304 7424 4334
rect 7439 4316 7469 4334
rect 7512 4304 7525 4334
rect 7555 4304 7568 4334
rect 7583 4316 7613 4334
rect 7656 4320 7670 4334
rect 7706 4320 7926 4334
rect 7657 4318 7670 4320
rect 7623 4306 7638 4318
rect 7620 4304 7642 4306
rect 7647 4304 7677 4318
rect 7738 4316 7891 4320
rect 7720 4304 7912 4316
rect 7955 4304 7985 4318
rect 7991 4304 8004 4334
rect 8019 4316 8049 4334
rect 8092 4304 8105 4334
rect 8135 4304 8148 4334
rect 8163 4316 8193 4334
rect 8236 4320 8250 4334
rect 8286 4320 8506 4334
rect 8237 4318 8250 4320
rect 8203 4306 8218 4318
rect 8200 4304 8222 4306
rect 8227 4304 8257 4318
rect 8318 4316 8471 4320
rect 8300 4304 8492 4316
rect 8535 4304 8565 4318
rect 8571 4304 8584 4334
rect 8599 4316 8629 4334
rect 8672 4304 8685 4334
rect 8715 4304 8728 4334
rect 8743 4316 8773 4334
rect 8816 4320 8830 4334
rect 8866 4320 9086 4334
rect 8817 4318 8830 4320
rect 8783 4306 8798 4318
rect 8780 4304 8802 4306
rect 8807 4304 8837 4318
rect 8898 4316 9051 4320
rect 8880 4304 9072 4316
rect 9115 4304 9145 4318
rect 9151 4304 9164 4334
rect 9179 4316 9209 4334
rect 9252 4304 9265 4334
rect 0 4290 9265 4304
rect 15 4186 28 4290
rect 73 4268 74 4278
rect 89 4268 102 4278
rect 73 4264 102 4268
rect 107 4264 137 4290
rect 155 4276 171 4278
rect 243 4276 296 4290
rect 244 4274 308 4276
rect 351 4274 366 4290
rect 415 4287 445 4290
rect 415 4284 451 4287
rect 381 4276 397 4278
rect 155 4264 170 4268
rect 73 4262 170 4264
rect 198 4262 366 4274
rect 382 4264 397 4268
rect 415 4265 454 4284
rect 473 4278 480 4279
rect 479 4271 480 4278
rect 463 4268 464 4271
rect 479 4268 492 4271
rect 415 4264 445 4265
rect 454 4264 460 4265
rect 463 4264 492 4268
rect 382 4263 492 4264
rect 382 4262 498 4263
rect 57 4254 108 4262
rect 57 4242 82 4254
rect 89 4242 108 4254
rect 139 4254 189 4262
rect 139 4246 155 4254
rect 162 4252 189 4254
rect 198 4252 419 4262
rect 162 4242 419 4252
rect 448 4254 498 4262
rect 448 4245 464 4254
rect 57 4234 108 4242
rect 155 4234 419 4242
rect 445 4242 464 4245
rect 471 4242 498 4254
rect 445 4234 498 4242
rect 73 4226 74 4234
rect 89 4226 102 4234
rect 73 4218 89 4226
rect 70 4211 89 4214
rect 70 4202 92 4211
rect 43 4192 92 4202
rect 43 4186 73 4192
rect 92 4187 97 4192
rect 15 4170 89 4186
rect 107 4178 137 4234
rect 172 4224 380 4234
rect 415 4230 460 4234
rect 463 4233 464 4234
rect 479 4233 492 4234
rect 198 4194 387 4224
rect 213 4191 387 4194
rect 206 4188 387 4191
rect 15 4168 28 4170
rect 43 4168 77 4170
rect 15 4152 89 4168
rect 116 4164 129 4178
rect 144 4164 160 4180
rect 206 4175 217 4188
rect -1 4130 0 4146
rect 15 4130 28 4152
rect 43 4130 73 4152
rect 116 4148 178 4164
rect 206 4157 217 4173
rect 222 4168 232 4188
rect 242 4168 256 4188
rect 259 4175 268 4188
rect 284 4175 293 4188
rect 222 4157 256 4168
rect 259 4157 268 4173
rect 284 4157 293 4173
rect 300 4168 310 4188
rect 320 4168 334 4188
rect 335 4175 346 4188
rect 300 4157 334 4168
rect 335 4157 346 4173
rect 392 4164 408 4180
rect 415 4178 445 4230
rect 479 4226 480 4233
rect 464 4218 480 4226
rect 451 4186 464 4205
rect 479 4186 509 4202
rect 451 4170 525 4186
rect 451 4168 464 4170
rect 479 4168 513 4170
rect 116 4146 129 4148
rect 144 4146 178 4148
rect 116 4130 178 4146
rect 222 4141 238 4144
rect 300 4141 330 4152
rect 378 4148 424 4164
rect 451 4152 525 4168
rect 378 4146 412 4148
rect 377 4130 424 4146
rect 451 4130 464 4152
rect 479 4130 509 4152
rect 536 4130 537 4146
rect 552 4130 565 4290
rect 595 4186 608 4290
rect 653 4268 654 4278
rect 669 4268 682 4278
rect 653 4264 682 4268
rect 687 4264 717 4290
rect 735 4276 751 4278
rect 823 4276 876 4290
rect 824 4274 888 4276
rect 931 4274 946 4290
rect 995 4287 1025 4290
rect 995 4284 1031 4287
rect 961 4276 977 4278
rect 735 4264 750 4268
rect 653 4262 750 4264
rect 778 4262 946 4274
rect 962 4264 977 4268
rect 995 4265 1034 4284
rect 1053 4278 1060 4279
rect 1059 4271 1060 4278
rect 1043 4268 1044 4271
rect 1059 4268 1072 4271
rect 995 4264 1025 4265
rect 1034 4264 1040 4265
rect 1043 4264 1072 4268
rect 962 4263 1072 4264
rect 962 4262 1078 4263
rect 637 4254 688 4262
rect 637 4242 662 4254
rect 669 4242 688 4254
rect 719 4254 769 4262
rect 719 4246 735 4254
rect 742 4252 769 4254
rect 778 4252 999 4262
rect 742 4242 999 4252
rect 1028 4254 1078 4262
rect 1028 4245 1044 4254
rect 637 4234 688 4242
rect 735 4234 999 4242
rect 1025 4242 1044 4245
rect 1051 4242 1078 4254
rect 1025 4234 1078 4242
rect 653 4226 654 4234
rect 669 4226 682 4234
rect 653 4218 669 4226
rect 650 4211 669 4214
rect 650 4202 672 4211
rect 623 4192 672 4202
rect 623 4186 653 4192
rect 672 4187 677 4192
rect 595 4170 669 4186
rect 687 4178 717 4234
rect 752 4224 960 4234
rect 995 4230 1040 4234
rect 1043 4233 1044 4234
rect 1059 4233 1072 4234
rect 778 4194 967 4224
rect 793 4191 967 4194
rect 786 4188 967 4191
rect 595 4168 608 4170
rect 623 4168 657 4170
rect 595 4152 669 4168
rect 696 4164 709 4178
rect 724 4164 740 4180
rect 786 4175 797 4188
rect 579 4130 580 4146
rect 595 4130 608 4152
rect 623 4130 653 4152
rect 696 4148 758 4164
rect 786 4157 797 4173
rect 802 4168 812 4188
rect 822 4168 836 4188
rect 839 4175 848 4188
rect 864 4175 873 4188
rect 802 4157 836 4168
rect 839 4157 848 4173
rect 864 4157 873 4173
rect 880 4168 890 4188
rect 900 4168 914 4188
rect 915 4175 926 4188
rect 880 4157 914 4168
rect 915 4157 926 4173
rect 972 4164 988 4180
rect 995 4178 1025 4230
rect 1059 4226 1060 4233
rect 1044 4218 1060 4226
rect 1031 4186 1044 4205
rect 1059 4186 1089 4202
rect 1031 4170 1105 4186
rect 1031 4168 1044 4170
rect 1059 4168 1093 4170
rect 696 4146 709 4148
rect 724 4146 758 4148
rect 696 4130 758 4146
rect 802 4141 818 4144
rect 880 4141 910 4152
rect 958 4148 1004 4164
rect 1031 4152 1105 4168
rect 958 4146 992 4148
rect 957 4130 1004 4146
rect 1031 4130 1044 4152
rect 1059 4130 1089 4152
rect 1116 4130 1117 4146
rect 1132 4130 1145 4290
rect 1175 4186 1188 4290
rect 1233 4268 1234 4278
rect 1249 4268 1262 4278
rect 1233 4264 1262 4268
rect 1267 4264 1297 4290
rect 1315 4276 1331 4278
rect 1403 4276 1456 4290
rect 1404 4274 1468 4276
rect 1511 4274 1526 4290
rect 1575 4287 1605 4290
rect 1575 4284 1611 4287
rect 1541 4276 1557 4278
rect 1315 4264 1330 4268
rect 1233 4262 1330 4264
rect 1358 4262 1526 4274
rect 1542 4264 1557 4268
rect 1575 4265 1614 4284
rect 1633 4278 1640 4279
rect 1639 4271 1640 4278
rect 1623 4268 1624 4271
rect 1639 4268 1652 4271
rect 1575 4264 1605 4265
rect 1614 4264 1620 4265
rect 1623 4264 1652 4268
rect 1542 4263 1652 4264
rect 1542 4262 1658 4263
rect 1217 4254 1268 4262
rect 1217 4242 1242 4254
rect 1249 4242 1268 4254
rect 1299 4254 1349 4262
rect 1299 4246 1315 4254
rect 1322 4252 1349 4254
rect 1358 4252 1579 4262
rect 1322 4242 1579 4252
rect 1608 4254 1658 4262
rect 1608 4245 1624 4254
rect 1217 4234 1268 4242
rect 1315 4234 1579 4242
rect 1605 4242 1624 4245
rect 1631 4242 1658 4254
rect 1605 4234 1658 4242
rect 1233 4226 1234 4234
rect 1249 4226 1262 4234
rect 1233 4218 1249 4226
rect 1230 4211 1249 4214
rect 1230 4202 1252 4211
rect 1203 4192 1252 4202
rect 1203 4186 1233 4192
rect 1252 4187 1257 4192
rect 1175 4170 1249 4186
rect 1267 4178 1297 4234
rect 1332 4224 1540 4234
rect 1575 4230 1620 4234
rect 1623 4233 1624 4234
rect 1639 4233 1652 4234
rect 1358 4194 1547 4224
rect 1373 4191 1547 4194
rect 1366 4188 1547 4191
rect 1175 4168 1188 4170
rect 1203 4168 1237 4170
rect 1175 4152 1249 4168
rect 1276 4164 1289 4178
rect 1304 4164 1320 4180
rect 1366 4175 1377 4188
rect 1159 4130 1160 4146
rect 1175 4130 1188 4152
rect 1203 4130 1233 4152
rect 1276 4148 1338 4164
rect 1366 4157 1377 4173
rect 1382 4168 1392 4188
rect 1402 4168 1416 4188
rect 1419 4175 1428 4188
rect 1444 4175 1453 4188
rect 1382 4157 1416 4168
rect 1419 4157 1428 4173
rect 1444 4157 1453 4173
rect 1460 4168 1470 4188
rect 1480 4168 1494 4188
rect 1495 4175 1506 4188
rect 1460 4157 1494 4168
rect 1495 4157 1506 4173
rect 1552 4164 1568 4180
rect 1575 4178 1605 4230
rect 1639 4226 1640 4233
rect 1624 4218 1640 4226
rect 1611 4186 1624 4205
rect 1639 4186 1669 4202
rect 1611 4170 1685 4186
rect 1611 4168 1624 4170
rect 1639 4168 1673 4170
rect 1276 4146 1289 4148
rect 1304 4146 1338 4148
rect 1276 4130 1338 4146
rect 1382 4141 1398 4144
rect 1460 4141 1490 4152
rect 1538 4148 1584 4164
rect 1611 4152 1685 4168
rect 1538 4146 1572 4148
rect 1537 4130 1584 4146
rect 1611 4130 1624 4152
rect 1639 4130 1669 4152
rect 1696 4130 1697 4146
rect 1712 4130 1725 4290
rect 1755 4186 1768 4290
rect 1813 4268 1814 4278
rect 1829 4268 1842 4278
rect 1813 4264 1842 4268
rect 1847 4264 1877 4290
rect 1895 4276 1911 4278
rect 1983 4276 2036 4290
rect 1984 4274 2048 4276
rect 2091 4274 2106 4290
rect 2155 4287 2185 4290
rect 2155 4284 2191 4287
rect 2121 4276 2137 4278
rect 1895 4264 1910 4268
rect 1813 4262 1910 4264
rect 1938 4262 2106 4274
rect 2122 4264 2137 4268
rect 2155 4265 2194 4284
rect 2213 4278 2220 4279
rect 2219 4271 2220 4278
rect 2203 4268 2204 4271
rect 2219 4268 2232 4271
rect 2155 4264 2185 4265
rect 2194 4264 2200 4265
rect 2203 4264 2232 4268
rect 2122 4263 2232 4264
rect 2122 4262 2238 4263
rect 1797 4254 1848 4262
rect 1797 4242 1822 4254
rect 1829 4242 1848 4254
rect 1879 4254 1929 4262
rect 1879 4246 1895 4254
rect 1902 4252 1929 4254
rect 1938 4252 2159 4262
rect 1902 4242 2159 4252
rect 2188 4254 2238 4262
rect 2188 4245 2204 4254
rect 1797 4234 1848 4242
rect 1895 4234 2159 4242
rect 2185 4242 2204 4245
rect 2211 4242 2238 4254
rect 2185 4234 2238 4242
rect 1813 4226 1814 4234
rect 1829 4226 1842 4234
rect 1813 4218 1829 4226
rect 1810 4211 1829 4214
rect 1810 4202 1832 4211
rect 1783 4192 1832 4202
rect 1783 4186 1813 4192
rect 1832 4187 1837 4192
rect 1755 4170 1829 4186
rect 1847 4178 1877 4234
rect 1912 4224 2120 4234
rect 2155 4230 2200 4234
rect 2203 4233 2204 4234
rect 2219 4233 2232 4234
rect 1938 4194 2127 4224
rect 1953 4191 2127 4194
rect 1946 4188 2127 4191
rect 1755 4168 1768 4170
rect 1783 4168 1817 4170
rect 1755 4152 1829 4168
rect 1856 4164 1869 4178
rect 1884 4164 1900 4180
rect 1946 4175 1957 4188
rect 1739 4130 1740 4146
rect 1755 4130 1768 4152
rect 1783 4130 1813 4152
rect 1856 4148 1918 4164
rect 1946 4157 1957 4173
rect 1962 4168 1972 4188
rect 1982 4168 1996 4188
rect 1999 4175 2008 4188
rect 2024 4175 2033 4188
rect 1962 4157 1996 4168
rect 1999 4157 2008 4173
rect 2024 4157 2033 4173
rect 2040 4168 2050 4188
rect 2060 4168 2074 4188
rect 2075 4175 2086 4188
rect 2040 4157 2074 4168
rect 2075 4157 2086 4173
rect 2132 4164 2148 4180
rect 2155 4178 2185 4230
rect 2219 4226 2220 4233
rect 2204 4218 2220 4226
rect 2191 4186 2204 4205
rect 2219 4186 2249 4202
rect 2191 4170 2265 4186
rect 2191 4168 2204 4170
rect 2219 4168 2253 4170
rect 1856 4146 1869 4148
rect 1884 4146 1918 4148
rect 1856 4130 1918 4146
rect 1962 4141 1976 4144
rect 2040 4141 2070 4152
rect 2118 4148 2164 4164
rect 2191 4152 2265 4168
rect 2118 4146 2152 4148
rect 2117 4130 2164 4146
rect 2191 4130 2204 4152
rect 2219 4130 2249 4152
rect 2276 4130 2277 4146
rect 2292 4130 2305 4290
rect 2335 4186 2348 4290
rect 2393 4268 2394 4278
rect 2409 4268 2422 4278
rect 2393 4264 2422 4268
rect 2427 4264 2457 4290
rect 2475 4276 2491 4278
rect 2563 4276 2616 4290
rect 2564 4274 2628 4276
rect 2671 4274 2686 4290
rect 2735 4287 2765 4290
rect 2735 4284 2771 4287
rect 2701 4276 2717 4278
rect 2475 4264 2490 4268
rect 2393 4262 2490 4264
rect 2518 4262 2686 4274
rect 2702 4264 2717 4268
rect 2735 4265 2774 4284
rect 2793 4278 2800 4279
rect 2799 4271 2800 4278
rect 2783 4268 2784 4271
rect 2799 4268 2812 4271
rect 2735 4264 2765 4265
rect 2774 4264 2780 4265
rect 2783 4264 2812 4268
rect 2702 4263 2812 4264
rect 2702 4262 2818 4263
rect 2377 4254 2428 4262
rect 2377 4242 2402 4254
rect 2409 4242 2428 4254
rect 2459 4254 2509 4262
rect 2459 4246 2475 4254
rect 2482 4252 2509 4254
rect 2518 4252 2739 4262
rect 2482 4242 2739 4252
rect 2768 4254 2818 4262
rect 2768 4245 2784 4254
rect 2377 4234 2428 4242
rect 2475 4234 2739 4242
rect 2765 4242 2784 4245
rect 2791 4242 2818 4254
rect 2765 4234 2818 4242
rect 2393 4226 2394 4234
rect 2409 4226 2422 4234
rect 2393 4218 2409 4226
rect 2390 4211 2409 4214
rect 2390 4202 2412 4211
rect 2363 4192 2412 4202
rect 2363 4186 2393 4192
rect 2412 4187 2417 4192
rect 2335 4170 2409 4186
rect 2427 4178 2457 4234
rect 2492 4224 2700 4234
rect 2735 4230 2780 4234
rect 2783 4233 2784 4234
rect 2799 4233 2812 4234
rect 2518 4194 2707 4224
rect 2533 4191 2707 4194
rect 2526 4188 2707 4191
rect 2335 4168 2348 4170
rect 2363 4168 2397 4170
rect 2335 4152 2409 4168
rect 2436 4164 2449 4178
rect 2464 4164 2480 4180
rect 2526 4175 2537 4188
rect 2319 4130 2320 4146
rect 2335 4130 2348 4152
rect 2363 4130 2393 4152
rect 2436 4148 2498 4164
rect 2526 4157 2537 4173
rect 2542 4168 2552 4188
rect 2562 4168 2576 4188
rect 2579 4175 2588 4188
rect 2604 4175 2613 4188
rect 2542 4157 2576 4168
rect 2579 4157 2588 4173
rect 2604 4157 2613 4173
rect 2620 4168 2630 4188
rect 2640 4168 2654 4188
rect 2655 4175 2666 4188
rect 2620 4157 2654 4168
rect 2655 4157 2666 4173
rect 2712 4164 2728 4180
rect 2735 4178 2765 4230
rect 2799 4226 2800 4233
rect 2784 4218 2800 4226
rect 2771 4186 2784 4205
rect 2799 4186 2829 4202
rect 2771 4170 2845 4186
rect 2771 4168 2784 4170
rect 2799 4168 2833 4170
rect 2436 4146 2449 4148
rect 2464 4146 2498 4148
rect 2436 4130 2498 4146
rect 2542 4141 2558 4144
rect 2620 4141 2650 4152
rect 2698 4148 2744 4164
rect 2771 4152 2845 4168
rect 2698 4146 2732 4148
rect 2697 4130 2744 4146
rect 2771 4130 2784 4152
rect 2799 4130 2829 4152
rect 2856 4130 2857 4146
rect 2872 4130 2885 4290
rect 2915 4186 2928 4290
rect 2973 4268 2974 4278
rect 2989 4268 3002 4278
rect 2973 4264 3002 4268
rect 3007 4264 3037 4290
rect 3055 4276 3071 4278
rect 3143 4276 3196 4290
rect 3144 4274 3208 4276
rect 3251 4274 3266 4290
rect 3315 4287 3345 4290
rect 3315 4284 3351 4287
rect 3281 4276 3297 4278
rect 3055 4264 3070 4268
rect 2973 4262 3070 4264
rect 3098 4262 3266 4274
rect 3282 4264 3297 4268
rect 3315 4265 3354 4284
rect 3373 4278 3380 4279
rect 3379 4271 3380 4278
rect 3363 4268 3364 4271
rect 3379 4268 3392 4271
rect 3315 4264 3345 4265
rect 3354 4264 3360 4265
rect 3363 4264 3392 4268
rect 3282 4263 3392 4264
rect 3282 4262 3398 4263
rect 2957 4254 3008 4262
rect 2957 4242 2982 4254
rect 2989 4242 3008 4254
rect 3039 4254 3089 4262
rect 3039 4246 3055 4254
rect 3062 4252 3089 4254
rect 3098 4252 3319 4262
rect 3062 4242 3319 4252
rect 3348 4254 3398 4262
rect 3348 4245 3364 4254
rect 2957 4234 3008 4242
rect 3055 4234 3319 4242
rect 3345 4242 3364 4245
rect 3371 4242 3398 4254
rect 3345 4234 3398 4242
rect 2973 4226 2974 4234
rect 2989 4226 3002 4234
rect 2973 4218 2989 4226
rect 2970 4211 2989 4214
rect 2970 4202 2992 4211
rect 2943 4192 2992 4202
rect 2943 4186 2973 4192
rect 2992 4187 2997 4192
rect 2915 4170 2989 4186
rect 3007 4178 3037 4234
rect 3072 4224 3280 4234
rect 3315 4230 3360 4234
rect 3363 4233 3364 4234
rect 3379 4233 3392 4234
rect 3098 4194 3287 4224
rect 3113 4191 3287 4194
rect 3106 4188 3287 4191
rect 2915 4168 2928 4170
rect 2943 4168 2977 4170
rect 2915 4152 2989 4168
rect 3016 4164 3029 4178
rect 3044 4164 3060 4180
rect 3106 4175 3117 4188
rect 2899 4130 2900 4146
rect 2915 4130 2928 4152
rect 2943 4130 2973 4152
rect 3016 4148 3078 4164
rect 3106 4157 3117 4173
rect 3122 4168 3132 4188
rect 3142 4168 3156 4188
rect 3159 4175 3168 4188
rect 3184 4175 3193 4188
rect 3122 4157 3156 4168
rect 3159 4157 3168 4173
rect 3184 4157 3193 4173
rect 3200 4168 3210 4188
rect 3220 4168 3234 4188
rect 3235 4175 3246 4188
rect 3200 4157 3234 4168
rect 3235 4157 3246 4173
rect 3292 4164 3308 4180
rect 3315 4178 3345 4230
rect 3379 4226 3380 4233
rect 3364 4218 3380 4226
rect 3351 4186 3364 4205
rect 3379 4186 3409 4202
rect 3351 4170 3425 4186
rect 3351 4168 3364 4170
rect 3379 4168 3413 4170
rect 3016 4146 3029 4148
rect 3044 4146 3078 4148
rect 3016 4130 3078 4146
rect 3122 4141 3138 4144
rect 3200 4141 3230 4152
rect 3278 4148 3324 4164
rect 3351 4152 3425 4168
rect 3278 4146 3312 4148
rect 3277 4130 3324 4146
rect 3351 4130 3364 4152
rect 3379 4130 3409 4152
rect 3436 4130 3437 4146
rect 3452 4130 3465 4290
rect 3495 4186 3508 4290
rect 3553 4268 3554 4278
rect 3569 4268 3582 4278
rect 3553 4264 3582 4268
rect 3587 4264 3617 4290
rect 3635 4276 3651 4278
rect 3723 4276 3776 4290
rect 3724 4274 3788 4276
rect 3831 4274 3846 4290
rect 3895 4287 3925 4290
rect 3895 4284 3931 4287
rect 3861 4276 3877 4278
rect 3635 4264 3650 4268
rect 3553 4262 3650 4264
rect 3678 4262 3846 4274
rect 3862 4264 3877 4268
rect 3895 4265 3934 4284
rect 3953 4278 3960 4279
rect 3959 4271 3960 4278
rect 3943 4268 3944 4271
rect 3959 4268 3972 4271
rect 3895 4264 3925 4265
rect 3934 4264 3940 4265
rect 3943 4264 3972 4268
rect 3862 4263 3972 4264
rect 3862 4262 3978 4263
rect 3537 4254 3588 4262
rect 3537 4242 3562 4254
rect 3569 4242 3588 4254
rect 3619 4254 3669 4262
rect 3619 4246 3635 4254
rect 3642 4252 3669 4254
rect 3678 4252 3899 4262
rect 3642 4242 3899 4252
rect 3928 4254 3978 4262
rect 3928 4245 3944 4254
rect 3537 4234 3588 4242
rect 3635 4234 3899 4242
rect 3925 4242 3944 4245
rect 3951 4242 3978 4254
rect 3925 4234 3978 4242
rect 3553 4226 3554 4234
rect 3569 4226 3582 4234
rect 3553 4218 3569 4226
rect 3550 4211 3569 4214
rect 3550 4202 3572 4211
rect 3523 4192 3572 4202
rect 3523 4186 3553 4192
rect 3572 4187 3577 4192
rect 3495 4170 3569 4186
rect 3587 4178 3617 4234
rect 3652 4224 3860 4234
rect 3895 4230 3940 4234
rect 3943 4233 3944 4234
rect 3959 4233 3972 4234
rect 3678 4194 3867 4224
rect 3693 4191 3867 4194
rect 3686 4188 3867 4191
rect 3495 4168 3508 4170
rect 3523 4168 3557 4170
rect 3495 4152 3569 4168
rect 3596 4164 3609 4178
rect 3624 4164 3640 4180
rect 3686 4175 3697 4188
rect 3479 4130 3480 4146
rect 3495 4130 3508 4152
rect 3523 4130 3553 4152
rect 3596 4148 3658 4164
rect 3686 4157 3697 4173
rect 3702 4168 3712 4188
rect 3722 4168 3736 4188
rect 3739 4175 3748 4188
rect 3764 4175 3773 4188
rect 3702 4157 3736 4168
rect 3739 4157 3748 4173
rect 3764 4157 3773 4173
rect 3780 4168 3790 4188
rect 3800 4168 3814 4188
rect 3815 4175 3826 4188
rect 3780 4157 3814 4168
rect 3815 4157 3826 4173
rect 3872 4164 3888 4180
rect 3895 4178 3925 4230
rect 3959 4226 3960 4233
rect 3944 4218 3960 4226
rect 3931 4186 3944 4205
rect 3959 4186 3989 4202
rect 3931 4170 4005 4186
rect 3931 4168 3944 4170
rect 3959 4168 3993 4170
rect 3596 4146 3609 4148
rect 3624 4146 3658 4148
rect 3596 4130 3658 4146
rect 3702 4141 3718 4144
rect 3780 4141 3810 4152
rect 3858 4148 3904 4164
rect 3931 4152 4005 4168
rect 3858 4146 3892 4148
rect 3857 4130 3904 4146
rect 3931 4130 3944 4152
rect 3959 4130 3989 4152
rect 4016 4130 4017 4146
rect 4032 4130 4045 4290
rect 4075 4186 4088 4290
rect 4133 4268 4134 4278
rect 4149 4268 4162 4278
rect 4133 4264 4162 4268
rect 4167 4264 4197 4290
rect 4215 4276 4231 4278
rect 4303 4276 4356 4290
rect 4304 4274 4368 4276
rect 4411 4274 4426 4290
rect 4475 4287 4505 4290
rect 4475 4284 4511 4287
rect 4441 4276 4457 4278
rect 4215 4264 4230 4268
rect 4133 4262 4230 4264
rect 4258 4262 4426 4274
rect 4442 4264 4457 4268
rect 4475 4265 4514 4284
rect 4533 4278 4540 4279
rect 4539 4271 4540 4278
rect 4523 4268 4524 4271
rect 4539 4268 4552 4271
rect 4475 4264 4505 4265
rect 4514 4264 4520 4265
rect 4523 4264 4552 4268
rect 4442 4263 4552 4264
rect 4442 4262 4558 4263
rect 4117 4254 4168 4262
rect 4117 4242 4142 4254
rect 4149 4242 4168 4254
rect 4199 4254 4249 4262
rect 4199 4246 4215 4254
rect 4222 4252 4249 4254
rect 4258 4252 4479 4262
rect 4222 4242 4479 4252
rect 4508 4254 4558 4262
rect 4508 4245 4524 4254
rect 4117 4234 4168 4242
rect 4215 4234 4479 4242
rect 4505 4242 4524 4245
rect 4531 4242 4558 4254
rect 4505 4234 4558 4242
rect 4133 4226 4134 4234
rect 4149 4226 4162 4234
rect 4133 4218 4149 4226
rect 4130 4211 4149 4214
rect 4130 4202 4152 4211
rect 4103 4192 4152 4202
rect 4103 4186 4133 4192
rect 4152 4187 4157 4192
rect 4075 4170 4149 4186
rect 4167 4178 4197 4234
rect 4232 4224 4440 4234
rect 4475 4230 4520 4234
rect 4523 4233 4524 4234
rect 4539 4233 4552 4234
rect 4258 4194 4447 4224
rect 4273 4191 4447 4194
rect 4266 4188 4447 4191
rect 4075 4168 4088 4170
rect 4103 4168 4137 4170
rect 4075 4152 4149 4168
rect 4176 4164 4189 4178
rect 4204 4164 4220 4180
rect 4266 4175 4277 4188
rect 4059 4130 4060 4146
rect 4075 4130 4088 4152
rect 4103 4130 4133 4152
rect 4176 4148 4238 4164
rect 4266 4157 4277 4173
rect 4282 4168 4292 4188
rect 4302 4168 4316 4188
rect 4319 4175 4328 4188
rect 4344 4175 4353 4188
rect 4282 4157 4316 4168
rect 4319 4157 4328 4173
rect 4344 4157 4353 4173
rect 4360 4168 4370 4188
rect 4380 4168 4394 4188
rect 4395 4175 4406 4188
rect 4360 4157 4394 4168
rect 4395 4157 4406 4173
rect 4452 4164 4468 4180
rect 4475 4178 4505 4230
rect 4539 4226 4540 4233
rect 4524 4218 4540 4226
rect 4511 4186 4524 4205
rect 4539 4186 4569 4202
rect 4511 4170 4585 4186
rect 4511 4168 4524 4170
rect 4539 4168 4573 4170
rect 4176 4146 4189 4148
rect 4204 4146 4238 4148
rect 4176 4130 4238 4146
rect 4282 4141 4298 4144
rect 4360 4141 4390 4152
rect 4438 4148 4484 4164
rect 4511 4152 4585 4168
rect 4438 4146 4472 4148
rect 4437 4130 4484 4146
rect 4511 4130 4524 4152
rect 4539 4130 4569 4152
rect 4596 4130 4597 4146
rect 4612 4130 4625 4290
rect 4655 4186 4668 4290
rect 4713 4268 4714 4278
rect 4729 4268 4742 4278
rect 4713 4264 4742 4268
rect 4747 4264 4777 4290
rect 4795 4276 4811 4278
rect 4883 4276 4936 4290
rect 4884 4274 4948 4276
rect 4991 4274 5006 4290
rect 5055 4287 5085 4290
rect 5055 4284 5091 4287
rect 5021 4276 5037 4278
rect 4795 4264 4810 4268
rect 4713 4262 4810 4264
rect 4838 4262 5006 4274
rect 5022 4264 5037 4268
rect 5055 4265 5094 4284
rect 5113 4278 5120 4279
rect 5119 4271 5120 4278
rect 5103 4268 5104 4271
rect 5119 4268 5132 4271
rect 5055 4264 5085 4265
rect 5094 4264 5100 4265
rect 5103 4264 5132 4268
rect 5022 4263 5132 4264
rect 5022 4262 5138 4263
rect 4697 4254 4748 4262
rect 4697 4242 4722 4254
rect 4729 4242 4748 4254
rect 4779 4254 4829 4262
rect 4779 4246 4795 4254
rect 4802 4252 4829 4254
rect 4838 4252 5059 4262
rect 4802 4242 5059 4252
rect 5088 4254 5138 4262
rect 5088 4245 5104 4254
rect 4697 4234 4748 4242
rect 4795 4234 5059 4242
rect 5085 4242 5104 4245
rect 5111 4242 5138 4254
rect 5085 4234 5138 4242
rect 4713 4226 4714 4234
rect 4729 4226 4742 4234
rect 4713 4218 4729 4226
rect 4710 4211 4729 4214
rect 4710 4202 4732 4211
rect 4683 4192 4732 4202
rect 4683 4186 4713 4192
rect 4732 4187 4737 4192
rect 4655 4170 4729 4186
rect 4747 4178 4777 4234
rect 4812 4224 5020 4234
rect 5055 4230 5100 4234
rect 5103 4233 5104 4234
rect 5119 4233 5132 4234
rect 4838 4194 5027 4224
rect 4853 4191 5027 4194
rect 4846 4188 5027 4191
rect 4655 4168 4668 4170
rect 4683 4168 4717 4170
rect 4655 4152 4729 4168
rect 4756 4164 4769 4178
rect 4784 4164 4800 4180
rect 4846 4175 4857 4188
rect 4639 4130 4640 4146
rect 4655 4130 4668 4152
rect 4683 4130 4713 4152
rect 4756 4148 4818 4164
rect 4846 4157 4857 4173
rect 4862 4168 4872 4188
rect 4882 4168 4896 4188
rect 4899 4175 4908 4188
rect 4924 4175 4933 4188
rect 4862 4157 4896 4168
rect 4899 4157 4908 4173
rect 4924 4157 4933 4173
rect 4940 4168 4950 4188
rect 4960 4168 4974 4188
rect 4975 4175 4986 4188
rect 4940 4157 4974 4168
rect 4975 4157 4986 4173
rect 5032 4164 5048 4180
rect 5055 4178 5085 4230
rect 5119 4226 5120 4233
rect 5104 4218 5120 4226
rect 5091 4186 5104 4205
rect 5119 4186 5149 4202
rect 5091 4170 5165 4186
rect 5091 4168 5104 4170
rect 5119 4168 5153 4170
rect 4756 4146 4769 4148
rect 4784 4146 4818 4148
rect 4756 4130 4818 4146
rect 4862 4141 4878 4144
rect 4940 4141 4970 4152
rect 5018 4148 5064 4164
rect 5091 4152 5165 4168
rect 5018 4146 5052 4148
rect 5017 4130 5064 4146
rect 5091 4130 5104 4152
rect 5119 4130 5149 4152
rect 5176 4130 5177 4146
rect 5192 4130 5205 4290
rect 5235 4186 5248 4290
rect 5293 4268 5294 4278
rect 5309 4268 5322 4278
rect 5293 4264 5322 4268
rect 5327 4264 5357 4290
rect 5375 4276 5391 4278
rect 5463 4276 5516 4290
rect 5464 4274 5528 4276
rect 5571 4274 5586 4290
rect 5635 4287 5665 4290
rect 5635 4284 5671 4287
rect 5601 4276 5617 4278
rect 5375 4264 5390 4268
rect 5293 4262 5390 4264
rect 5418 4262 5586 4274
rect 5602 4264 5617 4268
rect 5635 4265 5674 4284
rect 5693 4278 5700 4279
rect 5699 4271 5700 4278
rect 5683 4268 5684 4271
rect 5699 4268 5712 4271
rect 5635 4264 5665 4265
rect 5674 4264 5680 4265
rect 5683 4264 5712 4268
rect 5602 4263 5712 4264
rect 5602 4262 5718 4263
rect 5277 4254 5328 4262
rect 5277 4242 5302 4254
rect 5309 4242 5328 4254
rect 5359 4254 5409 4262
rect 5359 4246 5375 4254
rect 5382 4252 5409 4254
rect 5418 4252 5639 4262
rect 5382 4242 5639 4252
rect 5668 4254 5718 4262
rect 5668 4245 5684 4254
rect 5277 4234 5328 4242
rect 5375 4234 5639 4242
rect 5665 4242 5684 4245
rect 5691 4242 5718 4254
rect 5665 4234 5718 4242
rect 5293 4226 5294 4234
rect 5309 4226 5322 4234
rect 5293 4218 5309 4226
rect 5290 4211 5309 4214
rect 5290 4202 5312 4211
rect 5263 4192 5312 4202
rect 5263 4186 5293 4192
rect 5312 4187 5317 4192
rect 5235 4170 5309 4186
rect 5327 4178 5357 4234
rect 5392 4224 5600 4234
rect 5635 4230 5680 4234
rect 5683 4233 5684 4234
rect 5699 4233 5712 4234
rect 5418 4194 5607 4224
rect 5433 4191 5607 4194
rect 5426 4188 5607 4191
rect 5235 4168 5248 4170
rect 5263 4168 5297 4170
rect 5235 4152 5309 4168
rect 5336 4164 5349 4178
rect 5364 4164 5380 4180
rect 5426 4175 5437 4188
rect 5219 4130 5220 4146
rect 5235 4130 5248 4152
rect 5263 4130 5293 4152
rect 5336 4148 5398 4164
rect 5426 4157 5437 4173
rect 5442 4168 5452 4188
rect 5462 4168 5476 4188
rect 5479 4175 5488 4188
rect 5504 4175 5513 4188
rect 5442 4157 5476 4168
rect 5479 4157 5488 4173
rect 5504 4157 5513 4173
rect 5520 4168 5530 4188
rect 5540 4168 5554 4188
rect 5555 4175 5566 4188
rect 5520 4157 5554 4168
rect 5555 4157 5566 4173
rect 5612 4164 5628 4180
rect 5635 4178 5665 4230
rect 5699 4226 5700 4233
rect 5684 4218 5700 4226
rect 5671 4186 5684 4205
rect 5699 4186 5729 4202
rect 5671 4170 5745 4186
rect 5671 4168 5684 4170
rect 5699 4168 5733 4170
rect 5336 4146 5349 4148
rect 5364 4146 5398 4148
rect 5336 4130 5398 4146
rect 5442 4141 5458 4144
rect 5520 4141 5550 4152
rect 5598 4148 5644 4164
rect 5671 4152 5745 4168
rect 5598 4146 5632 4148
rect 5597 4130 5644 4146
rect 5671 4130 5684 4152
rect 5699 4130 5729 4152
rect 5756 4130 5757 4146
rect 5772 4130 5785 4290
rect 5815 4186 5828 4290
rect 5873 4268 5874 4278
rect 5889 4268 5902 4278
rect 5873 4264 5902 4268
rect 5907 4264 5937 4290
rect 5955 4276 5971 4278
rect 6043 4276 6096 4290
rect 6044 4274 6108 4276
rect 6151 4274 6166 4290
rect 6215 4287 6245 4290
rect 6215 4284 6251 4287
rect 6181 4276 6197 4278
rect 5955 4264 5970 4268
rect 5873 4262 5970 4264
rect 5998 4262 6166 4274
rect 6182 4264 6197 4268
rect 6215 4265 6254 4284
rect 6273 4278 6280 4279
rect 6279 4271 6280 4278
rect 6263 4268 6264 4271
rect 6279 4268 6292 4271
rect 6215 4264 6245 4265
rect 6254 4264 6260 4265
rect 6263 4264 6292 4268
rect 6182 4263 6292 4264
rect 6182 4262 6298 4263
rect 5857 4254 5908 4262
rect 5857 4242 5882 4254
rect 5889 4242 5908 4254
rect 5939 4254 5989 4262
rect 5939 4246 5955 4254
rect 5962 4252 5989 4254
rect 5998 4252 6219 4262
rect 5962 4242 6219 4252
rect 6248 4254 6298 4262
rect 6248 4245 6264 4254
rect 5857 4234 5908 4242
rect 5955 4234 6219 4242
rect 6245 4242 6264 4245
rect 6271 4242 6298 4254
rect 6245 4234 6298 4242
rect 5873 4226 5874 4234
rect 5889 4226 5902 4234
rect 5873 4218 5889 4226
rect 5870 4211 5889 4214
rect 5870 4202 5892 4211
rect 5843 4192 5892 4202
rect 5843 4186 5873 4192
rect 5892 4187 5897 4192
rect 5815 4170 5889 4186
rect 5907 4178 5937 4234
rect 5972 4224 6180 4234
rect 6215 4230 6260 4234
rect 6263 4233 6264 4234
rect 6279 4233 6292 4234
rect 5998 4194 6187 4224
rect 6013 4191 6187 4194
rect 6006 4188 6187 4191
rect 5815 4168 5828 4170
rect 5843 4168 5877 4170
rect 5815 4152 5889 4168
rect 5916 4164 5929 4178
rect 5944 4164 5960 4180
rect 6006 4175 6017 4188
rect 5799 4130 5800 4146
rect 5815 4130 5828 4152
rect 5843 4130 5873 4152
rect 5916 4148 5978 4164
rect 6006 4157 6017 4173
rect 6022 4168 6032 4188
rect 6042 4168 6056 4188
rect 6059 4175 6068 4188
rect 6084 4175 6093 4188
rect 6022 4157 6056 4168
rect 6059 4157 6068 4173
rect 6084 4157 6093 4173
rect 6100 4168 6110 4188
rect 6120 4168 6134 4188
rect 6135 4175 6146 4188
rect 6100 4157 6134 4168
rect 6135 4157 6146 4173
rect 6192 4164 6208 4180
rect 6215 4178 6245 4230
rect 6279 4226 6280 4233
rect 6264 4218 6280 4226
rect 6251 4186 6264 4205
rect 6279 4186 6309 4202
rect 6251 4170 6325 4186
rect 6251 4168 6264 4170
rect 6279 4168 6313 4170
rect 5916 4146 5929 4148
rect 5944 4146 5978 4148
rect 5916 4130 5978 4146
rect 6022 4141 6038 4144
rect 6100 4141 6130 4152
rect 6178 4148 6224 4164
rect 6251 4152 6325 4168
rect 6178 4146 6212 4148
rect 6177 4130 6224 4146
rect 6251 4130 6264 4152
rect 6279 4130 6309 4152
rect 6336 4130 6337 4146
rect 6352 4130 6365 4290
rect 6395 4186 6408 4290
rect 6453 4268 6454 4278
rect 6469 4268 6482 4278
rect 6453 4264 6482 4268
rect 6487 4264 6517 4290
rect 6535 4276 6551 4278
rect 6623 4276 6676 4290
rect 6624 4274 6688 4276
rect 6731 4274 6746 4290
rect 6795 4287 6825 4290
rect 6795 4284 6831 4287
rect 6761 4276 6777 4278
rect 6535 4264 6550 4268
rect 6453 4262 6550 4264
rect 6578 4262 6746 4274
rect 6762 4264 6777 4268
rect 6795 4265 6834 4284
rect 6853 4278 6860 4279
rect 6859 4271 6860 4278
rect 6843 4268 6844 4271
rect 6859 4268 6872 4271
rect 6795 4264 6825 4265
rect 6834 4264 6840 4265
rect 6843 4264 6872 4268
rect 6762 4263 6872 4264
rect 6762 4262 6878 4263
rect 6437 4254 6488 4262
rect 6437 4242 6462 4254
rect 6469 4242 6488 4254
rect 6519 4254 6569 4262
rect 6519 4246 6535 4254
rect 6542 4252 6569 4254
rect 6578 4252 6799 4262
rect 6542 4242 6799 4252
rect 6828 4254 6878 4262
rect 6828 4245 6844 4254
rect 6437 4234 6488 4242
rect 6535 4234 6799 4242
rect 6825 4242 6844 4245
rect 6851 4242 6878 4254
rect 6825 4234 6878 4242
rect 6453 4226 6454 4234
rect 6469 4226 6482 4234
rect 6453 4218 6469 4226
rect 6450 4211 6469 4214
rect 6450 4202 6472 4211
rect 6423 4192 6472 4202
rect 6423 4186 6453 4192
rect 6472 4187 6477 4192
rect 6395 4170 6469 4186
rect 6487 4178 6517 4234
rect 6552 4224 6760 4234
rect 6795 4230 6840 4234
rect 6843 4233 6844 4234
rect 6859 4233 6872 4234
rect 6578 4194 6767 4224
rect 6593 4191 6767 4194
rect 6586 4188 6767 4191
rect 6395 4168 6408 4170
rect 6423 4168 6457 4170
rect 6395 4152 6469 4168
rect 6496 4164 6509 4178
rect 6524 4164 6540 4180
rect 6586 4175 6597 4188
rect 6379 4130 6380 4146
rect 6395 4130 6408 4152
rect 6423 4130 6453 4152
rect 6496 4148 6558 4164
rect 6586 4157 6597 4173
rect 6602 4168 6612 4188
rect 6622 4168 6636 4188
rect 6639 4175 6648 4188
rect 6664 4175 6673 4188
rect 6602 4157 6636 4168
rect 6639 4157 6648 4173
rect 6664 4157 6673 4173
rect 6680 4168 6690 4188
rect 6700 4168 6714 4188
rect 6715 4175 6726 4188
rect 6680 4157 6714 4168
rect 6715 4157 6726 4173
rect 6772 4164 6788 4180
rect 6795 4178 6825 4230
rect 6859 4226 6860 4233
rect 6844 4218 6860 4226
rect 6831 4186 6844 4205
rect 6859 4186 6889 4202
rect 6831 4170 6905 4186
rect 6831 4168 6844 4170
rect 6859 4168 6893 4170
rect 6496 4146 6509 4148
rect 6524 4146 6558 4148
rect 6496 4130 6558 4146
rect 6602 4141 6618 4144
rect 6680 4141 6710 4152
rect 6758 4148 6804 4164
rect 6831 4152 6905 4168
rect 6758 4146 6792 4148
rect 6757 4130 6804 4146
rect 6831 4130 6844 4152
rect 6859 4130 6889 4152
rect 6916 4130 6917 4146
rect 6932 4130 6945 4290
rect 6975 4186 6988 4290
rect 7033 4268 7034 4278
rect 7049 4268 7062 4278
rect 7033 4264 7062 4268
rect 7067 4264 7097 4290
rect 7115 4276 7131 4278
rect 7203 4276 7256 4290
rect 7206 4274 7268 4276
rect 7311 4274 7326 4290
rect 7375 4287 7405 4290
rect 7375 4284 7411 4287
rect 7341 4276 7357 4278
rect 7115 4264 7130 4268
rect 7033 4262 7130 4264
rect 7158 4262 7326 4274
rect 7342 4264 7357 4268
rect 7375 4265 7414 4284
rect 7433 4278 7440 4279
rect 7439 4271 7440 4278
rect 7423 4268 7424 4271
rect 7439 4268 7452 4271
rect 7375 4264 7405 4265
rect 7414 4264 7420 4265
rect 7423 4264 7452 4268
rect 7342 4263 7452 4264
rect 7342 4262 7458 4263
rect 7017 4254 7068 4262
rect 7017 4242 7042 4254
rect 7049 4242 7068 4254
rect 7099 4254 7149 4262
rect 7099 4246 7115 4254
rect 7122 4252 7149 4254
rect 7158 4252 7379 4262
rect 7122 4242 7379 4252
rect 7408 4254 7458 4262
rect 7408 4245 7424 4254
rect 7017 4234 7068 4242
rect 7115 4234 7379 4242
rect 7405 4242 7424 4245
rect 7431 4242 7458 4254
rect 7405 4234 7458 4242
rect 7033 4226 7034 4234
rect 7049 4226 7062 4234
rect 7033 4218 7049 4226
rect 7030 4211 7049 4214
rect 7030 4202 7052 4211
rect 7003 4192 7052 4202
rect 7003 4186 7033 4192
rect 7052 4187 7057 4192
rect 6975 4170 7049 4186
rect 7067 4178 7097 4234
rect 7132 4224 7340 4234
rect 7375 4230 7420 4234
rect 7423 4233 7424 4234
rect 7439 4233 7452 4234
rect 7158 4194 7347 4224
rect 7173 4191 7347 4194
rect 7166 4188 7347 4191
rect 6975 4168 6988 4170
rect 7003 4168 7037 4170
rect 6975 4152 7049 4168
rect 7076 4164 7089 4178
rect 7104 4164 7120 4180
rect 7166 4175 7177 4188
rect 6959 4130 6960 4146
rect 6975 4130 6988 4152
rect 7003 4130 7033 4152
rect 7076 4148 7138 4164
rect 7166 4157 7177 4173
rect 7182 4168 7192 4188
rect 7202 4168 7216 4188
rect 7219 4175 7228 4188
rect 7244 4175 7253 4188
rect 7182 4157 7216 4168
rect 7219 4157 7228 4173
rect 7244 4157 7253 4173
rect 7260 4168 7270 4188
rect 7280 4168 7294 4188
rect 7295 4175 7306 4188
rect 7260 4157 7294 4168
rect 7295 4157 7306 4173
rect 7352 4164 7368 4180
rect 7375 4178 7405 4230
rect 7439 4226 7440 4233
rect 7424 4218 7440 4226
rect 7411 4186 7424 4205
rect 7439 4186 7469 4202
rect 7411 4170 7485 4186
rect 7411 4168 7424 4170
rect 7439 4168 7473 4170
rect 7076 4146 7089 4148
rect 7104 4146 7138 4148
rect 7076 4130 7138 4146
rect 7182 4141 7198 4144
rect 7260 4141 7290 4152
rect 7338 4148 7384 4164
rect 7411 4152 7485 4168
rect 7338 4146 7372 4148
rect 7337 4130 7384 4146
rect 7411 4130 7424 4152
rect 7439 4130 7469 4152
rect 7496 4130 7497 4146
rect 7512 4130 7525 4290
rect 7555 4186 7568 4290
rect 7613 4268 7614 4278
rect 7629 4268 7642 4278
rect 7613 4264 7642 4268
rect 7647 4264 7677 4290
rect 7695 4276 7711 4278
rect 7783 4276 7836 4290
rect 7784 4274 7848 4276
rect 7891 4274 7906 4290
rect 7955 4287 7985 4290
rect 7955 4284 7991 4287
rect 7921 4276 7937 4278
rect 7695 4264 7710 4268
rect 7613 4262 7710 4264
rect 7738 4262 7906 4274
rect 7922 4264 7937 4268
rect 7955 4265 7994 4284
rect 8013 4278 8020 4279
rect 8019 4271 8020 4278
rect 8003 4268 8004 4271
rect 8019 4268 8032 4271
rect 7955 4264 7985 4265
rect 7994 4264 8000 4265
rect 8003 4264 8032 4268
rect 7922 4263 8032 4264
rect 7922 4262 8038 4263
rect 7597 4254 7648 4262
rect 7597 4242 7622 4254
rect 7629 4242 7648 4254
rect 7679 4254 7729 4262
rect 7679 4246 7695 4254
rect 7702 4252 7729 4254
rect 7738 4252 7959 4262
rect 7702 4242 7959 4252
rect 7988 4254 8038 4262
rect 7988 4245 8004 4254
rect 7597 4234 7648 4242
rect 7695 4234 7959 4242
rect 7985 4242 8004 4245
rect 8011 4242 8038 4254
rect 7985 4234 8038 4242
rect 7613 4226 7614 4234
rect 7629 4226 7642 4234
rect 7613 4218 7629 4226
rect 7610 4211 7629 4214
rect 7610 4202 7632 4211
rect 7583 4192 7632 4202
rect 7583 4186 7613 4192
rect 7632 4187 7637 4192
rect 7555 4170 7629 4186
rect 7647 4178 7677 4234
rect 7712 4224 7920 4234
rect 7955 4230 8000 4234
rect 8003 4233 8004 4234
rect 8019 4233 8032 4234
rect 7738 4194 7927 4224
rect 7753 4191 7927 4194
rect 7746 4188 7927 4191
rect 7555 4168 7568 4170
rect 7583 4168 7617 4170
rect 7555 4152 7629 4168
rect 7656 4164 7669 4178
rect 7684 4164 7700 4180
rect 7746 4175 7757 4188
rect 7539 4130 7540 4146
rect 7555 4130 7568 4152
rect 7583 4130 7613 4152
rect 7656 4148 7718 4164
rect 7746 4157 7757 4173
rect 7762 4168 7772 4188
rect 7782 4168 7796 4188
rect 7799 4175 7808 4188
rect 7824 4175 7833 4188
rect 7762 4157 7796 4168
rect 7799 4157 7808 4173
rect 7824 4157 7833 4173
rect 7840 4168 7850 4188
rect 7860 4168 7874 4188
rect 7875 4175 7886 4188
rect 7840 4157 7874 4168
rect 7875 4157 7886 4173
rect 7932 4164 7948 4180
rect 7955 4178 7985 4230
rect 8019 4226 8020 4233
rect 8004 4218 8020 4226
rect 7991 4186 8004 4205
rect 8019 4186 8049 4202
rect 7991 4170 8065 4186
rect 7991 4168 8004 4170
rect 8019 4168 8053 4170
rect 7656 4146 7669 4148
rect 7684 4146 7718 4148
rect 7656 4130 7718 4146
rect 7762 4141 7778 4144
rect 7840 4141 7870 4152
rect 7918 4148 7964 4164
rect 7991 4152 8065 4168
rect 7918 4146 7952 4148
rect 7917 4130 7964 4146
rect 7991 4130 8004 4152
rect 8019 4130 8049 4152
rect 8076 4130 8077 4146
rect 8092 4130 8105 4290
rect 8135 4186 8148 4290
rect 8193 4268 8194 4278
rect 8209 4268 8222 4278
rect 8193 4264 8222 4268
rect 8227 4264 8257 4290
rect 8275 4276 8291 4278
rect 8363 4276 8416 4290
rect 8364 4274 8428 4276
rect 8471 4274 8486 4290
rect 8535 4287 8565 4290
rect 8535 4284 8571 4287
rect 8501 4276 8517 4278
rect 8275 4264 8290 4268
rect 8193 4262 8290 4264
rect 8318 4262 8486 4274
rect 8502 4264 8517 4268
rect 8535 4265 8574 4284
rect 8593 4278 8600 4279
rect 8599 4271 8600 4278
rect 8583 4268 8584 4271
rect 8599 4268 8612 4271
rect 8535 4264 8565 4265
rect 8574 4264 8580 4265
rect 8583 4264 8612 4268
rect 8502 4263 8612 4264
rect 8502 4262 8618 4263
rect 8177 4254 8228 4262
rect 8177 4242 8202 4254
rect 8209 4242 8228 4254
rect 8259 4254 8309 4262
rect 8259 4246 8275 4254
rect 8282 4252 8309 4254
rect 8318 4252 8539 4262
rect 8282 4242 8539 4252
rect 8568 4254 8618 4262
rect 8568 4245 8584 4254
rect 8177 4234 8228 4242
rect 8275 4234 8539 4242
rect 8565 4242 8584 4245
rect 8591 4242 8618 4254
rect 8565 4234 8618 4242
rect 8193 4226 8194 4234
rect 8209 4226 8222 4234
rect 8193 4218 8209 4226
rect 8190 4211 8209 4214
rect 8190 4202 8212 4211
rect 8163 4192 8212 4202
rect 8163 4186 8193 4192
rect 8212 4187 8217 4192
rect 8135 4170 8209 4186
rect 8227 4178 8257 4234
rect 8292 4224 8500 4234
rect 8535 4230 8580 4234
rect 8583 4233 8584 4234
rect 8599 4233 8612 4234
rect 8318 4194 8507 4224
rect 8333 4191 8507 4194
rect 8326 4188 8507 4191
rect 8135 4168 8148 4170
rect 8163 4168 8197 4170
rect 8135 4152 8209 4168
rect 8236 4164 8249 4178
rect 8264 4164 8280 4180
rect 8326 4175 8337 4188
rect 8119 4130 8120 4146
rect 8135 4130 8148 4152
rect 8163 4130 8193 4152
rect 8236 4148 8298 4164
rect 8326 4157 8337 4173
rect 8342 4168 8352 4188
rect 8362 4168 8376 4188
rect 8379 4175 8388 4188
rect 8404 4175 8413 4188
rect 8342 4157 8376 4168
rect 8379 4157 8388 4173
rect 8404 4157 8413 4173
rect 8420 4168 8430 4188
rect 8440 4168 8454 4188
rect 8455 4175 8466 4188
rect 8420 4157 8454 4168
rect 8455 4157 8466 4173
rect 8512 4164 8528 4180
rect 8535 4178 8565 4230
rect 8599 4226 8600 4233
rect 8584 4218 8600 4226
rect 8571 4186 8584 4205
rect 8599 4186 8629 4202
rect 8571 4170 8645 4186
rect 8571 4168 8584 4170
rect 8599 4168 8633 4170
rect 8236 4146 8249 4148
rect 8264 4146 8298 4148
rect 8236 4130 8298 4146
rect 8342 4141 8358 4144
rect 8420 4141 8450 4152
rect 8498 4148 8544 4164
rect 8571 4152 8645 4168
rect 8498 4146 8532 4148
rect 8497 4130 8544 4146
rect 8571 4130 8584 4152
rect 8599 4130 8629 4152
rect 8656 4130 8657 4146
rect 8672 4130 8685 4290
rect 8715 4186 8728 4290
rect 8773 4268 8774 4278
rect 8789 4268 8802 4278
rect 8773 4264 8802 4268
rect 8807 4264 8837 4290
rect 8855 4276 8871 4278
rect 8943 4276 8996 4290
rect 8944 4274 9008 4276
rect 9051 4274 9066 4290
rect 9115 4287 9145 4290
rect 9115 4284 9151 4287
rect 9081 4276 9097 4278
rect 8855 4264 8870 4268
rect 8773 4262 8870 4264
rect 8898 4262 9066 4274
rect 9082 4264 9097 4268
rect 9115 4265 9154 4284
rect 9173 4278 9180 4279
rect 9179 4271 9180 4278
rect 9163 4268 9164 4271
rect 9179 4268 9192 4271
rect 9115 4264 9145 4265
rect 9154 4264 9160 4265
rect 9163 4264 9192 4268
rect 9082 4263 9192 4264
rect 9082 4262 9198 4263
rect 8757 4254 8808 4262
rect 8757 4242 8782 4254
rect 8789 4242 8808 4254
rect 8839 4254 8889 4262
rect 8839 4246 8855 4254
rect 8862 4252 8889 4254
rect 8898 4252 9119 4262
rect 8862 4242 9119 4252
rect 9148 4254 9198 4262
rect 9148 4245 9164 4254
rect 8757 4234 8808 4242
rect 8855 4234 9119 4242
rect 9145 4242 9164 4245
rect 9171 4242 9198 4254
rect 9145 4234 9198 4242
rect 8773 4226 8774 4234
rect 8789 4226 8802 4234
rect 8773 4218 8789 4226
rect 8770 4211 8789 4214
rect 8770 4202 8792 4211
rect 8743 4192 8792 4202
rect 8743 4186 8773 4192
rect 8792 4187 8797 4192
rect 8715 4170 8789 4186
rect 8807 4178 8837 4234
rect 8872 4224 9080 4234
rect 9115 4230 9160 4234
rect 9163 4233 9164 4234
rect 9179 4233 9192 4234
rect 8898 4194 9087 4224
rect 8913 4191 9087 4194
rect 8906 4188 9087 4191
rect 8715 4168 8728 4170
rect 8743 4168 8777 4170
rect 8715 4152 8789 4168
rect 8816 4164 8829 4178
rect 8844 4164 8860 4180
rect 8906 4175 8917 4188
rect 8699 4130 8700 4146
rect 8715 4130 8728 4152
rect 8743 4130 8773 4152
rect 8816 4148 8878 4164
rect 8906 4157 8917 4173
rect 8922 4168 8932 4188
rect 8942 4168 8956 4188
rect 8959 4175 8968 4188
rect 8984 4175 8993 4188
rect 8922 4157 8956 4168
rect 8959 4157 8968 4173
rect 8984 4157 8993 4173
rect 9000 4168 9010 4188
rect 9020 4168 9034 4188
rect 9035 4175 9046 4188
rect 9000 4157 9034 4168
rect 9035 4157 9046 4173
rect 9092 4164 9108 4180
rect 9115 4178 9145 4230
rect 9179 4226 9180 4233
rect 9164 4218 9180 4226
rect 9151 4186 9164 4205
rect 9179 4186 9209 4202
rect 9151 4170 9225 4186
rect 9151 4168 9164 4170
rect 9179 4168 9213 4170
rect 8816 4146 8829 4148
rect 8844 4146 8878 4148
rect 8816 4130 8878 4146
rect 8922 4141 8938 4144
rect 9000 4141 9030 4152
rect 9078 4148 9124 4164
rect 9151 4152 9225 4168
rect 9078 4146 9112 4148
rect 9077 4130 9124 4146
rect 9151 4130 9164 4152
rect 9179 4130 9209 4152
rect 9236 4130 9237 4146
rect 9252 4130 9265 4290
rect -7 4122 34 4130
rect -7 4096 8 4122
rect 15 4096 34 4122
rect 98 4118 160 4130
rect 172 4118 247 4130
rect 305 4118 380 4130
rect 392 4118 423 4130
rect 429 4118 464 4130
rect 98 4116 260 4118
rect -7 4088 34 4096
rect 116 4092 129 4116
rect 144 4114 159 4116
rect -1 4078 0 4088
rect 15 4078 28 4088
rect 43 4078 73 4092
rect 116 4078 159 4092
rect 183 4089 190 4096
rect 193 4092 260 4116
rect 292 4116 464 4118
rect 262 4094 290 4098
rect 292 4094 372 4116
rect 393 4114 408 4116
rect 262 4092 372 4094
rect 193 4088 372 4092
rect 166 4078 196 4088
rect 198 4078 351 4088
rect 359 4078 389 4088
rect 393 4078 423 4092
rect 451 4078 464 4116
rect 536 4122 571 4130
rect 536 4096 537 4122
rect 544 4096 571 4122
rect 479 4078 509 4092
rect 536 4088 571 4096
rect 573 4122 614 4130
rect 573 4096 588 4122
rect 595 4096 614 4122
rect 678 4118 740 4130
rect 752 4118 827 4130
rect 885 4118 960 4130
rect 972 4118 1003 4130
rect 1009 4118 1044 4130
rect 678 4116 840 4118
rect 573 4088 614 4096
rect 696 4092 709 4116
rect 724 4114 739 4116
rect 536 4078 537 4088
rect 552 4078 565 4088
rect 579 4078 580 4088
rect 595 4078 608 4088
rect 623 4078 653 4092
rect 696 4078 739 4092
rect 763 4089 770 4096
rect 773 4092 840 4116
rect 872 4116 1044 4118
rect 842 4094 870 4098
rect 872 4094 952 4116
rect 973 4114 988 4116
rect 842 4092 952 4094
rect 773 4088 952 4092
rect 746 4078 776 4088
rect 778 4078 931 4088
rect 939 4078 969 4088
rect 973 4078 1003 4092
rect 1031 4078 1044 4116
rect 1116 4122 1151 4130
rect 1116 4096 1117 4122
rect 1124 4096 1151 4122
rect 1059 4078 1089 4092
rect 1116 4088 1151 4096
rect 1153 4122 1194 4130
rect 1153 4096 1168 4122
rect 1175 4096 1194 4122
rect 1258 4118 1320 4130
rect 1332 4118 1407 4130
rect 1465 4118 1540 4130
rect 1552 4118 1583 4130
rect 1589 4118 1624 4130
rect 1258 4116 1420 4118
rect 1153 4088 1194 4096
rect 1276 4092 1289 4116
rect 1304 4114 1319 4116
rect 1116 4078 1117 4088
rect 1132 4078 1145 4088
rect 1159 4078 1160 4088
rect 1175 4078 1188 4088
rect 1203 4078 1233 4092
rect 1276 4078 1319 4092
rect 1343 4089 1350 4096
rect 1353 4092 1420 4116
rect 1452 4116 1624 4118
rect 1422 4094 1450 4098
rect 1452 4094 1532 4116
rect 1553 4114 1568 4116
rect 1422 4092 1532 4094
rect 1353 4088 1532 4092
rect 1326 4078 1356 4088
rect 1358 4078 1511 4088
rect 1519 4078 1549 4088
rect 1553 4078 1583 4092
rect 1611 4078 1624 4116
rect 1696 4122 1731 4130
rect 1696 4096 1697 4122
rect 1704 4096 1731 4122
rect 1639 4078 1669 4092
rect 1696 4088 1731 4096
rect 1733 4122 1774 4130
rect 1733 4096 1748 4122
rect 1755 4096 1774 4122
rect 1838 4118 1900 4130
rect 1912 4118 1987 4130
rect 2045 4118 2120 4130
rect 2132 4118 2163 4130
rect 2169 4118 2204 4130
rect 1838 4116 2000 4118
rect 1733 4088 1774 4096
rect 1856 4092 1869 4116
rect 1884 4114 1899 4116
rect 1696 4078 1697 4088
rect 1712 4078 1725 4088
rect 1739 4078 1740 4088
rect 1755 4078 1768 4088
rect 1783 4078 1813 4092
rect 1856 4078 1899 4092
rect 1923 4089 1930 4096
rect 1933 4092 2000 4116
rect 2032 4116 2204 4118
rect 2002 4094 2030 4098
rect 2032 4094 2112 4116
rect 2133 4114 2148 4116
rect 2002 4092 2112 4094
rect 1933 4088 2112 4092
rect 1906 4078 1936 4088
rect 1938 4078 2091 4088
rect 2099 4078 2129 4088
rect 2133 4078 2163 4092
rect 2191 4078 2204 4116
rect 2276 4122 2311 4130
rect 2276 4096 2277 4122
rect 2284 4096 2311 4122
rect 2219 4078 2249 4092
rect 2276 4088 2311 4096
rect 2313 4122 2354 4130
rect 2313 4096 2328 4122
rect 2335 4096 2354 4122
rect 2418 4118 2480 4130
rect 2492 4118 2567 4130
rect 2625 4118 2700 4130
rect 2712 4118 2743 4130
rect 2749 4118 2784 4130
rect 2418 4116 2580 4118
rect 2313 4088 2354 4096
rect 2436 4092 2449 4116
rect 2464 4114 2479 4116
rect 2276 4078 2277 4088
rect 2292 4078 2305 4088
rect 2319 4078 2320 4088
rect 2335 4078 2348 4088
rect 2363 4078 2393 4092
rect 2436 4078 2479 4092
rect 2503 4089 2510 4096
rect 2513 4092 2580 4116
rect 2612 4116 2784 4118
rect 2582 4094 2610 4098
rect 2612 4094 2692 4116
rect 2713 4114 2728 4116
rect 2582 4092 2692 4094
rect 2513 4088 2692 4092
rect 2486 4078 2516 4088
rect 2518 4078 2671 4088
rect 2679 4078 2709 4088
rect 2713 4078 2743 4092
rect 2771 4078 2784 4116
rect 2856 4122 2891 4130
rect 2856 4096 2857 4122
rect 2864 4096 2891 4122
rect 2799 4078 2829 4092
rect 2856 4088 2891 4096
rect 2893 4122 2934 4130
rect 2893 4096 2908 4122
rect 2915 4096 2934 4122
rect 2998 4118 3060 4130
rect 3072 4118 3147 4130
rect 3205 4118 3280 4130
rect 3292 4118 3323 4130
rect 3329 4118 3364 4130
rect 2998 4116 3160 4118
rect 2893 4088 2934 4096
rect 3016 4092 3029 4116
rect 3044 4114 3059 4116
rect 2856 4078 2857 4088
rect 2872 4078 2885 4088
rect 2899 4078 2900 4088
rect 2915 4078 2928 4088
rect 2943 4078 2973 4092
rect 3016 4078 3059 4092
rect 3083 4089 3090 4096
rect 3093 4092 3160 4116
rect 3192 4116 3364 4118
rect 3162 4094 3190 4098
rect 3192 4094 3272 4116
rect 3293 4114 3308 4116
rect 3162 4092 3272 4094
rect 3093 4088 3272 4092
rect 3066 4078 3096 4088
rect 3098 4078 3251 4088
rect 3259 4078 3289 4088
rect 3293 4078 3323 4092
rect 3351 4078 3364 4116
rect 3436 4122 3471 4130
rect 3436 4096 3437 4122
rect 3444 4096 3471 4122
rect 3379 4078 3409 4092
rect 3436 4088 3471 4096
rect 3473 4122 3514 4130
rect 3473 4096 3488 4122
rect 3495 4096 3514 4122
rect 3578 4118 3640 4130
rect 3652 4118 3727 4130
rect 3785 4118 3860 4130
rect 3872 4118 3903 4130
rect 3909 4118 3944 4130
rect 3578 4116 3740 4118
rect 3473 4088 3514 4096
rect 3596 4092 3609 4116
rect 3624 4114 3639 4116
rect 3436 4078 3437 4088
rect 3452 4078 3465 4088
rect 3479 4078 3480 4088
rect 3495 4078 3508 4088
rect 3523 4078 3553 4092
rect 3596 4078 3639 4092
rect 3663 4089 3670 4096
rect 3673 4092 3740 4116
rect 3772 4116 3944 4118
rect 3742 4094 3770 4098
rect 3772 4094 3852 4116
rect 3873 4114 3888 4116
rect 3742 4092 3852 4094
rect 3673 4088 3852 4092
rect 3646 4078 3676 4088
rect 3678 4078 3831 4088
rect 3839 4078 3869 4088
rect 3873 4078 3903 4092
rect 3931 4078 3944 4116
rect 4016 4122 4051 4130
rect 4016 4096 4017 4122
rect 4024 4096 4051 4122
rect 3959 4078 3989 4092
rect 4016 4088 4051 4096
rect 4053 4122 4094 4130
rect 4053 4096 4068 4122
rect 4075 4096 4094 4122
rect 4158 4118 4220 4130
rect 4232 4118 4307 4130
rect 4365 4118 4440 4130
rect 4452 4118 4483 4130
rect 4489 4118 4524 4130
rect 4158 4116 4320 4118
rect 4053 4088 4094 4096
rect 4176 4092 4189 4116
rect 4204 4114 4219 4116
rect 4016 4078 4017 4088
rect 4032 4078 4045 4088
rect 4059 4078 4060 4088
rect 4075 4078 4088 4088
rect 4103 4078 4133 4092
rect 4176 4078 4219 4092
rect 4243 4089 4250 4096
rect 4253 4092 4320 4116
rect 4352 4116 4524 4118
rect 4322 4094 4350 4098
rect 4352 4094 4432 4116
rect 4453 4114 4468 4116
rect 4322 4092 4432 4094
rect 4253 4088 4432 4092
rect 4226 4078 4256 4088
rect 4258 4078 4411 4088
rect 4419 4078 4449 4088
rect 4453 4078 4483 4092
rect 4511 4078 4524 4116
rect 4596 4122 4631 4130
rect 4596 4096 4597 4122
rect 4604 4096 4631 4122
rect 4539 4078 4569 4092
rect 4596 4088 4631 4096
rect 4633 4122 4674 4130
rect 4633 4096 4648 4122
rect 4655 4096 4674 4122
rect 4738 4118 4800 4130
rect 4812 4118 4887 4130
rect 4945 4118 5020 4130
rect 5032 4118 5063 4130
rect 5069 4118 5104 4130
rect 4738 4116 4900 4118
rect 4633 4088 4674 4096
rect 4756 4092 4769 4116
rect 4784 4114 4799 4116
rect 4596 4078 4597 4088
rect 4612 4078 4625 4088
rect 4639 4078 4640 4088
rect 4655 4078 4668 4088
rect 4683 4078 4713 4092
rect 4756 4078 4799 4092
rect 4823 4089 4830 4096
rect 4833 4092 4900 4116
rect 4932 4116 5104 4118
rect 4902 4094 4930 4098
rect 4932 4094 5012 4116
rect 5033 4114 5048 4116
rect 4902 4092 5012 4094
rect 4833 4088 5012 4092
rect 4806 4078 4836 4088
rect 4838 4078 4991 4088
rect 4999 4078 5029 4088
rect 5033 4078 5063 4092
rect 5091 4078 5104 4116
rect 5176 4122 5211 4130
rect 5176 4096 5177 4122
rect 5184 4096 5211 4122
rect 5119 4078 5149 4092
rect 5176 4088 5211 4096
rect 5213 4122 5254 4130
rect 5213 4096 5228 4122
rect 5235 4096 5254 4122
rect 5318 4118 5380 4130
rect 5392 4118 5467 4130
rect 5525 4118 5600 4130
rect 5612 4118 5643 4130
rect 5649 4118 5684 4130
rect 5318 4116 5480 4118
rect 5213 4088 5254 4096
rect 5336 4092 5349 4116
rect 5364 4114 5379 4116
rect 5176 4078 5177 4088
rect 5192 4078 5205 4088
rect 5219 4078 5220 4088
rect 5235 4078 5248 4088
rect 5263 4078 5293 4092
rect 5336 4078 5379 4092
rect 5403 4089 5410 4096
rect 5413 4092 5480 4116
rect 5512 4116 5684 4118
rect 5482 4094 5510 4098
rect 5512 4094 5592 4116
rect 5613 4114 5628 4116
rect 5482 4092 5592 4094
rect 5413 4088 5592 4092
rect 5386 4078 5416 4088
rect 5418 4078 5571 4088
rect 5579 4078 5609 4088
rect 5613 4078 5643 4092
rect 5671 4078 5684 4116
rect 5756 4122 5791 4130
rect 5756 4096 5757 4122
rect 5764 4096 5791 4122
rect 5699 4078 5729 4092
rect 5756 4088 5791 4096
rect 5793 4122 5834 4130
rect 5793 4096 5808 4122
rect 5815 4096 5834 4122
rect 5898 4118 5960 4130
rect 5972 4118 6047 4130
rect 6105 4118 6180 4130
rect 6192 4118 6223 4130
rect 6229 4118 6264 4130
rect 5898 4116 6060 4118
rect 5793 4088 5834 4096
rect 5916 4092 5929 4116
rect 5944 4114 5959 4116
rect 5756 4078 5757 4088
rect 5772 4078 5785 4088
rect 5799 4078 5800 4088
rect 5815 4078 5828 4088
rect 5843 4078 5873 4092
rect 5916 4078 5959 4092
rect 5983 4089 5990 4096
rect 5993 4092 6060 4116
rect 6092 4116 6264 4118
rect 6062 4094 6090 4098
rect 6092 4094 6172 4116
rect 6193 4114 6208 4116
rect 6062 4092 6172 4094
rect 5993 4088 6172 4092
rect 5966 4078 5996 4088
rect 5998 4078 6151 4088
rect 6159 4078 6189 4088
rect 6193 4078 6223 4092
rect 6251 4078 6264 4116
rect 6336 4122 6371 4130
rect 6336 4096 6337 4122
rect 6344 4096 6371 4122
rect 6279 4078 6309 4092
rect 6336 4088 6371 4096
rect 6373 4122 6414 4130
rect 6373 4096 6388 4122
rect 6395 4096 6414 4122
rect 6478 4118 6540 4130
rect 6552 4118 6627 4130
rect 6685 4118 6760 4130
rect 6772 4118 6803 4130
rect 6809 4118 6844 4130
rect 6478 4116 6640 4118
rect 6373 4088 6414 4096
rect 6496 4092 6509 4116
rect 6524 4114 6539 4116
rect 6336 4078 6337 4088
rect 6352 4078 6365 4088
rect 6379 4078 6380 4088
rect 6395 4078 6408 4088
rect 6423 4078 6453 4092
rect 6496 4078 6539 4092
rect 6563 4089 6570 4096
rect 6573 4092 6640 4116
rect 6672 4116 6844 4118
rect 6642 4094 6670 4098
rect 6672 4094 6752 4116
rect 6773 4114 6788 4116
rect 6642 4092 6752 4094
rect 6573 4088 6752 4092
rect 6546 4078 6576 4088
rect 6578 4078 6731 4088
rect 6739 4078 6769 4088
rect 6773 4078 6803 4092
rect 6831 4078 6844 4116
rect 6916 4122 6951 4130
rect 6916 4096 6917 4122
rect 6924 4096 6951 4122
rect 6859 4078 6889 4092
rect 6916 4088 6951 4096
rect 6953 4122 6994 4130
rect 6953 4096 6968 4122
rect 6975 4096 6994 4122
rect 7058 4118 7120 4130
rect 7132 4118 7207 4130
rect 7265 4118 7340 4130
rect 7352 4118 7383 4130
rect 7389 4118 7424 4130
rect 7058 4116 7220 4118
rect 6953 4088 6994 4096
rect 7076 4092 7089 4116
rect 7104 4114 7119 4116
rect 6916 4078 6917 4088
rect 6932 4078 6945 4088
rect 6959 4078 6960 4088
rect 6975 4078 6988 4088
rect 7003 4078 7033 4092
rect 7076 4078 7119 4092
rect 7143 4089 7150 4096
rect 7153 4092 7220 4116
rect 7252 4116 7424 4118
rect 7222 4094 7250 4098
rect 7252 4094 7332 4116
rect 7353 4114 7368 4116
rect 7222 4092 7332 4094
rect 7153 4088 7332 4092
rect 7126 4078 7156 4088
rect 7158 4078 7311 4088
rect 7319 4078 7349 4088
rect 7353 4078 7383 4092
rect 7411 4078 7424 4116
rect 7496 4122 7531 4130
rect 7496 4096 7497 4122
rect 7504 4096 7531 4122
rect 7439 4078 7469 4092
rect 7496 4088 7531 4096
rect 7533 4122 7574 4130
rect 7533 4096 7548 4122
rect 7555 4096 7574 4122
rect 7638 4118 7700 4130
rect 7712 4118 7787 4130
rect 7845 4118 7920 4130
rect 7932 4118 7963 4130
rect 7969 4118 8004 4130
rect 7638 4116 7800 4118
rect 7533 4088 7574 4096
rect 7656 4092 7669 4116
rect 7684 4114 7699 4116
rect 7496 4078 7497 4088
rect 7512 4078 7525 4088
rect 7539 4078 7540 4088
rect 7555 4078 7568 4088
rect 7583 4078 7613 4092
rect 7656 4078 7699 4092
rect 7723 4089 7730 4096
rect 7733 4092 7800 4116
rect 7832 4116 8004 4118
rect 7802 4094 7830 4098
rect 7832 4094 7912 4116
rect 7933 4114 7948 4116
rect 7802 4092 7912 4094
rect 7733 4088 7912 4092
rect 7706 4078 7736 4088
rect 7738 4078 7891 4088
rect 7899 4078 7929 4088
rect 7933 4078 7963 4092
rect 7991 4078 8004 4116
rect 8076 4122 8111 4130
rect 8076 4096 8077 4122
rect 8084 4096 8111 4122
rect 8019 4078 8049 4092
rect 8076 4088 8111 4096
rect 8113 4122 8154 4130
rect 8113 4096 8128 4122
rect 8135 4096 8154 4122
rect 8218 4118 8280 4130
rect 8292 4118 8367 4130
rect 8425 4118 8500 4130
rect 8512 4118 8543 4130
rect 8549 4118 8584 4130
rect 8218 4116 8380 4118
rect 8113 4088 8154 4096
rect 8236 4092 8249 4116
rect 8264 4114 8279 4116
rect 8076 4078 8077 4088
rect 8092 4078 8105 4088
rect 8119 4078 8120 4088
rect 8135 4078 8148 4088
rect 8163 4078 8193 4092
rect 8236 4078 8279 4092
rect 8303 4089 8310 4096
rect 8313 4092 8380 4116
rect 8412 4116 8584 4118
rect 8382 4094 8410 4098
rect 8412 4094 8492 4116
rect 8513 4114 8528 4116
rect 8382 4092 8492 4094
rect 8313 4088 8492 4092
rect 8286 4078 8316 4088
rect 8318 4078 8471 4088
rect 8479 4078 8509 4088
rect 8513 4078 8543 4092
rect 8571 4078 8584 4116
rect 8656 4122 8691 4130
rect 8656 4096 8657 4122
rect 8664 4096 8691 4122
rect 8599 4078 8629 4092
rect 8656 4088 8691 4096
rect 8693 4122 8734 4130
rect 8693 4096 8708 4122
rect 8715 4096 8734 4122
rect 8798 4118 8860 4130
rect 8872 4118 8947 4130
rect 9005 4118 9080 4130
rect 9092 4118 9123 4130
rect 9129 4118 9164 4130
rect 8798 4116 8960 4118
rect 8693 4088 8734 4096
rect 8816 4092 8829 4116
rect 8844 4114 8859 4116
rect 8656 4078 8657 4088
rect 8672 4078 8685 4088
rect 8699 4078 8700 4088
rect 8715 4078 8728 4088
rect 8743 4078 8773 4092
rect 8816 4078 8859 4092
rect 8883 4089 8890 4096
rect 8893 4092 8960 4116
rect 8992 4116 9164 4118
rect 8962 4094 8990 4098
rect 8992 4094 9072 4116
rect 9093 4114 9108 4116
rect 8962 4092 9072 4094
rect 8893 4088 9072 4092
rect 8866 4078 8896 4088
rect 8898 4078 9051 4088
rect 9059 4078 9089 4088
rect 9093 4078 9123 4092
rect 9151 4078 9164 4116
rect 9236 4122 9271 4130
rect 9236 4096 9237 4122
rect 9244 4096 9271 4122
rect 9179 4078 9209 4092
rect 9236 4088 9271 4096
rect 9236 4078 9237 4088
rect 9252 4078 9265 4088
rect -1 4072 9265 4078
rect 0 4064 9265 4072
rect 15 4034 28 4064
rect 43 4046 73 4064
rect 116 4050 130 4064
rect 166 4050 386 4064
rect 117 4048 130 4050
rect 83 4036 98 4048
rect 80 4034 102 4036
rect 107 4034 137 4048
rect 198 4046 351 4050
rect 180 4034 372 4046
rect 415 4034 445 4048
rect 451 4034 464 4064
rect 479 4046 509 4064
rect 552 4034 565 4064
rect 595 4034 608 4064
rect 623 4046 653 4064
rect 696 4050 710 4064
rect 746 4050 966 4064
rect 697 4048 710 4050
rect 663 4036 678 4048
rect 660 4034 682 4036
rect 687 4034 717 4048
rect 778 4046 931 4050
rect 760 4034 952 4046
rect 995 4034 1025 4048
rect 1031 4034 1044 4064
rect 1059 4046 1089 4064
rect 1132 4034 1145 4064
rect 1175 4034 1188 4064
rect 1203 4046 1233 4064
rect 1276 4050 1290 4064
rect 1326 4050 1546 4064
rect 1277 4048 1290 4050
rect 1243 4036 1258 4048
rect 1240 4034 1262 4036
rect 1267 4034 1297 4048
rect 1358 4046 1511 4050
rect 1340 4034 1532 4046
rect 1575 4034 1605 4048
rect 1611 4034 1624 4064
rect 1639 4046 1669 4064
rect 1712 4034 1725 4064
rect 1755 4034 1768 4064
rect 1783 4046 1813 4064
rect 1856 4050 1870 4064
rect 1906 4050 2126 4064
rect 1857 4048 1870 4050
rect 1823 4036 1838 4048
rect 1820 4034 1842 4036
rect 1847 4034 1877 4048
rect 1938 4046 2091 4050
rect 1920 4034 2112 4046
rect 2155 4034 2185 4048
rect 2191 4034 2204 4064
rect 2219 4046 2249 4064
rect 2292 4034 2305 4064
rect 2335 4034 2348 4064
rect 2363 4046 2393 4064
rect 2436 4050 2450 4064
rect 2486 4050 2706 4064
rect 2437 4048 2450 4050
rect 2403 4036 2418 4048
rect 2400 4034 2422 4036
rect 2427 4034 2457 4048
rect 2518 4046 2671 4050
rect 2500 4034 2692 4046
rect 2735 4034 2765 4048
rect 2771 4034 2784 4064
rect 2799 4046 2829 4064
rect 2872 4034 2885 4064
rect 2915 4034 2928 4064
rect 2943 4046 2973 4064
rect 3016 4050 3030 4064
rect 3066 4050 3286 4064
rect 3017 4048 3030 4050
rect 2983 4036 2998 4048
rect 2980 4034 3002 4036
rect 3007 4034 3037 4048
rect 3098 4046 3251 4050
rect 3080 4034 3272 4046
rect 3315 4034 3345 4048
rect 3351 4034 3364 4064
rect 3379 4046 3409 4064
rect 3452 4034 3465 4064
rect 3495 4034 3508 4064
rect 3523 4046 3553 4064
rect 3596 4050 3610 4064
rect 3646 4050 3866 4064
rect 3597 4048 3610 4050
rect 3563 4036 3578 4048
rect 3560 4034 3582 4036
rect 3587 4034 3617 4048
rect 3678 4046 3831 4050
rect 3660 4034 3852 4046
rect 3895 4034 3925 4048
rect 3931 4034 3944 4064
rect 3959 4046 3989 4064
rect 4032 4034 4045 4064
rect 4075 4034 4088 4064
rect 4103 4046 4133 4064
rect 4176 4050 4190 4064
rect 4226 4050 4446 4064
rect 4177 4048 4190 4050
rect 4143 4036 4158 4048
rect 4140 4034 4162 4036
rect 4167 4034 4197 4048
rect 4258 4046 4411 4050
rect 4240 4034 4432 4046
rect 4475 4034 4505 4048
rect 4511 4034 4524 4064
rect 4539 4046 4569 4064
rect 4612 4034 4625 4064
rect 4655 4034 4668 4064
rect 4683 4046 4713 4064
rect 4756 4050 4770 4064
rect 4806 4050 5026 4064
rect 4757 4048 4770 4050
rect 4723 4036 4738 4048
rect 4720 4034 4742 4036
rect 4747 4034 4777 4048
rect 4838 4046 4991 4050
rect 4820 4034 5012 4046
rect 5055 4034 5085 4048
rect 5091 4034 5104 4064
rect 5119 4046 5149 4064
rect 5192 4034 5205 4064
rect 5235 4034 5248 4064
rect 5263 4046 5293 4064
rect 5336 4050 5350 4064
rect 5386 4050 5606 4064
rect 5337 4048 5350 4050
rect 5303 4036 5318 4048
rect 5300 4034 5322 4036
rect 5327 4034 5357 4048
rect 5418 4046 5571 4050
rect 5400 4034 5592 4046
rect 5635 4034 5665 4048
rect 5671 4034 5684 4064
rect 5699 4046 5729 4064
rect 5772 4034 5785 4064
rect 5815 4034 5828 4064
rect 5843 4046 5873 4064
rect 5916 4050 5930 4064
rect 5966 4050 6186 4064
rect 5917 4048 5930 4050
rect 5883 4036 5898 4048
rect 5880 4034 5902 4036
rect 5907 4034 5937 4048
rect 5998 4046 6151 4050
rect 5980 4034 6172 4046
rect 6215 4034 6245 4048
rect 6251 4034 6264 4064
rect 6279 4046 6309 4064
rect 6352 4034 6365 4064
rect 6395 4034 6408 4064
rect 6423 4046 6453 4064
rect 6496 4050 6510 4064
rect 6546 4050 6766 4064
rect 6497 4048 6510 4050
rect 6463 4036 6478 4048
rect 6460 4034 6482 4036
rect 6487 4034 6517 4048
rect 6578 4046 6731 4050
rect 6560 4034 6752 4046
rect 6795 4034 6825 4048
rect 6831 4034 6844 4064
rect 6859 4046 6889 4064
rect 6932 4034 6945 4064
rect 6975 4034 6988 4064
rect 7003 4046 7033 4064
rect 7076 4050 7090 4064
rect 7126 4050 7346 4064
rect 7077 4048 7090 4050
rect 7043 4036 7058 4048
rect 7040 4034 7062 4036
rect 7067 4034 7097 4048
rect 7158 4046 7311 4050
rect 7140 4034 7332 4046
rect 7375 4034 7405 4048
rect 7411 4034 7424 4064
rect 7439 4046 7469 4064
rect 7512 4034 7525 4064
rect 7555 4034 7568 4064
rect 7583 4046 7613 4064
rect 7656 4050 7670 4064
rect 7706 4050 7926 4064
rect 7657 4048 7670 4050
rect 7623 4036 7638 4048
rect 7620 4034 7642 4036
rect 7647 4034 7677 4048
rect 7738 4046 7891 4050
rect 7720 4034 7912 4046
rect 7955 4034 7985 4048
rect 7991 4034 8004 4064
rect 8019 4046 8049 4064
rect 8092 4034 8105 4064
rect 8135 4034 8148 4064
rect 8163 4046 8193 4064
rect 8236 4050 8250 4064
rect 8286 4050 8506 4064
rect 8237 4048 8250 4050
rect 8203 4036 8218 4048
rect 8200 4034 8222 4036
rect 8227 4034 8257 4048
rect 8318 4046 8471 4050
rect 8300 4034 8492 4046
rect 8535 4034 8565 4048
rect 8571 4034 8584 4064
rect 8599 4046 8629 4064
rect 8672 4034 8685 4064
rect 8715 4034 8728 4064
rect 8743 4046 8773 4064
rect 8816 4050 8830 4064
rect 8866 4050 9086 4064
rect 8817 4048 8830 4050
rect 8783 4036 8798 4048
rect 8780 4034 8802 4036
rect 8807 4034 8837 4048
rect 8898 4046 9051 4050
rect 8880 4034 9072 4046
rect 9115 4034 9145 4048
rect 9151 4034 9164 4064
rect 9179 4046 9209 4064
rect 9252 4034 9265 4064
rect 0 4020 9265 4034
rect 15 3916 28 4020
rect 73 3998 74 4008
rect 89 3998 102 4008
rect 73 3994 102 3998
rect 107 3994 137 4020
rect 155 4006 171 4008
rect 243 4006 296 4020
rect 244 4004 308 4006
rect 351 4004 366 4020
rect 415 4017 445 4020
rect 415 4014 451 4017
rect 381 4006 397 4008
rect 155 3994 170 3998
rect 73 3992 170 3994
rect 198 3992 366 4004
rect 382 3994 397 3998
rect 415 3995 454 4014
rect 473 4008 480 4009
rect 479 4001 480 4008
rect 463 3998 464 4001
rect 479 3998 492 4001
rect 415 3994 445 3995
rect 454 3994 460 3995
rect 463 3994 492 3998
rect 382 3993 492 3994
rect 382 3992 498 3993
rect 57 3984 108 3992
rect 57 3972 82 3984
rect 89 3972 108 3984
rect 139 3984 189 3992
rect 139 3976 155 3984
rect 162 3982 189 3984
rect 198 3982 419 3992
rect 162 3972 419 3982
rect 448 3984 498 3992
rect 448 3975 464 3984
rect 57 3964 108 3972
rect 155 3964 419 3972
rect 445 3972 464 3975
rect 471 3972 498 3984
rect 445 3964 498 3972
rect 73 3956 74 3964
rect 89 3956 102 3964
rect 73 3948 89 3956
rect 70 3941 89 3944
rect 70 3932 92 3941
rect 43 3922 92 3932
rect 43 3916 73 3922
rect 92 3917 97 3922
rect 15 3900 89 3916
rect 107 3908 137 3964
rect 172 3954 380 3964
rect 415 3960 460 3964
rect 463 3963 464 3964
rect 479 3963 492 3964
rect 198 3924 387 3954
rect 213 3921 387 3924
rect 206 3918 387 3921
rect 15 3898 28 3900
rect 43 3898 77 3900
rect 15 3882 89 3898
rect 116 3894 129 3908
rect 144 3894 160 3910
rect 206 3905 217 3918
rect -1 3860 0 3876
rect 15 3860 28 3882
rect 43 3860 73 3882
rect 116 3878 178 3894
rect 206 3887 217 3903
rect 222 3898 232 3918
rect 242 3898 256 3918
rect 259 3905 268 3918
rect 284 3905 293 3918
rect 222 3887 256 3898
rect 259 3887 268 3903
rect 284 3887 293 3903
rect 300 3898 310 3918
rect 320 3898 334 3918
rect 335 3905 346 3918
rect 300 3887 334 3898
rect 335 3887 346 3903
rect 392 3894 408 3910
rect 415 3908 445 3960
rect 479 3956 480 3963
rect 464 3948 480 3956
rect 451 3916 464 3935
rect 479 3916 509 3932
rect 451 3900 525 3916
rect 451 3898 464 3900
rect 479 3898 513 3900
rect 116 3876 129 3878
rect 144 3876 178 3878
rect 116 3860 178 3876
rect 222 3871 238 3874
rect 300 3871 330 3882
rect 378 3878 424 3894
rect 451 3882 525 3898
rect 378 3876 412 3878
rect 377 3860 424 3876
rect 451 3860 464 3882
rect 479 3860 509 3882
rect 536 3860 537 3876
rect 552 3860 565 4020
rect 595 3916 608 4020
rect 653 3998 654 4008
rect 669 3998 682 4008
rect 653 3994 682 3998
rect 687 3994 717 4020
rect 735 4006 751 4008
rect 823 4006 876 4020
rect 824 4004 888 4006
rect 931 4004 946 4020
rect 995 4017 1025 4020
rect 995 4014 1031 4017
rect 961 4006 977 4008
rect 735 3994 750 3998
rect 653 3992 750 3994
rect 778 3992 946 4004
rect 962 3994 977 3998
rect 995 3995 1034 4014
rect 1053 4008 1060 4009
rect 1059 4001 1060 4008
rect 1043 3998 1044 4001
rect 1059 3998 1072 4001
rect 995 3994 1025 3995
rect 1034 3994 1040 3995
rect 1043 3994 1072 3998
rect 962 3993 1072 3994
rect 962 3992 1078 3993
rect 637 3984 688 3992
rect 637 3972 662 3984
rect 669 3972 688 3984
rect 719 3984 769 3992
rect 719 3976 735 3984
rect 742 3982 769 3984
rect 778 3982 999 3992
rect 742 3972 999 3982
rect 1028 3984 1078 3992
rect 1028 3975 1044 3984
rect 637 3964 688 3972
rect 735 3964 999 3972
rect 1025 3972 1044 3975
rect 1051 3972 1078 3984
rect 1025 3964 1078 3972
rect 653 3956 654 3964
rect 669 3956 682 3964
rect 653 3948 669 3956
rect 650 3941 669 3944
rect 650 3932 672 3941
rect 623 3922 672 3932
rect 623 3916 653 3922
rect 672 3917 677 3922
rect 595 3900 669 3916
rect 687 3908 717 3964
rect 752 3954 960 3964
rect 995 3960 1040 3964
rect 1043 3963 1044 3964
rect 1059 3963 1072 3964
rect 778 3924 967 3954
rect 793 3921 967 3924
rect 786 3918 967 3921
rect 595 3898 608 3900
rect 623 3898 657 3900
rect 595 3882 669 3898
rect 696 3894 709 3908
rect 724 3894 740 3910
rect 786 3905 797 3918
rect 579 3860 580 3876
rect 595 3860 608 3882
rect 623 3860 653 3882
rect 696 3878 758 3894
rect 786 3887 797 3903
rect 802 3898 812 3918
rect 822 3898 836 3918
rect 839 3905 848 3918
rect 864 3905 873 3918
rect 802 3887 836 3898
rect 839 3887 848 3903
rect 864 3887 873 3903
rect 880 3898 890 3918
rect 900 3898 914 3918
rect 915 3905 926 3918
rect 880 3887 914 3898
rect 915 3887 926 3903
rect 972 3894 988 3910
rect 995 3908 1025 3960
rect 1059 3956 1060 3963
rect 1044 3948 1060 3956
rect 1031 3916 1044 3935
rect 1059 3916 1089 3932
rect 1031 3900 1105 3916
rect 1031 3898 1044 3900
rect 1059 3898 1093 3900
rect 696 3876 709 3878
rect 724 3876 758 3878
rect 696 3860 758 3876
rect 802 3871 818 3874
rect 880 3871 910 3882
rect 958 3878 1004 3894
rect 1031 3882 1105 3898
rect 958 3876 992 3878
rect 957 3860 1004 3876
rect 1031 3860 1044 3882
rect 1059 3860 1089 3882
rect 1116 3860 1117 3876
rect 1132 3860 1145 4020
rect 1175 3916 1188 4020
rect 1233 3998 1234 4008
rect 1249 3998 1262 4008
rect 1233 3994 1262 3998
rect 1267 3994 1297 4020
rect 1315 4006 1331 4008
rect 1403 4006 1456 4020
rect 1404 4004 1468 4006
rect 1511 4004 1526 4020
rect 1575 4017 1605 4020
rect 1575 4014 1611 4017
rect 1541 4006 1557 4008
rect 1315 3994 1330 3998
rect 1233 3992 1330 3994
rect 1358 3992 1526 4004
rect 1542 3994 1557 3998
rect 1575 3995 1614 4014
rect 1633 4008 1640 4009
rect 1639 4001 1640 4008
rect 1623 3998 1624 4001
rect 1639 3998 1652 4001
rect 1575 3994 1605 3995
rect 1614 3994 1620 3995
rect 1623 3994 1652 3998
rect 1542 3993 1652 3994
rect 1542 3992 1658 3993
rect 1217 3984 1268 3992
rect 1217 3972 1242 3984
rect 1249 3972 1268 3984
rect 1299 3984 1349 3992
rect 1299 3976 1315 3984
rect 1322 3982 1349 3984
rect 1358 3982 1579 3992
rect 1322 3972 1579 3982
rect 1608 3984 1658 3992
rect 1608 3975 1624 3984
rect 1217 3964 1268 3972
rect 1315 3964 1579 3972
rect 1605 3972 1624 3975
rect 1631 3972 1658 3984
rect 1605 3964 1658 3972
rect 1233 3956 1234 3964
rect 1249 3956 1262 3964
rect 1233 3948 1249 3956
rect 1230 3941 1249 3944
rect 1230 3932 1252 3941
rect 1203 3922 1252 3932
rect 1203 3916 1233 3922
rect 1252 3917 1257 3922
rect 1175 3900 1249 3916
rect 1267 3908 1297 3964
rect 1332 3954 1540 3964
rect 1575 3960 1620 3964
rect 1623 3963 1624 3964
rect 1639 3963 1652 3964
rect 1358 3924 1547 3954
rect 1373 3921 1547 3924
rect 1366 3918 1547 3921
rect 1175 3898 1188 3900
rect 1203 3898 1237 3900
rect 1175 3882 1249 3898
rect 1276 3894 1289 3908
rect 1304 3894 1320 3910
rect 1366 3905 1377 3918
rect 1159 3860 1160 3876
rect 1175 3860 1188 3882
rect 1203 3860 1233 3882
rect 1276 3878 1338 3894
rect 1366 3887 1377 3903
rect 1382 3898 1392 3918
rect 1402 3898 1416 3918
rect 1419 3905 1428 3918
rect 1444 3905 1453 3918
rect 1382 3887 1416 3898
rect 1419 3887 1428 3903
rect 1444 3887 1453 3903
rect 1460 3898 1470 3918
rect 1480 3898 1494 3918
rect 1495 3905 1506 3918
rect 1460 3887 1494 3898
rect 1495 3887 1506 3903
rect 1552 3894 1568 3910
rect 1575 3908 1605 3960
rect 1639 3956 1640 3963
rect 1624 3948 1640 3956
rect 1611 3916 1624 3935
rect 1639 3916 1669 3932
rect 1611 3900 1685 3916
rect 1611 3898 1624 3900
rect 1639 3898 1673 3900
rect 1276 3876 1289 3878
rect 1304 3876 1338 3878
rect 1276 3860 1338 3876
rect 1382 3871 1398 3874
rect 1460 3871 1490 3882
rect 1538 3878 1584 3894
rect 1611 3882 1685 3898
rect 1538 3876 1572 3878
rect 1537 3860 1584 3876
rect 1611 3860 1624 3882
rect 1639 3860 1669 3882
rect 1696 3860 1697 3876
rect 1712 3860 1725 4020
rect 1755 3916 1768 4020
rect 1813 3998 1814 4008
rect 1829 3998 1842 4008
rect 1813 3994 1842 3998
rect 1847 3994 1877 4020
rect 1895 4006 1911 4008
rect 1983 4006 2036 4020
rect 1984 4004 2048 4006
rect 2091 4004 2106 4020
rect 2155 4017 2185 4020
rect 2155 4014 2191 4017
rect 2121 4006 2137 4008
rect 1895 3994 1910 3998
rect 1813 3992 1910 3994
rect 1938 3992 2106 4004
rect 2122 3994 2137 3998
rect 2155 3995 2194 4014
rect 2213 4008 2220 4009
rect 2219 4001 2220 4008
rect 2203 3998 2204 4001
rect 2219 3998 2232 4001
rect 2155 3994 2185 3995
rect 2194 3994 2200 3995
rect 2203 3994 2232 3998
rect 2122 3993 2232 3994
rect 2122 3992 2238 3993
rect 1797 3984 1848 3992
rect 1797 3972 1822 3984
rect 1829 3972 1848 3984
rect 1879 3984 1929 3992
rect 1879 3976 1895 3984
rect 1902 3982 1929 3984
rect 1938 3982 2159 3992
rect 1902 3972 2159 3982
rect 2188 3984 2238 3992
rect 2188 3975 2204 3984
rect 1797 3964 1848 3972
rect 1895 3964 2159 3972
rect 2185 3972 2204 3975
rect 2211 3972 2238 3984
rect 2185 3964 2238 3972
rect 1813 3956 1814 3964
rect 1829 3956 1842 3964
rect 1813 3948 1829 3956
rect 1810 3941 1829 3944
rect 1810 3932 1832 3941
rect 1783 3922 1832 3932
rect 1783 3916 1813 3922
rect 1832 3917 1837 3922
rect 1755 3900 1829 3916
rect 1847 3908 1877 3964
rect 1912 3954 2120 3964
rect 2155 3960 2200 3964
rect 2203 3963 2204 3964
rect 2219 3963 2232 3964
rect 1938 3924 2127 3954
rect 1953 3921 2127 3924
rect 1946 3918 2127 3921
rect 1755 3898 1768 3900
rect 1783 3898 1817 3900
rect 1755 3882 1829 3898
rect 1856 3894 1869 3908
rect 1884 3894 1900 3910
rect 1946 3905 1957 3918
rect 1739 3860 1740 3876
rect 1755 3860 1768 3882
rect 1783 3860 1813 3882
rect 1856 3878 1918 3894
rect 1946 3887 1957 3903
rect 1962 3898 1972 3918
rect 1982 3898 1996 3918
rect 1999 3905 2008 3918
rect 2024 3905 2033 3918
rect 1962 3887 1996 3898
rect 1999 3887 2008 3903
rect 2024 3887 2033 3903
rect 2040 3898 2050 3918
rect 2060 3898 2074 3918
rect 2075 3905 2086 3918
rect 2040 3887 2074 3898
rect 2075 3887 2086 3903
rect 2132 3894 2148 3910
rect 2155 3908 2185 3960
rect 2219 3956 2220 3963
rect 2204 3948 2220 3956
rect 2191 3916 2204 3935
rect 2219 3916 2249 3932
rect 2191 3900 2265 3916
rect 2191 3898 2204 3900
rect 2219 3898 2253 3900
rect 1856 3876 1869 3878
rect 1884 3876 1918 3878
rect 1856 3860 1918 3876
rect 1962 3871 1976 3874
rect 2040 3871 2070 3882
rect 2118 3878 2164 3894
rect 2191 3882 2265 3898
rect 2118 3876 2152 3878
rect 2117 3860 2164 3876
rect 2191 3860 2204 3882
rect 2219 3860 2249 3882
rect 2276 3860 2277 3876
rect 2292 3860 2305 4020
rect 2335 3916 2348 4020
rect 2393 3998 2394 4008
rect 2409 3998 2422 4008
rect 2393 3994 2422 3998
rect 2427 3994 2457 4020
rect 2475 4006 2491 4008
rect 2563 4006 2616 4020
rect 2564 4004 2628 4006
rect 2671 4004 2686 4020
rect 2735 4017 2765 4020
rect 2735 4014 2771 4017
rect 2701 4006 2717 4008
rect 2475 3994 2490 3998
rect 2393 3992 2490 3994
rect 2518 3992 2686 4004
rect 2702 3994 2717 3998
rect 2735 3995 2774 4014
rect 2793 4008 2800 4009
rect 2799 4001 2800 4008
rect 2783 3998 2784 4001
rect 2799 3998 2812 4001
rect 2735 3994 2765 3995
rect 2774 3994 2780 3995
rect 2783 3994 2812 3998
rect 2702 3993 2812 3994
rect 2702 3992 2818 3993
rect 2377 3984 2428 3992
rect 2377 3972 2402 3984
rect 2409 3972 2428 3984
rect 2459 3984 2509 3992
rect 2459 3976 2475 3984
rect 2482 3982 2509 3984
rect 2518 3982 2739 3992
rect 2482 3972 2739 3982
rect 2768 3984 2818 3992
rect 2768 3975 2784 3984
rect 2377 3964 2428 3972
rect 2475 3964 2739 3972
rect 2765 3972 2784 3975
rect 2791 3972 2818 3984
rect 2765 3964 2818 3972
rect 2393 3956 2394 3964
rect 2409 3956 2422 3964
rect 2393 3948 2409 3956
rect 2390 3941 2409 3944
rect 2390 3932 2412 3941
rect 2363 3922 2412 3932
rect 2363 3916 2393 3922
rect 2412 3917 2417 3922
rect 2335 3900 2409 3916
rect 2427 3908 2457 3964
rect 2492 3954 2700 3964
rect 2735 3960 2780 3964
rect 2783 3963 2784 3964
rect 2799 3963 2812 3964
rect 2518 3924 2707 3954
rect 2533 3921 2707 3924
rect 2526 3918 2707 3921
rect 2335 3898 2348 3900
rect 2363 3898 2397 3900
rect 2335 3882 2409 3898
rect 2436 3894 2449 3908
rect 2464 3894 2480 3910
rect 2526 3905 2537 3918
rect 2319 3860 2320 3876
rect 2335 3860 2348 3882
rect 2363 3860 2393 3882
rect 2436 3878 2498 3894
rect 2526 3887 2537 3903
rect 2542 3898 2552 3918
rect 2562 3898 2576 3918
rect 2579 3905 2588 3918
rect 2604 3905 2613 3918
rect 2542 3887 2576 3898
rect 2579 3887 2588 3903
rect 2604 3887 2613 3903
rect 2620 3898 2630 3918
rect 2640 3898 2654 3918
rect 2655 3905 2666 3918
rect 2620 3887 2654 3898
rect 2655 3887 2666 3903
rect 2712 3894 2728 3910
rect 2735 3908 2765 3960
rect 2799 3956 2800 3963
rect 2784 3948 2800 3956
rect 2771 3916 2784 3935
rect 2799 3916 2829 3932
rect 2771 3900 2845 3916
rect 2771 3898 2784 3900
rect 2799 3898 2833 3900
rect 2436 3876 2449 3878
rect 2464 3876 2498 3878
rect 2436 3860 2498 3876
rect 2542 3871 2558 3874
rect 2620 3871 2650 3882
rect 2698 3878 2744 3894
rect 2771 3882 2845 3898
rect 2698 3876 2732 3878
rect 2697 3860 2744 3876
rect 2771 3860 2784 3882
rect 2799 3860 2829 3882
rect 2856 3860 2857 3876
rect 2872 3860 2885 4020
rect 2915 3916 2928 4020
rect 2973 3998 2974 4008
rect 2989 3998 3002 4008
rect 2973 3994 3002 3998
rect 3007 3994 3037 4020
rect 3055 4006 3071 4008
rect 3143 4006 3196 4020
rect 3144 4004 3208 4006
rect 3251 4004 3266 4020
rect 3315 4017 3345 4020
rect 3315 4014 3351 4017
rect 3281 4006 3297 4008
rect 3055 3994 3070 3998
rect 2973 3992 3070 3994
rect 3098 3992 3266 4004
rect 3282 3994 3297 3998
rect 3315 3995 3354 4014
rect 3373 4008 3380 4009
rect 3379 4001 3380 4008
rect 3363 3998 3364 4001
rect 3379 3998 3392 4001
rect 3315 3994 3345 3995
rect 3354 3994 3360 3995
rect 3363 3994 3392 3998
rect 3282 3993 3392 3994
rect 3282 3992 3398 3993
rect 2957 3984 3008 3992
rect 2957 3972 2982 3984
rect 2989 3972 3008 3984
rect 3039 3984 3089 3992
rect 3039 3976 3055 3984
rect 3062 3982 3089 3984
rect 3098 3982 3319 3992
rect 3062 3972 3319 3982
rect 3348 3984 3398 3992
rect 3348 3975 3364 3984
rect 2957 3964 3008 3972
rect 3055 3964 3319 3972
rect 3345 3972 3364 3975
rect 3371 3972 3398 3984
rect 3345 3964 3398 3972
rect 2973 3956 2974 3964
rect 2989 3956 3002 3964
rect 2973 3948 2989 3956
rect 2970 3941 2989 3944
rect 2970 3932 2992 3941
rect 2943 3922 2992 3932
rect 2943 3916 2973 3922
rect 2992 3917 2997 3922
rect 2915 3900 2989 3916
rect 3007 3908 3037 3964
rect 3072 3954 3280 3964
rect 3315 3960 3360 3964
rect 3363 3963 3364 3964
rect 3379 3963 3392 3964
rect 3098 3924 3287 3954
rect 3113 3921 3287 3924
rect 3106 3918 3287 3921
rect 2915 3898 2928 3900
rect 2943 3898 2977 3900
rect 2915 3882 2989 3898
rect 3016 3894 3029 3908
rect 3044 3894 3060 3910
rect 3106 3905 3117 3918
rect 2899 3860 2900 3876
rect 2915 3860 2928 3882
rect 2943 3860 2973 3882
rect 3016 3878 3078 3894
rect 3106 3887 3117 3903
rect 3122 3898 3132 3918
rect 3142 3898 3156 3918
rect 3159 3905 3168 3918
rect 3184 3905 3193 3918
rect 3122 3887 3156 3898
rect 3159 3887 3168 3903
rect 3184 3887 3193 3903
rect 3200 3898 3210 3918
rect 3220 3898 3234 3918
rect 3235 3905 3246 3918
rect 3200 3887 3234 3898
rect 3235 3887 3246 3903
rect 3292 3894 3308 3910
rect 3315 3908 3345 3960
rect 3379 3956 3380 3963
rect 3364 3948 3380 3956
rect 3351 3916 3364 3935
rect 3379 3916 3409 3932
rect 3351 3900 3425 3916
rect 3351 3898 3364 3900
rect 3379 3898 3413 3900
rect 3016 3876 3029 3878
rect 3044 3876 3078 3878
rect 3016 3860 3078 3876
rect 3122 3871 3138 3874
rect 3200 3871 3230 3882
rect 3278 3878 3324 3894
rect 3351 3882 3425 3898
rect 3278 3876 3312 3878
rect 3277 3860 3324 3876
rect 3351 3860 3364 3882
rect 3379 3860 3409 3882
rect 3436 3860 3437 3876
rect 3452 3860 3465 4020
rect 3495 3916 3508 4020
rect 3553 3998 3554 4008
rect 3569 3998 3582 4008
rect 3553 3994 3582 3998
rect 3587 3994 3617 4020
rect 3635 4006 3651 4008
rect 3723 4006 3776 4020
rect 3724 4004 3788 4006
rect 3831 4004 3846 4020
rect 3895 4017 3925 4020
rect 3895 4014 3931 4017
rect 3861 4006 3877 4008
rect 3635 3994 3650 3998
rect 3553 3992 3650 3994
rect 3678 3992 3846 4004
rect 3862 3994 3877 3998
rect 3895 3995 3934 4014
rect 3953 4008 3960 4009
rect 3959 4001 3960 4008
rect 3943 3998 3944 4001
rect 3959 3998 3972 4001
rect 3895 3994 3925 3995
rect 3934 3994 3940 3995
rect 3943 3994 3972 3998
rect 3862 3993 3972 3994
rect 3862 3992 3978 3993
rect 3537 3984 3588 3992
rect 3537 3972 3562 3984
rect 3569 3972 3588 3984
rect 3619 3984 3669 3992
rect 3619 3976 3635 3984
rect 3642 3982 3669 3984
rect 3678 3982 3899 3992
rect 3642 3972 3899 3982
rect 3928 3984 3978 3992
rect 3928 3975 3944 3984
rect 3537 3964 3588 3972
rect 3635 3964 3899 3972
rect 3925 3972 3944 3975
rect 3951 3972 3978 3984
rect 3925 3964 3978 3972
rect 3553 3956 3554 3964
rect 3569 3956 3582 3964
rect 3553 3948 3569 3956
rect 3550 3941 3569 3944
rect 3550 3932 3572 3941
rect 3523 3922 3572 3932
rect 3523 3916 3553 3922
rect 3572 3917 3577 3922
rect 3495 3900 3569 3916
rect 3587 3908 3617 3964
rect 3652 3954 3860 3964
rect 3895 3960 3940 3964
rect 3943 3963 3944 3964
rect 3959 3963 3972 3964
rect 3678 3924 3867 3954
rect 3693 3921 3867 3924
rect 3686 3918 3867 3921
rect 3495 3898 3508 3900
rect 3523 3898 3557 3900
rect 3495 3882 3569 3898
rect 3596 3894 3609 3908
rect 3624 3894 3640 3910
rect 3686 3905 3697 3918
rect 3479 3860 3480 3876
rect 3495 3860 3508 3882
rect 3523 3860 3553 3882
rect 3596 3878 3658 3894
rect 3686 3887 3697 3903
rect 3702 3898 3712 3918
rect 3722 3898 3736 3918
rect 3739 3905 3748 3918
rect 3764 3905 3773 3918
rect 3702 3887 3736 3898
rect 3739 3887 3748 3903
rect 3764 3887 3773 3903
rect 3780 3898 3790 3918
rect 3800 3898 3814 3918
rect 3815 3905 3826 3918
rect 3780 3887 3814 3898
rect 3815 3887 3826 3903
rect 3872 3894 3888 3910
rect 3895 3908 3925 3960
rect 3959 3956 3960 3963
rect 3944 3948 3960 3956
rect 3931 3916 3944 3935
rect 3959 3916 3989 3932
rect 3931 3900 4005 3916
rect 3931 3898 3944 3900
rect 3959 3898 3993 3900
rect 3596 3876 3609 3878
rect 3624 3876 3658 3878
rect 3596 3860 3658 3876
rect 3702 3871 3718 3874
rect 3780 3871 3810 3882
rect 3858 3878 3904 3894
rect 3931 3882 4005 3898
rect 3858 3876 3892 3878
rect 3857 3860 3904 3876
rect 3931 3860 3944 3882
rect 3959 3860 3989 3882
rect 4016 3860 4017 3876
rect 4032 3860 4045 4020
rect 4075 3916 4088 4020
rect 4133 3998 4134 4008
rect 4149 3998 4162 4008
rect 4133 3994 4162 3998
rect 4167 3994 4197 4020
rect 4215 4006 4231 4008
rect 4303 4006 4356 4020
rect 4304 4004 4368 4006
rect 4411 4004 4426 4020
rect 4475 4017 4505 4020
rect 4475 4014 4511 4017
rect 4441 4006 4457 4008
rect 4215 3994 4230 3998
rect 4133 3992 4230 3994
rect 4258 3992 4426 4004
rect 4442 3994 4457 3998
rect 4475 3995 4514 4014
rect 4533 4008 4540 4009
rect 4539 4001 4540 4008
rect 4523 3998 4524 4001
rect 4539 3998 4552 4001
rect 4475 3994 4505 3995
rect 4514 3994 4520 3995
rect 4523 3994 4552 3998
rect 4442 3993 4552 3994
rect 4442 3992 4558 3993
rect 4117 3984 4168 3992
rect 4117 3972 4142 3984
rect 4149 3972 4168 3984
rect 4199 3984 4249 3992
rect 4199 3976 4215 3984
rect 4222 3982 4249 3984
rect 4258 3982 4479 3992
rect 4222 3972 4479 3982
rect 4508 3984 4558 3992
rect 4508 3975 4524 3984
rect 4117 3964 4168 3972
rect 4215 3964 4479 3972
rect 4505 3972 4524 3975
rect 4531 3972 4558 3984
rect 4505 3964 4558 3972
rect 4133 3956 4134 3964
rect 4149 3956 4162 3964
rect 4133 3948 4149 3956
rect 4130 3941 4149 3944
rect 4130 3932 4152 3941
rect 4103 3922 4152 3932
rect 4103 3916 4133 3922
rect 4152 3917 4157 3922
rect 4075 3900 4149 3916
rect 4167 3908 4197 3964
rect 4232 3954 4440 3964
rect 4475 3960 4520 3964
rect 4523 3963 4524 3964
rect 4539 3963 4552 3964
rect 4258 3924 4447 3954
rect 4273 3921 4447 3924
rect 4266 3918 4447 3921
rect 4075 3898 4088 3900
rect 4103 3898 4137 3900
rect 4075 3882 4149 3898
rect 4176 3894 4189 3908
rect 4204 3894 4220 3910
rect 4266 3905 4277 3918
rect 4059 3860 4060 3876
rect 4075 3860 4088 3882
rect 4103 3860 4133 3882
rect 4176 3878 4238 3894
rect 4266 3887 4277 3903
rect 4282 3898 4292 3918
rect 4302 3898 4316 3918
rect 4319 3905 4328 3918
rect 4344 3905 4353 3918
rect 4282 3887 4316 3898
rect 4319 3887 4328 3903
rect 4344 3887 4353 3903
rect 4360 3898 4370 3918
rect 4380 3898 4394 3918
rect 4395 3905 4406 3918
rect 4360 3887 4394 3898
rect 4395 3887 4406 3903
rect 4452 3894 4468 3910
rect 4475 3908 4505 3960
rect 4539 3956 4540 3963
rect 4524 3948 4540 3956
rect 4511 3916 4524 3935
rect 4539 3916 4569 3932
rect 4511 3900 4585 3916
rect 4511 3898 4524 3900
rect 4539 3898 4573 3900
rect 4176 3876 4189 3878
rect 4204 3876 4238 3878
rect 4176 3860 4238 3876
rect 4282 3871 4298 3874
rect 4360 3871 4390 3882
rect 4438 3878 4484 3894
rect 4511 3882 4585 3898
rect 4438 3876 4472 3878
rect 4437 3860 4484 3876
rect 4511 3860 4524 3882
rect 4539 3860 4569 3882
rect 4596 3860 4597 3876
rect 4612 3860 4625 4020
rect 4655 3916 4668 4020
rect 4713 3998 4714 4008
rect 4729 3998 4742 4008
rect 4713 3994 4742 3998
rect 4747 3994 4777 4020
rect 4795 4006 4811 4008
rect 4883 4006 4936 4020
rect 4884 4004 4948 4006
rect 4991 4004 5006 4020
rect 5055 4017 5085 4020
rect 5055 4014 5091 4017
rect 5021 4006 5037 4008
rect 4795 3994 4810 3998
rect 4713 3992 4810 3994
rect 4838 3992 5006 4004
rect 5022 3994 5037 3998
rect 5055 3995 5094 4014
rect 5113 4008 5120 4009
rect 5119 4001 5120 4008
rect 5103 3998 5104 4001
rect 5119 3998 5132 4001
rect 5055 3994 5085 3995
rect 5094 3994 5100 3995
rect 5103 3994 5132 3998
rect 5022 3993 5132 3994
rect 5022 3992 5138 3993
rect 4697 3984 4748 3992
rect 4697 3972 4722 3984
rect 4729 3972 4748 3984
rect 4779 3984 4829 3992
rect 4779 3976 4795 3984
rect 4802 3982 4829 3984
rect 4838 3982 5059 3992
rect 4802 3972 5059 3982
rect 5088 3984 5138 3992
rect 5088 3975 5104 3984
rect 4697 3964 4748 3972
rect 4795 3964 5059 3972
rect 5085 3972 5104 3975
rect 5111 3972 5138 3984
rect 5085 3964 5138 3972
rect 4713 3956 4714 3964
rect 4729 3956 4742 3964
rect 4713 3948 4729 3956
rect 4710 3941 4729 3944
rect 4710 3932 4732 3941
rect 4683 3922 4732 3932
rect 4683 3916 4713 3922
rect 4732 3917 4737 3922
rect 4655 3900 4729 3916
rect 4747 3908 4777 3964
rect 4812 3954 5020 3964
rect 5055 3960 5100 3964
rect 5103 3963 5104 3964
rect 5119 3963 5132 3964
rect 4838 3924 5027 3954
rect 4853 3921 5027 3924
rect 4846 3918 5027 3921
rect 4655 3898 4668 3900
rect 4683 3898 4717 3900
rect 4655 3882 4729 3898
rect 4756 3894 4769 3908
rect 4784 3894 4800 3910
rect 4846 3905 4857 3918
rect 4639 3860 4640 3876
rect 4655 3860 4668 3882
rect 4683 3860 4713 3882
rect 4756 3878 4818 3894
rect 4846 3887 4857 3903
rect 4862 3898 4872 3918
rect 4882 3898 4896 3918
rect 4899 3905 4908 3918
rect 4924 3905 4933 3918
rect 4862 3887 4896 3898
rect 4899 3887 4908 3903
rect 4924 3887 4933 3903
rect 4940 3898 4950 3918
rect 4960 3898 4974 3918
rect 4975 3905 4986 3918
rect 4940 3887 4974 3898
rect 4975 3887 4986 3903
rect 5032 3894 5048 3910
rect 5055 3908 5085 3960
rect 5119 3956 5120 3963
rect 5104 3948 5120 3956
rect 5091 3916 5104 3935
rect 5119 3916 5149 3932
rect 5091 3900 5165 3916
rect 5091 3898 5104 3900
rect 5119 3898 5153 3900
rect 4756 3876 4769 3878
rect 4784 3876 4818 3878
rect 4756 3860 4818 3876
rect 4862 3871 4878 3874
rect 4940 3871 4970 3882
rect 5018 3878 5064 3894
rect 5091 3882 5165 3898
rect 5018 3876 5052 3878
rect 5017 3860 5064 3876
rect 5091 3860 5104 3882
rect 5119 3860 5149 3882
rect 5176 3860 5177 3876
rect 5192 3860 5205 4020
rect 5235 3916 5248 4020
rect 5293 3998 5294 4008
rect 5309 3998 5322 4008
rect 5293 3994 5322 3998
rect 5327 3994 5357 4020
rect 5375 4006 5391 4008
rect 5463 4006 5516 4020
rect 5464 4004 5528 4006
rect 5571 4004 5586 4020
rect 5635 4017 5665 4020
rect 5635 4014 5671 4017
rect 5601 4006 5617 4008
rect 5375 3994 5390 3998
rect 5293 3992 5390 3994
rect 5418 3992 5586 4004
rect 5602 3994 5617 3998
rect 5635 3995 5674 4014
rect 5693 4008 5700 4009
rect 5699 4001 5700 4008
rect 5683 3998 5684 4001
rect 5699 3998 5712 4001
rect 5635 3994 5665 3995
rect 5674 3994 5680 3995
rect 5683 3994 5712 3998
rect 5602 3993 5712 3994
rect 5602 3992 5718 3993
rect 5277 3984 5328 3992
rect 5277 3972 5302 3984
rect 5309 3972 5328 3984
rect 5359 3984 5409 3992
rect 5359 3976 5375 3984
rect 5382 3982 5409 3984
rect 5418 3982 5639 3992
rect 5382 3972 5639 3982
rect 5668 3984 5718 3992
rect 5668 3975 5684 3984
rect 5277 3964 5328 3972
rect 5375 3964 5639 3972
rect 5665 3972 5684 3975
rect 5691 3972 5718 3984
rect 5665 3964 5718 3972
rect 5293 3956 5294 3964
rect 5309 3956 5322 3964
rect 5293 3948 5309 3956
rect 5290 3941 5309 3944
rect 5290 3932 5312 3941
rect 5263 3922 5312 3932
rect 5263 3916 5293 3922
rect 5312 3917 5317 3922
rect 5235 3900 5309 3916
rect 5327 3908 5357 3964
rect 5392 3954 5600 3964
rect 5635 3960 5680 3964
rect 5683 3963 5684 3964
rect 5699 3963 5712 3964
rect 5418 3924 5607 3954
rect 5433 3921 5607 3924
rect 5426 3918 5607 3921
rect 5235 3898 5248 3900
rect 5263 3898 5297 3900
rect 5235 3882 5309 3898
rect 5336 3894 5349 3908
rect 5364 3894 5380 3910
rect 5426 3905 5437 3918
rect 5219 3860 5220 3876
rect 5235 3860 5248 3882
rect 5263 3860 5293 3882
rect 5336 3878 5398 3894
rect 5426 3887 5437 3903
rect 5442 3898 5452 3918
rect 5462 3898 5476 3918
rect 5479 3905 5488 3918
rect 5504 3905 5513 3918
rect 5442 3887 5476 3898
rect 5479 3887 5488 3903
rect 5504 3887 5513 3903
rect 5520 3898 5530 3918
rect 5540 3898 5554 3918
rect 5555 3905 5566 3918
rect 5520 3887 5554 3898
rect 5555 3887 5566 3903
rect 5612 3894 5628 3910
rect 5635 3908 5665 3960
rect 5699 3956 5700 3963
rect 5684 3948 5700 3956
rect 5671 3916 5684 3935
rect 5699 3916 5729 3932
rect 5671 3900 5745 3916
rect 5671 3898 5684 3900
rect 5699 3898 5733 3900
rect 5336 3876 5349 3878
rect 5364 3876 5398 3878
rect 5336 3860 5398 3876
rect 5442 3871 5458 3874
rect 5520 3871 5550 3882
rect 5598 3878 5644 3894
rect 5671 3882 5745 3898
rect 5598 3876 5632 3878
rect 5597 3860 5644 3876
rect 5671 3860 5684 3882
rect 5699 3860 5729 3882
rect 5756 3860 5757 3876
rect 5772 3860 5785 4020
rect 5815 3916 5828 4020
rect 5873 3998 5874 4008
rect 5889 3998 5902 4008
rect 5873 3994 5902 3998
rect 5907 3994 5937 4020
rect 5955 4006 5971 4008
rect 6043 4006 6096 4020
rect 6044 4004 6108 4006
rect 6151 4004 6166 4020
rect 6215 4017 6245 4020
rect 6215 4014 6251 4017
rect 6181 4006 6197 4008
rect 5955 3994 5970 3998
rect 5873 3992 5970 3994
rect 5998 3992 6166 4004
rect 6182 3994 6197 3998
rect 6215 3995 6254 4014
rect 6273 4008 6280 4009
rect 6279 4001 6280 4008
rect 6263 3998 6264 4001
rect 6279 3998 6292 4001
rect 6215 3994 6245 3995
rect 6254 3994 6260 3995
rect 6263 3994 6292 3998
rect 6182 3993 6292 3994
rect 6182 3992 6298 3993
rect 5857 3984 5908 3992
rect 5857 3972 5882 3984
rect 5889 3972 5908 3984
rect 5939 3984 5989 3992
rect 5939 3976 5955 3984
rect 5962 3982 5989 3984
rect 5998 3982 6219 3992
rect 5962 3972 6219 3982
rect 6248 3984 6298 3992
rect 6248 3975 6264 3984
rect 5857 3964 5908 3972
rect 5955 3964 6219 3972
rect 6245 3972 6264 3975
rect 6271 3972 6298 3984
rect 6245 3964 6298 3972
rect 5873 3956 5874 3964
rect 5889 3956 5902 3964
rect 5873 3948 5889 3956
rect 5870 3941 5889 3944
rect 5870 3932 5892 3941
rect 5843 3922 5892 3932
rect 5843 3916 5873 3922
rect 5892 3917 5897 3922
rect 5815 3900 5889 3916
rect 5907 3908 5937 3964
rect 5972 3954 6180 3964
rect 6215 3960 6260 3964
rect 6263 3963 6264 3964
rect 6279 3963 6292 3964
rect 5998 3924 6187 3954
rect 6013 3921 6187 3924
rect 6006 3918 6187 3921
rect 5815 3898 5828 3900
rect 5843 3898 5877 3900
rect 5815 3882 5889 3898
rect 5916 3894 5929 3908
rect 5944 3894 5960 3910
rect 6006 3905 6017 3918
rect 5799 3860 5800 3876
rect 5815 3860 5828 3882
rect 5843 3860 5873 3882
rect 5916 3878 5978 3894
rect 6006 3887 6017 3903
rect 6022 3898 6032 3918
rect 6042 3898 6056 3918
rect 6059 3905 6068 3918
rect 6084 3905 6093 3918
rect 6022 3887 6056 3898
rect 6059 3887 6068 3903
rect 6084 3887 6093 3903
rect 6100 3898 6110 3918
rect 6120 3898 6134 3918
rect 6135 3905 6146 3918
rect 6100 3887 6134 3898
rect 6135 3887 6146 3903
rect 6192 3894 6208 3910
rect 6215 3908 6245 3960
rect 6279 3956 6280 3963
rect 6264 3948 6280 3956
rect 6251 3916 6264 3935
rect 6279 3916 6309 3932
rect 6251 3900 6325 3916
rect 6251 3898 6264 3900
rect 6279 3898 6313 3900
rect 5916 3876 5929 3878
rect 5944 3876 5978 3878
rect 5916 3860 5978 3876
rect 6022 3871 6038 3874
rect 6100 3871 6130 3882
rect 6178 3878 6224 3894
rect 6251 3882 6325 3898
rect 6178 3876 6212 3878
rect 6177 3860 6224 3876
rect 6251 3860 6264 3882
rect 6279 3860 6309 3882
rect 6336 3860 6337 3876
rect 6352 3860 6365 4020
rect 6395 3916 6408 4020
rect 6453 3998 6454 4008
rect 6469 3998 6482 4008
rect 6453 3994 6482 3998
rect 6487 3994 6517 4020
rect 6535 4006 6551 4008
rect 6623 4006 6676 4020
rect 6624 4004 6688 4006
rect 6731 4004 6746 4020
rect 6795 4017 6825 4020
rect 6795 4014 6831 4017
rect 6761 4006 6777 4008
rect 6535 3994 6550 3998
rect 6453 3992 6550 3994
rect 6578 3992 6746 4004
rect 6762 3994 6777 3998
rect 6795 3995 6834 4014
rect 6853 4008 6860 4009
rect 6859 4001 6860 4008
rect 6843 3998 6844 4001
rect 6859 3998 6872 4001
rect 6795 3994 6825 3995
rect 6834 3994 6840 3995
rect 6843 3994 6872 3998
rect 6762 3993 6872 3994
rect 6762 3992 6878 3993
rect 6437 3984 6488 3992
rect 6437 3972 6462 3984
rect 6469 3972 6488 3984
rect 6519 3984 6569 3992
rect 6519 3976 6535 3984
rect 6542 3982 6569 3984
rect 6578 3982 6799 3992
rect 6542 3972 6799 3982
rect 6828 3984 6878 3992
rect 6828 3975 6844 3984
rect 6437 3964 6488 3972
rect 6535 3964 6799 3972
rect 6825 3972 6844 3975
rect 6851 3972 6878 3984
rect 6825 3964 6878 3972
rect 6453 3956 6454 3964
rect 6469 3956 6482 3964
rect 6453 3948 6469 3956
rect 6450 3941 6469 3944
rect 6450 3932 6472 3941
rect 6423 3922 6472 3932
rect 6423 3916 6453 3922
rect 6472 3917 6477 3922
rect 6395 3900 6469 3916
rect 6487 3908 6517 3964
rect 6552 3954 6760 3964
rect 6795 3960 6840 3964
rect 6843 3963 6844 3964
rect 6859 3963 6872 3964
rect 6578 3924 6767 3954
rect 6593 3921 6767 3924
rect 6586 3918 6767 3921
rect 6395 3898 6408 3900
rect 6423 3898 6457 3900
rect 6395 3882 6469 3898
rect 6496 3894 6509 3908
rect 6524 3894 6540 3910
rect 6586 3905 6597 3918
rect 6379 3860 6380 3876
rect 6395 3860 6408 3882
rect 6423 3860 6453 3882
rect 6496 3878 6558 3894
rect 6586 3887 6597 3903
rect 6602 3898 6612 3918
rect 6622 3898 6636 3918
rect 6639 3905 6648 3918
rect 6664 3905 6673 3918
rect 6602 3887 6636 3898
rect 6639 3887 6648 3903
rect 6664 3887 6673 3903
rect 6680 3898 6690 3918
rect 6700 3898 6714 3918
rect 6715 3905 6726 3918
rect 6680 3887 6714 3898
rect 6715 3887 6726 3903
rect 6772 3894 6788 3910
rect 6795 3908 6825 3960
rect 6859 3956 6860 3963
rect 6844 3948 6860 3956
rect 6831 3916 6844 3935
rect 6859 3916 6889 3932
rect 6831 3900 6905 3916
rect 6831 3898 6844 3900
rect 6859 3898 6893 3900
rect 6496 3876 6509 3878
rect 6524 3876 6558 3878
rect 6496 3860 6558 3876
rect 6602 3871 6618 3874
rect 6680 3871 6710 3882
rect 6758 3878 6804 3894
rect 6831 3882 6905 3898
rect 6758 3876 6792 3878
rect 6757 3860 6804 3876
rect 6831 3860 6844 3882
rect 6859 3860 6889 3882
rect 6916 3860 6917 3876
rect 6932 3860 6945 4020
rect 6975 3916 6988 4020
rect 7033 3998 7034 4008
rect 7049 3998 7062 4008
rect 7033 3994 7062 3998
rect 7067 3994 7097 4020
rect 7115 4006 7131 4008
rect 7203 4006 7256 4020
rect 7204 4004 7268 4006
rect 7311 4004 7326 4020
rect 7375 4017 7405 4020
rect 7375 4014 7411 4017
rect 7341 4006 7357 4008
rect 7115 3994 7130 3998
rect 7033 3992 7130 3994
rect 7158 3992 7326 4004
rect 7342 3994 7357 3998
rect 7375 3995 7414 4014
rect 7433 4008 7440 4009
rect 7439 4001 7440 4008
rect 7423 3998 7424 4001
rect 7439 3998 7452 4001
rect 7375 3994 7405 3995
rect 7414 3994 7420 3995
rect 7423 3994 7452 3998
rect 7342 3993 7452 3994
rect 7342 3992 7458 3993
rect 7017 3984 7068 3992
rect 7017 3972 7042 3984
rect 7049 3972 7068 3984
rect 7099 3984 7149 3992
rect 7099 3976 7115 3984
rect 7122 3982 7149 3984
rect 7158 3982 7379 3992
rect 7122 3972 7379 3982
rect 7408 3984 7458 3992
rect 7408 3975 7424 3984
rect 7017 3964 7068 3972
rect 7115 3964 7379 3972
rect 7405 3972 7424 3975
rect 7431 3972 7458 3984
rect 7405 3964 7458 3972
rect 7033 3956 7034 3964
rect 7049 3956 7062 3964
rect 7033 3948 7049 3956
rect 7030 3941 7049 3944
rect 7030 3932 7052 3941
rect 7003 3922 7052 3932
rect 7003 3916 7033 3922
rect 7052 3917 7057 3922
rect 6975 3900 7049 3916
rect 7067 3908 7097 3964
rect 7132 3954 7340 3964
rect 7375 3960 7420 3964
rect 7423 3963 7424 3964
rect 7439 3963 7452 3964
rect 7158 3924 7347 3954
rect 7173 3921 7347 3924
rect 7166 3918 7347 3921
rect 6975 3898 6988 3900
rect 7003 3898 7037 3900
rect 6975 3882 7049 3898
rect 7076 3894 7089 3908
rect 7104 3894 7120 3910
rect 7166 3905 7177 3918
rect 6959 3860 6960 3876
rect 6975 3860 6988 3882
rect 7003 3860 7033 3882
rect 7076 3878 7138 3894
rect 7166 3887 7177 3903
rect 7182 3898 7192 3918
rect 7202 3898 7216 3918
rect 7219 3905 7228 3918
rect 7244 3905 7253 3918
rect 7182 3887 7216 3898
rect 7219 3887 7228 3903
rect 7244 3887 7253 3903
rect 7260 3898 7270 3918
rect 7280 3898 7294 3918
rect 7295 3905 7306 3918
rect 7260 3887 7294 3898
rect 7295 3887 7306 3903
rect 7352 3894 7368 3910
rect 7375 3908 7405 3960
rect 7439 3956 7440 3963
rect 7424 3948 7440 3956
rect 7411 3916 7424 3935
rect 7439 3916 7469 3932
rect 7411 3900 7485 3916
rect 7411 3898 7424 3900
rect 7439 3898 7473 3900
rect 7076 3876 7089 3878
rect 7104 3876 7138 3878
rect 7076 3860 7138 3876
rect 7182 3871 7198 3874
rect 7260 3871 7290 3882
rect 7338 3878 7384 3894
rect 7411 3882 7485 3898
rect 7338 3876 7372 3878
rect 7337 3860 7384 3876
rect 7411 3860 7424 3882
rect 7439 3860 7469 3882
rect 7496 3860 7497 3876
rect 7512 3860 7525 4020
rect 7555 3916 7568 4020
rect 7613 3998 7614 4008
rect 7629 3998 7642 4008
rect 7613 3994 7642 3998
rect 7647 3994 7677 4020
rect 7695 4006 7711 4008
rect 7783 4006 7836 4020
rect 7784 4004 7848 4006
rect 7891 4004 7906 4020
rect 7955 4017 7985 4020
rect 7955 4014 7991 4017
rect 7921 4006 7937 4008
rect 7695 3994 7710 3998
rect 7613 3992 7710 3994
rect 7738 3992 7906 4004
rect 7922 3994 7937 3998
rect 7955 3995 7994 4014
rect 8013 4008 8020 4009
rect 8019 4001 8020 4008
rect 8003 3998 8004 4001
rect 8019 3998 8032 4001
rect 7955 3994 7985 3995
rect 7994 3994 8000 3995
rect 8003 3994 8032 3998
rect 7922 3993 8032 3994
rect 7922 3992 8038 3993
rect 7597 3984 7648 3992
rect 7597 3972 7622 3984
rect 7629 3972 7648 3984
rect 7679 3984 7729 3992
rect 7679 3976 7695 3984
rect 7702 3982 7729 3984
rect 7738 3982 7959 3992
rect 7702 3972 7959 3982
rect 7988 3984 8038 3992
rect 7988 3975 8004 3984
rect 7597 3964 7648 3972
rect 7695 3964 7959 3972
rect 7985 3972 8004 3975
rect 8011 3972 8038 3984
rect 7985 3964 8038 3972
rect 7613 3956 7614 3964
rect 7629 3956 7642 3964
rect 7613 3948 7629 3956
rect 7610 3941 7629 3944
rect 7610 3932 7632 3941
rect 7583 3922 7632 3932
rect 7583 3916 7613 3922
rect 7632 3917 7637 3922
rect 7555 3900 7629 3916
rect 7647 3908 7677 3964
rect 7712 3954 7920 3964
rect 7955 3960 8000 3964
rect 8003 3963 8004 3964
rect 8019 3963 8032 3964
rect 7738 3924 7927 3954
rect 7753 3921 7927 3924
rect 7746 3918 7927 3921
rect 7555 3898 7568 3900
rect 7583 3898 7617 3900
rect 7555 3882 7629 3898
rect 7656 3894 7669 3908
rect 7684 3894 7700 3910
rect 7746 3905 7757 3918
rect 7539 3860 7540 3876
rect 7555 3860 7568 3882
rect 7583 3860 7613 3882
rect 7656 3878 7718 3894
rect 7746 3887 7757 3903
rect 7762 3898 7772 3918
rect 7782 3898 7796 3918
rect 7799 3905 7808 3918
rect 7824 3905 7833 3918
rect 7762 3887 7796 3898
rect 7799 3887 7808 3903
rect 7824 3887 7833 3903
rect 7840 3898 7850 3918
rect 7860 3898 7874 3918
rect 7875 3905 7886 3918
rect 7840 3887 7874 3898
rect 7875 3887 7886 3903
rect 7932 3894 7948 3910
rect 7955 3908 7985 3960
rect 8019 3956 8020 3963
rect 8004 3948 8020 3956
rect 7991 3916 8004 3935
rect 8019 3916 8049 3932
rect 7991 3900 8065 3916
rect 7991 3898 8004 3900
rect 8019 3898 8053 3900
rect 7656 3876 7669 3878
rect 7684 3876 7718 3878
rect 7656 3860 7718 3876
rect 7762 3871 7778 3874
rect 7840 3871 7870 3882
rect 7918 3878 7964 3894
rect 7991 3882 8065 3898
rect 7918 3876 7952 3878
rect 7917 3860 7964 3876
rect 7991 3860 8004 3882
rect 8019 3860 8049 3882
rect 8076 3860 8077 3876
rect 8092 3860 8105 4020
rect 8135 3916 8148 4020
rect 8193 3998 8194 4008
rect 8209 3998 8222 4008
rect 8193 3994 8222 3998
rect 8227 3994 8257 4020
rect 8275 4006 8291 4008
rect 8363 4006 8416 4020
rect 8364 4004 8428 4006
rect 8471 4004 8486 4020
rect 8535 4017 8565 4020
rect 8535 4014 8571 4017
rect 8501 4006 8517 4008
rect 8275 3994 8290 3998
rect 8193 3992 8290 3994
rect 8318 3992 8486 4004
rect 8502 3994 8517 3998
rect 8535 3995 8574 4014
rect 8593 4008 8600 4009
rect 8599 4001 8600 4008
rect 8583 3998 8584 4001
rect 8599 3998 8612 4001
rect 8535 3994 8565 3995
rect 8574 3994 8580 3995
rect 8583 3994 8612 3998
rect 8502 3993 8612 3994
rect 8502 3992 8618 3993
rect 8177 3984 8228 3992
rect 8177 3972 8202 3984
rect 8209 3972 8228 3984
rect 8259 3984 8309 3992
rect 8259 3976 8275 3984
rect 8282 3982 8309 3984
rect 8318 3982 8539 3992
rect 8282 3972 8539 3982
rect 8568 3984 8618 3992
rect 8568 3975 8584 3984
rect 8177 3964 8228 3972
rect 8275 3964 8539 3972
rect 8565 3972 8584 3975
rect 8591 3972 8618 3984
rect 8565 3964 8618 3972
rect 8193 3956 8194 3964
rect 8209 3956 8222 3964
rect 8193 3948 8209 3956
rect 8190 3941 8209 3944
rect 8190 3932 8212 3941
rect 8163 3922 8212 3932
rect 8163 3916 8193 3922
rect 8212 3917 8217 3922
rect 8135 3900 8209 3916
rect 8227 3908 8257 3964
rect 8292 3954 8500 3964
rect 8535 3960 8580 3964
rect 8583 3963 8584 3964
rect 8599 3963 8612 3964
rect 8318 3924 8507 3954
rect 8333 3921 8507 3924
rect 8326 3918 8507 3921
rect 8135 3898 8148 3900
rect 8163 3898 8197 3900
rect 8135 3882 8209 3898
rect 8236 3894 8249 3908
rect 8264 3894 8280 3910
rect 8326 3905 8337 3918
rect 8119 3860 8120 3876
rect 8135 3860 8148 3882
rect 8163 3860 8193 3882
rect 8236 3878 8298 3894
rect 8326 3887 8337 3903
rect 8342 3898 8352 3918
rect 8362 3898 8376 3918
rect 8379 3905 8388 3918
rect 8404 3905 8413 3918
rect 8342 3887 8376 3898
rect 8379 3887 8388 3903
rect 8404 3887 8413 3903
rect 8420 3898 8430 3918
rect 8440 3898 8454 3918
rect 8455 3905 8466 3918
rect 8420 3887 8454 3898
rect 8455 3887 8466 3903
rect 8512 3894 8528 3910
rect 8535 3908 8565 3960
rect 8599 3956 8600 3963
rect 8584 3948 8600 3956
rect 8571 3916 8584 3935
rect 8599 3916 8629 3932
rect 8571 3900 8645 3916
rect 8571 3898 8584 3900
rect 8599 3898 8633 3900
rect 8236 3876 8249 3878
rect 8264 3876 8298 3878
rect 8236 3860 8298 3876
rect 8342 3871 8358 3874
rect 8420 3871 8450 3882
rect 8498 3878 8544 3894
rect 8571 3882 8645 3898
rect 8498 3876 8532 3878
rect 8497 3860 8544 3876
rect 8571 3860 8584 3882
rect 8599 3860 8629 3882
rect 8656 3860 8657 3876
rect 8672 3860 8685 4020
rect 8715 3916 8728 4020
rect 8773 3998 8774 4008
rect 8789 3998 8802 4008
rect 8773 3994 8802 3998
rect 8807 3994 8837 4020
rect 8855 4006 8871 4008
rect 8943 4006 8996 4020
rect 8944 4004 9008 4006
rect 9051 4004 9066 4020
rect 9115 4017 9145 4020
rect 9115 4014 9151 4017
rect 9081 4006 9097 4008
rect 8855 3994 8870 3998
rect 8773 3992 8870 3994
rect 8898 3992 9066 4004
rect 9082 3994 9097 3998
rect 9115 3995 9154 4014
rect 9173 4008 9180 4009
rect 9179 4001 9180 4008
rect 9163 3998 9164 4001
rect 9179 3998 9192 4001
rect 9115 3994 9145 3995
rect 9154 3994 9160 3995
rect 9163 3994 9192 3998
rect 9082 3993 9192 3994
rect 9082 3992 9198 3993
rect 8757 3984 8808 3992
rect 8757 3972 8782 3984
rect 8789 3972 8808 3984
rect 8839 3984 8889 3992
rect 8839 3976 8855 3984
rect 8862 3982 8889 3984
rect 8898 3982 9119 3992
rect 8862 3972 9119 3982
rect 9148 3984 9198 3992
rect 9148 3975 9164 3984
rect 8757 3964 8808 3972
rect 8855 3964 9119 3972
rect 9145 3972 9164 3975
rect 9171 3972 9198 3984
rect 9145 3964 9198 3972
rect 8773 3956 8774 3964
rect 8789 3956 8802 3964
rect 8773 3948 8789 3956
rect 8770 3941 8789 3944
rect 8770 3932 8792 3941
rect 8743 3922 8792 3932
rect 8743 3916 8773 3922
rect 8792 3917 8797 3922
rect 8715 3900 8789 3916
rect 8807 3908 8837 3964
rect 8872 3954 9080 3964
rect 9115 3960 9160 3964
rect 9163 3963 9164 3964
rect 9179 3963 9192 3964
rect 8898 3924 9087 3954
rect 8913 3921 9087 3924
rect 8906 3918 9087 3921
rect 8715 3898 8728 3900
rect 8743 3898 8777 3900
rect 8715 3882 8789 3898
rect 8816 3894 8829 3908
rect 8844 3894 8860 3910
rect 8906 3905 8917 3918
rect 8699 3860 8700 3876
rect 8715 3860 8728 3882
rect 8743 3860 8773 3882
rect 8816 3878 8878 3894
rect 8906 3887 8917 3903
rect 8922 3898 8932 3918
rect 8942 3898 8956 3918
rect 8959 3905 8968 3918
rect 8984 3905 8993 3918
rect 8922 3887 8956 3898
rect 8959 3887 8968 3903
rect 8984 3887 8993 3903
rect 9000 3898 9010 3918
rect 9020 3898 9034 3918
rect 9035 3905 9046 3918
rect 9000 3887 9034 3898
rect 9035 3887 9046 3903
rect 9092 3894 9108 3910
rect 9115 3908 9145 3960
rect 9179 3956 9180 3963
rect 9164 3948 9180 3956
rect 9151 3916 9164 3935
rect 9179 3916 9209 3932
rect 9151 3900 9225 3916
rect 9151 3898 9164 3900
rect 9179 3898 9213 3900
rect 8816 3876 8829 3878
rect 8844 3876 8878 3878
rect 8816 3860 8878 3876
rect 8922 3871 8938 3874
rect 9000 3871 9030 3882
rect 9078 3878 9124 3894
rect 9151 3882 9225 3898
rect 9078 3876 9112 3878
rect 9077 3860 9124 3876
rect 9151 3860 9164 3882
rect 9179 3860 9209 3882
rect 9236 3860 9237 3876
rect 9252 3860 9265 4020
rect -7 3852 34 3860
rect -7 3826 8 3852
rect 15 3826 34 3852
rect 98 3848 160 3860
rect 172 3848 247 3860
rect 305 3848 380 3860
rect 392 3848 423 3860
rect 429 3848 464 3860
rect 98 3846 260 3848
rect -7 3818 34 3826
rect 116 3822 129 3846
rect 144 3844 159 3846
rect -1 3808 0 3818
rect 15 3808 28 3818
rect 43 3808 73 3822
rect 116 3808 159 3822
rect 183 3819 190 3826
rect 193 3822 260 3846
rect 292 3846 464 3848
rect 262 3824 290 3828
rect 292 3824 372 3846
rect 393 3844 408 3846
rect 262 3822 372 3824
rect 193 3818 372 3822
rect 166 3808 196 3818
rect 198 3808 351 3818
rect 359 3808 389 3818
rect 393 3808 423 3822
rect 451 3808 464 3846
rect 536 3852 571 3860
rect 536 3826 537 3852
rect 544 3826 571 3852
rect 479 3808 509 3822
rect 536 3818 571 3826
rect 573 3852 614 3860
rect 573 3826 588 3852
rect 595 3826 614 3852
rect 678 3848 740 3860
rect 752 3848 827 3860
rect 885 3848 960 3860
rect 972 3848 1003 3860
rect 1009 3848 1044 3860
rect 678 3846 840 3848
rect 573 3818 614 3826
rect 696 3822 709 3846
rect 724 3844 739 3846
rect 536 3808 537 3818
rect 552 3808 565 3818
rect 579 3808 580 3818
rect 595 3808 608 3818
rect 623 3808 653 3822
rect 696 3808 739 3822
rect 763 3819 770 3826
rect 773 3822 840 3846
rect 872 3846 1044 3848
rect 842 3824 870 3828
rect 872 3824 952 3846
rect 973 3844 988 3846
rect 842 3822 952 3824
rect 773 3818 952 3822
rect 746 3808 776 3818
rect 778 3808 931 3818
rect 939 3808 969 3818
rect 973 3808 1003 3822
rect 1031 3808 1044 3846
rect 1116 3852 1151 3860
rect 1116 3826 1117 3852
rect 1124 3826 1151 3852
rect 1059 3808 1089 3822
rect 1116 3818 1151 3826
rect 1153 3852 1194 3860
rect 1153 3826 1168 3852
rect 1175 3826 1194 3852
rect 1258 3848 1320 3860
rect 1332 3848 1407 3860
rect 1465 3848 1540 3860
rect 1552 3848 1583 3860
rect 1589 3848 1624 3860
rect 1258 3846 1420 3848
rect 1153 3818 1194 3826
rect 1276 3822 1289 3846
rect 1304 3844 1319 3846
rect 1116 3808 1117 3818
rect 1132 3808 1145 3818
rect 1159 3808 1160 3818
rect 1175 3808 1188 3818
rect 1203 3808 1233 3822
rect 1276 3808 1319 3822
rect 1343 3819 1350 3826
rect 1353 3822 1420 3846
rect 1452 3846 1624 3848
rect 1422 3824 1450 3828
rect 1452 3824 1532 3846
rect 1553 3844 1568 3846
rect 1422 3822 1532 3824
rect 1353 3818 1532 3822
rect 1326 3808 1356 3818
rect 1358 3808 1511 3818
rect 1519 3808 1549 3818
rect 1553 3808 1583 3822
rect 1611 3808 1624 3846
rect 1696 3852 1731 3860
rect 1696 3826 1697 3852
rect 1704 3826 1731 3852
rect 1639 3808 1669 3822
rect 1696 3818 1731 3826
rect 1733 3852 1774 3860
rect 1733 3826 1748 3852
rect 1755 3826 1774 3852
rect 1838 3848 1900 3860
rect 1912 3848 1987 3860
rect 2045 3848 2120 3860
rect 2132 3848 2163 3860
rect 2169 3848 2204 3860
rect 1838 3846 2000 3848
rect 1733 3818 1774 3826
rect 1856 3822 1869 3846
rect 1884 3844 1899 3846
rect 1696 3808 1697 3818
rect 1712 3808 1725 3818
rect 1739 3808 1740 3818
rect 1755 3808 1768 3818
rect 1783 3808 1813 3822
rect 1856 3808 1899 3822
rect 1923 3819 1930 3826
rect 1933 3822 2000 3846
rect 2032 3846 2204 3848
rect 2002 3824 2030 3828
rect 2032 3824 2112 3846
rect 2133 3844 2148 3846
rect 2002 3822 2112 3824
rect 1933 3818 2112 3822
rect 1906 3808 1936 3818
rect 1938 3808 2091 3818
rect 2099 3808 2129 3818
rect 2133 3808 2163 3822
rect 2191 3808 2204 3846
rect 2276 3852 2311 3860
rect 2276 3826 2277 3852
rect 2284 3826 2311 3852
rect 2219 3808 2249 3822
rect 2276 3818 2311 3826
rect 2313 3852 2354 3860
rect 2313 3826 2328 3852
rect 2335 3826 2354 3852
rect 2418 3848 2480 3860
rect 2492 3848 2567 3860
rect 2625 3848 2700 3860
rect 2712 3848 2743 3860
rect 2749 3848 2784 3860
rect 2418 3846 2580 3848
rect 2313 3818 2354 3826
rect 2436 3822 2449 3846
rect 2464 3844 2479 3846
rect 2276 3808 2277 3818
rect 2292 3808 2305 3818
rect 2319 3808 2320 3818
rect 2335 3808 2348 3818
rect 2363 3808 2393 3822
rect 2436 3808 2479 3822
rect 2503 3819 2510 3826
rect 2513 3822 2580 3846
rect 2612 3846 2784 3848
rect 2582 3824 2610 3828
rect 2612 3824 2692 3846
rect 2713 3844 2728 3846
rect 2582 3822 2692 3824
rect 2513 3818 2692 3822
rect 2486 3808 2516 3818
rect 2518 3808 2671 3818
rect 2679 3808 2709 3818
rect 2713 3808 2743 3822
rect 2771 3808 2784 3846
rect 2856 3852 2891 3860
rect 2856 3826 2857 3852
rect 2864 3826 2891 3852
rect 2799 3808 2829 3822
rect 2856 3818 2891 3826
rect 2893 3852 2934 3860
rect 2893 3826 2908 3852
rect 2915 3826 2934 3852
rect 2998 3848 3060 3860
rect 3072 3848 3147 3860
rect 3205 3848 3280 3860
rect 3292 3848 3323 3860
rect 3329 3848 3364 3860
rect 2998 3846 3160 3848
rect 2893 3818 2934 3826
rect 3016 3822 3029 3846
rect 3044 3844 3059 3846
rect 2856 3808 2857 3818
rect 2872 3808 2885 3818
rect 2899 3808 2900 3818
rect 2915 3808 2928 3818
rect 2943 3808 2973 3822
rect 3016 3808 3059 3822
rect 3083 3819 3090 3826
rect 3093 3822 3160 3846
rect 3192 3846 3364 3848
rect 3162 3824 3190 3828
rect 3192 3824 3272 3846
rect 3293 3844 3308 3846
rect 3162 3822 3272 3824
rect 3093 3818 3272 3822
rect 3066 3808 3096 3818
rect 3098 3808 3251 3818
rect 3259 3808 3289 3818
rect 3293 3808 3323 3822
rect 3351 3808 3364 3846
rect 3436 3852 3471 3860
rect 3436 3826 3437 3852
rect 3444 3826 3471 3852
rect 3379 3808 3409 3822
rect 3436 3818 3471 3826
rect 3473 3852 3514 3860
rect 3473 3826 3488 3852
rect 3495 3826 3514 3852
rect 3578 3848 3640 3860
rect 3652 3848 3727 3860
rect 3785 3848 3860 3860
rect 3872 3848 3903 3860
rect 3909 3848 3944 3860
rect 3578 3846 3740 3848
rect 3473 3818 3514 3826
rect 3596 3822 3609 3846
rect 3624 3844 3639 3846
rect 3436 3808 3437 3818
rect 3452 3808 3465 3818
rect 3479 3808 3480 3818
rect 3495 3808 3508 3818
rect 3523 3808 3553 3822
rect 3596 3808 3639 3822
rect 3663 3819 3670 3826
rect 3673 3822 3740 3846
rect 3772 3846 3944 3848
rect 3742 3824 3770 3828
rect 3772 3824 3852 3846
rect 3873 3844 3888 3846
rect 3742 3822 3852 3824
rect 3673 3818 3852 3822
rect 3646 3808 3676 3818
rect 3678 3808 3831 3818
rect 3839 3808 3869 3818
rect 3873 3808 3903 3822
rect 3931 3808 3944 3846
rect 4016 3852 4051 3860
rect 4016 3826 4017 3852
rect 4024 3826 4051 3852
rect 3959 3808 3989 3822
rect 4016 3818 4051 3826
rect 4053 3852 4094 3860
rect 4053 3826 4068 3852
rect 4075 3826 4094 3852
rect 4158 3848 4220 3860
rect 4232 3848 4307 3860
rect 4365 3848 4440 3860
rect 4452 3848 4483 3860
rect 4489 3848 4524 3860
rect 4158 3846 4320 3848
rect 4053 3818 4094 3826
rect 4176 3822 4189 3846
rect 4204 3844 4219 3846
rect 4016 3808 4017 3818
rect 4032 3808 4045 3818
rect 4059 3808 4060 3818
rect 4075 3808 4088 3818
rect 4103 3808 4133 3822
rect 4176 3808 4219 3822
rect 4243 3819 4250 3826
rect 4253 3822 4320 3846
rect 4352 3846 4524 3848
rect 4322 3824 4350 3828
rect 4352 3824 4432 3846
rect 4453 3844 4468 3846
rect 4322 3822 4432 3824
rect 4253 3818 4432 3822
rect 4226 3808 4256 3818
rect 4258 3808 4411 3818
rect 4419 3808 4449 3818
rect 4453 3808 4483 3822
rect 4511 3808 4524 3846
rect 4596 3852 4631 3860
rect 4596 3826 4597 3852
rect 4604 3826 4631 3852
rect 4539 3808 4569 3822
rect 4596 3818 4631 3826
rect 4633 3852 4674 3860
rect 4633 3826 4648 3852
rect 4655 3826 4674 3852
rect 4738 3848 4800 3860
rect 4812 3848 4887 3860
rect 4945 3848 5020 3860
rect 5032 3848 5063 3860
rect 5069 3848 5104 3860
rect 4738 3846 4900 3848
rect 4633 3818 4674 3826
rect 4756 3822 4769 3846
rect 4784 3844 4799 3846
rect 4596 3808 4597 3818
rect 4612 3808 4625 3818
rect 4639 3808 4640 3818
rect 4655 3808 4668 3818
rect 4683 3808 4713 3822
rect 4756 3808 4799 3822
rect 4823 3819 4830 3826
rect 4833 3822 4900 3846
rect 4932 3846 5104 3848
rect 4902 3824 4930 3828
rect 4932 3824 5012 3846
rect 5033 3844 5048 3846
rect 4902 3822 5012 3824
rect 4833 3818 5012 3822
rect 4806 3808 4836 3818
rect 4838 3808 4991 3818
rect 4999 3808 5029 3818
rect 5033 3808 5063 3822
rect 5091 3808 5104 3846
rect 5176 3852 5211 3860
rect 5176 3826 5177 3852
rect 5184 3826 5211 3852
rect 5119 3808 5149 3822
rect 5176 3818 5211 3826
rect 5213 3852 5254 3860
rect 5213 3826 5228 3852
rect 5235 3826 5254 3852
rect 5318 3848 5380 3860
rect 5392 3848 5467 3860
rect 5525 3848 5600 3860
rect 5612 3848 5643 3860
rect 5649 3848 5684 3860
rect 5318 3846 5480 3848
rect 5213 3818 5254 3826
rect 5336 3822 5349 3846
rect 5364 3844 5379 3846
rect 5176 3808 5177 3818
rect 5192 3808 5205 3818
rect 5219 3808 5220 3818
rect 5235 3808 5248 3818
rect 5263 3808 5293 3822
rect 5336 3808 5379 3822
rect 5403 3819 5410 3826
rect 5413 3822 5480 3846
rect 5512 3846 5684 3848
rect 5482 3824 5510 3828
rect 5512 3824 5592 3846
rect 5613 3844 5628 3846
rect 5482 3822 5592 3824
rect 5413 3818 5592 3822
rect 5386 3808 5416 3818
rect 5418 3808 5571 3818
rect 5579 3808 5609 3818
rect 5613 3808 5643 3822
rect 5671 3808 5684 3846
rect 5756 3852 5791 3860
rect 5756 3826 5757 3852
rect 5764 3826 5791 3852
rect 5699 3808 5729 3822
rect 5756 3818 5791 3826
rect 5793 3852 5834 3860
rect 5793 3826 5808 3852
rect 5815 3826 5834 3852
rect 5898 3848 5960 3860
rect 5972 3848 6047 3860
rect 6105 3848 6180 3860
rect 6192 3848 6223 3860
rect 6229 3848 6264 3860
rect 5898 3846 6060 3848
rect 5793 3818 5834 3826
rect 5916 3822 5929 3846
rect 5944 3844 5959 3846
rect 5756 3808 5757 3818
rect 5772 3808 5785 3818
rect 5799 3808 5800 3818
rect 5815 3808 5828 3818
rect 5843 3808 5873 3822
rect 5916 3808 5959 3822
rect 5983 3819 5990 3826
rect 5993 3822 6060 3846
rect 6092 3846 6264 3848
rect 6062 3824 6090 3828
rect 6092 3824 6172 3846
rect 6193 3844 6208 3846
rect 6062 3822 6172 3824
rect 5993 3818 6172 3822
rect 5966 3808 5996 3818
rect 5998 3808 6151 3818
rect 6159 3808 6189 3818
rect 6193 3808 6223 3822
rect 6251 3808 6264 3846
rect 6336 3852 6371 3860
rect 6336 3826 6337 3852
rect 6344 3826 6371 3852
rect 6279 3808 6309 3822
rect 6336 3818 6371 3826
rect 6373 3852 6414 3860
rect 6373 3826 6388 3852
rect 6395 3826 6414 3852
rect 6478 3848 6540 3860
rect 6552 3848 6627 3860
rect 6685 3848 6760 3860
rect 6772 3848 6803 3860
rect 6809 3848 6844 3860
rect 6478 3846 6640 3848
rect 6373 3818 6414 3826
rect 6496 3822 6509 3846
rect 6524 3844 6539 3846
rect 6336 3808 6337 3818
rect 6352 3808 6365 3818
rect 6379 3808 6380 3818
rect 6395 3808 6408 3818
rect 6423 3808 6453 3822
rect 6496 3808 6539 3822
rect 6563 3819 6570 3826
rect 6573 3822 6640 3846
rect 6672 3846 6844 3848
rect 6642 3824 6670 3828
rect 6672 3824 6752 3846
rect 6773 3844 6788 3846
rect 6642 3822 6752 3824
rect 6573 3818 6752 3822
rect 6546 3808 6576 3818
rect 6578 3808 6731 3818
rect 6739 3808 6769 3818
rect 6773 3808 6803 3822
rect 6831 3808 6844 3846
rect 6916 3852 6951 3860
rect 6916 3826 6917 3852
rect 6924 3826 6951 3852
rect 6859 3808 6889 3822
rect 6916 3818 6951 3826
rect 6953 3852 6994 3860
rect 6953 3826 6968 3852
rect 6975 3826 6994 3852
rect 7058 3848 7120 3860
rect 7132 3848 7207 3860
rect 7265 3848 7340 3860
rect 7352 3848 7383 3860
rect 7389 3848 7424 3860
rect 7058 3846 7220 3848
rect 6953 3818 6994 3826
rect 7076 3822 7089 3846
rect 7104 3844 7119 3846
rect 6916 3808 6917 3818
rect 6932 3808 6945 3818
rect 6959 3808 6960 3818
rect 6975 3808 6988 3818
rect 7003 3808 7033 3822
rect 7076 3808 7119 3822
rect 7143 3819 7150 3826
rect 7153 3822 7220 3846
rect 7252 3846 7424 3848
rect 7222 3824 7250 3828
rect 7252 3824 7332 3846
rect 7353 3844 7368 3846
rect 7222 3822 7332 3824
rect 7153 3818 7332 3822
rect 7126 3808 7156 3818
rect 7158 3808 7311 3818
rect 7319 3808 7349 3818
rect 7353 3808 7383 3822
rect 7411 3808 7424 3846
rect 7496 3852 7531 3860
rect 7496 3826 7497 3852
rect 7504 3826 7531 3852
rect 7439 3808 7469 3822
rect 7496 3818 7531 3826
rect 7533 3852 7574 3860
rect 7533 3826 7548 3852
rect 7555 3826 7574 3852
rect 7638 3848 7700 3860
rect 7712 3848 7787 3860
rect 7845 3848 7920 3860
rect 7932 3848 7963 3860
rect 7969 3848 8004 3860
rect 7638 3846 7800 3848
rect 7533 3818 7574 3826
rect 7656 3822 7669 3846
rect 7684 3844 7699 3846
rect 7496 3808 7497 3818
rect 7512 3808 7525 3818
rect 7539 3808 7540 3818
rect 7555 3808 7568 3818
rect 7583 3808 7613 3822
rect 7656 3808 7699 3822
rect 7723 3819 7730 3826
rect 7733 3822 7800 3846
rect 7832 3846 8004 3848
rect 7802 3824 7830 3828
rect 7832 3824 7912 3846
rect 7933 3844 7948 3846
rect 7802 3822 7912 3824
rect 7733 3818 7912 3822
rect 7706 3808 7736 3818
rect 7738 3808 7891 3818
rect 7899 3808 7929 3818
rect 7933 3808 7963 3822
rect 7991 3808 8004 3846
rect 8076 3852 8111 3860
rect 8076 3826 8077 3852
rect 8084 3826 8111 3852
rect 8019 3808 8049 3822
rect 8076 3818 8111 3826
rect 8113 3852 8154 3860
rect 8113 3826 8128 3852
rect 8135 3826 8154 3852
rect 8218 3848 8280 3860
rect 8292 3848 8367 3860
rect 8425 3848 8500 3860
rect 8512 3848 8543 3860
rect 8549 3848 8584 3860
rect 8218 3846 8380 3848
rect 8113 3818 8154 3826
rect 8236 3822 8249 3846
rect 8264 3844 8279 3846
rect 8076 3808 8077 3818
rect 8092 3808 8105 3818
rect 8119 3808 8120 3818
rect 8135 3808 8148 3818
rect 8163 3808 8193 3822
rect 8236 3808 8279 3822
rect 8303 3819 8310 3826
rect 8313 3822 8380 3846
rect 8412 3846 8584 3848
rect 8382 3824 8410 3828
rect 8412 3824 8492 3846
rect 8513 3844 8528 3846
rect 8382 3822 8492 3824
rect 8313 3818 8492 3822
rect 8286 3808 8316 3818
rect 8318 3808 8471 3818
rect 8479 3808 8509 3818
rect 8513 3808 8543 3822
rect 8571 3808 8584 3846
rect 8656 3852 8691 3860
rect 8656 3826 8657 3852
rect 8664 3826 8691 3852
rect 8599 3808 8629 3822
rect 8656 3818 8691 3826
rect 8693 3852 8734 3860
rect 8693 3826 8708 3852
rect 8715 3826 8734 3852
rect 8798 3848 8860 3860
rect 8872 3848 8947 3860
rect 9005 3848 9080 3860
rect 9092 3848 9123 3860
rect 9129 3848 9164 3860
rect 8798 3846 8960 3848
rect 8693 3818 8734 3826
rect 8816 3822 8829 3846
rect 8844 3844 8859 3846
rect 8656 3808 8657 3818
rect 8672 3808 8685 3818
rect 8699 3808 8700 3818
rect 8715 3808 8728 3818
rect 8743 3808 8773 3822
rect 8816 3808 8859 3822
rect 8883 3819 8890 3826
rect 8893 3822 8960 3846
rect 8992 3846 9164 3848
rect 8962 3824 8990 3828
rect 8992 3824 9072 3846
rect 9093 3844 9108 3846
rect 8962 3822 9072 3824
rect 8893 3818 9072 3822
rect 8866 3808 8896 3818
rect 8898 3808 9051 3818
rect 9059 3808 9089 3818
rect 9093 3808 9123 3822
rect 9151 3808 9164 3846
rect 9236 3852 9271 3860
rect 9236 3826 9237 3852
rect 9244 3826 9271 3852
rect 9179 3808 9209 3822
rect 9236 3818 9271 3826
rect 9236 3808 9237 3818
rect 9252 3808 9265 3818
rect -1 3802 9265 3808
rect 0 3794 9265 3802
rect 15 3764 28 3794
rect 43 3776 73 3794
rect 116 3780 130 3794
rect 166 3780 386 3794
rect 117 3778 130 3780
rect 83 3766 98 3778
rect 80 3764 102 3766
rect 107 3764 137 3778
rect 198 3776 351 3780
rect 180 3764 372 3776
rect 415 3764 445 3778
rect 451 3764 464 3794
rect 479 3776 509 3794
rect 552 3764 565 3794
rect 595 3764 608 3794
rect 623 3776 653 3794
rect 696 3780 710 3794
rect 746 3780 966 3794
rect 697 3778 710 3780
rect 663 3766 678 3778
rect 660 3764 682 3766
rect 687 3764 717 3778
rect 778 3776 931 3780
rect 760 3764 952 3776
rect 995 3764 1025 3778
rect 1031 3764 1044 3794
rect 1059 3776 1089 3794
rect 1132 3764 1145 3794
rect 1175 3764 1188 3794
rect 1203 3776 1233 3794
rect 1276 3780 1290 3794
rect 1326 3780 1546 3794
rect 1277 3778 1290 3780
rect 1243 3766 1258 3778
rect 1240 3764 1262 3766
rect 1267 3764 1297 3778
rect 1358 3776 1511 3780
rect 1340 3764 1532 3776
rect 1575 3764 1605 3778
rect 1611 3764 1624 3794
rect 1639 3776 1669 3794
rect 1712 3764 1725 3794
rect 1755 3764 1768 3794
rect 1783 3776 1813 3794
rect 1856 3780 1870 3794
rect 1906 3780 2126 3794
rect 1857 3778 1870 3780
rect 1823 3766 1838 3778
rect 1820 3764 1842 3766
rect 1847 3764 1877 3778
rect 1938 3776 2091 3780
rect 1920 3764 2112 3776
rect 2155 3764 2185 3778
rect 2191 3764 2204 3794
rect 2219 3776 2249 3794
rect 2292 3764 2305 3794
rect 2335 3764 2348 3794
rect 2363 3776 2393 3794
rect 2436 3780 2450 3794
rect 2486 3780 2706 3794
rect 2437 3778 2450 3780
rect 2403 3766 2418 3778
rect 2400 3764 2422 3766
rect 2427 3764 2457 3778
rect 2518 3776 2671 3780
rect 2500 3764 2692 3776
rect 2735 3764 2765 3778
rect 2771 3764 2784 3794
rect 2799 3776 2829 3794
rect 2872 3764 2885 3794
rect 2915 3764 2928 3794
rect 2943 3776 2973 3794
rect 3016 3780 3030 3794
rect 3066 3780 3286 3794
rect 3017 3778 3030 3780
rect 2983 3766 2998 3778
rect 2980 3764 3002 3766
rect 3007 3764 3037 3778
rect 3098 3776 3251 3780
rect 3080 3764 3272 3776
rect 3315 3764 3345 3778
rect 3351 3764 3364 3794
rect 3379 3776 3409 3794
rect 3452 3764 3465 3794
rect 3495 3764 3508 3794
rect 3523 3776 3553 3794
rect 3596 3780 3610 3794
rect 3646 3780 3866 3794
rect 3597 3778 3610 3780
rect 3563 3766 3578 3778
rect 3560 3764 3582 3766
rect 3587 3764 3617 3778
rect 3678 3776 3831 3780
rect 3660 3764 3852 3776
rect 3895 3764 3925 3778
rect 3931 3764 3944 3794
rect 3959 3776 3989 3794
rect 4032 3764 4045 3794
rect 4075 3764 4088 3794
rect 4103 3776 4133 3794
rect 4176 3780 4190 3794
rect 4226 3780 4446 3794
rect 4177 3778 4190 3780
rect 4143 3766 4158 3778
rect 4140 3764 4162 3766
rect 4167 3764 4197 3778
rect 4258 3776 4411 3780
rect 4240 3764 4432 3776
rect 4475 3764 4505 3778
rect 4511 3764 4524 3794
rect 4539 3776 4569 3794
rect 4612 3764 4625 3794
rect 4655 3764 4668 3794
rect 4683 3776 4713 3794
rect 4756 3780 4770 3794
rect 4806 3780 5026 3794
rect 4757 3778 4770 3780
rect 4723 3766 4738 3778
rect 4720 3764 4742 3766
rect 4747 3764 4777 3778
rect 4838 3776 4991 3780
rect 4820 3764 5012 3776
rect 5055 3764 5085 3778
rect 5091 3764 5104 3794
rect 5119 3776 5149 3794
rect 5192 3764 5205 3794
rect 5235 3764 5248 3794
rect 5263 3776 5293 3794
rect 5336 3780 5350 3794
rect 5386 3780 5606 3794
rect 5337 3778 5350 3780
rect 5303 3766 5318 3778
rect 5300 3764 5322 3766
rect 5327 3764 5357 3778
rect 5418 3776 5571 3780
rect 5400 3764 5592 3776
rect 5635 3764 5665 3778
rect 5671 3764 5684 3794
rect 5699 3776 5729 3794
rect 5772 3764 5785 3794
rect 5815 3764 5828 3794
rect 5843 3776 5873 3794
rect 5916 3780 5930 3794
rect 5966 3780 6186 3794
rect 5917 3778 5930 3780
rect 5883 3766 5898 3778
rect 5880 3764 5902 3766
rect 5907 3764 5937 3778
rect 5998 3776 6151 3780
rect 5980 3764 6172 3776
rect 6215 3764 6245 3778
rect 6251 3764 6264 3794
rect 6279 3776 6309 3794
rect 6352 3764 6365 3794
rect 6395 3764 6408 3794
rect 6423 3776 6453 3794
rect 6496 3780 6510 3794
rect 6546 3780 6766 3794
rect 6497 3778 6510 3780
rect 6463 3766 6478 3778
rect 6460 3764 6482 3766
rect 6487 3764 6517 3778
rect 6578 3776 6731 3780
rect 6560 3764 6752 3776
rect 6795 3764 6825 3778
rect 6831 3764 6844 3794
rect 6859 3776 6889 3794
rect 6932 3764 6945 3794
rect 6975 3764 6988 3794
rect 7003 3776 7033 3794
rect 7076 3780 7090 3794
rect 7126 3780 7346 3794
rect 7077 3778 7090 3780
rect 7043 3766 7058 3778
rect 7040 3764 7062 3766
rect 7067 3764 7097 3778
rect 7158 3776 7311 3780
rect 7140 3764 7332 3776
rect 7375 3764 7405 3778
rect 7411 3764 7424 3794
rect 7439 3776 7469 3794
rect 7512 3764 7525 3794
rect 7555 3764 7568 3794
rect 7583 3776 7613 3794
rect 7656 3780 7670 3794
rect 7706 3780 7926 3794
rect 7657 3778 7670 3780
rect 7623 3766 7638 3778
rect 7620 3764 7642 3766
rect 7647 3764 7677 3778
rect 7738 3776 7891 3780
rect 7720 3764 7912 3776
rect 7955 3764 7985 3778
rect 7991 3764 8004 3794
rect 8019 3776 8049 3794
rect 8092 3764 8105 3794
rect 8135 3764 8148 3794
rect 8163 3776 8193 3794
rect 8236 3780 8250 3794
rect 8286 3780 8506 3794
rect 8237 3778 8250 3780
rect 8203 3766 8218 3778
rect 8200 3764 8222 3766
rect 8227 3764 8257 3778
rect 8318 3776 8471 3780
rect 8300 3764 8492 3776
rect 8535 3764 8565 3778
rect 8571 3764 8584 3794
rect 8599 3776 8629 3794
rect 8672 3764 8685 3794
rect 8715 3764 8728 3794
rect 8743 3776 8773 3794
rect 8816 3780 8830 3794
rect 8866 3780 9086 3794
rect 8817 3778 8830 3780
rect 8783 3766 8798 3778
rect 8780 3764 8802 3766
rect 8807 3764 8837 3778
rect 8898 3776 9051 3780
rect 8880 3764 9072 3776
rect 9115 3764 9145 3778
rect 9151 3764 9164 3794
rect 9179 3776 9209 3794
rect 9252 3764 9265 3794
rect 0 3750 9265 3764
rect 15 3646 28 3750
rect 73 3728 74 3738
rect 89 3728 102 3738
rect 73 3724 102 3728
rect 107 3724 137 3750
rect 155 3736 171 3738
rect 243 3736 296 3750
rect 244 3734 308 3736
rect 351 3734 366 3750
rect 415 3747 445 3750
rect 415 3744 451 3747
rect 381 3736 397 3738
rect 155 3724 170 3728
rect 73 3722 170 3724
rect 198 3722 366 3734
rect 382 3724 397 3728
rect 415 3725 454 3744
rect 473 3738 480 3739
rect 479 3731 480 3738
rect 463 3728 464 3731
rect 479 3728 492 3731
rect 415 3724 445 3725
rect 454 3724 460 3725
rect 463 3724 492 3728
rect 382 3723 492 3724
rect 382 3722 498 3723
rect 57 3714 108 3722
rect 57 3702 82 3714
rect 89 3702 108 3714
rect 139 3714 189 3722
rect 139 3706 155 3714
rect 162 3712 189 3714
rect 198 3712 419 3722
rect 162 3702 419 3712
rect 448 3714 498 3722
rect 448 3705 464 3714
rect 57 3694 108 3702
rect 155 3694 419 3702
rect 445 3702 464 3705
rect 471 3702 498 3714
rect 445 3694 498 3702
rect 73 3686 74 3694
rect 89 3686 102 3694
rect 73 3678 89 3686
rect 70 3671 89 3674
rect 70 3662 92 3671
rect 43 3652 92 3662
rect 43 3646 73 3652
rect 92 3647 97 3652
rect 15 3630 89 3646
rect 107 3638 137 3694
rect 172 3684 380 3694
rect 415 3690 460 3694
rect 463 3693 464 3694
rect 479 3693 492 3694
rect 198 3654 387 3684
rect 213 3651 387 3654
rect 206 3648 387 3651
rect 15 3628 28 3630
rect 43 3628 77 3630
rect 15 3612 89 3628
rect 116 3624 129 3638
rect 144 3624 160 3640
rect 206 3635 217 3648
rect -1 3590 0 3606
rect 15 3590 28 3612
rect 43 3590 73 3612
rect 116 3608 178 3624
rect 206 3617 217 3633
rect 222 3628 232 3648
rect 242 3628 256 3648
rect 259 3635 268 3648
rect 284 3635 293 3648
rect 222 3617 256 3628
rect 259 3617 268 3633
rect 284 3617 293 3633
rect 300 3628 310 3648
rect 320 3628 334 3648
rect 335 3635 346 3648
rect 300 3617 334 3628
rect 335 3617 346 3633
rect 392 3624 408 3640
rect 415 3638 445 3690
rect 479 3686 480 3693
rect 464 3678 480 3686
rect 451 3646 464 3665
rect 479 3646 509 3662
rect 451 3630 525 3646
rect 451 3628 464 3630
rect 479 3628 513 3630
rect 116 3606 129 3608
rect 144 3606 178 3608
rect 116 3590 178 3606
rect 222 3601 238 3604
rect 300 3601 330 3612
rect 378 3608 424 3624
rect 451 3612 525 3628
rect 378 3606 412 3608
rect 377 3590 424 3606
rect 451 3590 464 3612
rect 479 3590 509 3612
rect 536 3590 537 3606
rect 552 3590 565 3750
rect 595 3646 608 3750
rect 653 3728 654 3738
rect 669 3728 682 3738
rect 653 3724 682 3728
rect 687 3724 717 3750
rect 735 3736 751 3738
rect 823 3736 876 3750
rect 824 3734 888 3736
rect 931 3734 946 3750
rect 995 3747 1025 3750
rect 995 3744 1031 3747
rect 961 3736 977 3738
rect 735 3724 750 3728
rect 653 3722 750 3724
rect 778 3722 946 3734
rect 962 3724 977 3728
rect 995 3725 1034 3744
rect 1053 3738 1060 3739
rect 1059 3731 1060 3738
rect 1043 3728 1044 3731
rect 1059 3728 1072 3731
rect 995 3724 1025 3725
rect 1034 3724 1040 3725
rect 1043 3724 1072 3728
rect 962 3723 1072 3724
rect 962 3722 1078 3723
rect 637 3714 688 3722
rect 637 3702 662 3714
rect 669 3702 688 3714
rect 719 3714 769 3722
rect 719 3706 735 3714
rect 742 3712 769 3714
rect 778 3712 999 3722
rect 742 3702 999 3712
rect 1028 3714 1078 3722
rect 1028 3705 1044 3714
rect 637 3694 688 3702
rect 735 3694 999 3702
rect 1025 3702 1044 3705
rect 1051 3702 1078 3714
rect 1025 3694 1078 3702
rect 653 3686 654 3694
rect 669 3686 682 3694
rect 653 3678 669 3686
rect 650 3671 669 3674
rect 650 3662 672 3671
rect 623 3652 672 3662
rect 623 3646 653 3652
rect 672 3647 677 3652
rect 595 3630 669 3646
rect 687 3638 717 3694
rect 752 3684 960 3694
rect 995 3690 1040 3694
rect 1043 3693 1044 3694
rect 1059 3693 1072 3694
rect 778 3654 967 3684
rect 793 3651 967 3654
rect 786 3648 967 3651
rect 595 3628 608 3630
rect 623 3628 657 3630
rect 595 3612 669 3628
rect 696 3624 709 3638
rect 724 3624 740 3640
rect 786 3635 797 3648
rect 579 3590 580 3606
rect 595 3590 608 3612
rect 623 3590 653 3612
rect 696 3608 758 3624
rect 786 3617 797 3633
rect 802 3628 812 3648
rect 822 3628 836 3648
rect 839 3635 848 3648
rect 864 3635 873 3648
rect 802 3617 836 3628
rect 839 3617 848 3633
rect 864 3617 873 3633
rect 880 3628 890 3648
rect 900 3628 914 3648
rect 915 3635 926 3648
rect 880 3617 914 3628
rect 915 3617 926 3633
rect 972 3624 988 3640
rect 995 3638 1025 3690
rect 1059 3686 1060 3693
rect 1044 3678 1060 3686
rect 1031 3646 1044 3665
rect 1059 3646 1089 3662
rect 1031 3630 1105 3646
rect 1031 3628 1044 3630
rect 1059 3628 1093 3630
rect 696 3606 709 3608
rect 724 3606 758 3608
rect 696 3590 758 3606
rect 802 3601 818 3604
rect 880 3601 910 3612
rect 958 3608 1004 3624
rect 1031 3612 1105 3628
rect 958 3606 992 3608
rect 957 3590 1004 3606
rect 1031 3590 1044 3612
rect 1059 3590 1089 3612
rect 1116 3590 1117 3606
rect 1132 3590 1145 3750
rect 1175 3646 1188 3750
rect 1233 3728 1234 3738
rect 1249 3728 1262 3738
rect 1233 3724 1262 3728
rect 1267 3724 1297 3750
rect 1315 3736 1331 3738
rect 1403 3736 1456 3750
rect 1404 3734 1468 3736
rect 1511 3734 1526 3750
rect 1575 3747 1605 3750
rect 1575 3744 1611 3747
rect 1541 3736 1557 3738
rect 1315 3724 1330 3728
rect 1233 3722 1330 3724
rect 1358 3722 1526 3734
rect 1542 3724 1557 3728
rect 1575 3725 1614 3744
rect 1633 3738 1640 3739
rect 1639 3731 1640 3738
rect 1623 3728 1624 3731
rect 1639 3728 1652 3731
rect 1575 3724 1605 3725
rect 1614 3724 1620 3725
rect 1623 3724 1652 3728
rect 1542 3723 1652 3724
rect 1542 3722 1658 3723
rect 1217 3714 1268 3722
rect 1217 3702 1242 3714
rect 1249 3702 1268 3714
rect 1299 3714 1349 3722
rect 1299 3706 1315 3714
rect 1322 3712 1349 3714
rect 1358 3712 1579 3722
rect 1322 3702 1579 3712
rect 1608 3714 1658 3722
rect 1608 3705 1624 3714
rect 1217 3694 1268 3702
rect 1315 3694 1579 3702
rect 1605 3702 1624 3705
rect 1631 3702 1658 3714
rect 1605 3694 1658 3702
rect 1233 3686 1234 3694
rect 1249 3686 1262 3694
rect 1233 3678 1249 3686
rect 1230 3671 1249 3674
rect 1230 3662 1252 3671
rect 1203 3652 1252 3662
rect 1203 3646 1233 3652
rect 1252 3647 1257 3652
rect 1175 3630 1249 3646
rect 1267 3638 1297 3694
rect 1332 3684 1540 3694
rect 1575 3690 1620 3694
rect 1623 3693 1624 3694
rect 1639 3693 1652 3694
rect 1358 3654 1547 3684
rect 1373 3651 1547 3654
rect 1366 3648 1547 3651
rect 1175 3628 1188 3630
rect 1203 3628 1237 3630
rect 1175 3612 1249 3628
rect 1276 3624 1289 3638
rect 1304 3624 1320 3640
rect 1366 3635 1377 3648
rect 1159 3590 1160 3606
rect 1175 3590 1188 3612
rect 1203 3590 1233 3612
rect 1276 3608 1338 3624
rect 1366 3617 1377 3633
rect 1382 3628 1392 3648
rect 1402 3628 1416 3648
rect 1419 3635 1428 3648
rect 1444 3635 1453 3648
rect 1382 3617 1416 3628
rect 1419 3617 1428 3633
rect 1444 3617 1453 3633
rect 1460 3628 1470 3648
rect 1480 3628 1494 3648
rect 1495 3635 1506 3648
rect 1460 3617 1494 3628
rect 1495 3617 1506 3633
rect 1552 3624 1568 3640
rect 1575 3638 1605 3690
rect 1639 3686 1640 3693
rect 1624 3678 1640 3686
rect 1611 3646 1624 3665
rect 1639 3646 1669 3662
rect 1611 3630 1685 3646
rect 1611 3628 1624 3630
rect 1639 3628 1673 3630
rect 1276 3606 1289 3608
rect 1304 3606 1338 3608
rect 1276 3590 1338 3606
rect 1382 3601 1398 3604
rect 1460 3601 1490 3612
rect 1538 3608 1584 3624
rect 1611 3612 1685 3628
rect 1538 3606 1572 3608
rect 1537 3590 1584 3606
rect 1611 3590 1624 3612
rect 1639 3590 1669 3612
rect 1696 3590 1697 3606
rect 1712 3590 1725 3750
rect 1755 3646 1768 3750
rect 1813 3728 1814 3738
rect 1829 3728 1842 3738
rect 1813 3724 1842 3728
rect 1847 3724 1877 3750
rect 1895 3736 1911 3738
rect 1983 3736 2036 3750
rect 1984 3734 2048 3736
rect 2091 3734 2106 3750
rect 2155 3747 2185 3750
rect 2155 3744 2191 3747
rect 2121 3736 2137 3738
rect 1895 3724 1910 3728
rect 1813 3722 1910 3724
rect 1938 3722 2106 3734
rect 2122 3724 2137 3728
rect 2155 3725 2194 3744
rect 2213 3738 2220 3739
rect 2219 3731 2220 3738
rect 2203 3728 2204 3731
rect 2219 3728 2232 3731
rect 2155 3724 2185 3725
rect 2194 3724 2200 3725
rect 2203 3724 2232 3728
rect 2122 3723 2232 3724
rect 2122 3722 2238 3723
rect 1797 3714 1848 3722
rect 1797 3702 1822 3714
rect 1829 3702 1848 3714
rect 1879 3714 1929 3722
rect 1879 3706 1895 3714
rect 1902 3712 1929 3714
rect 1938 3712 2159 3722
rect 1902 3702 2159 3712
rect 2188 3714 2238 3722
rect 2188 3705 2204 3714
rect 1797 3694 1848 3702
rect 1895 3694 2159 3702
rect 2185 3702 2204 3705
rect 2211 3702 2238 3714
rect 2185 3694 2238 3702
rect 1813 3686 1814 3694
rect 1829 3686 1842 3694
rect 1813 3678 1829 3686
rect 1810 3671 1829 3674
rect 1810 3662 1832 3671
rect 1783 3652 1832 3662
rect 1783 3646 1813 3652
rect 1832 3647 1837 3652
rect 1755 3630 1829 3646
rect 1847 3638 1877 3694
rect 1912 3684 2120 3694
rect 2155 3690 2200 3694
rect 2203 3693 2204 3694
rect 2219 3693 2232 3694
rect 1938 3654 2127 3684
rect 1953 3651 2127 3654
rect 1946 3648 2127 3651
rect 1755 3628 1768 3630
rect 1783 3628 1817 3630
rect 1755 3612 1829 3628
rect 1856 3624 1869 3638
rect 1884 3624 1900 3640
rect 1946 3635 1957 3648
rect 1739 3590 1740 3606
rect 1755 3590 1768 3612
rect 1783 3590 1813 3612
rect 1856 3608 1918 3624
rect 1946 3617 1957 3633
rect 1962 3628 1972 3648
rect 1982 3628 1996 3648
rect 1999 3635 2008 3648
rect 2024 3635 2033 3648
rect 1962 3617 1996 3628
rect 1999 3617 2008 3633
rect 2024 3617 2033 3633
rect 2040 3628 2050 3648
rect 2060 3628 2074 3648
rect 2075 3635 2086 3648
rect 2040 3617 2074 3628
rect 2075 3617 2086 3633
rect 2132 3624 2148 3640
rect 2155 3638 2185 3690
rect 2219 3686 2220 3693
rect 2204 3678 2220 3686
rect 2191 3646 2204 3665
rect 2219 3646 2249 3662
rect 2191 3630 2265 3646
rect 2191 3628 2204 3630
rect 2219 3628 2253 3630
rect 1856 3606 1869 3608
rect 1884 3606 1918 3608
rect 1856 3590 1918 3606
rect 1962 3601 1976 3604
rect 2040 3601 2070 3612
rect 2118 3608 2164 3624
rect 2191 3612 2265 3628
rect 2118 3606 2152 3608
rect 2117 3590 2164 3606
rect 2191 3590 2204 3612
rect 2219 3590 2249 3612
rect 2276 3590 2277 3606
rect 2292 3590 2305 3750
rect 2335 3646 2348 3750
rect 2393 3728 2394 3738
rect 2409 3728 2422 3738
rect 2393 3724 2422 3728
rect 2427 3724 2457 3750
rect 2475 3736 2491 3738
rect 2563 3736 2616 3750
rect 2564 3734 2628 3736
rect 2671 3734 2686 3750
rect 2735 3747 2765 3750
rect 2735 3744 2771 3747
rect 2701 3736 2717 3738
rect 2475 3724 2490 3728
rect 2393 3722 2490 3724
rect 2518 3722 2686 3734
rect 2702 3724 2717 3728
rect 2735 3725 2774 3744
rect 2793 3738 2800 3739
rect 2799 3731 2800 3738
rect 2783 3728 2784 3731
rect 2799 3728 2812 3731
rect 2735 3724 2765 3725
rect 2774 3724 2780 3725
rect 2783 3724 2812 3728
rect 2702 3723 2812 3724
rect 2702 3722 2818 3723
rect 2377 3714 2428 3722
rect 2377 3702 2402 3714
rect 2409 3702 2428 3714
rect 2459 3714 2509 3722
rect 2459 3706 2475 3714
rect 2482 3712 2509 3714
rect 2518 3712 2739 3722
rect 2482 3702 2739 3712
rect 2768 3714 2818 3722
rect 2768 3705 2784 3714
rect 2377 3694 2428 3702
rect 2475 3694 2739 3702
rect 2765 3702 2784 3705
rect 2791 3702 2818 3714
rect 2765 3694 2818 3702
rect 2393 3686 2394 3694
rect 2409 3686 2422 3694
rect 2393 3678 2409 3686
rect 2390 3671 2409 3674
rect 2390 3662 2412 3671
rect 2363 3652 2412 3662
rect 2363 3646 2393 3652
rect 2412 3647 2417 3652
rect 2335 3630 2409 3646
rect 2427 3638 2457 3694
rect 2492 3684 2700 3694
rect 2735 3690 2780 3694
rect 2783 3693 2784 3694
rect 2799 3693 2812 3694
rect 2518 3654 2707 3684
rect 2533 3651 2707 3654
rect 2526 3648 2707 3651
rect 2335 3628 2348 3630
rect 2363 3628 2397 3630
rect 2335 3612 2409 3628
rect 2436 3624 2449 3638
rect 2464 3624 2480 3640
rect 2526 3635 2537 3648
rect 2319 3590 2320 3606
rect 2335 3590 2348 3612
rect 2363 3590 2393 3612
rect 2436 3608 2498 3624
rect 2526 3617 2537 3633
rect 2542 3628 2552 3648
rect 2562 3628 2576 3648
rect 2579 3635 2588 3648
rect 2604 3635 2613 3648
rect 2542 3617 2576 3628
rect 2579 3617 2588 3633
rect 2604 3617 2613 3633
rect 2620 3628 2630 3648
rect 2640 3628 2654 3648
rect 2655 3635 2666 3648
rect 2620 3617 2654 3628
rect 2655 3617 2666 3633
rect 2712 3624 2728 3640
rect 2735 3638 2765 3690
rect 2799 3686 2800 3693
rect 2784 3678 2800 3686
rect 2771 3646 2784 3665
rect 2799 3646 2829 3662
rect 2771 3630 2845 3646
rect 2771 3628 2784 3630
rect 2799 3628 2833 3630
rect 2436 3606 2449 3608
rect 2464 3606 2498 3608
rect 2436 3590 2498 3606
rect 2542 3601 2558 3604
rect 2620 3601 2650 3612
rect 2698 3608 2744 3624
rect 2771 3612 2845 3628
rect 2698 3606 2732 3608
rect 2697 3590 2744 3606
rect 2771 3590 2784 3612
rect 2799 3590 2829 3612
rect 2856 3590 2857 3606
rect 2872 3590 2885 3750
rect 2915 3646 2928 3750
rect 2973 3728 2974 3738
rect 2989 3728 3002 3738
rect 2973 3724 3002 3728
rect 3007 3724 3037 3750
rect 3055 3736 3071 3738
rect 3143 3736 3196 3750
rect 3144 3734 3208 3736
rect 3251 3734 3266 3750
rect 3315 3747 3345 3750
rect 3315 3744 3351 3747
rect 3281 3736 3297 3738
rect 3055 3724 3070 3728
rect 2973 3722 3070 3724
rect 3098 3722 3266 3734
rect 3282 3724 3297 3728
rect 3315 3725 3354 3744
rect 3373 3738 3380 3739
rect 3379 3731 3380 3738
rect 3363 3728 3364 3731
rect 3379 3728 3392 3731
rect 3315 3724 3345 3725
rect 3354 3724 3360 3725
rect 3363 3724 3392 3728
rect 3282 3723 3392 3724
rect 3282 3722 3398 3723
rect 2957 3714 3008 3722
rect 2957 3702 2982 3714
rect 2989 3702 3008 3714
rect 3039 3714 3089 3722
rect 3039 3706 3055 3714
rect 3062 3712 3089 3714
rect 3098 3712 3319 3722
rect 3062 3702 3319 3712
rect 3348 3714 3398 3722
rect 3348 3705 3364 3714
rect 2957 3694 3008 3702
rect 3055 3694 3319 3702
rect 3345 3702 3364 3705
rect 3371 3702 3398 3714
rect 3345 3694 3398 3702
rect 2973 3686 2974 3694
rect 2989 3686 3002 3694
rect 2973 3678 2989 3686
rect 2970 3671 2989 3674
rect 2970 3662 2992 3671
rect 2943 3652 2992 3662
rect 2943 3646 2973 3652
rect 2992 3647 2997 3652
rect 2915 3630 2989 3646
rect 3007 3638 3037 3694
rect 3072 3684 3280 3694
rect 3315 3690 3360 3694
rect 3363 3693 3364 3694
rect 3379 3693 3392 3694
rect 3098 3654 3287 3684
rect 3113 3651 3287 3654
rect 3106 3648 3287 3651
rect 2915 3628 2928 3630
rect 2943 3628 2977 3630
rect 2915 3612 2989 3628
rect 3016 3624 3029 3638
rect 3044 3624 3060 3640
rect 3106 3635 3117 3648
rect 2899 3590 2900 3606
rect 2915 3590 2928 3612
rect 2943 3590 2973 3612
rect 3016 3608 3078 3624
rect 3106 3617 3117 3633
rect 3122 3628 3132 3648
rect 3142 3628 3156 3648
rect 3159 3635 3168 3648
rect 3184 3635 3193 3648
rect 3122 3617 3156 3628
rect 3159 3617 3168 3633
rect 3184 3617 3193 3633
rect 3200 3628 3210 3648
rect 3220 3628 3234 3648
rect 3235 3635 3246 3648
rect 3200 3617 3234 3628
rect 3235 3617 3246 3633
rect 3292 3624 3308 3640
rect 3315 3638 3345 3690
rect 3379 3686 3380 3693
rect 3364 3678 3380 3686
rect 3351 3646 3364 3665
rect 3379 3646 3409 3662
rect 3351 3630 3425 3646
rect 3351 3628 3364 3630
rect 3379 3628 3413 3630
rect 3016 3606 3029 3608
rect 3044 3606 3078 3608
rect 3016 3590 3078 3606
rect 3122 3601 3138 3604
rect 3200 3601 3230 3612
rect 3278 3608 3324 3624
rect 3351 3612 3425 3628
rect 3278 3606 3312 3608
rect 3277 3590 3324 3606
rect 3351 3590 3364 3612
rect 3379 3590 3409 3612
rect 3436 3590 3437 3606
rect 3452 3590 3465 3750
rect 3495 3646 3508 3750
rect 3553 3728 3554 3738
rect 3569 3728 3582 3738
rect 3553 3724 3582 3728
rect 3587 3724 3617 3750
rect 3635 3736 3651 3738
rect 3723 3736 3776 3750
rect 3724 3734 3788 3736
rect 3831 3734 3846 3750
rect 3895 3747 3925 3750
rect 3895 3744 3931 3747
rect 3861 3736 3877 3738
rect 3635 3724 3650 3728
rect 3553 3722 3650 3724
rect 3678 3722 3846 3734
rect 3862 3724 3877 3728
rect 3895 3725 3934 3744
rect 3953 3738 3960 3739
rect 3959 3731 3960 3738
rect 3943 3728 3944 3731
rect 3959 3728 3972 3731
rect 3895 3724 3925 3725
rect 3934 3724 3940 3725
rect 3943 3724 3972 3728
rect 3862 3723 3972 3724
rect 3862 3722 3978 3723
rect 3537 3714 3588 3722
rect 3537 3702 3562 3714
rect 3569 3702 3588 3714
rect 3619 3714 3669 3722
rect 3619 3706 3635 3714
rect 3642 3712 3669 3714
rect 3678 3712 3899 3722
rect 3642 3702 3899 3712
rect 3928 3714 3978 3722
rect 3928 3705 3944 3714
rect 3537 3694 3588 3702
rect 3635 3694 3899 3702
rect 3925 3702 3944 3705
rect 3951 3702 3978 3714
rect 3925 3694 3978 3702
rect 3553 3686 3554 3694
rect 3569 3686 3582 3694
rect 3553 3678 3569 3686
rect 3550 3671 3569 3674
rect 3550 3662 3572 3671
rect 3523 3652 3572 3662
rect 3523 3646 3553 3652
rect 3572 3647 3577 3652
rect 3495 3630 3569 3646
rect 3587 3638 3617 3694
rect 3652 3684 3860 3694
rect 3895 3690 3940 3694
rect 3943 3693 3944 3694
rect 3959 3693 3972 3694
rect 3678 3654 3867 3684
rect 3693 3651 3867 3654
rect 3686 3648 3867 3651
rect 3495 3628 3508 3630
rect 3523 3628 3557 3630
rect 3495 3612 3569 3628
rect 3596 3624 3609 3638
rect 3624 3624 3640 3640
rect 3686 3635 3697 3648
rect 3479 3590 3480 3606
rect 3495 3590 3508 3612
rect 3523 3590 3553 3612
rect 3596 3608 3658 3624
rect 3686 3617 3697 3633
rect 3702 3628 3712 3648
rect 3722 3628 3736 3648
rect 3739 3635 3748 3648
rect 3764 3635 3773 3648
rect 3702 3617 3736 3628
rect 3739 3617 3748 3633
rect 3764 3617 3773 3633
rect 3780 3628 3790 3648
rect 3800 3628 3814 3648
rect 3815 3635 3826 3648
rect 3780 3617 3814 3628
rect 3815 3617 3826 3633
rect 3872 3624 3888 3640
rect 3895 3638 3925 3690
rect 3959 3686 3960 3693
rect 3944 3678 3960 3686
rect 3931 3646 3944 3665
rect 3959 3646 3989 3662
rect 3931 3630 4005 3646
rect 3931 3628 3944 3630
rect 3959 3628 3993 3630
rect 3596 3606 3609 3608
rect 3624 3606 3658 3608
rect 3596 3590 3658 3606
rect 3702 3601 3718 3604
rect 3780 3601 3810 3612
rect 3858 3608 3904 3624
rect 3931 3612 4005 3628
rect 3858 3606 3892 3608
rect 3857 3590 3904 3606
rect 3931 3590 3944 3612
rect 3959 3590 3989 3612
rect 4016 3590 4017 3606
rect 4032 3590 4045 3750
rect 4075 3646 4088 3750
rect 4133 3728 4134 3738
rect 4149 3728 4162 3738
rect 4133 3724 4162 3728
rect 4167 3724 4197 3750
rect 4215 3736 4231 3738
rect 4303 3736 4356 3750
rect 4304 3734 4368 3736
rect 4411 3734 4426 3750
rect 4475 3747 4505 3750
rect 4475 3744 4511 3747
rect 4441 3736 4457 3738
rect 4215 3724 4230 3728
rect 4133 3722 4230 3724
rect 4258 3722 4426 3734
rect 4442 3724 4457 3728
rect 4475 3725 4514 3744
rect 4533 3738 4540 3739
rect 4539 3731 4540 3738
rect 4523 3728 4524 3731
rect 4539 3728 4552 3731
rect 4475 3724 4505 3725
rect 4514 3724 4520 3725
rect 4523 3724 4552 3728
rect 4442 3723 4552 3724
rect 4442 3722 4558 3723
rect 4117 3714 4168 3722
rect 4117 3702 4142 3714
rect 4149 3702 4168 3714
rect 4199 3714 4249 3722
rect 4199 3706 4215 3714
rect 4222 3712 4249 3714
rect 4258 3712 4479 3722
rect 4222 3702 4479 3712
rect 4508 3714 4558 3722
rect 4508 3705 4524 3714
rect 4117 3694 4168 3702
rect 4215 3694 4479 3702
rect 4505 3702 4524 3705
rect 4531 3702 4558 3714
rect 4505 3694 4558 3702
rect 4133 3686 4134 3694
rect 4149 3686 4162 3694
rect 4133 3678 4149 3686
rect 4130 3671 4149 3674
rect 4130 3662 4152 3671
rect 4103 3652 4152 3662
rect 4103 3646 4133 3652
rect 4152 3647 4157 3652
rect 4075 3630 4149 3646
rect 4167 3638 4197 3694
rect 4232 3684 4440 3694
rect 4475 3690 4520 3694
rect 4523 3693 4524 3694
rect 4539 3693 4552 3694
rect 4258 3654 4447 3684
rect 4273 3651 4447 3654
rect 4266 3648 4447 3651
rect 4075 3628 4088 3630
rect 4103 3628 4137 3630
rect 4075 3612 4149 3628
rect 4176 3624 4189 3638
rect 4204 3624 4220 3640
rect 4266 3635 4277 3648
rect 4059 3590 4060 3606
rect 4075 3590 4088 3612
rect 4103 3590 4133 3612
rect 4176 3608 4238 3624
rect 4266 3617 4277 3633
rect 4282 3628 4292 3648
rect 4302 3628 4316 3648
rect 4319 3635 4328 3648
rect 4344 3635 4353 3648
rect 4282 3617 4316 3628
rect 4319 3617 4328 3633
rect 4344 3617 4353 3633
rect 4360 3628 4370 3648
rect 4380 3628 4394 3648
rect 4395 3635 4406 3648
rect 4360 3617 4394 3628
rect 4395 3617 4406 3633
rect 4452 3624 4468 3640
rect 4475 3638 4505 3690
rect 4539 3686 4540 3693
rect 4524 3678 4540 3686
rect 4511 3646 4524 3665
rect 4539 3646 4569 3662
rect 4511 3630 4585 3646
rect 4511 3628 4524 3630
rect 4539 3628 4573 3630
rect 4176 3606 4189 3608
rect 4204 3606 4238 3608
rect 4176 3590 4238 3606
rect 4282 3601 4298 3604
rect 4360 3601 4390 3612
rect 4438 3608 4484 3624
rect 4511 3612 4585 3628
rect 4438 3606 4472 3608
rect 4437 3590 4484 3606
rect 4511 3590 4524 3612
rect 4539 3590 4569 3612
rect 4596 3590 4597 3606
rect 4612 3590 4625 3750
rect 4655 3646 4668 3750
rect 4713 3728 4714 3738
rect 4729 3728 4742 3738
rect 4713 3724 4742 3728
rect 4747 3724 4777 3750
rect 4795 3736 4811 3738
rect 4883 3736 4936 3750
rect 4884 3734 4948 3736
rect 4991 3734 5006 3750
rect 5055 3747 5085 3750
rect 5055 3744 5091 3747
rect 5021 3736 5037 3738
rect 4795 3724 4810 3728
rect 4713 3722 4810 3724
rect 4838 3722 5006 3734
rect 5022 3724 5037 3728
rect 5055 3725 5094 3744
rect 5113 3738 5120 3739
rect 5119 3731 5120 3738
rect 5103 3728 5104 3731
rect 5119 3728 5132 3731
rect 5055 3724 5085 3725
rect 5094 3724 5100 3725
rect 5103 3724 5132 3728
rect 5022 3723 5132 3724
rect 5022 3722 5138 3723
rect 4697 3714 4748 3722
rect 4697 3702 4722 3714
rect 4729 3702 4748 3714
rect 4779 3714 4829 3722
rect 4779 3706 4795 3714
rect 4802 3712 4829 3714
rect 4838 3712 5059 3722
rect 4802 3702 5059 3712
rect 5088 3714 5138 3722
rect 5088 3705 5104 3714
rect 4697 3694 4748 3702
rect 4795 3694 5059 3702
rect 5085 3702 5104 3705
rect 5111 3702 5138 3714
rect 5085 3694 5138 3702
rect 4713 3686 4714 3694
rect 4729 3686 4742 3694
rect 4713 3678 4729 3686
rect 4710 3671 4729 3674
rect 4710 3662 4732 3671
rect 4683 3652 4732 3662
rect 4683 3646 4713 3652
rect 4732 3647 4737 3652
rect 4655 3630 4729 3646
rect 4747 3638 4777 3694
rect 4812 3684 5020 3694
rect 5055 3690 5100 3694
rect 5103 3693 5104 3694
rect 5119 3693 5132 3694
rect 4838 3654 5027 3684
rect 4853 3651 5027 3654
rect 4846 3648 5027 3651
rect 4655 3628 4668 3630
rect 4683 3628 4717 3630
rect 4655 3612 4729 3628
rect 4756 3624 4769 3638
rect 4784 3624 4800 3640
rect 4846 3635 4857 3648
rect 4639 3590 4640 3606
rect 4655 3590 4668 3612
rect 4683 3590 4713 3612
rect 4756 3608 4818 3624
rect 4846 3617 4857 3633
rect 4862 3628 4872 3648
rect 4882 3628 4896 3648
rect 4899 3635 4908 3648
rect 4924 3635 4933 3648
rect 4862 3617 4896 3628
rect 4899 3617 4908 3633
rect 4924 3617 4933 3633
rect 4940 3628 4950 3648
rect 4960 3628 4974 3648
rect 4975 3635 4986 3648
rect 4940 3617 4974 3628
rect 4975 3617 4986 3633
rect 5032 3624 5048 3640
rect 5055 3638 5085 3690
rect 5119 3686 5120 3693
rect 5104 3678 5120 3686
rect 5091 3646 5104 3665
rect 5119 3646 5149 3662
rect 5091 3630 5165 3646
rect 5091 3628 5104 3630
rect 5119 3628 5153 3630
rect 4756 3606 4769 3608
rect 4784 3606 4818 3608
rect 4756 3590 4818 3606
rect 4862 3601 4878 3604
rect 4940 3601 4970 3612
rect 5018 3608 5064 3624
rect 5091 3612 5165 3628
rect 5018 3606 5052 3608
rect 5017 3590 5064 3606
rect 5091 3590 5104 3612
rect 5119 3590 5149 3612
rect 5176 3590 5177 3606
rect 5192 3590 5205 3750
rect 5235 3646 5248 3750
rect 5293 3728 5294 3738
rect 5309 3728 5322 3738
rect 5293 3724 5322 3728
rect 5327 3724 5357 3750
rect 5375 3736 5391 3738
rect 5463 3736 5516 3750
rect 5464 3734 5528 3736
rect 5571 3734 5586 3750
rect 5635 3747 5665 3750
rect 5635 3744 5671 3747
rect 5601 3736 5617 3738
rect 5375 3724 5390 3728
rect 5293 3722 5390 3724
rect 5418 3722 5586 3734
rect 5602 3724 5617 3728
rect 5635 3725 5674 3744
rect 5693 3738 5700 3739
rect 5699 3731 5700 3738
rect 5683 3728 5684 3731
rect 5699 3728 5712 3731
rect 5635 3724 5665 3725
rect 5674 3724 5680 3725
rect 5683 3724 5712 3728
rect 5602 3723 5712 3724
rect 5602 3722 5718 3723
rect 5277 3714 5328 3722
rect 5277 3702 5302 3714
rect 5309 3702 5328 3714
rect 5359 3714 5409 3722
rect 5359 3706 5375 3714
rect 5382 3712 5409 3714
rect 5418 3712 5639 3722
rect 5382 3702 5639 3712
rect 5668 3714 5718 3722
rect 5668 3705 5684 3714
rect 5277 3694 5328 3702
rect 5375 3694 5639 3702
rect 5665 3702 5684 3705
rect 5691 3702 5718 3714
rect 5665 3694 5718 3702
rect 5293 3686 5294 3694
rect 5309 3686 5322 3694
rect 5293 3678 5309 3686
rect 5290 3671 5309 3674
rect 5290 3662 5312 3671
rect 5263 3652 5312 3662
rect 5263 3646 5293 3652
rect 5312 3647 5317 3652
rect 5235 3630 5309 3646
rect 5327 3638 5357 3694
rect 5392 3684 5600 3694
rect 5635 3690 5680 3694
rect 5683 3693 5684 3694
rect 5699 3693 5712 3694
rect 5418 3654 5607 3684
rect 5433 3651 5607 3654
rect 5426 3648 5607 3651
rect 5235 3628 5248 3630
rect 5263 3628 5297 3630
rect 5235 3612 5309 3628
rect 5336 3624 5349 3638
rect 5364 3624 5380 3640
rect 5426 3635 5437 3648
rect 5219 3590 5220 3606
rect 5235 3590 5248 3612
rect 5263 3590 5293 3612
rect 5336 3608 5398 3624
rect 5426 3617 5437 3633
rect 5442 3628 5452 3648
rect 5462 3628 5476 3648
rect 5479 3635 5488 3648
rect 5504 3635 5513 3648
rect 5442 3617 5476 3628
rect 5479 3617 5488 3633
rect 5504 3617 5513 3633
rect 5520 3628 5530 3648
rect 5540 3628 5554 3648
rect 5555 3635 5566 3648
rect 5520 3617 5554 3628
rect 5555 3617 5566 3633
rect 5612 3624 5628 3640
rect 5635 3638 5665 3690
rect 5699 3686 5700 3693
rect 5684 3678 5700 3686
rect 5671 3646 5684 3665
rect 5699 3646 5729 3662
rect 5671 3630 5745 3646
rect 5671 3628 5684 3630
rect 5699 3628 5733 3630
rect 5336 3606 5349 3608
rect 5364 3606 5398 3608
rect 5336 3590 5398 3606
rect 5442 3601 5458 3604
rect 5520 3601 5550 3612
rect 5598 3608 5644 3624
rect 5671 3612 5745 3628
rect 5598 3606 5632 3608
rect 5597 3590 5644 3606
rect 5671 3590 5684 3612
rect 5699 3590 5729 3612
rect 5756 3590 5757 3606
rect 5772 3590 5785 3750
rect 5815 3646 5828 3750
rect 5873 3728 5874 3738
rect 5889 3728 5902 3738
rect 5873 3724 5902 3728
rect 5907 3724 5937 3750
rect 5955 3736 5971 3738
rect 6043 3736 6096 3750
rect 6044 3734 6108 3736
rect 6151 3734 6166 3750
rect 6215 3747 6245 3750
rect 6215 3744 6251 3747
rect 6181 3736 6197 3738
rect 5955 3724 5970 3728
rect 5873 3722 5970 3724
rect 5998 3722 6166 3734
rect 6182 3724 6197 3728
rect 6215 3725 6254 3744
rect 6273 3738 6280 3739
rect 6279 3731 6280 3738
rect 6263 3728 6264 3731
rect 6279 3728 6292 3731
rect 6215 3724 6245 3725
rect 6254 3724 6260 3725
rect 6263 3724 6292 3728
rect 6182 3723 6292 3724
rect 6182 3722 6298 3723
rect 5857 3714 5908 3722
rect 5857 3702 5882 3714
rect 5889 3702 5908 3714
rect 5939 3714 5989 3722
rect 5939 3706 5955 3714
rect 5962 3712 5989 3714
rect 5998 3712 6219 3722
rect 5962 3702 6219 3712
rect 6248 3714 6298 3722
rect 6248 3705 6264 3714
rect 5857 3694 5908 3702
rect 5955 3694 6219 3702
rect 6245 3702 6264 3705
rect 6271 3702 6298 3714
rect 6245 3694 6298 3702
rect 5873 3686 5874 3694
rect 5889 3686 5902 3694
rect 5873 3678 5889 3686
rect 5870 3671 5889 3674
rect 5870 3662 5892 3671
rect 5843 3652 5892 3662
rect 5843 3646 5873 3652
rect 5892 3647 5897 3652
rect 5815 3630 5889 3646
rect 5907 3638 5937 3694
rect 5972 3684 6180 3694
rect 6215 3690 6260 3694
rect 6263 3693 6264 3694
rect 6279 3693 6292 3694
rect 5998 3654 6187 3684
rect 6013 3651 6187 3654
rect 6006 3648 6187 3651
rect 5815 3628 5828 3630
rect 5843 3628 5877 3630
rect 5815 3612 5889 3628
rect 5916 3624 5929 3638
rect 5944 3624 5960 3640
rect 6006 3635 6017 3648
rect 5799 3590 5800 3606
rect 5815 3590 5828 3612
rect 5843 3590 5873 3612
rect 5916 3608 5978 3624
rect 6006 3617 6017 3633
rect 6022 3628 6032 3648
rect 6042 3628 6056 3648
rect 6059 3635 6068 3648
rect 6084 3635 6093 3648
rect 6022 3617 6056 3628
rect 6059 3617 6068 3633
rect 6084 3617 6093 3633
rect 6100 3628 6110 3648
rect 6120 3628 6134 3648
rect 6135 3635 6146 3648
rect 6100 3617 6134 3628
rect 6135 3617 6146 3633
rect 6192 3624 6208 3640
rect 6215 3638 6245 3690
rect 6279 3686 6280 3693
rect 6264 3678 6280 3686
rect 6251 3646 6264 3665
rect 6279 3646 6309 3662
rect 6251 3630 6325 3646
rect 6251 3628 6264 3630
rect 6279 3628 6313 3630
rect 5916 3606 5929 3608
rect 5944 3606 5978 3608
rect 5916 3590 5978 3606
rect 6022 3601 6038 3604
rect 6100 3601 6130 3612
rect 6178 3608 6224 3624
rect 6251 3612 6325 3628
rect 6178 3606 6212 3608
rect 6177 3590 6224 3606
rect 6251 3590 6264 3612
rect 6279 3590 6309 3612
rect 6336 3590 6337 3606
rect 6352 3590 6365 3750
rect 6395 3646 6408 3750
rect 6453 3728 6454 3738
rect 6469 3728 6482 3738
rect 6453 3724 6482 3728
rect 6487 3724 6517 3750
rect 6535 3736 6551 3738
rect 6623 3736 6676 3750
rect 6624 3734 6688 3736
rect 6731 3734 6746 3750
rect 6795 3747 6825 3750
rect 6795 3744 6831 3747
rect 6761 3736 6777 3738
rect 6535 3724 6550 3728
rect 6453 3722 6550 3724
rect 6578 3722 6746 3734
rect 6762 3724 6777 3728
rect 6795 3725 6834 3744
rect 6853 3738 6860 3739
rect 6859 3731 6860 3738
rect 6843 3728 6844 3731
rect 6859 3728 6872 3731
rect 6795 3724 6825 3725
rect 6834 3724 6840 3725
rect 6843 3724 6872 3728
rect 6762 3723 6872 3724
rect 6762 3722 6878 3723
rect 6437 3714 6488 3722
rect 6437 3702 6462 3714
rect 6469 3702 6488 3714
rect 6519 3714 6569 3722
rect 6519 3706 6535 3714
rect 6542 3712 6569 3714
rect 6578 3712 6799 3722
rect 6542 3702 6799 3712
rect 6828 3714 6878 3722
rect 6828 3705 6844 3714
rect 6437 3694 6488 3702
rect 6535 3694 6799 3702
rect 6825 3702 6844 3705
rect 6851 3702 6878 3714
rect 6825 3694 6878 3702
rect 6453 3686 6454 3694
rect 6469 3686 6482 3694
rect 6453 3678 6469 3686
rect 6450 3671 6469 3674
rect 6450 3662 6472 3671
rect 6423 3652 6472 3662
rect 6423 3646 6453 3652
rect 6472 3647 6477 3652
rect 6395 3630 6469 3646
rect 6487 3638 6517 3694
rect 6552 3684 6760 3694
rect 6795 3690 6840 3694
rect 6843 3693 6844 3694
rect 6859 3693 6872 3694
rect 6578 3654 6767 3684
rect 6593 3651 6767 3654
rect 6586 3648 6767 3651
rect 6395 3628 6408 3630
rect 6423 3628 6457 3630
rect 6395 3612 6469 3628
rect 6496 3624 6509 3638
rect 6524 3624 6540 3640
rect 6586 3635 6597 3648
rect 6379 3590 6380 3606
rect 6395 3590 6408 3612
rect 6423 3590 6453 3612
rect 6496 3608 6558 3624
rect 6586 3617 6597 3633
rect 6602 3628 6612 3648
rect 6622 3628 6636 3648
rect 6639 3635 6648 3648
rect 6664 3635 6673 3648
rect 6602 3617 6636 3628
rect 6639 3617 6648 3633
rect 6664 3617 6673 3633
rect 6680 3628 6690 3648
rect 6700 3628 6714 3648
rect 6715 3635 6726 3648
rect 6680 3617 6714 3628
rect 6715 3617 6726 3633
rect 6772 3624 6788 3640
rect 6795 3638 6825 3690
rect 6859 3686 6860 3693
rect 6844 3678 6860 3686
rect 6831 3646 6844 3665
rect 6859 3646 6889 3662
rect 6831 3630 6905 3646
rect 6831 3628 6844 3630
rect 6859 3628 6893 3630
rect 6496 3606 6509 3608
rect 6524 3606 6558 3608
rect 6496 3590 6558 3606
rect 6602 3601 6618 3604
rect 6680 3601 6710 3612
rect 6758 3608 6804 3624
rect 6831 3612 6905 3628
rect 6758 3606 6792 3608
rect 6757 3590 6804 3606
rect 6831 3590 6844 3612
rect 6859 3590 6889 3612
rect 6916 3590 6917 3606
rect 6932 3590 6945 3750
rect 6975 3646 6988 3750
rect 7033 3728 7034 3738
rect 7049 3728 7062 3738
rect 7033 3724 7062 3728
rect 7067 3724 7097 3750
rect 7115 3736 7131 3738
rect 7203 3736 7256 3750
rect 7204 3734 7268 3736
rect 7311 3734 7326 3750
rect 7375 3747 7405 3750
rect 7375 3744 7411 3747
rect 7341 3736 7357 3738
rect 7115 3724 7130 3728
rect 7033 3722 7130 3724
rect 7158 3722 7326 3734
rect 7342 3724 7357 3728
rect 7375 3725 7414 3744
rect 7433 3738 7440 3739
rect 7439 3731 7440 3738
rect 7423 3728 7424 3731
rect 7439 3728 7452 3731
rect 7375 3724 7405 3725
rect 7414 3724 7420 3725
rect 7423 3724 7452 3728
rect 7342 3723 7452 3724
rect 7342 3722 7458 3723
rect 7017 3714 7068 3722
rect 7017 3702 7042 3714
rect 7049 3702 7068 3714
rect 7099 3714 7149 3722
rect 7099 3706 7115 3714
rect 7122 3712 7149 3714
rect 7158 3712 7379 3722
rect 7122 3702 7379 3712
rect 7408 3714 7458 3722
rect 7408 3705 7424 3714
rect 7017 3694 7068 3702
rect 7115 3694 7379 3702
rect 7405 3702 7424 3705
rect 7431 3702 7458 3714
rect 7405 3694 7458 3702
rect 7033 3686 7034 3694
rect 7049 3686 7062 3694
rect 7033 3678 7049 3686
rect 7030 3671 7049 3674
rect 7030 3662 7052 3671
rect 7003 3652 7052 3662
rect 7003 3646 7033 3652
rect 7052 3647 7057 3652
rect 6975 3630 7049 3646
rect 7067 3638 7097 3694
rect 7132 3684 7340 3694
rect 7375 3690 7420 3694
rect 7423 3693 7424 3694
rect 7439 3693 7452 3694
rect 7158 3654 7347 3684
rect 7173 3651 7347 3654
rect 7166 3648 7347 3651
rect 6975 3628 6988 3630
rect 7003 3628 7037 3630
rect 6975 3612 7049 3628
rect 7076 3624 7089 3638
rect 7104 3624 7120 3640
rect 7166 3635 7177 3648
rect 6959 3590 6960 3606
rect 6975 3590 6988 3612
rect 7003 3590 7033 3612
rect 7076 3608 7138 3624
rect 7166 3617 7177 3633
rect 7182 3628 7192 3648
rect 7202 3628 7216 3648
rect 7219 3635 7228 3648
rect 7244 3635 7253 3648
rect 7182 3617 7216 3628
rect 7219 3617 7228 3633
rect 7244 3617 7253 3633
rect 7260 3628 7270 3648
rect 7280 3628 7294 3648
rect 7295 3635 7306 3648
rect 7260 3617 7294 3628
rect 7295 3617 7306 3633
rect 7352 3624 7368 3640
rect 7375 3638 7405 3690
rect 7439 3686 7440 3693
rect 7424 3678 7440 3686
rect 7411 3646 7424 3665
rect 7439 3646 7469 3662
rect 7411 3630 7485 3646
rect 7411 3628 7424 3630
rect 7439 3628 7473 3630
rect 7076 3606 7089 3608
rect 7104 3606 7138 3608
rect 7076 3590 7138 3606
rect 7182 3601 7198 3604
rect 7260 3601 7290 3612
rect 7338 3608 7384 3624
rect 7411 3612 7485 3628
rect 7338 3606 7372 3608
rect 7337 3590 7384 3606
rect 7411 3590 7424 3612
rect 7439 3590 7469 3612
rect 7496 3590 7497 3606
rect 7512 3590 7525 3750
rect 7555 3646 7568 3750
rect 7613 3728 7614 3738
rect 7629 3728 7642 3738
rect 7613 3724 7642 3728
rect 7647 3724 7677 3750
rect 7695 3736 7711 3738
rect 7783 3736 7836 3750
rect 7784 3734 7848 3736
rect 7891 3734 7906 3750
rect 7955 3747 7985 3750
rect 7955 3744 7991 3747
rect 7921 3736 7937 3738
rect 7695 3724 7710 3728
rect 7613 3722 7710 3724
rect 7738 3722 7906 3734
rect 7922 3724 7937 3728
rect 7955 3725 7994 3744
rect 8013 3738 8020 3739
rect 8019 3731 8020 3738
rect 8003 3728 8004 3731
rect 8019 3728 8032 3731
rect 7955 3724 7985 3725
rect 7994 3724 8000 3725
rect 8003 3724 8032 3728
rect 7922 3723 8032 3724
rect 7922 3722 8038 3723
rect 7597 3714 7648 3722
rect 7597 3702 7622 3714
rect 7629 3702 7648 3714
rect 7679 3714 7729 3722
rect 7679 3706 7695 3714
rect 7702 3712 7729 3714
rect 7738 3712 7959 3722
rect 7702 3702 7959 3712
rect 7988 3714 8038 3722
rect 7988 3705 8004 3714
rect 7597 3694 7648 3702
rect 7695 3694 7959 3702
rect 7985 3702 8004 3705
rect 8011 3702 8038 3714
rect 7985 3694 8038 3702
rect 7613 3686 7614 3694
rect 7629 3686 7642 3694
rect 7613 3678 7629 3686
rect 7610 3671 7629 3674
rect 7610 3662 7632 3671
rect 7583 3652 7632 3662
rect 7583 3646 7613 3652
rect 7632 3647 7637 3652
rect 7555 3630 7629 3646
rect 7647 3638 7677 3694
rect 7712 3684 7920 3694
rect 7955 3690 8000 3694
rect 8003 3693 8004 3694
rect 8019 3693 8032 3694
rect 7738 3654 7927 3684
rect 7753 3651 7927 3654
rect 7746 3648 7927 3651
rect 7555 3628 7568 3630
rect 7583 3628 7617 3630
rect 7555 3612 7629 3628
rect 7656 3624 7669 3638
rect 7684 3624 7700 3640
rect 7746 3635 7757 3648
rect 7539 3590 7540 3606
rect 7555 3590 7568 3612
rect 7583 3590 7613 3612
rect 7656 3608 7718 3624
rect 7746 3617 7757 3633
rect 7762 3628 7772 3648
rect 7782 3628 7796 3648
rect 7799 3635 7808 3648
rect 7824 3635 7833 3648
rect 7762 3617 7796 3628
rect 7799 3617 7808 3633
rect 7824 3617 7833 3633
rect 7840 3628 7850 3648
rect 7860 3628 7874 3648
rect 7875 3635 7886 3648
rect 7840 3617 7874 3628
rect 7875 3617 7886 3633
rect 7932 3624 7948 3640
rect 7955 3638 7985 3690
rect 8019 3686 8020 3693
rect 8004 3678 8020 3686
rect 7991 3646 8004 3665
rect 8019 3646 8049 3662
rect 7991 3630 8065 3646
rect 7991 3628 8004 3630
rect 8019 3628 8053 3630
rect 7656 3606 7669 3608
rect 7684 3606 7718 3608
rect 7656 3590 7718 3606
rect 7762 3601 7778 3604
rect 7840 3601 7870 3612
rect 7918 3608 7964 3624
rect 7991 3612 8065 3628
rect 7918 3606 7952 3608
rect 7917 3590 7964 3606
rect 7991 3590 8004 3612
rect 8019 3590 8049 3612
rect 8076 3590 8077 3606
rect 8092 3590 8105 3750
rect 8135 3646 8148 3750
rect 8193 3728 8194 3738
rect 8209 3728 8222 3738
rect 8193 3724 8222 3728
rect 8227 3724 8257 3750
rect 8275 3736 8291 3738
rect 8363 3736 8416 3750
rect 8364 3734 8428 3736
rect 8471 3734 8486 3750
rect 8535 3747 8565 3750
rect 8535 3744 8571 3747
rect 8501 3736 8517 3738
rect 8275 3724 8290 3728
rect 8193 3722 8290 3724
rect 8318 3722 8486 3734
rect 8502 3724 8517 3728
rect 8535 3725 8574 3744
rect 8593 3738 8600 3739
rect 8599 3731 8600 3738
rect 8583 3728 8584 3731
rect 8599 3728 8612 3731
rect 8535 3724 8565 3725
rect 8574 3724 8580 3725
rect 8583 3724 8612 3728
rect 8502 3723 8612 3724
rect 8502 3722 8618 3723
rect 8177 3714 8228 3722
rect 8177 3702 8202 3714
rect 8209 3702 8228 3714
rect 8259 3714 8309 3722
rect 8259 3706 8275 3714
rect 8282 3712 8309 3714
rect 8318 3712 8539 3722
rect 8282 3702 8539 3712
rect 8568 3714 8618 3722
rect 8568 3705 8584 3714
rect 8177 3694 8228 3702
rect 8275 3694 8539 3702
rect 8565 3702 8584 3705
rect 8591 3702 8618 3714
rect 8565 3694 8618 3702
rect 8193 3686 8194 3694
rect 8209 3686 8222 3694
rect 8193 3678 8209 3686
rect 8190 3671 8209 3674
rect 8190 3662 8212 3671
rect 8163 3652 8212 3662
rect 8163 3646 8193 3652
rect 8212 3647 8217 3652
rect 8135 3630 8209 3646
rect 8227 3638 8257 3694
rect 8292 3684 8500 3694
rect 8535 3690 8580 3694
rect 8583 3693 8584 3694
rect 8599 3693 8612 3694
rect 8318 3654 8507 3684
rect 8333 3651 8507 3654
rect 8326 3648 8507 3651
rect 8135 3628 8148 3630
rect 8163 3628 8197 3630
rect 8135 3612 8209 3628
rect 8236 3624 8249 3638
rect 8264 3624 8280 3640
rect 8326 3635 8337 3648
rect 8119 3590 8120 3606
rect 8135 3590 8148 3612
rect 8163 3590 8193 3612
rect 8236 3608 8298 3624
rect 8326 3617 8337 3633
rect 8342 3628 8352 3648
rect 8362 3628 8376 3648
rect 8379 3635 8388 3648
rect 8404 3635 8413 3648
rect 8342 3617 8376 3628
rect 8379 3617 8388 3633
rect 8404 3617 8413 3633
rect 8420 3628 8430 3648
rect 8440 3628 8454 3648
rect 8455 3635 8466 3648
rect 8420 3617 8454 3628
rect 8455 3617 8466 3633
rect 8512 3624 8528 3640
rect 8535 3638 8565 3690
rect 8599 3686 8600 3693
rect 8584 3678 8600 3686
rect 8571 3646 8584 3665
rect 8599 3646 8629 3662
rect 8571 3630 8645 3646
rect 8571 3628 8584 3630
rect 8599 3628 8633 3630
rect 8236 3606 8249 3608
rect 8264 3606 8298 3608
rect 8236 3590 8298 3606
rect 8342 3601 8358 3604
rect 8420 3601 8450 3612
rect 8498 3608 8544 3624
rect 8571 3612 8645 3628
rect 8498 3606 8532 3608
rect 8497 3590 8544 3606
rect 8571 3590 8584 3612
rect 8599 3590 8629 3612
rect 8656 3590 8657 3606
rect 8672 3590 8685 3750
rect 8715 3646 8728 3750
rect 8773 3728 8774 3738
rect 8789 3728 8802 3738
rect 8773 3724 8802 3728
rect 8807 3724 8837 3750
rect 8855 3736 8871 3738
rect 8943 3736 8996 3750
rect 8944 3734 9008 3736
rect 9051 3734 9066 3750
rect 9115 3747 9145 3750
rect 9115 3744 9151 3747
rect 9081 3736 9097 3738
rect 8855 3724 8870 3728
rect 8773 3722 8870 3724
rect 8898 3722 9066 3734
rect 9082 3724 9097 3728
rect 9115 3725 9154 3744
rect 9173 3738 9180 3739
rect 9179 3731 9180 3738
rect 9163 3728 9164 3731
rect 9179 3728 9192 3731
rect 9115 3724 9145 3725
rect 9154 3724 9160 3725
rect 9163 3724 9192 3728
rect 9082 3723 9192 3724
rect 9082 3722 9198 3723
rect 8757 3714 8808 3722
rect 8757 3702 8782 3714
rect 8789 3702 8808 3714
rect 8839 3714 8889 3722
rect 8839 3706 8855 3714
rect 8862 3712 8889 3714
rect 8898 3712 9119 3722
rect 8862 3702 9119 3712
rect 9148 3714 9198 3722
rect 9148 3705 9164 3714
rect 8757 3694 8808 3702
rect 8855 3694 9119 3702
rect 9145 3702 9164 3705
rect 9171 3702 9198 3714
rect 9145 3694 9198 3702
rect 8773 3686 8774 3694
rect 8789 3686 8802 3694
rect 8773 3678 8789 3686
rect 8770 3671 8789 3674
rect 8770 3662 8792 3671
rect 8743 3652 8792 3662
rect 8743 3646 8773 3652
rect 8792 3647 8797 3652
rect 8715 3630 8789 3646
rect 8807 3638 8837 3694
rect 8872 3684 9080 3694
rect 9115 3690 9160 3694
rect 9163 3693 9164 3694
rect 9179 3693 9192 3694
rect 8898 3654 9087 3684
rect 8913 3651 9087 3654
rect 8906 3648 9087 3651
rect 8715 3628 8728 3630
rect 8743 3628 8777 3630
rect 8715 3612 8789 3628
rect 8816 3624 8829 3638
rect 8844 3624 8860 3640
rect 8906 3635 8917 3648
rect 8699 3590 8700 3606
rect 8715 3590 8728 3612
rect 8743 3590 8773 3612
rect 8816 3608 8878 3624
rect 8906 3617 8917 3633
rect 8922 3628 8932 3648
rect 8942 3628 8956 3648
rect 8959 3635 8968 3648
rect 8984 3635 8993 3648
rect 8922 3617 8956 3628
rect 8959 3617 8968 3633
rect 8984 3617 8993 3633
rect 9000 3628 9010 3648
rect 9020 3628 9034 3648
rect 9035 3635 9046 3648
rect 9000 3617 9034 3628
rect 9035 3617 9046 3633
rect 9092 3624 9108 3640
rect 9115 3638 9145 3690
rect 9179 3686 9180 3693
rect 9164 3678 9180 3686
rect 9151 3646 9164 3665
rect 9179 3646 9209 3662
rect 9151 3630 9225 3646
rect 9151 3628 9164 3630
rect 9179 3628 9213 3630
rect 8816 3606 8829 3608
rect 8844 3606 8878 3608
rect 8816 3590 8878 3606
rect 8922 3601 8938 3604
rect 9000 3601 9030 3612
rect 9078 3608 9124 3624
rect 9151 3612 9225 3628
rect 9078 3606 9112 3608
rect 9077 3590 9124 3606
rect 9151 3590 9164 3612
rect 9179 3590 9209 3612
rect 9236 3590 9237 3606
rect 9252 3590 9265 3750
rect -7 3582 34 3590
rect -7 3556 8 3582
rect 15 3556 34 3582
rect 98 3578 160 3590
rect 172 3578 247 3590
rect 305 3578 380 3590
rect 392 3578 423 3590
rect 429 3578 464 3590
rect 98 3576 260 3578
rect -7 3548 34 3556
rect 116 3552 129 3576
rect 144 3574 159 3576
rect -1 3538 0 3548
rect 15 3538 28 3548
rect 43 3538 73 3552
rect 116 3538 159 3552
rect 183 3549 190 3556
rect 193 3552 260 3576
rect 292 3576 464 3578
rect 262 3554 290 3558
rect 292 3554 372 3576
rect 393 3574 408 3576
rect 262 3552 372 3554
rect 193 3548 372 3552
rect 166 3538 196 3548
rect 198 3538 351 3548
rect 359 3538 389 3548
rect 393 3538 423 3552
rect 451 3538 464 3576
rect 536 3582 571 3590
rect 536 3556 537 3582
rect 544 3556 571 3582
rect 479 3538 509 3552
rect 536 3548 571 3556
rect 573 3582 614 3590
rect 573 3556 588 3582
rect 595 3556 614 3582
rect 678 3578 740 3590
rect 752 3578 827 3590
rect 885 3578 960 3590
rect 972 3578 1003 3590
rect 1009 3578 1044 3590
rect 678 3576 840 3578
rect 573 3548 614 3556
rect 696 3552 709 3576
rect 724 3574 739 3576
rect 536 3538 537 3548
rect 552 3538 565 3548
rect 579 3538 580 3548
rect 595 3538 608 3548
rect 623 3538 653 3552
rect 696 3538 739 3552
rect 763 3549 770 3556
rect 773 3552 840 3576
rect 872 3576 1044 3578
rect 842 3554 870 3558
rect 872 3554 952 3576
rect 973 3574 988 3576
rect 842 3552 952 3554
rect 773 3548 952 3552
rect 746 3538 776 3548
rect 778 3538 931 3548
rect 939 3538 969 3548
rect 973 3538 1003 3552
rect 1031 3538 1044 3576
rect 1116 3582 1151 3590
rect 1116 3556 1117 3582
rect 1124 3556 1151 3582
rect 1059 3538 1089 3552
rect 1116 3548 1151 3556
rect 1153 3582 1194 3590
rect 1153 3556 1168 3582
rect 1175 3556 1194 3582
rect 1258 3578 1320 3590
rect 1332 3578 1407 3590
rect 1465 3578 1540 3590
rect 1552 3578 1583 3590
rect 1589 3578 1624 3590
rect 1258 3576 1420 3578
rect 1153 3548 1194 3556
rect 1276 3552 1289 3576
rect 1304 3574 1319 3576
rect 1116 3538 1117 3548
rect 1132 3538 1145 3548
rect 1159 3538 1160 3548
rect 1175 3538 1188 3548
rect 1203 3538 1233 3552
rect 1276 3538 1319 3552
rect 1343 3549 1350 3556
rect 1353 3552 1420 3576
rect 1452 3576 1624 3578
rect 1422 3554 1450 3558
rect 1452 3554 1532 3576
rect 1553 3574 1568 3576
rect 1422 3552 1532 3554
rect 1353 3548 1532 3552
rect 1326 3538 1356 3548
rect 1358 3538 1511 3548
rect 1519 3538 1549 3548
rect 1553 3538 1583 3552
rect 1611 3538 1624 3576
rect 1696 3582 1731 3590
rect 1696 3556 1697 3582
rect 1704 3556 1731 3582
rect 1639 3538 1669 3552
rect 1696 3548 1731 3556
rect 1733 3582 1774 3590
rect 1733 3556 1748 3582
rect 1755 3556 1774 3582
rect 1838 3578 1900 3590
rect 1912 3578 1987 3590
rect 2045 3578 2120 3590
rect 2132 3578 2163 3590
rect 2169 3578 2204 3590
rect 1838 3576 2000 3578
rect 1733 3548 1774 3556
rect 1856 3552 1869 3576
rect 1884 3574 1899 3576
rect 1696 3538 1697 3548
rect 1712 3538 1725 3548
rect 1739 3538 1740 3548
rect 1755 3538 1768 3548
rect 1783 3538 1813 3552
rect 1856 3538 1899 3552
rect 1923 3549 1930 3556
rect 1933 3552 2000 3576
rect 2032 3576 2204 3578
rect 2002 3554 2030 3558
rect 2032 3554 2112 3576
rect 2133 3574 2148 3576
rect 2002 3552 2112 3554
rect 1933 3548 2112 3552
rect 1906 3538 1936 3548
rect 1938 3538 2091 3548
rect 2099 3538 2129 3548
rect 2133 3538 2163 3552
rect 2191 3538 2204 3576
rect 2276 3582 2311 3590
rect 2276 3556 2277 3582
rect 2284 3556 2311 3582
rect 2219 3538 2249 3552
rect 2276 3548 2311 3556
rect 2313 3582 2354 3590
rect 2313 3556 2328 3582
rect 2335 3556 2354 3582
rect 2418 3578 2480 3590
rect 2492 3578 2567 3590
rect 2625 3578 2700 3590
rect 2712 3578 2743 3590
rect 2749 3578 2784 3590
rect 2418 3576 2580 3578
rect 2313 3548 2354 3556
rect 2436 3552 2449 3576
rect 2464 3574 2479 3576
rect 2276 3538 2277 3548
rect 2292 3538 2305 3548
rect 2319 3538 2320 3548
rect 2335 3538 2348 3548
rect 2363 3538 2393 3552
rect 2436 3538 2479 3552
rect 2503 3549 2510 3556
rect 2513 3552 2580 3576
rect 2612 3576 2784 3578
rect 2582 3554 2610 3558
rect 2612 3554 2692 3576
rect 2713 3574 2728 3576
rect 2582 3552 2692 3554
rect 2513 3548 2692 3552
rect 2486 3538 2516 3548
rect 2518 3538 2671 3548
rect 2679 3538 2709 3548
rect 2713 3538 2743 3552
rect 2771 3538 2784 3576
rect 2856 3582 2891 3590
rect 2856 3556 2857 3582
rect 2864 3556 2891 3582
rect 2799 3538 2829 3552
rect 2856 3548 2891 3556
rect 2893 3582 2934 3590
rect 2893 3556 2908 3582
rect 2915 3556 2934 3582
rect 2998 3578 3060 3590
rect 3072 3578 3147 3590
rect 3205 3578 3280 3590
rect 3292 3578 3323 3590
rect 3329 3578 3364 3590
rect 2998 3576 3160 3578
rect 2893 3548 2934 3556
rect 3016 3552 3029 3576
rect 3044 3574 3059 3576
rect 2856 3538 2857 3548
rect 2872 3538 2885 3548
rect 2899 3538 2900 3548
rect 2915 3538 2928 3548
rect 2943 3538 2973 3552
rect 3016 3538 3059 3552
rect 3083 3549 3090 3556
rect 3093 3552 3160 3576
rect 3192 3576 3364 3578
rect 3162 3554 3190 3558
rect 3192 3554 3272 3576
rect 3293 3574 3308 3576
rect 3162 3552 3272 3554
rect 3093 3548 3272 3552
rect 3066 3538 3096 3548
rect 3098 3538 3251 3548
rect 3259 3538 3289 3548
rect 3293 3538 3323 3552
rect 3351 3538 3364 3576
rect 3436 3582 3471 3590
rect 3436 3556 3437 3582
rect 3444 3556 3471 3582
rect 3379 3538 3409 3552
rect 3436 3548 3471 3556
rect 3473 3582 3514 3590
rect 3473 3556 3488 3582
rect 3495 3556 3514 3582
rect 3578 3578 3640 3590
rect 3652 3578 3727 3590
rect 3785 3578 3860 3590
rect 3872 3578 3903 3590
rect 3909 3578 3944 3590
rect 3578 3576 3740 3578
rect 3473 3548 3514 3556
rect 3596 3552 3609 3576
rect 3624 3574 3639 3576
rect 3436 3538 3437 3548
rect 3452 3538 3465 3548
rect 3479 3538 3480 3548
rect 3495 3538 3508 3548
rect 3523 3538 3553 3552
rect 3596 3538 3639 3552
rect 3663 3549 3670 3556
rect 3673 3552 3740 3576
rect 3772 3576 3944 3578
rect 3742 3554 3770 3558
rect 3772 3554 3852 3576
rect 3873 3574 3888 3576
rect 3742 3552 3852 3554
rect 3673 3548 3852 3552
rect 3646 3538 3676 3548
rect 3678 3538 3831 3548
rect 3839 3538 3869 3548
rect 3873 3538 3903 3552
rect 3931 3538 3944 3576
rect 4016 3582 4051 3590
rect 4016 3556 4017 3582
rect 4024 3556 4051 3582
rect 3959 3538 3989 3552
rect 4016 3548 4051 3556
rect 4053 3582 4094 3590
rect 4053 3556 4068 3582
rect 4075 3556 4094 3582
rect 4158 3578 4220 3590
rect 4232 3578 4307 3590
rect 4365 3578 4440 3590
rect 4452 3578 4483 3590
rect 4489 3578 4524 3590
rect 4158 3576 4320 3578
rect 4053 3548 4094 3556
rect 4176 3552 4189 3576
rect 4204 3574 4219 3576
rect 4016 3538 4017 3548
rect 4032 3538 4045 3548
rect 4059 3538 4060 3548
rect 4075 3538 4088 3548
rect 4103 3538 4133 3552
rect 4176 3538 4219 3552
rect 4243 3549 4250 3556
rect 4253 3552 4320 3576
rect 4352 3576 4524 3578
rect 4322 3554 4350 3558
rect 4352 3554 4432 3576
rect 4453 3574 4468 3576
rect 4322 3552 4432 3554
rect 4253 3548 4432 3552
rect 4226 3538 4256 3548
rect 4258 3538 4411 3548
rect 4419 3538 4449 3548
rect 4453 3538 4483 3552
rect 4511 3538 4524 3576
rect 4596 3582 4631 3590
rect 4596 3556 4597 3582
rect 4604 3556 4631 3582
rect 4539 3538 4569 3552
rect 4596 3548 4631 3556
rect 4633 3582 4674 3590
rect 4633 3556 4648 3582
rect 4655 3556 4674 3582
rect 4738 3578 4800 3590
rect 4812 3578 4887 3590
rect 4945 3578 5020 3590
rect 5032 3578 5063 3590
rect 5069 3578 5104 3590
rect 4738 3576 4900 3578
rect 4633 3548 4674 3556
rect 4756 3552 4769 3576
rect 4784 3574 4799 3576
rect 4596 3538 4597 3548
rect 4612 3538 4625 3548
rect 4639 3538 4640 3548
rect 4655 3538 4668 3548
rect 4683 3538 4713 3552
rect 4756 3538 4799 3552
rect 4823 3549 4830 3556
rect 4833 3552 4900 3576
rect 4932 3576 5104 3578
rect 4902 3554 4930 3558
rect 4932 3554 5012 3576
rect 5033 3574 5048 3576
rect 4902 3552 5012 3554
rect 4833 3548 5012 3552
rect 4806 3538 4836 3548
rect 4838 3538 4991 3548
rect 4999 3538 5029 3548
rect 5033 3538 5063 3552
rect 5091 3538 5104 3576
rect 5176 3582 5211 3590
rect 5176 3556 5177 3582
rect 5184 3556 5211 3582
rect 5119 3538 5149 3552
rect 5176 3548 5211 3556
rect 5213 3582 5254 3590
rect 5213 3556 5228 3582
rect 5235 3556 5254 3582
rect 5318 3578 5380 3590
rect 5392 3578 5467 3590
rect 5525 3578 5600 3590
rect 5612 3578 5643 3590
rect 5649 3578 5684 3590
rect 5318 3576 5480 3578
rect 5213 3548 5254 3556
rect 5336 3552 5349 3576
rect 5364 3574 5379 3576
rect 5176 3538 5177 3548
rect 5192 3538 5205 3548
rect 5219 3538 5220 3548
rect 5235 3538 5248 3548
rect 5263 3538 5293 3552
rect 5336 3538 5379 3552
rect 5403 3549 5410 3556
rect 5413 3552 5480 3576
rect 5512 3576 5684 3578
rect 5482 3554 5510 3558
rect 5512 3554 5592 3576
rect 5613 3574 5628 3576
rect 5482 3552 5592 3554
rect 5413 3548 5592 3552
rect 5386 3538 5416 3548
rect 5418 3538 5571 3548
rect 5579 3538 5609 3548
rect 5613 3538 5643 3552
rect 5671 3538 5684 3576
rect 5756 3582 5791 3590
rect 5756 3556 5757 3582
rect 5764 3556 5791 3582
rect 5699 3538 5729 3552
rect 5756 3548 5791 3556
rect 5793 3582 5834 3590
rect 5793 3556 5808 3582
rect 5815 3556 5834 3582
rect 5898 3578 5960 3590
rect 5972 3578 6047 3590
rect 6105 3578 6180 3590
rect 6192 3578 6223 3590
rect 6229 3578 6264 3590
rect 5898 3576 6060 3578
rect 5793 3548 5834 3556
rect 5916 3552 5929 3576
rect 5944 3574 5959 3576
rect 5756 3538 5757 3548
rect 5772 3538 5785 3548
rect 5799 3538 5800 3548
rect 5815 3538 5828 3548
rect 5843 3538 5873 3552
rect 5916 3538 5959 3552
rect 5983 3549 5990 3556
rect 5993 3552 6060 3576
rect 6092 3576 6264 3578
rect 6062 3554 6090 3558
rect 6092 3554 6172 3576
rect 6193 3574 6208 3576
rect 6062 3552 6172 3554
rect 5993 3548 6172 3552
rect 5966 3538 5996 3548
rect 5998 3538 6151 3548
rect 6159 3538 6189 3548
rect 6193 3538 6223 3552
rect 6251 3538 6264 3576
rect 6336 3582 6371 3590
rect 6336 3556 6337 3582
rect 6344 3556 6371 3582
rect 6279 3538 6309 3552
rect 6336 3548 6371 3556
rect 6373 3582 6414 3590
rect 6373 3556 6388 3582
rect 6395 3556 6414 3582
rect 6478 3578 6540 3590
rect 6552 3578 6627 3590
rect 6685 3578 6760 3590
rect 6772 3578 6803 3590
rect 6809 3578 6844 3590
rect 6478 3576 6640 3578
rect 6373 3548 6414 3556
rect 6496 3552 6509 3576
rect 6524 3574 6539 3576
rect 6336 3538 6337 3548
rect 6352 3538 6365 3548
rect 6379 3538 6380 3548
rect 6395 3538 6408 3548
rect 6423 3538 6453 3552
rect 6496 3538 6539 3552
rect 6563 3549 6570 3556
rect 6573 3552 6640 3576
rect 6672 3576 6844 3578
rect 6642 3554 6670 3558
rect 6672 3554 6752 3576
rect 6773 3574 6788 3576
rect 6642 3552 6752 3554
rect 6573 3548 6752 3552
rect 6546 3538 6576 3548
rect 6578 3538 6731 3548
rect 6739 3538 6769 3548
rect 6773 3538 6803 3552
rect 6831 3538 6844 3576
rect 6916 3582 6951 3590
rect 6916 3556 6917 3582
rect 6924 3556 6951 3582
rect 6859 3538 6889 3552
rect 6916 3548 6951 3556
rect 6953 3582 6994 3590
rect 6953 3556 6968 3582
rect 6975 3556 6994 3582
rect 7058 3578 7120 3590
rect 7132 3578 7207 3590
rect 7265 3578 7340 3590
rect 7352 3578 7383 3590
rect 7389 3578 7424 3590
rect 7058 3576 7220 3578
rect 6953 3548 6994 3556
rect 7076 3552 7089 3576
rect 7104 3574 7119 3576
rect 6916 3538 6917 3548
rect 6932 3538 6945 3548
rect 6959 3538 6960 3548
rect 6975 3538 6988 3548
rect 7003 3538 7033 3552
rect 7076 3538 7119 3552
rect 7143 3549 7150 3556
rect 7153 3552 7220 3576
rect 7252 3576 7424 3578
rect 7222 3554 7250 3558
rect 7252 3554 7332 3576
rect 7353 3574 7368 3576
rect 7222 3552 7332 3554
rect 7153 3548 7332 3552
rect 7126 3538 7156 3548
rect 7158 3538 7311 3548
rect 7319 3538 7349 3548
rect 7353 3538 7383 3552
rect 7411 3538 7424 3576
rect 7496 3582 7531 3590
rect 7496 3556 7497 3582
rect 7504 3556 7531 3582
rect 7439 3538 7469 3552
rect 7496 3548 7531 3556
rect 7533 3582 7574 3590
rect 7533 3556 7548 3582
rect 7555 3556 7574 3582
rect 7638 3578 7700 3590
rect 7712 3578 7787 3590
rect 7845 3578 7920 3590
rect 7932 3578 7963 3590
rect 7969 3578 8004 3590
rect 7638 3576 7800 3578
rect 7533 3548 7574 3556
rect 7656 3552 7669 3576
rect 7684 3574 7699 3576
rect 7496 3538 7497 3548
rect 7512 3538 7525 3548
rect 7539 3538 7540 3548
rect 7555 3538 7568 3548
rect 7583 3538 7613 3552
rect 7656 3538 7699 3552
rect 7723 3549 7730 3556
rect 7733 3552 7800 3576
rect 7832 3576 8004 3578
rect 7802 3554 7830 3558
rect 7832 3554 7912 3576
rect 7933 3574 7948 3576
rect 7802 3552 7912 3554
rect 7733 3548 7912 3552
rect 7706 3538 7736 3548
rect 7738 3538 7891 3548
rect 7899 3538 7929 3548
rect 7933 3538 7963 3552
rect 7991 3538 8004 3576
rect 8076 3582 8111 3590
rect 8076 3556 8077 3582
rect 8084 3556 8111 3582
rect 8019 3538 8049 3552
rect 8076 3548 8111 3556
rect 8113 3582 8154 3590
rect 8113 3556 8128 3582
rect 8135 3556 8154 3582
rect 8218 3578 8280 3590
rect 8292 3578 8367 3590
rect 8425 3578 8500 3590
rect 8512 3578 8543 3590
rect 8549 3578 8584 3590
rect 8218 3576 8380 3578
rect 8113 3548 8154 3556
rect 8236 3552 8249 3576
rect 8264 3574 8279 3576
rect 8076 3538 8077 3548
rect 8092 3538 8105 3548
rect 8119 3538 8120 3548
rect 8135 3538 8148 3548
rect 8163 3538 8193 3552
rect 8236 3538 8279 3552
rect 8303 3549 8310 3556
rect 8313 3552 8380 3576
rect 8412 3576 8584 3578
rect 8382 3554 8410 3558
rect 8412 3554 8492 3576
rect 8513 3574 8528 3576
rect 8382 3552 8492 3554
rect 8313 3548 8492 3552
rect 8286 3538 8316 3548
rect 8318 3538 8471 3548
rect 8479 3538 8509 3548
rect 8513 3538 8543 3552
rect 8571 3538 8584 3576
rect 8656 3582 8691 3590
rect 8656 3556 8657 3582
rect 8664 3556 8691 3582
rect 8599 3538 8629 3552
rect 8656 3548 8691 3556
rect 8693 3582 8734 3590
rect 8693 3556 8708 3582
rect 8715 3556 8734 3582
rect 8798 3578 8860 3590
rect 8872 3578 8947 3590
rect 9005 3578 9080 3590
rect 9092 3578 9123 3590
rect 9129 3578 9164 3590
rect 8798 3576 8960 3578
rect 8693 3548 8734 3556
rect 8816 3552 8829 3576
rect 8844 3574 8859 3576
rect 8656 3538 8657 3548
rect 8672 3538 8685 3548
rect 8699 3538 8700 3548
rect 8715 3538 8728 3548
rect 8743 3538 8773 3552
rect 8816 3538 8859 3552
rect 8883 3549 8890 3556
rect 8893 3552 8960 3576
rect 8992 3576 9164 3578
rect 8962 3554 8990 3558
rect 8992 3554 9072 3576
rect 9093 3574 9108 3576
rect 8962 3552 9072 3554
rect 8893 3548 9072 3552
rect 8866 3538 8896 3548
rect 8898 3538 9051 3548
rect 9059 3538 9089 3548
rect 9093 3538 9123 3552
rect 9151 3538 9164 3576
rect 9236 3582 9271 3590
rect 9236 3556 9237 3582
rect 9244 3556 9271 3582
rect 9179 3538 9209 3552
rect 9236 3548 9271 3556
rect 9236 3538 9237 3548
rect 9252 3538 9265 3548
rect -1 3532 9265 3538
rect 0 3524 9265 3532
rect 15 3494 28 3524
rect 43 3506 73 3524
rect 116 3510 130 3524
rect 166 3510 386 3524
rect 117 3508 130 3510
rect 83 3496 98 3508
rect 80 3494 102 3496
rect 107 3494 137 3508
rect 198 3506 351 3510
rect 180 3494 372 3506
rect 415 3494 445 3508
rect 451 3494 464 3524
rect 479 3506 509 3524
rect 552 3494 565 3524
rect 595 3494 608 3524
rect 623 3506 653 3524
rect 696 3510 710 3524
rect 746 3510 966 3524
rect 697 3508 710 3510
rect 663 3496 678 3508
rect 660 3494 682 3496
rect 687 3494 717 3508
rect 778 3506 931 3510
rect 760 3494 952 3506
rect 995 3494 1025 3508
rect 1031 3494 1044 3524
rect 1059 3506 1089 3524
rect 1132 3494 1145 3524
rect 1175 3494 1188 3524
rect 1203 3506 1233 3524
rect 1276 3510 1290 3524
rect 1326 3510 1546 3524
rect 1277 3508 1290 3510
rect 1243 3496 1258 3508
rect 1240 3494 1262 3496
rect 1267 3494 1297 3508
rect 1358 3506 1511 3510
rect 1340 3494 1532 3506
rect 1575 3494 1605 3508
rect 1611 3494 1624 3524
rect 1639 3506 1669 3524
rect 1712 3494 1725 3524
rect 1755 3494 1768 3524
rect 1783 3506 1813 3524
rect 1856 3510 1870 3524
rect 1906 3510 2126 3524
rect 1857 3508 1870 3510
rect 1823 3496 1838 3508
rect 1820 3494 1842 3496
rect 1847 3494 1877 3508
rect 1938 3506 2091 3510
rect 1920 3494 2112 3506
rect 2155 3494 2185 3508
rect 2191 3494 2204 3524
rect 2219 3506 2249 3524
rect 2292 3494 2305 3524
rect 2335 3494 2348 3524
rect 2363 3506 2393 3524
rect 2436 3510 2450 3524
rect 2486 3510 2706 3524
rect 2437 3508 2450 3510
rect 2403 3496 2418 3508
rect 2400 3494 2422 3496
rect 2427 3494 2457 3508
rect 2518 3506 2671 3510
rect 2500 3494 2692 3506
rect 2735 3494 2765 3508
rect 2771 3494 2784 3524
rect 2799 3506 2829 3524
rect 2872 3494 2885 3524
rect 2915 3494 2928 3524
rect 2943 3506 2973 3524
rect 3016 3510 3030 3524
rect 3066 3510 3286 3524
rect 3017 3508 3030 3510
rect 2983 3496 2998 3508
rect 2980 3494 3002 3496
rect 3007 3494 3037 3508
rect 3098 3506 3251 3510
rect 3080 3494 3272 3506
rect 3315 3494 3345 3508
rect 3351 3494 3364 3524
rect 3379 3506 3409 3524
rect 3452 3494 3465 3524
rect 3495 3494 3508 3524
rect 3523 3506 3553 3524
rect 3596 3510 3610 3524
rect 3646 3510 3866 3524
rect 3597 3508 3610 3510
rect 3563 3496 3578 3508
rect 3560 3494 3582 3496
rect 3587 3494 3617 3508
rect 3678 3506 3831 3510
rect 3660 3494 3852 3506
rect 3895 3494 3925 3508
rect 3931 3494 3944 3524
rect 3959 3506 3989 3524
rect 4032 3494 4045 3524
rect 4075 3494 4088 3524
rect 4103 3506 4133 3524
rect 4176 3510 4190 3524
rect 4226 3510 4446 3524
rect 4177 3508 4190 3510
rect 4143 3496 4158 3508
rect 4140 3494 4162 3496
rect 4167 3494 4197 3508
rect 4258 3506 4411 3510
rect 4240 3494 4432 3506
rect 4475 3494 4505 3508
rect 4511 3494 4524 3524
rect 4539 3506 4569 3524
rect 4612 3494 4625 3524
rect 4655 3494 4668 3524
rect 4683 3506 4713 3524
rect 4756 3510 4770 3524
rect 4806 3510 5026 3524
rect 4757 3508 4770 3510
rect 4723 3496 4738 3508
rect 4720 3494 4742 3496
rect 4747 3494 4777 3508
rect 4838 3506 4991 3510
rect 4820 3494 5012 3506
rect 5055 3494 5085 3508
rect 5091 3494 5104 3524
rect 5119 3506 5149 3524
rect 5192 3494 5205 3524
rect 5235 3494 5248 3524
rect 5263 3506 5293 3524
rect 5336 3510 5350 3524
rect 5386 3510 5606 3524
rect 5337 3508 5350 3510
rect 5303 3496 5318 3508
rect 5300 3494 5322 3496
rect 5327 3494 5357 3508
rect 5418 3506 5571 3510
rect 5400 3494 5592 3506
rect 5635 3494 5665 3508
rect 5671 3494 5684 3524
rect 5699 3506 5729 3524
rect 5772 3494 5785 3524
rect 5815 3494 5828 3524
rect 5843 3506 5873 3524
rect 5916 3510 5930 3524
rect 5966 3510 6186 3524
rect 5917 3508 5930 3510
rect 5883 3496 5898 3508
rect 5880 3494 5902 3496
rect 5907 3494 5937 3508
rect 5998 3506 6151 3510
rect 5980 3494 6172 3506
rect 6215 3494 6245 3508
rect 6251 3494 6264 3524
rect 6279 3506 6309 3524
rect 6352 3494 6365 3524
rect 6395 3494 6408 3524
rect 6423 3506 6453 3524
rect 6496 3510 6510 3524
rect 6546 3510 6766 3524
rect 6497 3508 6510 3510
rect 6463 3496 6478 3508
rect 6460 3494 6482 3496
rect 6487 3494 6517 3508
rect 6578 3506 6731 3510
rect 6560 3494 6752 3506
rect 6795 3494 6825 3508
rect 6831 3494 6844 3524
rect 6859 3506 6889 3524
rect 6932 3494 6945 3524
rect 6975 3494 6988 3524
rect 7003 3506 7033 3524
rect 7076 3510 7090 3524
rect 7126 3510 7346 3524
rect 7077 3508 7090 3510
rect 7043 3496 7058 3508
rect 7040 3494 7062 3496
rect 7067 3494 7097 3508
rect 7158 3506 7311 3510
rect 7140 3494 7332 3506
rect 7375 3494 7405 3508
rect 7411 3494 7424 3524
rect 7439 3506 7469 3524
rect 7512 3494 7525 3524
rect 7555 3494 7568 3524
rect 7583 3506 7613 3524
rect 7656 3510 7670 3524
rect 7706 3510 7926 3524
rect 7657 3508 7670 3510
rect 7623 3496 7638 3508
rect 7620 3494 7642 3496
rect 7647 3494 7677 3508
rect 7738 3506 7891 3510
rect 7720 3494 7912 3506
rect 7955 3494 7985 3508
rect 7991 3494 8004 3524
rect 8019 3506 8049 3524
rect 8092 3494 8105 3524
rect 8135 3494 8148 3524
rect 8163 3506 8193 3524
rect 8236 3510 8250 3524
rect 8286 3510 8506 3524
rect 8237 3508 8250 3510
rect 8203 3496 8218 3508
rect 8200 3494 8222 3496
rect 8227 3494 8257 3508
rect 8318 3506 8471 3510
rect 8300 3494 8492 3506
rect 8535 3494 8565 3508
rect 8571 3494 8584 3524
rect 8599 3506 8629 3524
rect 8672 3494 8685 3524
rect 8715 3494 8728 3524
rect 8743 3506 8773 3524
rect 8816 3510 8830 3524
rect 8866 3510 9086 3524
rect 8817 3508 8830 3510
rect 8783 3496 8798 3508
rect 8780 3494 8802 3496
rect 8807 3494 8837 3508
rect 8898 3506 9051 3510
rect 8880 3494 9072 3506
rect 9115 3494 9145 3508
rect 9151 3494 9164 3524
rect 9179 3506 9209 3524
rect 9252 3494 9265 3524
rect 0 3480 9265 3494
rect 15 3376 28 3480
rect 73 3458 74 3468
rect 89 3458 102 3468
rect 73 3454 102 3458
rect 107 3454 137 3480
rect 155 3466 171 3468
rect 243 3466 296 3480
rect 244 3464 308 3466
rect 351 3464 366 3480
rect 415 3477 445 3480
rect 415 3474 451 3477
rect 381 3466 397 3468
rect 155 3454 170 3458
rect 73 3452 170 3454
rect 198 3452 366 3464
rect 382 3454 397 3458
rect 415 3455 454 3474
rect 473 3468 480 3469
rect 479 3461 480 3468
rect 463 3458 464 3461
rect 479 3458 492 3461
rect 415 3454 445 3455
rect 454 3454 460 3455
rect 463 3454 492 3458
rect 382 3453 492 3454
rect 382 3452 498 3453
rect 57 3444 108 3452
rect 57 3432 82 3444
rect 89 3432 108 3444
rect 139 3444 189 3452
rect 139 3436 155 3444
rect 162 3442 189 3444
rect 198 3442 419 3452
rect 162 3432 419 3442
rect 448 3444 498 3452
rect 448 3435 464 3444
rect 57 3424 108 3432
rect 155 3424 419 3432
rect 445 3432 464 3435
rect 471 3432 498 3444
rect 445 3424 498 3432
rect 73 3416 74 3424
rect 89 3416 102 3424
rect 73 3408 89 3416
rect 70 3401 89 3404
rect 70 3392 92 3401
rect 43 3382 92 3392
rect 43 3376 73 3382
rect 92 3377 97 3382
rect 15 3360 89 3376
rect 107 3368 137 3424
rect 172 3414 380 3424
rect 415 3420 460 3424
rect 463 3423 464 3424
rect 479 3423 492 3424
rect 198 3384 387 3414
rect 213 3381 387 3384
rect 206 3378 387 3381
rect 15 3358 28 3360
rect 43 3358 77 3360
rect 15 3342 89 3358
rect 116 3354 129 3368
rect 144 3354 160 3370
rect 206 3365 217 3378
rect -1 3320 0 3336
rect 15 3320 28 3342
rect 43 3320 73 3342
rect 116 3338 178 3354
rect 206 3347 217 3363
rect 222 3358 232 3378
rect 242 3358 256 3378
rect 259 3365 268 3378
rect 284 3365 293 3378
rect 222 3347 256 3358
rect 259 3347 268 3363
rect 284 3347 293 3363
rect 300 3358 310 3378
rect 320 3358 334 3378
rect 335 3365 346 3378
rect 300 3347 334 3358
rect 335 3347 346 3363
rect 392 3354 408 3370
rect 415 3368 445 3420
rect 479 3416 480 3423
rect 464 3408 480 3416
rect 451 3376 464 3395
rect 479 3376 509 3392
rect 451 3360 525 3376
rect 451 3358 464 3360
rect 479 3358 513 3360
rect 116 3336 129 3338
rect 144 3336 178 3338
rect 116 3320 178 3336
rect 222 3331 238 3334
rect 300 3331 330 3342
rect 378 3338 424 3354
rect 451 3342 525 3358
rect 378 3336 412 3338
rect 377 3320 424 3336
rect 451 3320 464 3342
rect 479 3320 509 3342
rect 536 3320 537 3336
rect 552 3320 565 3480
rect 595 3376 608 3480
rect 653 3458 654 3468
rect 669 3458 682 3468
rect 653 3454 682 3458
rect 687 3454 717 3480
rect 735 3466 751 3468
rect 823 3466 876 3480
rect 824 3464 888 3466
rect 931 3464 946 3480
rect 995 3477 1025 3480
rect 995 3474 1031 3477
rect 961 3466 977 3468
rect 735 3454 750 3458
rect 653 3452 750 3454
rect 778 3452 946 3464
rect 962 3454 977 3458
rect 995 3455 1034 3474
rect 1053 3468 1060 3469
rect 1059 3461 1060 3468
rect 1043 3458 1044 3461
rect 1059 3458 1072 3461
rect 995 3454 1025 3455
rect 1034 3454 1040 3455
rect 1043 3454 1072 3458
rect 962 3453 1072 3454
rect 962 3452 1078 3453
rect 637 3444 688 3452
rect 637 3432 662 3444
rect 669 3432 688 3444
rect 719 3444 769 3452
rect 719 3436 735 3444
rect 742 3442 769 3444
rect 778 3442 999 3452
rect 742 3432 999 3442
rect 1028 3444 1078 3452
rect 1028 3435 1044 3444
rect 637 3424 688 3432
rect 735 3424 999 3432
rect 1025 3432 1044 3435
rect 1051 3432 1078 3444
rect 1025 3424 1078 3432
rect 653 3416 654 3424
rect 669 3416 682 3424
rect 653 3408 669 3416
rect 650 3401 669 3404
rect 650 3392 672 3401
rect 623 3382 672 3392
rect 623 3376 653 3382
rect 672 3377 677 3382
rect 595 3360 669 3376
rect 687 3368 717 3424
rect 752 3414 960 3424
rect 995 3420 1040 3424
rect 1043 3423 1044 3424
rect 1059 3423 1072 3424
rect 778 3384 967 3414
rect 793 3381 967 3384
rect 786 3378 967 3381
rect 595 3358 608 3360
rect 623 3358 657 3360
rect 595 3342 669 3358
rect 696 3354 709 3368
rect 724 3354 740 3370
rect 786 3365 797 3378
rect 579 3320 580 3336
rect 595 3320 608 3342
rect 623 3320 653 3342
rect 696 3338 758 3354
rect 786 3347 797 3363
rect 802 3358 812 3378
rect 822 3358 836 3378
rect 839 3365 848 3378
rect 864 3365 873 3378
rect 802 3347 836 3358
rect 839 3347 848 3363
rect 864 3347 873 3363
rect 880 3358 890 3378
rect 900 3358 914 3378
rect 915 3365 926 3378
rect 880 3347 914 3358
rect 915 3347 926 3363
rect 972 3354 988 3370
rect 995 3368 1025 3420
rect 1059 3416 1060 3423
rect 1044 3408 1060 3416
rect 1031 3376 1044 3395
rect 1059 3376 1089 3392
rect 1031 3360 1105 3376
rect 1031 3358 1044 3360
rect 1059 3358 1093 3360
rect 696 3336 709 3338
rect 724 3336 758 3338
rect 696 3320 758 3336
rect 802 3331 818 3334
rect 880 3331 910 3342
rect 958 3338 1004 3354
rect 1031 3342 1105 3358
rect 958 3336 992 3338
rect 957 3320 1004 3336
rect 1031 3320 1044 3342
rect 1059 3320 1089 3342
rect 1116 3320 1117 3336
rect 1132 3320 1145 3480
rect 1175 3376 1188 3480
rect 1233 3458 1234 3468
rect 1249 3458 1262 3468
rect 1233 3454 1262 3458
rect 1267 3454 1297 3480
rect 1315 3466 1331 3468
rect 1403 3466 1456 3480
rect 1404 3464 1468 3466
rect 1511 3464 1526 3480
rect 1575 3477 1605 3480
rect 1575 3474 1611 3477
rect 1541 3466 1557 3468
rect 1315 3454 1330 3458
rect 1233 3452 1330 3454
rect 1358 3452 1526 3464
rect 1542 3454 1557 3458
rect 1575 3455 1614 3474
rect 1633 3468 1640 3469
rect 1639 3461 1640 3468
rect 1623 3458 1624 3461
rect 1639 3458 1652 3461
rect 1575 3454 1605 3455
rect 1614 3454 1620 3455
rect 1623 3454 1652 3458
rect 1542 3453 1652 3454
rect 1542 3452 1658 3453
rect 1217 3444 1268 3452
rect 1217 3432 1242 3444
rect 1249 3432 1268 3444
rect 1299 3444 1349 3452
rect 1299 3436 1315 3444
rect 1322 3442 1349 3444
rect 1358 3442 1579 3452
rect 1322 3432 1579 3442
rect 1608 3444 1658 3452
rect 1608 3435 1624 3444
rect 1217 3424 1268 3432
rect 1315 3424 1579 3432
rect 1605 3432 1624 3435
rect 1631 3432 1658 3444
rect 1605 3424 1658 3432
rect 1233 3416 1234 3424
rect 1249 3416 1262 3424
rect 1233 3408 1249 3416
rect 1230 3401 1249 3404
rect 1230 3392 1252 3401
rect 1203 3382 1252 3392
rect 1203 3376 1233 3382
rect 1252 3377 1257 3382
rect 1175 3360 1249 3376
rect 1267 3368 1297 3424
rect 1332 3414 1540 3424
rect 1575 3420 1620 3424
rect 1623 3423 1624 3424
rect 1639 3423 1652 3424
rect 1358 3384 1547 3414
rect 1373 3381 1547 3384
rect 1366 3378 1547 3381
rect 1175 3358 1188 3360
rect 1203 3358 1237 3360
rect 1175 3342 1249 3358
rect 1276 3354 1289 3368
rect 1304 3354 1320 3370
rect 1366 3365 1377 3378
rect 1159 3320 1160 3336
rect 1175 3320 1188 3342
rect 1203 3320 1233 3342
rect 1276 3338 1338 3354
rect 1366 3347 1377 3363
rect 1382 3358 1392 3378
rect 1402 3358 1416 3378
rect 1419 3365 1428 3378
rect 1444 3365 1453 3378
rect 1382 3347 1416 3358
rect 1419 3347 1428 3363
rect 1444 3347 1453 3363
rect 1460 3358 1470 3378
rect 1480 3358 1494 3378
rect 1495 3365 1506 3378
rect 1460 3347 1494 3358
rect 1495 3347 1506 3363
rect 1552 3354 1568 3370
rect 1575 3368 1605 3420
rect 1639 3416 1640 3423
rect 1624 3408 1640 3416
rect 1611 3376 1624 3395
rect 1639 3376 1669 3392
rect 1611 3360 1685 3376
rect 1611 3358 1624 3360
rect 1639 3358 1673 3360
rect 1276 3336 1289 3338
rect 1304 3336 1338 3338
rect 1276 3320 1338 3336
rect 1382 3331 1398 3334
rect 1460 3331 1490 3342
rect 1538 3338 1584 3354
rect 1611 3342 1685 3358
rect 1538 3336 1572 3338
rect 1537 3320 1584 3336
rect 1611 3320 1624 3342
rect 1639 3320 1669 3342
rect 1696 3320 1697 3336
rect 1712 3320 1725 3480
rect 1755 3376 1768 3480
rect 1813 3458 1814 3468
rect 1829 3458 1842 3468
rect 1813 3454 1842 3458
rect 1847 3454 1877 3480
rect 1895 3466 1911 3468
rect 1983 3466 2036 3480
rect 1984 3464 2048 3466
rect 2091 3464 2106 3480
rect 2155 3477 2185 3480
rect 2155 3474 2191 3477
rect 2121 3466 2137 3468
rect 1895 3454 1910 3458
rect 1813 3452 1910 3454
rect 1938 3452 2106 3464
rect 2122 3454 2137 3458
rect 2155 3455 2194 3474
rect 2213 3468 2220 3469
rect 2219 3461 2220 3468
rect 2203 3458 2204 3461
rect 2219 3458 2232 3461
rect 2155 3454 2185 3455
rect 2194 3454 2200 3455
rect 2203 3454 2232 3458
rect 2122 3453 2232 3454
rect 2122 3452 2238 3453
rect 1797 3444 1848 3452
rect 1797 3432 1822 3444
rect 1829 3432 1848 3444
rect 1879 3444 1929 3452
rect 1879 3436 1895 3444
rect 1902 3442 1929 3444
rect 1938 3442 2159 3452
rect 1902 3432 2159 3442
rect 2188 3444 2238 3452
rect 2188 3435 2204 3444
rect 1797 3424 1848 3432
rect 1895 3424 2159 3432
rect 2185 3432 2204 3435
rect 2211 3432 2238 3444
rect 2185 3424 2238 3432
rect 1813 3416 1814 3424
rect 1829 3416 1842 3424
rect 1813 3408 1829 3416
rect 1810 3401 1829 3404
rect 1810 3392 1832 3401
rect 1783 3382 1832 3392
rect 1783 3376 1813 3382
rect 1832 3377 1837 3382
rect 1755 3360 1829 3376
rect 1847 3368 1877 3424
rect 1912 3414 2120 3424
rect 2155 3420 2200 3424
rect 2203 3423 2204 3424
rect 2219 3423 2232 3424
rect 1938 3384 2127 3414
rect 1953 3381 2127 3384
rect 1946 3378 2127 3381
rect 1755 3358 1768 3360
rect 1783 3358 1817 3360
rect 1755 3342 1829 3358
rect 1856 3354 1869 3368
rect 1884 3354 1900 3370
rect 1946 3365 1957 3378
rect 1739 3320 1740 3336
rect 1755 3320 1768 3342
rect 1783 3320 1813 3342
rect 1856 3338 1918 3354
rect 1946 3347 1957 3363
rect 1962 3358 1972 3378
rect 1982 3358 1996 3378
rect 1999 3365 2008 3378
rect 2024 3365 2033 3378
rect 1962 3347 1996 3358
rect 1999 3347 2008 3363
rect 2024 3347 2033 3363
rect 2040 3358 2050 3378
rect 2060 3358 2074 3378
rect 2075 3365 2086 3378
rect 2040 3347 2074 3358
rect 2075 3347 2086 3363
rect 2132 3354 2148 3370
rect 2155 3368 2185 3420
rect 2219 3416 2220 3423
rect 2204 3408 2220 3416
rect 2191 3376 2204 3395
rect 2219 3376 2249 3392
rect 2191 3360 2265 3376
rect 2191 3358 2204 3360
rect 2219 3358 2253 3360
rect 1856 3336 1869 3338
rect 1884 3336 1918 3338
rect 1856 3320 1918 3336
rect 1962 3331 1976 3334
rect 2040 3331 2070 3342
rect 2118 3338 2164 3354
rect 2191 3342 2265 3358
rect 2118 3336 2152 3338
rect 2117 3320 2164 3336
rect 2191 3320 2204 3342
rect 2219 3320 2249 3342
rect 2276 3320 2277 3336
rect 2292 3320 2305 3480
rect 2335 3376 2348 3480
rect 2393 3458 2394 3468
rect 2409 3458 2422 3468
rect 2393 3454 2422 3458
rect 2427 3454 2457 3480
rect 2475 3466 2491 3468
rect 2563 3466 2616 3480
rect 2564 3464 2628 3466
rect 2671 3464 2686 3480
rect 2735 3477 2765 3480
rect 2735 3474 2771 3477
rect 2701 3466 2717 3468
rect 2475 3454 2490 3458
rect 2393 3452 2490 3454
rect 2518 3452 2686 3464
rect 2702 3454 2717 3458
rect 2735 3455 2774 3474
rect 2793 3468 2800 3469
rect 2799 3461 2800 3468
rect 2783 3458 2784 3461
rect 2799 3458 2812 3461
rect 2735 3454 2765 3455
rect 2774 3454 2780 3455
rect 2783 3454 2812 3458
rect 2702 3453 2812 3454
rect 2702 3452 2818 3453
rect 2377 3444 2428 3452
rect 2377 3432 2402 3444
rect 2409 3432 2428 3444
rect 2459 3444 2509 3452
rect 2459 3436 2475 3444
rect 2482 3442 2509 3444
rect 2518 3442 2739 3452
rect 2482 3432 2739 3442
rect 2768 3444 2818 3452
rect 2768 3435 2784 3444
rect 2377 3424 2428 3432
rect 2475 3424 2739 3432
rect 2765 3432 2784 3435
rect 2791 3432 2818 3444
rect 2765 3424 2818 3432
rect 2393 3416 2394 3424
rect 2409 3416 2422 3424
rect 2393 3408 2409 3416
rect 2390 3401 2409 3404
rect 2390 3392 2412 3401
rect 2363 3382 2412 3392
rect 2363 3376 2393 3382
rect 2412 3377 2417 3382
rect 2335 3360 2409 3376
rect 2427 3368 2457 3424
rect 2492 3414 2700 3424
rect 2735 3420 2780 3424
rect 2783 3423 2784 3424
rect 2799 3423 2812 3424
rect 2518 3384 2707 3414
rect 2533 3381 2707 3384
rect 2526 3378 2707 3381
rect 2335 3358 2348 3360
rect 2363 3358 2397 3360
rect 2335 3342 2409 3358
rect 2436 3354 2449 3368
rect 2464 3354 2480 3370
rect 2526 3365 2537 3378
rect 2319 3320 2320 3336
rect 2335 3320 2348 3342
rect 2363 3320 2393 3342
rect 2436 3338 2498 3354
rect 2526 3347 2537 3363
rect 2542 3358 2552 3378
rect 2562 3358 2576 3378
rect 2579 3365 2588 3378
rect 2604 3365 2613 3378
rect 2542 3347 2576 3358
rect 2579 3347 2588 3363
rect 2604 3347 2613 3363
rect 2620 3358 2630 3378
rect 2640 3358 2654 3378
rect 2655 3365 2666 3378
rect 2620 3347 2654 3358
rect 2655 3347 2666 3363
rect 2712 3354 2728 3370
rect 2735 3368 2765 3420
rect 2799 3416 2800 3423
rect 2784 3408 2800 3416
rect 2771 3376 2784 3395
rect 2799 3376 2829 3392
rect 2771 3360 2845 3376
rect 2771 3358 2784 3360
rect 2799 3358 2833 3360
rect 2436 3336 2449 3338
rect 2464 3336 2498 3338
rect 2436 3320 2498 3336
rect 2542 3331 2558 3334
rect 2620 3331 2650 3342
rect 2698 3338 2744 3354
rect 2771 3342 2845 3358
rect 2698 3336 2732 3338
rect 2697 3320 2744 3336
rect 2771 3320 2784 3342
rect 2799 3320 2829 3342
rect 2856 3320 2857 3336
rect 2872 3320 2885 3480
rect 2915 3376 2928 3480
rect 2973 3458 2974 3468
rect 2989 3458 3002 3468
rect 2973 3454 3002 3458
rect 3007 3454 3037 3480
rect 3055 3466 3071 3468
rect 3143 3466 3196 3480
rect 3144 3464 3208 3466
rect 3251 3464 3266 3480
rect 3315 3477 3345 3480
rect 3315 3474 3351 3477
rect 3281 3466 3297 3468
rect 3055 3454 3070 3458
rect 2973 3452 3070 3454
rect 3098 3452 3266 3464
rect 3282 3454 3297 3458
rect 3315 3455 3354 3474
rect 3373 3468 3380 3469
rect 3379 3461 3380 3468
rect 3363 3458 3364 3461
rect 3379 3458 3392 3461
rect 3315 3454 3345 3455
rect 3354 3454 3360 3455
rect 3363 3454 3392 3458
rect 3282 3453 3392 3454
rect 3282 3452 3398 3453
rect 2957 3444 3008 3452
rect 2957 3432 2982 3444
rect 2989 3432 3008 3444
rect 3039 3444 3089 3452
rect 3039 3436 3055 3444
rect 3062 3442 3089 3444
rect 3098 3442 3319 3452
rect 3062 3432 3319 3442
rect 3348 3444 3398 3452
rect 3348 3435 3364 3444
rect 2957 3424 3008 3432
rect 3055 3424 3319 3432
rect 3345 3432 3364 3435
rect 3371 3432 3398 3444
rect 3345 3424 3398 3432
rect 2973 3416 2974 3424
rect 2989 3416 3002 3424
rect 2973 3408 2989 3416
rect 2970 3401 2989 3404
rect 2970 3392 2992 3401
rect 2943 3382 2992 3392
rect 2943 3376 2973 3382
rect 2992 3377 2997 3382
rect 2915 3360 2989 3376
rect 3007 3368 3037 3424
rect 3072 3414 3280 3424
rect 3315 3420 3360 3424
rect 3363 3423 3364 3424
rect 3379 3423 3392 3424
rect 3098 3384 3287 3414
rect 3113 3381 3287 3384
rect 3106 3378 3287 3381
rect 2915 3358 2928 3360
rect 2943 3358 2977 3360
rect 2915 3342 2989 3358
rect 3016 3354 3029 3368
rect 3044 3354 3060 3370
rect 3106 3365 3117 3378
rect 2899 3320 2900 3336
rect 2915 3320 2928 3342
rect 2943 3320 2973 3342
rect 3016 3338 3078 3354
rect 3106 3347 3117 3363
rect 3122 3358 3132 3378
rect 3142 3358 3156 3378
rect 3159 3365 3168 3378
rect 3184 3365 3193 3378
rect 3122 3347 3156 3358
rect 3159 3347 3168 3363
rect 3184 3347 3193 3363
rect 3200 3358 3210 3378
rect 3220 3358 3234 3378
rect 3235 3365 3246 3378
rect 3200 3347 3234 3358
rect 3235 3347 3246 3363
rect 3292 3354 3308 3370
rect 3315 3368 3345 3420
rect 3379 3416 3380 3423
rect 3364 3408 3380 3416
rect 3351 3376 3364 3395
rect 3379 3376 3409 3392
rect 3351 3360 3425 3376
rect 3351 3358 3364 3360
rect 3379 3358 3413 3360
rect 3016 3336 3029 3338
rect 3044 3336 3078 3338
rect 3016 3320 3078 3336
rect 3122 3331 3138 3334
rect 3200 3331 3230 3342
rect 3278 3338 3324 3354
rect 3351 3342 3425 3358
rect 3278 3336 3312 3338
rect 3277 3320 3324 3336
rect 3351 3320 3364 3342
rect 3379 3320 3409 3342
rect 3436 3320 3437 3336
rect 3452 3320 3465 3480
rect 3495 3376 3508 3480
rect 3553 3458 3554 3468
rect 3569 3458 3582 3468
rect 3553 3454 3582 3458
rect 3587 3454 3617 3480
rect 3635 3466 3651 3468
rect 3723 3466 3776 3480
rect 3724 3464 3788 3466
rect 3831 3464 3846 3480
rect 3895 3477 3925 3480
rect 3895 3474 3931 3477
rect 3861 3466 3877 3468
rect 3635 3454 3650 3458
rect 3553 3452 3650 3454
rect 3678 3452 3846 3464
rect 3862 3454 3877 3458
rect 3895 3455 3934 3474
rect 3953 3468 3960 3469
rect 3959 3461 3960 3468
rect 3943 3458 3944 3461
rect 3959 3458 3972 3461
rect 3895 3454 3925 3455
rect 3934 3454 3940 3455
rect 3943 3454 3972 3458
rect 3862 3453 3972 3454
rect 3862 3452 3978 3453
rect 3537 3444 3588 3452
rect 3537 3432 3562 3444
rect 3569 3432 3588 3444
rect 3619 3444 3669 3452
rect 3619 3436 3635 3444
rect 3642 3442 3669 3444
rect 3678 3442 3899 3452
rect 3642 3432 3899 3442
rect 3928 3444 3978 3452
rect 3928 3435 3944 3444
rect 3537 3424 3588 3432
rect 3635 3424 3899 3432
rect 3925 3432 3944 3435
rect 3951 3432 3978 3444
rect 3925 3424 3978 3432
rect 3553 3416 3554 3424
rect 3569 3416 3582 3424
rect 3553 3408 3569 3416
rect 3550 3401 3569 3404
rect 3550 3392 3572 3401
rect 3523 3382 3572 3392
rect 3523 3376 3553 3382
rect 3572 3377 3577 3382
rect 3495 3360 3569 3376
rect 3587 3368 3617 3424
rect 3652 3414 3860 3424
rect 3895 3420 3940 3424
rect 3943 3423 3944 3424
rect 3959 3423 3972 3424
rect 3678 3384 3867 3414
rect 3693 3381 3867 3384
rect 3686 3378 3867 3381
rect 3495 3358 3508 3360
rect 3523 3358 3557 3360
rect 3495 3342 3569 3358
rect 3596 3354 3609 3368
rect 3624 3354 3640 3370
rect 3686 3365 3697 3378
rect 3479 3320 3480 3336
rect 3495 3320 3508 3342
rect 3523 3320 3553 3342
rect 3596 3338 3658 3354
rect 3686 3347 3697 3363
rect 3702 3358 3712 3378
rect 3722 3358 3736 3378
rect 3739 3365 3748 3378
rect 3764 3365 3773 3378
rect 3702 3347 3736 3358
rect 3739 3347 3748 3363
rect 3764 3347 3773 3363
rect 3780 3358 3790 3378
rect 3800 3358 3814 3378
rect 3815 3365 3826 3378
rect 3780 3347 3814 3358
rect 3815 3347 3826 3363
rect 3872 3354 3888 3370
rect 3895 3368 3925 3420
rect 3959 3416 3960 3423
rect 3944 3408 3960 3416
rect 3931 3376 3944 3395
rect 3959 3376 3989 3392
rect 3931 3360 4005 3376
rect 3931 3358 3944 3360
rect 3959 3358 3993 3360
rect 3596 3336 3609 3338
rect 3624 3336 3658 3338
rect 3596 3320 3658 3336
rect 3702 3331 3718 3334
rect 3780 3331 3810 3342
rect 3858 3338 3904 3354
rect 3931 3342 4005 3358
rect 3858 3336 3892 3338
rect 3857 3320 3904 3336
rect 3931 3320 3944 3342
rect 3959 3320 3989 3342
rect 4016 3320 4017 3336
rect 4032 3320 4045 3480
rect 4075 3376 4088 3480
rect 4133 3458 4134 3468
rect 4149 3458 4162 3468
rect 4133 3454 4162 3458
rect 4167 3454 4197 3480
rect 4215 3466 4231 3468
rect 4303 3466 4356 3480
rect 4304 3464 4368 3466
rect 4411 3464 4426 3480
rect 4475 3477 4505 3480
rect 4475 3474 4511 3477
rect 4441 3466 4457 3468
rect 4215 3454 4230 3458
rect 4133 3452 4230 3454
rect 4258 3452 4426 3464
rect 4442 3454 4457 3458
rect 4475 3455 4514 3474
rect 4533 3468 4540 3469
rect 4539 3461 4540 3468
rect 4523 3458 4524 3461
rect 4539 3458 4552 3461
rect 4475 3454 4505 3455
rect 4514 3454 4520 3455
rect 4523 3454 4552 3458
rect 4442 3453 4552 3454
rect 4442 3452 4558 3453
rect 4117 3444 4168 3452
rect 4117 3432 4142 3444
rect 4149 3432 4168 3444
rect 4199 3444 4249 3452
rect 4199 3436 4215 3444
rect 4222 3442 4249 3444
rect 4258 3442 4479 3452
rect 4222 3432 4479 3442
rect 4508 3444 4558 3452
rect 4508 3435 4524 3444
rect 4117 3424 4168 3432
rect 4215 3424 4479 3432
rect 4505 3432 4524 3435
rect 4531 3432 4558 3444
rect 4505 3424 4558 3432
rect 4133 3416 4134 3424
rect 4149 3416 4162 3424
rect 4133 3408 4149 3416
rect 4130 3401 4149 3404
rect 4130 3392 4152 3401
rect 4103 3382 4152 3392
rect 4103 3376 4133 3382
rect 4152 3377 4157 3382
rect 4075 3360 4149 3376
rect 4167 3368 4197 3424
rect 4232 3414 4440 3424
rect 4475 3420 4520 3424
rect 4523 3423 4524 3424
rect 4539 3423 4552 3424
rect 4258 3384 4447 3414
rect 4273 3381 4447 3384
rect 4266 3378 4447 3381
rect 4075 3358 4088 3360
rect 4103 3358 4137 3360
rect 4075 3342 4149 3358
rect 4176 3354 4189 3368
rect 4204 3354 4220 3370
rect 4266 3365 4277 3378
rect 4059 3320 4060 3336
rect 4075 3320 4088 3342
rect 4103 3320 4133 3342
rect 4176 3338 4238 3354
rect 4266 3347 4277 3363
rect 4282 3358 4292 3378
rect 4302 3358 4316 3378
rect 4319 3365 4328 3378
rect 4344 3365 4353 3378
rect 4282 3347 4316 3358
rect 4319 3347 4328 3363
rect 4344 3347 4353 3363
rect 4360 3358 4370 3378
rect 4380 3358 4394 3378
rect 4395 3365 4406 3378
rect 4360 3347 4394 3358
rect 4395 3347 4406 3363
rect 4452 3354 4468 3370
rect 4475 3368 4505 3420
rect 4539 3416 4540 3423
rect 4524 3408 4540 3416
rect 4511 3376 4524 3395
rect 4539 3376 4569 3392
rect 4511 3360 4585 3376
rect 4511 3358 4524 3360
rect 4539 3358 4573 3360
rect 4176 3336 4189 3338
rect 4204 3336 4238 3338
rect 4176 3320 4238 3336
rect 4282 3331 4298 3334
rect 4360 3331 4390 3342
rect 4438 3338 4484 3354
rect 4511 3342 4585 3358
rect 4438 3336 4472 3338
rect 4437 3320 4484 3336
rect 4511 3320 4524 3342
rect 4539 3320 4569 3342
rect 4596 3320 4597 3336
rect 4612 3320 4625 3480
rect 4655 3376 4668 3480
rect 4713 3458 4714 3468
rect 4729 3458 4742 3468
rect 4713 3454 4742 3458
rect 4747 3454 4777 3480
rect 4795 3466 4811 3468
rect 4883 3466 4936 3480
rect 4884 3464 4948 3466
rect 4991 3464 5006 3480
rect 5055 3477 5085 3480
rect 5055 3474 5091 3477
rect 5021 3466 5037 3468
rect 4795 3454 4810 3458
rect 4713 3452 4810 3454
rect 4838 3452 5006 3464
rect 5022 3454 5037 3458
rect 5055 3455 5094 3474
rect 5113 3468 5120 3469
rect 5119 3461 5120 3468
rect 5103 3458 5104 3461
rect 5119 3458 5132 3461
rect 5055 3454 5085 3455
rect 5094 3454 5100 3455
rect 5103 3454 5132 3458
rect 5022 3453 5132 3454
rect 5022 3452 5138 3453
rect 4697 3444 4748 3452
rect 4697 3432 4722 3444
rect 4729 3432 4748 3444
rect 4779 3444 4829 3452
rect 4779 3436 4795 3444
rect 4802 3442 4829 3444
rect 4838 3442 5059 3452
rect 4802 3432 5059 3442
rect 5088 3444 5138 3452
rect 5088 3435 5104 3444
rect 4697 3424 4748 3432
rect 4795 3424 5059 3432
rect 5085 3432 5104 3435
rect 5111 3432 5138 3444
rect 5085 3424 5138 3432
rect 4713 3416 4714 3424
rect 4729 3416 4742 3424
rect 4713 3408 4729 3416
rect 4710 3401 4729 3404
rect 4710 3392 4732 3401
rect 4683 3382 4732 3392
rect 4683 3376 4713 3382
rect 4732 3377 4737 3382
rect 4655 3360 4729 3376
rect 4747 3368 4777 3424
rect 4812 3414 5020 3424
rect 5055 3420 5100 3424
rect 5103 3423 5104 3424
rect 5119 3423 5132 3424
rect 4838 3384 5027 3414
rect 4853 3381 5027 3384
rect 4846 3378 5027 3381
rect 4655 3358 4668 3360
rect 4683 3358 4717 3360
rect 4655 3342 4729 3358
rect 4756 3354 4769 3368
rect 4784 3354 4800 3370
rect 4846 3365 4857 3378
rect 4639 3320 4640 3336
rect 4655 3320 4668 3342
rect 4683 3320 4713 3342
rect 4756 3338 4818 3354
rect 4846 3347 4857 3363
rect 4862 3358 4872 3378
rect 4882 3358 4896 3378
rect 4899 3365 4908 3378
rect 4924 3365 4933 3378
rect 4862 3347 4896 3358
rect 4899 3347 4908 3363
rect 4924 3347 4933 3363
rect 4940 3358 4950 3378
rect 4960 3358 4974 3378
rect 4975 3365 4986 3378
rect 4940 3347 4974 3358
rect 4975 3347 4986 3363
rect 5032 3354 5048 3370
rect 5055 3368 5085 3420
rect 5119 3416 5120 3423
rect 5104 3408 5120 3416
rect 5091 3376 5104 3395
rect 5119 3376 5149 3392
rect 5091 3360 5165 3376
rect 5091 3358 5104 3360
rect 5119 3358 5153 3360
rect 4756 3336 4769 3338
rect 4784 3336 4818 3338
rect 4756 3320 4818 3336
rect 4862 3331 4878 3334
rect 4940 3331 4970 3342
rect 5018 3338 5064 3354
rect 5091 3342 5165 3358
rect 5018 3336 5052 3338
rect 5017 3320 5064 3336
rect 5091 3320 5104 3342
rect 5119 3320 5149 3342
rect 5176 3320 5177 3336
rect 5192 3320 5205 3480
rect 5235 3376 5248 3480
rect 5293 3458 5294 3468
rect 5309 3458 5322 3468
rect 5293 3454 5322 3458
rect 5327 3454 5357 3480
rect 5375 3466 5391 3468
rect 5463 3466 5516 3480
rect 5464 3464 5528 3466
rect 5571 3464 5586 3480
rect 5635 3477 5665 3480
rect 5635 3474 5671 3477
rect 5601 3466 5617 3468
rect 5375 3454 5390 3458
rect 5293 3452 5390 3454
rect 5418 3452 5586 3464
rect 5602 3454 5617 3458
rect 5635 3455 5674 3474
rect 5693 3468 5700 3469
rect 5699 3461 5700 3468
rect 5683 3458 5684 3461
rect 5699 3458 5712 3461
rect 5635 3454 5665 3455
rect 5674 3454 5680 3455
rect 5683 3454 5712 3458
rect 5602 3453 5712 3454
rect 5602 3452 5718 3453
rect 5277 3444 5328 3452
rect 5277 3432 5302 3444
rect 5309 3432 5328 3444
rect 5359 3444 5409 3452
rect 5359 3436 5375 3444
rect 5382 3442 5409 3444
rect 5418 3442 5639 3452
rect 5382 3432 5639 3442
rect 5668 3444 5718 3452
rect 5668 3435 5684 3444
rect 5277 3424 5328 3432
rect 5375 3424 5639 3432
rect 5665 3432 5684 3435
rect 5691 3432 5718 3444
rect 5665 3424 5718 3432
rect 5293 3416 5294 3424
rect 5309 3416 5322 3424
rect 5293 3408 5309 3416
rect 5290 3401 5309 3404
rect 5290 3392 5312 3401
rect 5263 3382 5312 3392
rect 5263 3376 5293 3382
rect 5312 3377 5317 3382
rect 5235 3360 5309 3376
rect 5327 3368 5357 3424
rect 5392 3414 5600 3424
rect 5635 3420 5680 3424
rect 5683 3423 5684 3424
rect 5699 3423 5712 3424
rect 5418 3384 5607 3414
rect 5433 3381 5607 3384
rect 5426 3378 5607 3381
rect 5235 3358 5248 3360
rect 5263 3358 5297 3360
rect 5235 3342 5309 3358
rect 5336 3354 5349 3368
rect 5364 3354 5380 3370
rect 5426 3365 5437 3378
rect 5219 3320 5220 3336
rect 5235 3320 5248 3342
rect 5263 3320 5293 3342
rect 5336 3338 5398 3354
rect 5426 3347 5437 3363
rect 5442 3358 5452 3378
rect 5462 3358 5476 3378
rect 5479 3365 5488 3378
rect 5504 3365 5513 3378
rect 5442 3347 5476 3358
rect 5479 3347 5488 3363
rect 5504 3347 5513 3363
rect 5520 3358 5530 3378
rect 5540 3358 5554 3378
rect 5555 3365 5566 3378
rect 5520 3347 5554 3358
rect 5555 3347 5566 3363
rect 5612 3354 5628 3370
rect 5635 3368 5665 3420
rect 5699 3416 5700 3423
rect 5684 3408 5700 3416
rect 5671 3376 5684 3395
rect 5699 3376 5729 3392
rect 5671 3360 5745 3376
rect 5671 3358 5684 3360
rect 5699 3358 5733 3360
rect 5336 3336 5349 3338
rect 5364 3336 5398 3338
rect 5336 3320 5398 3336
rect 5442 3331 5458 3334
rect 5520 3331 5550 3342
rect 5598 3338 5644 3354
rect 5671 3342 5745 3358
rect 5598 3336 5632 3338
rect 5597 3320 5644 3336
rect 5671 3320 5684 3342
rect 5699 3320 5729 3342
rect 5756 3320 5757 3336
rect 5772 3320 5785 3480
rect 5815 3376 5828 3480
rect 5873 3458 5874 3468
rect 5889 3458 5902 3468
rect 5873 3454 5902 3458
rect 5907 3454 5937 3480
rect 5955 3466 5971 3468
rect 6043 3466 6096 3480
rect 6044 3464 6108 3466
rect 6151 3464 6166 3480
rect 6215 3477 6245 3480
rect 6215 3474 6251 3477
rect 6181 3466 6197 3468
rect 5955 3454 5970 3458
rect 5873 3452 5970 3454
rect 5998 3452 6166 3464
rect 6182 3454 6197 3458
rect 6215 3455 6254 3474
rect 6273 3468 6280 3469
rect 6279 3461 6280 3468
rect 6263 3458 6264 3461
rect 6279 3458 6292 3461
rect 6215 3454 6245 3455
rect 6254 3454 6260 3455
rect 6263 3454 6292 3458
rect 6182 3453 6292 3454
rect 6182 3452 6298 3453
rect 5857 3444 5908 3452
rect 5857 3432 5882 3444
rect 5889 3432 5908 3444
rect 5939 3444 5989 3452
rect 5939 3436 5955 3444
rect 5962 3442 5989 3444
rect 5998 3442 6219 3452
rect 5962 3432 6219 3442
rect 6248 3444 6298 3452
rect 6248 3435 6264 3444
rect 5857 3424 5908 3432
rect 5955 3424 6219 3432
rect 6245 3432 6264 3435
rect 6271 3432 6298 3444
rect 6245 3424 6298 3432
rect 5873 3416 5874 3424
rect 5889 3416 5902 3424
rect 5873 3408 5889 3416
rect 5870 3401 5889 3404
rect 5870 3392 5892 3401
rect 5843 3382 5892 3392
rect 5843 3376 5873 3382
rect 5892 3377 5897 3382
rect 5815 3360 5889 3376
rect 5907 3368 5937 3424
rect 5972 3414 6180 3424
rect 6215 3420 6260 3424
rect 6263 3423 6264 3424
rect 6279 3423 6292 3424
rect 5998 3384 6187 3414
rect 6013 3381 6187 3384
rect 6006 3378 6187 3381
rect 5815 3358 5828 3360
rect 5843 3358 5877 3360
rect 5815 3342 5889 3358
rect 5916 3354 5929 3368
rect 5944 3354 5960 3370
rect 6006 3365 6017 3378
rect 5799 3320 5800 3336
rect 5815 3320 5828 3342
rect 5843 3320 5873 3342
rect 5916 3338 5978 3354
rect 6006 3347 6017 3363
rect 6022 3358 6032 3378
rect 6042 3358 6056 3378
rect 6059 3365 6068 3378
rect 6084 3365 6093 3378
rect 6022 3347 6056 3358
rect 6059 3347 6068 3363
rect 6084 3347 6093 3363
rect 6100 3358 6110 3378
rect 6120 3358 6134 3378
rect 6135 3365 6146 3378
rect 6100 3347 6134 3358
rect 6135 3347 6146 3363
rect 6192 3354 6208 3370
rect 6215 3368 6245 3420
rect 6279 3416 6280 3423
rect 6264 3408 6280 3416
rect 6251 3376 6264 3395
rect 6279 3376 6309 3392
rect 6251 3360 6325 3376
rect 6251 3358 6264 3360
rect 6279 3358 6313 3360
rect 5916 3336 5929 3338
rect 5944 3336 5978 3338
rect 5916 3320 5978 3336
rect 6022 3331 6038 3334
rect 6100 3331 6130 3342
rect 6178 3338 6224 3354
rect 6251 3342 6325 3358
rect 6178 3336 6212 3338
rect 6177 3320 6224 3336
rect 6251 3320 6264 3342
rect 6279 3320 6309 3342
rect 6336 3320 6337 3336
rect 6352 3320 6365 3480
rect 6395 3376 6408 3480
rect 6453 3458 6454 3468
rect 6469 3458 6482 3468
rect 6453 3454 6482 3458
rect 6487 3454 6517 3480
rect 6535 3466 6551 3468
rect 6623 3466 6676 3480
rect 6624 3464 6688 3466
rect 6731 3464 6746 3480
rect 6795 3477 6825 3480
rect 6795 3474 6831 3477
rect 6761 3466 6777 3468
rect 6535 3454 6550 3458
rect 6453 3452 6550 3454
rect 6578 3452 6746 3464
rect 6762 3454 6777 3458
rect 6795 3455 6834 3474
rect 6853 3468 6860 3469
rect 6859 3461 6860 3468
rect 6843 3458 6844 3461
rect 6859 3458 6872 3461
rect 6795 3454 6825 3455
rect 6834 3454 6840 3455
rect 6843 3454 6872 3458
rect 6762 3453 6872 3454
rect 6762 3452 6878 3453
rect 6437 3444 6488 3452
rect 6437 3432 6462 3444
rect 6469 3432 6488 3444
rect 6519 3444 6569 3452
rect 6519 3436 6535 3444
rect 6542 3442 6569 3444
rect 6578 3442 6799 3452
rect 6542 3432 6799 3442
rect 6828 3444 6878 3452
rect 6828 3435 6844 3444
rect 6437 3424 6488 3432
rect 6535 3424 6799 3432
rect 6825 3432 6844 3435
rect 6851 3432 6878 3444
rect 6825 3424 6878 3432
rect 6453 3416 6454 3424
rect 6469 3416 6482 3424
rect 6453 3408 6469 3416
rect 6450 3401 6469 3404
rect 6450 3392 6472 3401
rect 6423 3382 6472 3392
rect 6423 3376 6453 3382
rect 6472 3377 6477 3382
rect 6395 3360 6469 3376
rect 6487 3368 6517 3424
rect 6552 3414 6760 3424
rect 6795 3420 6840 3424
rect 6843 3423 6844 3424
rect 6859 3423 6872 3424
rect 6578 3384 6767 3414
rect 6593 3381 6767 3384
rect 6586 3378 6767 3381
rect 6395 3358 6408 3360
rect 6423 3358 6457 3360
rect 6395 3342 6469 3358
rect 6496 3354 6509 3368
rect 6524 3354 6540 3370
rect 6586 3365 6597 3378
rect 6379 3320 6380 3336
rect 6395 3320 6408 3342
rect 6423 3320 6453 3342
rect 6496 3338 6558 3354
rect 6586 3347 6597 3363
rect 6602 3358 6612 3378
rect 6622 3358 6636 3378
rect 6639 3365 6648 3378
rect 6664 3365 6673 3378
rect 6602 3347 6636 3358
rect 6639 3347 6648 3363
rect 6664 3347 6673 3363
rect 6680 3358 6690 3378
rect 6700 3358 6714 3378
rect 6715 3365 6726 3378
rect 6680 3347 6714 3358
rect 6715 3347 6726 3363
rect 6772 3354 6788 3370
rect 6795 3368 6825 3420
rect 6859 3416 6860 3423
rect 6844 3408 6860 3416
rect 6831 3376 6844 3395
rect 6859 3376 6889 3392
rect 6831 3360 6905 3376
rect 6831 3358 6844 3360
rect 6859 3358 6893 3360
rect 6496 3336 6509 3338
rect 6524 3336 6558 3338
rect 6496 3320 6558 3336
rect 6602 3331 6618 3334
rect 6680 3331 6710 3342
rect 6758 3338 6804 3354
rect 6831 3342 6905 3358
rect 6758 3336 6792 3338
rect 6757 3320 6804 3336
rect 6831 3320 6844 3342
rect 6859 3320 6889 3342
rect 6916 3320 6917 3336
rect 6932 3320 6945 3480
rect 6975 3376 6988 3480
rect 7033 3458 7034 3468
rect 7049 3458 7062 3468
rect 7033 3454 7062 3458
rect 7067 3454 7097 3480
rect 7115 3466 7131 3468
rect 7203 3466 7256 3480
rect 7204 3464 7268 3466
rect 7311 3464 7326 3480
rect 7375 3477 7405 3480
rect 7375 3474 7411 3477
rect 7341 3466 7357 3468
rect 7115 3454 7130 3458
rect 7033 3452 7130 3454
rect 7158 3452 7326 3464
rect 7342 3454 7357 3458
rect 7375 3455 7414 3474
rect 7433 3468 7440 3469
rect 7439 3461 7440 3468
rect 7423 3458 7424 3461
rect 7439 3458 7452 3461
rect 7375 3454 7405 3455
rect 7414 3454 7420 3455
rect 7423 3454 7452 3458
rect 7342 3453 7452 3454
rect 7342 3452 7458 3453
rect 7017 3444 7068 3452
rect 7017 3432 7042 3444
rect 7049 3432 7068 3444
rect 7099 3444 7149 3452
rect 7099 3436 7115 3444
rect 7122 3442 7149 3444
rect 7158 3442 7379 3452
rect 7122 3432 7379 3442
rect 7408 3444 7458 3452
rect 7408 3435 7424 3444
rect 7017 3424 7068 3432
rect 7115 3424 7379 3432
rect 7405 3432 7424 3435
rect 7431 3432 7458 3444
rect 7405 3424 7458 3432
rect 7033 3416 7034 3424
rect 7049 3416 7062 3424
rect 7033 3408 7049 3416
rect 7030 3401 7049 3404
rect 7030 3392 7052 3401
rect 7003 3382 7052 3392
rect 7003 3376 7033 3382
rect 7052 3377 7057 3382
rect 6975 3360 7049 3376
rect 7067 3368 7097 3424
rect 7132 3414 7340 3424
rect 7375 3420 7420 3424
rect 7423 3423 7424 3424
rect 7439 3423 7452 3424
rect 7158 3384 7347 3414
rect 7173 3381 7347 3384
rect 7166 3378 7347 3381
rect 6975 3358 6988 3360
rect 7003 3358 7037 3360
rect 6975 3342 7049 3358
rect 7076 3354 7089 3368
rect 7104 3354 7120 3370
rect 7166 3365 7177 3378
rect 6959 3320 6960 3336
rect 6975 3320 6988 3342
rect 7003 3320 7033 3342
rect 7076 3338 7138 3354
rect 7166 3347 7177 3363
rect 7182 3358 7192 3378
rect 7202 3358 7216 3378
rect 7219 3365 7228 3378
rect 7244 3365 7253 3378
rect 7182 3347 7216 3358
rect 7219 3347 7228 3363
rect 7244 3347 7253 3363
rect 7260 3358 7270 3378
rect 7280 3358 7294 3378
rect 7295 3365 7306 3378
rect 7260 3347 7294 3358
rect 7295 3347 7306 3363
rect 7352 3354 7368 3370
rect 7375 3368 7405 3420
rect 7439 3416 7440 3423
rect 7424 3408 7440 3416
rect 7411 3376 7424 3395
rect 7439 3376 7469 3392
rect 7411 3360 7485 3376
rect 7411 3358 7424 3360
rect 7439 3358 7473 3360
rect 7076 3336 7089 3338
rect 7104 3336 7138 3338
rect 7076 3320 7138 3336
rect 7182 3331 7198 3334
rect 7260 3331 7290 3342
rect 7338 3338 7384 3354
rect 7411 3342 7485 3358
rect 7338 3336 7372 3338
rect 7337 3320 7384 3336
rect 7411 3320 7424 3342
rect 7439 3320 7469 3342
rect 7496 3320 7497 3336
rect 7512 3320 7525 3480
rect 7555 3376 7568 3480
rect 7613 3458 7614 3468
rect 7629 3458 7642 3468
rect 7613 3454 7642 3458
rect 7647 3454 7677 3480
rect 7695 3466 7711 3468
rect 7783 3466 7836 3480
rect 7784 3464 7848 3466
rect 7891 3464 7906 3480
rect 7955 3477 7985 3480
rect 7955 3474 7991 3477
rect 7921 3466 7937 3468
rect 7695 3454 7710 3458
rect 7613 3452 7710 3454
rect 7738 3452 7906 3464
rect 7922 3454 7937 3458
rect 7955 3455 7994 3474
rect 8013 3468 8020 3469
rect 8019 3461 8020 3468
rect 8003 3458 8004 3461
rect 8019 3458 8032 3461
rect 7955 3454 7985 3455
rect 7994 3454 8000 3455
rect 8003 3454 8032 3458
rect 7922 3453 8032 3454
rect 7922 3452 8038 3453
rect 7597 3444 7648 3452
rect 7597 3432 7622 3444
rect 7629 3432 7648 3444
rect 7679 3444 7729 3452
rect 7679 3436 7695 3444
rect 7702 3442 7729 3444
rect 7738 3442 7959 3452
rect 7702 3432 7959 3442
rect 7988 3444 8038 3452
rect 7988 3435 8004 3444
rect 7597 3424 7648 3432
rect 7695 3424 7959 3432
rect 7985 3432 8004 3435
rect 8011 3432 8038 3444
rect 7985 3424 8038 3432
rect 7613 3416 7614 3424
rect 7629 3416 7642 3424
rect 7613 3408 7629 3416
rect 7610 3401 7629 3404
rect 7610 3392 7632 3401
rect 7583 3382 7632 3392
rect 7583 3376 7613 3382
rect 7632 3377 7637 3382
rect 7555 3360 7629 3376
rect 7647 3368 7677 3424
rect 7712 3414 7920 3424
rect 7955 3420 8000 3424
rect 8003 3423 8004 3424
rect 8019 3423 8032 3424
rect 7738 3384 7927 3414
rect 7753 3381 7927 3384
rect 7746 3378 7927 3381
rect 7555 3358 7568 3360
rect 7583 3358 7617 3360
rect 7555 3342 7629 3358
rect 7656 3354 7669 3368
rect 7684 3354 7700 3370
rect 7746 3365 7757 3378
rect 7539 3320 7540 3336
rect 7555 3320 7568 3342
rect 7583 3320 7613 3342
rect 7656 3338 7718 3354
rect 7746 3347 7757 3363
rect 7762 3358 7772 3378
rect 7782 3358 7796 3378
rect 7799 3365 7808 3378
rect 7824 3365 7833 3378
rect 7762 3347 7796 3358
rect 7799 3347 7808 3363
rect 7824 3347 7833 3363
rect 7840 3358 7850 3378
rect 7860 3358 7874 3378
rect 7875 3365 7886 3378
rect 7840 3347 7874 3358
rect 7875 3347 7886 3363
rect 7932 3354 7948 3370
rect 7955 3368 7985 3420
rect 8019 3416 8020 3423
rect 8004 3408 8020 3416
rect 7991 3376 8004 3395
rect 8019 3376 8049 3392
rect 7991 3360 8065 3376
rect 7991 3358 8004 3360
rect 8019 3358 8053 3360
rect 7656 3336 7669 3338
rect 7684 3336 7718 3338
rect 7656 3320 7718 3336
rect 7762 3331 7778 3334
rect 7840 3331 7870 3342
rect 7918 3338 7964 3354
rect 7991 3342 8065 3358
rect 7918 3336 7952 3338
rect 7917 3320 7964 3336
rect 7991 3320 8004 3342
rect 8019 3320 8049 3342
rect 8076 3320 8077 3336
rect 8092 3320 8105 3480
rect 8135 3376 8148 3480
rect 8193 3458 8194 3468
rect 8209 3458 8222 3468
rect 8193 3454 8222 3458
rect 8227 3454 8257 3480
rect 8275 3466 8291 3468
rect 8363 3466 8416 3480
rect 8364 3464 8428 3466
rect 8471 3464 8486 3480
rect 8535 3477 8565 3480
rect 8535 3474 8571 3477
rect 8501 3466 8517 3468
rect 8275 3454 8290 3458
rect 8193 3452 8290 3454
rect 8318 3452 8486 3464
rect 8502 3454 8517 3458
rect 8535 3455 8574 3474
rect 8593 3468 8600 3469
rect 8599 3461 8600 3468
rect 8583 3458 8584 3461
rect 8599 3458 8612 3461
rect 8535 3454 8565 3455
rect 8574 3454 8580 3455
rect 8583 3454 8612 3458
rect 8502 3453 8612 3454
rect 8502 3452 8618 3453
rect 8177 3444 8228 3452
rect 8177 3432 8202 3444
rect 8209 3432 8228 3444
rect 8259 3444 8309 3452
rect 8259 3436 8275 3444
rect 8282 3442 8309 3444
rect 8318 3442 8539 3452
rect 8282 3432 8539 3442
rect 8568 3444 8618 3452
rect 8568 3435 8584 3444
rect 8177 3424 8228 3432
rect 8275 3424 8539 3432
rect 8565 3432 8584 3435
rect 8591 3432 8618 3444
rect 8565 3424 8618 3432
rect 8193 3416 8194 3424
rect 8209 3416 8222 3424
rect 8193 3408 8209 3416
rect 8190 3401 8209 3404
rect 8190 3392 8212 3401
rect 8163 3382 8212 3392
rect 8163 3376 8193 3382
rect 8212 3377 8217 3382
rect 8135 3360 8209 3376
rect 8227 3368 8257 3424
rect 8292 3414 8500 3424
rect 8535 3420 8580 3424
rect 8583 3423 8584 3424
rect 8599 3423 8612 3424
rect 8318 3384 8507 3414
rect 8333 3381 8507 3384
rect 8326 3378 8507 3381
rect 8135 3358 8148 3360
rect 8163 3358 8197 3360
rect 8135 3342 8209 3358
rect 8236 3354 8249 3368
rect 8264 3354 8280 3370
rect 8326 3365 8337 3378
rect 8119 3320 8120 3336
rect 8135 3320 8148 3342
rect 8163 3320 8193 3342
rect 8236 3338 8298 3354
rect 8326 3347 8337 3363
rect 8342 3358 8352 3378
rect 8362 3358 8376 3378
rect 8379 3365 8388 3378
rect 8404 3365 8413 3378
rect 8342 3347 8376 3358
rect 8379 3347 8388 3363
rect 8404 3347 8413 3363
rect 8420 3358 8430 3378
rect 8440 3358 8454 3378
rect 8455 3365 8466 3378
rect 8420 3347 8454 3358
rect 8455 3347 8466 3363
rect 8512 3354 8528 3370
rect 8535 3368 8565 3420
rect 8599 3416 8600 3423
rect 8584 3408 8600 3416
rect 8571 3376 8584 3395
rect 8599 3376 8629 3392
rect 8571 3360 8645 3376
rect 8571 3358 8584 3360
rect 8599 3358 8633 3360
rect 8236 3336 8249 3338
rect 8264 3336 8298 3338
rect 8236 3320 8298 3336
rect 8342 3331 8358 3334
rect 8420 3331 8450 3342
rect 8498 3338 8544 3354
rect 8571 3342 8645 3358
rect 8498 3336 8532 3338
rect 8497 3320 8544 3336
rect 8571 3320 8584 3342
rect 8599 3320 8629 3342
rect 8656 3320 8657 3336
rect 8672 3320 8685 3480
rect 8715 3376 8728 3480
rect 8773 3458 8774 3468
rect 8789 3458 8802 3468
rect 8773 3454 8802 3458
rect 8807 3454 8837 3480
rect 8855 3466 8871 3468
rect 8943 3466 8996 3480
rect 8944 3464 9008 3466
rect 9051 3464 9066 3480
rect 9115 3477 9145 3480
rect 9115 3474 9151 3477
rect 9081 3466 9097 3468
rect 8855 3454 8870 3458
rect 8773 3452 8870 3454
rect 8898 3452 9066 3464
rect 9082 3454 9097 3458
rect 9115 3455 9154 3474
rect 9173 3468 9180 3469
rect 9179 3461 9180 3468
rect 9163 3458 9164 3461
rect 9179 3458 9192 3461
rect 9115 3454 9145 3455
rect 9154 3454 9160 3455
rect 9163 3454 9192 3458
rect 9082 3453 9192 3454
rect 9082 3452 9198 3453
rect 8757 3444 8808 3452
rect 8757 3432 8782 3444
rect 8789 3432 8808 3444
rect 8839 3444 8889 3452
rect 8839 3436 8855 3444
rect 8862 3442 8889 3444
rect 8898 3442 9119 3452
rect 8862 3432 9119 3442
rect 9148 3444 9198 3452
rect 9148 3435 9164 3444
rect 8757 3424 8808 3432
rect 8855 3424 9119 3432
rect 9145 3432 9164 3435
rect 9171 3432 9198 3444
rect 9145 3424 9198 3432
rect 8773 3416 8774 3424
rect 8789 3416 8802 3424
rect 8773 3408 8789 3416
rect 8770 3401 8789 3404
rect 8770 3392 8792 3401
rect 8743 3382 8792 3392
rect 8743 3376 8773 3382
rect 8792 3377 8797 3382
rect 8715 3360 8789 3376
rect 8807 3368 8837 3424
rect 8872 3414 9080 3424
rect 9115 3420 9160 3424
rect 9163 3423 9164 3424
rect 9179 3423 9192 3424
rect 8898 3384 9087 3414
rect 8913 3381 9087 3384
rect 8906 3378 9087 3381
rect 8715 3358 8728 3360
rect 8743 3358 8777 3360
rect 8715 3342 8789 3358
rect 8816 3354 8829 3368
rect 8844 3354 8860 3370
rect 8906 3365 8917 3378
rect 8699 3320 8700 3336
rect 8715 3320 8728 3342
rect 8743 3320 8773 3342
rect 8816 3338 8878 3354
rect 8906 3347 8917 3363
rect 8922 3358 8932 3378
rect 8942 3358 8956 3378
rect 8959 3365 8968 3378
rect 8984 3365 8993 3378
rect 8922 3347 8956 3358
rect 8959 3347 8968 3363
rect 8984 3347 8993 3363
rect 9000 3358 9010 3378
rect 9020 3358 9034 3378
rect 9035 3365 9046 3378
rect 9000 3347 9034 3358
rect 9035 3347 9046 3363
rect 9092 3354 9108 3370
rect 9115 3368 9145 3420
rect 9179 3416 9180 3423
rect 9164 3408 9180 3416
rect 9151 3376 9164 3395
rect 9179 3376 9209 3392
rect 9151 3360 9225 3376
rect 9151 3358 9164 3360
rect 9179 3358 9213 3360
rect 8816 3336 8829 3338
rect 8844 3336 8878 3338
rect 8816 3320 8878 3336
rect 8922 3331 8938 3334
rect 9000 3331 9030 3342
rect 9078 3338 9124 3354
rect 9151 3342 9225 3358
rect 9078 3336 9112 3338
rect 9077 3320 9124 3336
rect 9151 3320 9164 3342
rect 9179 3320 9209 3342
rect 9236 3320 9237 3336
rect 9252 3320 9265 3480
rect -7 3312 34 3320
rect -7 3286 8 3312
rect 15 3286 34 3312
rect 98 3308 160 3320
rect 172 3308 247 3320
rect 305 3308 380 3320
rect 392 3308 423 3320
rect 429 3308 464 3320
rect 98 3306 260 3308
rect -7 3278 34 3286
rect 116 3282 129 3306
rect 144 3304 159 3306
rect -1 3268 0 3278
rect 15 3268 28 3278
rect 43 3268 73 3282
rect 116 3268 159 3282
rect 183 3279 190 3286
rect 193 3282 260 3306
rect 292 3306 464 3308
rect 262 3284 290 3288
rect 292 3284 372 3306
rect 393 3304 408 3306
rect 262 3282 372 3284
rect 193 3278 372 3282
rect 166 3268 196 3278
rect 198 3268 351 3278
rect 359 3268 389 3278
rect 393 3268 423 3282
rect 451 3268 464 3306
rect 536 3312 571 3320
rect 536 3286 537 3312
rect 544 3286 571 3312
rect 479 3268 509 3282
rect 536 3278 571 3286
rect 573 3312 614 3320
rect 573 3286 588 3312
rect 595 3286 614 3312
rect 678 3308 740 3320
rect 752 3308 827 3320
rect 885 3308 960 3320
rect 972 3308 1003 3320
rect 1009 3308 1044 3320
rect 678 3306 840 3308
rect 573 3278 614 3286
rect 696 3282 709 3306
rect 724 3304 739 3306
rect 536 3268 537 3278
rect 552 3268 565 3278
rect 579 3268 580 3278
rect 595 3268 608 3278
rect 623 3268 653 3282
rect 696 3268 739 3282
rect 763 3279 770 3286
rect 773 3282 840 3306
rect 872 3306 1044 3308
rect 842 3284 870 3288
rect 872 3284 952 3306
rect 973 3304 988 3306
rect 842 3282 952 3284
rect 773 3278 952 3282
rect 746 3268 776 3278
rect 778 3268 931 3278
rect 939 3268 969 3278
rect 973 3268 1003 3282
rect 1031 3268 1044 3306
rect 1116 3312 1151 3320
rect 1116 3286 1117 3312
rect 1124 3286 1151 3312
rect 1059 3268 1089 3282
rect 1116 3278 1151 3286
rect 1153 3312 1194 3320
rect 1153 3286 1168 3312
rect 1175 3286 1194 3312
rect 1258 3308 1320 3320
rect 1332 3308 1407 3320
rect 1465 3308 1540 3320
rect 1552 3308 1583 3320
rect 1589 3308 1624 3320
rect 1258 3306 1420 3308
rect 1153 3278 1194 3286
rect 1276 3282 1289 3306
rect 1304 3304 1319 3306
rect 1116 3268 1117 3278
rect 1132 3268 1145 3278
rect 1159 3268 1160 3278
rect 1175 3268 1188 3278
rect 1203 3268 1233 3282
rect 1276 3268 1319 3282
rect 1343 3279 1350 3286
rect 1353 3282 1420 3306
rect 1452 3306 1624 3308
rect 1422 3284 1450 3288
rect 1452 3284 1532 3306
rect 1553 3304 1568 3306
rect 1422 3282 1532 3284
rect 1353 3278 1532 3282
rect 1326 3268 1356 3278
rect 1358 3268 1511 3278
rect 1519 3268 1549 3278
rect 1553 3268 1583 3282
rect 1611 3268 1624 3306
rect 1696 3312 1731 3320
rect 1696 3286 1697 3312
rect 1704 3286 1731 3312
rect 1639 3268 1669 3282
rect 1696 3278 1731 3286
rect 1733 3312 1774 3320
rect 1733 3286 1748 3312
rect 1755 3286 1774 3312
rect 1838 3308 1900 3320
rect 1912 3308 1987 3320
rect 2045 3308 2120 3320
rect 2132 3308 2163 3320
rect 2169 3308 2204 3320
rect 1838 3306 2000 3308
rect 1733 3278 1774 3286
rect 1856 3282 1869 3306
rect 1884 3304 1899 3306
rect 1696 3268 1697 3278
rect 1712 3268 1725 3278
rect 1739 3268 1740 3278
rect 1755 3268 1768 3278
rect 1783 3268 1813 3282
rect 1856 3268 1899 3282
rect 1923 3279 1930 3286
rect 1933 3282 2000 3306
rect 2032 3306 2204 3308
rect 2002 3284 2030 3288
rect 2032 3284 2112 3306
rect 2133 3304 2148 3306
rect 2002 3282 2112 3284
rect 1933 3278 2112 3282
rect 1906 3268 1936 3278
rect 1938 3268 2091 3278
rect 2099 3268 2129 3278
rect 2133 3268 2163 3282
rect 2191 3268 2204 3306
rect 2276 3312 2311 3320
rect 2276 3286 2277 3312
rect 2284 3286 2311 3312
rect 2219 3268 2249 3282
rect 2276 3278 2311 3286
rect 2313 3312 2354 3320
rect 2313 3286 2328 3312
rect 2335 3286 2354 3312
rect 2418 3308 2480 3320
rect 2492 3308 2567 3320
rect 2625 3308 2700 3320
rect 2712 3308 2743 3320
rect 2749 3308 2784 3320
rect 2418 3306 2580 3308
rect 2313 3278 2354 3286
rect 2436 3282 2449 3306
rect 2464 3304 2479 3306
rect 2276 3268 2277 3278
rect 2292 3268 2305 3278
rect 2319 3268 2320 3278
rect 2335 3268 2348 3278
rect 2363 3268 2393 3282
rect 2436 3268 2479 3282
rect 2503 3279 2510 3286
rect 2513 3282 2580 3306
rect 2612 3306 2784 3308
rect 2582 3284 2610 3288
rect 2612 3284 2692 3306
rect 2713 3304 2728 3306
rect 2582 3282 2692 3284
rect 2513 3278 2692 3282
rect 2486 3268 2516 3278
rect 2518 3268 2671 3278
rect 2679 3268 2709 3278
rect 2713 3268 2743 3282
rect 2771 3268 2784 3306
rect 2856 3312 2891 3320
rect 2856 3286 2857 3312
rect 2864 3286 2891 3312
rect 2799 3268 2829 3282
rect 2856 3278 2891 3286
rect 2893 3312 2934 3320
rect 2893 3286 2908 3312
rect 2915 3286 2934 3312
rect 2998 3308 3060 3320
rect 3072 3308 3147 3320
rect 3205 3308 3280 3320
rect 3292 3308 3323 3320
rect 3329 3308 3364 3320
rect 2998 3306 3160 3308
rect 2893 3278 2934 3286
rect 3016 3282 3029 3306
rect 3044 3304 3059 3306
rect 2856 3268 2857 3278
rect 2872 3268 2885 3278
rect 2899 3268 2900 3278
rect 2915 3268 2928 3278
rect 2943 3268 2973 3282
rect 3016 3268 3059 3282
rect 3083 3279 3090 3286
rect 3093 3282 3160 3306
rect 3192 3306 3364 3308
rect 3162 3284 3190 3288
rect 3192 3284 3272 3306
rect 3293 3304 3308 3306
rect 3162 3282 3272 3284
rect 3093 3278 3272 3282
rect 3066 3268 3096 3278
rect 3098 3268 3251 3278
rect 3259 3268 3289 3278
rect 3293 3268 3323 3282
rect 3351 3268 3364 3306
rect 3436 3312 3471 3320
rect 3436 3286 3437 3312
rect 3444 3286 3471 3312
rect 3379 3268 3409 3282
rect 3436 3278 3471 3286
rect 3473 3312 3514 3320
rect 3473 3286 3488 3312
rect 3495 3286 3514 3312
rect 3578 3308 3640 3320
rect 3652 3308 3727 3320
rect 3785 3308 3860 3320
rect 3872 3308 3903 3320
rect 3909 3308 3944 3320
rect 3578 3306 3740 3308
rect 3473 3278 3514 3286
rect 3596 3282 3609 3306
rect 3624 3304 3639 3306
rect 3436 3268 3437 3278
rect 3452 3268 3465 3278
rect 3479 3268 3480 3278
rect 3495 3268 3508 3278
rect 3523 3268 3553 3282
rect 3596 3268 3639 3282
rect 3663 3279 3670 3286
rect 3673 3282 3740 3306
rect 3772 3306 3944 3308
rect 3742 3284 3770 3288
rect 3772 3284 3852 3306
rect 3873 3304 3888 3306
rect 3742 3282 3852 3284
rect 3673 3278 3852 3282
rect 3646 3268 3676 3278
rect 3678 3268 3831 3278
rect 3839 3268 3869 3278
rect 3873 3268 3903 3282
rect 3931 3268 3944 3306
rect 4016 3312 4051 3320
rect 4016 3286 4017 3312
rect 4024 3286 4051 3312
rect 3959 3268 3989 3282
rect 4016 3278 4051 3286
rect 4053 3312 4094 3320
rect 4053 3286 4068 3312
rect 4075 3286 4094 3312
rect 4158 3308 4220 3320
rect 4232 3308 4307 3320
rect 4365 3308 4440 3320
rect 4452 3308 4483 3320
rect 4489 3308 4524 3320
rect 4158 3306 4320 3308
rect 4053 3278 4094 3286
rect 4176 3282 4189 3306
rect 4204 3304 4219 3306
rect 4016 3268 4017 3278
rect 4032 3268 4045 3278
rect 4059 3268 4060 3278
rect 4075 3268 4088 3278
rect 4103 3268 4133 3282
rect 4176 3268 4219 3282
rect 4243 3279 4250 3286
rect 4253 3282 4320 3306
rect 4352 3306 4524 3308
rect 4322 3284 4350 3288
rect 4352 3284 4432 3306
rect 4453 3304 4468 3306
rect 4322 3282 4432 3284
rect 4253 3278 4432 3282
rect 4226 3268 4256 3278
rect 4258 3268 4411 3278
rect 4419 3268 4449 3278
rect 4453 3268 4483 3282
rect 4511 3268 4524 3306
rect 4596 3312 4631 3320
rect 4596 3286 4597 3312
rect 4604 3286 4631 3312
rect 4539 3268 4569 3282
rect 4596 3278 4631 3286
rect 4633 3312 4674 3320
rect 4633 3286 4648 3312
rect 4655 3286 4674 3312
rect 4738 3308 4800 3320
rect 4812 3308 4887 3320
rect 4945 3308 5020 3320
rect 5032 3308 5063 3320
rect 5069 3308 5104 3320
rect 4738 3306 4900 3308
rect 4633 3278 4674 3286
rect 4756 3282 4769 3306
rect 4784 3304 4799 3306
rect 4596 3268 4597 3278
rect 4612 3268 4625 3278
rect 4639 3268 4640 3278
rect 4655 3268 4668 3278
rect 4683 3268 4713 3282
rect 4756 3268 4799 3282
rect 4823 3279 4830 3286
rect 4833 3282 4900 3306
rect 4932 3306 5104 3308
rect 4902 3284 4930 3288
rect 4932 3284 5012 3306
rect 5033 3304 5048 3306
rect 4902 3282 5012 3284
rect 4833 3278 5012 3282
rect 4806 3268 4836 3278
rect 4838 3268 4991 3278
rect 4999 3268 5029 3278
rect 5033 3268 5063 3282
rect 5091 3268 5104 3306
rect 5176 3312 5211 3320
rect 5176 3286 5177 3312
rect 5184 3286 5211 3312
rect 5119 3268 5149 3282
rect 5176 3278 5211 3286
rect 5213 3312 5254 3320
rect 5213 3286 5228 3312
rect 5235 3286 5254 3312
rect 5318 3308 5380 3320
rect 5392 3308 5467 3320
rect 5525 3308 5600 3320
rect 5612 3308 5643 3320
rect 5649 3308 5684 3320
rect 5318 3306 5480 3308
rect 5213 3278 5254 3286
rect 5336 3282 5349 3306
rect 5364 3304 5379 3306
rect 5176 3268 5177 3278
rect 5192 3268 5205 3278
rect 5219 3268 5220 3278
rect 5235 3268 5248 3278
rect 5263 3268 5293 3282
rect 5336 3268 5379 3282
rect 5403 3279 5410 3286
rect 5413 3282 5480 3306
rect 5512 3306 5684 3308
rect 5482 3284 5510 3288
rect 5512 3284 5592 3306
rect 5613 3304 5628 3306
rect 5482 3282 5592 3284
rect 5413 3278 5592 3282
rect 5386 3268 5416 3278
rect 5418 3268 5571 3278
rect 5579 3268 5609 3278
rect 5613 3268 5643 3282
rect 5671 3268 5684 3306
rect 5756 3312 5791 3320
rect 5756 3286 5757 3312
rect 5764 3286 5791 3312
rect 5699 3268 5729 3282
rect 5756 3278 5791 3286
rect 5793 3312 5834 3320
rect 5793 3286 5808 3312
rect 5815 3286 5834 3312
rect 5898 3308 5960 3320
rect 5972 3308 6047 3320
rect 6105 3308 6180 3320
rect 6192 3308 6223 3320
rect 6229 3308 6264 3320
rect 5898 3306 6060 3308
rect 5793 3278 5834 3286
rect 5916 3282 5929 3306
rect 5944 3304 5959 3306
rect 5756 3268 5757 3278
rect 5772 3268 5785 3278
rect 5799 3268 5800 3278
rect 5815 3268 5828 3278
rect 5843 3268 5873 3282
rect 5916 3268 5959 3282
rect 5983 3279 5990 3286
rect 5993 3282 6060 3306
rect 6092 3306 6264 3308
rect 6062 3284 6090 3288
rect 6092 3284 6172 3306
rect 6193 3304 6208 3306
rect 6062 3282 6172 3284
rect 5993 3278 6172 3282
rect 5966 3268 5996 3278
rect 5998 3268 6151 3278
rect 6159 3268 6189 3278
rect 6193 3268 6223 3282
rect 6251 3268 6264 3306
rect 6336 3312 6371 3320
rect 6336 3286 6337 3312
rect 6344 3286 6371 3312
rect 6279 3268 6309 3282
rect 6336 3278 6371 3286
rect 6373 3312 6414 3320
rect 6373 3286 6388 3312
rect 6395 3286 6414 3312
rect 6478 3308 6540 3320
rect 6552 3308 6627 3320
rect 6685 3308 6760 3320
rect 6772 3308 6803 3320
rect 6809 3308 6844 3320
rect 6478 3306 6640 3308
rect 6373 3278 6414 3286
rect 6496 3282 6509 3306
rect 6524 3304 6539 3306
rect 6336 3268 6337 3278
rect 6352 3268 6365 3278
rect 6379 3268 6380 3278
rect 6395 3268 6408 3278
rect 6423 3268 6453 3282
rect 6496 3268 6539 3282
rect 6563 3279 6570 3286
rect 6573 3282 6640 3306
rect 6672 3306 6844 3308
rect 6642 3284 6670 3288
rect 6672 3284 6752 3306
rect 6773 3304 6788 3306
rect 6642 3282 6752 3284
rect 6573 3278 6752 3282
rect 6546 3268 6576 3278
rect 6578 3268 6731 3278
rect 6739 3268 6769 3278
rect 6773 3268 6803 3282
rect 6831 3268 6844 3306
rect 6916 3312 6951 3320
rect 6916 3286 6917 3312
rect 6924 3286 6951 3312
rect 6859 3268 6889 3282
rect 6916 3278 6951 3286
rect 6953 3312 6994 3320
rect 6953 3286 6968 3312
rect 6975 3286 6994 3312
rect 7058 3308 7120 3320
rect 7132 3308 7207 3320
rect 7265 3308 7340 3320
rect 7352 3308 7383 3320
rect 7389 3308 7424 3320
rect 7058 3306 7220 3308
rect 6953 3278 6994 3286
rect 7076 3282 7089 3306
rect 7104 3304 7119 3306
rect 6916 3268 6917 3278
rect 6932 3268 6945 3278
rect 6959 3268 6960 3278
rect 6975 3268 6988 3278
rect 7003 3268 7033 3282
rect 7076 3268 7119 3282
rect 7143 3279 7150 3286
rect 7153 3282 7220 3306
rect 7252 3306 7424 3308
rect 7222 3284 7250 3288
rect 7252 3284 7332 3306
rect 7353 3304 7368 3306
rect 7222 3282 7332 3284
rect 7153 3278 7332 3282
rect 7126 3268 7156 3278
rect 7158 3268 7311 3278
rect 7319 3268 7349 3278
rect 7353 3268 7383 3282
rect 7411 3268 7424 3306
rect 7496 3312 7531 3320
rect 7496 3286 7497 3312
rect 7504 3286 7531 3312
rect 7439 3268 7469 3282
rect 7496 3278 7531 3286
rect 7533 3312 7574 3320
rect 7533 3286 7548 3312
rect 7555 3286 7574 3312
rect 7638 3308 7700 3320
rect 7712 3308 7787 3320
rect 7845 3308 7920 3320
rect 7932 3308 7963 3320
rect 7969 3308 8004 3320
rect 7638 3306 7800 3308
rect 7533 3278 7574 3286
rect 7656 3282 7669 3306
rect 7684 3304 7699 3306
rect 7496 3268 7497 3278
rect 7512 3268 7525 3278
rect 7539 3268 7540 3278
rect 7555 3268 7568 3278
rect 7583 3268 7613 3282
rect 7656 3268 7699 3282
rect 7723 3279 7730 3286
rect 7733 3282 7800 3306
rect 7832 3306 8004 3308
rect 7802 3284 7830 3288
rect 7832 3284 7912 3306
rect 7933 3304 7948 3306
rect 7802 3282 7912 3284
rect 7733 3278 7912 3282
rect 7706 3268 7736 3278
rect 7738 3268 7891 3278
rect 7899 3268 7929 3278
rect 7933 3268 7963 3282
rect 7991 3268 8004 3306
rect 8076 3312 8111 3320
rect 8076 3286 8077 3312
rect 8084 3286 8111 3312
rect 8019 3268 8049 3282
rect 8076 3278 8111 3286
rect 8113 3312 8154 3320
rect 8113 3286 8128 3312
rect 8135 3286 8154 3312
rect 8218 3308 8280 3320
rect 8292 3308 8367 3320
rect 8425 3308 8500 3320
rect 8512 3308 8543 3320
rect 8549 3308 8584 3320
rect 8218 3306 8380 3308
rect 8113 3278 8154 3286
rect 8236 3282 8249 3306
rect 8264 3304 8279 3306
rect 8076 3268 8077 3278
rect 8092 3268 8105 3278
rect 8119 3268 8120 3278
rect 8135 3268 8148 3278
rect 8163 3268 8193 3282
rect 8236 3268 8279 3282
rect 8303 3279 8310 3286
rect 8313 3282 8380 3306
rect 8412 3306 8584 3308
rect 8382 3284 8410 3288
rect 8412 3284 8492 3306
rect 8513 3304 8528 3306
rect 8382 3282 8492 3284
rect 8313 3278 8492 3282
rect 8286 3268 8316 3278
rect 8318 3268 8471 3278
rect 8479 3268 8509 3278
rect 8513 3268 8543 3282
rect 8571 3268 8584 3306
rect 8656 3312 8691 3320
rect 8656 3286 8657 3312
rect 8664 3286 8691 3312
rect 8599 3268 8629 3282
rect 8656 3278 8691 3286
rect 8693 3312 8734 3320
rect 8693 3286 8708 3312
rect 8715 3286 8734 3312
rect 8798 3308 8860 3320
rect 8872 3308 8947 3320
rect 9005 3308 9080 3320
rect 9092 3308 9123 3320
rect 9129 3308 9164 3320
rect 8798 3306 8960 3308
rect 8693 3278 8734 3286
rect 8816 3282 8829 3306
rect 8844 3304 8859 3306
rect 8656 3268 8657 3278
rect 8672 3268 8685 3278
rect 8699 3268 8700 3278
rect 8715 3268 8728 3278
rect 8743 3268 8773 3282
rect 8816 3268 8859 3282
rect 8883 3279 8890 3286
rect 8893 3282 8960 3306
rect 8992 3306 9164 3308
rect 8962 3284 8990 3288
rect 8992 3284 9072 3306
rect 9093 3304 9108 3306
rect 8962 3282 9072 3284
rect 8893 3278 9072 3282
rect 8866 3268 8896 3278
rect 8898 3268 9051 3278
rect 9059 3268 9089 3278
rect 9093 3268 9123 3282
rect 9151 3268 9164 3306
rect 9236 3312 9271 3320
rect 9236 3286 9237 3312
rect 9244 3286 9271 3312
rect 9179 3268 9209 3282
rect 9236 3278 9271 3286
rect 9236 3268 9237 3278
rect 9252 3268 9265 3278
rect -1 3262 9265 3268
rect 0 3254 9265 3262
rect 15 3224 28 3254
rect 43 3236 73 3254
rect 116 3240 130 3254
rect 166 3240 386 3254
rect 117 3238 130 3240
rect 83 3226 98 3238
rect 80 3224 102 3226
rect 107 3224 137 3238
rect 198 3236 351 3240
rect 180 3224 372 3236
rect 415 3224 445 3238
rect 451 3224 464 3254
rect 479 3236 509 3254
rect 552 3224 565 3254
rect 595 3224 608 3254
rect 623 3236 653 3254
rect 696 3240 710 3254
rect 746 3240 966 3254
rect 697 3238 710 3240
rect 663 3226 678 3238
rect 660 3224 682 3226
rect 687 3224 717 3238
rect 778 3236 931 3240
rect 760 3224 952 3236
rect 995 3224 1025 3238
rect 1031 3224 1044 3254
rect 1059 3236 1089 3254
rect 1132 3224 1145 3254
rect 1175 3224 1188 3254
rect 1203 3236 1233 3254
rect 1276 3240 1290 3254
rect 1326 3240 1546 3254
rect 1277 3238 1290 3240
rect 1243 3226 1258 3238
rect 1240 3224 1262 3226
rect 1267 3224 1297 3238
rect 1358 3236 1511 3240
rect 1340 3224 1532 3236
rect 1575 3224 1605 3238
rect 1611 3224 1624 3254
rect 1639 3236 1669 3254
rect 1712 3224 1725 3254
rect 1755 3224 1768 3254
rect 1783 3236 1813 3254
rect 1856 3240 1870 3254
rect 1906 3240 2126 3254
rect 1857 3238 1870 3240
rect 1823 3226 1838 3238
rect 1820 3224 1842 3226
rect 1847 3224 1877 3238
rect 1938 3236 2091 3240
rect 1920 3224 2112 3236
rect 2155 3224 2185 3238
rect 2191 3224 2204 3254
rect 2219 3236 2249 3254
rect 2292 3224 2305 3254
rect 2335 3224 2348 3254
rect 2363 3236 2393 3254
rect 2436 3240 2450 3254
rect 2486 3240 2706 3254
rect 2437 3238 2450 3240
rect 2403 3226 2418 3238
rect 2400 3224 2422 3226
rect 2427 3224 2457 3238
rect 2518 3236 2671 3240
rect 2500 3224 2692 3236
rect 2735 3224 2765 3238
rect 2771 3224 2784 3254
rect 2799 3236 2829 3254
rect 2872 3224 2885 3254
rect 2915 3224 2928 3254
rect 2943 3236 2973 3254
rect 3016 3240 3030 3254
rect 3066 3240 3286 3254
rect 3017 3238 3030 3240
rect 2983 3226 2998 3238
rect 2980 3224 3002 3226
rect 3007 3224 3037 3238
rect 3098 3236 3251 3240
rect 3080 3224 3272 3236
rect 3315 3224 3345 3238
rect 3351 3224 3364 3254
rect 3379 3236 3409 3254
rect 3452 3224 3465 3254
rect 3495 3224 3508 3254
rect 3523 3236 3553 3254
rect 3596 3240 3610 3254
rect 3646 3240 3866 3254
rect 3597 3238 3610 3240
rect 3563 3226 3578 3238
rect 3560 3224 3582 3226
rect 3587 3224 3617 3238
rect 3678 3236 3831 3240
rect 3660 3224 3852 3236
rect 3895 3224 3925 3238
rect 3931 3224 3944 3254
rect 3959 3236 3989 3254
rect 4032 3224 4045 3254
rect 4075 3224 4088 3254
rect 4103 3236 4133 3254
rect 4176 3240 4190 3254
rect 4226 3240 4446 3254
rect 4177 3238 4190 3240
rect 4143 3226 4158 3238
rect 4140 3224 4162 3226
rect 4167 3224 4197 3238
rect 4258 3236 4411 3240
rect 4240 3224 4432 3236
rect 4475 3224 4505 3238
rect 4511 3224 4524 3254
rect 4539 3236 4569 3254
rect 4612 3224 4625 3254
rect 4655 3224 4668 3254
rect 4683 3236 4713 3254
rect 4756 3240 4770 3254
rect 4806 3240 5026 3254
rect 4757 3238 4770 3240
rect 4723 3226 4738 3238
rect 4720 3224 4742 3226
rect 4747 3224 4777 3238
rect 4838 3236 4991 3240
rect 4820 3224 5012 3236
rect 5055 3224 5085 3238
rect 5091 3224 5104 3254
rect 5119 3236 5149 3254
rect 5192 3224 5205 3254
rect 5235 3224 5248 3254
rect 5263 3236 5293 3254
rect 5336 3240 5350 3254
rect 5386 3240 5606 3254
rect 5337 3238 5350 3240
rect 5303 3226 5318 3238
rect 5300 3224 5322 3226
rect 5327 3224 5357 3238
rect 5418 3236 5571 3240
rect 5400 3224 5592 3236
rect 5635 3224 5665 3238
rect 5671 3224 5684 3254
rect 5699 3236 5729 3254
rect 5772 3224 5785 3254
rect 5815 3224 5828 3254
rect 5843 3236 5873 3254
rect 5916 3240 5930 3254
rect 5966 3240 6186 3254
rect 5917 3238 5930 3240
rect 5883 3226 5898 3238
rect 5880 3224 5902 3226
rect 5907 3224 5937 3238
rect 5998 3236 6151 3240
rect 5980 3224 6172 3236
rect 6215 3224 6245 3238
rect 6251 3224 6264 3254
rect 6279 3236 6309 3254
rect 6352 3224 6365 3254
rect 6395 3224 6408 3254
rect 6423 3236 6453 3254
rect 6496 3240 6510 3254
rect 6546 3240 6766 3254
rect 6497 3238 6510 3240
rect 6463 3226 6478 3238
rect 6460 3224 6482 3226
rect 6487 3224 6517 3238
rect 6578 3236 6731 3240
rect 6560 3224 6752 3236
rect 6795 3224 6825 3238
rect 6831 3224 6844 3254
rect 6859 3236 6889 3254
rect 6932 3224 6945 3254
rect 6975 3224 6988 3254
rect 7003 3236 7033 3254
rect 7076 3240 7090 3254
rect 7126 3240 7346 3254
rect 7077 3238 7090 3240
rect 7043 3226 7058 3238
rect 7040 3224 7062 3226
rect 7067 3224 7097 3238
rect 7158 3236 7311 3240
rect 7140 3224 7332 3236
rect 7375 3224 7405 3238
rect 7411 3224 7424 3254
rect 7439 3236 7469 3254
rect 7512 3224 7525 3254
rect 7555 3224 7568 3254
rect 7583 3236 7613 3254
rect 7656 3240 7670 3254
rect 7706 3240 7926 3254
rect 7657 3238 7670 3240
rect 7623 3226 7638 3238
rect 7620 3224 7642 3226
rect 7647 3224 7677 3238
rect 7738 3236 7891 3240
rect 7720 3224 7912 3236
rect 7955 3224 7985 3238
rect 7991 3224 8004 3254
rect 8019 3236 8049 3254
rect 8092 3224 8105 3254
rect 8135 3224 8148 3254
rect 8163 3236 8193 3254
rect 8236 3240 8250 3254
rect 8286 3240 8506 3254
rect 8237 3238 8250 3240
rect 8203 3226 8218 3238
rect 8200 3224 8222 3226
rect 8227 3224 8257 3238
rect 8318 3236 8471 3240
rect 8300 3224 8492 3236
rect 8535 3224 8565 3238
rect 8571 3224 8584 3254
rect 8599 3236 8629 3254
rect 8672 3224 8685 3254
rect 8715 3224 8728 3254
rect 8743 3236 8773 3254
rect 8816 3240 8830 3254
rect 8866 3240 9086 3254
rect 8817 3238 8830 3240
rect 8783 3226 8798 3238
rect 8780 3224 8802 3226
rect 8807 3224 8837 3238
rect 8898 3236 9051 3240
rect 8880 3224 9072 3236
rect 9115 3224 9145 3238
rect 9151 3224 9164 3254
rect 9179 3236 9209 3254
rect 9252 3224 9265 3254
rect 0 3210 9265 3224
rect 15 3106 28 3210
rect 73 3188 74 3198
rect 89 3188 102 3198
rect 73 3184 102 3188
rect 107 3184 137 3210
rect 155 3196 171 3198
rect 243 3196 296 3210
rect 244 3194 308 3196
rect 351 3194 366 3210
rect 415 3207 445 3210
rect 415 3204 451 3207
rect 381 3196 397 3198
rect 155 3184 170 3188
rect 73 3182 170 3184
rect 198 3182 366 3194
rect 382 3184 397 3188
rect 415 3185 454 3204
rect 473 3198 480 3199
rect 479 3191 480 3198
rect 463 3188 464 3191
rect 479 3188 492 3191
rect 415 3184 445 3185
rect 454 3184 460 3185
rect 463 3184 492 3188
rect 382 3183 492 3184
rect 382 3182 498 3183
rect 57 3174 108 3182
rect 57 3162 82 3174
rect 89 3162 108 3174
rect 139 3174 189 3182
rect 139 3166 155 3174
rect 162 3172 189 3174
rect 198 3172 419 3182
rect 162 3162 419 3172
rect 448 3174 498 3182
rect 448 3165 464 3174
rect 57 3154 108 3162
rect 155 3154 419 3162
rect 445 3162 464 3165
rect 471 3162 498 3174
rect 445 3154 498 3162
rect 73 3146 74 3154
rect 89 3146 102 3154
rect 73 3138 89 3146
rect 70 3131 89 3134
rect 70 3122 92 3131
rect 43 3112 92 3122
rect 43 3106 73 3112
rect 92 3107 97 3112
rect 15 3090 89 3106
rect 107 3098 137 3154
rect 172 3144 380 3154
rect 415 3150 460 3154
rect 463 3153 464 3154
rect 479 3153 492 3154
rect 198 3114 387 3144
rect 213 3111 387 3114
rect 206 3108 387 3111
rect 15 3088 28 3090
rect 43 3088 77 3090
rect 15 3072 89 3088
rect 116 3084 129 3098
rect 144 3084 160 3100
rect 206 3095 217 3108
rect -1 3050 0 3066
rect 15 3050 28 3072
rect 43 3050 73 3072
rect 116 3068 178 3084
rect 206 3077 217 3093
rect 222 3088 232 3108
rect 242 3088 256 3108
rect 259 3095 268 3108
rect 284 3095 293 3108
rect 222 3077 256 3088
rect 259 3077 268 3093
rect 284 3077 293 3093
rect 300 3088 310 3108
rect 320 3088 334 3108
rect 335 3095 346 3108
rect 300 3077 334 3088
rect 335 3077 346 3093
rect 392 3084 408 3100
rect 415 3098 445 3150
rect 479 3146 480 3153
rect 464 3138 480 3146
rect 451 3106 464 3125
rect 479 3106 509 3122
rect 451 3090 525 3106
rect 451 3088 464 3090
rect 479 3088 513 3090
rect 116 3066 129 3068
rect 144 3066 178 3068
rect 116 3050 178 3066
rect 222 3061 238 3064
rect 300 3061 330 3072
rect 378 3068 424 3084
rect 451 3072 525 3088
rect 378 3066 412 3068
rect 377 3050 424 3066
rect 451 3050 464 3072
rect 479 3050 509 3072
rect 536 3050 537 3066
rect 552 3050 565 3210
rect 595 3106 608 3210
rect 653 3188 654 3198
rect 669 3188 682 3198
rect 653 3184 682 3188
rect 687 3184 717 3210
rect 735 3196 751 3198
rect 823 3196 876 3210
rect 824 3194 888 3196
rect 931 3194 946 3210
rect 995 3207 1025 3210
rect 995 3204 1031 3207
rect 961 3196 977 3198
rect 735 3184 750 3188
rect 653 3182 750 3184
rect 778 3182 946 3194
rect 962 3184 977 3188
rect 995 3185 1034 3204
rect 1053 3198 1060 3199
rect 1059 3191 1060 3198
rect 1043 3188 1044 3191
rect 1059 3188 1072 3191
rect 995 3184 1025 3185
rect 1034 3184 1040 3185
rect 1043 3184 1072 3188
rect 962 3183 1072 3184
rect 962 3182 1078 3183
rect 637 3174 688 3182
rect 637 3162 662 3174
rect 669 3162 688 3174
rect 719 3174 769 3182
rect 719 3166 735 3174
rect 742 3172 769 3174
rect 778 3172 999 3182
rect 742 3162 999 3172
rect 1028 3174 1078 3182
rect 1028 3165 1044 3174
rect 637 3154 688 3162
rect 735 3154 999 3162
rect 1025 3162 1044 3165
rect 1051 3162 1078 3174
rect 1025 3154 1078 3162
rect 653 3146 654 3154
rect 669 3146 682 3154
rect 653 3138 669 3146
rect 650 3131 669 3134
rect 650 3122 672 3131
rect 623 3112 672 3122
rect 623 3106 653 3112
rect 672 3107 677 3112
rect 595 3090 669 3106
rect 687 3098 717 3154
rect 752 3144 960 3154
rect 995 3150 1040 3154
rect 1043 3153 1044 3154
rect 1059 3153 1072 3154
rect 778 3114 967 3144
rect 793 3111 967 3114
rect 786 3108 967 3111
rect 595 3088 608 3090
rect 623 3088 657 3090
rect 595 3072 669 3088
rect 696 3084 709 3098
rect 724 3084 740 3100
rect 786 3095 797 3108
rect 579 3050 580 3066
rect 595 3050 608 3072
rect 623 3050 653 3072
rect 696 3068 758 3084
rect 786 3077 797 3093
rect 802 3088 812 3108
rect 822 3088 836 3108
rect 839 3095 848 3108
rect 864 3095 873 3108
rect 802 3077 836 3088
rect 839 3077 848 3093
rect 864 3077 873 3093
rect 880 3088 890 3108
rect 900 3088 914 3108
rect 915 3095 926 3108
rect 880 3077 914 3088
rect 915 3077 926 3093
rect 972 3084 988 3100
rect 995 3098 1025 3150
rect 1059 3146 1060 3153
rect 1044 3138 1060 3146
rect 1031 3106 1044 3125
rect 1059 3106 1089 3122
rect 1031 3090 1105 3106
rect 1031 3088 1044 3090
rect 1059 3088 1093 3090
rect 696 3066 709 3068
rect 724 3066 758 3068
rect 696 3050 758 3066
rect 802 3061 818 3064
rect 880 3061 910 3072
rect 958 3068 1004 3084
rect 1031 3072 1105 3088
rect 958 3066 992 3068
rect 957 3050 1004 3066
rect 1031 3050 1044 3072
rect 1059 3050 1089 3072
rect 1116 3050 1117 3066
rect 1132 3050 1145 3210
rect 1175 3106 1188 3210
rect 1233 3188 1234 3198
rect 1249 3188 1262 3198
rect 1233 3184 1262 3188
rect 1267 3184 1297 3210
rect 1315 3196 1331 3198
rect 1403 3196 1456 3210
rect 1404 3194 1468 3196
rect 1511 3194 1526 3210
rect 1575 3207 1605 3210
rect 1575 3204 1611 3207
rect 1541 3196 1557 3198
rect 1315 3184 1330 3188
rect 1233 3182 1330 3184
rect 1358 3182 1526 3194
rect 1542 3184 1557 3188
rect 1575 3185 1614 3204
rect 1633 3198 1640 3199
rect 1639 3191 1640 3198
rect 1623 3188 1624 3191
rect 1639 3188 1652 3191
rect 1575 3184 1605 3185
rect 1614 3184 1620 3185
rect 1623 3184 1652 3188
rect 1542 3183 1652 3184
rect 1542 3182 1658 3183
rect 1217 3174 1268 3182
rect 1217 3162 1242 3174
rect 1249 3162 1268 3174
rect 1299 3174 1349 3182
rect 1299 3166 1315 3174
rect 1322 3172 1349 3174
rect 1358 3172 1579 3182
rect 1322 3162 1579 3172
rect 1608 3174 1658 3182
rect 1608 3165 1624 3174
rect 1217 3154 1268 3162
rect 1315 3154 1579 3162
rect 1605 3162 1624 3165
rect 1631 3162 1658 3174
rect 1605 3154 1658 3162
rect 1233 3146 1234 3154
rect 1249 3146 1262 3154
rect 1233 3138 1249 3146
rect 1230 3131 1249 3134
rect 1230 3122 1252 3131
rect 1203 3112 1252 3122
rect 1203 3106 1233 3112
rect 1252 3107 1257 3112
rect 1175 3090 1249 3106
rect 1267 3098 1297 3154
rect 1332 3144 1540 3154
rect 1575 3150 1620 3154
rect 1623 3153 1624 3154
rect 1639 3153 1652 3154
rect 1358 3114 1547 3144
rect 1373 3111 1547 3114
rect 1366 3108 1547 3111
rect 1175 3088 1188 3090
rect 1203 3088 1237 3090
rect 1175 3072 1249 3088
rect 1276 3084 1289 3098
rect 1304 3084 1320 3100
rect 1366 3095 1377 3108
rect 1159 3050 1160 3066
rect 1175 3050 1188 3072
rect 1203 3050 1233 3072
rect 1276 3068 1338 3084
rect 1366 3077 1377 3093
rect 1382 3088 1392 3108
rect 1402 3088 1416 3108
rect 1419 3095 1428 3108
rect 1444 3095 1453 3108
rect 1382 3077 1416 3088
rect 1419 3077 1428 3093
rect 1444 3077 1453 3093
rect 1460 3088 1470 3108
rect 1480 3088 1494 3108
rect 1495 3095 1506 3108
rect 1460 3077 1494 3088
rect 1495 3077 1506 3093
rect 1552 3084 1568 3100
rect 1575 3098 1605 3150
rect 1639 3146 1640 3153
rect 1624 3138 1640 3146
rect 1611 3106 1624 3125
rect 1639 3106 1669 3122
rect 1611 3090 1685 3106
rect 1611 3088 1624 3090
rect 1639 3088 1673 3090
rect 1276 3066 1289 3068
rect 1304 3066 1338 3068
rect 1276 3050 1338 3066
rect 1382 3061 1398 3064
rect 1460 3061 1490 3072
rect 1538 3068 1584 3084
rect 1611 3072 1685 3088
rect 1538 3066 1572 3068
rect 1537 3050 1584 3066
rect 1611 3050 1624 3072
rect 1639 3050 1669 3072
rect 1696 3050 1697 3066
rect 1712 3050 1725 3210
rect 1755 3106 1768 3210
rect 1813 3188 1814 3198
rect 1829 3188 1842 3198
rect 1813 3184 1842 3188
rect 1847 3184 1877 3210
rect 1895 3196 1911 3198
rect 1983 3196 2036 3210
rect 1984 3194 2048 3196
rect 2091 3194 2106 3210
rect 2155 3207 2185 3210
rect 2155 3204 2191 3207
rect 2121 3196 2137 3198
rect 1895 3184 1910 3188
rect 1813 3182 1910 3184
rect 1938 3182 2106 3194
rect 2122 3184 2137 3188
rect 2155 3185 2194 3204
rect 2213 3198 2220 3199
rect 2219 3191 2220 3198
rect 2203 3188 2204 3191
rect 2219 3188 2232 3191
rect 2155 3184 2185 3185
rect 2194 3184 2200 3185
rect 2203 3184 2232 3188
rect 2122 3183 2232 3184
rect 2122 3182 2238 3183
rect 1797 3174 1848 3182
rect 1797 3162 1822 3174
rect 1829 3162 1848 3174
rect 1879 3174 1929 3182
rect 1879 3166 1895 3174
rect 1902 3172 1929 3174
rect 1938 3172 2159 3182
rect 1902 3162 2159 3172
rect 2188 3174 2238 3182
rect 2188 3165 2204 3174
rect 1797 3154 1848 3162
rect 1895 3154 2159 3162
rect 2185 3162 2204 3165
rect 2211 3162 2238 3174
rect 2185 3154 2238 3162
rect 1813 3146 1814 3154
rect 1829 3146 1842 3154
rect 1813 3138 1829 3146
rect 1810 3131 1829 3134
rect 1810 3122 1832 3131
rect 1783 3112 1832 3122
rect 1783 3106 1813 3112
rect 1832 3107 1837 3112
rect 1755 3090 1829 3106
rect 1847 3098 1877 3154
rect 1912 3144 2120 3154
rect 2155 3150 2200 3154
rect 2203 3153 2204 3154
rect 2219 3153 2232 3154
rect 1938 3114 2127 3144
rect 1953 3111 2127 3114
rect 1946 3108 2127 3111
rect 1755 3088 1768 3090
rect 1783 3088 1817 3090
rect 1755 3072 1829 3088
rect 1856 3084 1869 3098
rect 1884 3084 1900 3100
rect 1946 3095 1957 3108
rect 1739 3050 1740 3066
rect 1755 3050 1768 3072
rect 1783 3050 1813 3072
rect 1856 3068 1918 3084
rect 1946 3077 1957 3093
rect 1962 3088 1972 3108
rect 1982 3088 1996 3108
rect 1999 3095 2008 3108
rect 2024 3095 2033 3108
rect 1962 3077 1996 3088
rect 1999 3077 2008 3093
rect 2024 3077 2033 3093
rect 2040 3088 2050 3108
rect 2060 3088 2074 3108
rect 2075 3095 2086 3108
rect 2040 3077 2074 3088
rect 2075 3077 2086 3093
rect 2132 3084 2148 3100
rect 2155 3098 2185 3150
rect 2219 3146 2220 3153
rect 2204 3138 2220 3146
rect 2191 3106 2204 3125
rect 2219 3106 2249 3122
rect 2191 3090 2265 3106
rect 2191 3088 2204 3090
rect 2219 3088 2253 3090
rect 1856 3066 1869 3068
rect 1884 3066 1918 3068
rect 1856 3050 1918 3066
rect 1962 3061 1976 3064
rect 2040 3061 2070 3072
rect 2118 3068 2164 3084
rect 2191 3072 2265 3088
rect 2118 3066 2152 3068
rect 2117 3050 2164 3066
rect 2191 3050 2204 3072
rect 2219 3050 2249 3072
rect 2276 3050 2277 3066
rect 2292 3050 2305 3210
rect 2335 3106 2348 3210
rect 2393 3188 2394 3198
rect 2409 3188 2422 3198
rect 2393 3184 2422 3188
rect 2427 3184 2457 3210
rect 2475 3196 2491 3198
rect 2563 3196 2616 3210
rect 2564 3194 2628 3196
rect 2671 3194 2686 3210
rect 2735 3207 2765 3210
rect 2735 3204 2771 3207
rect 2701 3196 2717 3198
rect 2475 3184 2490 3188
rect 2393 3182 2490 3184
rect 2518 3182 2686 3194
rect 2702 3184 2717 3188
rect 2735 3185 2774 3204
rect 2793 3198 2800 3199
rect 2799 3191 2800 3198
rect 2783 3188 2784 3191
rect 2799 3188 2812 3191
rect 2735 3184 2765 3185
rect 2774 3184 2780 3185
rect 2783 3184 2812 3188
rect 2702 3183 2812 3184
rect 2702 3182 2818 3183
rect 2377 3174 2428 3182
rect 2377 3162 2402 3174
rect 2409 3162 2428 3174
rect 2459 3174 2509 3182
rect 2459 3166 2475 3174
rect 2482 3172 2509 3174
rect 2518 3172 2739 3182
rect 2482 3162 2739 3172
rect 2768 3174 2818 3182
rect 2768 3165 2784 3174
rect 2377 3154 2428 3162
rect 2475 3154 2739 3162
rect 2765 3162 2784 3165
rect 2791 3162 2818 3174
rect 2765 3154 2818 3162
rect 2393 3146 2394 3154
rect 2409 3146 2422 3154
rect 2393 3138 2409 3146
rect 2390 3131 2409 3134
rect 2390 3122 2412 3131
rect 2363 3112 2412 3122
rect 2363 3106 2393 3112
rect 2412 3107 2417 3112
rect 2335 3090 2409 3106
rect 2427 3098 2457 3154
rect 2492 3144 2700 3154
rect 2735 3150 2780 3154
rect 2783 3153 2784 3154
rect 2799 3153 2812 3154
rect 2518 3114 2707 3144
rect 2533 3111 2707 3114
rect 2526 3108 2707 3111
rect 2335 3088 2348 3090
rect 2363 3088 2397 3090
rect 2335 3072 2409 3088
rect 2436 3084 2449 3098
rect 2464 3084 2480 3100
rect 2526 3095 2537 3108
rect 2319 3050 2320 3066
rect 2335 3050 2348 3072
rect 2363 3050 2393 3072
rect 2436 3068 2498 3084
rect 2526 3077 2537 3093
rect 2542 3088 2552 3108
rect 2562 3088 2576 3108
rect 2579 3095 2588 3108
rect 2604 3095 2613 3108
rect 2542 3077 2576 3088
rect 2579 3077 2588 3093
rect 2604 3077 2613 3093
rect 2620 3088 2630 3108
rect 2640 3088 2654 3108
rect 2655 3095 2666 3108
rect 2620 3077 2654 3088
rect 2655 3077 2666 3093
rect 2712 3084 2728 3100
rect 2735 3098 2765 3150
rect 2799 3146 2800 3153
rect 2784 3138 2800 3146
rect 2771 3106 2784 3125
rect 2799 3106 2829 3122
rect 2771 3090 2845 3106
rect 2771 3088 2784 3090
rect 2799 3088 2833 3090
rect 2436 3066 2449 3068
rect 2464 3066 2498 3068
rect 2436 3050 2498 3066
rect 2542 3061 2558 3064
rect 2620 3061 2650 3072
rect 2698 3068 2744 3084
rect 2771 3072 2845 3088
rect 2698 3066 2732 3068
rect 2697 3050 2744 3066
rect 2771 3050 2784 3072
rect 2799 3050 2829 3072
rect 2856 3050 2857 3066
rect 2872 3050 2885 3210
rect 2915 3106 2928 3210
rect 2973 3188 2974 3198
rect 2989 3188 3002 3198
rect 2973 3184 3002 3188
rect 3007 3184 3037 3210
rect 3055 3196 3071 3198
rect 3143 3196 3196 3210
rect 3144 3194 3208 3196
rect 3251 3194 3266 3210
rect 3315 3207 3345 3210
rect 3315 3204 3351 3207
rect 3281 3196 3297 3198
rect 3055 3184 3070 3188
rect 2973 3182 3070 3184
rect 3098 3182 3266 3194
rect 3282 3184 3297 3188
rect 3315 3185 3354 3204
rect 3373 3198 3380 3199
rect 3379 3191 3380 3198
rect 3363 3188 3364 3191
rect 3379 3188 3392 3191
rect 3315 3184 3345 3185
rect 3354 3184 3360 3185
rect 3363 3184 3392 3188
rect 3282 3183 3392 3184
rect 3282 3182 3398 3183
rect 2957 3174 3008 3182
rect 2957 3162 2982 3174
rect 2989 3162 3008 3174
rect 3039 3174 3089 3182
rect 3039 3166 3055 3174
rect 3062 3172 3089 3174
rect 3098 3172 3319 3182
rect 3062 3162 3319 3172
rect 3348 3174 3398 3182
rect 3348 3165 3364 3174
rect 2957 3154 3008 3162
rect 3055 3154 3319 3162
rect 3345 3162 3364 3165
rect 3371 3162 3398 3174
rect 3345 3154 3398 3162
rect 2973 3146 2974 3154
rect 2989 3146 3002 3154
rect 2973 3138 2989 3146
rect 2970 3131 2989 3134
rect 2970 3122 2992 3131
rect 2943 3112 2992 3122
rect 2943 3106 2973 3112
rect 2992 3107 2997 3112
rect 2915 3090 2989 3106
rect 3007 3098 3037 3154
rect 3072 3144 3280 3154
rect 3315 3150 3360 3154
rect 3363 3153 3364 3154
rect 3379 3153 3392 3154
rect 3098 3114 3287 3144
rect 3113 3111 3287 3114
rect 3106 3108 3287 3111
rect 2915 3088 2928 3090
rect 2943 3088 2977 3090
rect 2915 3072 2989 3088
rect 3016 3084 3029 3098
rect 3044 3084 3060 3100
rect 3106 3095 3117 3108
rect 2899 3050 2900 3066
rect 2915 3050 2928 3072
rect 2943 3050 2973 3072
rect 3016 3068 3078 3084
rect 3106 3077 3117 3093
rect 3122 3088 3132 3108
rect 3142 3088 3156 3108
rect 3159 3095 3168 3108
rect 3184 3095 3193 3108
rect 3122 3077 3156 3088
rect 3159 3077 3168 3093
rect 3184 3077 3193 3093
rect 3200 3088 3210 3108
rect 3220 3088 3234 3108
rect 3235 3095 3246 3108
rect 3200 3077 3234 3088
rect 3235 3077 3246 3093
rect 3292 3084 3308 3100
rect 3315 3098 3345 3150
rect 3379 3146 3380 3153
rect 3364 3138 3380 3146
rect 3351 3106 3364 3125
rect 3379 3106 3409 3122
rect 3351 3090 3425 3106
rect 3351 3088 3364 3090
rect 3379 3088 3413 3090
rect 3016 3066 3029 3068
rect 3044 3066 3078 3068
rect 3016 3050 3078 3066
rect 3122 3061 3138 3064
rect 3200 3061 3230 3072
rect 3278 3068 3324 3084
rect 3351 3072 3425 3088
rect 3278 3066 3312 3068
rect 3277 3050 3324 3066
rect 3351 3050 3364 3072
rect 3379 3050 3409 3072
rect 3436 3050 3437 3066
rect 3452 3050 3465 3210
rect 3495 3106 3508 3210
rect 3553 3188 3554 3198
rect 3569 3188 3582 3198
rect 3553 3184 3582 3188
rect 3587 3184 3617 3210
rect 3635 3196 3651 3198
rect 3723 3196 3776 3210
rect 3724 3194 3788 3196
rect 3831 3194 3846 3210
rect 3895 3207 3925 3210
rect 3895 3204 3931 3207
rect 3861 3196 3877 3198
rect 3635 3184 3650 3188
rect 3553 3182 3650 3184
rect 3678 3182 3846 3194
rect 3862 3184 3877 3188
rect 3895 3185 3934 3204
rect 3953 3198 3960 3199
rect 3959 3191 3960 3198
rect 3943 3188 3944 3191
rect 3959 3188 3972 3191
rect 3895 3184 3925 3185
rect 3934 3184 3940 3185
rect 3943 3184 3972 3188
rect 3862 3183 3972 3184
rect 3862 3182 3978 3183
rect 3537 3174 3588 3182
rect 3537 3162 3562 3174
rect 3569 3162 3588 3174
rect 3619 3174 3669 3182
rect 3619 3166 3635 3174
rect 3642 3172 3669 3174
rect 3678 3172 3899 3182
rect 3642 3162 3899 3172
rect 3928 3174 3978 3182
rect 3928 3165 3944 3174
rect 3537 3154 3588 3162
rect 3635 3154 3899 3162
rect 3925 3162 3944 3165
rect 3951 3162 3978 3174
rect 3925 3154 3978 3162
rect 3553 3146 3554 3154
rect 3569 3146 3582 3154
rect 3553 3138 3569 3146
rect 3550 3131 3569 3134
rect 3550 3122 3572 3131
rect 3523 3112 3572 3122
rect 3523 3106 3553 3112
rect 3572 3107 3577 3112
rect 3495 3090 3569 3106
rect 3587 3098 3617 3154
rect 3652 3144 3860 3154
rect 3895 3150 3940 3154
rect 3943 3153 3944 3154
rect 3959 3153 3972 3154
rect 3678 3114 3867 3144
rect 3693 3111 3867 3114
rect 3686 3108 3867 3111
rect 3495 3088 3508 3090
rect 3523 3088 3557 3090
rect 3495 3072 3569 3088
rect 3596 3084 3609 3098
rect 3624 3084 3640 3100
rect 3686 3095 3697 3108
rect 3479 3050 3480 3066
rect 3495 3050 3508 3072
rect 3523 3050 3553 3072
rect 3596 3068 3658 3084
rect 3686 3077 3697 3093
rect 3702 3088 3712 3108
rect 3722 3088 3736 3108
rect 3739 3095 3748 3108
rect 3764 3095 3773 3108
rect 3702 3077 3736 3088
rect 3739 3077 3748 3093
rect 3764 3077 3773 3093
rect 3780 3088 3790 3108
rect 3800 3088 3814 3108
rect 3815 3095 3826 3108
rect 3780 3077 3814 3088
rect 3815 3077 3826 3093
rect 3872 3084 3888 3100
rect 3895 3098 3925 3150
rect 3959 3146 3960 3153
rect 3944 3138 3960 3146
rect 3931 3106 3944 3125
rect 3959 3106 3989 3122
rect 3931 3090 4005 3106
rect 3931 3088 3944 3090
rect 3959 3088 3993 3090
rect 3596 3066 3609 3068
rect 3624 3066 3658 3068
rect 3596 3050 3658 3066
rect 3702 3061 3718 3064
rect 3780 3061 3810 3072
rect 3858 3068 3904 3084
rect 3931 3072 4005 3088
rect 3858 3066 3892 3068
rect 3857 3050 3904 3066
rect 3931 3050 3944 3072
rect 3959 3050 3989 3072
rect 4016 3050 4017 3066
rect 4032 3050 4045 3210
rect 4075 3106 4088 3210
rect 4133 3188 4134 3198
rect 4149 3188 4162 3198
rect 4133 3184 4162 3188
rect 4167 3184 4197 3210
rect 4215 3196 4231 3198
rect 4303 3196 4356 3210
rect 4304 3194 4368 3196
rect 4411 3194 4426 3210
rect 4475 3207 4505 3210
rect 4475 3204 4511 3207
rect 4441 3196 4457 3198
rect 4215 3184 4230 3188
rect 4133 3182 4230 3184
rect 4258 3182 4426 3194
rect 4442 3184 4457 3188
rect 4475 3185 4514 3204
rect 4533 3198 4540 3199
rect 4539 3191 4540 3198
rect 4523 3188 4524 3191
rect 4539 3188 4552 3191
rect 4475 3184 4505 3185
rect 4514 3184 4520 3185
rect 4523 3184 4552 3188
rect 4442 3183 4552 3184
rect 4442 3182 4558 3183
rect 4117 3174 4168 3182
rect 4117 3162 4142 3174
rect 4149 3162 4168 3174
rect 4199 3174 4249 3182
rect 4199 3166 4215 3174
rect 4222 3172 4249 3174
rect 4258 3172 4479 3182
rect 4222 3162 4479 3172
rect 4508 3174 4558 3182
rect 4508 3165 4524 3174
rect 4117 3154 4168 3162
rect 4215 3154 4479 3162
rect 4505 3162 4524 3165
rect 4531 3162 4558 3174
rect 4505 3154 4558 3162
rect 4133 3146 4134 3154
rect 4149 3146 4162 3154
rect 4133 3138 4149 3146
rect 4130 3131 4149 3134
rect 4130 3122 4152 3131
rect 4103 3112 4152 3122
rect 4103 3106 4133 3112
rect 4152 3107 4157 3112
rect 4075 3090 4149 3106
rect 4167 3098 4197 3154
rect 4232 3144 4440 3154
rect 4475 3150 4520 3154
rect 4523 3153 4524 3154
rect 4539 3153 4552 3154
rect 4258 3114 4447 3144
rect 4273 3111 4447 3114
rect 4266 3108 4447 3111
rect 4075 3088 4088 3090
rect 4103 3088 4137 3090
rect 4075 3072 4149 3088
rect 4176 3084 4189 3098
rect 4204 3084 4220 3100
rect 4266 3095 4277 3108
rect 4059 3050 4060 3066
rect 4075 3050 4088 3072
rect 4103 3050 4133 3072
rect 4176 3068 4238 3084
rect 4266 3077 4277 3093
rect 4282 3088 4292 3108
rect 4302 3088 4316 3108
rect 4319 3095 4328 3108
rect 4344 3095 4353 3108
rect 4282 3077 4316 3088
rect 4319 3077 4328 3093
rect 4344 3077 4353 3093
rect 4360 3088 4370 3108
rect 4380 3088 4394 3108
rect 4395 3095 4406 3108
rect 4360 3077 4394 3088
rect 4395 3077 4406 3093
rect 4452 3084 4468 3100
rect 4475 3098 4505 3150
rect 4539 3146 4540 3153
rect 4524 3138 4540 3146
rect 4511 3106 4524 3125
rect 4539 3106 4569 3122
rect 4511 3090 4585 3106
rect 4511 3088 4524 3090
rect 4539 3088 4573 3090
rect 4176 3066 4189 3068
rect 4204 3066 4238 3068
rect 4176 3050 4238 3066
rect 4282 3061 4298 3064
rect 4360 3061 4390 3072
rect 4438 3068 4484 3084
rect 4511 3072 4585 3088
rect 4438 3066 4472 3068
rect 4437 3050 4484 3066
rect 4511 3050 4524 3072
rect 4539 3050 4569 3072
rect 4596 3050 4597 3066
rect 4612 3050 4625 3210
rect 4655 3106 4668 3210
rect 4713 3188 4714 3198
rect 4729 3188 4742 3198
rect 4713 3184 4742 3188
rect 4747 3184 4777 3210
rect 4795 3196 4811 3198
rect 4883 3196 4936 3210
rect 4884 3194 4948 3196
rect 4991 3194 5006 3210
rect 5055 3207 5085 3210
rect 5055 3204 5091 3207
rect 5021 3196 5037 3198
rect 4795 3184 4810 3188
rect 4713 3182 4810 3184
rect 4838 3182 5006 3194
rect 5022 3184 5037 3188
rect 5055 3185 5094 3204
rect 5113 3198 5120 3199
rect 5119 3191 5120 3198
rect 5103 3188 5104 3191
rect 5119 3188 5132 3191
rect 5055 3184 5085 3185
rect 5094 3184 5100 3185
rect 5103 3184 5132 3188
rect 5022 3183 5132 3184
rect 5022 3182 5138 3183
rect 4697 3174 4748 3182
rect 4697 3162 4722 3174
rect 4729 3162 4748 3174
rect 4779 3174 4829 3182
rect 4779 3166 4795 3174
rect 4802 3172 4829 3174
rect 4838 3172 5059 3182
rect 4802 3162 5059 3172
rect 5088 3174 5138 3182
rect 5088 3165 5104 3174
rect 4697 3154 4748 3162
rect 4795 3154 5059 3162
rect 5085 3162 5104 3165
rect 5111 3162 5138 3174
rect 5085 3154 5138 3162
rect 4713 3146 4714 3154
rect 4729 3146 4742 3154
rect 4713 3138 4729 3146
rect 4710 3131 4729 3134
rect 4710 3122 4732 3131
rect 4683 3112 4732 3122
rect 4683 3106 4713 3112
rect 4732 3107 4737 3112
rect 4655 3090 4729 3106
rect 4747 3098 4777 3154
rect 4812 3144 5020 3154
rect 5055 3150 5100 3154
rect 5103 3153 5104 3154
rect 5119 3153 5132 3154
rect 4838 3114 5027 3144
rect 4853 3111 5027 3114
rect 4846 3108 5027 3111
rect 4655 3088 4668 3090
rect 4683 3088 4717 3090
rect 4655 3072 4729 3088
rect 4756 3084 4769 3098
rect 4784 3084 4800 3100
rect 4846 3095 4857 3108
rect 4639 3050 4640 3066
rect 4655 3050 4668 3072
rect 4683 3050 4713 3072
rect 4756 3068 4818 3084
rect 4846 3077 4857 3093
rect 4862 3088 4872 3108
rect 4882 3088 4896 3108
rect 4899 3095 4908 3108
rect 4924 3095 4933 3108
rect 4862 3077 4896 3088
rect 4899 3077 4908 3093
rect 4924 3077 4933 3093
rect 4940 3088 4950 3108
rect 4960 3088 4974 3108
rect 4975 3095 4986 3108
rect 4940 3077 4974 3088
rect 4975 3077 4986 3093
rect 5032 3084 5048 3100
rect 5055 3098 5085 3150
rect 5119 3146 5120 3153
rect 5104 3138 5120 3146
rect 5091 3106 5104 3125
rect 5119 3106 5149 3122
rect 5091 3090 5165 3106
rect 5091 3088 5104 3090
rect 5119 3088 5153 3090
rect 4756 3066 4769 3068
rect 4784 3066 4818 3068
rect 4756 3050 4818 3066
rect 4862 3061 4878 3064
rect 4940 3061 4970 3072
rect 5018 3068 5064 3084
rect 5091 3072 5165 3088
rect 5018 3066 5052 3068
rect 5017 3050 5064 3066
rect 5091 3050 5104 3072
rect 5119 3050 5149 3072
rect 5176 3050 5177 3066
rect 5192 3050 5205 3210
rect 5235 3106 5248 3210
rect 5293 3188 5294 3198
rect 5309 3188 5322 3198
rect 5293 3184 5322 3188
rect 5327 3184 5357 3210
rect 5375 3196 5391 3198
rect 5463 3196 5516 3210
rect 5464 3194 5528 3196
rect 5571 3194 5586 3210
rect 5635 3207 5665 3210
rect 5635 3204 5671 3207
rect 5601 3196 5617 3198
rect 5375 3184 5390 3188
rect 5293 3182 5390 3184
rect 5418 3182 5586 3194
rect 5602 3184 5617 3188
rect 5635 3185 5674 3204
rect 5693 3198 5700 3199
rect 5699 3191 5700 3198
rect 5683 3188 5684 3191
rect 5699 3188 5712 3191
rect 5635 3184 5665 3185
rect 5674 3184 5680 3185
rect 5683 3184 5712 3188
rect 5602 3183 5712 3184
rect 5602 3182 5718 3183
rect 5277 3174 5328 3182
rect 5277 3162 5302 3174
rect 5309 3162 5328 3174
rect 5359 3174 5409 3182
rect 5359 3166 5375 3174
rect 5382 3172 5409 3174
rect 5418 3172 5639 3182
rect 5382 3162 5639 3172
rect 5668 3174 5718 3182
rect 5668 3165 5684 3174
rect 5277 3154 5328 3162
rect 5375 3154 5639 3162
rect 5665 3162 5684 3165
rect 5691 3162 5718 3174
rect 5665 3154 5718 3162
rect 5293 3146 5294 3154
rect 5309 3146 5322 3154
rect 5293 3138 5309 3146
rect 5290 3131 5309 3134
rect 5290 3122 5312 3131
rect 5263 3112 5312 3122
rect 5263 3106 5293 3112
rect 5312 3107 5317 3112
rect 5235 3090 5309 3106
rect 5327 3098 5357 3154
rect 5392 3144 5600 3154
rect 5635 3150 5680 3154
rect 5683 3153 5684 3154
rect 5699 3153 5712 3154
rect 5418 3114 5607 3144
rect 5433 3111 5607 3114
rect 5426 3108 5607 3111
rect 5235 3088 5248 3090
rect 5263 3088 5297 3090
rect 5235 3072 5309 3088
rect 5336 3084 5349 3098
rect 5364 3084 5380 3100
rect 5426 3095 5437 3108
rect 5219 3050 5220 3066
rect 5235 3050 5248 3072
rect 5263 3050 5293 3072
rect 5336 3068 5398 3084
rect 5426 3077 5437 3093
rect 5442 3088 5452 3108
rect 5462 3088 5476 3108
rect 5479 3095 5488 3108
rect 5504 3095 5513 3108
rect 5442 3077 5476 3088
rect 5479 3077 5488 3093
rect 5504 3077 5513 3093
rect 5520 3088 5530 3108
rect 5540 3088 5554 3108
rect 5555 3095 5566 3108
rect 5520 3077 5554 3088
rect 5555 3077 5566 3093
rect 5612 3084 5628 3100
rect 5635 3098 5665 3150
rect 5699 3146 5700 3153
rect 5684 3138 5700 3146
rect 5671 3106 5684 3125
rect 5699 3106 5729 3122
rect 5671 3090 5745 3106
rect 5671 3088 5684 3090
rect 5699 3088 5733 3090
rect 5336 3066 5349 3068
rect 5364 3066 5398 3068
rect 5336 3050 5398 3066
rect 5442 3061 5458 3064
rect 5520 3061 5550 3072
rect 5598 3068 5644 3084
rect 5671 3072 5745 3088
rect 5598 3066 5632 3068
rect 5597 3050 5644 3066
rect 5671 3050 5684 3072
rect 5699 3050 5729 3072
rect 5756 3050 5757 3066
rect 5772 3050 5785 3210
rect 5815 3106 5828 3210
rect 5873 3188 5874 3198
rect 5889 3188 5902 3198
rect 5873 3184 5902 3188
rect 5907 3184 5937 3210
rect 5955 3196 5971 3198
rect 6043 3196 6096 3210
rect 6044 3194 6108 3196
rect 6151 3194 6166 3210
rect 6215 3207 6245 3210
rect 6215 3204 6251 3207
rect 6181 3196 6197 3198
rect 5955 3184 5970 3188
rect 5873 3182 5970 3184
rect 5998 3182 6166 3194
rect 6182 3184 6197 3188
rect 6215 3185 6254 3204
rect 6273 3198 6280 3199
rect 6279 3191 6280 3198
rect 6263 3188 6264 3191
rect 6279 3188 6292 3191
rect 6215 3184 6245 3185
rect 6254 3184 6260 3185
rect 6263 3184 6292 3188
rect 6182 3183 6292 3184
rect 6182 3182 6298 3183
rect 5857 3174 5908 3182
rect 5857 3162 5882 3174
rect 5889 3162 5908 3174
rect 5939 3174 5989 3182
rect 5939 3166 5955 3174
rect 5962 3172 5989 3174
rect 5998 3172 6219 3182
rect 5962 3162 6219 3172
rect 6248 3174 6298 3182
rect 6248 3165 6264 3174
rect 5857 3154 5908 3162
rect 5955 3154 6219 3162
rect 6245 3162 6264 3165
rect 6271 3162 6298 3174
rect 6245 3154 6298 3162
rect 5873 3146 5874 3154
rect 5889 3146 5902 3154
rect 5873 3138 5889 3146
rect 5870 3131 5889 3134
rect 5870 3122 5892 3131
rect 5843 3112 5892 3122
rect 5843 3106 5873 3112
rect 5892 3107 5897 3112
rect 5815 3090 5889 3106
rect 5907 3098 5937 3154
rect 5972 3144 6180 3154
rect 6215 3150 6260 3154
rect 6263 3153 6264 3154
rect 6279 3153 6292 3154
rect 5998 3114 6187 3144
rect 6013 3111 6187 3114
rect 6006 3108 6187 3111
rect 5815 3088 5828 3090
rect 5843 3088 5877 3090
rect 5815 3072 5889 3088
rect 5916 3084 5929 3098
rect 5944 3084 5960 3100
rect 6006 3095 6017 3108
rect 5799 3050 5800 3066
rect 5815 3050 5828 3072
rect 5843 3050 5873 3072
rect 5916 3068 5978 3084
rect 6006 3077 6017 3093
rect 6022 3088 6032 3108
rect 6042 3088 6056 3108
rect 6059 3095 6068 3108
rect 6084 3095 6093 3108
rect 6022 3077 6056 3088
rect 6059 3077 6068 3093
rect 6084 3077 6093 3093
rect 6100 3088 6110 3108
rect 6120 3088 6134 3108
rect 6135 3095 6146 3108
rect 6100 3077 6134 3088
rect 6135 3077 6146 3093
rect 6192 3084 6208 3100
rect 6215 3098 6245 3150
rect 6279 3146 6280 3153
rect 6264 3138 6280 3146
rect 6251 3106 6264 3125
rect 6279 3106 6309 3122
rect 6251 3090 6325 3106
rect 6251 3088 6264 3090
rect 6279 3088 6313 3090
rect 5916 3066 5929 3068
rect 5944 3066 5978 3068
rect 5916 3050 5978 3066
rect 6022 3061 6038 3064
rect 6100 3061 6130 3072
rect 6178 3068 6224 3084
rect 6251 3072 6325 3088
rect 6178 3066 6212 3068
rect 6177 3050 6224 3066
rect 6251 3050 6264 3072
rect 6279 3050 6309 3072
rect 6336 3050 6337 3066
rect 6352 3050 6365 3210
rect 6395 3106 6408 3210
rect 6453 3188 6454 3198
rect 6469 3188 6482 3198
rect 6453 3184 6482 3188
rect 6487 3184 6517 3210
rect 6535 3196 6551 3198
rect 6623 3196 6676 3210
rect 6624 3194 6688 3196
rect 6731 3194 6746 3210
rect 6795 3207 6825 3210
rect 6795 3204 6831 3207
rect 6761 3196 6777 3198
rect 6535 3184 6550 3188
rect 6453 3182 6550 3184
rect 6578 3182 6746 3194
rect 6762 3184 6777 3188
rect 6795 3185 6834 3204
rect 6853 3198 6860 3199
rect 6859 3191 6860 3198
rect 6843 3188 6844 3191
rect 6859 3188 6872 3191
rect 6795 3184 6825 3185
rect 6834 3184 6840 3185
rect 6843 3184 6872 3188
rect 6762 3183 6872 3184
rect 6762 3182 6878 3183
rect 6437 3174 6488 3182
rect 6437 3162 6462 3174
rect 6469 3162 6488 3174
rect 6519 3174 6569 3182
rect 6519 3166 6535 3174
rect 6542 3172 6569 3174
rect 6578 3172 6799 3182
rect 6542 3162 6799 3172
rect 6828 3174 6878 3182
rect 6828 3165 6844 3174
rect 6437 3154 6488 3162
rect 6535 3154 6799 3162
rect 6825 3162 6844 3165
rect 6851 3162 6878 3174
rect 6825 3154 6878 3162
rect 6453 3146 6454 3154
rect 6469 3146 6482 3154
rect 6453 3138 6469 3146
rect 6450 3131 6469 3134
rect 6450 3122 6472 3131
rect 6423 3112 6472 3122
rect 6423 3106 6453 3112
rect 6472 3107 6477 3112
rect 6395 3090 6469 3106
rect 6487 3098 6517 3154
rect 6552 3144 6760 3154
rect 6795 3150 6840 3154
rect 6843 3153 6844 3154
rect 6859 3153 6872 3154
rect 6578 3114 6767 3144
rect 6593 3111 6767 3114
rect 6586 3108 6767 3111
rect 6395 3088 6408 3090
rect 6423 3088 6457 3090
rect 6395 3072 6469 3088
rect 6496 3084 6509 3098
rect 6524 3084 6540 3100
rect 6586 3095 6597 3108
rect 6379 3050 6380 3066
rect 6395 3050 6408 3072
rect 6423 3050 6453 3072
rect 6496 3068 6558 3084
rect 6586 3077 6597 3093
rect 6602 3088 6612 3108
rect 6622 3088 6636 3108
rect 6639 3095 6648 3108
rect 6664 3095 6673 3108
rect 6602 3077 6636 3088
rect 6639 3077 6648 3093
rect 6664 3077 6673 3093
rect 6680 3088 6690 3108
rect 6700 3088 6714 3108
rect 6715 3095 6726 3108
rect 6680 3077 6714 3088
rect 6715 3077 6726 3093
rect 6772 3084 6788 3100
rect 6795 3098 6825 3150
rect 6859 3146 6860 3153
rect 6844 3138 6860 3146
rect 6831 3106 6844 3125
rect 6859 3106 6889 3122
rect 6831 3090 6905 3106
rect 6831 3088 6844 3090
rect 6859 3088 6893 3090
rect 6496 3066 6509 3068
rect 6524 3066 6558 3068
rect 6496 3050 6558 3066
rect 6602 3061 6618 3064
rect 6680 3061 6710 3072
rect 6758 3068 6804 3084
rect 6831 3072 6905 3088
rect 6758 3066 6792 3068
rect 6757 3050 6804 3066
rect 6831 3050 6844 3072
rect 6859 3050 6889 3072
rect 6916 3050 6917 3066
rect 6932 3050 6945 3210
rect 6975 3106 6988 3210
rect 7033 3188 7034 3198
rect 7049 3188 7062 3198
rect 7033 3184 7062 3188
rect 7067 3184 7097 3210
rect 7115 3196 7131 3198
rect 7203 3196 7256 3210
rect 7204 3194 7268 3196
rect 7311 3194 7326 3210
rect 7375 3207 7405 3210
rect 7375 3204 7411 3207
rect 7341 3196 7357 3198
rect 7115 3184 7130 3188
rect 7033 3182 7130 3184
rect 7158 3182 7326 3194
rect 7342 3184 7357 3188
rect 7375 3185 7414 3204
rect 7433 3198 7440 3199
rect 7439 3191 7440 3198
rect 7423 3188 7424 3191
rect 7439 3188 7452 3191
rect 7375 3184 7405 3185
rect 7414 3184 7420 3185
rect 7423 3184 7452 3188
rect 7342 3183 7452 3184
rect 7342 3182 7458 3183
rect 7017 3174 7068 3182
rect 7017 3162 7042 3174
rect 7049 3162 7068 3174
rect 7099 3174 7149 3182
rect 7099 3166 7115 3174
rect 7122 3172 7149 3174
rect 7158 3172 7379 3182
rect 7122 3162 7379 3172
rect 7408 3174 7458 3182
rect 7408 3165 7424 3174
rect 7017 3154 7068 3162
rect 7115 3154 7379 3162
rect 7405 3162 7424 3165
rect 7431 3162 7458 3174
rect 7405 3154 7458 3162
rect 7033 3146 7034 3154
rect 7049 3146 7062 3154
rect 7033 3138 7049 3146
rect 7030 3131 7049 3134
rect 7030 3122 7052 3131
rect 7003 3112 7052 3122
rect 7003 3106 7033 3112
rect 7052 3107 7057 3112
rect 6975 3090 7049 3106
rect 7067 3098 7097 3154
rect 7132 3144 7340 3154
rect 7375 3150 7420 3154
rect 7423 3153 7424 3154
rect 7439 3153 7452 3154
rect 7158 3114 7347 3144
rect 7173 3111 7347 3114
rect 7166 3108 7347 3111
rect 6975 3088 6988 3090
rect 7003 3088 7037 3090
rect 6975 3072 7049 3088
rect 7076 3084 7089 3098
rect 7104 3084 7120 3100
rect 7166 3095 7177 3108
rect 6959 3050 6960 3066
rect 6975 3050 6988 3072
rect 7003 3050 7033 3072
rect 7076 3068 7138 3084
rect 7166 3077 7177 3093
rect 7182 3088 7192 3108
rect 7202 3088 7216 3108
rect 7219 3095 7228 3108
rect 7244 3095 7253 3108
rect 7182 3077 7216 3088
rect 7219 3077 7228 3093
rect 7244 3077 7253 3093
rect 7260 3088 7270 3108
rect 7280 3088 7294 3108
rect 7295 3095 7306 3108
rect 7260 3077 7294 3088
rect 7295 3077 7306 3093
rect 7352 3084 7368 3100
rect 7375 3098 7405 3150
rect 7439 3146 7440 3153
rect 7424 3138 7440 3146
rect 7411 3106 7424 3125
rect 7439 3106 7469 3122
rect 7411 3090 7485 3106
rect 7411 3088 7424 3090
rect 7439 3088 7473 3090
rect 7076 3066 7089 3068
rect 7104 3066 7138 3068
rect 7076 3050 7138 3066
rect 7182 3061 7198 3064
rect 7260 3061 7290 3072
rect 7338 3068 7384 3084
rect 7411 3072 7485 3088
rect 7338 3066 7372 3068
rect 7337 3050 7384 3066
rect 7411 3050 7424 3072
rect 7439 3050 7469 3072
rect 7496 3050 7497 3066
rect 7512 3050 7525 3210
rect 7555 3106 7568 3210
rect 7613 3188 7614 3198
rect 7629 3188 7642 3198
rect 7613 3184 7642 3188
rect 7647 3184 7677 3210
rect 7695 3196 7711 3198
rect 7783 3196 7836 3210
rect 7784 3194 7848 3196
rect 7891 3194 7906 3210
rect 7955 3207 7985 3210
rect 7955 3204 7991 3207
rect 7921 3196 7937 3198
rect 7695 3184 7710 3188
rect 7613 3182 7710 3184
rect 7738 3182 7906 3194
rect 7922 3184 7937 3188
rect 7955 3185 7994 3204
rect 8013 3198 8020 3199
rect 8019 3191 8020 3198
rect 8003 3188 8004 3191
rect 8019 3188 8032 3191
rect 7955 3184 7985 3185
rect 7994 3184 8000 3185
rect 8003 3184 8032 3188
rect 7922 3183 8032 3184
rect 7922 3182 8038 3183
rect 7597 3174 7648 3182
rect 7597 3162 7622 3174
rect 7629 3162 7648 3174
rect 7679 3174 7729 3182
rect 7679 3166 7695 3174
rect 7702 3172 7729 3174
rect 7738 3172 7959 3182
rect 7702 3162 7959 3172
rect 7988 3174 8038 3182
rect 7988 3165 8004 3174
rect 7597 3154 7648 3162
rect 7695 3154 7959 3162
rect 7985 3162 8004 3165
rect 8011 3162 8038 3174
rect 7985 3154 8038 3162
rect 7613 3146 7614 3154
rect 7629 3146 7642 3154
rect 7613 3138 7629 3146
rect 7610 3131 7629 3134
rect 7610 3122 7632 3131
rect 7583 3112 7632 3122
rect 7583 3106 7613 3112
rect 7632 3107 7637 3112
rect 7555 3090 7629 3106
rect 7647 3098 7677 3154
rect 7712 3144 7920 3154
rect 7955 3150 8000 3154
rect 8003 3153 8004 3154
rect 8019 3153 8032 3154
rect 7738 3114 7927 3144
rect 7753 3111 7927 3114
rect 7746 3108 7927 3111
rect 7555 3088 7568 3090
rect 7583 3088 7617 3090
rect 7555 3072 7629 3088
rect 7656 3084 7669 3098
rect 7684 3084 7700 3100
rect 7746 3095 7757 3108
rect 7539 3050 7540 3066
rect 7555 3050 7568 3072
rect 7583 3050 7613 3072
rect 7656 3068 7718 3084
rect 7746 3077 7757 3093
rect 7762 3088 7772 3108
rect 7782 3088 7796 3108
rect 7799 3095 7808 3108
rect 7824 3095 7833 3108
rect 7762 3077 7796 3088
rect 7799 3077 7808 3093
rect 7824 3077 7833 3093
rect 7840 3088 7850 3108
rect 7860 3088 7874 3108
rect 7875 3095 7886 3108
rect 7840 3077 7874 3088
rect 7875 3077 7886 3093
rect 7932 3084 7948 3100
rect 7955 3098 7985 3150
rect 8019 3146 8020 3153
rect 8004 3138 8020 3146
rect 7991 3106 8004 3125
rect 8019 3106 8049 3122
rect 7991 3090 8065 3106
rect 7991 3088 8004 3090
rect 8019 3088 8053 3090
rect 7656 3066 7669 3068
rect 7684 3066 7718 3068
rect 7656 3050 7718 3066
rect 7762 3061 7778 3064
rect 7840 3061 7870 3072
rect 7918 3068 7964 3084
rect 7991 3072 8065 3088
rect 7918 3066 7952 3068
rect 7917 3050 7964 3066
rect 7991 3050 8004 3072
rect 8019 3050 8049 3072
rect 8076 3050 8077 3066
rect 8092 3050 8105 3210
rect 8135 3106 8148 3210
rect 8193 3188 8194 3198
rect 8209 3188 8222 3198
rect 8193 3184 8222 3188
rect 8227 3184 8257 3210
rect 8275 3196 8291 3198
rect 8363 3196 8416 3210
rect 8364 3194 8428 3196
rect 8471 3194 8486 3210
rect 8535 3207 8565 3210
rect 8535 3204 8571 3207
rect 8501 3196 8517 3198
rect 8275 3184 8290 3188
rect 8193 3182 8290 3184
rect 8318 3182 8486 3194
rect 8502 3184 8517 3188
rect 8535 3185 8574 3204
rect 8593 3198 8600 3199
rect 8599 3191 8600 3198
rect 8583 3188 8584 3191
rect 8599 3188 8612 3191
rect 8535 3184 8565 3185
rect 8574 3184 8580 3185
rect 8583 3184 8612 3188
rect 8502 3183 8612 3184
rect 8502 3182 8618 3183
rect 8177 3174 8228 3182
rect 8177 3162 8202 3174
rect 8209 3162 8228 3174
rect 8259 3174 8309 3182
rect 8259 3166 8275 3174
rect 8282 3172 8309 3174
rect 8318 3172 8539 3182
rect 8282 3162 8539 3172
rect 8568 3174 8618 3182
rect 8568 3165 8584 3174
rect 8177 3154 8228 3162
rect 8275 3154 8539 3162
rect 8565 3162 8584 3165
rect 8591 3162 8618 3174
rect 8565 3154 8618 3162
rect 8193 3146 8194 3154
rect 8209 3146 8222 3154
rect 8193 3138 8209 3146
rect 8190 3131 8209 3134
rect 8190 3122 8212 3131
rect 8163 3112 8212 3122
rect 8163 3106 8193 3112
rect 8212 3107 8217 3112
rect 8135 3090 8209 3106
rect 8227 3098 8257 3154
rect 8292 3144 8500 3154
rect 8535 3150 8580 3154
rect 8583 3153 8584 3154
rect 8599 3153 8612 3154
rect 8318 3114 8507 3144
rect 8333 3111 8507 3114
rect 8326 3108 8507 3111
rect 8135 3088 8148 3090
rect 8163 3088 8197 3090
rect 8135 3072 8209 3088
rect 8236 3084 8249 3098
rect 8264 3084 8280 3100
rect 8326 3095 8337 3108
rect 8119 3050 8120 3066
rect 8135 3050 8148 3072
rect 8163 3050 8193 3072
rect 8236 3068 8298 3084
rect 8326 3077 8337 3093
rect 8342 3088 8352 3108
rect 8362 3088 8376 3108
rect 8379 3095 8388 3108
rect 8404 3095 8413 3108
rect 8342 3077 8376 3088
rect 8379 3077 8388 3093
rect 8404 3077 8413 3093
rect 8420 3088 8430 3108
rect 8440 3088 8454 3108
rect 8455 3095 8466 3108
rect 8420 3077 8454 3088
rect 8455 3077 8466 3093
rect 8512 3084 8528 3100
rect 8535 3098 8565 3150
rect 8599 3146 8600 3153
rect 8584 3138 8600 3146
rect 8571 3106 8584 3125
rect 8599 3106 8629 3122
rect 8571 3090 8645 3106
rect 8571 3088 8584 3090
rect 8599 3088 8633 3090
rect 8236 3066 8249 3068
rect 8264 3066 8298 3068
rect 8236 3050 8298 3066
rect 8342 3061 8358 3064
rect 8420 3061 8450 3072
rect 8498 3068 8544 3084
rect 8571 3072 8645 3088
rect 8498 3066 8532 3068
rect 8497 3050 8544 3066
rect 8571 3050 8584 3072
rect 8599 3050 8629 3072
rect 8656 3050 8657 3066
rect 8672 3050 8685 3210
rect 8715 3106 8728 3210
rect 8773 3188 8774 3198
rect 8789 3188 8802 3198
rect 8773 3184 8802 3188
rect 8807 3184 8837 3210
rect 8855 3196 8871 3198
rect 8943 3196 8996 3210
rect 8944 3194 9008 3196
rect 9051 3194 9066 3210
rect 9115 3207 9145 3210
rect 9115 3204 9151 3207
rect 9081 3196 9097 3198
rect 8855 3184 8870 3188
rect 8773 3182 8870 3184
rect 8898 3182 9066 3194
rect 9082 3184 9097 3188
rect 9115 3185 9154 3204
rect 9173 3198 9180 3199
rect 9179 3191 9180 3198
rect 9163 3188 9164 3191
rect 9179 3188 9192 3191
rect 9115 3184 9145 3185
rect 9154 3184 9160 3185
rect 9163 3184 9192 3188
rect 9082 3183 9192 3184
rect 9082 3182 9198 3183
rect 8757 3174 8808 3182
rect 8757 3162 8782 3174
rect 8789 3162 8808 3174
rect 8839 3174 8889 3182
rect 8839 3166 8855 3174
rect 8862 3172 8889 3174
rect 8898 3172 9119 3182
rect 8862 3162 9119 3172
rect 9148 3174 9198 3182
rect 9148 3165 9164 3174
rect 8757 3154 8808 3162
rect 8855 3154 9119 3162
rect 9145 3162 9164 3165
rect 9171 3162 9198 3174
rect 9145 3154 9198 3162
rect 8773 3146 8774 3154
rect 8789 3146 8802 3154
rect 8773 3138 8789 3146
rect 8770 3131 8789 3134
rect 8770 3122 8792 3131
rect 8743 3112 8792 3122
rect 8743 3106 8773 3112
rect 8792 3107 8797 3112
rect 8715 3090 8789 3106
rect 8807 3098 8837 3154
rect 8872 3144 9080 3154
rect 9115 3150 9160 3154
rect 9163 3153 9164 3154
rect 9179 3153 9192 3154
rect 8898 3114 9087 3144
rect 8913 3111 9087 3114
rect 8906 3108 9087 3111
rect 8715 3088 8728 3090
rect 8743 3088 8777 3090
rect 8715 3072 8789 3088
rect 8816 3084 8829 3098
rect 8844 3084 8860 3100
rect 8906 3095 8917 3108
rect 8699 3050 8700 3066
rect 8715 3050 8728 3072
rect 8743 3050 8773 3072
rect 8816 3068 8878 3084
rect 8906 3077 8917 3093
rect 8922 3088 8932 3108
rect 8942 3088 8956 3108
rect 8959 3095 8968 3108
rect 8984 3095 8993 3108
rect 8922 3077 8956 3088
rect 8959 3077 8968 3093
rect 8984 3077 8993 3093
rect 9000 3088 9010 3108
rect 9020 3088 9034 3108
rect 9035 3095 9046 3108
rect 9000 3077 9034 3088
rect 9035 3077 9046 3093
rect 9092 3084 9108 3100
rect 9115 3098 9145 3150
rect 9179 3146 9180 3153
rect 9164 3138 9180 3146
rect 9151 3106 9164 3125
rect 9179 3106 9209 3122
rect 9151 3090 9225 3106
rect 9151 3088 9164 3090
rect 9179 3088 9213 3090
rect 8816 3066 8829 3068
rect 8844 3066 8878 3068
rect 8816 3050 8878 3066
rect 8922 3061 8938 3064
rect 9000 3061 9030 3072
rect 9078 3068 9124 3084
rect 9151 3072 9225 3088
rect 9078 3066 9112 3068
rect 9077 3050 9124 3066
rect 9151 3050 9164 3072
rect 9179 3050 9209 3072
rect 9236 3050 9237 3066
rect 9252 3050 9265 3210
rect -7 3042 34 3050
rect -7 3016 8 3042
rect 15 3016 34 3042
rect 98 3038 160 3050
rect 172 3038 247 3050
rect 305 3038 380 3050
rect 392 3038 423 3050
rect 429 3038 464 3050
rect 98 3036 260 3038
rect -7 3008 34 3016
rect 116 3012 129 3036
rect 144 3034 159 3036
rect -1 2998 0 3008
rect 15 2998 28 3008
rect 43 2998 73 3012
rect 116 2998 159 3012
rect 183 3009 190 3016
rect 193 3012 260 3036
rect 292 3036 464 3038
rect 262 3014 290 3018
rect 292 3014 372 3036
rect 393 3034 408 3036
rect 262 3012 372 3014
rect 193 3008 372 3012
rect 166 2998 196 3008
rect 198 2998 351 3008
rect 359 2998 389 3008
rect 393 2998 423 3012
rect 451 2998 464 3036
rect 536 3042 571 3050
rect 536 3016 537 3042
rect 544 3016 571 3042
rect 479 2998 509 3012
rect 536 3008 571 3016
rect 573 3042 614 3050
rect 573 3016 588 3042
rect 595 3016 614 3042
rect 678 3038 740 3050
rect 752 3038 827 3050
rect 885 3038 960 3050
rect 972 3038 1003 3050
rect 1009 3038 1044 3050
rect 678 3036 840 3038
rect 573 3008 614 3016
rect 696 3012 709 3036
rect 724 3034 739 3036
rect 536 2998 537 3008
rect 552 2998 565 3008
rect 579 2998 580 3008
rect 595 2998 608 3008
rect 623 2998 653 3012
rect 696 2998 739 3012
rect 763 3009 770 3016
rect 773 3012 840 3036
rect 872 3036 1044 3038
rect 842 3014 870 3018
rect 872 3014 952 3036
rect 973 3034 988 3036
rect 842 3012 952 3014
rect 773 3008 952 3012
rect 746 2998 776 3008
rect 778 2998 931 3008
rect 939 2998 969 3008
rect 973 2998 1003 3012
rect 1031 2998 1044 3036
rect 1116 3042 1151 3050
rect 1116 3016 1117 3042
rect 1124 3016 1151 3042
rect 1059 2998 1089 3012
rect 1116 3008 1151 3016
rect 1153 3042 1194 3050
rect 1153 3016 1168 3042
rect 1175 3016 1194 3042
rect 1258 3038 1320 3050
rect 1332 3038 1407 3050
rect 1465 3038 1540 3050
rect 1552 3038 1583 3050
rect 1589 3038 1624 3050
rect 1258 3036 1420 3038
rect 1153 3008 1194 3016
rect 1276 3012 1289 3036
rect 1304 3034 1319 3036
rect 1116 2998 1117 3008
rect 1132 2998 1145 3008
rect 1159 2998 1160 3008
rect 1175 2998 1188 3008
rect 1203 2998 1233 3012
rect 1276 2998 1319 3012
rect 1343 3009 1350 3016
rect 1353 3012 1420 3036
rect 1452 3036 1624 3038
rect 1422 3014 1450 3018
rect 1452 3014 1532 3036
rect 1553 3034 1568 3036
rect 1422 3012 1532 3014
rect 1353 3008 1532 3012
rect 1326 2998 1356 3008
rect 1358 2998 1511 3008
rect 1519 2998 1549 3008
rect 1553 2998 1583 3012
rect 1611 2998 1624 3036
rect 1696 3042 1731 3050
rect 1696 3016 1697 3042
rect 1704 3016 1731 3042
rect 1639 2998 1669 3012
rect 1696 3008 1731 3016
rect 1733 3042 1774 3050
rect 1733 3016 1748 3042
rect 1755 3016 1774 3042
rect 1838 3038 1900 3050
rect 1912 3038 1987 3050
rect 2045 3038 2120 3050
rect 2132 3038 2163 3050
rect 2169 3038 2204 3050
rect 1838 3036 2000 3038
rect 1733 3008 1774 3016
rect 1856 3012 1869 3036
rect 1884 3034 1899 3036
rect 1696 2998 1697 3008
rect 1712 2998 1725 3008
rect 1739 2998 1740 3008
rect 1755 2998 1768 3008
rect 1783 2998 1813 3012
rect 1856 2998 1899 3012
rect 1923 3009 1930 3016
rect 1933 3012 2000 3036
rect 2032 3036 2204 3038
rect 2002 3014 2030 3018
rect 2032 3014 2112 3036
rect 2133 3034 2148 3036
rect 2002 3012 2112 3014
rect 1933 3008 2112 3012
rect 1906 2998 1936 3008
rect 1938 2998 2091 3008
rect 2099 2998 2129 3008
rect 2133 2998 2163 3012
rect 2191 2998 2204 3036
rect 2276 3042 2311 3050
rect 2276 3016 2277 3042
rect 2284 3016 2311 3042
rect 2219 2998 2249 3012
rect 2276 3008 2311 3016
rect 2313 3042 2354 3050
rect 2313 3016 2328 3042
rect 2335 3016 2354 3042
rect 2418 3038 2480 3050
rect 2492 3038 2567 3050
rect 2625 3038 2700 3050
rect 2712 3038 2743 3050
rect 2749 3038 2784 3050
rect 2418 3036 2580 3038
rect 2313 3008 2354 3016
rect 2436 3012 2449 3036
rect 2464 3034 2479 3036
rect 2276 2998 2277 3008
rect 2292 2998 2305 3008
rect 2319 2998 2320 3008
rect 2335 2998 2348 3008
rect 2363 2998 2393 3012
rect 2436 2998 2479 3012
rect 2503 3009 2510 3016
rect 2513 3012 2580 3036
rect 2612 3036 2784 3038
rect 2582 3014 2610 3018
rect 2612 3014 2692 3036
rect 2713 3034 2728 3036
rect 2582 3012 2692 3014
rect 2513 3008 2692 3012
rect 2486 2998 2516 3008
rect 2518 2998 2671 3008
rect 2679 2998 2709 3008
rect 2713 2998 2743 3012
rect 2771 2998 2784 3036
rect 2856 3042 2891 3050
rect 2856 3016 2857 3042
rect 2864 3016 2891 3042
rect 2799 2998 2829 3012
rect 2856 3008 2891 3016
rect 2893 3042 2934 3050
rect 2893 3016 2908 3042
rect 2915 3016 2934 3042
rect 2998 3038 3060 3050
rect 3072 3038 3147 3050
rect 3205 3038 3280 3050
rect 3292 3038 3323 3050
rect 3329 3038 3364 3050
rect 2998 3036 3160 3038
rect 2893 3008 2934 3016
rect 3016 3012 3029 3036
rect 3044 3034 3059 3036
rect 2856 2998 2857 3008
rect 2872 2998 2885 3008
rect 2899 2998 2900 3008
rect 2915 2998 2928 3008
rect 2943 2998 2973 3012
rect 3016 2998 3059 3012
rect 3083 3009 3090 3016
rect 3093 3012 3160 3036
rect 3192 3036 3364 3038
rect 3162 3014 3190 3018
rect 3192 3014 3272 3036
rect 3293 3034 3308 3036
rect 3162 3012 3272 3014
rect 3093 3008 3272 3012
rect 3066 2998 3096 3008
rect 3098 2998 3251 3008
rect 3259 2998 3289 3008
rect 3293 2998 3323 3012
rect 3351 2998 3364 3036
rect 3436 3042 3471 3050
rect 3436 3016 3437 3042
rect 3444 3016 3471 3042
rect 3379 2998 3409 3012
rect 3436 3008 3471 3016
rect 3473 3042 3514 3050
rect 3473 3016 3488 3042
rect 3495 3016 3514 3042
rect 3578 3038 3640 3050
rect 3652 3038 3727 3050
rect 3785 3038 3860 3050
rect 3872 3038 3903 3050
rect 3909 3038 3944 3050
rect 3578 3036 3740 3038
rect 3473 3008 3514 3016
rect 3596 3012 3609 3036
rect 3624 3034 3639 3036
rect 3436 2998 3437 3008
rect 3452 2998 3465 3008
rect 3479 2998 3480 3008
rect 3495 2998 3508 3008
rect 3523 2998 3553 3012
rect 3596 2998 3639 3012
rect 3663 3009 3670 3016
rect 3673 3012 3740 3036
rect 3772 3036 3944 3038
rect 3742 3014 3770 3018
rect 3772 3014 3852 3036
rect 3873 3034 3888 3036
rect 3742 3012 3852 3014
rect 3673 3008 3852 3012
rect 3646 2998 3676 3008
rect 3678 2998 3831 3008
rect 3839 2998 3869 3008
rect 3873 2998 3903 3012
rect 3931 2998 3944 3036
rect 4016 3042 4051 3050
rect 4016 3016 4017 3042
rect 4024 3016 4051 3042
rect 3959 2998 3989 3012
rect 4016 3008 4051 3016
rect 4053 3042 4094 3050
rect 4053 3016 4068 3042
rect 4075 3016 4094 3042
rect 4158 3038 4220 3050
rect 4232 3038 4307 3050
rect 4365 3038 4440 3050
rect 4452 3038 4483 3050
rect 4489 3038 4524 3050
rect 4158 3036 4320 3038
rect 4053 3008 4094 3016
rect 4176 3012 4189 3036
rect 4204 3034 4219 3036
rect 4016 2998 4017 3008
rect 4032 2998 4045 3008
rect 4059 2998 4060 3008
rect 4075 2998 4088 3008
rect 4103 2998 4133 3012
rect 4176 2998 4219 3012
rect 4243 3009 4250 3016
rect 4253 3012 4320 3036
rect 4352 3036 4524 3038
rect 4322 3014 4350 3018
rect 4352 3014 4432 3036
rect 4453 3034 4468 3036
rect 4322 3012 4432 3014
rect 4253 3008 4432 3012
rect 4226 2998 4256 3008
rect 4258 2998 4411 3008
rect 4419 2998 4449 3008
rect 4453 2998 4483 3012
rect 4511 2998 4524 3036
rect 4596 3042 4631 3050
rect 4596 3016 4597 3042
rect 4604 3016 4631 3042
rect 4539 2998 4569 3012
rect 4596 3008 4631 3016
rect 4633 3042 4674 3050
rect 4633 3016 4648 3042
rect 4655 3016 4674 3042
rect 4738 3038 4800 3050
rect 4812 3038 4887 3050
rect 4945 3038 5020 3050
rect 5032 3038 5063 3050
rect 5069 3038 5104 3050
rect 4738 3036 4900 3038
rect 4633 3008 4674 3016
rect 4756 3012 4769 3036
rect 4784 3034 4799 3036
rect 4596 2998 4597 3008
rect 4612 2998 4625 3008
rect 4639 2998 4640 3008
rect 4655 2998 4668 3008
rect 4683 2998 4713 3012
rect 4756 2998 4799 3012
rect 4823 3009 4830 3016
rect 4833 3012 4900 3036
rect 4932 3036 5104 3038
rect 4902 3014 4930 3018
rect 4932 3014 5012 3036
rect 5033 3034 5048 3036
rect 4902 3012 5012 3014
rect 4833 3008 5012 3012
rect 4806 2998 4836 3008
rect 4838 2998 4991 3008
rect 4999 2998 5029 3008
rect 5033 2998 5063 3012
rect 5091 2998 5104 3036
rect 5176 3042 5211 3050
rect 5176 3016 5177 3042
rect 5184 3016 5211 3042
rect 5119 2998 5149 3012
rect 5176 3008 5211 3016
rect 5213 3042 5254 3050
rect 5213 3016 5228 3042
rect 5235 3016 5254 3042
rect 5318 3038 5380 3050
rect 5392 3038 5467 3050
rect 5525 3038 5600 3050
rect 5612 3038 5643 3050
rect 5649 3038 5684 3050
rect 5318 3036 5480 3038
rect 5213 3008 5254 3016
rect 5336 3012 5349 3036
rect 5364 3034 5379 3036
rect 5176 2998 5177 3008
rect 5192 2998 5205 3008
rect 5219 2998 5220 3008
rect 5235 2998 5248 3008
rect 5263 2998 5293 3012
rect 5336 2998 5379 3012
rect 5403 3009 5410 3016
rect 5413 3012 5480 3036
rect 5512 3036 5684 3038
rect 5482 3014 5510 3018
rect 5512 3014 5592 3036
rect 5613 3034 5628 3036
rect 5482 3012 5592 3014
rect 5413 3008 5592 3012
rect 5386 2998 5416 3008
rect 5418 2998 5571 3008
rect 5579 2998 5609 3008
rect 5613 2998 5643 3012
rect 5671 2998 5684 3036
rect 5756 3042 5791 3050
rect 5756 3016 5757 3042
rect 5764 3016 5791 3042
rect 5699 2998 5729 3012
rect 5756 3008 5791 3016
rect 5793 3042 5834 3050
rect 5793 3016 5808 3042
rect 5815 3016 5834 3042
rect 5898 3038 5960 3050
rect 5972 3038 6047 3050
rect 6105 3038 6180 3050
rect 6192 3038 6223 3050
rect 6229 3038 6264 3050
rect 5898 3036 6060 3038
rect 5793 3008 5834 3016
rect 5916 3012 5929 3036
rect 5944 3034 5959 3036
rect 5756 2998 5757 3008
rect 5772 2998 5785 3008
rect 5799 2998 5800 3008
rect 5815 2998 5828 3008
rect 5843 2998 5873 3012
rect 5916 2998 5959 3012
rect 5983 3009 5990 3016
rect 5993 3012 6060 3036
rect 6092 3036 6264 3038
rect 6062 3014 6090 3018
rect 6092 3014 6172 3036
rect 6193 3034 6208 3036
rect 6062 3012 6172 3014
rect 5993 3008 6172 3012
rect 5966 2998 5996 3008
rect 5998 2998 6151 3008
rect 6159 2998 6189 3008
rect 6193 2998 6223 3012
rect 6251 2998 6264 3036
rect 6336 3042 6371 3050
rect 6336 3016 6337 3042
rect 6344 3016 6371 3042
rect 6279 2998 6309 3012
rect 6336 3008 6371 3016
rect 6373 3042 6414 3050
rect 6373 3016 6388 3042
rect 6395 3016 6414 3042
rect 6478 3038 6540 3050
rect 6552 3038 6627 3050
rect 6685 3038 6760 3050
rect 6772 3038 6803 3050
rect 6809 3038 6844 3050
rect 6478 3036 6640 3038
rect 6373 3008 6414 3016
rect 6496 3012 6509 3036
rect 6524 3034 6539 3036
rect 6336 2998 6337 3008
rect 6352 2998 6365 3008
rect 6379 2998 6380 3008
rect 6395 2998 6408 3008
rect 6423 2998 6453 3012
rect 6496 2998 6539 3012
rect 6563 3009 6570 3016
rect 6573 3012 6640 3036
rect 6672 3036 6844 3038
rect 6642 3014 6670 3018
rect 6672 3014 6752 3036
rect 6773 3034 6788 3036
rect 6642 3012 6752 3014
rect 6573 3008 6752 3012
rect 6546 2998 6576 3008
rect 6578 2998 6731 3008
rect 6739 2998 6769 3008
rect 6773 2998 6803 3012
rect 6831 2998 6844 3036
rect 6916 3042 6951 3050
rect 6916 3016 6917 3042
rect 6924 3016 6951 3042
rect 6859 2998 6889 3012
rect 6916 3008 6951 3016
rect 6953 3042 6994 3050
rect 6953 3016 6968 3042
rect 6975 3016 6994 3042
rect 7058 3038 7120 3050
rect 7132 3038 7207 3050
rect 7265 3038 7340 3050
rect 7352 3038 7383 3050
rect 7389 3038 7424 3050
rect 7058 3036 7220 3038
rect 6953 3008 6994 3016
rect 7076 3012 7089 3036
rect 7104 3034 7119 3036
rect 6916 2998 6917 3008
rect 6932 2998 6945 3008
rect 6959 2998 6960 3008
rect 6975 2998 6988 3008
rect 7003 2998 7033 3012
rect 7076 2998 7119 3012
rect 7143 3009 7150 3016
rect 7153 3012 7220 3036
rect 7252 3036 7424 3038
rect 7222 3014 7250 3018
rect 7252 3014 7332 3036
rect 7353 3034 7368 3036
rect 7222 3012 7332 3014
rect 7153 3008 7332 3012
rect 7126 2998 7156 3008
rect 7158 2998 7311 3008
rect 7319 2998 7349 3008
rect 7353 2998 7383 3012
rect 7411 2998 7424 3036
rect 7496 3042 7531 3050
rect 7496 3016 7497 3042
rect 7504 3016 7531 3042
rect 7439 2998 7469 3012
rect 7496 3008 7531 3016
rect 7533 3042 7574 3050
rect 7533 3016 7548 3042
rect 7555 3016 7574 3042
rect 7638 3038 7700 3050
rect 7712 3038 7787 3050
rect 7845 3038 7920 3050
rect 7932 3038 7963 3050
rect 7969 3038 8004 3050
rect 7638 3036 7800 3038
rect 7533 3008 7574 3016
rect 7656 3012 7669 3036
rect 7684 3034 7699 3036
rect 7496 2998 7497 3008
rect 7512 2998 7525 3008
rect 7539 2998 7540 3008
rect 7555 2998 7568 3008
rect 7583 2998 7613 3012
rect 7656 2998 7699 3012
rect 7723 3009 7730 3016
rect 7733 3012 7800 3036
rect 7832 3036 8004 3038
rect 7802 3014 7830 3018
rect 7832 3014 7912 3036
rect 7933 3034 7948 3036
rect 7802 3012 7912 3014
rect 7733 3008 7912 3012
rect 7706 2998 7736 3008
rect 7738 2998 7891 3008
rect 7899 2998 7929 3008
rect 7933 2998 7963 3012
rect 7991 2998 8004 3036
rect 8076 3042 8111 3050
rect 8076 3016 8077 3042
rect 8084 3016 8111 3042
rect 8019 2998 8049 3012
rect 8076 3008 8111 3016
rect 8113 3042 8154 3050
rect 8113 3016 8128 3042
rect 8135 3016 8154 3042
rect 8218 3038 8280 3050
rect 8292 3038 8367 3050
rect 8425 3038 8500 3050
rect 8512 3038 8543 3050
rect 8549 3038 8584 3050
rect 8218 3036 8380 3038
rect 8113 3008 8154 3016
rect 8236 3012 8249 3036
rect 8264 3034 8279 3036
rect 8076 2998 8077 3008
rect 8092 2998 8105 3008
rect 8119 2998 8120 3008
rect 8135 2998 8148 3008
rect 8163 2998 8193 3012
rect 8236 2998 8279 3012
rect 8303 3009 8310 3016
rect 8313 3012 8380 3036
rect 8412 3036 8584 3038
rect 8382 3014 8410 3018
rect 8412 3014 8492 3036
rect 8513 3034 8528 3036
rect 8382 3012 8492 3014
rect 8313 3008 8492 3012
rect 8286 2998 8316 3008
rect 8318 2998 8471 3008
rect 8479 2998 8509 3008
rect 8513 2998 8543 3012
rect 8571 2998 8584 3036
rect 8656 3042 8691 3050
rect 8656 3016 8657 3042
rect 8664 3016 8691 3042
rect 8599 2998 8629 3012
rect 8656 3008 8691 3016
rect 8693 3042 8734 3050
rect 8693 3016 8708 3042
rect 8715 3016 8734 3042
rect 8798 3038 8860 3050
rect 8872 3038 8947 3050
rect 9005 3038 9080 3050
rect 9092 3038 9123 3050
rect 9129 3038 9164 3050
rect 8798 3036 8960 3038
rect 8693 3008 8734 3016
rect 8816 3012 8829 3036
rect 8844 3034 8859 3036
rect 8656 2998 8657 3008
rect 8672 2998 8685 3008
rect 8699 2998 8700 3008
rect 8715 2998 8728 3008
rect 8743 2998 8773 3012
rect 8816 2998 8859 3012
rect 8883 3009 8890 3016
rect 8893 3012 8960 3036
rect 8992 3036 9164 3038
rect 8962 3014 8990 3018
rect 8992 3014 9072 3036
rect 9093 3034 9108 3036
rect 8962 3012 9072 3014
rect 8893 3008 9072 3012
rect 8866 2998 8896 3008
rect 8898 2998 9051 3008
rect 9059 2998 9089 3008
rect 9093 2998 9123 3012
rect 9151 2998 9164 3036
rect 9236 3042 9271 3050
rect 9236 3016 9237 3042
rect 9244 3016 9271 3042
rect 9179 2998 9209 3012
rect 9236 3008 9271 3016
rect 9236 2998 9237 3008
rect 9252 2998 9265 3008
rect -1 2992 9265 2998
rect 0 2984 9265 2992
rect 15 2954 28 2984
rect 43 2966 73 2984
rect 116 2970 130 2984
rect 166 2970 386 2984
rect 117 2968 130 2970
rect 83 2956 98 2968
rect 80 2954 102 2956
rect 107 2954 137 2968
rect 198 2966 351 2970
rect 180 2954 372 2966
rect 415 2954 445 2968
rect 451 2954 464 2984
rect 479 2966 509 2984
rect 552 2954 565 2984
rect 595 2954 608 2984
rect 623 2966 653 2984
rect 696 2970 710 2984
rect 746 2970 966 2984
rect 697 2968 710 2970
rect 663 2956 678 2968
rect 660 2954 682 2956
rect 687 2954 717 2968
rect 778 2966 931 2970
rect 760 2954 952 2966
rect 995 2954 1025 2968
rect 1031 2954 1044 2984
rect 1059 2966 1089 2984
rect 1132 2954 1145 2984
rect 1175 2954 1188 2984
rect 1203 2966 1233 2984
rect 1276 2970 1290 2984
rect 1326 2970 1546 2984
rect 1277 2968 1290 2970
rect 1243 2956 1258 2968
rect 1240 2954 1262 2956
rect 1267 2954 1297 2968
rect 1358 2966 1511 2970
rect 1340 2954 1532 2966
rect 1575 2954 1605 2968
rect 1611 2954 1624 2984
rect 1639 2966 1669 2984
rect 1712 2954 1725 2984
rect 1755 2954 1768 2984
rect 1783 2966 1813 2984
rect 1856 2970 1870 2984
rect 1906 2970 2126 2984
rect 1857 2968 1870 2970
rect 1823 2956 1838 2968
rect 1820 2954 1842 2956
rect 1847 2954 1877 2968
rect 1938 2966 2091 2970
rect 1920 2954 2112 2966
rect 2155 2954 2185 2968
rect 2191 2954 2204 2984
rect 2219 2966 2249 2984
rect 2292 2954 2305 2984
rect 2335 2954 2348 2984
rect 2363 2966 2393 2984
rect 2436 2970 2450 2984
rect 2486 2970 2706 2984
rect 2437 2968 2450 2970
rect 2403 2956 2418 2968
rect 2400 2954 2422 2956
rect 2427 2954 2457 2968
rect 2518 2966 2671 2970
rect 2500 2954 2692 2966
rect 2735 2954 2765 2968
rect 2771 2954 2784 2984
rect 2799 2966 2829 2984
rect 2872 2954 2885 2984
rect 2915 2954 2928 2984
rect 2943 2966 2973 2984
rect 3016 2970 3030 2984
rect 3066 2970 3286 2984
rect 3017 2968 3030 2970
rect 2983 2956 2998 2968
rect 2980 2954 3002 2956
rect 3007 2954 3037 2968
rect 3098 2966 3251 2970
rect 3080 2954 3272 2966
rect 3315 2954 3345 2968
rect 3351 2954 3364 2984
rect 3379 2966 3409 2984
rect 3452 2954 3465 2984
rect 3495 2954 3508 2984
rect 3523 2966 3553 2984
rect 3596 2970 3610 2984
rect 3646 2970 3866 2984
rect 3597 2968 3610 2970
rect 3563 2956 3578 2968
rect 3560 2954 3582 2956
rect 3587 2954 3617 2968
rect 3678 2966 3831 2970
rect 3660 2954 3852 2966
rect 3895 2954 3925 2968
rect 3931 2954 3944 2984
rect 3959 2966 3989 2984
rect 4032 2954 4045 2984
rect 4075 2954 4088 2984
rect 4103 2966 4133 2984
rect 4176 2970 4190 2984
rect 4226 2970 4446 2984
rect 4177 2968 4190 2970
rect 4143 2956 4158 2968
rect 4140 2954 4162 2956
rect 4167 2954 4197 2968
rect 4258 2966 4411 2970
rect 4240 2954 4432 2966
rect 4475 2954 4505 2968
rect 4511 2954 4524 2984
rect 4539 2966 4569 2984
rect 4612 2954 4625 2984
rect 4655 2954 4668 2984
rect 4683 2966 4713 2984
rect 4756 2970 4770 2984
rect 4806 2970 5026 2984
rect 4757 2968 4770 2970
rect 4723 2956 4738 2968
rect 4720 2954 4742 2956
rect 4747 2954 4777 2968
rect 4838 2966 4991 2970
rect 4820 2954 5012 2966
rect 5055 2954 5085 2968
rect 5091 2954 5104 2984
rect 5119 2966 5149 2984
rect 5192 2954 5205 2984
rect 5235 2954 5248 2984
rect 5263 2966 5293 2984
rect 5336 2970 5350 2984
rect 5386 2970 5606 2984
rect 5337 2968 5350 2970
rect 5303 2956 5318 2968
rect 5300 2954 5322 2956
rect 5327 2954 5357 2968
rect 5418 2966 5571 2970
rect 5400 2954 5592 2966
rect 5635 2954 5665 2968
rect 5671 2954 5684 2984
rect 5699 2966 5729 2984
rect 5772 2954 5785 2984
rect 5815 2954 5828 2984
rect 5843 2966 5873 2984
rect 5916 2970 5930 2984
rect 5966 2970 6186 2984
rect 5917 2968 5930 2970
rect 5883 2956 5898 2968
rect 5880 2954 5902 2956
rect 5907 2954 5937 2968
rect 5998 2966 6151 2970
rect 5980 2954 6172 2966
rect 6215 2954 6245 2968
rect 6251 2954 6264 2984
rect 6279 2966 6309 2984
rect 6352 2954 6365 2984
rect 6395 2954 6408 2984
rect 6423 2966 6453 2984
rect 6496 2970 6510 2984
rect 6546 2970 6766 2984
rect 6497 2968 6510 2970
rect 6463 2956 6478 2968
rect 6460 2954 6482 2956
rect 6487 2954 6517 2968
rect 6578 2966 6731 2970
rect 6560 2954 6752 2966
rect 6795 2954 6825 2968
rect 6831 2954 6844 2984
rect 6859 2966 6889 2984
rect 6932 2954 6945 2984
rect 6975 2954 6988 2984
rect 7003 2966 7033 2984
rect 7076 2970 7090 2984
rect 7126 2970 7346 2984
rect 7077 2968 7090 2970
rect 7043 2956 7058 2968
rect 7040 2954 7062 2956
rect 7067 2954 7097 2968
rect 7158 2966 7311 2970
rect 7140 2954 7332 2966
rect 7375 2954 7405 2968
rect 7411 2954 7424 2984
rect 7439 2966 7469 2984
rect 7512 2954 7525 2984
rect 7555 2954 7568 2984
rect 7583 2966 7613 2984
rect 7656 2970 7670 2984
rect 7706 2970 7926 2984
rect 7657 2968 7670 2970
rect 7623 2956 7638 2968
rect 7620 2954 7642 2956
rect 7647 2954 7677 2968
rect 7738 2966 7891 2970
rect 7720 2954 7912 2966
rect 7955 2954 7985 2968
rect 7991 2954 8004 2984
rect 8019 2966 8049 2984
rect 8092 2954 8105 2984
rect 8135 2954 8148 2984
rect 8163 2966 8193 2984
rect 8236 2970 8250 2984
rect 8286 2970 8506 2984
rect 8237 2968 8250 2970
rect 8203 2956 8218 2968
rect 8200 2954 8222 2956
rect 8227 2954 8257 2968
rect 8318 2966 8471 2970
rect 8300 2954 8492 2966
rect 8535 2954 8565 2968
rect 8571 2954 8584 2984
rect 8599 2966 8629 2984
rect 8672 2954 8685 2984
rect 8715 2954 8728 2984
rect 8743 2966 8773 2984
rect 8816 2970 8830 2984
rect 8866 2970 9086 2984
rect 8817 2968 8830 2970
rect 8783 2956 8798 2968
rect 8780 2954 8802 2956
rect 8807 2954 8837 2968
rect 8898 2966 9051 2970
rect 8880 2954 9072 2966
rect 9115 2954 9145 2968
rect 9151 2954 9164 2984
rect 9179 2966 9209 2984
rect 9252 2954 9265 2984
rect 0 2940 9265 2954
rect 15 2836 28 2940
rect 73 2918 74 2928
rect 89 2918 102 2928
rect 73 2914 102 2918
rect 107 2914 137 2940
rect 155 2926 171 2928
rect 243 2926 296 2940
rect 244 2924 308 2926
rect 351 2924 366 2940
rect 415 2937 445 2940
rect 415 2934 451 2937
rect 381 2926 397 2928
rect 155 2914 170 2918
rect 73 2912 170 2914
rect 198 2912 366 2924
rect 382 2914 397 2918
rect 415 2915 454 2934
rect 473 2928 480 2929
rect 479 2921 480 2928
rect 463 2918 464 2921
rect 479 2918 492 2921
rect 415 2914 445 2915
rect 454 2914 460 2915
rect 463 2914 492 2918
rect 382 2913 492 2914
rect 382 2912 498 2913
rect 57 2904 108 2912
rect 57 2892 82 2904
rect 89 2892 108 2904
rect 139 2904 189 2912
rect 139 2896 155 2904
rect 162 2902 189 2904
rect 198 2902 419 2912
rect 162 2892 419 2902
rect 448 2904 498 2912
rect 448 2895 464 2904
rect 57 2884 108 2892
rect 155 2884 419 2892
rect 445 2892 464 2895
rect 471 2892 498 2904
rect 445 2884 498 2892
rect 73 2876 74 2884
rect 89 2876 102 2884
rect 73 2868 89 2876
rect 70 2861 89 2864
rect 70 2852 92 2861
rect 43 2842 92 2852
rect 43 2836 73 2842
rect 92 2837 97 2842
rect 15 2820 89 2836
rect 107 2828 137 2884
rect 172 2874 380 2884
rect 415 2880 460 2884
rect 463 2883 464 2884
rect 479 2883 492 2884
rect 198 2844 387 2874
rect 213 2841 387 2844
rect 206 2838 387 2841
rect 15 2818 28 2820
rect 43 2818 77 2820
rect 15 2802 89 2818
rect 116 2814 129 2828
rect 144 2814 160 2830
rect 206 2825 217 2838
rect -1 2780 0 2796
rect 15 2780 28 2802
rect 43 2780 73 2802
rect 116 2798 178 2814
rect 206 2807 217 2823
rect 222 2818 232 2838
rect 242 2818 256 2838
rect 259 2825 268 2838
rect 284 2825 293 2838
rect 222 2807 256 2818
rect 259 2807 268 2823
rect 284 2807 293 2823
rect 300 2818 310 2838
rect 320 2818 334 2838
rect 335 2825 346 2838
rect 300 2807 334 2818
rect 335 2807 346 2823
rect 392 2814 408 2830
rect 415 2828 445 2880
rect 479 2876 480 2883
rect 464 2868 480 2876
rect 451 2836 464 2855
rect 479 2836 509 2852
rect 451 2820 525 2836
rect 451 2818 464 2820
rect 479 2818 513 2820
rect 116 2796 129 2798
rect 144 2796 178 2798
rect 116 2780 178 2796
rect 222 2791 238 2794
rect 300 2791 330 2802
rect 378 2798 424 2814
rect 451 2802 525 2818
rect 378 2796 412 2798
rect 377 2780 424 2796
rect 451 2780 464 2802
rect 479 2780 509 2802
rect 536 2780 537 2796
rect 552 2780 565 2940
rect 595 2836 608 2940
rect 653 2918 654 2928
rect 669 2918 682 2928
rect 653 2914 682 2918
rect 687 2914 717 2940
rect 735 2926 751 2928
rect 823 2926 876 2940
rect 824 2924 888 2926
rect 931 2924 946 2940
rect 995 2937 1025 2940
rect 995 2934 1031 2937
rect 961 2926 977 2928
rect 735 2914 750 2918
rect 653 2912 750 2914
rect 778 2912 946 2924
rect 962 2914 977 2918
rect 995 2915 1034 2934
rect 1053 2928 1060 2929
rect 1059 2921 1060 2928
rect 1043 2918 1044 2921
rect 1059 2918 1072 2921
rect 995 2914 1025 2915
rect 1034 2914 1040 2915
rect 1043 2914 1072 2918
rect 962 2913 1072 2914
rect 962 2912 1078 2913
rect 637 2904 688 2912
rect 637 2892 662 2904
rect 669 2892 688 2904
rect 719 2904 769 2912
rect 719 2896 735 2904
rect 742 2902 769 2904
rect 778 2902 999 2912
rect 742 2892 999 2902
rect 1028 2904 1078 2912
rect 1028 2895 1044 2904
rect 637 2884 688 2892
rect 735 2884 999 2892
rect 1025 2892 1044 2895
rect 1051 2892 1078 2904
rect 1025 2884 1078 2892
rect 653 2876 654 2884
rect 669 2876 682 2884
rect 653 2868 669 2876
rect 650 2861 669 2864
rect 650 2852 672 2861
rect 623 2842 672 2852
rect 623 2836 653 2842
rect 672 2837 677 2842
rect 595 2820 669 2836
rect 687 2828 717 2884
rect 752 2874 960 2884
rect 995 2880 1040 2884
rect 1043 2883 1044 2884
rect 1059 2883 1072 2884
rect 778 2844 967 2874
rect 793 2841 967 2844
rect 786 2838 967 2841
rect 595 2818 608 2820
rect 623 2818 657 2820
rect 595 2802 669 2818
rect 696 2814 709 2828
rect 724 2814 740 2830
rect 786 2825 797 2838
rect 579 2780 580 2796
rect 595 2780 608 2802
rect 623 2780 653 2802
rect 696 2798 758 2814
rect 786 2807 797 2823
rect 802 2818 812 2838
rect 822 2818 836 2838
rect 839 2825 848 2838
rect 864 2825 873 2838
rect 802 2807 836 2818
rect 839 2807 848 2823
rect 864 2807 873 2823
rect 880 2818 890 2838
rect 900 2818 914 2838
rect 915 2825 926 2838
rect 880 2807 914 2818
rect 915 2807 926 2823
rect 972 2814 988 2830
rect 995 2828 1025 2880
rect 1059 2876 1060 2883
rect 1044 2868 1060 2876
rect 1031 2836 1044 2855
rect 1059 2836 1089 2852
rect 1031 2820 1105 2836
rect 1031 2818 1044 2820
rect 1059 2818 1093 2820
rect 696 2796 709 2798
rect 724 2796 758 2798
rect 696 2780 758 2796
rect 802 2791 818 2794
rect 880 2791 910 2802
rect 958 2798 1004 2814
rect 1031 2802 1105 2818
rect 958 2796 992 2798
rect 957 2780 1004 2796
rect 1031 2780 1044 2802
rect 1059 2780 1089 2802
rect 1116 2780 1117 2796
rect 1132 2780 1145 2940
rect 1175 2836 1188 2940
rect 1233 2918 1234 2928
rect 1249 2918 1262 2928
rect 1233 2914 1262 2918
rect 1267 2914 1297 2940
rect 1315 2926 1331 2928
rect 1403 2926 1456 2940
rect 1404 2924 1468 2926
rect 1511 2924 1526 2940
rect 1575 2937 1605 2940
rect 1575 2934 1611 2937
rect 1541 2926 1557 2928
rect 1315 2914 1330 2918
rect 1233 2912 1330 2914
rect 1358 2912 1526 2924
rect 1542 2914 1557 2918
rect 1575 2915 1614 2934
rect 1633 2928 1640 2929
rect 1639 2921 1640 2928
rect 1623 2918 1624 2921
rect 1639 2918 1652 2921
rect 1575 2914 1605 2915
rect 1614 2914 1620 2915
rect 1623 2914 1652 2918
rect 1542 2913 1652 2914
rect 1542 2912 1658 2913
rect 1217 2904 1268 2912
rect 1217 2892 1242 2904
rect 1249 2892 1268 2904
rect 1299 2904 1349 2912
rect 1299 2896 1315 2904
rect 1322 2902 1349 2904
rect 1358 2902 1579 2912
rect 1322 2892 1579 2902
rect 1608 2904 1658 2912
rect 1608 2895 1624 2904
rect 1217 2884 1268 2892
rect 1315 2884 1579 2892
rect 1605 2892 1624 2895
rect 1631 2892 1658 2904
rect 1605 2884 1658 2892
rect 1233 2876 1234 2884
rect 1249 2876 1262 2884
rect 1233 2868 1249 2876
rect 1230 2861 1249 2864
rect 1230 2852 1252 2861
rect 1203 2842 1252 2852
rect 1203 2836 1233 2842
rect 1252 2837 1257 2842
rect 1175 2820 1249 2836
rect 1267 2828 1297 2884
rect 1332 2874 1540 2884
rect 1575 2880 1620 2884
rect 1623 2883 1624 2884
rect 1639 2883 1652 2884
rect 1358 2844 1547 2874
rect 1373 2841 1547 2844
rect 1366 2838 1547 2841
rect 1175 2818 1188 2820
rect 1203 2818 1237 2820
rect 1175 2802 1249 2818
rect 1276 2814 1289 2828
rect 1304 2814 1320 2830
rect 1366 2825 1377 2838
rect 1159 2780 1160 2796
rect 1175 2780 1188 2802
rect 1203 2780 1233 2802
rect 1276 2798 1338 2814
rect 1366 2807 1377 2823
rect 1382 2818 1392 2838
rect 1402 2818 1416 2838
rect 1419 2825 1428 2838
rect 1444 2825 1453 2838
rect 1382 2807 1416 2818
rect 1419 2807 1428 2823
rect 1444 2807 1453 2823
rect 1460 2818 1470 2838
rect 1480 2818 1494 2838
rect 1495 2825 1506 2838
rect 1460 2807 1494 2818
rect 1495 2807 1506 2823
rect 1552 2814 1568 2830
rect 1575 2828 1605 2880
rect 1639 2876 1640 2883
rect 1624 2868 1640 2876
rect 1611 2836 1624 2855
rect 1639 2836 1669 2852
rect 1611 2820 1685 2836
rect 1611 2818 1624 2820
rect 1639 2818 1673 2820
rect 1276 2796 1289 2798
rect 1304 2796 1338 2798
rect 1276 2780 1338 2796
rect 1382 2791 1398 2794
rect 1460 2791 1490 2802
rect 1538 2798 1584 2814
rect 1611 2802 1685 2818
rect 1538 2796 1572 2798
rect 1537 2780 1584 2796
rect 1611 2780 1624 2802
rect 1639 2780 1669 2802
rect 1696 2780 1697 2796
rect 1712 2780 1725 2940
rect 1755 2836 1768 2940
rect 1813 2918 1814 2928
rect 1829 2918 1842 2928
rect 1813 2914 1842 2918
rect 1847 2914 1877 2940
rect 1895 2926 1911 2928
rect 1983 2926 2036 2940
rect 1984 2924 2048 2926
rect 2091 2924 2106 2940
rect 2155 2937 2185 2940
rect 2155 2934 2191 2937
rect 2121 2926 2137 2928
rect 1895 2914 1910 2918
rect 1813 2912 1910 2914
rect 1938 2912 2106 2924
rect 2122 2914 2137 2918
rect 2155 2915 2194 2934
rect 2213 2928 2220 2929
rect 2219 2921 2220 2928
rect 2203 2918 2204 2921
rect 2219 2918 2232 2921
rect 2155 2914 2185 2915
rect 2194 2914 2200 2915
rect 2203 2914 2232 2918
rect 2122 2913 2232 2914
rect 2122 2912 2238 2913
rect 1797 2904 1848 2912
rect 1797 2892 1822 2904
rect 1829 2892 1848 2904
rect 1879 2904 1929 2912
rect 1879 2896 1895 2904
rect 1902 2902 1929 2904
rect 1938 2902 2159 2912
rect 1902 2892 2159 2902
rect 2188 2904 2238 2912
rect 2188 2895 2204 2904
rect 1797 2884 1848 2892
rect 1895 2884 2159 2892
rect 2185 2892 2204 2895
rect 2211 2892 2238 2904
rect 2185 2884 2238 2892
rect 1813 2876 1814 2884
rect 1829 2876 1842 2884
rect 1813 2868 1829 2876
rect 1810 2861 1829 2864
rect 1810 2852 1832 2861
rect 1783 2842 1832 2852
rect 1783 2836 1813 2842
rect 1832 2837 1837 2842
rect 1755 2820 1829 2836
rect 1847 2828 1877 2884
rect 1912 2874 2120 2884
rect 2155 2880 2200 2884
rect 2203 2883 2204 2884
rect 2219 2883 2232 2884
rect 1938 2844 2127 2874
rect 1953 2841 2127 2844
rect 1946 2838 2127 2841
rect 1755 2818 1768 2820
rect 1783 2818 1817 2820
rect 1755 2802 1829 2818
rect 1856 2814 1869 2828
rect 1884 2814 1900 2830
rect 1946 2825 1957 2838
rect 1739 2780 1740 2796
rect 1755 2780 1768 2802
rect 1783 2780 1813 2802
rect 1856 2798 1918 2814
rect 1946 2807 1957 2823
rect 1962 2818 1972 2838
rect 1982 2818 1996 2838
rect 1999 2825 2008 2838
rect 2024 2825 2033 2838
rect 1962 2807 1996 2818
rect 1999 2807 2008 2823
rect 2024 2807 2033 2823
rect 2040 2818 2050 2838
rect 2060 2818 2074 2838
rect 2075 2825 2086 2838
rect 2040 2807 2074 2818
rect 2075 2807 2086 2823
rect 2132 2814 2148 2830
rect 2155 2828 2185 2880
rect 2219 2876 2220 2883
rect 2204 2868 2220 2876
rect 2191 2836 2204 2855
rect 2219 2836 2249 2852
rect 2191 2820 2265 2836
rect 2191 2818 2204 2820
rect 2219 2818 2253 2820
rect 1856 2796 1869 2798
rect 1884 2796 1918 2798
rect 1856 2780 1918 2796
rect 1962 2791 1976 2794
rect 2040 2791 2070 2802
rect 2118 2798 2164 2814
rect 2191 2802 2265 2818
rect 2118 2796 2152 2798
rect 2117 2780 2164 2796
rect 2191 2780 2204 2802
rect 2219 2780 2249 2802
rect 2276 2780 2277 2796
rect 2292 2780 2305 2940
rect 2335 2836 2348 2940
rect 2393 2918 2394 2928
rect 2409 2918 2422 2928
rect 2393 2914 2422 2918
rect 2427 2914 2457 2940
rect 2475 2926 2491 2928
rect 2563 2926 2616 2940
rect 2564 2924 2628 2926
rect 2671 2924 2686 2940
rect 2735 2937 2765 2940
rect 2735 2934 2771 2937
rect 2701 2926 2717 2928
rect 2475 2914 2490 2918
rect 2393 2912 2490 2914
rect 2518 2912 2686 2924
rect 2702 2914 2717 2918
rect 2735 2915 2774 2934
rect 2793 2928 2800 2929
rect 2799 2921 2800 2928
rect 2783 2918 2784 2921
rect 2799 2918 2812 2921
rect 2735 2914 2765 2915
rect 2774 2914 2780 2915
rect 2783 2914 2812 2918
rect 2702 2913 2812 2914
rect 2702 2912 2818 2913
rect 2377 2904 2428 2912
rect 2377 2892 2402 2904
rect 2409 2892 2428 2904
rect 2459 2904 2509 2912
rect 2459 2896 2475 2904
rect 2482 2902 2509 2904
rect 2518 2902 2739 2912
rect 2482 2892 2739 2902
rect 2768 2904 2818 2912
rect 2768 2895 2784 2904
rect 2377 2884 2428 2892
rect 2475 2884 2739 2892
rect 2765 2892 2784 2895
rect 2791 2892 2818 2904
rect 2765 2884 2818 2892
rect 2393 2876 2394 2884
rect 2409 2876 2422 2884
rect 2393 2868 2409 2876
rect 2390 2861 2409 2864
rect 2390 2852 2412 2861
rect 2363 2842 2412 2852
rect 2363 2836 2393 2842
rect 2412 2837 2417 2842
rect 2335 2820 2409 2836
rect 2427 2828 2457 2884
rect 2492 2874 2700 2884
rect 2735 2880 2780 2884
rect 2783 2883 2784 2884
rect 2799 2883 2812 2884
rect 2518 2844 2707 2874
rect 2533 2841 2707 2844
rect 2526 2838 2707 2841
rect 2335 2818 2348 2820
rect 2363 2818 2397 2820
rect 2335 2802 2409 2818
rect 2436 2814 2449 2828
rect 2464 2814 2480 2830
rect 2526 2825 2537 2838
rect 2319 2780 2320 2796
rect 2335 2780 2348 2802
rect 2363 2780 2393 2802
rect 2436 2798 2498 2814
rect 2526 2807 2537 2823
rect 2542 2818 2552 2838
rect 2562 2818 2576 2838
rect 2579 2825 2588 2838
rect 2604 2825 2613 2838
rect 2542 2807 2576 2818
rect 2579 2807 2588 2823
rect 2604 2807 2613 2823
rect 2620 2818 2630 2838
rect 2640 2818 2654 2838
rect 2655 2825 2666 2838
rect 2620 2807 2654 2818
rect 2655 2807 2666 2823
rect 2712 2814 2728 2830
rect 2735 2828 2765 2880
rect 2799 2876 2800 2883
rect 2784 2868 2800 2876
rect 2771 2836 2784 2855
rect 2799 2836 2829 2852
rect 2771 2820 2845 2836
rect 2771 2818 2784 2820
rect 2799 2818 2833 2820
rect 2436 2796 2449 2798
rect 2464 2796 2498 2798
rect 2436 2780 2498 2796
rect 2542 2791 2558 2794
rect 2620 2791 2650 2802
rect 2698 2798 2744 2814
rect 2771 2802 2845 2818
rect 2698 2796 2732 2798
rect 2697 2780 2744 2796
rect 2771 2780 2784 2802
rect 2799 2780 2829 2802
rect 2856 2780 2857 2796
rect 2872 2780 2885 2940
rect 2915 2836 2928 2940
rect 2973 2918 2974 2928
rect 2989 2918 3002 2928
rect 2973 2914 3002 2918
rect 3007 2914 3037 2940
rect 3055 2926 3071 2928
rect 3143 2926 3196 2940
rect 3144 2924 3208 2926
rect 3251 2924 3266 2940
rect 3315 2937 3345 2940
rect 3315 2934 3351 2937
rect 3281 2926 3297 2928
rect 3055 2914 3070 2918
rect 2973 2912 3070 2914
rect 3098 2912 3266 2924
rect 3282 2914 3297 2918
rect 3315 2915 3354 2934
rect 3373 2928 3380 2929
rect 3379 2921 3380 2928
rect 3363 2918 3364 2921
rect 3379 2918 3392 2921
rect 3315 2914 3345 2915
rect 3354 2914 3360 2915
rect 3363 2914 3392 2918
rect 3282 2913 3392 2914
rect 3282 2912 3398 2913
rect 2957 2904 3008 2912
rect 2957 2892 2982 2904
rect 2989 2892 3008 2904
rect 3039 2904 3089 2912
rect 3039 2896 3055 2904
rect 3062 2902 3089 2904
rect 3098 2902 3319 2912
rect 3062 2892 3319 2902
rect 3348 2904 3398 2912
rect 3348 2895 3364 2904
rect 2957 2884 3008 2892
rect 3055 2884 3319 2892
rect 3345 2892 3364 2895
rect 3371 2892 3398 2904
rect 3345 2884 3398 2892
rect 2973 2876 2974 2884
rect 2989 2876 3002 2884
rect 2973 2868 2989 2876
rect 2970 2861 2989 2864
rect 2970 2852 2992 2861
rect 2943 2842 2992 2852
rect 2943 2836 2973 2842
rect 2992 2837 2997 2842
rect 2915 2820 2989 2836
rect 3007 2828 3037 2884
rect 3072 2874 3280 2884
rect 3315 2880 3360 2884
rect 3363 2883 3364 2884
rect 3379 2883 3392 2884
rect 3098 2844 3287 2874
rect 3113 2841 3287 2844
rect 3106 2838 3287 2841
rect 2915 2818 2928 2820
rect 2943 2818 2977 2820
rect 2915 2802 2989 2818
rect 3016 2814 3029 2828
rect 3044 2814 3060 2830
rect 3106 2825 3117 2838
rect 2899 2780 2900 2796
rect 2915 2780 2928 2802
rect 2943 2780 2973 2802
rect 3016 2798 3078 2814
rect 3106 2807 3117 2823
rect 3122 2818 3132 2838
rect 3142 2818 3156 2838
rect 3159 2825 3168 2838
rect 3184 2825 3193 2838
rect 3122 2807 3156 2818
rect 3159 2807 3168 2823
rect 3184 2807 3193 2823
rect 3200 2818 3210 2838
rect 3220 2818 3234 2838
rect 3235 2825 3246 2838
rect 3200 2807 3234 2818
rect 3235 2807 3246 2823
rect 3292 2814 3308 2830
rect 3315 2828 3345 2880
rect 3379 2876 3380 2883
rect 3364 2868 3380 2876
rect 3351 2836 3364 2855
rect 3379 2836 3409 2852
rect 3351 2820 3425 2836
rect 3351 2818 3364 2820
rect 3379 2818 3413 2820
rect 3016 2796 3029 2798
rect 3044 2796 3078 2798
rect 3016 2780 3078 2796
rect 3122 2791 3138 2794
rect 3200 2791 3230 2802
rect 3278 2798 3324 2814
rect 3351 2802 3425 2818
rect 3278 2796 3312 2798
rect 3277 2780 3324 2796
rect 3351 2780 3364 2802
rect 3379 2780 3409 2802
rect 3436 2780 3437 2796
rect 3452 2780 3465 2940
rect 3495 2836 3508 2940
rect 3553 2918 3554 2928
rect 3569 2918 3582 2928
rect 3553 2914 3582 2918
rect 3587 2914 3617 2940
rect 3635 2926 3651 2928
rect 3723 2926 3776 2940
rect 3724 2924 3788 2926
rect 3831 2924 3846 2940
rect 3895 2937 3925 2940
rect 3895 2934 3931 2937
rect 3861 2926 3877 2928
rect 3635 2914 3650 2918
rect 3553 2912 3650 2914
rect 3678 2912 3846 2924
rect 3862 2914 3877 2918
rect 3895 2915 3934 2934
rect 3953 2928 3960 2929
rect 3959 2921 3960 2928
rect 3943 2918 3944 2921
rect 3959 2918 3972 2921
rect 3895 2914 3925 2915
rect 3934 2914 3940 2915
rect 3943 2914 3972 2918
rect 3862 2913 3972 2914
rect 3862 2912 3978 2913
rect 3537 2904 3588 2912
rect 3537 2892 3562 2904
rect 3569 2892 3588 2904
rect 3619 2904 3669 2912
rect 3619 2896 3635 2904
rect 3642 2902 3669 2904
rect 3678 2902 3899 2912
rect 3642 2892 3899 2902
rect 3928 2904 3978 2912
rect 3928 2895 3944 2904
rect 3537 2884 3588 2892
rect 3635 2884 3899 2892
rect 3925 2892 3944 2895
rect 3951 2892 3978 2904
rect 3925 2884 3978 2892
rect 3553 2876 3554 2884
rect 3569 2876 3582 2884
rect 3553 2868 3569 2876
rect 3550 2861 3569 2864
rect 3550 2852 3572 2861
rect 3523 2842 3572 2852
rect 3523 2836 3553 2842
rect 3572 2837 3577 2842
rect 3495 2820 3569 2836
rect 3587 2828 3617 2884
rect 3652 2874 3860 2884
rect 3895 2880 3940 2884
rect 3943 2883 3944 2884
rect 3959 2883 3972 2884
rect 3678 2844 3867 2874
rect 3693 2841 3867 2844
rect 3686 2838 3867 2841
rect 3495 2818 3508 2820
rect 3523 2818 3557 2820
rect 3495 2802 3569 2818
rect 3596 2814 3609 2828
rect 3624 2814 3640 2830
rect 3686 2825 3697 2838
rect 3479 2780 3480 2796
rect 3495 2780 3508 2802
rect 3523 2780 3553 2802
rect 3596 2798 3658 2814
rect 3686 2807 3697 2823
rect 3702 2818 3712 2838
rect 3722 2818 3736 2838
rect 3739 2825 3748 2838
rect 3764 2825 3773 2838
rect 3702 2807 3736 2818
rect 3739 2807 3748 2823
rect 3764 2807 3773 2823
rect 3780 2818 3790 2838
rect 3800 2818 3814 2838
rect 3815 2825 3826 2838
rect 3780 2807 3814 2818
rect 3815 2807 3826 2823
rect 3872 2814 3888 2830
rect 3895 2828 3925 2880
rect 3959 2876 3960 2883
rect 3944 2868 3960 2876
rect 3931 2836 3944 2855
rect 3959 2836 3989 2852
rect 3931 2820 4005 2836
rect 3931 2818 3944 2820
rect 3959 2818 3993 2820
rect 3596 2796 3609 2798
rect 3624 2796 3658 2798
rect 3596 2780 3658 2796
rect 3702 2791 3718 2794
rect 3780 2791 3810 2802
rect 3858 2798 3904 2814
rect 3931 2802 4005 2818
rect 3858 2796 3892 2798
rect 3857 2780 3904 2796
rect 3931 2780 3944 2802
rect 3959 2780 3989 2802
rect 4016 2780 4017 2796
rect 4032 2780 4045 2940
rect 4075 2836 4088 2940
rect 4133 2918 4134 2928
rect 4149 2918 4162 2928
rect 4133 2914 4162 2918
rect 4167 2914 4197 2940
rect 4215 2926 4231 2928
rect 4303 2926 4356 2940
rect 4304 2924 4368 2926
rect 4411 2924 4426 2940
rect 4475 2937 4505 2940
rect 4475 2934 4511 2937
rect 4441 2926 4457 2928
rect 4215 2914 4230 2918
rect 4133 2912 4230 2914
rect 4258 2912 4426 2924
rect 4442 2914 4457 2918
rect 4475 2915 4514 2934
rect 4533 2928 4540 2929
rect 4539 2921 4540 2928
rect 4523 2918 4524 2921
rect 4539 2918 4552 2921
rect 4475 2914 4505 2915
rect 4514 2914 4520 2915
rect 4523 2914 4552 2918
rect 4442 2913 4552 2914
rect 4442 2912 4558 2913
rect 4117 2904 4168 2912
rect 4117 2892 4142 2904
rect 4149 2892 4168 2904
rect 4199 2904 4249 2912
rect 4199 2896 4215 2904
rect 4222 2902 4249 2904
rect 4258 2902 4479 2912
rect 4222 2892 4479 2902
rect 4508 2904 4558 2912
rect 4508 2895 4524 2904
rect 4117 2884 4168 2892
rect 4215 2884 4479 2892
rect 4505 2892 4524 2895
rect 4531 2892 4558 2904
rect 4505 2884 4558 2892
rect 4133 2876 4134 2884
rect 4149 2876 4162 2884
rect 4133 2868 4149 2876
rect 4130 2861 4149 2864
rect 4130 2852 4152 2861
rect 4103 2842 4152 2852
rect 4103 2836 4133 2842
rect 4152 2837 4157 2842
rect 4075 2820 4149 2836
rect 4167 2828 4197 2884
rect 4232 2874 4440 2884
rect 4475 2880 4520 2884
rect 4523 2883 4524 2884
rect 4539 2883 4552 2884
rect 4258 2844 4447 2874
rect 4273 2841 4447 2844
rect 4266 2838 4447 2841
rect 4075 2818 4088 2820
rect 4103 2818 4137 2820
rect 4075 2802 4149 2818
rect 4176 2814 4189 2828
rect 4204 2814 4220 2830
rect 4266 2825 4277 2838
rect 4059 2780 4060 2796
rect 4075 2780 4088 2802
rect 4103 2780 4133 2802
rect 4176 2798 4238 2814
rect 4266 2807 4277 2823
rect 4282 2818 4292 2838
rect 4302 2818 4316 2838
rect 4319 2825 4328 2838
rect 4344 2825 4353 2838
rect 4282 2807 4316 2818
rect 4319 2807 4328 2823
rect 4344 2807 4353 2823
rect 4360 2818 4370 2838
rect 4380 2818 4394 2838
rect 4395 2825 4406 2838
rect 4360 2807 4394 2818
rect 4395 2807 4406 2823
rect 4452 2814 4468 2830
rect 4475 2828 4505 2880
rect 4539 2876 4540 2883
rect 4524 2868 4540 2876
rect 4511 2836 4524 2855
rect 4539 2836 4569 2852
rect 4511 2820 4585 2836
rect 4511 2818 4524 2820
rect 4539 2818 4573 2820
rect 4176 2796 4189 2798
rect 4204 2796 4238 2798
rect 4176 2780 4238 2796
rect 4282 2791 4298 2794
rect 4360 2791 4390 2802
rect 4438 2798 4484 2814
rect 4511 2802 4585 2818
rect 4438 2796 4472 2798
rect 4437 2780 4484 2796
rect 4511 2780 4524 2802
rect 4539 2780 4569 2802
rect 4596 2780 4597 2796
rect 4612 2780 4625 2940
rect 4655 2836 4668 2940
rect 4713 2918 4714 2928
rect 4729 2918 4742 2928
rect 4713 2914 4742 2918
rect 4747 2914 4777 2940
rect 4795 2926 4811 2928
rect 4883 2926 4936 2940
rect 4884 2924 4948 2926
rect 4991 2924 5006 2940
rect 5055 2937 5085 2940
rect 5055 2934 5091 2937
rect 5021 2926 5037 2928
rect 4795 2914 4810 2918
rect 4713 2912 4810 2914
rect 4838 2912 5006 2924
rect 5022 2914 5037 2918
rect 5055 2915 5094 2934
rect 5113 2928 5120 2929
rect 5119 2921 5120 2928
rect 5103 2918 5104 2921
rect 5119 2918 5132 2921
rect 5055 2914 5085 2915
rect 5094 2914 5100 2915
rect 5103 2914 5132 2918
rect 5022 2913 5132 2914
rect 5022 2912 5138 2913
rect 4697 2904 4748 2912
rect 4697 2892 4722 2904
rect 4729 2892 4748 2904
rect 4779 2904 4829 2912
rect 4779 2896 4795 2904
rect 4802 2902 4829 2904
rect 4838 2902 5059 2912
rect 4802 2892 5059 2902
rect 5088 2904 5138 2912
rect 5088 2895 5104 2904
rect 4697 2884 4748 2892
rect 4795 2884 5059 2892
rect 5085 2892 5104 2895
rect 5111 2892 5138 2904
rect 5085 2884 5138 2892
rect 4713 2876 4714 2884
rect 4729 2876 4742 2884
rect 4713 2868 4729 2876
rect 4710 2861 4729 2864
rect 4710 2852 4732 2861
rect 4683 2842 4732 2852
rect 4683 2836 4713 2842
rect 4732 2837 4737 2842
rect 4655 2820 4729 2836
rect 4747 2828 4777 2884
rect 4812 2874 5020 2884
rect 5055 2880 5100 2884
rect 5103 2883 5104 2884
rect 5119 2883 5132 2884
rect 4838 2844 5027 2874
rect 4853 2841 5027 2844
rect 4846 2838 5027 2841
rect 4655 2818 4668 2820
rect 4683 2818 4717 2820
rect 4655 2802 4729 2818
rect 4756 2814 4769 2828
rect 4784 2814 4800 2830
rect 4846 2825 4857 2838
rect 4639 2780 4640 2796
rect 4655 2780 4668 2802
rect 4683 2780 4713 2802
rect 4756 2798 4818 2814
rect 4846 2807 4857 2823
rect 4862 2818 4872 2838
rect 4882 2818 4896 2838
rect 4899 2825 4908 2838
rect 4924 2825 4933 2838
rect 4862 2807 4896 2818
rect 4899 2807 4908 2823
rect 4924 2807 4933 2823
rect 4940 2818 4950 2838
rect 4960 2818 4974 2838
rect 4975 2825 4986 2838
rect 4940 2807 4974 2818
rect 4975 2807 4986 2823
rect 5032 2814 5048 2830
rect 5055 2828 5085 2880
rect 5119 2876 5120 2883
rect 5104 2868 5120 2876
rect 5091 2836 5104 2855
rect 5119 2836 5149 2852
rect 5091 2820 5165 2836
rect 5091 2818 5104 2820
rect 5119 2818 5153 2820
rect 4756 2796 4769 2798
rect 4784 2796 4818 2798
rect 4756 2780 4818 2796
rect 4862 2791 4878 2794
rect 4940 2791 4970 2802
rect 5018 2798 5064 2814
rect 5091 2802 5165 2818
rect 5018 2796 5052 2798
rect 5017 2780 5064 2796
rect 5091 2780 5104 2802
rect 5119 2780 5149 2802
rect 5176 2780 5177 2796
rect 5192 2780 5205 2940
rect 5235 2836 5248 2940
rect 5293 2918 5294 2928
rect 5309 2918 5322 2928
rect 5293 2914 5322 2918
rect 5327 2914 5357 2940
rect 5375 2926 5391 2928
rect 5463 2926 5516 2940
rect 5464 2924 5528 2926
rect 5571 2924 5586 2940
rect 5635 2937 5665 2940
rect 5635 2934 5671 2937
rect 5601 2926 5617 2928
rect 5375 2914 5390 2918
rect 5293 2912 5390 2914
rect 5418 2912 5586 2924
rect 5602 2914 5617 2918
rect 5635 2915 5674 2934
rect 5693 2928 5700 2929
rect 5699 2921 5700 2928
rect 5683 2918 5684 2921
rect 5699 2918 5712 2921
rect 5635 2914 5665 2915
rect 5674 2914 5680 2915
rect 5683 2914 5712 2918
rect 5602 2913 5712 2914
rect 5602 2912 5718 2913
rect 5277 2904 5328 2912
rect 5277 2892 5302 2904
rect 5309 2892 5328 2904
rect 5359 2904 5409 2912
rect 5359 2896 5375 2904
rect 5382 2902 5409 2904
rect 5418 2902 5639 2912
rect 5382 2892 5639 2902
rect 5668 2904 5718 2912
rect 5668 2895 5684 2904
rect 5277 2884 5328 2892
rect 5375 2884 5639 2892
rect 5665 2892 5684 2895
rect 5691 2892 5718 2904
rect 5665 2884 5718 2892
rect 5293 2876 5294 2884
rect 5309 2876 5322 2884
rect 5293 2868 5309 2876
rect 5290 2861 5309 2864
rect 5290 2852 5312 2861
rect 5263 2842 5312 2852
rect 5263 2836 5293 2842
rect 5312 2837 5317 2842
rect 5235 2820 5309 2836
rect 5327 2828 5357 2884
rect 5392 2874 5600 2884
rect 5635 2880 5680 2884
rect 5683 2883 5684 2884
rect 5699 2883 5712 2884
rect 5418 2844 5607 2874
rect 5433 2841 5607 2844
rect 5426 2838 5607 2841
rect 5235 2818 5248 2820
rect 5263 2818 5297 2820
rect 5235 2802 5309 2818
rect 5336 2814 5349 2828
rect 5364 2814 5380 2830
rect 5426 2825 5437 2838
rect 5219 2780 5220 2796
rect 5235 2780 5248 2802
rect 5263 2780 5293 2802
rect 5336 2798 5398 2814
rect 5426 2807 5437 2823
rect 5442 2818 5452 2838
rect 5462 2818 5476 2838
rect 5479 2825 5488 2838
rect 5504 2825 5513 2838
rect 5442 2807 5476 2818
rect 5479 2807 5488 2823
rect 5504 2807 5513 2823
rect 5520 2818 5530 2838
rect 5540 2818 5554 2838
rect 5555 2825 5566 2838
rect 5520 2807 5554 2818
rect 5555 2807 5566 2823
rect 5612 2814 5628 2830
rect 5635 2828 5665 2880
rect 5699 2876 5700 2883
rect 5684 2868 5700 2876
rect 5671 2836 5684 2855
rect 5699 2836 5729 2852
rect 5671 2820 5745 2836
rect 5671 2818 5684 2820
rect 5699 2818 5733 2820
rect 5336 2796 5349 2798
rect 5364 2796 5398 2798
rect 5336 2780 5398 2796
rect 5442 2791 5458 2794
rect 5520 2791 5550 2802
rect 5598 2798 5644 2814
rect 5671 2802 5745 2818
rect 5598 2796 5632 2798
rect 5597 2780 5644 2796
rect 5671 2780 5684 2802
rect 5699 2780 5729 2802
rect 5756 2780 5757 2796
rect 5772 2780 5785 2940
rect 5815 2836 5828 2940
rect 5873 2918 5874 2928
rect 5889 2918 5902 2928
rect 5873 2914 5902 2918
rect 5907 2914 5937 2940
rect 5955 2926 5971 2928
rect 6043 2926 6096 2940
rect 6044 2924 6108 2926
rect 6151 2924 6166 2940
rect 6215 2937 6245 2940
rect 6215 2934 6251 2937
rect 6181 2926 6197 2928
rect 5955 2914 5970 2918
rect 5873 2912 5970 2914
rect 5998 2912 6166 2924
rect 6182 2914 6197 2918
rect 6215 2915 6254 2934
rect 6273 2928 6280 2929
rect 6279 2921 6280 2928
rect 6263 2918 6264 2921
rect 6279 2918 6292 2921
rect 6215 2914 6245 2915
rect 6254 2914 6260 2915
rect 6263 2914 6292 2918
rect 6182 2913 6292 2914
rect 6182 2912 6298 2913
rect 5857 2904 5908 2912
rect 5857 2892 5882 2904
rect 5889 2892 5908 2904
rect 5939 2904 5989 2912
rect 5939 2896 5955 2904
rect 5962 2902 5989 2904
rect 5998 2902 6219 2912
rect 5962 2892 6219 2902
rect 6248 2904 6298 2912
rect 6248 2895 6264 2904
rect 5857 2884 5908 2892
rect 5955 2884 6219 2892
rect 6245 2892 6264 2895
rect 6271 2892 6298 2904
rect 6245 2884 6298 2892
rect 5873 2876 5874 2884
rect 5889 2876 5902 2884
rect 5873 2868 5889 2876
rect 5870 2861 5889 2864
rect 5870 2852 5892 2861
rect 5843 2842 5892 2852
rect 5843 2836 5873 2842
rect 5892 2837 5897 2842
rect 5815 2820 5889 2836
rect 5907 2828 5937 2884
rect 5972 2874 6180 2884
rect 6215 2880 6260 2884
rect 6263 2883 6264 2884
rect 6279 2883 6292 2884
rect 5998 2844 6187 2874
rect 6013 2841 6187 2844
rect 6006 2838 6187 2841
rect 5815 2818 5828 2820
rect 5843 2818 5877 2820
rect 5815 2802 5889 2818
rect 5916 2814 5929 2828
rect 5944 2814 5960 2830
rect 6006 2825 6017 2838
rect 5799 2780 5800 2796
rect 5815 2780 5828 2802
rect 5843 2780 5873 2802
rect 5916 2798 5978 2814
rect 6006 2807 6017 2823
rect 6022 2818 6032 2838
rect 6042 2818 6056 2838
rect 6059 2825 6068 2838
rect 6084 2825 6093 2838
rect 6022 2807 6056 2818
rect 6059 2807 6068 2823
rect 6084 2807 6093 2823
rect 6100 2818 6110 2838
rect 6120 2818 6134 2838
rect 6135 2825 6146 2838
rect 6100 2807 6134 2818
rect 6135 2807 6146 2823
rect 6192 2814 6208 2830
rect 6215 2828 6245 2880
rect 6279 2876 6280 2883
rect 6264 2868 6280 2876
rect 6251 2836 6264 2855
rect 6279 2836 6309 2852
rect 6251 2820 6325 2836
rect 6251 2818 6264 2820
rect 6279 2818 6313 2820
rect 5916 2796 5929 2798
rect 5944 2796 5978 2798
rect 5916 2780 5978 2796
rect 6022 2791 6038 2794
rect 6100 2791 6130 2802
rect 6178 2798 6224 2814
rect 6251 2802 6325 2818
rect 6178 2796 6212 2798
rect 6177 2780 6224 2796
rect 6251 2780 6264 2802
rect 6279 2780 6309 2802
rect 6336 2780 6337 2796
rect 6352 2780 6365 2940
rect 6395 2836 6408 2940
rect 6453 2918 6454 2928
rect 6469 2918 6482 2928
rect 6453 2914 6482 2918
rect 6487 2914 6517 2940
rect 6535 2926 6551 2928
rect 6623 2926 6676 2940
rect 6624 2924 6688 2926
rect 6731 2924 6746 2940
rect 6795 2937 6825 2940
rect 6795 2934 6831 2937
rect 6761 2926 6777 2928
rect 6535 2914 6550 2918
rect 6453 2912 6550 2914
rect 6578 2912 6746 2924
rect 6762 2914 6777 2918
rect 6795 2915 6834 2934
rect 6853 2928 6860 2929
rect 6859 2921 6860 2928
rect 6843 2918 6844 2921
rect 6859 2918 6872 2921
rect 6795 2914 6825 2915
rect 6834 2914 6840 2915
rect 6843 2914 6872 2918
rect 6762 2913 6872 2914
rect 6762 2912 6878 2913
rect 6437 2904 6488 2912
rect 6437 2892 6462 2904
rect 6469 2892 6488 2904
rect 6519 2904 6569 2912
rect 6519 2896 6535 2904
rect 6542 2902 6569 2904
rect 6578 2902 6799 2912
rect 6542 2892 6799 2902
rect 6828 2904 6878 2912
rect 6828 2895 6844 2904
rect 6437 2884 6488 2892
rect 6535 2884 6799 2892
rect 6825 2892 6844 2895
rect 6851 2892 6878 2904
rect 6825 2884 6878 2892
rect 6453 2876 6454 2884
rect 6469 2876 6482 2884
rect 6453 2868 6469 2876
rect 6450 2861 6469 2864
rect 6450 2852 6472 2861
rect 6423 2842 6472 2852
rect 6423 2836 6453 2842
rect 6472 2837 6477 2842
rect 6395 2820 6469 2836
rect 6487 2828 6517 2884
rect 6552 2874 6760 2884
rect 6795 2880 6840 2884
rect 6843 2883 6844 2884
rect 6859 2883 6872 2884
rect 6578 2844 6767 2874
rect 6593 2841 6767 2844
rect 6586 2838 6767 2841
rect 6395 2818 6408 2820
rect 6423 2818 6457 2820
rect 6395 2802 6469 2818
rect 6496 2814 6509 2828
rect 6524 2814 6540 2830
rect 6586 2825 6597 2838
rect 6379 2780 6380 2796
rect 6395 2780 6408 2802
rect 6423 2780 6453 2802
rect 6496 2798 6558 2814
rect 6586 2807 6597 2823
rect 6602 2818 6612 2838
rect 6622 2818 6636 2838
rect 6639 2825 6648 2838
rect 6664 2825 6673 2838
rect 6602 2807 6636 2818
rect 6639 2807 6648 2823
rect 6664 2807 6673 2823
rect 6680 2818 6690 2838
rect 6700 2818 6714 2838
rect 6715 2825 6726 2838
rect 6680 2807 6714 2818
rect 6715 2807 6726 2823
rect 6772 2814 6788 2830
rect 6795 2828 6825 2880
rect 6859 2876 6860 2883
rect 6844 2868 6860 2876
rect 6831 2836 6844 2855
rect 6859 2836 6889 2852
rect 6831 2820 6905 2836
rect 6831 2818 6844 2820
rect 6859 2818 6893 2820
rect 6496 2796 6509 2798
rect 6524 2796 6558 2798
rect 6496 2780 6558 2796
rect 6602 2791 6618 2794
rect 6680 2791 6710 2802
rect 6758 2798 6804 2814
rect 6831 2802 6905 2818
rect 6758 2796 6792 2798
rect 6757 2780 6804 2796
rect 6831 2780 6844 2802
rect 6859 2780 6889 2802
rect 6916 2780 6917 2796
rect 6932 2780 6945 2940
rect 6975 2836 6988 2940
rect 7033 2918 7034 2928
rect 7049 2918 7062 2928
rect 7033 2914 7062 2918
rect 7067 2914 7097 2940
rect 7115 2926 7131 2928
rect 7203 2926 7256 2940
rect 7204 2924 7268 2926
rect 7311 2924 7326 2940
rect 7375 2937 7405 2940
rect 7375 2934 7411 2937
rect 7341 2926 7357 2928
rect 7115 2914 7130 2918
rect 7033 2912 7130 2914
rect 7158 2912 7326 2924
rect 7342 2914 7357 2918
rect 7375 2915 7414 2934
rect 7433 2928 7440 2929
rect 7439 2921 7440 2928
rect 7423 2918 7424 2921
rect 7439 2918 7452 2921
rect 7375 2914 7405 2915
rect 7414 2914 7420 2915
rect 7423 2914 7452 2918
rect 7342 2913 7452 2914
rect 7342 2912 7458 2913
rect 7017 2904 7068 2912
rect 7017 2892 7042 2904
rect 7049 2892 7068 2904
rect 7099 2904 7149 2912
rect 7099 2896 7115 2904
rect 7122 2902 7149 2904
rect 7158 2902 7379 2912
rect 7122 2892 7379 2902
rect 7408 2904 7458 2912
rect 7408 2895 7424 2904
rect 7017 2884 7068 2892
rect 7115 2884 7379 2892
rect 7405 2892 7424 2895
rect 7431 2892 7458 2904
rect 7405 2884 7458 2892
rect 7033 2876 7034 2884
rect 7049 2876 7062 2884
rect 7033 2868 7049 2876
rect 7030 2861 7049 2864
rect 7030 2852 7052 2861
rect 7003 2842 7052 2852
rect 7003 2836 7033 2842
rect 7052 2837 7057 2842
rect 6975 2820 7049 2836
rect 7067 2828 7097 2884
rect 7132 2874 7340 2884
rect 7375 2880 7420 2884
rect 7423 2883 7424 2884
rect 7439 2883 7452 2884
rect 7158 2844 7347 2874
rect 7173 2841 7347 2844
rect 7166 2838 7347 2841
rect 6975 2818 6988 2820
rect 7003 2818 7037 2820
rect 6975 2802 7049 2818
rect 7076 2814 7089 2828
rect 7104 2814 7120 2830
rect 7166 2825 7177 2838
rect 6959 2780 6960 2796
rect 6975 2780 6988 2802
rect 7003 2780 7033 2802
rect 7076 2798 7138 2814
rect 7166 2807 7177 2823
rect 7182 2818 7192 2838
rect 7202 2818 7216 2838
rect 7219 2825 7228 2838
rect 7244 2825 7253 2838
rect 7182 2807 7216 2818
rect 7219 2807 7228 2823
rect 7244 2807 7253 2823
rect 7260 2818 7270 2838
rect 7280 2818 7294 2838
rect 7295 2825 7306 2838
rect 7260 2807 7294 2818
rect 7295 2807 7306 2823
rect 7352 2814 7368 2830
rect 7375 2828 7405 2880
rect 7439 2876 7440 2883
rect 7424 2868 7440 2876
rect 7411 2836 7424 2855
rect 7439 2836 7469 2852
rect 7411 2820 7485 2836
rect 7411 2818 7424 2820
rect 7439 2818 7473 2820
rect 7076 2796 7089 2798
rect 7104 2796 7138 2798
rect 7076 2780 7138 2796
rect 7182 2791 7198 2794
rect 7260 2791 7290 2802
rect 7338 2798 7384 2814
rect 7411 2802 7485 2818
rect 7338 2796 7372 2798
rect 7337 2780 7384 2796
rect 7411 2780 7424 2802
rect 7439 2780 7469 2802
rect 7496 2780 7497 2796
rect 7512 2780 7525 2940
rect 7555 2836 7568 2940
rect 7613 2918 7614 2928
rect 7629 2918 7642 2928
rect 7613 2914 7642 2918
rect 7647 2914 7677 2940
rect 7695 2926 7711 2928
rect 7783 2926 7836 2940
rect 7784 2924 7848 2926
rect 7891 2924 7906 2940
rect 7955 2937 7985 2940
rect 7955 2934 7991 2937
rect 7921 2926 7937 2928
rect 7695 2914 7710 2918
rect 7613 2912 7710 2914
rect 7738 2912 7906 2924
rect 7922 2914 7937 2918
rect 7955 2915 7994 2934
rect 8013 2928 8020 2929
rect 8019 2921 8020 2928
rect 8003 2918 8004 2921
rect 8019 2918 8032 2921
rect 7955 2914 7985 2915
rect 7994 2914 8000 2915
rect 8003 2914 8032 2918
rect 7922 2913 8032 2914
rect 7922 2912 8038 2913
rect 7597 2904 7648 2912
rect 7597 2892 7622 2904
rect 7629 2892 7648 2904
rect 7679 2904 7729 2912
rect 7679 2896 7695 2904
rect 7702 2902 7729 2904
rect 7738 2902 7959 2912
rect 7702 2892 7959 2902
rect 7988 2904 8038 2912
rect 7988 2895 8004 2904
rect 7597 2884 7648 2892
rect 7695 2884 7959 2892
rect 7985 2892 8004 2895
rect 8011 2892 8038 2904
rect 7985 2884 8038 2892
rect 7613 2876 7614 2884
rect 7629 2876 7642 2884
rect 7613 2868 7629 2876
rect 7610 2861 7629 2864
rect 7610 2852 7632 2861
rect 7583 2842 7632 2852
rect 7583 2836 7613 2842
rect 7632 2837 7637 2842
rect 7555 2820 7629 2836
rect 7647 2828 7677 2884
rect 7712 2874 7920 2884
rect 7955 2880 8000 2884
rect 8003 2883 8004 2884
rect 8019 2883 8032 2884
rect 7738 2844 7927 2874
rect 7753 2841 7927 2844
rect 7746 2838 7927 2841
rect 7555 2818 7568 2820
rect 7583 2818 7617 2820
rect 7555 2802 7629 2818
rect 7656 2814 7669 2828
rect 7684 2814 7700 2830
rect 7746 2825 7757 2838
rect 7539 2780 7540 2796
rect 7555 2780 7568 2802
rect 7583 2780 7613 2802
rect 7656 2798 7718 2814
rect 7746 2807 7757 2823
rect 7762 2818 7772 2838
rect 7782 2818 7796 2838
rect 7799 2825 7808 2838
rect 7824 2825 7833 2838
rect 7762 2807 7796 2818
rect 7799 2807 7808 2823
rect 7824 2807 7833 2823
rect 7840 2818 7850 2838
rect 7860 2818 7874 2838
rect 7875 2825 7886 2838
rect 7840 2807 7874 2818
rect 7875 2807 7886 2823
rect 7932 2814 7948 2830
rect 7955 2828 7985 2880
rect 8019 2876 8020 2883
rect 8004 2868 8020 2876
rect 7991 2836 8004 2855
rect 8019 2836 8049 2852
rect 7991 2820 8065 2836
rect 7991 2818 8004 2820
rect 8019 2818 8053 2820
rect 7656 2796 7669 2798
rect 7684 2796 7718 2798
rect 7656 2780 7718 2796
rect 7762 2791 7778 2794
rect 7840 2791 7870 2802
rect 7918 2798 7964 2814
rect 7991 2802 8065 2818
rect 7918 2796 7952 2798
rect 7917 2780 7964 2796
rect 7991 2780 8004 2802
rect 8019 2780 8049 2802
rect 8076 2780 8077 2796
rect 8092 2780 8105 2940
rect 8135 2836 8148 2940
rect 8193 2918 8194 2928
rect 8209 2918 8222 2928
rect 8193 2914 8222 2918
rect 8227 2914 8257 2940
rect 8275 2926 8291 2928
rect 8363 2926 8416 2940
rect 8364 2924 8428 2926
rect 8471 2924 8486 2940
rect 8535 2937 8565 2940
rect 8535 2934 8571 2937
rect 8501 2926 8517 2928
rect 8275 2914 8290 2918
rect 8193 2912 8290 2914
rect 8318 2912 8486 2924
rect 8502 2914 8517 2918
rect 8535 2915 8574 2934
rect 8593 2928 8600 2929
rect 8599 2921 8600 2928
rect 8583 2918 8584 2921
rect 8599 2918 8612 2921
rect 8535 2914 8565 2915
rect 8574 2914 8580 2915
rect 8583 2914 8612 2918
rect 8502 2913 8612 2914
rect 8502 2912 8618 2913
rect 8177 2904 8228 2912
rect 8177 2892 8202 2904
rect 8209 2892 8228 2904
rect 8259 2904 8309 2912
rect 8259 2896 8275 2904
rect 8282 2902 8309 2904
rect 8318 2902 8539 2912
rect 8282 2892 8539 2902
rect 8568 2904 8618 2912
rect 8568 2895 8584 2904
rect 8177 2884 8228 2892
rect 8275 2884 8539 2892
rect 8565 2892 8584 2895
rect 8591 2892 8618 2904
rect 8565 2884 8618 2892
rect 8193 2876 8194 2884
rect 8209 2876 8222 2884
rect 8193 2868 8209 2876
rect 8190 2861 8209 2864
rect 8190 2852 8212 2861
rect 8163 2842 8212 2852
rect 8163 2836 8193 2842
rect 8212 2837 8217 2842
rect 8135 2820 8209 2836
rect 8227 2828 8257 2884
rect 8292 2874 8500 2884
rect 8535 2880 8580 2884
rect 8583 2883 8584 2884
rect 8599 2883 8612 2884
rect 8318 2844 8507 2874
rect 8333 2841 8507 2844
rect 8326 2838 8507 2841
rect 8135 2818 8148 2820
rect 8163 2818 8197 2820
rect 8135 2802 8209 2818
rect 8236 2814 8249 2828
rect 8264 2814 8280 2830
rect 8326 2825 8337 2838
rect 8119 2780 8120 2796
rect 8135 2780 8148 2802
rect 8163 2780 8193 2802
rect 8236 2798 8298 2814
rect 8326 2807 8337 2823
rect 8342 2818 8352 2838
rect 8362 2818 8376 2838
rect 8379 2825 8388 2838
rect 8404 2825 8413 2838
rect 8342 2807 8376 2818
rect 8379 2807 8388 2823
rect 8404 2807 8413 2823
rect 8420 2818 8430 2838
rect 8440 2818 8454 2838
rect 8455 2825 8466 2838
rect 8420 2807 8454 2818
rect 8455 2807 8466 2823
rect 8512 2814 8528 2830
rect 8535 2828 8565 2880
rect 8599 2876 8600 2883
rect 8584 2868 8600 2876
rect 8571 2836 8584 2855
rect 8599 2836 8629 2852
rect 8571 2820 8645 2836
rect 8571 2818 8584 2820
rect 8599 2818 8633 2820
rect 8236 2796 8249 2798
rect 8264 2796 8298 2798
rect 8236 2780 8298 2796
rect 8342 2791 8358 2794
rect 8420 2791 8450 2802
rect 8498 2798 8544 2814
rect 8571 2802 8645 2818
rect 8498 2796 8532 2798
rect 8497 2780 8544 2796
rect 8571 2780 8584 2802
rect 8599 2780 8629 2802
rect 8656 2780 8657 2796
rect 8672 2780 8685 2940
rect 8715 2836 8728 2940
rect 8773 2918 8774 2928
rect 8789 2918 8802 2928
rect 8773 2914 8802 2918
rect 8807 2914 8837 2940
rect 8855 2926 8871 2928
rect 8943 2926 8996 2940
rect 8944 2924 9008 2926
rect 9051 2924 9066 2940
rect 9115 2937 9145 2940
rect 9115 2934 9151 2937
rect 9081 2926 9097 2928
rect 8855 2914 8870 2918
rect 8773 2912 8870 2914
rect 8898 2912 9066 2924
rect 9082 2914 9097 2918
rect 9115 2915 9154 2934
rect 9173 2928 9180 2929
rect 9179 2921 9180 2928
rect 9163 2918 9164 2921
rect 9179 2918 9192 2921
rect 9115 2914 9145 2915
rect 9154 2914 9160 2915
rect 9163 2914 9192 2918
rect 9082 2913 9192 2914
rect 9082 2912 9198 2913
rect 8757 2904 8808 2912
rect 8757 2892 8782 2904
rect 8789 2892 8808 2904
rect 8839 2904 8889 2912
rect 8839 2896 8855 2904
rect 8862 2902 8889 2904
rect 8898 2902 9119 2912
rect 8862 2892 9119 2902
rect 9148 2904 9198 2912
rect 9148 2895 9164 2904
rect 8757 2884 8808 2892
rect 8855 2884 9119 2892
rect 9145 2892 9164 2895
rect 9171 2892 9198 2904
rect 9145 2884 9198 2892
rect 8773 2876 8774 2884
rect 8789 2876 8802 2884
rect 8773 2868 8789 2876
rect 8770 2861 8789 2864
rect 8770 2852 8792 2861
rect 8743 2842 8792 2852
rect 8743 2836 8773 2842
rect 8792 2837 8797 2842
rect 8715 2820 8789 2836
rect 8807 2828 8837 2884
rect 8872 2874 9080 2884
rect 9115 2880 9160 2884
rect 9163 2883 9164 2884
rect 9179 2883 9192 2884
rect 8898 2844 9087 2874
rect 8913 2841 9087 2844
rect 8906 2838 9087 2841
rect 8715 2818 8728 2820
rect 8743 2818 8777 2820
rect 8715 2802 8789 2818
rect 8816 2814 8829 2828
rect 8844 2814 8860 2830
rect 8906 2825 8917 2838
rect 8699 2780 8700 2796
rect 8715 2780 8728 2802
rect 8743 2780 8773 2802
rect 8816 2798 8878 2814
rect 8906 2807 8917 2823
rect 8922 2818 8932 2838
rect 8942 2818 8956 2838
rect 8959 2825 8968 2838
rect 8984 2825 8993 2838
rect 8922 2807 8956 2818
rect 8959 2807 8968 2823
rect 8984 2807 8993 2823
rect 9000 2818 9010 2838
rect 9020 2818 9034 2838
rect 9035 2825 9046 2838
rect 9000 2807 9034 2818
rect 9035 2807 9046 2823
rect 9092 2814 9108 2830
rect 9115 2828 9145 2880
rect 9179 2876 9180 2883
rect 9164 2868 9180 2876
rect 9151 2836 9164 2855
rect 9179 2836 9209 2852
rect 9151 2820 9225 2836
rect 9151 2818 9164 2820
rect 9179 2818 9213 2820
rect 8816 2796 8829 2798
rect 8844 2796 8878 2798
rect 8816 2780 8878 2796
rect 8922 2791 8938 2794
rect 9000 2791 9030 2802
rect 9078 2798 9124 2814
rect 9151 2802 9225 2818
rect 9078 2796 9112 2798
rect 9077 2780 9124 2796
rect 9151 2780 9164 2802
rect 9179 2780 9209 2802
rect 9236 2780 9237 2796
rect 9252 2780 9265 2940
rect -7 2772 34 2780
rect -7 2746 8 2772
rect 15 2746 34 2772
rect 98 2768 160 2780
rect 172 2768 247 2780
rect 305 2768 380 2780
rect 392 2768 423 2780
rect 429 2768 464 2780
rect 98 2766 260 2768
rect -7 2738 34 2746
rect 116 2742 129 2766
rect 144 2764 159 2766
rect -1 2728 0 2738
rect 15 2728 28 2738
rect 43 2728 73 2742
rect 116 2728 159 2742
rect 183 2739 190 2746
rect 193 2742 260 2766
rect 292 2766 464 2768
rect 262 2744 290 2748
rect 292 2744 372 2766
rect 393 2764 408 2766
rect 262 2742 372 2744
rect 193 2738 372 2742
rect 166 2728 196 2738
rect 198 2728 351 2738
rect 359 2728 389 2738
rect 393 2728 423 2742
rect 451 2728 464 2766
rect 536 2772 571 2780
rect 536 2746 537 2772
rect 544 2746 571 2772
rect 479 2728 509 2742
rect 536 2738 571 2746
rect 573 2772 614 2780
rect 573 2746 588 2772
rect 595 2746 614 2772
rect 678 2768 740 2780
rect 752 2768 827 2780
rect 885 2768 960 2780
rect 972 2768 1003 2780
rect 1009 2768 1044 2780
rect 678 2766 840 2768
rect 573 2738 614 2746
rect 696 2742 709 2766
rect 724 2764 739 2766
rect 536 2728 537 2738
rect 552 2728 565 2738
rect 579 2728 580 2738
rect 595 2728 608 2738
rect 623 2728 653 2742
rect 696 2728 739 2742
rect 763 2739 770 2746
rect 773 2742 840 2766
rect 872 2766 1044 2768
rect 842 2744 870 2748
rect 872 2744 952 2766
rect 973 2764 988 2766
rect 842 2742 952 2744
rect 773 2738 952 2742
rect 746 2728 776 2738
rect 778 2728 931 2738
rect 939 2728 969 2738
rect 973 2728 1003 2742
rect 1031 2728 1044 2766
rect 1116 2772 1151 2780
rect 1116 2746 1117 2772
rect 1124 2746 1151 2772
rect 1059 2728 1089 2742
rect 1116 2738 1151 2746
rect 1153 2772 1194 2780
rect 1153 2746 1168 2772
rect 1175 2746 1194 2772
rect 1258 2768 1320 2780
rect 1332 2768 1407 2780
rect 1465 2768 1540 2780
rect 1552 2768 1583 2780
rect 1589 2768 1624 2780
rect 1258 2766 1420 2768
rect 1153 2738 1194 2746
rect 1276 2742 1289 2766
rect 1304 2764 1319 2766
rect 1116 2728 1117 2738
rect 1132 2728 1145 2738
rect 1159 2728 1160 2738
rect 1175 2728 1188 2738
rect 1203 2728 1233 2742
rect 1276 2728 1319 2742
rect 1343 2739 1350 2746
rect 1353 2742 1420 2766
rect 1452 2766 1624 2768
rect 1422 2744 1450 2748
rect 1452 2744 1532 2766
rect 1553 2764 1568 2766
rect 1422 2742 1532 2744
rect 1353 2738 1532 2742
rect 1326 2728 1356 2738
rect 1358 2728 1511 2738
rect 1519 2728 1549 2738
rect 1553 2728 1583 2742
rect 1611 2728 1624 2766
rect 1696 2772 1731 2780
rect 1696 2746 1697 2772
rect 1704 2746 1731 2772
rect 1639 2728 1669 2742
rect 1696 2738 1731 2746
rect 1733 2772 1774 2780
rect 1733 2746 1748 2772
rect 1755 2746 1774 2772
rect 1838 2768 1900 2780
rect 1912 2768 1987 2780
rect 2045 2768 2120 2780
rect 2132 2768 2163 2780
rect 2169 2768 2204 2780
rect 1838 2766 2000 2768
rect 1733 2738 1774 2746
rect 1856 2742 1869 2766
rect 1884 2764 1899 2766
rect 1696 2728 1697 2738
rect 1712 2728 1725 2738
rect 1739 2728 1740 2738
rect 1755 2728 1768 2738
rect 1783 2728 1813 2742
rect 1856 2728 1899 2742
rect 1923 2739 1930 2746
rect 1933 2742 2000 2766
rect 2032 2766 2204 2768
rect 2002 2744 2030 2748
rect 2032 2744 2112 2766
rect 2133 2764 2148 2766
rect 2002 2742 2112 2744
rect 1933 2738 2112 2742
rect 1906 2728 1936 2738
rect 1938 2728 2091 2738
rect 2099 2728 2129 2738
rect 2133 2728 2163 2742
rect 2191 2728 2204 2766
rect 2276 2772 2311 2780
rect 2276 2746 2277 2772
rect 2284 2746 2311 2772
rect 2219 2728 2249 2742
rect 2276 2738 2311 2746
rect 2313 2772 2354 2780
rect 2313 2746 2328 2772
rect 2335 2746 2354 2772
rect 2418 2768 2480 2780
rect 2492 2768 2567 2780
rect 2625 2768 2700 2780
rect 2712 2768 2743 2780
rect 2749 2768 2784 2780
rect 2418 2766 2580 2768
rect 2313 2738 2354 2746
rect 2436 2742 2449 2766
rect 2464 2764 2479 2766
rect 2276 2728 2277 2738
rect 2292 2728 2305 2738
rect 2319 2728 2320 2738
rect 2335 2728 2348 2738
rect 2363 2728 2393 2742
rect 2436 2728 2479 2742
rect 2503 2739 2510 2746
rect 2513 2742 2580 2766
rect 2612 2766 2784 2768
rect 2582 2744 2610 2748
rect 2612 2744 2692 2766
rect 2713 2764 2728 2766
rect 2582 2742 2692 2744
rect 2513 2738 2692 2742
rect 2486 2728 2516 2738
rect 2518 2728 2671 2738
rect 2679 2728 2709 2738
rect 2713 2728 2743 2742
rect 2771 2728 2784 2766
rect 2856 2772 2891 2780
rect 2856 2746 2857 2772
rect 2864 2746 2891 2772
rect 2799 2728 2829 2742
rect 2856 2738 2891 2746
rect 2893 2772 2934 2780
rect 2893 2746 2908 2772
rect 2915 2746 2934 2772
rect 2998 2768 3060 2780
rect 3072 2768 3147 2780
rect 3205 2768 3280 2780
rect 3292 2768 3323 2780
rect 3329 2768 3364 2780
rect 2998 2766 3160 2768
rect 2893 2738 2934 2746
rect 3016 2742 3029 2766
rect 3044 2764 3059 2766
rect 2856 2728 2857 2738
rect 2872 2728 2885 2738
rect 2899 2728 2900 2738
rect 2915 2728 2928 2738
rect 2943 2728 2973 2742
rect 3016 2728 3059 2742
rect 3083 2739 3090 2746
rect 3093 2742 3160 2766
rect 3192 2766 3364 2768
rect 3162 2744 3190 2748
rect 3192 2744 3272 2766
rect 3293 2764 3308 2766
rect 3162 2742 3272 2744
rect 3093 2738 3272 2742
rect 3066 2728 3096 2738
rect 3098 2728 3251 2738
rect 3259 2728 3289 2738
rect 3293 2728 3323 2742
rect 3351 2728 3364 2766
rect 3436 2772 3471 2780
rect 3436 2746 3437 2772
rect 3444 2746 3471 2772
rect 3379 2728 3409 2742
rect 3436 2738 3471 2746
rect 3473 2772 3514 2780
rect 3473 2746 3488 2772
rect 3495 2746 3514 2772
rect 3578 2768 3640 2780
rect 3652 2768 3727 2780
rect 3785 2768 3860 2780
rect 3872 2768 3903 2780
rect 3909 2768 3944 2780
rect 3578 2766 3740 2768
rect 3473 2738 3514 2746
rect 3596 2742 3609 2766
rect 3624 2764 3639 2766
rect 3436 2728 3437 2738
rect 3452 2728 3465 2738
rect 3479 2728 3480 2738
rect 3495 2728 3508 2738
rect 3523 2728 3553 2742
rect 3596 2728 3639 2742
rect 3663 2739 3670 2746
rect 3673 2742 3740 2766
rect 3772 2766 3944 2768
rect 3742 2744 3770 2748
rect 3772 2744 3852 2766
rect 3873 2764 3888 2766
rect 3742 2742 3852 2744
rect 3673 2738 3852 2742
rect 3646 2728 3676 2738
rect 3678 2728 3831 2738
rect 3839 2728 3869 2738
rect 3873 2728 3903 2742
rect 3931 2728 3944 2766
rect 4016 2772 4051 2780
rect 4016 2746 4017 2772
rect 4024 2746 4051 2772
rect 3959 2728 3989 2742
rect 4016 2738 4051 2746
rect 4053 2772 4094 2780
rect 4053 2746 4068 2772
rect 4075 2746 4094 2772
rect 4158 2768 4220 2780
rect 4232 2768 4307 2780
rect 4365 2768 4440 2780
rect 4452 2768 4483 2780
rect 4489 2768 4524 2780
rect 4158 2766 4320 2768
rect 4053 2738 4094 2746
rect 4176 2742 4189 2766
rect 4204 2764 4219 2766
rect 4016 2728 4017 2738
rect 4032 2728 4045 2738
rect 4059 2728 4060 2738
rect 4075 2728 4088 2738
rect 4103 2728 4133 2742
rect 4176 2728 4219 2742
rect 4243 2739 4250 2746
rect 4253 2742 4320 2766
rect 4352 2766 4524 2768
rect 4322 2744 4350 2748
rect 4352 2744 4432 2766
rect 4453 2764 4468 2766
rect 4322 2742 4432 2744
rect 4253 2738 4432 2742
rect 4226 2728 4256 2738
rect 4258 2728 4411 2738
rect 4419 2728 4449 2738
rect 4453 2728 4483 2742
rect 4511 2728 4524 2766
rect 4596 2772 4631 2780
rect 4596 2746 4597 2772
rect 4604 2746 4631 2772
rect 4539 2728 4569 2742
rect 4596 2738 4631 2746
rect 4633 2772 4674 2780
rect 4633 2746 4648 2772
rect 4655 2746 4674 2772
rect 4738 2768 4800 2780
rect 4812 2768 4887 2780
rect 4945 2768 5020 2780
rect 5032 2768 5063 2780
rect 5069 2768 5104 2780
rect 4738 2766 4900 2768
rect 4633 2738 4674 2746
rect 4756 2742 4769 2766
rect 4784 2764 4799 2766
rect 4596 2728 4597 2738
rect 4612 2728 4625 2738
rect 4639 2728 4640 2738
rect 4655 2728 4668 2738
rect 4683 2728 4713 2742
rect 4756 2728 4799 2742
rect 4823 2739 4830 2746
rect 4833 2742 4900 2766
rect 4932 2766 5104 2768
rect 4902 2744 4930 2748
rect 4932 2744 5012 2766
rect 5033 2764 5048 2766
rect 4902 2742 5012 2744
rect 4833 2738 5012 2742
rect 4806 2728 4836 2738
rect 4838 2728 4991 2738
rect 4999 2728 5029 2738
rect 5033 2728 5063 2742
rect 5091 2728 5104 2766
rect 5176 2772 5211 2780
rect 5176 2746 5177 2772
rect 5184 2746 5211 2772
rect 5119 2728 5149 2742
rect 5176 2738 5211 2746
rect 5213 2772 5254 2780
rect 5213 2746 5228 2772
rect 5235 2746 5254 2772
rect 5318 2768 5380 2780
rect 5392 2768 5467 2780
rect 5525 2768 5600 2780
rect 5612 2768 5643 2780
rect 5649 2768 5684 2780
rect 5318 2766 5480 2768
rect 5213 2738 5254 2746
rect 5336 2742 5349 2766
rect 5364 2764 5379 2766
rect 5176 2728 5177 2738
rect 5192 2728 5205 2738
rect 5219 2728 5220 2738
rect 5235 2728 5248 2738
rect 5263 2728 5293 2742
rect 5336 2728 5379 2742
rect 5403 2739 5410 2746
rect 5413 2742 5480 2766
rect 5512 2766 5684 2768
rect 5482 2744 5510 2748
rect 5512 2744 5592 2766
rect 5613 2764 5628 2766
rect 5482 2742 5592 2744
rect 5413 2738 5592 2742
rect 5386 2728 5416 2738
rect 5418 2728 5571 2738
rect 5579 2728 5609 2738
rect 5613 2728 5643 2742
rect 5671 2728 5684 2766
rect 5756 2772 5791 2780
rect 5756 2746 5757 2772
rect 5764 2746 5791 2772
rect 5699 2728 5729 2742
rect 5756 2738 5791 2746
rect 5793 2772 5834 2780
rect 5793 2746 5808 2772
rect 5815 2746 5834 2772
rect 5898 2768 5960 2780
rect 5972 2768 6047 2780
rect 6105 2768 6180 2780
rect 6192 2768 6223 2780
rect 6229 2768 6264 2780
rect 5898 2766 6060 2768
rect 5793 2738 5834 2746
rect 5916 2742 5929 2766
rect 5944 2764 5959 2766
rect 5756 2728 5757 2738
rect 5772 2728 5785 2738
rect 5799 2728 5800 2738
rect 5815 2728 5828 2738
rect 5843 2728 5873 2742
rect 5916 2728 5959 2742
rect 5983 2739 5990 2746
rect 5993 2742 6060 2766
rect 6092 2766 6264 2768
rect 6062 2744 6090 2748
rect 6092 2744 6172 2766
rect 6193 2764 6208 2766
rect 6062 2742 6172 2744
rect 5993 2738 6172 2742
rect 5966 2728 5996 2738
rect 5998 2728 6151 2738
rect 6159 2728 6189 2738
rect 6193 2728 6223 2742
rect 6251 2728 6264 2766
rect 6336 2772 6371 2780
rect 6336 2746 6337 2772
rect 6344 2746 6371 2772
rect 6279 2728 6309 2742
rect 6336 2738 6371 2746
rect 6373 2772 6414 2780
rect 6373 2746 6388 2772
rect 6395 2746 6414 2772
rect 6478 2768 6540 2780
rect 6552 2768 6627 2780
rect 6685 2768 6760 2780
rect 6772 2768 6803 2780
rect 6809 2768 6844 2780
rect 6478 2766 6640 2768
rect 6373 2738 6414 2746
rect 6496 2742 6509 2766
rect 6524 2764 6539 2766
rect 6336 2728 6337 2738
rect 6352 2728 6365 2738
rect 6379 2728 6380 2738
rect 6395 2728 6408 2738
rect 6423 2728 6453 2742
rect 6496 2728 6539 2742
rect 6563 2739 6570 2746
rect 6573 2742 6640 2766
rect 6672 2766 6844 2768
rect 6642 2744 6670 2748
rect 6672 2744 6752 2766
rect 6773 2764 6788 2766
rect 6642 2742 6752 2744
rect 6573 2738 6752 2742
rect 6546 2728 6576 2738
rect 6578 2728 6731 2738
rect 6739 2728 6769 2738
rect 6773 2728 6803 2742
rect 6831 2728 6844 2766
rect 6916 2772 6951 2780
rect 6916 2746 6917 2772
rect 6924 2746 6951 2772
rect 6859 2728 6889 2742
rect 6916 2738 6951 2746
rect 6953 2772 6994 2780
rect 6953 2746 6968 2772
rect 6975 2746 6994 2772
rect 7058 2768 7120 2780
rect 7132 2768 7207 2780
rect 7265 2768 7340 2780
rect 7352 2768 7383 2780
rect 7389 2768 7424 2780
rect 7058 2766 7220 2768
rect 6953 2738 6994 2746
rect 7076 2742 7089 2766
rect 7104 2764 7119 2766
rect 6916 2728 6917 2738
rect 6932 2728 6945 2738
rect 6959 2728 6960 2738
rect 6975 2728 6988 2738
rect 7003 2728 7033 2742
rect 7076 2728 7119 2742
rect 7143 2739 7150 2746
rect 7153 2742 7220 2766
rect 7252 2766 7424 2768
rect 7222 2744 7250 2748
rect 7252 2744 7332 2766
rect 7353 2764 7368 2766
rect 7222 2742 7332 2744
rect 7153 2738 7332 2742
rect 7126 2728 7156 2738
rect 7158 2728 7311 2738
rect 7319 2728 7349 2738
rect 7353 2728 7383 2742
rect 7411 2728 7424 2766
rect 7496 2772 7531 2780
rect 7496 2746 7497 2772
rect 7504 2746 7531 2772
rect 7439 2728 7469 2742
rect 7496 2738 7531 2746
rect 7533 2772 7574 2780
rect 7533 2746 7548 2772
rect 7555 2746 7574 2772
rect 7638 2768 7700 2780
rect 7712 2768 7787 2780
rect 7845 2768 7920 2780
rect 7932 2768 7963 2780
rect 7969 2768 8004 2780
rect 7638 2766 7800 2768
rect 7533 2738 7574 2746
rect 7656 2742 7669 2766
rect 7684 2764 7699 2766
rect 7496 2728 7497 2738
rect 7512 2728 7525 2738
rect 7539 2728 7540 2738
rect 7555 2728 7568 2738
rect 7583 2728 7613 2742
rect 7656 2728 7699 2742
rect 7723 2739 7730 2746
rect 7733 2742 7800 2766
rect 7832 2766 8004 2768
rect 7802 2744 7830 2748
rect 7832 2744 7912 2766
rect 7933 2764 7948 2766
rect 7802 2742 7912 2744
rect 7733 2738 7912 2742
rect 7706 2728 7736 2738
rect 7738 2728 7891 2738
rect 7899 2728 7929 2738
rect 7933 2728 7963 2742
rect 7991 2728 8004 2766
rect 8076 2772 8111 2780
rect 8076 2746 8077 2772
rect 8084 2746 8111 2772
rect 8019 2728 8049 2742
rect 8076 2738 8111 2746
rect 8113 2772 8154 2780
rect 8113 2746 8128 2772
rect 8135 2746 8154 2772
rect 8218 2768 8280 2780
rect 8292 2768 8367 2780
rect 8425 2768 8500 2780
rect 8512 2768 8543 2780
rect 8549 2768 8584 2780
rect 8218 2766 8380 2768
rect 8113 2738 8154 2746
rect 8236 2742 8249 2766
rect 8264 2764 8279 2766
rect 8076 2728 8077 2738
rect 8092 2728 8105 2738
rect 8119 2728 8120 2738
rect 8135 2728 8148 2738
rect 8163 2728 8193 2742
rect 8236 2728 8279 2742
rect 8303 2739 8310 2746
rect 8313 2742 8380 2766
rect 8412 2766 8584 2768
rect 8382 2744 8410 2748
rect 8412 2744 8492 2766
rect 8513 2764 8528 2766
rect 8382 2742 8492 2744
rect 8313 2738 8492 2742
rect 8286 2728 8316 2738
rect 8318 2728 8471 2738
rect 8479 2728 8509 2738
rect 8513 2728 8543 2742
rect 8571 2728 8584 2766
rect 8656 2772 8691 2780
rect 8656 2746 8657 2772
rect 8664 2746 8691 2772
rect 8599 2728 8629 2742
rect 8656 2738 8691 2746
rect 8693 2772 8734 2780
rect 8693 2746 8708 2772
rect 8715 2746 8734 2772
rect 8798 2768 8860 2780
rect 8872 2768 8947 2780
rect 9005 2768 9080 2780
rect 9092 2768 9123 2780
rect 9129 2768 9164 2780
rect 8798 2766 8960 2768
rect 8693 2738 8734 2746
rect 8816 2742 8829 2766
rect 8844 2764 8859 2766
rect 8656 2728 8657 2738
rect 8672 2728 8685 2738
rect 8699 2728 8700 2738
rect 8715 2728 8728 2738
rect 8743 2728 8773 2742
rect 8816 2728 8859 2742
rect 8883 2739 8890 2746
rect 8893 2742 8960 2766
rect 8992 2766 9164 2768
rect 8962 2744 8990 2748
rect 8992 2744 9072 2766
rect 9093 2764 9108 2766
rect 8962 2742 9072 2744
rect 8893 2738 9072 2742
rect 8866 2728 8896 2738
rect 8898 2728 9051 2738
rect 9059 2728 9089 2738
rect 9093 2728 9123 2742
rect 9151 2728 9164 2766
rect 9236 2772 9271 2780
rect 9236 2746 9237 2772
rect 9244 2746 9271 2772
rect 9179 2728 9209 2742
rect 9236 2738 9271 2746
rect 9236 2728 9237 2738
rect 9252 2728 9265 2738
rect -1 2722 9265 2728
rect 0 2714 9265 2722
rect 15 2684 28 2714
rect 43 2696 73 2714
rect 116 2700 130 2714
rect 166 2700 386 2714
rect 117 2698 130 2700
rect 83 2686 98 2698
rect 80 2684 102 2686
rect 107 2684 137 2698
rect 198 2696 351 2700
rect 180 2684 372 2696
rect 415 2684 445 2698
rect 451 2684 464 2714
rect 479 2696 509 2714
rect 552 2684 565 2714
rect 595 2684 608 2714
rect 623 2696 653 2714
rect 696 2700 710 2714
rect 746 2700 966 2714
rect 697 2698 710 2700
rect 663 2686 678 2698
rect 660 2684 682 2686
rect 687 2684 717 2698
rect 778 2696 931 2700
rect 760 2684 952 2696
rect 995 2684 1025 2698
rect 1031 2684 1044 2714
rect 1059 2696 1089 2714
rect 1132 2684 1145 2714
rect 1175 2684 1188 2714
rect 1203 2696 1233 2714
rect 1276 2700 1290 2714
rect 1326 2700 1546 2714
rect 1277 2698 1290 2700
rect 1243 2686 1258 2698
rect 1240 2684 1262 2686
rect 1267 2684 1297 2698
rect 1358 2696 1511 2700
rect 1340 2684 1532 2696
rect 1575 2684 1605 2698
rect 1611 2684 1624 2714
rect 1639 2696 1669 2714
rect 1712 2684 1725 2714
rect 1755 2684 1768 2714
rect 1783 2696 1813 2714
rect 1856 2700 1870 2714
rect 1906 2700 2126 2714
rect 1857 2698 1870 2700
rect 1823 2686 1838 2698
rect 1820 2684 1842 2686
rect 1847 2684 1877 2698
rect 1938 2696 2091 2700
rect 1920 2684 2112 2696
rect 2155 2684 2185 2698
rect 2191 2684 2204 2714
rect 2219 2696 2249 2714
rect 2292 2684 2305 2714
rect 2335 2684 2348 2714
rect 2363 2696 2393 2714
rect 2436 2700 2450 2714
rect 2486 2700 2706 2714
rect 2437 2698 2450 2700
rect 2403 2686 2418 2698
rect 2400 2684 2422 2686
rect 2427 2684 2457 2698
rect 2518 2696 2671 2700
rect 2500 2684 2692 2696
rect 2735 2684 2765 2698
rect 2771 2684 2784 2714
rect 2799 2696 2829 2714
rect 2872 2684 2885 2714
rect 2915 2684 2928 2714
rect 2943 2696 2973 2714
rect 3016 2700 3030 2714
rect 3066 2700 3286 2714
rect 3017 2698 3030 2700
rect 2983 2686 2998 2698
rect 2980 2684 3002 2686
rect 3007 2684 3037 2698
rect 3098 2696 3251 2700
rect 3080 2684 3272 2696
rect 3315 2684 3345 2698
rect 3351 2684 3364 2714
rect 3379 2696 3409 2714
rect 3452 2684 3465 2714
rect 3495 2684 3508 2714
rect 3523 2696 3553 2714
rect 3596 2700 3610 2714
rect 3646 2700 3866 2714
rect 3597 2698 3610 2700
rect 3563 2686 3578 2698
rect 3560 2684 3582 2686
rect 3587 2684 3617 2698
rect 3678 2696 3831 2700
rect 3660 2684 3852 2696
rect 3895 2684 3925 2698
rect 3931 2684 3944 2714
rect 3959 2696 3989 2714
rect 4032 2684 4045 2714
rect 4075 2684 4088 2714
rect 4103 2696 4133 2714
rect 4176 2700 4190 2714
rect 4226 2700 4446 2714
rect 4177 2698 4190 2700
rect 4143 2686 4158 2698
rect 4140 2684 4162 2686
rect 4167 2684 4197 2698
rect 4258 2696 4411 2700
rect 4240 2684 4432 2696
rect 4475 2684 4505 2698
rect 4511 2684 4524 2714
rect 4539 2696 4569 2714
rect 4612 2684 4625 2714
rect 4655 2684 4668 2714
rect 4683 2696 4713 2714
rect 4756 2700 4770 2714
rect 4806 2700 5026 2714
rect 4757 2698 4770 2700
rect 4723 2686 4738 2698
rect 4720 2684 4742 2686
rect 4747 2684 4777 2698
rect 4838 2696 4991 2700
rect 4820 2684 5012 2696
rect 5055 2684 5085 2698
rect 5091 2684 5104 2714
rect 5119 2696 5149 2714
rect 5192 2684 5205 2714
rect 5235 2684 5248 2714
rect 5263 2696 5293 2714
rect 5336 2700 5350 2714
rect 5386 2700 5606 2714
rect 5337 2698 5350 2700
rect 5303 2686 5318 2698
rect 5300 2684 5322 2686
rect 5327 2684 5357 2698
rect 5418 2696 5571 2700
rect 5400 2684 5592 2696
rect 5635 2684 5665 2698
rect 5671 2684 5684 2714
rect 5699 2696 5729 2714
rect 5772 2684 5785 2714
rect 5815 2684 5828 2714
rect 5843 2696 5873 2714
rect 5916 2700 5930 2714
rect 5966 2700 6186 2714
rect 5917 2698 5930 2700
rect 5883 2686 5898 2698
rect 5880 2684 5902 2686
rect 5907 2684 5937 2698
rect 5998 2696 6151 2700
rect 5980 2684 6172 2696
rect 6215 2684 6245 2698
rect 6251 2684 6264 2714
rect 6279 2696 6309 2714
rect 6352 2684 6365 2714
rect 6395 2684 6408 2714
rect 6423 2696 6453 2714
rect 6496 2700 6510 2714
rect 6546 2700 6766 2714
rect 6497 2698 6510 2700
rect 6463 2686 6478 2698
rect 6460 2684 6482 2686
rect 6487 2684 6517 2698
rect 6578 2696 6731 2700
rect 6560 2684 6752 2696
rect 6795 2684 6825 2698
rect 6831 2684 6844 2714
rect 6859 2696 6889 2714
rect 6932 2684 6945 2714
rect 6975 2684 6988 2714
rect 7003 2696 7033 2714
rect 7076 2700 7090 2714
rect 7126 2700 7346 2714
rect 7077 2698 7090 2700
rect 7043 2686 7058 2698
rect 7040 2684 7062 2686
rect 7067 2684 7097 2698
rect 7158 2696 7311 2700
rect 7140 2684 7332 2696
rect 7375 2684 7405 2698
rect 7411 2684 7424 2714
rect 7439 2696 7469 2714
rect 7512 2684 7525 2714
rect 7555 2684 7568 2714
rect 7583 2696 7613 2714
rect 7656 2700 7670 2714
rect 7706 2700 7926 2714
rect 7657 2698 7670 2700
rect 7623 2686 7638 2698
rect 7620 2684 7642 2686
rect 7647 2684 7677 2698
rect 7738 2696 7891 2700
rect 7720 2684 7912 2696
rect 7955 2684 7985 2698
rect 7991 2684 8004 2714
rect 8019 2696 8049 2714
rect 8092 2684 8105 2714
rect 8135 2684 8148 2714
rect 8163 2696 8193 2714
rect 8236 2700 8250 2714
rect 8286 2700 8506 2714
rect 8237 2698 8250 2700
rect 8203 2686 8218 2698
rect 8200 2684 8222 2686
rect 8227 2684 8257 2698
rect 8318 2696 8471 2700
rect 8300 2684 8492 2696
rect 8535 2684 8565 2698
rect 8571 2684 8584 2714
rect 8599 2696 8629 2714
rect 8672 2684 8685 2714
rect 8715 2684 8728 2714
rect 8743 2696 8773 2714
rect 8816 2700 8830 2714
rect 8866 2700 9086 2714
rect 8817 2698 8830 2700
rect 8783 2686 8798 2698
rect 8780 2684 8802 2686
rect 8807 2684 8837 2698
rect 8898 2696 9051 2700
rect 8880 2684 9072 2696
rect 9115 2684 9145 2698
rect 9151 2684 9164 2714
rect 9179 2696 9209 2714
rect 9252 2684 9265 2714
rect 0 2670 9265 2684
rect 15 2566 28 2670
rect 73 2648 74 2658
rect 89 2648 102 2658
rect 73 2644 102 2648
rect 107 2644 137 2670
rect 155 2656 171 2658
rect 243 2656 296 2670
rect 244 2654 308 2656
rect 351 2654 366 2670
rect 415 2667 445 2670
rect 415 2664 451 2667
rect 381 2656 397 2658
rect 155 2644 170 2648
rect 73 2642 170 2644
rect 198 2642 366 2654
rect 382 2644 397 2648
rect 415 2645 454 2664
rect 473 2658 480 2659
rect 479 2651 480 2658
rect 463 2648 464 2651
rect 479 2648 492 2651
rect 415 2644 445 2645
rect 454 2644 460 2645
rect 463 2644 492 2648
rect 382 2643 492 2644
rect 382 2642 498 2643
rect 57 2634 108 2642
rect 57 2622 82 2634
rect 89 2622 108 2634
rect 139 2634 189 2642
rect 139 2626 155 2634
rect 162 2632 189 2634
rect 198 2632 419 2642
rect 162 2622 419 2632
rect 448 2634 498 2642
rect 448 2625 464 2634
rect 57 2614 108 2622
rect 155 2614 419 2622
rect 445 2622 464 2625
rect 471 2622 498 2634
rect 445 2614 498 2622
rect 73 2606 74 2614
rect 89 2606 102 2614
rect 73 2598 89 2606
rect 70 2591 89 2594
rect 70 2582 92 2591
rect 43 2572 92 2582
rect 43 2566 73 2572
rect 92 2567 97 2572
rect 15 2550 89 2566
rect 107 2558 137 2614
rect 172 2604 380 2614
rect 415 2610 460 2614
rect 463 2613 464 2614
rect 479 2613 492 2614
rect 198 2574 387 2604
rect 213 2571 387 2574
rect 206 2568 387 2571
rect 15 2548 28 2550
rect 43 2548 77 2550
rect 15 2532 89 2548
rect 116 2544 129 2558
rect 144 2544 160 2560
rect 206 2555 217 2568
rect -1 2510 0 2526
rect 15 2510 28 2532
rect 43 2510 73 2532
rect 116 2528 178 2544
rect 206 2537 217 2553
rect 222 2548 232 2568
rect 242 2548 256 2568
rect 259 2555 268 2568
rect 284 2555 293 2568
rect 222 2537 256 2548
rect 259 2537 268 2553
rect 284 2537 293 2553
rect 300 2548 310 2568
rect 320 2548 334 2568
rect 335 2555 346 2568
rect 300 2537 334 2548
rect 335 2537 346 2553
rect 392 2544 408 2560
rect 415 2558 445 2610
rect 479 2606 480 2613
rect 464 2598 480 2606
rect 451 2566 464 2585
rect 479 2566 509 2582
rect 451 2550 525 2566
rect 451 2548 464 2550
rect 479 2548 513 2550
rect 116 2526 129 2528
rect 144 2526 178 2528
rect 116 2510 178 2526
rect 222 2521 238 2524
rect 300 2521 330 2532
rect 378 2528 424 2544
rect 451 2532 525 2548
rect 378 2526 412 2528
rect 377 2510 424 2526
rect 451 2510 464 2532
rect 479 2510 509 2532
rect 536 2510 537 2526
rect 552 2510 565 2670
rect 595 2566 608 2670
rect 653 2648 654 2658
rect 669 2648 682 2658
rect 653 2644 682 2648
rect 687 2644 717 2670
rect 735 2656 751 2658
rect 823 2656 876 2670
rect 824 2654 888 2656
rect 931 2654 946 2670
rect 995 2667 1025 2670
rect 995 2664 1031 2667
rect 961 2656 977 2658
rect 735 2644 750 2648
rect 653 2642 750 2644
rect 778 2642 946 2654
rect 962 2644 977 2648
rect 995 2645 1034 2664
rect 1053 2658 1060 2659
rect 1059 2651 1060 2658
rect 1043 2648 1044 2651
rect 1059 2648 1072 2651
rect 995 2644 1025 2645
rect 1034 2644 1040 2645
rect 1043 2644 1072 2648
rect 962 2643 1072 2644
rect 962 2642 1078 2643
rect 637 2634 688 2642
rect 637 2622 662 2634
rect 669 2622 688 2634
rect 719 2634 769 2642
rect 719 2626 735 2634
rect 742 2632 769 2634
rect 778 2632 999 2642
rect 742 2622 999 2632
rect 1028 2634 1078 2642
rect 1028 2625 1044 2634
rect 637 2614 688 2622
rect 735 2614 999 2622
rect 1025 2622 1044 2625
rect 1051 2622 1078 2634
rect 1025 2614 1078 2622
rect 653 2606 654 2614
rect 669 2606 682 2614
rect 653 2598 669 2606
rect 650 2591 669 2594
rect 650 2582 672 2591
rect 623 2572 672 2582
rect 623 2566 653 2572
rect 672 2567 677 2572
rect 595 2550 669 2566
rect 687 2558 717 2614
rect 752 2604 960 2614
rect 995 2610 1040 2614
rect 1043 2613 1044 2614
rect 1059 2613 1072 2614
rect 778 2574 967 2604
rect 793 2571 967 2574
rect 786 2568 967 2571
rect 595 2548 608 2550
rect 623 2548 657 2550
rect 595 2532 669 2548
rect 696 2544 709 2558
rect 724 2544 740 2560
rect 786 2555 797 2568
rect 579 2510 580 2526
rect 595 2510 608 2532
rect 623 2510 653 2532
rect 696 2528 758 2544
rect 786 2537 797 2553
rect 802 2548 812 2568
rect 822 2548 836 2568
rect 839 2555 848 2568
rect 864 2555 873 2568
rect 802 2537 836 2548
rect 839 2537 848 2553
rect 864 2537 873 2553
rect 880 2548 890 2568
rect 900 2548 914 2568
rect 915 2555 926 2568
rect 880 2537 914 2548
rect 915 2537 926 2553
rect 972 2544 988 2560
rect 995 2558 1025 2610
rect 1059 2606 1060 2613
rect 1044 2598 1060 2606
rect 1031 2566 1044 2585
rect 1059 2566 1089 2582
rect 1031 2550 1105 2566
rect 1031 2548 1044 2550
rect 1059 2548 1093 2550
rect 696 2526 709 2528
rect 724 2526 758 2528
rect 696 2510 758 2526
rect 802 2521 818 2524
rect 880 2521 910 2532
rect 958 2528 1004 2544
rect 1031 2532 1105 2548
rect 958 2526 992 2528
rect 957 2510 1004 2526
rect 1031 2510 1044 2532
rect 1059 2510 1089 2532
rect 1116 2510 1117 2526
rect 1132 2510 1145 2670
rect 1175 2566 1188 2670
rect 1233 2648 1234 2658
rect 1249 2648 1262 2658
rect 1233 2644 1262 2648
rect 1267 2644 1297 2670
rect 1315 2656 1331 2658
rect 1403 2656 1456 2670
rect 1404 2654 1468 2656
rect 1511 2654 1526 2670
rect 1575 2667 1605 2670
rect 1575 2664 1611 2667
rect 1541 2656 1557 2658
rect 1315 2644 1330 2648
rect 1233 2642 1330 2644
rect 1358 2642 1526 2654
rect 1542 2644 1557 2648
rect 1575 2645 1614 2664
rect 1633 2658 1640 2659
rect 1639 2651 1640 2658
rect 1623 2648 1624 2651
rect 1639 2648 1652 2651
rect 1575 2644 1605 2645
rect 1614 2644 1620 2645
rect 1623 2644 1652 2648
rect 1542 2643 1652 2644
rect 1542 2642 1658 2643
rect 1217 2634 1268 2642
rect 1217 2622 1242 2634
rect 1249 2622 1268 2634
rect 1299 2634 1349 2642
rect 1299 2626 1315 2634
rect 1322 2632 1349 2634
rect 1358 2632 1579 2642
rect 1322 2622 1579 2632
rect 1608 2634 1658 2642
rect 1608 2625 1624 2634
rect 1217 2614 1268 2622
rect 1315 2614 1579 2622
rect 1605 2622 1624 2625
rect 1631 2622 1658 2634
rect 1605 2614 1658 2622
rect 1233 2606 1234 2614
rect 1249 2606 1262 2614
rect 1233 2598 1249 2606
rect 1230 2591 1249 2594
rect 1230 2582 1252 2591
rect 1203 2572 1252 2582
rect 1203 2566 1233 2572
rect 1252 2567 1257 2572
rect 1175 2550 1249 2566
rect 1267 2558 1297 2614
rect 1332 2604 1540 2614
rect 1575 2610 1620 2614
rect 1623 2613 1624 2614
rect 1639 2613 1652 2614
rect 1358 2574 1547 2604
rect 1373 2571 1547 2574
rect 1366 2568 1547 2571
rect 1175 2548 1188 2550
rect 1203 2548 1237 2550
rect 1175 2532 1249 2548
rect 1276 2544 1289 2558
rect 1304 2544 1320 2560
rect 1366 2555 1377 2568
rect 1159 2510 1160 2526
rect 1175 2510 1188 2532
rect 1203 2510 1233 2532
rect 1276 2528 1338 2544
rect 1366 2537 1377 2553
rect 1382 2548 1392 2568
rect 1402 2548 1416 2568
rect 1419 2555 1428 2568
rect 1444 2555 1453 2568
rect 1382 2537 1416 2548
rect 1419 2537 1428 2553
rect 1444 2537 1453 2553
rect 1460 2548 1470 2568
rect 1480 2548 1494 2568
rect 1495 2555 1506 2568
rect 1460 2537 1494 2548
rect 1495 2537 1506 2553
rect 1552 2544 1568 2560
rect 1575 2558 1605 2610
rect 1639 2606 1640 2613
rect 1624 2598 1640 2606
rect 1611 2566 1624 2585
rect 1639 2566 1669 2582
rect 1611 2550 1685 2566
rect 1611 2548 1624 2550
rect 1639 2548 1673 2550
rect 1276 2526 1289 2528
rect 1304 2526 1338 2528
rect 1276 2510 1338 2526
rect 1382 2521 1398 2524
rect 1460 2521 1490 2532
rect 1538 2528 1584 2544
rect 1611 2532 1685 2548
rect 1538 2526 1572 2528
rect 1537 2510 1584 2526
rect 1611 2510 1624 2532
rect 1639 2510 1669 2532
rect 1696 2510 1697 2526
rect 1712 2510 1725 2670
rect 1755 2566 1768 2670
rect 1813 2648 1814 2658
rect 1829 2648 1842 2658
rect 1813 2644 1842 2648
rect 1847 2644 1877 2670
rect 1895 2656 1911 2658
rect 1983 2656 2036 2670
rect 1984 2654 2048 2656
rect 2091 2654 2106 2670
rect 2155 2667 2185 2670
rect 2155 2664 2191 2667
rect 2121 2656 2137 2658
rect 1895 2644 1910 2648
rect 1813 2642 1910 2644
rect 1938 2642 2106 2654
rect 2122 2644 2137 2648
rect 2155 2645 2194 2664
rect 2213 2658 2220 2659
rect 2219 2651 2220 2658
rect 2203 2648 2204 2651
rect 2219 2648 2232 2651
rect 2155 2644 2185 2645
rect 2194 2644 2200 2645
rect 2203 2644 2232 2648
rect 2122 2643 2232 2644
rect 2122 2642 2238 2643
rect 1797 2634 1848 2642
rect 1797 2622 1822 2634
rect 1829 2622 1848 2634
rect 1879 2634 1929 2642
rect 1879 2626 1895 2634
rect 1902 2632 1929 2634
rect 1938 2632 2159 2642
rect 1902 2622 2159 2632
rect 2188 2634 2238 2642
rect 2188 2625 2204 2634
rect 1797 2614 1848 2622
rect 1895 2614 2159 2622
rect 2185 2622 2204 2625
rect 2211 2622 2238 2634
rect 2185 2614 2238 2622
rect 1813 2606 1814 2614
rect 1829 2606 1842 2614
rect 1813 2598 1829 2606
rect 1810 2591 1829 2594
rect 1810 2582 1832 2591
rect 1783 2572 1832 2582
rect 1783 2566 1813 2572
rect 1832 2567 1837 2572
rect 1755 2550 1829 2566
rect 1847 2558 1877 2614
rect 1912 2604 2120 2614
rect 2155 2610 2200 2614
rect 2203 2613 2204 2614
rect 2219 2613 2232 2614
rect 1938 2574 2127 2604
rect 1953 2571 2127 2574
rect 1946 2568 2127 2571
rect 1755 2548 1768 2550
rect 1783 2548 1817 2550
rect 1755 2532 1829 2548
rect 1856 2544 1869 2558
rect 1884 2544 1900 2560
rect 1946 2555 1957 2568
rect 1739 2510 1740 2526
rect 1755 2510 1768 2532
rect 1783 2510 1813 2532
rect 1856 2528 1918 2544
rect 1946 2537 1957 2553
rect 1962 2548 1972 2568
rect 1982 2548 1996 2568
rect 1999 2555 2008 2568
rect 2024 2555 2033 2568
rect 1962 2537 1996 2548
rect 1999 2537 2008 2553
rect 2024 2537 2033 2553
rect 2040 2548 2050 2568
rect 2060 2548 2074 2568
rect 2075 2555 2086 2568
rect 2040 2537 2074 2548
rect 2075 2537 2086 2553
rect 2132 2544 2148 2560
rect 2155 2558 2185 2610
rect 2219 2606 2220 2613
rect 2204 2598 2220 2606
rect 2191 2566 2204 2585
rect 2219 2566 2249 2582
rect 2191 2550 2265 2566
rect 2191 2548 2204 2550
rect 2219 2548 2253 2550
rect 1856 2526 1869 2528
rect 1884 2526 1918 2528
rect 1856 2510 1918 2526
rect 1962 2521 1976 2524
rect 2040 2521 2070 2532
rect 2118 2528 2164 2544
rect 2191 2532 2265 2548
rect 2118 2526 2152 2528
rect 2117 2510 2164 2526
rect 2191 2510 2204 2532
rect 2219 2510 2249 2532
rect 2276 2510 2277 2526
rect 2292 2510 2305 2670
rect 2335 2566 2348 2670
rect 2393 2648 2394 2658
rect 2409 2648 2422 2658
rect 2393 2644 2422 2648
rect 2427 2644 2457 2670
rect 2475 2656 2491 2658
rect 2563 2656 2616 2670
rect 2564 2654 2628 2656
rect 2671 2654 2686 2670
rect 2735 2667 2765 2670
rect 2735 2664 2771 2667
rect 2701 2656 2717 2658
rect 2475 2644 2490 2648
rect 2393 2642 2490 2644
rect 2518 2642 2686 2654
rect 2702 2644 2717 2648
rect 2735 2645 2774 2664
rect 2793 2658 2800 2659
rect 2799 2651 2800 2658
rect 2783 2648 2784 2651
rect 2799 2648 2812 2651
rect 2735 2644 2765 2645
rect 2774 2644 2780 2645
rect 2783 2644 2812 2648
rect 2702 2643 2812 2644
rect 2702 2642 2818 2643
rect 2377 2634 2428 2642
rect 2377 2622 2402 2634
rect 2409 2622 2428 2634
rect 2459 2634 2509 2642
rect 2459 2626 2475 2634
rect 2482 2632 2509 2634
rect 2518 2632 2739 2642
rect 2482 2622 2739 2632
rect 2768 2634 2818 2642
rect 2768 2625 2784 2634
rect 2377 2614 2428 2622
rect 2475 2614 2739 2622
rect 2765 2622 2784 2625
rect 2791 2622 2818 2634
rect 2765 2614 2818 2622
rect 2393 2606 2394 2614
rect 2409 2606 2422 2614
rect 2393 2598 2409 2606
rect 2390 2591 2409 2594
rect 2390 2582 2412 2591
rect 2363 2572 2412 2582
rect 2363 2566 2393 2572
rect 2412 2567 2417 2572
rect 2335 2550 2409 2566
rect 2427 2558 2457 2614
rect 2492 2604 2700 2614
rect 2735 2610 2780 2614
rect 2783 2613 2784 2614
rect 2799 2613 2812 2614
rect 2518 2574 2707 2604
rect 2533 2571 2707 2574
rect 2526 2568 2707 2571
rect 2335 2548 2348 2550
rect 2363 2548 2397 2550
rect 2335 2532 2409 2548
rect 2436 2544 2449 2558
rect 2464 2544 2480 2560
rect 2526 2555 2537 2568
rect 2319 2510 2320 2526
rect 2335 2510 2348 2532
rect 2363 2510 2393 2532
rect 2436 2528 2498 2544
rect 2526 2537 2537 2553
rect 2542 2548 2552 2568
rect 2562 2548 2576 2568
rect 2579 2555 2588 2568
rect 2604 2555 2613 2568
rect 2542 2537 2576 2548
rect 2579 2537 2588 2553
rect 2604 2537 2613 2553
rect 2620 2548 2630 2568
rect 2640 2548 2654 2568
rect 2655 2555 2666 2568
rect 2620 2537 2654 2548
rect 2655 2537 2666 2553
rect 2712 2544 2728 2560
rect 2735 2558 2765 2610
rect 2799 2606 2800 2613
rect 2784 2598 2800 2606
rect 2771 2566 2784 2585
rect 2799 2566 2829 2582
rect 2771 2550 2845 2566
rect 2771 2548 2784 2550
rect 2799 2548 2833 2550
rect 2436 2526 2449 2528
rect 2464 2526 2498 2528
rect 2436 2510 2498 2526
rect 2542 2521 2558 2524
rect 2620 2521 2650 2532
rect 2698 2528 2744 2544
rect 2771 2532 2845 2548
rect 2698 2526 2732 2528
rect 2697 2510 2744 2526
rect 2771 2510 2784 2532
rect 2799 2510 2829 2532
rect 2856 2510 2857 2526
rect 2872 2510 2885 2670
rect 2915 2566 2928 2670
rect 2973 2648 2974 2658
rect 2989 2648 3002 2658
rect 2973 2644 3002 2648
rect 3007 2644 3037 2670
rect 3055 2656 3071 2658
rect 3143 2656 3196 2670
rect 3144 2654 3208 2656
rect 3251 2654 3266 2670
rect 3315 2667 3345 2670
rect 3315 2664 3351 2667
rect 3281 2656 3297 2658
rect 3055 2644 3070 2648
rect 2973 2642 3070 2644
rect 3098 2642 3266 2654
rect 3282 2644 3297 2648
rect 3315 2645 3354 2664
rect 3373 2658 3380 2659
rect 3379 2651 3380 2658
rect 3363 2648 3364 2651
rect 3379 2648 3392 2651
rect 3315 2644 3345 2645
rect 3354 2644 3360 2645
rect 3363 2644 3392 2648
rect 3282 2643 3392 2644
rect 3282 2642 3398 2643
rect 2957 2634 3008 2642
rect 2957 2622 2982 2634
rect 2989 2622 3008 2634
rect 3039 2634 3089 2642
rect 3039 2626 3055 2634
rect 3062 2632 3089 2634
rect 3098 2632 3319 2642
rect 3062 2622 3319 2632
rect 3348 2634 3398 2642
rect 3348 2625 3364 2634
rect 2957 2614 3008 2622
rect 3055 2614 3319 2622
rect 3345 2622 3364 2625
rect 3371 2622 3398 2634
rect 3345 2614 3398 2622
rect 2973 2606 2974 2614
rect 2989 2606 3002 2614
rect 2973 2598 2989 2606
rect 2970 2591 2989 2594
rect 2970 2582 2992 2591
rect 2943 2572 2992 2582
rect 2943 2566 2973 2572
rect 2992 2567 2997 2572
rect 2915 2550 2989 2566
rect 3007 2558 3037 2614
rect 3072 2604 3280 2614
rect 3315 2610 3360 2614
rect 3363 2613 3364 2614
rect 3379 2613 3392 2614
rect 3098 2574 3287 2604
rect 3113 2571 3287 2574
rect 3106 2568 3287 2571
rect 2915 2548 2928 2550
rect 2943 2548 2977 2550
rect 2915 2532 2989 2548
rect 3016 2544 3029 2558
rect 3044 2544 3060 2560
rect 3106 2555 3117 2568
rect 2899 2510 2900 2526
rect 2915 2510 2928 2532
rect 2943 2510 2973 2532
rect 3016 2528 3078 2544
rect 3106 2537 3117 2553
rect 3122 2548 3132 2568
rect 3142 2548 3156 2568
rect 3159 2555 3168 2568
rect 3184 2555 3193 2568
rect 3122 2537 3156 2548
rect 3159 2537 3168 2553
rect 3184 2537 3193 2553
rect 3200 2548 3210 2568
rect 3220 2548 3234 2568
rect 3235 2555 3246 2568
rect 3200 2537 3234 2548
rect 3235 2537 3246 2553
rect 3292 2544 3308 2560
rect 3315 2558 3345 2610
rect 3379 2606 3380 2613
rect 3364 2598 3380 2606
rect 3351 2566 3364 2585
rect 3379 2566 3409 2582
rect 3351 2550 3425 2566
rect 3351 2548 3364 2550
rect 3379 2548 3413 2550
rect 3016 2526 3029 2528
rect 3044 2526 3078 2528
rect 3016 2510 3078 2526
rect 3122 2521 3138 2524
rect 3200 2521 3230 2532
rect 3278 2528 3324 2544
rect 3351 2532 3425 2548
rect 3278 2526 3312 2528
rect 3277 2510 3324 2526
rect 3351 2510 3364 2532
rect 3379 2510 3409 2532
rect 3436 2510 3437 2526
rect 3452 2510 3465 2670
rect 3495 2566 3508 2670
rect 3553 2648 3554 2658
rect 3569 2648 3582 2658
rect 3553 2644 3582 2648
rect 3587 2644 3617 2670
rect 3635 2656 3651 2658
rect 3723 2656 3776 2670
rect 3724 2654 3788 2656
rect 3831 2654 3846 2670
rect 3895 2667 3925 2670
rect 3895 2664 3931 2667
rect 3861 2656 3877 2658
rect 3635 2644 3650 2648
rect 3553 2642 3650 2644
rect 3678 2642 3846 2654
rect 3862 2644 3877 2648
rect 3895 2645 3934 2664
rect 3953 2658 3960 2659
rect 3959 2651 3960 2658
rect 3943 2648 3944 2651
rect 3959 2648 3972 2651
rect 3895 2644 3925 2645
rect 3934 2644 3940 2645
rect 3943 2644 3972 2648
rect 3862 2643 3972 2644
rect 3862 2642 3978 2643
rect 3537 2634 3588 2642
rect 3537 2622 3562 2634
rect 3569 2622 3588 2634
rect 3619 2634 3669 2642
rect 3619 2626 3635 2634
rect 3642 2632 3669 2634
rect 3678 2632 3899 2642
rect 3642 2622 3899 2632
rect 3928 2634 3978 2642
rect 3928 2625 3944 2634
rect 3537 2614 3588 2622
rect 3635 2614 3899 2622
rect 3925 2622 3944 2625
rect 3951 2622 3978 2634
rect 3925 2614 3978 2622
rect 3553 2606 3554 2614
rect 3569 2606 3582 2614
rect 3553 2598 3569 2606
rect 3550 2591 3569 2594
rect 3550 2582 3572 2591
rect 3523 2572 3572 2582
rect 3523 2566 3553 2572
rect 3572 2567 3577 2572
rect 3495 2550 3569 2566
rect 3587 2558 3617 2614
rect 3652 2604 3860 2614
rect 3895 2610 3940 2614
rect 3943 2613 3944 2614
rect 3959 2613 3972 2614
rect 3678 2574 3867 2604
rect 3693 2571 3867 2574
rect 3686 2568 3867 2571
rect 3495 2548 3508 2550
rect 3523 2548 3557 2550
rect 3495 2532 3569 2548
rect 3596 2544 3609 2558
rect 3624 2544 3640 2560
rect 3686 2555 3697 2568
rect 3479 2510 3480 2526
rect 3495 2510 3508 2532
rect 3523 2510 3553 2532
rect 3596 2528 3658 2544
rect 3686 2537 3697 2553
rect 3702 2548 3712 2568
rect 3722 2548 3736 2568
rect 3739 2555 3748 2568
rect 3764 2555 3773 2568
rect 3702 2537 3736 2548
rect 3739 2537 3748 2553
rect 3764 2537 3773 2553
rect 3780 2548 3790 2568
rect 3800 2548 3814 2568
rect 3815 2555 3826 2568
rect 3780 2537 3814 2548
rect 3815 2537 3826 2553
rect 3872 2544 3888 2560
rect 3895 2558 3925 2610
rect 3959 2606 3960 2613
rect 3944 2598 3960 2606
rect 3931 2566 3944 2585
rect 3959 2566 3989 2582
rect 3931 2550 4005 2566
rect 3931 2548 3944 2550
rect 3959 2548 3993 2550
rect 3596 2526 3609 2528
rect 3624 2526 3658 2528
rect 3596 2510 3658 2526
rect 3702 2521 3718 2524
rect 3780 2521 3810 2532
rect 3858 2528 3904 2544
rect 3931 2532 4005 2548
rect 3858 2526 3892 2528
rect 3857 2510 3904 2526
rect 3931 2510 3944 2532
rect 3959 2510 3989 2532
rect 4016 2510 4017 2526
rect 4032 2510 4045 2670
rect 4075 2566 4088 2670
rect 4133 2648 4134 2658
rect 4149 2648 4162 2658
rect 4133 2644 4162 2648
rect 4167 2644 4197 2670
rect 4215 2656 4231 2658
rect 4303 2656 4356 2670
rect 4304 2654 4368 2656
rect 4411 2654 4426 2670
rect 4475 2667 4505 2670
rect 4475 2664 4511 2667
rect 4441 2656 4457 2658
rect 4215 2644 4230 2648
rect 4133 2642 4230 2644
rect 4258 2642 4426 2654
rect 4442 2644 4457 2648
rect 4475 2645 4514 2664
rect 4533 2658 4540 2659
rect 4539 2651 4540 2658
rect 4523 2648 4524 2651
rect 4539 2648 4552 2651
rect 4475 2644 4505 2645
rect 4514 2644 4520 2645
rect 4523 2644 4552 2648
rect 4442 2643 4552 2644
rect 4442 2642 4558 2643
rect 4117 2634 4168 2642
rect 4117 2622 4142 2634
rect 4149 2622 4168 2634
rect 4199 2634 4249 2642
rect 4199 2626 4215 2634
rect 4222 2632 4249 2634
rect 4258 2632 4479 2642
rect 4222 2622 4479 2632
rect 4508 2634 4558 2642
rect 4508 2625 4524 2634
rect 4117 2614 4168 2622
rect 4215 2614 4479 2622
rect 4505 2622 4524 2625
rect 4531 2622 4558 2634
rect 4505 2614 4558 2622
rect 4133 2606 4134 2614
rect 4149 2606 4162 2614
rect 4133 2598 4149 2606
rect 4130 2591 4149 2594
rect 4130 2582 4152 2591
rect 4103 2572 4152 2582
rect 4103 2566 4133 2572
rect 4152 2567 4157 2572
rect 4075 2550 4149 2566
rect 4167 2558 4197 2614
rect 4232 2604 4440 2614
rect 4475 2610 4520 2614
rect 4523 2613 4524 2614
rect 4539 2613 4552 2614
rect 4258 2574 4447 2604
rect 4273 2571 4447 2574
rect 4266 2568 4447 2571
rect 4075 2548 4088 2550
rect 4103 2548 4137 2550
rect 4075 2532 4149 2548
rect 4176 2544 4189 2558
rect 4204 2544 4220 2560
rect 4266 2555 4277 2568
rect 4059 2510 4060 2526
rect 4075 2510 4088 2532
rect 4103 2510 4133 2532
rect 4176 2528 4238 2544
rect 4266 2537 4277 2553
rect 4282 2548 4292 2568
rect 4302 2548 4316 2568
rect 4319 2555 4328 2568
rect 4344 2555 4353 2568
rect 4282 2537 4316 2548
rect 4319 2537 4328 2553
rect 4344 2537 4353 2553
rect 4360 2548 4370 2568
rect 4380 2548 4394 2568
rect 4395 2555 4406 2568
rect 4360 2537 4394 2548
rect 4395 2537 4406 2553
rect 4452 2544 4468 2560
rect 4475 2558 4505 2610
rect 4539 2606 4540 2613
rect 4524 2598 4540 2606
rect 4511 2566 4524 2585
rect 4539 2566 4569 2582
rect 4511 2550 4585 2566
rect 4511 2548 4524 2550
rect 4539 2548 4573 2550
rect 4176 2526 4189 2528
rect 4204 2526 4238 2528
rect 4176 2510 4238 2526
rect 4282 2521 4298 2524
rect 4360 2521 4390 2532
rect 4438 2528 4484 2544
rect 4511 2532 4585 2548
rect 4438 2526 4472 2528
rect 4437 2510 4484 2526
rect 4511 2510 4524 2532
rect 4539 2510 4569 2532
rect 4596 2510 4597 2526
rect 4612 2510 4625 2670
rect 4655 2566 4668 2670
rect 4713 2648 4714 2658
rect 4729 2648 4742 2658
rect 4713 2644 4742 2648
rect 4747 2644 4777 2670
rect 4795 2656 4811 2658
rect 4883 2656 4936 2670
rect 4884 2654 4948 2656
rect 4991 2654 5006 2670
rect 5055 2667 5085 2670
rect 5055 2664 5091 2667
rect 5021 2656 5037 2658
rect 4795 2644 4810 2648
rect 4713 2642 4810 2644
rect 4838 2642 5006 2654
rect 5022 2644 5037 2648
rect 5055 2645 5094 2664
rect 5113 2658 5120 2659
rect 5119 2651 5120 2658
rect 5103 2648 5104 2651
rect 5119 2648 5132 2651
rect 5055 2644 5085 2645
rect 5094 2644 5100 2645
rect 5103 2644 5132 2648
rect 5022 2643 5132 2644
rect 5022 2642 5138 2643
rect 4697 2634 4748 2642
rect 4697 2622 4722 2634
rect 4729 2622 4748 2634
rect 4779 2634 4829 2642
rect 4779 2626 4795 2634
rect 4802 2632 4829 2634
rect 4838 2632 5059 2642
rect 4802 2622 5059 2632
rect 5088 2634 5138 2642
rect 5088 2625 5104 2634
rect 4697 2614 4748 2622
rect 4795 2614 5059 2622
rect 5085 2622 5104 2625
rect 5111 2622 5138 2634
rect 5085 2614 5138 2622
rect 4713 2606 4714 2614
rect 4729 2606 4742 2614
rect 4713 2598 4729 2606
rect 4710 2591 4729 2594
rect 4710 2582 4732 2591
rect 4683 2572 4732 2582
rect 4683 2566 4713 2572
rect 4732 2567 4737 2572
rect 4655 2550 4729 2566
rect 4747 2558 4777 2614
rect 4812 2604 5020 2614
rect 5055 2610 5100 2614
rect 5103 2613 5104 2614
rect 5119 2613 5132 2614
rect 4838 2574 5027 2604
rect 4853 2571 5027 2574
rect 4846 2568 5027 2571
rect 4655 2548 4668 2550
rect 4683 2548 4717 2550
rect 4655 2532 4729 2548
rect 4756 2544 4769 2558
rect 4784 2544 4800 2560
rect 4846 2555 4857 2568
rect 4639 2510 4640 2526
rect 4655 2510 4668 2532
rect 4683 2510 4713 2532
rect 4756 2528 4818 2544
rect 4846 2537 4857 2553
rect 4862 2548 4872 2568
rect 4882 2548 4896 2568
rect 4899 2555 4908 2568
rect 4924 2555 4933 2568
rect 4862 2537 4896 2548
rect 4899 2537 4908 2553
rect 4924 2537 4933 2553
rect 4940 2548 4950 2568
rect 4960 2548 4974 2568
rect 4975 2555 4986 2568
rect 4940 2537 4974 2548
rect 4975 2537 4986 2553
rect 5032 2544 5048 2560
rect 5055 2558 5085 2610
rect 5119 2606 5120 2613
rect 5104 2598 5120 2606
rect 5091 2566 5104 2585
rect 5119 2566 5149 2582
rect 5091 2550 5165 2566
rect 5091 2548 5104 2550
rect 5119 2548 5153 2550
rect 4756 2526 4769 2528
rect 4784 2526 4818 2528
rect 4756 2510 4818 2526
rect 4862 2521 4878 2524
rect 4940 2521 4970 2532
rect 5018 2528 5064 2544
rect 5091 2532 5165 2548
rect 5018 2526 5052 2528
rect 5017 2510 5064 2526
rect 5091 2510 5104 2532
rect 5119 2510 5149 2532
rect 5176 2510 5177 2526
rect 5192 2510 5205 2670
rect 5235 2566 5248 2670
rect 5293 2648 5294 2658
rect 5309 2648 5322 2658
rect 5293 2644 5322 2648
rect 5327 2644 5357 2670
rect 5375 2656 5391 2658
rect 5463 2656 5516 2670
rect 5464 2654 5528 2656
rect 5571 2654 5586 2670
rect 5635 2667 5665 2670
rect 5635 2664 5671 2667
rect 5601 2656 5617 2658
rect 5375 2644 5390 2648
rect 5293 2642 5390 2644
rect 5418 2642 5586 2654
rect 5602 2644 5617 2648
rect 5635 2645 5674 2664
rect 5693 2658 5700 2659
rect 5699 2651 5700 2658
rect 5683 2648 5684 2651
rect 5699 2648 5712 2651
rect 5635 2644 5665 2645
rect 5674 2644 5680 2645
rect 5683 2644 5712 2648
rect 5602 2643 5712 2644
rect 5602 2642 5718 2643
rect 5277 2634 5328 2642
rect 5277 2622 5302 2634
rect 5309 2622 5328 2634
rect 5359 2634 5409 2642
rect 5359 2626 5375 2634
rect 5382 2632 5409 2634
rect 5418 2632 5639 2642
rect 5382 2622 5639 2632
rect 5668 2634 5718 2642
rect 5668 2625 5684 2634
rect 5277 2614 5328 2622
rect 5375 2614 5639 2622
rect 5665 2622 5684 2625
rect 5691 2622 5718 2634
rect 5665 2614 5718 2622
rect 5293 2606 5294 2614
rect 5309 2606 5322 2614
rect 5293 2598 5309 2606
rect 5290 2591 5309 2594
rect 5290 2582 5312 2591
rect 5263 2572 5312 2582
rect 5263 2566 5293 2572
rect 5312 2567 5317 2572
rect 5235 2550 5309 2566
rect 5327 2558 5357 2614
rect 5392 2604 5600 2614
rect 5635 2610 5680 2614
rect 5683 2613 5684 2614
rect 5699 2613 5712 2614
rect 5418 2574 5607 2604
rect 5433 2571 5607 2574
rect 5426 2568 5607 2571
rect 5235 2548 5248 2550
rect 5263 2548 5297 2550
rect 5235 2532 5309 2548
rect 5336 2544 5349 2558
rect 5364 2544 5380 2560
rect 5426 2555 5437 2568
rect 5219 2510 5220 2526
rect 5235 2510 5248 2532
rect 5263 2510 5293 2532
rect 5336 2528 5398 2544
rect 5426 2537 5437 2553
rect 5442 2548 5452 2568
rect 5462 2548 5476 2568
rect 5479 2555 5488 2568
rect 5504 2555 5513 2568
rect 5442 2537 5476 2548
rect 5479 2537 5488 2553
rect 5504 2537 5513 2553
rect 5520 2548 5530 2568
rect 5540 2548 5554 2568
rect 5555 2555 5566 2568
rect 5520 2537 5554 2548
rect 5555 2537 5566 2553
rect 5612 2544 5628 2560
rect 5635 2558 5665 2610
rect 5699 2606 5700 2613
rect 5684 2598 5700 2606
rect 5671 2566 5684 2585
rect 5699 2566 5729 2582
rect 5671 2550 5745 2566
rect 5671 2548 5684 2550
rect 5699 2548 5733 2550
rect 5336 2526 5349 2528
rect 5364 2526 5398 2528
rect 5336 2510 5398 2526
rect 5442 2521 5458 2524
rect 5520 2521 5550 2532
rect 5598 2528 5644 2544
rect 5671 2532 5745 2548
rect 5598 2526 5632 2528
rect 5597 2510 5644 2526
rect 5671 2510 5684 2532
rect 5699 2510 5729 2532
rect 5756 2510 5757 2526
rect 5772 2510 5785 2670
rect 5815 2566 5828 2670
rect 5873 2648 5874 2658
rect 5889 2648 5902 2658
rect 5873 2644 5902 2648
rect 5907 2644 5937 2670
rect 5955 2656 5971 2658
rect 6043 2656 6096 2670
rect 6044 2654 6108 2656
rect 6151 2654 6166 2670
rect 6215 2667 6245 2670
rect 6215 2664 6251 2667
rect 6181 2656 6197 2658
rect 5955 2644 5970 2648
rect 5873 2642 5970 2644
rect 5998 2642 6166 2654
rect 6182 2644 6197 2648
rect 6215 2645 6254 2664
rect 6273 2658 6280 2659
rect 6279 2651 6280 2658
rect 6263 2648 6264 2651
rect 6279 2648 6292 2651
rect 6215 2644 6245 2645
rect 6254 2644 6260 2645
rect 6263 2644 6292 2648
rect 6182 2643 6292 2644
rect 6182 2642 6298 2643
rect 5857 2634 5908 2642
rect 5857 2622 5882 2634
rect 5889 2622 5908 2634
rect 5939 2634 5989 2642
rect 5939 2626 5955 2634
rect 5962 2632 5989 2634
rect 5998 2632 6219 2642
rect 5962 2622 6219 2632
rect 6248 2634 6298 2642
rect 6248 2625 6264 2634
rect 5857 2614 5908 2622
rect 5955 2614 6219 2622
rect 6245 2622 6264 2625
rect 6271 2622 6298 2634
rect 6245 2614 6298 2622
rect 5873 2606 5874 2614
rect 5889 2606 5902 2614
rect 5873 2598 5889 2606
rect 5870 2591 5889 2594
rect 5870 2582 5892 2591
rect 5843 2572 5892 2582
rect 5843 2566 5873 2572
rect 5892 2567 5897 2572
rect 5815 2550 5889 2566
rect 5907 2558 5937 2614
rect 5972 2604 6180 2614
rect 6215 2610 6260 2614
rect 6263 2613 6264 2614
rect 6279 2613 6292 2614
rect 5998 2574 6187 2604
rect 6013 2571 6187 2574
rect 6006 2568 6187 2571
rect 5815 2548 5828 2550
rect 5843 2548 5877 2550
rect 5815 2532 5889 2548
rect 5916 2544 5929 2558
rect 5944 2544 5960 2560
rect 6006 2555 6017 2568
rect 5799 2510 5800 2526
rect 5815 2510 5828 2532
rect 5843 2510 5873 2532
rect 5916 2528 5978 2544
rect 6006 2537 6017 2553
rect 6022 2548 6032 2568
rect 6042 2548 6056 2568
rect 6059 2555 6068 2568
rect 6084 2555 6093 2568
rect 6022 2537 6056 2548
rect 6059 2537 6068 2553
rect 6084 2537 6093 2553
rect 6100 2548 6110 2568
rect 6120 2548 6134 2568
rect 6135 2555 6146 2568
rect 6100 2537 6134 2548
rect 6135 2537 6146 2553
rect 6192 2544 6208 2560
rect 6215 2558 6245 2610
rect 6279 2606 6280 2613
rect 6264 2598 6280 2606
rect 6251 2566 6264 2585
rect 6279 2566 6309 2582
rect 6251 2550 6325 2566
rect 6251 2548 6264 2550
rect 6279 2548 6313 2550
rect 5916 2526 5929 2528
rect 5944 2526 5978 2528
rect 5916 2510 5978 2526
rect 6022 2521 6038 2524
rect 6100 2521 6130 2532
rect 6178 2528 6224 2544
rect 6251 2532 6325 2548
rect 6178 2526 6212 2528
rect 6177 2510 6224 2526
rect 6251 2510 6264 2532
rect 6279 2510 6309 2532
rect 6336 2510 6337 2526
rect 6352 2510 6365 2670
rect 6395 2566 6408 2670
rect 6453 2648 6454 2658
rect 6469 2648 6482 2658
rect 6453 2644 6482 2648
rect 6487 2644 6517 2670
rect 6535 2656 6551 2658
rect 6623 2656 6676 2670
rect 6624 2654 6688 2656
rect 6731 2654 6746 2670
rect 6795 2667 6825 2670
rect 6795 2664 6831 2667
rect 6761 2656 6777 2658
rect 6535 2644 6550 2648
rect 6453 2642 6550 2644
rect 6578 2642 6746 2654
rect 6762 2644 6777 2648
rect 6795 2645 6834 2664
rect 6853 2658 6860 2659
rect 6859 2651 6860 2658
rect 6843 2648 6844 2651
rect 6859 2648 6872 2651
rect 6795 2644 6825 2645
rect 6834 2644 6840 2645
rect 6843 2644 6872 2648
rect 6762 2643 6872 2644
rect 6762 2642 6878 2643
rect 6437 2634 6488 2642
rect 6437 2622 6462 2634
rect 6469 2622 6488 2634
rect 6519 2634 6569 2642
rect 6519 2626 6535 2634
rect 6542 2632 6569 2634
rect 6578 2632 6799 2642
rect 6542 2622 6799 2632
rect 6828 2634 6878 2642
rect 6828 2625 6844 2634
rect 6437 2614 6488 2622
rect 6535 2614 6799 2622
rect 6825 2622 6844 2625
rect 6851 2622 6878 2634
rect 6825 2614 6878 2622
rect 6453 2606 6454 2614
rect 6469 2606 6482 2614
rect 6453 2598 6469 2606
rect 6450 2591 6469 2594
rect 6450 2582 6472 2591
rect 6423 2572 6472 2582
rect 6423 2566 6453 2572
rect 6472 2567 6477 2572
rect 6395 2550 6469 2566
rect 6487 2558 6517 2614
rect 6552 2604 6760 2614
rect 6795 2610 6840 2614
rect 6843 2613 6844 2614
rect 6859 2613 6872 2614
rect 6578 2574 6767 2604
rect 6593 2571 6767 2574
rect 6586 2568 6767 2571
rect 6395 2548 6408 2550
rect 6423 2548 6457 2550
rect 6395 2532 6469 2548
rect 6496 2544 6509 2558
rect 6524 2544 6540 2560
rect 6586 2555 6597 2568
rect 6379 2510 6380 2526
rect 6395 2510 6408 2532
rect 6423 2510 6453 2532
rect 6496 2528 6558 2544
rect 6586 2537 6597 2553
rect 6602 2548 6612 2568
rect 6622 2548 6636 2568
rect 6639 2555 6648 2568
rect 6664 2555 6673 2568
rect 6602 2537 6636 2548
rect 6639 2537 6648 2553
rect 6664 2537 6673 2553
rect 6680 2548 6690 2568
rect 6700 2548 6714 2568
rect 6715 2555 6726 2568
rect 6680 2537 6714 2548
rect 6715 2537 6726 2553
rect 6772 2544 6788 2560
rect 6795 2558 6825 2610
rect 6859 2606 6860 2613
rect 6844 2598 6860 2606
rect 6831 2566 6844 2585
rect 6859 2566 6889 2582
rect 6831 2550 6905 2566
rect 6831 2548 6844 2550
rect 6859 2548 6893 2550
rect 6496 2526 6509 2528
rect 6524 2526 6558 2528
rect 6496 2510 6558 2526
rect 6602 2521 6618 2524
rect 6680 2521 6710 2532
rect 6758 2528 6804 2544
rect 6831 2532 6905 2548
rect 6758 2526 6792 2528
rect 6757 2510 6804 2526
rect 6831 2510 6844 2532
rect 6859 2510 6889 2532
rect 6916 2510 6917 2526
rect 6932 2510 6945 2670
rect 6975 2566 6988 2670
rect 7033 2648 7034 2658
rect 7049 2648 7062 2658
rect 7033 2644 7062 2648
rect 7067 2644 7097 2670
rect 7115 2656 7131 2658
rect 7203 2656 7256 2670
rect 7204 2654 7268 2656
rect 7311 2654 7326 2670
rect 7375 2667 7405 2670
rect 7375 2664 7411 2667
rect 7341 2656 7357 2658
rect 7115 2644 7130 2648
rect 7033 2642 7130 2644
rect 7158 2642 7326 2654
rect 7342 2644 7357 2648
rect 7375 2645 7414 2664
rect 7433 2658 7440 2659
rect 7439 2651 7440 2658
rect 7423 2648 7424 2651
rect 7439 2648 7452 2651
rect 7375 2644 7405 2645
rect 7414 2644 7420 2645
rect 7423 2644 7452 2648
rect 7342 2643 7452 2644
rect 7342 2642 7458 2643
rect 7017 2634 7068 2642
rect 7017 2622 7042 2634
rect 7049 2622 7068 2634
rect 7099 2634 7149 2642
rect 7099 2626 7115 2634
rect 7122 2632 7149 2634
rect 7158 2632 7379 2642
rect 7122 2622 7379 2632
rect 7408 2634 7458 2642
rect 7408 2625 7424 2634
rect 7017 2614 7068 2622
rect 7115 2614 7379 2622
rect 7405 2622 7424 2625
rect 7431 2622 7458 2634
rect 7405 2614 7458 2622
rect 7033 2606 7034 2614
rect 7049 2606 7062 2614
rect 7033 2598 7049 2606
rect 7030 2591 7049 2594
rect 7030 2582 7052 2591
rect 7003 2572 7052 2582
rect 7003 2566 7033 2572
rect 7052 2567 7057 2572
rect 6975 2550 7049 2566
rect 7067 2558 7097 2614
rect 7132 2604 7340 2614
rect 7375 2610 7420 2614
rect 7423 2613 7424 2614
rect 7439 2613 7452 2614
rect 7158 2574 7347 2604
rect 7173 2571 7347 2574
rect 7166 2568 7347 2571
rect 6975 2548 6988 2550
rect 7003 2548 7037 2550
rect 6975 2532 7049 2548
rect 7076 2544 7089 2558
rect 7104 2544 7120 2560
rect 7166 2555 7177 2568
rect 6959 2510 6960 2526
rect 6975 2510 6988 2532
rect 7003 2510 7033 2532
rect 7076 2528 7138 2544
rect 7166 2537 7177 2553
rect 7182 2548 7192 2568
rect 7202 2548 7216 2568
rect 7219 2555 7228 2568
rect 7244 2555 7253 2568
rect 7182 2537 7216 2548
rect 7219 2537 7228 2553
rect 7244 2537 7253 2553
rect 7260 2548 7270 2568
rect 7280 2548 7294 2568
rect 7295 2555 7306 2568
rect 7260 2537 7294 2548
rect 7295 2537 7306 2553
rect 7352 2544 7368 2560
rect 7375 2558 7405 2610
rect 7439 2606 7440 2613
rect 7424 2598 7440 2606
rect 7411 2566 7424 2585
rect 7439 2566 7469 2582
rect 7411 2550 7485 2566
rect 7411 2548 7424 2550
rect 7439 2548 7473 2550
rect 7076 2526 7089 2528
rect 7104 2526 7138 2528
rect 7076 2510 7138 2526
rect 7182 2521 7198 2524
rect 7260 2521 7290 2532
rect 7338 2528 7384 2544
rect 7411 2532 7485 2548
rect 7338 2526 7372 2528
rect 7337 2510 7384 2526
rect 7411 2510 7424 2532
rect 7439 2510 7469 2532
rect 7496 2510 7497 2526
rect 7512 2510 7525 2670
rect 7555 2566 7568 2670
rect 7613 2648 7614 2658
rect 7629 2648 7642 2658
rect 7613 2644 7642 2648
rect 7647 2644 7677 2670
rect 7695 2656 7711 2658
rect 7783 2656 7836 2670
rect 7784 2654 7848 2656
rect 7891 2654 7906 2670
rect 7955 2667 7985 2670
rect 7955 2664 7991 2667
rect 7921 2656 7937 2658
rect 7695 2644 7710 2648
rect 7613 2642 7710 2644
rect 7738 2642 7906 2654
rect 7922 2644 7937 2648
rect 7955 2645 7994 2664
rect 8013 2658 8020 2659
rect 8019 2651 8020 2658
rect 8003 2648 8004 2651
rect 8019 2648 8032 2651
rect 7955 2644 7985 2645
rect 7994 2644 8000 2645
rect 8003 2644 8032 2648
rect 7922 2643 8032 2644
rect 7922 2642 8038 2643
rect 7597 2634 7648 2642
rect 7597 2622 7622 2634
rect 7629 2622 7648 2634
rect 7679 2634 7729 2642
rect 7679 2626 7695 2634
rect 7702 2632 7729 2634
rect 7738 2632 7959 2642
rect 7702 2622 7959 2632
rect 7988 2634 8038 2642
rect 7988 2625 8004 2634
rect 7597 2614 7648 2622
rect 7695 2614 7959 2622
rect 7985 2622 8004 2625
rect 8011 2622 8038 2634
rect 7985 2614 8038 2622
rect 7613 2606 7614 2614
rect 7629 2606 7642 2614
rect 7613 2598 7629 2606
rect 7610 2591 7629 2594
rect 7610 2582 7632 2591
rect 7583 2572 7632 2582
rect 7583 2566 7613 2572
rect 7632 2567 7637 2572
rect 7555 2550 7629 2566
rect 7647 2558 7677 2614
rect 7712 2604 7920 2614
rect 7955 2610 8000 2614
rect 8003 2613 8004 2614
rect 8019 2613 8032 2614
rect 7738 2574 7927 2604
rect 7753 2571 7927 2574
rect 7746 2568 7927 2571
rect 7555 2548 7568 2550
rect 7583 2548 7617 2550
rect 7555 2532 7629 2548
rect 7656 2544 7669 2558
rect 7684 2544 7700 2560
rect 7746 2555 7757 2568
rect 7539 2510 7540 2526
rect 7555 2510 7568 2532
rect 7583 2510 7613 2532
rect 7656 2528 7718 2544
rect 7746 2537 7757 2553
rect 7762 2548 7772 2568
rect 7782 2548 7796 2568
rect 7799 2555 7808 2568
rect 7824 2555 7833 2568
rect 7762 2537 7796 2548
rect 7799 2537 7808 2553
rect 7824 2537 7833 2553
rect 7840 2548 7850 2568
rect 7860 2548 7874 2568
rect 7875 2555 7886 2568
rect 7840 2537 7874 2548
rect 7875 2537 7886 2553
rect 7932 2544 7948 2560
rect 7955 2558 7985 2610
rect 8019 2606 8020 2613
rect 8004 2598 8020 2606
rect 7991 2566 8004 2585
rect 8019 2566 8049 2582
rect 7991 2550 8065 2566
rect 7991 2548 8004 2550
rect 8019 2548 8053 2550
rect 7656 2526 7669 2528
rect 7684 2526 7718 2528
rect 7656 2510 7718 2526
rect 7762 2521 7778 2524
rect 7840 2521 7870 2532
rect 7918 2528 7964 2544
rect 7991 2532 8065 2548
rect 7918 2526 7952 2528
rect 7917 2510 7964 2526
rect 7991 2510 8004 2532
rect 8019 2510 8049 2532
rect 8076 2510 8077 2526
rect 8092 2510 8105 2670
rect 8135 2566 8148 2670
rect 8193 2648 8194 2658
rect 8209 2648 8222 2658
rect 8193 2644 8222 2648
rect 8227 2644 8257 2670
rect 8275 2656 8291 2658
rect 8363 2656 8416 2670
rect 8364 2654 8428 2656
rect 8471 2654 8486 2670
rect 8535 2667 8565 2670
rect 8535 2664 8571 2667
rect 8501 2656 8517 2658
rect 8275 2644 8290 2648
rect 8193 2642 8290 2644
rect 8318 2642 8486 2654
rect 8502 2644 8517 2648
rect 8535 2645 8574 2664
rect 8593 2658 8600 2659
rect 8599 2651 8600 2658
rect 8583 2648 8584 2651
rect 8599 2648 8612 2651
rect 8535 2644 8565 2645
rect 8574 2644 8580 2645
rect 8583 2644 8612 2648
rect 8502 2643 8612 2644
rect 8502 2642 8618 2643
rect 8177 2634 8228 2642
rect 8177 2622 8202 2634
rect 8209 2622 8228 2634
rect 8259 2634 8309 2642
rect 8259 2626 8275 2634
rect 8282 2632 8309 2634
rect 8318 2632 8539 2642
rect 8282 2622 8539 2632
rect 8568 2634 8618 2642
rect 8568 2625 8584 2634
rect 8177 2614 8228 2622
rect 8275 2614 8539 2622
rect 8565 2622 8584 2625
rect 8591 2622 8618 2634
rect 8565 2614 8618 2622
rect 8193 2606 8194 2614
rect 8209 2606 8222 2614
rect 8193 2598 8209 2606
rect 8190 2591 8209 2594
rect 8190 2582 8212 2591
rect 8163 2572 8212 2582
rect 8163 2566 8193 2572
rect 8212 2567 8217 2572
rect 8135 2550 8209 2566
rect 8227 2558 8257 2614
rect 8292 2604 8500 2614
rect 8535 2610 8580 2614
rect 8583 2613 8584 2614
rect 8599 2613 8612 2614
rect 8318 2574 8507 2604
rect 8333 2571 8507 2574
rect 8326 2568 8507 2571
rect 8135 2548 8148 2550
rect 8163 2548 8197 2550
rect 8135 2532 8209 2548
rect 8236 2544 8249 2558
rect 8264 2544 8280 2560
rect 8326 2555 8337 2568
rect 8119 2510 8120 2526
rect 8135 2510 8148 2532
rect 8163 2510 8193 2532
rect 8236 2528 8298 2544
rect 8326 2537 8337 2553
rect 8342 2548 8352 2568
rect 8362 2548 8376 2568
rect 8379 2555 8388 2568
rect 8404 2555 8413 2568
rect 8342 2537 8376 2548
rect 8379 2537 8388 2553
rect 8404 2537 8413 2553
rect 8420 2548 8430 2568
rect 8440 2548 8454 2568
rect 8455 2555 8466 2568
rect 8420 2537 8454 2548
rect 8455 2537 8466 2553
rect 8512 2544 8528 2560
rect 8535 2558 8565 2610
rect 8599 2606 8600 2613
rect 8584 2598 8600 2606
rect 8571 2566 8584 2585
rect 8599 2566 8629 2582
rect 8571 2550 8645 2566
rect 8571 2548 8584 2550
rect 8599 2548 8633 2550
rect 8236 2526 8249 2528
rect 8264 2526 8298 2528
rect 8236 2510 8298 2526
rect 8342 2521 8358 2524
rect 8420 2521 8450 2532
rect 8498 2528 8544 2544
rect 8571 2532 8645 2548
rect 8498 2526 8532 2528
rect 8497 2510 8544 2526
rect 8571 2510 8584 2532
rect 8599 2510 8629 2532
rect 8656 2510 8657 2526
rect 8672 2510 8685 2670
rect 8715 2566 8728 2670
rect 8773 2648 8774 2658
rect 8789 2648 8802 2658
rect 8773 2644 8802 2648
rect 8807 2644 8837 2670
rect 8855 2656 8871 2658
rect 8943 2656 8996 2670
rect 8944 2654 9008 2656
rect 9051 2654 9066 2670
rect 9115 2667 9145 2670
rect 9115 2664 9151 2667
rect 9081 2656 9097 2658
rect 8855 2644 8870 2648
rect 8773 2642 8870 2644
rect 8898 2642 9066 2654
rect 9082 2644 9097 2648
rect 9115 2645 9154 2664
rect 9173 2658 9180 2659
rect 9179 2651 9180 2658
rect 9163 2648 9164 2651
rect 9179 2648 9192 2651
rect 9115 2644 9145 2645
rect 9154 2644 9160 2645
rect 9163 2644 9192 2648
rect 9082 2643 9192 2644
rect 9082 2642 9198 2643
rect 8757 2634 8808 2642
rect 8757 2622 8782 2634
rect 8789 2622 8808 2634
rect 8839 2634 8889 2642
rect 8839 2626 8855 2634
rect 8862 2632 8889 2634
rect 8898 2632 9119 2642
rect 8862 2622 9119 2632
rect 9148 2634 9198 2642
rect 9148 2625 9164 2634
rect 8757 2614 8808 2622
rect 8855 2614 9119 2622
rect 9145 2622 9164 2625
rect 9171 2622 9198 2634
rect 9145 2614 9198 2622
rect 8773 2606 8774 2614
rect 8789 2606 8802 2614
rect 8773 2598 8789 2606
rect 8770 2591 8789 2594
rect 8770 2582 8792 2591
rect 8743 2572 8792 2582
rect 8743 2566 8773 2572
rect 8792 2567 8797 2572
rect 8715 2550 8789 2566
rect 8807 2558 8837 2614
rect 8872 2604 9080 2614
rect 9115 2610 9160 2614
rect 9163 2613 9164 2614
rect 9179 2613 9192 2614
rect 8898 2574 9087 2604
rect 8913 2571 9087 2574
rect 8906 2568 9087 2571
rect 8715 2548 8728 2550
rect 8743 2548 8777 2550
rect 8715 2532 8789 2548
rect 8816 2544 8829 2558
rect 8844 2544 8860 2560
rect 8906 2555 8917 2568
rect 8699 2510 8700 2526
rect 8715 2510 8728 2532
rect 8743 2510 8773 2532
rect 8816 2528 8878 2544
rect 8906 2537 8917 2553
rect 8922 2548 8932 2568
rect 8942 2548 8956 2568
rect 8959 2555 8968 2568
rect 8984 2555 8993 2568
rect 8922 2537 8956 2548
rect 8959 2537 8968 2553
rect 8984 2537 8993 2553
rect 9000 2548 9010 2568
rect 9020 2548 9034 2568
rect 9035 2555 9046 2568
rect 9000 2537 9034 2548
rect 9035 2537 9046 2553
rect 9092 2544 9108 2560
rect 9115 2558 9145 2610
rect 9179 2606 9180 2613
rect 9164 2598 9180 2606
rect 9151 2566 9164 2585
rect 9179 2566 9209 2582
rect 9151 2550 9225 2566
rect 9151 2548 9164 2550
rect 9179 2548 9213 2550
rect 8816 2526 8829 2528
rect 8844 2526 8878 2528
rect 8816 2510 8878 2526
rect 8922 2521 8938 2524
rect 9000 2521 9030 2532
rect 9078 2528 9124 2544
rect 9151 2532 9225 2548
rect 9078 2526 9112 2528
rect 9077 2510 9124 2526
rect 9151 2510 9164 2532
rect 9179 2510 9209 2532
rect 9236 2510 9237 2526
rect 9252 2510 9265 2670
rect -7 2502 34 2510
rect -7 2476 8 2502
rect 15 2476 34 2502
rect 98 2498 160 2510
rect 172 2498 247 2510
rect 305 2498 380 2510
rect 392 2498 423 2510
rect 429 2498 464 2510
rect 98 2496 260 2498
rect -7 2468 34 2476
rect 116 2472 129 2496
rect 144 2494 159 2496
rect -1 2458 0 2468
rect 15 2458 28 2468
rect 43 2458 73 2472
rect 116 2458 159 2472
rect 183 2469 190 2476
rect 193 2472 260 2496
rect 292 2496 464 2498
rect 262 2474 290 2478
rect 292 2474 372 2496
rect 393 2494 408 2496
rect 262 2472 372 2474
rect 193 2468 372 2472
rect 166 2458 196 2468
rect 198 2458 351 2468
rect 359 2458 389 2468
rect 393 2458 423 2472
rect 451 2458 464 2496
rect 536 2502 571 2510
rect 536 2476 537 2502
rect 544 2476 571 2502
rect 479 2458 509 2472
rect 536 2468 571 2476
rect 573 2502 614 2510
rect 573 2476 588 2502
rect 595 2476 614 2502
rect 678 2498 740 2510
rect 752 2498 827 2510
rect 885 2498 960 2510
rect 972 2498 1003 2510
rect 1009 2498 1044 2510
rect 678 2496 840 2498
rect 573 2468 614 2476
rect 696 2472 709 2496
rect 724 2494 739 2496
rect 536 2458 537 2468
rect 552 2458 565 2468
rect 579 2458 580 2468
rect 595 2458 608 2468
rect 623 2458 653 2472
rect 696 2458 739 2472
rect 763 2469 770 2476
rect 773 2472 840 2496
rect 872 2496 1044 2498
rect 842 2474 870 2478
rect 872 2474 952 2496
rect 973 2494 988 2496
rect 842 2472 952 2474
rect 773 2468 952 2472
rect 746 2458 776 2468
rect 778 2458 931 2468
rect 939 2458 969 2468
rect 973 2458 1003 2472
rect 1031 2458 1044 2496
rect 1116 2502 1151 2510
rect 1116 2476 1117 2502
rect 1124 2476 1151 2502
rect 1059 2458 1089 2472
rect 1116 2468 1151 2476
rect 1153 2502 1194 2510
rect 1153 2476 1168 2502
rect 1175 2476 1194 2502
rect 1258 2498 1320 2510
rect 1332 2498 1407 2510
rect 1465 2498 1540 2510
rect 1552 2498 1583 2510
rect 1589 2498 1624 2510
rect 1258 2496 1420 2498
rect 1153 2468 1194 2476
rect 1276 2472 1289 2496
rect 1304 2494 1319 2496
rect 1116 2458 1117 2468
rect 1132 2458 1145 2468
rect 1159 2458 1160 2468
rect 1175 2458 1188 2468
rect 1203 2458 1233 2472
rect 1276 2458 1319 2472
rect 1343 2469 1350 2476
rect 1353 2472 1420 2496
rect 1452 2496 1624 2498
rect 1422 2474 1450 2478
rect 1452 2474 1532 2496
rect 1553 2494 1568 2496
rect 1422 2472 1532 2474
rect 1353 2468 1532 2472
rect 1326 2458 1356 2468
rect 1358 2458 1511 2468
rect 1519 2458 1549 2468
rect 1553 2458 1583 2472
rect 1611 2458 1624 2496
rect 1696 2502 1731 2510
rect 1696 2476 1697 2502
rect 1704 2476 1731 2502
rect 1639 2458 1669 2472
rect 1696 2468 1731 2476
rect 1733 2502 1774 2510
rect 1733 2476 1748 2502
rect 1755 2476 1774 2502
rect 1838 2498 1900 2510
rect 1912 2498 1987 2510
rect 2045 2498 2120 2510
rect 2132 2498 2163 2510
rect 2169 2498 2204 2510
rect 1838 2496 2000 2498
rect 1733 2468 1774 2476
rect 1856 2472 1869 2496
rect 1884 2494 1899 2496
rect 1696 2458 1697 2468
rect 1712 2458 1725 2468
rect 1739 2458 1740 2468
rect 1755 2458 1768 2468
rect 1783 2458 1813 2472
rect 1856 2458 1899 2472
rect 1923 2469 1930 2476
rect 1933 2472 2000 2496
rect 2032 2496 2204 2498
rect 2002 2474 2030 2478
rect 2032 2474 2112 2496
rect 2133 2494 2148 2496
rect 2002 2472 2112 2474
rect 1933 2468 2112 2472
rect 1906 2458 1936 2468
rect 1938 2458 2091 2468
rect 2099 2458 2129 2468
rect 2133 2458 2163 2472
rect 2191 2458 2204 2496
rect 2276 2502 2311 2510
rect 2276 2476 2277 2502
rect 2284 2476 2311 2502
rect 2219 2458 2249 2472
rect 2276 2468 2311 2476
rect 2313 2502 2354 2510
rect 2313 2476 2328 2502
rect 2335 2476 2354 2502
rect 2418 2498 2480 2510
rect 2492 2498 2567 2510
rect 2625 2498 2700 2510
rect 2712 2498 2743 2510
rect 2749 2498 2784 2510
rect 2418 2496 2580 2498
rect 2313 2468 2354 2476
rect 2436 2472 2449 2496
rect 2464 2494 2479 2496
rect 2276 2458 2277 2468
rect 2292 2458 2305 2468
rect 2319 2458 2320 2468
rect 2335 2458 2348 2468
rect 2363 2458 2393 2472
rect 2436 2458 2479 2472
rect 2503 2469 2510 2476
rect 2513 2472 2580 2496
rect 2612 2496 2784 2498
rect 2582 2474 2610 2478
rect 2612 2474 2692 2496
rect 2713 2494 2728 2496
rect 2582 2472 2692 2474
rect 2513 2468 2692 2472
rect 2486 2458 2516 2468
rect 2518 2458 2671 2468
rect 2679 2458 2709 2468
rect 2713 2458 2743 2472
rect 2771 2458 2784 2496
rect 2856 2502 2891 2510
rect 2856 2476 2857 2502
rect 2864 2476 2891 2502
rect 2799 2458 2829 2472
rect 2856 2468 2891 2476
rect 2893 2502 2934 2510
rect 2893 2476 2908 2502
rect 2915 2476 2934 2502
rect 2998 2498 3060 2510
rect 3072 2498 3147 2510
rect 3205 2498 3280 2510
rect 3292 2498 3323 2510
rect 3329 2498 3364 2510
rect 2998 2496 3160 2498
rect 2893 2468 2934 2476
rect 3016 2472 3029 2496
rect 3044 2494 3059 2496
rect 2856 2458 2857 2468
rect 2872 2458 2885 2468
rect 2899 2458 2900 2468
rect 2915 2458 2928 2468
rect 2943 2458 2973 2472
rect 3016 2458 3059 2472
rect 3083 2469 3090 2476
rect 3093 2472 3160 2496
rect 3192 2496 3364 2498
rect 3162 2474 3190 2478
rect 3192 2474 3272 2496
rect 3293 2494 3308 2496
rect 3162 2472 3272 2474
rect 3093 2468 3272 2472
rect 3066 2458 3096 2468
rect 3098 2458 3251 2468
rect 3259 2458 3289 2468
rect 3293 2458 3323 2472
rect 3351 2458 3364 2496
rect 3436 2502 3471 2510
rect 3436 2476 3437 2502
rect 3444 2476 3471 2502
rect 3379 2458 3409 2472
rect 3436 2468 3471 2476
rect 3473 2502 3514 2510
rect 3473 2476 3488 2502
rect 3495 2476 3514 2502
rect 3578 2498 3640 2510
rect 3652 2498 3727 2510
rect 3785 2498 3860 2510
rect 3872 2498 3903 2510
rect 3909 2498 3944 2510
rect 3578 2496 3740 2498
rect 3473 2468 3514 2476
rect 3596 2472 3609 2496
rect 3624 2494 3639 2496
rect 3436 2458 3437 2468
rect 3452 2458 3465 2468
rect 3479 2458 3480 2468
rect 3495 2458 3508 2468
rect 3523 2458 3553 2472
rect 3596 2458 3639 2472
rect 3663 2469 3670 2476
rect 3673 2472 3740 2496
rect 3772 2496 3944 2498
rect 3742 2474 3770 2478
rect 3772 2474 3852 2496
rect 3873 2494 3888 2496
rect 3742 2472 3852 2474
rect 3673 2468 3852 2472
rect 3646 2458 3676 2468
rect 3678 2458 3831 2468
rect 3839 2458 3869 2468
rect 3873 2458 3903 2472
rect 3931 2458 3944 2496
rect 4016 2502 4051 2510
rect 4016 2476 4017 2502
rect 4024 2476 4051 2502
rect 3959 2458 3989 2472
rect 4016 2468 4051 2476
rect 4053 2502 4094 2510
rect 4053 2476 4068 2502
rect 4075 2476 4094 2502
rect 4158 2498 4220 2510
rect 4232 2498 4307 2510
rect 4365 2498 4440 2510
rect 4452 2498 4483 2510
rect 4489 2498 4524 2510
rect 4158 2496 4320 2498
rect 4053 2468 4094 2476
rect 4176 2472 4189 2496
rect 4204 2494 4219 2496
rect 4016 2458 4017 2468
rect 4032 2458 4045 2468
rect 4059 2458 4060 2468
rect 4075 2458 4088 2468
rect 4103 2458 4133 2472
rect 4176 2458 4219 2472
rect 4243 2469 4250 2476
rect 4253 2472 4320 2496
rect 4352 2496 4524 2498
rect 4322 2474 4350 2478
rect 4352 2474 4432 2496
rect 4453 2494 4468 2496
rect 4322 2472 4432 2474
rect 4253 2468 4432 2472
rect 4226 2458 4256 2468
rect 4258 2458 4411 2468
rect 4419 2458 4449 2468
rect 4453 2458 4483 2472
rect 4511 2458 4524 2496
rect 4596 2502 4631 2510
rect 4596 2476 4597 2502
rect 4604 2476 4631 2502
rect 4539 2458 4569 2472
rect 4596 2468 4631 2476
rect 4633 2502 4674 2510
rect 4633 2476 4648 2502
rect 4655 2476 4674 2502
rect 4738 2498 4800 2510
rect 4812 2498 4887 2510
rect 4945 2498 5020 2510
rect 5032 2498 5063 2510
rect 5069 2498 5104 2510
rect 4738 2496 4900 2498
rect 4633 2468 4674 2476
rect 4756 2472 4769 2496
rect 4784 2494 4799 2496
rect 4596 2458 4597 2468
rect 4612 2458 4625 2468
rect 4639 2458 4640 2468
rect 4655 2458 4668 2468
rect 4683 2458 4713 2472
rect 4756 2458 4799 2472
rect 4823 2469 4830 2476
rect 4833 2472 4900 2496
rect 4932 2496 5104 2498
rect 4902 2474 4930 2478
rect 4932 2474 5012 2496
rect 5033 2494 5048 2496
rect 4902 2472 5012 2474
rect 4833 2468 5012 2472
rect 4806 2458 4836 2468
rect 4838 2458 4991 2468
rect 4999 2458 5029 2468
rect 5033 2458 5063 2472
rect 5091 2458 5104 2496
rect 5176 2502 5211 2510
rect 5176 2476 5177 2502
rect 5184 2476 5211 2502
rect 5119 2458 5149 2472
rect 5176 2468 5211 2476
rect 5213 2502 5254 2510
rect 5213 2476 5228 2502
rect 5235 2476 5254 2502
rect 5318 2498 5380 2510
rect 5392 2498 5467 2510
rect 5525 2498 5600 2510
rect 5612 2498 5643 2510
rect 5649 2498 5684 2510
rect 5318 2496 5480 2498
rect 5213 2468 5254 2476
rect 5336 2472 5349 2496
rect 5364 2494 5379 2496
rect 5176 2458 5177 2468
rect 5192 2458 5205 2468
rect 5219 2458 5220 2468
rect 5235 2458 5248 2468
rect 5263 2458 5293 2472
rect 5336 2458 5379 2472
rect 5403 2469 5410 2476
rect 5413 2472 5480 2496
rect 5512 2496 5684 2498
rect 5482 2474 5510 2478
rect 5512 2474 5592 2496
rect 5613 2494 5628 2496
rect 5482 2472 5592 2474
rect 5413 2468 5592 2472
rect 5386 2458 5416 2468
rect 5418 2458 5571 2468
rect 5579 2458 5609 2468
rect 5613 2458 5643 2472
rect 5671 2458 5684 2496
rect 5756 2502 5791 2510
rect 5756 2476 5757 2502
rect 5764 2476 5791 2502
rect 5699 2458 5729 2472
rect 5756 2468 5791 2476
rect 5793 2502 5834 2510
rect 5793 2476 5808 2502
rect 5815 2476 5834 2502
rect 5898 2498 5960 2510
rect 5972 2498 6047 2510
rect 6105 2498 6180 2510
rect 6192 2498 6223 2510
rect 6229 2498 6264 2510
rect 5898 2496 6060 2498
rect 5793 2468 5834 2476
rect 5916 2472 5929 2496
rect 5944 2494 5959 2496
rect 5756 2458 5757 2468
rect 5772 2458 5785 2468
rect 5799 2458 5800 2468
rect 5815 2458 5828 2468
rect 5843 2458 5873 2472
rect 5916 2458 5959 2472
rect 5983 2469 5990 2476
rect 5993 2472 6060 2496
rect 6092 2496 6264 2498
rect 6062 2474 6090 2478
rect 6092 2474 6172 2496
rect 6193 2494 6208 2496
rect 6062 2472 6172 2474
rect 5993 2468 6172 2472
rect 5966 2458 5996 2468
rect 5998 2458 6151 2468
rect 6159 2458 6189 2468
rect 6193 2458 6223 2472
rect 6251 2458 6264 2496
rect 6336 2502 6371 2510
rect 6336 2476 6337 2502
rect 6344 2476 6371 2502
rect 6279 2458 6309 2472
rect 6336 2468 6371 2476
rect 6373 2502 6414 2510
rect 6373 2476 6388 2502
rect 6395 2476 6414 2502
rect 6478 2498 6540 2510
rect 6552 2498 6627 2510
rect 6685 2498 6760 2510
rect 6772 2498 6803 2510
rect 6809 2498 6844 2510
rect 6478 2496 6640 2498
rect 6373 2468 6414 2476
rect 6496 2472 6509 2496
rect 6524 2494 6539 2496
rect 6336 2458 6337 2468
rect 6352 2458 6365 2468
rect 6379 2458 6380 2468
rect 6395 2458 6408 2468
rect 6423 2458 6453 2472
rect 6496 2458 6539 2472
rect 6563 2469 6570 2476
rect 6573 2472 6640 2496
rect 6672 2496 6844 2498
rect 6642 2474 6670 2478
rect 6672 2474 6752 2496
rect 6773 2494 6788 2496
rect 6642 2472 6752 2474
rect 6573 2468 6752 2472
rect 6546 2458 6576 2468
rect 6578 2458 6731 2468
rect 6739 2458 6769 2468
rect 6773 2458 6803 2472
rect 6831 2458 6844 2496
rect 6916 2502 6951 2510
rect 6916 2476 6917 2502
rect 6924 2476 6951 2502
rect 6859 2458 6889 2472
rect 6916 2468 6951 2476
rect 6953 2502 6994 2510
rect 6953 2476 6968 2502
rect 6975 2476 6994 2502
rect 7058 2498 7120 2510
rect 7132 2498 7207 2510
rect 7265 2498 7340 2510
rect 7352 2498 7383 2510
rect 7389 2498 7424 2510
rect 7058 2496 7220 2498
rect 6953 2468 6994 2476
rect 7076 2472 7089 2496
rect 7104 2494 7119 2496
rect 6916 2458 6917 2468
rect 6932 2458 6945 2468
rect 6959 2458 6960 2468
rect 6975 2458 6988 2468
rect 7003 2458 7033 2472
rect 7076 2458 7119 2472
rect 7143 2469 7150 2476
rect 7153 2472 7220 2496
rect 7252 2496 7424 2498
rect 7222 2474 7250 2478
rect 7252 2474 7332 2496
rect 7353 2494 7368 2496
rect 7222 2472 7332 2474
rect 7153 2468 7332 2472
rect 7126 2458 7156 2468
rect 7158 2458 7311 2468
rect 7319 2458 7349 2468
rect 7353 2458 7383 2472
rect 7411 2458 7424 2496
rect 7496 2502 7531 2510
rect 7496 2476 7497 2502
rect 7504 2476 7531 2502
rect 7439 2458 7469 2472
rect 7496 2468 7531 2476
rect 7533 2502 7574 2510
rect 7533 2476 7548 2502
rect 7555 2476 7574 2502
rect 7638 2498 7700 2510
rect 7712 2498 7787 2510
rect 7845 2498 7920 2510
rect 7932 2498 7963 2510
rect 7969 2498 8004 2510
rect 7638 2496 7800 2498
rect 7533 2468 7574 2476
rect 7656 2472 7669 2496
rect 7684 2494 7699 2496
rect 7496 2458 7497 2468
rect 7512 2458 7525 2468
rect 7539 2458 7540 2468
rect 7555 2458 7568 2468
rect 7583 2458 7613 2472
rect 7656 2458 7699 2472
rect 7723 2469 7730 2476
rect 7733 2472 7800 2496
rect 7832 2496 8004 2498
rect 7802 2474 7830 2478
rect 7832 2474 7912 2496
rect 7933 2494 7948 2496
rect 7802 2472 7912 2474
rect 7733 2468 7912 2472
rect 7706 2458 7736 2468
rect 7738 2458 7891 2468
rect 7899 2458 7929 2468
rect 7933 2458 7963 2472
rect 7991 2458 8004 2496
rect 8076 2502 8111 2510
rect 8076 2476 8077 2502
rect 8084 2476 8111 2502
rect 8019 2458 8049 2472
rect 8076 2468 8111 2476
rect 8113 2502 8154 2510
rect 8113 2476 8128 2502
rect 8135 2476 8154 2502
rect 8218 2498 8280 2510
rect 8292 2498 8367 2510
rect 8425 2498 8500 2510
rect 8512 2498 8543 2510
rect 8549 2498 8584 2510
rect 8218 2496 8380 2498
rect 8113 2468 8154 2476
rect 8236 2472 8249 2496
rect 8264 2494 8279 2496
rect 8076 2458 8077 2468
rect 8092 2458 8105 2468
rect 8119 2458 8120 2468
rect 8135 2458 8148 2468
rect 8163 2458 8193 2472
rect 8236 2458 8279 2472
rect 8303 2469 8310 2476
rect 8313 2472 8380 2496
rect 8412 2496 8584 2498
rect 8382 2474 8410 2478
rect 8412 2474 8492 2496
rect 8513 2494 8528 2496
rect 8382 2472 8492 2474
rect 8313 2468 8492 2472
rect 8286 2458 8316 2468
rect 8318 2458 8471 2468
rect 8479 2458 8509 2468
rect 8513 2458 8543 2472
rect 8571 2458 8584 2496
rect 8656 2502 8691 2510
rect 8656 2476 8657 2502
rect 8664 2476 8691 2502
rect 8599 2458 8629 2472
rect 8656 2468 8691 2476
rect 8693 2502 8734 2510
rect 8693 2476 8708 2502
rect 8715 2476 8734 2502
rect 8798 2498 8860 2510
rect 8872 2498 8947 2510
rect 9005 2498 9080 2510
rect 9092 2498 9123 2510
rect 9129 2498 9164 2510
rect 8798 2496 8960 2498
rect 8693 2468 8734 2476
rect 8816 2472 8829 2496
rect 8844 2494 8859 2496
rect 8656 2458 8657 2468
rect 8672 2458 8685 2468
rect 8699 2458 8700 2468
rect 8715 2458 8728 2468
rect 8743 2458 8773 2472
rect 8816 2458 8859 2472
rect 8883 2469 8890 2476
rect 8893 2472 8960 2496
rect 8992 2496 9164 2498
rect 8962 2474 8990 2478
rect 8992 2474 9072 2496
rect 9093 2494 9108 2496
rect 8962 2472 9072 2474
rect 8893 2468 9072 2472
rect 8866 2458 8896 2468
rect 8898 2458 9051 2468
rect 9059 2458 9089 2468
rect 9093 2458 9123 2472
rect 9151 2458 9164 2496
rect 9236 2502 9271 2510
rect 9236 2476 9237 2502
rect 9244 2476 9271 2502
rect 9179 2458 9209 2472
rect 9236 2468 9271 2476
rect 9236 2458 9237 2468
rect 9252 2458 9265 2468
rect -1 2452 9265 2458
rect 0 2444 9265 2452
rect 15 2414 28 2444
rect 43 2426 73 2444
rect 116 2430 130 2444
rect 166 2430 386 2444
rect 117 2428 130 2430
rect 83 2416 98 2428
rect 80 2414 102 2416
rect 107 2414 137 2428
rect 198 2426 351 2430
rect 180 2414 372 2426
rect 415 2414 445 2428
rect 451 2414 464 2444
rect 479 2426 509 2444
rect 552 2414 565 2444
rect 595 2414 608 2444
rect 623 2426 653 2444
rect 696 2430 710 2444
rect 746 2430 966 2444
rect 697 2428 710 2430
rect 663 2416 678 2428
rect 660 2414 682 2416
rect 687 2414 717 2428
rect 778 2426 931 2430
rect 760 2414 952 2426
rect 995 2414 1025 2428
rect 1031 2414 1044 2444
rect 1059 2426 1089 2444
rect 1132 2414 1145 2444
rect 1175 2414 1188 2444
rect 1203 2426 1233 2444
rect 1276 2430 1290 2444
rect 1326 2430 1546 2444
rect 1277 2428 1290 2430
rect 1243 2416 1258 2428
rect 1240 2414 1262 2416
rect 1267 2414 1297 2428
rect 1358 2426 1511 2430
rect 1340 2414 1532 2426
rect 1575 2414 1605 2428
rect 1611 2414 1624 2444
rect 1639 2426 1669 2444
rect 1712 2414 1725 2444
rect 1755 2414 1768 2444
rect 1783 2426 1813 2444
rect 1856 2430 1870 2444
rect 1906 2430 2126 2444
rect 1857 2428 1870 2430
rect 1823 2416 1838 2428
rect 1820 2414 1842 2416
rect 1847 2414 1877 2428
rect 1938 2426 2091 2430
rect 1920 2414 2112 2426
rect 2155 2414 2185 2428
rect 2191 2414 2204 2444
rect 2219 2426 2249 2444
rect 2292 2414 2305 2444
rect 2335 2414 2348 2444
rect 2363 2426 2393 2444
rect 2436 2430 2450 2444
rect 2486 2430 2706 2444
rect 2437 2428 2450 2430
rect 2403 2416 2418 2428
rect 2400 2414 2422 2416
rect 2427 2414 2457 2428
rect 2518 2426 2671 2430
rect 2500 2414 2692 2426
rect 2735 2414 2765 2428
rect 2771 2414 2784 2444
rect 2799 2426 2829 2444
rect 2872 2414 2885 2444
rect 2915 2414 2928 2444
rect 2943 2426 2973 2444
rect 3016 2430 3030 2444
rect 3066 2430 3286 2444
rect 3017 2428 3030 2430
rect 2983 2416 2998 2428
rect 2980 2414 3002 2416
rect 3007 2414 3037 2428
rect 3098 2426 3251 2430
rect 3080 2414 3272 2426
rect 3315 2414 3345 2428
rect 3351 2414 3364 2444
rect 3379 2426 3409 2444
rect 3452 2414 3465 2444
rect 3495 2414 3508 2444
rect 3523 2426 3553 2444
rect 3596 2430 3610 2444
rect 3646 2430 3866 2444
rect 3597 2428 3610 2430
rect 3563 2416 3578 2428
rect 3560 2414 3582 2416
rect 3587 2414 3617 2428
rect 3678 2426 3831 2430
rect 3660 2414 3852 2426
rect 3895 2414 3925 2428
rect 3931 2414 3944 2444
rect 3959 2426 3989 2444
rect 4032 2414 4045 2444
rect 4075 2414 4088 2444
rect 4103 2426 4133 2444
rect 4176 2430 4190 2444
rect 4226 2430 4446 2444
rect 4177 2428 4190 2430
rect 4143 2416 4158 2428
rect 4140 2414 4162 2416
rect 4167 2414 4197 2428
rect 4258 2426 4411 2430
rect 4240 2414 4432 2426
rect 4475 2414 4505 2428
rect 4511 2414 4524 2444
rect 4539 2426 4569 2444
rect 4612 2414 4625 2444
rect 4655 2414 4668 2444
rect 4683 2426 4713 2444
rect 4756 2430 4770 2444
rect 4806 2430 5026 2444
rect 4757 2428 4770 2430
rect 4723 2416 4738 2428
rect 4720 2414 4742 2416
rect 4747 2414 4777 2428
rect 4838 2426 4991 2430
rect 4820 2414 5012 2426
rect 5055 2414 5085 2428
rect 5091 2414 5104 2444
rect 5119 2426 5149 2444
rect 5192 2414 5205 2444
rect 5235 2414 5248 2444
rect 5263 2426 5293 2444
rect 5336 2430 5350 2444
rect 5386 2430 5606 2444
rect 5337 2428 5350 2430
rect 5303 2416 5318 2428
rect 5300 2414 5322 2416
rect 5327 2414 5357 2428
rect 5418 2426 5571 2430
rect 5400 2414 5592 2426
rect 5635 2414 5665 2428
rect 5671 2414 5684 2444
rect 5699 2426 5729 2444
rect 5772 2414 5785 2444
rect 5815 2414 5828 2444
rect 5843 2426 5873 2444
rect 5916 2430 5930 2444
rect 5966 2430 6186 2444
rect 5917 2428 5930 2430
rect 5883 2416 5898 2428
rect 5880 2414 5902 2416
rect 5907 2414 5937 2428
rect 5998 2426 6151 2430
rect 5980 2414 6172 2426
rect 6215 2414 6245 2428
rect 6251 2414 6264 2444
rect 6279 2426 6309 2444
rect 6352 2414 6365 2444
rect 6395 2414 6408 2444
rect 6423 2426 6453 2444
rect 6496 2430 6510 2444
rect 6546 2430 6766 2444
rect 6497 2428 6510 2430
rect 6463 2416 6478 2428
rect 6460 2414 6482 2416
rect 6487 2414 6517 2428
rect 6578 2426 6731 2430
rect 6560 2414 6752 2426
rect 6795 2414 6825 2428
rect 6831 2414 6844 2444
rect 6859 2426 6889 2444
rect 6932 2414 6945 2444
rect 6975 2414 6988 2444
rect 7003 2426 7033 2444
rect 7076 2430 7090 2444
rect 7126 2430 7346 2444
rect 7077 2428 7090 2430
rect 7043 2416 7058 2428
rect 7040 2414 7062 2416
rect 7067 2414 7097 2428
rect 7158 2426 7311 2430
rect 7140 2414 7332 2426
rect 7375 2414 7405 2428
rect 7411 2414 7424 2444
rect 7439 2426 7469 2444
rect 7512 2414 7525 2444
rect 7555 2414 7568 2444
rect 7583 2426 7613 2444
rect 7656 2430 7670 2444
rect 7706 2430 7926 2444
rect 7657 2428 7670 2430
rect 7623 2416 7638 2428
rect 7620 2414 7642 2416
rect 7647 2414 7677 2428
rect 7738 2426 7891 2430
rect 7720 2414 7912 2426
rect 7955 2414 7985 2428
rect 7991 2414 8004 2444
rect 8019 2426 8049 2444
rect 8092 2414 8105 2444
rect 8135 2414 8148 2444
rect 8163 2426 8193 2444
rect 8236 2430 8250 2444
rect 8286 2430 8506 2444
rect 8237 2428 8250 2430
rect 8203 2416 8218 2428
rect 8200 2414 8222 2416
rect 8227 2414 8257 2428
rect 8318 2426 8471 2430
rect 8300 2414 8492 2426
rect 8535 2414 8565 2428
rect 8571 2414 8584 2444
rect 8599 2426 8629 2444
rect 8672 2414 8685 2444
rect 8715 2414 8728 2444
rect 8743 2426 8773 2444
rect 8816 2430 8830 2444
rect 8866 2430 9086 2444
rect 8817 2428 8830 2430
rect 8783 2416 8798 2428
rect 8780 2414 8802 2416
rect 8807 2414 8837 2428
rect 8898 2426 9051 2430
rect 8880 2414 9072 2426
rect 9115 2414 9145 2428
rect 9151 2414 9164 2444
rect 9179 2426 9209 2444
rect 9252 2414 9265 2444
rect 0 2400 9265 2414
rect 15 2296 28 2400
rect 73 2378 74 2388
rect 89 2378 102 2388
rect 73 2374 102 2378
rect 107 2374 137 2400
rect 155 2386 171 2388
rect 243 2386 296 2400
rect 244 2384 308 2386
rect 351 2384 366 2400
rect 415 2397 445 2400
rect 415 2394 451 2397
rect 381 2386 397 2388
rect 155 2374 170 2378
rect 73 2372 170 2374
rect 198 2372 366 2384
rect 382 2374 397 2378
rect 415 2375 454 2394
rect 473 2388 480 2389
rect 479 2381 480 2388
rect 463 2378 464 2381
rect 479 2378 492 2381
rect 415 2374 445 2375
rect 454 2374 460 2375
rect 463 2374 492 2378
rect 382 2373 492 2374
rect 382 2372 498 2373
rect 57 2364 108 2372
rect 57 2352 82 2364
rect 89 2352 108 2364
rect 139 2364 189 2372
rect 139 2356 155 2364
rect 162 2362 189 2364
rect 198 2362 419 2372
rect 162 2352 419 2362
rect 448 2364 498 2372
rect 448 2355 464 2364
rect 57 2344 108 2352
rect 155 2344 419 2352
rect 445 2352 464 2355
rect 471 2352 498 2364
rect 445 2344 498 2352
rect 73 2336 74 2344
rect 89 2336 102 2344
rect 73 2328 89 2336
rect 70 2321 89 2324
rect 70 2312 92 2321
rect 43 2302 92 2312
rect 43 2296 73 2302
rect 92 2297 97 2302
rect 15 2280 89 2296
rect 107 2288 137 2344
rect 172 2334 380 2344
rect 415 2340 460 2344
rect 463 2343 464 2344
rect 479 2343 492 2344
rect 198 2304 387 2334
rect 213 2301 387 2304
rect 206 2298 387 2301
rect 15 2278 28 2280
rect 43 2278 77 2280
rect 15 2262 89 2278
rect 116 2274 129 2288
rect 144 2274 160 2290
rect 206 2285 217 2298
rect -1 2240 0 2256
rect 15 2240 28 2262
rect 43 2240 73 2262
rect 116 2258 178 2274
rect 206 2267 217 2283
rect 222 2278 232 2298
rect 242 2278 256 2298
rect 259 2285 268 2298
rect 284 2285 293 2298
rect 222 2267 256 2278
rect 259 2267 268 2283
rect 284 2267 293 2283
rect 300 2278 310 2298
rect 320 2278 334 2298
rect 335 2285 346 2298
rect 300 2267 334 2278
rect 335 2267 346 2283
rect 392 2274 408 2290
rect 415 2288 445 2340
rect 479 2336 480 2343
rect 464 2328 480 2336
rect 451 2296 464 2315
rect 479 2296 509 2312
rect 451 2280 525 2296
rect 451 2278 464 2280
rect 479 2278 513 2280
rect 116 2256 129 2258
rect 144 2256 178 2258
rect 116 2240 178 2256
rect 222 2251 238 2254
rect 300 2251 330 2262
rect 378 2258 424 2274
rect 451 2262 525 2278
rect 378 2256 412 2258
rect 377 2240 424 2256
rect 451 2240 464 2262
rect 479 2240 509 2262
rect 536 2240 537 2256
rect 552 2240 565 2400
rect 595 2296 608 2400
rect 653 2378 654 2388
rect 669 2378 682 2388
rect 653 2374 682 2378
rect 687 2374 717 2400
rect 735 2386 751 2388
rect 823 2386 876 2400
rect 824 2384 888 2386
rect 931 2384 946 2400
rect 995 2397 1025 2400
rect 995 2394 1031 2397
rect 961 2386 977 2388
rect 735 2374 750 2378
rect 653 2372 750 2374
rect 778 2372 946 2384
rect 962 2374 977 2378
rect 995 2375 1034 2394
rect 1053 2388 1060 2389
rect 1059 2381 1060 2388
rect 1043 2378 1044 2381
rect 1059 2378 1072 2381
rect 995 2374 1025 2375
rect 1034 2374 1040 2375
rect 1043 2374 1072 2378
rect 962 2373 1072 2374
rect 962 2372 1078 2373
rect 637 2364 688 2372
rect 637 2352 662 2364
rect 669 2352 688 2364
rect 719 2364 769 2372
rect 719 2356 735 2364
rect 742 2362 769 2364
rect 778 2362 999 2372
rect 742 2352 999 2362
rect 1028 2364 1078 2372
rect 1028 2355 1044 2364
rect 637 2344 688 2352
rect 735 2344 999 2352
rect 1025 2352 1044 2355
rect 1051 2352 1078 2364
rect 1025 2344 1078 2352
rect 653 2336 654 2344
rect 669 2336 682 2344
rect 653 2328 669 2336
rect 650 2321 669 2324
rect 650 2312 672 2321
rect 623 2302 672 2312
rect 623 2296 653 2302
rect 672 2297 677 2302
rect 595 2280 669 2296
rect 687 2288 717 2344
rect 752 2334 960 2344
rect 995 2340 1040 2344
rect 1043 2343 1044 2344
rect 1059 2343 1072 2344
rect 778 2304 967 2334
rect 793 2301 967 2304
rect 786 2298 967 2301
rect 595 2278 608 2280
rect 623 2278 657 2280
rect 595 2262 669 2278
rect 696 2274 709 2288
rect 724 2274 740 2290
rect 786 2285 797 2298
rect 579 2240 580 2256
rect 595 2240 608 2262
rect 623 2240 653 2262
rect 696 2258 758 2274
rect 786 2267 797 2283
rect 802 2278 812 2298
rect 822 2278 836 2298
rect 839 2285 848 2298
rect 864 2285 873 2298
rect 802 2267 836 2278
rect 839 2267 848 2283
rect 864 2267 873 2283
rect 880 2278 890 2298
rect 900 2278 914 2298
rect 915 2285 926 2298
rect 880 2267 914 2278
rect 915 2267 926 2283
rect 972 2274 988 2290
rect 995 2288 1025 2340
rect 1059 2336 1060 2343
rect 1044 2328 1060 2336
rect 1031 2296 1044 2315
rect 1059 2296 1089 2312
rect 1031 2280 1105 2296
rect 1031 2278 1044 2280
rect 1059 2278 1093 2280
rect 696 2256 709 2258
rect 724 2256 758 2258
rect 696 2240 758 2256
rect 802 2251 818 2254
rect 880 2251 910 2262
rect 958 2258 1004 2274
rect 1031 2262 1105 2278
rect 958 2256 992 2258
rect 957 2240 1004 2256
rect 1031 2240 1044 2262
rect 1059 2240 1089 2262
rect 1116 2240 1117 2256
rect 1132 2240 1145 2400
rect 1175 2296 1188 2400
rect 1233 2378 1234 2388
rect 1249 2378 1262 2388
rect 1233 2374 1262 2378
rect 1267 2374 1297 2400
rect 1315 2386 1331 2388
rect 1403 2386 1456 2400
rect 1404 2384 1468 2386
rect 1511 2384 1526 2400
rect 1575 2397 1605 2400
rect 1575 2394 1611 2397
rect 1541 2386 1557 2388
rect 1315 2374 1330 2378
rect 1233 2372 1330 2374
rect 1358 2372 1526 2384
rect 1542 2374 1557 2378
rect 1575 2375 1614 2394
rect 1633 2388 1640 2389
rect 1639 2381 1640 2388
rect 1623 2378 1624 2381
rect 1639 2378 1652 2381
rect 1575 2374 1605 2375
rect 1614 2374 1620 2375
rect 1623 2374 1652 2378
rect 1542 2373 1652 2374
rect 1542 2372 1658 2373
rect 1217 2364 1268 2372
rect 1217 2352 1242 2364
rect 1249 2352 1268 2364
rect 1299 2364 1349 2372
rect 1299 2356 1315 2364
rect 1322 2362 1349 2364
rect 1358 2362 1579 2372
rect 1322 2352 1579 2362
rect 1608 2364 1658 2372
rect 1608 2355 1624 2364
rect 1217 2344 1268 2352
rect 1315 2344 1579 2352
rect 1605 2352 1624 2355
rect 1631 2352 1658 2364
rect 1605 2344 1658 2352
rect 1233 2336 1234 2344
rect 1249 2336 1262 2344
rect 1233 2328 1249 2336
rect 1230 2321 1249 2324
rect 1230 2312 1252 2321
rect 1203 2302 1252 2312
rect 1203 2296 1233 2302
rect 1252 2297 1257 2302
rect 1175 2280 1249 2296
rect 1267 2288 1297 2344
rect 1332 2334 1540 2344
rect 1575 2340 1620 2344
rect 1623 2343 1624 2344
rect 1639 2343 1652 2344
rect 1358 2304 1547 2334
rect 1373 2301 1547 2304
rect 1366 2298 1547 2301
rect 1175 2278 1188 2280
rect 1203 2278 1237 2280
rect 1175 2262 1249 2278
rect 1276 2274 1289 2288
rect 1304 2274 1320 2290
rect 1366 2285 1377 2298
rect 1159 2240 1160 2256
rect 1175 2240 1188 2262
rect 1203 2240 1233 2262
rect 1276 2258 1338 2274
rect 1366 2267 1377 2283
rect 1382 2278 1392 2298
rect 1402 2278 1416 2298
rect 1419 2285 1428 2298
rect 1444 2285 1453 2298
rect 1382 2267 1416 2278
rect 1419 2267 1428 2283
rect 1444 2267 1453 2283
rect 1460 2278 1470 2298
rect 1480 2278 1494 2298
rect 1495 2285 1506 2298
rect 1460 2267 1494 2278
rect 1495 2267 1506 2283
rect 1552 2274 1568 2290
rect 1575 2288 1605 2340
rect 1639 2336 1640 2343
rect 1624 2328 1640 2336
rect 1611 2296 1624 2315
rect 1639 2296 1669 2312
rect 1611 2280 1685 2296
rect 1611 2278 1624 2280
rect 1639 2278 1673 2280
rect 1276 2256 1289 2258
rect 1304 2256 1338 2258
rect 1276 2240 1338 2256
rect 1382 2251 1398 2254
rect 1460 2251 1490 2262
rect 1538 2258 1584 2274
rect 1611 2262 1685 2278
rect 1538 2256 1572 2258
rect 1537 2240 1584 2256
rect 1611 2240 1624 2262
rect 1639 2240 1669 2262
rect 1696 2240 1697 2256
rect 1712 2240 1725 2400
rect 1755 2296 1768 2400
rect 1813 2378 1814 2388
rect 1829 2378 1842 2388
rect 1813 2374 1842 2378
rect 1847 2374 1877 2400
rect 1895 2386 1911 2388
rect 1983 2386 2036 2400
rect 1984 2384 2048 2386
rect 2091 2384 2106 2400
rect 2155 2397 2185 2400
rect 2155 2394 2191 2397
rect 2121 2386 2137 2388
rect 1895 2374 1910 2378
rect 1813 2372 1910 2374
rect 1938 2372 2106 2384
rect 2122 2374 2137 2378
rect 2155 2375 2194 2394
rect 2213 2388 2220 2389
rect 2219 2381 2220 2388
rect 2203 2378 2204 2381
rect 2219 2378 2232 2381
rect 2155 2374 2185 2375
rect 2194 2374 2200 2375
rect 2203 2374 2232 2378
rect 2122 2373 2232 2374
rect 2122 2372 2238 2373
rect 1797 2364 1848 2372
rect 1797 2352 1822 2364
rect 1829 2352 1848 2364
rect 1879 2364 1929 2372
rect 1879 2356 1895 2364
rect 1902 2362 1929 2364
rect 1938 2362 2159 2372
rect 1902 2352 2159 2362
rect 2188 2364 2238 2372
rect 2188 2355 2204 2364
rect 1797 2344 1848 2352
rect 1895 2344 2159 2352
rect 2185 2352 2204 2355
rect 2211 2352 2238 2364
rect 2185 2344 2238 2352
rect 1813 2336 1814 2344
rect 1829 2336 1842 2344
rect 1813 2328 1829 2336
rect 1810 2321 1829 2324
rect 1810 2312 1832 2321
rect 1783 2302 1832 2312
rect 1783 2296 1813 2302
rect 1832 2297 1837 2302
rect 1755 2280 1829 2296
rect 1847 2288 1877 2344
rect 1912 2334 2120 2344
rect 2155 2340 2200 2344
rect 2203 2343 2204 2344
rect 2219 2343 2232 2344
rect 1938 2304 2127 2334
rect 1953 2301 2127 2304
rect 1946 2298 2127 2301
rect 1755 2278 1768 2280
rect 1783 2278 1817 2280
rect 1755 2262 1829 2278
rect 1856 2274 1869 2288
rect 1884 2274 1900 2290
rect 1946 2285 1957 2298
rect 1739 2240 1740 2256
rect 1755 2240 1768 2262
rect 1783 2240 1813 2262
rect 1856 2258 1918 2274
rect 1946 2267 1957 2283
rect 1962 2278 1972 2298
rect 1982 2278 1996 2298
rect 1999 2285 2008 2298
rect 2024 2285 2033 2298
rect 1962 2267 1996 2278
rect 1999 2267 2008 2283
rect 2024 2267 2033 2283
rect 2040 2278 2050 2298
rect 2060 2278 2074 2298
rect 2075 2285 2086 2298
rect 2040 2267 2074 2278
rect 2075 2267 2086 2283
rect 2132 2274 2148 2290
rect 2155 2288 2185 2340
rect 2219 2336 2220 2343
rect 2204 2328 2220 2336
rect 2191 2296 2204 2315
rect 2219 2296 2249 2312
rect 2191 2280 2265 2296
rect 2191 2278 2204 2280
rect 2219 2278 2253 2280
rect 1856 2256 1869 2258
rect 1884 2256 1918 2258
rect 1856 2240 1918 2256
rect 1962 2251 1976 2254
rect 2040 2251 2070 2262
rect 2118 2258 2164 2274
rect 2191 2262 2265 2278
rect 2118 2256 2152 2258
rect 2117 2240 2164 2256
rect 2191 2240 2204 2262
rect 2219 2240 2249 2262
rect 2276 2240 2277 2256
rect 2292 2240 2305 2400
rect 2335 2296 2348 2400
rect 2393 2378 2394 2388
rect 2409 2378 2422 2388
rect 2393 2374 2422 2378
rect 2427 2374 2457 2400
rect 2475 2386 2491 2388
rect 2563 2386 2616 2400
rect 2564 2384 2628 2386
rect 2671 2384 2686 2400
rect 2735 2397 2765 2400
rect 2735 2394 2771 2397
rect 2701 2386 2717 2388
rect 2475 2374 2490 2378
rect 2393 2372 2490 2374
rect 2518 2372 2686 2384
rect 2702 2374 2717 2378
rect 2735 2375 2774 2394
rect 2793 2388 2800 2389
rect 2799 2381 2800 2388
rect 2783 2378 2784 2381
rect 2799 2378 2812 2381
rect 2735 2374 2765 2375
rect 2774 2374 2780 2375
rect 2783 2374 2812 2378
rect 2702 2373 2812 2374
rect 2702 2372 2818 2373
rect 2377 2364 2428 2372
rect 2377 2352 2402 2364
rect 2409 2352 2428 2364
rect 2459 2364 2509 2372
rect 2459 2356 2475 2364
rect 2482 2362 2509 2364
rect 2518 2362 2739 2372
rect 2482 2352 2739 2362
rect 2768 2364 2818 2372
rect 2768 2355 2784 2364
rect 2377 2344 2428 2352
rect 2475 2344 2739 2352
rect 2765 2352 2784 2355
rect 2791 2352 2818 2364
rect 2765 2344 2818 2352
rect 2393 2336 2394 2344
rect 2409 2336 2422 2344
rect 2393 2328 2409 2336
rect 2390 2321 2409 2324
rect 2390 2312 2412 2321
rect 2363 2302 2412 2312
rect 2363 2296 2393 2302
rect 2412 2297 2417 2302
rect 2335 2280 2409 2296
rect 2427 2288 2457 2344
rect 2492 2334 2700 2344
rect 2735 2340 2780 2344
rect 2783 2343 2784 2344
rect 2799 2343 2812 2344
rect 2518 2304 2707 2334
rect 2533 2301 2707 2304
rect 2526 2298 2707 2301
rect 2335 2278 2348 2280
rect 2363 2278 2397 2280
rect 2335 2262 2409 2278
rect 2436 2274 2449 2288
rect 2464 2274 2480 2290
rect 2526 2285 2537 2298
rect 2319 2240 2320 2256
rect 2335 2240 2348 2262
rect 2363 2240 2393 2262
rect 2436 2258 2498 2274
rect 2526 2267 2537 2283
rect 2542 2278 2552 2298
rect 2562 2278 2576 2298
rect 2579 2285 2588 2298
rect 2604 2285 2613 2298
rect 2542 2267 2576 2278
rect 2579 2267 2588 2283
rect 2604 2267 2613 2283
rect 2620 2278 2630 2298
rect 2640 2278 2654 2298
rect 2655 2285 2666 2298
rect 2620 2267 2654 2278
rect 2655 2267 2666 2283
rect 2712 2274 2728 2290
rect 2735 2288 2765 2340
rect 2799 2336 2800 2343
rect 2784 2328 2800 2336
rect 2771 2296 2784 2315
rect 2799 2296 2829 2312
rect 2771 2280 2845 2296
rect 2771 2278 2784 2280
rect 2799 2278 2833 2280
rect 2436 2256 2449 2258
rect 2464 2256 2498 2258
rect 2436 2240 2498 2256
rect 2542 2251 2558 2254
rect 2620 2251 2650 2262
rect 2698 2258 2744 2274
rect 2771 2262 2845 2278
rect 2698 2256 2732 2258
rect 2697 2240 2744 2256
rect 2771 2240 2784 2262
rect 2799 2240 2829 2262
rect 2856 2240 2857 2256
rect 2872 2240 2885 2400
rect 2915 2296 2928 2400
rect 2973 2378 2974 2388
rect 2989 2378 3002 2388
rect 2973 2374 3002 2378
rect 3007 2374 3037 2400
rect 3055 2386 3071 2388
rect 3143 2386 3196 2400
rect 3144 2384 3208 2386
rect 3251 2384 3266 2400
rect 3315 2397 3345 2400
rect 3315 2394 3351 2397
rect 3281 2386 3297 2388
rect 3055 2374 3070 2378
rect 2973 2372 3070 2374
rect 3098 2372 3266 2384
rect 3282 2374 3297 2378
rect 3315 2375 3354 2394
rect 3373 2388 3380 2389
rect 3379 2381 3380 2388
rect 3363 2378 3364 2381
rect 3379 2378 3392 2381
rect 3315 2374 3345 2375
rect 3354 2374 3360 2375
rect 3363 2374 3392 2378
rect 3282 2373 3392 2374
rect 3282 2372 3398 2373
rect 2957 2364 3008 2372
rect 2957 2352 2982 2364
rect 2989 2352 3008 2364
rect 3039 2364 3089 2372
rect 3039 2356 3055 2364
rect 3062 2362 3089 2364
rect 3098 2362 3319 2372
rect 3062 2352 3319 2362
rect 3348 2364 3398 2372
rect 3348 2355 3364 2364
rect 2957 2344 3008 2352
rect 3055 2344 3319 2352
rect 3345 2352 3364 2355
rect 3371 2352 3398 2364
rect 3345 2344 3398 2352
rect 2973 2336 2974 2344
rect 2989 2336 3002 2344
rect 2973 2328 2989 2336
rect 2970 2321 2989 2324
rect 2970 2312 2992 2321
rect 2943 2302 2992 2312
rect 2943 2296 2973 2302
rect 2992 2297 2997 2302
rect 2915 2280 2989 2296
rect 3007 2288 3037 2344
rect 3072 2334 3280 2344
rect 3315 2340 3360 2344
rect 3363 2343 3364 2344
rect 3379 2343 3392 2344
rect 3098 2304 3287 2334
rect 3113 2301 3287 2304
rect 3106 2298 3287 2301
rect 2915 2278 2928 2280
rect 2943 2278 2977 2280
rect 2915 2262 2989 2278
rect 3016 2274 3029 2288
rect 3044 2274 3060 2290
rect 3106 2285 3117 2298
rect 2899 2240 2900 2256
rect 2915 2240 2928 2262
rect 2943 2240 2973 2262
rect 3016 2258 3078 2274
rect 3106 2267 3117 2283
rect 3122 2278 3132 2298
rect 3142 2278 3156 2298
rect 3159 2285 3168 2298
rect 3184 2285 3193 2298
rect 3122 2267 3156 2278
rect 3159 2267 3168 2283
rect 3184 2267 3193 2283
rect 3200 2278 3210 2298
rect 3220 2278 3234 2298
rect 3235 2285 3246 2298
rect 3200 2267 3234 2278
rect 3235 2267 3246 2283
rect 3292 2274 3308 2290
rect 3315 2288 3345 2340
rect 3379 2336 3380 2343
rect 3364 2328 3380 2336
rect 3351 2296 3364 2315
rect 3379 2296 3409 2312
rect 3351 2280 3425 2296
rect 3351 2278 3364 2280
rect 3379 2278 3413 2280
rect 3016 2256 3029 2258
rect 3044 2256 3078 2258
rect 3016 2240 3078 2256
rect 3122 2251 3138 2254
rect 3200 2251 3230 2262
rect 3278 2258 3324 2274
rect 3351 2262 3425 2278
rect 3278 2256 3312 2258
rect 3277 2240 3324 2256
rect 3351 2240 3364 2262
rect 3379 2240 3409 2262
rect 3436 2240 3437 2256
rect 3452 2240 3465 2400
rect 3495 2296 3508 2400
rect 3553 2378 3554 2388
rect 3569 2378 3582 2388
rect 3553 2374 3582 2378
rect 3587 2374 3617 2400
rect 3635 2386 3651 2388
rect 3723 2386 3776 2400
rect 3724 2384 3788 2386
rect 3831 2384 3846 2400
rect 3895 2397 3925 2400
rect 3895 2394 3931 2397
rect 3861 2386 3877 2388
rect 3635 2374 3650 2378
rect 3553 2372 3650 2374
rect 3678 2372 3846 2384
rect 3862 2374 3877 2378
rect 3895 2375 3934 2394
rect 3953 2388 3960 2389
rect 3959 2381 3960 2388
rect 3943 2378 3944 2381
rect 3959 2378 3972 2381
rect 3895 2374 3925 2375
rect 3934 2374 3940 2375
rect 3943 2374 3972 2378
rect 3862 2373 3972 2374
rect 3862 2372 3978 2373
rect 3537 2364 3588 2372
rect 3537 2352 3562 2364
rect 3569 2352 3588 2364
rect 3619 2364 3669 2372
rect 3619 2356 3635 2364
rect 3642 2362 3669 2364
rect 3678 2362 3899 2372
rect 3642 2352 3899 2362
rect 3928 2364 3978 2372
rect 3928 2355 3944 2364
rect 3537 2344 3588 2352
rect 3635 2344 3899 2352
rect 3925 2352 3944 2355
rect 3951 2352 3978 2364
rect 3925 2344 3978 2352
rect 3553 2336 3554 2344
rect 3569 2336 3582 2344
rect 3553 2328 3569 2336
rect 3550 2321 3569 2324
rect 3550 2312 3572 2321
rect 3523 2302 3572 2312
rect 3523 2296 3553 2302
rect 3572 2297 3577 2302
rect 3495 2280 3569 2296
rect 3587 2288 3617 2344
rect 3652 2334 3860 2344
rect 3895 2340 3940 2344
rect 3943 2343 3944 2344
rect 3959 2343 3972 2344
rect 3678 2304 3867 2334
rect 3693 2301 3867 2304
rect 3686 2298 3867 2301
rect 3495 2278 3508 2280
rect 3523 2278 3557 2280
rect 3495 2262 3569 2278
rect 3596 2274 3609 2288
rect 3624 2274 3640 2290
rect 3686 2285 3697 2298
rect 3479 2240 3480 2256
rect 3495 2240 3508 2262
rect 3523 2240 3553 2262
rect 3596 2258 3658 2274
rect 3686 2267 3697 2283
rect 3702 2278 3712 2298
rect 3722 2278 3736 2298
rect 3739 2285 3748 2298
rect 3764 2285 3773 2298
rect 3702 2267 3736 2278
rect 3739 2267 3748 2283
rect 3764 2267 3773 2283
rect 3780 2278 3790 2298
rect 3800 2278 3814 2298
rect 3815 2285 3826 2298
rect 3780 2267 3814 2278
rect 3815 2267 3826 2283
rect 3872 2274 3888 2290
rect 3895 2288 3925 2340
rect 3959 2336 3960 2343
rect 3944 2328 3960 2336
rect 3931 2296 3944 2315
rect 3959 2296 3989 2312
rect 3931 2280 4005 2296
rect 3931 2278 3944 2280
rect 3959 2278 3993 2280
rect 3596 2256 3609 2258
rect 3624 2256 3658 2258
rect 3596 2240 3658 2256
rect 3702 2251 3718 2254
rect 3780 2251 3810 2262
rect 3858 2258 3904 2274
rect 3931 2262 4005 2278
rect 3858 2256 3892 2258
rect 3857 2240 3904 2256
rect 3931 2240 3944 2262
rect 3959 2240 3989 2262
rect 4016 2240 4017 2256
rect 4032 2240 4045 2400
rect 4075 2296 4088 2400
rect 4133 2378 4134 2388
rect 4149 2378 4162 2388
rect 4133 2374 4162 2378
rect 4167 2374 4197 2400
rect 4215 2386 4231 2388
rect 4303 2386 4356 2400
rect 4304 2384 4368 2386
rect 4411 2384 4426 2400
rect 4475 2397 4505 2400
rect 4475 2394 4511 2397
rect 4441 2386 4457 2388
rect 4215 2374 4230 2378
rect 4133 2372 4230 2374
rect 4258 2372 4426 2384
rect 4442 2374 4457 2378
rect 4475 2375 4514 2394
rect 4533 2388 4540 2389
rect 4539 2381 4540 2388
rect 4523 2378 4524 2381
rect 4539 2378 4552 2381
rect 4475 2374 4505 2375
rect 4514 2374 4520 2375
rect 4523 2374 4552 2378
rect 4442 2373 4552 2374
rect 4442 2372 4558 2373
rect 4117 2364 4168 2372
rect 4117 2352 4142 2364
rect 4149 2352 4168 2364
rect 4199 2364 4249 2372
rect 4199 2356 4215 2364
rect 4222 2362 4249 2364
rect 4258 2362 4479 2372
rect 4222 2352 4479 2362
rect 4508 2364 4558 2372
rect 4508 2355 4524 2364
rect 4117 2344 4168 2352
rect 4215 2344 4479 2352
rect 4505 2352 4524 2355
rect 4531 2352 4558 2364
rect 4505 2344 4558 2352
rect 4133 2336 4134 2344
rect 4149 2336 4162 2344
rect 4133 2328 4149 2336
rect 4130 2321 4149 2324
rect 4130 2312 4152 2321
rect 4103 2302 4152 2312
rect 4103 2296 4133 2302
rect 4152 2297 4157 2302
rect 4075 2280 4149 2296
rect 4167 2288 4197 2344
rect 4232 2334 4440 2344
rect 4475 2340 4520 2344
rect 4523 2343 4524 2344
rect 4539 2343 4552 2344
rect 4258 2304 4447 2334
rect 4273 2301 4447 2304
rect 4266 2298 4447 2301
rect 4075 2278 4088 2280
rect 4103 2278 4137 2280
rect 4075 2262 4149 2278
rect 4176 2274 4189 2288
rect 4204 2274 4220 2290
rect 4266 2285 4277 2298
rect 4059 2240 4060 2256
rect 4075 2240 4088 2262
rect 4103 2240 4133 2262
rect 4176 2258 4238 2274
rect 4266 2267 4277 2283
rect 4282 2278 4292 2298
rect 4302 2278 4316 2298
rect 4319 2285 4328 2298
rect 4344 2285 4353 2298
rect 4282 2267 4316 2278
rect 4319 2267 4328 2283
rect 4344 2267 4353 2283
rect 4360 2278 4370 2298
rect 4380 2278 4394 2298
rect 4395 2285 4406 2298
rect 4360 2267 4394 2278
rect 4395 2267 4406 2283
rect 4452 2274 4468 2290
rect 4475 2288 4505 2340
rect 4539 2336 4540 2343
rect 4524 2328 4540 2336
rect 4511 2296 4524 2315
rect 4539 2296 4569 2312
rect 4511 2280 4585 2296
rect 4511 2278 4524 2280
rect 4539 2278 4573 2280
rect 4176 2256 4189 2258
rect 4204 2256 4238 2258
rect 4176 2240 4238 2256
rect 4282 2251 4298 2254
rect 4360 2251 4390 2262
rect 4438 2258 4484 2274
rect 4511 2262 4585 2278
rect 4438 2256 4472 2258
rect 4437 2240 4484 2256
rect 4511 2240 4524 2262
rect 4539 2240 4569 2262
rect 4596 2240 4597 2256
rect 4612 2240 4625 2400
rect 4655 2296 4668 2400
rect 4713 2378 4714 2388
rect 4729 2378 4742 2388
rect 4713 2374 4742 2378
rect 4747 2374 4777 2400
rect 4795 2386 4811 2388
rect 4883 2386 4936 2400
rect 4884 2384 4948 2386
rect 4991 2384 5006 2400
rect 5055 2397 5085 2400
rect 5055 2394 5091 2397
rect 5021 2386 5037 2388
rect 4795 2374 4810 2378
rect 4713 2372 4810 2374
rect 4838 2372 5006 2384
rect 5022 2374 5037 2378
rect 5055 2375 5094 2394
rect 5113 2388 5120 2389
rect 5119 2381 5120 2388
rect 5103 2378 5104 2381
rect 5119 2378 5132 2381
rect 5055 2374 5085 2375
rect 5094 2374 5100 2375
rect 5103 2374 5132 2378
rect 5022 2373 5132 2374
rect 5022 2372 5138 2373
rect 4697 2364 4748 2372
rect 4697 2352 4722 2364
rect 4729 2352 4748 2364
rect 4779 2364 4829 2372
rect 4779 2356 4795 2364
rect 4802 2362 4829 2364
rect 4838 2362 5059 2372
rect 4802 2352 5059 2362
rect 5088 2364 5138 2372
rect 5088 2355 5104 2364
rect 4697 2344 4748 2352
rect 4795 2344 5059 2352
rect 5085 2352 5104 2355
rect 5111 2352 5138 2364
rect 5085 2344 5138 2352
rect 4713 2336 4714 2344
rect 4729 2336 4742 2344
rect 4713 2328 4729 2336
rect 4710 2321 4729 2324
rect 4710 2312 4732 2321
rect 4683 2302 4732 2312
rect 4683 2296 4713 2302
rect 4732 2297 4737 2302
rect 4655 2280 4729 2296
rect 4747 2288 4777 2344
rect 4812 2334 5020 2344
rect 5055 2340 5100 2344
rect 5103 2343 5104 2344
rect 5119 2343 5132 2344
rect 4838 2304 5027 2334
rect 4853 2301 5027 2304
rect 4846 2298 5027 2301
rect 4655 2278 4668 2280
rect 4683 2278 4717 2280
rect 4655 2262 4729 2278
rect 4756 2274 4769 2288
rect 4784 2274 4800 2290
rect 4846 2285 4857 2298
rect 4639 2240 4640 2256
rect 4655 2240 4668 2262
rect 4683 2240 4713 2262
rect 4756 2258 4818 2274
rect 4846 2267 4857 2283
rect 4862 2278 4872 2298
rect 4882 2278 4896 2298
rect 4899 2285 4908 2298
rect 4924 2285 4933 2298
rect 4862 2267 4896 2278
rect 4899 2267 4908 2283
rect 4924 2267 4933 2283
rect 4940 2278 4950 2298
rect 4960 2278 4974 2298
rect 4975 2285 4986 2298
rect 4940 2267 4974 2278
rect 4975 2267 4986 2283
rect 5032 2274 5048 2290
rect 5055 2288 5085 2340
rect 5119 2336 5120 2343
rect 5104 2328 5120 2336
rect 5091 2296 5104 2315
rect 5119 2296 5149 2312
rect 5091 2280 5165 2296
rect 5091 2278 5104 2280
rect 5119 2278 5153 2280
rect 4756 2256 4769 2258
rect 4784 2256 4818 2258
rect 4756 2240 4818 2256
rect 4862 2251 4878 2254
rect 4940 2251 4970 2262
rect 5018 2258 5064 2274
rect 5091 2262 5165 2278
rect 5018 2256 5052 2258
rect 5017 2240 5064 2256
rect 5091 2240 5104 2262
rect 5119 2240 5149 2262
rect 5176 2240 5177 2256
rect 5192 2240 5205 2400
rect 5235 2296 5248 2400
rect 5293 2378 5294 2388
rect 5309 2378 5322 2388
rect 5293 2374 5322 2378
rect 5327 2374 5357 2400
rect 5375 2386 5391 2388
rect 5463 2386 5516 2400
rect 5464 2384 5528 2386
rect 5571 2384 5586 2400
rect 5635 2397 5665 2400
rect 5635 2394 5671 2397
rect 5601 2386 5617 2388
rect 5375 2374 5390 2378
rect 5293 2372 5390 2374
rect 5418 2372 5586 2384
rect 5602 2374 5617 2378
rect 5635 2375 5674 2394
rect 5693 2388 5700 2389
rect 5699 2381 5700 2388
rect 5683 2378 5684 2381
rect 5699 2378 5712 2381
rect 5635 2374 5665 2375
rect 5674 2374 5680 2375
rect 5683 2374 5712 2378
rect 5602 2373 5712 2374
rect 5602 2372 5718 2373
rect 5277 2364 5328 2372
rect 5277 2352 5302 2364
rect 5309 2352 5328 2364
rect 5359 2364 5409 2372
rect 5359 2356 5375 2364
rect 5382 2362 5409 2364
rect 5418 2362 5639 2372
rect 5382 2352 5639 2362
rect 5668 2364 5718 2372
rect 5668 2355 5684 2364
rect 5277 2344 5328 2352
rect 5375 2344 5639 2352
rect 5665 2352 5684 2355
rect 5691 2352 5718 2364
rect 5665 2344 5718 2352
rect 5293 2336 5294 2344
rect 5309 2336 5322 2344
rect 5293 2328 5309 2336
rect 5290 2321 5309 2324
rect 5290 2312 5312 2321
rect 5263 2302 5312 2312
rect 5263 2296 5293 2302
rect 5312 2297 5317 2302
rect 5235 2280 5309 2296
rect 5327 2288 5357 2344
rect 5392 2334 5600 2344
rect 5635 2340 5680 2344
rect 5683 2343 5684 2344
rect 5699 2343 5712 2344
rect 5418 2304 5607 2334
rect 5433 2301 5607 2304
rect 5426 2298 5607 2301
rect 5235 2278 5248 2280
rect 5263 2278 5297 2280
rect 5235 2262 5309 2278
rect 5336 2274 5349 2288
rect 5364 2274 5380 2290
rect 5426 2285 5437 2298
rect 5219 2240 5220 2256
rect 5235 2240 5248 2262
rect 5263 2240 5293 2262
rect 5336 2258 5398 2274
rect 5426 2267 5437 2283
rect 5442 2278 5452 2298
rect 5462 2278 5476 2298
rect 5479 2285 5488 2298
rect 5504 2285 5513 2298
rect 5442 2267 5476 2278
rect 5479 2267 5488 2283
rect 5504 2267 5513 2283
rect 5520 2278 5530 2298
rect 5540 2278 5554 2298
rect 5555 2285 5566 2298
rect 5520 2267 5554 2278
rect 5555 2267 5566 2283
rect 5612 2274 5628 2290
rect 5635 2288 5665 2340
rect 5699 2336 5700 2343
rect 5684 2328 5700 2336
rect 5671 2296 5684 2315
rect 5699 2296 5729 2312
rect 5671 2280 5745 2296
rect 5671 2278 5684 2280
rect 5699 2278 5733 2280
rect 5336 2256 5349 2258
rect 5364 2256 5398 2258
rect 5336 2240 5398 2256
rect 5442 2251 5458 2254
rect 5520 2251 5550 2262
rect 5598 2258 5644 2274
rect 5671 2262 5745 2278
rect 5598 2256 5632 2258
rect 5597 2240 5644 2256
rect 5671 2240 5684 2262
rect 5699 2240 5729 2262
rect 5756 2240 5757 2256
rect 5772 2240 5785 2400
rect 5815 2296 5828 2400
rect 5873 2378 5874 2388
rect 5889 2378 5902 2388
rect 5873 2374 5902 2378
rect 5907 2374 5937 2400
rect 5955 2386 5971 2388
rect 6043 2386 6096 2400
rect 6044 2384 6108 2386
rect 6151 2384 6166 2400
rect 6215 2397 6245 2400
rect 6215 2394 6251 2397
rect 6181 2386 6197 2388
rect 5955 2374 5970 2378
rect 5873 2372 5970 2374
rect 5998 2372 6166 2384
rect 6182 2374 6197 2378
rect 6215 2375 6254 2394
rect 6273 2388 6280 2389
rect 6279 2381 6280 2388
rect 6263 2378 6264 2381
rect 6279 2378 6292 2381
rect 6215 2374 6245 2375
rect 6254 2374 6260 2375
rect 6263 2374 6292 2378
rect 6182 2373 6292 2374
rect 6182 2372 6298 2373
rect 5857 2364 5908 2372
rect 5857 2352 5882 2364
rect 5889 2352 5908 2364
rect 5939 2364 5989 2372
rect 5939 2356 5955 2364
rect 5962 2362 5989 2364
rect 5998 2362 6219 2372
rect 5962 2352 6219 2362
rect 6248 2364 6298 2372
rect 6248 2355 6264 2364
rect 5857 2344 5908 2352
rect 5955 2344 6219 2352
rect 6245 2352 6264 2355
rect 6271 2352 6298 2364
rect 6245 2344 6298 2352
rect 5873 2336 5874 2344
rect 5889 2336 5902 2344
rect 5873 2328 5889 2336
rect 5870 2321 5889 2324
rect 5870 2312 5892 2321
rect 5843 2302 5892 2312
rect 5843 2296 5873 2302
rect 5892 2297 5897 2302
rect 5815 2280 5889 2296
rect 5907 2288 5937 2344
rect 5972 2334 6180 2344
rect 6215 2340 6260 2344
rect 6263 2343 6264 2344
rect 6279 2343 6292 2344
rect 5998 2304 6187 2334
rect 6013 2301 6187 2304
rect 6006 2298 6187 2301
rect 5815 2278 5828 2280
rect 5843 2278 5877 2280
rect 5815 2262 5889 2278
rect 5916 2274 5929 2288
rect 5944 2274 5960 2290
rect 6006 2285 6017 2298
rect 5799 2240 5800 2256
rect 5815 2240 5828 2262
rect 5843 2240 5873 2262
rect 5916 2258 5978 2274
rect 6006 2267 6017 2283
rect 6022 2278 6032 2298
rect 6042 2278 6056 2298
rect 6059 2285 6068 2298
rect 6084 2285 6093 2298
rect 6022 2267 6056 2278
rect 6059 2267 6068 2283
rect 6084 2267 6093 2283
rect 6100 2278 6110 2298
rect 6120 2278 6134 2298
rect 6135 2285 6146 2298
rect 6100 2267 6134 2278
rect 6135 2267 6146 2283
rect 6192 2274 6208 2290
rect 6215 2288 6245 2340
rect 6279 2336 6280 2343
rect 6264 2328 6280 2336
rect 6251 2296 6264 2315
rect 6279 2296 6309 2312
rect 6251 2280 6325 2296
rect 6251 2278 6264 2280
rect 6279 2278 6313 2280
rect 5916 2256 5929 2258
rect 5944 2256 5978 2258
rect 5916 2240 5978 2256
rect 6022 2251 6038 2254
rect 6100 2251 6130 2262
rect 6178 2258 6224 2274
rect 6251 2262 6325 2278
rect 6178 2256 6212 2258
rect 6177 2240 6224 2256
rect 6251 2240 6264 2262
rect 6279 2240 6309 2262
rect 6336 2240 6337 2256
rect 6352 2240 6365 2400
rect 6395 2296 6408 2400
rect 6453 2378 6454 2388
rect 6469 2378 6482 2388
rect 6453 2374 6482 2378
rect 6487 2374 6517 2400
rect 6535 2386 6551 2388
rect 6623 2386 6676 2400
rect 6624 2384 6688 2386
rect 6731 2384 6746 2400
rect 6795 2397 6825 2400
rect 6795 2394 6831 2397
rect 6761 2386 6777 2388
rect 6535 2374 6550 2378
rect 6453 2372 6550 2374
rect 6578 2372 6746 2384
rect 6762 2374 6777 2378
rect 6795 2375 6834 2394
rect 6853 2388 6860 2389
rect 6859 2381 6860 2388
rect 6843 2378 6844 2381
rect 6859 2378 6872 2381
rect 6795 2374 6825 2375
rect 6834 2374 6840 2375
rect 6843 2374 6872 2378
rect 6762 2373 6872 2374
rect 6762 2372 6878 2373
rect 6437 2364 6488 2372
rect 6437 2352 6462 2364
rect 6469 2352 6488 2364
rect 6519 2364 6569 2372
rect 6519 2356 6535 2364
rect 6542 2362 6569 2364
rect 6578 2362 6799 2372
rect 6542 2352 6799 2362
rect 6828 2364 6878 2372
rect 6828 2355 6844 2364
rect 6437 2344 6488 2352
rect 6535 2344 6799 2352
rect 6825 2352 6844 2355
rect 6851 2352 6878 2364
rect 6825 2344 6878 2352
rect 6453 2336 6454 2344
rect 6469 2336 6482 2344
rect 6453 2328 6469 2336
rect 6450 2321 6469 2324
rect 6450 2312 6472 2321
rect 6423 2302 6472 2312
rect 6423 2296 6453 2302
rect 6472 2297 6477 2302
rect 6395 2280 6469 2296
rect 6487 2288 6517 2344
rect 6552 2334 6760 2344
rect 6795 2340 6840 2344
rect 6843 2343 6844 2344
rect 6859 2343 6872 2344
rect 6578 2304 6767 2334
rect 6593 2301 6767 2304
rect 6586 2298 6767 2301
rect 6395 2278 6408 2280
rect 6423 2278 6457 2280
rect 6395 2262 6469 2278
rect 6496 2274 6509 2288
rect 6524 2274 6540 2290
rect 6586 2285 6597 2298
rect 6379 2240 6380 2256
rect 6395 2240 6408 2262
rect 6423 2240 6453 2262
rect 6496 2258 6558 2274
rect 6586 2267 6597 2283
rect 6602 2278 6612 2298
rect 6622 2278 6636 2298
rect 6639 2285 6648 2298
rect 6664 2285 6673 2298
rect 6602 2267 6636 2278
rect 6639 2267 6648 2283
rect 6664 2267 6673 2283
rect 6680 2278 6690 2298
rect 6700 2278 6714 2298
rect 6715 2285 6726 2298
rect 6680 2267 6714 2278
rect 6715 2267 6726 2283
rect 6772 2274 6788 2290
rect 6795 2288 6825 2340
rect 6859 2336 6860 2343
rect 6844 2328 6860 2336
rect 6831 2296 6844 2315
rect 6859 2296 6889 2312
rect 6831 2280 6905 2296
rect 6831 2278 6844 2280
rect 6859 2278 6893 2280
rect 6496 2256 6509 2258
rect 6524 2256 6558 2258
rect 6496 2240 6558 2256
rect 6602 2251 6618 2254
rect 6680 2251 6710 2262
rect 6758 2258 6804 2274
rect 6831 2262 6905 2278
rect 6758 2256 6792 2258
rect 6757 2240 6804 2256
rect 6831 2240 6844 2262
rect 6859 2240 6889 2262
rect 6916 2240 6917 2256
rect 6932 2240 6945 2400
rect 6975 2296 6988 2400
rect 7033 2378 7034 2388
rect 7049 2378 7062 2388
rect 7033 2374 7062 2378
rect 7067 2374 7097 2400
rect 7115 2386 7131 2388
rect 7203 2386 7256 2400
rect 7204 2384 7268 2386
rect 7311 2384 7326 2400
rect 7375 2397 7405 2400
rect 7375 2394 7411 2397
rect 7341 2386 7357 2388
rect 7115 2374 7130 2378
rect 7033 2372 7130 2374
rect 7158 2372 7326 2384
rect 7342 2374 7357 2378
rect 7375 2375 7414 2394
rect 7433 2388 7440 2389
rect 7439 2381 7440 2388
rect 7423 2378 7424 2381
rect 7439 2378 7452 2381
rect 7375 2374 7405 2375
rect 7414 2374 7420 2375
rect 7423 2374 7452 2378
rect 7342 2373 7452 2374
rect 7342 2372 7458 2373
rect 7017 2364 7068 2372
rect 7017 2352 7042 2364
rect 7049 2352 7068 2364
rect 7099 2364 7149 2372
rect 7099 2356 7115 2364
rect 7122 2362 7149 2364
rect 7158 2362 7379 2372
rect 7122 2352 7379 2362
rect 7408 2364 7458 2372
rect 7408 2355 7424 2364
rect 7017 2344 7068 2352
rect 7115 2344 7379 2352
rect 7405 2352 7424 2355
rect 7431 2352 7458 2364
rect 7405 2344 7458 2352
rect 7033 2336 7034 2344
rect 7049 2336 7062 2344
rect 7033 2328 7049 2336
rect 7030 2321 7049 2324
rect 7030 2312 7052 2321
rect 7003 2302 7052 2312
rect 7003 2296 7033 2302
rect 7052 2297 7057 2302
rect 6975 2280 7049 2296
rect 7067 2288 7097 2344
rect 7132 2334 7340 2344
rect 7375 2340 7420 2344
rect 7423 2343 7424 2344
rect 7439 2343 7452 2344
rect 7158 2304 7347 2334
rect 7173 2301 7347 2304
rect 7166 2298 7347 2301
rect 6975 2278 6988 2280
rect 7003 2278 7037 2280
rect 6975 2262 7049 2278
rect 7076 2274 7089 2288
rect 7104 2274 7120 2290
rect 7166 2285 7177 2298
rect 6959 2240 6960 2256
rect 6975 2240 6988 2262
rect 7003 2240 7033 2262
rect 7076 2258 7138 2274
rect 7166 2267 7177 2283
rect 7182 2278 7192 2298
rect 7202 2278 7216 2298
rect 7219 2285 7228 2298
rect 7244 2285 7253 2298
rect 7182 2267 7216 2278
rect 7219 2267 7228 2283
rect 7244 2267 7253 2283
rect 7260 2278 7270 2298
rect 7280 2278 7294 2298
rect 7295 2285 7306 2298
rect 7260 2267 7294 2278
rect 7295 2267 7306 2283
rect 7352 2274 7368 2290
rect 7375 2288 7405 2340
rect 7439 2336 7440 2343
rect 7424 2328 7440 2336
rect 7411 2296 7424 2315
rect 7439 2296 7469 2312
rect 7411 2280 7485 2296
rect 7411 2278 7424 2280
rect 7439 2278 7473 2280
rect 7076 2256 7089 2258
rect 7104 2256 7138 2258
rect 7076 2240 7138 2256
rect 7182 2251 7198 2254
rect 7260 2251 7290 2262
rect 7338 2258 7384 2274
rect 7411 2262 7485 2278
rect 7338 2256 7372 2258
rect 7337 2240 7384 2256
rect 7411 2240 7424 2262
rect 7439 2240 7469 2262
rect 7496 2240 7497 2256
rect 7512 2240 7525 2400
rect 7555 2296 7568 2400
rect 7613 2378 7614 2388
rect 7629 2378 7642 2388
rect 7613 2374 7642 2378
rect 7647 2374 7677 2400
rect 7695 2386 7711 2388
rect 7783 2386 7836 2400
rect 7784 2384 7848 2386
rect 7891 2384 7906 2400
rect 7955 2397 7985 2400
rect 7955 2394 7991 2397
rect 7921 2386 7937 2388
rect 7695 2374 7710 2378
rect 7613 2372 7710 2374
rect 7738 2372 7906 2384
rect 7922 2374 7937 2378
rect 7955 2375 7994 2394
rect 8013 2388 8020 2389
rect 8019 2381 8020 2388
rect 8003 2378 8004 2381
rect 8019 2378 8032 2381
rect 7955 2374 7985 2375
rect 7994 2374 8000 2375
rect 8003 2374 8032 2378
rect 7922 2373 8032 2374
rect 7922 2372 8038 2373
rect 7597 2364 7648 2372
rect 7597 2352 7622 2364
rect 7629 2352 7648 2364
rect 7679 2364 7729 2372
rect 7679 2356 7695 2364
rect 7702 2362 7729 2364
rect 7738 2362 7959 2372
rect 7702 2352 7959 2362
rect 7988 2364 8038 2372
rect 7988 2355 8004 2364
rect 7597 2344 7648 2352
rect 7695 2344 7959 2352
rect 7985 2352 8004 2355
rect 8011 2352 8038 2364
rect 7985 2344 8038 2352
rect 7613 2336 7614 2344
rect 7629 2336 7642 2344
rect 7613 2328 7629 2336
rect 7610 2321 7629 2324
rect 7610 2312 7632 2321
rect 7583 2302 7632 2312
rect 7583 2296 7613 2302
rect 7632 2297 7637 2302
rect 7555 2280 7629 2296
rect 7647 2288 7677 2344
rect 7712 2334 7920 2344
rect 7955 2340 8000 2344
rect 8003 2343 8004 2344
rect 8019 2343 8032 2344
rect 7738 2304 7927 2334
rect 7753 2301 7927 2304
rect 7746 2298 7927 2301
rect 7555 2278 7568 2280
rect 7583 2278 7617 2280
rect 7555 2262 7629 2278
rect 7656 2274 7669 2288
rect 7684 2274 7700 2290
rect 7746 2285 7757 2298
rect 7539 2240 7540 2256
rect 7555 2240 7568 2262
rect 7583 2240 7613 2262
rect 7656 2258 7718 2274
rect 7746 2267 7757 2283
rect 7762 2278 7772 2298
rect 7782 2278 7796 2298
rect 7799 2285 7808 2298
rect 7824 2285 7833 2298
rect 7762 2267 7796 2278
rect 7799 2267 7808 2283
rect 7824 2267 7833 2283
rect 7840 2278 7850 2298
rect 7860 2278 7874 2298
rect 7875 2285 7886 2298
rect 7840 2267 7874 2278
rect 7875 2267 7886 2283
rect 7932 2274 7948 2290
rect 7955 2288 7985 2340
rect 8019 2336 8020 2343
rect 8004 2328 8020 2336
rect 7991 2296 8004 2315
rect 8019 2296 8049 2312
rect 7991 2280 8065 2296
rect 7991 2278 8004 2280
rect 8019 2278 8053 2280
rect 7656 2256 7669 2258
rect 7684 2256 7718 2258
rect 7656 2240 7718 2256
rect 7762 2251 7778 2254
rect 7840 2251 7870 2262
rect 7918 2258 7964 2274
rect 7991 2262 8065 2278
rect 7918 2256 7952 2258
rect 7917 2240 7964 2256
rect 7991 2240 8004 2262
rect 8019 2240 8049 2262
rect 8076 2240 8077 2256
rect 8092 2240 8105 2400
rect 8135 2296 8148 2400
rect 8193 2378 8194 2388
rect 8209 2378 8222 2388
rect 8193 2374 8222 2378
rect 8227 2374 8257 2400
rect 8275 2386 8291 2388
rect 8363 2386 8416 2400
rect 8364 2384 8428 2386
rect 8471 2384 8486 2400
rect 8535 2397 8565 2400
rect 8535 2394 8571 2397
rect 8501 2386 8517 2388
rect 8275 2374 8290 2378
rect 8193 2372 8290 2374
rect 8318 2372 8486 2384
rect 8502 2374 8517 2378
rect 8535 2375 8574 2394
rect 8593 2388 8600 2389
rect 8599 2381 8600 2388
rect 8583 2378 8584 2381
rect 8599 2378 8612 2381
rect 8535 2374 8565 2375
rect 8574 2374 8580 2375
rect 8583 2374 8612 2378
rect 8502 2373 8612 2374
rect 8502 2372 8618 2373
rect 8177 2364 8228 2372
rect 8177 2352 8202 2364
rect 8209 2352 8228 2364
rect 8259 2364 8309 2372
rect 8259 2356 8275 2364
rect 8282 2362 8309 2364
rect 8318 2362 8539 2372
rect 8282 2352 8539 2362
rect 8568 2364 8618 2372
rect 8568 2355 8584 2364
rect 8177 2344 8228 2352
rect 8275 2344 8539 2352
rect 8565 2352 8584 2355
rect 8591 2352 8618 2364
rect 8565 2344 8618 2352
rect 8193 2336 8194 2344
rect 8209 2336 8222 2344
rect 8193 2328 8209 2336
rect 8190 2321 8209 2324
rect 8190 2312 8212 2321
rect 8163 2302 8212 2312
rect 8163 2296 8193 2302
rect 8212 2297 8217 2302
rect 8135 2280 8209 2296
rect 8227 2288 8257 2344
rect 8292 2334 8500 2344
rect 8535 2340 8580 2344
rect 8583 2343 8584 2344
rect 8599 2343 8612 2344
rect 8318 2304 8507 2334
rect 8333 2301 8507 2304
rect 8326 2298 8507 2301
rect 8135 2278 8148 2280
rect 8163 2278 8197 2280
rect 8135 2262 8209 2278
rect 8236 2274 8249 2288
rect 8264 2274 8280 2290
rect 8326 2285 8337 2298
rect 8119 2240 8120 2256
rect 8135 2240 8148 2262
rect 8163 2240 8193 2262
rect 8236 2258 8298 2274
rect 8326 2267 8337 2283
rect 8342 2278 8352 2298
rect 8362 2278 8376 2298
rect 8379 2285 8388 2298
rect 8404 2285 8413 2298
rect 8342 2267 8376 2278
rect 8379 2267 8388 2283
rect 8404 2267 8413 2283
rect 8420 2278 8430 2298
rect 8440 2278 8454 2298
rect 8455 2285 8466 2298
rect 8420 2267 8454 2278
rect 8455 2267 8466 2283
rect 8512 2274 8528 2290
rect 8535 2288 8565 2340
rect 8599 2336 8600 2343
rect 8584 2328 8600 2336
rect 8571 2296 8584 2315
rect 8599 2296 8629 2312
rect 8571 2280 8645 2296
rect 8571 2278 8584 2280
rect 8599 2278 8633 2280
rect 8236 2256 8249 2258
rect 8264 2256 8298 2258
rect 8236 2240 8298 2256
rect 8342 2251 8358 2254
rect 8420 2251 8450 2262
rect 8498 2258 8544 2274
rect 8571 2262 8645 2278
rect 8498 2256 8532 2258
rect 8497 2240 8544 2256
rect 8571 2240 8584 2262
rect 8599 2240 8629 2262
rect 8656 2240 8657 2256
rect 8672 2240 8685 2400
rect 8715 2296 8728 2400
rect 8773 2378 8774 2388
rect 8789 2378 8802 2388
rect 8773 2374 8802 2378
rect 8807 2374 8837 2400
rect 8855 2386 8871 2388
rect 8943 2386 8996 2400
rect 8944 2384 9008 2386
rect 9051 2384 9066 2400
rect 9115 2397 9145 2400
rect 9115 2394 9151 2397
rect 9081 2386 9097 2388
rect 8855 2374 8870 2378
rect 8773 2372 8870 2374
rect 8898 2372 9066 2384
rect 9082 2374 9097 2378
rect 9115 2375 9154 2394
rect 9173 2388 9180 2389
rect 9179 2381 9180 2388
rect 9163 2378 9164 2381
rect 9179 2378 9192 2381
rect 9115 2374 9145 2375
rect 9154 2374 9160 2375
rect 9163 2374 9192 2378
rect 9082 2373 9192 2374
rect 9082 2372 9198 2373
rect 8757 2364 8808 2372
rect 8757 2352 8782 2364
rect 8789 2352 8808 2364
rect 8839 2364 8889 2372
rect 8839 2356 8855 2364
rect 8862 2362 8889 2364
rect 8898 2362 9119 2372
rect 8862 2352 9119 2362
rect 9148 2364 9198 2372
rect 9148 2355 9164 2364
rect 8757 2344 8808 2352
rect 8855 2344 9119 2352
rect 9145 2352 9164 2355
rect 9171 2352 9198 2364
rect 9145 2344 9198 2352
rect 8773 2336 8774 2344
rect 8789 2336 8802 2344
rect 8773 2328 8789 2336
rect 8770 2321 8789 2324
rect 8770 2312 8792 2321
rect 8743 2302 8792 2312
rect 8743 2296 8773 2302
rect 8792 2297 8797 2302
rect 8715 2280 8789 2296
rect 8807 2288 8837 2344
rect 8872 2334 9080 2344
rect 9115 2340 9160 2344
rect 9163 2343 9164 2344
rect 9179 2343 9192 2344
rect 8898 2304 9087 2334
rect 8913 2301 9087 2304
rect 8906 2298 9087 2301
rect 8715 2278 8728 2280
rect 8743 2278 8777 2280
rect 8715 2262 8789 2278
rect 8816 2274 8829 2288
rect 8844 2274 8860 2290
rect 8906 2285 8917 2298
rect 8699 2240 8700 2256
rect 8715 2240 8728 2262
rect 8743 2240 8773 2262
rect 8816 2258 8878 2274
rect 8906 2267 8917 2283
rect 8922 2278 8932 2298
rect 8942 2278 8956 2298
rect 8959 2285 8968 2298
rect 8984 2285 8993 2298
rect 8922 2267 8956 2278
rect 8959 2267 8968 2283
rect 8984 2267 8993 2283
rect 9000 2278 9010 2298
rect 9020 2278 9034 2298
rect 9035 2285 9046 2298
rect 9000 2267 9034 2278
rect 9035 2267 9046 2283
rect 9092 2274 9108 2290
rect 9115 2288 9145 2340
rect 9179 2336 9180 2343
rect 9164 2328 9180 2336
rect 9151 2296 9164 2315
rect 9179 2296 9209 2312
rect 9151 2280 9225 2296
rect 9151 2278 9164 2280
rect 9179 2278 9213 2280
rect 8816 2256 8829 2258
rect 8844 2256 8878 2258
rect 8816 2240 8878 2256
rect 8922 2251 8938 2254
rect 9000 2251 9030 2262
rect 9078 2258 9124 2274
rect 9151 2262 9225 2278
rect 9078 2256 9112 2258
rect 9077 2240 9124 2256
rect 9151 2240 9164 2262
rect 9179 2240 9209 2262
rect 9236 2240 9237 2256
rect 9252 2240 9265 2400
rect -7 2232 34 2240
rect -7 2206 8 2232
rect 15 2206 34 2232
rect 98 2228 160 2240
rect 172 2228 247 2240
rect 305 2228 380 2240
rect 392 2228 423 2240
rect 429 2228 464 2240
rect 98 2226 260 2228
rect -7 2198 34 2206
rect 116 2202 129 2226
rect 144 2224 159 2226
rect -1 2188 0 2198
rect 15 2188 28 2198
rect 43 2188 73 2202
rect 116 2188 159 2202
rect 183 2199 190 2206
rect 193 2202 260 2226
rect 292 2226 464 2228
rect 262 2204 290 2208
rect 292 2204 372 2226
rect 393 2224 408 2226
rect 262 2202 372 2204
rect 193 2198 372 2202
rect 166 2188 196 2198
rect 198 2188 351 2198
rect 359 2188 389 2198
rect 393 2188 423 2202
rect 451 2188 464 2226
rect 536 2232 571 2240
rect 536 2206 537 2232
rect 544 2206 571 2232
rect 479 2188 509 2202
rect 536 2198 571 2206
rect 573 2232 614 2240
rect 573 2206 588 2232
rect 595 2206 614 2232
rect 678 2228 740 2240
rect 752 2228 827 2240
rect 885 2228 960 2240
rect 972 2228 1003 2240
rect 1009 2228 1044 2240
rect 678 2226 840 2228
rect 573 2198 614 2206
rect 696 2202 709 2226
rect 724 2224 739 2226
rect 536 2188 537 2198
rect 552 2188 565 2198
rect 579 2188 580 2198
rect 595 2188 608 2198
rect 623 2188 653 2202
rect 696 2188 739 2202
rect 763 2199 770 2206
rect 773 2202 840 2226
rect 872 2226 1044 2228
rect 842 2204 870 2208
rect 872 2204 952 2226
rect 973 2224 988 2226
rect 842 2202 952 2204
rect 773 2198 952 2202
rect 746 2188 776 2198
rect 778 2188 931 2198
rect 939 2188 969 2198
rect 973 2188 1003 2202
rect 1031 2188 1044 2226
rect 1116 2232 1151 2240
rect 1116 2206 1117 2232
rect 1124 2206 1151 2232
rect 1059 2188 1089 2202
rect 1116 2198 1151 2206
rect 1153 2232 1194 2240
rect 1153 2206 1168 2232
rect 1175 2206 1194 2232
rect 1258 2228 1320 2240
rect 1332 2228 1407 2240
rect 1465 2228 1540 2240
rect 1552 2228 1583 2240
rect 1589 2228 1624 2240
rect 1258 2226 1420 2228
rect 1153 2198 1194 2206
rect 1276 2202 1289 2226
rect 1304 2224 1319 2226
rect 1116 2188 1117 2198
rect 1132 2188 1145 2198
rect 1159 2188 1160 2198
rect 1175 2188 1188 2198
rect 1203 2188 1233 2202
rect 1276 2188 1319 2202
rect 1343 2199 1350 2206
rect 1353 2202 1420 2226
rect 1452 2226 1624 2228
rect 1422 2204 1450 2208
rect 1452 2204 1532 2226
rect 1553 2224 1568 2226
rect 1422 2202 1532 2204
rect 1353 2198 1532 2202
rect 1326 2188 1356 2198
rect 1358 2188 1511 2198
rect 1519 2188 1549 2198
rect 1553 2188 1583 2202
rect 1611 2188 1624 2226
rect 1696 2232 1731 2240
rect 1696 2206 1697 2232
rect 1704 2206 1731 2232
rect 1639 2188 1669 2202
rect 1696 2198 1731 2206
rect 1733 2232 1774 2240
rect 1733 2206 1748 2232
rect 1755 2206 1774 2232
rect 1838 2228 1900 2240
rect 1912 2228 1987 2240
rect 2045 2228 2120 2240
rect 2132 2228 2163 2240
rect 2169 2228 2204 2240
rect 1838 2226 2000 2228
rect 1733 2198 1774 2206
rect 1856 2202 1869 2226
rect 1884 2224 1899 2226
rect 1696 2188 1697 2198
rect 1712 2188 1725 2198
rect 1739 2188 1740 2198
rect 1755 2188 1768 2198
rect 1783 2188 1813 2202
rect 1856 2188 1899 2202
rect 1923 2199 1930 2206
rect 1933 2202 2000 2226
rect 2032 2226 2204 2228
rect 2002 2204 2030 2208
rect 2032 2204 2112 2226
rect 2133 2224 2148 2226
rect 2002 2202 2112 2204
rect 1933 2198 2112 2202
rect 1906 2188 1936 2198
rect 1938 2188 2091 2198
rect 2099 2188 2129 2198
rect 2133 2188 2163 2202
rect 2191 2188 2204 2226
rect 2276 2232 2311 2240
rect 2276 2206 2277 2232
rect 2284 2206 2311 2232
rect 2219 2188 2249 2202
rect 2276 2198 2311 2206
rect 2313 2232 2354 2240
rect 2313 2206 2328 2232
rect 2335 2206 2354 2232
rect 2418 2228 2480 2240
rect 2492 2228 2567 2240
rect 2625 2228 2700 2240
rect 2712 2228 2743 2240
rect 2749 2228 2784 2240
rect 2418 2226 2580 2228
rect 2313 2198 2354 2206
rect 2436 2202 2449 2226
rect 2464 2224 2479 2226
rect 2276 2188 2277 2198
rect 2292 2188 2305 2198
rect 2319 2188 2320 2198
rect 2335 2188 2348 2198
rect 2363 2188 2393 2202
rect 2436 2188 2479 2202
rect 2503 2199 2510 2206
rect 2513 2202 2580 2226
rect 2612 2226 2784 2228
rect 2582 2204 2610 2208
rect 2612 2204 2692 2226
rect 2713 2224 2728 2226
rect 2582 2202 2692 2204
rect 2513 2198 2692 2202
rect 2486 2188 2516 2198
rect 2518 2188 2671 2198
rect 2679 2188 2709 2198
rect 2713 2188 2743 2202
rect 2771 2188 2784 2226
rect 2856 2232 2891 2240
rect 2856 2206 2857 2232
rect 2864 2206 2891 2232
rect 2799 2188 2829 2202
rect 2856 2198 2891 2206
rect 2893 2232 2934 2240
rect 2893 2206 2908 2232
rect 2915 2206 2934 2232
rect 2998 2228 3060 2240
rect 3072 2228 3147 2240
rect 3205 2228 3280 2240
rect 3292 2228 3323 2240
rect 3329 2228 3364 2240
rect 2998 2226 3160 2228
rect 2893 2198 2934 2206
rect 3016 2202 3029 2226
rect 3044 2224 3059 2226
rect 2856 2188 2857 2198
rect 2872 2188 2885 2198
rect 2899 2188 2900 2198
rect 2915 2188 2928 2198
rect 2943 2188 2973 2202
rect 3016 2188 3059 2202
rect 3083 2199 3090 2206
rect 3093 2202 3160 2226
rect 3192 2226 3364 2228
rect 3162 2204 3190 2208
rect 3192 2204 3272 2226
rect 3293 2224 3308 2226
rect 3162 2202 3272 2204
rect 3093 2198 3272 2202
rect 3066 2188 3096 2198
rect 3098 2188 3251 2198
rect 3259 2188 3289 2198
rect 3293 2188 3323 2202
rect 3351 2188 3364 2226
rect 3436 2232 3471 2240
rect 3436 2206 3437 2232
rect 3444 2206 3471 2232
rect 3379 2188 3409 2202
rect 3436 2198 3471 2206
rect 3473 2232 3514 2240
rect 3473 2206 3488 2232
rect 3495 2206 3514 2232
rect 3578 2228 3640 2240
rect 3652 2228 3727 2240
rect 3785 2228 3860 2240
rect 3872 2228 3903 2240
rect 3909 2228 3944 2240
rect 3578 2226 3740 2228
rect 3473 2198 3514 2206
rect 3596 2202 3609 2226
rect 3624 2224 3639 2226
rect 3436 2188 3437 2198
rect 3452 2188 3465 2198
rect 3479 2188 3480 2198
rect 3495 2188 3508 2198
rect 3523 2188 3553 2202
rect 3596 2188 3639 2202
rect 3663 2199 3670 2206
rect 3673 2202 3740 2226
rect 3772 2226 3944 2228
rect 3742 2204 3770 2208
rect 3772 2204 3852 2226
rect 3873 2224 3888 2226
rect 3742 2202 3852 2204
rect 3673 2198 3852 2202
rect 3646 2188 3676 2198
rect 3678 2188 3831 2198
rect 3839 2188 3869 2198
rect 3873 2188 3903 2202
rect 3931 2188 3944 2226
rect 4016 2232 4051 2240
rect 4016 2206 4017 2232
rect 4024 2206 4051 2232
rect 3959 2188 3989 2202
rect 4016 2198 4051 2206
rect 4053 2232 4094 2240
rect 4053 2206 4068 2232
rect 4075 2206 4094 2232
rect 4158 2228 4220 2240
rect 4232 2228 4307 2240
rect 4365 2228 4440 2240
rect 4452 2228 4483 2240
rect 4489 2228 4524 2240
rect 4158 2226 4320 2228
rect 4053 2198 4094 2206
rect 4176 2202 4189 2226
rect 4204 2224 4219 2226
rect 4016 2188 4017 2198
rect 4032 2188 4045 2198
rect 4059 2188 4060 2198
rect 4075 2188 4088 2198
rect 4103 2188 4133 2202
rect 4176 2188 4219 2202
rect 4243 2199 4250 2206
rect 4253 2202 4320 2226
rect 4352 2226 4524 2228
rect 4322 2204 4350 2208
rect 4352 2204 4432 2226
rect 4453 2224 4468 2226
rect 4322 2202 4432 2204
rect 4253 2198 4432 2202
rect 4226 2188 4256 2198
rect 4258 2188 4411 2198
rect 4419 2188 4449 2198
rect 4453 2188 4483 2202
rect 4511 2188 4524 2226
rect 4596 2232 4631 2240
rect 4596 2206 4597 2232
rect 4604 2206 4631 2232
rect 4539 2188 4569 2202
rect 4596 2198 4631 2206
rect 4633 2232 4674 2240
rect 4633 2206 4648 2232
rect 4655 2206 4674 2232
rect 4738 2228 4800 2240
rect 4812 2228 4887 2240
rect 4945 2228 5020 2240
rect 5032 2228 5063 2240
rect 5069 2228 5104 2240
rect 4738 2226 4900 2228
rect 4633 2198 4674 2206
rect 4756 2202 4769 2226
rect 4784 2224 4799 2226
rect 4596 2188 4597 2198
rect 4612 2188 4625 2198
rect 4639 2188 4640 2198
rect 4655 2188 4668 2198
rect 4683 2188 4713 2202
rect 4756 2188 4799 2202
rect 4823 2199 4830 2206
rect 4833 2202 4900 2226
rect 4932 2226 5104 2228
rect 4902 2204 4930 2208
rect 4932 2204 5012 2226
rect 5033 2224 5048 2226
rect 4902 2202 5012 2204
rect 4833 2198 5012 2202
rect 4806 2188 4836 2198
rect 4838 2188 4991 2198
rect 4999 2188 5029 2198
rect 5033 2188 5063 2202
rect 5091 2188 5104 2226
rect 5176 2232 5211 2240
rect 5176 2206 5177 2232
rect 5184 2206 5211 2232
rect 5119 2188 5149 2202
rect 5176 2198 5211 2206
rect 5213 2232 5254 2240
rect 5213 2206 5228 2232
rect 5235 2206 5254 2232
rect 5318 2228 5380 2240
rect 5392 2228 5467 2240
rect 5525 2228 5600 2240
rect 5612 2228 5643 2240
rect 5649 2228 5684 2240
rect 5318 2226 5480 2228
rect 5213 2198 5254 2206
rect 5336 2202 5349 2226
rect 5364 2224 5379 2226
rect 5176 2188 5177 2198
rect 5192 2188 5205 2198
rect 5219 2188 5220 2198
rect 5235 2188 5248 2198
rect 5263 2188 5293 2202
rect 5336 2188 5379 2202
rect 5403 2199 5410 2206
rect 5413 2202 5480 2226
rect 5512 2226 5684 2228
rect 5482 2204 5510 2208
rect 5512 2204 5592 2226
rect 5613 2224 5628 2226
rect 5482 2202 5592 2204
rect 5413 2198 5592 2202
rect 5386 2188 5416 2198
rect 5418 2188 5571 2198
rect 5579 2188 5609 2198
rect 5613 2188 5643 2202
rect 5671 2188 5684 2226
rect 5756 2232 5791 2240
rect 5756 2206 5757 2232
rect 5764 2206 5791 2232
rect 5699 2188 5729 2202
rect 5756 2198 5791 2206
rect 5793 2232 5834 2240
rect 5793 2206 5808 2232
rect 5815 2206 5834 2232
rect 5898 2228 5960 2240
rect 5972 2228 6047 2240
rect 6105 2228 6180 2240
rect 6192 2228 6223 2240
rect 6229 2228 6264 2240
rect 5898 2226 6060 2228
rect 5793 2198 5834 2206
rect 5916 2202 5929 2226
rect 5944 2224 5959 2226
rect 5756 2188 5757 2198
rect 5772 2188 5785 2198
rect 5799 2188 5800 2198
rect 5815 2188 5828 2198
rect 5843 2188 5873 2202
rect 5916 2188 5959 2202
rect 5983 2199 5990 2206
rect 5993 2202 6060 2226
rect 6092 2226 6264 2228
rect 6062 2204 6090 2208
rect 6092 2204 6172 2226
rect 6193 2224 6208 2226
rect 6062 2202 6172 2204
rect 5993 2198 6172 2202
rect 5966 2188 5996 2198
rect 5998 2188 6151 2198
rect 6159 2188 6189 2198
rect 6193 2188 6223 2202
rect 6251 2188 6264 2226
rect 6336 2232 6371 2240
rect 6336 2206 6337 2232
rect 6344 2206 6371 2232
rect 6279 2188 6309 2202
rect 6336 2198 6371 2206
rect 6373 2232 6414 2240
rect 6373 2206 6388 2232
rect 6395 2206 6414 2232
rect 6478 2228 6540 2240
rect 6552 2228 6627 2240
rect 6685 2228 6760 2240
rect 6772 2228 6803 2240
rect 6809 2228 6844 2240
rect 6478 2226 6640 2228
rect 6373 2198 6414 2206
rect 6496 2202 6509 2226
rect 6524 2224 6539 2226
rect 6336 2188 6337 2198
rect 6352 2188 6365 2198
rect 6379 2188 6380 2198
rect 6395 2188 6408 2198
rect 6423 2188 6453 2202
rect 6496 2188 6539 2202
rect 6563 2199 6570 2206
rect 6573 2202 6640 2226
rect 6672 2226 6844 2228
rect 6642 2204 6670 2208
rect 6672 2204 6752 2226
rect 6773 2224 6788 2226
rect 6642 2202 6752 2204
rect 6573 2198 6752 2202
rect 6546 2188 6576 2198
rect 6578 2188 6731 2198
rect 6739 2188 6769 2198
rect 6773 2188 6803 2202
rect 6831 2188 6844 2226
rect 6916 2232 6951 2240
rect 6916 2206 6917 2232
rect 6924 2206 6951 2232
rect 6859 2188 6889 2202
rect 6916 2198 6951 2206
rect 6953 2232 6994 2240
rect 6953 2206 6968 2232
rect 6975 2206 6994 2232
rect 7058 2228 7120 2240
rect 7132 2228 7207 2240
rect 7265 2228 7340 2240
rect 7352 2228 7383 2240
rect 7389 2228 7424 2240
rect 7058 2226 7220 2228
rect 6953 2198 6994 2206
rect 7076 2202 7089 2226
rect 7104 2224 7119 2226
rect 6916 2188 6917 2198
rect 6932 2188 6945 2198
rect 6959 2188 6960 2198
rect 6975 2188 6988 2198
rect 7003 2188 7033 2202
rect 7076 2188 7119 2202
rect 7143 2199 7150 2206
rect 7153 2202 7220 2226
rect 7252 2226 7424 2228
rect 7222 2204 7250 2208
rect 7252 2204 7332 2226
rect 7353 2224 7368 2226
rect 7222 2202 7332 2204
rect 7153 2198 7332 2202
rect 7126 2188 7156 2198
rect 7158 2188 7311 2198
rect 7319 2188 7349 2198
rect 7353 2188 7383 2202
rect 7411 2188 7424 2226
rect 7496 2232 7531 2240
rect 7496 2206 7497 2232
rect 7504 2206 7531 2232
rect 7439 2188 7469 2202
rect 7496 2198 7531 2206
rect 7533 2232 7574 2240
rect 7533 2206 7548 2232
rect 7555 2206 7574 2232
rect 7638 2228 7700 2240
rect 7712 2228 7787 2240
rect 7845 2228 7920 2240
rect 7932 2228 7963 2240
rect 7969 2228 8004 2240
rect 7638 2226 7800 2228
rect 7533 2198 7574 2206
rect 7656 2202 7669 2226
rect 7684 2224 7699 2226
rect 7496 2188 7497 2198
rect 7512 2188 7525 2198
rect 7539 2188 7540 2198
rect 7555 2188 7568 2198
rect 7583 2188 7613 2202
rect 7656 2188 7699 2202
rect 7723 2199 7730 2206
rect 7733 2202 7800 2226
rect 7832 2226 8004 2228
rect 7802 2204 7830 2208
rect 7832 2204 7912 2226
rect 7933 2224 7948 2226
rect 7802 2202 7912 2204
rect 7733 2198 7912 2202
rect 7706 2188 7736 2198
rect 7738 2188 7891 2198
rect 7899 2188 7929 2198
rect 7933 2188 7963 2202
rect 7991 2188 8004 2226
rect 8076 2232 8111 2240
rect 8076 2206 8077 2232
rect 8084 2206 8111 2232
rect 8019 2188 8049 2202
rect 8076 2198 8111 2206
rect 8113 2232 8154 2240
rect 8113 2206 8128 2232
rect 8135 2206 8154 2232
rect 8218 2228 8280 2240
rect 8292 2228 8367 2240
rect 8425 2228 8500 2240
rect 8512 2228 8543 2240
rect 8549 2228 8584 2240
rect 8218 2226 8380 2228
rect 8113 2198 8154 2206
rect 8236 2202 8249 2226
rect 8264 2224 8279 2226
rect 8076 2188 8077 2198
rect 8092 2188 8105 2198
rect 8119 2188 8120 2198
rect 8135 2188 8148 2198
rect 8163 2188 8193 2202
rect 8236 2188 8279 2202
rect 8303 2199 8310 2206
rect 8313 2202 8380 2226
rect 8412 2226 8584 2228
rect 8382 2204 8410 2208
rect 8412 2204 8492 2226
rect 8513 2224 8528 2226
rect 8382 2202 8492 2204
rect 8313 2198 8492 2202
rect 8286 2188 8316 2198
rect 8318 2188 8471 2198
rect 8479 2188 8509 2198
rect 8513 2188 8543 2202
rect 8571 2188 8584 2226
rect 8656 2232 8691 2240
rect 8656 2206 8657 2232
rect 8664 2206 8691 2232
rect 8599 2188 8629 2202
rect 8656 2198 8691 2206
rect 8693 2232 8734 2240
rect 8693 2206 8708 2232
rect 8715 2206 8734 2232
rect 8798 2228 8860 2240
rect 8872 2228 8947 2240
rect 9005 2228 9080 2240
rect 9092 2228 9123 2240
rect 9129 2228 9164 2240
rect 8798 2226 8960 2228
rect 8693 2198 8734 2206
rect 8816 2202 8829 2226
rect 8844 2224 8859 2226
rect 8656 2188 8657 2198
rect 8672 2188 8685 2198
rect 8699 2188 8700 2198
rect 8715 2188 8728 2198
rect 8743 2188 8773 2202
rect 8816 2188 8859 2202
rect 8883 2199 8890 2206
rect 8893 2202 8960 2226
rect 8992 2226 9164 2228
rect 8962 2204 8990 2208
rect 8992 2204 9072 2226
rect 9093 2224 9108 2226
rect 8962 2202 9072 2204
rect 8893 2198 9072 2202
rect 8866 2188 8896 2198
rect 8898 2188 9051 2198
rect 9059 2188 9089 2198
rect 9093 2188 9123 2202
rect 9151 2188 9164 2226
rect 9236 2232 9271 2240
rect 9236 2206 9237 2232
rect 9244 2206 9271 2232
rect 9179 2188 9209 2202
rect 9236 2198 9271 2206
rect 9236 2188 9237 2198
rect 9252 2188 9265 2198
rect -1 2182 9265 2188
rect 0 2174 9265 2182
rect 15 2144 28 2174
rect 43 2156 73 2174
rect 116 2160 130 2174
rect 166 2160 386 2174
rect 117 2158 130 2160
rect 83 2146 98 2158
rect 80 2144 102 2146
rect 107 2144 137 2158
rect 198 2156 351 2160
rect 180 2144 372 2156
rect 415 2144 445 2158
rect 451 2144 464 2174
rect 479 2156 509 2174
rect 552 2144 565 2174
rect 595 2144 608 2174
rect 623 2156 653 2174
rect 696 2160 710 2174
rect 746 2160 966 2174
rect 697 2158 710 2160
rect 663 2146 678 2158
rect 660 2144 682 2146
rect 687 2144 717 2158
rect 778 2156 931 2160
rect 760 2144 952 2156
rect 995 2144 1025 2158
rect 1031 2144 1044 2174
rect 1059 2156 1089 2174
rect 1132 2144 1145 2174
rect 1175 2144 1188 2174
rect 1203 2156 1233 2174
rect 1276 2160 1290 2174
rect 1326 2160 1546 2174
rect 1277 2158 1290 2160
rect 1243 2146 1258 2158
rect 1240 2144 1262 2146
rect 1267 2144 1297 2158
rect 1358 2156 1511 2160
rect 1340 2144 1532 2156
rect 1575 2144 1605 2158
rect 1611 2144 1624 2174
rect 1639 2156 1669 2174
rect 1712 2144 1725 2174
rect 1755 2144 1768 2174
rect 1783 2156 1813 2174
rect 1856 2160 1870 2174
rect 1906 2160 2126 2174
rect 1857 2158 1870 2160
rect 1823 2146 1838 2158
rect 1820 2144 1842 2146
rect 1847 2144 1877 2158
rect 1938 2156 2091 2160
rect 1920 2144 2112 2156
rect 2155 2144 2185 2158
rect 2191 2144 2204 2174
rect 2219 2156 2249 2174
rect 2292 2144 2305 2174
rect 2335 2144 2348 2174
rect 2363 2156 2393 2174
rect 2436 2160 2450 2174
rect 2486 2160 2706 2174
rect 2437 2158 2450 2160
rect 2403 2146 2418 2158
rect 2400 2144 2422 2146
rect 2427 2144 2457 2158
rect 2518 2156 2671 2160
rect 2500 2144 2692 2156
rect 2735 2144 2765 2158
rect 2771 2144 2784 2174
rect 2799 2156 2829 2174
rect 2872 2144 2885 2174
rect 2915 2144 2928 2174
rect 2943 2156 2973 2174
rect 3016 2160 3030 2174
rect 3066 2160 3286 2174
rect 3017 2158 3030 2160
rect 2983 2146 2998 2158
rect 2980 2144 3002 2146
rect 3007 2144 3037 2158
rect 3098 2156 3251 2160
rect 3080 2144 3272 2156
rect 3315 2144 3345 2158
rect 3351 2144 3364 2174
rect 3379 2156 3409 2174
rect 3452 2144 3465 2174
rect 3495 2144 3508 2174
rect 3523 2156 3553 2174
rect 3596 2160 3610 2174
rect 3646 2160 3866 2174
rect 3597 2158 3610 2160
rect 3563 2146 3578 2158
rect 3560 2144 3582 2146
rect 3587 2144 3617 2158
rect 3678 2156 3831 2160
rect 3660 2144 3852 2156
rect 3895 2144 3925 2158
rect 3931 2144 3944 2174
rect 3959 2156 3989 2174
rect 4032 2144 4045 2174
rect 4075 2144 4088 2174
rect 4103 2156 4133 2174
rect 4176 2160 4190 2174
rect 4226 2160 4446 2174
rect 4177 2158 4190 2160
rect 4143 2146 4158 2158
rect 4140 2144 4162 2146
rect 4167 2144 4197 2158
rect 4258 2156 4411 2160
rect 4240 2144 4432 2156
rect 4475 2144 4505 2158
rect 4511 2144 4524 2174
rect 4539 2156 4569 2174
rect 4612 2144 4625 2174
rect 4655 2144 4668 2174
rect 4683 2156 4713 2174
rect 4756 2160 4770 2174
rect 4806 2160 5026 2174
rect 4757 2158 4770 2160
rect 4723 2146 4738 2158
rect 4720 2144 4742 2146
rect 4747 2144 4777 2158
rect 4838 2156 4991 2160
rect 4820 2144 5012 2156
rect 5055 2144 5085 2158
rect 5091 2144 5104 2174
rect 5119 2156 5149 2174
rect 5192 2144 5205 2174
rect 5235 2144 5248 2174
rect 5263 2156 5293 2174
rect 5336 2160 5350 2174
rect 5386 2160 5606 2174
rect 5337 2158 5350 2160
rect 5303 2146 5318 2158
rect 5300 2144 5322 2146
rect 5327 2144 5357 2158
rect 5418 2156 5571 2160
rect 5400 2144 5592 2156
rect 5635 2144 5665 2158
rect 5671 2144 5684 2174
rect 5699 2156 5729 2174
rect 5772 2144 5785 2174
rect 5815 2144 5828 2174
rect 5843 2156 5873 2174
rect 5916 2160 5930 2174
rect 5966 2160 6186 2174
rect 5917 2158 5930 2160
rect 5883 2146 5898 2158
rect 5880 2144 5902 2146
rect 5907 2144 5937 2158
rect 5998 2156 6151 2160
rect 5980 2144 6172 2156
rect 6215 2144 6245 2158
rect 6251 2144 6264 2174
rect 6279 2156 6309 2174
rect 6352 2144 6365 2174
rect 6395 2144 6408 2174
rect 6423 2156 6453 2174
rect 6496 2160 6510 2174
rect 6546 2160 6766 2174
rect 6497 2158 6510 2160
rect 6463 2146 6478 2158
rect 6460 2144 6482 2146
rect 6487 2144 6517 2158
rect 6578 2156 6731 2160
rect 6560 2144 6752 2156
rect 6795 2144 6825 2158
rect 6831 2144 6844 2174
rect 6859 2156 6889 2174
rect 6932 2144 6945 2174
rect 6975 2144 6988 2174
rect 7003 2156 7033 2174
rect 7076 2160 7090 2174
rect 7126 2160 7346 2174
rect 7077 2158 7090 2160
rect 7043 2146 7058 2158
rect 7040 2144 7062 2146
rect 7067 2144 7097 2158
rect 7158 2156 7311 2160
rect 7140 2144 7332 2156
rect 7375 2144 7405 2158
rect 7411 2144 7424 2174
rect 7439 2156 7469 2174
rect 7512 2144 7525 2174
rect 7555 2144 7568 2174
rect 7583 2156 7613 2174
rect 7656 2160 7670 2174
rect 7706 2160 7926 2174
rect 7657 2158 7670 2160
rect 7623 2146 7638 2158
rect 7620 2144 7642 2146
rect 7647 2144 7677 2158
rect 7738 2156 7891 2160
rect 7720 2144 7912 2156
rect 7955 2144 7985 2158
rect 7991 2144 8004 2174
rect 8019 2156 8049 2174
rect 8092 2144 8105 2174
rect 8135 2144 8148 2174
rect 8163 2156 8193 2174
rect 8236 2160 8250 2174
rect 8286 2160 8506 2174
rect 8237 2158 8250 2160
rect 8203 2146 8218 2158
rect 8200 2144 8222 2146
rect 8227 2144 8257 2158
rect 8318 2156 8471 2160
rect 8300 2144 8492 2156
rect 8535 2144 8565 2158
rect 8571 2144 8584 2174
rect 8599 2156 8629 2174
rect 8672 2144 8685 2174
rect 8715 2144 8728 2174
rect 8743 2156 8773 2174
rect 8816 2160 8830 2174
rect 8866 2160 9086 2174
rect 8817 2158 8830 2160
rect 8783 2146 8798 2158
rect 8780 2144 8802 2146
rect 8807 2144 8837 2158
rect 8898 2156 9051 2160
rect 8880 2144 9072 2156
rect 9115 2144 9145 2158
rect 9151 2144 9164 2174
rect 9179 2156 9209 2174
rect 9252 2144 9265 2174
rect 0 2130 9265 2144
rect 15 2026 28 2130
rect 73 2108 74 2118
rect 89 2108 102 2118
rect 73 2104 102 2108
rect 107 2104 137 2130
rect 155 2116 171 2118
rect 243 2116 296 2130
rect 244 2114 308 2116
rect 351 2114 366 2130
rect 415 2127 445 2130
rect 415 2124 451 2127
rect 381 2116 397 2118
rect 155 2104 170 2108
rect 73 2102 170 2104
rect 198 2102 366 2114
rect 382 2104 397 2108
rect 415 2105 454 2124
rect 473 2118 480 2119
rect 479 2111 480 2118
rect 463 2108 464 2111
rect 479 2108 492 2111
rect 415 2104 445 2105
rect 454 2104 460 2105
rect 463 2104 492 2108
rect 382 2103 492 2104
rect 382 2102 498 2103
rect 57 2094 108 2102
rect 57 2082 82 2094
rect 89 2082 108 2094
rect 139 2094 189 2102
rect 139 2086 155 2094
rect 162 2092 189 2094
rect 198 2092 419 2102
rect 162 2082 419 2092
rect 448 2094 498 2102
rect 448 2085 464 2094
rect 57 2074 108 2082
rect 155 2074 419 2082
rect 445 2082 464 2085
rect 471 2082 498 2094
rect 445 2074 498 2082
rect 73 2066 74 2074
rect 89 2066 102 2074
rect 73 2058 89 2066
rect 70 2051 89 2054
rect 70 2042 92 2051
rect 43 2032 92 2042
rect 43 2026 73 2032
rect 92 2027 97 2032
rect 15 2010 89 2026
rect 107 2018 137 2074
rect 172 2064 380 2074
rect 415 2070 460 2074
rect 463 2073 464 2074
rect 479 2073 492 2074
rect 198 2034 387 2064
rect 213 2031 387 2034
rect 206 2028 387 2031
rect 15 2008 28 2010
rect 43 2008 77 2010
rect 15 1992 89 2008
rect 116 2004 129 2018
rect 144 2004 160 2020
rect 206 2015 217 2028
rect -1 1970 0 1986
rect 15 1970 28 1992
rect 43 1970 73 1992
rect 116 1988 178 2004
rect 206 1997 217 2013
rect 222 2008 232 2028
rect 242 2008 256 2028
rect 259 2015 268 2028
rect 284 2015 293 2028
rect 222 1997 256 2008
rect 259 1997 268 2013
rect 284 1997 293 2013
rect 300 2008 310 2028
rect 320 2008 334 2028
rect 335 2015 346 2028
rect 300 1997 334 2008
rect 335 1997 346 2013
rect 392 2004 408 2020
rect 415 2018 445 2070
rect 479 2066 480 2073
rect 464 2058 480 2066
rect 451 2026 464 2045
rect 479 2026 509 2042
rect 451 2010 525 2026
rect 451 2008 464 2010
rect 479 2008 513 2010
rect 116 1986 129 1988
rect 144 1986 178 1988
rect 116 1970 178 1986
rect 222 1981 238 1984
rect 300 1981 330 1992
rect 378 1988 424 2004
rect 451 1992 525 2008
rect 378 1986 412 1988
rect 377 1970 424 1986
rect 451 1970 464 1992
rect 479 1970 509 1992
rect 536 1970 537 1986
rect 552 1970 565 2130
rect 595 2026 608 2130
rect 653 2108 654 2118
rect 669 2108 682 2118
rect 653 2104 682 2108
rect 687 2104 717 2130
rect 735 2116 751 2118
rect 823 2116 876 2130
rect 824 2114 888 2116
rect 931 2114 946 2130
rect 995 2127 1025 2130
rect 995 2124 1031 2127
rect 961 2116 977 2118
rect 735 2104 750 2108
rect 653 2102 750 2104
rect 778 2102 946 2114
rect 962 2104 977 2108
rect 995 2105 1034 2124
rect 1053 2118 1060 2119
rect 1059 2111 1060 2118
rect 1043 2108 1044 2111
rect 1059 2108 1072 2111
rect 995 2104 1025 2105
rect 1034 2104 1040 2105
rect 1043 2104 1072 2108
rect 962 2103 1072 2104
rect 962 2102 1078 2103
rect 637 2094 688 2102
rect 637 2082 662 2094
rect 669 2082 688 2094
rect 719 2094 769 2102
rect 719 2086 735 2094
rect 742 2092 769 2094
rect 778 2092 999 2102
rect 742 2082 999 2092
rect 1028 2094 1078 2102
rect 1028 2085 1044 2094
rect 637 2074 688 2082
rect 735 2074 999 2082
rect 1025 2082 1044 2085
rect 1051 2082 1078 2094
rect 1025 2074 1078 2082
rect 653 2066 654 2074
rect 669 2066 682 2074
rect 653 2058 669 2066
rect 650 2051 669 2054
rect 650 2042 672 2051
rect 623 2032 672 2042
rect 623 2026 653 2032
rect 672 2027 677 2032
rect 595 2010 669 2026
rect 687 2018 717 2074
rect 752 2064 960 2074
rect 995 2070 1040 2074
rect 1043 2073 1044 2074
rect 1059 2073 1072 2074
rect 778 2034 967 2064
rect 793 2031 967 2034
rect 786 2028 967 2031
rect 595 2008 608 2010
rect 623 2008 657 2010
rect 595 1992 669 2008
rect 696 2004 709 2018
rect 724 2004 740 2020
rect 786 2015 797 2028
rect 579 1970 580 1986
rect 595 1970 608 1992
rect 623 1970 653 1992
rect 696 1988 758 2004
rect 786 1997 797 2013
rect 802 2008 812 2028
rect 822 2008 836 2028
rect 839 2015 848 2028
rect 864 2015 873 2028
rect 802 1997 836 2008
rect 839 1997 848 2013
rect 864 1997 873 2013
rect 880 2008 890 2028
rect 900 2008 914 2028
rect 915 2015 926 2028
rect 880 1997 914 2008
rect 915 1997 926 2013
rect 972 2004 988 2020
rect 995 2018 1025 2070
rect 1059 2066 1060 2073
rect 1044 2058 1060 2066
rect 1031 2026 1044 2045
rect 1059 2026 1089 2042
rect 1031 2010 1105 2026
rect 1031 2008 1044 2010
rect 1059 2008 1093 2010
rect 696 1986 709 1988
rect 724 1986 758 1988
rect 696 1970 758 1986
rect 802 1981 818 1984
rect 880 1981 910 1992
rect 958 1988 1004 2004
rect 1031 1992 1105 2008
rect 958 1986 992 1988
rect 957 1970 1004 1986
rect 1031 1970 1044 1992
rect 1059 1970 1089 1992
rect 1116 1970 1117 1986
rect 1132 1970 1145 2130
rect 1175 2026 1188 2130
rect 1233 2108 1234 2118
rect 1249 2108 1262 2118
rect 1233 2104 1262 2108
rect 1267 2104 1297 2130
rect 1315 2116 1331 2118
rect 1403 2116 1456 2130
rect 1404 2114 1468 2116
rect 1511 2114 1526 2130
rect 1575 2127 1605 2130
rect 1575 2124 1611 2127
rect 1541 2116 1557 2118
rect 1315 2104 1330 2108
rect 1233 2102 1330 2104
rect 1358 2102 1526 2114
rect 1542 2104 1557 2108
rect 1575 2105 1614 2124
rect 1633 2118 1640 2119
rect 1639 2111 1640 2118
rect 1623 2108 1624 2111
rect 1639 2108 1652 2111
rect 1575 2104 1605 2105
rect 1614 2104 1620 2105
rect 1623 2104 1652 2108
rect 1542 2103 1652 2104
rect 1542 2102 1658 2103
rect 1217 2094 1268 2102
rect 1217 2082 1242 2094
rect 1249 2082 1268 2094
rect 1299 2094 1349 2102
rect 1299 2086 1315 2094
rect 1322 2092 1349 2094
rect 1358 2092 1579 2102
rect 1322 2082 1579 2092
rect 1608 2094 1658 2102
rect 1608 2085 1624 2094
rect 1217 2074 1268 2082
rect 1315 2074 1579 2082
rect 1605 2082 1624 2085
rect 1631 2082 1658 2094
rect 1605 2074 1658 2082
rect 1233 2066 1234 2074
rect 1249 2066 1262 2074
rect 1233 2058 1249 2066
rect 1230 2051 1249 2054
rect 1230 2042 1252 2051
rect 1203 2032 1252 2042
rect 1203 2026 1233 2032
rect 1252 2027 1257 2032
rect 1175 2010 1249 2026
rect 1267 2018 1297 2074
rect 1332 2064 1540 2074
rect 1575 2070 1620 2074
rect 1623 2073 1624 2074
rect 1639 2073 1652 2074
rect 1358 2034 1547 2064
rect 1373 2031 1547 2034
rect 1366 2028 1547 2031
rect 1175 2008 1188 2010
rect 1203 2008 1237 2010
rect 1175 1992 1249 2008
rect 1276 2004 1289 2018
rect 1304 2004 1320 2020
rect 1366 2015 1377 2028
rect 1159 1970 1160 1986
rect 1175 1970 1188 1992
rect 1203 1970 1233 1992
rect 1276 1988 1338 2004
rect 1366 1997 1377 2013
rect 1382 2008 1392 2028
rect 1402 2008 1416 2028
rect 1419 2015 1428 2028
rect 1444 2015 1453 2028
rect 1382 1997 1416 2008
rect 1419 1997 1428 2013
rect 1444 1997 1453 2013
rect 1460 2008 1470 2028
rect 1480 2008 1494 2028
rect 1495 2015 1506 2028
rect 1460 1997 1494 2008
rect 1495 1997 1506 2013
rect 1552 2004 1568 2020
rect 1575 2018 1605 2070
rect 1639 2066 1640 2073
rect 1624 2058 1640 2066
rect 1611 2026 1624 2045
rect 1639 2026 1669 2042
rect 1611 2010 1685 2026
rect 1611 2008 1624 2010
rect 1639 2008 1673 2010
rect 1276 1986 1289 1988
rect 1304 1986 1338 1988
rect 1276 1970 1338 1986
rect 1382 1981 1398 1984
rect 1460 1981 1490 1992
rect 1538 1988 1584 2004
rect 1611 1992 1685 2008
rect 1538 1986 1572 1988
rect 1537 1970 1584 1986
rect 1611 1970 1624 1992
rect 1639 1970 1669 1992
rect 1696 1970 1697 1986
rect 1712 1970 1725 2130
rect 1755 2026 1768 2130
rect 1813 2108 1814 2118
rect 1829 2108 1842 2118
rect 1813 2104 1842 2108
rect 1847 2104 1877 2130
rect 1895 2116 1911 2118
rect 1983 2116 2036 2130
rect 1984 2114 2048 2116
rect 2091 2114 2106 2130
rect 2155 2127 2185 2130
rect 2155 2124 2191 2127
rect 2121 2116 2137 2118
rect 1895 2104 1910 2108
rect 1813 2102 1910 2104
rect 1938 2102 2106 2114
rect 2122 2104 2137 2108
rect 2155 2105 2194 2124
rect 2213 2118 2220 2119
rect 2219 2111 2220 2118
rect 2203 2108 2204 2111
rect 2219 2108 2232 2111
rect 2155 2104 2185 2105
rect 2194 2104 2200 2105
rect 2203 2104 2232 2108
rect 2122 2103 2232 2104
rect 2122 2102 2238 2103
rect 1797 2094 1848 2102
rect 1797 2082 1822 2094
rect 1829 2082 1848 2094
rect 1879 2094 1929 2102
rect 1879 2086 1895 2094
rect 1902 2092 1929 2094
rect 1938 2092 2159 2102
rect 1902 2082 2159 2092
rect 2188 2094 2238 2102
rect 2188 2085 2204 2094
rect 1797 2074 1848 2082
rect 1895 2074 2159 2082
rect 2185 2082 2204 2085
rect 2211 2082 2238 2094
rect 2185 2074 2238 2082
rect 1813 2066 1814 2074
rect 1829 2066 1842 2074
rect 1813 2058 1829 2066
rect 1810 2051 1829 2054
rect 1810 2042 1832 2051
rect 1783 2032 1832 2042
rect 1783 2026 1813 2032
rect 1832 2027 1837 2032
rect 1755 2010 1829 2026
rect 1847 2018 1877 2074
rect 1912 2064 2120 2074
rect 2155 2070 2200 2074
rect 2203 2073 2204 2074
rect 2219 2073 2232 2074
rect 1938 2034 2127 2064
rect 1953 2031 2127 2034
rect 1946 2028 2127 2031
rect 1755 2008 1768 2010
rect 1783 2008 1817 2010
rect 1755 1992 1829 2008
rect 1856 2004 1869 2018
rect 1884 2004 1900 2020
rect 1946 2015 1957 2028
rect 1739 1970 1740 1986
rect 1755 1970 1768 1992
rect 1783 1970 1813 1992
rect 1856 1988 1918 2004
rect 1946 1997 1957 2013
rect 1962 2008 1972 2028
rect 1982 2008 1996 2028
rect 1999 2015 2008 2028
rect 2024 2015 2033 2028
rect 1962 1997 1996 2008
rect 1999 1997 2008 2013
rect 2024 1997 2033 2013
rect 2040 2008 2050 2028
rect 2060 2008 2074 2028
rect 2075 2015 2086 2028
rect 2040 1997 2074 2008
rect 2075 1997 2086 2013
rect 2132 2004 2148 2020
rect 2155 2018 2185 2070
rect 2219 2066 2220 2073
rect 2204 2058 2220 2066
rect 2191 2026 2204 2045
rect 2219 2026 2249 2042
rect 2191 2010 2265 2026
rect 2191 2008 2204 2010
rect 2219 2008 2253 2010
rect 1856 1986 1869 1988
rect 1884 1986 1918 1988
rect 1856 1970 1918 1986
rect 1962 1981 1976 1984
rect 2040 1981 2070 1992
rect 2118 1988 2164 2004
rect 2191 1992 2265 2008
rect 2118 1986 2152 1988
rect 2117 1970 2164 1986
rect 2191 1970 2204 1992
rect 2219 1970 2249 1992
rect 2276 1970 2277 1986
rect 2292 1970 2305 2130
rect 2335 2026 2348 2130
rect 2393 2108 2394 2118
rect 2409 2108 2422 2118
rect 2393 2104 2422 2108
rect 2427 2104 2457 2130
rect 2475 2116 2491 2118
rect 2563 2116 2616 2130
rect 2564 2114 2628 2116
rect 2671 2114 2686 2130
rect 2735 2127 2765 2130
rect 2735 2124 2771 2127
rect 2701 2116 2717 2118
rect 2475 2104 2490 2108
rect 2393 2102 2490 2104
rect 2518 2102 2686 2114
rect 2702 2104 2717 2108
rect 2735 2105 2774 2124
rect 2793 2118 2800 2119
rect 2799 2111 2800 2118
rect 2783 2108 2784 2111
rect 2799 2108 2812 2111
rect 2735 2104 2765 2105
rect 2774 2104 2780 2105
rect 2783 2104 2812 2108
rect 2702 2103 2812 2104
rect 2702 2102 2818 2103
rect 2377 2094 2428 2102
rect 2377 2082 2402 2094
rect 2409 2082 2428 2094
rect 2459 2094 2509 2102
rect 2459 2086 2475 2094
rect 2482 2092 2509 2094
rect 2518 2092 2739 2102
rect 2482 2082 2739 2092
rect 2768 2094 2818 2102
rect 2768 2085 2784 2094
rect 2377 2074 2428 2082
rect 2475 2074 2739 2082
rect 2765 2082 2784 2085
rect 2791 2082 2818 2094
rect 2765 2074 2818 2082
rect 2393 2066 2394 2074
rect 2409 2066 2422 2074
rect 2393 2058 2409 2066
rect 2390 2051 2409 2054
rect 2390 2042 2412 2051
rect 2363 2032 2412 2042
rect 2363 2026 2393 2032
rect 2412 2027 2417 2032
rect 2335 2010 2409 2026
rect 2427 2018 2457 2074
rect 2492 2064 2700 2074
rect 2735 2070 2780 2074
rect 2783 2073 2784 2074
rect 2799 2073 2812 2074
rect 2518 2034 2707 2064
rect 2533 2031 2707 2034
rect 2526 2028 2707 2031
rect 2335 2008 2348 2010
rect 2363 2008 2397 2010
rect 2335 1992 2409 2008
rect 2436 2004 2449 2018
rect 2464 2004 2480 2020
rect 2526 2015 2537 2028
rect 2319 1970 2320 1986
rect 2335 1970 2348 1992
rect 2363 1970 2393 1992
rect 2436 1988 2498 2004
rect 2526 1997 2537 2013
rect 2542 2008 2552 2028
rect 2562 2008 2576 2028
rect 2579 2015 2588 2028
rect 2604 2015 2613 2028
rect 2542 1997 2576 2008
rect 2579 1997 2588 2013
rect 2604 1997 2613 2013
rect 2620 2008 2630 2028
rect 2640 2008 2654 2028
rect 2655 2015 2666 2028
rect 2620 1997 2654 2008
rect 2655 1997 2666 2013
rect 2712 2004 2728 2020
rect 2735 2018 2765 2070
rect 2799 2066 2800 2073
rect 2784 2058 2800 2066
rect 2771 2026 2784 2045
rect 2799 2026 2829 2042
rect 2771 2010 2845 2026
rect 2771 2008 2784 2010
rect 2799 2008 2833 2010
rect 2436 1986 2449 1988
rect 2464 1986 2498 1988
rect 2436 1970 2498 1986
rect 2542 1981 2558 1984
rect 2620 1981 2650 1992
rect 2698 1988 2744 2004
rect 2771 1992 2845 2008
rect 2698 1986 2732 1988
rect 2697 1970 2744 1986
rect 2771 1970 2784 1992
rect 2799 1970 2829 1992
rect 2856 1970 2857 1986
rect 2872 1970 2885 2130
rect 2915 2026 2928 2130
rect 2973 2108 2974 2118
rect 2989 2108 3002 2118
rect 2973 2104 3002 2108
rect 3007 2104 3037 2130
rect 3055 2116 3071 2118
rect 3143 2116 3196 2130
rect 3144 2114 3208 2116
rect 3251 2114 3266 2130
rect 3315 2127 3345 2130
rect 3315 2124 3351 2127
rect 3281 2116 3297 2118
rect 3055 2104 3070 2108
rect 2973 2102 3070 2104
rect 3098 2102 3266 2114
rect 3282 2104 3297 2108
rect 3315 2105 3354 2124
rect 3373 2118 3380 2119
rect 3379 2111 3380 2118
rect 3363 2108 3364 2111
rect 3379 2108 3392 2111
rect 3315 2104 3345 2105
rect 3354 2104 3360 2105
rect 3363 2104 3392 2108
rect 3282 2103 3392 2104
rect 3282 2102 3398 2103
rect 2957 2094 3008 2102
rect 2957 2082 2982 2094
rect 2989 2082 3008 2094
rect 3039 2094 3089 2102
rect 3039 2086 3055 2094
rect 3062 2092 3089 2094
rect 3098 2092 3319 2102
rect 3062 2082 3319 2092
rect 3348 2094 3398 2102
rect 3348 2085 3364 2094
rect 2957 2074 3008 2082
rect 3055 2074 3319 2082
rect 3345 2082 3364 2085
rect 3371 2082 3398 2094
rect 3345 2074 3398 2082
rect 2973 2066 2974 2074
rect 2989 2066 3002 2074
rect 2973 2058 2989 2066
rect 2970 2051 2989 2054
rect 2970 2042 2992 2051
rect 2943 2032 2992 2042
rect 2943 2026 2973 2032
rect 2992 2027 2997 2032
rect 2915 2010 2989 2026
rect 3007 2018 3037 2074
rect 3072 2064 3280 2074
rect 3315 2070 3360 2074
rect 3363 2073 3364 2074
rect 3379 2073 3392 2074
rect 3098 2034 3287 2064
rect 3113 2031 3287 2034
rect 3106 2028 3287 2031
rect 2915 2008 2928 2010
rect 2943 2008 2977 2010
rect 2915 1992 2989 2008
rect 3016 2004 3029 2018
rect 3044 2004 3060 2020
rect 3106 2015 3117 2028
rect 2899 1970 2900 1986
rect 2915 1970 2928 1992
rect 2943 1970 2973 1992
rect 3016 1988 3078 2004
rect 3106 1997 3117 2013
rect 3122 2008 3132 2028
rect 3142 2008 3156 2028
rect 3159 2015 3168 2028
rect 3184 2015 3193 2028
rect 3122 1997 3156 2008
rect 3159 1997 3168 2013
rect 3184 1997 3193 2013
rect 3200 2008 3210 2028
rect 3220 2008 3234 2028
rect 3235 2015 3246 2028
rect 3200 1997 3234 2008
rect 3235 1997 3246 2013
rect 3292 2004 3308 2020
rect 3315 2018 3345 2070
rect 3379 2066 3380 2073
rect 3364 2058 3380 2066
rect 3351 2026 3364 2045
rect 3379 2026 3409 2042
rect 3351 2010 3425 2026
rect 3351 2008 3364 2010
rect 3379 2008 3413 2010
rect 3016 1986 3029 1988
rect 3044 1986 3078 1988
rect 3016 1970 3078 1986
rect 3122 1981 3138 1984
rect 3200 1981 3230 1992
rect 3278 1988 3324 2004
rect 3351 1992 3425 2008
rect 3278 1986 3312 1988
rect 3277 1970 3324 1986
rect 3351 1970 3364 1992
rect 3379 1970 3409 1992
rect 3436 1970 3437 1986
rect 3452 1970 3465 2130
rect 3495 2026 3508 2130
rect 3553 2108 3554 2118
rect 3569 2108 3582 2118
rect 3553 2104 3582 2108
rect 3587 2104 3617 2130
rect 3635 2116 3651 2118
rect 3723 2116 3776 2130
rect 3724 2114 3788 2116
rect 3831 2114 3846 2130
rect 3895 2127 3925 2130
rect 3895 2124 3931 2127
rect 3861 2116 3877 2118
rect 3635 2104 3650 2108
rect 3553 2102 3650 2104
rect 3678 2102 3846 2114
rect 3862 2104 3877 2108
rect 3895 2105 3934 2124
rect 3953 2118 3960 2119
rect 3959 2111 3960 2118
rect 3943 2108 3944 2111
rect 3959 2108 3972 2111
rect 3895 2104 3925 2105
rect 3934 2104 3940 2105
rect 3943 2104 3972 2108
rect 3862 2103 3972 2104
rect 3862 2102 3978 2103
rect 3537 2094 3588 2102
rect 3537 2082 3562 2094
rect 3569 2082 3588 2094
rect 3619 2094 3669 2102
rect 3619 2086 3635 2094
rect 3642 2092 3669 2094
rect 3678 2092 3899 2102
rect 3642 2082 3899 2092
rect 3928 2094 3978 2102
rect 3928 2085 3944 2094
rect 3537 2074 3588 2082
rect 3635 2074 3899 2082
rect 3925 2082 3944 2085
rect 3951 2082 3978 2094
rect 3925 2074 3978 2082
rect 3553 2066 3554 2074
rect 3569 2066 3582 2074
rect 3553 2058 3569 2066
rect 3550 2051 3569 2054
rect 3550 2042 3572 2051
rect 3523 2032 3572 2042
rect 3523 2026 3553 2032
rect 3572 2027 3577 2032
rect 3495 2010 3569 2026
rect 3587 2018 3617 2074
rect 3652 2064 3860 2074
rect 3895 2070 3940 2074
rect 3943 2073 3944 2074
rect 3959 2073 3972 2074
rect 3678 2034 3867 2064
rect 3693 2031 3867 2034
rect 3686 2028 3867 2031
rect 3495 2008 3508 2010
rect 3523 2008 3557 2010
rect 3495 1992 3569 2008
rect 3596 2004 3609 2018
rect 3624 2004 3640 2020
rect 3686 2015 3697 2028
rect 3479 1970 3480 1986
rect 3495 1970 3508 1992
rect 3523 1970 3553 1992
rect 3596 1988 3658 2004
rect 3686 1997 3697 2013
rect 3702 2008 3712 2028
rect 3722 2008 3736 2028
rect 3739 2015 3748 2028
rect 3764 2015 3773 2028
rect 3702 1997 3736 2008
rect 3739 1997 3748 2013
rect 3764 1997 3773 2013
rect 3780 2008 3790 2028
rect 3800 2008 3814 2028
rect 3815 2015 3826 2028
rect 3780 1997 3814 2008
rect 3815 1997 3826 2013
rect 3872 2004 3888 2020
rect 3895 2018 3925 2070
rect 3959 2066 3960 2073
rect 3944 2058 3960 2066
rect 3931 2026 3944 2045
rect 3959 2026 3989 2042
rect 3931 2010 4005 2026
rect 3931 2008 3944 2010
rect 3959 2008 3993 2010
rect 3596 1986 3609 1988
rect 3624 1986 3658 1988
rect 3596 1970 3658 1986
rect 3702 1981 3718 1984
rect 3780 1981 3810 1992
rect 3858 1988 3904 2004
rect 3931 1992 4005 2008
rect 3858 1986 3892 1988
rect 3857 1970 3904 1986
rect 3931 1970 3944 1992
rect 3959 1970 3989 1992
rect 4016 1970 4017 1986
rect 4032 1970 4045 2130
rect 4075 2026 4088 2130
rect 4133 2108 4134 2118
rect 4149 2108 4162 2118
rect 4133 2104 4162 2108
rect 4167 2104 4197 2130
rect 4215 2116 4231 2118
rect 4303 2116 4356 2130
rect 4304 2114 4368 2116
rect 4411 2114 4426 2130
rect 4475 2127 4505 2130
rect 4475 2124 4511 2127
rect 4441 2116 4457 2118
rect 4215 2104 4230 2108
rect 4133 2102 4230 2104
rect 4258 2102 4426 2114
rect 4442 2104 4457 2108
rect 4475 2105 4514 2124
rect 4533 2118 4540 2119
rect 4539 2111 4540 2118
rect 4523 2108 4524 2111
rect 4539 2108 4552 2111
rect 4475 2104 4505 2105
rect 4514 2104 4520 2105
rect 4523 2104 4552 2108
rect 4442 2103 4552 2104
rect 4442 2102 4558 2103
rect 4117 2094 4168 2102
rect 4117 2082 4142 2094
rect 4149 2082 4168 2094
rect 4199 2094 4249 2102
rect 4199 2086 4215 2094
rect 4222 2092 4249 2094
rect 4258 2092 4479 2102
rect 4222 2082 4479 2092
rect 4508 2094 4558 2102
rect 4508 2085 4524 2094
rect 4117 2074 4168 2082
rect 4215 2074 4479 2082
rect 4505 2082 4524 2085
rect 4531 2082 4558 2094
rect 4505 2074 4558 2082
rect 4133 2066 4134 2074
rect 4149 2066 4162 2074
rect 4133 2058 4149 2066
rect 4130 2051 4149 2054
rect 4130 2042 4152 2051
rect 4103 2032 4152 2042
rect 4103 2026 4133 2032
rect 4152 2027 4157 2032
rect 4075 2010 4149 2026
rect 4167 2018 4197 2074
rect 4232 2064 4440 2074
rect 4475 2070 4520 2074
rect 4523 2073 4524 2074
rect 4539 2073 4552 2074
rect 4258 2034 4447 2064
rect 4273 2031 4447 2034
rect 4266 2028 4447 2031
rect 4075 2008 4088 2010
rect 4103 2008 4137 2010
rect 4075 1992 4149 2008
rect 4176 2004 4189 2018
rect 4204 2004 4220 2020
rect 4266 2015 4277 2028
rect 4059 1970 4060 1986
rect 4075 1970 4088 1992
rect 4103 1970 4133 1992
rect 4176 1988 4238 2004
rect 4266 1997 4277 2013
rect 4282 2008 4292 2028
rect 4302 2008 4316 2028
rect 4319 2015 4328 2028
rect 4344 2015 4353 2028
rect 4282 1997 4316 2008
rect 4319 1997 4328 2013
rect 4344 1997 4353 2013
rect 4360 2008 4370 2028
rect 4380 2008 4394 2028
rect 4395 2015 4406 2028
rect 4360 1997 4394 2008
rect 4395 1997 4406 2013
rect 4452 2004 4468 2020
rect 4475 2018 4505 2070
rect 4539 2066 4540 2073
rect 4524 2058 4540 2066
rect 4511 2026 4524 2045
rect 4539 2026 4569 2042
rect 4511 2010 4585 2026
rect 4511 2008 4524 2010
rect 4539 2008 4573 2010
rect 4176 1986 4189 1988
rect 4204 1986 4238 1988
rect 4176 1970 4238 1986
rect 4282 1981 4298 1984
rect 4360 1981 4390 1992
rect 4438 1988 4484 2004
rect 4511 1992 4585 2008
rect 4438 1986 4472 1988
rect 4437 1970 4484 1986
rect 4511 1970 4524 1992
rect 4539 1970 4569 1992
rect 4596 1970 4597 1986
rect 4612 1970 4625 2130
rect 4655 2026 4668 2130
rect 4713 2108 4714 2118
rect 4729 2108 4742 2118
rect 4713 2104 4742 2108
rect 4747 2104 4777 2130
rect 4795 2116 4811 2118
rect 4883 2116 4936 2130
rect 4884 2114 4948 2116
rect 4991 2114 5006 2130
rect 5055 2127 5085 2130
rect 5055 2124 5091 2127
rect 5021 2116 5037 2118
rect 4795 2104 4810 2108
rect 4713 2102 4810 2104
rect 4838 2102 5006 2114
rect 5022 2104 5037 2108
rect 5055 2105 5094 2124
rect 5113 2118 5120 2119
rect 5119 2111 5120 2118
rect 5103 2108 5104 2111
rect 5119 2108 5132 2111
rect 5055 2104 5085 2105
rect 5094 2104 5100 2105
rect 5103 2104 5132 2108
rect 5022 2103 5132 2104
rect 5022 2102 5138 2103
rect 4697 2094 4748 2102
rect 4697 2082 4722 2094
rect 4729 2082 4748 2094
rect 4779 2094 4829 2102
rect 4779 2086 4795 2094
rect 4802 2092 4829 2094
rect 4838 2092 5059 2102
rect 4802 2082 5059 2092
rect 5088 2094 5138 2102
rect 5088 2085 5104 2094
rect 4697 2074 4748 2082
rect 4795 2074 5059 2082
rect 5085 2082 5104 2085
rect 5111 2082 5138 2094
rect 5085 2074 5138 2082
rect 4713 2066 4714 2074
rect 4729 2066 4742 2074
rect 4713 2058 4729 2066
rect 4710 2051 4729 2054
rect 4710 2042 4732 2051
rect 4683 2032 4732 2042
rect 4683 2026 4713 2032
rect 4732 2027 4737 2032
rect 4655 2010 4729 2026
rect 4747 2018 4777 2074
rect 4812 2064 5020 2074
rect 5055 2070 5100 2074
rect 5103 2073 5104 2074
rect 5119 2073 5132 2074
rect 4838 2034 5027 2064
rect 4853 2031 5027 2034
rect 4846 2028 5027 2031
rect 4655 2008 4668 2010
rect 4683 2008 4717 2010
rect 4655 1992 4729 2008
rect 4756 2004 4769 2018
rect 4784 2004 4800 2020
rect 4846 2015 4857 2028
rect 4639 1970 4640 1986
rect 4655 1970 4668 1992
rect 4683 1970 4713 1992
rect 4756 1988 4818 2004
rect 4846 1997 4857 2013
rect 4862 2008 4872 2028
rect 4882 2008 4896 2028
rect 4899 2015 4908 2028
rect 4924 2015 4933 2028
rect 4862 1997 4896 2008
rect 4899 1997 4908 2013
rect 4924 1997 4933 2013
rect 4940 2008 4950 2028
rect 4960 2008 4974 2028
rect 4975 2015 4986 2028
rect 4940 1997 4974 2008
rect 4975 1997 4986 2013
rect 5032 2004 5048 2020
rect 5055 2018 5085 2070
rect 5119 2066 5120 2073
rect 5104 2058 5120 2066
rect 5091 2026 5104 2045
rect 5119 2026 5149 2042
rect 5091 2010 5165 2026
rect 5091 2008 5104 2010
rect 5119 2008 5153 2010
rect 4756 1986 4769 1988
rect 4784 1986 4818 1988
rect 4756 1970 4818 1986
rect 4862 1981 4878 1984
rect 4940 1981 4970 1992
rect 5018 1988 5064 2004
rect 5091 1992 5165 2008
rect 5018 1986 5052 1988
rect 5017 1970 5064 1986
rect 5091 1970 5104 1992
rect 5119 1970 5149 1992
rect 5176 1970 5177 1986
rect 5192 1970 5205 2130
rect 5235 2026 5248 2130
rect 5293 2108 5294 2118
rect 5309 2108 5322 2118
rect 5293 2104 5322 2108
rect 5327 2104 5357 2130
rect 5375 2116 5391 2118
rect 5463 2116 5516 2130
rect 5464 2114 5528 2116
rect 5571 2114 5586 2130
rect 5635 2127 5665 2130
rect 5635 2124 5671 2127
rect 5601 2116 5617 2118
rect 5375 2104 5390 2108
rect 5293 2102 5390 2104
rect 5418 2102 5586 2114
rect 5602 2104 5617 2108
rect 5635 2105 5674 2124
rect 5693 2118 5700 2119
rect 5699 2111 5700 2118
rect 5683 2108 5684 2111
rect 5699 2108 5712 2111
rect 5635 2104 5665 2105
rect 5674 2104 5680 2105
rect 5683 2104 5712 2108
rect 5602 2103 5712 2104
rect 5602 2102 5718 2103
rect 5277 2094 5328 2102
rect 5277 2082 5302 2094
rect 5309 2082 5328 2094
rect 5359 2094 5409 2102
rect 5359 2086 5375 2094
rect 5382 2092 5409 2094
rect 5418 2092 5639 2102
rect 5382 2082 5639 2092
rect 5668 2094 5718 2102
rect 5668 2085 5684 2094
rect 5277 2074 5328 2082
rect 5375 2074 5639 2082
rect 5665 2082 5684 2085
rect 5691 2082 5718 2094
rect 5665 2074 5718 2082
rect 5293 2066 5294 2074
rect 5309 2066 5322 2074
rect 5293 2058 5309 2066
rect 5290 2051 5309 2054
rect 5290 2042 5312 2051
rect 5263 2032 5312 2042
rect 5263 2026 5293 2032
rect 5312 2027 5317 2032
rect 5235 2010 5309 2026
rect 5327 2018 5357 2074
rect 5392 2064 5600 2074
rect 5635 2070 5680 2074
rect 5683 2073 5684 2074
rect 5699 2073 5712 2074
rect 5418 2034 5607 2064
rect 5433 2031 5607 2034
rect 5426 2028 5607 2031
rect 5235 2008 5248 2010
rect 5263 2008 5297 2010
rect 5235 1992 5309 2008
rect 5336 2004 5349 2018
rect 5364 2004 5380 2020
rect 5426 2015 5437 2028
rect 5219 1970 5220 1986
rect 5235 1970 5248 1992
rect 5263 1970 5293 1992
rect 5336 1988 5398 2004
rect 5426 1997 5437 2013
rect 5442 2008 5452 2028
rect 5462 2008 5476 2028
rect 5479 2015 5488 2028
rect 5504 2015 5513 2028
rect 5442 1997 5476 2008
rect 5479 1997 5488 2013
rect 5504 1997 5513 2013
rect 5520 2008 5530 2028
rect 5540 2008 5554 2028
rect 5555 2015 5566 2028
rect 5520 1997 5554 2008
rect 5555 1997 5566 2013
rect 5612 2004 5628 2020
rect 5635 2018 5665 2070
rect 5699 2066 5700 2073
rect 5684 2058 5700 2066
rect 5671 2026 5684 2045
rect 5699 2026 5729 2042
rect 5671 2010 5745 2026
rect 5671 2008 5684 2010
rect 5699 2008 5733 2010
rect 5336 1986 5349 1988
rect 5364 1986 5398 1988
rect 5336 1970 5398 1986
rect 5442 1981 5458 1984
rect 5520 1981 5550 1992
rect 5598 1988 5644 2004
rect 5671 1992 5745 2008
rect 5598 1986 5632 1988
rect 5597 1970 5644 1986
rect 5671 1970 5684 1992
rect 5699 1970 5729 1992
rect 5756 1970 5757 1986
rect 5772 1970 5785 2130
rect 5815 2026 5828 2130
rect 5873 2108 5874 2118
rect 5889 2108 5902 2118
rect 5873 2104 5902 2108
rect 5907 2104 5937 2130
rect 5955 2116 5971 2118
rect 6043 2116 6096 2130
rect 6044 2114 6108 2116
rect 6151 2114 6166 2130
rect 6215 2127 6245 2130
rect 6215 2124 6251 2127
rect 6181 2116 6197 2118
rect 5955 2104 5970 2108
rect 5873 2102 5970 2104
rect 5998 2102 6166 2114
rect 6182 2104 6197 2108
rect 6215 2105 6254 2124
rect 6273 2118 6280 2119
rect 6279 2111 6280 2118
rect 6263 2108 6264 2111
rect 6279 2108 6292 2111
rect 6215 2104 6245 2105
rect 6254 2104 6260 2105
rect 6263 2104 6292 2108
rect 6182 2103 6292 2104
rect 6182 2102 6298 2103
rect 5857 2094 5908 2102
rect 5857 2082 5882 2094
rect 5889 2082 5908 2094
rect 5939 2094 5989 2102
rect 5939 2086 5955 2094
rect 5962 2092 5989 2094
rect 5998 2092 6219 2102
rect 5962 2082 6219 2092
rect 6248 2094 6298 2102
rect 6248 2085 6264 2094
rect 5857 2074 5908 2082
rect 5955 2074 6219 2082
rect 6245 2082 6264 2085
rect 6271 2082 6298 2094
rect 6245 2074 6298 2082
rect 5873 2066 5874 2074
rect 5889 2066 5902 2074
rect 5873 2058 5889 2066
rect 5870 2051 5889 2054
rect 5870 2042 5892 2051
rect 5843 2032 5892 2042
rect 5843 2026 5873 2032
rect 5892 2027 5897 2032
rect 5815 2010 5889 2026
rect 5907 2018 5937 2074
rect 5972 2064 6180 2074
rect 6215 2070 6260 2074
rect 6263 2073 6264 2074
rect 6279 2073 6292 2074
rect 5998 2034 6187 2064
rect 6013 2031 6187 2034
rect 6006 2028 6187 2031
rect 5815 2008 5828 2010
rect 5843 2008 5877 2010
rect 5815 1992 5889 2008
rect 5916 2004 5929 2018
rect 5944 2004 5960 2020
rect 6006 2015 6017 2028
rect 5799 1970 5800 1986
rect 5815 1970 5828 1992
rect 5843 1970 5873 1992
rect 5916 1988 5978 2004
rect 6006 1997 6017 2013
rect 6022 2008 6032 2028
rect 6042 2008 6056 2028
rect 6059 2015 6068 2028
rect 6084 2015 6093 2028
rect 6022 1997 6056 2008
rect 6059 1997 6068 2013
rect 6084 1997 6093 2013
rect 6100 2008 6110 2028
rect 6120 2008 6134 2028
rect 6135 2015 6146 2028
rect 6100 1997 6134 2008
rect 6135 1997 6146 2013
rect 6192 2004 6208 2020
rect 6215 2018 6245 2070
rect 6279 2066 6280 2073
rect 6264 2058 6280 2066
rect 6251 2026 6264 2045
rect 6279 2026 6309 2042
rect 6251 2010 6325 2026
rect 6251 2008 6264 2010
rect 6279 2008 6313 2010
rect 5916 1986 5929 1988
rect 5944 1986 5978 1988
rect 5916 1970 5978 1986
rect 6022 1981 6038 1984
rect 6100 1981 6130 1992
rect 6178 1988 6224 2004
rect 6251 1992 6325 2008
rect 6178 1986 6212 1988
rect 6177 1970 6224 1986
rect 6251 1970 6264 1992
rect 6279 1970 6309 1992
rect 6336 1970 6337 1986
rect 6352 1970 6365 2130
rect 6395 2026 6408 2130
rect 6453 2108 6454 2118
rect 6469 2108 6482 2118
rect 6453 2104 6482 2108
rect 6487 2104 6517 2130
rect 6535 2116 6551 2118
rect 6623 2116 6676 2130
rect 6624 2114 6688 2116
rect 6731 2114 6746 2130
rect 6795 2127 6825 2130
rect 6795 2124 6831 2127
rect 6761 2116 6777 2118
rect 6535 2104 6550 2108
rect 6453 2102 6550 2104
rect 6578 2102 6746 2114
rect 6762 2104 6777 2108
rect 6795 2105 6834 2124
rect 6853 2118 6860 2119
rect 6859 2111 6860 2118
rect 6843 2108 6844 2111
rect 6859 2108 6872 2111
rect 6795 2104 6825 2105
rect 6834 2104 6840 2105
rect 6843 2104 6872 2108
rect 6762 2103 6872 2104
rect 6762 2102 6878 2103
rect 6437 2094 6488 2102
rect 6437 2082 6462 2094
rect 6469 2082 6488 2094
rect 6519 2094 6569 2102
rect 6519 2086 6535 2094
rect 6542 2092 6569 2094
rect 6578 2092 6799 2102
rect 6542 2082 6799 2092
rect 6828 2094 6878 2102
rect 6828 2085 6844 2094
rect 6437 2074 6488 2082
rect 6535 2074 6799 2082
rect 6825 2082 6844 2085
rect 6851 2082 6878 2094
rect 6825 2074 6878 2082
rect 6453 2066 6454 2074
rect 6469 2066 6482 2074
rect 6453 2058 6469 2066
rect 6450 2051 6469 2054
rect 6450 2042 6472 2051
rect 6423 2032 6472 2042
rect 6423 2026 6453 2032
rect 6472 2027 6477 2032
rect 6395 2010 6469 2026
rect 6487 2018 6517 2074
rect 6552 2064 6760 2074
rect 6795 2070 6840 2074
rect 6843 2073 6844 2074
rect 6859 2073 6872 2074
rect 6578 2034 6767 2064
rect 6593 2031 6767 2034
rect 6586 2028 6767 2031
rect 6395 2008 6408 2010
rect 6423 2008 6457 2010
rect 6395 1992 6469 2008
rect 6496 2004 6509 2018
rect 6524 2004 6540 2020
rect 6586 2015 6597 2028
rect 6379 1970 6380 1986
rect 6395 1970 6408 1992
rect 6423 1970 6453 1992
rect 6496 1988 6558 2004
rect 6586 1997 6597 2013
rect 6602 2008 6612 2028
rect 6622 2008 6636 2028
rect 6639 2015 6648 2028
rect 6664 2015 6673 2028
rect 6602 1997 6636 2008
rect 6639 1997 6648 2013
rect 6664 1997 6673 2013
rect 6680 2008 6690 2028
rect 6700 2008 6714 2028
rect 6715 2015 6726 2028
rect 6680 1997 6714 2008
rect 6715 1997 6726 2013
rect 6772 2004 6788 2020
rect 6795 2018 6825 2070
rect 6859 2066 6860 2073
rect 6844 2058 6860 2066
rect 6831 2026 6844 2045
rect 6859 2026 6889 2042
rect 6831 2010 6905 2026
rect 6831 2008 6844 2010
rect 6859 2008 6893 2010
rect 6496 1986 6509 1988
rect 6524 1986 6558 1988
rect 6496 1970 6558 1986
rect 6602 1981 6618 1984
rect 6680 1981 6710 1992
rect 6758 1988 6804 2004
rect 6831 1992 6905 2008
rect 6758 1986 6792 1988
rect 6757 1970 6804 1986
rect 6831 1970 6844 1992
rect 6859 1970 6889 1992
rect 6916 1970 6917 1986
rect 6932 1970 6945 2130
rect 6975 2026 6988 2130
rect 7033 2108 7034 2118
rect 7049 2108 7062 2118
rect 7033 2104 7062 2108
rect 7067 2104 7097 2130
rect 7115 2116 7131 2118
rect 7203 2116 7256 2130
rect 7204 2114 7268 2116
rect 7311 2114 7326 2130
rect 7375 2127 7405 2130
rect 7375 2124 7411 2127
rect 7341 2116 7357 2118
rect 7115 2104 7130 2108
rect 7033 2102 7130 2104
rect 7158 2102 7326 2114
rect 7342 2104 7357 2108
rect 7375 2105 7414 2124
rect 7433 2118 7440 2119
rect 7439 2111 7440 2118
rect 7423 2108 7424 2111
rect 7439 2108 7452 2111
rect 7375 2104 7405 2105
rect 7414 2104 7420 2105
rect 7423 2104 7452 2108
rect 7342 2103 7452 2104
rect 7342 2102 7458 2103
rect 7017 2094 7068 2102
rect 7017 2082 7042 2094
rect 7049 2082 7068 2094
rect 7099 2094 7149 2102
rect 7099 2086 7115 2094
rect 7122 2092 7149 2094
rect 7158 2092 7379 2102
rect 7122 2082 7379 2092
rect 7408 2094 7458 2102
rect 7408 2085 7424 2094
rect 7017 2074 7068 2082
rect 7115 2074 7379 2082
rect 7405 2082 7424 2085
rect 7431 2082 7458 2094
rect 7405 2074 7458 2082
rect 7033 2066 7034 2074
rect 7049 2066 7062 2074
rect 7033 2058 7049 2066
rect 7030 2051 7049 2054
rect 7030 2042 7052 2051
rect 7003 2032 7052 2042
rect 7003 2026 7033 2032
rect 7052 2027 7057 2032
rect 6975 2010 7049 2026
rect 7067 2018 7097 2074
rect 7132 2064 7340 2074
rect 7375 2070 7420 2074
rect 7423 2073 7424 2074
rect 7439 2073 7452 2074
rect 7158 2034 7347 2064
rect 7173 2031 7347 2034
rect 7166 2028 7347 2031
rect 6975 2008 6988 2010
rect 7003 2008 7037 2010
rect 6975 1992 7049 2008
rect 7076 2004 7089 2018
rect 7104 2004 7120 2020
rect 7166 2015 7177 2028
rect 6959 1970 6960 1986
rect 6975 1970 6988 1992
rect 7003 1970 7033 1992
rect 7076 1988 7138 2004
rect 7166 1997 7177 2013
rect 7182 2008 7192 2028
rect 7202 2008 7216 2028
rect 7219 2015 7228 2028
rect 7244 2015 7253 2028
rect 7182 1997 7216 2008
rect 7219 1997 7228 2013
rect 7244 1997 7253 2013
rect 7260 2008 7270 2028
rect 7280 2008 7294 2028
rect 7295 2015 7306 2028
rect 7260 1997 7294 2008
rect 7295 1997 7306 2013
rect 7352 2004 7368 2020
rect 7375 2018 7405 2070
rect 7439 2066 7440 2073
rect 7424 2058 7440 2066
rect 7411 2026 7424 2045
rect 7439 2026 7469 2042
rect 7411 2010 7485 2026
rect 7411 2008 7424 2010
rect 7439 2008 7473 2010
rect 7076 1986 7089 1988
rect 7104 1986 7138 1988
rect 7076 1970 7138 1986
rect 7182 1981 7198 1984
rect 7260 1981 7290 1992
rect 7338 1988 7384 2004
rect 7411 1992 7485 2008
rect 7338 1986 7372 1988
rect 7337 1970 7384 1986
rect 7411 1970 7424 1992
rect 7439 1970 7469 1992
rect 7496 1970 7497 1986
rect 7512 1970 7525 2130
rect 7555 2026 7568 2130
rect 7613 2108 7614 2118
rect 7629 2108 7642 2118
rect 7613 2104 7642 2108
rect 7647 2104 7677 2130
rect 7695 2116 7711 2118
rect 7783 2116 7836 2130
rect 7784 2114 7848 2116
rect 7891 2114 7906 2130
rect 7955 2127 7985 2130
rect 7955 2124 7991 2127
rect 7921 2116 7937 2118
rect 7695 2104 7710 2108
rect 7613 2102 7710 2104
rect 7738 2102 7906 2114
rect 7922 2104 7937 2108
rect 7955 2105 7994 2124
rect 8013 2118 8020 2119
rect 8019 2111 8020 2118
rect 8003 2108 8004 2111
rect 8019 2108 8032 2111
rect 7955 2104 7985 2105
rect 7994 2104 8000 2105
rect 8003 2104 8032 2108
rect 7922 2103 8032 2104
rect 7922 2102 8038 2103
rect 7597 2094 7648 2102
rect 7597 2082 7622 2094
rect 7629 2082 7648 2094
rect 7679 2094 7729 2102
rect 7679 2086 7695 2094
rect 7702 2092 7729 2094
rect 7738 2092 7959 2102
rect 7702 2082 7959 2092
rect 7988 2094 8038 2102
rect 7988 2085 8004 2094
rect 7597 2074 7648 2082
rect 7695 2074 7959 2082
rect 7985 2082 8004 2085
rect 8011 2082 8038 2094
rect 7985 2074 8038 2082
rect 7613 2066 7614 2074
rect 7629 2066 7642 2074
rect 7613 2058 7629 2066
rect 7610 2051 7629 2054
rect 7610 2042 7632 2051
rect 7583 2032 7632 2042
rect 7583 2026 7613 2032
rect 7632 2027 7637 2032
rect 7555 2010 7629 2026
rect 7647 2018 7677 2074
rect 7712 2064 7920 2074
rect 7955 2070 8000 2074
rect 8003 2073 8004 2074
rect 8019 2073 8032 2074
rect 7738 2034 7927 2064
rect 7753 2031 7927 2034
rect 7746 2028 7927 2031
rect 7555 2008 7568 2010
rect 7583 2008 7617 2010
rect 7555 1992 7629 2008
rect 7656 2004 7669 2018
rect 7684 2004 7700 2020
rect 7746 2015 7757 2028
rect 7539 1970 7540 1986
rect 7555 1970 7568 1992
rect 7583 1970 7613 1992
rect 7656 1988 7718 2004
rect 7746 1997 7757 2013
rect 7762 2008 7772 2028
rect 7782 2008 7796 2028
rect 7799 2015 7808 2028
rect 7824 2015 7833 2028
rect 7762 1997 7796 2008
rect 7799 1997 7808 2013
rect 7824 1997 7833 2013
rect 7840 2008 7850 2028
rect 7860 2008 7874 2028
rect 7875 2015 7886 2028
rect 7840 1997 7874 2008
rect 7875 1997 7886 2013
rect 7932 2004 7948 2020
rect 7955 2018 7985 2070
rect 8019 2066 8020 2073
rect 8004 2058 8020 2066
rect 7991 2026 8004 2045
rect 8019 2026 8049 2042
rect 7991 2010 8065 2026
rect 7991 2008 8004 2010
rect 8019 2008 8053 2010
rect 7656 1986 7669 1988
rect 7684 1986 7718 1988
rect 7656 1970 7718 1986
rect 7762 1981 7778 1984
rect 7840 1981 7870 1992
rect 7918 1988 7964 2004
rect 7991 1992 8065 2008
rect 7918 1986 7952 1988
rect 7917 1970 7964 1986
rect 7991 1970 8004 1992
rect 8019 1970 8049 1992
rect 8076 1970 8077 1986
rect 8092 1970 8105 2130
rect 8135 2026 8148 2130
rect 8193 2108 8194 2118
rect 8209 2108 8222 2118
rect 8193 2104 8222 2108
rect 8227 2104 8257 2130
rect 8275 2116 8291 2118
rect 8363 2116 8416 2130
rect 8364 2114 8428 2116
rect 8471 2114 8486 2130
rect 8535 2127 8565 2130
rect 8535 2124 8571 2127
rect 8501 2116 8517 2118
rect 8275 2104 8290 2108
rect 8193 2102 8290 2104
rect 8318 2102 8486 2114
rect 8502 2104 8517 2108
rect 8535 2105 8574 2124
rect 8593 2118 8600 2119
rect 8599 2111 8600 2118
rect 8583 2108 8584 2111
rect 8599 2108 8612 2111
rect 8535 2104 8565 2105
rect 8574 2104 8580 2105
rect 8583 2104 8612 2108
rect 8502 2103 8612 2104
rect 8502 2102 8618 2103
rect 8177 2094 8228 2102
rect 8177 2082 8202 2094
rect 8209 2082 8228 2094
rect 8259 2094 8309 2102
rect 8259 2086 8275 2094
rect 8282 2092 8309 2094
rect 8318 2092 8539 2102
rect 8282 2082 8539 2092
rect 8568 2094 8618 2102
rect 8568 2085 8584 2094
rect 8177 2074 8228 2082
rect 8275 2074 8539 2082
rect 8565 2082 8584 2085
rect 8591 2082 8618 2094
rect 8565 2074 8618 2082
rect 8193 2066 8194 2074
rect 8209 2066 8222 2074
rect 8193 2058 8209 2066
rect 8190 2051 8209 2054
rect 8190 2042 8212 2051
rect 8163 2032 8212 2042
rect 8163 2026 8193 2032
rect 8212 2027 8217 2032
rect 8135 2010 8209 2026
rect 8227 2018 8257 2074
rect 8292 2064 8500 2074
rect 8535 2070 8580 2074
rect 8583 2073 8584 2074
rect 8599 2073 8612 2074
rect 8318 2034 8507 2064
rect 8333 2031 8507 2034
rect 8326 2028 8507 2031
rect 8135 2008 8148 2010
rect 8163 2008 8197 2010
rect 8135 1992 8209 2008
rect 8236 2004 8249 2018
rect 8264 2004 8280 2020
rect 8326 2015 8337 2028
rect 8119 1970 8120 1986
rect 8135 1970 8148 1992
rect 8163 1970 8193 1992
rect 8236 1988 8298 2004
rect 8326 1997 8337 2013
rect 8342 2008 8352 2028
rect 8362 2008 8376 2028
rect 8379 2015 8388 2028
rect 8404 2015 8413 2028
rect 8342 1997 8376 2008
rect 8379 1997 8388 2013
rect 8404 1997 8413 2013
rect 8420 2008 8430 2028
rect 8440 2008 8454 2028
rect 8455 2015 8466 2028
rect 8420 1997 8454 2008
rect 8455 1997 8466 2013
rect 8512 2004 8528 2020
rect 8535 2018 8565 2070
rect 8599 2066 8600 2073
rect 8584 2058 8600 2066
rect 8571 2026 8584 2045
rect 8599 2026 8629 2042
rect 8571 2010 8645 2026
rect 8571 2008 8584 2010
rect 8599 2008 8633 2010
rect 8236 1986 8249 1988
rect 8264 1986 8298 1988
rect 8236 1970 8298 1986
rect 8342 1981 8358 1984
rect 8420 1981 8450 1992
rect 8498 1988 8544 2004
rect 8571 1992 8645 2008
rect 8498 1986 8532 1988
rect 8497 1970 8544 1986
rect 8571 1970 8584 1992
rect 8599 1970 8629 1992
rect 8656 1970 8657 1986
rect 8672 1970 8685 2130
rect 8715 2026 8728 2130
rect 8773 2108 8774 2118
rect 8789 2108 8802 2118
rect 8773 2104 8802 2108
rect 8807 2104 8837 2130
rect 8855 2116 8871 2118
rect 8943 2116 8996 2130
rect 8944 2114 9008 2116
rect 9051 2114 9066 2130
rect 9115 2127 9145 2130
rect 9115 2124 9151 2127
rect 9081 2116 9097 2118
rect 8855 2104 8870 2108
rect 8773 2102 8870 2104
rect 8898 2102 9066 2114
rect 9082 2104 9097 2108
rect 9115 2105 9154 2124
rect 9173 2118 9180 2119
rect 9179 2111 9180 2118
rect 9163 2108 9164 2111
rect 9179 2108 9192 2111
rect 9115 2104 9145 2105
rect 9154 2104 9160 2105
rect 9163 2104 9192 2108
rect 9082 2103 9192 2104
rect 9082 2102 9198 2103
rect 8757 2094 8808 2102
rect 8757 2082 8782 2094
rect 8789 2082 8808 2094
rect 8839 2094 8889 2102
rect 8839 2086 8855 2094
rect 8862 2092 8889 2094
rect 8898 2092 9119 2102
rect 8862 2082 9119 2092
rect 9148 2094 9198 2102
rect 9148 2085 9164 2094
rect 8757 2074 8808 2082
rect 8855 2074 9119 2082
rect 9145 2082 9164 2085
rect 9171 2082 9198 2094
rect 9145 2074 9198 2082
rect 8773 2066 8774 2074
rect 8789 2066 8802 2074
rect 8773 2058 8789 2066
rect 8770 2051 8789 2054
rect 8770 2042 8792 2051
rect 8743 2032 8792 2042
rect 8743 2026 8773 2032
rect 8792 2027 8797 2032
rect 8715 2010 8789 2026
rect 8807 2018 8837 2074
rect 8872 2064 9080 2074
rect 9115 2070 9160 2074
rect 9163 2073 9164 2074
rect 9179 2073 9192 2074
rect 8898 2034 9087 2064
rect 8913 2031 9087 2034
rect 8906 2028 9087 2031
rect 8715 2008 8728 2010
rect 8743 2008 8777 2010
rect 8715 1992 8789 2008
rect 8816 2004 8829 2018
rect 8844 2004 8860 2020
rect 8906 2015 8917 2028
rect 8699 1970 8700 1986
rect 8715 1970 8728 1992
rect 8743 1970 8773 1992
rect 8816 1988 8878 2004
rect 8906 1997 8917 2013
rect 8922 2008 8932 2028
rect 8942 2008 8956 2028
rect 8959 2015 8968 2028
rect 8984 2015 8993 2028
rect 8922 1997 8956 2008
rect 8959 1997 8968 2013
rect 8984 1997 8993 2013
rect 9000 2008 9010 2028
rect 9020 2008 9034 2028
rect 9035 2015 9046 2028
rect 9000 1997 9034 2008
rect 9035 1997 9046 2013
rect 9092 2004 9108 2020
rect 9115 2018 9145 2070
rect 9179 2066 9180 2073
rect 9164 2058 9180 2066
rect 9151 2026 9164 2045
rect 9179 2026 9209 2042
rect 9151 2010 9225 2026
rect 9151 2008 9164 2010
rect 9179 2008 9213 2010
rect 8816 1986 8829 1988
rect 8844 1986 8878 1988
rect 8816 1970 8878 1986
rect 8922 1981 8938 1984
rect 9000 1981 9030 1992
rect 9078 1988 9124 2004
rect 9151 1992 9225 2008
rect 9078 1986 9112 1988
rect 9077 1970 9124 1986
rect 9151 1970 9164 1992
rect 9179 1970 9209 1992
rect 9236 1970 9237 1986
rect 9252 1970 9265 2130
rect -7 1962 34 1970
rect -7 1936 8 1962
rect 15 1936 34 1962
rect 98 1958 160 1970
rect 172 1958 247 1970
rect 305 1958 380 1970
rect 392 1958 423 1970
rect 429 1958 464 1970
rect 98 1956 260 1958
rect -7 1928 34 1936
rect 116 1932 129 1956
rect 144 1954 159 1956
rect -1 1918 0 1928
rect 15 1918 28 1928
rect 43 1918 73 1932
rect 116 1918 159 1932
rect 183 1929 190 1936
rect 193 1932 260 1956
rect 292 1956 464 1958
rect 262 1934 290 1938
rect 292 1934 372 1956
rect 393 1954 408 1956
rect 262 1932 372 1934
rect 193 1928 372 1932
rect 166 1918 196 1928
rect 198 1918 351 1928
rect 359 1918 389 1928
rect 393 1918 423 1932
rect 451 1918 464 1956
rect 536 1962 571 1970
rect 536 1936 537 1962
rect 544 1936 571 1962
rect 479 1918 509 1932
rect 536 1928 571 1936
rect 573 1962 614 1970
rect 573 1936 588 1962
rect 595 1936 614 1962
rect 678 1958 740 1970
rect 752 1958 827 1970
rect 885 1958 960 1970
rect 972 1958 1003 1970
rect 1009 1958 1044 1970
rect 678 1956 840 1958
rect 573 1928 614 1936
rect 696 1932 709 1956
rect 724 1954 739 1956
rect 536 1918 537 1928
rect 552 1918 565 1928
rect 579 1918 580 1928
rect 595 1918 608 1928
rect 623 1918 653 1932
rect 696 1918 739 1932
rect 763 1929 770 1936
rect 773 1932 840 1956
rect 872 1956 1044 1958
rect 842 1934 870 1938
rect 872 1934 952 1956
rect 973 1954 988 1956
rect 842 1932 952 1934
rect 773 1928 952 1932
rect 746 1918 776 1928
rect 778 1918 931 1928
rect 939 1918 969 1928
rect 973 1918 1003 1932
rect 1031 1918 1044 1956
rect 1116 1962 1151 1970
rect 1116 1936 1117 1962
rect 1124 1936 1151 1962
rect 1059 1918 1089 1932
rect 1116 1928 1151 1936
rect 1153 1962 1194 1970
rect 1153 1936 1168 1962
rect 1175 1936 1194 1962
rect 1258 1958 1320 1970
rect 1332 1958 1407 1970
rect 1465 1958 1540 1970
rect 1552 1958 1583 1970
rect 1589 1958 1624 1970
rect 1258 1956 1420 1958
rect 1153 1928 1194 1936
rect 1276 1932 1289 1956
rect 1304 1954 1319 1956
rect 1116 1918 1117 1928
rect 1132 1918 1145 1928
rect 1159 1918 1160 1928
rect 1175 1918 1188 1928
rect 1203 1918 1233 1932
rect 1276 1918 1319 1932
rect 1343 1929 1350 1936
rect 1353 1932 1420 1956
rect 1452 1956 1624 1958
rect 1422 1934 1450 1938
rect 1452 1934 1532 1956
rect 1553 1954 1568 1956
rect 1422 1932 1532 1934
rect 1353 1928 1532 1932
rect 1326 1918 1356 1928
rect 1358 1918 1511 1928
rect 1519 1918 1549 1928
rect 1553 1918 1583 1932
rect 1611 1918 1624 1956
rect 1696 1962 1731 1970
rect 1696 1936 1697 1962
rect 1704 1936 1731 1962
rect 1639 1918 1669 1932
rect 1696 1928 1731 1936
rect 1733 1962 1774 1970
rect 1733 1936 1748 1962
rect 1755 1936 1774 1962
rect 1838 1958 1900 1970
rect 1912 1958 1987 1970
rect 2045 1958 2120 1970
rect 2132 1958 2163 1970
rect 2169 1958 2204 1970
rect 1838 1956 2000 1958
rect 1733 1928 1774 1936
rect 1856 1932 1869 1956
rect 1884 1954 1899 1956
rect 1696 1918 1697 1928
rect 1712 1918 1725 1928
rect 1739 1918 1740 1928
rect 1755 1918 1768 1928
rect 1783 1918 1813 1932
rect 1856 1918 1899 1932
rect 1923 1929 1930 1936
rect 1933 1932 2000 1956
rect 2032 1956 2204 1958
rect 2002 1934 2030 1938
rect 2032 1934 2112 1956
rect 2133 1954 2148 1956
rect 2002 1932 2112 1934
rect 1933 1928 2112 1932
rect 1906 1918 1936 1928
rect 1938 1918 2091 1928
rect 2099 1918 2129 1928
rect 2133 1918 2163 1932
rect 2191 1918 2204 1956
rect 2276 1962 2311 1970
rect 2276 1936 2277 1962
rect 2284 1936 2311 1962
rect 2219 1918 2249 1932
rect 2276 1928 2311 1936
rect 2313 1962 2354 1970
rect 2313 1936 2328 1962
rect 2335 1936 2354 1962
rect 2418 1958 2480 1970
rect 2492 1958 2567 1970
rect 2625 1958 2700 1970
rect 2712 1958 2743 1970
rect 2749 1958 2784 1970
rect 2418 1956 2580 1958
rect 2313 1928 2354 1936
rect 2436 1932 2449 1956
rect 2464 1954 2479 1956
rect 2276 1918 2277 1928
rect 2292 1918 2305 1928
rect 2319 1918 2320 1928
rect 2335 1918 2348 1928
rect 2363 1918 2393 1932
rect 2436 1918 2479 1932
rect 2503 1929 2510 1936
rect 2513 1932 2580 1956
rect 2612 1956 2784 1958
rect 2582 1934 2610 1938
rect 2612 1934 2692 1956
rect 2713 1954 2728 1956
rect 2582 1932 2692 1934
rect 2513 1928 2692 1932
rect 2486 1918 2516 1928
rect 2518 1918 2671 1928
rect 2679 1918 2709 1928
rect 2713 1918 2743 1932
rect 2771 1918 2784 1956
rect 2856 1962 2891 1970
rect 2856 1936 2857 1962
rect 2864 1936 2891 1962
rect 2799 1918 2829 1932
rect 2856 1928 2891 1936
rect 2893 1962 2934 1970
rect 2893 1936 2908 1962
rect 2915 1936 2934 1962
rect 2998 1958 3060 1970
rect 3072 1958 3147 1970
rect 3205 1958 3280 1970
rect 3292 1958 3323 1970
rect 3329 1958 3364 1970
rect 2998 1956 3160 1958
rect 2893 1928 2934 1936
rect 3016 1932 3029 1956
rect 3044 1954 3059 1956
rect 2856 1918 2857 1928
rect 2872 1918 2885 1928
rect 2899 1918 2900 1928
rect 2915 1918 2928 1928
rect 2943 1918 2973 1932
rect 3016 1918 3059 1932
rect 3083 1929 3090 1936
rect 3093 1932 3160 1956
rect 3192 1956 3364 1958
rect 3162 1934 3190 1938
rect 3192 1934 3272 1956
rect 3293 1954 3308 1956
rect 3162 1932 3272 1934
rect 3093 1928 3272 1932
rect 3066 1918 3096 1928
rect 3098 1918 3251 1928
rect 3259 1918 3289 1928
rect 3293 1918 3323 1932
rect 3351 1918 3364 1956
rect 3436 1962 3471 1970
rect 3436 1936 3437 1962
rect 3444 1936 3471 1962
rect 3379 1918 3409 1932
rect 3436 1928 3471 1936
rect 3473 1962 3514 1970
rect 3473 1936 3488 1962
rect 3495 1936 3514 1962
rect 3578 1958 3640 1970
rect 3652 1958 3727 1970
rect 3785 1958 3860 1970
rect 3872 1958 3903 1970
rect 3909 1958 3944 1970
rect 3578 1956 3740 1958
rect 3473 1928 3514 1936
rect 3596 1932 3609 1956
rect 3624 1954 3639 1956
rect 3436 1918 3437 1928
rect 3452 1918 3465 1928
rect 3479 1918 3480 1928
rect 3495 1918 3508 1928
rect 3523 1918 3553 1932
rect 3596 1918 3639 1932
rect 3663 1929 3670 1936
rect 3673 1932 3740 1956
rect 3772 1956 3944 1958
rect 3742 1934 3770 1938
rect 3772 1934 3852 1956
rect 3873 1954 3888 1956
rect 3742 1932 3852 1934
rect 3673 1928 3852 1932
rect 3646 1918 3676 1928
rect 3678 1918 3831 1928
rect 3839 1918 3869 1928
rect 3873 1918 3903 1932
rect 3931 1918 3944 1956
rect 4016 1962 4051 1970
rect 4016 1936 4017 1962
rect 4024 1936 4051 1962
rect 3959 1918 3989 1932
rect 4016 1928 4051 1936
rect 4053 1962 4094 1970
rect 4053 1936 4068 1962
rect 4075 1936 4094 1962
rect 4158 1958 4220 1970
rect 4232 1958 4307 1970
rect 4365 1958 4440 1970
rect 4452 1958 4483 1970
rect 4489 1958 4524 1970
rect 4158 1956 4320 1958
rect 4053 1928 4094 1936
rect 4176 1932 4189 1956
rect 4204 1954 4219 1956
rect 4016 1918 4017 1928
rect 4032 1918 4045 1928
rect 4059 1918 4060 1928
rect 4075 1918 4088 1928
rect 4103 1918 4133 1932
rect 4176 1918 4219 1932
rect 4243 1929 4250 1936
rect 4253 1932 4320 1956
rect 4352 1956 4524 1958
rect 4322 1934 4350 1938
rect 4352 1934 4432 1956
rect 4453 1954 4468 1956
rect 4322 1932 4432 1934
rect 4253 1928 4432 1932
rect 4226 1918 4256 1928
rect 4258 1918 4411 1928
rect 4419 1918 4449 1928
rect 4453 1918 4483 1932
rect 4511 1918 4524 1956
rect 4596 1962 4631 1970
rect 4596 1936 4597 1962
rect 4604 1936 4631 1962
rect 4539 1918 4569 1932
rect 4596 1928 4631 1936
rect 4633 1962 4674 1970
rect 4633 1936 4648 1962
rect 4655 1936 4674 1962
rect 4738 1958 4800 1970
rect 4812 1958 4887 1970
rect 4945 1958 5020 1970
rect 5032 1958 5063 1970
rect 5069 1958 5104 1970
rect 4738 1956 4900 1958
rect 4633 1928 4674 1936
rect 4756 1932 4769 1956
rect 4784 1954 4799 1956
rect 4596 1918 4597 1928
rect 4612 1918 4625 1928
rect 4639 1918 4640 1928
rect 4655 1918 4668 1928
rect 4683 1918 4713 1932
rect 4756 1918 4799 1932
rect 4823 1929 4830 1936
rect 4833 1932 4900 1956
rect 4932 1956 5104 1958
rect 4902 1934 4930 1938
rect 4932 1934 5012 1956
rect 5033 1954 5048 1956
rect 4902 1932 5012 1934
rect 4833 1928 5012 1932
rect 4806 1918 4836 1928
rect 4838 1918 4991 1928
rect 4999 1918 5029 1928
rect 5033 1918 5063 1932
rect 5091 1918 5104 1956
rect 5176 1962 5211 1970
rect 5176 1936 5177 1962
rect 5184 1936 5211 1962
rect 5119 1918 5149 1932
rect 5176 1928 5211 1936
rect 5213 1962 5254 1970
rect 5213 1936 5228 1962
rect 5235 1936 5254 1962
rect 5318 1958 5380 1970
rect 5392 1958 5467 1970
rect 5525 1958 5600 1970
rect 5612 1958 5643 1970
rect 5649 1958 5684 1970
rect 5318 1956 5480 1958
rect 5213 1928 5254 1936
rect 5336 1932 5349 1956
rect 5364 1954 5379 1956
rect 5176 1918 5177 1928
rect 5192 1918 5205 1928
rect 5219 1918 5220 1928
rect 5235 1918 5248 1928
rect 5263 1918 5293 1932
rect 5336 1918 5379 1932
rect 5403 1929 5410 1936
rect 5413 1932 5480 1956
rect 5512 1956 5684 1958
rect 5482 1934 5510 1938
rect 5512 1934 5592 1956
rect 5613 1954 5628 1956
rect 5482 1932 5592 1934
rect 5413 1928 5592 1932
rect 5386 1918 5416 1928
rect 5418 1918 5571 1928
rect 5579 1918 5609 1928
rect 5613 1918 5643 1932
rect 5671 1918 5684 1956
rect 5756 1962 5791 1970
rect 5756 1936 5757 1962
rect 5764 1936 5791 1962
rect 5699 1918 5729 1932
rect 5756 1928 5791 1936
rect 5793 1962 5834 1970
rect 5793 1936 5808 1962
rect 5815 1936 5834 1962
rect 5898 1958 5960 1970
rect 5972 1958 6047 1970
rect 6105 1958 6180 1970
rect 6192 1958 6223 1970
rect 6229 1958 6264 1970
rect 5898 1956 6060 1958
rect 5793 1928 5834 1936
rect 5916 1932 5929 1956
rect 5944 1954 5959 1956
rect 5756 1918 5757 1928
rect 5772 1918 5785 1928
rect 5799 1918 5800 1928
rect 5815 1918 5828 1928
rect 5843 1918 5873 1932
rect 5916 1918 5959 1932
rect 5983 1929 5990 1936
rect 5993 1932 6060 1956
rect 6092 1956 6264 1958
rect 6062 1934 6090 1938
rect 6092 1934 6172 1956
rect 6193 1954 6208 1956
rect 6062 1932 6172 1934
rect 5993 1928 6172 1932
rect 5966 1918 5996 1928
rect 5998 1918 6151 1928
rect 6159 1918 6189 1928
rect 6193 1918 6223 1932
rect 6251 1918 6264 1956
rect 6336 1962 6371 1970
rect 6336 1936 6337 1962
rect 6344 1936 6371 1962
rect 6279 1918 6309 1932
rect 6336 1928 6371 1936
rect 6373 1962 6414 1970
rect 6373 1936 6388 1962
rect 6395 1936 6414 1962
rect 6478 1958 6540 1970
rect 6552 1958 6627 1970
rect 6685 1958 6760 1970
rect 6772 1958 6803 1970
rect 6809 1958 6844 1970
rect 6478 1956 6640 1958
rect 6373 1928 6414 1936
rect 6496 1932 6509 1956
rect 6524 1954 6539 1956
rect 6336 1918 6337 1928
rect 6352 1918 6365 1928
rect 6379 1918 6380 1928
rect 6395 1918 6408 1928
rect 6423 1918 6453 1932
rect 6496 1918 6539 1932
rect 6563 1929 6570 1936
rect 6573 1932 6640 1956
rect 6672 1956 6844 1958
rect 6642 1934 6670 1938
rect 6672 1934 6752 1956
rect 6773 1954 6788 1956
rect 6642 1932 6752 1934
rect 6573 1928 6752 1932
rect 6546 1918 6576 1928
rect 6578 1918 6731 1928
rect 6739 1918 6769 1928
rect 6773 1918 6803 1932
rect 6831 1918 6844 1956
rect 6916 1962 6951 1970
rect 6916 1936 6917 1962
rect 6924 1936 6951 1962
rect 6859 1918 6889 1932
rect 6916 1928 6951 1936
rect 6953 1962 6994 1970
rect 6953 1936 6968 1962
rect 6975 1936 6994 1962
rect 7058 1958 7120 1970
rect 7132 1958 7207 1970
rect 7265 1958 7340 1970
rect 7352 1958 7383 1970
rect 7389 1958 7424 1970
rect 7058 1956 7220 1958
rect 6953 1928 6994 1936
rect 7076 1932 7089 1956
rect 7104 1954 7119 1956
rect 6916 1918 6917 1928
rect 6932 1918 6945 1928
rect 6959 1918 6960 1928
rect 6975 1918 6988 1928
rect 7003 1918 7033 1932
rect 7076 1918 7119 1932
rect 7143 1929 7150 1936
rect 7153 1932 7220 1956
rect 7252 1956 7424 1958
rect 7222 1934 7250 1938
rect 7252 1934 7332 1956
rect 7353 1954 7368 1956
rect 7222 1932 7332 1934
rect 7153 1928 7332 1932
rect 7126 1918 7156 1928
rect 7158 1918 7311 1928
rect 7319 1918 7349 1928
rect 7353 1918 7383 1932
rect 7411 1918 7424 1956
rect 7496 1962 7531 1970
rect 7496 1936 7497 1962
rect 7504 1936 7531 1962
rect 7439 1918 7469 1932
rect 7496 1928 7531 1936
rect 7533 1962 7574 1970
rect 7533 1936 7548 1962
rect 7555 1936 7574 1962
rect 7638 1958 7700 1970
rect 7712 1958 7787 1970
rect 7845 1958 7920 1970
rect 7932 1958 7963 1970
rect 7969 1958 8004 1970
rect 7638 1956 7800 1958
rect 7533 1928 7574 1936
rect 7656 1932 7669 1956
rect 7684 1954 7699 1956
rect 7496 1918 7497 1928
rect 7512 1918 7525 1928
rect 7539 1918 7540 1928
rect 7555 1918 7568 1928
rect 7583 1918 7613 1932
rect 7656 1918 7699 1932
rect 7723 1929 7730 1936
rect 7733 1932 7800 1956
rect 7832 1956 8004 1958
rect 7802 1934 7830 1938
rect 7832 1934 7912 1956
rect 7933 1954 7948 1956
rect 7802 1932 7912 1934
rect 7733 1928 7912 1932
rect 7706 1918 7736 1928
rect 7738 1918 7891 1928
rect 7899 1918 7929 1928
rect 7933 1918 7963 1932
rect 7991 1918 8004 1956
rect 8076 1962 8111 1970
rect 8076 1936 8077 1962
rect 8084 1936 8111 1962
rect 8019 1918 8049 1932
rect 8076 1928 8111 1936
rect 8113 1962 8154 1970
rect 8113 1936 8128 1962
rect 8135 1936 8154 1962
rect 8218 1958 8280 1970
rect 8292 1958 8367 1970
rect 8425 1958 8500 1970
rect 8512 1958 8543 1970
rect 8549 1958 8584 1970
rect 8218 1956 8380 1958
rect 8113 1928 8154 1936
rect 8236 1932 8249 1956
rect 8264 1954 8279 1956
rect 8076 1918 8077 1928
rect 8092 1918 8105 1928
rect 8119 1918 8120 1928
rect 8135 1918 8148 1928
rect 8163 1918 8193 1932
rect 8236 1918 8279 1932
rect 8303 1929 8310 1936
rect 8313 1932 8380 1956
rect 8412 1956 8584 1958
rect 8382 1934 8410 1938
rect 8412 1934 8492 1956
rect 8513 1954 8528 1956
rect 8382 1932 8492 1934
rect 8313 1928 8492 1932
rect 8286 1918 8316 1928
rect 8318 1918 8471 1928
rect 8479 1918 8509 1928
rect 8513 1918 8543 1932
rect 8571 1918 8584 1956
rect 8656 1962 8691 1970
rect 8656 1936 8657 1962
rect 8664 1936 8691 1962
rect 8599 1918 8629 1932
rect 8656 1928 8691 1936
rect 8693 1962 8734 1970
rect 8693 1936 8708 1962
rect 8715 1936 8734 1962
rect 8798 1958 8860 1970
rect 8872 1958 8947 1970
rect 9005 1958 9080 1970
rect 9092 1958 9123 1970
rect 9129 1958 9164 1970
rect 8798 1956 8960 1958
rect 8693 1928 8734 1936
rect 8816 1932 8829 1956
rect 8844 1954 8859 1956
rect 8656 1918 8657 1928
rect 8672 1918 8685 1928
rect 8699 1918 8700 1928
rect 8715 1918 8728 1928
rect 8743 1918 8773 1932
rect 8816 1918 8859 1932
rect 8883 1929 8890 1936
rect 8893 1932 8960 1956
rect 8992 1956 9164 1958
rect 8962 1934 8990 1938
rect 8992 1934 9072 1956
rect 9093 1954 9108 1956
rect 8962 1932 9072 1934
rect 8893 1928 9072 1932
rect 8866 1918 8896 1928
rect 8898 1918 9051 1928
rect 9059 1918 9089 1928
rect 9093 1918 9123 1932
rect 9151 1918 9164 1956
rect 9236 1962 9271 1970
rect 9236 1936 9237 1962
rect 9244 1936 9271 1962
rect 9179 1918 9209 1932
rect 9236 1928 9271 1936
rect 9236 1918 9237 1928
rect 9252 1918 9265 1928
rect -1 1912 9265 1918
rect 0 1904 9265 1912
rect 15 1874 28 1904
rect 43 1886 73 1904
rect 116 1890 130 1904
rect 166 1890 386 1904
rect 117 1888 130 1890
rect 83 1876 98 1888
rect 80 1874 102 1876
rect 107 1874 137 1888
rect 198 1886 351 1890
rect 180 1874 372 1886
rect 415 1874 445 1888
rect 451 1874 464 1904
rect 479 1886 509 1904
rect 552 1874 565 1904
rect 595 1874 608 1904
rect 623 1886 653 1904
rect 696 1890 710 1904
rect 746 1890 966 1904
rect 697 1888 710 1890
rect 663 1876 678 1888
rect 660 1874 682 1876
rect 687 1874 717 1888
rect 778 1886 931 1890
rect 760 1874 952 1886
rect 995 1874 1025 1888
rect 1031 1874 1044 1904
rect 1059 1886 1089 1904
rect 1132 1874 1145 1904
rect 1175 1874 1188 1904
rect 1203 1886 1233 1904
rect 1276 1890 1290 1904
rect 1326 1890 1546 1904
rect 1277 1888 1290 1890
rect 1243 1876 1258 1888
rect 1240 1874 1262 1876
rect 1267 1874 1297 1888
rect 1358 1886 1511 1890
rect 1340 1874 1532 1886
rect 1575 1874 1605 1888
rect 1611 1874 1624 1904
rect 1639 1886 1669 1904
rect 1712 1874 1725 1904
rect 1755 1874 1768 1904
rect 1783 1886 1813 1904
rect 1856 1890 1870 1904
rect 1906 1890 2126 1904
rect 1857 1888 1870 1890
rect 1823 1876 1838 1888
rect 1820 1874 1842 1876
rect 1847 1874 1877 1888
rect 1938 1886 2091 1890
rect 1920 1874 2112 1886
rect 2155 1874 2185 1888
rect 2191 1874 2204 1904
rect 2219 1886 2249 1904
rect 2292 1874 2305 1904
rect 2335 1874 2348 1904
rect 2363 1886 2393 1904
rect 2436 1890 2450 1904
rect 2486 1890 2706 1904
rect 2437 1888 2450 1890
rect 2403 1876 2418 1888
rect 2400 1874 2422 1876
rect 2427 1874 2457 1888
rect 2518 1886 2671 1890
rect 2500 1874 2692 1886
rect 2735 1874 2765 1888
rect 2771 1874 2784 1904
rect 2799 1886 2829 1904
rect 2872 1874 2885 1904
rect 2915 1874 2928 1904
rect 2943 1886 2973 1904
rect 3016 1890 3030 1904
rect 3066 1890 3286 1904
rect 3017 1888 3030 1890
rect 2983 1876 2998 1888
rect 2980 1874 3002 1876
rect 3007 1874 3037 1888
rect 3098 1886 3251 1890
rect 3080 1874 3272 1886
rect 3315 1874 3345 1888
rect 3351 1874 3364 1904
rect 3379 1886 3409 1904
rect 3452 1874 3465 1904
rect 3495 1874 3508 1904
rect 3523 1886 3553 1904
rect 3596 1890 3610 1904
rect 3646 1890 3866 1904
rect 3597 1888 3610 1890
rect 3563 1876 3578 1888
rect 3560 1874 3582 1876
rect 3587 1874 3617 1888
rect 3678 1886 3831 1890
rect 3660 1874 3852 1886
rect 3895 1874 3925 1888
rect 3931 1874 3944 1904
rect 3959 1886 3989 1904
rect 4032 1874 4045 1904
rect 4075 1874 4088 1904
rect 4103 1886 4133 1904
rect 4176 1890 4190 1904
rect 4226 1890 4446 1904
rect 4177 1888 4190 1890
rect 4143 1876 4158 1888
rect 4140 1874 4162 1876
rect 4167 1874 4197 1888
rect 4258 1886 4411 1890
rect 4240 1874 4432 1886
rect 4475 1874 4505 1888
rect 4511 1874 4524 1904
rect 4539 1886 4569 1904
rect 4612 1874 4625 1904
rect 4655 1874 4668 1904
rect 4683 1886 4713 1904
rect 4756 1890 4770 1904
rect 4806 1890 5026 1904
rect 4757 1888 4770 1890
rect 4723 1876 4738 1888
rect 4720 1874 4742 1876
rect 4747 1874 4777 1888
rect 4838 1886 4991 1890
rect 4820 1874 5012 1886
rect 5055 1874 5085 1888
rect 5091 1874 5104 1904
rect 5119 1886 5149 1904
rect 5192 1874 5205 1904
rect 5235 1874 5248 1904
rect 5263 1886 5293 1904
rect 5336 1890 5350 1904
rect 5386 1890 5606 1904
rect 5337 1888 5350 1890
rect 5303 1876 5318 1888
rect 5300 1874 5322 1876
rect 5327 1874 5357 1888
rect 5418 1886 5571 1890
rect 5400 1874 5592 1886
rect 5635 1874 5665 1888
rect 5671 1874 5684 1904
rect 5699 1886 5729 1904
rect 5772 1874 5785 1904
rect 5815 1874 5828 1904
rect 5843 1886 5873 1904
rect 5916 1890 5930 1904
rect 5966 1890 6186 1904
rect 5917 1888 5930 1890
rect 5883 1876 5898 1888
rect 5880 1874 5902 1876
rect 5907 1874 5937 1888
rect 5998 1886 6151 1890
rect 5980 1874 6172 1886
rect 6215 1874 6245 1888
rect 6251 1874 6264 1904
rect 6279 1886 6309 1904
rect 6352 1874 6365 1904
rect 6395 1874 6408 1904
rect 6423 1886 6453 1904
rect 6496 1890 6510 1904
rect 6546 1890 6766 1904
rect 6497 1888 6510 1890
rect 6463 1876 6478 1888
rect 6460 1874 6482 1876
rect 6487 1874 6517 1888
rect 6578 1886 6731 1890
rect 6560 1874 6752 1886
rect 6795 1874 6825 1888
rect 6831 1874 6844 1904
rect 6859 1886 6889 1904
rect 6932 1874 6945 1904
rect 6975 1874 6988 1904
rect 7003 1886 7033 1904
rect 7076 1890 7090 1904
rect 7126 1890 7346 1904
rect 7077 1888 7090 1890
rect 7043 1876 7058 1888
rect 7040 1874 7062 1876
rect 7067 1874 7097 1888
rect 7158 1886 7311 1890
rect 7140 1874 7332 1886
rect 7375 1874 7405 1888
rect 7411 1874 7424 1904
rect 7439 1886 7469 1904
rect 7512 1874 7525 1904
rect 7555 1874 7568 1904
rect 7583 1886 7613 1904
rect 7656 1890 7670 1904
rect 7706 1890 7926 1904
rect 7657 1888 7670 1890
rect 7623 1876 7638 1888
rect 7620 1874 7642 1876
rect 7647 1874 7677 1888
rect 7738 1886 7891 1890
rect 7720 1874 7912 1886
rect 7955 1874 7985 1888
rect 7991 1874 8004 1904
rect 8019 1886 8049 1904
rect 8092 1874 8105 1904
rect 8135 1874 8148 1904
rect 8163 1886 8193 1904
rect 8236 1890 8250 1904
rect 8286 1890 8506 1904
rect 8237 1888 8250 1890
rect 8203 1876 8218 1888
rect 8200 1874 8222 1876
rect 8227 1874 8257 1888
rect 8318 1886 8471 1890
rect 8300 1874 8492 1886
rect 8535 1874 8565 1888
rect 8571 1874 8584 1904
rect 8599 1886 8629 1904
rect 8672 1874 8685 1904
rect 8715 1874 8728 1904
rect 8743 1886 8773 1904
rect 8816 1890 8830 1904
rect 8866 1890 9086 1904
rect 8817 1888 8830 1890
rect 8783 1876 8798 1888
rect 8780 1874 8802 1876
rect 8807 1874 8837 1888
rect 8898 1886 9051 1890
rect 8880 1874 9072 1886
rect 9115 1874 9145 1888
rect 9151 1874 9164 1904
rect 9179 1886 9209 1904
rect 9252 1874 9265 1904
rect 0 1860 9265 1874
rect 15 1756 28 1860
rect 73 1838 74 1848
rect 89 1838 102 1848
rect 73 1834 102 1838
rect 107 1834 137 1860
rect 155 1846 171 1848
rect 243 1846 296 1860
rect 244 1844 308 1846
rect 351 1844 366 1860
rect 415 1857 445 1860
rect 415 1854 451 1857
rect 381 1846 397 1848
rect 155 1834 170 1838
rect 73 1832 170 1834
rect 198 1832 366 1844
rect 382 1834 397 1838
rect 415 1835 454 1854
rect 473 1848 480 1849
rect 479 1841 480 1848
rect 463 1838 464 1841
rect 479 1838 492 1841
rect 415 1834 445 1835
rect 454 1834 460 1835
rect 463 1834 492 1838
rect 382 1833 492 1834
rect 382 1832 498 1833
rect 57 1824 108 1832
rect 57 1812 82 1824
rect 89 1812 108 1824
rect 139 1824 189 1832
rect 139 1816 155 1824
rect 162 1822 189 1824
rect 198 1822 419 1832
rect 162 1812 419 1822
rect 448 1824 498 1832
rect 448 1815 464 1824
rect 57 1804 108 1812
rect 155 1804 419 1812
rect 445 1812 464 1815
rect 471 1812 498 1824
rect 445 1804 498 1812
rect 73 1796 74 1804
rect 89 1796 102 1804
rect 73 1788 89 1796
rect 70 1781 89 1784
rect 70 1772 92 1781
rect 43 1762 92 1772
rect 43 1756 73 1762
rect 92 1757 97 1762
rect 15 1740 89 1756
rect 107 1748 137 1804
rect 172 1794 380 1804
rect 415 1800 460 1804
rect 463 1803 464 1804
rect 479 1803 492 1804
rect 198 1764 387 1794
rect 213 1761 387 1764
rect 206 1758 387 1761
rect 15 1738 28 1740
rect 43 1738 77 1740
rect 15 1722 89 1738
rect 116 1734 129 1748
rect 144 1734 160 1750
rect 206 1745 217 1758
rect -1 1700 0 1716
rect 15 1700 28 1722
rect 43 1700 73 1722
rect 116 1718 178 1734
rect 206 1727 217 1743
rect 222 1738 232 1758
rect 242 1738 256 1758
rect 259 1745 268 1758
rect 284 1745 293 1758
rect 222 1727 256 1738
rect 259 1727 268 1743
rect 284 1727 293 1743
rect 300 1738 310 1758
rect 320 1738 334 1758
rect 335 1745 346 1758
rect 300 1727 334 1738
rect 335 1727 346 1743
rect 392 1734 408 1750
rect 415 1748 445 1800
rect 479 1796 480 1803
rect 464 1788 480 1796
rect 451 1756 464 1775
rect 479 1756 509 1772
rect 451 1740 525 1756
rect 451 1738 464 1740
rect 479 1738 513 1740
rect 116 1716 129 1718
rect 144 1716 178 1718
rect 116 1700 178 1716
rect 222 1711 238 1714
rect 300 1711 330 1722
rect 378 1718 424 1734
rect 451 1722 525 1738
rect 378 1716 412 1718
rect 377 1700 424 1716
rect 451 1700 464 1722
rect 479 1700 509 1722
rect 536 1700 537 1716
rect 552 1700 565 1860
rect 595 1756 608 1860
rect 653 1838 654 1848
rect 669 1838 682 1848
rect 653 1834 682 1838
rect 687 1834 717 1860
rect 735 1846 751 1848
rect 823 1846 876 1860
rect 824 1844 888 1846
rect 931 1844 946 1860
rect 995 1857 1025 1860
rect 995 1854 1031 1857
rect 961 1846 977 1848
rect 735 1834 750 1838
rect 653 1832 750 1834
rect 778 1832 946 1844
rect 962 1834 977 1838
rect 995 1835 1034 1854
rect 1053 1848 1060 1849
rect 1059 1841 1060 1848
rect 1043 1838 1044 1841
rect 1059 1838 1072 1841
rect 995 1834 1025 1835
rect 1034 1834 1040 1835
rect 1043 1834 1072 1838
rect 962 1833 1072 1834
rect 962 1832 1078 1833
rect 637 1824 688 1832
rect 637 1812 662 1824
rect 669 1812 688 1824
rect 719 1824 769 1832
rect 719 1816 735 1824
rect 742 1822 769 1824
rect 778 1822 999 1832
rect 742 1812 999 1822
rect 1028 1824 1078 1832
rect 1028 1815 1044 1824
rect 637 1804 688 1812
rect 735 1804 999 1812
rect 1025 1812 1044 1815
rect 1051 1812 1078 1824
rect 1025 1804 1078 1812
rect 653 1796 654 1804
rect 669 1796 682 1804
rect 653 1788 669 1796
rect 650 1781 669 1784
rect 650 1772 672 1781
rect 623 1762 672 1772
rect 623 1756 653 1762
rect 672 1757 677 1762
rect 595 1740 669 1756
rect 687 1748 717 1804
rect 752 1794 960 1804
rect 995 1800 1040 1804
rect 1043 1803 1044 1804
rect 1059 1803 1072 1804
rect 778 1764 967 1794
rect 793 1761 967 1764
rect 786 1758 967 1761
rect 595 1738 608 1740
rect 623 1738 657 1740
rect 595 1722 669 1738
rect 696 1734 709 1748
rect 724 1734 740 1750
rect 786 1745 797 1758
rect 579 1700 580 1716
rect 595 1700 608 1722
rect 623 1700 653 1722
rect 696 1718 758 1734
rect 786 1727 797 1743
rect 802 1738 812 1758
rect 822 1738 836 1758
rect 839 1745 848 1758
rect 864 1745 873 1758
rect 802 1727 836 1738
rect 839 1727 848 1743
rect 864 1727 873 1743
rect 880 1738 890 1758
rect 900 1738 914 1758
rect 915 1745 926 1758
rect 880 1727 914 1738
rect 915 1727 926 1743
rect 972 1734 988 1750
rect 995 1748 1025 1800
rect 1059 1796 1060 1803
rect 1044 1788 1060 1796
rect 1031 1756 1044 1775
rect 1059 1756 1089 1772
rect 1031 1740 1105 1756
rect 1031 1738 1044 1740
rect 1059 1738 1093 1740
rect 696 1716 709 1718
rect 724 1716 758 1718
rect 696 1700 758 1716
rect 802 1711 818 1714
rect 880 1711 910 1722
rect 958 1718 1004 1734
rect 1031 1722 1105 1738
rect 958 1716 992 1718
rect 957 1700 1004 1716
rect 1031 1700 1044 1722
rect 1059 1700 1089 1722
rect 1116 1700 1117 1716
rect 1132 1700 1145 1860
rect 1175 1756 1188 1860
rect 1233 1838 1234 1848
rect 1249 1838 1262 1848
rect 1233 1834 1262 1838
rect 1267 1834 1297 1860
rect 1315 1846 1331 1848
rect 1403 1846 1456 1860
rect 1404 1844 1468 1846
rect 1511 1844 1526 1860
rect 1575 1857 1605 1860
rect 1575 1854 1611 1857
rect 1541 1846 1557 1848
rect 1315 1834 1330 1838
rect 1233 1832 1330 1834
rect 1358 1832 1526 1844
rect 1542 1834 1557 1838
rect 1575 1835 1614 1854
rect 1633 1848 1640 1849
rect 1639 1841 1640 1848
rect 1623 1838 1624 1841
rect 1639 1838 1652 1841
rect 1575 1834 1605 1835
rect 1614 1834 1620 1835
rect 1623 1834 1652 1838
rect 1542 1833 1652 1834
rect 1542 1832 1658 1833
rect 1217 1824 1268 1832
rect 1217 1812 1242 1824
rect 1249 1812 1268 1824
rect 1299 1824 1349 1832
rect 1299 1816 1315 1824
rect 1322 1822 1349 1824
rect 1358 1822 1579 1832
rect 1322 1812 1579 1822
rect 1608 1824 1658 1832
rect 1608 1815 1624 1824
rect 1217 1804 1268 1812
rect 1315 1804 1579 1812
rect 1605 1812 1624 1815
rect 1631 1812 1658 1824
rect 1605 1804 1658 1812
rect 1233 1796 1234 1804
rect 1249 1796 1262 1804
rect 1233 1788 1249 1796
rect 1230 1781 1249 1784
rect 1230 1772 1252 1781
rect 1203 1762 1252 1772
rect 1203 1756 1233 1762
rect 1252 1757 1257 1762
rect 1175 1740 1249 1756
rect 1267 1748 1297 1804
rect 1332 1794 1540 1804
rect 1575 1800 1620 1804
rect 1623 1803 1624 1804
rect 1639 1803 1652 1804
rect 1358 1764 1547 1794
rect 1373 1761 1547 1764
rect 1366 1758 1547 1761
rect 1175 1738 1188 1740
rect 1203 1738 1237 1740
rect 1175 1722 1249 1738
rect 1276 1734 1289 1748
rect 1304 1734 1320 1750
rect 1366 1745 1377 1758
rect 1159 1700 1160 1716
rect 1175 1700 1188 1722
rect 1203 1700 1233 1722
rect 1276 1718 1338 1734
rect 1366 1727 1377 1743
rect 1382 1738 1392 1758
rect 1402 1738 1416 1758
rect 1419 1745 1428 1758
rect 1444 1745 1453 1758
rect 1382 1727 1416 1738
rect 1419 1727 1428 1743
rect 1444 1727 1453 1743
rect 1460 1738 1470 1758
rect 1480 1738 1494 1758
rect 1495 1745 1506 1758
rect 1460 1727 1494 1738
rect 1495 1727 1506 1743
rect 1552 1734 1568 1750
rect 1575 1748 1605 1800
rect 1639 1796 1640 1803
rect 1624 1788 1640 1796
rect 1611 1756 1624 1775
rect 1639 1756 1669 1772
rect 1611 1740 1685 1756
rect 1611 1738 1624 1740
rect 1639 1738 1673 1740
rect 1276 1716 1289 1718
rect 1304 1716 1338 1718
rect 1276 1700 1338 1716
rect 1382 1711 1398 1714
rect 1460 1711 1490 1722
rect 1538 1718 1584 1734
rect 1611 1722 1685 1738
rect 1538 1716 1572 1718
rect 1537 1700 1584 1716
rect 1611 1700 1624 1722
rect 1639 1700 1669 1722
rect 1696 1700 1697 1716
rect 1712 1700 1725 1860
rect 1755 1756 1768 1860
rect 1813 1838 1814 1848
rect 1829 1838 1842 1848
rect 1813 1834 1842 1838
rect 1847 1834 1877 1860
rect 1895 1846 1911 1848
rect 1983 1846 2036 1860
rect 1984 1844 2048 1846
rect 2091 1844 2106 1860
rect 2155 1857 2185 1860
rect 2155 1854 2191 1857
rect 2121 1846 2137 1848
rect 1895 1834 1910 1838
rect 1813 1832 1910 1834
rect 1938 1832 2106 1844
rect 2122 1834 2137 1838
rect 2155 1835 2194 1854
rect 2213 1848 2220 1849
rect 2219 1841 2220 1848
rect 2203 1838 2204 1841
rect 2219 1838 2232 1841
rect 2155 1834 2185 1835
rect 2194 1834 2200 1835
rect 2203 1834 2232 1838
rect 2122 1833 2232 1834
rect 2122 1832 2238 1833
rect 1797 1824 1848 1832
rect 1797 1812 1822 1824
rect 1829 1812 1848 1824
rect 1879 1824 1929 1832
rect 1879 1816 1895 1824
rect 1902 1822 1929 1824
rect 1938 1822 2159 1832
rect 1902 1812 2159 1822
rect 2188 1824 2238 1832
rect 2188 1815 2204 1824
rect 1797 1804 1848 1812
rect 1895 1804 2159 1812
rect 2185 1812 2204 1815
rect 2211 1812 2238 1824
rect 2185 1804 2238 1812
rect 1813 1796 1814 1804
rect 1829 1796 1842 1804
rect 1813 1788 1829 1796
rect 1810 1781 1829 1784
rect 1810 1772 1832 1781
rect 1783 1762 1832 1772
rect 1783 1756 1813 1762
rect 1832 1757 1837 1762
rect 1755 1740 1829 1756
rect 1847 1748 1877 1804
rect 1912 1794 2120 1804
rect 2155 1800 2200 1804
rect 2203 1803 2204 1804
rect 2219 1803 2232 1804
rect 1938 1764 2127 1794
rect 1953 1761 2127 1764
rect 1946 1758 2127 1761
rect 1755 1738 1768 1740
rect 1783 1738 1817 1740
rect 1755 1722 1829 1738
rect 1856 1734 1869 1748
rect 1884 1734 1900 1750
rect 1946 1745 1957 1758
rect 1739 1700 1740 1716
rect 1755 1700 1768 1722
rect 1783 1700 1813 1722
rect 1856 1718 1918 1734
rect 1946 1727 1957 1743
rect 1962 1738 1972 1758
rect 1982 1738 1996 1758
rect 1999 1745 2008 1758
rect 2024 1745 2033 1758
rect 1962 1727 1996 1738
rect 1999 1727 2008 1743
rect 2024 1727 2033 1743
rect 2040 1738 2050 1758
rect 2060 1738 2074 1758
rect 2075 1745 2086 1758
rect 2040 1727 2074 1738
rect 2075 1727 2086 1743
rect 2132 1734 2148 1750
rect 2155 1748 2185 1800
rect 2219 1796 2220 1803
rect 2204 1788 2220 1796
rect 2191 1756 2204 1775
rect 2219 1756 2249 1772
rect 2191 1740 2265 1756
rect 2191 1738 2204 1740
rect 2219 1738 2253 1740
rect 1856 1716 1869 1718
rect 1884 1716 1918 1718
rect 1856 1700 1918 1716
rect 1962 1711 1976 1714
rect 2040 1711 2070 1722
rect 2118 1718 2164 1734
rect 2191 1722 2265 1738
rect 2118 1716 2152 1718
rect 2117 1700 2164 1716
rect 2191 1700 2204 1722
rect 2219 1700 2249 1722
rect 2276 1700 2277 1716
rect 2292 1700 2305 1860
rect 2335 1756 2348 1860
rect 2393 1838 2394 1848
rect 2409 1838 2422 1848
rect 2393 1834 2422 1838
rect 2427 1834 2457 1860
rect 2475 1846 2491 1848
rect 2563 1846 2616 1860
rect 2564 1844 2628 1846
rect 2671 1844 2686 1860
rect 2735 1857 2765 1860
rect 2735 1854 2771 1857
rect 2701 1846 2717 1848
rect 2475 1834 2490 1838
rect 2393 1832 2490 1834
rect 2518 1832 2686 1844
rect 2702 1834 2717 1838
rect 2735 1835 2774 1854
rect 2793 1848 2800 1849
rect 2799 1841 2800 1848
rect 2783 1838 2784 1841
rect 2799 1838 2812 1841
rect 2735 1834 2765 1835
rect 2774 1834 2780 1835
rect 2783 1834 2812 1838
rect 2702 1833 2812 1834
rect 2702 1832 2818 1833
rect 2377 1824 2428 1832
rect 2377 1812 2402 1824
rect 2409 1812 2428 1824
rect 2459 1824 2509 1832
rect 2459 1816 2475 1824
rect 2482 1822 2509 1824
rect 2518 1822 2739 1832
rect 2482 1812 2739 1822
rect 2768 1824 2818 1832
rect 2768 1815 2784 1824
rect 2377 1804 2428 1812
rect 2475 1804 2739 1812
rect 2765 1812 2784 1815
rect 2791 1812 2818 1824
rect 2765 1804 2818 1812
rect 2393 1796 2394 1804
rect 2409 1796 2422 1804
rect 2393 1788 2409 1796
rect 2390 1781 2409 1784
rect 2390 1772 2412 1781
rect 2363 1762 2412 1772
rect 2363 1756 2393 1762
rect 2412 1757 2417 1762
rect 2335 1740 2409 1756
rect 2427 1748 2457 1804
rect 2492 1794 2700 1804
rect 2735 1800 2780 1804
rect 2783 1803 2784 1804
rect 2799 1803 2812 1804
rect 2518 1764 2707 1794
rect 2533 1761 2707 1764
rect 2526 1758 2707 1761
rect 2335 1738 2348 1740
rect 2363 1738 2397 1740
rect 2335 1722 2409 1738
rect 2436 1734 2449 1748
rect 2464 1734 2480 1750
rect 2526 1745 2537 1758
rect 2319 1700 2320 1716
rect 2335 1700 2348 1722
rect 2363 1700 2393 1722
rect 2436 1718 2498 1734
rect 2526 1727 2537 1743
rect 2542 1738 2552 1758
rect 2562 1738 2576 1758
rect 2579 1745 2588 1758
rect 2604 1745 2613 1758
rect 2542 1727 2576 1738
rect 2579 1727 2588 1743
rect 2604 1727 2613 1743
rect 2620 1738 2630 1758
rect 2640 1738 2654 1758
rect 2655 1745 2666 1758
rect 2620 1727 2654 1738
rect 2655 1727 2666 1743
rect 2712 1734 2728 1750
rect 2735 1748 2765 1800
rect 2799 1796 2800 1803
rect 2784 1788 2800 1796
rect 2771 1756 2784 1775
rect 2799 1756 2829 1772
rect 2771 1740 2845 1756
rect 2771 1738 2784 1740
rect 2799 1738 2833 1740
rect 2436 1716 2449 1718
rect 2464 1716 2498 1718
rect 2436 1700 2498 1716
rect 2542 1711 2558 1714
rect 2620 1711 2650 1722
rect 2698 1718 2744 1734
rect 2771 1722 2845 1738
rect 2698 1716 2732 1718
rect 2697 1700 2744 1716
rect 2771 1700 2784 1722
rect 2799 1700 2829 1722
rect 2856 1700 2857 1716
rect 2872 1700 2885 1860
rect 2915 1756 2928 1860
rect 2973 1838 2974 1848
rect 2989 1838 3002 1848
rect 2973 1834 3002 1838
rect 3007 1834 3037 1860
rect 3055 1846 3071 1848
rect 3143 1846 3196 1860
rect 3144 1844 3208 1846
rect 3251 1844 3266 1860
rect 3315 1857 3345 1860
rect 3315 1854 3351 1857
rect 3281 1846 3297 1848
rect 3055 1834 3070 1838
rect 2973 1832 3070 1834
rect 3098 1832 3266 1844
rect 3282 1834 3297 1838
rect 3315 1835 3354 1854
rect 3373 1848 3380 1849
rect 3379 1841 3380 1848
rect 3363 1838 3364 1841
rect 3379 1838 3392 1841
rect 3315 1834 3345 1835
rect 3354 1834 3360 1835
rect 3363 1834 3392 1838
rect 3282 1833 3392 1834
rect 3282 1832 3398 1833
rect 2957 1824 3008 1832
rect 2957 1812 2982 1824
rect 2989 1812 3008 1824
rect 3039 1824 3089 1832
rect 3039 1816 3055 1824
rect 3062 1822 3089 1824
rect 3098 1822 3319 1832
rect 3062 1812 3319 1822
rect 3348 1824 3398 1832
rect 3348 1815 3364 1824
rect 2957 1804 3008 1812
rect 3055 1804 3319 1812
rect 3345 1812 3364 1815
rect 3371 1812 3398 1824
rect 3345 1804 3398 1812
rect 2973 1796 2974 1804
rect 2989 1796 3002 1804
rect 2973 1788 2989 1796
rect 2970 1781 2989 1784
rect 2970 1772 2992 1781
rect 2943 1762 2992 1772
rect 2943 1756 2973 1762
rect 2992 1757 2997 1762
rect 2915 1740 2989 1756
rect 3007 1748 3037 1804
rect 3072 1794 3280 1804
rect 3315 1800 3360 1804
rect 3363 1803 3364 1804
rect 3379 1803 3392 1804
rect 3098 1764 3287 1794
rect 3113 1761 3287 1764
rect 3106 1758 3287 1761
rect 2915 1738 2928 1740
rect 2943 1738 2977 1740
rect 2915 1722 2989 1738
rect 3016 1734 3029 1748
rect 3044 1734 3060 1750
rect 3106 1745 3117 1758
rect 2899 1700 2900 1716
rect 2915 1700 2928 1722
rect 2943 1700 2973 1722
rect 3016 1718 3078 1734
rect 3106 1727 3117 1743
rect 3122 1738 3132 1758
rect 3142 1738 3156 1758
rect 3159 1745 3168 1758
rect 3184 1745 3193 1758
rect 3122 1727 3156 1738
rect 3159 1727 3168 1743
rect 3184 1727 3193 1743
rect 3200 1738 3210 1758
rect 3220 1738 3234 1758
rect 3235 1745 3246 1758
rect 3200 1727 3234 1738
rect 3235 1727 3246 1743
rect 3292 1734 3308 1750
rect 3315 1748 3345 1800
rect 3379 1796 3380 1803
rect 3364 1788 3380 1796
rect 3351 1756 3364 1775
rect 3379 1756 3409 1772
rect 3351 1740 3425 1756
rect 3351 1738 3364 1740
rect 3379 1738 3413 1740
rect 3016 1716 3029 1718
rect 3044 1716 3078 1718
rect 3016 1700 3078 1716
rect 3122 1711 3138 1714
rect 3200 1711 3230 1722
rect 3278 1718 3324 1734
rect 3351 1722 3425 1738
rect 3278 1716 3312 1718
rect 3277 1700 3324 1716
rect 3351 1700 3364 1722
rect 3379 1700 3409 1722
rect 3436 1700 3437 1716
rect 3452 1700 3465 1860
rect 3495 1756 3508 1860
rect 3553 1838 3554 1848
rect 3569 1838 3582 1848
rect 3553 1834 3582 1838
rect 3587 1834 3617 1860
rect 3635 1846 3651 1848
rect 3723 1846 3776 1860
rect 3724 1844 3788 1846
rect 3831 1844 3846 1860
rect 3895 1857 3925 1860
rect 3895 1854 3931 1857
rect 3861 1846 3877 1848
rect 3635 1834 3650 1838
rect 3553 1832 3650 1834
rect 3678 1832 3846 1844
rect 3862 1834 3877 1838
rect 3895 1835 3934 1854
rect 3953 1848 3960 1849
rect 3959 1841 3960 1848
rect 3943 1838 3944 1841
rect 3959 1838 3972 1841
rect 3895 1834 3925 1835
rect 3934 1834 3940 1835
rect 3943 1834 3972 1838
rect 3862 1833 3972 1834
rect 3862 1832 3978 1833
rect 3537 1824 3588 1832
rect 3537 1812 3562 1824
rect 3569 1812 3588 1824
rect 3619 1824 3669 1832
rect 3619 1816 3635 1824
rect 3642 1822 3669 1824
rect 3678 1822 3899 1832
rect 3642 1812 3899 1822
rect 3928 1824 3978 1832
rect 3928 1815 3944 1824
rect 3537 1804 3588 1812
rect 3635 1804 3899 1812
rect 3925 1812 3944 1815
rect 3951 1812 3978 1824
rect 3925 1804 3978 1812
rect 3553 1796 3554 1804
rect 3569 1796 3582 1804
rect 3553 1788 3569 1796
rect 3550 1781 3569 1784
rect 3550 1772 3572 1781
rect 3523 1762 3572 1772
rect 3523 1756 3553 1762
rect 3572 1757 3577 1762
rect 3495 1740 3569 1756
rect 3587 1748 3617 1804
rect 3652 1794 3860 1804
rect 3895 1800 3940 1804
rect 3943 1803 3944 1804
rect 3959 1803 3972 1804
rect 3678 1764 3867 1794
rect 3693 1761 3867 1764
rect 3686 1758 3867 1761
rect 3495 1738 3508 1740
rect 3523 1738 3557 1740
rect 3495 1722 3569 1738
rect 3596 1734 3609 1748
rect 3624 1734 3640 1750
rect 3686 1745 3697 1758
rect 3479 1700 3480 1716
rect 3495 1700 3508 1722
rect 3523 1700 3553 1722
rect 3596 1718 3658 1734
rect 3686 1727 3697 1743
rect 3702 1738 3712 1758
rect 3722 1738 3736 1758
rect 3739 1745 3748 1758
rect 3764 1745 3773 1758
rect 3702 1727 3736 1738
rect 3739 1727 3748 1743
rect 3764 1727 3773 1743
rect 3780 1738 3790 1758
rect 3800 1738 3814 1758
rect 3815 1745 3826 1758
rect 3780 1727 3814 1738
rect 3815 1727 3826 1743
rect 3872 1734 3888 1750
rect 3895 1748 3925 1800
rect 3959 1796 3960 1803
rect 3944 1788 3960 1796
rect 3931 1756 3944 1775
rect 3959 1756 3989 1772
rect 3931 1740 4005 1756
rect 3931 1738 3944 1740
rect 3959 1738 3993 1740
rect 3596 1716 3609 1718
rect 3624 1716 3658 1718
rect 3596 1700 3658 1716
rect 3702 1711 3718 1714
rect 3780 1711 3810 1722
rect 3858 1718 3904 1734
rect 3931 1722 4005 1738
rect 3858 1716 3892 1718
rect 3857 1700 3904 1716
rect 3931 1700 3944 1722
rect 3959 1700 3989 1722
rect 4016 1700 4017 1716
rect 4032 1700 4045 1860
rect 4075 1756 4088 1860
rect 4133 1838 4134 1848
rect 4149 1838 4162 1848
rect 4133 1834 4162 1838
rect 4167 1834 4197 1860
rect 4215 1846 4231 1848
rect 4303 1846 4356 1860
rect 4304 1844 4368 1846
rect 4411 1844 4426 1860
rect 4475 1857 4505 1860
rect 4475 1854 4511 1857
rect 4441 1846 4457 1848
rect 4215 1834 4230 1838
rect 4133 1832 4230 1834
rect 4258 1832 4426 1844
rect 4442 1834 4457 1838
rect 4475 1835 4514 1854
rect 4533 1848 4540 1849
rect 4539 1841 4540 1848
rect 4523 1838 4524 1841
rect 4539 1838 4552 1841
rect 4475 1834 4505 1835
rect 4514 1834 4520 1835
rect 4523 1834 4552 1838
rect 4442 1833 4552 1834
rect 4442 1832 4558 1833
rect 4117 1824 4168 1832
rect 4117 1812 4142 1824
rect 4149 1812 4168 1824
rect 4199 1824 4249 1832
rect 4199 1816 4215 1824
rect 4222 1822 4249 1824
rect 4258 1822 4479 1832
rect 4222 1812 4479 1822
rect 4508 1824 4558 1832
rect 4508 1815 4524 1824
rect 4117 1804 4168 1812
rect 4215 1804 4479 1812
rect 4505 1812 4524 1815
rect 4531 1812 4558 1824
rect 4505 1804 4558 1812
rect 4133 1796 4134 1804
rect 4149 1796 4162 1804
rect 4133 1788 4149 1796
rect 4130 1781 4149 1784
rect 4130 1772 4152 1781
rect 4103 1762 4152 1772
rect 4103 1756 4133 1762
rect 4152 1757 4157 1762
rect 4075 1740 4149 1756
rect 4167 1748 4197 1804
rect 4232 1794 4440 1804
rect 4475 1800 4520 1804
rect 4523 1803 4524 1804
rect 4539 1803 4552 1804
rect 4258 1764 4447 1794
rect 4273 1761 4447 1764
rect 4266 1758 4447 1761
rect 4075 1738 4088 1740
rect 4103 1738 4137 1740
rect 4075 1722 4149 1738
rect 4176 1734 4189 1748
rect 4204 1734 4220 1750
rect 4266 1745 4277 1758
rect 4059 1700 4060 1716
rect 4075 1700 4088 1722
rect 4103 1700 4133 1722
rect 4176 1718 4238 1734
rect 4266 1727 4277 1743
rect 4282 1738 4292 1758
rect 4302 1738 4316 1758
rect 4319 1745 4328 1758
rect 4344 1745 4353 1758
rect 4282 1727 4316 1738
rect 4319 1727 4328 1743
rect 4344 1727 4353 1743
rect 4360 1738 4370 1758
rect 4380 1738 4394 1758
rect 4395 1745 4406 1758
rect 4360 1727 4394 1738
rect 4395 1727 4406 1743
rect 4452 1734 4468 1750
rect 4475 1748 4505 1800
rect 4539 1796 4540 1803
rect 4524 1788 4540 1796
rect 4511 1756 4524 1775
rect 4539 1756 4569 1772
rect 4511 1740 4585 1756
rect 4511 1738 4524 1740
rect 4539 1738 4573 1740
rect 4176 1716 4189 1718
rect 4204 1716 4238 1718
rect 4176 1700 4238 1716
rect 4282 1711 4298 1714
rect 4360 1711 4390 1722
rect 4438 1718 4484 1734
rect 4511 1722 4585 1738
rect 4438 1716 4472 1718
rect 4437 1700 4484 1716
rect 4511 1700 4524 1722
rect 4539 1700 4569 1722
rect 4596 1700 4597 1716
rect 4612 1700 4625 1860
rect 4655 1756 4668 1860
rect 4713 1838 4714 1848
rect 4729 1838 4742 1848
rect 4713 1834 4742 1838
rect 4747 1834 4777 1860
rect 4795 1846 4811 1848
rect 4883 1846 4936 1860
rect 4884 1844 4948 1846
rect 4991 1844 5006 1860
rect 5055 1857 5085 1860
rect 5055 1854 5091 1857
rect 5021 1846 5037 1848
rect 4795 1834 4810 1838
rect 4713 1832 4810 1834
rect 4838 1832 5006 1844
rect 5022 1834 5037 1838
rect 5055 1835 5094 1854
rect 5113 1848 5120 1849
rect 5119 1841 5120 1848
rect 5103 1838 5104 1841
rect 5119 1838 5132 1841
rect 5055 1834 5085 1835
rect 5094 1834 5100 1835
rect 5103 1834 5132 1838
rect 5022 1833 5132 1834
rect 5022 1832 5138 1833
rect 4697 1824 4748 1832
rect 4697 1812 4722 1824
rect 4729 1812 4748 1824
rect 4779 1824 4829 1832
rect 4779 1816 4795 1824
rect 4802 1822 4829 1824
rect 4838 1822 5059 1832
rect 4802 1812 5059 1822
rect 5088 1824 5138 1832
rect 5088 1815 5104 1824
rect 4697 1804 4748 1812
rect 4795 1804 5059 1812
rect 5085 1812 5104 1815
rect 5111 1812 5138 1824
rect 5085 1804 5138 1812
rect 4713 1796 4714 1804
rect 4729 1796 4742 1804
rect 4713 1788 4729 1796
rect 4710 1781 4729 1784
rect 4710 1772 4732 1781
rect 4683 1762 4732 1772
rect 4683 1756 4713 1762
rect 4732 1757 4737 1762
rect 4655 1740 4729 1756
rect 4747 1748 4777 1804
rect 4812 1794 5020 1804
rect 5055 1800 5100 1804
rect 5103 1803 5104 1804
rect 5119 1803 5132 1804
rect 4838 1764 5027 1794
rect 4853 1761 5027 1764
rect 4846 1758 5027 1761
rect 4655 1738 4668 1740
rect 4683 1738 4717 1740
rect 4655 1722 4729 1738
rect 4756 1734 4769 1748
rect 4784 1734 4800 1750
rect 4846 1745 4857 1758
rect 4639 1700 4640 1716
rect 4655 1700 4668 1722
rect 4683 1700 4713 1722
rect 4756 1718 4818 1734
rect 4846 1727 4857 1743
rect 4862 1738 4872 1758
rect 4882 1738 4896 1758
rect 4899 1745 4908 1758
rect 4924 1745 4933 1758
rect 4862 1727 4896 1738
rect 4899 1727 4908 1743
rect 4924 1727 4933 1743
rect 4940 1738 4950 1758
rect 4960 1738 4974 1758
rect 4975 1745 4986 1758
rect 4940 1727 4974 1738
rect 4975 1727 4986 1743
rect 5032 1734 5048 1750
rect 5055 1748 5085 1800
rect 5119 1796 5120 1803
rect 5104 1788 5120 1796
rect 5091 1756 5104 1775
rect 5119 1756 5149 1772
rect 5091 1740 5165 1756
rect 5091 1738 5104 1740
rect 5119 1738 5153 1740
rect 4756 1716 4769 1718
rect 4784 1716 4818 1718
rect 4756 1700 4818 1716
rect 4862 1711 4878 1714
rect 4940 1711 4970 1722
rect 5018 1718 5064 1734
rect 5091 1722 5165 1738
rect 5018 1716 5052 1718
rect 5017 1700 5064 1716
rect 5091 1700 5104 1722
rect 5119 1700 5149 1722
rect 5176 1700 5177 1716
rect 5192 1700 5205 1860
rect 5235 1756 5248 1860
rect 5293 1838 5294 1848
rect 5309 1838 5322 1848
rect 5293 1834 5322 1838
rect 5327 1834 5357 1860
rect 5375 1846 5391 1848
rect 5463 1846 5516 1860
rect 5464 1844 5528 1846
rect 5571 1844 5586 1860
rect 5635 1857 5665 1860
rect 5635 1854 5671 1857
rect 5601 1846 5617 1848
rect 5375 1834 5390 1838
rect 5293 1832 5390 1834
rect 5418 1832 5586 1844
rect 5602 1834 5617 1838
rect 5635 1835 5674 1854
rect 5693 1848 5700 1849
rect 5699 1841 5700 1848
rect 5683 1838 5684 1841
rect 5699 1838 5712 1841
rect 5635 1834 5665 1835
rect 5674 1834 5680 1835
rect 5683 1834 5712 1838
rect 5602 1833 5712 1834
rect 5602 1832 5718 1833
rect 5277 1824 5328 1832
rect 5277 1812 5302 1824
rect 5309 1812 5328 1824
rect 5359 1824 5409 1832
rect 5359 1816 5375 1824
rect 5382 1822 5409 1824
rect 5418 1822 5639 1832
rect 5382 1812 5639 1822
rect 5668 1824 5718 1832
rect 5668 1815 5684 1824
rect 5277 1804 5328 1812
rect 5375 1804 5639 1812
rect 5665 1812 5684 1815
rect 5691 1812 5718 1824
rect 5665 1804 5718 1812
rect 5293 1796 5294 1804
rect 5309 1796 5322 1804
rect 5293 1788 5309 1796
rect 5290 1781 5309 1784
rect 5290 1772 5312 1781
rect 5263 1762 5312 1772
rect 5263 1756 5293 1762
rect 5312 1757 5317 1762
rect 5235 1740 5309 1756
rect 5327 1748 5357 1804
rect 5392 1794 5600 1804
rect 5635 1800 5680 1804
rect 5683 1803 5684 1804
rect 5699 1803 5712 1804
rect 5418 1764 5607 1794
rect 5433 1761 5607 1764
rect 5426 1758 5607 1761
rect 5235 1738 5248 1740
rect 5263 1738 5297 1740
rect 5235 1722 5309 1738
rect 5336 1734 5349 1748
rect 5364 1734 5380 1750
rect 5426 1745 5437 1758
rect 5219 1700 5220 1716
rect 5235 1700 5248 1722
rect 5263 1700 5293 1722
rect 5336 1718 5398 1734
rect 5426 1727 5437 1743
rect 5442 1738 5452 1758
rect 5462 1738 5476 1758
rect 5479 1745 5488 1758
rect 5504 1745 5513 1758
rect 5442 1727 5476 1738
rect 5479 1727 5488 1743
rect 5504 1727 5513 1743
rect 5520 1738 5530 1758
rect 5540 1738 5554 1758
rect 5555 1745 5566 1758
rect 5520 1727 5554 1738
rect 5555 1727 5566 1743
rect 5612 1734 5628 1750
rect 5635 1748 5665 1800
rect 5699 1796 5700 1803
rect 5684 1788 5700 1796
rect 5671 1756 5684 1775
rect 5699 1756 5729 1772
rect 5671 1740 5745 1756
rect 5671 1738 5684 1740
rect 5699 1738 5733 1740
rect 5336 1716 5349 1718
rect 5364 1716 5398 1718
rect 5336 1700 5398 1716
rect 5442 1711 5458 1714
rect 5520 1711 5550 1722
rect 5598 1718 5644 1734
rect 5671 1722 5745 1738
rect 5598 1716 5632 1718
rect 5597 1700 5644 1716
rect 5671 1700 5684 1722
rect 5699 1700 5729 1722
rect 5756 1700 5757 1716
rect 5772 1700 5785 1860
rect 5815 1756 5828 1860
rect 5873 1838 5874 1848
rect 5889 1838 5902 1848
rect 5873 1834 5902 1838
rect 5907 1834 5937 1860
rect 5955 1846 5971 1848
rect 6043 1846 6096 1860
rect 6044 1844 6108 1846
rect 6151 1844 6166 1860
rect 6215 1857 6245 1860
rect 6215 1854 6251 1857
rect 6181 1846 6197 1848
rect 5955 1834 5970 1838
rect 5873 1832 5970 1834
rect 5998 1832 6166 1844
rect 6182 1834 6197 1838
rect 6215 1835 6254 1854
rect 6273 1848 6280 1849
rect 6279 1841 6280 1848
rect 6263 1838 6264 1841
rect 6279 1838 6292 1841
rect 6215 1834 6245 1835
rect 6254 1834 6260 1835
rect 6263 1834 6292 1838
rect 6182 1833 6292 1834
rect 6182 1832 6298 1833
rect 5857 1824 5908 1832
rect 5857 1812 5882 1824
rect 5889 1812 5908 1824
rect 5939 1824 5989 1832
rect 5939 1816 5955 1824
rect 5962 1822 5989 1824
rect 5998 1822 6219 1832
rect 5962 1812 6219 1822
rect 6248 1824 6298 1832
rect 6248 1815 6264 1824
rect 5857 1804 5908 1812
rect 5955 1804 6219 1812
rect 6245 1812 6264 1815
rect 6271 1812 6298 1824
rect 6245 1804 6298 1812
rect 5873 1796 5874 1804
rect 5889 1796 5902 1804
rect 5873 1788 5889 1796
rect 5870 1781 5889 1784
rect 5870 1772 5892 1781
rect 5843 1762 5892 1772
rect 5843 1756 5873 1762
rect 5892 1757 5897 1762
rect 5815 1740 5889 1756
rect 5907 1748 5937 1804
rect 5972 1794 6180 1804
rect 6215 1800 6260 1804
rect 6263 1803 6264 1804
rect 6279 1803 6292 1804
rect 5998 1764 6187 1794
rect 6013 1761 6187 1764
rect 6006 1758 6187 1761
rect 5815 1738 5828 1740
rect 5843 1738 5877 1740
rect 5815 1722 5889 1738
rect 5916 1734 5929 1748
rect 5944 1734 5960 1750
rect 6006 1745 6017 1758
rect 5799 1700 5800 1716
rect 5815 1700 5828 1722
rect 5843 1700 5873 1722
rect 5916 1718 5978 1734
rect 6006 1727 6017 1743
rect 6022 1738 6032 1758
rect 6042 1738 6056 1758
rect 6059 1745 6068 1758
rect 6084 1745 6093 1758
rect 6022 1727 6056 1738
rect 6059 1727 6068 1743
rect 6084 1727 6093 1743
rect 6100 1738 6110 1758
rect 6120 1738 6134 1758
rect 6135 1745 6146 1758
rect 6100 1727 6134 1738
rect 6135 1727 6146 1743
rect 6192 1734 6208 1750
rect 6215 1748 6245 1800
rect 6279 1796 6280 1803
rect 6264 1788 6280 1796
rect 6251 1756 6264 1775
rect 6279 1756 6309 1772
rect 6251 1740 6325 1756
rect 6251 1738 6264 1740
rect 6279 1738 6313 1740
rect 5916 1716 5929 1718
rect 5944 1716 5978 1718
rect 5916 1700 5978 1716
rect 6022 1711 6038 1714
rect 6100 1711 6130 1722
rect 6178 1718 6224 1734
rect 6251 1722 6325 1738
rect 6178 1716 6212 1718
rect 6177 1700 6224 1716
rect 6251 1700 6264 1722
rect 6279 1700 6309 1722
rect 6336 1700 6337 1716
rect 6352 1700 6365 1860
rect 6395 1756 6408 1860
rect 6453 1838 6454 1848
rect 6469 1838 6482 1848
rect 6453 1834 6482 1838
rect 6487 1834 6517 1860
rect 6535 1846 6551 1848
rect 6623 1846 6676 1860
rect 6624 1844 6688 1846
rect 6731 1844 6746 1860
rect 6795 1857 6825 1860
rect 6795 1854 6831 1857
rect 6761 1846 6777 1848
rect 6535 1834 6550 1838
rect 6453 1832 6550 1834
rect 6578 1832 6746 1844
rect 6762 1834 6777 1838
rect 6795 1835 6834 1854
rect 6853 1848 6860 1849
rect 6859 1841 6860 1848
rect 6843 1838 6844 1841
rect 6859 1838 6872 1841
rect 6795 1834 6825 1835
rect 6834 1834 6840 1835
rect 6843 1834 6872 1838
rect 6762 1833 6872 1834
rect 6762 1832 6878 1833
rect 6437 1824 6488 1832
rect 6437 1812 6462 1824
rect 6469 1812 6488 1824
rect 6519 1824 6569 1832
rect 6519 1816 6535 1824
rect 6542 1822 6569 1824
rect 6578 1822 6799 1832
rect 6542 1812 6799 1822
rect 6828 1824 6878 1832
rect 6828 1815 6844 1824
rect 6437 1804 6488 1812
rect 6535 1804 6799 1812
rect 6825 1812 6844 1815
rect 6851 1812 6878 1824
rect 6825 1804 6878 1812
rect 6453 1796 6454 1804
rect 6469 1796 6482 1804
rect 6453 1788 6469 1796
rect 6450 1781 6469 1784
rect 6450 1772 6472 1781
rect 6423 1762 6472 1772
rect 6423 1756 6453 1762
rect 6472 1757 6477 1762
rect 6395 1740 6469 1756
rect 6487 1748 6517 1804
rect 6552 1794 6760 1804
rect 6795 1800 6840 1804
rect 6843 1803 6844 1804
rect 6859 1803 6872 1804
rect 6578 1764 6767 1794
rect 6593 1761 6767 1764
rect 6586 1758 6767 1761
rect 6395 1738 6408 1740
rect 6423 1738 6457 1740
rect 6395 1722 6469 1738
rect 6496 1734 6509 1748
rect 6524 1734 6540 1750
rect 6586 1745 6597 1758
rect 6379 1700 6380 1716
rect 6395 1700 6408 1722
rect 6423 1700 6453 1722
rect 6496 1718 6558 1734
rect 6586 1727 6597 1743
rect 6602 1738 6612 1758
rect 6622 1738 6636 1758
rect 6639 1745 6648 1758
rect 6664 1745 6673 1758
rect 6602 1727 6636 1738
rect 6639 1727 6648 1743
rect 6664 1727 6673 1743
rect 6680 1738 6690 1758
rect 6700 1738 6714 1758
rect 6715 1745 6726 1758
rect 6680 1727 6714 1738
rect 6715 1727 6726 1743
rect 6772 1734 6788 1750
rect 6795 1748 6825 1800
rect 6859 1796 6860 1803
rect 6844 1788 6860 1796
rect 6831 1756 6844 1775
rect 6859 1756 6889 1772
rect 6831 1740 6905 1756
rect 6831 1738 6844 1740
rect 6859 1738 6893 1740
rect 6496 1716 6509 1718
rect 6524 1716 6558 1718
rect 6496 1700 6558 1716
rect 6602 1711 6618 1714
rect 6680 1711 6710 1722
rect 6758 1718 6804 1734
rect 6831 1722 6905 1738
rect 6758 1716 6792 1718
rect 6757 1700 6804 1716
rect 6831 1700 6844 1722
rect 6859 1700 6889 1722
rect 6916 1700 6917 1716
rect 6932 1700 6945 1860
rect 6975 1756 6988 1860
rect 7033 1838 7034 1848
rect 7049 1838 7062 1848
rect 7033 1834 7062 1838
rect 7067 1834 7097 1860
rect 7115 1846 7131 1848
rect 7203 1846 7256 1860
rect 7204 1844 7268 1846
rect 7311 1844 7326 1860
rect 7375 1857 7405 1860
rect 7375 1854 7411 1857
rect 7341 1846 7357 1848
rect 7115 1834 7130 1838
rect 7033 1832 7130 1834
rect 7158 1832 7326 1844
rect 7342 1834 7357 1838
rect 7375 1835 7414 1854
rect 7433 1848 7440 1849
rect 7439 1841 7440 1848
rect 7423 1838 7424 1841
rect 7439 1838 7452 1841
rect 7375 1834 7405 1835
rect 7414 1834 7420 1835
rect 7423 1834 7452 1838
rect 7342 1833 7452 1834
rect 7342 1832 7458 1833
rect 7017 1824 7068 1832
rect 7017 1812 7042 1824
rect 7049 1812 7068 1824
rect 7099 1824 7149 1832
rect 7099 1816 7115 1824
rect 7122 1822 7149 1824
rect 7158 1822 7379 1832
rect 7122 1812 7379 1822
rect 7408 1824 7458 1832
rect 7408 1815 7424 1824
rect 7017 1804 7068 1812
rect 7115 1804 7379 1812
rect 7405 1812 7424 1815
rect 7431 1812 7458 1824
rect 7405 1804 7458 1812
rect 7033 1796 7034 1804
rect 7049 1796 7062 1804
rect 7033 1788 7049 1796
rect 7030 1781 7049 1784
rect 7030 1772 7052 1781
rect 7003 1762 7052 1772
rect 7003 1756 7033 1762
rect 7052 1757 7057 1762
rect 6975 1740 7049 1756
rect 7067 1748 7097 1804
rect 7132 1794 7340 1804
rect 7375 1800 7420 1804
rect 7423 1803 7424 1804
rect 7439 1803 7452 1804
rect 7158 1764 7347 1794
rect 7173 1761 7347 1764
rect 7166 1758 7347 1761
rect 6975 1738 6988 1740
rect 7003 1738 7037 1740
rect 6975 1722 7049 1738
rect 7076 1734 7089 1748
rect 7104 1734 7120 1750
rect 7166 1745 7177 1758
rect 6959 1700 6960 1716
rect 6975 1700 6988 1722
rect 7003 1700 7033 1722
rect 7076 1718 7138 1734
rect 7166 1727 7177 1743
rect 7182 1738 7192 1758
rect 7202 1738 7216 1758
rect 7219 1745 7228 1758
rect 7244 1745 7253 1758
rect 7182 1727 7216 1738
rect 7219 1727 7228 1743
rect 7244 1727 7253 1743
rect 7260 1738 7270 1758
rect 7280 1738 7294 1758
rect 7295 1745 7306 1758
rect 7260 1727 7294 1738
rect 7295 1727 7306 1743
rect 7352 1734 7368 1750
rect 7375 1748 7405 1800
rect 7439 1796 7440 1803
rect 7424 1788 7440 1796
rect 7411 1756 7424 1775
rect 7439 1756 7469 1772
rect 7411 1740 7485 1756
rect 7411 1738 7424 1740
rect 7439 1738 7473 1740
rect 7076 1716 7089 1718
rect 7104 1716 7138 1718
rect 7076 1700 7138 1716
rect 7182 1711 7198 1714
rect 7260 1711 7290 1722
rect 7338 1718 7384 1734
rect 7411 1722 7485 1738
rect 7338 1716 7372 1718
rect 7337 1700 7384 1716
rect 7411 1700 7424 1722
rect 7439 1700 7469 1722
rect 7496 1700 7497 1716
rect 7512 1700 7525 1860
rect 7555 1756 7568 1860
rect 7613 1838 7614 1848
rect 7629 1838 7642 1848
rect 7613 1834 7642 1838
rect 7647 1834 7677 1860
rect 7695 1846 7711 1848
rect 7783 1846 7836 1860
rect 7784 1844 7848 1846
rect 7891 1844 7906 1860
rect 7955 1857 7985 1860
rect 7955 1854 7991 1857
rect 7921 1846 7937 1848
rect 7695 1834 7710 1838
rect 7613 1832 7710 1834
rect 7738 1832 7906 1844
rect 7922 1834 7937 1838
rect 7955 1835 7994 1854
rect 8013 1848 8020 1849
rect 8019 1841 8020 1848
rect 8003 1838 8004 1841
rect 8019 1838 8032 1841
rect 7955 1834 7985 1835
rect 7994 1834 8000 1835
rect 8003 1834 8032 1838
rect 7922 1833 8032 1834
rect 7922 1832 8038 1833
rect 7597 1824 7648 1832
rect 7597 1812 7622 1824
rect 7629 1812 7648 1824
rect 7679 1824 7729 1832
rect 7679 1816 7695 1824
rect 7702 1822 7729 1824
rect 7738 1822 7959 1832
rect 7702 1812 7959 1822
rect 7988 1824 8038 1832
rect 7988 1815 8004 1824
rect 7597 1804 7648 1812
rect 7695 1804 7959 1812
rect 7985 1812 8004 1815
rect 8011 1812 8038 1824
rect 7985 1804 8038 1812
rect 7613 1796 7614 1804
rect 7629 1796 7642 1804
rect 7613 1788 7629 1796
rect 7610 1781 7629 1784
rect 7610 1772 7632 1781
rect 7583 1762 7632 1772
rect 7583 1756 7613 1762
rect 7632 1757 7637 1762
rect 7555 1740 7629 1756
rect 7647 1748 7677 1804
rect 7712 1794 7920 1804
rect 7955 1800 8000 1804
rect 8003 1803 8004 1804
rect 8019 1803 8032 1804
rect 7738 1764 7927 1794
rect 7753 1761 7927 1764
rect 7746 1758 7927 1761
rect 7555 1738 7568 1740
rect 7583 1738 7617 1740
rect 7555 1722 7629 1738
rect 7656 1734 7669 1748
rect 7684 1734 7700 1750
rect 7746 1745 7757 1758
rect 7539 1700 7540 1716
rect 7555 1700 7568 1722
rect 7583 1700 7613 1722
rect 7656 1718 7718 1734
rect 7746 1727 7757 1743
rect 7762 1738 7772 1758
rect 7782 1738 7796 1758
rect 7799 1745 7808 1758
rect 7824 1745 7833 1758
rect 7762 1727 7796 1738
rect 7799 1727 7808 1743
rect 7824 1727 7833 1743
rect 7840 1738 7850 1758
rect 7860 1738 7874 1758
rect 7875 1745 7886 1758
rect 7840 1727 7874 1738
rect 7875 1727 7886 1743
rect 7932 1734 7948 1750
rect 7955 1748 7985 1800
rect 8019 1796 8020 1803
rect 8004 1788 8020 1796
rect 7991 1756 8004 1775
rect 8019 1756 8049 1772
rect 7991 1740 8065 1756
rect 7991 1738 8004 1740
rect 8019 1738 8053 1740
rect 7656 1716 7669 1718
rect 7684 1716 7718 1718
rect 7656 1700 7718 1716
rect 7762 1711 7778 1714
rect 7840 1711 7870 1722
rect 7918 1718 7964 1734
rect 7991 1722 8065 1738
rect 7918 1716 7952 1718
rect 7917 1700 7964 1716
rect 7991 1700 8004 1722
rect 8019 1700 8049 1722
rect 8076 1700 8077 1716
rect 8092 1700 8105 1860
rect 8135 1756 8148 1860
rect 8193 1838 8194 1848
rect 8209 1838 8222 1848
rect 8193 1834 8222 1838
rect 8227 1834 8257 1860
rect 8275 1846 8291 1848
rect 8363 1846 8416 1860
rect 8364 1844 8428 1846
rect 8471 1844 8486 1860
rect 8535 1857 8565 1860
rect 8535 1854 8571 1857
rect 8501 1846 8517 1848
rect 8275 1834 8290 1838
rect 8193 1832 8290 1834
rect 8318 1832 8486 1844
rect 8502 1834 8517 1838
rect 8535 1835 8574 1854
rect 8593 1848 8600 1849
rect 8599 1841 8600 1848
rect 8583 1838 8584 1841
rect 8599 1838 8612 1841
rect 8535 1834 8565 1835
rect 8574 1834 8580 1835
rect 8583 1834 8612 1838
rect 8502 1833 8612 1834
rect 8502 1832 8618 1833
rect 8177 1824 8228 1832
rect 8177 1812 8202 1824
rect 8209 1812 8228 1824
rect 8259 1824 8309 1832
rect 8259 1816 8275 1824
rect 8282 1822 8309 1824
rect 8318 1822 8539 1832
rect 8282 1812 8539 1822
rect 8568 1824 8618 1832
rect 8568 1815 8584 1824
rect 8177 1804 8228 1812
rect 8275 1804 8539 1812
rect 8565 1812 8584 1815
rect 8591 1812 8618 1824
rect 8565 1804 8618 1812
rect 8193 1796 8194 1804
rect 8209 1796 8222 1804
rect 8193 1788 8209 1796
rect 8190 1781 8209 1784
rect 8190 1772 8212 1781
rect 8163 1762 8212 1772
rect 8163 1756 8193 1762
rect 8212 1757 8217 1762
rect 8135 1740 8209 1756
rect 8227 1748 8257 1804
rect 8292 1794 8500 1804
rect 8535 1800 8580 1804
rect 8583 1803 8584 1804
rect 8599 1803 8612 1804
rect 8318 1764 8507 1794
rect 8333 1761 8507 1764
rect 8326 1758 8507 1761
rect 8135 1738 8148 1740
rect 8163 1738 8197 1740
rect 8135 1722 8209 1738
rect 8236 1734 8249 1748
rect 8264 1734 8280 1750
rect 8326 1745 8337 1758
rect 8119 1700 8120 1716
rect 8135 1700 8148 1722
rect 8163 1700 8193 1722
rect 8236 1718 8298 1734
rect 8326 1727 8337 1743
rect 8342 1738 8352 1758
rect 8362 1738 8376 1758
rect 8379 1745 8388 1758
rect 8404 1745 8413 1758
rect 8342 1727 8376 1738
rect 8379 1727 8388 1743
rect 8404 1727 8413 1743
rect 8420 1738 8430 1758
rect 8440 1738 8454 1758
rect 8455 1745 8466 1758
rect 8420 1727 8454 1738
rect 8455 1727 8466 1743
rect 8512 1734 8528 1750
rect 8535 1748 8565 1800
rect 8599 1796 8600 1803
rect 8584 1788 8600 1796
rect 8571 1756 8584 1775
rect 8599 1756 8629 1772
rect 8571 1740 8645 1756
rect 8571 1738 8584 1740
rect 8599 1738 8633 1740
rect 8236 1716 8249 1718
rect 8264 1716 8298 1718
rect 8236 1700 8298 1716
rect 8342 1711 8358 1714
rect 8420 1711 8450 1722
rect 8498 1718 8544 1734
rect 8571 1722 8645 1738
rect 8498 1716 8532 1718
rect 8497 1700 8544 1716
rect 8571 1700 8584 1722
rect 8599 1700 8629 1722
rect 8656 1700 8657 1716
rect 8672 1700 8685 1860
rect 8715 1756 8728 1860
rect 8773 1838 8774 1848
rect 8789 1838 8802 1848
rect 8773 1834 8802 1838
rect 8807 1834 8837 1860
rect 8855 1846 8871 1848
rect 8943 1846 8996 1860
rect 8944 1844 9008 1846
rect 9051 1844 9066 1860
rect 9115 1857 9145 1860
rect 9115 1854 9151 1857
rect 9081 1846 9097 1848
rect 8855 1834 8870 1838
rect 8773 1832 8870 1834
rect 8898 1832 9066 1844
rect 9082 1834 9097 1838
rect 9115 1835 9154 1854
rect 9173 1848 9180 1849
rect 9179 1841 9180 1848
rect 9163 1838 9164 1841
rect 9179 1838 9192 1841
rect 9115 1834 9145 1835
rect 9154 1834 9160 1835
rect 9163 1834 9192 1838
rect 9082 1833 9192 1834
rect 9082 1832 9198 1833
rect 8757 1824 8808 1832
rect 8757 1812 8782 1824
rect 8789 1812 8808 1824
rect 8839 1824 8889 1832
rect 8839 1816 8855 1824
rect 8862 1822 8889 1824
rect 8898 1822 9119 1832
rect 8862 1812 9119 1822
rect 9148 1824 9198 1832
rect 9148 1815 9164 1824
rect 8757 1804 8808 1812
rect 8855 1804 9119 1812
rect 9145 1812 9164 1815
rect 9171 1812 9198 1824
rect 9145 1804 9198 1812
rect 8773 1796 8774 1804
rect 8789 1796 8802 1804
rect 8773 1788 8789 1796
rect 8770 1781 8789 1784
rect 8770 1772 8792 1781
rect 8743 1762 8792 1772
rect 8743 1756 8773 1762
rect 8792 1757 8797 1762
rect 8715 1740 8789 1756
rect 8807 1748 8837 1804
rect 8872 1794 9080 1804
rect 9115 1800 9160 1804
rect 9163 1803 9164 1804
rect 9179 1803 9192 1804
rect 8898 1764 9087 1794
rect 8913 1761 9087 1764
rect 8906 1758 9087 1761
rect 8715 1738 8728 1740
rect 8743 1738 8777 1740
rect 8715 1722 8789 1738
rect 8816 1734 8829 1748
rect 8844 1734 8860 1750
rect 8906 1745 8917 1758
rect 8699 1700 8700 1716
rect 8715 1700 8728 1722
rect 8743 1700 8773 1722
rect 8816 1718 8878 1734
rect 8906 1727 8917 1743
rect 8922 1738 8932 1758
rect 8942 1738 8956 1758
rect 8959 1745 8968 1758
rect 8984 1745 8993 1758
rect 8922 1727 8956 1738
rect 8959 1727 8968 1743
rect 8984 1727 8993 1743
rect 9000 1738 9010 1758
rect 9020 1738 9034 1758
rect 9035 1745 9046 1758
rect 9000 1727 9034 1738
rect 9035 1727 9046 1743
rect 9092 1734 9108 1750
rect 9115 1748 9145 1800
rect 9179 1796 9180 1803
rect 9164 1788 9180 1796
rect 9151 1756 9164 1775
rect 9179 1756 9209 1772
rect 9151 1740 9225 1756
rect 9151 1738 9164 1740
rect 9179 1738 9213 1740
rect 8816 1716 8829 1718
rect 8844 1716 8878 1718
rect 8816 1700 8878 1716
rect 8922 1711 8938 1714
rect 9000 1711 9030 1722
rect 9078 1718 9124 1734
rect 9151 1722 9225 1738
rect 9078 1716 9112 1718
rect 9077 1700 9124 1716
rect 9151 1700 9164 1722
rect 9179 1700 9209 1722
rect 9236 1700 9237 1716
rect 9252 1700 9265 1860
rect -7 1692 34 1700
rect -7 1666 8 1692
rect 15 1666 34 1692
rect 98 1688 160 1700
rect 172 1688 247 1700
rect 305 1688 380 1700
rect 392 1688 423 1700
rect 429 1688 464 1700
rect 98 1686 260 1688
rect -7 1658 34 1666
rect 116 1662 129 1686
rect 144 1684 159 1686
rect -1 1648 0 1658
rect 15 1648 28 1658
rect 43 1648 73 1662
rect 116 1648 159 1662
rect 183 1659 190 1666
rect 193 1662 260 1686
rect 292 1686 464 1688
rect 262 1664 290 1668
rect 292 1664 372 1686
rect 393 1684 408 1686
rect 262 1662 372 1664
rect 193 1658 372 1662
rect 166 1648 196 1658
rect 198 1648 351 1658
rect 359 1648 389 1658
rect 393 1648 423 1662
rect 451 1648 464 1686
rect 536 1692 571 1700
rect 536 1666 537 1692
rect 544 1666 571 1692
rect 479 1648 509 1662
rect 536 1658 571 1666
rect 573 1692 614 1700
rect 573 1666 588 1692
rect 595 1666 614 1692
rect 678 1688 740 1700
rect 752 1688 827 1700
rect 885 1688 960 1700
rect 972 1688 1003 1700
rect 1009 1688 1044 1700
rect 678 1686 840 1688
rect 573 1658 614 1666
rect 696 1662 709 1686
rect 724 1684 739 1686
rect 536 1648 537 1658
rect 552 1648 565 1658
rect 579 1648 580 1658
rect 595 1648 608 1658
rect 623 1648 653 1662
rect 696 1648 739 1662
rect 763 1659 770 1666
rect 773 1662 840 1686
rect 872 1686 1044 1688
rect 842 1664 870 1668
rect 872 1664 952 1686
rect 973 1684 988 1686
rect 842 1662 952 1664
rect 773 1658 952 1662
rect 746 1648 776 1658
rect 778 1648 931 1658
rect 939 1648 969 1658
rect 973 1648 1003 1662
rect 1031 1648 1044 1686
rect 1116 1692 1151 1700
rect 1116 1666 1117 1692
rect 1124 1666 1151 1692
rect 1059 1648 1089 1662
rect 1116 1658 1151 1666
rect 1153 1692 1194 1700
rect 1153 1666 1168 1692
rect 1175 1666 1194 1692
rect 1258 1688 1320 1700
rect 1332 1688 1407 1700
rect 1465 1688 1540 1700
rect 1552 1688 1583 1700
rect 1589 1688 1624 1700
rect 1258 1686 1420 1688
rect 1153 1658 1194 1666
rect 1276 1662 1289 1686
rect 1304 1684 1319 1686
rect 1116 1648 1117 1658
rect 1132 1648 1145 1658
rect 1159 1648 1160 1658
rect 1175 1648 1188 1658
rect 1203 1648 1233 1662
rect 1276 1648 1319 1662
rect 1343 1659 1350 1666
rect 1353 1662 1420 1686
rect 1452 1686 1624 1688
rect 1422 1664 1450 1668
rect 1452 1664 1532 1686
rect 1553 1684 1568 1686
rect 1422 1662 1532 1664
rect 1353 1658 1532 1662
rect 1326 1648 1356 1658
rect 1358 1648 1511 1658
rect 1519 1648 1549 1658
rect 1553 1648 1583 1662
rect 1611 1648 1624 1686
rect 1696 1692 1731 1700
rect 1696 1666 1697 1692
rect 1704 1666 1731 1692
rect 1639 1648 1669 1662
rect 1696 1658 1731 1666
rect 1733 1692 1774 1700
rect 1733 1666 1748 1692
rect 1755 1666 1774 1692
rect 1838 1688 1900 1700
rect 1912 1688 1987 1700
rect 2045 1688 2120 1700
rect 2132 1688 2163 1700
rect 2169 1688 2204 1700
rect 1838 1686 2000 1688
rect 1733 1658 1774 1666
rect 1856 1662 1869 1686
rect 1884 1684 1899 1686
rect 1696 1648 1697 1658
rect 1712 1648 1725 1658
rect 1739 1648 1740 1658
rect 1755 1648 1768 1658
rect 1783 1648 1813 1662
rect 1856 1648 1899 1662
rect 1923 1659 1930 1666
rect 1933 1662 2000 1686
rect 2032 1686 2204 1688
rect 2002 1664 2030 1668
rect 2032 1664 2112 1686
rect 2133 1684 2148 1686
rect 2002 1662 2112 1664
rect 1933 1658 2112 1662
rect 1906 1648 1936 1658
rect 1938 1648 2091 1658
rect 2099 1648 2129 1658
rect 2133 1648 2163 1662
rect 2191 1648 2204 1686
rect 2276 1692 2311 1700
rect 2276 1666 2277 1692
rect 2284 1666 2311 1692
rect 2219 1648 2249 1662
rect 2276 1658 2311 1666
rect 2313 1692 2354 1700
rect 2313 1666 2328 1692
rect 2335 1666 2354 1692
rect 2418 1688 2480 1700
rect 2492 1688 2567 1700
rect 2625 1688 2700 1700
rect 2712 1688 2743 1700
rect 2749 1688 2784 1700
rect 2418 1686 2580 1688
rect 2313 1658 2354 1666
rect 2436 1662 2449 1686
rect 2464 1684 2479 1686
rect 2276 1648 2277 1658
rect 2292 1648 2305 1658
rect 2319 1648 2320 1658
rect 2335 1648 2348 1658
rect 2363 1648 2393 1662
rect 2436 1648 2479 1662
rect 2503 1659 2510 1666
rect 2513 1662 2580 1686
rect 2612 1686 2784 1688
rect 2582 1664 2610 1668
rect 2612 1664 2692 1686
rect 2713 1684 2728 1686
rect 2582 1662 2692 1664
rect 2513 1658 2692 1662
rect 2486 1648 2516 1658
rect 2518 1648 2671 1658
rect 2679 1648 2709 1658
rect 2713 1648 2743 1662
rect 2771 1648 2784 1686
rect 2856 1692 2891 1700
rect 2856 1666 2857 1692
rect 2864 1666 2891 1692
rect 2799 1648 2829 1662
rect 2856 1658 2891 1666
rect 2893 1692 2934 1700
rect 2893 1666 2908 1692
rect 2915 1666 2934 1692
rect 2998 1688 3060 1700
rect 3072 1688 3147 1700
rect 3205 1688 3280 1700
rect 3292 1688 3323 1700
rect 3329 1688 3364 1700
rect 2998 1686 3160 1688
rect 2893 1658 2934 1666
rect 3016 1662 3029 1686
rect 3044 1684 3059 1686
rect 2856 1648 2857 1658
rect 2872 1648 2885 1658
rect 2899 1648 2900 1658
rect 2915 1648 2928 1658
rect 2943 1648 2973 1662
rect 3016 1648 3059 1662
rect 3083 1659 3090 1666
rect 3093 1662 3160 1686
rect 3192 1686 3364 1688
rect 3162 1664 3190 1668
rect 3192 1664 3272 1686
rect 3293 1684 3308 1686
rect 3162 1662 3272 1664
rect 3093 1658 3272 1662
rect 3066 1648 3096 1658
rect 3098 1648 3251 1658
rect 3259 1648 3289 1658
rect 3293 1648 3323 1662
rect 3351 1648 3364 1686
rect 3436 1692 3471 1700
rect 3436 1666 3437 1692
rect 3444 1666 3471 1692
rect 3379 1648 3409 1662
rect 3436 1658 3471 1666
rect 3473 1692 3514 1700
rect 3473 1666 3488 1692
rect 3495 1666 3514 1692
rect 3578 1688 3640 1700
rect 3652 1688 3727 1700
rect 3785 1688 3860 1700
rect 3872 1688 3903 1700
rect 3909 1688 3944 1700
rect 3578 1686 3740 1688
rect 3473 1658 3514 1666
rect 3596 1662 3609 1686
rect 3624 1684 3639 1686
rect 3436 1648 3437 1658
rect 3452 1648 3465 1658
rect 3479 1648 3480 1658
rect 3495 1648 3508 1658
rect 3523 1648 3553 1662
rect 3596 1648 3639 1662
rect 3663 1659 3670 1666
rect 3673 1662 3740 1686
rect 3772 1686 3944 1688
rect 3742 1664 3770 1668
rect 3772 1664 3852 1686
rect 3873 1684 3888 1686
rect 3742 1662 3852 1664
rect 3673 1658 3852 1662
rect 3646 1648 3676 1658
rect 3678 1648 3831 1658
rect 3839 1648 3869 1658
rect 3873 1648 3903 1662
rect 3931 1648 3944 1686
rect 4016 1692 4051 1700
rect 4016 1666 4017 1692
rect 4024 1666 4051 1692
rect 3959 1648 3989 1662
rect 4016 1658 4051 1666
rect 4053 1692 4094 1700
rect 4053 1666 4068 1692
rect 4075 1666 4094 1692
rect 4158 1688 4220 1700
rect 4232 1688 4307 1700
rect 4365 1688 4440 1700
rect 4452 1688 4483 1700
rect 4489 1688 4524 1700
rect 4158 1686 4320 1688
rect 4053 1658 4094 1666
rect 4176 1662 4189 1686
rect 4204 1684 4219 1686
rect 4016 1648 4017 1658
rect 4032 1648 4045 1658
rect 4059 1648 4060 1658
rect 4075 1648 4088 1658
rect 4103 1648 4133 1662
rect 4176 1648 4219 1662
rect 4243 1659 4250 1666
rect 4253 1662 4320 1686
rect 4352 1686 4524 1688
rect 4322 1664 4350 1668
rect 4352 1664 4432 1686
rect 4453 1684 4468 1686
rect 4322 1662 4432 1664
rect 4253 1658 4432 1662
rect 4226 1648 4256 1658
rect 4258 1648 4411 1658
rect 4419 1648 4449 1658
rect 4453 1648 4483 1662
rect 4511 1648 4524 1686
rect 4596 1692 4631 1700
rect 4596 1666 4597 1692
rect 4604 1666 4631 1692
rect 4539 1648 4569 1662
rect 4596 1658 4631 1666
rect 4633 1692 4674 1700
rect 4633 1666 4648 1692
rect 4655 1666 4674 1692
rect 4738 1688 4800 1700
rect 4812 1688 4887 1700
rect 4945 1688 5020 1700
rect 5032 1688 5063 1700
rect 5069 1688 5104 1700
rect 4738 1686 4900 1688
rect 4633 1658 4674 1666
rect 4756 1662 4769 1686
rect 4784 1684 4799 1686
rect 4596 1648 4597 1658
rect 4612 1648 4625 1658
rect 4639 1648 4640 1658
rect 4655 1648 4668 1658
rect 4683 1648 4713 1662
rect 4756 1648 4799 1662
rect 4823 1659 4830 1666
rect 4833 1662 4900 1686
rect 4932 1686 5104 1688
rect 4902 1664 4930 1668
rect 4932 1664 5012 1686
rect 5033 1684 5048 1686
rect 4902 1662 5012 1664
rect 4833 1658 5012 1662
rect 4806 1648 4836 1658
rect 4838 1648 4991 1658
rect 4999 1648 5029 1658
rect 5033 1648 5063 1662
rect 5091 1648 5104 1686
rect 5176 1692 5211 1700
rect 5176 1666 5177 1692
rect 5184 1666 5211 1692
rect 5119 1648 5149 1662
rect 5176 1658 5211 1666
rect 5213 1692 5254 1700
rect 5213 1666 5228 1692
rect 5235 1666 5254 1692
rect 5318 1688 5380 1700
rect 5392 1688 5467 1700
rect 5525 1688 5600 1700
rect 5612 1688 5643 1700
rect 5649 1688 5684 1700
rect 5318 1686 5480 1688
rect 5213 1658 5254 1666
rect 5336 1662 5349 1686
rect 5364 1684 5379 1686
rect 5176 1648 5177 1658
rect 5192 1648 5205 1658
rect 5219 1648 5220 1658
rect 5235 1648 5248 1658
rect 5263 1648 5293 1662
rect 5336 1648 5379 1662
rect 5403 1659 5410 1666
rect 5413 1662 5480 1686
rect 5512 1686 5684 1688
rect 5482 1664 5510 1668
rect 5512 1664 5592 1686
rect 5613 1684 5628 1686
rect 5482 1662 5592 1664
rect 5413 1658 5592 1662
rect 5386 1648 5416 1658
rect 5418 1648 5571 1658
rect 5579 1648 5609 1658
rect 5613 1648 5643 1662
rect 5671 1648 5684 1686
rect 5756 1692 5791 1700
rect 5756 1666 5757 1692
rect 5764 1666 5791 1692
rect 5699 1648 5729 1662
rect 5756 1658 5791 1666
rect 5793 1692 5834 1700
rect 5793 1666 5808 1692
rect 5815 1666 5834 1692
rect 5898 1688 5960 1700
rect 5972 1688 6047 1700
rect 6105 1688 6180 1700
rect 6192 1688 6223 1700
rect 6229 1688 6264 1700
rect 5898 1686 6060 1688
rect 5793 1658 5834 1666
rect 5916 1662 5929 1686
rect 5944 1684 5959 1686
rect 5756 1648 5757 1658
rect 5772 1648 5785 1658
rect 5799 1648 5800 1658
rect 5815 1648 5828 1658
rect 5843 1648 5873 1662
rect 5916 1648 5959 1662
rect 5983 1659 5990 1666
rect 5993 1662 6060 1686
rect 6092 1686 6264 1688
rect 6062 1664 6090 1668
rect 6092 1664 6172 1686
rect 6193 1684 6208 1686
rect 6062 1662 6172 1664
rect 5993 1658 6172 1662
rect 5966 1648 5996 1658
rect 5998 1648 6151 1658
rect 6159 1648 6189 1658
rect 6193 1648 6223 1662
rect 6251 1648 6264 1686
rect 6336 1692 6371 1700
rect 6336 1666 6337 1692
rect 6344 1666 6371 1692
rect 6279 1648 6309 1662
rect 6336 1658 6371 1666
rect 6373 1692 6414 1700
rect 6373 1666 6388 1692
rect 6395 1666 6414 1692
rect 6478 1688 6540 1700
rect 6552 1688 6627 1700
rect 6685 1688 6760 1700
rect 6772 1688 6803 1700
rect 6809 1688 6844 1700
rect 6478 1686 6640 1688
rect 6373 1658 6414 1666
rect 6496 1662 6509 1686
rect 6524 1684 6539 1686
rect 6336 1648 6337 1658
rect 6352 1648 6365 1658
rect 6379 1648 6380 1658
rect 6395 1648 6408 1658
rect 6423 1648 6453 1662
rect 6496 1648 6539 1662
rect 6563 1659 6570 1666
rect 6573 1662 6640 1686
rect 6672 1686 6844 1688
rect 6642 1664 6670 1668
rect 6672 1664 6752 1686
rect 6773 1684 6788 1686
rect 6642 1662 6752 1664
rect 6573 1658 6752 1662
rect 6546 1648 6576 1658
rect 6578 1648 6731 1658
rect 6739 1648 6769 1658
rect 6773 1648 6803 1662
rect 6831 1648 6844 1686
rect 6916 1692 6951 1700
rect 6916 1666 6917 1692
rect 6924 1666 6951 1692
rect 6859 1648 6889 1662
rect 6916 1658 6951 1666
rect 6953 1692 6994 1700
rect 6953 1666 6968 1692
rect 6975 1666 6994 1692
rect 7058 1688 7120 1700
rect 7132 1688 7207 1700
rect 7265 1688 7340 1700
rect 7352 1688 7383 1700
rect 7389 1688 7424 1700
rect 7058 1686 7220 1688
rect 6953 1658 6994 1666
rect 7076 1662 7089 1686
rect 7104 1684 7119 1686
rect 6916 1648 6917 1658
rect 6932 1648 6945 1658
rect 6959 1648 6960 1658
rect 6975 1648 6988 1658
rect 7003 1648 7033 1662
rect 7076 1648 7119 1662
rect 7143 1659 7150 1666
rect 7153 1662 7220 1686
rect 7252 1686 7424 1688
rect 7222 1664 7250 1668
rect 7252 1664 7332 1686
rect 7353 1684 7368 1686
rect 7222 1662 7332 1664
rect 7153 1658 7332 1662
rect 7126 1648 7156 1658
rect 7158 1648 7311 1658
rect 7319 1648 7349 1658
rect 7353 1648 7383 1662
rect 7411 1648 7424 1686
rect 7496 1692 7531 1700
rect 7496 1666 7497 1692
rect 7504 1666 7531 1692
rect 7439 1648 7469 1662
rect 7496 1658 7531 1666
rect 7533 1692 7574 1700
rect 7533 1666 7548 1692
rect 7555 1666 7574 1692
rect 7638 1688 7700 1700
rect 7712 1688 7787 1700
rect 7845 1688 7920 1700
rect 7932 1688 7963 1700
rect 7969 1688 8004 1700
rect 7638 1686 7800 1688
rect 7533 1658 7574 1666
rect 7656 1662 7669 1686
rect 7684 1684 7699 1686
rect 7496 1648 7497 1658
rect 7512 1648 7525 1658
rect 7539 1648 7540 1658
rect 7555 1648 7568 1658
rect 7583 1648 7613 1662
rect 7656 1648 7699 1662
rect 7723 1659 7730 1666
rect 7733 1662 7800 1686
rect 7832 1686 8004 1688
rect 7802 1664 7830 1668
rect 7832 1664 7912 1686
rect 7933 1684 7948 1686
rect 7802 1662 7912 1664
rect 7733 1658 7912 1662
rect 7706 1648 7736 1658
rect 7738 1648 7891 1658
rect 7899 1648 7929 1658
rect 7933 1648 7963 1662
rect 7991 1648 8004 1686
rect 8076 1692 8111 1700
rect 8076 1666 8077 1692
rect 8084 1666 8111 1692
rect 8019 1648 8049 1662
rect 8076 1658 8111 1666
rect 8113 1692 8154 1700
rect 8113 1666 8128 1692
rect 8135 1666 8154 1692
rect 8218 1688 8280 1700
rect 8292 1688 8367 1700
rect 8425 1688 8500 1700
rect 8512 1688 8543 1700
rect 8549 1688 8584 1700
rect 8218 1686 8380 1688
rect 8113 1658 8154 1666
rect 8236 1662 8249 1686
rect 8264 1684 8279 1686
rect 8076 1648 8077 1658
rect 8092 1648 8105 1658
rect 8119 1648 8120 1658
rect 8135 1648 8148 1658
rect 8163 1648 8193 1662
rect 8236 1648 8279 1662
rect 8303 1659 8310 1666
rect 8313 1662 8380 1686
rect 8412 1686 8584 1688
rect 8382 1664 8410 1668
rect 8412 1664 8492 1686
rect 8513 1684 8528 1686
rect 8382 1662 8492 1664
rect 8313 1658 8492 1662
rect 8286 1648 8316 1658
rect 8318 1648 8471 1658
rect 8479 1648 8509 1658
rect 8513 1648 8543 1662
rect 8571 1648 8584 1686
rect 8656 1692 8691 1700
rect 8656 1666 8657 1692
rect 8664 1666 8691 1692
rect 8599 1648 8629 1662
rect 8656 1658 8691 1666
rect 8693 1692 8734 1700
rect 8693 1666 8708 1692
rect 8715 1666 8734 1692
rect 8798 1688 8860 1700
rect 8872 1688 8947 1700
rect 9005 1688 9080 1700
rect 9092 1688 9123 1700
rect 9129 1688 9164 1700
rect 8798 1686 8960 1688
rect 8693 1658 8734 1666
rect 8816 1662 8829 1686
rect 8844 1684 8859 1686
rect 8656 1648 8657 1658
rect 8672 1648 8685 1658
rect 8699 1648 8700 1658
rect 8715 1648 8728 1658
rect 8743 1648 8773 1662
rect 8816 1648 8859 1662
rect 8883 1659 8890 1666
rect 8893 1662 8960 1686
rect 8992 1686 9164 1688
rect 8962 1664 8990 1668
rect 8992 1664 9072 1686
rect 9093 1684 9108 1686
rect 8962 1662 9072 1664
rect 8893 1658 9072 1662
rect 8866 1648 8896 1658
rect 8898 1648 9051 1658
rect 9059 1648 9089 1658
rect 9093 1648 9123 1662
rect 9151 1648 9164 1686
rect 9236 1692 9271 1700
rect 9236 1666 9237 1692
rect 9244 1666 9271 1692
rect 9179 1648 9209 1662
rect 9236 1658 9271 1666
rect 9236 1648 9237 1658
rect 9252 1648 9265 1658
rect -1 1642 9265 1648
rect 0 1634 9265 1642
rect 15 1604 28 1634
rect 43 1616 73 1634
rect 116 1620 130 1634
rect 166 1620 386 1634
rect 117 1618 130 1620
rect 83 1606 98 1618
rect 80 1604 102 1606
rect 107 1604 137 1618
rect 198 1616 351 1620
rect 180 1604 372 1616
rect 415 1604 445 1618
rect 451 1604 464 1634
rect 479 1616 509 1634
rect 552 1604 565 1634
rect 595 1604 608 1634
rect 623 1616 653 1634
rect 696 1620 710 1634
rect 746 1620 966 1634
rect 697 1618 710 1620
rect 663 1606 678 1618
rect 660 1604 682 1606
rect 687 1604 717 1618
rect 778 1616 931 1620
rect 760 1604 952 1616
rect 995 1604 1025 1618
rect 1031 1604 1044 1634
rect 1059 1616 1089 1634
rect 1132 1604 1145 1634
rect 1175 1604 1188 1634
rect 1203 1616 1233 1634
rect 1276 1620 1290 1634
rect 1326 1620 1546 1634
rect 1277 1618 1290 1620
rect 1243 1606 1258 1618
rect 1240 1604 1262 1606
rect 1267 1604 1297 1618
rect 1358 1616 1511 1620
rect 1340 1604 1532 1616
rect 1575 1604 1605 1618
rect 1611 1604 1624 1634
rect 1639 1616 1669 1634
rect 1712 1604 1725 1634
rect 1755 1604 1768 1634
rect 1783 1616 1813 1634
rect 1856 1620 1870 1634
rect 1906 1620 2126 1634
rect 1857 1618 1870 1620
rect 1823 1606 1838 1618
rect 1820 1604 1842 1606
rect 1847 1604 1877 1618
rect 1938 1616 2091 1620
rect 1920 1604 2112 1616
rect 2155 1604 2185 1618
rect 2191 1604 2204 1634
rect 2219 1616 2249 1634
rect 2292 1604 2305 1634
rect 2335 1604 2348 1634
rect 2363 1616 2393 1634
rect 2436 1620 2450 1634
rect 2486 1620 2706 1634
rect 2437 1618 2450 1620
rect 2403 1606 2418 1618
rect 2400 1604 2422 1606
rect 2427 1604 2457 1618
rect 2518 1616 2671 1620
rect 2500 1604 2692 1616
rect 2735 1604 2765 1618
rect 2771 1604 2784 1634
rect 2799 1616 2829 1634
rect 2872 1604 2885 1634
rect 2915 1604 2928 1634
rect 2943 1616 2973 1634
rect 3016 1620 3030 1634
rect 3066 1620 3286 1634
rect 3017 1618 3030 1620
rect 2983 1606 2998 1618
rect 2980 1604 3002 1606
rect 3007 1604 3037 1618
rect 3098 1616 3251 1620
rect 3080 1604 3272 1616
rect 3315 1604 3345 1618
rect 3351 1604 3364 1634
rect 3379 1616 3409 1634
rect 3452 1604 3465 1634
rect 3495 1604 3508 1634
rect 3523 1616 3553 1634
rect 3596 1620 3610 1634
rect 3646 1620 3866 1634
rect 3597 1618 3610 1620
rect 3563 1606 3578 1618
rect 3560 1604 3582 1606
rect 3587 1604 3617 1618
rect 3678 1616 3831 1620
rect 3660 1604 3852 1616
rect 3895 1604 3925 1618
rect 3931 1604 3944 1634
rect 3959 1616 3989 1634
rect 4032 1604 4045 1634
rect 4075 1604 4088 1634
rect 4103 1616 4133 1634
rect 4176 1620 4190 1634
rect 4226 1620 4446 1634
rect 4177 1618 4190 1620
rect 4143 1606 4158 1618
rect 4140 1604 4162 1606
rect 4167 1604 4197 1618
rect 4258 1616 4411 1620
rect 4240 1604 4432 1616
rect 4475 1604 4505 1618
rect 4511 1604 4524 1634
rect 4539 1616 4569 1634
rect 4612 1604 4625 1634
rect 4655 1604 4668 1634
rect 4683 1616 4713 1634
rect 4756 1620 4770 1634
rect 4806 1620 5026 1634
rect 4757 1618 4770 1620
rect 4723 1606 4738 1618
rect 4720 1604 4742 1606
rect 4747 1604 4777 1618
rect 4838 1616 4991 1620
rect 4820 1604 5012 1616
rect 5055 1604 5085 1618
rect 5091 1604 5104 1634
rect 5119 1616 5149 1634
rect 5192 1604 5205 1634
rect 5235 1604 5248 1634
rect 5263 1616 5293 1634
rect 5336 1620 5350 1634
rect 5386 1620 5606 1634
rect 5337 1618 5350 1620
rect 5303 1606 5318 1618
rect 5300 1604 5322 1606
rect 5327 1604 5357 1618
rect 5418 1616 5571 1620
rect 5400 1604 5592 1616
rect 5635 1604 5665 1618
rect 5671 1604 5684 1634
rect 5699 1616 5729 1634
rect 5772 1604 5785 1634
rect 5815 1604 5828 1634
rect 5843 1616 5873 1634
rect 5916 1620 5930 1634
rect 5966 1620 6186 1634
rect 5917 1618 5930 1620
rect 5883 1606 5898 1618
rect 5880 1604 5902 1606
rect 5907 1604 5937 1618
rect 5998 1616 6151 1620
rect 5980 1604 6172 1616
rect 6215 1604 6245 1618
rect 6251 1604 6264 1634
rect 6279 1616 6309 1634
rect 6352 1604 6365 1634
rect 6395 1604 6408 1634
rect 6423 1616 6453 1634
rect 6496 1620 6510 1634
rect 6546 1620 6766 1634
rect 6497 1618 6510 1620
rect 6463 1606 6478 1618
rect 6460 1604 6482 1606
rect 6487 1604 6517 1618
rect 6578 1616 6731 1620
rect 6560 1604 6752 1616
rect 6795 1604 6825 1618
rect 6831 1604 6844 1634
rect 6859 1616 6889 1634
rect 6932 1604 6945 1634
rect 6975 1604 6988 1634
rect 7003 1616 7033 1634
rect 7076 1620 7090 1634
rect 7126 1620 7346 1634
rect 7077 1618 7090 1620
rect 7043 1606 7058 1618
rect 7040 1604 7062 1606
rect 7067 1604 7097 1618
rect 7158 1616 7311 1620
rect 7140 1604 7332 1616
rect 7375 1604 7405 1618
rect 7411 1604 7424 1634
rect 7439 1616 7469 1634
rect 7512 1604 7525 1634
rect 7555 1604 7568 1634
rect 7583 1616 7613 1634
rect 7656 1620 7670 1634
rect 7706 1620 7926 1634
rect 7657 1618 7670 1620
rect 7623 1606 7638 1618
rect 7620 1604 7642 1606
rect 7647 1604 7677 1618
rect 7738 1616 7891 1620
rect 7720 1604 7912 1616
rect 7955 1604 7985 1618
rect 7991 1604 8004 1634
rect 8019 1616 8049 1634
rect 8092 1604 8105 1634
rect 8135 1604 8148 1634
rect 8163 1616 8193 1634
rect 8236 1620 8250 1634
rect 8286 1620 8506 1634
rect 8237 1618 8250 1620
rect 8203 1606 8218 1618
rect 8200 1604 8222 1606
rect 8227 1604 8257 1618
rect 8318 1616 8471 1620
rect 8300 1604 8492 1616
rect 8535 1604 8565 1618
rect 8571 1604 8584 1634
rect 8599 1616 8629 1634
rect 8672 1604 8685 1634
rect 8715 1604 8728 1634
rect 8743 1616 8773 1634
rect 8816 1620 8830 1634
rect 8866 1620 9086 1634
rect 8817 1618 8830 1620
rect 8783 1606 8798 1618
rect 8780 1604 8802 1606
rect 8807 1604 8837 1618
rect 8898 1616 9051 1620
rect 8880 1604 9072 1616
rect 9115 1604 9145 1618
rect 9151 1604 9164 1634
rect 9179 1616 9209 1634
rect 9252 1604 9265 1634
rect 0 1590 9265 1604
rect 15 1486 28 1590
rect 73 1568 74 1578
rect 89 1568 102 1578
rect 73 1564 102 1568
rect 107 1564 137 1590
rect 155 1576 171 1578
rect 243 1576 296 1590
rect 244 1574 308 1576
rect 351 1574 366 1590
rect 415 1587 445 1590
rect 415 1584 451 1587
rect 381 1576 397 1578
rect 155 1564 170 1568
rect 73 1562 170 1564
rect 198 1562 366 1574
rect 382 1564 397 1568
rect 415 1565 454 1584
rect 473 1578 480 1579
rect 479 1571 480 1578
rect 463 1568 464 1571
rect 479 1568 492 1571
rect 415 1564 445 1565
rect 454 1564 460 1565
rect 463 1564 492 1568
rect 382 1563 492 1564
rect 382 1562 498 1563
rect 57 1554 108 1562
rect 57 1542 82 1554
rect 89 1542 108 1554
rect 139 1554 189 1562
rect 139 1546 155 1554
rect 162 1552 189 1554
rect 198 1552 419 1562
rect 162 1542 419 1552
rect 448 1554 498 1562
rect 448 1545 464 1554
rect 57 1534 108 1542
rect 155 1534 419 1542
rect 445 1542 464 1545
rect 471 1542 498 1554
rect 445 1534 498 1542
rect 73 1526 74 1534
rect 89 1526 102 1534
rect 73 1518 89 1526
rect 70 1511 89 1514
rect 70 1502 92 1511
rect 43 1492 92 1502
rect 43 1486 73 1492
rect 92 1487 97 1492
rect 15 1470 89 1486
rect 107 1478 137 1534
rect 172 1524 380 1534
rect 415 1530 460 1534
rect 463 1533 464 1534
rect 479 1533 492 1534
rect 198 1494 387 1524
rect 213 1491 387 1494
rect 206 1488 387 1491
rect 15 1468 28 1470
rect 43 1468 77 1470
rect 15 1452 89 1468
rect 116 1464 129 1478
rect 144 1464 160 1480
rect 206 1475 217 1488
rect -1 1430 0 1446
rect 15 1430 28 1452
rect 43 1430 73 1452
rect 116 1448 178 1464
rect 206 1457 217 1473
rect 222 1468 232 1488
rect 242 1468 256 1488
rect 259 1475 268 1488
rect 284 1475 293 1488
rect 222 1457 256 1468
rect 259 1457 268 1473
rect 284 1457 293 1473
rect 300 1468 310 1488
rect 320 1468 334 1488
rect 335 1475 346 1488
rect 300 1457 334 1468
rect 335 1457 346 1473
rect 392 1464 408 1480
rect 415 1478 445 1530
rect 479 1526 480 1533
rect 464 1518 480 1526
rect 451 1486 464 1505
rect 479 1486 509 1502
rect 451 1470 525 1486
rect 451 1468 464 1470
rect 479 1468 513 1470
rect 116 1446 129 1448
rect 144 1446 178 1448
rect 116 1430 178 1446
rect 222 1441 238 1444
rect 300 1441 330 1452
rect 378 1448 424 1464
rect 451 1452 525 1468
rect 378 1446 412 1448
rect 377 1430 424 1446
rect 451 1430 464 1452
rect 479 1430 509 1452
rect 536 1430 537 1446
rect 552 1430 565 1590
rect 595 1486 608 1590
rect 653 1568 654 1578
rect 669 1568 682 1578
rect 653 1564 682 1568
rect 687 1564 717 1590
rect 735 1576 751 1578
rect 823 1576 876 1590
rect 824 1574 888 1576
rect 931 1574 946 1590
rect 995 1587 1025 1590
rect 995 1584 1031 1587
rect 961 1576 977 1578
rect 735 1564 750 1568
rect 653 1562 750 1564
rect 778 1562 946 1574
rect 962 1564 977 1568
rect 995 1565 1034 1584
rect 1053 1578 1060 1579
rect 1059 1571 1060 1578
rect 1043 1568 1044 1571
rect 1059 1568 1072 1571
rect 995 1564 1025 1565
rect 1034 1564 1040 1565
rect 1043 1564 1072 1568
rect 962 1563 1072 1564
rect 962 1562 1078 1563
rect 637 1554 688 1562
rect 637 1542 662 1554
rect 669 1542 688 1554
rect 719 1554 769 1562
rect 719 1546 735 1554
rect 742 1552 769 1554
rect 778 1552 999 1562
rect 742 1542 999 1552
rect 1028 1554 1078 1562
rect 1028 1545 1044 1554
rect 637 1534 688 1542
rect 735 1534 999 1542
rect 1025 1542 1044 1545
rect 1051 1542 1078 1554
rect 1025 1534 1078 1542
rect 653 1526 654 1534
rect 669 1526 682 1534
rect 653 1518 669 1526
rect 650 1511 669 1514
rect 650 1502 672 1511
rect 623 1492 672 1502
rect 623 1486 653 1492
rect 672 1487 677 1492
rect 595 1470 669 1486
rect 687 1478 717 1534
rect 752 1524 960 1534
rect 995 1530 1040 1534
rect 1043 1533 1044 1534
rect 1059 1533 1072 1534
rect 778 1494 967 1524
rect 793 1491 967 1494
rect 786 1488 967 1491
rect 595 1468 608 1470
rect 623 1468 657 1470
rect 595 1452 669 1468
rect 696 1464 709 1478
rect 724 1464 740 1480
rect 786 1475 797 1488
rect 579 1430 580 1446
rect 595 1430 608 1452
rect 623 1430 653 1452
rect 696 1448 758 1464
rect 786 1457 797 1473
rect 802 1468 812 1488
rect 822 1468 836 1488
rect 839 1475 848 1488
rect 864 1475 873 1488
rect 802 1457 836 1468
rect 839 1457 848 1473
rect 864 1457 873 1473
rect 880 1468 890 1488
rect 900 1468 914 1488
rect 915 1475 926 1488
rect 880 1457 914 1468
rect 915 1457 926 1473
rect 972 1464 988 1480
rect 995 1478 1025 1530
rect 1059 1526 1060 1533
rect 1044 1518 1060 1526
rect 1031 1486 1044 1505
rect 1059 1486 1089 1502
rect 1031 1470 1105 1486
rect 1031 1468 1044 1470
rect 1059 1468 1093 1470
rect 696 1446 709 1448
rect 724 1446 758 1448
rect 696 1430 758 1446
rect 802 1441 818 1444
rect 880 1441 910 1452
rect 958 1448 1004 1464
rect 1031 1452 1105 1468
rect 958 1446 992 1448
rect 957 1430 1004 1446
rect 1031 1430 1044 1452
rect 1059 1430 1089 1452
rect 1116 1430 1117 1446
rect 1132 1430 1145 1590
rect 1175 1486 1188 1590
rect 1233 1568 1234 1578
rect 1249 1568 1262 1578
rect 1233 1564 1262 1568
rect 1267 1564 1297 1590
rect 1315 1576 1331 1578
rect 1403 1576 1456 1590
rect 1404 1574 1468 1576
rect 1511 1574 1526 1590
rect 1575 1587 1605 1590
rect 1575 1584 1611 1587
rect 1541 1576 1557 1578
rect 1315 1564 1330 1568
rect 1233 1562 1330 1564
rect 1358 1562 1526 1574
rect 1542 1564 1557 1568
rect 1575 1565 1614 1584
rect 1633 1578 1640 1579
rect 1639 1571 1640 1578
rect 1623 1568 1624 1571
rect 1639 1568 1652 1571
rect 1575 1564 1605 1565
rect 1614 1564 1620 1565
rect 1623 1564 1652 1568
rect 1542 1563 1652 1564
rect 1542 1562 1658 1563
rect 1217 1554 1268 1562
rect 1217 1542 1242 1554
rect 1249 1542 1268 1554
rect 1299 1554 1349 1562
rect 1299 1546 1315 1554
rect 1322 1552 1349 1554
rect 1358 1552 1579 1562
rect 1322 1542 1579 1552
rect 1608 1554 1658 1562
rect 1608 1545 1624 1554
rect 1217 1534 1268 1542
rect 1315 1534 1579 1542
rect 1605 1542 1624 1545
rect 1631 1542 1658 1554
rect 1605 1534 1658 1542
rect 1233 1526 1234 1534
rect 1249 1526 1262 1534
rect 1233 1518 1249 1526
rect 1230 1511 1249 1514
rect 1230 1502 1252 1511
rect 1203 1492 1252 1502
rect 1203 1486 1233 1492
rect 1252 1487 1257 1492
rect 1175 1470 1249 1486
rect 1267 1478 1297 1534
rect 1332 1524 1540 1534
rect 1575 1530 1620 1534
rect 1623 1533 1624 1534
rect 1639 1533 1652 1534
rect 1358 1494 1547 1524
rect 1373 1491 1547 1494
rect 1366 1488 1547 1491
rect 1175 1468 1188 1470
rect 1203 1468 1237 1470
rect 1175 1452 1249 1468
rect 1276 1464 1289 1478
rect 1304 1464 1320 1480
rect 1366 1475 1377 1488
rect 1159 1430 1160 1446
rect 1175 1430 1188 1452
rect 1203 1430 1233 1452
rect 1276 1448 1338 1464
rect 1366 1457 1377 1473
rect 1382 1468 1392 1488
rect 1402 1468 1416 1488
rect 1419 1475 1428 1488
rect 1444 1475 1453 1488
rect 1382 1457 1416 1468
rect 1419 1457 1428 1473
rect 1444 1457 1453 1473
rect 1460 1468 1470 1488
rect 1480 1468 1494 1488
rect 1495 1475 1506 1488
rect 1460 1457 1494 1468
rect 1495 1457 1506 1473
rect 1552 1464 1568 1480
rect 1575 1478 1605 1530
rect 1639 1526 1640 1533
rect 1624 1518 1640 1526
rect 1611 1486 1624 1505
rect 1639 1486 1669 1502
rect 1611 1470 1685 1486
rect 1611 1468 1624 1470
rect 1639 1468 1673 1470
rect 1276 1446 1289 1448
rect 1304 1446 1338 1448
rect 1276 1430 1338 1446
rect 1382 1441 1398 1444
rect 1460 1441 1490 1452
rect 1538 1448 1584 1464
rect 1611 1452 1685 1468
rect 1538 1446 1572 1448
rect 1537 1430 1584 1446
rect 1611 1430 1624 1452
rect 1639 1430 1669 1452
rect 1696 1430 1697 1446
rect 1712 1430 1725 1590
rect 1755 1486 1768 1590
rect 1813 1568 1814 1578
rect 1829 1568 1842 1578
rect 1813 1564 1842 1568
rect 1847 1564 1877 1590
rect 1895 1576 1911 1578
rect 1983 1576 2036 1590
rect 1984 1574 2048 1576
rect 2091 1574 2106 1590
rect 2155 1587 2185 1590
rect 2155 1584 2191 1587
rect 2121 1576 2137 1578
rect 1895 1564 1910 1568
rect 1813 1562 1910 1564
rect 1938 1562 2106 1574
rect 2122 1564 2137 1568
rect 2155 1565 2194 1584
rect 2213 1578 2220 1579
rect 2219 1571 2220 1578
rect 2203 1568 2204 1571
rect 2219 1568 2232 1571
rect 2155 1564 2185 1565
rect 2194 1564 2200 1565
rect 2203 1564 2232 1568
rect 2122 1563 2232 1564
rect 2122 1562 2238 1563
rect 1797 1554 1848 1562
rect 1797 1542 1822 1554
rect 1829 1542 1848 1554
rect 1879 1554 1929 1562
rect 1879 1546 1895 1554
rect 1902 1552 1929 1554
rect 1938 1552 2159 1562
rect 1902 1542 2159 1552
rect 2188 1554 2238 1562
rect 2188 1545 2204 1554
rect 1797 1534 1848 1542
rect 1895 1534 2159 1542
rect 2185 1542 2204 1545
rect 2211 1542 2238 1554
rect 2185 1534 2238 1542
rect 1813 1526 1814 1534
rect 1829 1526 1842 1534
rect 1813 1518 1829 1526
rect 1810 1511 1829 1514
rect 1810 1502 1832 1511
rect 1783 1492 1832 1502
rect 1783 1486 1813 1492
rect 1832 1487 1837 1492
rect 1755 1470 1829 1486
rect 1847 1478 1877 1534
rect 1912 1524 2120 1534
rect 2155 1530 2200 1534
rect 2203 1533 2204 1534
rect 2219 1533 2232 1534
rect 1938 1494 2127 1524
rect 1953 1491 2127 1494
rect 1946 1488 2127 1491
rect 1755 1468 1768 1470
rect 1783 1468 1817 1470
rect 1755 1452 1829 1468
rect 1856 1464 1869 1478
rect 1884 1464 1900 1480
rect 1946 1475 1957 1488
rect 1739 1430 1740 1446
rect 1755 1430 1768 1452
rect 1783 1430 1813 1452
rect 1856 1448 1918 1464
rect 1946 1457 1957 1473
rect 1962 1468 1972 1488
rect 1982 1468 1996 1488
rect 1999 1475 2008 1488
rect 2024 1475 2033 1488
rect 1962 1457 1996 1468
rect 1999 1457 2008 1473
rect 2024 1457 2033 1473
rect 2040 1468 2050 1488
rect 2060 1468 2074 1488
rect 2075 1475 2086 1488
rect 2040 1457 2074 1468
rect 2075 1457 2086 1473
rect 2132 1464 2148 1480
rect 2155 1478 2185 1530
rect 2219 1526 2220 1533
rect 2204 1518 2220 1526
rect 2191 1486 2204 1505
rect 2219 1486 2249 1502
rect 2191 1470 2265 1486
rect 2191 1468 2204 1470
rect 2219 1468 2253 1470
rect 1856 1446 1869 1448
rect 1884 1446 1918 1448
rect 1856 1430 1918 1446
rect 1962 1441 1976 1444
rect 2040 1441 2070 1452
rect 2118 1448 2164 1464
rect 2191 1452 2265 1468
rect 2118 1446 2152 1448
rect 2117 1430 2164 1446
rect 2191 1430 2204 1452
rect 2219 1430 2249 1452
rect 2276 1430 2277 1446
rect 2292 1430 2305 1590
rect 2335 1486 2348 1590
rect 2393 1568 2394 1578
rect 2409 1568 2422 1578
rect 2393 1564 2422 1568
rect 2427 1564 2457 1590
rect 2475 1576 2491 1578
rect 2563 1576 2616 1590
rect 2564 1574 2628 1576
rect 2671 1574 2686 1590
rect 2735 1587 2765 1590
rect 2735 1584 2771 1587
rect 2701 1576 2717 1578
rect 2475 1564 2490 1568
rect 2393 1562 2490 1564
rect 2518 1562 2686 1574
rect 2702 1564 2717 1568
rect 2735 1565 2774 1584
rect 2793 1578 2800 1579
rect 2799 1571 2800 1578
rect 2783 1568 2784 1571
rect 2799 1568 2812 1571
rect 2735 1564 2765 1565
rect 2774 1564 2780 1565
rect 2783 1564 2812 1568
rect 2702 1563 2812 1564
rect 2702 1562 2818 1563
rect 2377 1554 2428 1562
rect 2377 1542 2402 1554
rect 2409 1542 2428 1554
rect 2459 1554 2509 1562
rect 2459 1546 2475 1554
rect 2482 1552 2509 1554
rect 2518 1552 2739 1562
rect 2482 1542 2739 1552
rect 2768 1554 2818 1562
rect 2768 1545 2784 1554
rect 2377 1534 2428 1542
rect 2475 1534 2739 1542
rect 2765 1542 2784 1545
rect 2791 1542 2818 1554
rect 2765 1534 2818 1542
rect 2393 1526 2394 1534
rect 2409 1526 2422 1534
rect 2393 1518 2409 1526
rect 2390 1511 2409 1514
rect 2390 1502 2412 1511
rect 2363 1492 2412 1502
rect 2363 1486 2393 1492
rect 2412 1487 2417 1492
rect 2335 1470 2409 1486
rect 2427 1478 2457 1534
rect 2492 1524 2700 1534
rect 2735 1530 2780 1534
rect 2783 1533 2784 1534
rect 2799 1533 2812 1534
rect 2518 1494 2707 1524
rect 2533 1491 2707 1494
rect 2526 1488 2707 1491
rect 2335 1468 2348 1470
rect 2363 1468 2397 1470
rect 2335 1452 2409 1468
rect 2436 1464 2449 1478
rect 2464 1464 2480 1480
rect 2526 1475 2537 1488
rect 2319 1430 2320 1446
rect 2335 1430 2348 1452
rect 2363 1430 2393 1452
rect 2436 1448 2498 1464
rect 2526 1457 2537 1473
rect 2542 1468 2552 1488
rect 2562 1468 2576 1488
rect 2579 1475 2588 1488
rect 2604 1475 2613 1488
rect 2542 1457 2576 1468
rect 2579 1457 2588 1473
rect 2604 1457 2613 1473
rect 2620 1468 2630 1488
rect 2640 1468 2654 1488
rect 2655 1475 2666 1488
rect 2620 1457 2654 1468
rect 2655 1457 2666 1473
rect 2712 1464 2728 1480
rect 2735 1478 2765 1530
rect 2799 1526 2800 1533
rect 2784 1518 2800 1526
rect 2771 1486 2784 1505
rect 2799 1486 2829 1502
rect 2771 1470 2845 1486
rect 2771 1468 2784 1470
rect 2799 1468 2833 1470
rect 2436 1446 2449 1448
rect 2464 1446 2498 1448
rect 2436 1430 2498 1446
rect 2542 1441 2558 1444
rect 2620 1441 2650 1452
rect 2698 1448 2744 1464
rect 2771 1452 2845 1468
rect 2698 1446 2732 1448
rect 2697 1430 2744 1446
rect 2771 1430 2784 1452
rect 2799 1430 2829 1452
rect 2856 1430 2857 1446
rect 2872 1430 2885 1590
rect 2915 1486 2928 1590
rect 2973 1568 2974 1578
rect 2989 1568 3002 1578
rect 2973 1564 3002 1568
rect 3007 1564 3037 1590
rect 3055 1576 3071 1578
rect 3143 1576 3196 1590
rect 3144 1574 3208 1576
rect 3251 1574 3266 1590
rect 3315 1587 3345 1590
rect 3315 1584 3351 1587
rect 3281 1576 3297 1578
rect 3055 1564 3070 1568
rect 2973 1562 3070 1564
rect 3098 1562 3266 1574
rect 3282 1564 3297 1568
rect 3315 1565 3354 1584
rect 3373 1578 3380 1579
rect 3379 1571 3380 1578
rect 3363 1568 3364 1571
rect 3379 1568 3392 1571
rect 3315 1564 3345 1565
rect 3354 1564 3360 1565
rect 3363 1564 3392 1568
rect 3282 1563 3392 1564
rect 3282 1562 3398 1563
rect 2957 1554 3008 1562
rect 2957 1542 2982 1554
rect 2989 1542 3008 1554
rect 3039 1554 3089 1562
rect 3039 1546 3055 1554
rect 3062 1552 3089 1554
rect 3098 1552 3319 1562
rect 3062 1542 3319 1552
rect 3348 1554 3398 1562
rect 3348 1545 3364 1554
rect 2957 1534 3008 1542
rect 3055 1534 3319 1542
rect 3345 1542 3364 1545
rect 3371 1542 3398 1554
rect 3345 1534 3398 1542
rect 2973 1526 2974 1534
rect 2989 1526 3002 1534
rect 2973 1518 2989 1526
rect 2970 1511 2989 1514
rect 2970 1502 2992 1511
rect 2943 1492 2992 1502
rect 2943 1486 2973 1492
rect 2992 1487 2997 1492
rect 2915 1470 2989 1486
rect 3007 1478 3037 1534
rect 3072 1524 3280 1534
rect 3315 1530 3360 1534
rect 3363 1533 3364 1534
rect 3379 1533 3392 1534
rect 3098 1494 3287 1524
rect 3113 1491 3287 1494
rect 3106 1488 3287 1491
rect 2915 1468 2928 1470
rect 2943 1468 2977 1470
rect 2915 1452 2989 1468
rect 3016 1464 3029 1478
rect 3044 1464 3060 1480
rect 3106 1475 3117 1488
rect 2899 1430 2900 1446
rect 2915 1430 2928 1452
rect 2943 1430 2973 1452
rect 3016 1448 3078 1464
rect 3106 1457 3117 1473
rect 3122 1468 3132 1488
rect 3142 1468 3156 1488
rect 3159 1475 3168 1488
rect 3184 1475 3193 1488
rect 3122 1457 3156 1468
rect 3159 1457 3168 1473
rect 3184 1457 3193 1473
rect 3200 1468 3210 1488
rect 3220 1468 3234 1488
rect 3235 1475 3246 1488
rect 3200 1457 3234 1468
rect 3235 1457 3246 1473
rect 3292 1464 3308 1480
rect 3315 1478 3345 1530
rect 3379 1526 3380 1533
rect 3364 1518 3380 1526
rect 3351 1486 3364 1505
rect 3379 1486 3409 1502
rect 3351 1470 3425 1486
rect 3351 1468 3364 1470
rect 3379 1468 3413 1470
rect 3016 1446 3029 1448
rect 3044 1446 3078 1448
rect 3016 1430 3078 1446
rect 3122 1441 3138 1444
rect 3200 1441 3230 1452
rect 3278 1448 3324 1464
rect 3351 1452 3425 1468
rect 3278 1446 3312 1448
rect 3277 1430 3324 1446
rect 3351 1430 3364 1452
rect 3379 1430 3409 1452
rect 3436 1430 3437 1446
rect 3452 1430 3465 1590
rect 3495 1486 3508 1590
rect 3553 1568 3554 1578
rect 3569 1568 3582 1578
rect 3553 1564 3582 1568
rect 3587 1564 3617 1590
rect 3635 1576 3651 1578
rect 3723 1576 3776 1590
rect 3724 1574 3788 1576
rect 3831 1574 3846 1590
rect 3895 1587 3925 1590
rect 3895 1584 3931 1587
rect 3861 1576 3877 1578
rect 3635 1564 3650 1568
rect 3553 1562 3650 1564
rect 3678 1562 3846 1574
rect 3862 1564 3877 1568
rect 3895 1565 3934 1584
rect 3953 1578 3960 1579
rect 3959 1571 3960 1578
rect 3943 1568 3944 1571
rect 3959 1568 3972 1571
rect 3895 1564 3925 1565
rect 3934 1564 3940 1565
rect 3943 1564 3972 1568
rect 3862 1563 3972 1564
rect 3862 1562 3978 1563
rect 3537 1554 3588 1562
rect 3537 1542 3562 1554
rect 3569 1542 3588 1554
rect 3619 1554 3669 1562
rect 3619 1546 3635 1554
rect 3642 1552 3669 1554
rect 3678 1552 3899 1562
rect 3642 1542 3899 1552
rect 3928 1554 3978 1562
rect 3928 1545 3944 1554
rect 3537 1534 3588 1542
rect 3635 1534 3899 1542
rect 3925 1542 3944 1545
rect 3951 1542 3978 1554
rect 3925 1534 3978 1542
rect 3553 1526 3554 1534
rect 3569 1526 3582 1534
rect 3553 1518 3569 1526
rect 3550 1511 3569 1514
rect 3550 1502 3572 1511
rect 3523 1492 3572 1502
rect 3523 1486 3553 1492
rect 3572 1487 3577 1492
rect 3495 1470 3569 1486
rect 3587 1478 3617 1534
rect 3652 1524 3860 1534
rect 3895 1530 3940 1534
rect 3943 1533 3944 1534
rect 3959 1533 3972 1534
rect 3678 1494 3867 1524
rect 3693 1491 3867 1494
rect 3686 1488 3867 1491
rect 3495 1468 3508 1470
rect 3523 1468 3557 1470
rect 3495 1452 3569 1468
rect 3596 1464 3609 1478
rect 3624 1464 3640 1480
rect 3686 1475 3697 1488
rect 3479 1430 3480 1446
rect 3495 1430 3508 1452
rect 3523 1430 3553 1452
rect 3596 1448 3658 1464
rect 3686 1457 3697 1473
rect 3702 1468 3712 1488
rect 3722 1468 3736 1488
rect 3739 1475 3748 1488
rect 3764 1475 3773 1488
rect 3702 1457 3736 1468
rect 3739 1457 3748 1473
rect 3764 1457 3773 1473
rect 3780 1468 3790 1488
rect 3800 1468 3814 1488
rect 3815 1475 3826 1488
rect 3780 1457 3814 1468
rect 3815 1457 3826 1473
rect 3872 1464 3888 1480
rect 3895 1478 3925 1530
rect 3959 1526 3960 1533
rect 3944 1518 3960 1526
rect 3931 1486 3944 1505
rect 3959 1486 3989 1502
rect 3931 1470 4005 1486
rect 3931 1468 3944 1470
rect 3959 1468 3993 1470
rect 3596 1446 3609 1448
rect 3624 1446 3658 1448
rect 3596 1430 3658 1446
rect 3702 1441 3718 1444
rect 3780 1441 3810 1452
rect 3858 1448 3904 1464
rect 3931 1452 4005 1468
rect 3858 1446 3892 1448
rect 3857 1430 3904 1446
rect 3931 1430 3944 1452
rect 3959 1430 3989 1452
rect 4016 1430 4017 1446
rect 4032 1430 4045 1590
rect 4075 1486 4088 1590
rect 4133 1568 4134 1578
rect 4149 1568 4162 1578
rect 4133 1564 4162 1568
rect 4167 1564 4197 1590
rect 4215 1576 4231 1578
rect 4303 1576 4356 1590
rect 4304 1574 4368 1576
rect 4411 1574 4426 1590
rect 4475 1587 4505 1590
rect 4475 1584 4511 1587
rect 4441 1576 4457 1578
rect 4215 1564 4230 1568
rect 4133 1562 4230 1564
rect 4258 1562 4426 1574
rect 4442 1564 4457 1568
rect 4475 1565 4514 1584
rect 4533 1578 4540 1579
rect 4539 1571 4540 1578
rect 4523 1568 4524 1571
rect 4539 1568 4552 1571
rect 4475 1564 4505 1565
rect 4514 1564 4520 1565
rect 4523 1564 4552 1568
rect 4442 1563 4552 1564
rect 4442 1562 4558 1563
rect 4117 1554 4168 1562
rect 4117 1542 4142 1554
rect 4149 1542 4168 1554
rect 4199 1554 4249 1562
rect 4199 1546 4215 1554
rect 4222 1552 4249 1554
rect 4258 1552 4479 1562
rect 4222 1542 4479 1552
rect 4508 1554 4558 1562
rect 4508 1545 4524 1554
rect 4117 1534 4168 1542
rect 4215 1534 4479 1542
rect 4505 1542 4524 1545
rect 4531 1542 4558 1554
rect 4505 1534 4558 1542
rect 4133 1526 4134 1534
rect 4149 1526 4162 1534
rect 4133 1518 4149 1526
rect 4130 1511 4149 1514
rect 4130 1502 4152 1511
rect 4103 1492 4152 1502
rect 4103 1486 4133 1492
rect 4152 1487 4157 1492
rect 4075 1470 4149 1486
rect 4167 1478 4197 1534
rect 4232 1524 4440 1534
rect 4475 1530 4520 1534
rect 4523 1533 4524 1534
rect 4539 1533 4552 1534
rect 4258 1494 4447 1524
rect 4273 1491 4447 1494
rect 4266 1488 4447 1491
rect 4075 1468 4088 1470
rect 4103 1468 4137 1470
rect 4075 1452 4149 1468
rect 4176 1464 4189 1478
rect 4204 1464 4220 1480
rect 4266 1475 4277 1488
rect 4059 1430 4060 1446
rect 4075 1430 4088 1452
rect 4103 1430 4133 1452
rect 4176 1448 4238 1464
rect 4266 1457 4277 1473
rect 4282 1468 4292 1488
rect 4302 1468 4316 1488
rect 4319 1475 4328 1488
rect 4344 1475 4353 1488
rect 4282 1457 4316 1468
rect 4319 1457 4328 1473
rect 4344 1457 4353 1473
rect 4360 1468 4370 1488
rect 4380 1468 4394 1488
rect 4395 1475 4406 1488
rect 4360 1457 4394 1468
rect 4395 1457 4406 1473
rect 4452 1464 4468 1480
rect 4475 1478 4505 1530
rect 4539 1526 4540 1533
rect 4524 1518 4540 1526
rect 4511 1486 4524 1505
rect 4539 1486 4569 1502
rect 4511 1470 4585 1486
rect 4511 1468 4524 1470
rect 4539 1468 4573 1470
rect 4176 1446 4189 1448
rect 4204 1446 4238 1448
rect 4176 1430 4238 1446
rect 4282 1441 4298 1444
rect 4360 1441 4390 1452
rect 4438 1448 4484 1464
rect 4511 1452 4585 1468
rect 4438 1446 4472 1448
rect 4437 1430 4484 1446
rect 4511 1430 4524 1452
rect 4539 1430 4569 1452
rect 4596 1430 4597 1446
rect 4612 1430 4625 1590
rect 4655 1486 4668 1590
rect 4713 1568 4714 1578
rect 4729 1568 4742 1578
rect 4713 1564 4742 1568
rect 4747 1564 4777 1590
rect 4795 1576 4811 1578
rect 4883 1576 4936 1590
rect 4884 1574 4948 1576
rect 4991 1574 5006 1590
rect 5055 1587 5085 1590
rect 5055 1584 5091 1587
rect 5021 1576 5037 1578
rect 4795 1564 4810 1568
rect 4713 1562 4810 1564
rect 4838 1562 5006 1574
rect 5022 1564 5037 1568
rect 5055 1565 5094 1584
rect 5113 1578 5120 1579
rect 5119 1571 5120 1578
rect 5103 1568 5104 1571
rect 5119 1568 5132 1571
rect 5055 1564 5085 1565
rect 5094 1564 5100 1565
rect 5103 1564 5132 1568
rect 5022 1563 5132 1564
rect 5022 1562 5138 1563
rect 4697 1554 4748 1562
rect 4697 1542 4722 1554
rect 4729 1542 4748 1554
rect 4779 1554 4829 1562
rect 4779 1546 4795 1554
rect 4802 1552 4829 1554
rect 4838 1552 5059 1562
rect 4802 1542 5059 1552
rect 5088 1554 5138 1562
rect 5088 1545 5104 1554
rect 4697 1534 4748 1542
rect 4795 1534 5059 1542
rect 5085 1542 5104 1545
rect 5111 1542 5138 1554
rect 5085 1534 5138 1542
rect 4713 1526 4714 1534
rect 4729 1526 4742 1534
rect 4713 1518 4729 1526
rect 4710 1511 4729 1514
rect 4710 1502 4732 1511
rect 4683 1492 4732 1502
rect 4683 1486 4713 1492
rect 4732 1487 4737 1492
rect 4655 1470 4729 1486
rect 4747 1478 4777 1534
rect 4812 1524 5020 1534
rect 5055 1530 5100 1534
rect 5103 1533 5104 1534
rect 5119 1533 5132 1534
rect 4838 1494 5027 1524
rect 4853 1491 5027 1494
rect 4846 1488 5027 1491
rect 4655 1468 4668 1470
rect 4683 1468 4717 1470
rect 4655 1452 4729 1468
rect 4756 1464 4769 1478
rect 4784 1464 4800 1480
rect 4846 1475 4857 1488
rect 4639 1430 4640 1446
rect 4655 1430 4668 1452
rect 4683 1430 4713 1452
rect 4756 1448 4818 1464
rect 4846 1457 4857 1473
rect 4862 1468 4872 1488
rect 4882 1468 4896 1488
rect 4899 1475 4908 1488
rect 4924 1475 4933 1488
rect 4862 1457 4896 1468
rect 4899 1457 4908 1473
rect 4924 1457 4933 1473
rect 4940 1468 4950 1488
rect 4960 1468 4974 1488
rect 4975 1475 4986 1488
rect 4940 1457 4974 1468
rect 4975 1457 4986 1473
rect 5032 1464 5048 1480
rect 5055 1478 5085 1530
rect 5119 1526 5120 1533
rect 5104 1518 5120 1526
rect 5091 1486 5104 1505
rect 5119 1486 5149 1502
rect 5091 1470 5165 1486
rect 5091 1468 5104 1470
rect 5119 1468 5153 1470
rect 4756 1446 4769 1448
rect 4784 1446 4818 1448
rect 4756 1430 4818 1446
rect 4862 1441 4878 1444
rect 4940 1441 4970 1452
rect 5018 1448 5064 1464
rect 5091 1452 5165 1468
rect 5018 1446 5052 1448
rect 5017 1430 5064 1446
rect 5091 1430 5104 1452
rect 5119 1430 5149 1452
rect 5176 1430 5177 1446
rect 5192 1430 5205 1590
rect 5235 1486 5248 1590
rect 5293 1568 5294 1578
rect 5309 1568 5322 1578
rect 5293 1564 5322 1568
rect 5327 1564 5357 1590
rect 5375 1576 5391 1578
rect 5463 1576 5516 1590
rect 5464 1574 5528 1576
rect 5571 1574 5586 1590
rect 5635 1587 5665 1590
rect 5635 1584 5671 1587
rect 5601 1576 5617 1578
rect 5375 1564 5390 1568
rect 5293 1562 5390 1564
rect 5418 1562 5586 1574
rect 5602 1564 5617 1568
rect 5635 1565 5674 1584
rect 5693 1578 5700 1579
rect 5699 1571 5700 1578
rect 5683 1568 5684 1571
rect 5699 1568 5712 1571
rect 5635 1564 5665 1565
rect 5674 1564 5680 1565
rect 5683 1564 5712 1568
rect 5602 1563 5712 1564
rect 5602 1562 5718 1563
rect 5277 1554 5328 1562
rect 5277 1542 5302 1554
rect 5309 1542 5328 1554
rect 5359 1554 5409 1562
rect 5359 1546 5375 1554
rect 5382 1552 5409 1554
rect 5418 1552 5639 1562
rect 5382 1542 5639 1552
rect 5668 1554 5718 1562
rect 5668 1545 5684 1554
rect 5277 1534 5328 1542
rect 5375 1534 5639 1542
rect 5665 1542 5684 1545
rect 5691 1542 5718 1554
rect 5665 1534 5718 1542
rect 5293 1526 5294 1534
rect 5309 1526 5322 1534
rect 5293 1518 5309 1526
rect 5290 1511 5309 1514
rect 5290 1502 5312 1511
rect 5263 1492 5312 1502
rect 5263 1486 5293 1492
rect 5312 1487 5317 1492
rect 5235 1470 5309 1486
rect 5327 1478 5357 1534
rect 5392 1524 5600 1534
rect 5635 1530 5680 1534
rect 5683 1533 5684 1534
rect 5699 1533 5712 1534
rect 5418 1494 5607 1524
rect 5433 1491 5607 1494
rect 5426 1488 5607 1491
rect 5235 1468 5248 1470
rect 5263 1468 5297 1470
rect 5235 1452 5309 1468
rect 5336 1464 5349 1478
rect 5364 1464 5380 1480
rect 5426 1475 5437 1488
rect 5219 1430 5220 1446
rect 5235 1430 5248 1452
rect 5263 1430 5293 1452
rect 5336 1448 5398 1464
rect 5426 1457 5437 1473
rect 5442 1468 5452 1488
rect 5462 1468 5476 1488
rect 5479 1475 5488 1488
rect 5504 1475 5513 1488
rect 5442 1457 5476 1468
rect 5479 1457 5488 1473
rect 5504 1457 5513 1473
rect 5520 1468 5530 1488
rect 5540 1468 5554 1488
rect 5555 1475 5566 1488
rect 5520 1457 5554 1468
rect 5555 1457 5566 1473
rect 5612 1464 5628 1480
rect 5635 1478 5665 1530
rect 5699 1526 5700 1533
rect 5684 1518 5700 1526
rect 5671 1486 5684 1505
rect 5699 1486 5729 1502
rect 5671 1470 5745 1486
rect 5671 1468 5684 1470
rect 5699 1468 5733 1470
rect 5336 1446 5349 1448
rect 5364 1446 5398 1448
rect 5336 1430 5398 1446
rect 5442 1441 5458 1444
rect 5520 1441 5550 1452
rect 5598 1448 5644 1464
rect 5671 1452 5745 1468
rect 5598 1446 5632 1448
rect 5597 1430 5644 1446
rect 5671 1430 5684 1452
rect 5699 1430 5729 1452
rect 5756 1430 5757 1446
rect 5772 1430 5785 1590
rect 5815 1486 5828 1590
rect 5873 1568 5874 1578
rect 5889 1568 5902 1578
rect 5873 1564 5902 1568
rect 5907 1564 5937 1590
rect 5955 1576 5971 1578
rect 6043 1576 6096 1590
rect 6044 1574 6108 1576
rect 6151 1574 6166 1590
rect 6215 1587 6245 1590
rect 6215 1584 6251 1587
rect 6181 1576 6197 1578
rect 5955 1564 5970 1568
rect 5873 1562 5970 1564
rect 5998 1562 6166 1574
rect 6182 1564 6197 1568
rect 6215 1565 6254 1584
rect 6273 1578 6280 1579
rect 6279 1571 6280 1578
rect 6263 1568 6264 1571
rect 6279 1568 6292 1571
rect 6215 1564 6245 1565
rect 6254 1564 6260 1565
rect 6263 1564 6292 1568
rect 6182 1563 6292 1564
rect 6182 1562 6298 1563
rect 5857 1554 5908 1562
rect 5857 1542 5882 1554
rect 5889 1542 5908 1554
rect 5939 1554 5989 1562
rect 5939 1546 5955 1554
rect 5962 1552 5989 1554
rect 5998 1552 6219 1562
rect 5962 1542 6219 1552
rect 6248 1554 6298 1562
rect 6248 1545 6264 1554
rect 5857 1534 5908 1542
rect 5955 1534 6219 1542
rect 6245 1542 6264 1545
rect 6271 1542 6298 1554
rect 6245 1534 6298 1542
rect 5873 1526 5874 1534
rect 5889 1526 5902 1534
rect 5873 1518 5889 1526
rect 5870 1511 5889 1514
rect 5870 1502 5892 1511
rect 5843 1492 5892 1502
rect 5843 1486 5873 1492
rect 5892 1487 5897 1492
rect 5815 1470 5889 1486
rect 5907 1478 5937 1534
rect 5972 1524 6180 1534
rect 6215 1530 6260 1534
rect 6263 1533 6264 1534
rect 6279 1533 6292 1534
rect 5998 1494 6187 1524
rect 6013 1491 6187 1494
rect 6006 1488 6187 1491
rect 5815 1468 5828 1470
rect 5843 1468 5877 1470
rect 5815 1452 5889 1468
rect 5916 1464 5929 1478
rect 5944 1464 5960 1480
rect 6006 1475 6017 1488
rect 5799 1430 5800 1446
rect 5815 1430 5828 1452
rect 5843 1430 5873 1452
rect 5916 1448 5978 1464
rect 6006 1457 6017 1473
rect 6022 1468 6032 1488
rect 6042 1468 6056 1488
rect 6059 1475 6068 1488
rect 6084 1475 6093 1488
rect 6022 1457 6056 1468
rect 6059 1457 6068 1473
rect 6084 1457 6093 1473
rect 6100 1468 6110 1488
rect 6120 1468 6134 1488
rect 6135 1475 6146 1488
rect 6100 1457 6134 1468
rect 6135 1457 6146 1473
rect 6192 1464 6208 1480
rect 6215 1478 6245 1530
rect 6279 1526 6280 1533
rect 6264 1518 6280 1526
rect 6251 1486 6264 1505
rect 6279 1486 6309 1502
rect 6251 1470 6325 1486
rect 6251 1468 6264 1470
rect 6279 1468 6313 1470
rect 5916 1446 5929 1448
rect 5944 1446 5978 1448
rect 5916 1430 5978 1446
rect 6022 1441 6038 1444
rect 6100 1441 6130 1452
rect 6178 1448 6224 1464
rect 6251 1452 6325 1468
rect 6178 1446 6212 1448
rect 6177 1430 6224 1446
rect 6251 1430 6264 1452
rect 6279 1430 6309 1452
rect 6336 1430 6337 1446
rect 6352 1430 6365 1590
rect 6395 1486 6408 1590
rect 6453 1568 6454 1578
rect 6469 1568 6482 1578
rect 6453 1564 6482 1568
rect 6487 1564 6517 1590
rect 6535 1576 6551 1578
rect 6623 1576 6676 1590
rect 6624 1574 6688 1576
rect 6731 1574 6746 1590
rect 6795 1587 6825 1590
rect 6795 1584 6831 1587
rect 6761 1576 6777 1578
rect 6535 1564 6550 1568
rect 6453 1562 6550 1564
rect 6578 1562 6746 1574
rect 6762 1564 6777 1568
rect 6795 1565 6834 1584
rect 6853 1578 6860 1579
rect 6859 1571 6860 1578
rect 6843 1568 6844 1571
rect 6859 1568 6872 1571
rect 6795 1564 6825 1565
rect 6834 1564 6840 1565
rect 6843 1564 6872 1568
rect 6762 1563 6872 1564
rect 6762 1562 6878 1563
rect 6437 1554 6488 1562
rect 6437 1542 6462 1554
rect 6469 1542 6488 1554
rect 6519 1554 6569 1562
rect 6519 1546 6535 1554
rect 6542 1552 6569 1554
rect 6578 1552 6799 1562
rect 6542 1542 6799 1552
rect 6828 1554 6878 1562
rect 6828 1545 6844 1554
rect 6437 1534 6488 1542
rect 6535 1534 6799 1542
rect 6825 1542 6844 1545
rect 6851 1542 6878 1554
rect 6825 1534 6878 1542
rect 6453 1526 6454 1534
rect 6469 1526 6482 1534
rect 6453 1518 6469 1526
rect 6450 1511 6469 1514
rect 6450 1502 6472 1511
rect 6423 1492 6472 1502
rect 6423 1486 6453 1492
rect 6472 1487 6477 1492
rect 6395 1470 6469 1486
rect 6487 1478 6517 1534
rect 6552 1524 6760 1534
rect 6795 1530 6840 1534
rect 6843 1533 6844 1534
rect 6859 1533 6872 1534
rect 6578 1494 6767 1524
rect 6593 1491 6767 1494
rect 6586 1488 6767 1491
rect 6395 1468 6408 1470
rect 6423 1468 6457 1470
rect 6395 1452 6469 1468
rect 6496 1464 6509 1478
rect 6524 1464 6540 1480
rect 6586 1475 6597 1488
rect 6379 1430 6380 1446
rect 6395 1430 6408 1452
rect 6423 1430 6453 1452
rect 6496 1448 6558 1464
rect 6586 1457 6597 1473
rect 6602 1468 6612 1488
rect 6622 1468 6636 1488
rect 6639 1475 6648 1488
rect 6664 1475 6673 1488
rect 6602 1457 6636 1468
rect 6639 1457 6648 1473
rect 6664 1457 6673 1473
rect 6680 1468 6690 1488
rect 6700 1468 6714 1488
rect 6715 1475 6726 1488
rect 6680 1457 6714 1468
rect 6715 1457 6726 1473
rect 6772 1464 6788 1480
rect 6795 1478 6825 1530
rect 6859 1526 6860 1533
rect 6844 1518 6860 1526
rect 6831 1486 6844 1505
rect 6859 1486 6889 1502
rect 6831 1470 6905 1486
rect 6831 1468 6844 1470
rect 6859 1468 6893 1470
rect 6496 1446 6509 1448
rect 6524 1446 6558 1448
rect 6496 1430 6558 1446
rect 6602 1441 6618 1444
rect 6680 1441 6710 1452
rect 6758 1448 6804 1464
rect 6831 1452 6905 1468
rect 6758 1446 6792 1448
rect 6757 1430 6804 1446
rect 6831 1430 6844 1452
rect 6859 1430 6889 1452
rect 6916 1430 6917 1446
rect 6932 1430 6945 1590
rect 6975 1486 6988 1590
rect 7033 1568 7034 1578
rect 7049 1568 7062 1578
rect 7033 1564 7062 1568
rect 7067 1564 7097 1590
rect 7115 1576 7131 1578
rect 7203 1576 7256 1590
rect 7204 1574 7268 1576
rect 7311 1574 7326 1590
rect 7375 1587 7405 1590
rect 7375 1584 7411 1587
rect 7341 1576 7357 1578
rect 7115 1564 7130 1568
rect 7033 1562 7130 1564
rect 7158 1562 7326 1574
rect 7342 1564 7357 1568
rect 7375 1565 7414 1584
rect 7433 1578 7440 1579
rect 7439 1571 7440 1578
rect 7423 1568 7424 1571
rect 7439 1568 7452 1571
rect 7375 1564 7405 1565
rect 7414 1564 7420 1565
rect 7423 1564 7452 1568
rect 7342 1563 7452 1564
rect 7342 1562 7458 1563
rect 7017 1554 7068 1562
rect 7017 1542 7042 1554
rect 7049 1542 7068 1554
rect 7099 1554 7149 1562
rect 7099 1546 7115 1554
rect 7122 1552 7149 1554
rect 7158 1552 7379 1562
rect 7122 1542 7379 1552
rect 7408 1554 7458 1562
rect 7408 1545 7424 1554
rect 7017 1534 7068 1542
rect 7115 1534 7379 1542
rect 7405 1542 7424 1545
rect 7431 1542 7458 1554
rect 7405 1534 7458 1542
rect 7033 1526 7034 1534
rect 7049 1526 7062 1534
rect 7033 1518 7049 1526
rect 7030 1511 7049 1514
rect 7030 1502 7052 1511
rect 7003 1492 7052 1502
rect 7003 1486 7033 1492
rect 7052 1487 7057 1492
rect 6975 1470 7049 1486
rect 7067 1478 7097 1534
rect 7132 1524 7340 1534
rect 7375 1530 7420 1534
rect 7423 1533 7424 1534
rect 7439 1533 7452 1534
rect 7158 1494 7347 1524
rect 7173 1491 7347 1494
rect 7166 1488 7347 1491
rect 6975 1468 6988 1470
rect 7003 1468 7037 1470
rect 6975 1452 7049 1468
rect 7076 1464 7089 1478
rect 7104 1464 7120 1480
rect 7166 1475 7177 1488
rect 6959 1430 6960 1446
rect 6975 1430 6988 1452
rect 7003 1430 7033 1452
rect 7076 1448 7138 1464
rect 7166 1457 7177 1473
rect 7182 1468 7192 1488
rect 7202 1468 7216 1488
rect 7219 1475 7228 1488
rect 7244 1475 7253 1488
rect 7182 1457 7216 1468
rect 7219 1457 7228 1473
rect 7244 1457 7253 1473
rect 7260 1468 7270 1488
rect 7280 1468 7294 1488
rect 7295 1475 7306 1488
rect 7260 1457 7294 1468
rect 7295 1457 7306 1473
rect 7352 1464 7368 1480
rect 7375 1478 7405 1530
rect 7439 1526 7440 1533
rect 7424 1518 7440 1526
rect 7411 1486 7424 1505
rect 7439 1486 7469 1502
rect 7411 1470 7485 1486
rect 7411 1468 7424 1470
rect 7439 1468 7473 1470
rect 7076 1446 7089 1448
rect 7104 1446 7138 1448
rect 7076 1430 7138 1446
rect 7182 1441 7198 1444
rect 7260 1441 7290 1452
rect 7338 1448 7384 1464
rect 7411 1452 7485 1468
rect 7338 1446 7372 1448
rect 7337 1430 7384 1446
rect 7411 1430 7424 1452
rect 7439 1430 7469 1452
rect 7496 1430 7497 1446
rect 7512 1430 7525 1590
rect 7555 1486 7568 1590
rect 7613 1568 7614 1578
rect 7629 1568 7642 1578
rect 7613 1564 7642 1568
rect 7647 1564 7677 1590
rect 7695 1576 7711 1578
rect 7783 1576 7836 1590
rect 7784 1574 7848 1576
rect 7891 1574 7906 1590
rect 7955 1587 7985 1590
rect 7955 1584 7991 1587
rect 7921 1576 7937 1578
rect 7695 1564 7710 1568
rect 7613 1562 7710 1564
rect 7738 1562 7906 1574
rect 7922 1564 7937 1568
rect 7955 1565 7994 1584
rect 8013 1578 8020 1579
rect 8019 1571 8020 1578
rect 8003 1568 8004 1571
rect 8019 1568 8032 1571
rect 7955 1564 7985 1565
rect 7994 1564 8000 1565
rect 8003 1564 8032 1568
rect 7922 1563 8032 1564
rect 7922 1562 8038 1563
rect 7597 1554 7648 1562
rect 7597 1542 7622 1554
rect 7629 1542 7648 1554
rect 7679 1554 7729 1562
rect 7679 1546 7695 1554
rect 7702 1552 7729 1554
rect 7738 1552 7959 1562
rect 7702 1542 7959 1552
rect 7988 1554 8038 1562
rect 7988 1545 8004 1554
rect 7597 1534 7648 1542
rect 7695 1534 7959 1542
rect 7985 1542 8004 1545
rect 8011 1542 8038 1554
rect 7985 1534 8038 1542
rect 7613 1526 7614 1534
rect 7629 1526 7642 1534
rect 7613 1518 7629 1526
rect 7610 1511 7629 1514
rect 7610 1502 7632 1511
rect 7583 1492 7632 1502
rect 7583 1486 7613 1492
rect 7632 1487 7637 1492
rect 7555 1470 7629 1486
rect 7647 1478 7677 1534
rect 7712 1524 7920 1534
rect 7955 1530 8000 1534
rect 8003 1533 8004 1534
rect 8019 1533 8032 1534
rect 7738 1494 7927 1524
rect 7753 1491 7927 1494
rect 7746 1488 7927 1491
rect 7555 1468 7568 1470
rect 7583 1468 7617 1470
rect 7555 1452 7629 1468
rect 7656 1464 7669 1478
rect 7684 1464 7700 1480
rect 7746 1475 7757 1488
rect 7539 1430 7540 1446
rect 7555 1430 7568 1452
rect 7583 1430 7613 1452
rect 7656 1448 7718 1464
rect 7746 1457 7757 1473
rect 7762 1468 7772 1488
rect 7782 1468 7796 1488
rect 7799 1475 7808 1488
rect 7824 1475 7833 1488
rect 7762 1457 7796 1468
rect 7799 1457 7808 1473
rect 7824 1457 7833 1473
rect 7840 1468 7850 1488
rect 7860 1468 7874 1488
rect 7875 1475 7886 1488
rect 7840 1457 7874 1468
rect 7875 1457 7886 1473
rect 7932 1464 7948 1480
rect 7955 1478 7985 1530
rect 8019 1526 8020 1533
rect 8004 1518 8020 1526
rect 7991 1486 8004 1505
rect 8019 1486 8049 1502
rect 7991 1470 8065 1486
rect 7991 1468 8004 1470
rect 8019 1468 8053 1470
rect 7656 1446 7669 1448
rect 7684 1446 7718 1448
rect 7656 1430 7718 1446
rect 7762 1441 7778 1444
rect 7840 1441 7870 1452
rect 7918 1448 7964 1464
rect 7991 1452 8065 1468
rect 7918 1446 7952 1448
rect 7917 1430 7964 1446
rect 7991 1430 8004 1452
rect 8019 1430 8049 1452
rect 8076 1430 8077 1446
rect 8092 1430 8105 1590
rect 8135 1486 8148 1590
rect 8193 1568 8194 1578
rect 8209 1568 8222 1578
rect 8193 1564 8222 1568
rect 8227 1564 8257 1590
rect 8275 1576 8291 1578
rect 8363 1576 8416 1590
rect 8364 1574 8428 1576
rect 8471 1574 8486 1590
rect 8535 1587 8565 1590
rect 8535 1584 8571 1587
rect 8501 1576 8517 1578
rect 8275 1564 8290 1568
rect 8193 1562 8290 1564
rect 8318 1562 8486 1574
rect 8502 1564 8517 1568
rect 8535 1565 8574 1584
rect 8593 1578 8600 1579
rect 8599 1571 8600 1578
rect 8583 1568 8584 1571
rect 8599 1568 8612 1571
rect 8535 1564 8565 1565
rect 8574 1564 8580 1565
rect 8583 1564 8612 1568
rect 8502 1563 8612 1564
rect 8502 1562 8618 1563
rect 8177 1554 8228 1562
rect 8177 1542 8202 1554
rect 8209 1542 8228 1554
rect 8259 1554 8309 1562
rect 8259 1546 8275 1554
rect 8282 1552 8309 1554
rect 8318 1552 8539 1562
rect 8282 1542 8539 1552
rect 8568 1554 8618 1562
rect 8568 1545 8584 1554
rect 8177 1534 8228 1542
rect 8275 1534 8539 1542
rect 8565 1542 8584 1545
rect 8591 1542 8618 1554
rect 8565 1534 8618 1542
rect 8193 1526 8194 1534
rect 8209 1526 8222 1534
rect 8193 1518 8209 1526
rect 8190 1511 8209 1514
rect 8190 1502 8212 1511
rect 8163 1492 8212 1502
rect 8163 1486 8193 1492
rect 8212 1487 8217 1492
rect 8135 1470 8209 1486
rect 8227 1478 8257 1534
rect 8292 1524 8500 1534
rect 8535 1530 8580 1534
rect 8583 1533 8584 1534
rect 8599 1533 8612 1534
rect 8318 1494 8507 1524
rect 8333 1491 8507 1494
rect 8326 1488 8507 1491
rect 8135 1468 8148 1470
rect 8163 1468 8197 1470
rect 8135 1452 8209 1468
rect 8236 1464 8249 1478
rect 8264 1464 8280 1480
rect 8326 1475 8337 1488
rect 8119 1430 8120 1446
rect 8135 1430 8148 1452
rect 8163 1430 8193 1452
rect 8236 1448 8298 1464
rect 8326 1457 8337 1473
rect 8342 1468 8352 1488
rect 8362 1468 8376 1488
rect 8379 1475 8388 1488
rect 8404 1475 8413 1488
rect 8342 1457 8376 1468
rect 8379 1457 8388 1473
rect 8404 1457 8413 1473
rect 8420 1468 8430 1488
rect 8440 1468 8454 1488
rect 8455 1475 8466 1488
rect 8420 1457 8454 1468
rect 8455 1457 8466 1473
rect 8512 1464 8528 1480
rect 8535 1478 8565 1530
rect 8599 1526 8600 1533
rect 8584 1518 8600 1526
rect 8571 1486 8584 1505
rect 8599 1486 8629 1502
rect 8571 1470 8645 1486
rect 8571 1468 8584 1470
rect 8599 1468 8633 1470
rect 8236 1446 8249 1448
rect 8264 1446 8298 1448
rect 8236 1430 8298 1446
rect 8342 1441 8358 1444
rect 8420 1441 8450 1452
rect 8498 1448 8544 1464
rect 8571 1452 8645 1468
rect 8498 1446 8532 1448
rect 8497 1430 8544 1446
rect 8571 1430 8584 1452
rect 8599 1430 8629 1452
rect 8656 1430 8657 1446
rect 8672 1430 8685 1590
rect 8715 1486 8728 1590
rect 8773 1568 8774 1578
rect 8789 1568 8802 1578
rect 8773 1564 8802 1568
rect 8807 1564 8837 1590
rect 8855 1576 8871 1578
rect 8943 1576 8996 1590
rect 8944 1574 9008 1576
rect 9051 1574 9066 1590
rect 9115 1587 9145 1590
rect 9115 1584 9151 1587
rect 9081 1576 9097 1578
rect 8855 1564 8870 1568
rect 8773 1562 8870 1564
rect 8898 1562 9066 1574
rect 9082 1564 9097 1568
rect 9115 1565 9154 1584
rect 9173 1578 9180 1579
rect 9179 1571 9180 1578
rect 9163 1568 9164 1571
rect 9179 1568 9192 1571
rect 9115 1564 9145 1565
rect 9154 1564 9160 1565
rect 9163 1564 9192 1568
rect 9082 1563 9192 1564
rect 9082 1562 9198 1563
rect 8757 1554 8808 1562
rect 8757 1542 8782 1554
rect 8789 1542 8808 1554
rect 8839 1554 8889 1562
rect 8839 1546 8855 1554
rect 8862 1552 8889 1554
rect 8898 1552 9119 1562
rect 8862 1542 9119 1552
rect 9148 1554 9198 1562
rect 9148 1545 9164 1554
rect 8757 1534 8808 1542
rect 8855 1534 9119 1542
rect 9145 1542 9164 1545
rect 9171 1542 9198 1554
rect 9145 1534 9198 1542
rect 8773 1526 8774 1534
rect 8789 1526 8802 1534
rect 8773 1518 8789 1526
rect 8770 1511 8789 1514
rect 8770 1502 8792 1511
rect 8743 1492 8792 1502
rect 8743 1486 8773 1492
rect 8792 1487 8797 1492
rect 8715 1470 8789 1486
rect 8807 1478 8837 1534
rect 8872 1524 9080 1534
rect 9115 1530 9160 1534
rect 9163 1533 9164 1534
rect 9179 1533 9192 1534
rect 8898 1494 9087 1524
rect 8913 1491 9087 1494
rect 8906 1488 9087 1491
rect 8715 1468 8728 1470
rect 8743 1468 8777 1470
rect 8715 1452 8789 1468
rect 8816 1464 8829 1478
rect 8844 1464 8860 1480
rect 8906 1475 8917 1488
rect 8699 1430 8700 1446
rect 8715 1430 8728 1452
rect 8743 1430 8773 1452
rect 8816 1448 8878 1464
rect 8906 1457 8917 1473
rect 8922 1468 8932 1488
rect 8942 1468 8956 1488
rect 8959 1475 8968 1488
rect 8984 1475 8993 1488
rect 8922 1457 8956 1468
rect 8959 1457 8968 1473
rect 8984 1457 8993 1473
rect 9000 1468 9010 1488
rect 9020 1468 9034 1488
rect 9035 1475 9046 1488
rect 9000 1457 9034 1468
rect 9035 1457 9046 1473
rect 9092 1464 9108 1480
rect 9115 1478 9145 1530
rect 9179 1526 9180 1533
rect 9164 1518 9180 1526
rect 9151 1486 9164 1505
rect 9179 1486 9209 1502
rect 9151 1470 9225 1486
rect 9151 1468 9164 1470
rect 9179 1468 9213 1470
rect 8816 1446 8829 1448
rect 8844 1446 8878 1448
rect 8816 1430 8878 1446
rect 8922 1441 8938 1444
rect 9000 1441 9030 1452
rect 9078 1448 9124 1464
rect 9151 1452 9225 1468
rect 9078 1446 9112 1448
rect 9077 1430 9124 1446
rect 9151 1430 9164 1452
rect 9179 1430 9209 1452
rect 9236 1430 9237 1446
rect 9252 1430 9265 1590
rect -7 1422 34 1430
rect -7 1396 8 1422
rect 15 1396 34 1422
rect 98 1418 160 1430
rect 172 1418 247 1430
rect 305 1418 380 1430
rect 392 1418 423 1430
rect 429 1418 464 1430
rect 98 1416 260 1418
rect -7 1388 34 1396
rect 116 1392 129 1416
rect 144 1414 159 1416
rect -1 1378 0 1388
rect 15 1378 28 1388
rect 43 1378 73 1392
rect 116 1378 159 1392
rect 183 1389 190 1396
rect 193 1392 260 1416
rect 292 1416 464 1418
rect 262 1394 290 1398
rect 292 1394 372 1416
rect 393 1414 408 1416
rect 262 1392 372 1394
rect 193 1388 372 1392
rect 166 1378 196 1388
rect 198 1378 351 1388
rect 359 1378 389 1388
rect 393 1378 423 1392
rect 451 1378 464 1416
rect 536 1422 571 1430
rect 536 1396 537 1422
rect 544 1396 571 1422
rect 479 1378 509 1392
rect 536 1388 571 1396
rect 573 1422 614 1430
rect 573 1396 588 1422
rect 595 1396 614 1422
rect 678 1418 740 1430
rect 752 1418 827 1430
rect 885 1418 960 1430
rect 972 1418 1003 1430
rect 1009 1418 1044 1430
rect 678 1416 840 1418
rect 573 1388 614 1396
rect 696 1392 709 1416
rect 724 1414 739 1416
rect 536 1378 537 1388
rect 552 1378 565 1388
rect 579 1378 580 1388
rect 595 1378 608 1388
rect 623 1378 653 1392
rect 696 1378 739 1392
rect 763 1389 770 1396
rect 773 1392 840 1416
rect 872 1416 1044 1418
rect 842 1394 870 1398
rect 872 1394 952 1416
rect 973 1414 988 1416
rect 842 1392 952 1394
rect 773 1388 952 1392
rect 746 1378 776 1388
rect 778 1378 931 1388
rect 939 1378 969 1388
rect 973 1378 1003 1392
rect 1031 1378 1044 1416
rect 1116 1422 1151 1430
rect 1116 1396 1117 1422
rect 1124 1396 1151 1422
rect 1059 1378 1089 1392
rect 1116 1388 1151 1396
rect 1153 1422 1194 1430
rect 1153 1396 1168 1422
rect 1175 1396 1194 1422
rect 1258 1418 1320 1430
rect 1332 1418 1407 1430
rect 1465 1418 1540 1430
rect 1552 1418 1583 1430
rect 1589 1418 1624 1430
rect 1258 1416 1420 1418
rect 1153 1388 1194 1396
rect 1276 1392 1289 1416
rect 1304 1414 1319 1416
rect 1116 1378 1117 1388
rect 1132 1378 1145 1388
rect 1159 1378 1160 1388
rect 1175 1378 1188 1388
rect 1203 1378 1233 1392
rect 1276 1378 1319 1392
rect 1343 1389 1350 1396
rect 1353 1392 1420 1416
rect 1452 1416 1624 1418
rect 1422 1394 1450 1398
rect 1452 1394 1532 1416
rect 1553 1414 1568 1416
rect 1422 1392 1532 1394
rect 1353 1388 1532 1392
rect 1326 1378 1356 1388
rect 1358 1378 1511 1388
rect 1519 1378 1549 1388
rect 1553 1378 1583 1392
rect 1611 1378 1624 1416
rect 1696 1422 1731 1430
rect 1696 1396 1697 1422
rect 1704 1396 1731 1422
rect 1639 1378 1669 1392
rect 1696 1388 1731 1396
rect 1733 1422 1774 1430
rect 1733 1396 1748 1422
rect 1755 1396 1774 1422
rect 1838 1418 1900 1430
rect 1912 1418 1987 1430
rect 2045 1418 2120 1430
rect 2132 1418 2163 1430
rect 2169 1418 2204 1430
rect 1838 1416 2000 1418
rect 1733 1388 1774 1396
rect 1856 1392 1869 1416
rect 1884 1414 1899 1416
rect 1696 1378 1697 1388
rect 1712 1378 1725 1388
rect 1739 1378 1740 1388
rect 1755 1378 1768 1388
rect 1783 1378 1813 1392
rect 1856 1378 1899 1392
rect 1923 1389 1930 1396
rect 1933 1392 2000 1416
rect 2032 1416 2204 1418
rect 2002 1394 2030 1398
rect 2032 1394 2112 1416
rect 2133 1414 2148 1416
rect 2002 1392 2112 1394
rect 1933 1388 2112 1392
rect 1906 1378 1936 1388
rect 1938 1378 2091 1388
rect 2099 1378 2129 1388
rect 2133 1378 2163 1392
rect 2191 1378 2204 1416
rect 2276 1422 2311 1430
rect 2276 1396 2277 1422
rect 2284 1396 2311 1422
rect 2219 1378 2249 1392
rect 2276 1388 2311 1396
rect 2313 1422 2354 1430
rect 2313 1396 2328 1422
rect 2335 1396 2354 1422
rect 2418 1418 2480 1430
rect 2492 1418 2567 1430
rect 2625 1418 2700 1430
rect 2712 1418 2743 1430
rect 2749 1418 2784 1430
rect 2418 1416 2580 1418
rect 2313 1388 2354 1396
rect 2436 1392 2449 1416
rect 2464 1414 2479 1416
rect 2276 1378 2277 1388
rect 2292 1378 2305 1388
rect 2319 1378 2320 1388
rect 2335 1378 2348 1388
rect 2363 1378 2393 1392
rect 2436 1378 2479 1392
rect 2503 1389 2510 1396
rect 2513 1392 2580 1416
rect 2612 1416 2784 1418
rect 2582 1394 2610 1398
rect 2612 1394 2692 1416
rect 2713 1414 2728 1416
rect 2582 1392 2692 1394
rect 2513 1388 2692 1392
rect 2486 1378 2516 1388
rect 2518 1378 2671 1388
rect 2679 1378 2709 1388
rect 2713 1378 2743 1392
rect 2771 1378 2784 1416
rect 2856 1422 2891 1430
rect 2856 1396 2857 1422
rect 2864 1396 2891 1422
rect 2799 1378 2829 1392
rect 2856 1388 2891 1396
rect 2893 1422 2934 1430
rect 2893 1396 2908 1422
rect 2915 1396 2934 1422
rect 2998 1418 3060 1430
rect 3072 1418 3147 1430
rect 3205 1418 3280 1430
rect 3292 1418 3323 1430
rect 3329 1418 3364 1430
rect 2998 1416 3160 1418
rect 2893 1388 2934 1396
rect 3016 1392 3029 1416
rect 3044 1414 3059 1416
rect 2856 1378 2857 1388
rect 2872 1378 2885 1388
rect 2899 1378 2900 1388
rect 2915 1378 2928 1388
rect 2943 1378 2973 1392
rect 3016 1378 3059 1392
rect 3083 1389 3090 1396
rect 3093 1392 3160 1416
rect 3192 1416 3364 1418
rect 3162 1394 3190 1398
rect 3192 1394 3272 1416
rect 3293 1414 3308 1416
rect 3162 1392 3272 1394
rect 3093 1388 3272 1392
rect 3066 1378 3096 1388
rect 3098 1378 3251 1388
rect 3259 1378 3289 1388
rect 3293 1378 3323 1392
rect 3351 1378 3364 1416
rect 3436 1422 3471 1430
rect 3436 1396 3437 1422
rect 3444 1396 3471 1422
rect 3379 1378 3409 1392
rect 3436 1388 3471 1396
rect 3473 1422 3514 1430
rect 3473 1396 3488 1422
rect 3495 1396 3514 1422
rect 3578 1418 3640 1430
rect 3652 1418 3727 1430
rect 3785 1418 3860 1430
rect 3872 1418 3903 1430
rect 3909 1418 3944 1430
rect 3578 1416 3740 1418
rect 3473 1388 3514 1396
rect 3596 1392 3609 1416
rect 3624 1414 3639 1416
rect 3436 1378 3437 1388
rect 3452 1378 3465 1388
rect 3479 1378 3480 1388
rect 3495 1378 3508 1388
rect 3523 1378 3553 1392
rect 3596 1378 3639 1392
rect 3663 1389 3670 1396
rect 3673 1392 3740 1416
rect 3772 1416 3944 1418
rect 3742 1394 3770 1398
rect 3772 1394 3852 1416
rect 3873 1414 3888 1416
rect 3742 1392 3852 1394
rect 3673 1388 3852 1392
rect 3646 1378 3676 1388
rect 3678 1378 3831 1388
rect 3839 1378 3869 1388
rect 3873 1378 3903 1392
rect 3931 1378 3944 1416
rect 4016 1422 4051 1430
rect 4016 1396 4017 1422
rect 4024 1396 4051 1422
rect 3959 1378 3989 1392
rect 4016 1388 4051 1396
rect 4053 1422 4094 1430
rect 4053 1396 4068 1422
rect 4075 1396 4094 1422
rect 4158 1418 4220 1430
rect 4232 1418 4307 1430
rect 4365 1418 4440 1430
rect 4452 1418 4483 1430
rect 4489 1418 4524 1430
rect 4158 1416 4320 1418
rect 4053 1388 4094 1396
rect 4176 1392 4189 1416
rect 4204 1414 4219 1416
rect 4016 1378 4017 1388
rect 4032 1378 4045 1388
rect 4059 1378 4060 1388
rect 4075 1378 4088 1388
rect 4103 1378 4133 1392
rect 4176 1378 4219 1392
rect 4243 1389 4250 1396
rect 4253 1392 4320 1416
rect 4352 1416 4524 1418
rect 4322 1394 4350 1398
rect 4352 1394 4432 1416
rect 4453 1414 4468 1416
rect 4322 1392 4432 1394
rect 4253 1388 4432 1392
rect 4226 1378 4256 1388
rect 4258 1378 4411 1388
rect 4419 1378 4449 1388
rect 4453 1378 4483 1392
rect 4511 1378 4524 1416
rect 4596 1422 4631 1430
rect 4596 1396 4597 1422
rect 4604 1396 4631 1422
rect 4539 1378 4569 1392
rect 4596 1388 4631 1396
rect 4633 1422 4674 1430
rect 4633 1396 4648 1422
rect 4655 1396 4674 1422
rect 4738 1418 4800 1430
rect 4812 1418 4887 1430
rect 4945 1418 5020 1430
rect 5032 1418 5063 1430
rect 5069 1418 5104 1430
rect 4738 1416 4900 1418
rect 4633 1388 4674 1396
rect 4756 1392 4769 1416
rect 4784 1414 4799 1416
rect 4596 1378 4597 1388
rect 4612 1378 4625 1388
rect 4639 1378 4640 1388
rect 4655 1378 4668 1388
rect 4683 1378 4713 1392
rect 4756 1378 4799 1392
rect 4823 1389 4830 1396
rect 4833 1392 4900 1416
rect 4932 1416 5104 1418
rect 4902 1394 4930 1398
rect 4932 1394 5012 1416
rect 5033 1414 5048 1416
rect 4902 1392 5012 1394
rect 4833 1388 5012 1392
rect 4806 1378 4836 1388
rect 4838 1378 4991 1388
rect 4999 1378 5029 1388
rect 5033 1378 5063 1392
rect 5091 1378 5104 1416
rect 5176 1422 5211 1430
rect 5176 1396 5177 1422
rect 5184 1396 5211 1422
rect 5119 1378 5149 1392
rect 5176 1388 5211 1396
rect 5213 1422 5254 1430
rect 5213 1396 5228 1422
rect 5235 1396 5254 1422
rect 5318 1418 5380 1430
rect 5392 1418 5467 1430
rect 5525 1418 5600 1430
rect 5612 1418 5643 1430
rect 5649 1418 5684 1430
rect 5318 1416 5480 1418
rect 5213 1388 5254 1396
rect 5336 1392 5349 1416
rect 5364 1414 5379 1416
rect 5176 1378 5177 1388
rect 5192 1378 5205 1388
rect 5219 1378 5220 1388
rect 5235 1378 5248 1388
rect 5263 1378 5293 1392
rect 5336 1378 5379 1392
rect 5403 1389 5410 1396
rect 5413 1392 5480 1416
rect 5512 1416 5684 1418
rect 5482 1394 5510 1398
rect 5512 1394 5592 1416
rect 5613 1414 5628 1416
rect 5482 1392 5592 1394
rect 5413 1388 5592 1392
rect 5386 1378 5416 1388
rect 5418 1378 5571 1388
rect 5579 1378 5609 1388
rect 5613 1378 5643 1392
rect 5671 1378 5684 1416
rect 5756 1422 5791 1430
rect 5756 1396 5757 1422
rect 5764 1396 5791 1422
rect 5699 1378 5729 1392
rect 5756 1388 5791 1396
rect 5793 1422 5834 1430
rect 5793 1396 5808 1422
rect 5815 1396 5834 1422
rect 5898 1418 5960 1430
rect 5972 1418 6047 1430
rect 6105 1418 6180 1430
rect 6192 1418 6223 1430
rect 6229 1418 6264 1430
rect 5898 1416 6060 1418
rect 5793 1388 5834 1396
rect 5916 1392 5929 1416
rect 5944 1414 5959 1416
rect 5756 1378 5757 1388
rect 5772 1378 5785 1388
rect 5799 1378 5800 1388
rect 5815 1378 5828 1388
rect 5843 1378 5873 1392
rect 5916 1378 5959 1392
rect 5983 1389 5990 1396
rect 5993 1392 6060 1416
rect 6092 1416 6264 1418
rect 6062 1394 6090 1398
rect 6092 1394 6172 1416
rect 6193 1414 6208 1416
rect 6062 1392 6172 1394
rect 5993 1388 6172 1392
rect 5966 1378 5996 1388
rect 5998 1378 6151 1388
rect 6159 1378 6189 1388
rect 6193 1378 6223 1392
rect 6251 1378 6264 1416
rect 6336 1422 6371 1430
rect 6336 1396 6337 1422
rect 6344 1396 6371 1422
rect 6279 1378 6309 1392
rect 6336 1388 6371 1396
rect 6373 1422 6414 1430
rect 6373 1396 6388 1422
rect 6395 1396 6414 1422
rect 6478 1418 6540 1430
rect 6552 1418 6627 1430
rect 6685 1418 6760 1430
rect 6772 1418 6803 1430
rect 6809 1418 6844 1430
rect 6478 1416 6640 1418
rect 6373 1388 6414 1396
rect 6496 1392 6509 1416
rect 6524 1414 6539 1416
rect 6336 1378 6337 1388
rect 6352 1378 6365 1388
rect 6379 1378 6380 1388
rect 6395 1378 6408 1388
rect 6423 1378 6453 1392
rect 6496 1378 6539 1392
rect 6563 1389 6570 1396
rect 6573 1392 6640 1416
rect 6672 1416 6844 1418
rect 6642 1394 6670 1398
rect 6672 1394 6752 1416
rect 6773 1414 6788 1416
rect 6642 1392 6752 1394
rect 6573 1388 6752 1392
rect 6546 1378 6576 1388
rect 6578 1378 6731 1388
rect 6739 1378 6769 1388
rect 6773 1378 6803 1392
rect 6831 1378 6844 1416
rect 6916 1422 6951 1430
rect 6916 1396 6917 1422
rect 6924 1396 6951 1422
rect 6859 1378 6889 1392
rect 6916 1388 6951 1396
rect 6953 1422 6994 1430
rect 6953 1396 6968 1422
rect 6975 1396 6994 1422
rect 7058 1418 7120 1430
rect 7132 1418 7207 1430
rect 7265 1418 7340 1430
rect 7352 1418 7383 1430
rect 7389 1418 7424 1430
rect 7058 1416 7220 1418
rect 6953 1388 6994 1396
rect 7076 1392 7089 1416
rect 7104 1414 7119 1416
rect 6916 1378 6917 1388
rect 6932 1378 6945 1388
rect 6959 1378 6960 1388
rect 6975 1378 6988 1388
rect 7003 1378 7033 1392
rect 7076 1378 7119 1392
rect 7143 1389 7150 1396
rect 7153 1392 7220 1416
rect 7252 1416 7424 1418
rect 7222 1394 7250 1398
rect 7252 1394 7332 1416
rect 7353 1414 7368 1416
rect 7222 1392 7332 1394
rect 7153 1388 7332 1392
rect 7126 1378 7156 1388
rect 7158 1378 7311 1388
rect 7319 1378 7349 1388
rect 7353 1378 7383 1392
rect 7411 1378 7424 1416
rect 7496 1422 7531 1430
rect 7496 1396 7497 1422
rect 7504 1396 7531 1422
rect 7439 1378 7469 1392
rect 7496 1388 7531 1396
rect 7533 1422 7574 1430
rect 7533 1396 7548 1422
rect 7555 1396 7574 1422
rect 7638 1418 7700 1430
rect 7712 1418 7787 1430
rect 7845 1418 7920 1430
rect 7932 1418 7963 1430
rect 7969 1418 8004 1430
rect 7638 1416 7800 1418
rect 7533 1388 7574 1396
rect 7656 1392 7669 1416
rect 7684 1414 7699 1416
rect 7496 1378 7497 1388
rect 7512 1378 7525 1388
rect 7539 1378 7540 1388
rect 7555 1378 7568 1388
rect 7583 1378 7613 1392
rect 7656 1378 7699 1392
rect 7723 1389 7730 1396
rect 7733 1392 7800 1416
rect 7832 1416 8004 1418
rect 7802 1394 7830 1398
rect 7832 1394 7912 1416
rect 7933 1414 7948 1416
rect 7802 1392 7912 1394
rect 7733 1388 7912 1392
rect 7706 1378 7736 1388
rect 7738 1378 7891 1388
rect 7899 1378 7929 1388
rect 7933 1378 7963 1392
rect 7991 1378 8004 1416
rect 8076 1422 8111 1430
rect 8076 1396 8077 1422
rect 8084 1396 8111 1422
rect 8019 1378 8049 1392
rect 8076 1388 8111 1396
rect 8113 1422 8154 1430
rect 8113 1396 8128 1422
rect 8135 1396 8154 1422
rect 8218 1418 8280 1430
rect 8292 1418 8367 1430
rect 8425 1418 8500 1430
rect 8512 1418 8543 1430
rect 8549 1418 8584 1430
rect 8218 1416 8380 1418
rect 8113 1388 8154 1396
rect 8236 1392 8249 1416
rect 8264 1414 8279 1416
rect 8076 1378 8077 1388
rect 8092 1378 8105 1388
rect 8119 1378 8120 1388
rect 8135 1378 8148 1388
rect 8163 1378 8193 1392
rect 8236 1378 8279 1392
rect 8303 1389 8310 1396
rect 8313 1392 8380 1416
rect 8412 1416 8584 1418
rect 8382 1394 8410 1398
rect 8412 1394 8492 1416
rect 8513 1414 8528 1416
rect 8382 1392 8492 1394
rect 8313 1388 8492 1392
rect 8286 1378 8316 1388
rect 8318 1378 8471 1388
rect 8479 1378 8509 1388
rect 8513 1378 8543 1392
rect 8571 1378 8584 1416
rect 8656 1422 8691 1430
rect 8656 1396 8657 1422
rect 8664 1396 8691 1422
rect 8599 1378 8629 1392
rect 8656 1388 8691 1396
rect 8693 1422 8734 1430
rect 8693 1396 8708 1422
rect 8715 1396 8734 1422
rect 8798 1418 8860 1430
rect 8872 1418 8947 1430
rect 9005 1418 9080 1430
rect 9092 1418 9123 1430
rect 9129 1418 9164 1430
rect 8798 1416 8960 1418
rect 8693 1388 8734 1396
rect 8816 1392 8829 1416
rect 8844 1414 8859 1416
rect 8656 1378 8657 1388
rect 8672 1378 8685 1388
rect 8699 1378 8700 1388
rect 8715 1378 8728 1388
rect 8743 1378 8773 1392
rect 8816 1378 8859 1392
rect 8883 1389 8890 1396
rect 8893 1392 8960 1416
rect 8992 1416 9164 1418
rect 8962 1394 8990 1398
rect 8992 1394 9072 1416
rect 9093 1414 9108 1416
rect 8962 1392 9072 1394
rect 8893 1388 9072 1392
rect 8866 1378 8896 1388
rect 8898 1378 9051 1388
rect 9059 1378 9089 1388
rect 9093 1378 9123 1392
rect 9151 1378 9164 1416
rect 9236 1422 9271 1430
rect 9236 1396 9237 1422
rect 9244 1396 9271 1422
rect 9179 1378 9209 1392
rect 9236 1388 9271 1396
rect 9236 1378 9237 1388
rect 9252 1378 9265 1388
rect -1 1372 9265 1378
rect 0 1364 9265 1372
rect 15 1334 28 1364
rect 43 1346 73 1364
rect 116 1350 130 1364
rect 166 1350 386 1364
rect 117 1348 130 1350
rect 83 1336 98 1348
rect 80 1334 102 1336
rect 107 1334 137 1348
rect 198 1346 351 1350
rect 180 1334 372 1346
rect 415 1334 445 1348
rect 451 1334 464 1364
rect 479 1346 509 1364
rect 552 1334 565 1364
rect 595 1334 608 1364
rect 623 1346 653 1364
rect 696 1350 710 1364
rect 746 1350 966 1364
rect 697 1348 710 1350
rect 663 1336 678 1348
rect 660 1334 682 1336
rect 687 1334 717 1348
rect 778 1346 931 1350
rect 760 1334 952 1346
rect 995 1334 1025 1348
rect 1031 1334 1044 1364
rect 1059 1346 1089 1364
rect 1132 1334 1145 1364
rect 1175 1334 1188 1364
rect 1203 1346 1233 1364
rect 1276 1350 1290 1364
rect 1326 1350 1546 1364
rect 1277 1348 1290 1350
rect 1243 1336 1258 1348
rect 1240 1334 1262 1336
rect 1267 1334 1297 1348
rect 1358 1346 1511 1350
rect 1340 1334 1532 1346
rect 1575 1334 1605 1348
rect 1611 1334 1624 1364
rect 1639 1346 1669 1364
rect 1712 1334 1725 1364
rect 1755 1334 1768 1364
rect 1783 1346 1813 1364
rect 1856 1350 1870 1364
rect 1906 1350 2126 1364
rect 1857 1348 1870 1350
rect 1823 1336 1838 1348
rect 1820 1334 1842 1336
rect 1847 1334 1877 1348
rect 1938 1346 2091 1350
rect 1920 1334 2112 1346
rect 2155 1334 2185 1348
rect 2191 1334 2204 1364
rect 2219 1346 2249 1364
rect 2292 1334 2305 1364
rect 2335 1334 2348 1364
rect 2363 1346 2393 1364
rect 2436 1350 2450 1364
rect 2486 1350 2706 1364
rect 2437 1348 2450 1350
rect 2403 1336 2418 1348
rect 2400 1334 2422 1336
rect 2427 1334 2457 1348
rect 2518 1346 2671 1350
rect 2500 1334 2692 1346
rect 2735 1334 2765 1348
rect 2771 1334 2784 1364
rect 2799 1346 2829 1364
rect 2872 1334 2885 1364
rect 2915 1334 2928 1364
rect 2943 1346 2973 1364
rect 3016 1350 3030 1364
rect 3066 1350 3286 1364
rect 3017 1348 3030 1350
rect 2983 1336 2998 1348
rect 2980 1334 3002 1336
rect 3007 1334 3037 1348
rect 3098 1346 3251 1350
rect 3080 1334 3272 1346
rect 3315 1334 3345 1348
rect 3351 1334 3364 1364
rect 3379 1346 3409 1364
rect 3452 1334 3465 1364
rect 3495 1334 3508 1364
rect 3523 1346 3553 1364
rect 3596 1350 3610 1364
rect 3646 1350 3866 1364
rect 3597 1348 3610 1350
rect 3563 1336 3578 1348
rect 3560 1334 3582 1336
rect 3587 1334 3617 1348
rect 3678 1346 3831 1350
rect 3660 1334 3852 1346
rect 3895 1334 3925 1348
rect 3931 1334 3944 1364
rect 3959 1346 3989 1364
rect 4032 1334 4045 1364
rect 4075 1334 4088 1364
rect 4103 1346 4133 1364
rect 4176 1350 4190 1364
rect 4226 1350 4446 1364
rect 4177 1348 4190 1350
rect 4143 1336 4158 1348
rect 4140 1334 4162 1336
rect 4167 1334 4197 1348
rect 4258 1346 4411 1350
rect 4240 1334 4432 1346
rect 4475 1334 4505 1348
rect 4511 1334 4524 1364
rect 4539 1346 4569 1364
rect 4612 1334 4625 1364
rect 4655 1334 4668 1364
rect 4683 1346 4713 1364
rect 4756 1350 4770 1364
rect 4806 1350 5026 1364
rect 4757 1348 4770 1350
rect 4723 1336 4738 1348
rect 4720 1334 4742 1336
rect 4747 1334 4777 1348
rect 4838 1346 4991 1350
rect 4820 1334 5012 1346
rect 5055 1334 5085 1348
rect 5091 1334 5104 1364
rect 5119 1346 5149 1364
rect 5192 1334 5205 1364
rect 5235 1334 5248 1364
rect 5263 1346 5293 1364
rect 5336 1350 5350 1364
rect 5386 1350 5606 1364
rect 5337 1348 5350 1350
rect 5303 1336 5318 1348
rect 5300 1334 5322 1336
rect 5327 1334 5357 1348
rect 5418 1346 5571 1350
rect 5400 1334 5592 1346
rect 5635 1334 5665 1348
rect 5671 1334 5684 1364
rect 5699 1346 5729 1364
rect 5772 1334 5785 1364
rect 5815 1334 5828 1364
rect 5843 1346 5873 1364
rect 5916 1350 5930 1364
rect 5966 1350 6186 1364
rect 5917 1348 5930 1350
rect 5883 1336 5898 1348
rect 5880 1334 5902 1336
rect 5907 1334 5937 1348
rect 5998 1346 6151 1350
rect 5980 1334 6172 1346
rect 6215 1334 6245 1348
rect 6251 1334 6264 1364
rect 6279 1346 6309 1364
rect 6352 1334 6365 1364
rect 6395 1334 6408 1364
rect 6423 1346 6453 1364
rect 6496 1350 6510 1364
rect 6546 1350 6766 1364
rect 6497 1348 6510 1350
rect 6463 1336 6478 1348
rect 6460 1334 6482 1336
rect 6487 1334 6517 1348
rect 6578 1346 6731 1350
rect 6560 1334 6752 1346
rect 6795 1334 6825 1348
rect 6831 1334 6844 1364
rect 6859 1346 6889 1364
rect 6932 1334 6945 1364
rect 6975 1334 6988 1364
rect 7003 1346 7033 1364
rect 7076 1350 7090 1364
rect 7126 1350 7346 1364
rect 7077 1348 7090 1350
rect 7043 1336 7058 1348
rect 7040 1334 7062 1336
rect 7067 1334 7097 1348
rect 7158 1346 7311 1350
rect 7140 1334 7332 1346
rect 7375 1334 7405 1348
rect 7411 1334 7424 1364
rect 7439 1346 7469 1364
rect 7512 1334 7525 1364
rect 7555 1334 7568 1364
rect 7583 1346 7613 1364
rect 7656 1350 7670 1364
rect 7706 1350 7926 1364
rect 7657 1348 7670 1350
rect 7623 1336 7638 1348
rect 7620 1334 7642 1336
rect 7647 1334 7677 1348
rect 7738 1346 7891 1350
rect 7720 1334 7912 1346
rect 7955 1334 7985 1348
rect 7991 1334 8004 1364
rect 8019 1346 8049 1364
rect 8092 1334 8105 1364
rect 8135 1334 8148 1364
rect 8163 1346 8193 1364
rect 8236 1350 8250 1364
rect 8286 1350 8506 1364
rect 8237 1348 8250 1350
rect 8203 1336 8218 1348
rect 8200 1334 8222 1336
rect 8227 1334 8257 1348
rect 8318 1346 8471 1350
rect 8300 1334 8492 1346
rect 8535 1334 8565 1348
rect 8571 1334 8584 1364
rect 8599 1346 8629 1364
rect 8672 1334 8685 1364
rect 8715 1334 8728 1364
rect 8743 1346 8773 1364
rect 8816 1350 8830 1364
rect 8866 1350 9086 1364
rect 8817 1348 8830 1350
rect 8783 1336 8798 1348
rect 8780 1334 8802 1336
rect 8807 1334 8837 1348
rect 8898 1346 9051 1350
rect 8880 1334 9072 1346
rect 9115 1334 9145 1348
rect 9151 1334 9164 1364
rect 9179 1346 9209 1364
rect 9252 1334 9265 1364
rect 0 1320 9265 1334
rect 15 1216 28 1320
rect 73 1298 74 1308
rect 89 1298 102 1308
rect 73 1294 102 1298
rect 107 1294 137 1320
rect 155 1306 171 1308
rect 243 1306 296 1320
rect 244 1304 308 1306
rect 351 1304 366 1320
rect 415 1317 445 1320
rect 415 1314 451 1317
rect 381 1306 397 1308
rect 155 1294 170 1298
rect 73 1292 170 1294
rect 198 1292 366 1304
rect 382 1294 397 1298
rect 415 1295 454 1314
rect 473 1308 480 1309
rect 479 1301 480 1308
rect 463 1298 464 1301
rect 479 1298 492 1301
rect 415 1294 445 1295
rect 454 1294 460 1295
rect 463 1294 492 1298
rect 382 1293 492 1294
rect 382 1292 498 1293
rect 57 1284 108 1292
rect 57 1272 82 1284
rect 89 1272 108 1284
rect 139 1284 189 1292
rect 139 1276 155 1284
rect 162 1282 189 1284
rect 198 1282 419 1292
rect 162 1272 419 1282
rect 448 1284 498 1292
rect 448 1275 464 1284
rect 57 1264 108 1272
rect 155 1264 419 1272
rect 445 1272 464 1275
rect 471 1272 498 1284
rect 445 1264 498 1272
rect 73 1256 74 1264
rect 89 1256 102 1264
rect 73 1248 89 1256
rect 70 1241 89 1244
rect 70 1232 92 1241
rect 43 1222 92 1232
rect 43 1216 73 1222
rect 92 1217 97 1222
rect 15 1200 89 1216
rect 107 1208 137 1264
rect 172 1254 380 1264
rect 415 1260 460 1264
rect 463 1263 464 1264
rect 479 1263 492 1264
rect 198 1224 387 1254
rect 213 1221 387 1224
rect 206 1218 387 1221
rect 15 1198 28 1200
rect 43 1198 77 1200
rect 15 1182 89 1198
rect 116 1194 129 1208
rect 144 1194 160 1210
rect 206 1205 217 1218
rect -1 1160 0 1176
rect 15 1160 28 1182
rect 43 1160 73 1182
rect 116 1178 178 1194
rect 206 1187 217 1203
rect 222 1198 232 1218
rect 242 1198 256 1218
rect 259 1205 268 1218
rect 284 1205 293 1218
rect 222 1187 256 1198
rect 259 1187 268 1203
rect 284 1187 293 1203
rect 300 1198 310 1218
rect 320 1198 334 1218
rect 335 1205 346 1218
rect 300 1187 334 1198
rect 335 1187 346 1203
rect 392 1194 408 1210
rect 415 1208 445 1260
rect 479 1256 480 1263
rect 464 1248 480 1256
rect 451 1216 464 1235
rect 479 1216 509 1232
rect 451 1200 525 1216
rect 451 1198 464 1200
rect 479 1198 513 1200
rect 116 1176 129 1178
rect 144 1176 178 1178
rect 116 1160 178 1176
rect 222 1171 238 1174
rect 300 1171 330 1182
rect 378 1178 424 1194
rect 451 1182 525 1198
rect 378 1176 412 1178
rect 377 1160 424 1176
rect 451 1160 464 1182
rect 479 1160 509 1182
rect 536 1160 537 1176
rect 552 1160 565 1320
rect 595 1216 608 1320
rect 653 1298 654 1308
rect 669 1298 682 1308
rect 653 1294 682 1298
rect 687 1294 717 1320
rect 735 1306 751 1308
rect 823 1306 876 1320
rect 824 1304 888 1306
rect 931 1304 946 1320
rect 995 1317 1025 1320
rect 995 1314 1031 1317
rect 961 1306 977 1308
rect 735 1294 750 1298
rect 653 1292 750 1294
rect 778 1292 946 1304
rect 962 1294 977 1298
rect 995 1295 1034 1314
rect 1053 1308 1060 1309
rect 1059 1301 1060 1308
rect 1043 1298 1044 1301
rect 1059 1298 1072 1301
rect 995 1294 1025 1295
rect 1034 1294 1040 1295
rect 1043 1294 1072 1298
rect 962 1293 1072 1294
rect 962 1292 1078 1293
rect 637 1284 688 1292
rect 637 1272 662 1284
rect 669 1272 688 1284
rect 719 1284 769 1292
rect 719 1276 735 1284
rect 742 1282 769 1284
rect 778 1282 999 1292
rect 742 1272 999 1282
rect 1028 1284 1078 1292
rect 1028 1275 1044 1284
rect 637 1264 688 1272
rect 735 1264 999 1272
rect 1025 1272 1044 1275
rect 1051 1272 1078 1284
rect 1025 1264 1078 1272
rect 653 1256 654 1264
rect 669 1256 682 1264
rect 653 1248 669 1256
rect 650 1241 669 1244
rect 650 1232 672 1241
rect 623 1222 672 1232
rect 623 1216 653 1222
rect 672 1217 677 1222
rect 595 1200 669 1216
rect 687 1208 717 1264
rect 752 1254 960 1264
rect 995 1260 1040 1264
rect 1043 1263 1044 1264
rect 1059 1263 1072 1264
rect 778 1224 967 1254
rect 793 1221 967 1224
rect 786 1218 967 1221
rect 595 1198 608 1200
rect 623 1198 657 1200
rect 595 1182 669 1198
rect 696 1194 709 1208
rect 724 1194 740 1210
rect 786 1205 797 1218
rect 579 1160 580 1176
rect 595 1160 608 1182
rect 623 1160 653 1182
rect 696 1178 758 1194
rect 786 1187 797 1203
rect 802 1198 812 1218
rect 822 1198 836 1218
rect 839 1205 848 1218
rect 864 1205 873 1218
rect 802 1187 836 1198
rect 839 1187 848 1203
rect 864 1187 873 1203
rect 880 1198 890 1218
rect 900 1198 914 1218
rect 915 1205 926 1218
rect 880 1187 914 1198
rect 915 1187 926 1203
rect 972 1194 988 1210
rect 995 1208 1025 1260
rect 1059 1256 1060 1263
rect 1044 1248 1060 1256
rect 1031 1216 1044 1235
rect 1059 1216 1089 1232
rect 1031 1200 1105 1216
rect 1031 1198 1044 1200
rect 1059 1198 1093 1200
rect 696 1176 709 1178
rect 724 1176 758 1178
rect 696 1160 758 1176
rect 802 1171 818 1174
rect 880 1171 910 1182
rect 958 1178 1004 1194
rect 1031 1182 1105 1198
rect 958 1176 992 1178
rect 957 1160 1004 1176
rect 1031 1160 1044 1182
rect 1059 1160 1089 1182
rect 1116 1160 1117 1176
rect 1132 1160 1145 1320
rect 1175 1216 1188 1320
rect 1233 1298 1234 1308
rect 1249 1298 1262 1308
rect 1233 1294 1262 1298
rect 1267 1294 1297 1320
rect 1315 1306 1331 1308
rect 1403 1306 1456 1320
rect 1404 1304 1468 1306
rect 1511 1304 1526 1320
rect 1575 1317 1605 1320
rect 1575 1314 1611 1317
rect 1541 1306 1557 1308
rect 1315 1294 1330 1298
rect 1233 1292 1330 1294
rect 1358 1292 1526 1304
rect 1542 1294 1557 1298
rect 1575 1295 1614 1314
rect 1633 1308 1640 1309
rect 1639 1301 1640 1308
rect 1623 1298 1624 1301
rect 1639 1298 1652 1301
rect 1575 1294 1605 1295
rect 1614 1294 1620 1295
rect 1623 1294 1652 1298
rect 1542 1293 1652 1294
rect 1542 1292 1658 1293
rect 1217 1284 1268 1292
rect 1217 1272 1242 1284
rect 1249 1272 1268 1284
rect 1299 1284 1349 1292
rect 1299 1276 1315 1284
rect 1322 1282 1349 1284
rect 1358 1282 1579 1292
rect 1322 1272 1579 1282
rect 1608 1284 1658 1292
rect 1608 1275 1624 1284
rect 1217 1264 1268 1272
rect 1315 1264 1579 1272
rect 1605 1272 1624 1275
rect 1631 1272 1658 1284
rect 1605 1264 1658 1272
rect 1233 1256 1234 1264
rect 1249 1256 1262 1264
rect 1233 1248 1249 1256
rect 1230 1241 1249 1244
rect 1230 1232 1252 1241
rect 1203 1222 1252 1232
rect 1203 1216 1233 1222
rect 1252 1217 1257 1222
rect 1175 1200 1249 1216
rect 1267 1208 1297 1264
rect 1332 1254 1540 1264
rect 1575 1260 1620 1264
rect 1623 1263 1624 1264
rect 1639 1263 1652 1264
rect 1358 1224 1547 1254
rect 1373 1221 1547 1224
rect 1366 1218 1547 1221
rect 1175 1198 1188 1200
rect 1203 1198 1237 1200
rect 1175 1182 1249 1198
rect 1276 1194 1289 1208
rect 1304 1194 1320 1210
rect 1366 1205 1377 1218
rect 1159 1160 1160 1176
rect 1175 1160 1188 1182
rect 1203 1160 1233 1182
rect 1276 1178 1338 1194
rect 1366 1187 1377 1203
rect 1382 1198 1392 1218
rect 1402 1198 1416 1218
rect 1419 1205 1428 1218
rect 1444 1205 1453 1218
rect 1382 1187 1416 1198
rect 1419 1187 1428 1203
rect 1444 1187 1453 1203
rect 1460 1198 1470 1218
rect 1480 1198 1494 1218
rect 1495 1205 1506 1218
rect 1460 1187 1494 1198
rect 1495 1187 1506 1203
rect 1552 1194 1568 1210
rect 1575 1208 1605 1260
rect 1639 1256 1640 1263
rect 1624 1248 1640 1256
rect 1611 1216 1624 1235
rect 1639 1216 1669 1232
rect 1611 1200 1685 1216
rect 1611 1198 1624 1200
rect 1639 1198 1673 1200
rect 1276 1176 1289 1178
rect 1304 1176 1338 1178
rect 1276 1160 1338 1176
rect 1382 1171 1398 1174
rect 1460 1171 1490 1182
rect 1538 1178 1584 1194
rect 1611 1182 1685 1198
rect 1538 1176 1572 1178
rect 1537 1160 1584 1176
rect 1611 1160 1624 1182
rect 1639 1160 1669 1182
rect 1696 1160 1697 1176
rect 1712 1160 1725 1320
rect 1755 1216 1768 1320
rect 1813 1298 1814 1308
rect 1829 1298 1842 1308
rect 1813 1294 1842 1298
rect 1847 1294 1877 1320
rect 1895 1306 1911 1308
rect 1983 1306 2036 1320
rect 1984 1304 2048 1306
rect 2091 1304 2106 1320
rect 2155 1317 2185 1320
rect 2155 1314 2191 1317
rect 2121 1306 2137 1308
rect 1895 1294 1910 1298
rect 1813 1292 1910 1294
rect 1938 1292 2106 1304
rect 2122 1294 2137 1298
rect 2155 1295 2194 1314
rect 2213 1308 2220 1309
rect 2219 1301 2220 1308
rect 2203 1298 2204 1301
rect 2219 1298 2232 1301
rect 2155 1294 2185 1295
rect 2194 1294 2200 1295
rect 2203 1294 2232 1298
rect 2122 1293 2232 1294
rect 2122 1292 2238 1293
rect 1797 1284 1848 1292
rect 1797 1272 1822 1284
rect 1829 1272 1848 1284
rect 1879 1284 1929 1292
rect 1879 1276 1895 1284
rect 1902 1282 1929 1284
rect 1938 1282 2159 1292
rect 1902 1272 2159 1282
rect 2188 1284 2238 1292
rect 2188 1275 2204 1284
rect 1797 1264 1848 1272
rect 1895 1264 2159 1272
rect 2185 1272 2204 1275
rect 2211 1272 2238 1284
rect 2185 1264 2238 1272
rect 1813 1256 1814 1264
rect 1829 1256 1842 1264
rect 1813 1248 1829 1256
rect 1810 1241 1829 1244
rect 1810 1232 1832 1241
rect 1783 1222 1832 1232
rect 1783 1216 1813 1222
rect 1832 1217 1837 1222
rect 1755 1200 1829 1216
rect 1847 1208 1877 1264
rect 1912 1254 2120 1264
rect 2155 1260 2200 1264
rect 2203 1263 2204 1264
rect 2219 1263 2232 1264
rect 1938 1224 2127 1254
rect 1953 1221 2127 1224
rect 1946 1218 2127 1221
rect 1755 1198 1768 1200
rect 1783 1198 1817 1200
rect 1755 1182 1829 1198
rect 1856 1194 1869 1208
rect 1884 1194 1900 1210
rect 1946 1205 1957 1218
rect 1739 1160 1740 1176
rect 1755 1160 1768 1182
rect 1783 1160 1813 1182
rect 1856 1178 1918 1194
rect 1946 1187 1957 1203
rect 1962 1198 1972 1218
rect 1982 1198 1996 1218
rect 1999 1205 2008 1218
rect 2024 1205 2033 1218
rect 1962 1187 1996 1198
rect 1999 1187 2008 1203
rect 2024 1187 2033 1203
rect 2040 1198 2050 1218
rect 2060 1198 2074 1218
rect 2075 1205 2086 1218
rect 2040 1187 2074 1198
rect 2075 1187 2086 1203
rect 2132 1194 2148 1210
rect 2155 1208 2185 1260
rect 2219 1256 2220 1263
rect 2204 1248 2220 1256
rect 2191 1216 2204 1235
rect 2219 1216 2249 1232
rect 2191 1200 2265 1216
rect 2191 1198 2204 1200
rect 2219 1198 2253 1200
rect 1856 1176 1869 1178
rect 1884 1176 1918 1178
rect 1856 1160 1918 1176
rect 1962 1171 1976 1174
rect 2040 1171 2070 1182
rect 2118 1178 2164 1194
rect 2191 1182 2265 1198
rect 2118 1176 2152 1178
rect 2117 1160 2164 1176
rect 2191 1160 2204 1182
rect 2219 1160 2249 1182
rect 2276 1160 2277 1176
rect 2292 1160 2305 1320
rect 2335 1216 2348 1320
rect 2393 1298 2394 1308
rect 2409 1298 2422 1308
rect 2393 1294 2422 1298
rect 2427 1294 2457 1320
rect 2475 1306 2491 1308
rect 2563 1306 2616 1320
rect 2564 1304 2628 1306
rect 2671 1304 2686 1320
rect 2735 1317 2765 1320
rect 2735 1314 2771 1317
rect 2701 1306 2717 1308
rect 2475 1294 2490 1298
rect 2393 1292 2490 1294
rect 2518 1292 2686 1304
rect 2702 1294 2717 1298
rect 2735 1295 2774 1314
rect 2793 1308 2800 1309
rect 2799 1301 2800 1308
rect 2783 1298 2784 1301
rect 2799 1298 2812 1301
rect 2735 1294 2765 1295
rect 2774 1294 2780 1295
rect 2783 1294 2812 1298
rect 2702 1293 2812 1294
rect 2702 1292 2818 1293
rect 2377 1284 2428 1292
rect 2377 1272 2402 1284
rect 2409 1272 2428 1284
rect 2459 1284 2509 1292
rect 2459 1276 2475 1284
rect 2482 1282 2509 1284
rect 2518 1282 2739 1292
rect 2482 1272 2739 1282
rect 2768 1284 2818 1292
rect 2768 1275 2784 1284
rect 2377 1264 2428 1272
rect 2475 1264 2739 1272
rect 2765 1272 2784 1275
rect 2791 1272 2818 1284
rect 2765 1264 2818 1272
rect 2393 1256 2394 1264
rect 2409 1256 2422 1264
rect 2393 1248 2409 1256
rect 2390 1241 2409 1244
rect 2390 1232 2412 1241
rect 2363 1222 2412 1232
rect 2363 1216 2393 1222
rect 2412 1217 2417 1222
rect 2335 1200 2409 1216
rect 2427 1208 2457 1264
rect 2492 1254 2700 1264
rect 2735 1260 2780 1264
rect 2783 1263 2784 1264
rect 2799 1263 2812 1264
rect 2518 1224 2707 1254
rect 2533 1221 2707 1224
rect 2526 1218 2707 1221
rect 2335 1198 2348 1200
rect 2363 1198 2397 1200
rect 2335 1182 2409 1198
rect 2436 1194 2449 1208
rect 2464 1194 2480 1210
rect 2526 1205 2537 1218
rect 2319 1160 2320 1176
rect 2335 1160 2348 1182
rect 2363 1160 2393 1182
rect 2436 1178 2498 1194
rect 2526 1187 2537 1203
rect 2542 1198 2552 1218
rect 2562 1198 2576 1218
rect 2579 1205 2588 1218
rect 2604 1205 2613 1218
rect 2542 1187 2576 1198
rect 2579 1187 2588 1203
rect 2604 1187 2613 1203
rect 2620 1198 2630 1218
rect 2640 1198 2654 1218
rect 2655 1205 2666 1218
rect 2620 1187 2654 1198
rect 2655 1187 2666 1203
rect 2712 1194 2728 1210
rect 2735 1208 2765 1260
rect 2799 1256 2800 1263
rect 2784 1248 2800 1256
rect 2771 1216 2784 1235
rect 2799 1216 2829 1232
rect 2771 1200 2845 1216
rect 2771 1198 2784 1200
rect 2799 1198 2833 1200
rect 2436 1176 2449 1178
rect 2464 1176 2498 1178
rect 2436 1160 2498 1176
rect 2542 1171 2558 1174
rect 2620 1171 2650 1182
rect 2698 1178 2744 1194
rect 2771 1182 2845 1198
rect 2698 1176 2732 1178
rect 2697 1160 2744 1176
rect 2771 1160 2784 1182
rect 2799 1160 2829 1182
rect 2856 1160 2857 1176
rect 2872 1160 2885 1320
rect 2915 1216 2928 1320
rect 2973 1298 2974 1308
rect 2989 1298 3002 1308
rect 2973 1294 3002 1298
rect 3007 1294 3037 1320
rect 3055 1306 3071 1308
rect 3143 1306 3196 1320
rect 3144 1304 3208 1306
rect 3251 1304 3266 1320
rect 3315 1317 3345 1320
rect 3315 1314 3351 1317
rect 3281 1306 3297 1308
rect 3055 1294 3070 1298
rect 2973 1292 3070 1294
rect 3098 1292 3266 1304
rect 3282 1294 3297 1298
rect 3315 1295 3354 1314
rect 3373 1308 3380 1309
rect 3379 1301 3380 1308
rect 3363 1298 3364 1301
rect 3379 1298 3392 1301
rect 3315 1294 3345 1295
rect 3354 1294 3360 1295
rect 3363 1294 3392 1298
rect 3282 1293 3392 1294
rect 3282 1292 3398 1293
rect 2957 1284 3008 1292
rect 2957 1272 2982 1284
rect 2989 1272 3008 1284
rect 3039 1284 3089 1292
rect 3039 1276 3055 1284
rect 3062 1282 3089 1284
rect 3098 1282 3319 1292
rect 3062 1272 3319 1282
rect 3348 1284 3398 1292
rect 3348 1275 3364 1284
rect 2957 1264 3008 1272
rect 3055 1264 3319 1272
rect 3345 1272 3364 1275
rect 3371 1272 3398 1284
rect 3345 1264 3398 1272
rect 2973 1256 2974 1264
rect 2989 1256 3002 1264
rect 2973 1248 2989 1256
rect 2970 1241 2989 1244
rect 2970 1232 2992 1241
rect 2943 1222 2992 1232
rect 2943 1216 2973 1222
rect 2992 1217 2997 1222
rect 2915 1200 2989 1216
rect 3007 1208 3037 1264
rect 3072 1254 3280 1264
rect 3315 1260 3360 1264
rect 3363 1263 3364 1264
rect 3379 1263 3392 1264
rect 3098 1224 3287 1254
rect 3113 1221 3287 1224
rect 3106 1218 3287 1221
rect 2915 1198 2928 1200
rect 2943 1198 2977 1200
rect 2915 1182 2989 1198
rect 3016 1194 3029 1208
rect 3044 1194 3060 1210
rect 3106 1205 3117 1218
rect 2899 1160 2900 1176
rect 2915 1160 2928 1182
rect 2943 1160 2973 1182
rect 3016 1178 3078 1194
rect 3106 1187 3117 1203
rect 3122 1198 3132 1218
rect 3142 1198 3156 1218
rect 3159 1205 3168 1218
rect 3184 1205 3193 1218
rect 3122 1187 3156 1198
rect 3159 1187 3168 1203
rect 3184 1187 3193 1203
rect 3200 1198 3210 1218
rect 3220 1198 3234 1218
rect 3235 1205 3246 1218
rect 3200 1187 3234 1198
rect 3235 1187 3246 1203
rect 3292 1194 3308 1210
rect 3315 1208 3345 1260
rect 3379 1256 3380 1263
rect 3364 1248 3380 1256
rect 3351 1216 3364 1235
rect 3379 1216 3409 1232
rect 3351 1200 3425 1216
rect 3351 1198 3364 1200
rect 3379 1198 3413 1200
rect 3016 1176 3029 1178
rect 3044 1176 3078 1178
rect 3016 1160 3078 1176
rect 3122 1171 3138 1174
rect 3200 1171 3230 1182
rect 3278 1178 3324 1194
rect 3351 1182 3425 1198
rect 3278 1176 3312 1178
rect 3277 1160 3324 1176
rect 3351 1160 3364 1182
rect 3379 1160 3409 1182
rect 3436 1160 3437 1176
rect 3452 1160 3465 1320
rect 3495 1216 3508 1320
rect 3553 1298 3554 1308
rect 3569 1298 3582 1308
rect 3553 1294 3582 1298
rect 3587 1294 3617 1320
rect 3635 1306 3651 1308
rect 3723 1306 3776 1320
rect 3724 1304 3788 1306
rect 3831 1304 3846 1320
rect 3895 1317 3925 1320
rect 3895 1314 3931 1317
rect 3861 1306 3877 1308
rect 3635 1294 3650 1298
rect 3553 1292 3650 1294
rect 3678 1292 3846 1304
rect 3862 1294 3877 1298
rect 3895 1295 3934 1314
rect 3953 1308 3960 1309
rect 3959 1301 3960 1308
rect 3943 1298 3944 1301
rect 3959 1298 3972 1301
rect 3895 1294 3925 1295
rect 3934 1294 3940 1295
rect 3943 1294 3972 1298
rect 3862 1293 3972 1294
rect 3862 1292 3978 1293
rect 3537 1284 3588 1292
rect 3537 1272 3562 1284
rect 3569 1272 3588 1284
rect 3619 1284 3669 1292
rect 3619 1276 3635 1284
rect 3642 1282 3669 1284
rect 3678 1282 3899 1292
rect 3642 1272 3899 1282
rect 3928 1284 3978 1292
rect 3928 1275 3944 1284
rect 3537 1264 3588 1272
rect 3635 1264 3899 1272
rect 3925 1272 3944 1275
rect 3951 1272 3978 1284
rect 3925 1264 3978 1272
rect 3553 1256 3554 1264
rect 3569 1256 3582 1264
rect 3553 1248 3569 1256
rect 3550 1241 3569 1244
rect 3550 1232 3572 1241
rect 3523 1222 3572 1232
rect 3523 1216 3553 1222
rect 3572 1217 3577 1222
rect 3495 1200 3569 1216
rect 3587 1208 3617 1264
rect 3652 1254 3860 1264
rect 3895 1260 3940 1264
rect 3943 1263 3944 1264
rect 3959 1263 3972 1264
rect 3678 1224 3867 1254
rect 3693 1221 3867 1224
rect 3686 1218 3867 1221
rect 3495 1198 3508 1200
rect 3523 1198 3557 1200
rect 3495 1182 3569 1198
rect 3596 1194 3609 1208
rect 3624 1194 3640 1210
rect 3686 1205 3697 1218
rect 3479 1160 3480 1176
rect 3495 1160 3508 1182
rect 3523 1160 3553 1182
rect 3596 1178 3658 1194
rect 3686 1187 3697 1203
rect 3702 1198 3712 1218
rect 3722 1198 3736 1218
rect 3739 1205 3748 1218
rect 3764 1205 3773 1218
rect 3702 1187 3736 1198
rect 3739 1187 3748 1203
rect 3764 1187 3773 1203
rect 3780 1198 3790 1218
rect 3800 1198 3814 1218
rect 3815 1205 3826 1218
rect 3780 1187 3814 1198
rect 3815 1187 3826 1203
rect 3872 1194 3888 1210
rect 3895 1208 3925 1260
rect 3959 1256 3960 1263
rect 3944 1248 3960 1256
rect 3931 1216 3944 1235
rect 3959 1216 3989 1232
rect 3931 1200 4005 1216
rect 3931 1198 3944 1200
rect 3959 1198 3993 1200
rect 3596 1176 3609 1178
rect 3624 1176 3658 1178
rect 3596 1160 3658 1176
rect 3702 1171 3718 1174
rect 3780 1171 3810 1182
rect 3858 1178 3904 1194
rect 3931 1182 4005 1198
rect 3858 1176 3892 1178
rect 3857 1160 3904 1176
rect 3931 1160 3944 1182
rect 3959 1160 3989 1182
rect 4016 1160 4017 1176
rect 4032 1160 4045 1320
rect 4075 1216 4088 1320
rect 4133 1298 4134 1308
rect 4149 1298 4162 1308
rect 4133 1294 4162 1298
rect 4167 1294 4197 1320
rect 4215 1306 4231 1308
rect 4303 1306 4356 1320
rect 4304 1304 4368 1306
rect 4411 1304 4426 1320
rect 4475 1317 4505 1320
rect 4475 1314 4511 1317
rect 4441 1306 4457 1308
rect 4215 1294 4230 1298
rect 4133 1292 4230 1294
rect 4258 1292 4426 1304
rect 4442 1294 4457 1298
rect 4475 1295 4514 1314
rect 4533 1308 4540 1309
rect 4539 1301 4540 1308
rect 4523 1298 4524 1301
rect 4539 1298 4552 1301
rect 4475 1294 4505 1295
rect 4514 1294 4520 1295
rect 4523 1294 4552 1298
rect 4442 1293 4552 1294
rect 4442 1292 4558 1293
rect 4117 1284 4168 1292
rect 4117 1272 4142 1284
rect 4149 1272 4168 1284
rect 4199 1284 4249 1292
rect 4199 1276 4215 1284
rect 4222 1282 4249 1284
rect 4258 1282 4479 1292
rect 4222 1272 4479 1282
rect 4508 1284 4558 1292
rect 4508 1275 4524 1284
rect 4117 1264 4168 1272
rect 4215 1264 4479 1272
rect 4505 1272 4524 1275
rect 4531 1272 4558 1284
rect 4505 1264 4558 1272
rect 4133 1256 4134 1264
rect 4149 1256 4162 1264
rect 4133 1248 4149 1256
rect 4130 1241 4149 1244
rect 4130 1232 4152 1241
rect 4103 1222 4152 1232
rect 4103 1216 4133 1222
rect 4152 1217 4157 1222
rect 4075 1200 4149 1216
rect 4167 1208 4197 1264
rect 4232 1254 4440 1264
rect 4475 1260 4520 1264
rect 4523 1263 4524 1264
rect 4539 1263 4552 1264
rect 4258 1224 4447 1254
rect 4273 1221 4447 1224
rect 4266 1218 4447 1221
rect 4075 1198 4088 1200
rect 4103 1198 4137 1200
rect 4075 1182 4149 1198
rect 4176 1194 4189 1208
rect 4204 1194 4220 1210
rect 4266 1205 4277 1218
rect 4059 1160 4060 1176
rect 4075 1160 4088 1182
rect 4103 1160 4133 1182
rect 4176 1178 4238 1194
rect 4266 1187 4277 1203
rect 4282 1198 4292 1218
rect 4302 1198 4316 1218
rect 4319 1205 4328 1218
rect 4344 1205 4353 1218
rect 4282 1187 4316 1198
rect 4319 1187 4328 1203
rect 4344 1187 4353 1203
rect 4360 1198 4370 1218
rect 4380 1198 4394 1218
rect 4395 1205 4406 1218
rect 4360 1187 4394 1198
rect 4395 1187 4406 1203
rect 4452 1194 4468 1210
rect 4475 1208 4505 1260
rect 4539 1256 4540 1263
rect 4524 1248 4540 1256
rect 4511 1216 4524 1235
rect 4539 1216 4569 1232
rect 4511 1200 4585 1216
rect 4511 1198 4524 1200
rect 4539 1198 4573 1200
rect 4176 1176 4189 1178
rect 4204 1176 4238 1178
rect 4176 1160 4238 1176
rect 4282 1171 4298 1174
rect 4360 1171 4390 1182
rect 4438 1178 4484 1194
rect 4511 1182 4585 1198
rect 4438 1176 4472 1178
rect 4437 1160 4484 1176
rect 4511 1160 4524 1182
rect 4539 1160 4569 1182
rect 4596 1160 4597 1176
rect 4612 1160 4625 1320
rect 4655 1216 4668 1320
rect 4713 1298 4714 1308
rect 4729 1298 4742 1308
rect 4713 1294 4742 1298
rect 4747 1294 4777 1320
rect 4795 1306 4811 1308
rect 4883 1306 4936 1320
rect 4884 1304 4948 1306
rect 4991 1304 5006 1320
rect 5055 1317 5085 1320
rect 5055 1314 5091 1317
rect 5021 1306 5037 1308
rect 4795 1294 4810 1298
rect 4713 1292 4810 1294
rect 4838 1292 5006 1304
rect 5022 1294 5037 1298
rect 5055 1295 5094 1314
rect 5113 1308 5120 1309
rect 5119 1301 5120 1308
rect 5103 1298 5104 1301
rect 5119 1298 5132 1301
rect 5055 1294 5085 1295
rect 5094 1294 5100 1295
rect 5103 1294 5132 1298
rect 5022 1293 5132 1294
rect 5022 1292 5138 1293
rect 4697 1284 4748 1292
rect 4697 1272 4722 1284
rect 4729 1272 4748 1284
rect 4779 1284 4829 1292
rect 4779 1276 4795 1284
rect 4802 1282 4829 1284
rect 4838 1282 5059 1292
rect 4802 1272 5059 1282
rect 5088 1284 5138 1292
rect 5088 1275 5104 1284
rect 4697 1264 4748 1272
rect 4795 1264 5059 1272
rect 5085 1272 5104 1275
rect 5111 1272 5138 1284
rect 5085 1264 5138 1272
rect 4713 1256 4714 1264
rect 4729 1256 4742 1264
rect 4713 1248 4729 1256
rect 4710 1241 4729 1244
rect 4710 1232 4732 1241
rect 4683 1222 4732 1232
rect 4683 1216 4713 1222
rect 4732 1217 4737 1222
rect 4655 1200 4729 1216
rect 4747 1208 4777 1264
rect 4812 1254 5020 1264
rect 5055 1260 5100 1264
rect 5103 1263 5104 1264
rect 5119 1263 5132 1264
rect 4838 1224 5027 1254
rect 4853 1221 5027 1224
rect 4846 1218 5027 1221
rect 4655 1198 4668 1200
rect 4683 1198 4717 1200
rect 4655 1182 4729 1198
rect 4756 1194 4769 1208
rect 4784 1194 4800 1210
rect 4846 1205 4857 1218
rect 4639 1160 4640 1176
rect 4655 1160 4668 1182
rect 4683 1160 4713 1182
rect 4756 1178 4818 1194
rect 4846 1187 4857 1203
rect 4862 1198 4872 1218
rect 4882 1198 4896 1218
rect 4899 1205 4908 1218
rect 4924 1205 4933 1218
rect 4862 1187 4896 1198
rect 4899 1187 4908 1203
rect 4924 1187 4933 1203
rect 4940 1198 4950 1218
rect 4960 1198 4974 1218
rect 4975 1205 4986 1218
rect 4940 1187 4974 1198
rect 4975 1187 4986 1203
rect 5032 1194 5048 1210
rect 5055 1208 5085 1260
rect 5119 1256 5120 1263
rect 5104 1248 5120 1256
rect 5091 1216 5104 1235
rect 5119 1216 5149 1232
rect 5091 1200 5165 1216
rect 5091 1198 5104 1200
rect 5119 1198 5153 1200
rect 4756 1176 4769 1178
rect 4784 1176 4818 1178
rect 4756 1160 4818 1176
rect 4862 1171 4878 1174
rect 4940 1171 4970 1182
rect 5018 1178 5064 1194
rect 5091 1182 5165 1198
rect 5018 1176 5052 1178
rect 5017 1160 5064 1176
rect 5091 1160 5104 1182
rect 5119 1160 5149 1182
rect 5176 1160 5177 1176
rect 5192 1160 5205 1320
rect 5235 1216 5248 1320
rect 5293 1298 5294 1308
rect 5309 1298 5322 1308
rect 5293 1294 5322 1298
rect 5327 1294 5357 1320
rect 5375 1306 5391 1308
rect 5463 1306 5516 1320
rect 5464 1304 5528 1306
rect 5571 1304 5586 1320
rect 5635 1317 5665 1320
rect 5635 1314 5671 1317
rect 5601 1306 5617 1308
rect 5375 1294 5390 1298
rect 5293 1292 5390 1294
rect 5418 1292 5586 1304
rect 5602 1294 5617 1298
rect 5635 1295 5674 1314
rect 5693 1308 5700 1309
rect 5699 1301 5700 1308
rect 5683 1298 5684 1301
rect 5699 1298 5712 1301
rect 5635 1294 5665 1295
rect 5674 1294 5680 1295
rect 5683 1294 5712 1298
rect 5602 1293 5712 1294
rect 5602 1292 5718 1293
rect 5277 1284 5328 1292
rect 5277 1272 5302 1284
rect 5309 1272 5328 1284
rect 5359 1284 5409 1292
rect 5359 1276 5375 1284
rect 5382 1282 5409 1284
rect 5418 1282 5639 1292
rect 5382 1272 5639 1282
rect 5668 1284 5718 1292
rect 5668 1275 5684 1284
rect 5277 1264 5328 1272
rect 5375 1264 5639 1272
rect 5665 1272 5684 1275
rect 5691 1272 5718 1284
rect 5665 1264 5718 1272
rect 5293 1256 5294 1264
rect 5309 1256 5322 1264
rect 5293 1248 5309 1256
rect 5290 1241 5309 1244
rect 5290 1232 5312 1241
rect 5263 1222 5312 1232
rect 5263 1216 5293 1222
rect 5312 1217 5317 1222
rect 5235 1200 5309 1216
rect 5327 1208 5357 1264
rect 5392 1254 5600 1264
rect 5635 1260 5680 1264
rect 5683 1263 5684 1264
rect 5699 1263 5712 1264
rect 5418 1224 5607 1254
rect 5433 1221 5607 1224
rect 5426 1218 5607 1221
rect 5235 1198 5248 1200
rect 5263 1198 5297 1200
rect 5235 1182 5309 1198
rect 5336 1194 5349 1208
rect 5364 1194 5380 1210
rect 5426 1205 5437 1218
rect 5219 1160 5220 1176
rect 5235 1160 5248 1182
rect 5263 1160 5293 1182
rect 5336 1178 5398 1194
rect 5426 1187 5437 1203
rect 5442 1198 5452 1218
rect 5462 1198 5476 1218
rect 5479 1205 5488 1218
rect 5504 1205 5513 1218
rect 5442 1187 5476 1198
rect 5479 1187 5488 1203
rect 5504 1187 5513 1203
rect 5520 1198 5530 1218
rect 5540 1198 5554 1218
rect 5555 1205 5566 1218
rect 5520 1187 5554 1198
rect 5555 1187 5566 1203
rect 5612 1194 5628 1210
rect 5635 1208 5665 1260
rect 5699 1256 5700 1263
rect 5684 1248 5700 1256
rect 5671 1216 5684 1235
rect 5699 1216 5729 1232
rect 5671 1200 5745 1216
rect 5671 1198 5684 1200
rect 5699 1198 5733 1200
rect 5336 1176 5349 1178
rect 5364 1176 5398 1178
rect 5336 1160 5398 1176
rect 5442 1171 5458 1174
rect 5520 1171 5550 1182
rect 5598 1178 5644 1194
rect 5671 1182 5745 1198
rect 5598 1176 5632 1178
rect 5597 1160 5644 1176
rect 5671 1160 5684 1182
rect 5699 1160 5729 1182
rect 5756 1160 5757 1176
rect 5772 1160 5785 1320
rect 5815 1216 5828 1320
rect 5873 1298 5874 1308
rect 5889 1298 5902 1308
rect 5873 1294 5902 1298
rect 5907 1294 5937 1320
rect 5955 1306 5971 1308
rect 6043 1306 6096 1320
rect 6044 1304 6108 1306
rect 6151 1304 6166 1320
rect 6215 1317 6245 1320
rect 6215 1314 6251 1317
rect 6181 1306 6197 1308
rect 5955 1294 5970 1298
rect 5873 1292 5970 1294
rect 5998 1292 6166 1304
rect 6182 1294 6197 1298
rect 6215 1295 6254 1314
rect 6273 1308 6280 1309
rect 6279 1301 6280 1308
rect 6263 1298 6264 1301
rect 6279 1298 6292 1301
rect 6215 1294 6245 1295
rect 6254 1294 6260 1295
rect 6263 1294 6292 1298
rect 6182 1293 6292 1294
rect 6182 1292 6298 1293
rect 5857 1284 5908 1292
rect 5857 1272 5882 1284
rect 5889 1272 5908 1284
rect 5939 1284 5989 1292
rect 5939 1276 5955 1284
rect 5962 1282 5989 1284
rect 5998 1282 6219 1292
rect 5962 1272 6219 1282
rect 6248 1284 6298 1292
rect 6248 1275 6264 1284
rect 5857 1264 5908 1272
rect 5955 1264 6219 1272
rect 6245 1272 6264 1275
rect 6271 1272 6298 1284
rect 6245 1264 6298 1272
rect 5873 1256 5874 1264
rect 5889 1256 5902 1264
rect 5873 1248 5889 1256
rect 5870 1241 5889 1244
rect 5870 1232 5892 1241
rect 5843 1222 5892 1232
rect 5843 1216 5873 1222
rect 5892 1217 5897 1222
rect 5815 1200 5889 1216
rect 5907 1208 5937 1264
rect 5972 1254 6180 1264
rect 6215 1260 6260 1264
rect 6263 1263 6264 1264
rect 6279 1263 6292 1264
rect 5998 1224 6187 1254
rect 6013 1221 6187 1224
rect 6006 1218 6187 1221
rect 5815 1198 5828 1200
rect 5843 1198 5877 1200
rect 5815 1182 5889 1198
rect 5916 1194 5929 1208
rect 5944 1194 5960 1210
rect 6006 1205 6017 1218
rect 5799 1160 5800 1176
rect 5815 1160 5828 1182
rect 5843 1160 5873 1182
rect 5916 1178 5978 1194
rect 6006 1187 6017 1203
rect 6022 1198 6032 1218
rect 6042 1198 6056 1218
rect 6059 1205 6068 1218
rect 6084 1205 6093 1218
rect 6022 1187 6056 1198
rect 6059 1187 6068 1203
rect 6084 1187 6093 1203
rect 6100 1198 6110 1218
rect 6120 1198 6134 1218
rect 6135 1205 6146 1218
rect 6100 1187 6134 1198
rect 6135 1187 6146 1203
rect 6192 1194 6208 1210
rect 6215 1208 6245 1260
rect 6279 1256 6280 1263
rect 6264 1248 6280 1256
rect 6251 1216 6264 1235
rect 6279 1216 6309 1232
rect 6251 1200 6325 1216
rect 6251 1198 6264 1200
rect 6279 1198 6313 1200
rect 5916 1176 5929 1178
rect 5944 1176 5978 1178
rect 5916 1160 5978 1176
rect 6022 1171 6038 1174
rect 6100 1171 6130 1182
rect 6178 1178 6224 1194
rect 6251 1182 6325 1198
rect 6178 1176 6212 1178
rect 6177 1160 6224 1176
rect 6251 1160 6264 1182
rect 6279 1160 6309 1182
rect 6336 1160 6337 1176
rect 6352 1160 6365 1320
rect 6395 1216 6408 1320
rect 6453 1298 6454 1308
rect 6469 1298 6482 1308
rect 6453 1294 6482 1298
rect 6487 1294 6517 1320
rect 6535 1306 6551 1308
rect 6623 1306 6676 1320
rect 6624 1304 6688 1306
rect 6731 1304 6746 1320
rect 6795 1317 6825 1320
rect 6795 1314 6831 1317
rect 6761 1306 6777 1308
rect 6535 1294 6550 1298
rect 6453 1292 6550 1294
rect 6578 1292 6746 1304
rect 6762 1294 6777 1298
rect 6795 1295 6834 1314
rect 6853 1308 6860 1309
rect 6859 1301 6860 1308
rect 6843 1298 6844 1301
rect 6859 1298 6872 1301
rect 6795 1294 6825 1295
rect 6834 1294 6840 1295
rect 6843 1294 6872 1298
rect 6762 1293 6872 1294
rect 6762 1292 6878 1293
rect 6437 1284 6488 1292
rect 6437 1272 6462 1284
rect 6469 1272 6488 1284
rect 6519 1284 6569 1292
rect 6519 1276 6535 1284
rect 6542 1282 6569 1284
rect 6578 1282 6799 1292
rect 6542 1272 6799 1282
rect 6828 1284 6878 1292
rect 6828 1275 6844 1284
rect 6437 1264 6488 1272
rect 6535 1264 6799 1272
rect 6825 1272 6844 1275
rect 6851 1272 6878 1284
rect 6825 1264 6878 1272
rect 6453 1256 6454 1264
rect 6469 1256 6482 1264
rect 6453 1248 6469 1256
rect 6450 1241 6469 1244
rect 6450 1232 6472 1241
rect 6423 1222 6472 1232
rect 6423 1216 6453 1222
rect 6472 1217 6477 1222
rect 6395 1200 6469 1216
rect 6487 1208 6517 1264
rect 6552 1254 6760 1264
rect 6795 1260 6840 1264
rect 6843 1263 6844 1264
rect 6859 1263 6872 1264
rect 6578 1224 6767 1254
rect 6593 1221 6767 1224
rect 6586 1218 6767 1221
rect 6395 1198 6408 1200
rect 6423 1198 6457 1200
rect 6395 1182 6469 1198
rect 6496 1194 6509 1208
rect 6524 1194 6540 1210
rect 6586 1205 6597 1218
rect 6379 1160 6380 1176
rect 6395 1160 6408 1182
rect 6423 1160 6453 1182
rect 6496 1178 6558 1194
rect 6586 1187 6597 1203
rect 6602 1198 6612 1218
rect 6622 1198 6636 1218
rect 6639 1205 6648 1218
rect 6664 1205 6673 1218
rect 6602 1187 6636 1198
rect 6639 1187 6648 1203
rect 6664 1187 6673 1203
rect 6680 1198 6690 1218
rect 6700 1198 6714 1218
rect 6715 1205 6726 1218
rect 6680 1187 6714 1198
rect 6715 1187 6726 1203
rect 6772 1194 6788 1210
rect 6795 1208 6825 1260
rect 6859 1256 6860 1263
rect 6844 1248 6860 1256
rect 6831 1216 6844 1235
rect 6859 1216 6889 1232
rect 6831 1200 6905 1216
rect 6831 1198 6844 1200
rect 6859 1198 6893 1200
rect 6496 1176 6509 1178
rect 6524 1176 6558 1178
rect 6496 1160 6558 1176
rect 6602 1171 6618 1174
rect 6680 1171 6710 1182
rect 6758 1178 6804 1194
rect 6831 1182 6905 1198
rect 6758 1176 6792 1178
rect 6757 1160 6804 1176
rect 6831 1160 6844 1182
rect 6859 1160 6889 1182
rect 6916 1160 6917 1176
rect 6932 1160 6945 1320
rect 6975 1216 6988 1320
rect 7033 1298 7034 1308
rect 7049 1298 7062 1308
rect 7033 1294 7062 1298
rect 7067 1294 7097 1320
rect 7115 1306 7131 1308
rect 7203 1306 7256 1320
rect 7204 1304 7268 1306
rect 7311 1304 7326 1320
rect 7375 1317 7405 1320
rect 7375 1314 7411 1317
rect 7341 1306 7357 1308
rect 7115 1294 7130 1298
rect 7033 1292 7130 1294
rect 7158 1292 7326 1304
rect 7342 1294 7357 1298
rect 7375 1295 7414 1314
rect 7433 1308 7440 1309
rect 7439 1301 7440 1308
rect 7423 1298 7424 1301
rect 7439 1298 7452 1301
rect 7375 1294 7405 1295
rect 7414 1294 7420 1295
rect 7423 1294 7452 1298
rect 7342 1293 7452 1294
rect 7342 1292 7458 1293
rect 7017 1284 7068 1292
rect 7017 1272 7042 1284
rect 7049 1272 7068 1284
rect 7099 1284 7149 1292
rect 7099 1276 7115 1284
rect 7122 1282 7149 1284
rect 7158 1282 7379 1292
rect 7122 1272 7379 1282
rect 7408 1284 7458 1292
rect 7408 1275 7424 1284
rect 7017 1264 7068 1272
rect 7115 1264 7379 1272
rect 7405 1272 7424 1275
rect 7431 1272 7458 1284
rect 7405 1264 7458 1272
rect 7033 1256 7034 1264
rect 7049 1256 7062 1264
rect 7033 1248 7049 1256
rect 7030 1241 7049 1244
rect 7030 1232 7052 1241
rect 7003 1222 7052 1232
rect 7003 1216 7033 1222
rect 7052 1217 7057 1222
rect 6975 1200 7049 1216
rect 7067 1208 7097 1264
rect 7132 1254 7340 1264
rect 7375 1260 7420 1264
rect 7423 1263 7424 1264
rect 7439 1263 7452 1264
rect 7158 1224 7347 1254
rect 7173 1221 7347 1224
rect 7166 1218 7347 1221
rect 6975 1198 6988 1200
rect 7003 1198 7037 1200
rect 6975 1182 7049 1198
rect 7076 1194 7089 1208
rect 7104 1194 7120 1210
rect 7166 1205 7177 1218
rect 6959 1160 6960 1176
rect 6975 1160 6988 1182
rect 7003 1160 7033 1182
rect 7076 1178 7138 1194
rect 7166 1187 7177 1203
rect 7182 1198 7192 1218
rect 7202 1198 7216 1218
rect 7219 1205 7228 1218
rect 7244 1205 7253 1218
rect 7182 1187 7216 1198
rect 7219 1187 7228 1203
rect 7244 1187 7253 1203
rect 7260 1198 7270 1218
rect 7280 1198 7294 1218
rect 7295 1205 7306 1218
rect 7260 1187 7294 1198
rect 7295 1187 7306 1203
rect 7352 1194 7368 1210
rect 7375 1208 7405 1260
rect 7439 1256 7440 1263
rect 7424 1248 7440 1256
rect 7411 1216 7424 1235
rect 7439 1216 7469 1232
rect 7411 1200 7485 1216
rect 7411 1198 7424 1200
rect 7439 1198 7473 1200
rect 7076 1176 7089 1178
rect 7104 1176 7138 1178
rect 7076 1160 7138 1176
rect 7182 1171 7198 1174
rect 7260 1171 7290 1182
rect 7338 1178 7384 1194
rect 7411 1182 7485 1198
rect 7338 1176 7372 1178
rect 7337 1160 7384 1176
rect 7411 1160 7424 1182
rect 7439 1160 7469 1182
rect 7496 1160 7497 1176
rect 7512 1160 7525 1320
rect 7555 1216 7568 1320
rect 7613 1298 7614 1308
rect 7629 1298 7642 1308
rect 7613 1294 7642 1298
rect 7647 1294 7677 1320
rect 7695 1306 7711 1308
rect 7783 1306 7836 1320
rect 7784 1304 7848 1306
rect 7891 1304 7906 1320
rect 7955 1317 7985 1320
rect 7955 1314 7991 1317
rect 7921 1306 7937 1308
rect 7695 1294 7710 1298
rect 7613 1292 7710 1294
rect 7738 1292 7906 1304
rect 7922 1294 7937 1298
rect 7955 1295 7994 1314
rect 8013 1308 8020 1309
rect 8019 1301 8020 1308
rect 8003 1298 8004 1301
rect 8019 1298 8032 1301
rect 7955 1294 7985 1295
rect 7994 1294 8000 1295
rect 8003 1294 8032 1298
rect 7922 1293 8032 1294
rect 7922 1292 8038 1293
rect 7597 1284 7648 1292
rect 7597 1272 7622 1284
rect 7629 1272 7648 1284
rect 7679 1284 7729 1292
rect 7679 1276 7695 1284
rect 7702 1282 7729 1284
rect 7738 1282 7959 1292
rect 7702 1272 7959 1282
rect 7988 1284 8038 1292
rect 7988 1275 8004 1284
rect 7597 1264 7648 1272
rect 7695 1264 7959 1272
rect 7985 1272 8004 1275
rect 8011 1272 8038 1284
rect 7985 1264 8038 1272
rect 7613 1256 7614 1264
rect 7629 1256 7642 1264
rect 7613 1248 7629 1256
rect 7610 1241 7629 1244
rect 7610 1232 7632 1241
rect 7583 1222 7632 1232
rect 7583 1216 7613 1222
rect 7632 1217 7637 1222
rect 7555 1200 7629 1216
rect 7647 1208 7677 1264
rect 7712 1254 7920 1264
rect 7955 1260 8000 1264
rect 8003 1263 8004 1264
rect 8019 1263 8032 1264
rect 7738 1224 7927 1254
rect 7753 1221 7927 1224
rect 7746 1218 7927 1221
rect 7555 1198 7568 1200
rect 7583 1198 7617 1200
rect 7555 1182 7629 1198
rect 7656 1194 7669 1208
rect 7684 1194 7700 1210
rect 7746 1205 7757 1218
rect 7539 1160 7540 1176
rect 7555 1160 7568 1182
rect 7583 1160 7613 1182
rect 7656 1178 7718 1194
rect 7746 1187 7757 1203
rect 7762 1198 7772 1218
rect 7782 1198 7796 1218
rect 7799 1205 7808 1218
rect 7824 1205 7833 1218
rect 7762 1187 7796 1198
rect 7799 1187 7808 1203
rect 7824 1187 7833 1203
rect 7840 1198 7850 1218
rect 7860 1198 7874 1218
rect 7875 1205 7886 1218
rect 7840 1187 7874 1198
rect 7875 1187 7886 1203
rect 7932 1194 7948 1210
rect 7955 1208 7985 1260
rect 8019 1256 8020 1263
rect 8004 1248 8020 1256
rect 7991 1216 8004 1235
rect 8019 1216 8049 1232
rect 7991 1200 8065 1216
rect 7991 1198 8004 1200
rect 8019 1198 8053 1200
rect 7656 1176 7669 1178
rect 7684 1176 7718 1178
rect 7656 1160 7718 1176
rect 7762 1171 7778 1174
rect 7840 1171 7870 1182
rect 7918 1178 7964 1194
rect 7991 1182 8065 1198
rect 7918 1176 7952 1178
rect 7917 1160 7964 1176
rect 7991 1160 8004 1182
rect 8019 1160 8049 1182
rect 8076 1160 8077 1176
rect 8092 1160 8105 1320
rect 8135 1216 8148 1320
rect 8193 1298 8194 1308
rect 8209 1298 8222 1308
rect 8193 1294 8222 1298
rect 8227 1294 8257 1320
rect 8275 1306 8291 1308
rect 8363 1306 8416 1320
rect 8364 1304 8428 1306
rect 8471 1304 8486 1320
rect 8535 1317 8565 1320
rect 8535 1314 8571 1317
rect 8501 1306 8517 1308
rect 8275 1294 8290 1298
rect 8193 1292 8290 1294
rect 8318 1292 8486 1304
rect 8502 1294 8517 1298
rect 8535 1295 8574 1314
rect 8593 1308 8600 1309
rect 8599 1301 8600 1308
rect 8583 1298 8584 1301
rect 8599 1298 8612 1301
rect 8535 1294 8565 1295
rect 8574 1294 8580 1295
rect 8583 1294 8612 1298
rect 8502 1293 8612 1294
rect 8502 1292 8618 1293
rect 8177 1284 8228 1292
rect 8177 1272 8202 1284
rect 8209 1272 8228 1284
rect 8259 1284 8309 1292
rect 8259 1276 8275 1284
rect 8282 1282 8309 1284
rect 8318 1282 8539 1292
rect 8282 1272 8539 1282
rect 8568 1284 8618 1292
rect 8568 1275 8584 1284
rect 8177 1264 8228 1272
rect 8275 1264 8539 1272
rect 8565 1272 8584 1275
rect 8591 1272 8618 1284
rect 8565 1264 8618 1272
rect 8193 1256 8194 1264
rect 8209 1256 8222 1264
rect 8193 1248 8209 1256
rect 8190 1241 8209 1244
rect 8190 1232 8212 1241
rect 8163 1222 8212 1232
rect 8163 1216 8193 1222
rect 8212 1217 8217 1222
rect 8135 1200 8209 1216
rect 8227 1208 8257 1264
rect 8292 1254 8500 1264
rect 8535 1260 8580 1264
rect 8583 1263 8584 1264
rect 8599 1263 8612 1264
rect 8318 1224 8507 1254
rect 8333 1221 8507 1224
rect 8326 1218 8507 1221
rect 8135 1198 8148 1200
rect 8163 1198 8197 1200
rect 8135 1182 8209 1198
rect 8236 1194 8249 1208
rect 8264 1194 8280 1210
rect 8326 1205 8337 1218
rect 8119 1160 8120 1176
rect 8135 1160 8148 1182
rect 8163 1160 8193 1182
rect 8236 1178 8298 1194
rect 8326 1187 8337 1203
rect 8342 1198 8352 1218
rect 8362 1198 8376 1218
rect 8379 1205 8388 1218
rect 8404 1205 8413 1218
rect 8342 1187 8376 1198
rect 8379 1187 8388 1203
rect 8404 1187 8413 1203
rect 8420 1198 8430 1218
rect 8440 1198 8454 1218
rect 8455 1205 8466 1218
rect 8420 1187 8454 1198
rect 8455 1187 8466 1203
rect 8512 1194 8528 1210
rect 8535 1208 8565 1260
rect 8599 1256 8600 1263
rect 8584 1248 8600 1256
rect 8571 1216 8584 1235
rect 8599 1216 8629 1232
rect 8571 1200 8645 1216
rect 8571 1198 8584 1200
rect 8599 1198 8633 1200
rect 8236 1176 8249 1178
rect 8264 1176 8298 1178
rect 8236 1160 8298 1176
rect 8342 1171 8358 1174
rect 8420 1171 8450 1182
rect 8498 1178 8544 1194
rect 8571 1182 8645 1198
rect 8498 1176 8532 1178
rect 8497 1160 8544 1176
rect 8571 1160 8584 1182
rect 8599 1160 8629 1182
rect 8656 1160 8657 1176
rect 8672 1160 8685 1320
rect 8715 1216 8728 1320
rect 8773 1298 8774 1308
rect 8789 1298 8802 1308
rect 8773 1294 8802 1298
rect 8807 1294 8837 1320
rect 8855 1306 8871 1308
rect 8943 1306 8996 1320
rect 8944 1304 9008 1306
rect 9051 1304 9066 1320
rect 9115 1317 9145 1320
rect 9115 1314 9151 1317
rect 9081 1306 9097 1308
rect 8855 1294 8870 1298
rect 8773 1292 8870 1294
rect 8898 1292 9066 1304
rect 9082 1294 9097 1298
rect 9115 1295 9154 1314
rect 9173 1308 9180 1309
rect 9179 1301 9180 1308
rect 9163 1298 9164 1301
rect 9179 1298 9192 1301
rect 9115 1294 9145 1295
rect 9154 1294 9160 1295
rect 9163 1294 9192 1298
rect 9082 1293 9192 1294
rect 9082 1292 9198 1293
rect 8757 1284 8808 1292
rect 8757 1272 8782 1284
rect 8789 1272 8808 1284
rect 8839 1284 8889 1292
rect 8839 1276 8855 1284
rect 8862 1282 8889 1284
rect 8898 1282 9119 1292
rect 8862 1272 9119 1282
rect 9148 1284 9198 1292
rect 9148 1275 9164 1284
rect 8757 1264 8808 1272
rect 8855 1264 9119 1272
rect 9145 1272 9164 1275
rect 9171 1272 9198 1284
rect 9145 1264 9198 1272
rect 8773 1256 8774 1264
rect 8789 1256 8802 1264
rect 8773 1248 8789 1256
rect 8770 1241 8789 1244
rect 8770 1232 8792 1241
rect 8743 1222 8792 1232
rect 8743 1216 8773 1222
rect 8792 1217 8797 1222
rect 8715 1200 8789 1216
rect 8807 1208 8837 1264
rect 8872 1254 9080 1264
rect 9115 1260 9160 1264
rect 9163 1263 9164 1264
rect 9179 1263 9192 1264
rect 8898 1224 9087 1254
rect 8913 1221 9087 1224
rect 8906 1218 9087 1221
rect 8715 1198 8728 1200
rect 8743 1198 8777 1200
rect 8715 1182 8789 1198
rect 8816 1194 8829 1208
rect 8844 1194 8860 1210
rect 8906 1205 8917 1218
rect 8699 1160 8700 1176
rect 8715 1160 8728 1182
rect 8743 1160 8773 1182
rect 8816 1178 8878 1194
rect 8906 1187 8917 1203
rect 8922 1198 8932 1218
rect 8942 1198 8956 1218
rect 8959 1205 8968 1218
rect 8984 1205 8993 1218
rect 8922 1187 8956 1198
rect 8959 1187 8968 1203
rect 8984 1187 8993 1203
rect 9000 1198 9010 1218
rect 9020 1198 9034 1218
rect 9035 1205 9046 1218
rect 9000 1187 9034 1198
rect 9035 1187 9046 1203
rect 9092 1194 9108 1210
rect 9115 1208 9145 1260
rect 9179 1256 9180 1263
rect 9164 1248 9180 1256
rect 9151 1216 9164 1235
rect 9179 1216 9209 1232
rect 9151 1200 9225 1216
rect 9151 1198 9164 1200
rect 9179 1198 9213 1200
rect 8816 1176 8829 1178
rect 8844 1176 8878 1178
rect 8816 1160 8878 1176
rect 8922 1171 8938 1174
rect 9000 1171 9030 1182
rect 9078 1178 9124 1194
rect 9151 1182 9225 1198
rect 9078 1176 9112 1178
rect 9077 1160 9124 1176
rect 9151 1160 9164 1182
rect 9179 1160 9209 1182
rect 9236 1160 9237 1176
rect 9252 1160 9265 1320
rect -7 1152 34 1160
rect -7 1126 8 1152
rect 15 1126 34 1152
rect 98 1148 160 1160
rect 172 1148 247 1160
rect 305 1148 380 1160
rect 392 1148 423 1160
rect 429 1148 464 1160
rect 98 1146 260 1148
rect -7 1118 34 1126
rect 116 1122 129 1146
rect 144 1144 159 1146
rect -1 1108 0 1118
rect 15 1108 28 1118
rect 43 1108 73 1122
rect 116 1108 159 1122
rect 183 1119 190 1126
rect 193 1122 260 1146
rect 292 1146 464 1148
rect 262 1124 290 1128
rect 292 1124 372 1146
rect 393 1144 408 1146
rect 262 1122 372 1124
rect 193 1118 372 1122
rect 166 1108 196 1118
rect 198 1108 351 1118
rect 359 1108 389 1118
rect 393 1108 423 1122
rect 451 1108 464 1146
rect 536 1152 571 1160
rect 536 1126 537 1152
rect 544 1126 571 1152
rect 479 1108 509 1122
rect 536 1118 571 1126
rect 573 1152 614 1160
rect 573 1126 588 1152
rect 595 1126 614 1152
rect 678 1148 740 1160
rect 752 1148 827 1160
rect 885 1148 960 1160
rect 972 1148 1003 1160
rect 1009 1148 1044 1160
rect 678 1146 840 1148
rect 573 1118 614 1126
rect 696 1122 709 1146
rect 724 1144 739 1146
rect 536 1108 537 1118
rect 552 1108 565 1118
rect 579 1108 580 1118
rect 595 1108 608 1118
rect 623 1108 653 1122
rect 696 1108 739 1122
rect 763 1119 770 1126
rect 773 1122 840 1146
rect 872 1146 1044 1148
rect 842 1124 870 1128
rect 872 1124 952 1146
rect 973 1144 988 1146
rect 842 1122 952 1124
rect 773 1118 952 1122
rect 746 1108 776 1118
rect 778 1108 931 1118
rect 939 1108 969 1118
rect 973 1108 1003 1122
rect 1031 1108 1044 1146
rect 1116 1152 1151 1160
rect 1116 1126 1117 1152
rect 1124 1126 1151 1152
rect 1059 1108 1089 1122
rect 1116 1118 1151 1126
rect 1153 1152 1194 1160
rect 1153 1126 1168 1152
rect 1175 1126 1194 1152
rect 1258 1148 1320 1160
rect 1332 1148 1407 1160
rect 1465 1148 1540 1160
rect 1552 1148 1583 1160
rect 1589 1148 1624 1160
rect 1258 1146 1420 1148
rect 1153 1118 1194 1126
rect 1276 1122 1289 1146
rect 1304 1144 1319 1146
rect 1116 1108 1117 1118
rect 1132 1108 1145 1118
rect 1159 1108 1160 1118
rect 1175 1108 1188 1118
rect 1203 1108 1233 1122
rect 1276 1108 1319 1122
rect 1343 1119 1350 1126
rect 1353 1122 1420 1146
rect 1452 1146 1624 1148
rect 1422 1124 1450 1128
rect 1452 1124 1532 1146
rect 1553 1144 1568 1146
rect 1422 1122 1532 1124
rect 1353 1118 1532 1122
rect 1326 1108 1356 1118
rect 1358 1108 1511 1118
rect 1519 1108 1549 1118
rect 1553 1108 1583 1122
rect 1611 1108 1624 1146
rect 1696 1152 1731 1160
rect 1696 1126 1697 1152
rect 1704 1126 1731 1152
rect 1639 1108 1669 1122
rect 1696 1118 1731 1126
rect 1733 1152 1774 1160
rect 1733 1126 1748 1152
rect 1755 1126 1774 1152
rect 1838 1148 1900 1160
rect 1912 1148 1987 1160
rect 2045 1148 2120 1160
rect 2132 1148 2163 1160
rect 2169 1148 2204 1160
rect 1838 1146 2000 1148
rect 1733 1118 1774 1126
rect 1856 1122 1869 1146
rect 1884 1144 1899 1146
rect 1696 1108 1697 1118
rect 1712 1108 1725 1118
rect 1739 1108 1740 1118
rect 1755 1108 1768 1118
rect 1783 1108 1813 1122
rect 1856 1108 1899 1122
rect 1923 1119 1930 1126
rect 1933 1122 2000 1146
rect 2032 1146 2204 1148
rect 2002 1124 2030 1128
rect 2032 1124 2112 1146
rect 2133 1144 2148 1146
rect 2002 1122 2112 1124
rect 1933 1118 2112 1122
rect 1906 1108 1936 1118
rect 1938 1108 2091 1118
rect 2099 1108 2129 1118
rect 2133 1108 2163 1122
rect 2191 1108 2204 1146
rect 2276 1152 2311 1160
rect 2276 1126 2277 1152
rect 2284 1126 2311 1152
rect 2219 1108 2249 1122
rect 2276 1118 2311 1126
rect 2313 1152 2354 1160
rect 2313 1126 2328 1152
rect 2335 1126 2354 1152
rect 2418 1148 2480 1160
rect 2492 1148 2567 1160
rect 2625 1148 2700 1160
rect 2712 1148 2743 1160
rect 2749 1148 2784 1160
rect 2418 1146 2580 1148
rect 2313 1118 2354 1126
rect 2436 1122 2449 1146
rect 2464 1144 2479 1146
rect 2276 1108 2277 1118
rect 2292 1108 2305 1118
rect 2319 1108 2320 1118
rect 2335 1108 2348 1118
rect 2363 1108 2393 1122
rect 2436 1108 2479 1122
rect 2503 1119 2510 1126
rect 2513 1122 2580 1146
rect 2612 1146 2784 1148
rect 2582 1124 2610 1128
rect 2612 1124 2692 1146
rect 2713 1144 2728 1146
rect 2582 1122 2692 1124
rect 2513 1118 2692 1122
rect 2486 1108 2516 1118
rect 2518 1108 2671 1118
rect 2679 1108 2709 1118
rect 2713 1108 2743 1122
rect 2771 1108 2784 1146
rect 2856 1152 2891 1160
rect 2856 1126 2857 1152
rect 2864 1126 2891 1152
rect 2799 1108 2829 1122
rect 2856 1118 2891 1126
rect 2893 1152 2934 1160
rect 2893 1126 2908 1152
rect 2915 1126 2934 1152
rect 2998 1148 3060 1160
rect 3072 1148 3147 1160
rect 3205 1148 3280 1160
rect 3292 1148 3323 1160
rect 3329 1148 3364 1160
rect 2998 1146 3160 1148
rect 2893 1118 2934 1126
rect 3016 1122 3029 1146
rect 3044 1144 3059 1146
rect 2856 1108 2857 1118
rect 2872 1108 2885 1118
rect 2899 1108 2900 1118
rect 2915 1108 2928 1118
rect 2943 1108 2973 1122
rect 3016 1108 3059 1122
rect 3083 1119 3090 1126
rect 3093 1122 3160 1146
rect 3192 1146 3364 1148
rect 3162 1124 3190 1128
rect 3192 1124 3272 1146
rect 3293 1144 3308 1146
rect 3162 1122 3272 1124
rect 3093 1118 3272 1122
rect 3066 1108 3096 1118
rect 3098 1108 3251 1118
rect 3259 1108 3289 1118
rect 3293 1108 3323 1122
rect 3351 1108 3364 1146
rect 3436 1152 3471 1160
rect 3436 1126 3437 1152
rect 3444 1126 3471 1152
rect 3379 1108 3409 1122
rect 3436 1118 3471 1126
rect 3473 1152 3514 1160
rect 3473 1126 3488 1152
rect 3495 1126 3514 1152
rect 3578 1148 3640 1160
rect 3652 1148 3727 1160
rect 3785 1148 3860 1160
rect 3872 1148 3903 1160
rect 3909 1148 3944 1160
rect 3578 1146 3740 1148
rect 3473 1118 3514 1126
rect 3596 1122 3609 1146
rect 3624 1144 3639 1146
rect 3436 1108 3437 1118
rect 3452 1108 3465 1118
rect 3479 1108 3480 1118
rect 3495 1108 3508 1118
rect 3523 1108 3553 1122
rect 3596 1108 3639 1122
rect 3663 1119 3670 1126
rect 3673 1122 3740 1146
rect 3772 1146 3944 1148
rect 3742 1124 3770 1128
rect 3772 1124 3852 1146
rect 3873 1144 3888 1146
rect 3742 1122 3852 1124
rect 3673 1118 3852 1122
rect 3646 1108 3676 1118
rect 3678 1108 3831 1118
rect 3839 1108 3869 1118
rect 3873 1108 3903 1122
rect 3931 1108 3944 1146
rect 4016 1152 4051 1160
rect 4016 1126 4017 1152
rect 4024 1126 4051 1152
rect 3959 1108 3989 1122
rect 4016 1118 4051 1126
rect 4053 1152 4094 1160
rect 4053 1126 4068 1152
rect 4075 1126 4094 1152
rect 4158 1148 4220 1160
rect 4232 1148 4307 1160
rect 4365 1148 4440 1160
rect 4452 1148 4483 1160
rect 4489 1148 4524 1160
rect 4158 1146 4320 1148
rect 4053 1118 4094 1126
rect 4176 1122 4189 1146
rect 4204 1144 4219 1146
rect 4016 1108 4017 1118
rect 4032 1108 4045 1118
rect 4059 1108 4060 1118
rect 4075 1108 4088 1118
rect 4103 1108 4133 1122
rect 4176 1108 4219 1122
rect 4243 1119 4250 1126
rect 4253 1122 4320 1146
rect 4352 1146 4524 1148
rect 4322 1124 4350 1128
rect 4352 1124 4432 1146
rect 4453 1144 4468 1146
rect 4322 1122 4432 1124
rect 4253 1118 4432 1122
rect 4226 1108 4256 1118
rect 4258 1108 4411 1118
rect 4419 1108 4449 1118
rect 4453 1108 4483 1122
rect 4511 1108 4524 1146
rect 4596 1152 4631 1160
rect 4596 1126 4597 1152
rect 4604 1126 4631 1152
rect 4539 1108 4569 1122
rect 4596 1118 4631 1126
rect 4633 1152 4674 1160
rect 4633 1126 4648 1152
rect 4655 1126 4674 1152
rect 4738 1148 4800 1160
rect 4812 1148 4887 1160
rect 4945 1148 5020 1160
rect 5032 1148 5063 1160
rect 5069 1148 5104 1160
rect 4738 1146 4900 1148
rect 4633 1118 4674 1126
rect 4756 1122 4769 1146
rect 4784 1144 4799 1146
rect 4596 1108 4597 1118
rect 4612 1108 4625 1118
rect 4639 1108 4640 1118
rect 4655 1108 4668 1118
rect 4683 1108 4713 1122
rect 4756 1108 4799 1122
rect 4823 1119 4830 1126
rect 4833 1122 4900 1146
rect 4932 1146 5104 1148
rect 4902 1124 4930 1128
rect 4932 1124 5012 1146
rect 5033 1144 5048 1146
rect 4902 1122 5012 1124
rect 4833 1118 5012 1122
rect 4806 1108 4836 1118
rect 4838 1108 4991 1118
rect 4999 1108 5029 1118
rect 5033 1108 5063 1122
rect 5091 1108 5104 1146
rect 5176 1152 5211 1160
rect 5176 1126 5177 1152
rect 5184 1126 5211 1152
rect 5119 1108 5149 1122
rect 5176 1118 5211 1126
rect 5213 1152 5254 1160
rect 5213 1126 5228 1152
rect 5235 1126 5254 1152
rect 5318 1148 5380 1160
rect 5392 1148 5467 1160
rect 5525 1148 5600 1160
rect 5612 1148 5643 1160
rect 5649 1148 5684 1160
rect 5318 1146 5480 1148
rect 5213 1118 5254 1126
rect 5336 1122 5349 1146
rect 5364 1144 5379 1146
rect 5176 1108 5177 1118
rect 5192 1108 5205 1118
rect 5219 1108 5220 1118
rect 5235 1108 5248 1118
rect 5263 1108 5293 1122
rect 5336 1108 5379 1122
rect 5403 1119 5410 1126
rect 5413 1122 5480 1146
rect 5512 1146 5684 1148
rect 5482 1124 5510 1128
rect 5512 1124 5592 1146
rect 5613 1144 5628 1146
rect 5482 1122 5592 1124
rect 5413 1118 5592 1122
rect 5386 1108 5416 1118
rect 5418 1108 5571 1118
rect 5579 1108 5609 1118
rect 5613 1108 5643 1122
rect 5671 1108 5684 1146
rect 5756 1152 5791 1160
rect 5756 1126 5757 1152
rect 5764 1126 5791 1152
rect 5699 1108 5729 1122
rect 5756 1118 5791 1126
rect 5793 1152 5834 1160
rect 5793 1126 5808 1152
rect 5815 1126 5834 1152
rect 5898 1148 5960 1160
rect 5972 1148 6047 1160
rect 6105 1148 6180 1160
rect 6192 1148 6223 1160
rect 6229 1148 6264 1160
rect 5898 1146 6060 1148
rect 5793 1118 5834 1126
rect 5916 1122 5929 1146
rect 5944 1144 5959 1146
rect 5756 1108 5757 1118
rect 5772 1108 5785 1118
rect 5799 1108 5800 1118
rect 5815 1108 5828 1118
rect 5843 1108 5873 1122
rect 5916 1108 5959 1122
rect 5983 1119 5990 1126
rect 5993 1122 6060 1146
rect 6092 1146 6264 1148
rect 6062 1124 6090 1128
rect 6092 1124 6172 1146
rect 6193 1144 6208 1146
rect 6062 1122 6172 1124
rect 5993 1118 6172 1122
rect 5966 1108 5996 1118
rect 5998 1108 6151 1118
rect 6159 1108 6189 1118
rect 6193 1108 6223 1122
rect 6251 1108 6264 1146
rect 6336 1152 6371 1160
rect 6336 1126 6337 1152
rect 6344 1126 6371 1152
rect 6279 1108 6309 1122
rect 6336 1118 6371 1126
rect 6373 1152 6414 1160
rect 6373 1126 6388 1152
rect 6395 1126 6414 1152
rect 6478 1148 6540 1160
rect 6552 1148 6627 1160
rect 6685 1148 6760 1160
rect 6772 1148 6803 1160
rect 6809 1148 6844 1160
rect 6478 1146 6640 1148
rect 6373 1118 6414 1126
rect 6496 1122 6509 1146
rect 6524 1144 6539 1146
rect 6336 1108 6337 1118
rect 6352 1108 6365 1118
rect 6379 1108 6380 1118
rect 6395 1108 6408 1118
rect 6423 1108 6453 1122
rect 6496 1108 6539 1122
rect 6563 1119 6570 1126
rect 6573 1122 6640 1146
rect 6672 1146 6844 1148
rect 6642 1124 6670 1128
rect 6672 1124 6752 1146
rect 6773 1144 6788 1146
rect 6642 1122 6752 1124
rect 6573 1118 6752 1122
rect 6546 1108 6576 1118
rect 6578 1108 6731 1118
rect 6739 1108 6769 1118
rect 6773 1108 6803 1122
rect 6831 1108 6844 1146
rect 6916 1152 6951 1160
rect 6916 1126 6917 1152
rect 6924 1126 6951 1152
rect 6859 1108 6889 1122
rect 6916 1118 6951 1126
rect 6953 1152 6994 1160
rect 6953 1126 6968 1152
rect 6975 1126 6994 1152
rect 7058 1148 7120 1160
rect 7132 1148 7207 1160
rect 7265 1148 7340 1160
rect 7352 1148 7383 1160
rect 7389 1148 7424 1160
rect 7058 1146 7220 1148
rect 6953 1118 6994 1126
rect 7076 1122 7089 1146
rect 7104 1144 7119 1146
rect 6916 1108 6917 1118
rect 6932 1108 6945 1118
rect 6959 1108 6960 1118
rect 6975 1108 6988 1118
rect 7003 1108 7033 1122
rect 7076 1108 7119 1122
rect 7143 1119 7150 1126
rect 7153 1122 7220 1146
rect 7252 1146 7424 1148
rect 7222 1124 7250 1128
rect 7252 1124 7332 1146
rect 7353 1144 7368 1146
rect 7222 1122 7332 1124
rect 7153 1118 7332 1122
rect 7126 1108 7156 1118
rect 7158 1108 7311 1118
rect 7319 1108 7349 1118
rect 7353 1108 7383 1122
rect 7411 1108 7424 1146
rect 7496 1152 7531 1160
rect 7496 1126 7497 1152
rect 7504 1126 7531 1152
rect 7439 1108 7469 1122
rect 7496 1118 7531 1126
rect 7533 1152 7574 1160
rect 7533 1126 7548 1152
rect 7555 1126 7574 1152
rect 7638 1148 7700 1160
rect 7712 1148 7787 1160
rect 7845 1148 7920 1160
rect 7932 1148 7963 1160
rect 7969 1148 8004 1160
rect 7638 1146 7800 1148
rect 7533 1118 7574 1126
rect 7656 1122 7669 1146
rect 7684 1144 7699 1146
rect 7496 1108 7497 1118
rect 7512 1108 7525 1118
rect 7539 1108 7540 1118
rect 7555 1108 7568 1118
rect 7583 1108 7613 1122
rect 7656 1108 7699 1122
rect 7723 1119 7730 1126
rect 7733 1122 7800 1146
rect 7832 1146 8004 1148
rect 7802 1124 7830 1128
rect 7832 1124 7912 1146
rect 7933 1144 7948 1146
rect 7802 1122 7912 1124
rect 7733 1118 7912 1122
rect 7706 1108 7736 1118
rect 7738 1108 7891 1118
rect 7899 1108 7929 1118
rect 7933 1108 7963 1122
rect 7991 1108 8004 1146
rect 8076 1152 8111 1160
rect 8076 1126 8077 1152
rect 8084 1126 8111 1152
rect 8019 1108 8049 1122
rect 8076 1118 8111 1126
rect 8113 1152 8154 1160
rect 8113 1126 8128 1152
rect 8135 1126 8154 1152
rect 8218 1148 8280 1160
rect 8292 1148 8367 1160
rect 8425 1148 8500 1160
rect 8512 1148 8543 1160
rect 8549 1148 8584 1160
rect 8218 1146 8380 1148
rect 8113 1118 8154 1126
rect 8236 1122 8249 1146
rect 8264 1144 8279 1146
rect 8076 1108 8077 1118
rect 8092 1108 8105 1118
rect 8119 1108 8120 1118
rect 8135 1108 8148 1118
rect 8163 1108 8193 1122
rect 8236 1108 8279 1122
rect 8303 1119 8310 1126
rect 8313 1122 8380 1146
rect 8412 1146 8584 1148
rect 8382 1124 8410 1128
rect 8412 1124 8492 1146
rect 8513 1144 8528 1146
rect 8382 1122 8492 1124
rect 8313 1118 8492 1122
rect 8286 1108 8316 1118
rect 8318 1108 8471 1118
rect 8479 1108 8509 1118
rect 8513 1108 8543 1122
rect 8571 1108 8584 1146
rect 8656 1152 8691 1160
rect 8656 1126 8657 1152
rect 8664 1126 8691 1152
rect 8599 1108 8629 1122
rect 8656 1118 8691 1126
rect 8693 1152 8734 1160
rect 8693 1126 8708 1152
rect 8715 1126 8734 1152
rect 8798 1148 8860 1160
rect 8872 1148 8947 1160
rect 9005 1148 9080 1160
rect 9092 1148 9123 1160
rect 9129 1148 9164 1160
rect 8798 1146 8960 1148
rect 8693 1118 8734 1126
rect 8816 1122 8829 1146
rect 8844 1144 8859 1146
rect 8656 1108 8657 1118
rect 8672 1108 8685 1118
rect 8699 1108 8700 1118
rect 8715 1108 8728 1118
rect 8743 1108 8773 1122
rect 8816 1108 8859 1122
rect 8883 1119 8890 1126
rect 8893 1122 8960 1146
rect 8992 1146 9164 1148
rect 8962 1124 8990 1128
rect 8992 1124 9072 1146
rect 9093 1144 9108 1146
rect 8962 1122 9072 1124
rect 8893 1118 9072 1122
rect 8866 1108 8896 1118
rect 8898 1108 9051 1118
rect 9059 1108 9089 1118
rect 9093 1108 9123 1122
rect 9151 1108 9164 1146
rect 9236 1152 9271 1160
rect 9236 1126 9237 1152
rect 9244 1126 9271 1152
rect 9179 1108 9209 1122
rect 9236 1118 9271 1126
rect 9236 1108 9237 1118
rect 9252 1108 9265 1118
rect -1 1102 9265 1108
rect 0 1094 9265 1102
rect 15 1064 28 1094
rect 43 1076 73 1094
rect 116 1080 130 1094
rect 166 1080 386 1094
rect 117 1078 130 1080
rect 83 1066 98 1078
rect 80 1064 102 1066
rect 107 1064 137 1078
rect 198 1076 351 1080
rect 180 1064 372 1076
rect 415 1064 445 1078
rect 451 1064 464 1094
rect 479 1076 509 1094
rect 552 1064 565 1094
rect 595 1064 608 1094
rect 623 1076 653 1094
rect 696 1080 710 1094
rect 746 1080 966 1094
rect 697 1078 710 1080
rect 663 1066 678 1078
rect 660 1064 682 1066
rect 687 1064 717 1078
rect 778 1076 931 1080
rect 760 1064 952 1076
rect 995 1064 1025 1078
rect 1031 1064 1044 1094
rect 1059 1076 1089 1094
rect 1132 1064 1145 1094
rect 1175 1064 1188 1094
rect 1203 1076 1233 1094
rect 1276 1080 1290 1094
rect 1326 1080 1546 1094
rect 1277 1078 1290 1080
rect 1243 1066 1258 1078
rect 1240 1064 1262 1066
rect 1267 1064 1297 1078
rect 1358 1076 1511 1080
rect 1340 1064 1532 1076
rect 1575 1064 1605 1078
rect 1611 1064 1624 1094
rect 1639 1076 1669 1094
rect 1712 1064 1725 1094
rect 1755 1064 1768 1094
rect 1783 1076 1813 1094
rect 1856 1080 1870 1094
rect 1906 1080 2126 1094
rect 1857 1078 1870 1080
rect 1823 1066 1838 1078
rect 1820 1064 1842 1066
rect 1847 1064 1877 1078
rect 1938 1076 2091 1080
rect 1920 1064 2112 1076
rect 2155 1064 2185 1078
rect 2191 1064 2204 1094
rect 2219 1076 2249 1094
rect 2292 1064 2305 1094
rect 2335 1064 2348 1094
rect 2363 1076 2393 1094
rect 2436 1080 2450 1094
rect 2486 1080 2706 1094
rect 2437 1078 2450 1080
rect 2403 1066 2418 1078
rect 2400 1064 2422 1066
rect 2427 1064 2457 1078
rect 2518 1076 2671 1080
rect 2500 1064 2692 1076
rect 2735 1064 2765 1078
rect 2771 1064 2784 1094
rect 2799 1076 2829 1094
rect 2872 1064 2885 1094
rect 2915 1064 2928 1094
rect 2943 1076 2973 1094
rect 3016 1080 3030 1094
rect 3066 1080 3286 1094
rect 3017 1078 3030 1080
rect 2983 1066 2998 1078
rect 2980 1064 3002 1066
rect 3007 1064 3037 1078
rect 3098 1076 3251 1080
rect 3080 1064 3272 1076
rect 3315 1064 3345 1078
rect 3351 1064 3364 1094
rect 3379 1076 3409 1094
rect 3452 1064 3465 1094
rect 3495 1064 3508 1094
rect 3523 1076 3553 1094
rect 3596 1080 3610 1094
rect 3646 1080 3866 1094
rect 3597 1078 3610 1080
rect 3563 1066 3578 1078
rect 3560 1064 3582 1066
rect 3587 1064 3617 1078
rect 3678 1076 3831 1080
rect 3660 1064 3852 1076
rect 3895 1064 3925 1078
rect 3931 1064 3944 1094
rect 3959 1076 3989 1094
rect 4032 1064 4045 1094
rect 4075 1064 4088 1094
rect 4103 1076 4133 1094
rect 4176 1080 4190 1094
rect 4226 1080 4446 1094
rect 4177 1078 4190 1080
rect 4143 1066 4158 1078
rect 4140 1064 4162 1066
rect 4167 1064 4197 1078
rect 4258 1076 4411 1080
rect 4240 1064 4432 1076
rect 4475 1064 4505 1078
rect 4511 1064 4524 1094
rect 4539 1076 4569 1094
rect 4612 1064 4625 1094
rect 4655 1064 4668 1094
rect 4683 1076 4713 1094
rect 4756 1080 4770 1094
rect 4806 1080 5026 1094
rect 4757 1078 4770 1080
rect 4723 1066 4738 1078
rect 4720 1064 4742 1066
rect 4747 1064 4777 1078
rect 4838 1076 4991 1080
rect 4820 1064 5012 1076
rect 5055 1064 5085 1078
rect 5091 1064 5104 1094
rect 5119 1076 5149 1094
rect 5192 1064 5205 1094
rect 5235 1064 5248 1094
rect 5263 1076 5293 1094
rect 5336 1080 5350 1094
rect 5386 1080 5606 1094
rect 5337 1078 5350 1080
rect 5303 1066 5318 1078
rect 5300 1064 5322 1066
rect 5327 1064 5357 1078
rect 5418 1076 5571 1080
rect 5400 1064 5592 1076
rect 5635 1064 5665 1078
rect 5671 1064 5684 1094
rect 5699 1076 5729 1094
rect 5772 1064 5785 1094
rect 5815 1064 5828 1094
rect 5843 1076 5873 1094
rect 5916 1080 5930 1094
rect 5966 1080 6186 1094
rect 5917 1078 5930 1080
rect 5883 1066 5898 1078
rect 5880 1064 5902 1066
rect 5907 1064 5937 1078
rect 5998 1076 6151 1080
rect 5980 1064 6172 1076
rect 6215 1064 6245 1078
rect 6251 1064 6264 1094
rect 6279 1076 6309 1094
rect 6352 1064 6365 1094
rect 6395 1064 6408 1094
rect 6423 1076 6453 1094
rect 6496 1080 6510 1094
rect 6546 1080 6766 1094
rect 6497 1078 6510 1080
rect 6463 1066 6478 1078
rect 6460 1064 6482 1066
rect 6487 1064 6517 1078
rect 6578 1076 6731 1080
rect 6560 1064 6752 1076
rect 6795 1064 6825 1078
rect 6831 1064 6844 1094
rect 6859 1076 6889 1094
rect 6932 1064 6945 1094
rect 6975 1064 6988 1094
rect 7003 1076 7033 1094
rect 7076 1080 7090 1094
rect 7126 1080 7346 1094
rect 7077 1078 7090 1080
rect 7043 1066 7058 1078
rect 7040 1064 7062 1066
rect 7067 1064 7097 1078
rect 7158 1076 7311 1080
rect 7140 1064 7332 1076
rect 7375 1064 7405 1078
rect 7411 1064 7424 1094
rect 7439 1076 7469 1094
rect 7512 1064 7525 1094
rect 7555 1064 7568 1094
rect 7583 1076 7613 1094
rect 7656 1080 7670 1094
rect 7706 1080 7926 1094
rect 7657 1078 7670 1080
rect 7623 1066 7638 1078
rect 7620 1064 7642 1066
rect 7647 1064 7677 1078
rect 7738 1076 7891 1080
rect 7720 1064 7912 1076
rect 7955 1064 7985 1078
rect 7991 1064 8004 1094
rect 8019 1076 8049 1094
rect 8092 1064 8105 1094
rect 8135 1064 8148 1094
rect 8163 1076 8193 1094
rect 8236 1080 8250 1094
rect 8286 1080 8506 1094
rect 8237 1078 8250 1080
rect 8203 1066 8218 1078
rect 8200 1064 8222 1066
rect 8227 1064 8257 1078
rect 8318 1076 8471 1080
rect 8300 1064 8492 1076
rect 8535 1064 8565 1078
rect 8571 1064 8584 1094
rect 8599 1076 8629 1094
rect 8672 1064 8685 1094
rect 8715 1064 8728 1094
rect 8743 1076 8773 1094
rect 8816 1080 8830 1094
rect 8866 1080 9086 1094
rect 8817 1078 8830 1080
rect 8783 1066 8798 1078
rect 8780 1064 8802 1066
rect 8807 1064 8837 1078
rect 8898 1076 9051 1080
rect 8880 1064 9072 1076
rect 9115 1064 9145 1078
rect 9151 1064 9164 1094
rect 9179 1076 9209 1094
rect 9252 1064 9265 1094
rect 0 1050 9265 1064
rect 15 946 28 1050
rect 73 1028 74 1038
rect 89 1028 102 1038
rect 73 1024 102 1028
rect 107 1024 137 1050
rect 155 1036 171 1038
rect 243 1036 296 1050
rect 244 1034 308 1036
rect 351 1034 366 1050
rect 415 1047 445 1050
rect 415 1044 451 1047
rect 381 1036 397 1038
rect 155 1024 170 1028
rect 73 1022 170 1024
rect 198 1022 366 1034
rect 382 1024 397 1028
rect 415 1025 454 1044
rect 473 1038 480 1039
rect 479 1031 480 1038
rect 463 1028 464 1031
rect 479 1028 492 1031
rect 415 1024 445 1025
rect 454 1024 460 1025
rect 463 1024 492 1028
rect 382 1023 492 1024
rect 382 1022 498 1023
rect 57 1014 108 1022
rect 57 1002 82 1014
rect 89 1002 108 1014
rect 139 1014 189 1022
rect 139 1006 155 1014
rect 162 1012 189 1014
rect 198 1012 419 1022
rect 162 1002 419 1012
rect 448 1014 498 1022
rect 448 1005 464 1014
rect 57 994 108 1002
rect 155 994 419 1002
rect 445 1002 464 1005
rect 471 1002 498 1014
rect 445 994 498 1002
rect 73 986 74 994
rect 89 986 102 994
rect 73 978 89 986
rect 70 971 89 974
rect 70 962 92 971
rect 43 952 92 962
rect 43 946 73 952
rect 92 947 97 952
rect 15 930 89 946
rect 107 938 137 994
rect 172 984 380 994
rect 415 990 460 994
rect 463 993 464 994
rect 479 993 492 994
rect 198 954 387 984
rect 213 951 387 954
rect 206 948 387 951
rect 15 928 28 930
rect 43 928 77 930
rect 15 912 89 928
rect 116 924 129 938
rect 144 924 160 940
rect 206 935 217 948
rect -1 890 0 906
rect 15 890 28 912
rect 43 890 73 912
rect 116 908 178 924
rect 206 917 217 933
rect 222 928 232 948
rect 242 928 256 948
rect 259 935 268 948
rect 284 935 293 948
rect 222 917 256 928
rect 259 917 268 933
rect 284 917 293 933
rect 300 928 310 948
rect 320 928 334 948
rect 335 935 346 948
rect 300 917 334 928
rect 335 917 346 933
rect 392 924 408 940
rect 415 938 445 990
rect 479 986 480 993
rect 464 978 480 986
rect 451 946 464 965
rect 479 946 509 962
rect 451 930 525 946
rect 451 928 464 930
rect 479 928 513 930
rect 116 906 129 908
rect 144 906 178 908
rect 116 890 178 906
rect 222 901 238 904
rect 300 901 330 912
rect 378 908 424 924
rect 451 912 525 928
rect 378 906 412 908
rect 377 890 424 906
rect 451 890 464 912
rect 479 890 509 912
rect 536 890 537 906
rect 552 890 565 1050
rect 595 946 608 1050
rect 653 1028 654 1038
rect 669 1028 682 1038
rect 653 1024 682 1028
rect 687 1024 717 1050
rect 735 1036 751 1038
rect 823 1036 876 1050
rect 824 1034 888 1036
rect 931 1034 946 1050
rect 995 1047 1025 1050
rect 995 1044 1031 1047
rect 961 1036 977 1038
rect 735 1024 750 1028
rect 653 1022 750 1024
rect 778 1022 946 1034
rect 962 1024 977 1028
rect 995 1025 1034 1044
rect 1053 1038 1060 1039
rect 1059 1031 1060 1038
rect 1043 1028 1044 1031
rect 1059 1028 1072 1031
rect 995 1024 1025 1025
rect 1034 1024 1040 1025
rect 1043 1024 1072 1028
rect 962 1023 1072 1024
rect 962 1022 1078 1023
rect 637 1014 688 1022
rect 637 1002 662 1014
rect 669 1002 688 1014
rect 719 1014 769 1022
rect 719 1006 735 1014
rect 742 1012 769 1014
rect 778 1012 999 1022
rect 742 1002 999 1012
rect 1028 1014 1078 1022
rect 1028 1005 1044 1014
rect 637 994 688 1002
rect 735 994 999 1002
rect 1025 1002 1044 1005
rect 1051 1002 1078 1014
rect 1025 994 1078 1002
rect 653 986 654 994
rect 669 986 682 994
rect 653 978 669 986
rect 650 971 669 974
rect 650 962 672 971
rect 623 952 672 962
rect 623 946 653 952
rect 672 947 677 952
rect 595 930 669 946
rect 687 938 717 994
rect 752 984 960 994
rect 995 990 1040 994
rect 1043 993 1044 994
rect 1059 993 1072 994
rect 778 954 967 984
rect 793 951 967 954
rect 786 948 967 951
rect 595 928 608 930
rect 623 928 657 930
rect 595 912 669 928
rect 696 924 709 938
rect 724 924 740 940
rect 786 935 797 948
rect 579 890 580 906
rect 595 890 608 912
rect 623 890 653 912
rect 696 908 758 924
rect 786 917 797 933
rect 802 928 812 948
rect 822 928 836 948
rect 839 935 848 948
rect 864 935 873 948
rect 802 917 836 928
rect 839 917 848 933
rect 864 917 873 933
rect 880 928 890 948
rect 900 928 914 948
rect 915 935 926 948
rect 880 917 914 928
rect 915 917 926 933
rect 972 924 988 940
rect 995 938 1025 990
rect 1059 986 1060 993
rect 1044 978 1060 986
rect 1031 946 1044 965
rect 1059 946 1089 962
rect 1031 930 1105 946
rect 1031 928 1044 930
rect 1059 928 1093 930
rect 696 906 709 908
rect 724 906 758 908
rect 696 890 758 906
rect 802 901 818 904
rect 880 901 910 912
rect 958 908 1004 924
rect 1031 912 1105 928
rect 958 906 992 908
rect 957 890 1004 906
rect 1031 890 1044 912
rect 1059 890 1089 912
rect 1116 890 1117 906
rect 1132 890 1145 1050
rect 1175 946 1188 1050
rect 1233 1028 1234 1038
rect 1249 1028 1262 1038
rect 1233 1024 1262 1028
rect 1267 1024 1297 1050
rect 1315 1036 1331 1038
rect 1403 1036 1456 1050
rect 1404 1034 1468 1036
rect 1511 1034 1526 1050
rect 1575 1047 1605 1050
rect 1575 1044 1611 1047
rect 1541 1036 1557 1038
rect 1315 1024 1330 1028
rect 1233 1022 1330 1024
rect 1358 1022 1526 1034
rect 1542 1024 1557 1028
rect 1575 1025 1614 1044
rect 1633 1038 1640 1039
rect 1639 1031 1640 1038
rect 1623 1028 1624 1031
rect 1639 1028 1652 1031
rect 1575 1024 1605 1025
rect 1614 1024 1620 1025
rect 1623 1024 1652 1028
rect 1542 1023 1652 1024
rect 1542 1022 1658 1023
rect 1217 1014 1268 1022
rect 1217 1002 1242 1014
rect 1249 1002 1268 1014
rect 1299 1014 1349 1022
rect 1299 1006 1315 1014
rect 1322 1012 1349 1014
rect 1358 1012 1579 1022
rect 1322 1002 1579 1012
rect 1608 1014 1658 1022
rect 1608 1005 1624 1014
rect 1217 994 1268 1002
rect 1315 994 1579 1002
rect 1605 1002 1624 1005
rect 1631 1002 1658 1014
rect 1605 994 1658 1002
rect 1233 986 1234 994
rect 1249 986 1262 994
rect 1233 978 1249 986
rect 1230 971 1249 974
rect 1230 962 1252 971
rect 1203 952 1252 962
rect 1203 946 1233 952
rect 1252 947 1257 952
rect 1175 930 1249 946
rect 1267 938 1297 994
rect 1332 984 1540 994
rect 1575 990 1620 994
rect 1623 993 1624 994
rect 1639 993 1652 994
rect 1358 954 1547 984
rect 1373 951 1547 954
rect 1366 948 1547 951
rect 1175 928 1188 930
rect 1203 928 1237 930
rect 1175 912 1249 928
rect 1276 924 1289 938
rect 1304 924 1320 940
rect 1366 935 1377 948
rect 1159 890 1160 906
rect 1175 890 1188 912
rect 1203 890 1233 912
rect 1276 908 1338 924
rect 1366 917 1377 933
rect 1382 928 1392 948
rect 1402 928 1416 948
rect 1419 935 1428 948
rect 1444 935 1453 948
rect 1382 917 1416 928
rect 1419 917 1428 933
rect 1444 917 1453 933
rect 1460 928 1470 948
rect 1480 928 1494 948
rect 1495 935 1506 948
rect 1460 917 1494 928
rect 1495 917 1506 933
rect 1552 924 1568 940
rect 1575 938 1605 990
rect 1639 986 1640 993
rect 1624 978 1640 986
rect 1611 946 1624 965
rect 1639 946 1669 962
rect 1611 930 1685 946
rect 1611 928 1624 930
rect 1639 928 1673 930
rect 1276 906 1289 908
rect 1304 906 1338 908
rect 1276 890 1338 906
rect 1382 901 1398 904
rect 1460 901 1490 912
rect 1538 908 1584 924
rect 1611 912 1685 928
rect 1538 906 1572 908
rect 1537 890 1584 906
rect 1611 890 1624 912
rect 1639 890 1669 912
rect 1696 890 1697 906
rect 1712 890 1725 1050
rect 1755 946 1768 1050
rect 1813 1028 1814 1038
rect 1829 1028 1842 1038
rect 1813 1024 1842 1028
rect 1847 1024 1877 1050
rect 1895 1036 1911 1038
rect 1983 1036 2036 1050
rect 1984 1034 2048 1036
rect 2091 1034 2106 1050
rect 2155 1047 2185 1050
rect 2155 1044 2191 1047
rect 2121 1036 2137 1038
rect 1895 1024 1910 1028
rect 1813 1022 1910 1024
rect 1938 1022 2106 1034
rect 2122 1024 2137 1028
rect 2155 1025 2194 1044
rect 2213 1038 2220 1039
rect 2219 1031 2220 1038
rect 2203 1028 2204 1031
rect 2219 1028 2232 1031
rect 2155 1024 2185 1025
rect 2194 1024 2200 1025
rect 2203 1024 2232 1028
rect 2122 1023 2232 1024
rect 2122 1022 2238 1023
rect 1797 1014 1848 1022
rect 1797 1002 1822 1014
rect 1829 1002 1848 1014
rect 1879 1014 1929 1022
rect 1879 1006 1895 1014
rect 1902 1012 1929 1014
rect 1938 1012 2159 1022
rect 1902 1002 2159 1012
rect 2188 1014 2238 1022
rect 2188 1005 2204 1014
rect 1797 994 1848 1002
rect 1895 994 2159 1002
rect 2185 1002 2204 1005
rect 2211 1002 2238 1014
rect 2185 994 2238 1002
rect 1813 986 1814 994
rect 1829 986 1842 994
rect 1813 978 1829 986
rect 1810 971 1829 974
rect 1810 962 1832 971
rect 1783 952 1832 962
rect 1783 946 1813 952
rect 1832 947 1837 952
rect 1755 930 1829 946
rect 1847 938 1877 994
rect 1912 984 2120 994
rect 2155 990 2200 994
rect 2203 993 2204 994
rect 2219 993 2232 994
rect 1938 954 2127 984
rect 1953 951 2127 954
rect 1946 948 2127 951
rect 1755 928 1768 930
rect 1783 928 1817 930
rect 1755 912 1829 928
rect 1856 924 1869 938
rect 1884 924 1900 940
rect 1946 935 1957 948
rect 1739 890 1740 906
rect 1755 890 1768 912
rect 1783 890 1813 912
rect 1856 908 1918 924
rect 1946 917 1957 933
rect 1962 928 1972 948
rect 1982 928 1996 948
rect 1999 935 2008 948
rect 2024 935 2033 948
rect 1962 917 1996 928
rect 1999 917 2008 933
rect 2024 917 2033 933
rect 2040 928 2050 948
rect 2060 928 2074 948
rect 2075 935 2086 948
rect 2040 917 2074 928
rect 2075 917 2086 933
rect 2132 924 2148 940
rect 2155 938 2185 990
rect 2219 986 2220 993
rect 2204 978 2220 986
rect 2191 946 2204 965
rect 2219 946 2249 962
rect 2191 930 2265 946
rect 2191 928 2204 930
rect 2219 928 2253 930
rect 1856 906 1869 908
rect 1884 906 1918 908
rect 1856 890 1918 906
rect 1962 901 1976 904
rect 2040 901 2070 912
rect 2118 908 2164 924
rect 2191 912 2265 928
rect 2118 906 2152 908
rect 2117 890 2164 906
rect 2191 890 2204 912
rect 2219 890 2249 912
rect 2276 890 2277 906
rect 2292 890 2305 1050
rect 2335 946 2348 1050
rect 2393 1028 2394 1038
rect 2409 1028 2422 1038
rect 2393 1024 2422 1028
rect 2427 1024 2457 1050
rect 2475 1036 2491 1038
rect 2563 1036 2616 1050
rect 2564 1034 2628 1036
rect 2671 1034 2686 1050
rect 2735 1047 2765 1050
rect 2735 1044 2771 1047
rect 2701 1036 2717 1038
rect 2475 1024 2490 1028
rect 2393 1022 2490 1024
rect 2518 1022 2686 1034
rect 2702 1024 2717 1028
rect 2735 1025 2774 1044
rect 2793 1038 2800 1039
rect 2799 1031 2800 1038
rect 2783 1028 2784 1031
rect 2799 1028 2812 1031
rect 2735 1024 2765 1025
rect 2774 1024 2780 1025
rect 2783 1024 2812 1028
rect 2702 1023 2812 1024
rect 2702 1022 2818 1023
rect 2377 1014 2428 1022
rect 2377 1002 2402 1014
rect 2409 1002 2428 1014
rect 2459 1014 2509 1022
rect 2459 1006 2475 1014
rect 2482 1012 2509 1014
rect 2518 1012 2739 1022
rect 2482 1002 2739 1012
rect 2768 1014 2818 1022
rect 2768 1005 2784 1014
rect 2377 994 2428 1002
rect 2475 994 2739 1002
rect 2765 1002 2784 1005
rect 2791 1002 2818 1014
rect 2765 994 2818 1002
rect 2393 986 2394 994
rect 2409 986 2422 994
rect 2393 978 2409 986
rect 2390 971 2409 974
rect 2390 962 2412 971
rect 2363 952 2412 962
rect 2363 946 2393 952
rect 2412 947 2417 952
rect 2335 930 2409 946
rect 2427 938 2457 994
rect 2492 984 2700 994
rect 2735 990 2780 994
rect 2783 993 2784 994
rect 2799 993 2812 994
rect 2518 954 2707 984
rect 2533 951 2707 954
rect 2526 948 2707 951
rect 2335 928 2348 930
rect 2363 928 2397 930
rect 2335 912 2409 928
rect 2436 924 2449 938
rect 2464 924 2480 940
rect 2526 935 2537 948
rect 2319 890 2320 906
rect 2335 890 2348 912
rect 2363 890 2393 912
rect 2436 908 2498 924
rect 2526 917 2537 933
rect 2542 928 2552 948
rect 2562 928 2576 948
rect 2579 935 2588 948
rect 2604 935 2613 948
rect 2542 917 2576 928
rect 2579 917 2588 933
rect 2604 917 2613 933
rect 2620 928 2630 948
rect 2640 928 2654 948
rect 2655 935 2666 948
rect 2620 917 2654 928
rect 2655 917 2666 933
rect 2712 924 2728 940
rect 2735 938 2765 990
rect 2799 986 2800 993
rect 2784 978 2800 986
rect 2771 946 2784 965
rect 2799 946 2829 962
rect 2771 930 2845 946
rect 2771 928 2784 930
rect 2799 928 2833 930
rect 2436 906 2449 908
rect 2464 906 2498 908
rect 2436 890 2498 906
rect 2542 901 2558 904
rect 2620 901 2650 912
rect 2698 908 2744 924
rect 2771 912 2845 928
rect 2698 906 2732 908
rect 2697 890 2744 906
rect 2771 890 2784 912
rect 2799 890 2829 912
rect 2856 890 2857 906
rect 2872 890 2885 1050
rect 2915 946 2928 1050
rect 2973 1028 2974 1038
rect 2989 1028 3002 1038
rect 2973 1024 3002 1028
rect 3007 1024 3037 1050
rect 3055 1036 3071 1038
rect 3143 1036 3196 1050
rect 3144 1034 3208 1036
rect 3251 1034 3266 1050
rect 3315 1047 3345 1050
rect 3315 1044 3351 1047
rect 3281 1036 3297 1038
rect 3055 1024 3070 1028
rect 2973 1022 3070 1024
rect 3098 1022 3266 1034
rect 3282 1024 3297 1028
rect 3315 1025 3354 1044
rect 3373 1038 3380 1039
rect 3379 1031 3380 1038
rect 3363 1028 3364 1031
rect 3379 1028 3392 1031
rect 3315 1024 3345 1025
rect 3354 1024 3360 1025
rect 3363 1024 3392 1028
rect 3282 1023 3392 1024
rect 3282 1022 3398 1023
rect 2957 1014 3008 1022
rect 2957 1002 2982 1014
rect 2989 1002 3008 1014
rect 3039 1014 3089 1022
rect 3039 1006 3055 1014
rect 3062 1012 3089 1014
rect 3098 1012 3319 1022
rect 3062 1002 3319 1012
rect 3348 1014 3398 1022
rect 3348 1005 3364 1014
rect 2957 994 3008 1002
rect 3055 994 3319 1002
rect 3345 1002 3364 1005
rect 3371 1002 3398 1014
rect 3345 994 3398 1002
rect 2973 986 2974 994
rect 2989 986 3002 994
rect 2973 978 2989 986
rect 2970 971 2989 974
rect 2970 962 2992 971
rect 2943 952 2992 962
rect 2943 946 2973 952
rect 2992 947 2997 952
rect 2915 930 2989 946
rect 3007 938 3037 994
rect 3072 984 3280 994
rect 3315 990 3360 994
rect 3363 993 3364 994
rect 3379 993 3392 994
rect 3098 954 3287 984
rect 3113 951 3287 954
rect 3106 948 3287 951
rect 2915 928 2928 930
rect 2943 928 2977 930
rect 2915 912 2989 928
rect 3016 924 3029 938
rect 3044 924 3060 940
rect 3106 935 3117 948
rect 2899 890 2900 906
rect 2915 890 2928 912
rect 2943 890 2973 912
rect 3016 908 3078 924
rect 3106 917 3117 933
rect 3122 928 3132 948
rect 3142 928 3156 948
rect 3159 935 3168 948
rect 3184 935 3193 948
rect 3122 917 3156 928
rect 3159 917 3168 933
rect 3184 917 3193 933
rect 3200 928 3210 948
rect 3220 928 3234 948
rect 3235 935 3246 948
rect 3200 917 3234 928
rect 3235 917 3246 933
rect 3292 924 3308 940
rect 3315 938 3345 990
rect 3379 986 3380 993
rect 3364 978 3380 986
rect 3351 946 3364 965
rect 3379 946 3409 962
rect 3351 930 3425 946
rect 3351 928 3364 930
rect 3379 928 3413 930
rect 3016 906 3029 908
rect 3044 906 3078 908
rect 3016 890 3078 906
rect 3122 901 3138 904
rect 3200 901 3230 912
rect 3278 908 3324 924
rect 3351 912 3425 928
rect 3278 906 3312 908
rect 3277 890 3324 906
rect 3351 890 3364 912
rect 3379 890 3409 912
rect 3436 890 3437 906
rect 3452 890 3465 1050
rect 3495 946 3508 1050
rect 3553 1028 3554 1038
rect 3569 1028 3582 1038
rect 3553 1024 3582 1028
rect 3587 1024 3617 1050
rect 3635 1036 3651 1038
rect 3723 1036 3776 1050
rect 3724 1034 3788 1036
rect 3831 1034 3846 1050
rect 3895 1047 3925 1050
rect 3895 1044 3931 1047
rect 3861 1036 3877 1038
rect 3635 1024 3650 1028
rect 3553 1022 3650 1024
rect 3678 1022 3846 1034
rect 3862 1024 3877 1028
rect 3895 1025 3934 1044
rect 3953 1038 3960 1039
rect 3959 1031 3960 1038
rect 3943 1028 3944 1031
rect 3959 1028 3972 1031
rect 3895 1024 3925 1025
rect 3934 1024 3940 1025
rect 3943 1024 3972 1028
rect 3862 1023 3972 1024
rect 3862 1022 3978 1023
rect 3537 1014 3588 1022
rect 3537 1002 3562 1014
rect 3569 1002 3588 1014
rect 3619 1014 3669 1022
rect 3619 1006 3635 1014
rect 3642 1012 3669 1014
rect 3678 1012 3899 1022
rect 3642 1002 3899 1012
rect 3928 1014 3978 1022
rect 3928 1005 3944 1014
rect 3537 994 3588 1002
rect 3635 994 3899 1002
rect 3925 1002 3944 1005
rect 3951 1002 3978 1014
rect 3925 994 3978 1002
rect 3553 986 3554 994
rect 3569 986 3582 994
rect 3553 978 3569 986
rect 3550 971 3569 974
rect 3550 962 3572 971
rect 3523 952 3572 962
rect 3523 946 3553 952
rect 3572 947 3577 952
rect 3495 930 3569 946
rect 3587 938 3617 994
rect 3652 984 3860 994
rect 3895 990 3940 994
rect 3943 993 3944 994
rect 3959 993 3972 994
rect 3678 954 3867 984
rect 3693 951 3867 954
rect 3686 948 3867 951
rect 3495 928 3508 930
rect 3523 928 3557 930
rect 3495 912 3569 928
rect 3596 924 3609 938
rect 3624 924 3640 940
rect 3686 935 3697 948
rect 3479 890 3480 906
rect 3495 890 3508 912
rect 3523 890 3553 912
rect 3596 908 3658 924
rect 3686 917 3697 933
rect 3702 928 3712 948
rect 3722 928 3736 948
rect 3739 935 3748 948
rect 3764 935 3773 948
rect 3702 917 3736 928
rect 3739 917 3748 933
rect 3764 917 3773 933
rect 3780 928 3790 948
rect 3800 928 3814 948
rect 3815 935 3826 948
rect 3780 917 3814 928
rect 3815 917 3826 933
rect 3872 924 3888 940
rect 3895 938 3925 990
rect 3959 986 3960 993
rect 3944 978 3960 986
rect 3931 946 3944 965
rect 3959 946 3989 962
rect 3931 930 4005 946
rect 3931 928 3944 930
rect 3959 928 3993 930
rect 3596 906 3609 908
rect 3624 906 3658 908
rect 3596 890 3658 906
rect 3702 901 3718 904
rect 3780 901 3810 912
rect 3858 908 3904 924
rect 3931 912 4005 928
rect 3858 906 3892 908
rect 3857 890 3904 906
rect 3931 890 3944 912
rect 3959 890 3989 912
rect 4016 890 4017 906
rect 4032 890 4045 1050
rect 4075 946 4088 1050
rect 4133 1028 4134 1038
rect 4149 1028 4162 1038
rect 4133 1024 4162 1028
rect 4167 1024 4197 1050
rect 4215 1036 4231 1038
rect 4303 1036 4356 1050
rect 4304 1034 4368 1036
rect 4411 1034 4426 1050
rect 4475 1047 4505 1050
rect 4475 1044 4511 1047
rect 4441 1036 4457 1038
rect 4215 1024 4230 1028
rect 4133 1022 4230 1024
rect 4258 1022 4426 1034
rect 4442 1024 4457 1028
rect 4475 1025 4514 1044
rect 4533 1038 4540 1039
rect 4539 1031 4540 1038
rect 4523 1028 4524 1031
rect 4539 1028 4552 1031
rect 4475 1024 4505 1025
rect 4514 1024 4520 1025
rect 4523 1024 4552 1028
rect 4442 1023 4552 1024
rect 4442 1022 4558 1023
rect 4117 1014 4168 1022
rect 4117 1002 4142 1014
rect 4149 1002 4168 1014
rect 4199 1014 4249 1022
rect 4199 1006 4215 1014
rect 4222 1012 4249 1014
rect 4258 1012 4479 1022
rect 4222 1002 4479 1012
rect 4508 1014 4558 1022
rect 4508 1005 4524 1014
rect 4117 994 4168 1002
rect 4215 994 4479 1002
rect 4505 1002 4524 1005
rect 4531 1002 4558 1014
rect 4505 994 4558 1002
rect 4133 986 4134 994
rect 4149 986 4162 994
rect 4133 978 4149 986
rect 4130 971 4149 974
rect 4130 962 4152 971
rect 4103 952 4152 962
rect 4103 946 4133 952
rect 4152 947 4157 952
rect 4075 930 4149 946
rect 4167 938 4197 994
rect 4232 984 4440 994
rect 4475 990 4520 994
rect 4523 993 4524 994
rect 4539 993 4552 994
rect 4258 954 4447 984
rect 4273 951 4447 954
rect 4266 948 4447 951
rect 4075 928 4088 930
rect 4103 928 4137 930
rect 4075 912 4149 928
rect 4176 924 4189 938
rect 4204 924 4220 940
rect 4266 935 4277 948
rect 4059 890 4060 906
rect 4075 890 4088 912
rect 4103 890 4133 912
rect 4176 908 4238 924
rect 4266 917 4277 933
rect 4282 928 4292 948
rect 4302 928 4316 948
rect 4319 935 4328 948
rect 4344 935 4353 948
rect 4282 917 4316 928
rect 4319 917 4328 933
rect 4344 917 4353 933
rect 4360 928 4370 948
rect 4380 928 4394 948
rect 4395 935 4406 948
rect 4360 917 4394 928
rect 4395 917 4406 933
rect 4452 924 4468 940
rect 4475 938 4505 990
rect 4539 986 4540 993
rect 4524 978 4540 986
rect 4511 946 4524 965
rect 4539 946 4569 962
rect 4511 930 4585 946
rect 4511 928 4524 930
rect 4539 928 4573 930
rect 4176 906 4189 908
rect 4204 906 4238 908
rect 4176 890 4238 906
rect 4282 901 4298 904
rect 4360 901 4390 912
rect 4438 908 4484 924
rect 4511 912 4585 928
rect 4438 906 4472 908
rect 4437 890 4484 906
rect 4511 890 4524 912
rect 4539 890 4569 912
rect 4596 890 4597 906
rect 4612 890 4625 1050
rect 4655 946 4668 1050
rect 4713 1028 4714 1038
rect 4729 1028 4742 1038
rect 4713 1024 4742 1028
rect 4747 1024 4777 1050
rect 4795 1036 4811 1038
rect 4883 1036 4936 1050
rect 4884 1034 4948 1036
rect 4991 1034 5006 1050
rect 5055 1047 5085 1050
rect 5055 1044 5091 1047
rect 5021 1036 5037 1038
rect 4795 1024 4810 1028
rect 4713 1022 4810 1024
rect 4838 1022 5006 1034
rect 5022 1024 5037 1028
rect 5055 1025 5094 1044
rect 5113 1038 5120 1039
rect 5119 1031 5120 1038
rect 5103 1028 5104 1031
rect 5119 1028 5132 1031
rect 5055 1024 5085 1025
rect 5094 1024 5100 1025
rect 5103 1024 5132 1028
rect 5022 1023 5132 1024
rect 5022 1022 5138 1023
rect 4697 1014 4748 1022
rect 4697 1002 4722 1014
rect 4729 1002 4748 1014
rect 4779 1014 4829 1022
rect 4779 1006 4795 1014
rect 4802 1012 4829 1014
rect 4838 1012 5059 1022
rect 4802 1002 5059 1012
rect 5088 1014 5138 1022
rect 5088 1005 5104 1014
rect 4697 994 4748 1002
rect 4795 994 5059 1002
rect 5085 1002 5104 1005
rect 5111 1002 5138 1014
rect 5085 994 5138 1002
rect 4713 986 4714 994
rect 4729 986 4742 994
rect 4713 978 4729 986
rect 4710 971 4729 974
rect 4710 962 4732 971
rect 4683 952 4732 962
rect 4683 946 4713 952
rect 4732 947 4737 952
rect 4655 930 4729 946
rect 4747 938 4777 994
rect 4812 984 5020 994
rect 5055 990 5100 994
rect 5103 993 5104 994
rect 5119 993 5132 994
rect 4838 954 5027 984
rect 4853 951 5027 954
rect 4846 948 5027 951
rect 4655 928 4668 930
rect 4683 928 4717 930
rect 4655 912 4729 928
rect 4756 924 4769 938
rect 4784 924 4800 940
rect 4846 935 4857 948
rect 4639 890 4640 906
rect 4655 890 4668 912
rect 4683 890 4713 912
rect 4756 908 4818 924
rect 4846 917 4857 933
rect 4862 928 4872 948
rect 4882 928 4896 948
rect 4899 935 4908 948
rect 4924 935 4933 948
rect 4862 917 4896 928
rect 4899 917 4908 933
rect 4924 917 4933 933
rect 4940 928 4950 948
rect 4960 928 4974 948
rect 4975 935 4986 948
rect 4940 917 4974 928
rect 4975 917 4986 933
rect 5032 924 5048 940
rect 5055 938 5085 990
rect 5119 986 5120 993
rect 5104 978 5120 986
rect 5091 946 5104 965
rect 5119 946 5149 962
rect 5091 930 5165 946
rect 5091 928 5104 930
rect 5119 928 5153 930
rect 4756 906 4769 908
rect 4784 906 4818 908
rect 4756 890 4818 906
rect 4862 901 4878 904
rect 4940 901 4970 912
rect 5018 908 5064 924
rect 5091 912 5165 928
rect 5018 906 5052 908
rect 5017 890 5064 906
rect 5091 890 5104 912
rect 5119 890 5149 912
rect 5176 890 5177 906
rect 5192 890 5205 1050
rect 5235 946 5248 1050
rect 5293 1028 5294 1038
rect 5309 1028 5322 1038
rect 5293 1024 5322 1028
rect 5327 1024 5357 1050
rect 5375 1036 5391 1038
rect 5463 1036 5516 1050
rect 5464 1034 5528 1036
rect 5571 1034 5586 1050
rect 5635 1047 5665 1050
rect 5635 1044 5671 1047
rect 5601 1036 5617 1038
rect 5375 1024 5390 1028
rect 5293 1022 5390 1024
rect 5418 1022 5586 1034
rect 5602 1024 5617 1028
rect 5635 1025 5674 1044
rect 5693 1038 5700 1039
rect 5699 1031 5700 1038
rect 5683 1028 5684 1031
rect 5699 1028 5712 1031
rect 5635 1024 5665 1025
rect 5674 1024 5680 1025
rect 5683 1024 5712 1028
rect 5602 1023 5712 1024
rect 5602 1022 5718 1023
rect 5277 1014 5328 1022
rect 5277 1002 5302 1014
rect 5309 1002 5328 1014
rect 5359 1014 5409 1022
rect 5359 1006 5375 1014
rect 5382 1012 5409 1014
rect 5418 1012 5639 1022
rect 5382 1002 5639 1012
rect 5668 1014 5718 1022
rect 5668 1005 5684 1014
rect 5277 994 5328 1002
rect 5375 994 5639 1002
rect 5665 1002 5684 1005
rect 5691 1002 5718 1014
rect 5665 994 5718 1002
rect 5293 986 5294 994
rect 5309 986 5322 994
rect 5293 978 5309 986
rect 5290 971 5309 974
rect 5290 962 5312 971
rect 5263 952 5312 962
rect 5263 946 5293 952
rect 5312 947 5317 952
rect 5235 930 5309 946
rect 5327 938 5357 994
rect 5392 984 5600 994
rect 5635 990 5680 994
rect 5683 993 5684 994
rect 5699 993 5712 994
rect 5418 954 5607 984
rect 5433 951 5607 954
rect 5426 948 5607 951
rect 5235 928 5248 930
rect 5263 928 5297 930
rect 5235 912 5309 928
rect 5336 924 5349 938
rect 5364 924 5380 940
rect 5426 935 5437 948
rect 5219 890 5220 906
rect 5235 890 5248 912
rect 5263 890 5293 912
rect 5336 908 5398 924
rect 5426 917 5437 933
rect 5442 928 5452 948
rect 5462 928 5476 948
rect 5479 935 5488 948
rect 5504 935 5513 948
rect 5442 917 5476 928
rect 5479 917 5488 933
rect 5504 917 5513 933
rect 5520 928 5530 948
rect 5540 928 5554 948
rect 5555 935 5566 948
rect 5520 917 5554 928
rect 5555 917 5566 933
rect 5612 924 5628 940
rect 5635 938 5665 990
rect 5699 986 5700 993
rect 5684 978 5700 986
rect 5671 946 5684 965
rect 5699 946 5729 962
rect 5671 930 5745 946
rect 5671 928 5684 930
rect 5699 928 5733 930
rect 5336 906 5349 908
rect 5364 906 5398 908
rect 5336 890 5398 906
rect 5442 901 5458 904
rect 5520 901 5550 912
rect 5598 908 5644 924
rect 5671 912 5745 928
rect 5598 906 5632 908
rect 5597 890 5644 906
rect 5671 890 5684 912
rect 5699 890 5729 912
rect 5756 890 5757 906
rect 5772 890 5785 1050
rect 5815 946 5828 1050
rect 5873 1028 5874 1038
rect 5889 1028 5902 1038
rect 5873 1024 5902 1028
rect 5907 1024 5937 1050
rect 5955 1036 5971 1038
rect 6043 1036 6096 1050
rect 6044 1034 6108 1036
rect 6151 1034 6166 1050
rect 6215 1047 6245 1050
rect 6215 1044 6251 1047
rect 6181 1036 6197 1038
rect 5955 1024 5970 1028
rect 5873 1022 5970 1024
rect 5998 1022 6166 1034
rect 6182 1024 6197 1028
rect 6215 1025 6254 1044
rect 6273 1038 6280 1039
rect 6279 1031 6280 1038
rect 6263 1028 6264 1031
rect 6279 1028 6292 1031
rect 6215 1024 6245 1025
rect 6254 1024 6260 1025
rect 6263 1024 6292 1028
rect 6182 1023 6292 1024
rect 6182 1022 6298 1023
rect 5857 1014 5908 1022
rect 5857 1002 5882 1014
rect 5889 1002 5908 1014
rect 5939 1014 5989 1022
rect 5939 1006 5955 1014
rect 5962 1012 5989 1014
rect 5998 1012 6219 1022
rect 5962 1002 6219 1012
rect 6248 1014 6298 1022
rect 6248 1005 6264 1014
rect 5857 994 5908 1002
rect 5955 994 6219 1002
rect 6245 1002 6264 1005
rect 6271 1002 6298 1014
rect 6245 994 6298 1002
rect 5873 986 5874 994
rect 5889 986 5902 994
rect 5873 978 5889 986
rect 5870 971 5889 974
rect 5870 962 5892 971
rect 5843 952 5892 962
rect 5843 946 5873 952
rect 5892 947 5897 952
rect 5815 930 5889 946
rect 5907 938 5937 994
rect 5972 984 6180 994
rect 6215 990 6260 994
rect 6263 993 6264 994
rect 6279 993 6292 994
rect 5998 954 6187 984
rect 6013 951 6187 954
rect 6006 948 6187 951
rect 5815 928 5828 930
rect 5843 928 5877 930
rect 5815 912 5889 928
rect 5916 924 5929 938
rect 5944 924 5960 940
rect 6006 935 6017 948
rect 5799 890 5800 906
rect 5815 890 5828 912
rect 5843 890 5873 912
rect 5916 908 5978 924
rect 6006 917 6017 933
rect 6022 928 6032 948
rect 6042 928 6056 948
rect 6059 935 6068 948
rect 6084 935 6093 948
rect 6022 917 6056 928
rect 6059 917 6068 933
rect 6084 917 6093 933
rect 6100 928 6110 948
rect 6120 928 6134 948
rect 6135 935 6146 948
rect 6100 917 6134 928
rect 6135 917 6146 933
rect 6192 924 6208 940
rect 6215 938 6245 990
rect 6279 986 6280 993
rect 6264 978 6280 986
rect 6251 946 6264 965
rect 6279 946 6309 962
rect 6251 930 6325 946
rect 6251 928 6264 930
rect 6279 928 6313 930
rect 5916 906 5929 908
rect 5944 906 5978 908
rect 5916 890 5978 906
rect 6022 901 6038 904
rect 6100 901 6130 912
rect 6178 908 6224 924
rect 6251 912 6325 928
rect 6178 906 6212 908
rect 6177 890 6224 906
rect 6251 890 6264 912
rect 6279 890 6309 912
rect 6336 890 6337 906
rect 6352 890 6365 1050
rect 6395 946 6408 1050
rect 6453 1028 6454 1038
rect 6469 1028 6482 1038
rect 6453 1024 6482 1028
rect 6487 1024 6517 1050
rect 6535 1036 6551 1038
rect 6623 1036 6676 1050
rect 6624 1034 6688 1036
rect 6731 1034 6746 1050
rect 6795 1047 6825 1050
rect 6795 1044 6831 1047
rect 6761 1036 6777 1038
rect 6535 1024 6550 1028
rect 6453 1022 6550 1024
rect 6578 1022 6746 1034
rect 6762 1024 6777 1028
rect 6795 1025 6834 1044
rect 6853 1038 6860 1039
rect 6859 1031 6860 1038
rect 6843 1028 6844 1031
rect 6859 1028 6872 1031
rect 6795 1024 6825 1025
rect 6834 1024 6840 1025
rect 6843 1024 6872 1028
rect 6762 1023 6872 1024
rect 6762 1022 6878 1023
rect 6437 1014 6488 1022
rect 6437 1002 6462 1014
rect 6469 1002 6488 1014
rect 6519 1014 6569 1022
rect 6519 1006 6535 1014
rect 6542 1012 6569 1014
rect 6578 1012 6799 1022
rect 6542 1002 6799 1012
rect 6828 1014 6878 1022
rect 6828 1005 6844 1014
rect 6437 994 6488 1002
rect 6535 994 6799 1002
rect 6825 1002 6844 1005
rect 6851 1002 6878 1014
rect 6825 994 6878 1002
rect 6453 986 6454 994
rect 6469 986 6482 994
rect 6453 978 6469 986
rect 6450 971 6469 974
rect 6450 962 6472 971
rect 6423 952 6472 962
rect 6423 946 6453 952
rect 6472 947 6477 952
rect 6395 930 6469 946
rect 6487 938 6517 994
rect 6552 984 6760 994
rect 6795 990 6840 994
rect 6843 993 6844 994
rect 6859 993 6872 994
rect 6578 954 6767 984
rect 6593 951 6767 954
rect 6586 948 6767 951
rect 6395 928 6408 930
rect 6423 928 6457 930
rect 6395 912 6469 928
rect 6496 924 6509 938
rect 6524 924 6540 940
rect 6586 935 6597 948
rect 6379 890 6380 906
rect 6395 890 6408 912
rect 6423 890 6453 912
rect 6496 908 6558 924
rect 6586 917 6597 933
rect 6602 928 6612 948
rect 6622 928 6636 948
rect 6639 935 6648 948
rect 6664 935 6673 948
rect 6602 917 6636 928
rect 6639 917 6648 933
rect 6664 917 6673 933
rect 6680 928 6690 948
rect 6700 928 6714 948
rect 6715 935 6726 948
rect 6680 917 6714 928
rect 6715 917 6726 933
rect 6772 924 6788 940
rect 6795 938 6825 990
rect 6859 986 6860 993
rect 6844 978 6860 986
rect 6831 946 6844 965
rect 6859 946 6889 962
rect 6831 930 6905 946
rect 6831 928 6844 930
rect 6859 928 6893 930
rect 6496 906 6509 908
rect 6524 906 6558 908
rect 6496 890 6558 906
rect 6602 901 6618 904
rect 6680 901 6710 912
rect 6758 908 6804 924
rect 6831 912 6905 928
rect 6758 906 6792 908
rect 6757 890 6804 906
rect 6831 890 6844 912
rect 6859 890 6889 912
rect 6916 890 6917 906
rect 6932 890 6945 1050
rect 6975 946 6988 1050
rect 7033 1028 7034 1038
rect 7049 1028 7062 1038
rect 7033 1024 7062 1028
rect 7067 1024 7097 1050
rect 7115 1036 7131 1038
rect 7203 1036 7256 1050
rect 7204 1034 7268 1036
rect 7311 1034 7326 1050
rect 7375 1047 7405 1050
rect 7375 1044 7411 1047
rect 7341 1036 7357 1038
rect 7115 1024 7130 1028
rect 7033 1022 7130 1024
rect 7158 1022 7326 1034
rect 7342 1024 7357 1028
rect 7375 1025 7414 1044
rect 7433 1038 7440 1039
rect 7439 1031 7440 1038
rect 7423 1028 7424 1031
rect 7439 1028 7452 1031
rect 7375 1024 7405 1025
rect 7414 1024 7420 1025
rect 7423 1024 7452 1028
rect 7342 1023 7452 1024
rect 7342 1022 7458 1023
rect 7017 1014 7068 1022
rect 7017 1002 7042 1014
rect 7049 1002 7068 1014
rect 7099 1014 7149 1022
rect 7099 1006 7115 1014
rect 7122 1012 7149 1014
rect 7158 1012 7379 1022
rect 7122 1002 7379 1012
rect 7408 1014 7458 1022
rect 7408 1005 7424 1014
rect 7017 994 7068 1002
rect 7115 994 7379 1002
rect 7405 1002 7424 1005
rect 7431 1002 7458 1014
rect 7405 994 7458 1002
rect 7033 986 7034 994
rect 7049 986 7062 994
rect 7033 978 7049 986
rect 7030 971 7049 974
rect 7030 962 7052 971
rect 7003 952 7052 962
rect 7003 946 7033 952
rect 7052 947 7057 952
rect 6975 930 7049 946
rect 7067 938 7097 994
rect 7132 984 7340 994
rect 7375 990 7420 994
rect 7423 993 7424 994
rect 7439 993 7452 994
rect 7158 954 7347 984
rect 7173 951 7347 954
rect 7166 948 7347 951
rect 6975 928 6988 930
rect 7003 928 7037 930
rect 6975 912 7049 928
rect 7076 924 7089 938
rect 7104 924 7120 940
rect 7166 935 7177 948
rect 6959 890 6960 906
rect 6975 890 6988 912
rect 7003 890 7033 912
rect 7076 908 7138 924
rect 7166 917 7177 933
rect 7182 928 7192 948
rect 7202 928 7216 948
rect 7219 935 7228 948
rect 7244 935 7253 948
rect 7182 917 7216 928
rect 7219 917 7228 933
rect 7244 917 7253 933
rect 7260 928 7270 948
rect 7280 928 7294 948
rect 7295 935 7306 948
rect 7260 917 7294 928
rect 7295 917 7306 933
rect 7352 924 7368 940
rect 7375 938 7405 990
rect 7439 986 7440 993
rect 7424 978 7440 986
rect 7411 946 7424 965
rect 7439 946 7469 962
rect 7411 930 7485 946
rect 7411 928 7424 930
rect 7439 928 7473 930
rect 7076 906 7089 908
rect 7104 906 7138 908
rect 7076 890 7138 906
rect 7182 901 7198 904
rect 7260 901 7290 912
rect 7338 908 7384 924
rect 7411 912 7485 928
rect 7338 906 7372 908
rect 7337 890 7384 906
rect 7411 890 7424 912
rect 7439 890 7469 912
rect 7496 890 7497 906
rect 7512 890 7525 1050
rect 7555 946 7568 1050
rect 7613 1028 7614 1038
rect 7629 1028 7642 1038
rect 7613 1024 7642 1028
rect 7647 1024 7677 1050
rect 7695 1036 7711 1038
rect 7783 1036 7836 1050
rect 7784 1034 7848 1036
rect 7891 1034 7906 1050
rect 7955 1047 7985 1050
rect 7955 1044 7991 1047
rect 7921 1036 7937 1038
rect 7695 1024 7710 1028
rect 7613 1022 7710 1024
rect 7738 1022 7906 1034
rect 7922 1024 7937 1028
rect 7955 1025 7994 1044
rect 8013 1038 8020 1039
rect 8019 1031 8020 1038
rect 8003 1028 8004 1031
rect 8019 1028 8032 1031
rect 7955 1024 7985 1025
rect 7994 1024 8000 1025
rect 8003 1024 8032 1028
rect 7922 1023 8032 1024
rect 7922 1022 8038 1023
rect 7597 1014 7648 1022
rect 7597 1002 7622 1014
rect 7629 1002 7648 1014
rect 7679 1014 7729 1022
rect 7679 1006 7695 1014
rect 7702 1012 7729 1014
rect 7738 1012 7959 1022
rect 7702 1002 7959 1012
rect 7988 1014 8038 1022
rect 7988 1005 8004 1014
rect 7597 994 7648 1002
rect 7695 994 7959 1002
rect 7985 1002 8004 1005
rect 8011 1002 8038 1014
rect 7985 994 8038 1002
rect 7613 986 7614 994
rect 7629 986 7642 994
rect 7613 978 7629 986
rect 7610 971 7629 974
rect 7610 962 7632 971
rect 7583 952 7632 962
rect 7583 946 7613 952
rect 7632 947 7637 952
rect 7555 930 7629 946
rect 7647 938 7677 994
rect 7712 984 7920 994
rect 7955 990 8000 994
rect 8003 993 8004 994
rect 8019 993 8032 994
rect 7738 954 7927 984
rect 7753 951 7927 954
rect 7746 948 7927 951
rect 7555 928 7568 930
rect 7583 928 7617 930
rect 7555 912 7629 928
rect 7656 924 7669 938
rect 7684 924 7700 940
rect 7746 935 7757 948
rect 7539 890 7540 906
rect 7555 890 7568 912
rect 7583 890 7613 912
rect 7656 908 7718 924
rect 7746 917 7757 933
rect 7762 928 7772 948
rect 7782 928 7796 948
rect 7799 935 7808 948
rect 7824 935 7833 948
rect 7762 917 7796 928
rect 7799 917 7808 933
rect 7824 917 7833 933
rect 7840 928 7850 948
rect 7860 928 7874 948
rect 7875 935 7886 948
rect 7840 917 7874 928
rect 7875 917 7886 933
rect 7932 924 7948 940
rect 7955 938 7985 990
rect 8019 986 8020 993
rect 8004 978 8020 986
rect 7991 946 8004 965
rect 8019 946 8049 962
rect 7991 930 8065 946
rect 7991 928 8004 930
rect 8019 928 8053 930
rect 7656 906 7669 908
rect 7684 906 7718 908
rect 7656 890 7718 906
rect 7762 901 7778 904
rect 7840 901 7870 912
rect 7918 908 7964 924
rect 7991 912 8065 928
rect 7918 906 7952 908
rect 7917 890 7964 906
rect 7991 890 8004 912
rect 8019 890 8049 912
rect 8076 890 8077 906
rect 8092 890 8105 1050
rect 8135 946 8148 1050
rect 8193 1028 8194 1038
rect 8209 1028 8222 1038
rect 8193 1024 8222 1028
rect 8227 1024 8257 1050
rect 8275 1036 8291 1038
rect 8363 1036 8416 1050
rect 8364 1034 8428 1036
rect 8471 1034 8486 1050
rect 8535 1047 8565 1050
rect 8535 1044 8571 1047
rect 8501 1036 8517 1038
rect 8275 1024 8290 1028
rect 8193 1022 8290 1024
rect 8318 1022 8486 1034
rect 8502 1024 8517 1028
rect 8535 1025 8574 1044
rect 8593 1038 8600 1039
rect 8599 1031 8600 1038
rect 8583 1028 8584 1031
rect 8599 1028 8612 1031
rect 8535 1024 8565 1025
rect 8574 1024 8580 1025
rect 8583 1024 8612 1028
rect 8502 1023 8612 1024
rect 8502 1022 8618 1023
rect 8177 1014 8228 1022
rect 8177 1002 8202 1014
rect 8209 1002 8228 1014
rect 8259 1014 8309 1022
rect 8259 1006 8275 1014
rect 8282 1012 8309 1014
rect 8318 1012 8539 1022
rect 8282 1002 8539 1012
rect 8568 1014 8618 1022
rect 8568 1005 8584 1014
rect 8177 994 8228 1002
rect 8275 994 8539 1002
rect 8565 1002 8584 1005
rect 8591 1002 8618 1014
rect 8565 994 8618 1002
rect 8193 986 8194 994
rect 8209 986 8222 994
rect 8193 978 8209 986
rect 8190 971 8209 974
rect 8190 962 8212 971
rect 8163 952 8212 962
rect 8163 946 8193 952
rect 8212 947 8217 952
rect 8135 930 8209 946
rect 8227 938 8257 994
rect 8292 984 8500 994
rect 8535 990 8580 994
rect 8583 993 8584 994
rect 8599 993 8612 994
rect 8318 954 8507 984
rect 8333 951 8507 954
rect 8326 948 8507 951
rect 8135 928 8148 930
rect 8163 928 8197 930
rect 8135 912 8209 928
rect 8236 924 8249 938
rect 8264 924 8280 940
rect 8326 935 8337 948
rect 8119 890 8120 906
rect 8135 890 8148 912
rect 8163 890 8193 912
rect 8236 908 8298 924
rect 8326 917 8337 933
rect 8342 928 8352 948
rect 8362 928 8376 948
rect 8379 935 8388 948
rect 8404 935 8413 948
rect 8342 917 8376 928
rect 8379 917 8388 933
rect 8404 917 8413 933
rect 8420 928 8430 948
rect 8440 928 8454 948
rect 8455 935 8466 948
rect 8420 917 8454 928
rect 8455 917 8466 933
rect 8512 924 8528 940
rect 8535 938 8565 990
rect 8599 986 8600 993
rect 8584 978 8600 986
rect 8571 946 8584 965
rect 8599 946 8629 962
rect 8571 930 8645 946
rect 8571 928 8584 930
rect 8599 928 8633 930
rect 8236 906 8249 908
rect 8264 906 8298 908
rect 8236 890 8298 906
rect 8342 901 8358 904
rect 8420 901 8450 912
rect 8498 908 8544 924
rect 8571 912 8645 928
rect 8498 906 8532 908
rect 8497 890 8544 906
rect 8571 890 8584 912
rect 8599 890 8629 912
rect 8656 890 8657 906
rect 8672 890 8685 1050
rect 8715 946 8728 1050
rect 8773 1028 8774 1038
rect 8789 1028 8802 1038
rect 8773 1024 8802 1028
rect 8807 1024 8837 1050
rect 8855 1036 8871 1038
rect 8943 1036 8996 1050
rect 8944 1034 9008 1036
rect 9051 1034 9066 1050
rect 9115 1047 9145 1050
rect 9115 1044 9151 1047
rect 9081 1036 9097 1038
rect 8855 1024 8870 1028
rect 8773 1022 8870 1024
rect 8898 1022 9066 1034
rect 9082 1024 9097 1028
rect 9115 1025 9154 1044
rect 9173 1038 9180 1039
rect 9179 1031 9180 1038
rect 9163 1028 9164 1031
rect 9179 1028 9192 1031
rect 9115 1024 9145 1025
rect 9154 1024 9160 1025
rect 9163 1024 9192 1028
rect 9082 1023 9192 1024
rect 9082 1022 9198 1023
rect 8757 1014 8808 1022
rect 8757 1002 8782 1014
rect 8789 1002 8808 1014
rect 8839 1014 8889 1022
rect 8839 1006 8855 1014
rect 8862 1012 8889 1014
rect 8898 1012 9119 1022
rect 8862 1002 9119 1012
rect 9148 1014 9198 1022
rect 9148 1005 9164 1014
rect 8757 994 8808 1002
rect 8855 994 9119 1002
rect 9145 1002 9164 1005
rect 9171 1002 9198 1014
rect 9145 994 9198 1002
rect 8773 986 8774 994
rect 8789 986 8802 994
rect 8773 978 8789 986
rect 8770 971 8789 974
rect 8770 962 8792 971
rect 8743 952 8792 962
rect 8743 946 8773 952
rect 8792 947 8797 952
rect 8715 930 8789 946
rect 8807 938 8837 994
rect 8872 984 9080 994
rect 9115 990 9160 994
rect 9163 993 9164 994
rect 9179 993 9192 994
rect 8898 954 9087 984
rect 8913 951 9087 954
rect 8906 948 9087 951
rect 8715 928 8728 930
rect 8743 928 8777 930
rect 8715 912 8789 928
rect 8816 924 8829 938
rect 8844 924 8860 940
rect 8906 935 8917 948
rect 8699 890 8700 906
rect 8715 890 8728 912
rect 8743 890 8773 912
rect 8816 908 8878 924
rect 8906 917 8917 933
rect 8922 928 8932 948
rect 8942 928 8956 948
rect 8959 935 8968 948
rect 8984 935 8993 948
rect 8922 917 8956 928
rect 8959 917 8968 933
rect 8984 917 8993 933
rect 9000 928 9010 948
rect 9020 928 9034 948
rect 9035 935 9046 948
rect 9000 917 9034 928
rect 9035 917 9046 933
rect 9092 924 9108 940
rect 9115 938 9145 990
rect 9179 986 9180 993
rect 9164 978 9180 986
rect 9151 946 9164 965
rect 9179 946 9209 962
rect 9151 930 9225 946
rect 9151 928 9164 930
rect 9179 928 9213 930
rect 8816 906 8829 908
rect 8844 906 8878 908
rect 8816 890 8878 906
rect 8922 901 8938 904
rect 9000 901 9030 912
rect 9078 908 9124 924
rect 9151 912 9225 928
rect 9078 906 9112 908
rect 9077 890 9124 906
rect 9151 890 9164 912
rect 9179 890 9209 912
rect 9236 890 9237 906
rect 9252 890 9265 1050
rect -7 882 34 890
rect -7 856 8 882
rect 15 856 34 882
rect 98 878 160 890
rect 172 878 247 890
rect 305 878 380 890
rect 392 878 423 890
rect 429 878 464 890
rect 98 876 260 878
rect -7 848 34 856
rect 116 852 129 876
rect 144 874 159 876
rect -1 838 0 848
rect 15 838 28 848
rect 43 838 73 852
rect 116 838 159 852
rect 183 849 190 856
rect 193 852 260 876
rect 292 876 464 878
rect 262 854 290 858
rect 292 854 372 876
rect 393 874 408 876
rect 262 852 372 854
rect 193 848 372 852
rect 166 838 196 848
rect 198 838 351 848
rect 359 838 389 848
rect 393 838 423 852
rect 451 838 464 876
rect 536 882 571 890
rect 536 856 537 882
rect 544 856 571 882
rect 479 838 509 852
rect 536 848 571 856
rect 573 882 614 890
rect 573 856 588 882
rect 595 856 614 882
rect 678 878 740 890
rect 752 878 827 890
rect 885 878 960 890
rect 972 878 1003 890
rect 1009 878 1044 890
rect 678 876 840 878
rect 573 848 614 856
rect 696 852 709 876
rect 724 874 739 876
rect 536 838 537 848
rect 552 838 565 848
rect 579 838 580 848
rect 595 838 608 848
rect 623 838 653 852
rect 696 838 739 852
rect 763 849 770 856
rect 773 852 840 876
rect 872 876 1044 878
rect 842 854 870 858
rect 872 854 952 876
rect 973 874 988 876
rect 842 852 952 854
rect 773 848 952 852
rect 746 838 776 848
rect 778 838 931 848
rect 939 838 969 848
rect 973 838 1003 852
rect 1031 838 1044 876
rect 1116 882 1151 890
rect 1116 856 1117 882
rect 1124 856 1151 882
rect 1059 838 1089 852
rect 1116 848 1151 856
rect 1153 882 1194 890
rect 1153 856 1168 882
rect 1175 856 1194 882
rect 1258 878 1320 890
rect 1332 878 1407 890
rect 1465 878 1540 890
rect 1552 878 1583 890
rect 1589 878 1624 890
rect 1258 876 1420 878
rect 1153 848 1194 856
rect 1276 852 1289 876
rect 1304 874 1319 876
rect 1116 838 1117 848
rect 1132 838 1145 848
rect 1159 838 1160 848
rect 1175 838 1188 848
rect 1203 838 1233 852
rect 1276 838 1319 852
rect 1343 849 1350 856
rect 1353 852 1420 876
rect 1452 876 1624 878
rect 1422 854 1450 858
rect 1452 854 1532 876
rect 1553 874 1568 876
rect 1422 852 1532 854
rect 1353 848 1532 852
rect 1326 838 1356 848
rect 1358 838 1511 848
rect 1519 838 1549 848
rect 1553 838 1583 852
rect 1611 838 1624 876
rect 1696 882 1731 890
rect 1696 856 1697 882
rect 1704 856 1731 882
rect 1639 838 1669 852
rect 1696 848 1731 856
rect 1733 882 1774 890
rect 1733 856 1748 882
rect 1755 856 1774 882
rect 1838 878 1900 890
rect 1912 878 1987 890
rect 2045 878 2120 890
rect 2132 878 2163 890
rect 2169 878 2204 890
rect 1838 876 2000 878
rect 1733 848 1774 856
rect 1856 852 1869 876
rect 1884 874 1899 876
rect 1696 838 1697 848
rect 1712 838 1725 848
rect 1739 838 1740 848
rect 1755 838 1768 848
rect 1783 838 1813 852
rect 1856 838 1899 852
rect 1923 849 1930 856
rect 1933 852 2000 876
rect 2032 876 2204 878
rect 2002 854 2030 858
rect 2032 854 2112 876
rect 2133 874 2148 876
rect 2002 852 2112 854
rect 1933 848 2112 852
rect 1906 838 1936 848
rect 1938 838 2091 848
rect 2099 838 2129 848
rect 2133 838 2163 852
rect 2191 838 2204 876
rect 2276 882 2311 890
rect 2276 856 2277 882
rect 2284 856 2311 882
rect 2219 838 2249 852
rect 2276 848 2311 856
rect 2313 882 2354 890
rect 2313 856 2328 882
rect 2335 856 2354 882
rect 2418 878 2480 890
rect 2492 878 2567 890
rect 2625 878 2700 890
rect 2712 878 2743 890
rect 2749 878 2784 890
rect 2418 876 2580 878
rect 2313 848 2354 856
rect 2436 852 2449 876
rect 2464 874 2479 876
rect 2276 838 2277 848
rect 2292 838 2305 848
rect 2319 838 2320 848
rect 2335 838 2348 848
rect 2363 838 2393 852
rect 2436 838 2479 852
rect 2503 849 2510 856
rect 2513 852 2580 876
rect 2612 876 2784 878
rect 2582 854 2610 858
rect 2612 854 2692 876
rect 2713 874 2728 876
rect 2582 852 2692 854
rect 2513 848 2692 852
rect 2486 838 2516 848
rect 2518 838 2671 848
rect 2679 838 2709 848
rect 2713 838 2743 852
rect 2771 838 2784 876
rect 2856 882 2891 890
rect 2856 856 2857 882
rect 2864 856 2891 882
rect 2799 838 2829 852
rect 2856 848 2891 856
rect 2893 882 2934 890
rect 2893 856 2908 882
rect 2915 856 2934 882
rect 2998 878 3060 890
rect 3072 878 3147 890
rect 3205 878 3280 890
rect 3292 878 3323 890
rect 3329 878 3364 890
rect 2998 876 3160 878
rect 2893 848 2934 856
rect 3016 852 3029 876
rect 3044 874 3059 876
rect 2856 838 2857 848
rect 2872 838 2885 848
rect 2899 838 2900 848
rect 2915 838 2928 848
rect 2943 838 2973 852
rect 3016 838 3059 852
rect 3083 849 3090 856
rect 3093 852 3160 876
rect 3192 876 3364 878
rect 3162 854 3190 858
rect 3192 854 3272 876
rect 3293 874 3308 876
rect 3162 852 3272 854
rect 3093 848 3272 852
rect 3066 838 3096 848
rect 3098 838 3251 848
rect 3259 838 3289 848
rect 3293 838 3323 852
rect 3351 838 3364 876
rect 3436 882 3471 890
rect 3436 856 3437 882
rect 3444 856 3471 882
rect 3379 838 3409 852
rect 3436 848 3471 856
rect 3473 882 3514 890
rect 3473 856 3488 882
rect 3495 856 3514 882
rect 3578 878 3640 890
rect 3652 878 3727 890
rect 3785 878 3860 890
rect 3872 878 3903 890
rect 3909 878 3944 890
rect 3578 876 3740 878
rect 3473 848 3514 856
rect 3596 852 3609 876
rect 3624 874 3639 876
rect 3436 838 3437 848
rect 3452 838 3465 848
rect 3479 838 3480 848
rect 3495 838 3508 848
rect 3523 838 3553 852
rect 3596 838 3639 852
rect 3663 849 3670 856
rect 3673 852 3740 876
rect 3772 876 3944 878
rect 3742 854 3770 858
rect 3772 854 3852 876
rect 3873 874 3888 876
rect 3742 852 3852 854
rect 3673 848 3852 852
rect 3646 838 3676 848
rect 3678 838 3831 848
rect 3839 838 3869 848
rect 3873 838 3903 852
rect 3931 838 3944 876
rect 4016 882 4051 890
rect 4016 856 4017 882
rect 4024 856 4051 882
rect 3959 838 3989 852
rect 4016 848 4051 856
rect 4053 882 4094 890
rect 4053 856 4068 882
rect 4075 856 4094 882
rect 4158 878 4220 890
rect 4232 878 4307 890
rect 4365 878 4440 890
rect 4452 878 4483 890
rect 4489 878 4524 890
rect 4158 876 4320 878
rect 4053 848 4094 856
rect 4176 852 4189 876
rect 4204 874 4219 876
rect 4016 838 4017 848
rect 4032 838 4045 848
rect 4059 838 4060 848
rect 4075 838 4088 848
rect 4103 838 4133 852
rect 4176 838 4219 852
rect 4243 849 4250 856
rect 4253 852 4320 876
rect 4352 876 4524 878
rect 4322 854 4350 858
rect 4352 854 4432 876
rect 4453 874 4468 876
rect 4322 852 4432 854
rect 4253 848 4432 852
rect 4226 838 4256 848
rect 4258 838 4411 848
rect 4419 838 4449 848
rect 4453 838 4483 852
rect 4511 838 4524 876
rect 4596 882 4631 890
rect 4596 856 4597 882
rect 4604 856 4631 882
rect 4539 838 4569 852
rect 4596 848 4631 856
rect 4633 882 4674 890
rect 4633 856 4648 882
rect 4655 856 4674 882
rect 4738 878 4800 890
rect 4812 878 4887 890
rect 4945 878 5020 890
rect 5032 878 5063 890
rect 5069 878 5104 890
rect 4738 876 4900 878
rect 4633 848 4674 856
rect 4756 852 4769 876
rect 4784 874 4799 876
rect 4596 838 4597 848
rect 4612 838 4625 848
rect 4639 838 4640 848
rect 4655 838 4668 848
rect 4683 838 4713 852
rect 4756 838 4799 852
rect 4823 849 4830 856
rect 4833 852 4900 876
rect 4932 876 5104 878
rect 4902 854 4930 858
rect 4932 854 5012 876
rect 5033 874 5048 876
rect 4902 852 5012 854
rect 4833 848 5012 852
rect 4806 838 4836 848
rect 4838 838 4991 848
rect 4999 838 5029 848
rect 5033 838 5063 852
rect 5091 838 5104 876
rect 5176 882 5211 890
rect 5176 856 5177 882
rect 5184 856 5211 882
rect 5119 838 5149 852
rect 5176 848 5211 856
rect 5213 882 5254 890
rect 5213 856 5228 882
rect 5235 856 5254 882
rect 5318 878 5380 890
rect 5392 878 5467 890
rect 5525 878 5600 890
rect 5612 878 5643 890
rect 5649 878 5684 890
rect 5318 876 5480 878
rect 5213 848 5254 856
rect 5336 852 5349 876
rect 5364 874 5379 876
rect 5176 838 5177 848
rect 5192 838 5205 848
rect 5219 838 5220 848
rect 5235 838 5248 848
rect 5263 838 5293 852
rect 5336 838 5379 852
rect 5403 849 5410 856
rect 5413 852 5480 876
rect 5512 876 5684 878
rect 5482 854 5510 858
rect 5512 854 5592 876
rect 5613 874 5628 876
rect 5482 852 5592 854
rect 5413 848 5592 852
rect 5386 838 5416 848
rect 5418 838 5571 848
rect 5579 838 5609 848
rect 5613 838 5643 852
rect 5671 838 5684 876
rect 5756 882 5791 890
rect 5756 856 5757 882
rect 5764 856 5791 882
rect 5699 838 5729 852
rect 5756 848 5791 856
rect 5793 882 5834 890
rect 5793 856 5808 882
rect 5815 856 5834 882
rect 5898 878 5960 890
rect 5972 878 6047 890
rect 6105 878 6180 890
rect 6192 878 6223 890
rect 6229 878 6264 890
rect 5898 876 6060 878
rect 5793 848 5834 856
rect 5916 852 5929 876
rect 5944 874 5959 876
rect 5756 838 5757 848
rect 5772 838 5785 848
rect 5799 838 5800 848
rect 5815 838 5828 848
rect 5843 838 5873 852
rect 5916 838 5959 852
rect 5983 849 5990 856
rect 5993 852 6060 876
rect 6092 876 6264 878
rect 6062 854 6090 858
rect 6092 854 6172 876
rect 6193 874 6208 876
rect 6062 852 6172 854
rect 5993 848 6172 852
rect 5966 838 5996 848
rect 5998 838 6151 848
rect 6159 838 6189 848
rect 6193 838 6223 852
rect 6251 838 6264 876
rect 6336 882 6371 890
rect 6336 856 6337 882
rect 6344 856 6371 882
rect 6279 838 6309 852
rect 6336 848 6371 856
rect 6373 882 6414 890
rect 6373 856 6388 882
rect 6395 856 6414 882
rect 6478 878 6540 890
rect 6552 878 6627 890
rect 6685 878 6760 890
rect 6772 878 6803 890
rect 6809 878 6844 890
rect 6478 876 6640 878
rect 6373 848 6414 856
rect 6496 852 6509 876
rect 6524 874 6539 876
rect 6336 838 6337 848
rect 6352 838 6365 848
rect 6379 838 6380 848
rect 6395 838 6408 848
rect 6423 838 6453 852
rect 6496 838 6539 852
rect 6563 849 6570 856
rect 6573 852 6640 876
rect 6672 876 6844 878
rect 6642 854 6670 858
rect 6672 854 6752 876
rect 6773 874 6788 876
rect 6642 852 6752 854
rect 6573 848 6752 852
rect 6546 838 6576 848
rect 6578 838 6731 848
rect 6739 838 6769 848
rect 6773 838 6803 852
rect 6831 838 6844 876
rect 6916 882 6951 890
rect 6916 856 6917 882
rect 6924 856 6951 882
rect 6859 838 6889 852
rect 6916 848 6951 856
rect 6953 882 6994 890
rect 6953 856 6968 882
rect 6975 856 6994 882
rect 7058 878 7120 890
rect 7132 878 7207 890
rect 7265 878 7340 890
rect 7352 878 7383 890
rect 7389 878 7424 890
rect 7058 876 7220 878
rect 6953 848 6994 856
rect 7076 852 7089 876
rect 7104 874 7119 876
rect 6916 838 6917 848
rect 6932 838 6945 848
rect 6959 838 6960 848
rect 6975 838 6988 848
rect 7003 838 7033 852
rect 7076 838 7119 852
rect 7143 849 7150 856
rect 7153 852 7220 876
rect 7252 876 7424 878
rect 7222 854 7250 858
rect 7252 854 7332 876
rect 7353 874 7368 876
rect 7222 852 7332 854
rect 7153 848 7332 852
rect 7126 838 7156 848
rect 7158 838 7311 848
rect 7319 838 7349 848
rect 7353 838 7383 852
rect 7411 838 7424 876
rect 7496 882 7531 890
rect 7496 856 7497 882
rect 7504 856 7531 882
rect 7439 838 7469 852
rect 7496 848 7531 856
rect 7533 882 7574 890
rect 7533 856 7548 882
rect 7555 856 7574 882
rect 7638 878 7700 890
rect 7712 878 7787 890
rect 7845 878 7920 890
rect 7932 878 7963 890
rect 7969 878 8004 890
rect 7638 876 7800 878
rect 7533 848 7574 856
rect 7656 852 7669 876
rect 7684 874 7699 876
rect 7496 838 7497 848
rect 7512 838 7525 848
rect 7539 838 7540 848
rect 7555 838 7568 848
rect 7583 838 7613 852
rect 7656 838 7699 852
rect 7723 849 7730 856
rect 7733 852 7800 876
rect 7832 876 8004 878
rect 7802 854 7830 858
rect 7832 854 7912 876
rect 7933 874 7948 876
rect 7802 852 7912 854
rect 7733 848 7912 852
rect 7706 838 7736 848
rect 7738 838 7891 848
rect 7899 838 7929 848
rect 7933 838 7963 852
rect 7991 838 8004 876
rect 8076 882 8111 890
rect 8076 856 8077 882
rect 8084 856 8111 882
rect 8019 838 8049 852
rect 8076 848 8111 856
rect 8113 882 8154 890
rect 8113 856 8128 882
rect 8135 856 8154 882
rect 8218 878 8280 890
rect 8292 878 8367 890
rect 8425 878 8500 890
rect 8512 878 8543 890
rect 8549 878 8584 890
rect 8218 876 8380 878
rect 8113 848 8154 856
rect 8236 852 8249 876
rect 8264 874 8279 876
rect 8076 838 8077 848
rect 8092 838 8105 848
rect 8119 838 8120 848
rect 8135 838 8148 848
rect 8163 838 8193 852
rect 8236 838 8279 852
rect 8303 849 8310 856
rect 8313 852 8380 876
rect 8412 876 8584 878
rect 8382 854 8410 858
rect 8412 854 8492 876
rect 8513 874 8528 876
rect 8382 852 8492 854
rect 8313 848 8492 852
rect 8286 838 8316 848
rect 8318 838 8471 848
rect 8479 838 8509 848
rect 8513 838 8543 852
rect 8571 838 8584 876
rect 8656 882 8691 890
rect 8656 856 8657 882
rect 8664 856 8691 882
rect 8599 838 8629 852
rect 8656 848 8691 856
rect 8693 882 8734 890
rect 8693 856 8708 882
rect 8715 856 8734 882
rect 8798 878 8860 890
rect 8872 878 8947 890
rect 9005 878 9080 890
rect 9092 878 9123 890
rect 9129 878 9164 890
rect 8798 876 8960 878
rect 8693 848 8734 856
rect 8816 852 8829 876
rect 8844 874 8859 876
rect 8656 838 8657 848
rect 8672 838 8685 848
rect 8699 838 8700 848
rect 8715 838 8728 848
rect 8743 838 8773 852
rect 8816 838 8859 852
rect 8883 849 8890 856
rect 8893 852 8960 876
rect 8992 876 9164 878
rect 8962 854 8990 858
rect 8992 854 9072 876
rect 9093 874 9108 876
rect 8962 852 9072 854
rect 8893 848 9072 852
rect 8866 838 8896 848
rect 8898 838 9051 848
rect 9059 838 9089 848
rect 9093 838 9123 852
rect 9151 838 9164 876
rect 9236 882 9271 890
rect 9236 856 9237 882
rect 9244 856 9271 882
rect 9179 838 9209 852
rect 9236 848 9271 856
rect 9236 838 9237 848
rect 9252 838 9265 848
rect -1 832 9265 838
rect 0 824 9265 832
rect 15 794 28 824
rect 43 806 73 824
rect 116 810 130 824
rect 166 810 386 824
rect 117 808 130 810
rect 83 796 98 808
rect 80 794 102 796
rect 107 794 137 808
rect 198 806 351 810
rect 180 794 372 806
rect 415 794 445 808
rect 451 794 464 824
rect 479 806 509 824
rect 552 794 565 824
rect 595 794 608 824
rect 623 806 653 824
rect 696 810 710 824
rect 746 810 966 824
rect 697 808 710 810
rect 663 796 678 808
rect 660 794 682 796
rect 687 794 717 808
rect 778 806 931 810
rect 760 794 952 806
rect 995 794 1025 808
rect 1031 794 1044 824
rect 1059 806 1089 824
rect 1132 794 1145 824
rect 1175 794 1188 824
rect 1203 806 1233 824
rect 1276 810 1290 824
rect 1326 810 1546 824
rect 1277 808 1290 810
rect 1243 796 1258 808
rect 1240 794 1262 796
rect 1267 794 1297 808
rect 1358 806 1511 810
rect 1340 794 1532 806
rect 1575 794 1605 808
rect 1611 794 1624 824
rect 1639 806 1669 824
rect 1712 794 1725 824
rect 1755 794 1768 824
rect 1783 806 1813 824
rect 1856 810 1870 824
rect 1906 810 2126 824
rect 1857 808 1870 810
rect 1823 796 1838 808
rect 1820 794 1842 796
rect 1847 794 1877 808
rect 1938 806 2091 810
rect 1920 794 2112 806
rect 2155 794 2185 808
rect 2191 794 2204 824
rect 2219 806 2249 824
rect 2292 794 2305 824
rect 2335 794 2348 824
rect 2363 806 2393 824
rect 2436 810 2450 824
rect 2486 810 2706 824
rect 2437 808 2450 810
rect 2403 796 2418 808
rect 2400 794 2422 796
rect 2427 794 2457 808
rect 2518 806 2671 810
rect 2500 794 2692 806
rect 2735 794 2765 808
rect 2771 794 2784 824
rect 2799 806 2829 824
rect 2872 794 2885 824
rect 2915 794 2928 824
rect 2943 806 2973 824
rect 3016 810 3030 824
rect 3066 810 3286 824
rect 3017 808 3030 810
rect 2983 796 2998 808
rect 2980 794 3002 796
rect 3007 794 3037 808
rect 3098 806 3251 810
rect 3080 794 3272 806
rect 3315 794 3345 808
rect 3351 794 3364 824
rect 3379 806 3409 824
rect 3452 794 3465 824
rect 3495 794 3508 824
rect 3523 806 3553 824
rect 3596 810 3610 824
rect 3646 810 3866 824
rect 3597 808 3610 810
rect 3563 796 3578 808
rect 3560 794 3582 796
rect 3587 794 3617 808
rect 3678 806 3831 810
rect 3660 794 3852 806
rect 3895 794 3925 808
rect 3931 794 3944 824
rect 3959 806 3989 824
rect 4032 794 4045 824
rect 4075 794 4088 824
rect 4103 806 4133 824
rect 4176 810 4190 824
rect 4226 810 4446 824
rect 4177 808 4190 810
rect 4143 796 4158 808
rect 4140 794 4162 796
rect 4167 794 4197 808
rect 4258 806 4411 810
rect 4240 794 4432 806
rect 4475 794 4505 808
rect 4511 794 4524 824
rect 4539 806 4569 824
rect 4612 794 4625 824
rect 4655 794 4668 824
rect 4683 806 4713 824
rect 4756 810 4770 824
rect 4806 810 5026 824
rect 4757 808 4770 810
rect 4723 796 4738 808
rect 4720 794 4742 796
rect 4747 794 4777 808
rect 4838 806 4991 810
rect 4820 794 5012 806
rect 5055 794 5085 808
rect 5091 794 5104 824
rect 5119 806 5149 824
rect 5192 794 5205 824
rect 5235 794 5248 824
rect 5263 806 5293 824
rect 5336 810 5350 824
rect 5386 810 5606 824
rect 5337 808 5350 810
rect 5303 796 5318 808
rect 5300 794 5322 796
rect 5327 794 5357 808
rect 5418 806 5571 810
rect 5400 794 5592 806
rect 5635 794 5665 808
rect 5671 794 5684 824
rect 5699 806 5729 824
rect 5772 794 5785 824
rect 5815 794 5828 824
rect 5843 806 5873 824
rect 5916 810 5930 824
rect 5966 810 6186 824
rect 5917 808 5930 810
rect 5883 796 5898 808
rect 5880 794 5902 796
rect 5907 794 5937 808
rect 5998 806 6151 810
rect 5980 794 6172 806
rect 6215 794 6245 808
rect 6251 794 6264 824
rect 6279 806 6309 824
rect 6352 794 6365 824
rect 6395 794 6408 824
rect 6423 806 6453 824
rect 6496 810 6510 824
rect 6546 810 6766 824
rect 6497 808 6510 810
rect 6463 796 6478 808
rect 6460 794 6482 796
rect 6487 794 6517 808
rect 6578 806 6731 810
rect 6560 794 6752 806
rect 6795 794 6825 808
rect 6831 794 6844 824
rect 6859 806 6889 824
rect 6932 794 6945 824
rect 6975 794 6988 824
rect 7003 806 7033 824
rect 7076 810 7090 824
rect 7126 810 7346 824
rect 7077 808 7090 810
rect 7043 796 7058 808
rect 7040 794 7062 796
rect 7067 794 7097 808
rect 7158 806 7311 810
rect 7140 794 7332 806
rect 7375 794 7405 808
rect 7411 794 7424 824
rect 7439 806 7469 824
rect 7512 794 7525 824
rect 7555 794 7568 824
rect 7583 806 7613 824
rect 7656 810 7670 824
rect 7706 810 7926 824
rect 7657 808 7670 810
rect 7623 796 7638 808
rect 7620 794 7642 796
rect 7647 794 7677 808
rect 7738 806 7891 810
rect 7720 794 7912 806
rect 7955 794 7985 808
rect 7991 794 8004 824
rect 8019 806 8049 824
rect 8092 794 8105 824
rect 8135 794 8148 824
rect 8163 806 8193 824
rect 8236 810 8250 824
rect 8286 810 8506 824
rect 8237 808 8250 810
rect 8203 796 8218 808
rect 8200 794 8222 796
rect 8227 794 8257 808
rect 8318 806 8471 810
rect 8300 794 8492 806
rect 8535 794 8565 808
rect 8571 794 8584 824
rect 8599 806 8629 824
rect 8672 794 8685 824
rect 8715 794 8728 824
rect 8743 806 8773 824
rect 8816 810 8830 824
rect 8866 810 9086 824
rect 8817 808 8830 810
rect 8783 796 8798 808
rect 8780 794 8802 796
rect 8807 794 8837 808
rect 8898 806 9051 810
rect 8880 794 9072 806
rect 9115 794 9145 808
rect 9151 794 9164 824
rect 9179 806 9209 824
rect 9252 794 9265 824
rect 0 780 9265 794
rect 15 676 28 780
rect 73 758 74 768
rect 89 758 102 768
rect 73 754 102 758
rect 107 754 137 780
rect 155 766 171 768
rect 243 766 296 780
rect 244 764 308 766
rect 351 764 366 780
rect 415 777 445 780
rect 415 774 451 777
rect 381 766 397 768
rect 155 754 170 758
rect 73 752 170 754
rect 198 752 366 764
rect 382 754 397 758
rect 415 755 454 774
rect 473 768 480 769
rect 479 761 480 768
rect 463 758 464 761
rect 479 758 492 761
rect 415 754 445 755
rect 454 754 460 755
rect 463 754 492 758
rect 382 753 492 754
rect 382 752 498 753
rect 57 744 108 752
rect 57 732 82 744
rect 89 732 108 744
rect 139 744 189 752
rect 139 736 155 744
rect 162 742 189 744
rect 198 742 419 752
rect 162 732 419 742
rect 448 744 498 752
rect 448 735 464 744
rect 57 724 108 732
rect 155 724 419 732
rect 445 732 464 735
rect 471 732 498 744
rect 445 724 498 732
rect 73 716 74 724
rect 89 716 102 724
rect 73 708 89 716
rect 70 701 89 704
rect 70 692 92 701
rect 43 682 92 692
rect 43 676 73 682
rect 92 677 97 682
rect 15 660 89 676
rect 107 668 137 724
rect 172 714 380 724
rect 415 720 460 724
rect 463 723 464 724
rect 479 723 492 724
rect 198 684 387 714
rect 213 681 387 684
rect 206 678 387 681
rect 15 658 28 660
rect 43 658 77 660
rect 15 642 89 658
rect 116 654 129 668
rect 144 654 160 670
rect 206 665 217 678
rect -1 620 0 636
rect 15 620 28 642
rect 43 620 73 642
rect 116 638 178 654
rect 206 647 217 663
rect 222 658 232 678
rect 242 658 256 678
rect 259 665 268 678
rect 284 665 293 678
rect 222 647 256 658
rect 259 647 268 663
rect 284 647 293 663
rect 300 658 310 678
rect 320 658 334 678
rect 335 665 346 678
rect 300 647 334 658
rect 335 647 346 663
rect 392 654 408 670
rect 415 668 445 720
rect 479 716 480 723
rect 464 708 480 716
rect 451 676 464 695
rect 479 676 509 692
rect 451 660 525 676
rect 451 658 464 660
rect 479 658 513 660
rect 116 636 129 638
rect 144 636 178 638
rect 116 620 178 636
rect 222 631 238 634
rect 300 631 330 642
rect 378 638 424 654
rect 451 642 525 658
rect 378 636 412 638
rect 377 620 424 636
rect 451 620 464 642
rect 479 620 509 642
rect 536 620 537 636
rect 552 620 565 780
rect 595 676 608 780
rect 653 758 654 768
rect 669 758 682 768
rect 653 754 682 758
rect 687 754 717 780
rect 735 766 751 768
rect 823 766 876 780
rect 824 764 888 766
rect 931 764 946 780
rect 995 777 1025 780
rect 995 774 1031 777
rect 961 766 977 768
rect 735 754 750 758
rect 653 752 750 754
rect 778 752 946 764
rect 962 754 977 758
rect 995 755 1034 774
rect 1053 768 1060 769
rect 1059 761 1060 768
rect 1043 758 1044 761
rect 1059 758 1072 761
rect 995 754 1025 755
rect 1034 754 1040 755
rect 1043 754 1072 758
rect 962 753 1072 754
rect 962 752 1078 753
rect 637 744 688 752
rect 637 732 662 744
rect 669 732 688 744
rect 719 744 769 752
rect 719 736 735 744
rect 742 742 769 744
rect 778 742 999 752
rect 742 732 999 742
rect 1028 744 1078 752
rect 1028 735 1044 744
rect 637 724 688 732
rect 735 724 999 732
rect 1025 732 1044 735
rect 1051 732 1078 744
rect 1025 724 1078 732
rect 653 716 654 724
rect 669 716 682 724
rect 653 708 669 716
rect 650 701 669 704
rect 650 692 672 701
rect 623 682 672 692
rect 623 676 653 682
rect 672 677 677 682
rect 595 660 669 676
rect 687 668 717 724
rect 752 714 960 724
rect 995 720 1040 724
rect 1043 723 1044 724
rect 1059 723 1072 724
rect 778 684 967 714
rect 793 681 967 684
rect 786 678 967 681
rect 595 658 608 660
rect 623 658 657 660
rect 595 642 669 658
rect 696 654 709 668
rect 724 654 740 670
rect 786 665 797 678
rect 579 620 580 636
rect 595 620 608 642
rect 623 620 653 642
rect 696 638 758 654
rect 786 647 797 663
rect 802 658 812 678
rect 822 658 836 678
rect 839 665 848 678
rect 864 665 873 678
rect 802 647 836 658
rect 839 647 848 663
rect 864 647 873 663
rect 880 658 890 678
rect 900 658 914 678
rect 915 665 926 678
rect 880 647 914 658
rect 915 647 926 663
rect 972 654 988 670
rect 995 668 1025 720
rect 1059 716 1060 723
rect 1044 708 1060 716
rect 1031 676 1044 695
rect 1059 676 1089 692
rect 1031 660 1105 676
rect 1031 658 1044 660
rect 1059 658 1093 660
rect 696 636 709 638
rect 724 636 758 638
rect 696 620 758 636
rect 802 631 818 634
rect 880 631 910 642
rect 958 638 1004 654
rect 1031 642 1105 658
rect 958 636 992 638
rect 957 620 1004 636
rect 1031 620 1044 642
rect 1059 620 1089 642
rect 1116 620 1117 636
rect 1132 620 1145 780
rect 1175 676 1188 780
rect 1233 758 1234 768
rect 1249 758 1262 768
rect 1233 754 1262 758
rect 1267 754 1297 780
rect 1315 766 1331 768
rect 1403 766 1456 780
rect 1404 764 1468 766
rect 1511 764 1526 780
rect 1575 777 1605 780
rect 1575 774 1611 777
rect 1541 766 1557 768
rect 1315 754 1330 758
rect 1233 752 1330 754
rect 1358 752 1526 764
rect 1542 754 1557 758
rect 1575 755 1614 774
rect 1633 768 1640 769
rect 1639 761 1640 768
rect 1623 758 1624 761
rect 1639 758 1652 761
rect 1575 754 1605 755
rect 1614 754 1620 755
rect 1623 754 1652 758
rect 1542 753 1652 754
rect 1542 752 1658 753
rect 1217 744 1268 752
rect 1217 732 1242 744
rect 1249 732 1268 744
rect 1299 744 1349 752
rect 1299 736 1315 744
rect 1322 742 1349 744
rect 1358 742 1579 752
rect 1322 732 1579 742
rect 1608 744 1658 752
rect 1608 735 1624 744
rect 1217 724 1268 732
rect 1315 724 1579 732
rect 1605 732 1624 735
rect 1631 732 1658 744
rect 1605 724 1658 732
rect 1233 716 1234 724
rect 1249 716 1262 724
rect 1233 708 1249 716
rect 1230 701 1249 704
rect 1230 692 1252 701
rect 1203 682 1252 692
rect 1203 676 1233 682
rect 1252 677 1257 682
rect 1175 660 1249 676
rect 1267 668 1297 724
rect 1332 714 1540 724
rect 1575 720 1620 724
rect 1623 723 1624 724
rect 1639 723 1652 724
rect 1358 684 1547 714
rect 1373 681 1547 684
rect 1366 678 1547 681
rect 1175 658 1188 660
rect 1203 658 1237 660
rect 1175 642 1249 658
rect 1276 654 1289 668
rect 1304 654 1320 670
rect 1366 665 1377 678
rect 1159 620 1160 636
rect 1175 620 1188 642
rect 1203 620 1233 642
rect 1276 638 1338 654
rect 1366 647 1377 663
rect 1382 658 1392 678
rect 1402 658 1416 678
rect 1419 665 1428 678
rect 1444 665 1453 678
rect 1382 647 1416 658
rect 1419 647 1428 663
rect 1444 647 1453 663
rect 1460 658 1470 678
rect 1480 658 1494 678
rect 1495 665 1506 678
rect 1460 647 1494 658
rect 1495 647 1506 663
rect 1552 654 1568 670
rect 1575 668 1605 720
rect 1639 716 1640 723
rect 1624 708 1640 716
rect 1611 676 1624 695
rect 1639 676 1669 692
rect 1611 660 1685 676
rect 1611 658 1624 660
rect 1639 658 1673 660
rect 1276 636 1289 638
rect 1304 636 1338 638
rect 1276 620 1338 636
rect 1382 631 1398 634
rect 1460 631 1490 642
rect 1538 638 1584 654
rect 1611 642 1685 658
rect 1538 636 1572 638
rect 1537 620 1584 636
rect 1611 620 1624 642
rect 1639 620 1669 642
rect 1696 620 1697 636
rect 1712 620 1725 780
rect 1755 676 1768 780
rect 1813 758 1814 768
rect 1829 758 1842 768
rect 1813 754 1842 758
rect 1847 754 1877 780
rect 1895 766 1911 768
rect 1983 766 2036 780
rect 1984 764 2048 766
rect 2091 764 2106 780
rect 2155 777 2185 780
rect 2155 774 2191 777
rect 2121 766 2137 768
rect 1895 754 1910 758
rect 1813 752 1910 754
rect 1938 752 2106 764
rect 2122 754 2137 758
rect 2155 755 2194 774
rect 2213 768 2220 769
rect 2219 761 2220 768
rect 2203 758 2204 761
rect 2219 758 2232 761
rect 2155 754 2185 755
rect 2194 754 2200 755
rect 2203 754 2232 758
rect 2122 753 2232 754
rect 2122 752 2238 753
rect 1797 744 1848 752
rect 1797 732 1822 744
rect 1829 732 1848 744
rect 1879 744 1929 752
rect 1879 736 1895 744
rect 1902 742 1929 744
rect 1938 742 2159 752
rect 1902 732 2159 742
rect 2188 744 2238 752
rect 2188 735 2204 744
rect 1797 724 1848 732
rect 1895 724 2159 732
rect 2185 732 2204 735
rect 2211 732 2238 744
rect 2185 724 2238 732
rect 1813 716 1814 724
rect 1829 716 1842 724
rect 1813 708 1829 716
rect 1810 701 1829 704
rect 1810 692 1832 701
rect 1783 682 1832 692
rect 1783 676 1813 682
rect 1832 677 1837 682
rect 1755 660 1829 676
rect 1847 668 1877 724
rect 1912 714 2120 724
rect 2155 720 2200 724
rect 2203 723 2204 724
rect 2219 723 2232 724
rect 1938 684 2127 714
rect 1953 681 2127 684
rect 1946 678 2127 681
rect 1755 658 1768 660
rect 1783 658 1817 660
rect 1755 642 1829 658
rect 1856 654 1869 668
rect 1884 654 1900 670
rect 1946 665 1957 678
rect 1739 620 1740 636
rect 1755 620 1768 642
rect 1783 620 1813 642
rect 1856 638 1918 654
rect 1946 647 1957 663
rect 1962 658 1972 678
rect 1982 658 1996 678
rect 1999 665 2008 678
rect 2024 665 2033 678
rect 1962 647 1996 658
rect 1999 647 2008 663
rect 2024 647 2033 663
rect 2040 658 2050 678
rect 2060 658 2074 678
rect 2075 665 2086 678
rect 2040 647 2074 658
rect 2075 647 2086 663
rect 2132 654 2148 670
rect 2155 668 2185 720
rect 2219 716 2220 723
rect 2204 708 2220 716
rect 2191 676 2204 695
rect 2219 676 2249 692
rect 2191 660 2265 676
rect 2191 658 2204 660
rect 2219 658 2253 660
rect 1856 636 1869 638
rect 1884 636 1918 638
rect 1856 620 1918 636
rect 1962 631 1977 634
rect 2040 631 2070 642
rect 2118 638 2164 654
rect 2191 642 2265 658
rect 2118 636 2152 638
rect 2117 620 2164 636
rect 2191 620 2204 642
rect 2219 620 2249 642
rect 2276 620 2277 636
rect 2292 620 2305 780
rect 2335 676 2348 780
rect 2393 758 2394 768
rect 2409 758 2422 768
rect 2393 754 2422 758
rect 2427 754 2457 780
rect 2475 766 2491 768
rect 2563 766 2616 780
rect 2564 764 2628 766
rect 2671 764 2686 780
rect 2735 777 2765 780
rect 2735 774 2771 777
rect 2701 766 2717 768
rect 2475 754 2490 758
rect 2393 752 2490 754
rect 2518 752 2686 764
rect 2702 754 2717 758
rect 2735 755 2774 774
rect 2793 768 2800 769
rect 2799 761 2800 768
rect 2783 758 2784 761
rect 2799 758 2812 761
rect 2735 754 2765 755
rect 2774 754 2780 755
rect 2783 754 2812 758
rect 2702 753 2812 754
rect 2702 752 2818 753
rect 2377 744 2428 752
rect 2377 732 2402 744
rect 2409 732 2428 744
rect 2459 744 2509 752
rect 2459 736 2475 744
rect 2482 742 2509 744
rect 2518 742 2739 752
rect 2482 732 2739 742
rect 2768 744 2818 752
rect 2768 735 2784 744
rect 2377 724 2428 732
rect 2475 724 2739 732
rect 2765 732 2784 735
rect 2791 732 2818 744
rect 2765 724 2818 732
rect 2393 716 2394 724
rect 2409 716 2422 724
rect 2393 708 2409 716
rect 2390 701 2409 704
rect 2390 692 2412 701
rect 2363 682 2412 692
rect 2363 676 2393 682
rect 2412 677 2417 682
rect 2335 660 2409 676
rect 2427 668 2457 724
rect 2492 714 2700 724
rect 2735 720 2780 724
rect 2783 723 2784 724
rect 2799 723 2812 724
rect 2518 684 2707 714
rect 2533 681 2707 684
rect 2526 678 2707 681
rect 2335 658 2348 660
rect 2363 658 2397 660
rect 2335 642 2409 658
rect 2436 654 2449 668
rect 2464 654 2480 670
rect 2526 665 2537 678
rect 2319 620 2320 636
rect 2335 620 2348 642
rect 2363 620 2393 642
rect 2436 638 2498 654
rect 2526 647 2537 663
rect 2542 658 2552 678
rect 2562 658 2576 678
rect 2579 665 2588 678
rect 2604 665 2613 678
rect 2542 647 2576 658
rect 2579 647 2588 663
rect 2604 647 2613 663
rect 2620 658 2630 678
rect 2640 658 2654 678
rect 2655 665 2666 678
rect 2620 647 2654 658
rect 2655 647 2666 663
rect 2712 654 2728 670
rect 2735 668 2765 720
rect 2799 716 2800 723
rect 2784 708 2800 716
rect 2771 676 2784 695
rect 2799 676 2829 692
rect 2771 660 2845 676
rect 2771 658 2784 660
rect 2799 658 2833 660
rect 2436 636 2449 638
rect 2464 636 2498 638
rect 2436 620 2498 636
rect 2542 631 2558 634
rect 2620 631 2650 642
rect 2698 638 2744 654
rect 2771 642 2845 658
rect 2698 636 2732 638
rect 2697 620 2744 636
rect 2771 620 2784 642
rect 2799 620 2829 642
rect 2856 620 2857 636
rect 2872 620 2885 780
rect 2915 676 2928 780
rect 2973 758 2974 768
rect 2989 758 3002 768
rect 2973 754 3002 758
rect 3007 754 3037 780
rect 3055 766 3071 768
rect 3143 766 3196 780
rect 3144 764 3208 766
rect 3251 764 3266 780
rect 3315 777 3345 780
rect 3315 774 3351 777
rect 3281 766 3297 768
rect 3055 754 3070 758
rect 2973 752 3070 754
rect 3098 752 3266 764
rect 3282 754 3297 758
rect 3315 755 3354 774
rect 3373 768 3380 769
rect 3379 761 3380 768
rect 3363 758 3364 761
rect 3379 758 3392 761
rect 3315 754 3345 755
rect 3354 754 3360 755
rect 3363 754 3392 758
rect 3282 753 3392 754
rect 3282 752 3398 753
rect 2957 744 3008 752
rect 2957 732 2982 744
rect 2989 732 3008 744
rect 3039 744 3089 752
rect 3039 736 3055 744
rect 3062 742 3089 744
rect 3098 742 3319 752
rect 3062 732 3319 742
rect 3348 744 3398 752
rect 3348 735 3364 744
rect 2957 724 3008 732
rect 3055 724 3319 732
rect 3345 732 3364 735
rect 3371 732 3398 744
rect 3345 724 3398 732
rect 2973 716 2974 724
rect 2989 716 3002 724
rect 2973 708 2989 716
rect 2970 701 2989 704
rect 2970 692 2992 701
rect 2943 682 2992 692
rect 2943 676 2973 682
rect 2992 677 2997 682
rect 2915 660 2989 676
rect 3007 668 3037 724
rect 3072 714 3280 724
rect 3315 720 3360 724
rect 3363 723 3364 724
rect 3379 723 3392 724
rect 3098 684 3287 714
rect 3113 681 3287 684
rect 3106 678 3287 681
rect 2915 658 2928 660
rect 2943 658 2977 660
rect 2915 642 2989 658
rect 3016 654 3029 668
rect 3044 654 3060 670
rect 3106 665 3117 678
rect 2899 620 2900 636
rect 2915 620 2928 642
rect 2943 620 2973 642
rect 3016 638 3078 654
rect 3106 647 3117 663
rect 3122 658 3132 678
rect 3142 658 3156 678
rect 3159 665 3168 678
rect 3184 665 3193 678
rect 3122 647 3156 658
rect 3159 647 3168 663
rect 3184 647 3193 663
rect 3200 658 3210 678
rect 3220 658 3234 678
rect 3235 665 3246 678
rect 3200 647 3234 658
rect 3235 647 3246 663
rect 3292 654 3308 670
rect 3315 668 3345 720
rect 3379 716 3380 723
rect 3364 708 3380 716
rect 3351 676 3364 695
rect 3379 676 3409 692
rect 3351 660 3425 676
rect 3351 658 3364 660
rect 3379 658 3413 660
rect 3016 636 3029 638
rect 3044 636 3078 638
rect 3016 620 3078 636
rect 3122 631 3138 634
rect 3200 631 3230 642
rect 3278 638 3324 654
rect 3351 642 3425 658
rect 3278 636 3312 638
rect 3277 620 3324 636
rect 3351 620 3364 642
rect 3379 620 3409 642
rect 3436 620 3437 636
rect 3452 620 3465 780
rect 3495 676 3508 780
rect 3553 758 3554 768
rect 3569 758 3582 768
rect 3553 754 3582 758
rect 3587 754 3617 780
rect 3635 766 3651 768
rect 3723 766 3776 780
rect 3724 764 3788 766
rect 3831 764 3846 780
rect 3895 777 3925 780
rect 3895 774 3931 777
rect 3861 766 3877 768
rect 3635 754 3650 758
rect 3553 752 3650 754
rect 3678 752 3846 764
rect 3862 754 3877 758
rect 3895 755 3934 774
rect 3953 768 3960 769
rect 3959 761 3960 768
rect 3943 758 3944 761
rect 3959 758 3972 761
rect 3895 754 3925 755
rect 3934 754 3940 755
rect 3943 754 3972 758
rect 3862 753 3972 754
rect 3862 752 3978 753
rect 3537 744 3588 752
rect 3537 732 3562 744
rect 3569 732 3588 744
rect 3619 744 3669 752
rect 3619 736 3635 744
rect 3642 742 3669 744
rect 3678 742 3899 752
rect 3642 732 3899 742
rect 3928 744 3978 752
rect 3928 735 3944 744
rect 3537 724 3588 732
rect 3635 724 3899 732
rect 3925 732 3944 735
rect 3951 732 3978 744
rect 3925 724 3978 732
rect 3553 716 3554 724
rect 3569 716 3582 724
rect 3553 708 3569 716
rect 3550 701 3569 704
rect 3550 692 3572 701
rect 3523 682 3572 692
rect 3523 676 3553 682
rect 3572 677 3577 682
rect 3495 660 3569 676
rect 3587 668 3617 724
rect 3652 714 3860 724
rect 3895 720 3940 724
rect 3943 723 3944 724
rect 3959 723 3972 724
rect 3678 684 3867 714
rect 3693 681 3867 684
rect 3686 678 3867 681
rect 3495 658 3508 660
rect 3523 658 3557 660
rect 3495 642 3569 658
rect 3596 654 3609 668
rect 3624 654 3640 670
rect 3686 665 3697 678
rect 3479 620 3480 636
rect 3495 620 3508 642
rect 3523 620 3553 642
rect 3596 638 3658 654
rect 3686 647 3697 663
rect 3702 658 3712 678
rect 3722 658 3736 678
rect 3739 665 3748 678
rect 3764 665 3773 678
rect 3702 647 3736 658
rect 3739 647 3748 663
rect 3764 647 3773 663
rect 3780 658 3790 678
rect 3800 658 3814 678
rect 3815 665 3826 678
rect 3780 647 3814 658
rect 3815 647 3826 663
rect 3872 654 3888 670
rect 3895 668 3925 720
rect 3959 716 3960 723
rect 3944 708 3960 716
rect 3931 676 3944 695
rect 3959 676 3989 692
rect 3931 660 4005 676
rect 3931 658 3944 660
rect 3959 658 3993 660
rect 3596 636 3609 638
rect 3624 636 3658 638
rect 3596 620 3658 636
rect 3702 631 3718 634
rect 3780 631 3810 642
rect 3858 638 3904 654
rect 3931 642 4005 658
rect 3858 636 3892 638
rect 3857 620 3904 636
rect 3931 620 3944 642
rect 3959 620 3989 642
rect 4016 620 4017 636
rect 4032 620 4045 780
rect 4075 676 4088 780
rect 4133 758 4134 768
rect 4149 758 4162 768
rect 4133 754 4162 758
rect 4167 754 4197 780
rect 4215 766 4231 768
rect 4303 766 4356 780
rect 4304 764 4368 766
rect 4411 764 4426 780
rect 4475 777 4505 780
rect 4475 774 4511 777
rect 4441 766 4457 768
rect 4215 754 4230 758
rect 4133 752 4230 754
rect 4258 752 4426 764
rect 4442 754 4457 758
rect 4475 755 4514 774
rect 4533 768 4540 769
rect 4539 761 4540 768
rect 4523 758 4524 761
rect 4539 758 4552 761
rect 4475 754 4505 755
rect 4514 754 4520 755
rect 4523 754 4552 758
rect 4442 753 4552 754
rect 4442 752 4558 753
rect 4117 744 4168 752
rect 4117 732 4142 744
rect 4149 732 4168 744
rect 4199 744 4249 752
rect 4199 736 4215 744
rect 4222 742 4249 744
rect 4258 742 4479 752
rect 4222 732 4479 742
rect 4508 744 4558 752
rect 4508 735 4524 744
rect 4117 724 4168 732
rect 4215 724 4479 732
rect 4505 732 4524 735
rect 4531 732 4558 744
rect 4505 724 4558 732
rect 4133 716 4134 724
rect 4149 716 4162 724
rect 4133 708 4149 716
rect 4130 701 4149 704
rect 4130 692 4152 701
rect 4103 682 4152 692
rect 4103 676 4133 682
rect 4152 677 4157 682
rect 4075 660 4149 676
rect 4167 668 4197 724
rect 4232 714 4440 724
rect 4475 720 4520 724
rect 4523 723 4524 724
rect 4539 723 4552 724
rect 4258 684 4447 714
rect 4273 681 4447 684
rect 4266 678 4447 681
rect 4075 658 4088 660
rect 4103 658 4137 660
rect 4075 642 4149 658
rect 4176 654 4189 668
rect 4204 654 4220 670
rect 4266 665 4277 678
rect 4059 620 4060 636
rect 4075 620 4088 642
rect 4103 620 4133 642
rect 4176 638 4238 654
rect 4266 647 4277 663
rect 4282 658 4292 678
rect 4302 658 4316 678
rect 4319 665 4328 678
rect 4344 665 4353 678
rect 4282 647 4316 658
rect 4319 647 4328 663
rect 4344 647 4353 663
rect 4360 658 4370 678
rect 4380 658 4394 678
rect 4395 665 4406 678
rect 4360 647 4394 658
rect 4395 647 4406 663
rect 4452 654 4468 670
rect 4475 668 4505 720
rect 4539 716 4540 723
rect 4524 708 4540 716
rect 4511 676 4524 695
rect 4539 676 4569 692
rect 4511 660 4585 676
rect 4511 658 4524 660
rect 4539 658 4573 660
rect 4176 636 4189 638
rect 4204 636 4238 638
rect 4176 620 4238 636
rect 4282 631 4298 634
rect 4360 631 4390 642
rect 4438 638 4484 654
rect 4511 642 4585 658
rect 4438 636 4472 638
rect 4437 620 4484 636
rect 4511 620 4524 642
rect 4539 620 4569 642
rect 4596 620 4597 636
rect 4612 620 4625 780
rect 4655 676 4668 780
rect 4713 758 4714 768
rect 4729 758 4742 768
rect 4713 754 4742 758
rect 4747 754 4777 780
rect 4795 766 4811 768
rect 4883 766 4936 780
rect 4884 764 4948 766
rect 4991 764 5006 780
rect 5055 777 5085 780
rect 5055 774 5091 777
rect 5021 766 5037 768
rect 4795 754 4810 758
rect 4713 752 4810 754
rect 4838 752 5006 764
rect 5022 754 5037 758
rect 5055 755 5094 774
rect 5113 768 5120 769
rect 5119 761 5120 768
rect 5103 758 5104 761
rect 5119 758 5132 761
rect 5055 754 5085 755
rect 5094 754 5100 755
rect 5103 754 5132 758
rect 5022 753 5132 754
rect 5022 752 5138 753
rect 4697 744 4748 752
rect 4697 732 4722 744
rect 4729 732 4748 744
rect 4779 744 4829 752
rect 4779 736 4795 744
rect 4802 742 4829 744
rect 4838 742 5059 752
rect 4802 732 5059 742
rect 5088 744 5138 752
rect 5088 735 5104 744
rect 4697 724 4748 732
rect 4795 724 5059 732
rect 5085 732 5104 735
rect 5111 732 5138 744
rect 5085 724 5138 732
rect 4713 716 4714 724
rect 4729 716 4742 724
rect 4713 708 4729 716
rect 4710 701 4729 704
rect 4710 692 4732 701
rect 4683 682 4732 692
rect 4683 676 4713 682
rect 4732 677 4737 682
rect 4655 660 4729 676
rect 4747 668 4777 724
rect 4812 714 5020 724
rect 5055 720 5100 724
rect 5103 723 5104 724
rect 5119 723 5132 724
rect 4838 684 5027 714
rect 4853 681 5027 684
rect 4846 678 5027 681
rect 4655 658 4668 660
rect 4683 658 4717 660
rect 4655 642 4729 658
rect 4756 654 4769 668
rect 4784 654 4800 670
rect 4846 665 4857 678
rect 4639 620 4640 636
rect 4655 620 4668 642
rect 4683 620 4713 642
rect 4756 638 4818 654
rect 4846 647 4857 663
rect 4862 658 4872 678
rect 4882 658 4896 678
rect 4899 665 4908 678
rect 4924 665 4933 678
rect 4862 647 4896 658
rect 4899 647 4908 663
rect 4924 647 4933 663
rect 4940 658 4950 678
rect 4960 658 4974 678
rect 4975 665 4986 678
rect 4940 647 4974 658
rect 4975 647 4986 663
rect 5032 654 5048 670
rect 5055 668 5085 720
rect 5119 716 5120 723
rect 5104 708 5120 716
rect 5091 676 5104 695
rect 5119 676 5149 692
rect 5091 660 5165 676
rect 5091 658 5104 660
rect 5119 658 5153 660
rect 4756 636 4769 638
rect 4784 636 4818 638
rect 4756 620 4818 636
rect 4862 631 4878 634
rect 4940 631 4970 642
rect 5018 638 5064 654
rect 5091 642 5165 658
rect 5018 636 5052 638
rect 5017 620 5064 636
rect 5091 620 5104 642
rect 5119 620 5149 642
rect 5176 620 5177 636
rect 5192 620 5205 780
rect 5235 676 5248 780
rect 5293 758 5294 768
rect 5309 758 5322 768
rect 5293 754 5322 758
rect 5327 754 5357 780
rect 5375 766 5391 768
rect 5463 766 5516 780
rect 5464 764 5528 766
rect 5571 764 5586 780
rect 5635 777 5665 780
rect 5635 774 5671 777
rect 5601 766 5617 768
rect 5375 754 5390 758
rect 5293 752 5390 754
rect 5418 752 5586 764
rect 5602 754 5617 758
rect 5635 755 5674 774
rect 5693 768 5700 769
rect 5699 761 5700 768
rect 5683 758 5684 761
rect 5699 758 5712 761
rect 5635 754 5665 755
rect 5674 754 5680 755
rect 5683 754 5712 758
rect 5602 753 5712 754
rect 5602 752 5718 753
rect 5277 744 5328 752
rect 5277 732 5302 744
rect 5309 732 5328 744
rect 5359 744 5409 752
rect 5359 736 5375 744
rect 5382 742 5409 744
rect 5418 742 5639 752
rect 5382 732 5639 742
rect 5668 744 5718 752
rect 5668 735 5684 744
rect 5277 724 5328 732
rect 5375 724 5639 732
rect 5665 732 5684 735
rect 5691 732 5718 744
rect 5665 724 5718 732
rect 5293 716 5294 724
rect 5309 716 5322 724
rect 5293 708 5309 716
rect 5290 701 5309 704
rect 5290 692 5312 701
rect 5263 682 5312 692
rect 5263 676 5293 682
rect 5312 677 5317 682
rect 5235 660 5309 676
rect 5327 668 5357 724
rect 5392 714 5600 724
rect 5635 720 5680 724
rect 5683 723 5684 724
rect 5699 723 5712 724
rect 5418 684 5607 714
rect 5433 681 5607 684
rect 5426 678 5607 681
rect 5235 658 5248 660
rect 5263 658 5297 660
rect 5235 642 5309 658
rect 5336 654 5349 668
rect 5364 654 5380 670
rect 5426 665 5437 678
rect 5219 620 5220 636
rect 5235 620 5248 642
rect 5263 620 5293 642
rect 5336 638 5398 654
rect 5426 647 5437 663
rect 5442 658 5452 678
rect 5462 658 5476 678
rect 5479 665 5488 678
rect 5504 665 5513 678
rect 5442 647 5476 658
rect 5479 647 5488 663
rect 5504 647 5513 663
rect 5520 658 5530 678
rect 5540 658 5554 678
rect 5555 665 5566 678
rect 5520 647 5554 658
rect 5555 647 5566 663
rect 5612 654 5628 670
rect 5635 668 5665 720
rect 5699 716 5700 723
rect 5684 708 5700 716
rect 5671 676 5684 695
rect 5699 676 5729 692
rect 5671 660 5745 676
rect 5671 658 5684 660
rect 5699 658 5733 660
rect 5336 636 5349 638
rect 5364 636 5398 638
rect 5336 620 5398 636
rect 5442 631 5458 634
rect 5520 631 5550 642
rect 5598 638 5644 654
rect 5671 642 5745 658
rect 5598 636 5632 638
rect 5597 620 5644 636
rect 5671 620 5684 642
rect 5699 620 5729 642
rect 5756 620 5757 636
rect 5772 620 5785 780
rect 5815 676 5828 780
rect 5873 758 5874 768
rect 5889 758 5902 768
rect 5873 754 5902 758
rect 5907 754 5937 780
rect 5955 766 5971 768
rect 6043 766 6096 780
rect 6044 764 6108 766
rect 6151 764 6166 780
rect 6215 777 6245 780
rect 6215 774 6251 777
rect 6181 766 6197 768
rect 5955 754 5970 758
rect 5873 752 5970 754
rect 5998 752 6166 764
rect 6182 754 6197 758
rect 6215 755 6254 774
rect 6273 768 6280 769
rect 6279 761 6280 768
rect 6263 758 6264 761
rect 6279 758 6292 761
rect 6215 754 6245 755
rect 6254 754 6260 755
rect 6263 754 6292 758
rect 6182 753 6292 754
rect 6182 752 6298 753
rect 5857 744 5908 752
rect 5857 732 5882 744
rect 5889 732 5908 744
rect 5939 744 5989 752
rect 5939 736 5955 744
rect 5962 742 5989 744
rect 5998 742 6219 752
rect 5962 732 6219 742
rect 6248 744 6298 752
rect 6248 735 6264 744
rect 5857 724 5908 732
rect 5955 724 6219 732
rect 6245 732 6264 735
rect 6271 732 6298 744
rect 6245 724 6298 732
rect 5873 716 5874 724
rect 5889 716 5902 724
rect 5873 708 5889 716
rect 5870 701 5889 704
rect 5870 692 5892 701
rect 5843 682 5892 692
rect 5843 676 5873 682
rect 5892 677 5897 682
rect 5815 660 5889 676
rect 5907 668 5937 724
rect 5972 714 6180 724
rect 6215 720 6260 724
rect 6263 723 6264 724
rect 6279 723 6292 724
rect 5998 684 6187 714
rect 6013 681 6187 684
rect 6006 678 6187 681
rect 5815 658 5828 660
rect 5843 658 5877 660
rect 5815 642 5889 658
rect 5916 654 5929 668
rect 5944 654 5960 670
rect 6006 665 6017 678
rect 5799 620 5800 636
rect 5815 620 5828 642
rect 5843 620 5873 642
rect 5916 638 5978 654
rect 6006 647 6017 663
rect 6022 658 6032 678
rect 6042 658 6056 678
rect 6059 665 6068 678
rect 6084 665 6093 678
rect 6022 647 6056 658
rect 6059 647 6068 663
rect 6084 647 6093 663
rect 6100 658 6110 678
rect 6120 658 6134 678
rect 6135 665 6146 678
rect 6100 647 6134 658
rect 6135 647 6146 663
rect 6192 654 6208 670
rect 6215 668 6245 720
rect 6279 716 6280 723
rect 6264 708 6280 716
rect 6251 676 6264 695
rect 6279 676 6309 692
rect 6251 660 6325 676
rect 6251 658 6264 660
rect 6279 658 6313 660
rect 5916 636 5929 638
rect 5944 636 5978 638
rect 5916 620 5978 636
rect 6022 631 6038 634
rect 6100 631 6130 642
rect 6178 638 6224 654
rect 6251 642 6325 658
rect 6178 636 6212 638
rect 6177 620 6224 636
rect 6251 620 6264 642
rect 6279 620 6309 642
rect 6336 620 6337 636
rect 6352 620 6365 780
rect 6395 676 6408 780
rect 6453 758 6454 768
rect 6469 758 6482 768
rect 6453 754 6482 758
rect 6487 754 6517 780
rect 6535 766 6551 768
rect 6623 766 6676 780
rect 6624 764 6688 766
rect 6731 764 6746 780
rect 6795 777 6825 780
rect 6795 774 6831 777
rect 6761 766 6777 768
rect 6535 754 6550 758
rect 6453 752 6550 754
rect 6578 752 6746 764
rect 6762 754 6777 758
rect 6795 755 6834 774
rect 6853 768 6860 769
rect 6859 761 6860 768
rect 6843 758 6844 761
rect 6859 758 6872 761
rect 6795 754 6825 755
rect 6834 754 6840 755
rect 6843 754 6872 758
rect 6762 753 6872 754
rect 6762 752 6878 753
rect 6437 744 6488 752
rect 6437 732 6462 744
rect 6469 732 6488 744
rect 6519 744 6569 752
rect 6519 736 6535 744
rect 6542 742 6569 744
rect 6578 742 6799 752
rect 6542 732 6799 742
rect 6828 744 6878 752
rect 6828 735 6844 744
rect 6437 724 6488 732
rect 6535 724 6799 732
rect 6825 732 6844 735
rect 6851 732 6878 744
rect 6825 724 6878 732
rect 6453 716 6454 724
rect 6469 716 6482 724
rect 6453 708 6469 716
rect 6450 701 6469 704
rect 6450 692 6472 701
rect 6423 682 6472 692
rect 6423 676 6453 682
rect 6472 677 6477 682
rect 6395 660 6469 676
rect 6487 668 6517 724
rect 6552 714 6760 724
rect 6795 720 6840 724
rect 6843 723 6844 724
rect 6859 723 6872 724
rect 6578 684 6767 714
rect 6593 681 6767 684
rect 6586 678 6767 681
rect 6395 658 6408 660
rect 6423 658 6457 660
rect 6395 642 6469 658
rect 6496 654 6509 668
rect 6524 654 6540 670
rect 6586 665 6597 678
rect 6379 620 6380 636
rect 6395 620 6408 642
rect 6423 620 6453 642
rect 6496 638 6558 654
rect 6586 647 6597 663
rect 6602 658 6612 678
rect 6622 658 6636 678
rect 6639 665 6648 678
rect 6664 665 6673 678
rect 6602 647 6636 658
rect 6639 647 6648 663
rect 6664 647 6673 663
rect 6680 658 6690 678
rect 6700 658 6714 678
rect 6715 665 6726 678
rect 6680 647 6714 658
rect 6715 647 6726 663
rect 6772 654 6788 670
rect 6795 668 6825 720
rect 6859 716 6860 723
rect 6844 708 6860 716
rect 6831 676 6844 695
rect 6859 676 6889 692
rect 6831 660 6905 676
rect 6831 658 6844 660
rect 6859 658 6893 660
rect 6496 636 6509 638
rect 6524 636 6558 638
rect 6496 620 6558 636
rect 6602 631 6618 634
rect 6680 631 6710 642
rect 6758 638 6804 654
rect 6831 642 6905 658
rect 6758 636 6792 638
rect 6757 620 6804 636
rect 6831 620 6844 642
rect 6859 620 6889 642
rect 6916 620 6917 636
rect 6932 620 6945 780
rect 6975 676 6988 780
rect 7033 758 7034 768
rect 7049 758 7062 768
rect 7033 754 7062 758
rect 7067 754 7097 780
rect 7115 766 7131 768
rect 7203 766 7256 780
rect 7204 764 7268 766
rect 7311 764 7326 780
rect 7375 777 7405 780
rect 7375 774 7411 777
rect 7341 766 7357 768
rect 7115 754 7130 758
rect 7033 752 7130 754
rect 7158 752 7326 764
rect 7342 754 7357 758
rect 7375 755 7414 774
rect 7433 768 7440 769
rect 7439 761 7440 768
rect 7423 758 7424 761
rect 7439 758 7452 761
rect 7375 754 7405 755
rect 7414 754 7420 755
rect 7423 754 7452 758
rect 7342 753 7452 754
rect 7342 752 7458 753
rect 7017 744 7068 752
rect 7017 732 7042 744
rect 7049 732 7068 744
rect 7099 744 7149 752
rect 7099 736 7115 744
rect 7122 742 7149 744
rect 7158 742 7379 752
rect 7122 732 7379 742
rect 7408 744 7458 752
rect 7408 735 7424 744
rect 7017 724 7068 732
rect 7115 724 7379 732
rect 7405 732 7424 735
rect 7431 732 7458 744
rect 7405 724 7458 732
rect 7033 716 7034 724
rect 7049 716 7062 724
rect 7033 708 7049 716
rect 7030 701 7049 704
rect 7030 692 7052 701
rect 7003 682 7052 692
rect 7003 676 7033 682
rect 7052 677 7057 682
rect 6975 660 7049 676
rect 7067 668 7097 724
rect 7132 714 7340 724
rect 7375 720 7420 724
rect 7423 723 7424 724
rect 7439 723 7452 724
rect 7158 684 7347 714
rect 7173 681 7347 684
rect 7166 678 7347 681
rect 6975 658 6988 660
rect 7003 658 7037 660
rect 6975 642 7049 658
rect 7076 654 7089 668
rect 7104 654 7120 670
rect 7166 665 7177 678
rect 6959 620 6960 636
rect 6975 620 6988 642
rect 7003 620 7033 642
rect 7076 638 7138 654
rect 7166 647 7177 663
rect 7182 658 7192 678
rect 7202 658 7216 678
rect 7219 665 7228 678
rect 7244 665 7253 678
rect 7182 647 7216 658
rect 7219 647 7228 663
rect 7244 647 7253 663
rect 7260 658 7270 678
rect 7280 658 7294 678
rect 7295 665 7306 678
rect 7260 647 7294 658
rect 7295 647 7306 663
rect 7352 654 7368 670
rect 7375 668 7405 720
rect 7439 716 7440 723
rect 7424 708 7440 716
rect 7411 676 7424 695
rect 7439 676 7469 692
rect 7411 660 7485 676
rect 7411 658 7424 660
rect 7439 658 7473 660
rect 7076 636 7089 638
rect 7104 636 7138 638
rect 7076 620 7138 636
rect 7182 631 7198 634
rect 7260 631 7290 642
rect 7338 638 7384 654
rect 7411 642 7485 658
rect 7338 636 7372 638
rect 7337 620 7384 636
rect 7411 620 7424 642
rect 7439 620 7469 642
rect 7496 620 7497 636
rect 7512 620 7525 780
rect 7555 676 7568 780
rect 7613 758 7614 768
rect 7629 758 7642 768
rect 7613 754 7642 758
rect 7647 754 7677 780
rect 7695 766 7711 768
rect 7783 766 7836 780
rect 7784 764 7848 766
rect 7891 764 7906 780
rect 7955 777 7985 780
rect 7955 774 7991 777
rect 7921 766 7937 768
rect 7695 754 7710 758
rect 7613 752 7710 754
rect 7738 752 7906 764
rect 7922 754 7937 758
rect 7955 755 7994 774
rect 8013 768 8020 769
rect 8019 761 8020 768
rect 8003 758 8004 761
rect 8019 758 8032 761
rect 7955 754 7985 755
rect 7994 754 8000 755
rect 8003 754 8032 758
rect 7922 753 8032 754
rect 7922 752 8038 753
rect 7597 744 7648 752
rect 7597 732 7622 744
rect 7629 732 7648 744
rect 7679 744 7729 752
rect 7679 736 7695 744
rect 7702 742 7729 744
rect 7738 742 7959 752
rect 7702 732 7959 742
rect 7988 744 8038 752
rect 7988 735 8004 744
rect 7597 724 7648 732
rect 7695 724 7959 732
rect 7985 732 8004 735
rect 8011 732 8038 744
rect 7985 724 8038 732
rect 7613 716 7614 724
rect 7629 716 7642 724
rect 7613 708 7629 716
rect 7610 701 7629 704
rect 7610 692 7632 701
rect 7583 682 7632 692
rect 7583 676 7613 682
rect 7632 677 7637 682
rect 7555 660 7629 676
rect 7647 668 7677 724
rect 7712 714 7920 724
rect 7955 720 8000 724
rect 8003 723 8004 724
rect 8019 723 8032 724
rect 7738 684 7927 714
rect 7753 681 7927 684
rect 7746 678 7927 681
rect 7555 658 7568 660
rect 7583 658 7617 660
rect 7555 642 7629 658
rect 7656 654 7669 668
rect 7684 654 7700 670
rect 7746 665 7757 678
rect 7539 620 7540 636
rect 7555 620 7568 642
rect 7583 620 7613 642
rect 7656 638 7718 654
rect 7746 647 7757 663
rect 7762 658 7772 678
rect 7782 658 7796 678
rect 7799 665 7808 678
rect 7824 665 7833 678
rect 7762 647 7796 658
rect 7799 647 7808 663
rect 7824 647 7833 663
rect 7840 658 7850 678
rect 7860 658 7874 678
rect 7875 665 7886 678
rect 7840 647 7874 658
rect 7875 647 7886 663
rect 7932 654 7948 670
rect 7955 668 7985 720
rect 8019 716 8020 723
rect 8004 708 8020 716
rect 7991 676 8004 695
rect 8019 676 8049 692
rect 7991 660 8065 676
rect 7991 658 8004 660
rect 8019 658 8053 660
rect 7656 636 7669 638
rect 7684 636 7718 638
rect 7656 620 7718 636
rect 7762 631 7778 634
rect 7840 631 7870 642
rect 7918 638 7964 654
rect 7991 642 8065 658
rect 7918 636 7952 638
rect 7917 620 7964 636
rect 7991 620 8004 642
rect 8019 620 8049 642
rect 8076 620 8077 636
rect 8092 620 8105 780
rect 8135 676 8148 780
rect 8193 758 8194 768
rect 8209 758 8222 768
rect 8193 754 8222 758
rect 8227 754 8257 780
rect 8275 766 8291 768
rect 8363 766 8416 780
rect 8364 764 8428 766
rect 8471 764 8486 780
rect 8535 777 8565 780
rect 8535 774 8571 777
rect 8501 766 8517 768
rect 8275 754 8290 758
rect 8193 752 8290 754
rect 8318 752 8486 764
rect 8502 754 8517 758
rect 8535 755 8574 774
rect 8593 768 8600 769
rect 8599 761 8600 768
rect 8583 758 8584 761
rect 8599 758 8612 761
rect 8535 754 8565 755
rect 8574 754 8580 755
rect 8583 754 8612 758
rect 8502 753 8612 754
rect 8502 752 8618 753
rect 8177 744 8228 752
rect 8177 732 8202 744
rect 8209 732 8228 744
rect 8259 744 8309 752
rect 8259 736 8275 744
rect 8282 742 8309 744
rect 8318 742 8539 752
rect 8282 732 8539 742
rect 8568 744 8618 752
rect 8568 735 8584 744
rect 8177 724 8228 732
rect 8275 724 8539 732
rect 8565 732 8584 735
rect 8591 732 8618 744
rect 8565 724 8618 732
rect 8193 716 8194 724
rect 8209 716 8222 724
rect 8193 708 8209 716
rect 8190 701 8209 704
rect 8190 692 8212 701
rect 8163 682 8212 692
rect 8163 676 8193 682
rect 8212 677 8217 682
rect 8135 660 8209 676
rect 8227 668 8257 724
rect 8292 714 8500 724
rect 8535 720 8580 724
rect 8583 723 8584 724
rect 8599 723 8612 724
rect 8318 684 8507 714
rect 8333 681 8507 684
rect 8326 678 8507 681
rect 8135 658 8148 660
rect 8163 658 8197 660
rect 8135 642 8209 658
rect 8236 654 8249 668
rect 8264 654 8280 670
rect 8326 665 8337 678
rect 8119 620 8120 636
rect 8135 620 8148 642
rect 8163 620 8193 642
rect 8236 638 8298 654
rect 8326 647 8337 663
rect 8342 658 8352 678
rect 8362 658 8376 678
rect 8379 665 8388 678
rect 8404 665 8413 678
rect 8342 647 8376 658
rect 8379 647 8388 663
rect 8404 647 8413 663
rect 8420 658 8430 678
rect 8440 658 8454 678
rect 8455 665 8466 678
rect 8420 647 8454 658
rect 8455 647 8466 663
rect 8512 654 8528 670
rect 8535 668 8565 720
rect 8599 716 8600 723
rect 8584 708 8600 716
rect 8571 676 8584 695
rect 8599 676 8629 692
rect 8571 660 8645 676
rect 8571 658 8584 660
rect 8599 658 8633 660
rect 8236 636 8249 638
rect 8264 636 8298 638
rect 8236 620 8298 636
rect 8342 631 8358 634
rect 8420 631 8450 642
rect 8498 638 8544 654
rect 8571 642 8645 658
rect 8498 636 8532 638
rect 8497 620 8544 636
rect 8571 620 8584 642
rect 8599 620 8629 642
rect 8656 620 8657 636
rect 8672 620 8685 780
rect 8715 676 8728 780
rect 8773 758 8774 768
rect 8789 758 8802 768
rect 8773 754 8802 758
rect 8807 754 8837 780
rect 8855 766 8871 768
rect 8943 766 8996 780
rect 8944 764 9008 766
rect 9051 764 9066 780
rect 9115 777 9145 780
rect 9115 774 9151 777
rect 9081 766 9097 768
rect 8855 754 8870 758
rect 8773 752 8870 754
rect 8898 752 9066 764
rect 9082 754 9097 758
rect 9115 755 9154 774
rect 9173 768 9180 769
rect 9179 761 9180 768
rect 9163 758 9164 761
rect 9179 758 9192 761
rect 9115 754 9145 755
rect 9154 754 9160 755
rect 9163 754 9192 758
rect 9082 753 9192 754
rect 9082 752 9198 753
rect 8757 744 8808 752
rect 8757 732 8782 744
rect 8789 732 8808 744
rect 8839 744 8889 752
rect 8839 736 8855 744
rect 8862 742 8889 744
rect 8898 742 9119 752
rect 8862 732 9119 742
rect 9148 744 9198 752
rect 9148 735 9164 744
rect 8757 724 8808 732
rect 8855 724 9119 732
rect 9145 732 9164 735
rect 9171 732 9198 744
rect 9145 724 9198 732
rect 8773 716 8774 724
rect 8789 716 8802 724
rect 8773 708 8789 716
rect 8770 701 8789 704
rect 8770 692 8792 701
rect 8743 682 8792 692
rect 8743 676 8773 682
rect 8792 677 8797 682
rect 8715 660 8789 676
rect 8807 668 8837 724
rect 8872 714 9080 724
rect 9115 720 9160 724
rect 9163 723 9164 724
rect 9179 723 9192 724
rect 8898 684 9087 714
rect 8913 681 9087 684
rect 8906 678 9087 681
rect 8715 658 8728 660
rect 8743 658 8777 660
rect 8715 642 8789 658
rect 8816 654 8829 668
rect 8844 654 8860 670
rect 8906 665 8917 678
rect 8699 620 8700 636
rect 8715 620 8728 642
rect 8743 620 8773 642
rect 8816 638 8878 654
rect 8906 647 8917 663
rect 8922 658 8932 678
rect 8942 658 8956 678
rect 8959 665 8968 678
rect 8984 665 8993 678
rect 8922 647 8956 658
rect 8959 647 8968 663
rect 8984 647 8993 663
rect 9000 658 9010 678
rect 9020 658 9034 678
rect 9035 665 9046 678
rect 9000 647 9034 658
rect 9035 647 9046 663
rect 9092 654 9108 670
rect 9115 668 9145 720
rect 9179 716 9180 723
rect 9164 708 9180 716
rect 9151 676 9164 695
rect 9179 676 9209 692
rect 9151 660 9225 676
rect 9151 658 9164 660
rect 9179 658 9213 660
rect 8816 636 8829 638
rect 8844 636 8878 638
rect 8816 620 8878 636
rect 8922 631 8938 634
rect 9000 631 9030 642
rect 9078 638 9124 654
rect 9151 642 9225 658
rect 9078 636 9112 638
rect 9077 620 9124 636
rect 9151 620 9164 642
rect 9179 620 9209 642
rect 9236 620 9237 636
rect 9252 620 9265 780
rect -7 612 34 620
rect -7 586 8 612
rect 15 586 34 612
rect 98 608 160 620
rect 172 608 247 620
rect 305 608 380 620
rect 392 608 423 620
rect 429 608 464 620
rect 98 606 260 608
rect -7 578 34 586
rect 116 582 129 606
rect 144 604 159 606
rect -1 568 0 578
rect 15 568 28 578
rect 43 568 73 582
rect 116 568 159 582
rect 183 579 190 586
rect 193 582 260 606
rect 292 606 464 608
rect 262 584 290 588
rect 292 584 372 606
rect 393 604 408 606
rect 262 582 372 584
rect 193 578 372 582
rect 166 568 196 578
rect 198 568 351 578
rect 359 568 389 578
rect 393 568 423 582
rect 451 568 464 606
rect 536 612 571 620
rect 536 586 537 612
rect 544 586 571 612
rect 479 568 509 582
rect 536 578 571 586
rect 573 612 614 620
rect 573 586 588 612
rect 595 586 614 612
rect 678 608 740 620
rect 752 608 827 620
rect 885 608 960 620
rect 972 608 1003 620
rect 1009 608 1044 620
rect 678 606 840 608
rect 573 578 614 586
rect 696 582 709 606
rect 724 604 739 606
rect 536 568 537 578
rect 552 568 565 578
rect 579 568 580 578
rect 595 568 608 578
rect 623 568 653 582
rect 696 568 739 582
rect 763 579 770 586
rect 773 582 840 606
rect 872 606 1044 608
rect 842 584 870 588
rect 872 584 952 606
rect 973 604 988 606
rect 842 582 952 584
rect 773 578 952 582
rect 746 568 776 578
rect 778 568 931 578
rect 939 568 969 578
rect 973 568 1003 582
rect 1031 568 1044 606
rect 1116 612 1151 620
rect 1116 586 1117 612
rect 1124 586 1151 612
rect 1059 568 1089 582
rect 1116 578 1151 586
rect 1153 612 1194 620
rect 1153 586 1168 612
rect 1175 586 1194 612
rect 1258 608 1320 620
rect 1332 608 1407 620
rect 1465 608 1540 620
rect 1552 608 1583 620
rect 1589 608 1624 620
rect 1258 606 1420 608
rect 1153 578 1194 586
rect 1276 582 1289 606
rect 1304 604 1319 606
rect 1116 568 1117 578
rect 1132 568 1145 578
rect 1159 568 1160 578
rect 1175 568 1188 578
rect 1203 568 1233 582
rect 1276 568 1319 582
rect 1343 579 1350 586
rect 1353 582 1420 606
rect 1452 606 1624 608
rect 1422 584 1450 588
rect 1452 584 1532 606
rect 1553 604 1568 606
rect 1422 582 1532 584
rect 1353 578 1532 582
rect 1326 568 1356 578
rect 1358 568 1511 578
rect 1519 568 1549 578
rect 1553 568 1583 582
rect 1611 568 1624 606
rect 1696 612 1731 620
rect 1696 586 1697 612
rect 1704 586 1731 612
rect 1639 568 1669 582
rect 1696 578 1731 586
rect 1733 612 1774 620
rect 1733 586 1748 612
rect 1755 586 1774 612
rect 1838 608 1900 620
rect 1912 608 1987 620
rect 2045 608 2120 620
rect 2132 608 2163 620
rect 2169 608 2204 620
rect 1838 606 2000 608
rect 1733 578 1774 586
rect 1856 582 1869 606
rect 1884 604 1899 606
rect 1696 568 1697 578
rect 1712 568 1725 578
rect 1739 568 1740 578
rect 1755 568 1768 578
rect 1783 568 1813 582
rect 1856 568 1899 582
rect 1923 579 1930 586
rect 1933 582 2000 606
rect 2032 606 2204 608
rect 2002 584 2030 588
rect 2032 584 2112 606
rect 2133 604 2148 606
rect 2002 582 2112 584
rect 1933 578 2112 582
rect 1906 568 1936 578
rect 1938 568 2091 578
rect 2099 568 2129 578
rect 2133 568 2163 582
rect 2191 568 2204 606
rect 2276 612 2311 620
rect 2276 586 2277 612
rect 2284 586 2311 612
rect 2219 568 2249 582
rect 2276 578 2311 586
rect 2313 612 2354 620
rect 2313 586 2328 612
rect 2335 586 2354 612
rect 2418 608 2480 620
rect 2492 608 2567 620
rect 2625 608 2700 620
rect 2712 608 2743 620
rect 2749 608 2784 620
rect 2418 606 2580 608
rect 2313 578 2354 586
rect 2436 582 2449 606
rect 2464 604 2479 606
rect 2276 568 2277 578
rect 2292 568 2305 578
rect 2319 568 2320 578
rect 2335 568 2348 578
rect 2363 568 2393 582
rect 2436 568 2479 582
rect 2503 579 2510 586
rect 2513 582 2580 606
rect 2612 606 2784 608
rect 2582 584 2610 588
rect 2612 584 2692 606
rect 2713 604 2728 606
rect 2582 582 2692 584
rect 2513 578 2692 582
rect 2486 568 2516 578
rect 2518 568 2671 578
rect 2679 568 2709 578
rect 2713 568 2743 582
rect 2771 568 2784 606
rect 2856 612 2891 620
rect 2856 586 2857 612
rect 2864 586 2891 612
rect 2799 568 2829 582
rect 2856 578 2891 586
rect 2893 612 2934 620
rect 2893 586 2908 612
rect 2915 586 2934 612
rect 2998 608 3060 620
rect 3072 608 3147 620
rect 3205 608 3280 620
rect 3292 608 3323 620
rect 3329 608 3364 620
rect 2998 606 3160 608
rect 2893 578 2934 586
rect 3016 582 3029 606
rect 3044 604 3059 606
rect 2856 568 2857 578
rect 2872 568 2885 578
rect 2899 568 2900 578
rect 2915 568 2928 578
rect 2943 568 2973 582
rect 3016 568 3059 582
rect 3083 579 3090 586
rect 3093 582 3160 606
rect 3192 606 3364 608
rect 3162 584 3190 588
rect 3192 584 3272 606
rect 3293 604 3308 606
rect 3162 582 3272 584
rect 3093 578 3272 582
rect 3066 568 3096 578
rect 3098 568 3251 578
rect 3259 568 3289 578
rect 3293 568 3323 582
rect 3351 568 3364 606
rect 3436 612 3471 620
rect 3436 586 3437 612
rect 3444 586 3471 612
rect 3379 568 3409 582
rect 3436 578 3471 586
rect 3473 612 3514 620
rect 3473 586 3488 612
rect 3495 586 3514 612
rect 3578 608 3640 620
rect 3652 608 3727 620
rect 3785 608 3860 620
rect 3872 608 3903 620
rect 3909 608 3944 620
rect 3578 606 3740 608
rect 3473 578 3514 586
rect 3596 582 3609 606
rect 3624 604 3639 606
rect 3436 568 3437 578
rect 3452 568 3465 578
rect 3479 568 3480 578
rect 3495 568 3508 578
rect 3523 568 3553 582
rect 3596 568 3639 582
rect 3663 579 3670 586
rect 3673 582 3740 606
rect 3772 606 3944 608
rect 3742 584 3770 588
rect 3772 584 3852 606
rect 3873 604 3888 606
rect 3742 582 3852 584
rect 3673 578 3852 582
rect 3646 568 3676 578
rect 3678 568 3831 578
rect 3839 568 3869 578
rect 3873 568 3903 582
rect 3931 568 3944 606
rect 4016 612 4051 620
rect 4016 586 4017 612
rect 4024 586 4051 612
rect 3959 568 3989 582
rect 4016 578 4051 586
rect 4053 612 4094 620
rect 4053 586 4068 612
rect 4075 586 4094 612
rect 4158 608 4220 620
rect 4232 608 4307 620
rect 4365 608 4440 620
rect 4452 608 4483 620
rect 4489 608 4524 620
rect 4158 606 4320 608
rect 4053 578 4094 586
rect 4176 582 4189 606
rect 4204 604 4219 606
rect 4016 568 4017 578
rect 4032 568 4045 578
rect 4059 568 4060 578
rect 4075 568 4088 578
rect 4103 568 4133 582
rect 4176 568 4219 582
rect 4243 579 4250 586
rect 4253 582 4320 606
rect 4352 606 4524 608
rect 4322 584 4350 588
rect 4352 584 4432 606
rect 4453 604 4468 606
rect 4322 582 4432 584
rect 4253 578 4432 582
rect 4226 568 4256 578
rect 4258 568 4411 578
rect 4419 568 4449 578
rect 4453 568 4483 582
rect 4511 568 4524 606
rect 4596 612 4631 620
rect 4596 586 4597 612
rect 4604 586 4631 612
rect 4539 568 4569 582
rect 4596 578 4631 586
rect 4633 612 4674 620
rect 4633 586 4648 612
rect 4655 586 4674 612
rect 4738 608 4800 620
rect 4812 608 4887 620
rect 4945 608 5020 620
rect 5032 608 5063 620
rect 5069 608 5104 620
rect 4738 606 4900 608
rect 4633 578 4674 586
rect 4756 582 4769 606
rect 4784 604 4799 606
rect 4596 568 4597 578
rect 4612 568 4625 578
rect 4639 568 4640 578
rect 4655 568 4668 578
rect 4683 568 4713 582
rect 4756 568 4799 582
rect 4823 579 4830 586
rect 4833 582 4900 606
rect 4932 606 5104 608
rect 4902 584 4930 588
rect 4932 584 5012 606
rect 5033 604 5048 606
rect 4902 582 5012 584
rect 4833 578 5012 582
rect 4806 568 4836 578
rect 4838 568 4991 578
rect 4999 568 5029 578
rect 5033 568 5063 582
rect 5091 568 5104 606
rect 5176 612 5211 620
rect 5176 586 5177 612
rect 5184 586 5211 612
rect 5119 568 5149 582
rect 5176 578 5211 586
rect 5213 612 5254 620
rect 5213 586 5228 612
rect 5235 586 5254 612
rect 5318 608 5380 620
rect 5392 608 5467 620
rect 5525 608 5600 620
rect 5612 608 5643 620
rect 5649 608 5684 620
rect 5318 606 5480 608
rect 5213 578 5254 586
rect 5336 582 5349 606
rect 5364 604 5379 606
rect 5176 568 5177 578
rect 5192 568 5205 578
rect 5219 568 5220 578
rect 5235 568 5248 578
rect 5263 568 5293 582
rect 5336 568 5379 582
rect 5403 579 5410 586
rect 5413 582 5480 606
rect 5512 606 5684 608
rect 5482 584 5510 588
rect 5512 584 5592 606
rect 5613 604 5628 606
rect 5482 582 5592 584
rect 5413 578 5592 582
rect 5386 568 5416 578
rect 5418 568 5571 578
rect 5579 568 5609 578
rect 5613 568 5643 582
rect 5671 568 5684 606
rect 5756 612 5791 620
rect 5756 586 5757 612
rect 5764 586 5791 612
rect 5699 568 5729 582
rect 5756 578 5791 586
rect 5793 612 5834 620
rect 5793 586 5808 612
rect 5815 586 5834 612
rect 5898 608 5960 620
rect 5972 608 6047 620
rect 6105 608 6180 620
rect 6192 608 6223 620
rect 6229 608 6264 620
rect 5898 606 6060 608
rect 5793 578 5834 586
rect 5916 582 5929 606
rect 5944 604 5959 606
rect 5756 568 5757 578
rect 5772 568 5785 578
rect 5799 568 5800 578
rect 5815 568 5828 578
rect 5843 568 5873 582
rect 5916 568 5959 582
rect 5983 579 5990 586
rect 5993 582 6060 606
rect 6092 606 6264 608
rect 6062 584 6090 588
rect 6092 584 6172 606
rect 6193 604 6208 606
rect 6062 582 6172 584
rect 5993 578 6172 582
rect 5966 568 5996 578
rect 5998 568 6151 578
rect 6159 568 6189 578
rect 6193 568 6223 582
rect 6251 568 6264 606
rect 6336 612 6371 620
rect 6336 586 6337 612
rect 6344 586 6371 612
rect 6279 568 6309 582
rect 6336 578 6371 586
rect 6373 612 6414 620
rect 6373 586 6388 612
rect 6395 586 6414 612
rect 6478 608 6540 620
rect 6552 608 6627 620
rect 6685 608 6760 620
rect 6772 608 6803 620
rect 6809 608 6844 620
rect 6478 606 6640 608
rect 6373 578 6414 586
rect 6496 582 6509 606
rect 6524 604 6539 606
rect 6336 568 6337 578
rect 6352 568 6365 578
rect 6379 568 6380 578
rect 6395 568 6408 578
rect 6423 568 6453 582
rect 6496 568 6539 582
rect 6563 579 6570 586
rect 6573 582 6640 606
rect 6672 606 6844 608
rect 6642 584 6670 588
rect 6672 584 6752 606
rect 6773 604 6788 606
rect 6642 582 6752 584
rect 6573 578 6752 582
rect 6546 568 6576 578
rect 6578 568 6731 578
rect 6739 568 6769 578
rect 6773 568 6803 582
rect 6831 568 6844 606
rect 6916 612 6951 620
rect 6916 586 6917 612
rect 6924 586 6951 612
rect 6859 568 6889 582
rect 6916 578 6951 586
rect 6953 612 6994 620
rect 6953 586 6968 612
rect 6975 586 6994 612
rect 7058 608 7120 620
rect 7132 608 7207 620
rect 7265 608 7340 620
rect 7352 608 7383 620
rect 7389 608 7424 620
rect 7058 606 7220 608
rect 6953 578 6994 586
rect 7076 582 7089 606
rect 7104 604 7119 606
rect 6916 568 6917 578
rect 6932 568 6945 578
rect 6959 568 6960 578
rect 6975 568 6988 578
rect 7003 568 7033 582
rect 7076 568 7119 582
rect 7143 579 7150 586
rect 7153 582 7220 606
rect 7252 606 7424 608
rect 7222 584 7250 588
rect 7252 584 7332 606
rect 7353 604 7368 606
rect 7222 582 7332 584
rect 7153 578 7332 582
rect 7126 568 7156 578
rect 7158 568 7311 578
rect 7319 568 7349 578
rect 7353 568 7383 582
rect 7411 568 7424 606
rect 7496 612 7531 620
rect 7496 586 7497 612
rect 7504 586 7531 612
rect 7439 568 7469 582
rect 7496 578 7531 586
rect 7533 612 7574 620
rect 7533 586 7548 612
rect 7555 586 7574 612
rect 7638 608 7700 620
rect 7712 608 7787 620
rect 7845 608 7920 620
rect 7932 608 7963 620
rect 7969 608 8004 620
rect 7638 606 7800 608
rect 7533 578 7574 586
rect 7656 582 7669 606
rect 7684 604 7699 606
rect 7496 568 7497 578
rect 7512 568 7525 578
rect 7539 568 7540 578
rect 7555 568 7568 578
rect 7583 568 7613 582
rect 7656 568 7699 582
rect 7723 579 7730 586
rect 7733 582 7800 606
rect 7832 606 8004 608
rect 7802 584 7830 588
rect 7832 584 7912 606
rect 7933 604 7948 606
rect 7802 582 7912 584
rect 7733 578 7912 582
rect 7706 568 7736 578
rect 7738 568 7891 578
rect 7899 568 7929 578
rect 7933 568 7963 582
rect 7991 568 8004 606
rect 8076 612 8111 620
rect 8076 586 8077 612
rect 8084 586 8111 612
rect 8019 568 8049 582
rect 8076 578 8111 586
rect 8113 612 8154 620
rect 8113 586 8128 612
rect 8135 586 8154 612
rect 8218 608 8280 620
rect 8292 608 8367 620
rect 8425 608 8500 620
rect 8512 608 8543 620
rect 8549 608 8584 620
rect 8218 606 8380 608
rect 8113 578 8154 586
rect 8236 582 8249 606
rect 8264 604 8279 606
rect 8076 568 8077 578
rect 8092 568 8105 578
rect 8119 568 8120 578
rect 8135 568 8148 578
rect 8163 568 8193 582
rect 8236 568 8279 582
rect 8303 579 8310 586
rect 8313 582 8380 606
rect 8412 606 8584 608
rect 8382 584 8410 588
rect 8412 584 8492 606
rect 8513 604 8528 606
rect 8382 582 8492 584
rect 8313 578 8492 582
rect 8286 568 8316 578
rect 8318 568 8471 578
rect 8479 568 8509 578
rect 8513 568 8543 582
rect 8571 568 8584 606
rect 8656 612 8691 620
rect 8656 586 8657 612
rect 8664 586 8691 612
rect 8599 568 8629 582
rect 8656 578 8691 586
rect 8693 612 8734 620
rect 8693 586 8708 612
rect 8715 586 8734 612
rect 8798 608 8860 620
rect 8872 608 8947 620
rect 9005 608 9080 620
rect 9092 608 9123 620
rect 9129 608 9164 620
rect 8798 606 8960 608
rect 8693 578 8734 586
rect 8816 582 8829 606
rect 8844 604 8859 606
rect 8656 568 8657 578
rect 8672 568 8685 578
rect 8699 568 8700 578
rect 8715 568 8728 578
rect 8743 568 8773 582
rect 8816 568 8859 582
rect 8883 579 8890 586
rect 8893 582 8960 606
rect 8992 606 9164 608
rect 8962 584 8990 588
rect 8992 584 9072 606
rect 9093 604 9108 606
rect 8962 582 9072 584
rect 8893 578 9072 582
rect 8866 568 8896 578
rect 8898 568 9051 578
rect 9059 568 9089 578
rect 9093 568 9123 582
rect 9151 568 9164 606
rect 9236 612 9271 620
rect 9236 586 9237 612
rect 9244 586 9271 612
rect 9179 568 9209 582
rect 9236 578 9271 586
rect 9236 568 9237 578
rect 9252 568 9265 578
rect -1 562 9265 568
rect 0 554 9265 562
rect 15 524 28 554
rect 43 536 73 554
rect 116 540 130 554
rect 166 540 386 554
rect 117 538 130 540
rect 83 526 98 538
rect 80 524 102 526
rect 107 524 137 538
rect 198 536 351 540
rect 180 524 372 536
rect 415 524 445 538
rect 451 524 464 554
rect 479 536 509 554
rect 552 524 565 554
rect 595 524 608 554
rect 623 536 653 554
rect 696 540 710 554
rect 746 540 966 554
rect 697 538 710 540
rect 663 526 678 538
rect 660 524 682 526
rect 687 524 717 538
rect 778 536 931 540
rect 760 524 952 536
rect 995 524 1025 538
rect 1031 524 1044 554
rect 1059 536 1089 554
rect 1132 524 1145 554
rect 1175 524 1188 554
rect 1203 536 1233 554
rect 1276 540 1290 554
rect 1326 540 1546 554
rect 1277 538 1290 540
rect 1243 526 1258 538
rect 1240 524 1262 526
rect 1267 524 1297 538
rect 1358 536 1511 540
rect 1340 524 1532 536
rect 1575 524 1605 538
rect 1611 524 1624 554
rect 1639 536 1669 554
rect 1712 524 1725 554
rect 1755 524 1768 554
rect 1783 536 1813 554
rect 1856 540 1870 554
rect 1906 540 2126 554
rect 1857 538 1870 540
rect 1823 526 1838 538
rect 1820 524 1842 526
rect 1847 524 1877 538
rect 1938 536 2091 540
rect 1920 524 2112 536
rect 2155 524 2185 538
rect 2191 524 2204 554
rect 2219 536 2249 554
rect 2292 524 2305 554
rect 2335 524 2348 554
rect 2363 536 2393 554
rect 2436 540 2450 554
rect 2486 540 2706 554
rect 2437 538 2450 540
rect 2403 526 2418 538
rect 2400 524 2422 526
rect 2427 524 2457 538
rect 2518 536 2671 540
rect 2500 524 2692 536
rect 2735 524 2765 538
rect 2771 524 2784 554
rect 2799 536 2829 554
rect 2872 524 2885 554
rect 2915 524 2928 554
rect 2943 536 2973 554
rect 3016 540 3030 554
rect 3066 540 3286 554
rect 3017 538 3030 540
rect 2983 526 2998 538
rect 2980 524 3002 526
rect 3007 524 3037 538
rect 3098 536 3251 540
rect 3080 524 3272 536
rect 3315 524 3345 538
rect 3351 524 3364 554
rect 3379 536 3409 554
rect 3452 524 3465 554
rect 3495 524 3508 554
rect 3523 536 3553 554
rect 3596 540 3610 554
rect 3646 540 3866 554
rect 3597 538 3610 540
rect 3563 526 3578 538
rect 3560 524 3582 526
rect 3587 524 3617 538
rect 3678 536 3831 540
rect 3660 524 3852 536
rect 3895 524 3925 538
rect 3931 524 3944 554
rect 3959 536 3989 554
rect 4032 524 4045 554
rect 4075 524 4088 554
rect 4103 536 4133 554
rect 4176 540 4190 554
rect 4226 540 4446 554
rect 4177 538 4190 540
rect 4143 526 4158 538
rect 4140 524 4162 526
rect 4167 524 4197 538
rect 4258 536 4411 540
rect 4240 524 4432 536
rect 4475 524 4505 538
rect 4511 524 4524 554
rect 4539 536 4569 554
rect 4612 524 4625 554
rect 4655 524 4668 554
rect 4683 536 4713 554
rect 4756 540 4770 554
rect 4806 540 5026 554
rect 4757 538 4770 540
rect 4723 526 4738 538
rect 4720 524 4742 526
rect 4747 524 4777 538
rect 4838 536 4991 540
rect 4820 524 5012 536
rect 5055 524 5085 538
rect 5091 524 5104 554
rect 5119 536 5149 554
rect 5192 524 5205 554
rect 5235 524 5248 554
rect 5263 536 5293 554
rect 5336 540 5350 554
rect 5386 540 5606 554
rect 5337 538 5350 540
rect 5303 526 5318 538
rect 5300 524 5322 526
rect 5327 524 5357 538
rect 5418 536 5571 540
rect 5400 524 5592 536
rect 5635 524 5665 538
rect 5671 524 5684 554
rect 5699 536 5729 554
rect 5772 524 5785 554
rect 5815 524 5828 554
rect 5843 536 5873 554
rect 5916 540 5930 554
rect 5966 540 6186 554
rect 5917 538 5930 540
rect 5883 526 5898 538
rect 5880 524 5902 526
rect 5907 524 5937 538
rect 5998 536 6151 540
rect 5980 524 6172 536
rect 6215 524 6245 538
rect 6251 524 6264 554
rect 6279 536 6309 554
rect 6352 524 6365 554
rect 6395 524 6408 554
rect 6423 536 6453 554
rect 6496 540 6510 554
rect 6546 540 6766 554
rect 6497 538 6510 540
rect 6463 526 6478 538
rect 6460 524 6482 526
rect 6487 524 6517 538
rect 6578 536 6731 540
rect 6560 524 6752 536
rect 6795 524 6825 538
rect 6831 524 6844 554
rect 6859 536 6889 554
rect 6932 524 6945 554
rect 6975 524 6988 554
rect 7003 536 7033 554
rect 7076 540 7090 554
rect 7126 540 7346 554
rect 7077 538 7090 540
rect 7043 526 7058 538
rect 7040 524 7062 526
rect 7067 524 7097 538
rect 7158 536 7311 540
rect 7140 524 7332 536
rect 7375 524 7405 538
rect 7411 524 7424 554
rect 7439 536 7469 554
rect 7512 524 7525 554
rect 7555 524 7568 554
rect 7583 536 7613 554
rect 7656 540 7670 554
rect 7706 540 7926 554
rect 7657 538 7670 540
rect 7623 526 7638 538
rect 7620 524 7642 526
rect 7647 524 7677 538
rect 7738 536 7891 540
rect 7720 524 7912 536
rect 7955 524 7985 538
rect 7991 524 8004 554
rect 8019 536 8049 554
rect 8092 524 8105 554
rect 8135 524 8148 554
rect 8163 536 8193 554
rect 8236 540 8250 554
rect 8286 540 8506 554
rect 8237 538 8250 540
rect 8203 526 8218 538
rect 8200 524 8222 526
rect 8227 524 8257 538
rect 8318 536 8471 540
rect 8300 524 8492 536
rect 8535 524 8565 538
rect 8571 524 8584 554
rect 8599 536 8629 554
rect 8672 524 8685 554
rect 8715 524 8728 554
rect 8743 536 8773 554
rect 8816 540 8830 554
rect 8866 540 9086 554
rect 8817 538 8830 540
rect 8783 526 8798 538
rect 8780 524 8802 526
rect 8807 524 8837 538
rect 8898 536 9051 540
rect 8880 524 9072 536
rect 9115 524 9145 538
rect 9151 524 9164 554
rect 9179 536 9209 554
rect 9252 524 9265 554
rect 0 510 9265 524
rect 15 406 28 510
rect 73 488 74 498
rect 89 488 102 498
rect 73 484 102 488
rect 107 484 137 510
rect 155 496 171 498
rect 243 496 296 510
rect 244 494 308 496
rect 351 494 366 510
rect 415 507 445 510
rect 415 504 451 507
rect 381 496 397 498
rect 155 484 170 488
rect 73 482 170 484
rect 198 482 366 494
rect 382 484 397 488
rect 415 485 454 504
rect 473 498 480 499
rect 479 491 480 498
rect 463 488 464 491
rect 479 488 492 491
rect 415 484 445 485
rect 454 484 460 485
rect 463 484 492 488
rect 382 483 492 484
rect 382 482 498 483
rect 57 474 108 482
rect 57 462 82 474
rect 89 462 108 474
rect 139 474 189 482
rect 139 466 155 474
rect 162 472 189 474
rect 198 472 419 482
rect 162 462 419 472
rect 448 474 498 482
rect 448 465 464 474
rect 57 454 108 462
rect 155 454 419 462
rect 445 462 464 465
rect 471 462 498 474
rect 445 454 498 462
rect 73 446 74 454
rect 89 446 102 454
rect 73 438 89 446
rect 70 431 89 434
rect 70 422 92 431
rect 43 412 92 422
rect 43 406 73 412
rect 92 407 97 412
rect 15 390 89 406
rect 107 398 137 454
rect 172 444 380 454
rect 415 450 460 454
rect 463 453 464 454
rect 479 453 492 454
rect 198 414 387 444
rect 213 411 387 414
rect 206 408 387 411
rect 15 388 28 390
rect 43 388 77 390
rect 15 372 89 388
rect 116 384 129 398
rect 144 384 160 400
rect 206 395 217 408
rect -1 350 0 366
rect 15 350 28 372
rect 43 350 73 372
rect 116 368 178 384
rect 206 377 217 393
rect 222 388 232 408
rect 242 388 256 408
rect 259 395 268 408
rect 284 395 293 408
rect 222 377 256 388
rect 259 377 268 393
rect 284 377 293 393
rect 300 388 310 408
rect 320 388 334 408
rect 335 395 346 408
rect 300 377 334 388
rect 335 377 346 393
rect 392 384 408 400
rect 415 398 445 450
rect 479 446 480 453
rect 464 438 480 446
rect 451 406 464 425
rect 479 406 509 422
rect 451 390 525 406
rect 451 388 464 390
rect 479 388 513 390
rect 116 366 129 368
rect 144 366 178 368
rect 116 350 178 366
rect 222 361 238 364
rect 300 361 330 372
rect 378 368 424 384
rect 451 372 525 388
rect 378 366 412 368
rect 377 350 424 366
rect 451 350 464 372
rect 479 350 509 372
rect 536 350 537 366
rect 552 350 565 510
rect 595 406 608 510
rect 653 488 654 498
rect 669 488 682 498
rect 653 484 682 488
rect 687 484 717 510
rect 735 496 751 498
rect 823 496 876 510
rect 824 494 888 496
rect 931 494 946 510
rect 995 507 1025 510
rect 995 504 1031 507
rect 961 496 977 498
rect 735 484 750 488
rect 653 482 750 484
rect 778 482 946 494
rect 962 484 977 488
rect 995 485 1034 504
rect 1053 498 1060 499
rect 1059 491 1060 498
rect 1043 488 1044 491
rect 1059 488 1072 491
rect 995 484 1025 485
rect 1034 484 1040 485
rect 1043 484 1072 488
rect 962 483 1072 484
rect 962 482 1078 483
rect 637 474 688 482
rect 637 462 662 474
rect 669 462 688 474
rect 719 474 769 482
rect 719 466 735 474
rect 742 472 769 474
rect 778 472 999 482
rect 742 462 999 472
rect 1028 474 1078 482
rect 1028 465 1044 474
rect 637 454 688 462
rect 735 454 999 462
rect 1025 462 1044 465
rect 1051 462 1078 474
rect 1025 454 1078 462
rect 653 446 654 454
rect 669 446 682 454
rect 653 438 669 446
rect 650 431 669 434
rect 650 422 672 431
rect 623 412 672 422
rect 623 406 653 412
rect 672 407 677 412
rect 595 390 669 406
rect 687 398 717 454
rect 752 444 960 454
rect 995 450 1040 454
rect 1043 453 1044 454
rect 1059 453 1072 454
rect 778 414 967 444
rect 793 411 967 414
rect 786 408 967 411
rect 595 388 608 390
rect 623 388 657 390
rect 595 372 669 388
rect 696 384 709 398
rect 724 384 740 400
rect 786 395 797 408
rect 579 350 580 366
rect 595 350 608 372
rect 623 350 653 372
rect 696 368 758 384
rect 786 377 797 393
rect 802 388 812 408
rect 822 388 836 408
rect 839 395 848 408
rect 864 395 873 408
rect 802 377 836 388
rect 839 377 848 393
rect 864 377 873 393
rect 880 388 890 408
rect 900 388 914 408
rect 915 395 926 408
rect 880 377 914 388
rect 915 377 926 393
rect 972 384 988 400
rect 995 398 1025 450
rect 1059 446 1060 453
rect 1044 438 1060 446
rect 1031 406 1044 425
rect 1059 406 1089 422
rect 1031 390 1105 406
rect 1031 388 1044 390
rect 1059 388 1093 390
rect 696 366 709 368
rect 724 366 758 368
rect 696 350 758 366
rect 802 361 818 364
rect 880 361 910 372
rect 958 368 1004 384
rect 1031 372 1105 388
rect 958 366 992 368
rect 957 350 1004 366
rect 1031 350 1044 372
rect 1059 350 1089 372
rect 1116 350 1117 366
rect 1132 350 1145 510
rect 1175 406 1188 510
rect 1233 488 1234 498
rect 1249 488 1262 498
rect 1233 484 1262 488
rect 1267 484 1297 510
rect 1315 496 1331 498
rect 1403 496 1456 510
rect 1404 494 1468 496
rect 1511 494 1526 510
rect 1575 507 1605 510
rect 1575 504 1611 507
rect 1541 496 1557 498
rect 1315 484 1330 488
rect 1233 482 1330 484
rect 1358 482 1526 494
rect 1542 484 1557 488
rect 1575 485 1614 504
rect 1633 498 1640 499
rect 1639 491 1640 498
rect 1623 488 1624 491
rect 1639 488 1652 491
rect 1575 484 1605 485
rect 1614 484 1620 485
rect 1623 484 1652 488
rect 1542 483 1652 484
rect 1542 482 1658 483
rect 1217 474 1268 482
rect 1217 462 1242 474
rect 1249 462 1268 474
rect 1299 474 1349 482
rect 1299 466 1315 474
rect 1322 472 1349 474
rect 1358 472 1579 482
rect 1322 462 1579 472
rect 1608 474 1658 482
rect 1608 465 1624 474
rect 1217 454 1268 462
rect 1315 454 1579 462
rect 1605 462 1624 465
rect 1631 462 1658 474
rect 1605 454 1658 462
rect 1233 446 1234 454
rect 1249 446 1262 454
rect 1233 438 1249 446
rect 1230 431 1249 434
rect 1230 422 1252 431
rect 1203 412 1252 422
rect 1203 406 1233 412
rect 1252 407 1257 412
rect 1175 390 1249 406
rect 1267 398 1297 454
rect 1332 444 1540 454
rect 1575 450 1620 454
rect 1623 453 1624 454
rect 1639 453 1652 454
rect 1358 414 1547 444
rect 1373 411 1547 414
rect 1366 408 1547 411
rect 1175 388 1188 390
rect 1203 388 1237 390
rect 1175 372 1249 388
rect 1276 384 1289 398
rect 1304 384 1320 400
rect 1366 395 1377 408
rect 1159 350 1160 366
rect 1175 350 1188 372
rect 1203 350 1233 372
rect 1276 368 1338 384
rect 1366 377 1377 393
rect 1382 388 1392 408
rect 1402 388 1416 408
rect 1419 395 1428 408
rect 1444 395 1453 408
rect 1382 377 1416 388
rect 1419 377 1428 393
rect 1444 377 1453 393
rect 1460 388 1470 408
rect 1480 388 1494 408
rect 1495 395 1506 408
rect 1460 377 1494 388
rect 1495 377 1506 393
rect 1552 384 1568 400
rect 1575 398 1605 450
rect 1639 446 1640 453
rect 1624 438 1640 446
rect 1611 406 1624 425
rect 1639 406 1669 422
rect 1611 390 1685 406
rect 1611 388 1624 390
rect 1639 388 1673 390
rect 1276 366 1289 368
rect 1304 366 1338 368
rect 1276 350 1338 366
rect 1382 361 1398 364
rect 1460 361 1490 372
rect 1538 368 1584 384
rect 1611 372 1685 388
rect 1538 366 1572 368
rect 1537 350 1584 366
rect 1611 350 1624 372
rect 1639 350 1669 372
rect 1696 350 1697 366
rect 1712 350 1725 510
rect 1755 406 1768 510
rect 1813 488 1814 498
rect 1829 488 1842 498
rect 1813 484 1842 488
rect 1847 484 1877 510
rect 1895 496 1911 498
rect 1983 496 2036 510
rect 1984 494 2048 496
rect 2091 494 2106 510
rect 2155 507 2185 510
rect 2155 504 2191 507
rect 2121 496 2137 498
rect 1895 484 1910 488
rect 1813 482 1910 484
rect 1938 482 2106 494
rect 2122 484 2137 488
rect 2155 485 2194 504
rect 2213 498 2220 499
rect 2219 491 2220 498
rect 2203 488 2204 491
rect 2219 488 2232 491
rect 2155 484 2185 485
rect 2194 484 2200 485
rect 2203 484 2232 488
rect 2122 483 2232 484
rect 2122 482 2238 483
rect 1797 474 1848 482
rect 1797 462 1822 474
rect 1829 462 1848 474
rect 1879 474 1929 482
rect 1879 466 1895 474
rect 1902 472 1929 474
rect 1938 472 2159 482
rect 1902 462 2159 472
rect 2188 474 2238 482
rect 2188 465 2204 474
rect 1797 454 1848 462
rect 1895 454 2159 462
rect 2185 462 2204 465
rect 2211 462 2238 474
rect 2185 454 2238 462
rect 1813 446 1814 454
rect 1829 446 1842 454
rect 1813 438 1829 446
rect 1810 431 1829 434
rect 1810 422 1832 431
rect 1783 412 1832 422
rect 1783 406 1813 412
rect 1832 407 1837 412
rect 1755 390 1829 406
rect 1847 398 1877 454
rect 1912 444 2120 454
rect 2155 450 2200 454
rect 2203 453 2204 454
rect 2219 453 2232 454
rect 1938 414 2127 444
rect 1953 411 2127 414
rect 1946 408 2127 411
rect 1755 388 1768 390
rect 1783 388 1817 390
rect 1755 372 1829 388
rect 1856 384 1869 398
rect 1884 384 1900 400
rect 1946 395 1957 408
rect 1739 350 1740 366
rect 1755 350 1768 372
rect 1783 350 1813 372
rect 1856 368 1918 384
rect 1946 377 1957 393
rect 1962 388 1972 408
rect 1982 388 1996 408
rect 1999 395 2008 408
rect 2024 395 2033 408
rect 1962 377 1996 388
rect 1999 377 2008 393
rect 2024 377 2033 393
rect 2040 388 2050 408
rect 2060 388 2074 408
rect 2075 395 2086 408
rect 2040 377 2074 388
rect 2075 377 2086 393
rect 2132 384 2148 400
rect 2155 398 2185 450
rect 2219 446 2220 453
rect 2204 438 2220 446
rect 2191 406 2204 425
rect 2219 406 2249 422
rect 2191 390 2265 406
rect 2191 388 2204 390
rect 2219 388 2253 390
rect 1856 366 1869 368
rect 1884 366 1918 368
rect 1856 350 1918 366
rect 1962 361 1977 364
rect 2040 361 2070 372
rect 2118 368 2164 384
rect 2191 372 2265 388
rect 2118 366 2152 368
rect 2117 350 2164 366
rect 2191 350 2204 372
rect 2219 350 2249 372
rect 2276 350 2277 366
rect 2292 350 2305 510
rect 2335 406 2348 510
rect 2393 488 2394 498
rect 2409 488 2422 498
rect 2393 484 2422 488
rect 2427 484 2457 510
rect 2475 496 2491 498
rect 2563 496 2616 510
rect 2564 494 2628 496
rect 2671 494 2686 510
rect 2735 507 2765 510
rect 2735 504 2771 507
rect 2701 496 2717 498
rect 2475 484 2490 488
rect 2393 482 2490 484
rect 2518 482 2686 494
rect 2702 484 2717 488
rect 2735 485 2774 504
rect 2793 498 2800 499
rect 2799 491 2800 498
rect 2783 488 2784 491
rect 2799 488 2812 491
rect 2735 484 2765 485
rect 2774 484 2780 485
rect 2783 484 2812 488
rect 2702 483 2812 484
rect 2702 482 2818 483
rect 2377 474 2428 482
rect 2377 462 2402 474
rect 2409 462 2428 474
rect 2459 474 2509 482
rect 2459 466 2475 474
rect 2482 472 2509 474
rect 2518 472 2739 482
rect 2482 462 2739 472
rect 2768 474 2818 482
rect 2768 465 2784 474
rect 2377 454 2428 462
rect 2475 454 2739 462
rect 2765 462 2784 465
rect 2791 462 2818 474
rect 2765 454 2818 462
rect 2393 446 2394 454
rect 2409 446 2422 454
rect 2393 438 2409 446
rect 2390 431 2409 434
rect 2390 422 2412 431
rect 2363 412 2412 422
rect 2363 406 2393 412
rect 2412 407 2417 412
rect 2335 390 2409 406
rect 2427 398 2457 454
rect 2492 444 2700 454
rect 2735 450 2780 454
rect 2783 453 2784 454
rect 2799 453 2812 454
rect 2518 414 2707 444
rect 2533 411 2707 414
rect 2526 408 2707 411
rect 2335 388 2348 390
rect 2363 388 2397 390
rect 2335 372 2409 388
rect 2436 384 2449 398
rect 2464 384 2480 400
rect 2526 395 2537 408
rect 2319 350 2320 366
rect 2335 350 2348 372
rect 2363 350 2393 372
rect 2436 368 2498 384
rect 2526 377 2537 393
rect 2542 388 2552 408
rect 2562 388 2576 408
rect 2579 395 2588 408
rect 2604 395 2613 408
rect 2542 377 2576 388
rect 2579 377 2588 393
rect 2604 377 2613 393
rect 2620 388 2630 408
rect 2640 388 2654 408
rect 2655 395 2666 408
rect 2620 377 2654 388
rect 2655 377 2666 393
rect 2712 384 2728 400
rect 2735 398 2765 450
rect 2799 446 2800 453
rect 2784 438 2800 446
rect 2771 406 2784 425
rect 2799 406 2829 422
rect 2771 390 2845 406
rect 2771 388 2784 390
rect 2799 388 2833 390
rect 2436 366 2449 368
rect 2464 366 2498 368
rect 2436 350 2498 366
rect 2542 361 2558 364
rect 2620 361 2650 372
rect 2698 368 2744 384
rect 2771 372 2845 388
rect 2698 366 2732 368
rect 2697 350 2744 366
rect 2771 350 2784 372
rect 2799 350 2829 372
rect 2856 350 2857 366
rect 2872 350 2885 510
rect 2915 406 2928 510
rect 2973 488 2974 498
rect 2989 488 3002 498
rect 2973 484 3002 488
rect 3007 484 3037 510
rect 3055 496 3071 498
rect 3143 496 3196 510
rect 3144 494 3208 496
rect 3251 494 3266 510
rect 3315 507 3345 510
rect 3315 504 3351 507
rect 3281 496 3297 498
rect 3055 484 3070 488
rect 2973 482 3070 484
rect 3098 482 3266 494
rect 3282 484 3297 488
rect 3315 485 3354 504
rect 3373 498 3380 499
rect 3379 491 3380 498
rect 3363 488 3364 491
rect 3379 488 3392 491
rect 3315 484 3345 485
rect 3354 484 3360 485
rect 3363 484 3392 488
rect 3282 483 3392 484
rect 3282 482 3398 483
rect 2957 474 3008 482
rect 2957 462 2982 474
rect 2989 462 3008 474
rect 3039 474 3089 482
rect 3039 466 3055 474
rect 3062 472 3089 474
rect 3098 472 3319 482
rect 3062 462 3319 472
rect 3348 474 3398 482
rect 3348 465 3364 474
rect 2957 454 3008 462
rect 3055 454 3319 462
rect 3345 462 3364 465
rect 3371 462 3398 474
rect 3345 454 3398 462
rect 2973 446 2974 454
rect 2989 446 3002 454
rect 2973 438 2989 446
rect 2970 431 2989 434
rect 2970 422 2992 431
rect 2943 412 2992 422
rect 2943 406 2973 412
rect 2992 407 2997 412
rect 2915 390 2989 406
rect 3007 398 3037 454
rect 3072 444 3280 454
rect 3315 450 3360 454
rect 3363 453 3364 454
rect 3379 453 3392 454
rect 3098 414 3287 444
rect 3113 411 3287 414
rect 3106 408 3287 411
rect 2915 388 2928 390
rect 2943 388 2977 390
rect 2915 372 2989 388
rect 3016 384 3029 398
rect 3044 384 3060 400
rect 3106 395 3117 408
rect 2899 350 2900 366
rect 2915 350 2928 372
rect 2943 350 2973 372
rect 3016 368 3078 384
rect 3106 377 3117 393
rect 3122 388 3132 408
rect 3142 388 3156 408
rect 3159 395 3168 408
rect 3184 395 3193 408
rect 3122 377 3156 388
rect 3159 377 3168 393
rect 3184 377 3193 393
rect 3200 388 3210 408
rect 3220 388 3234 408
rect 3235 395 3246 408
rect 3200 377 3234 388
rect 3235 377 3246 393
rect 3292 384 3308 400
rect 3315 398 3345 450
rect 3379 446 3380 453
rect 3364 438 3380 446
rect 3351 406 3364 425
rect 3379 406 3409 422
rect 3351 390 3425 406
rect 3351 388 3364 390
rect 3379 388 3413 390
rect 3016 366 3029 368
rect 3044 366 3078 368
rect 3016 350 3078 366
rect 3122 361 3138 364
rect 3200 361 3230 372
rect 3278 368 3324 384
rect 3351 372 3425 388
rect 3278 366 3312 368
rect 3277 350 3324 366
rect 3351 350 3364 372
rect 3379 350 3409 372
rect 3436 350 3437 366
rect 3452 350 3465 510
rect 3495 406 3508 510
rect 3553 488 3554 498
rect 3569 488 3582 498
rect 3553 484 3582 488
rect 3587 484 3617 510
rect 3635 496 3651 498
rect 3723 496 3776 510
rect 3724 494 3788 496
rect 3831 494 3846 510
rect 3895 507 3925 510
rect 3895 504 3931 507
rect 3861 496 3877 498
rect 3635 484 3650 488
rect 3553 482 3650 484
rect 3678 482 3846 494
rect 3862 484 3877 488
rect 3895 485 3934 504
rect 3953 498 3960 499
rect 3959 491 3960 498
rect 3943 488 3944 491
rect 3959 488 3972 491
rect 3895 484 3925 485
rect 3934 484 3940 485
rect 3943 484 3972 488
rect 3862 483 3972 484
rect 3862 482 3978 483
rect 3537 474 3588 482
rect 3537 462 3562 474
rect 3569 462 3588 474
rect 3619 474 3669 482
rect 3619 466 3635 474
rect 3642 472 3669 474
rect 3678 472 3899 482
rect 3642 462 3899 472
rect 3928 474 3978 482
rect 3928 465 3944 474
rect 3537 454 3588 462
rect 3635 454 3899 462
rect 3925 462 3944 465
rect 3951 462 3978 474
rect 3925 454 3978 462
rect 3553 446 3554 454
rect 3569 446 3582 454
rect 3553 438 3569 446
rect 3550 431 3569 434
rect 3550 422 3572 431
rect 3523 412 3572 422
rect 3523 406 3553 412
rect 3572 407 3577 412
rect 3495 390 3569 406
rect 3587 398 3617 454
rect 3652 444 3860 454
rect 3895 450 3940 454
rect 3943 453 3944 454
rect 3959 453 3972 454
rect 3678 414 3867 444
rect 3693 411 3867 414
rect 3686 408 3867 411
rect 3495 388 3508 390
rect 3523 388 3557 390
rect 3495 372 3569 388
rect 3596 384 3609 398
rect 3624 384 3640 400
rect 3686 395 3697 408
rect 3479 350 3480 366
rect 3495 350 3508 372
rect 3523 350 3553 372
rect 3596 368 3658 384
rect 3686 377 3697 393
rect 3702 388 3712 408
rect 3722 388 3736 408
rect 3739 395 3748 408
rect 3764 395 3773 408
rect 3702 377 3736 388
rect 3739 377 3748 393
rect 3764 377 3773 393
rect 3780 388 3790 408
rect 3800 388 3814 408
rect 3815 395 3826 408
rect 3780 377 3814 388
rect 3815 377 3826 393
rect 3872 384 3888 400
rect 3895 398 3925 450
rect 3959 446 3960 453
rect 3944 438 3960 446
rect 3931 406 3944 425
rect 3959 406 3989 422
rect 3931 390 4005 406
rect 3931 388 3944 390
rect 3959 388 3993 390
rect 3596 366 3609 368
rect 3624 366 3658 368
rect 3596 350 3658 366
rect 3702 361 3718 364
rect 3780 361 3810 372
rect 3858 368 3904 384
rect 3931 372 4005 388
rect 3858 366 3892 368
rect 3857 350 3904 366
rect 3931 350 3944 372
rect 3959 350 3989 372
rect 4016 350 4017 366
rect 4032 350 4045 510
rect 4075 406 4088 510
rect 4133 488 4134 498
rect 4149 488 4162 498
rect 4133 484 4162 488
rect 4167 484 4197 510
rect 4215 496 4231 498
rect 4303 496 4356 510
rect 4304 494 4368 496
rect 4411 494 4426 510
rect 4475 507 4505 510
rect 4475 504 4511 507
rect 4441 496 4457 498
rect 4215 484 4230 488
rect 4133 482 4230 484
rect 4258 482 4426 494
rect 4442 484 4457 488
rect 4475 485 4514 504
rect 4533 498 4540 499
rect 4539 491 4540 498
rect 4523 488 4524 491
rect 4539 488 4552 491
rect 4475 484 4505 485
rect 4514 484 4520 485
rect 4523 484 4552 488
rect 4442 483 4552 484
rect 4442 482 4558 483
rect 4117 474 4168 482
rect 4117 462 4142 474
rect 4149 462 4168 474
rect 4199 474 4249 482
rect 4199 466 4215 474
rect 4222 472 4249 474
rect 4258 472 4479 482
rect 4222 462 4479 472
rect 4508 474 4558 482
rect 4508 465 4524 474
rect 4117 454 4168 462
rect 4215 454 4479 462
rect 4505 462 4524 465
rect 4531 462 4558 474
rect 4505 454 4558 462
rect 4133 446 4134 454
rect 4149 446 4162 454
rect 4133 438 4149 446
rect 4130 431 4149 434
rect 4130 422 4152 431
rect 4103 412 4152 422
rect 4103 406 4133 412
rect 4152 407 4157 412
rect 4075 390 4149 406
rect 4167 398 4197 454
rect 4232 444 4440 454
rect 4475 450 4520 454
rect 4523 453 4524 454
rect 4539 453 4552 454
rect 4258 414 4447 444
rect 4273 411 4447 414
rect 4266 408 4447 411
rect 4075 388 4088 390
rect 4103 388 4137 390
rect 4075 372 4149 388
rect 4176 384 4189 398
rect 4204 384 4220 400
rect 4266 395 4277 408
rect 4059 350 4060 366
rect 4075 350 4088 372
rect 4103 350 4133 372
rect 4176 368 4238 384
rect 4266 377 4277 393
rect 4282 388 4292 408
rect 4302 388 4316 408
rect 4319 395 4328 408
rect 4344 395 4353 408
rect 4282 377 4316 388
rect 4319 377 4328 393
rect 4344 377 4353 393
rect 4360 388 4370 408
rect 4380 388 4394 408
rect 4395 395 4406 408
rect 4360 377 4394 388
rect 4395 377 4406 393
rect 4452 384 4468 400
rect 4475 398 4505 450
rect 4539 446 4540 453
rect 4524 438 4540 446
rect 4511 406 4524 425
rect 4539 406 4569 422
rect 4511 390 4585 406
rect 4511 388 4524 390
rect 4539 388 4573 390
rect 4176 366 4189 368
rect 4204 366 4238 368
rect 4176 350 4238 366
rect 4282 361 4298 364
rect 4360 361 4390 372
rect 4438 368 4484 384
rect 4511 372 4585 388
rect 4438 366 4472 368
rect 4437 350 4484 366
rect 4511 350 4524 372
rect 4539 350 4569 372
rect 4596 350 4597 366
rect 4612 350 4625 510
rect 4655 406 4668 510
rect 4713 488 4714 498
rect 4729 488 4742 498
rect 4713 484 4742 488
rect 4747 484 4777 510
rect 4795 496 4811 498
rect 4883 496 4936 510
rect 4884 494 4948 496
rect 4991 494 5006 510
rect 5055 507 5085 510
rect 5055 504 5091 507
rect 5021 496 5037 498
rect 4795 484 4810 488
rect 4713 482 4810 484
rect 4838 482 5006 494
rect 5022 484 5037 488
rect 5055 485 5094 504
rect 5113 498 5120 499
rect 5119 491 5120 498
rect 5103 488 5104 491
rect 5119 488 5132 491
rect 5055 484 5085 485
rect 5094 484 5100 485
rect 5103 484 5132 488
rect 5022 483 5132 484
rect 5022 482 5138 483
rect 4697 474 4748 482
rect 4697 462 4722 474
rect 4729 462 4748 474
rect 4779 474 4829 482
rect 4779 466 4795 474
rect 4802 472 4829 474
rect 4838 472 5059 482
rect 4802 462 5059 472
rect 5088 474 5138 482
rect 5088 465 5104 474
rect 4697 454 4748 462
rect 4795 454 5059 462
rect 5085 462 5104 465
rect 5111 462 5138 474
rect 5085 454 5138 462
rect 4713 446 4714 454
rect 4729 446 4742 454
rect 4713 438 4729 446
rect 4710 431 4729 434
rect 4710 422 4732 431
rect 4683 412 4732 422
rect 4683 406 4713 412
rect 4732 407 4737 412
rect 4655 390 4729 406
rect 4747 398 4777 454
rect 4812 444 5020 454
rect 5055 450 5100 454
rect 5103 453 5104 454
rect 5119 453 5132 454
rect 4838 414 5027 444
rect 4853 411 5027 414
rect 4846 408 5027 411
rect 4655 388 4668 390
rect 4683 388 4717 390
rect 4655 372 4729 388
rect 4756 384 4769 398
rect 4784 384 4800 400
rect 4846 395 4857 408
rect 4639 350 4640 366
rect 4655 350 4668 372
rect 4683 350 4713 372
rect 4756 368 4818 384
rect 4846 377 4857 393
rect 4862 388 4872 408
rect 4882 388 4896 408
rect 4899 395 4908 408
rect 4924 395 4933 408
rect 4862 377 4896 388
rect 4899 377 4908 393
rect 4924 377 4933 393
rect 4940 388 4950 408
rect 4960 388 4974 408
rect 4975 395 4986 408
rect 4940 377 4974 388
rect 4975 377 4986 393
rect 5032 384 5048 400
rect 5055 398 5085 450
rect 5119 446 5120 453
rect 5104 438 5120 446
rect 5091 406 5104 425
rect 5119 406 5149 422
rect 5091 390 5165 406
rect 5091 388 5104 390
rect 5119 388 5153 390
rect 4756 366 4769 368
rect 4784 366 4818 368
rect 4756 350 4818 366
rect 4862 361 4878 364
rect 4940 361 4970 372
rect 5018 368 5064 384
rect 5091 372 5165 388
rect 5018 366 5052 368
rect 5017 350 5064 366
rect 5091 350 5104 372
rect 5119 350 5149 372
rect 5176 350 5177 366
rect 5192 350 5205 510
rect 5235 406 5248 510
rect 5293 488 5294 498
rect 5309 488 5322 498
rect 5293 484 5322 488
rect 5327 484 5357 510
rect 5375 496 5391 498
rect 5463 496 5516 510
rect 5464 494 5528 496
rect 5571 494 5586 510
rect 5635 507 5665 510
rect 5635 504 5671 507
rect 5601 496 5617 498
rect 5375 484 5390 488
rect 5293 482 5390 484
rect 5418 482 5586 494
rect 5602 484 5617 488
rect 5635 485 5674 504
rect 5693 498 5700 499
rect 5699 491 5700 498
rect 5683 488 5684 491
rect 5699 488 5712 491
rect 5635 484 5665 485
rect 5674 484 5680 485
rect 5683 484 5712 488
rect 5602 483 5712 484
rect 5602 482 5718 483
rect 5277 474 5328 482
rect 5277 462 5302 474
rect 5309 462 5328 474
rect 5359 474 5409 482
rect 5359 466 5375 474
rect 5382 472 5409 474
rect 5418 472 5639 482
rect 5382 462 5639 472
rect 5668 474 5718 482
rect 5668 465 5684 474
rect 5277 454 5328 462
rect 5375 454 5639 462
rect 5665 462 5684 465
rect 5691 462 5718 474
rect 5665 454 5718 462
rect 5293 446 5294 454
rect 5309 446 5322 454
rect 5293 438 5309 446
rect 5290 431 5309 434
rect 5290 422 5312 431
rect 5263 412 5312 422
rect 5263 406 5293 412
rect 5312 407 5317 412
rect 5235 390 5309 406
rect 5327 398 5357 454
rect 5392 444 5600 454
rect 5635 450 5680 454
rect 5683 453 5684 454
rect 5699 453 5712 454
rect 5418 414 5607 444
rect 5433 411 5607 414
rect 5426 408 5607 411
rect 5235 388 5248 390
rect 5263 388 5297 390
rect 5235 372 5309 388
rect 5336 384 5349 398
rect 5364 384 5380 400
rect 5426 395 5437 408
rect 5219 350 5220 366
rect 5235 350 5248 372
rect 5263 350 5293 372
rect 5336 368 5398 384
rect 5426 377 5437 393
rect 5442 388 5452 408
rect 5462 388 5476 408
rect 5479 395 5488 408
rect 5504 395 5513 408
rect 5442 377 5476 388
rect 5479 377 5488 393
rect 5504 377 5513 393
rect 5520 388 5530 408
rect 5540 388 5554 408
rect 5555 395 5566 408
rect 5520 377 5554 388
rect 5555 377 5566 393
rect 5612 384 5628 400
rect 5635 398 5665 450
rect 5699 446 5700 453
rect 5684 438 5700 446
rect 5671 406 5684 425
rect 5699 406 5729 422
rect 5671 390 5745 406
rect 5671 388 5684 390
rect 5699 388 5733 390
rect 5336 366 5349 368
rect 5364 366 5398 368
rect 5336 350 5398 366
rect 5442 361 5458 364
rect 5520 361 5550 372
rect 5598 368 5644 384
rect 5671 372 5745 388
rect 5598 366 5632 368
rect 5597 350 5644 366
rect 5671 350 5684 372
rect 5699 350 5729 372
rect 5756 350 5757 366
rect 5772 350 5785 510
rect 5815 406 5828 510
rect 5873 488 5874 498
rect 5889 488 5902 498
rect 5873 484 5902 488
rect 5907 484 5937 510
rect 5955 496 5971 498
rect 6043 496 6096 510
rect 6044 494 6108 496
rect 6151 494 6166 510
rect 6215 507 6245 510
rect 6215 504 6251 507
rect 6181 496 6197 498
rect 5955 484 5970 488
rect 5873 482 5970 484
rect 5998 482 6166 494
rect 6182 484 6197 488
rect 6215 485 6254 504
rect 6273 498 6280 499
rect 6279 491 6280 498
rect 6263 488 6264 491
rect 6279 488 6292 491
rect 6215 484 6245 485
rect 6254 484 6260 485
rect 6263 484 6292 488
rect 6182 483 6292 484
rect 6182 482 6298 483
rect 5857 474 5908 482
rect 5857 462 5882 474
rect 5889 462 5908 474
rect 5939 474 5989 482
rect 5939 466 5955 474
rect 5962 472 5989 474
rect 5998 472 6219 482
rect 5962 462 6219 472
rect 6248 474 6298 482
rect 6248 465 6264 474
rect 5857 454 5908 462
rect 5955 454 6219 462
rect 6245 462 6264 465
rect 6271 462 6298 474
rect 6245 454 6298 462
rect 5873 446 5874 454
rect 5889 446 5902 454
rect 5873 438 5889 446
rect 5870 431 5889 434
rect 5870 422 5892 431
rect 5843 412 5892 422
rect 5843 406 5873 412
rect 5892 407 5897 412
rect 5815 390 5889 406
rect 5907 398 5937 454
rect 5972 444 6180 454
rect 6215 450 6260 454
rect 6263 453 6264 454
rect 6279 453 6292 454
rect 5998 414 6187 444
rect 6013 411 6187 414
rect 6006 408 6187 411
rect 5815 388 5828 390
rect 5843 388 5877 390
rect 5815 372 5889 388
rect 5916 384 5929 398
rect 5944 384 5960 400
rect 6006 395 6017 408
rect 5799 350 5800 366
rect 5815 350 5828 372
rect 5843 350 5873 372
rect 5916 368 5978 384
rect 6006 377 6017 393
rect 6022 388 6032 408
rect 6042 388 6056 408
rect 6059 395 6068 408
rect 6084 395 6093 408
rect 6022 377 6056 388
rect 6059 377 6068 393
rect 6084 377 6093 393
rect 6100 388 6110 408
rect 6120 388 6134 408
rect 6135 395 6146 408
rect 6100 377 6134 388
rect 6135 377 6146 393
rect 6192 384 6208 400
rect 6215 398 6245 450
rect 6279 446 6280 453
rect 6264 438 6280 446
rect 6251 406 6264 425
rect 6279 406 6309 422
rect 6251 390 6325 406
rect 6251 388 6264 390
rect 6279 388 6313 390
rect 5916 366 5929 368
rect 5944 366 5978 368
rect 5916 350 5978 366
rect 6022 361 6038 364
rect 6100 361 6130 372
rect 6178 368 6224 384
rect 6251 372 6325 388
rect 6178 366 6212 368
rect 6177 350 6224 366
rect 6251 350 6264 372
rect 6279 350 6309 372
rect 6336 350 6337 366
rect 6352 350 6365 510
rect 6395 406 6408 510
rect 6453 488 6454 498
rect 6469 488 6482 498
rect 6453 484 6482 488
rect 6487 484 6517 510
rect 6535 496 6551 498
rect 6623 496 6676 510
rect 6624 494 6688 496
rect 6731 494 6746 510
rect 6795 507 6825 510
rect 6795 504 6831 507
rect 6761 496 6777 498
rect 6535 484 6550 488
rect 6453 482 6550 484
rect 6578 482 6746 494
rect 6762 484 6777 488
rect 6795 485 6834 504
rect 6853 498 6860 499
rect 6859 491 6860 498
rect 6843 488 6844 491
rect 6859 488 6872 491
rect 6795 484 6825 485
rect 6834 484 6840 485
rect 6843 484 6872 488
rect 6762 483 6872 484
rect 6762 482 6878 483
rect 6437 474 6488 482
rect 6437 462 6462 474
rect 6469 462 6488 474
rect 6519 474 6569 482
rect 6519 466 6535 474
rect 6542 472 6569 474
rect 6578 472 6799 482
rect 6542 462 6799 472
rect 6828 474 6878 482
rect 6828 465 6844 474
rect 6437 454 6488 462
rect 6535 454 6799 462
rect 6825 462 6844 465
rect 6851 462 6878 474
rect 6825 454 6878 462
rect 6453 446 6454 454
rect 6469 446 6482 454
rect 6453 438 6469 446
rect 6450 431 6469 434
rect 6450 422 6472 431
rect 6423 412 6472 422
rect 6423 406 6453 412
rect 6472 407 6477 412
rect 6395 390 6469 406
rect 6487 398 6517 454
rect 6552 444 6760 454
rect 6795 450 6840 454
rect 6843 453 6844 454
rect 6859 453 6872 454
rect 6578 414 6767 444
rect 6593 411 6767 414
rect 6586 408 6767 411
rect 6395 388 6408 390
rect 6423 388 6457 390
rect 6395 372 6469 388
rect 6496 384 6509 398
rect 6524 384 6540 400
rect 6586 395 6597 408
rect 6379 350 6380 366
rect 6395 350 6408 372
rect 6423 350 6453 372
rect 6496 368 6558 384
rect 6586 377 6597 393
rect 6602 388 6612 408
rect 6622 388 6636 408
rect 6639 395 6648 408
rect 6664 395 6673 408
rect 6602 377 6636 388
rect 6639 377 6648 393
rect 6664 377 6673 393
rect 6680 388 6690 408
rect 6700 388 6714 408
rect 6715 395 6726 408
rect 6680 377 6714 388
rect 6715 377 6726 393
rect 6772 384 6788 400
rect 6795 398 6825 450
rect 6859 446 6860 453
rect 6844 438 6860 446
rect 6831 406 6844 425
rect 6859 406 6889 422
rect 6831 390 6905 406
rect 6831 388 6844 390
rect 6859 388 6893 390
rect 6496 366 6509 368
rect 6524 366 6558 368
rect 6496 350 6558 366
rect 6602 361 6618 364
rect 6680 361 6710 372
rect 6758 368 6804 384
rect 6831 372 6905 388
rect 6758 366 6792 368
rect 6757 350 6804 366
rect 6831 350 6844 372
rect 6859 350 6889 372
rect 6916 350 6917 366
rect 6932 350 6945 510
rect 6975 406 6988 510
rect 7033 488 7034 498
rect 7049 488 7062 498
rect 7033 484 7062 488
rect 7067 484 7097 510
rect 7115 496 7131 498
rect 7203 496 7256 510
rect 7204 494 7268 496
rect 7311 494 7326 510
rect 7375 507 7405 510
rect 7375 504 7411 507
rect 7341 496 7357 498
rect 7115 484 7130 488
rect 7033 482 7130 484
rect 7158 482 7326 494
rect 7342 484 7357 488
rect 7375 485 7414 504
rect 7433 498 7440 499
rect 7439 491 7440 498
rect 7423 488 7424 491
rect 7439 488 7452 491
rect 7375 484 7405 485
rect 7414 484 7420 485
rect 7423 484 7452 488
rect 7342 483 7452 484
rect 7342 482 7458 483
rect 7017 474 7068 482
rect 7017 462 7042 474
rect 7049 462 7068 474
rect 7099 474 7149 482
rect 7099 466 7115 474
rect 7122 472 7149 474
rect 7158 472 7379 482
rect 7122 462 7379 472
rect 7408 474 7458 482
rect 7408 465 7424 474
rect 7017 454 7068 462
rect 7115 454 7379 462
rect 7405 462 7424 465
rect 7431 462 7458 474
rect 7405 454 7458 462
rect 7033 446 7034 454
rect 7049 446 7062 454
rect 7033 438 7049 446
rect 7030 431 7049 434
rect 7030 422 7052 431
rect 7003 412 7052 422
rect 7003 406 7033 412
rect 7052 407 7057 412
rect 6975 390 7049 406
rect 7067 398 7097 454
rect 7132 444 7340 454
rect 7375 450 7420 454
rect 7423 453 7424 454
rect 7439 453 7452 454
rect 7158 414 7347 444
rect 7173 411 7347 414
rect 7166 408 7347 411
rect 6975 388 6988 390
rect 7003 388 7037 390
rect 6975 372 7049 388
rect 7076 384 7089 398
rect 7104 384 7120 400
rect 7166 395 7177 408
rect 6959 350 6960 366
rect 6975 350 6988 372
rect 7003 350 7033 372
rect 7076 368 7138 384
rect 7166 377 7177 393
rect 7182 388 7192 408
rect 7202 388 7216 408
rect 7219 395 7228 408
rect 7244 395 7253 408
rect 7182 377 7216 388
rect 7219 377 7228 393
rect 7244 377 7253 393
rect 7260 388 7270 408
rect 7280 388 7294 408
rect 7295 395 7306 408
rect 7260 377 7294 388
rect 7295 377 7306 393
rect 7352 384 7368 400
rect 7375 398 7405 450
rect 7439 446 7440 453
rect 7424 438 7440 446
rect 7411 406 7424 425
rect 7439 406 7469 422
rect 7411 390 7485 406
rect 7411 388 7424 390
rect 7439 388 7473 390
rect 7076 366 7089 368
rect 7104 366 7138 368
rect 7076 350 7138 366
rect 7182 361 7198 364
rect 7260 361 7290 372
rect 7338 368 7384 384
rect 7411 372 7485 388
rect 7338 366 7372 368
rect 7337 350 7384 366
rect 7411 350 7424 372
rect 7439 350 7469 372
rect 7496 350 7497 366
rect 7512 350 7525 510
rect 7555 406 7568 510
rect 7613 488 7614 498
rect 7629 488 7642 498
rect 7613 484 7642 488
rect 7647 484 7677 510
rect 7695 496 7711 498
rect 7783 496 7836 510
rect 7784 494 7848 496
rect 7891 494 7906 510
rect 7955 507 7985 510
rect 7955 504 7991 507
rect 7921 496 7937 498
rect 7695 484 7710 488
rect 7613 482 7710 484
rect 7738 482 7906 494
rect 7922 484 7937 488
rect 7955 485 7994 504
rect 8013 498 8020 499
rect 8019 491 8020 498
rect 8003 488 8004 491
rect 8019 488 8032 491
rect 7955 484 7985 485
rect 7994 484 8000 485
rect 8003 484 8032 488
rect 7922 483 8032 484
rect 7922 482 8038 483
rect 7597 474 7648 482
rect 7597 462 7622 474
rect 7629 462 7648 474
rect 7679 474 7729 482
rect 7679 466 7695 474
rect 7702 472 7729 474
rect 7738 472 7959 482
rect 7702 462 7959 472
rect 7988 474 8038 482
rect 7988 465 8004 474
rect 7597 454 7648 462
rect 7695 454 7959 462
rect 7985 462 8004 465
rect 8011 462 8038 474
rect 7985 454 8038 462
rect 7613 446 7614 454
rect 7629 446 7642 454
rect 7613 438 7629 446
rect 7610 431 7629 434
rect 7610 422 7632 431
rect 7583 412 7632 422
rect 7583 406 7613 412
rect 7632 407 7637 412
rect 7555 390 7629 406
rect 7647 398 7677 454
rect 7712 444 7920 454
rect 7955 450 8000 454
rect 8003 453 8004 454
rect 8019 453 8032 454
rect 7738 414 7927 444
rect 7753 411 7927 414
rect 7746 408 7927 411
rect 7555 388 7568 390
rect 7583 388 7617 390
rect 7555 372 7629 388
rect 7656 384 7669 398
rect 7684 384 7700 400
rect 7746 395 7757 408
rect 7539 350 7540 366
rect 7555 350 7568 372
rect 7583 350 7613 372
rect 7656 368 7718 384
rect 7746 377 7757 393
rect 7762 388 7772 408
rect 7782 388 7796 408
rect 7799 395 7808 408
rect 7824 395 7833 408
rect 7762 377 7796 388
rect 7799 377 7808 393
rect 7824 377 7833 393
rect 7840 388 7850 408
rect 7860 388 7874 408
rect 7875 395 7886 408
rect 7840 377 7874 388
rect 7875 377 7886 393
rect 7932 384 7948 400
rect 7955 398 7985 450
rect 8019 446 8020 453
rect 8004 438 8020 446
rect 7991 406 8004 425
rect 8019 406 8049 422
rect 7991 390 8065 406
rect 7991 388 8004 390
rect 8019 388 8053 390
rect 7656 366 7669 368
rect 7684 366 7718 368
rect 7656 350 7718 366
rect 7762 361 7778 364
rect 7840 361 7870 372
rect 7918 368 7964 384
rect 7991 372 8065 388
rect 7918 366 7952 368
rect 7917 350 7964 366
rect 7991 350 8004 372
rect 8019 350 8049 372
rect 8076 350 8077 366
rect 8092 350 8105 510
rect 8135 406 8148 510
rect 8193 488 8194 498
rect 8209 488 8222 498
rect 8193 484 8222 488
rect 8227 484 8257 510
rect 8275 496 8291 498
rect 8363 496 8416 510
rect 8364 494 8428 496
rect 8471 494 8486 510
rect 8535 507 8565 510
rect 8535 504 8571 507
rect 8501 496 8517 498
rect 8275 484 8290 488
rect 8193 482 8290 484
rect 8318 482 8486 494
rect 8502 484 8517 488
rect 8535 485 8574 504
rect 8593 498 8600 499
rect 8599 491 8600 498
rect 8583 488 8584 491
rect 8599 488 8612 491
rect 8535 484 8565 485
rect 8574 484 8580 485
rect 8583 484 8612 488
rect 8502 483 8612 484
rect 8502 482 8618 483
rect 8177 474 8228 482
rect 8177 462 8202 474
rect 8209 462 8228 474
rect 8259 474 8309 482
rect 8259 466 8275 474
rect 8282 472 8309 474
rect 8318 472 8539 482
rect 8282 462 8539 472
rect 8568 474 8618 482
rect 8568 465 8584 474
rect 8177 454 8228 462
rect 8275 454 8539 462
rect 8565 462 8584 465
rect 8591 462 8618 474
rect 8565 454 8618 462
rect 8193 446 8194 454
rect 8209 446 8222 454
rect 8193 438 8209 446
rect 8190 431 8209 434
rect 8190 422 8212 431
rect 8163 412 8212 422
rect 8163 406 8193 412
rect 8212 407 8217 412
rect 8135 390 8209 406
rect 8227 398 8257 454
rect 8292 444 8500 454
rect 8535 450 8580 454
rect 8583 453 8584 454
rect 8599 453 8612 454
rect 8318 414 8507 444
rect 8333 411 8507 414
rect 8326 408 8507 411
rect 8135 388 8148 390
rect 8163 388 8197 390
rect 8135 372 8209 388
rect 8236 384 8249 398
rect 8264 384 8280 400
rect 8326 395 8337 408
rect 8119 350 8120 366
rect 8135 350 8148 372
rect 8163 350 8193 372
rect 8236 368 8298 384
rect 8326 377 8337 393
rect 8342 388 8352 408
rect 8362 388 8376 408
rect 8379 395 8388 408
rect 8404 395 8413 408
rect 8342 377 8376 388
rect 8379 377 8388 393
rect 8404 377 8413 393
rect 8420 388 8430 408
rect 8440 388 8454 408
rect 8455 395 8466 408
rect 8420 377 8454 388
rect 8455 377 8466 393
rect 8512 384 8528 400
rect 8535 398 8565 450
rect 8599 446 8600 453
rect 8584 438 8600 446
rect 8571 406 8584 425
rect 8599 406 8629 422
rect 8571 390 8645 406
rect 8571 388 8584 390
rect 8599 388 8633 390
rect 8236 366 8249 368
rect 8264 366 8298 368
rect 8236 350 8298 366
rect 8342 361 8358 364
rect 8420 361 8450 372
rect 8498 368 8544 384
rect 8571 372 8645 388
rect 8498 366 8532 368
rect 8497 350 8544 366
rect 8571 350 8584 372
rect 8599 350 8629 372
rect 8656 350 8657 366
rect 8672 350 8685 510
rect 8715 406 8728 510
rect 8773 488 8774 498
rect 8789 488 8802 498
rect 8773 484 8802 488
rect 8807 484 8837 510
rect 8855 496 8871 498
rect 8943 496 8996 510
rect 8944 494 9008 496
rect 9051 494 9066 510
rect 9115 507 9145 510
rect 9115 504 9151 507
rect 9081 496 9097 498
rect 8855 484 8870 488
rect 8773 482 8870 484
rect 8898 482 9066 494
rect 9082 484 9097 488
rect 9115 485 9154 504
rect 9173 498 9180 499
rect 9179 491 9180 498
rect 9163 488 9164 491
rect 9179 488 9192 491
rect 9115 484 9145 485
rect 9154 484 9160 485
rect 9163 484 9192 488
rect 9082 483 9192 484
rect 9082 482 9198 483
rect 8757 474 8808 482
rect 8757 462 8782 474
rect 8789 462 8808 474
rect 8839 474 8889 482
rect 8839 466 8855 474
rect 8862 472 8889 474
rect 8898 472 9119 482
rect 8862 462 9119 472
rect 9148 474 9198 482
rect 9148 465 9164 474
rect 8757 454 8808 462
rect 8855 454 9119 462
rect 9145 462 9164 465
rect 9171 462 9198 474
rect 9145 454 9198 462
rect 8773 446 8774 454
rect 8789 446 8802 454
rect 8773 438 8789 446
rect 8770 431 8789 434
rect 8770 422 8792 431
rect 8743 412 8792 422
rect 8743 406 8773 412
rect 8792 407 8797 412
rect 8715 390 8789 406
rect 8807 398 8837 454
rect 8872 444 9080 454
rect 9115 450 9160 454
rect 9163 453 9164 454
rect 9179 453 9192 454
rect 8898 414 9087 444
rect 8913 411 9087 414
rect 8906 408 9087 411
rect 8715 388 8728 390
rect 8743 388 8777 390
rect 8715 372 8789 388
rect 8816 384 8829 398
rect 8844 384 8860 400
rect 8906 395 8917 408
rect 8699 350 8700 366
rect 8715 350 8728 372
rect 8743 350 8773 372
rect 8816 368 8878 384
rect 8906 377 8917 393
rect 8922 388 8932 408
rect 8942 388 8956 408
rect 8959 395 8968 408
rect 8984 395 8993 408
rect 8922 377 8956 388
rect 8959 377 8968 393
rect 8984 377 8993 393
rect 9000 388 9010 408
rect 9020 388 9034 408
rect 9035 395 9046 408
rect 9000 377 9034 388
rect 9035 377 9046 393
rect 9092 384 9108 400
rect 9115 398 9145 450
rect 9179 446 9180 453
rect 9164 438 9180 446
rect 9151 406 9164 425
rect 9179 406 9209 422
rect 9151 390 9225 406
rect 9151 388 9164 390
rect 9179 388 9213 390
rect 8816 366 8829 368
rect 8844 366 8878 368
rect 8816 350 8878 366
rect 8922 361 8938 364
rect 9000 361 9030 372
rect 9078 368 9124 384
rect 9151 372 9225 388
rect 9078 366 9112 368
rect 9077 350 9124 366
rect 9151 350 9164 372
rect 9179 350 9209 372
rect 9236 350 9237 366
rect 9252 350 9265 510
rect -7 342 34 350
rect -7 316 8 342
rect 15 316 34 342
rect 98 338 160 350
rect 172 338 247 350
rect 305 338 380 350
rect 392 338 423 350
rect 429 338 464 350
rect 98 336 260 338
rect -7 308 34 316
rect 116 312 129 336
rect 144 334 159 336
rect -1 298 0 308
rect 15 298 28 308
rect 43 298 73 312
rect 116 298 159 312
rect 183 309 190 316
rect 193 312 260 336
rect 292 336 464 338
rect 262 314 290 318
rect 292 314 372 336
rect 393 334 408 336
rect 262 312 372 314
rect 193 308 372 312
rect 166 298 196 308
rect 198 298 351 308
rect 359 298 389 308
rect 393 298 423 312
rect 451 298 464 336
rect 536 342 571 350
rect 536 316 537 342
rect 544 316 571 342
rect 479 298 509 312
rect 536 308 571 316
rect 573 342 614 350
rect 573 316 588 342
rect 595 316 614 342
rect 678 338 740 350
rect 752 338 827 350
rect 885 338 960 350
rect 972 338 1003 350
rect 1009 338 1044 350
rect 678 336 840 338
rect 573 308 614 316
rect 696 312 709 336
rect 724 334 739 336
rect 536 298 537 308
rect 552 298 565 308
rect 579 298 580 308
rect 595 298 608 308
rect 623 298 653 312
rect 696 298 739 312
rect 763 309 770 316
rect 773 312 840 336
rect 872 336 1044 338
rect 842 314 870 318
rect 872 314 952 336
rect 973 334 988 336
rect 842 312 952 314
rect 773 308 952 312
rect 746 298 776 308
rect 778 298 931 308
rect 939 298 969 308
rect 973 298 1003 312
rect 1031 298 1044 336
rect 1116 342 1151 350
rect 1116 316 1117 342
rect 1124 316 1151 342
rect 1059 298 1089 312
rect 1116 308 1151 316
rect 1153 342 1194 350
rect 1153 316 1168 342
rect 1175 316 1194 342
rect 1258 338 1320 350
rect 1332 338 1407 350
rect 1465 338 1540 350
rect 1552 338 1583 350
rect 1589 338 1624 350
rect 1258 336 1420 338
rect 1153 308 1194 316
rect 1276 312 1289 336
rect 1304 334 1319 336
rect 1116 298 1117 308
rect 1132 298 1145 308
rect 1159 298 1160 308
rect 1175 298 1188 308
rect 1203 298 1233 312
rect 1276 298 1319 312
rect 1343 309 1350 316
rect 1353 312 1420 336
rect 1452 336 1624 338
rect 1422 314 1450 318
rect 1452 314 1532 336
rect 1553 334 1568 336
rect 1422 312 1532 314
rect 1353 308 1532 312
rect 1326 298 1356 308
rect 1358 298 1511 308
rect 1519 298 1549 308
rect 1553 298 1583 312
rect 1611 298 1624 336
rect 1696 342 1731 350
rect 1696 316 1697 342
rect 1704 316 1731 342
rect 1639 298 1669 312
rect 1696 308 1731 316
rect 1733 342 1774 350
rect 1733 316 1748 342
rect 1755 316 1774 342
rect 1838 338 1900 350
rect 1912 338 1987 350
rect 2045 338 2120 350
rect 2132 338 2163 350
rect 2169 338 2204 350
rect 1838 336 2000 338
rect 1733 308 1774 316
rect 1856 312 1869 336
rect 1884 334 1899 336
rect 1696 298 1697 308
rect 1712 298 1725 308
rect 1739 298 1740 308
rect 1755 298 1768 308
rect 1783 298 1813 312
rect 1856 298 1899 312
rect 1923 309 1930 316
rect 1933 312 2000 336
rect 2032 336 2204 338
rect 2002 314 2030 318
rect 2032 314 2112 336
rect 2133 334 2148 336
rect 2002 312 2112 314
rect 1933 308 2112 312
rect 1906 298 1936 308
rect 1938 298 2091 308
rect 2099 298 2129 308
rect 2133 298 2163 312
rect 2191 298 2204 336
rect 2276 342 2311 350
rect 2276 316 2277 342
rect 2284 316 2311 342
rect 2219 298 2249 312
rect 2276 308 2311 316
rect 2313 342 2354 350
rect 2313 316 2328 342
rect 2335 316 2354 342
rect 2418 338 2480 350
rect 2492 338 2567 350
rect 2625 338 2700 350
rect 2712 338 2743 350
rect 2749 338 2784 350
rect 2418 336 2580 338
rect 2313 308 2354 316
rect 2436 312 2449 336
rect 2464 334 2479 336
rect 2276 298 2277 308
rect 2292 298 2305 308
rect 2319 298 2320 308
rect 2335 298 2348 308
rect 2363 298 2393 312
rect 2436 298 2479 312
rect 2503 309 2510 316
rect 2513 312 2580 336
rect 2612 336 2784 338
rect 2582 314 2610 318
rect 2612 314 2692 336
rect 2713 334 2728 336
rect 2582 312 2692 314
rect 2513 308 2692 312
rect 2486 298 2516 308
rect 2518 298 2671 308
rect 2679 298 2709 308
rect 2713 298 2743 312
rect 2771 298 2784 336
rect 2856 342 2891 350
rect 2856 316 2857 342
rect 2864 316 2891 342
rect 2799 298 2829 312
rect 2856 308 2891 316
rect 2893 342 2934 350
rect 2893 316 2908 342
rect 2915 316 2934 342
rect 2998 338 3060 350
rect 3072 338 3147 350
rect 3205 338 3280 350
rect 3292 338 3323 350
rect 3329 338 3364 350
rect 2998 336 3160 338
rect 2893 308 2934 316
rect 3016 312 3029 336
rect 3044 334 3059 336
rect 2856 298 2857 308
rect 2872 298 2885 308
rect 2899 298 2900 308
rect 2915 298 2928 308
rect 2943 298 2973 312
rect 3016 298 3059 312
rect 3083 309 3090 316
rect 3093 312 3160 336
rect 3192 336 3364 338
rect 3162 314 3190 318
rect 3192 314 3272 336
rect 3293 334 3308 336
rect 3162 312 3272 314
rect 3093 308 3272 312
rect 3066 298 3096 308
rect 3098 298 3251 308
rect 3259 298 3289 308
rect 3293 298 3323 312
rect 3351 298 3364 336
rect 3436 342 3471 350
rect 3436 316 3437 342
rect 3444 316 3471 342
rect 3379 298 3409 312
rect 3436 308 3471 316
rect 3473 342 3514 350
rect 3473 316 3488 342
rect 3495 316 3514 342
rect 3578 338 3640 350
rect 3652 338 3727 350
rect 3785 338 3860 350
rect 3872 338 3903 350
rect 3909 338 3944 350
rect 3578 336 3740 338
rect 3473 308 3514 316
rect 3596 312 3609 336
rect 3624 334 3639 336
rect 3436 298 3437 308
rect 3452 298 3465 308
rect 3479 298 3480 308
rect 3495 298 3508 308
rect 3523 298 3553 312
rect 3596 298 3639 312
rect 3663 309 3670 316
rect 3673 312 3740 336
rect 3772 336 3944 338
rect 3742 314 3770 318
rect 3772 314 3852 336
rect 3873 334 3888 336
rect 3742 312 3852 314
rect 3673 308 3852 312
rect 3646 298 3676 308
rect 3678 298 3831 308
rect 3839 298 3869 308
rect 3873 298 3903 312
rect 3931 298 3944 336
rect 4016 342 4051 350
rect 4016 316 4017 342
rect 4024 316 4051 342
rect 3959 298 3989 312
rect 4016 308 4051 316
rect 4053 342 4094 350
rect 4053 316 4068 342
rect 4075 316 4094 342
rect 4158 338 4220 350
rect 4232 338 4307 350
rect 4365 338 4440 350
rect 4452 338 4483 350
rect 4489 338 4524 350
rect 4158 336 4320 338
rect 4053 308 4094 316
rect 4176 312 4189 336
rect 4204 334 4219 336
rect 4016 298 4017 308
rect 4032 298 4045 308
rect 4059 298 4060 308
rect 4075 298 4088 308
rect 4103 298 4133 312
rect 4176 298 4219 312
rect 4243 309 4250 316
rect 4253 312 4320 336
rect 4352 336 4524 338
rect 4322 314 4350 318
rect 4352 314 4432 336
rect 4453 334 4468 336
rect 4322 312 4432 314
rect 4253 308 4432 312
rect 4226 298 4256 308
rect 4258 298 4411 308
rect 4419 298 4449 308
rect 4453 298 4483 312
rect 4511 298 4524 336
rect 4596 342 4631 350
rect 4596 316 4597 342
rect 4604 316 4631 342
rect 4539 298 4569 312
rect 4596 308 4631 316
rect 4633 342 4674 350
rect 4633 316 4648 342
rect 4655 316 4674 342
rect 4738 338 4800 350
rect 4812 338 4887 350
rect 4945 338 5020 350
rect 5032 338 5063 350
rect 5069 338 5104 350
rect 4738 336 4900 338
rect 4633 308 4674 316
rect 4756 312 4769 336
rect 4784 334 4799 336
rect 4596 298 4597 308
rect 4612 298 4625 308
rect 4639 298 4640 308
rect 4655 298 4668 308
rect 4683 298 4713 312
rect 4756 298 4799 312
rect 4823 309 4830 316
rect 4833 312 4900 336
rect 4932 336 5104 338
rect 4902 314 4930 318
rect 4932 314 5012 336
rect 5033 334 5048 336
rect 4902 312 5012 314
rect 4833 308 5012 312
rect 4806 298 4836 308
rect 4838 298 4991 308
rect 4999 298 5029 308
rect 5033 298 5063 312
rect 5091 298 5104 336
rect 5176 342 5211 350
rect 5176 316 5177 342
rect 5184 316 5211 342
rect 5119 298 5149 312
rect 5176 308 5211 316
rect 5213 342 5254 350
rect 5213 316 5228 342
rect 5235 316 5254 342
rect 5318 338 5380 350
rect 5392 338 5467 350
rect 5525 338 5600 350
rect 5612 338 5643 350
rect 5649 338 5684 350
rect 5318 336 5480 338
rect 5213 308 5254 316
rect 5336 312 5349 336
rect 5364 334 5379 336
rect 5176 298 5177 308
rect 5192 298 5205 308
rect 5219 298 5220 308
rect 5235 298 5248 308
rect 5263 298 5293 312
rect 5336 298 5379 312
rect 5403 309 5410 316
rect 5413 312 5480 336
rect 5512 336 5684 338
rect 5482 314 5510 318
rect 5512 314 5592 336
rect 5613 334 5628 336
rect 5482 312 5592 314
rect 5413 308 5592 312
rect 5386 298 5416 308
rect 5418 298 5571 308
rect 5579 298 5609 308
rect 5613 298 5643 312
rect 5671 298 5684 336
rect 5756 342 5791 350
rect 5756 316 5757 342
rect 5764 316 5791 342
rect 5699 298 5729 312
rect 5756 308 5791 316
rect 5793 342 5834 350
rect 5793 316 5808 342
rect 5815 316 5834 342
rect 5898 338 5960 350
rect 5972 338 6047 350
rect 6105 338 6180 350
rect 6192 338 6223 350
rect 6229 338 6264 350
rect 5898 336 6060 338
rect 5793 308 5834 316
rect 5916 312 5929 336
rect 5944 334 5959 336
rect 5756 298 5757 308
rect 5772 298 5785 308
rect 5799 298 5800 308
rect 5815 298 5828 308
rect 5843 298 5873 312
rect 5916 298 5959 312
rect 5983 309 5990 316
rect 5993 312 6060 336
rect 6092 336 6264 338
rect 6062 314 6090 318
rect 6092 314 6172 336
rect 6193 334 6208 336
rect 6062 312 6172 314
rect 5993 308 6172 312
rect 5966 298 5996 308
rect 5998 298 6151 308
rect 6159 298 6189 308
rect 6193 298 6223 312
rect 6251 298 6264 336
rect 6336 342 6371 350
rect 6336 316 6337 342
rect 6344 316 6371 342
rect 6279 298 6309 312
rect 6336 308 6371 316
rect 6373 342 6414 350
rect 6373 316 6388 342
rect 6395 316 6414 342
rect 6478 338 6540 350
rect 6552 338 6627 350
rect 6685 338 6760 350
rect 6772 338 6803 350
rect 6809 338 6844 350
rect 6478 336 6640 338
rect 6373 308 6414 316
rect 6496 312 6509 336
rect 6524 334 6539 336
rect 6336 298 6337 308
rect 6352 298 6365 308
rect 6379 298 6380 308
rect 6395 298 6408 308
rect 6423 298 6453 312
rect 6496 298 6539 312
rect 6563 309 6570 316
rect 6573 312 6640 336
rect 6672 336 6844 338
rect 6642 314 6670 318
rect 6672 314 6752 336
rect 6773 334 6788 336
rect 6642 312 6752 314
rect 6573 308 6752 312
rect 6546 298 6576 308
rect 6578 298 6731 308
rect 6739 298 6769 308
rect 6773 298 6803 312
rect 6831 298 6844 336
rect 6916 342 6951 350
rect 6916 316 6917 342
rect 6924 316 6951 342
rect 6859 298 6889 312
rect 6916 308 6951 316
rect 6953 342 6994 350
rect 6953 316 6968 342
rect 6975 316 6994 342
rect 7058 338 7120 350
rect 7132 338 7207 350
rect 7265 338 7340 350
rect 7352 338 7383 350
rect 7389 338 7424 350
rect 7058 336 7220 338
rect 6953 308 6994 316
rect 7076 312 7089 336
rect 7104 334 7119 336
rect 6916 298 6917 308
rect 6932 298 6945 308
rect 6959 298 6960 308
rect 6975 298 6988 308
rect 7003 298 7033 312
rect 7076 298 7119 312
rect 7143 309 7150 316
rect 7153 312 7220 336
rect 7252 336 7424 338
rect 7222 314 7250 318
rect 7252 314 7332 336
rect 7353 334 7368 336
rect 7222 312 7332 314
rect 7153 308 7332 312
rect 7126 298 7156 308
rect 7158 298 7311 308
rect 7319 298 7349 308
rect 7353 298 7383 312
rect 7411 298 7424 336
rect 7496 342 7531 350
rect 7496 316 7497 342
rect 7504 316 7531 342
rect 7439 298 7469 312
rect 7496 308 7531 316
rect 7533 342 7574 350
rect 7533 316 7548 342
rect 7555 316 7574 342
rect 7638 338 7700 350
rect 7712 338 7787 350
rect 7845 338 7920 350
rect 7932 338 7963 350
rect 7969 338 8004 350
rect 7638 336 7800 338
rect 7533 308 7574 316
rect 7656 312 7669 336
rect 7684 334 7699 336
rect 7496 298 7497 308
rect 7512 298 7525 308
rect 7539 298 7540 308
rect 7555 298 7568 308
rect 7583 298 7613 312
rect 7656 298 7699 312
rect 7723 309 7730 316
rect 7733 312 7800 336
rect 7832 336 8004 338
rect 7802 314 7830 318
rect 7832 314 7912 336
rect 7933 334 7948 336
rect 7802 312 7912 314
rect 7733 308 7912 312
rect 7706 298 7736 308
rect 7738 298 7891 308
rect 7899 298 7929 308
rect 7933 298 7963 312
rect 7991 298 8004 336
rect 8076 342 8111 350
rect 8076 316 8077 342
rect 8084 316 8111 342
rect 8019 298 8049 312
rect 8076 308 8111 316
rect 8113 342 8154 350
rect 8113 316 8128 342
rect 8135 316 8154 342
rect 8218 338 8280 350
rect 8292 338 8367 350
rect 8425 338 8500 350
rect 8512 338 8543 350
rect 8549 338 8584 350
rect 8218 336 8380 338
rect 8113 308 8154 316
rect 8236 312 8249 336
rect 8264 334 8279 336
rect 8076 298 8077 308
rect 8092 298 8105 308
rect 8119 298 8120 308
rect 8135 298 8148 308
rect 8163 298 8193 312
rect 8236 298 8279 312
rect 8303 309 8310 316
rect 8313 312 8380 336
rect 8412 336 8584 338
rect 8382 314 8410 318
rect 8412 314 8492 336
rect 8513 334 8528 336
rect 8382 312 8492 314
rect 8313 308 8492 312
rect 8286 298 8316 308
rect 8318 298 8471 308
rect 8479 298 8509 308
rect 8513 298 8543 312
rect 8571 298 8584 336
rect 8656 342 8691 350
rect 8656 316 8657 342
rect 8664 316 8691 342
rect 8599 298 8629 312
rect 8656 308 8691 316
rect 8693 342 8734 350
rect 8693 316 8708 342
rect 8715 316 8734 342
rect 8798 338 8860 350
rect 8872 338 8947 350
rect 9005 338 9080 350
rect 9092 338 9123 350
rect 9129 338 9164 350
rect 8798 336 8960 338
rect 8693 308 8734 316
rect 8816 312 8829 336
rect 8844 334 8859 336
rect 8656 298 8657 308
rect 8672 298 8685 308
rect 8699 298 8700 308
rect 8715 298 8728 308
rect 8743 298 8773 312
rect 8816 298 8859 312
rect 8883 309 8890 316
rect 8893 312 8960 336
rect 8992 336 9164 338
rect 8962 314 8990 318
rect 8992 314 9072 336
rect 9093 334 9108 336
rect 8962 312 9072 314
rect 8893 308 9072 312
rect 8866 298 8896 308
rect 8898 298 9051 308
rect 9059 298 9089 308
rect 9093 298 9123 312
rect 9151 298 9164 336
rect 9236 342 9271 350
rect 9236 316 9237 342
rect 9244 316 9271 342
rect 9179 298 9209 312
rect 9236 308 9271 316
rect 9236 298 9237 308
rect 9252 298 9265 308
rect -1 292 9265 298
rect 0 284 9265 292
rect 15 254 28 284
rect 43 266 73 284
rect 116 270 130 284
rect 166 270 386 284
rect 117 268 130 270
rect 83 256 98 268
rect 80 254 102 256
rect 107 254 137 268
rect 198 266 351 270
rect 180 254 372 266
rect 415 254 445 268
rect 451 254 464 284
rect 479 266 509 284
rect 552 254 565 284
rect 595 254 608 284
rect 623 266 653 284
rect 696 270 710 284
rect 746 270 966 284
rect 697 268 710 270
rect 663 256 678 268
rect 660 254 682 256
rect 687 254 717 268
rect 778 266 931 270
rect 760 254 952 266
rect 995 254 1025 268
rect 1031 254 1044 284
rect 1059 266 1089 284
rect 1132 254 1145 284
rect 1175 254 1188 284
rect 1203 266 1233 284
rect 1276 270 1290 284
rect 1326 270 1546 284
rect 1277 268 1290 270
rect 1243 256 1258 268
rect 1240 254 1262 256
rect 1267 254 1297 268
rect 1358 266 1511 270
rect 1340 254 1532 266
rect 1575 254 1605 268
rect 1611 254 1624 284
rect 1639 266 1669 284
rect 1712 254 1725 284
rect 1755 254 1768 284
rect 1783 266 1813 284
rect 1856 270 1870 284
rect 1906 270 2126 284
rect 1857 268 1870 270
rect 1823 256 1838 268
rect 1820 254 1842 256
rect 1847 254 1877 268
rect 1938 266 2091 270
rect 1920 254 2112 266
rect 2155 254 2185 268
rect 2191 254 2204 284
rect 2219 266 2249 284
rect 2292 254 2305 284
rect 2335 254 2348 284
rect 2363 266 2393 284
rect 2436 270 2450 284
rect 2486 270 2706 284
rect 2437 268 2450 270
rect 2403 256 2418 268
rect 2400 254 2422 256
rect 2427 254 2457 268
rect 2518 266 2671 270
rect 2500 254 2692 266
rect 2735 254 2765 268
rect 2771 254 2784 284
rect 2799 266 2829 284
rect 2872 254 2885 284
rect 2915 254 2928 284
rect 2943 266 2973 284
rect 3016 270 3030 284
rect 3066 270 3286 284
rect 3017 268 3030 270
rect 2983 256 2998 268
rect 2980 254 3002 256
rect 3007 254 3037 268
rect 3098 266 3251 270
rect 3080 254 3272 266
rect 3315 254 3345 268
rect 3351 254 3364 284
rect 3379 266 3409 284
rect 3452 254 3465 284
rect 3495 254 3508 284
rect 3523 266 3553 284
rect 3596 270 3610 284
rect 3646 270 3866 284
rect 3597 268 3610 270
rect 3563 256 3578 268
rect 3560 254 3582 256
rect 3587 254 3617 268
rect 3678 266 3831 270
rect 3660 254 3852 266
rect 3895 254 3925 268
rect 3931 254 3944 284
rect 3959 266 3989 284
rect 4032 254 4045 284
rect 4075 254 4088 284
rect 4103 266 4133 284
rect 4176 270 4190 284
rect 4226 270 4446 284
rect 4177 268 4190 270
rect 4143 256 4158 268
rect 4140 254 4162 256
rect 4167 254 4197 268
rect 4258 266 4411 270
rect 4240 254 4432 266
rect 4475 254 4505 268
rect 4511 254 4524 284
rect 4539 266 4569 284
rect 4612 254 4625 284
rect 4655 254 4668 284
rect 4683 266 4713 284
rect 4756 270 4770 284
rect 4806 270 5026 284
rect 4757 268 4770 270
rect 4723 256 4738 268
rect 4720 254 4742 256
rect 4747 254 4777 268
rect 4838 266 4991 270
rect 4820 254 5012 266
rect 5055 254 5085 268
rect 5091 254 5104 284
rect 5119 266 5149 284
rect 5192 254 5205 284
rect 5235 254 5248 284
rect 5263 266 5293 284
rect 5336 270 5350 284
rect 5386 270 5606 284
rect 5337 268 5350 270
rect 5303 256 5318 268
rect 5300 254 5322 256
rect 5327 254 5357 268
rect 5418 266 5571 270
rect 5400 254 5592 266
rect 5635 254 5665 268
rect 5671 254 5684 284
rect 5699 266 5729 284
rect 5772 254 5785 284
rect 5815 254 5828 284
rect 5843 266 5873 284
rect 5916 270 5930 284
rect 5966 270 6186 284
rect 5917 268 5930 270
rect 5883 256 5898 268
rect 5880 254 5902 256
rect 5907 254 5937 268
rect 5998 266 6151 270
rect 5980 254 6172 266
rect 6215 254 6245 268
rect 6251 254 6264 284
rect 6279 266 6309 284
rect 6352 254 6365 284
rect 6395 254 6408 284
rect 6423 266 6453 284
rect 6496 270 6510 284
rect 6546 270 6766 284
rect 6497 268 6510 270
rect 6463 256 6478 268
rect 6460 254 6482 256
rect 6487 254 6517 268
rect 6578 266 6731 270
rect 6560 254 6752 266
rect 6795 254 6825 268
rect 6831 254 6844 284
rect 6859 266 6889 284
rect 6932 254 6945 284
rect 6975 254 6988 284
rect 7003 266 7033 284
rect 7076 270 7090 284
rect 7126 270 7346 284
rect 7077 268 7090 270
rect 7043 256 7058 268
rect 7040 254 7062 256
rect 7067 254 7097 268
rect 7158 266 7311 270
rect 7140 254 7332 266
rect 7375 254 7405 268
rect 7411 254 7424 284
rect 7439 266 7469 284
rect 7512 254 7525 284
rect 7555 254 7568 284
rect 7583 266 7613 284
rect 7656 270 7670 284
rect 7706 270 7926 284
rect 7657 268 7670 270
rect 7623 256 7638 268
rect 7620 254 7642 256
rect 7647 254 7677 268
rect 7738 266 7891 270
rect 7720 254 7912 266
rect 7955 254 7985 268
rect 7991 254 8004 284
rect 8019 266 8049 284
rect 8092 254 8105 284
rect 8135 254 8148 284
rect 8163 266 8193 284
rect 8236 270 8250 284
rect 8286 270 8506 284
rect 8237 268 8250 270
rect 8203 256 8218 268
rect 8200 254 8222 256
rect 8227 254 8257 268
rect 8318 266 8471 270
rect 8300 254 8492 266
rect 8535 254 8565 268
rect 8571 254 8584 284
rect 8599 266 8629 284
rect 8672 254 8685 284
rect 8715 254 8728 284
rect 8743 266 8773 284
rect 8816 270 8830 284
rect 8866 270 9086 284
rect 8817 268 8830 270
rect 8783 256 8798 268
rect 8780 254 8802 256
rect 8807 254 8837 268
rect 8898 266 9051 270
rect 8880 254 9072 266
rect 9115 254 9145 268
rect 9151 254 9164 284
rect 9179 266 9209 284
rect 9252 254 9265 284
rect 0 240 9265 254
rect 15 136 28 240
rect 73 218 74 228
rect 89 218 102 228
rect 73 214 102 218
rect 107 214 137 240
rect 155 226 171 228
rect 243 226 296 240
rect 244 224 308 226
rect 155 214 170 218
rect 73 212 170 214
rect 57 204 108 212
rect 57 192 82 204
rect 89 192 108 204
rect 139 204 189 212
rect 139 196 155 204
rect 162 202 189 204
rect 198 204 213 208
rect 260 204 292 224
rect 351 212 366 240
rect 415 237 445 240
rect 415 234 451 237
rect 381 226 397 228
rect 382 214 397 218
rect 415 215 454 234
rect 473 228 480 229
rect 479 221 480 228
rect 463 218 464 221
rect 479 218 492 221
rect 415 214 445 215
rect 454 214 460 215
rect 463 214 492 218
rect 382 213 492 214
rect 382 212 498 213
rect 351 204 419 212
rect 198 202 267 204
rect 285 202 419 204
rect 162 198 234 202
rect 162 196 287 198
rect 162 192 234 196
rect 57 184 108 192
rect 155 188 234 192
rect 315 188 419 202
rect 448 204 498 212
rect 448 195 464 204
rect 155 184 419 188
rect 445 192 464 195
rect 471 192 498 204
rect 445 184 498 192
rect 73 176 74 184
rect 89 176 102 184
rect 73 168 89 176
rect 70 161 89 164
rect 70 152 92 161
rect 43 142 92 152
rect 43 136 73 142
rect 92 137 97 142
rect 15 120 89 136
rect 107 128 137 184
rect 172 174 380 184
rect 415 180 460 184
rect 463 183 464 184
rect 479 183 492 184
rect 339 170 387 174
rect 222 148 252 157
rect 315 150 330 157
rect 351 148 387 170
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 15 118 28 120
rect 43 118 77 120
rect 15 102 89 118
rect 116 114 129 128
rect 144 114 160 130
rect 206 125 217 138
rect -1 80 0 96
rect 15 80 28 102
rect 43 80 73 102
rect 116 98 178 114
rect 206 107 217 123
rect 222 118 232 138
rect 242 118 256 138
rect 259 125 268 138
rect 284 125 293 138
rect 222 107 256 118
rect 259 107 267 123
rect 284 107 293 123
rect 300 118 310 138
rect 320 118 334 138
rect 335 125 346 138
rect 300 107 334 118
rect 335 107 346 123
rect 392 114 408 130
rect 415 128 445 180
rect 479 176 480 183
rect 464 168 480 176
rect 451 136 464 155
rect 479 136 509 152
rect 451 120 525 136
rect 451 118 464 120
rect 479 118 513 120
rect 116 96 129 98
rect 144 96 178 98
rect 116 80 178 96
rect 222 91 235 94
rect 300 91 330 102
rect 378 98 424 114
rect 451 102 525 118
rect 378 96 412 98
rect 377 80 424 96
rect 451 80 464 102
rect 479 80 509 102
rect 536 80 537 96
rect 552 80 565 240
rect 595 136 608 240
rect 653 218 654 228
rect 669 218 682 228
rect 653 214 682 218
rect 687 214 717 240
rect 735 226 751 228
rect 823 226 876 240
rect 824 224 888 226
rect 735 214 750 218
rect 653 212 750 214
rect 637 204 688 212
rect 637 192 662 204
rect 669 192 688 204
rect 719 204 769 212
rect 719 196 735 204
rect 742 202 769 204
rect 778 204 793 208
rect 840 204 872 224
rect 931 212 946 240
rect 995 237 1025 240
rect 995 234 1031 237
rect 961 226 977 228
rect 962 214 977 218
rect 995 215 1034 234
rect 1053 228 1060 229
rect 1059 221 1060 228
rect 1043 218 1044 221
rect 1059 218 1072 221
rect 995 214 1025 215
rect 1034 214 1040 215
rect 1043 214 1072 218
rect 962 213 1072 214
rect 962 212 1078 213
rect 931 204 999 212
rect 778 202 847 204
rect 865 202 999 204
rect 742 198 814 202
rect 742 196 867 198
rect 742 192 814 196
rect 637 184 688 192
rect 735 188 814 192
rect 895 188 999 202
rect 1028 204 1078 212
rect 1028 195 1044 204
rect 735 184 999 188
rect 1025 192 1044 195
rect 1051 192 1078 204
rect 1025 184 1078 192
rect 653 176 654 184
rect 669 176 682 184
rect 653 168 669 176
rect 650 161 669 164
rect 650 152 672 161
rect 623 142 672 152
rect 623 136 653 142
rect 672 137 677 142
rect 595 120 669 136
rect 687 128 717 184
rect 752 174 960 184
rect 995 180 1040 184
rect 1043 183 1044 184
rect 1059 183 1072 184
rect 919 170 967 174
rect 802 148 832 157
rect 895 150 910 157
rect 931 148 967 170
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 595 118 608 120
rect 623 118 657 120
rect 595 102 669 118
rect 696 114 709 128
rect 724 114 740 130
rect 786 125 797 138
rect 579 80 580 96
rect 595 80 608 102
rect 623 80 653 102
rect 696 98 758 114
rect 786 107 797 123
rect 802 118 812 138
rect 822 118 836 138
rect 839 125 848 138
rect 864 125 873 138
rect 802 107 836 118
rect 839 107 847 123
rect 864 107 873 123
rect 880 118 890 138
rect 900 118 914 138
rect 915 125 926 138
rect 880 107 914 118
rect 915 107 926 123
rect 972 114 988 130
rect 995 128 1025 180
rect 1059 176 1060 183
rect 1044 168 1060 176
rect 1031 136 1044 155
rect 1059 136 1089 152
rect 1031 120 1105 136
rect 1031 118 1044 120
rect 1059 118 1093 120
rect 696 96 709 98
rect 724 96 758 98
rect 696 80 758 96
rect 802 91 815 94
rect 880 91 910 102
rect 958 98 1004 114
rect 1031 102 1105 118
rect 958 96 992 98
rect 957 80 1004 96
rect 1031 80 1044 102
rect 1059 80 1089 102
rect 1116 80 1117 96
rect 1132 80 1145 240
rect 1175 136 1188 240
rect 1233 218 1234 228
rect 1249 218 1262 228
rect 1233 214 1262 218
rect 1267 214 1297 240
rect 1315 226 1331 228
rect 1403 226 1456 240
rect 1404 224 1468 226
rect 1315 214 1330 218
rect 1233 212 1330 214
rect 1217 204 1268 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1299 204 1349 212
rect 1299 196 1315 204
rect 1322 202 1349 204
rect 1358 204 1373 208
rect 1420 204 1452 224
rect 1511 212 1526 240
rect 1575 237 1605 240
rect 1575 234 1611 237
rect 1541 226 1557 228
rect 1542 214 1557 218
rect 1575 215 1614 234
rect 1633 228 1640 229
rect 1639 221 1640 228
rect 1623 218 1624 221
rect 1639 218 1652 221
rect 1575 214 1605 215
rect 1614 214 1620 215
rect 1623 214 1652 218
rect 1542 213 1652 214
rect 1542 212 1658 213
rect 1511 204 1579 212
rect 1358 202 1427 204
rect 1445 202 1579 204
rect 1322 198 1394 202
rect 1322 196 1447 198
rect 1322 192 1394 196
rect 1217 184 1268 192
rect 1315 188 1394 192
rect 1475 188 1579 202
rect 1608 204 1658 212
rect 1608 195 1624 204
rect 1315 184 1579 188
rect 1605 192 1624 195
rect 1631 192 1658 204
rect 1605 184 1658 192
rect 1233 176 1234 184
rect 1249 176 1262 184
rect 1233 168 1249 176
rect 1230 161 1249 164
rect 1230 152 1252 161
rect 1203 142 1252 152
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1175 120 1249 136
rect 1267 128 1297 184
rect 1332 174 1540 184
rect 1575 180 1620 184
rect 1623 183 1624 184
rect 1639 183 1652 184
rect 1499 170 1547 174
rect 1382 148 1412 157
rect 1475 150 1490 157
rect 1511 148 1547 170
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1175 118 1188 120
rect 1203 118 1237 120
rect 1175 102 1249 118
rect 1276 114 1289 128
rect 1304 114 1320 130
rect 1366 125 1377 138
rect 1159 80 1160 96
rect 1175 80 1188 102
rect 1203 80 1233 102
rect 1276 98 1338 114
rect 1366 107 1377 123
rect 1382 118 1392 138
rect 1402 118 1416 138
rect 1419 125 1428 138
rect 1444 125 1453 138
rect 1382 107 1416 118
rect 1419 107 1427 123
rect 1444 107 1453 123
rect 1460 118 1470 138
rect 1480 118 1494 138
rect 1495 125 1506 138
rect 1460 107 1494 118
rect 1495 107 1506 123
rect 1552 114 1568 130
rect 1575 128 1605 180
rect 1639 176 1640 183
rect 1624 168 1640 176
rect 1611 136 1624 155
rect 1639 136 1669 152
rect 1611 120 1685 136
rect 1611 118 1624 120
rect 1639 118 1673 120
rect 1276 96 1289 98
rect 1304 96 1338 98
rect 1276 80 1338 96
rect 1382 91 1395 94
rect 1460 91 1490 102
rect 1538 98 1584 114
rect 1611 102 1685 118
rect 1538 96 1572 98
rect 1537 80 1584 96
rect 1611 80 1624 102
rect 1639 80 1669 102
rect 1696 80 1697 96
rect 1712 80 1725 240
rect 1755 136 1768 240
rect 1813 218 1814 228
rect 1829 218 1842 228
rect 1813 214 1842 218
rect 1847 214 1877 240
rect 1895 226 1911 228
rect 1983 226 2036 240
rect 1984 224 2048 226
rect 1895 214 1910 218
rect 1813 212 1910 214
rect 1797 204 1848 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1879 204 1929 212
rect 1879 196 1895 204
rect 1902 202 1929 204
rect 1938 204 1953 208
rect 2000 204 2032 224
rect 2091 212 2106 240
rect 2155 237 2185 240
rect 2155 234 2191 237
rect 2121 226 2137 228
rect 2122 214 2137 218
rect 2155 215 2194 234
rect 2213 228 2220 229
rect 2219 221 2220 228
rect 2203 218 2204 221
rect 2219 218 2232 221
rect 2155 214 2185 215
rect 2194 214 2200 215
rect 2203 214 2232 218
rect 2122 213 2232 214
rect 2122 212 2238 213
rect 2091 204 2159 212
rect 1938 202 2007 204
rect 2025 202 2159 204
rect 1902 198 1974 202
rect 1902 196 2027 198
rect 1902 192 1974 196
rect 1797 184 1848 192
rect 1895 188 1974 192
rect 2055 188 2159 202
rect 2188 204 2238 212
rect 2188 195 2204 204
rect 1895 184 2159 188
rect 2185 192 2204 195
rect 2211 192 2238 204
rect 2185 184 2238 192
rect 1813 176 1814 184
rect 1829 176 1842 184
rect 1813 168 1829 176
rect 1810 161 1829 164
rect 1810 152 1832 161
rect 1783 142 1832 152
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1755 120 1829 136
rect 1847 128 1877 184
rect 1912 174 2120 184
rect 2155 180 2200 184
rect 2203 183 2204 184
rect 2219 183 2232 184
rect 2079 170 2127 174
rect 1962 148 1992 157
rect 2055 150 2070 157
rect 2091 148 2127 170
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 1755 118 1768 120
rect 1783 118 1817 120
rect 1755 102 1829 118
rect 1856 114 1869 128
rect 1884 114 1900 130
rect 1946 125 1957 138
rect 1739 80 1740 96
rect 1755 80 1768 102
rect 1783 80 1813 102
rect 1856 98 1918 114
rect 1946 107 1957 123
rect 1962 118 1972 138
rect 1982 118 1996 138
rect 1999 125 2008 138
rect 2024 125 2033 138
rect 1962 107 1996 118
rect 1999 107 2007 123
rect 2024 107 2033 123
rect 2040 118 2050 138
rect 2060 118 2074 138
rect 2075 125 2086 138
rect 2040 107 2074 118
rect 2075 107 2086 123
rect 2132 114 2148 130
rect 2155 128 2185 180
rect 2219 176 2220 183
rect 2204 168 2220 176
rect 2191 136 2204 155
rect 2219 136 2249 152
rect 2191 120 2265 136
rect 2191 118 2204 120
rect 2219 118 2253 120
rect 1856 96 1869 98
rect 1884 96 1918 98
rect 1856 80 1918 96
rect 1962 91 1975 94
rect 2040 91 2070 102
rect 2118 98 2164 114
rect 2191 102 2265 118
rect 2118 96 2152 98
rect 2117 80 2164 96
rect 2191 80 2204 102
rect 2219 80 2249 102
rect 2276 80 2277 96
rect 2292 80 2305 240
rect 2335 136 2348 240
rect 2393 218 2394 228
rect 2409 218 2422 228
rect 2393 214 2422 218
rect 2427 214 2457 240
rect 2475 226 2491 228
rect 2563 226 2616 240
rect 2564 224 2628 226
rect 2475 214 2490 218
rect 2393 212 2490 214
rect 2377 204 2428 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2459 204 2509 212
rect 2459 196 2475 204
rect 2482 202 2509 204
rect 2518 204 2533 208
rect 2580 204 2612 224
rect 2671 212 2686 240
rect 2735 237 2765 240
rect 2735 234 2771 237
rect 2701 226 2717 228
rect 2702 214 2717 218
rect 2735 215 2774 234
rect 2793 228 2800 229
rect 2799 221 2800 228
rect 2783 218 2784 221
rect 2799 218 2812 221
rect 2735 214 2765 215
rect 2774 214 2780 215
rect 2783 214 2812 218
rect 2702 213 2812 214
rect 2702 212 2818 213
rect 2671 204 2739 212
rect 2518 202 2587 204
rect 2605 202 2739 204
rect 2482 198 2554 202
rect 2482 196 2607 198
rect 2482 192 2554 196
rect 2377 184 2428 192
rect 2475 188 2554 192
rect 2635 188 2739 202
rect 2768 204 2818 212
rect 2768 195 2784 204
rect 2475 184 2739 188
rect 2765 192 2784 195
rect 2791 192 2818 204
rect 2765 184 2818 192
rect 2393 176 2394 184
rect 2409 176 2422 184
rect 2393 168 2409 176
rect 2390 161 2409 164
rect 2390 152 2412 161
rect 2363 142 2412 152
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2335 120 2409 136
rect 2427 128 2457 184
rect 2492 174 2700 184
rect 2735 180 2780 184
rect 2783 183 2784 184
rect 2799 183 2812 184
rect 2659 170 2707 174
rect 2542 148 2572 157
rect 2635 150 2650 157
rect 2671 148 2707 170
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2335 118 2348 120
rect 2363 118 2397 120
rect 2335 102 2409 118
rect 2436 114 2449 128
rect 2464 114 2480 130
rect 2526 125 2537 138
rect 2319 80 2320 96
rect 2335 80 2348 102
rect 2363 80 2393 102
rect 2436 98 2498 114
rect 2526 107 2537 123
rect 2542 118 2552 138
rect 2562 118 2576 138
rect 2579 125 2588 138
rect 2604 125 2613 138
rect 2542 107 2576 118
rect 2579 107 2587 123
rect 2604 107 2613 123
rect 2620 118 2630 138
rect 2640 118 2654 138
rect 2655 125 2666 138
rect 2620 107 2654 118
rect 2655 107 2666 123
rect 2712 114 2728 130
rect 2735 128 2765 180
rect 2799 176 2800 183
rect 2784 168 2800 176
rect 2771 136 2784 155
rect 2799 136 2829 152
rect 2771 120 2845 136
rect 2771 118 2784 120
rect 2799 118 2833 120
rect 2436 96 2449 98
rect 2464 96 2498 98
rect 2436 80 2498 96
rect 2542 91 2555 94
rect 2620 91 2650 102
rect 2698 98 2744 114
rect 2771 102 2845 118
rect 2698 96 2732 98
rect 2697 80 2744 96
rect 2771 80 2784 102
rect 2799 80 2829 102
rect 2856 80 2857 96
rect 2872 80 2885 240
rect 2915 136 2928 240
rect 2973 218 2974 228
rect 2989 218 3002 228
rect 2973 214 3002 218
rect 3007 214 3037 240
rect 3055 226 3071 228
rect 3143 226 3196 240
rect 3144 224 3208 226
rect 3055 214 3070 218
rect 2973 212 3070 214
rect 2957 204 3008 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3039 204 3089 212
rect 3039 196 3055 204
rect 3062 202 3089 204
rect 3098 204 3113 208
rect 3160 204 3192 224
rect 3251 212 3266 240
rect 3315 237 3345 240
rect 3315 234 3351 237
rect 3281 226 3297 228
rect 3282 214 3297 218
rect 3315 215 3354 234
rect 3373 228 3380 229
rect 3379 221 3380 228
rect 3363 218 3364 221
rect 3379 218 3392 221
rect 3315 214 3345 215
rect 3354 214 3360 215
rect 3363 214 3392 218
rect 3282 213 3392 214
rect 3282 212 3398 213
rect 3251 204 3319 212
rect 3098 202 3167 204
rect 3185 202 3319 204
rect 3062 198 3134 202
rect 3062 196 3187 198
rect 3062 192 3134 196
rect 2957 184 3008 192
rect 3055 188 3134 192
rect 3215 188 3319 202
rect 3348 204 3398 212
rect 3348 195 3364 204
rect 3055 184 3319 188
rect 3345 192 3364 195
rect 3371 192 3398 204
rect 3345 184 3398 192
rect 2973 176 2974 184
rect 2989 176 3002 184
rect 2973 168 2989 176
rect 2970 161 2989 164
rect 2970 152 2992 161
rect 2943 142 2992 152
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2915 120 2989 136
rect 3007 128 3037 184
rect 3072 174 3280 184
rect 3315 180 3360 184
rect 3363 183 3364 184
rect 3379 183 3392 184
rect 3239 170 3287 174
rect 3122 148 3152 157
rect 3215 150 3230 157
rect 3251 148 3287 170
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 2915 118 2928 120
rect 2943 118 2977 120
rect 2915 102 2989 118
rect 3016 114 3029 128
rect 3044 114 3060 130
rect 3106 125 3117 138
rect 2899 80 2900 96
rect 2915 80 2928 102
rect 2943 80 2973 102
rect 3016 98 3078 114
rect 3106 107 3117 123
rect 3122 118 3132 138
rect 3142 118 3156 138
rect 3159 125 3168 138
rect 3184 125 3193 138
rect 3122 107 3156 118
rect 3159 107 3167 123
rect 3184 107 3193 123
rect 3200 118 3210 138
rect 3220 118 3234 138
rect 3235 125 3246 138
rect 3200 107 3234 118
rect 3235 107 3246 123
rect 3292 114 3308 130
rect 3315 128 3345 180
rect 3379 176 3380 183
rect 3364 168 3380 176
rect 3351 136 3364 155
rect 3379 136 3409 152
rect 3351 120 3425 136
rect 3351 118 3364 120
rect 3379 118 3413 120
rect 3016 96 3029 98
rect 3044 96 3078 98
rect 3016 80 3078 96
rect 3122 91 3135 94
rect 3200 91 3230 102
rect 3278 98 3324 114
rect 3351 102 3425 118
rect 3278 96 3312 98
rect 3277 80 3324 96
rect 3351 80 3364 102
rect 3379 80 3409 102
rect 3436 80 3437 96
rect 3452 80 3465 240
rect 3495 136 3508 240
rect 3553 218 3554 228
rect 3569 218 3582 228
rect 3553 214 3582 218
rect 3587 214 3617 240
rect 3635 226 3651 228
rect 3723 226 3776 240
rect 3724 224 3788 226
rect 3635 214 3650 218
rect 3553 212 3650 214
rect 3537 204 3588 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3619 204 3669 212
rect 3619 196 3635 204
rect 3642 202 3669 204
rect 3678 204 3693 208
rect 3740 204 3772 224
rect 3831 212 3846 240
rect 3895 237 3925 240
rect 3895 234 3931 237
rect 3861 226 3877 228
rect 3862 214 3877 218
rect 3895 215 3934 234
rect 3953 228 3960 229
rect 3959 221 3960 228
rect 3943 218 3944 221
rect 3959 218 3972 221
rect 3895 214 3925 215
rect 3934 214 3940 215
rect 3943 214 3972 218
rect 3862 213 3972 214
rect 3862 212 3978 213
rect 3831 204 3899 212
rect 3678 202 3747 204
rect 3765 202 3899 204
rect 3642 198 3714 202
rect 3642 196 3767 198
rect 3642 192 3714 196
rect 3537 184 3588 192
rect 3635 188 3714 192
rect 3795 188 3899 202
rect 3928 204 3978 212
rect 3928 195 3944 204
rect 3635 184 3899 188
rect 3925 192 3944 195
rect 3951 192 3978 204
rect 3925 184 3978 192
rect 3553 176 3554 184
rect 3569 176 3582 184
rect 3553 168 3569 176
rect 3550 161 3569 164
rect 3550 152 3572 161
rect 3523 142 3572 152
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3495 120 3569 136
rect 3587 128 3617 184
rect 3652 174 3860 184
rect 3895 180 3940 184
rect 3943 183 3944 184
rect 3959 183 3972 184
rect 3819 170 3867 174
rect 3702 148 3732 157
rect 3795 150 3810 157
rect 3831 148 3867 170
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3495 118 3508 120
rect 3523 118 3557 120
rect 3495 102 3569 118
rect 3596 114 3609 128
rect 3624 114 3640 130
rect 3686 125 3697 138
rect 3479 80 3480 96
rect 3495 80 3508 102
rect 3523 80 3553 102
rect 3596 98 3658 114
rect 3686 107 3697 123
rect 3702 118 3712 138
rect 3722 118 3736 138
rect 3739 125 3748 138
rect 3764 125 3773 138
rect 3702 107 3736 118
rect 3739 107 3747 123
rect 3764 107 3773 123
rect 3780 118 3790 138
rect 3800 118 3814 138
rect 3815 125 3826 138
rect 3780 107 3814 118
rect 3815 107 3826 123
rect 3872 114 3888 130
rect 3895 128 3925 180
rect 3959 176 3960 183
rect 3944 168 3960 176
rect 3931 136 3944 155
rect 3959 136 3989 152
rect 3931 120 4005 136
rect 3931 118 3944 120
rect 3959 118 3993 120
rect 3596 96 3609 98
rect 3624 96 3658 98
rect 3596 80 3658 96
rect 3702 91 3715 94
rect 3780 91 3810 102
rect 3858 98 3904 114
rect 3931 102 4005 118
rect 3858 96 3892 98
rect 3857 80 3904 96
rect 3931 80 3944 102
rect 3959 80 3989 102
rect 4016 80 4017 96
rect 4032 80 4045 240
rect 4075 136 4088 240
rect 4133 218 4134 228
rect 4149 218 4162 228
rect 4133 214 4162 218
rect 4167 214 4197 240
rect 4215 226 4231 228
rect 4303 226 4356 240
rect 4304 224 4368 226
rect 4215 214 4230 218
rect 4133 212 4230 214
rect 4117 204 4168 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4199 204 4249 212
rect 4199 196 4215 204
rect 4222 202 4249 204
rect 4258 204 4273 208
rect 4320 204 4352 224
rect 4411 212 4426 240
rect 4475 237 4505 240
rect 4475 234 4511 237
rect 4441 226 4457 228
rect 4442 214 4457 218
rect 4475 215 4514 234
rect 4533 228 4540 229
rect 4539 221 4540 228
rect 4523 218 4524 221
rect 4539 218 4552 221
rect 4475 214 4505 215
rect 4514 214 4520 215
rect 4523 214 4552 218
rect 4442 213 4552 214
rect 4442 212 4558 213
rect 4411 204 4479 212
rect 4258 202 4327 204
rect 4345 202 4479 204
rect 4222 198 4294 202
rect 4222 196 4347 198
rect 4222 192 4294 196
rect 4117 184 4168 192
rect 4215 188 4294 192
rect 4375 188 4479 202
rect 4508 204 4558 212
rect 4508 195 4524 204
rect 4215 184 4479 188
rect 4505 192 4524 195
rect 4531 192 4558 204
rect 4505 184 4558 192
rect 4133 176 4134 184
rect 4149 176 4162 184
rect 4133 168 4149 176
rect 4130 161 4149 164
rect 4130 152 4152 161
rect 4103 142 4152 152
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4075 120 4149 136
rect 4167 128 4197 184
rect 4232 174 4440 184
rect 4475 180 4520 184
rect 4523 183 4524 184
rect 4539 183 4552 184
rect 4399 170 4447 174
rect 4282 148 4312 157
rect 4375 150 4390 157
rect 4411 148 4447 170
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4075 118 4088 120
rect 4103 118 4137 120
rect 4075 102 4149 118
rect 4176 114 4189 128
rect 4204 114 4220 130
rect 4266 125 4277 138
rect 4059 80 4060 96
rect 4075 80 4088 102
rect 4103 80 4133 102
rect 4176 98 4238 114
rect 4266 107 4277 123
rect 4282 118 4292 138
rect 4302 118 4316 138
rect 4319 125 4328 138
rect 4344 125 4353 138
rect 4282 107 4316 118
rect 4319 107 4327 123
rect 4344 107 4353 123
rect 4360 118 4370 138
rect 4380 118 4394 138
rect 4395 125 4406 138
rect 4360 107 4394 118
rect 4395 107 4406 123
rect 4452 114 4468 130
rect 4475 128 4505 180
rect 4539 176 4540 183
rect 4524 168 4540 176
rect 4511 136 4524 155
rect 4539 136 4569 152
rect 4511 120 4585 136
rect 4511 118 4524 120
rect 4539 118 4573 120
rect 4176 96 4189 98
rect 4204 96 4238 98
rect 4176 80 4238 96
rect 4282 91 4295 94
rect 4360 91 4390 102
rect 4438 98 4484 114
rect 4511 102 4585 118
rect 4438 96 4472 98
rect 4437 80 4484 96
rect 4511 80 4524 102
rect 4539 80 4569 102
rect 4596 80 4597 96
rect 4612 80 4625 240
rect 4655 136 4668 240
rect 4713 218 4714 228
rect 4729 218 4742 228
rect 4713 214 4742 218
rect 4747 214 4777 240
rect 4795 226 4811 228
rect 4883 226 4936 240
rect 4884 224 4948 226
rect 4795 214 4810 218
rect 4713 212 4810 214
rect 4697 204 4748 212
rect 4697 192 4722 204
rect 4729 192 4748 204
rect 4779 204 4829 212
rect 4779 196 4795 204
rect 4802 202 4829 204
rect 4838 204 4853 208
rect 4900 204 4932 224
rect 4991 212 5006 240
rect 5055 237 5085 240
rect 5055 234 5091 237
rect 5021 226 5037 228
rect 5022 214 5037 218
rect 5055 215 5094 234
rect 5113 228 5120 229
rect 5119 221 5120 228
rect 5103 218 5104 221
rect 5119 218 5132 221
rect 5055 214 5085 215
rect 5094 214 5100 215
rect 5103 214 5132 218
rect 5022 213 5132 214
rect 5022 212 5138 213
rect 4991 204 5059 212
rect 4838 202 4907 204
rect 4925 202 5059 204
rect 4802 198 4874 202
rect 4802 196 4927 198
rect 4802 192 4874 196
rect 4697 184 4748 192
rect 4795 188 4874 192
rect 4955 188 5059 202
rect 5088 204 5138 212
rect 5088 195 5104 204
rect 4795 184 5059 188
rect 5085 192 5104 195
rect 5111 192 5138 204
rect 5085 184 5138 192
rect 4713 176 4714 184
rect 4729 176 4742 184
rect 4713 168 4729 176
rect 4710 161 4729 164
rect 4710 152 4732 161
rect 4683 142 4732 152
rect 4683 136 4713 142
rect 4732 137 4737 142
rect 4655 120 4729 136
rect 4747 128 4777 184
rect 4812 174 5020 184
rect 5055 180 5100 184
rect 5103 183 5104 184
rect 5119 183 5132 184
rect 4979 170 5027 174
rect 4862 148 4892 157
rect 4955 150 4970 157
rect 4991 148 5027 170
rect 4838 144 5027 148
rect 4853 141 5027 144
rect 4846 138 5027 141
rect 4655 118 4668 120
rect 4683 118 4717 120
rect 4655 102 4729 118
rect 4756 114 4769 128
rect 4784 114 4800 130
rect 4846 125 4857 138
rect 4639 80 4640 96
rect 4655 80 4668 102
rect 4683 80 4713 102
rect 4756 98 4818 114
rect 4846 107 4857 123
rect 4862 118 4872 138
rect 4882 118 4896 138
rect 4899 125 4908 138
rect 4924 125 4933 138
rect 4862 107 4896 118
rect 4899 107 4907 123
rect 4924 107 4933 123
rect 4940 118 4950 138
rect 4960 118 4974 138
rect 4975 125 4986 138
rect 4940 107 4974 118
rect 4975 107 4986 123
rect 5032 114 5048 130
rect 5055 128 5085 180
rect 5119 176 5120 183
rect 5104 168 5120 176
rect 5091 136 5104 155
rect 5119 136 5149 152
rect 5091 120 5165 136
rect 5091 118 5104 120
rect 5119 118 5153 120
rect 4756 96 4769 98
rect 4784 96 4818 98
rect 4756 80 4818 96
rect 4862 91 4875 94
rect 4940 91 4970 102
rect 5018 98 5064 114
rect 5091 102 5165 118
rect 5018 96 5052 98
rect 5017 80 5064 96
rect 5091 80 5104 102
rect 5119 80 5149 102
rect 5176 80 5177 96
rect 5192 80 5205 240
rect 5235 136 5248 240
rect 5293 218 5294 228
rect 5309 218 5322 228
rect 5293 214 5322 218
rect 5327 214 5357 240
rect 5375 226 5391 228
rect 5463 226 5516 240
rect 5464 224 5528 226
rect 5375 214 5390 218
rect 5293 212 5390 214
rect 5277 204 5328 212
rect 5277 192 5302 204
rect 5309 192 5328 204
rect 5359 204 5409 212
rect 5359 196 5375 204
rect 5382 202 5409 204
rect 5418 204 5433 208
rect 5480 204 5512 224
rect 5571 212 5586 240
rect 5635 237 5665 240
rect 5635 234 5671 237
rect 5601 226 5617 228
rect 5602 214 5617 218
rect 5635 215 5674 234
rect 5693 228 5700 229
rect 5699 221 5700 228
rect 5683 218 5684 221
rect 5699 218 5712 221
rect 5635 214 5665 215
rect 5674 214 5680 215
rect 5683 214 5712 218
rect 5602 213 5712 214
rect 5602 212 5718 213
rect 5571 204 5639 212
rect 5418 202 5487 204
rect 5505 202 5639 204
rect 5382 198 5454 202
rect 5382 196 5507 198
rect 5382 192 5454 196
rect 5277 184 5328 192
rect 5375 188 5454 192
rect 5535 188 5639 202
rect 5668 204 5718 212
rect 5668 195 5684 204
rect 5375 184 5639 188
rect 5665 192 5684 195
rect 5691 192 5718 204
rect 5665 184 5718 192
rect 5293 176 5294 184
rect 5309 176 5322 184
rect 5293 168 5309 176
rect 5290 161 5309 164
rect 5290 152 5312 161
rect 5263 142 5312 152
rect 5263 136 5293 142
rect 5312 137 5317 142
rect 5235 120 5309 136
rect 5327 128 5357 184
rect 5392 174 5600 184
rect 5635 180 5680 184
rect 5683 183 5684 184
rect 5699 183 5712 184
rect 5559 170 5607 174
rect 5442 148 5472 157
rect 5535 150 5550 157
rect 5571 148 5607 170
rect 5418 144 5607 148
rect 5433 141 5607 144
rect 5426 138 5607 141
rect 5235 118 5248 120
rect 5263 118 5297 120
rect 5235 102 5309 118
rect 5336 114 5349 128
rect 5364 114 5380 130
rect 5426 125 5437 138
rect 5219 80 5220 96
rect 5235 80 5248 102
rect 5263 80 5293 102
rect 5336 98 5398 114
rect 5426 107 5437 123
rect 5442 118 5452 138
rect 5462 118 5476 138
rect 5479 125 5488 138
rect 5504 125 5513 138
rect 5442 107 5476 118
rect 5479 107 5487 123
rect 5504 107 5513 123
rect 5520 118 5530 138
rect 5540 118 5554 138
rect 5555 125 5566 138
rect 5520 107 5554 118
rect 5555 107 5566 123
rect 5612 114 5628 130
rect 5635 128 5665 180
rect 5699 176 5700 183
rect 5684 168 5700 176
rect 5671 136 5684 155
rect 5699 136 5729 152
rect 5671 120 5745 136
rect 5671 118 5684 120
rect 5699 118 5733 120
rect 5336 96 5349 98
rect 5364 96 5398 98
rect 5336 80 5398 96
rect 5442 91 5455 94
rect 5520 91 5550 102
rect 5598 98 5644 114
rect 5671 102 5745 118
rect 5598 96 5632 98
rect 5597 80 5644 96
rect 5671 80 5684 102
rect 5699 80 5729 102
rect 5756 80 5757 96
rect 5772 80 5785 240
rect 5815 136 5828 240
rect 5873 218 5874 228
rect 5889 218 5902 228
rect 5873 214 5902 218
rect 5907 214 5937 240
rect 5955 226 5971 228
rect 6043 226 6096 240
rect 6044 224 6108 226
rect 5955 214 5970 218
rect 5873 212 5970 214
rect 5857 204 5908 212
rect 5857 192 5882 204
rect 5889 192 5908 204
rect 5939 204 5989 212
rect 5939 196 5955 204
rect 5962 202 5989 204
rect 5998 204 6013 208
rect 6060 204 6092 224
rect 6151 212 6166 240
rect 6215 237 6245 240
rect 6215 234 6251 237
rect 6181 226 6197 228
rect 6182 214 6197 218
rect 6215 215 6254 234
rect 6273 228 6280 229
rect 6279 221 6280 228
rect 6263 218 6264 221
rect 6279 218 6292 221
rect 6215 214 6245 215
rect 6254 214 6260 215
rect 6263 214 6292 218
rect 6182 213 6292 214
rect 6182 212 6298 213
rect 6151 204 6219 212
rect 5998 202 6067 204
rect 6085 202 6219 204
rect 5962 198 6034 202
rect 5962 196 6087 198
rect 5962 192 6034 196
rect 5857 184 5908 192
rect 5955 188 6034 192
rect 6115 188 6219 202
rect 6248 204 6298 212
rect 6248 195 6264 204
rect 5955 184 6219 188
rect 6245 192 6264 195
rect 6271 192 6298 204
rect 6245 184 6298 192
rect 5873 176 5874 184
rect 5889 176 5902 184
rect 5873 168 5889 176
rect 5870 161 5889 164
rect 5870 152 5892 161
rect 5843 142 5892 152
rect 5843 136 5873 142
rect 5892 137 5897 142
rect 5815 120 5889 136
rect 5907 128 5937 184
rect 5972 174 6180 184
rect 6215 180 6260 184
rect 6263 183 6264 184
rect 6279 183 6292 184
rect 6139 170 6187 174
rect 6022 148 6052 157
rect 6115 150 6130 157
rect 6151 148 6187 170
rect 5998 144 6187 148
rect 6013 141 6187 144
rect 6006 138 6187 141
rect 5815 118 5828 120
rect 5843 118 5877 120
rect 5815 102 5889 118
rect 5916 114 5929 128
rect 5944 114 5960 130
rect 6006 125 6017 138
rect 5799 80 5800 96
rect 5815 80 5828 102
rect 5843 80 5873 102
rect 5916 98 5978 114
rect 6006 107 6017 123
rect 6022 118 6032 138
rect 6042 118 6056 138
rect 6059 125 6068 138
rect 6084 125 6093 138
rect 6022 107 6056 118
rect 6059 107 6067 123
rect 6084 107 6093 123
rect 6100 118 6110 138
rect 6120 118 6134 138
rect 6135 125 6146 138
rect 6100 107 6134 118
rect 6135 107 6146 123
rect 6192 114 6208 130
rect 6215 128 6245 180
rect 6279 176 6280 183
rect 6264 168 6280 176
rect 6251 136 6264 155
rect 6279 136 6309 152
rect 6251 120 6325 136
rect 6251 118 6264 120
rect 6279 118 6313 120
rect 5916 96 5929 98
rect 5944 96 5978 98
rect 5916 80 5978 96
rect 6022 91 6035 94
rect 6100 91 6130 102
rect 6178 98 6224 114
rect 6251 102 6325 118
rect 6178 96 6212 98
rect 6177 80 6224 96
rect 6251 80 6264 102
rect 6279 80 6309 102
rect 6336 80 6337 96
rect 6352 80 6365 240
rect 6395 136 6408 240
rect 6453 218 6454 228
rect 6469 218 6482 228
rect 6453 214 6482 218
rect 6487 214 6517 240
rect 6535 226 6551 228
rect 6623 226 6676 240
rect 6624 224 6688 226
rect 6535 214 6550 218
rect 6453 212 6550 214
rect 6437 204 6488 212
rect 6437 192 6462 204
rect 6469 192 6488 204
rect 6519 204 6569 212
rect 6519 196 6535 204
rect 6542 202 6569 204
rect 6578 204 6593 208
rect 6640 204 6672 224
rect 6731 212 6746 240
rect 6795 237 6825 240
rect 6795 234 6831 237
rect 6761 226 6777 228
rect 6762 214 6777 218
rect 6795 215 6834 234
rect 6853 228 6860 229
rect 6859 221 6860 228
rect 6843 218 6844 221
rect 6859 218 6872 221
rect 6795 214 6825 215
rect 6834 214 6840 215
rect 6843 214 6872 218
rect 6762 213 6872 214
rect 6762 212 6878 213
rect 6731 204 6799 212
rect 6578 202 6647 204
rect 6665 202 6799 204
rect 6542 198 6614 202
rect 6542 196 6667 198
rect 6542 192 6614 196
rect 6437 184 6488 192
rect 6535 188 6614 192
rect 6695 188 6799 202
rect 6828 204 6878 212
rect 6828 195 6844 204
rect 6535 184 6799 188
rect 6825 192 6844 195
rect 6851 192 6878 204
rect 6825 184 6878 192
rect 6453 176 6454 184
rect 6469 176 6482 184
rect 6453 168 6469 176
rect 6450 161 6469 164
rect 6450 152 6472 161
rect 6423 142 6472 152
rect 6423 136 6453 142
rect 6472 137 6477 142
rect 6395 120 6469 136
rect 6487 128 6517 184
rect 6552 174 6760 184
rect 6795 180 6840 184
rect 6843 183 6844 184
rect 6859 183 6872 184
rect 6719 170 6767 174
rect 6602 148 6632 157
rect 6695 150 6710 157
rect 6731 148 6767 170
rect 6578 144 6767 148
rect 6593 141 6767 144
rect 6586 138 6767 141
rect 6395 118 6408 120
rect 6423 118 6457 120
rect 6395 102 6469 118
rect 6496 114 6509 128
rect 6524 114 6540 130
rect 6586 125 6597 138
rect 6379 80 6380 96
rect 6395 80 6408 102
rect 6423 80 6453 102
rect 6496 98 6558 114
rect 6586 107 6597 123
rect 6602 118 6612 138
rect 6622 118 6636 138
rect 6639 125 6648 138
rect 6664 125 6673 138
rect 6602 107 6636 118
rect 6639 107 6647 123
rect 6664 107 6673 123
rect 6680 118 6690 138
rect 6700 118 6714 138
rect 6715 125 6726 138
rect 6680 107 6714 118
rect 6715 107 6726 123
rect 6772 114 6788 130
rect 6795 128 6825 180
rect 6859 176 6860 183
rect 6844 168 6860 176
rect 6831 136 6844 155
rect 6859 136 6889 152
rect 6831 120 6905 136
rect 6831 118 6844 120
rect 6859 118 6893 120
rect 6496 96 6509 98
rect 6524 96 6558 98
rect 6496 80 6558 96
rect 6602 91 6615 94
rect 6680 91 6710 102
rect 6758 98 6804 114
rect 6831 102 6905 118
rect 6758 96 6792 98
rect 6757 80 6804 96
rect 6831 80 6844 102
rect 6859 80 6889 102
rect 6916 80 6917 96
rect 6932 80 6945 240
rect 6975 136 6988 240
rect 7033 218 7034 228
rect 7049 218 7062 228
rect 7033 214 7062 218
rect 7067 214 7097 240
rect 7115 226 7131 228
rect 7203 226 7256 240
rect 7204 224 7268 226
rect 7115 214 7130 218
rect 7033 212 7130 214
rect 7017 204 7068 212
rect 7017 192 7042 204
rect 7049 192 7068 204
rect 7099 204 7149 212
rect 7099 196 7115 204
rect 7122 202 7149 204
rect 7158 204 7173 208
rect 7220 204 7252 224
rect 7311 212 7326 240
rect 7375 237 7405 240
rect 7375 234 7411 237
rect 7341 226 7357 228
rect 7342 214 7357 218
rect 7375 215 7414 234
rect 7433 228 7440 229
rect 7439 221 7440 228
rect 7423 218 7424 221
rect 7439 218 7452 221
rect 7375 214 7405 215
rect 7414 214 7420 215
rect 7423 214 7452 218
rect 7342 213 7452 214
rect 7342 212 7458 213
rect 7311 204 7379 212
rect 7158 202 7227 204
rect 7245 202 7379 204
rect 7122 198 7194 202
rect 7122 196 7247 198
rect 7122 192 7194 196
rect 7017 184 7068 192
rect 7115 188 7194 192
rect 7275 188 7379 202
rect 7408 204 7458 212
rect 7408 195 7424 204
rect 7115 184 7379 188
rect 7405 192 7424 195
rect 7431 192 7458 204
rect 7405 184 7458 192
rect 7033 176 7034 184
rect 7049 176 7062 184
rect 7033 168 7049 176
rect 7030 161 7049 164
rect 7030 152 7052 161
rect 7003 142 7052 152
rect 7003 136 7033 142
rect 7052 137 7057 142
rect 6975 120 7049 136
rect 7067 128 7097 184
rect 7132 174 7340 184
rect 7375 180 7420 184
rect 7423 183 7424 184
rect 7439 183 7452 184
rect 7299 170 7347 174
rect 7182 148 7212 157
rect 7275 150 7290 157
rect 7311 148 7347 170
rect 7158 144 7347 148
rect 7173 141 7347 144
rect 7166 138 7347 141
rect 6975 118 6988 120
rect 7003 118 7037 120
rect 6975 102 7049 118
rect 7076 114 7089 128
rect 7104 114 7120 130
rect 7166 125 7177 138
rect 6959 80 6960 96
rect 6975 80 6988 102
rect 7003 80 7033 102
rect 7076 98 7138 114
rect 7166 107 7177 123
rect 7182 118 7192 138
rect 7202 118 7216 138
rect 7219 125 7228 138
rect 7244 125 7253 138
rect 7182 107 7216 118
rect 7219 107 7227 123
rect 7244 107 7253 123
rect 7260 118 7270 138
rect 7280 118 7294 138
rect 7295 125 7306 138
rect 7260 107 7294 118
rect 7295 107 7306 123
rect 7352 114 7368 130
rect 7375 128 7405 180
rect 7439 176 7440 183
rect 7424 168 7440 176
rect 7411 136 7424 155
rect 7439 136 7469 152
rect 7411 120 7485 136
rect 7411 118 7424 120
rect 7439 118 7473 120
rect 7076 96 7089 98
rect 7104 96 7138 98
rect 7076 80 7138 96
rect 7182 91 7195 94
rect 7260 91 7290 102
rect 7338 98 7384 114
rect 7411 102 7485 118
rect 7338 96 7372 98
rect 7337 80 7384 96
rect 7411 80 7424 102
rect 7439 80 7469 102
rect 7496 80 7497 96
rect 7512 80 7525 240
rect 7555 136 7568 240
rect 7613 218 7614 228
rect 7629 218 7642 228
rect 7613 214 7642 218
rect 7647 214 7677 240
rect 7695 226 7711 228
rect 7783 226 7836 240
rect 7784 224 7848 226
rect 7695 214 7710 218
rect 7613 212 7710 214
rect 7597 204 7648 212
rect 7597 192 7622 204
rect 7629 192 7648 204
rect 7679 204 7729 212
rect 7679 196 7695 204
rect 7702 202 7729 204
rect 7738 204 7753 208
rect 7800 204 7832 224
rect 7891 212 7906 240
rect 7955 237 7985 240
rect 7955 234 7991 237
rect 7921 226 7937 228
rect 7922 214 7937 218
rect 7955 215 7994 234
rect 8013 228 8020 229
rect 8019 221 8020 228
rect 8003 218 8004 221
rect 8019 218 8032 221
rect 7955 214 7985 215
rect 7994 214 8000 215
rect 8003 214 8032 218
rect 7922 213 8032 214
rect 7922 212 8038 213
rect 7891 204 7959 212
rect 7738 202 7807 204
rect 7825 202 7959 204
rect 7702 198 7774 202
rect 7702 196 7827 198
rect 7702 192 7774 196
rect 7597 184 7648 192
rect 7695 188 7774 192
rect 7855 188 7959 202
rect 7988 204 8038 212
rect 7988 195 8004 204
rect 7695 184 7959 188
rect 7985 192 8004 195
rect 8011 192 8038 204
rect 7985 184 8038 192
rect 7613 176 7614 184
rect 7629 176 7642 184
rect 7613 168 7629 176
rect 7610 161 7629 164
rect 7610 152 7632 161
rect 7583 142 7632 152
rect 7583 136 7613 142
rect 7632 137 7637 142
rect 7555 120 7629 136
rect 7647 128 7677 184
rect 7712 174 7920 184
rect 7955 180 8000 184
rect 8003 183 8004 184
rect 8019 183 8032 184
rect 7879 170 7927 174
rect 7762 148 7792 157
rect 7855 150 7870 157
rect 7891 148 7927 170
rect 7738 144 7927 148
rect 7753 141 7927 144
rect 7746 138 7927 141
rect 7555 118 7568 120
rect 7583 118 7617 120
rect 7555 102 7629 118
rect 7656 114 7669 128
rect 7684 114 7700 130
rect 7746 125 7757 138
rect 7539 80 7540 96
rect 7555 80 7568 102
rect 7583 80 7613 102
rect 7656 98 7718 114
rect 7746 107 7757 123
rect 7762 118 7772 138
rect 7782 118 7796 138
rect 7799 125 7808 138
rect 7824 125 7833 138
rect 7762 107 7796 118
rect 7799 107 7807 123
rect 7824 107 7833 123
rect 7840 118 7850 138
rect 7860 118 7874 138
rect 7875 125 7886 138
rect 7840 107 7874 118
rect 7875 107 7886 123
rect 7932 114 7948 130
rect 7955 128 7985 180
rect 8019 176 8020 183
rect 8004 168 8020 176
rect 7991 136 8004 155
rect 8019 136 8049 152
rect 7991 120 8065 136
rect 7991 118 8004 120
rect 8019 118 8053 120
rect 7656 96 7669 98
rect 7684 96 7718 98
rect 7656 80 7718 96
rect 7762 91 7775 94
rect 7840 91 7870 102
rect 7918 98 7964 114
rect 7991 102 8065 118
rect 7918 96 7952 98
rect 7917 80 7964 96
rect 7991 80 8004 102
rect 8019 80 8049 102
rect 8076 80 8077 96
rect 8092 80 8105 240
rect 8135 136 8148 240
rect 8193 218 8194 228
rect 8209 218 8222 228
rect 8193 214 8222 218
rect 8227 214 8257 240
rect 8275 226 8291 228
rect 8363 226 8416 240
rect 8364 224 8428 226
rect 8275 214 8290 218
rect 8193 212 8290 214
rect 8177 204 8228 212
rect 8177 192 8202 204
rect 8209 192 8228 204
rect 8259 204 8309 212
rect 8259 196 8275 204
rect 8282 202 8309 204
rect 8318 204 8333 208
rect 8380 204 8412 224
rect 8471 212 8486 240
rect 8535 237 8565 240
rect 8535 234 8571 237
rect 8501 226 8517 228
rect 8502 214 8517 218
rect 8535 215 8574 234
rect 8593 228 8600 229
rect 8599 221 8600 228
rect 8583 218 8584 221
rect 8599 218 8612 221
rect 8535 214 8565 215
rect 8574 214 8580 215
rect 8583 214 8612 218
rect 8502 213 8612 214
rect 8502 212 8618 213
rect 8471 204 8539 212
rect 8318 202 8387 204
rect 8405 202 8539 204
rect 8282 198 8354 202
rect 8282 196 8407 198
rect 8282 192 8354 196
rect 8177 184 8228 192
rect 8275 188 8354 192
rect 8435 188 8539 202
rect 8568 204 8618 212
rect 8568 195 8584 204
rect 8275 184 8539 188
rect 8565 192 8584 195
rect 8591 192 8618 204
rect 8565 184 8618 192
rect 8193 176 8194 184
rect 8209 176 8222 184
rect 8193 168 8209 176
rect 8190 161 8209 164
rect 8190 152 8212 161
rect 8163 142 8212 152
rect 8163 136 8193 142
rect 8212 137 8217 142
rect 8135 120 8209 136
rect 8227 128 8257 184
rect 8292 174 8500 184
rect 8535 180 8580 184
rect 8583 183 8584 184
rect 8599 183 8612 184
rect 8459 170 8507 174
rect 8342 148 8372 157
rect 8435 150 8450 157
rect 8471 148 8507 170
rect 8318 144 8507 148
rect 8333 141 8507 144
rect 8326 138 8507 141
rect 8135 118 8148 120
rect 8163 118 8197 120
rect 8135 102 8209 118
rect 8236 114 8249 128
rect 8264 114 8280 130
rect 8326 125 8337 138
rect 8119 80 8120 96
rect 8135 80 8148 102
rect 8163 80 8193 102
rect 8236 98 8298 114
rect 8326 107 8337 123
rect 8342 118 8352 138
rect 8362 118 8376 138
rect 8379 125 8388 138
rect 8404 125 8413 138
rect 8342 107 8376 118
rect 8379 107 8387 123
rect 8404 107 8413 123
rect 8420 118 8430 138
rect 8440 118 8454 138
rect 8455 125 8466 138
rect 8420 107 8454 118
rect 8455 107 8466 123
rect 8512 114 8528 130
rect 8535 128 8565 180
rect 8599 176 8600 183
rect 8584 168 8600 176
rect 8571 136 8584 155
rect 8599 136 8629 152
rect 8571 120 8645 136
rect 8571 118 8584 120
rect 8599 118 8633 120
rect 8236 96 8249 98
rect 8264 96 8298 98
rect 8236 80 8298 96
rect 8342 91 8355 94
rect 8420 91 8450 102
rect 8498 98 8544 114
rect 8571 102 8645 118
rect 8498 96 8532 98
rect 8497 80 8544 96
rect 8571 80 8584 102
rect 8599 80 8629 102
rect 8656 80 8657 96
rect 8672 80 8685 240
rect 8715 136 8728 240
rect 8773 218 8774 228
rect 8789 218 8802 228
rect 8773 214 8802 218
rect 8807 214 8837 240
rect 8855 226 8871 228
rect 8943 226 8996 240
rect 8944 224 9008 226
rect 8855 214 8870 218
rect 8773 212 8870 214
rect 8757 204 8808 212
rect 8757 192 8782 204
rect 8789 192 8808 204
rect 8839 204 8889 212
rect 8839 196 8855 204
rect 8862 202 8889 204
rect 8898 204 8913 208
rect 8960 204 8992 224
rect 9051 212 9066 240
rect 9115 237 9145 240
rect 9115 234 9151 237
rect 9081 226 9097 228
rect 9082 214 9097 218
rect 9115 215 9154 234
rect 9173 228 9180 229
rect 9179 221 9180 228
rect 9163 218 9164 221
rect 9179 218 9192 221
rect 9115 214 9145 215
rect 9154 214 9160 215
rect 9163 214 9192 218
rect 9082 213 9192 214
rect 9082 212 9198 213
rect 9051 204 9119 212
rect 8898 202 8967 204
rect 8985 202 9119 204
rect 8862 198 8934 202
rect 8862 196 8987 198
rect 8862 192 8934 196
rect 8757 184 8808 192
rect 8855 188 8934 192
rect 9015 188 9119 202
rect 9148 204 9198 212
rect 9148 195 9164 204
rect 8855 184 9119 188
rect 9145 192 9164 195
rect 9171 192 9198 204
rect 9145 184 9198 192
rect 8773 176 8774 184
rect 8789 176 8802 184
rect 8773 168 8789 176
rect 8770 161 8789 164
rect 8770 152 8792 161
rect 8743 142 8792 152
rect 8743 136 8773 142
rect 8792 137 8797 142
rect 8715 120 8789 136
rect 8807 128 8837 184
rect 8872 174 9080 184
rect 9115 180 9160 184
rect 9163 183 9164 184
rect 9179 183 9192 184
rect 9039 170 9087 174
rect 8922 148 8952 157
rect 9015 150 9030 157
rect 9051 148 9087 170
rect 8898 144 9087 148
rect 8913 141 9087 144
rect 8906 138 9087 141
rect 8715 118 8728 120
rect 8743 118 8777 120
rect 8715 102 8789 118
rect 8816 114 8829 128
rect 8844 114 8860 130
rect 8906 125 8917 138
rect 8699 80 8700 96
rect 8715 80 8728 102
rect 8743 80 8773 102
rect 8816 98 8878 114
rect 8906 107 8917 123
rect 8922 118 8932 138
rect 8942 118 8956 138
rect 8959 125 8968 138
rect 8984 125 8993 138
rect 8922 107 8956 118
rect 8959 107 8967 123
rect 8984 107 8993 123
rect 9000 118 9010 138
rect 9020 118 9034 138
rect 9035 125 9046 138
rect 9000 107 9034 118
rect 9035 107 9046 123
rect 9092 114 9108 130
rect 9115 128 9145 180
rect 9179 176 9180 183
rect 9164 168 9180 176
rect 9151 136 9164 155
rect 9179 136 9209 152
rect 9151 120 9225 136
rect 9151 118 9164 120
rect 9179 118 9213 120
rect 8816 96 8829 98
rect 8844 96 8878 98
rect 8816 80 8878 96
rect 8922 91 8935 94
rect 9000 91 9030 102
rect 9078 98 9124 114
rect 9151 102 9225 118
rect 9078 96 9112 98
rect 9077 80 9124 96
rect 9151 80 9164 102
rect 9179 80 9209 102
rect 9236 80 9237 96
rect 9252 80 9265 240
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 160 80
rect 172 68 247 80
rect 305 68 380 80
rect 392 68 423 80
rect 429 68 464 80
rect 98 66 260 68
rect -7 38 34 46
rect 116 38 129 66
rect 144 64 159 66
rect 183 39 190 46
rect 193 38 260 66
rect 292 66 464 68
rect 262 44 290 48
rect 292 44 372 66
rect 393 64 408 66
rect 262 42 372 44
rect 262 38 290 42
rect 292 38 372 42
rect -1 28 0 38
rect 15 28 28 38
rect 43 28 73 38
rect 116 28 159 38
rect 166 28 174 38
rect 193 30 196 38
rect 260 30 292 38
rect 193 28 359 30
rect 378 28 389 38
rect 393 28 423 38
rect 451 28 464 66
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 740 80
rect 752 68 827 80
rect 885 68 960 80
rect 972 68 1003 80
rect 1009 68 1044 80
rect 678 66 840 68
rect 573 38 614 46
rect 696 38 709 66
rect 724 64 739 66
rect 763 39 770 46
rect 773 38 840 66
rect 872 66 1044 68
rect 842 44 870 48
rect 872 44 952 66
rect 973 64 988 66
rect 842 42 952 44
rect 842 38 870 42
rect 872 38 952 42
rect 479 28 509 38
rect 536 28 537 38
rect 552 28 565 38
rect 579 28 580 38
rect 595 28 608 38
rect 623 28 653 38
rect 696 28 739 38
rect 746 28 754 38
rect 773 30 776 38
rect 840 30 872 38
rect 773 28 939 30
rect 958 28 969 38
rect 973 28 1003 38
rect 1031 28 1044 66
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1320 80
rect 1332 68 1407 80
rect 1465 68 1540 80
rect 1552 68 1583 80
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1153 38 1194 46
rect 1276 38 1289 66
rect 1304 64 1319 66
rect 1343 39 1350 46
rect 1353 38 1420 66
rect 1452 66 1624 68
rect 1422 44 1450 48
rect 1452 44 1532 66
rect 1553 64 1568 66
rect 1422 42 1532 44
rect 1422 38 1450 42
rect 1452 38 1532 42
rect 1059 28 1089 38
rect 1116 28 1117 38
rect 1132 28 1145 38
rect 1159 28 1160 38
rect 1175 28 1188 38
rect 1203 28 1233 38
rect 1276 28 1319 38
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1420 30 1452 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1553 28 1583 38
rect 1611 28 1624 66
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1900 80
rect 1912 68 1987 80
rect 2045 68 2120 80
rect 2132 68 2163 80
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1733 38 1774 46
rect 1856 38 1869 66
rect 1884 64 1899 66
rect 1923 39 1930 46
rect 1933 38 2000 66
rect 2032 66 2204 68
rect 2002 44 2030 48
rect 2032 44 2112 66
rect 2133 64 2148 66
rect 2002 42 2112 44
rect 2002 38 2030 42
rect 2032 38 2112 42
rect 1639 28 1669 38
rect 1696 28 1697 38
rect 1712 28 1725 38
rect 1739 28 1740 38
rect 1755 28 1768 38
rect 1783 28 1813 38
rect 1856 28 1899 38
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 2000 30 2032 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2133 28 2163 38
rect 2191 28 2204 66
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2480 80
rect 2492 68 2567 80
rect 2625 68 2700 80
rect 2712 68 2743 80
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2313 38 2354 46
rect 2436 38 2449 66
rect 2464 64 2479 66
rect 2503 39 2510 46
rect 2513 38 2580 66
rect 2612 66 2784 68
rect 2582 44 2610 48
rect 2612 44 2692 66
rect 2713 64 2728 66
rect 2582 42 2692 44
rect 2582 38 2610 42
rect 2612 38 2692 42
rect 2219 28 2249 38
rect 2276 28 2277 38
rect 2292 28 2305 38
rect 2319 28 2320 38
rect 2335 28 2348 38
rect 2363 28 2393 38
rect 2436 28 2479 38
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2580 30 2612 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2713 28 2743 38
rect 2771 28 2784 66
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3060 80
rect 3072 68 3147 80
rect 3205 68 3280 80
rect 3292 68 3323 80
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 2893 38 2934 46
rect 3016 38 3029 66
rect 3044 64 3059 66
rect 3083 39 3090 46
rect 3093 38 3160 66
rect 3192 66 3364 68
rect 3162 44 3190 48
rect 3192 44 3272 66
rect 3293 64 3308 66
rect 3162 42 3272 44
rect 3162 38 3190 42
rect 3192 38 3272 42
rect 2799 28 2829 38
rect 2856 28 2857 38
rect 2872 28 2885 38
rect 2899 28 2900 38
rect 2915 28 2928 38
rect 2943 28 2973 38
rect 3016 28 3059 38
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3160 30 3192 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3293 28 3323 38
rect 3351 28 3364 66
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3640 80
rect 3652 68 3727 80
rect 3785 68 3860 80
rect 3872 68 3903 80
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3473 38 3514 46
rect 3596 38 3609 66
rect 3624 64 3639 66
rect 3663 39 3670 46
rect 3673 38 3740 66
rect 3772 66 3944 68
rect 3742 44 3770 48
rect 3772 44 3852 66
rect 3873 64 3888 66
rect 3742 42 3852 44
rect 3742 38 3770 42
rect 3772 38 3852 42
rect 3379 28 3409 38
rect 3436 28 3437 38
rect 3452 28 3465 38
rect 3479 28 3480 38
rect 3495 28 3508 38
rect 3523 28 3553 38
rect 3596 28 3639 38
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3740 30 3772 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3873 28 3903 38
rect 3931 28 3944 66
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4220 80
rect 4232 68 4307 80
rect 4365 68 4440 80
rect 4452 68 4483 80
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4053 38 4094 46
rect 4176 38 4189 66
rect 4204 64 4219 66
rect 4243 39 4250 46
rect 4253 38 4320 66
rect 4352 66 4524 68
rect 4322 44 4350 48
rect 4352 44 4432 66
rect 4453 64 4468 66
rect 4322 42 4432 44
rect 4322 38 4350 42
rect 4352 38 4432 42
rect 3959 28 3989 38
rect 4016 28 4017 38
rect 4032 28 4045 38
rect 4059 28 4060 38
rect 4075 28 4088 38
rect 4103 28 4133 38
rect 4176 28 4219 38
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4320 30 4352 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4453 28 4483 38
rect 4511 28 4524 66
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4633 72 4674 80
rect 4633 46 4648 72
rect 4655 46 4674 72
rect 4738 68 4800 80
rect 4812 68 4887 80
rect 4945 68 5020 80
rect 5032 68 5063 80
rect 5069 68 5104 80
rect 4738 66 4900 68
rect 4633 38 4674 46
rect 4756 38 4769 66
rect 4784 64 4799 66
rect 4823 39 4830 46
rect 4833 38 4900 66
rect 4932 66 5104 68
rect 4902 44 4930 48
rect 4932 44 5012 66
rect 5033 64 5048 66
rect 4902 42 5012 44
rect 4902 38 4930 42
rect 4932 38 5012 42
rect 4539 28 4569 38
rect 4596 28 4597 38
rect 4612 28 4625 38
rect 4639 28 4640 38
rect 4655 28 4668 38
rect 4683 28 4713 38
rect 4756 28 4799 38
rect 4806 28 4814 38
rect 4833 30 4836 38
rect 4900 30 4932 38
rect 4833 28 4999 30
rect 5018 28 5029 38
rect 5033 28 5063 38
rect 5091 28 5104 66
rect 5176 72 5211 80
rect 5176 46 5177 72
rect 5184 46 5211 72
rect 5176 38 5211 46
rect 5213 72 5254 80
rect 5213 46 5228 72
rect 5235 46 5254 72
rect 5318 68 5380 80
rect 5392 68 5467 80
rect 5525 68 5600 80
rect 5612 68 5643 80
rect 5649 68 5684 80
rect 5318 66 5480 68
rect 5213 38 5254 46
rect 5336 38 5349 66
rect 5364 64 5379 66
rect 5403 39 5410 46
rect 5413 38 5480 66
rect 5512 66 5684 68
rect 5482 44 5510 48
rect 5512 44 5592 66
rect 5613 64 5628 66
rect 5482 42 5592 44
rect 5482 38 5510 42
rect 5512 38 5592 42
rect 5119 28 5149 38
rect 5176 28 5177 38
rect 5192 28 5205 38
rect 5219 28 5220 38
rect 5235 28 5248 38
rect 5263 28 5293 38
rect 5336 28 5379 38
rect 5386 28 5394 38
rect 5413 30 5416 38
rect 5480 30 5512 38
rect 5413 28 5579 30
rect 5598 28 5609 38
rect 5613 28 5643 38
rect 5671 28 5684 66
rect 5756 72 5791 80
rect 5756 46 5757 72
rect 5764 46 5791 72
rect 5756 38 5791 46
rect 5793 72 5834 80
rect 5793 46 5808 72
rect 5815 46 5834 72
rect 5898 68 5960 80
rect 5972 68 6047 80
rect 6105 68 6180 80
rect 6192 68 6223 80
rect 6229 68 6264 80
rect 5898 66 6060 68
rect 5793 38 5834 46
rect 5916 38 5929 66
rect 5944 64 5959 66
rect 5983 39 5990 46
rect 5993 38 6060 66
rect 6092 66 6264 68
rect 6062 44 6090 48
rect 6092 44 6172 66
rect 6193 64 6208 66
rect 6062 42 6172 44
rect 6062 38 6090 42
rect 6092 38 6172 42
rect 5699 28 5729 38
rect 5756 28 5757 38
rect 5772 28 5785 38
rect 5799 28 5800 38
rect 5815 28 5828 38
rect 5843 28 5873 38
rect 5916 28 5959 38
rect 5966 28 5974 38
rect 5993 30 5996 38
rect 6060 30 6092 38
rect 5993 28 6159 30
rect 6178 28 6189 38
rect 6193 28 6223 38
rect 6251 28 6264 66
rect 6336 72 6371 80
rect 6336 46 6337 72
rect 6344 46 6371 72
rect 6336 38 6371 46
rect 6373 72 6414 80
rect 6373 46 6388 72
rect 6395 46 6414 72
rect 6478 68 6540 80
rect 6552 68 6627 80
rect 6685 68 6760 80
rect 6772 68 6803 80
rect 6809 68 6844 80
rect 6478 66 6640 68
rect 6373 38 6414 46
rect 6496 38 6509 66
rect 6524 64 6539 66
rect 6563 39 6570 46
rect 6573 38 6640 66
rect 6672 66 6844 68
rect 6642 44 6670 48
rect 6672 44 6752 66
rect 6773 64 6788 66
rect 6642 42 6752 44
rect 6642 38 6670 42
rect 6672 38 6752 42
rect 6279 28 6309 38
rect 6336 28 6337 38
rect 6352 28 6365 38
rect 6379 28 6380 38
rect 6395 28 6408 38
rect 6423 28 6453 38
rect 6496 28 6539 38
rect 6546 28 6554 38
rect 6573 30 6576 38
rect 6640 30 6672 38
rect 6573 28 6739 30
rect 6758 28 6769 38
rect 6773 28 6803 38
rect 6831 28 6844 66
rect 6916 72 6951 80
rect 6916 46 6917 72
rect 6924 46 6951 72
rect 6916 38 6951 46
rect 6953 72 6994 80
rect 6953 46 6968 72
rect 6975 46 6994 72
rect 7058 68 7120 80
rect 7132 68 7207 80
rect 7265 68 7340 80
rect 7352 68 7383 80
rect 7389 68 7424 80
rect 7058 66 7220 68
rect 6953 38 6994 46
rect 7076 38 7089 66
rect 7104 64 7119 66
rect 7143 39 7150 46
rect 7153 38 7220 66
rect 7252 66 7424 68
rect 7222 44 7250 48
rect 7252 44 7332 66
rect 7353 64 7368 66
rect 7222 42 7332 44
rect 7222 38 7250 42
rect 7252 38 7332 42
rect 6859 28 6889 38
rect 6916 28 6917 38
rect 6932 28 6945 38
rect 6959 28 6960 38
rect 6975 28 6988 38
rect 7003 28 7033 38
rect 7076 28 7119 38
rect 7126 28 7134 38
rect 7153 30 7156 38
rect 7220 30 7252 38
rect 7153 28 7319 30
rect 7338 28 7349 38
rect 7353 28 7383 38
rect 7411 28 7424 66
rect 7496 72 7531 80
rect 7496 46 7497 72
rect 7504 46 7531 72
rect 7496 38 7531 46
rect 7533 72 7574 80
rect 7533 46 7548 72
rect 7555 46 7574 72
rect 7638 68 7700 80
rect 7712 68 7787 80
rect 7845 68 7920 80
rect 7932 68 7963 80
rect 7969 68 8004 80
rect 7638 66 7800 68
rect 7533 38 7574 46
rect 7656 38 7669 66
rect 7684 64 7699 66
rect 7723 39 7730 46
rect 7733 38 7800 66
rect 7832 66 8004 68
rect 7802 44 7830 48
rect 7832 44 7912 66
rect 7933 64 7948 66
rect 7802 42 7912 44
rect 7802 38 7830 42
rect 7832 38 7912 42
rect 7439 28 7469 38
rect 7496 28 7497 38
rect 7512 28 7525 38
rect 7539 28 7540 38
rect 7555 28 7568 38
rect 7583 28 7613 38
rect 7656 28 7699 38
rect 7706 28 7714 38
rect 7733 30 7736 38
rect 7800 30 7832 38
rect 7733 28 7899 30
rect 7918 28 7929 38
rect 7933 28 7963 38
rect 7991 28 8004 66
rect 8076 72 8111 80
rect 8076 46 8077 72
rect 8084 46 8111 72
rect 8076 38 8111 46
rect 8113 72 8154 80
rect 8113 46 8128 72
rect 8135 46 8154 72
rect 8218 68 8280 80
rect 8292 68 8367 80
rect 8425 68 8500 80
rect 8512 68 8543 80
rect 8549 68 8584 80
rect 8218 66 8380 68
rect 8113 38 8154 46
rect 8236 38 8249 66
rect 8264 64 8279 66
rect 8303 39 8310 46
rect 8313 38 8380 66
rect 8412 66 8584 68
rect 8382 44 8410 48
rect 8412 44 8492 66
rect 8513 64 8528 66
rect 8382 42 8492 44
rect 8382 38 8410 42
rect 8412 38 8492 42
rect 8019 28 8049 38
rect 8076 28 8077 38
rect 8092 28 8105 38
rect 8119 28 8120 38
rect 8135 28 8148 38
rect 8163 28 8193 38
rect 8236 28 8279 38
rect 8286 28 8294 38
rect 8313 30 8316 38
rect 8380 30 8412 38
rect 8313 28 8479 30
rect 8498 28 8509 38
rect 8513 28 8543 38
rect 8571 28 8584 66
rect 8656 72 8691 80
rect 8656 46 8657 72
rect 8664 46 8691 72
rect 8656 38 8691 46
rect 8693 72 8734 80
rect 8693 46 8708 72
rect 8715 46 8734 72
rect 8798 68 8860 80
rect 8872 68 8947 80
rect 9005 68 9080 80
rect 9092 68 9123 80
rect 9129 68 9164 80
rect 8798 66 8960 68
rect 8693 38 8734 46
rect 8816 38 8829 66
rect 8844 64 8859 66
rect 8883 39 8890 46
rect 8893 38 8960 66
rect 8992 66 9164 68
rect 8962 44 8990 48
rect 8992 44 9072 66
rect 9093 64 9108 66
rect 8962 42 9072 44
rect 8962 38 8990 42
rect 8992 38 9072 42
rect 8599 28 8629 38
rect 8656 28 8657 38
rect 8672 28 8685 38
rect 8699 28 8700 38
rect 8715 28 8728 38
rect 8743 28 8773 38
rect 8816 28 8859 38
rect 8866 28 8874 38
rect 8893 30 8896 38
rect 8960 30 8992 38
rect 8893 28 9059 30
rect 9078 28 9089 38
rect 9093 28 9123 38
rect 9151 28 9164 66
rect 9236 72 9271 80
rect 9236 46 9237 72
rect 9244 46 9271 72
rect 9236 38 9271 46
rect 9179 28 9209 38
rect 9236 28 9237 38
rect 9252 28 9265 38
rect -1 22 9265 28
rect 0 14 9265 22
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 129 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 243 0 294 1
rect 451 0 464 14
rect 244 -2 308 0
rect 479 -4 509 14
rect 552 0 565 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 709 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 823 0 874 1
rect 1031 0 1044 14
rect 824 -2 888 0
rect 1059 -4 1089 14
rect 1132 0 1145 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1289 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1403 0 1454 1
rect 1611 0 1624 14
rect 1404 -2 1468 0
rect 1639 -4 1669 14
rect 1712 0 1725 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1869 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1983 0 2034 1
rect 2191 0 2204 14
rect 1984 -2 2048 0
rect 2219 -4 2249 14
rect 2292 0 2305 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2449 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2563 0 2614 1
rect 2771 0 2784 14
rect 2564 -2 2628 0
rect 2799 -4 2829 14
rect 2872 0 2885 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3029 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3143 0 3194 1
rect 3351 0 3364 14
rect 3144 -2 3208 0
rect 3379 -4 3409 14
rect 3452 0 3465 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3609 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3723 0 3774 1
rect 3931 0 3944 14
rect 3724 -2 3788 0
rect 3959 -4 3989 14
rect 4032 0 4045 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4189 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4303 0 4354 1
rect 4511 0 4524 14
rect 4304 -2 4368 0
rect 4539 -4 4569 14
rect 4612 0 4625 14
rect 4655 0 4668 14
rect 4683 -4 4713 14
rect 4756 0 4769 14
rect 4806 1 4814 14
rect 4847 1 4985 14
rect 5018 1 5026 14
rect 4883 0 4934 1
rect 5091 0 5104 14
rect 4884 -2 4948 0
rect 5119 -4 5149 14
rect 5192 0 5205 14
rect 5235 0 5248 14
rect 5263 -4 5293 14
rect 5336 0 5349 14
rect 5386 1 5394 14
rect 5427 1 5565 14
rect 5598 1 5606 14
rect 5463 0 5514 1
rect 5671 0 5684 14
rect 5464 -2 5528 0
rect 5699 -4 5729 14
rect 5772 0 5785 14
rect 5815 0 5828 14
rect 5843 -4 5873 14
rect 5916 0 5929 14
rect 5966 1 5974 14
rect 6007 1 6145 14
rect 6178 1 6186 14
rect 6043 0 6094 1
rect 6251 0 6264 14
rect 6044 -2 6108 0
rect 6279 -4 6309 14
rect 6352 0 6365 14
rect 6395 0 6408 14
rect 6423 -4 6453 14
rect 6496 0 6509 14
rect 6546 1 6554 14
rect 6587 1 6725 14
rect 6758 1 6766 14
rect 6623 0 6674 1
rect 6831 0 6844 14
rect 6624 -2 6688 0
rect 6859 -4 6889 14
rect 6932 0 6945 14
rect 6975 0 6988 14
rect 7003 -4 7033 14
rect 7076 0 7089 14
rect 7126 1 7134 14
rect 7167 1 7305 14
rect 7338 1 7346 14
rect 7203 0 7254 1
rect 7411 0 7424 14
rect 7204 -2 7268 0
rect 7439 -4 7469 14
rect 7512 0 7525 14
rect 7555 0 7568 14
rect 7583 -4 7613 14
rect 7656 0 7669 14
rect 7706 1 7714 14
rect 7747 1 7885 14
rect 7918 1 7926 14
rect 7783 0 7834 1
rect 7991 0 8004 14
rect 7784 -2 7848 0
rect 8019 -4 8049 14
rect 8092 0 8105 14
rect 8135 0 8148 14
rect 8163 -4 8193 14
rect 8236 0 8249 14
rect 8286 1 8294 14
rect 8327 1 8465 14
rect 8498 1 8506 14
rect 8363 0 8414 1
rect 8571 0 8584 14
rect 8364 -2 8428 0
rect 8599 -4 8629 14
rect 8672 0 8685 14
rect 8715 0 8728 14
rect 8743 -4 8773 14
rect 8816 0 8829 14
rect 8866 1 8874 14
rect 8907 1 9045 14
rect 9078 1 9086 14
rect 8943 0 8994 1
rect 9151 0 9164 14
rect 8944 -2 9008 0
rect 9179 -4 9209 14
rect 9252 0 9265 14
<< pwell >>
rect 4612 7560 4640 7574
rect 4612 7516 4640 7530
rect 4612 7290 4640 7304
rect 4612 7246 4640 7260
rect 4612 7020 4640 7034
rect 4612 6976 4640 6990
rect 4612 6750 4640 6764
rect 4612 6706 4640 6720
rect 4612 6480 4640 6494
rect 4612 6436 4640 6450
rect 4612 6210 4640 6224
rect 4612 6166 4640 6180
rect 4612 5940 4640 5954
rect 4612 5896 4640 5910
rect 4612 5670 4640 5684
rect 4612 5626 4640 5640
rect 4612 5400 4640 5414
rect 4612 5356 4640 5370
rect 4612 5130 4640 5144
rect 4612 5086 4640 5100
rect 4612 4860 4640 4874
rect 4612 4816 4640 4830
rect 4612 4590 4640 4604
rect 4612 4546 4640 4560
rect 4612 4320 4640 4334
rect 4612 4276 4640 4290
rect 4612 4050 4640 4064
rect 4612 4006 4640 4020
rect 4612 3780 4640 3794
rect 4612 3736 4640 3750
rect 4612 3510 4640 3524
rect 4612 3466 4640 3480
rect 4612 3240 4640 3254
rect 4612 3196 4640 3210
rect 4612 2970 4640 2984
rect 4612 2926 4640 2940
rect 4612 2700 4640 2714
rect 4612 2656 4640 2670
rect 4612 2430 4640 2444
rect 4612 2386 4640 2400
rect 4612 2160 4640 2174
rect 4612 2116 4640 2130
rect 4612 1890 4640 1904
rect 4612 1846 4640 1860
rect 4612 1620 4640 1634
rect 4612 1576 4640 1590
rect 4612 1350 4640 1364
rect 4612 1306 4640 1320
rect 4612 1080 4640 1094
rect 4612 1036 4640 1050
rect 4612 810 4640 824
rect 4612 766 4640 780
rect 4612 540 4640 554
rect 4612 496 4640 510
rect 4612 270 4640 284
rect 4612 226 4640 240
rect 74 184 89 212
rect 464 184 479 213
rect 4714 184 4729 212
rect 5104 184 5119 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 4640 38 4655 80
rect 5177 38 5192 80
rect 5220 38 5235 80
rect 4612 0 4640 14
<< ndiffc >>
rect 74 184 89 212
rect 464 184 479 213
rect 654 184 669 212
rect 1044 184 1059 213
rect 1234 184 1249 212
rect 1624 184 1639 213
rect 1814 184 1829 212
rect 2204 184 2219 213
rect 2394 184 2409 212
rect 2784 184 2799 213
rect 2974 184 2989 212
rect 3364 184 3379 213
rect 3554 184 3569 212
rect 3944 184 3959 213
rect 4134 184 4149 212
rect 4524 184 4539 213
rect 4714 184 4729 212
rect 5104 184 5119 213
rect 5294 184 5309 212
rect 5684 184 5699 213
rect 5874 184 5889 212
rect 6264 184 6279 213
rect 6454 184 6469 212
rect 6844 184 6859 213
rect 7034 184 7049 212
rect 7424 184 7439 213
rect 7614 184 7629 212
rect 8004 184 8019 213
rect 8194 184 8209 212
rect 8584 184 8599 213
rect 8774 184 8789 212
rect 9164 184 9179 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 1117 38 1132 80
rect 1160 38 1175 80
rect 1697 38 1712 80
rect 1740 38 1755 80
rect 2277 38 2292 80
rect 2320 38 2335 80
rect 2857 38 2872 80
rect 2900 38 2915 80
rect 3437 38 3452 80
rect 3480 38 3495 80
rect 4017 38 4032 80
rect 4060 38 4075 80
rect 4597 38 4612 80
rect 4640 38 4655 80
rect 5177 38 5192 80
rect 5220 38 5235 80
rect 5757 38 5772 80
rect 5800 38 5815 80
rect 6337 38 6352 80
rect 6380 38 6395 80
rect 6917 38 6932 80
rect 6960 38 6975 80
rect 7497 38 7512 80
rect 7540 38 7555 80
rect 8077 38 8092 80
rect 8120 38 8135 80
rect 8657 38 8672 80
rect 8700 38 8715 80
rect 9237 38 9252 80
<< poly >>
rect 0 8610 30 8640
rect 4561 8610 4708 8640
rect 0 8340 30 8370
rect 4567 8340 4701 8370
rect 0 8070 30 8100
rect 4571 8070 4694 8100
rect 0 7800 30 7830
rect 4574 7800 4724 7830
rect 0 7530 30 7560
rect 4558 7530 4711 7560
rect 0 7260 30 7290
rect 4556 7260 4739 7290
rect 0 6990 30 7020
rect 4554 6990 4707 7020
rect 0 6720 30 6750
rect 4563 6720 4759 6750
rect 0 6450 30 6480
rect 4572 6450 4700 6480
rect 0 6180 30 6210
rect 4575 6180 4747 6210
rect 0 5910 30 5940
rect 4563 5910 4729 5940
rect 0 5640 30 5670
rect 4560 5640 4732 5670
rect 0 5370 30 5400
rect 4563 5370 4700 5400
rect 0 5100 30 5130
rect 4572 5100 4706 5130
rect 0 4830 30 4860
rect 4544 4830 4694 4860
rect 0 4560 30 4590
rect 4561 4560 4714 4590
rect 0 4290 30 4320
rect 4568 4290 4703 4320
rect 0 4020 30 4050
rect 4566 4020 4736 4050
rect 0 3750 30 3780
rect 4563 3750 4719 3780
rect 0 3480 30 3510
rect 4561 3480 4713 3510
rect 0 3210 30 3240
rect 4563 3210 4714 3240
rect 0 2940 30 2970
rect 4565 2940 4704 2970
rect 0 2670 30 2700
rect 4553 2670 4697 2700
rect 0 2400 30 2430
rect 4553 2400 4701 2430
rect 0 2130 30 2160
rect 4562 2130 4697 2160
rect 0 1860 30 1890
rect 4564 1860 4695 1890
rect 0 1590 30 1620
rect 4566 1590 4721 1620
rect 0 1320 30 1350
rect 4569 1320 4706 1350
rect 0 1050 30 1080
rect 4549 1050 4695 1080
rect 0 780 30 810
rect 4564 780 4713 810
rect 0 510 30 540
rect 4577 510 4701 540
rect 0 240 30 270
rect 4570 240 4698 270
<< metal1 >>
rect 0 8596 15 8610
rect 4576 8596 4671 8610
rect 0 8472 15 8506
rect 4505 8472 4691 8506
rect 0 8370 15 8384
rect 4573 8370 4670 8384
rect 0 8326 15 8340
rect 4578 8326 4678 8340
rect 0 8202 15 8236
rect 4502 8202 4701 8236
rect 0 8100 15 8114
rect 4578 8100 4688 8114
rect 0 8056 15 8070
rect 4581 8056 4663 8070
rect 0 7932 15 7966
rect 4505 7932 4727 7966
rect 0 7830 15 7844
rect 4582 7830 4666 7844
rect 0 7786 15 7800
rect 4575 7786 4685 7800
rect 0 7662 15 7696
rect 4640 7662 4655 7696
rect 0 7560 15 7574
rect 4612 7560 4655 7574
rect 0 7516 15 7530
rect 4612 7516 4655 7530
rect 0 7392 15 7426
rect 4504 7392 4727 7426
rect 0 7290 15 7304
rect 4612 7290 4655 7304
rect 0 7246 15 7260
rect 4612 7246 4655 7260
rect 0 7122 15 7156
rect 4496 7122 4683 7156
rect 0 7020 15 7034
rect 4612 7020 4655 7034
rect 0 6976 15 6990
rect 4612 6976 4655 6990
rect 0 6852 15 6886
rect 4505 6852 4734 6886
rect 0 6750 15 6764
rect 4612 6750 4655 6764
rect 0 6706 15 6720
rect 4612 6706 4655 6720
rect 0 6582 15 6616
rect 4502 6582 4705 6616
rect 0 6480 15 6494
rect 4612 6480 4655 6494
rect 0 6436 15 6450
rect 4612 6436 4655 6450
rect 0 6312 15 6346
rect 4505 6312 4722 6346
rect 0 6210 15 6224
rect 4612 6210 4655 6224
rect 0 6166 15 6180
rect 4612 6166 4655 6180
rect 0 6042 15 6076
rect 4499 6042 4731 6076
rect 0 5940 15 5954
rect 4612 5940 4655 5954
rect 0 5896 15 5910
rect 4612 5896 4655 5910
rect 0 5772 15 5806
rect 4505 5772 4740 5806
rect 0 5670 15 5684
rect 4612 5670 4655 5684
rect 0 5626 15 5640
rect 4612 5626 4655 5640
rect 0 5502 15 5536
rect 4505 5502 4728 5536
rect 0 5400 15 5414
rect 4612 5400 4655 5414
rect 0 5356 15 5370
rect 4612 5356 4655 5370
rect 0 5232 15 5266
rect 4496 5232 4728 5266
rect 0 5130 15 5144
rect 4612 5130 4655 5144
rect 0 5086 15 5100
rect 4612 5086 4655 5100
rect 0 4962 15 4996
rect 4502 4962 4746 4996
rect 0 4860 15 4874
rect 4612 4860 4655 4874
rect 0 4816 15 4830
rect 4612 4816 4655 4830
rect 0 4692 15 4726
rect 4505 4692 4716 4726
rect 0 4590 15 4604
rect 4612 4590 4655 4604
rect 0 4546 15 4560
rect 4612 4546 4655 4560
rect 0 4422 15 4456
rect 4503 4422 4753 4456
rect 0 4320 15 4334
rect 4612 4320 4655 4334
rect 0 4276 15 4290
rect 4612 4276 4655 4290
rect 0 4152 15 4186
rect 4505 4152 4724 4186
rect 0 4050 15 4064
rect 4612 4050 4655 4064
rect 0 4006 15 4020
rect 4612 4006 4655 4020
rect 0 3882 15 3916
rect 4503 3882 4731 3916
rect 0 3780 15 3794
rect 4612 3780 4655 3794
rect 0 3736 15 3750
rect 4612 3736 4655 3750
rect 0 3612 15 3646
rect 4505 3612 4736 3646
rect 0 3510 15 3524
rect 4612 3510 4655 3524
rect 0 3466 15 3480
rect 4612 3466 4655 3480
rect 0 3342 15 3376
rect 4496 3342 4727 3376
rect 0 3240 15 3254
rect 4612 3240 4655 3254
rect 0 3196 15 3210
rect 4612 3196 4655 3210
rect 0 3072 15 3106
rect 4502 3072 4741 3106
rect 0 2970 15 2984
rect 4612 2970 4655 2984
rect 0 2926 15 2940
rect 4612 2926 4655 2940
rect 0 2802 15 2836
rect 4502 2802 4734 2836
rect 0 2700 15 2714
rect 4612 2700 4655 2714
rect 0 2656 15 2670
rect 4612 2656 4655 2670
rect 0 2532 15 2566
rect 4505 2532 4736 2566
rect 0 2430 15 2444
rect 4612 2430 4655 2444
rect 0 2386 15 2400
rect 4612 2386 4655 2400
rect 0 2262 15 2296
rect 4497 2262 4740 2296
rect 0 2160 15 2174
rect 4612 2160 4655 2174
rect 0 2116 15 2130
rect 4612 2116 4655 2130
rect 0 1992 15 2026
rect 4505 1992 4710 2026
rect 0 1890 15 1904
rect 4612 1890 4655 1904
rect 0 1846 15 1860
rect 4612 1846 4655 1860
rect 0 1722 15 1756
rect 4505 1722 4688 1756
rect 0 1620 15 1634
rect 4612 1620 4655 1634
rect 0 1576 15 1590
rect 4612 1576 4655 1590
rect 0 1452 15 1486
rect 4501 1452 4708 1486
rect 0 1350 15 1364
rect 4612 1350 4655 1364
rect 0 1306 15 1320
rect 4612 1306 4655 1320
rect 0 1182 15 1216
rect 4505 1182 4701 1216
rect 0 1080 15 1094
rect 4612 1080 4655 1094
rect 0 1036 15 1050
rect 4612 1036 4655 1050
rect 0 912 15 946
rect 4505 912 4725 946
rect 0 810 15 824
rect 4612 810 4655 824
rect 0 766 15 780
rect 4612 766 4655 780
rect 0 642 15 676
rect 4505 642 4741 676
rect 0 540 15 554
rect 4612 540 4655 554
rect 0 496 15 510
rect 4612 496 4655 510
rect 0 372 15 406
rect 4505 372 4683 406
rect 0 270 15 284
rect 4612 270 4655 284
rect 0 226 15 240
rect 4612 226 4655 240
rect 0 102 15 136
rect 4505 102 4705 136
rect 0 0 15 14
rect 4612 0 4655 14
use 10T_1x8_magic  10T_1x8_magic_16
timestamp 1656019537
transform 1 0 0 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_18
timestamp 1656019537
transform 1 0 0 0 1 270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_17
timestamp 1656019537
transform 1 0 0 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_20
timestamp 1656019537
transform 1 0 0 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_19
timestamp 1656019537
transform 1 0 0 0 1 1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_37
timestamp 1656019537
transform 1 0 4640 0 1 1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_35
timestamp 1656019537
transform 1 0 4640 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_34
timestamp 1656019537
transform 1 0 4640 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_33
timestamp 1656019537
transform 1 0 4640 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_32
timestamp 1656019537
transform 1 0 4640 0 1 270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_22
timestamp 1656019537
transform 1 0 0 0 1 1350
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_21
timestamp 1656019537
transform 1 0 0 0 1 1620
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_24
timestamp 1656019537
transform 1 0 0 0 1 1890
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_23
timestamp 1656019537
transform 1 0 0 0 1 2160
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_39
timestamp 1656019537
transform 1 0 4640 0 1 2160
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_40
timestamp 1656019537
transform 1 0 4640 0 1 1620
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_38
timestamp 1656019537
transform 1 0 4640 0 1 1890
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_36
timestamp 1656019537
transform 1 0 4640 0 1 1350
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_26
timestamp 1656019537
transform 1 0 0 0 1 2430
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_25
timestamp 1656019537
transform 1 0 0 0 1 2700
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_28
timestamp 1656019537
transform 1 0 0 0 1 2970
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_27
timestamp 1656019537
transform 1 0 0 0 1 3240
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_42
timestamp 1656019537
transform 1 0 4640 0 1 2700
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_44
timestamp 1656019537
transform 1 0 4640 0 1 3240
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_43
timestamp 1656019537
transform 1 0 4640 0 1 2970
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_41
timestamp 1656019537
transform 1 0 4640 0 1 2430
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_29
timestamp 1656019537
transform 1 0 0 0 1 3780
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_30
timestamp 1656019537
transform 1 0 0 0 1 3510
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_31
timestamp 1656019537
transform 1 0 0 0 1 4050
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_9
timestamp 1656019537
transform 1 0 0 0 1 4320
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_48
timestamp 1656019537
transform 1 0 4640 0 1 4320
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_47
timestamp 1656019537
transform 1 0 4640 0 1 4050
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_46
timestamp 1656019537
transform 1 0 4640 0 1 3510
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_45
timestamp 1656019537
transform 1 0 4640 0 1 3780
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_8
timestamp 1656019537
transform 1 0 0 0 1 4590
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_10
timestamp 1656019537
transform 1 0 0 0 1 4860
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_11
timestamp 1656019537
transform 1 0 0 0 1 5130
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_12
timestamp 1656019537
transform 1 0 0 0 1 5400
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_52
timestamp 1656019537
transform 1 0 4640 0 1 5400
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_51
timestamp 1656019537
transform 1 0 4640 0 1 5130
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_50
timestamp 1656019537
transform 1 0 4640 0 1 4860
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_49
timestamp 1656019537
transform 1 0 4640 0 1 4590
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_13
timestamp 1656019537
transform 1 0 0 0 1 5670
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_15
timestamp 1656019537
transform 1 0 0 0 1 5940
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_14
timestamp 1656019537
transform 1 0 0 0 1 6210
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1656019537
transform 1 0 0 0 1 6480
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_56
timestamp 1656019537
transform 1 0 4640 0 1 6480
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_55
timestamp 1656019537
transform 1 0 4640 0 1 6210
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_54
timestamp 1656019537
transform 1 0 4640 0 1 5940
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_53
timestamp 1656019537
transform 1 0 4640 0 1 5670
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1656019537
transform 1 0 0 0 1 6750
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1656019537
transform 1 0 0 0 1 7020
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1656019537
transform 1 0 0 0 1 7290
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1656019537
transform 1 0 0 0 1 7560
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_60
timestamp 1656019537
transform 1 0 4640 0 1 7560
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_59
timestamp 1656019537
transform 1 0 4640 0 1 7290
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_58
timestamp 1656019537
transform 1 0 4640 0 1 7020
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_57
timestamp 1656019537
transform 1 0 4640 0 1 6750
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1656019537
transform 1 0 0 0 1 7830
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1656019537
transform 1 0 0 0 1 8100
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1656019537
transform 1 0 0 0 1 8370
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_63
timestamp 1656019537
transform 1 0 4640 0 1 8370
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_62
timestamp 1656019537
transform 1 0 4640 0 1 8100
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_61
timestamp 1656019537
transform 1 0 4640 0 1 7830
box -7 -4 4631 312
<< labels >>
rlabel locali 4640 38 4655 80 1 RBL1_0
port 1 ns signal output
rlabel locali 5177 38 5192 80 1 RBL0_0
port 2 ns signal output
rlabel locali 5220 38 5235 80 1 RBL1_1
port 3 ns signal output
rlabel locali 5757 38 5772 80 1 RBL0_1
port 4 ns signal output
rlabel locali 5800 38 5815 80 1 RBL1_2
port 5 ns signal output
rlabel locali 6337 38 6352 80 1 RBL0_2
port 6 ns signal output
rlabel locali 6380 38 6395 80 1 RBL1_3
port 7 ns signal output
rlabel locali 6917 38 6932 80 1 RBL0_3
port 8 ns signal output
rlabel locali 6960 38 6975 80 1 RBL1_4
port 9 ns signal output
rlabel locali 7497 38 7512 80 1 RBL0_4
port 10 ns signal output
rlabel locali 7540 38 7555 80 1 RBL1_5
port 11 ns signal output
rlabel locali 8077 38 8092 80 1 RBL0_5
port 12 ns signal output
rlabel locali 8120 38 8135 80 1 RBL1_6
port 13 ns signal output
rlabel locali 8657 38 8672 80 1 RBL0_6
port 14 ns signal output
rlabel locali 8700 38 8715 80 1 RBL1_7
port 15 ns signal output
rlabel locali 9237 38 9252 80 1 RBL0_7
port 16 ns signal output
rlabel locali 5104 184 5119 213 1 WBL_0
port 17 ns signal input
rlabel locali 4714 184 4729 212 1 WBLb_0
port 18 ns signal input
rlabel locali 5684 184 5699 213 1 WBL_1
port 19 ns signal input
rlabel locali 5294 184 5309 212 1 WBLb_1
port 20 ns signal input
rlabel locali 6264 184 6279 213 1 WBL_2
port 21 ns signal input
rlabel locali 5874 184 5889 212 1 WBLb_2
port 22 ns signal input
rlabel locali 6844 184 6859 213 1 WBL_3
port 23 ns signal input
rlabel locali 6454 184 6469 212 1 WBLb_3
port 24 ns signal input
rlabel locali 7424 184 7439 213 1 WBL_4
port 25 ns signal input
rlabel locali 7034 184 7049 212 1 WBLb_4
port 26 ns signal input
rlabel locali 8004 184 8019 213 1 WBL_5
port 27 ns signal input
rlabel locali 7614 184 7629 212 1 WBLb_5
port 28 ns signal input
rlabel locali 8584 184 8599 213 1 WBL_6
port 29 ns signal input
rlabel locali 8194 184 8209 212 1 WBLb_6
port 30 ns signal input
rlabel locali 9164 184 9179 213 1 WBL_7
port 31 ns signal input
rlabel locali 8774 184 8789 212 1 WBLb_7
port 32 ns signal input
rlabel metal1 0 4422 15 4456 1 RWL_15
port 64 ew signal input
rlabel poly 0 4560 30 4590 1 WWL_15
port 63 ew signal input
rlabel metal1 0 4692 15 4726 1 RWL_14
port 62 ew signal input
rlabel poly 0 4830 30 4860 1 WWL_14
port 61 ew signal input
rlabel metal1 0 4962 15 4996 1 RWL_13
port 60 ew signal input
rlabel poly 0 5100 30 5130 1 WWL_13
port 59 ew signal input
rlabel metal1 0 5232 15 5266 1 RWL_12
port 58 ew signal input
rlabel poly 0 5370 30 5400 1 WWL_12
port 57 ew signal input
rlabel metal1 0 5502 15 5536 1 RWL_11
port 56 ew signal input
rlabel poly 0 5640 30 5670 1 WWL_11
port 55 ew signal input
rlabel metal1 0 5772 15 5806 1 RWL_10
port 54 ew signal input
rlabel poly 0 5910 30 5940 1 WWL_10
port 53 ew signal input
rlabel metal1 0 6042 15 6076 1 RWL_9
port 52 ew signal input
rlabel poly 0 6180 30 6210 1 WWL_9
port 51 ew signal input
rlabel metal1 0 6312 15 6346 1 RWL_8
port 50 ew signal input
rlabel poly 0 6450 30 6480 1 WWL_8
port 49 ew signal input
rlabel metal1 0 6436 15 6450 1 VDD
rlabel metal1 0 6210 15 6224 1 GND
rlabel metal1 0 5896 15 5910 1 VDD
rlabel metal1 0 5626 15 5640 1 VDD
rlabel metal1 0 6166 15 6180 1 VDD
rlabel metal1 0 5356 15 5370 1 VDD
rlabel metal1 0 4816 15 4830 1 VDD
rlabel metal1 0 4546 15 4560 1 VDD
rlabel metal1 0 5086 15 5100 1 VDD
rlabel metal1 0 5400 15 5414 1 GND
rlabel metal1 0 5670 15 5684 1 GND
rlabel metal1 0 5940 15 5954 1 GND
rlabel metal1 0 5130 15 5144 1 GND
rlabel metal1 0 4320 15 4334 1 GND
rlabel metal1 0 4590 15 4604 1 GND
rlabel metal1 0 4860 15 4874 1 GND
rlabel poly 0 8610 30 8640 1 WWL_0
port 33 ew signal input
rlabel metal1 0 7020 15 7034 1 GND
rlabel metal1 0 6750 15 6764 1 GND
rlabel metal1 0 6480 15 6494 1 GND
rlabel metal1 0 7290 15 7304 1 GND
rlabel metal1 0 8100 15 8114 1 GND
rlabel metal1 0 7830 15 7844 1 GND
rlabel metal1 0 7560 15 7574 1 GND
rlabel metal1 0 7246 15 7260 1 VDD
rlabel metal1 0 6706 15 6720 1 VDD
rlabel metal1 0 6976 15 6990 1 VDD
rlabel metal1 0 7516 15 7530 1 VDD
rlabel metal1 0 8326 15 8340 1 VDD
rlabel metal1 0 7786 15 7800 1 VDD
rlabel metal1 0 8056 15 8070 1 VDD
rlabel metal1 0 8370 15 8384 1 GND
port 98 ew ground bidirectional abutment
rlabel metal1 0 8596 15 8610 1 VDD
port 97 ew power bidirectional abutment
rlabel metal1 0 6582 15 6616 1 RWL_7
port 48 ew signal input
rlabel poly 0 6720 30 6750 1 WWL_7
port 47 ew signal input
rlabel metal1 0 6852 15 6886 1 RWL_6
port 46 ew signal input
rlabel poly 0 6990 30 7020 1 WWL_6
port 45 ew signal input
rlabel metal1 0 7122 15 7156 1 RWL_5
port 44 ew signal input
rlabel poly 0 7260 30 7290 1 WWL_5
port 43 ew signal input
rlabel metal1 0 7392 15 7426 1 RWL_4
port 42 ew signal input
rlabel poly 0 7530 30 7560 1 WWL_4
port 41 ew signal input
rlabel metal1 0 7662 15 7696 1 RWL_3
port 40 ew signal input
rlabel poly 0 7800 30 7830 1 WWL_3
port 39 ew signal input
rlabel metal1 0 7932 15 7966 1 RWL_2
port 38 ew signal input
rlabel poly 0 8070 30 8100 1 WWL_2
port 37 ew signal input
rlabel metal1 0 8202 15 8236 1 RWL_1
port 36 ew signal input
rlabel poly 0 8340 30 8370 1 WWL_1
port 35 ew signal input
rlabel metal1 0 8472 15 8506 1 RWL_0
port 34 ew signal input
rlabel locali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel locali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel locali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel locali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel locali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel locali 2320 38 2335 80 1 RBL1_4
port 9 ns signal output
rlabel locali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel locali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel locali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel locali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel locali 464 184 479 213 1 WBL_0
port 17 ns signal input
rlabel locali 74 184 89 212 1 WBLb_0
port 18 ns signal input
rlabel locali 1044 184 1059 213 1 WBL_1
port 19 ns signal input
rlabel locali 654 184 669 212 1 WBLb_1
port 20 ns signal input
rlabel locali 1624 184 1639 213 1 WBL_2
port 21 ns signal input
rlabel locali 1234 184 1249 212 1 WBLb_2
port 22 ns signal input
rlabel locali 2204 184 2219 213 1 WBL_3
port 23 ns signal input
rlabel locali 1814 184 1829 212 1 WBLb_3
port 24 ns signal input
rlabel locali 2784 184 2799 213 1 WBL_4
port 25 ns signal input
rlabel locali 2394 184 2409 212 1 WBLb_4
port 26 ns signal input
rlabel locali 3364 184 3379 213 1 WBL_5
port 27 ns signal input
rlabel locali 2974 184 2989 212 1 WBLb_5
port 28 ns signal input
rlabel locali 3944 184 3959 213 1 WBL_6
port 29 ns signal input
rlabel locali 3554 184 3569 212 1 WBLb_6
port 30 ns signal input
rlabel locali 4524 184 4539 213 1 WBL_7
port 31 ns signal input
rlabel locali 4134 184 4149 212 1 WBLb_7
port 32 ns signal input
rlabel metal1 0 2116 15 2130 1 VDD
rlabel metal1 0 1890 15 1904 1 GND
rlabel metal1 0 1576 15 1590 1 VDD
rlabel metal1 0 1306 15 1320 1 VDD
rlabel metal1 0 1846 15 1860 1 VDD
rlabel metal1 0 1036 15 1050 1 VDD
rlabel metal1 0 496 15 510 1 VDD
rlabel metal1 0 226 15 240 1 VDD
rlabel metal1 0 766 15 780 1 VDD
rlabel metal1 0 1080 15 1094 1 GND
rlabel metal1 0 1350 15 1364 1 GND
rlabel metal1 0 1620 15 1634 1 GND
rlabel metal1 0 810 15 824 1 GND
rlabel metal1 0 0 15 14 1 GND
rlabel metal1 0 270 15 284 1 GND
rlabel metal1 0 540 15 554 1 GND
rlabel metal1 0 2700 15 2714 1 GND
rlabel metal1 0 2430 15 2444 1 GND
rlabel metal1 0 2160 15 2174 1 GND
rlabel metal1 0 2970 15 2984 1 GND
rlabel metal1 0 3780 15 3794 1 GND
rlabel metal1 0 3510 15 3524 1 GND
rlabel metal1 0 3240 15 3254 1 GND
rlabel metal1 0 2926 15 2940 1 VDD
rlabel metal1 0 2386 15 2400 1 VDD
rlabel metal1 0 2656 15 2670 1 VDD
rlabel metal1 0 3196 15 3210 1 VDD
rlabel metal1 0 4006 15 4020 1 VDD
rlabel metal1 0 3466 15 3480 1 VDD
rlabel metal1 0 3736 15 3750 1 VDD
rlabel metal1 0 4050 15 4064 1 GND
port 98 ew ground bidirectional abutment
rlabel metal1 0 4276 15 4290 1 VDD
port 97 ew power bidirectional abutment
rlabel poly 0 4290 30 4320 1 WWL_16
port 65 ew signal input
rlabel metal1 0 4152 15 4186 1 RWL_16
port 66 ew signal input
rlabel poly 0 4020 30 4050 1 WWL_17
port 67 ew signal input
rlabel metal1 0 3882 15 3916 1 RWL_17
port 68 ew signal input
rlabel poly 0 3750 30 3780 1 WWL_18
port 69 ew signal input
rlabel metal1 0 3612 15 3646 1 RWL_18
port 70 ew signal input
rlabel poly 0 3480 30 3510 1 WWL_19
port 71 ew signal input
rlabel metal1 0 3342 15 3376 1 RWL_19
port 72 ew signal input
rlabel poly 0 3210 30 3240 1 WWL_20
port 73 ew signal input
rlabel metal1 0 3072 15 3106 1 RWL_20
port 74 ew signal input
rlabel poly 0 2940 30 2970 1 WWL_21
port 75 ew signal input
rlabel metal1 0 2802 15 2836 1 RWL_21
port 76 ew signal input
rlabel poly 0 2670 30 2700 1 WWL_22
port 77 ew signal input
rlabel metal1 0 2532 15 2566 1 RWL_22
port 78 ew signal input
rlabel poly 0 2400 30 2430 1 WWL_23
port 79 ew signal input
rlabel metal1 0 2262 15 2296 1 RWL_23
port 80 ew signal input
rlabel poly 0 2130 30 2160 1 WWL_24
port 81 ew signal input
rlabel metal1 0 1992 15 2026 1 RWL_24
port 82 ew signal input
rlabel poly 0 1860 30 1890 1 WWL_25
port 83 ew signal input
rlabel metal1 0 1722 15 1756 1 RWL_25
port 84 ew signal input
rlabel poly 0 1590 30 1620 1 WWL_26
port 85 ew signal input
rlabel metal1 0 1452 15 1486 1 RWL_26
port 86 ew signal input
rlabel poly 0 1320 30 1350 1 WWL_27
port 87 ew signal input
rlabel metal1 0 1182 15 1216 1 RWL_27
port 88 ew signal input
rlabel poly 0 1050 30 1080 1 WWL_28
port 89 ew signal input
rlabel metal1 0 912 15 946 1 RWL_28
port 90 ew signal input
rlabel poly 0 780 30 810 1 WWL_29
port 91 ew signal input
rlabel metal1 0 642 15 676 1 RWL_29
port 92 ew signal input
rlabel poly 0 510 30 540 1 WWL_30
port 93 ew signal input
rlabel metal1 0 372 15 406 1 RWL_30
port 94 ew signal input
rlabel poly 0 240 30 270 1 WWL_31
port 95 ew signal input
rlabel metal1 0 102 15 136 1 RWL_31
port 96 ew signal input
rlabel metal1 4640 4422 4655 4456 1 RWL_15
port 64 ew signal input
rlabel poly 4640 4560 4670 4590 1 WWL_15
port 63 ew signal input
rlabel metal1 4640 4692 4655 4726 1 RWL_14
port 62 ew signal input
rlabel poly 4640 4830 4670 4860 1 WWL_14
port 61 ew signal input
rlabel metal1 4640 4962 4655 4996 1 RWL_13
port 60 ew signal input
rlabel poly 4640 5100 4670 5130 1 WWL_13
port 59 ew signal input
rlabel metal1 4640 5232 4655 5266 1 RWL_12
port 58 ew signal input
rlabel poly 4640 5370 4670 5400 1 WWL_12
port 57 ew signal input
rlabel metal1 4640 5502 4655 5536 1 RWL_11
port 56 ew signal input
rlabel poly 4640 5640 4670 5670 1 WWL_11
port 55 ew signal input
rlabel metal1 4640 5772 4655 5806 1 RWL_10
port 54 ew signal input
rlabel poly 4640 5910 4670 5940 1 WWL_10
port 53 ew signal input
rlabel metal1 4640 6042 4655 6076 1 RWL_9
port 52 ew signal input
rlabel poly 4640 6180 4670 6210 1 WWL_9
port 51 ew signal input
rlabel metal1 4640 6312 4655 6346 1 RWL_8
port 50 ew signal input
rlabel poly 4640 6450 4670 6480 1 WWL_8
port 49 ew signal input
rlabel metal1 4640 6436 4655 6450 1 VDD
rlabel metal1 4640 6210 4655 6224 1 GND
rlabel metal1 4640 5896 4655 5910 1 VDD
rlabel metal1 4640 5626 4655 5640 1 VDD
rlabel metal1 4640 6166 4655 6180 1 VDD
rlabel metal1 4640 5356 4655 5370 1 VDD
rlabel metal1 4640 4816 4655 4830 1 VDD
rlabel metal1 4640 4546 4655 4560 1 VDD
rlabel metal1 4640 5086 4655 5100 1 VDD
rlabel metal1 4640 5400 4655 5414 1 GND
rlabel metal1 4640 5670 4655 5684 1 GND
rlabel metal1 4640 5940 4655 5954 1 GND
rlabel metal1 4640 5130 4655 5144 1 GND
rlabel metal1 4640 4320 4655 4334 1 GND
rlabel metal1 4640 4590 4655 4604 1 GND
rlabel metal1 4640 4860 4655 4874 1 GND
rlabel poly 4640 8610 4670 8640 1 WWL_0
port 33 ew signal input
rlabel metal1 4640 7020 4655 7034 1 GND
rlabel metal1 4640 6750 4655 6764 1 GND
rlabel metal1 4640 6480 4655 6494 1 GND
rlabel metal1 4640 7290 4655 7304 1 GND
rlabel metal1 4640 8100 4655 8114 1 GND
rlabel metal1 4640 7830 4655 7844 1 GND
rlabel metal1 4640 7560 4655 7574 1 GND
rlabel metal1 4640 7246 4655 7260 1 VDD
rlabel metal1 4640 6706 4655 6720 1 VDD
rlabel metal1 4640 6976 4655 6990 1 VDD
rlabel metal1 4640 7516 4655 7530 1 VDD
rlabel metal1 4640 8326 4655 8340 1 VDD
rlabel metal1 4640 7786 4655 7800 1 VDD
rlabel metal1 4640 8056 4655 8070 1 VDD
rlabel metal1 4640 8370 4655 8384 1 GND
port 98 ew ground bidirectional abutment
rlabel metal1 4640 8596 4655 8610 1 VDD
port 97 ew power bidirectional abutment
rlabel metal1 4640 6582 4655 6616 1 RWL_7
port 48 ew signal input
rlabel poly 4640 6720 4670 6750 1 WWL_7
port 47 ew signal input
rlabel metal1 4640 6852 4655 6886 1 RWL_6
port 46 ew signal input
rlabel poly 4640 6990 4670 7020 1 WWL_6
port 45 ew signal input
rlabel metal1 4640 7122 4655 7156 1 RWL_5
port 44 ew signal input
rlabel poly 4640 7260 4670 7290 1 WWL_5
port 43 ew signal input
rlabel metal1 4640 7392 4655 7426 1 RWL_4
port 42 ew signal input
rlabel poly 4640 7530 4670 7560 1 WWL_4
port 41 ew signal input
rlabel metal1 4640 7662 4655 7696 1 RWL_3
port 40 ew signal input
rlabel poly 4640 7800 4670 7830 1 WWL_3
port 39 ew signal input
rlabel metal1 4640 7932 4655 7966 1 RWL_2
port 38 ew signal input
rlabel poly 4640 8070 4670 8100 1 WWL_2
port 37 ew signal input
rlabel metal1 4640 8202 4655 8236 1 RWL_1
port 36 ew signal input
rlabel poly 4640 8340 4670 8370 1 WWL_1
port 35 ew signal input
rlabel metal1 4640 8472 4655 8506 1 RWL_0
port 34 ew signal input
rlabel poly 4640 4290 4670 4320 1 WWL_16
port 65 ew signal input
rlabel metal1 4640 4152 4655 4186 1 RWL_16
port 66 ew signal input
rlabel poly 4640 4020 4670 4050 1 WWL_17
port 67 ew signal input
rlabel metal1 4640 3882 4655 3916 1 RWL_17
port 68 ew signal input
rlabel poly 4640 3750 4670 3780 1 WWL_18
port 69 ew signal input
rlabel metal1 4640 3612 4655 3646 1 RWL_18
port 70 ew signal input
rlabel poly 4640 3480 4670 3510 1 WWL_19
port 71 ew signal input
rlabel metal1 4640 3342 4655 3376 1 RWL_19
port 72 ew signal input
rlabel poly 4640 3210 4670 3240 1 WWL_20
port 73 ew signal input
rlabel metal1 4640 3072 4655 3106 1 RWL_20
port 74 ew signal input
rlabel poly 4640 2940 4670 2970 1 WWL_21
port 75 ew signal input
rlabel metal1 4640 2802 4655 2836 1 RWL_21
port 76 ew signal input
rlabel poly 4640 2670 4670 2700 1 WWL_22
port 77 ew signal input
rlabel metal1 4640 2532 4655 2566 1 RWL_22
port 78 ew signal input
rlabel poly 4640 2400 4670 2430 1 WWL_23
port 79 ew signal input
rlabel metal1 4640 2262 4655 2296 1 RWL_23
port 80 ew signal input
rlabel poly 4640 2130 4670 2160 1 WWL_24
port 81 ew signal input
rlabel metal1 4640 1992 4655 2026 1 RWL_24
port 82 ew signal input
rlabel poly 4640 1860 4670 1890 1 WWL_25
port 83 ew signal input
rlabel metal1 4640 1722 4655 1756 1 RWL_25
port 84 ew signal input
rlabel poly 4640 1590 4670 1620 1 WWL_26
port 85 ew signal input
rlabel metal1 4640 1452 4655 1486 1 RWL_26
port 86 ew signal input
rlabel poly 4640 1320 4670 1350 1 WWL_27
port 87 ew signal input
rlabel metal1 4640 1182 4655 1216 1 RWL_27
port 88 ew signal input
rlabel poly 4640 1050 4670 1080 1 WWL_28
port 89 ew signal input
rlabel metal1 4640 912 4655 946 1 RWL_28
port 90 ew signal input
rlabel poly 4640 780 4670 810 1 WWL_29
port 91 ew signal input
rlabel metal1 4640 642 4655 676 1 RWL_29
port 92 ew signal input
rlabel poly 4640 510 4670 540 1 WWL_30
port 93 ew signal input
rlabel metal1 4640 372 4655 406 1 RWL_30
port 94 ew signal input
rlabel poly 4640 240 4670 270 1 WWL_31
port 95 ew signal input
rlabel metal1 4640 102 4655 136 1 RWL_31
port 96 ew signal input
rlabel metal1 4640 4276 4655 4290 1 VDD
port 97 ew power bidirectional abutment
rlabel metal1 4640 4050 4655 4064 1 GND
port 98 ew ground bidirectional abutment
rlabel metal1 4640 2116 4655 2130 1 VDD
rlabel metal1 4640 1890 4655 1904 1 GND
rlabel metal1 4640 1576 4655 1590 1 VDD
rlabel metal1 4640 1306 4655 1320 1 VDD
rlabel metal1 4640 1846 4655 1860 1 VDD
rlabel metal1 4640 1036 4655 1050 1 VDD
rlabel metal1 4640 496 4655 510 1 VDD
rlabel metal1 4640 226 4655 240 1 VDD
rlabel metal1 4640 766 4655 780 1 VDD
rlabel metal1 4640 1080 4655 1094 1 GND
rlabel metal1 4640 1350 4655 1364 1 GND
rlabel metal1 4640 1620 4655 1634 1 GND
rlabel metal1 4640 810 4655 824 1 GND
rlabel metal1 4640 0 4655 14 1 GND
rlabel metal1 4640 270 4655 284 1 GND
rlabel metal1 4640 540 4655 554 1 GND
rlabel metal1 4640 2700 4655 2714 1 GND
rlabel metal1 4640 2430 4655 2444 1 GND
rlabel metal1 4640 2160 4655 2174 1 GND
rlabel metal1 4640 2970 4655 2984 1 GND
rlabel metal1 4640 3780 4655 3794 1 GND
rlabel metal1 4640 3510 4655 3524 1 GND
rlabel metal1 4640 3240 4655 3254 1 GND
rlabel metal1 4640 2926 4655 2940 1 VDD
rlabel metal1 4640 2386 4655 2400 1 VDD
rlabel metal1 4640 2656 4655 2670 1 VDD
rlabel metal1 4640 3196 4655 3210 1 VDD
rlabel metal1 4640 4006 4655 4020 1 VDD
rlabel metal1 4640 3466 4655 3480 1 VDD
rlabel metal1 4640 3736 4655 3750 1 VDD
<< end >>
