magic
tech sky130A
magscale 1 2
timestamp 1656029294
<< error_s >>
rect 15 8624 28 8640
rect 117 8638 130 8640
rect 83 8624 98 8638
rect 107 8624 137 8638
rect 198 8636 351 8682
rect 180 8624 372 8636
rect 415 8624 445 8638
rect 451 8624 464 8640
rect 552 8624 565 8640
rect 595 8624 608 8640
rect 697 8638 710 8640
rect 663 8624 678 8638
rect 687 8624 717 8638
rect 778 8636 931 8682
rect 760 8624 952 8636
rect 995 8624 1025 8638
rect 1031 8624 1044 8640
rect 1132 8624 1145 8640
rect 1175 8624 1188 8640
rect 1277 8638 1290 8640
rect 1243 8624 1258 8638
rect 1267 8624 1297 8638
rect 1358 8636 1511 8682
rect 1340 8624 1532 8636
rect 1575 8624 1605 8638
rect 1611 8624 1624 8640
rect 1712 8624 1725 8640
rect 1755 8624 1768 8640
rect 1857 8638 1870 8640
rect 1823 8624 1838 8638
rect 1847 8624 1877 8638
rect 1938 8636 2091 8682
rect 1920 8624 2112 8636
rect 2155 8624 2185 8638
rect 2191 8624 2204 8640
rect 2292 8624 2305 8640
rect 2335 8624 2348 8640
rect 2437 8638 2450 8640
rect 2403 8624 2418 8638
rect 2427 8624 2457 8638
rect 2518 8636 2671 8682
rect 2500 8624 2692 8636
rect 2735 8624 2765 8638
rect 2771 8624 2784 8640
rect 2872 8624 2885 8640
rect 2915 8624 2928 8640
rect 3017 8638 3030 8640
rect 2983 8624 2998 8638
rect 3007 8624 3037 8638
rect 3098 8636 3251 8682
rect 3080 8624 3272 8636
rect 3315 8624 3345 8638
rect 3351 8624 3364 8640
rect 3452 8624 3465 8640
rect 3495 8624 3508 8640
rect 3597 8638 3610 8640
rect 3563 8624 3578 8638
rect 3587 8624 3617 8638
rect 3678 8636 3831 8682
rect 3660 8624 3852 8636
rect 3895 8624 3925 8638
rect 3931 8624 3944 8640
rect 4032 8624 4045 8640
rect 4075 8624 4088 8640
rect 4177 8638 4190 8640
rect 4143 8624 4158 8638
rect 4167 8624 4197 8638
rect 4258 8636 4411 8682
rect 4240 8624 4432 8636
rect 4475 8624 4505 8638
rect 4511 8624 4524 8640
rect 4612 8624 4625 8640
rect 0 8610 4625 8624
rect 15 8506 28 8610
rect 73 8588 74 8598
rect 89 8588 102 8598
rect 73 8584 102 8588
rect 107 8584 137 8610
rect 155 8596 171 8598
rect 243 8596 296 8610
rect 244 8594 308 8596
rect 351 8594 366 8610
rect 415 8607 445 8610
rect 415 8604 451 8607
rect 381 8596 397 8598
rect 155 8584 170 8588
rect 73 8582 170 8584
rect 198 8582 366 8594
rect 382 8584 397 8588
rect 415 8585 454 8604
rect 473 8598 480 8599
rect 479 8591 480 8598
rect 463 8588 464 8591
rect 479 8588 492 8591
rect 415 8584 445 8585
rect 454 8584 460 8585
rect 463 8584 492 8588
rect 382 8583 492 8584
rect 382 8582 498 8583
rect 57 8574 108 8582
rect 57 8562 82 8574
rect 89 8562 108 8574
rect 139 8574 189 8582
rect 139 8566 155 8574
rect 162 8572 189 8574
rect 198 8572 419 8582
rect 162 8562 419 8572
rect 448 8574 498 8582
rect 448 8565 464 8574
rect 57 8554 108 8562
rect 155 8554 419 8562
rect 445 8562 464 8565
rect 471 8562 498 8574
rect 445 8554 498 8562
rect 73 8546 74 8554
rect 89 8546 102 8554
rect 73 8538 89 8546
rect 70 8531 89 8534
rect 70 8522 92 8531
rect 43 8512 92 8522
rect 43 8506 73 8512
rect 92 8507 97 8512
rect 15 8490 89 8506
rect 107 8498 137 8554
rect 172 8544 380 8554
rect 415 8550 460 8554
rect 463 8553 464 8554
rect 479 8553 492 8554
rect 198 8514 387 8544
rect 213 8511 387 8514
rect 206 8508 387 8511
rect 15 8488 28 8490
rect 43 8488 77 8490
rect 15 8472 89 8488
rect 116 8484 129 8498
rect 144 8484 160 8500
rect 206 8495 217 8508
rect -1 8450 0 8466
rect 15 8450 28 8472
rect 43 8450 73 8472
rect 116 8468 178 8484
rect 206 8477 217 8493
rect 222 8488 232 8508
rect 242 8488 256 8508
rect 259 8495 268 8508
rect 284 8495 293 8508
rect 222 8477 256 8488
rect 259 8477 268 8493
rect 284 8477 293 8493
rect 300 8488 310 8508
rect 320 8488 334 8508
rect 335 8495 346 8508
rect 300 8477 334 8488
rect 335 8477 346 8493
rect 392 8484 408 8500
rect 415 8498 445 8550
rect 479 8546 480 8553
rect 464 8538 480 8546
rect 451 8506 464 8525
rect 479 8506 509 8522
rect 451 8490 525 8506
rect 451 8488 464 8490
rect 479 8488 513 8490
rect 116 8466 129 8468
rect 144 8466 178 8468
rect 116 8450 178 8466
rect 222 8461 238 8464
rect 300 8461 330 8472
rect 378 8468 424 8484
rect 451 8472 525 8488
rect 378 8466 412 8468
rect 377 8450 424 8466
rect 451 8450 464 8472
rect 479 8450 509 8472
rect 536 8450 537 8466
rect 552 8450 565 8610
rect 595 8506 608 8610
rect 653 8588 654 8598
rect 669 8588 682 8598
rect 653 8584 682 8588
rect 687 8584 717 8610
rect 735 8596 751 8598
rect 823 8596 876 8610
rect 824 8594 888 8596
rect 931 8594 946 8610
rect 995 8607 1025 8610
rect 995 8604 1031 8607
rect 961 8596 977 8598
rect 735 8584 750 8588
rect 653 8582 750 8584
rect 778 8582 946 8594
rect 962 8584 977 8588
rect 995 8585 1034 8604
rect 1053 8598 1060 8599
rect 1059 8591 1060 8598
rect 1043 8588 1044 8591
rect 1059 8588 1072 8591
rect 995 8584 1025 8585
rect 1034 8584 1040 8585
rect 1043 8584 1072 8588
rect 962 8583 1072 8584
rect 962 8582 1078 8583
rect 637 8574 688 8582
rect 637 8562 662 8574
rect 669 8562 688 8574
rect 719 8574 769 8582
rect 719 8566 735 8574
rect 742 8572 769 8574
rect 778 8572 999 8582
rect 742 8562 999 8572
rect 1028 8574 1078 8582
rect 1028 8565 1044 8574
rect 637 8554 688 8562
rect 735 8554 999 8562
rect 1025 8562 1044 8565
rect 1051 8562 1078 8574
rect 1025 8554 1078 8562
rect 653 8546 654 8554
rect 669 8546 682 8554
rect 653 8538 669 8546
rect 650 8531 669 8534
rect 650 8522 672 8531
rect 623 8512 672 8522
rect 623 8506 653 8512
rect 672 8507 677 8512
rect 595 8490 669 8506
rect 687 8498 717 8554
rect 752 8544 960 8554
rect 995 8550 1040 8554
rect 1043 8553 1044 8554
rect 1059 8553 1072 8554
rect 778 8514 967 8544
rect 793 8511 967 8514
rect 786 8508 967 8511
rect 595 8488 608 8490
rect 623 8488 657 8490
rect 595 8472 669 8488
rect 696 8484 709 8498
rect 724 8484 740 8500
rect 786 8495 797 8508
rect 579 8450 580 8466
rect 595 8450 608 8472
rect 623 8450 653 8472
rect 696 8468 758 8484
rect 786 8477 797 8493
rect 802 8488 812 8508
rect 822 8488 836 8508
rect 839 8495 848 8508
rect 864 8495 873 8508
rect 802 8477 836 8488
rect 839 8477 848 8493
rect 864 8477 873 8493
rect 880 8488 890 8508
rect 900 8488 914 8508
rect 915 8495 926 8508
rect 880 8477 914 8488
rect 915 8477 926 8493
rect 972 8484 988 8500
rect 995 8498 1025 8550
rect 1059 8546 1060 8553
rect 1044 8538 1060 8546
rect 1031 8506 1044 8525
rect 1059 8506 1089 8522
rect 1031 8490 1105 8506
rect 1031 8488 1044 8490
rect 1059 8488 1093 8490
rect 696 8466 709 8468
rect 724 8466 758 8468
rect 696 8450 758 8466
rect 802 8461 818 8464
rect 880 8461 910 8472
rect 958 8468 1004 8484
rect 1031 8472 1105 8488
rect 958 8466 992 8468
rect 957 8450 1004 8466
rect 1031 8450 1044 8472
rect 1059 8450 1089 8472
rect 1116 8450 1117 8466
rect 1132 8450 1145 8610
rect 1175 8506 1188 8610
rect 1233 8588 1234 8598
rect 1249 8588 1262 8598
rect 1233 8584 1262 8588
rect 1267 8584 1297 8610
rect 1315 8596 1331 8598
rect 1403 8596 1456 8610
rect 1404 8594 1468 8596
rect 1511 8594 1526 8610
rect 1575 8607 1605 8610
rect 1575 8604 1611 8607
rect 1541 8596 1557 8598
rect 1315 8584 1330 8588
rect 1233 8582 1330 8584
rect 1358 8582 1526 8594
rect 1542 8584 1557 8588
rect 1575 8585 1614 8604
rect 1633 8598 1640 8599
rect 1639 8591 1640 8598
rect 1623 8588 1624 8591
rect 1639 8588 1652 8591
rect 1575 8584 1605 8585
rect 1614 8584 1620 8585
rect 1623 8584 1652 8588
rect 1542 8583 1652 8584
rect 1542 8582 1658 8583
rect 1217 8574 1268 8582
rect 1217 8562 1242 8574
rect 1249 8562 1268 8574
rect 1299 8574 1349 8582
rect 1299 8566 1315 8574
rect 1322 8572 1349 8574
rect 1358 8572 1579 8582
rect 1322 8562 1579 8572
rect 1608 8574 1658 8582
rect 1608 8565 1624 8574
rect 1217 8554 1268 8562
rect 1315 8554 1579 8562
rect 1605 8562 1624 8565
rect 1631 8562 1658 8574
rect 1605 8554 1658 8562
rect 1233 8546 1234 8554
rect 1249 8546 1262 8554
rect 1233 8538 1249 8546
rect 1230 8531 1249 8534
rect 1230 8522 1252 8531
rect 1203 8512 1252 8522
rect 1203 8506 1233 8512
rect 1252 8507 1257 8512
rect 1175 8490 1249 8506
rect 1267 8498 1297 8554
rect 1332 8544 1540 8554
rect 1575 8550 1620 8554
rect 1623 8553 1624 8554
rect 1639 8553 1652 8554
rect 1358 8514 1547 8544
rect 1373 8511 1547 8514
rect 1366 8508 1547 8511
rect 1175 8488 1188 8490
rect 1203 8488 1237 8490
rect 1175 8472 1249 8488
rect 1276 8484 1289 8498
rect 1304 8484 1320 8500
rect 1366 8495 1377 8508
rect 1159 8450 1160 8466
rect 1175 8450 1188 8472
rect 1203 8450 1233 8472
rect 1276 8468 1338 8484
rect 1366 8477 1377 8493
rect 1382 8488 1392 8508
rect 1402 8488 1416 8508
rect 1419 8495 1428 8508
rect 1444 8495 1453 8508
rect 1382 8477 1416 8488
rect 1419 8477 1428 8493
rect 1444 8477 1453 8493
rect 1460 8488 1470 8508
rect 1480 8488 1494 8508
rect 1495 8495 1506 8508
rect 1460 8477 1494 8488
rect 1495 8477 1506 8493
rect 1552 8484 1568 8500
rect 1575 8498 1605 8550
rect 1639 8546 1640 8553
rect 1624 8538 1640 8546
rect 1611 8506 1624 8525
rect 1639 8506 1669 8522
rect 1611 8490 1685 8506
rect 1611 8488 1624 8490
rect 1639 8488 1673 8490
rect 1276 8466 1289 8468
rect 1304 8466 1338 8468
rect 1276 8450 1338 8466
rect 1382 8461 1398 8464
rect 1460 8461 1490 8472
rect 1538 8468 1584 8484
rect 1611 8472 1685 8488
rect 1538 8466 1572 8468
rect 1537 8450 1584 8466
rect 1611 8450 1624 8472
rect 1639 8450 1669 8472
rect 1696 8450 1697 8466
rect 1712 8450 1725 8610
rect 1755 8506 1768 8610
rect 1813 8588 1814 8598
rect 1829 8588 1842 8598
rect 1813 8584 1842 8588
rect 1847 8584 1877 8610
rect 1895 8596 1911 8598
rect 1983 8596 2036 8610
rect 1984 8594 2048 8596
rect 2091 8594 2106 8610
rect 2155 8607 2185 8610
rect 2155 8604 2191 8607
rect 2121 8596 2137 8598
rect 1895 8584 1910 8588
rect 1813 8582 1910 8584
rect 1938 8582 2106 8594
rect 2122 8584 2137 8588
rect 2155 8585 2194 8604
rect 2213 8598 2220 8599
rect 2219 8591 2220 8598
rect 2203 8588 2204 8591
rect 2219 8588 2232 8591
rect 2155 8584 2185 8585
rect 2194 8584 2200 8585
rect 2203 8584 2232 8588
rect 2122 8583 2232 8584
rect 2122 8582 2238 8583
rect 1797 8574 1848 8582
rect 1797 8562 1822 8574
rect 1829 8562 1848 8574
rect 1879 8574 1929 8582
rect 1879 8566 1895 8574
rect 1902 8572 1929 8574
rect 1938 8572 2159 8582
rect 1902 8562 2159 8572
rect 2188 8574 2238 8582
rect 2188 8565 2204 8574
rect 1797 8554 1848 8562
rect 1895 8554 2159 8562
rect 2185 8562 2204 8565
rect 2211 8562 2238 8574
rect 2185 8554 2238 8562
rect 1813 8546 1814 8554
rect 1829 8546 1842 8554
rect 1813 8538 1829 8546
rect 1810 8531 1829 8534
rect 1810 8522 1832 8531
rect 1783 8512 1832 8522
rect 1783 8506 1813 8512
rect 1832 8507 1837 8512
rect 1755 8490 1829 8506
rect 1847 8498 1877 8554
rect 1912 8544 2120 8554
rect 2155 8550 2200 8554
rect 2203 8553 2204 8554
rect 2219 8553 2232 8554
rect 1938 8514 2127 8544
rect 1953 8511 2127 8514
rect 1946 8508 2127 8511
rect 1755 8488 1768 8490
rect 1783 8488 1817 8490
rect 1755 8472 1829 8488
rect 1856 8484 1869 8498
rect 1884 8484 1900 8500
rect 1946 8495 1957 8508
rect 1739 8450 1740 8466
rect 1755 8450 1768 8472
rect 1783 8450 1813 8472
rect 1856 8468 1918 8484
rect 1946 8477 1957 8493
rect 1962 8488 1972 8508
rect 1982 8488 1996 8508
rect 1999 8495 2008 8508
rect 2024 8495 2033 8508
rect 1962 8477 1996 8488
rect 1999 8477 2008 8493
rect 2024 8477 2033 8493
rect 2040 8488 2050 8508
rect 2060 8488 2074 8508
rect 2075 8495 2086 8508
rect 2040 8477 2074 8488
rect 2075 8477 2086 8493
rect 2132 8484 2148 8500
rect 2155 8498 2185 8550
rect 2219 8546 2220 8553
rect 2204 8538 2220 8546
rect 2191 8506 2204 8525
rect 2219 8506 2249 8522
rect 2191 8490 2265 8506
rect 2191 8488 2204 8490
rect 2219 8488 2253 8490
rect 1856 8466 1869 8468
rect 1884 8466 1918 8468
rect 1856 8450 1918 8466
rect 1962 8461 1978 8464
rect 2040 8461 2070 8472
rect 2118 8468 2164 8484
rect 2191 8472 2265 8488
rect 2118 8466 2152 8468
rect 2117 8450 2164 8466
rect 2191 8450 2204 8472
rect 2219 8450 2249 8472
rect 2276 8450 2277 8466
rect 2292 8450 2305 8610
rect 2335 8506 2348 8610
rect 2393 8588 2394 8598
rect 2409 8588 2422 8598
rect 2393 8584 2422 8588
rect 2427 8584 2457 8610
rect 2475 8596 2491 8598
rect 2563 8596 2616 8610
rect 2564 8594 2628 8596
rect 2671 8594 2686 8610
rect 2735 8607 2765 8610
rect 2735 8604 2771 8607
rect 2701 8596 2717 8598
rect 2475 8584 2490 8588
rect 2393 8582 2490 8584
rect 2518 8582 2686 8594
rect 2702 8584 2717 8588
rect 2735 8585 2774 8604
rect 2793 8598 2800 8599
rect 2799 8591 2800 8598
rect 2783 8588 2784 8591
rect 2799 8588 2812 8591
rect 2735 8584 2765 8585
rect 2774 8584 2780 8585
rect 2783 8584 2812 8588
rect 2702 8583 2812 8584
rect 2702 8582 2818 8583
rect 2377 8574 2428 8582
rect 2377 8562 2402 8574
rect 2409 8562 2428 8574
rect 2459 8574 2509 8582
rect 2459 8566 2475 8574
rect 2482 8572 2509 8574
rect 2518 8572 2739 8582
rect 2482 8562 2739 8572
rect 2768 8574 2818 8582
rect 2768 8565 2784 8574
rect 2377 8554 2428 8562
rect 2475 8554 2739 8562
rect 2765 8562 2784 8565
rect 2791 8562 2818 8574
rect 2765 8554 2818 8562
rect 2393 8546 2394 8554
rect 2409 8546 2422 8554
rect 2393 8538 2409 8546
rect 2390 8531 2409 8534
rect 2390 8522 2412 8531
rect 2363 8512 2412 8522
rect 2363 8506 2393 8512
rect 2412 8507 2417 8512
rect 2335 8490 2409 8506
rect 2427 8498 2457 8554
rect 2492 8544 2700 8554
rect 2735 8550 2780 8554
rect 2783 8553 2784 8554
rect 2799 8553 2812 8554
rect 2518 8514 2707 8544
rect 2533 8511 2707 8514
rect 2526 8508 2707 8511
rect 2335 8488 2348 8490
rect 2363 8488 2397 8490
rect 2335 8472 2409 8488
rect 2436 8484 2449 8498
rect 2464 8484 2480 8500
rect 2526 8495 2537 8508
rect 2319 8450 2320 8466
rect 2335 8450 2348 8472
rect 2363 8450 2393 8472
rect 2436 8468 2498 8484
rect 2526 8477 2537 8493
rect 2542 8488 2552 8508
rect 2562 8488 2576 8508
rect 2579 8495 2588 8508
rect 2604 8495 2613 8508
rect 2542 8477 2576 8488
rect 2579 8477 2588 8493
rect 2604 8477 2613 8493
rect 2620 8488 2630 8508
rect 2640 8488 2654 8508
rect 2655 8495 2666 8508
rect 2620 8477 2654 8488
rect 2655 8477 2666 8493
rect 2712 8484 2728 8500
rect 2735 8498 2765 8550
rect 2799 8546 2800 8553
rect 2784 8538 2800 8546
rect 2771 8506 2784 8525
rect 2799 8506 2829 8522
rect 2771 8490 2845 8506
rect 2771 8488 2784 8490
rect 2799 8488 2833 8490
rect 2436 8466 2449 8468
rect 2464 8466 2498 8468
rect 2436 8450 2498 8466
rect 2542 8461 2558 8464
rect 2620 8461 2650 8472
rect 2698 8468 2744 8484
rect 2771 8472 2845 8488
rect 2698 8466 2732 8468
rect 2697 8450 2744 8466
rect 2771 8450 2784 8472
rect 2799 8450 2829 8472
rect 2856 8450 2857 8466
rect 2872 8450 2885 8610
rect 2915 8506 2928 8610
rect 2973 8588 2974 8598
rect 2989 8588 3002 8598
rect 2973 8584 3002 8588
rect 3007 8584 3037 8610
rect 3055 8596 3071 8598
rect 3143 8596 3196 8610
rect 3144 8594 3208 8596
rect 3251 8594 3266 8610
rect 3315 8607 3345 8610
rect 3315 8604 3351 8607
rect 3281 8596 3297 8598
rect 3055 8584 3070 8588
rect 2973 8582 3070 8584
rect 3098 8582 3266 8594
rect 3282 8584 3297 8588
rect 3315 8585 3354 8604
rect 3373 8598 3380 8599
rect 3379 8591 3380 8598
rect 3363 8588 3364 8591
rect 3379 8588 3392 8591
rect 3315 8584 3345 8585
rect 3354 8584 3360 8585
rect 3363 8584 3392 8588
rect 3282 8583 3392 8584
rect 3282 8582 3398 8583
rect 2957 8574 3008 8582
rect 2957 8562 2982 8574
rect 2989 8562 3008 8574
rect 3039 8574 3089 8582
rect 3039 8566 3055 8574
rect 3062 8572 3089 8574
rect 3098 8572 3319 8582
rect 3062 8562 3319 8572
rect 3348 8574 3398 8582
rect 3348 8565 3364 8574
rect 2957 8554 3008 8562
rect 3055 8554 3319 8562
rect 3345 8562 3364 8565
rect 3371 8562 3398 8574
rect 3345 8554 3398 8562
rect 2973 8546 2974 8554
rect 2989 8546 3002 8554
rect 2973 8538 2989 8546
rect 2970 8531 2989 8534
rect 2970 8522 2992 8531
rect 2943 8512 2992 8522
rect 2943 8506 2973 8512
rect 2992 8507 2997 8512
rect 2915 8490 2989 8506
rect 3007 8498 3037 8554
rect 3072 8544 3280 8554
rect 3315 8550 3360 8554
rect 3363 8553 3364 8554
rect 3379 8553 3392 8554
rect 3098 8514 3287 8544
rect 3113 8511 3287 8514
rect 3106 8508 3287 8511
rect 2915 8488 2928 8490
rect 2943 8488 2977 8490
rect 2915 8472 2989 8488
rect 3016 8484 3029 8498
rect 3044 8484 3060 8500
rect 3106 8495 3117 8508
rect 2899 8450 2900 8466
rect 2915 8450 2928 8472
rect 2943 8450 2973 8472
rect 3016 8468 3078 8484
rect 3106 8477 3117 8493
rect 3122 8488 3132 8508
rect 3142 8488 3156 8508
rect 3159 8495 3168 8508
rect 3184 8495 3193 8508
rect 3122 8477 3156 8488
rect 3159 8477 3168 8493
rect 3184 8477 3193 8493
rect 3200 8488 3210 8508
rect 3220 8488 3234 8508
rect 3235 8495 3246 8508
rect 3200 8477 3234 8488
rect 3235 8477 3246 8493
rect 3292 8484 3308 8500
rect 3315 8498 3345 8550
rect 3379 8546 3380 8553
rect 3364 8538 3380 8546
rect 3351 8506 3364 8525
rect 3379 8506 3409 8522
rect 3351 8490 3425 8506
rect 3351 8488 3364 8490
rect 3379 8488 3413 8490
rect 3016 8466 3029 8468
rect 3044 8466 3078 8468
rect 3016 8450 3078 8466
rect 3122 8461 3138 8464
rect 3200 8461 3230 8472
rect 3278 8468 3324 8484
rect 3351 8472 3425 8488
rect 3278 8466 3312 8468
rect 3277 8450 3324 8466
rect 3351 8450 3364 8472
rect 3379 8450 3409 8472
rect 3436 8450 3437 8466
rect 3452 8450 3465 8610
rect 3495 8506 3508 8610
rect 3553 8588 3554 8598
rect 3569 8588 3582 8598
rect 3553 8584 3582 8588
rect 3587 8584 3617 8610
rect 3635 8596 3651 8598
rect 3723 8596 3776 8610
rect 3724 8594 3788 8596
rect 3831 8594 3846 8610
rect 3895 8607 3925 8610
rect 3895 8604 3931 8607
rect 3861 8596 3877 8598
rect 3635 8584 3650 8588
rect 3553 8582 3650 8584
rect 3678 8582 3846 8594
rect 3862 8584 3877 8588
rect 3895 8585 3934 8604
rect 3953 8598 3960 8599
rect 3959 8591 3960 8598
rect 3943 8588 3944 8591
rect 3959 8588 3972 8591
rect 3895 8584 3925 8585
rect 3934 8584 3940 8585
rect 3943 8584 3972 8588
rect 3862 8583 3972 8584
rect 3862 8582 3978 8583
rect 3537 8574 3588 8582
rect 3537 8562 3562 8574
rect 3569 8562 3588 8574
rect 3619 8574 3669 8582
rect 3619 8566 3635 8574
rect 3642 8572 3669 8574
rect 3678 8572 3899 8582
rect 3642 8562 3899 8572
rect 3928 8574 3978 8582
rect 3928 8565 3944 8574
rect 3537 8554 3588 8562
rect 3635 8554 3899 8562
rect 3925 8562 3944 8565
rect 3951 8562 3978 8574
rect 3925 8554 3978 8562
rect 3553 8546 3554 8554
rect 3569 8546 3582 8554
rect 3553 8538 3569 8546
rect 3550 8531 3569 8534
rect 3550 8522 3572 8531
rect 3523 8512 3572 8522
rect 3523 8506 3553 8512
rect 3572 8507 3577 8512
rect 3495 8490 3569 8506
rect 3587 8498 3617 8554
rect 3652 8544 3860 8554
rect 3895 8550 3940 8554
rect 3943 8553 3944 8554
rect 3959 8553 3972 8554
rect 3678 8514 3867 8544
rect 3693 8511 3867 8514
rect 3686 8508 3867 8511
rect 3495 8488 3508 8490
rect 3523 8488 3557 8490
rect 3495 8472 3569 8488
rect 3596 8484 3609 8498
rect 3624 8484 3640 8500
rect 3686 8495 3697 8508
rect 3479 8450 3480 8466
rect 3495 8450 3508 8472
rect 3523 8450 3553 8472
rect 3596 8468 3658 8484
rect 3686 8477 3697 8493
rect 3702 8488 3712 8508
rect 3722 8488 3736 8508
rect 3739 8495 3748 8508
rect 3764 8495 3773 8508
rect 3702 8477 3736 8488
rect 3739 8477 3748 8493
rect 3764 8477 3773 8493
rect 3780 8488 3790 8508
rect 3800 8488 3814 8508
rect 3815 8495 3826 8508
rect 3780 8477 3814 8488
rect 3815 8477 3826 8493
rect 3872 8484 3888 8500
rect 3895 8498 3925 8550
rect 3959 8546 3960 8553
rect 3944 8538 3960 8546
rect 3931 8506 3944 8525
rect 3959 8506 3989 8522
rect 3931 8490 4005 8506
rect 3931 8488 3944 8490
rect 3959 8488 3993 8490
rect 3596 8466 3609 8468
rect 3624 8466 3658 8468
rect 3596 8450 3658 8466
rect 3702 8461 3718 8464
rect 3780 8461 3810 8472
rect 3858 8468 3904 8484
rect 3931 8472 4005 8488
rect 3858 8466 3892 8468
rect 3857 8450 3904 8466
rect 3931 8450 3944 8472
rect 3959 8450 3989 8472
rect 4016 8450 4017 8466
rect 4032 8450 4045 8610
rect 4075 8506 4088 8610
rect 4133 8588 4134 8598
rect 4149 8588 4162 8598
rect 4133 8584 4162 8588
rect 4167 8584 4197 8610
rect 4215 8596 4231 8598
rect 4303 8596 4356 8610
rect 4304 8594 4368 8596
rect 4411 8594 4426 8610
rect 4475 8607 4505 8610
rect 4475 8604 4511 8607
rect 4441 8596 4457 8598
rect 4215 8584 4230 8588
rect 4133 8582 4230 8584
rect 4258 8582 4426 8594
rect 4442 8584 4457 8588
rect 4475 8585 4514 8604
rect 4533 8598 4540 8599
rect 4539 8591 4540 8598
rect 4523 8588 4524 8591
rect 4539 8588 4552 8591
rect 4475 8584 4505 8585
rect 4514 8584 4520 8585
rect 4523 8584 4552 8588
rect 4442 8583 4552 8584
rect 4442 8582 4558 8583
rect 4117 8574 4168 8582
rect 4117 8562 4142 8574
rect 4149 8562 4168 8574
rect 4199 8574 4249 8582
rect 4199 8566 4215 8574
rect 4222 8572 4249 8574
rect 4258 8572 4479 8582
rect 4222 8562 4479 8572
rect 4508 8574 4558 8582
rect 4508 8565 4524 8574
rect 4117 8554 4168 8562
rect 4215 8554 4479 8562
rect 4505 8562 4524 8565
rect 4531 8562 4558 8574
rect 4505 8554 4558 8562
rect 4133 8546 4134 8554
rect 4149 8546 4162 8554
rect 4133 8538 4149 8546
rect 4130 8531 4149 8534
rect 4130 8522 4152 8531
rect 4103 8512 4152 8522
rect 4103 8506 4133 8512
rect 4152 8507 4157 8512
rect 4075 8490 4149 8506
rect 4167 8498 4197 8554
rect 4232 8544 4440 8554
rect 4475 8550 4520 8554
rect 4523 8553 4524 8554
rect 4539 8553 4552 8554
rect 4258 8514 4447 8544
rect 4273 8511 4447 8514
rect 4266 8508 4447 8511
rect 4075 8488 4088 8490
rect 4103 8488 4137 8490
rect 4075 8472 4149 8488
rect 4176 8484 4189 8498
rect 4204 8484 4220 8500
rect 4266 8495 4277 8508
rect 4059 8450 4060 8466
rect 4075 8450 4088 8472
rect 4103 8450 4133 8472
rect 4176 8468 4238 8484
rect 4266 8477 4277 8493
rect 4282 8488 4292 8508
rect 4302 8488 4316 8508
rect 4319 8495 4328 8508
rect 4344 8495 4353 8508
rect 4282 8477 4316 8488
rect 4319 8477 4328 8493
rect 4344 8477 4353 8493
rect 4360 8488 4370 8508
rect 4380 8488 4394 8508
rect 4395 8495 4406 8508
rect 4360 8477 4394 8488
rect 4395 8477 4406 8493
rect 4452 8484 4468 8500
rect 4475 8498 4505 8550
rect 4539 8546 4540 8553
rect 4524 8538 4540 8546
rect 4511 8506 4524 8525
rect 4539 8506 4569 8522
rect 4511 8490 4585 8506
rect 4511 8488 4524 8490
rect 4539 8488 4573 8490
rect 4176 8466 4189 8468
rect 4204 8466 4238 8468
rect 4176 8450 4238 8466
rect 4282 8461 4298 8464
rect 4360 8461 4390 8472
rect 4438 8468 4484 8484
rect 4511 8472 4585 8488
rect 4438 8466 4472 8468
rect 4437 8450 4484 8466
rect 4511 8450 4524 8472
rect 4539 8450 4569 8472
rect 4596 8450 4597 8466
rect 4612 8450 4625 8610
rect -7 8442 34 8450
rect -7 8416 8 8442
rect 15 8416 34 8442
rect 98 8438 160 8450
rect 172 8438 247 8450
rect 305 8438 380 8450
rect 392 8438 423 8450
rect 429 8438 464 8450
rect 98 8436 260 8438
rect -7 8408 34 8416
rect 116 8412 129 8436
rect 144 8434 159 8436
rect -1 8398 0 8408
rect 15 8398 28 8408
rect 43 8398 73 8412
rect 116 8398 159 8412
rect 183 8409 190 8416
rect 193 8412 260 8436
rect 292 8436 464 8438
rect 262 8414 290 8418
rect 292 8414 372 8436
rect 393 8434 408 8436
rect 262 8412 372 8414
rect 193 8408 372 8412
rect 166 8398 196 8408
rect 198 8398 351 8408
rect 359 8398 389 8408
rect 393 8398 423 8412
rect 451 8398 464 8436
rect 536 8442 571 8450
rect 536 8416 537 8442
rect 544 8416 571 8442
rect 479 8398 509 8412
rect 536 8408 571 8416
rect 573 8442 614 8450
rect 573 8416 588 8442
rect 595 8416 614 8442
rect 678 8438 740 8450
rect 752 8438 827 8450
rect 885 8438 960 8450
rect 972 8438 1003 8450
rect 1009 8438 1044 8450
rect 678 8436 840 8438
rect 573 8408 614 8416
rect 696 8412 709 8436
rect 724 8434 739 8436
rect 536 8398 537 8408
rect 552 8398 565 8408
rect 579 8398 580 8408
rect 595 8398 608 8408
rect 623 8398 653 8412
rect 696 8398 739 8412
rect 763 8409 770 8416
rect 773 8412 840 8436
rect 872 8436 1044 8438
rect 842 8414 870 8418
rect 872 8414 952 8436
rect 973 8434 988 8436
rect 842 8412 952 8414
rect 773 8408 952 8412
rect 746 8398 776 8408
rect 778 8398 931 8408
rect 939 8398 969 8408
rect 973 8398 1003 8412
rect 1031 8398 1044 8436
rect 1116 8442 1151 8450
rect 1116 8416 1117 8442
rect 1124 8416 1151 8442
rect 1059 8398 1089 8412
rect 1116 8408 1151 8416
rect 1153 8442 1194 8450
rect 1153 8416 1168 8442
rect 1175 8416 1194 8442
rect 1258 8438 1320 8450
rect 1332 8438 1407 8450
rect 1465 8438 1540 8450
rect 1552 8438 1583 8450
rect 1589 8438 1624 8450
rect 1258 8436 1420 8438
rect 1153 8408 1194 8416
rect 1276 8412 1289 8436
rect 1304 8434 1319 8436
rect 1116 8398 1117 8408
rect 1132 8398 1145 8408
rect 1159 8398 1160 8408
rect 1175 8398 1188 8408
rect 1203 8398 1233 8412
rect 1276 8398 1319 8412
rect 1343 8409 1350 8416
rect 1353 8412 1420 8436
rect 1452 8436 1624 8438
rect 1422 8414 1450 8418
rect 1452 8414 1532 8436
rect 1553 8434 1568 8436
rect 1422 8412 1532 8414
rect 1353 8408 1532 8412
rect 1326 8398 1356 8408
rect 1358 8398 1511 8408
rect 1519 8398 1549 8408
rect 1553 8398 1583 8412
rect 1611 8398 1624 8436
rect 1696 8442 1731 8450
rect 1696 8416 1697 8442
rect 1704 8416 1731 8442
rect 1639 8398 1669 8412
rect 1696 8408 1731 8416
rect 1733 8442 1774 8450
rect 1733 8416 1748 8442
rect 1755 8416 1774 8442
rect 1838 8438 1900 8450
rect 1912 8438 1987 8450
rect 2045 8438 2120 8450
rect 2132 8438 2163 8450
rect 2169 8438 2204 8450
rect 1838 8436 2000 8438
rect 1733 8408 1774 8416
rect 1856 8412 1869 8436
rect 1884 8434 1899 8436
rect 1696 8398 1697 8408
rect 1712 8398 1725 8408
rect 1739 8398 1740 8408
rect 1755 8398 1768 8408
rect 1783 8398 1813 8412
rect 1856 8398 1899 8412
rect 1923 8409 1930 8416
rect 1933 8412 2000 8436
rect 2032 8436 2204 8438
rect 2002 8414 2030 8418
rect 2032 8414 2112 8436
rect 2133 8434 2148 8436
rect 2002 8412 2112 8414
rect 1933 8408 2112 8412
rect 1906 8398 1936 8408
rect 1938 8398 2091 8408
rect 2099 8398 2129 8408
rect 2133 8398 2163 8412
rect 2191 8398 2204 8436
rect 2276 8442 2311 8450
rect 2276 8416 2277 8442
rect 2284 8416 2311 8442
rect 2219 8398 2249 8412
rect 2276 8408 2311 8416
rect 2313 8442 2354 8450
rect 2313 8416 2328 8442
rect 2335 8416 2354 8442
rect 2418 8438 2480 8450
rect 2492 8438 2567 8450
rect 2625 8438 2700 8450
rect 2712 8438 2743 8450
rect 2749 8438 2784 8450
rect 2418 8436 2580 8438
rect 2313 8408 2354 8416
rect 2436 8412 2449 8436
rect 2464 8434 2479 8436
rect 2276 8398 2277 8408
rect 2292 8398 2305 8408
rect 2319 8398 2320 8408
rect 2335 8398 2348 8408
rect 2363 8398 2393 8412
rect 2436 8398 2479 8412
rect 2503 8409 2510 8416
rect 2513 8412 2580 8436
rect 2612 8436 2784 8438
rect 2582 8414 2610 8418
rect 2612 8414 2692 8436
rect 2713 8434 2728 8436
rect 2582 8412 2692 8414
rect 2513 8408 2692 8412
rect 2486 8398 2516 8408
rect 2518 8398 2671 8408
rect 2679 8398 2709 8408
rect 2713 8398 2743 8412
rect 2771 8398 2784 8436
rect 2856 8442 2891 8450
rect 2856 8416 2857 8442
rect 2864 8416 2891 8442
rect 2799 8398 2829 8412
rect 2856 8408 2891 8416
rect 2893 8442 2934 8450
rect 2893 8416 2908 8442
rect 2915 8416 2934 8442
rect 2998 8438 3060 8450
rect 3072 8438 3147 8450
rect 3205 8438 3280 8450
rect 3292 8438 3323 8450
rect 3329 8438 3364 8450
rect 2998 8436 3160 8438
rect 2893 8408 2934 8416
rect 3016 8412 3029 8436
rect 3044 8434 3059 8436
rect 2856 8398 2857 8408
rect 2872 8398 2885 8408
rect 2899 8398 2900 8408
rect 2915 8398 2928 8408
rect 2943 8398 2973 8412
rect 3016 8398 3059 8412
rect 3083 8409 3090 8416
rect 3093 8412 3160 8436
rect 3192 8436 3364 8438
rect 3162 8414 3190 8418
rect 3192 8414 3272 8436
rect 3293 8434 3308 8436
rect 3162 8412 3272 8414
rect 3093 8408 3272 8412
rect 3066 8398 3096 8408
rect 3098 8398 3251 8408
rect 3259 8398 3289 8408
rect 3293 8398 3323 8412
rect 3351 8398 3364 8436
rect 3436 8442 3471 8450
rect 3436 8416 3437 8442
rect 3444 8416 3471 8442
rect 3379 8398 3409 8412
rect 3436 8408 3471 8416
rect 3473 8442 3514 8450
rect 3473 8416 3488 8442
rect 3495 8416 3514 8442
rect 3578 8438 3640 8450
rect 3652 8438 3727 8450
rect 3785 8438 3860 8450
rect 3872 8438 3903 8450
rect 3909 8438 3944 8450
rect 3578 8436 3740 8438
rect 3473 8408 3514 8416
rect 3596 8412 3609 8436
rect 3624 8434 3639 8436
rect 3436 8398 3437 8408
rect 3452 8398 3465 8408
rect 3479 8398 3480 8408
rect 3495 8398 3508 8408
rect 3523 8398 3553 8412
rect 3596 8398 3639 8412
rect 3663 8409 3670 8416
rect 3673 8412 3740 8436
rect 3772 8436 3944 8438
rect 3742 8414 3770 8418
rect 3772 8414 3852 8436
rect 3873 8434 3888 8436
rect 3742 8412 3852 8414
rect 3673 8408 3852 8412
rect 3646 8398 3676 8408
rect 3678 8398 3831 8408
rect 3839 8398 3869 8408
rect 3873 8398 3903 8412
rect 3931 8398 3944 8436
rect 4016 8442 4051 8450
rect 4016 8416 4017 8442
rect 4024 8416 4051 8442
rect 3959 8398 3989 8412
rect 4016 8408 4051 8416
rect 4053 8442 4094 8450
rect 4053 8416 4068 8442
rect 4075 8416 4094 8442
rect 4158 8438 4220 8450
rect 4232 8438 4307 8450
rect 4365 8438 4440 8450
rect 4452 8438 4483 8450
rect 4489 8438 4524 8450
rect 4158 8436 4320 8438
rect 4053 8408 4094 8416
rect 4176 8412 4189 8436
rect 4204 8434 4219 8436
rect 4016 8398 4017 8408
rect 4032 8398 4045 8408
rect 4059 8398 4060 8408
rect 4075 8398 4088 8408
rect 4103 8398 4133 8412
rect 4176 8398 4219 8412
rect 4243 8409 4250 8416
rect 4253 8412 4320 8436
rect 4352 8436 4524 8438
rect 4322 8414 4350 8418
rect 4352 8414 4432 8436
rect 4453 8434 4468 8436
rect 4322 8412 4432 8414
rect 4253 8408 4432 8412
rect 4226 8398 4256 8408
rect 4258 8398 4411 8408
rect 4419 8398 4449 8408
rect 4453 8398 4483 8412
rect 4511 8398 4524 8436
rect 4596 8442 4631 8450
rect 4596 8416 4597 8442
rect 4604 8416 4631 8442
rect 4539 8398 4569 8412
rect 4596 8408 4631 8416
rect 4596 8398 4597 8408
rect 4612 8398 4625 8408
rect -1 8392 4625 8398
rect 0 8384 4625 8392
rect 15 8354 28 8384
rect 43 8366 73 8384
rect 116 8370 130 8384
rect 166 8370 386 8384
rect 117 8368 130 8370
rect 83 8356 98 8368
rect 80 8354 102 8356
rect 107 8354 137 8368
rect 198 8366 351 8370
rect 180 8354 372 8366
rect 415 8354 445 8368
rect 451 8354 464 8384
rect 479 8366 509 8384
rect 552 8354 565 8384
rect 595 8354 608 8384
rect 623 8366 653 8384
rect 696 8370 710 8384
rect 746 8370 966 8384
rect 697 8368 710 8370
rect 663 8356 678 8368
rect 660 8354 682 8356
rect 687 8354 717 8368
rect 778 8366 931 8370
rect 760 8354 952 8366
rect 995 8354 1025 8368
rect 1031 8354 1044 8384
rect 1059 8366 1089 8384
rect 1132 8354 1145 8384
rect 1175 8354 1188 8384
rect 1203 8366 1233 8384
rect 1276 8370 1290 8384
rect 1326 8370 1546 8384
rect 1277 8368 1290 8370
rect 1243 8356 1258 8368
rect 1240 8354 1262 8356
rect 1267 8354 1297 8368
rect 1358 8366 1511 8370
rect 1340 8354 1532 8366
rect 1575 8354 1605 8368
rect 1611 8354 1624 8384
rect 1639 8366 1669 8384
rect 1712 8354 1725 8384
rect 1755 8354 1768 8384
rect 1783 8366 1813 8384
rect 1856 8370 1870 8384
rect 1906 8370 2126 8384
rect 1857 8368 1870 8370
rect 1823 8356 1838 8368
rect 1820 8354 1842 8356
rect 1847 8354 1877 8368
rect 1938 8366 2091 8370
rect 1920 8354 2112 8366
rect 2155 8354 2185 8368
rect 2191 8354 2204 8384
rect 2219 8366 2249 8384
rect 2292 8354 2305 8384
rect 2335 8354 2348 8384
rect 2363 8366 2393 8384
rect 2436 8370 2450 8384
rect 2486 8370 2706 8384
rect 2437 8368 2450 8370
rect 2403 8356 2418 8368
rect 2400 8354 2422 8356
rect 2427 8354 2457 8368
rect 2518 8366 2671 8370
rect 2500 8354 2692 8366
rect 2735 8354 2765 8368
rect 2771 8354 2784 8384
rect 2799 8366 2829 8384
rect 2872 8354 2885 8384
rect 2915 8354 2928 8384
rect 2943 8366 2973 8384
rect 3016 8370 3030 8384
rect 3066 8370 3286 8384
rect 3017 8368 3030 8370
rect 2983 8356 2998 8368
rect 2980 8354 3002 8356
rect 3007 8354 3037 8368
rect 3098 8366 3251 8370
rect 3080 8354 3272 8366
rect 3315 8354 3345 8368
rect 3351 8354 3364 8384
rect 3379 8366 3409 8384
rect 3452 8354 3465 8384
rect 3495 8354 3508 8384
rect 3523 8366 3553 8384
rect 3596 8370 3610 8384
rect 3646 8370 3866 8384
rect 3597 8368 3610 8370
rect 3563 8356 3578 8368
rect 3560 8354 3582 8356
rect 3587 8354 3617 8368
rect 3678 8366 3831 8370
rect 3660 8354 3852 8366
rect 3895 8354 3925 8368
rect 3931 8354 3944 8384
rect 3959 8366 3989 8384
rect 4032 8354 4045 8384
rect 4075 8354 4088 8384
rect 4103 8366 4133 8384
rect 4176 8370 4190 8384
rect 4226 8370 4446 8384
rect 4177 8368 4190 8370
rect 4143 8356 4158 8368
rect 4140 8354 4162 8356
rect 4167 8354 4197 8368
rect 4258 8366 4411 8370
rect 4240 8354 4432 8366
rect 4475 8354 4505 8368
rect 4511 8354 4524 8384
rect 4539 8366 4569 8384
rect 4612 8354 4625 8384
rect 0 8340 4625 8354
rect 15 8236 28 8340
rect 73 8318 74 8328
rect 89 8318 102 8328
rect 73 8314 102 8318
rect 107 8314 137 8340
rect 155 8326 171 8328
rect 243 8326 296 8340
rect 244 8324 308 8326
rect 351 8324 366 8340
rect 415 8337 445 8340
rect 415 8334 451 8337
rect 381 8326 397 8328
rect 155 8314 170 8318
rect 73 8312 170 8314
rect 198 8312 366 8324
rect 382 8314 397 8318
rect 415 8315 454 8334
rect 473 8328 480 8329
rect 479 8321 480 8328
rect 463 8318 464 8321
rect 479 8318 492 8321
rect 415 8314 445 8315
rect 454 8314 460 8315
rect 463 8314 492 8318
rect 382 8313 492 8314
rect 382 8312 498 8313
rect 57 8304 108 8312
rect 57 8292 82 8304
rect 89 8292 108 8304
rect 139 8304 189 8312
rect 139 8296 155 8304
rect 162 8302 189 8304
rect 198 8302 419 8312
rect 162 8292 419 8302
rect 448 8304 498 8312
rect 448 8295 464 8304
rect 57 8284 108 8292
rect 155 8284 419 8292
rect 445 8292 464 8295
rect 471 8292 498 8304
rect 445 8284 498 8292
rect 73 8276 74 8284
rect 89 8276 102 8284
rect 73 8268 89 8276
rect 70 8261 89 8264
rect 70 8252 92 8261
rect 43 8242 92 8252
rect 43 8236 73 8242
rect 92 8237 97 8242
rect 15 8220 89 8236
rect 107 8228 137 8284
rect 172 8274 380 8284
rect 415 8280 460 8284
rect 463 8283 464 8284
rect 479 8283 492 8284
rect 198 8244 387 8274
rect 213 8241 387 8244
rect 206 8238 387 8241
rect 15 8218 28 8220
rect 43 8218 77 8220
rect 15 8202 89 8218
rect 116 8214 129 8228
rect 144 8214 160 8230
rect 206 8225 217 8238
rect -1 8180 0 8196
rect 15 8180 28 8202
rect 43 8180 73 8202
rect 116 8198 178 8214
rect 206 8207 217 8223
rect 222 8218 232 8238
rect 242 8218 256 8238
rect 259 8225 268 8238
rect 284 8225 293 8238
rect 222 8207 256 8218
rect 259 8207 268 8223
rect 284 8207 293 8223
rect 300 8218 310 8238
rect 320 8218 334 8238
rect 335 8225 346 8238
rect 300 8207 334 8218
rect 335 8207 346 8223
rect 392 8214 408 8230
rect 415 8228 445 8280
rect 479 8276 480 8283
rect 464 8268 480 8276
rect 451 8236 464 8255
rect 479 8236 509 8252
rect 451 8220 525 8236
rect 451 8218 464 8220
rect 479 8218 513 8220
rect 116 8196 129 8198
rect 144 8196 178 8198
rect 116 8180 178 8196
rect 222 8191 238 8194
rect 300 8191 330 8202
rect 378 8198 424 8214
rect 451 8202 525 8218
rect 378 8196 412 8198
rect 377 8180 424 8196
rect 451 8180 464 8202
rect 479 8180 509 8202
rect 536 8180 537 8196
rect 552 8180 565 8340
rect 595 8236 608 8340
rect 653 8318 654 8328
rect 669 8318 682 8328
rect 653 8314 682 8318
rect 687 8314 717 8340
rect 735 8326 751 8328
rect 823 8326 876 8340
rect 824 8324 888 8326
rect 931 8324 946 8340
rect 995 8337 1025 8340
rect 995 8334 1031 8337
rect 961 8326 977 8328
rect 735 8314 750 8318
rect 653 8312 750 8314
rect 778 8312 946 8324
rect 962 8314 977 8318
rect 995 8315 1034 8334
rect 1053 8328 1060 8329
rect 1059 8321 1060 8328
rect 1043 8318 1044 8321
rect 1059 8318 1072 8321
rect 995 8314 1025 8315
rect 1034 8314 1040 8315
rect 1043 8314 1072 8318
rect 962 8313 1072 8314
rect 962 8312 1078 8313
rect 637 8304 688 8312
rect 637 8292 662 8304
rect 669 8292 688 8304
rect 719 8304 769 8312
rect 719 8296 735 8304
rect 742 8302 769 8304
rect 778 8302 999 8312
rect 742 8292 999 8302
rect 1028 8304 1078 8312
rect 1028 8295 1044 8304
rect 637 8284 688 8292
rect 735 8284 999 8292
rect 1025 8292 1044 8295
rect 1051 8292 1078 8304
rect 1025 8284 1078 8292
rect 653 8276 654 8284
rect 669 8276 682 8284
rect 653 8268 669 8276
rect 650 8261 669 8264
rect 650 8252 672 8261
rect 623 8242 672 8252
rect 623 8236 653 8242
rect 672 8237 677 8242
rect 595 8220 669 8236
rect 687 8228 717 8284
rect 752 8274 960 8284
rect 995 8280 1040 8284
rect 1043 8283 1044 8284
rect 1059 8283 1072 8284
rect 778 8244 967 8274
rect 793 8241 967 8244
rect 786 8238 967 8241
rect 595 8218 608 8220
rect 623 8218 657 8220
rect 595 8202 669 8218
rect 696 8214 709 8228
rect 724 8214 740 8230
rect 786 8225 797 8238
rect 579 8180 580 8196
rect 595 8180 608 8202
rect 623 8180 653 8202
rect 696 8198 758 8214
rect 786 8207 797 8223
rect 802 8218 812 8238
rect 822 8218 836 8238
rect 839 8225 848 8238
rect 864 8225 873 8238
rect 802 8207 836 8218
rect 839 8207 848 8223
rect 864 8207 873 8223
rect 880 8218 890 8238
rect 900 8218 914 8238
rect 915 8225 926 8238
rect 880 8207 914 8218
rect 915 8207 926 8223
rect 972 8214 988 8230
rect 995 8228 1025 8280
rect 1059 8276 1060 8283
rect 1044 8268 1060 8276
rect 1031 8236 1044 8255
rect 1059 8236 1089 8252
rect 1031 8220 1105 8236
rect 1031 8218 1044 8220
rect 1059 8218 1093 8220
rect 696 8196 709 8198
rect 724 8196 758 8198
rect 696 8180 758 8196
rect 802 8191 818 8194
rect 880 8191 910 8202
rect 958 8198 1004 8214
rect 1031 8202 1105 8218
rect 958 8196 992 8198
rect 957 8180 1004 8196
rect 1031 8180 1044 8202
rect 1059 8180 1089 8202
rect 1116 8180 1117 8196
rect 1132 8180 1145 8340
rect 1175 8236 1188 8340
rect 1233 8318 1234 8328
rect 1249 8318 1262 8328
rect 1233 8314 1262 8318
rect 1267 8314 1297 8340
rect 1315 8326 1331 8328
rect 1403 8326 1456 8340
rect 1404 8324 1468 8326
rect 1511 8324 1526 8340
rect 1575 8337 1605 8340
rect 1575 8334 1611 8337
rect 1541 8326 1557 8328
rect 1315 8314 1330 8318
rect 1233 8312 1330 8314
rect 1358 8312 1526 8324
rect 1542 8314 1557 8318
rect 1575 8315 1614 8334
rect 1633 8328 1640 8329
rect 1639 8321 1640 8328
rect 1623 8318 1624 8321
rect 1639 8318 1652 8321
rect 1575 8314 1605 8315
rect 1614 8314 1620 8315
rect 1623 8314 1652 8318
rect 1542 8313 1652 8314
rect 1542 8312 1658 8313
rect 1217 8304 1268 8312
rect 1217 8292 1242 8304
rect 1249 8292 1268 8304
rect 1299 8304 1349 8312
rect 1299 8296 1315 8304
rect 1322 8302 1349 8304
rect 1358 8302 1579 8312
rect 1322 8292 1579 8302
rect 1608 8304 1658 8312
rect 1608 8295 1624 8304
rect 1217 8284 1268 8292
rect 1315 8284 1579 8292
rect 1605 8292 1624 8295
rect 1631 8292 1658 8304
rect 1605 8284 1658 8292
rect 1233 8276 1234 8284
rect 1249 8276 1262 8284
rect 1233 8268 1249 8276
rect 1230 8261 1249 8264
rect 1230 8252 1252 8261
rect 1203 8242 1252 8252
rect 1203 8236 1233 8242
rect 1252 8237 1257 8242
rect 1175 8220 1249 8236
rect 1267 8228 1297 8284
rect 1332 8274 1540 8284
rect 1575 8280 1620 8284
rect 1623 8283 1624 8284
rect 1639 8283 1652 8284
rect 1358 8244 1547 8274
rect 1373 8241 1547 8244
rect 1366 8238 1547 8241
rect 1175 8218 1188 8220
rect 1203 8218 1237 8220
rect 1175 8202 1249 8218
rect 1276 8214 1289 8228
rect 1304 8214 1320 8230
rect 1366 8225 1377 8238
rect 1159 8180 1160 8196
rect 1175 8180 1188 8202
rect 1203 8180 1233 8202
rect 1276 8198 1338 8214
rect 1366 8207 1377 8223
rect 1382 8218 1392 8238
rect 1402 8218 1416 8238
rect 1419 8225 1428 8238
rect 1444 8225 1453 8238
rect 1382 8207 1416 8218
rect 1419 8207 1428 8223
rect 1444 8207 1453 8223
rect 1460 8218 1470 8238
rect 1480 8218 1494 8238
rect 1495 8225 1506 8238
rect 1460 8207 1494 8218
rect 1495 8207 1506 8223
rect 1552 8214 1568 8230
rect 1575 8228 1605 8280
rect 1639 8276 1640 8283
rect 1624 8268 1640 8276
rect 1611 8236 1624 8255
rect 1639 8236 1669 8252
rect 1611 8220 1685 8236
rect 1611 8218 1624 8220
rect 1639 8218 1673 8220
rect 1276 8196 1289 8198
rect 1304 8196 1338 8198
rect 1276 8180 1338 8196
rect 1382 8191 1398 8194
rect 1460 8191 1490 8202
rect 1538 8198 1584 8214
rect 1611 8202 1685 8218
rect 1538 8196 1572 8198
rect 1537 8180 1584 8196
rect 1611 8180 1624 8202
rect 1639 8180 1669 8202
rect 1696 8180 1697 8196
rect 1712 8180 1725 8340
rect 1755 8236 1768 8340
rect 1813 8318 1814 8328
rect 1829 8318 1842 8328
rect 1813 8314 1842 8318
rect 1847 8314 1877 8340
rect 1895 8326 1911 8328
rect 1983 8326 2036 8340
rect 1984 8324 2048 8326
rect 2091 8324 2106 8340
rect 2155 8337 2185 8340
rect 2155 8334 2191 8337
rect 2121 8326 2137 8328
rect 1895 8314 1910 8318
rect 1813 8312 1910 8314
rect 1938 8312 2106 8324
rect 2122 8314 2137 8318
rect 2155 8315 2194 8334
rect 2213 8328 2220 8329
rect 2219 8321 2220 8328
rect 2203 8318 2204 8321
rect 2219 8318 2232 8321
rect 2155 8314 2185 8315
rect 2194 8314 2200 8315
rect 2203 8314 2232 8318
rect 2122 8313 2232 8314
rect 2122 8312 2238 8313
rect 1797 8304 1848 8312
rect 1797 8292 1822 8304
rect 1829 8292 1848 8304
rect 1879 8304 1929 8312
rect 1879 8296 1895 8304
rect 1902 8302 1929 8304
rect 1938 8302 2159 8312
rect 1902 8292 2159 8302
rect 2188 8304 2238 8312
rect 2188 8295 2204 8304
rect 1797 8284 1848 8292
rect 1895 8284 2159 8292
rect 2185 8292 2204 8295
rect 2211 8292 2238 8304
rect 2185 8284 2238 8292
rect 1813 8276 1814 8284
rect 1829 8276 1842 8284
rect 1813 8268 1829 8276
rect 1810 8261 1829 8264
rect 1810 8252 1832 8261
rect 1783 8242 1832 8252
rect 1783 8236 1813 8242
rect 1832 8237 1837 8242
rect 1755 8220 1829 8236
rect 1847 8228 1877 8284
rect 1912 8274 2120 8284
rect 2155 8280 2200 8284
rect 2203 8283 2204 8284
rect 2219 8283 2232 8284
rect 1938 8244 2127 8274
rect 1953 8241 2127 8244
rect 1946 8238 2127 8241
rect 1755 8218 1768 8220
rect 1783 8218 1817 8220
rect 1755 8202 1829 8218
rect 1856 8214 1869 8228
rect 1884 8214 1900 8230
rect 1946 8225 1957 8238
rect 1739 8180 1740 8196
rect 1755 8180 1768 8202
rect 1783 8180 1813 8202
rect 1856 8198 1918 8214
rect 1946 8207 1957 8223
rect 1962 8218 1972 8238
rect 1982 8218 1996 8238
rect 1999 8225 2008 8238
rect 2024 8225 2033 8238
rect 1962 8207 1996 8218
rect 1999 8207 2008 8223
rect 2024 8207 2033 8223
rect 2040 8218 2050 8238
rect 2060 8218 2074 8238
rect 2075 8225 2086 8238
rect 2040 8207 2074 8218
rect 2075 8207 2086 8223
rect 2132 8214 2148 8230
rect 2155 8228 2185 8280
rect 2219 8276 2220 8283
rect 2204 8268 2220 8276
rect 2191 8236 2204 8255
rect 2219 8236 2249 8252
rect 2191 8220 2265 8236
rect 2191 8218 2204 8220
rect 2219 8218 2253 8220
rect 1856 8196 1869 8198
rect 1884 8196 1918 8198
rect 1856 8180 1918 8196
rect 1962 8191 1978 8194
rect 2040 8191 2070 8202
rect 2118 8198 2164 8214
rect 2191 8202 2265 8218
rect 2118 8196 2152 8198
rect 2117 8180 2164 8196
rect 2191 8180 2204 8202
rect 2219 8180 2249 8202
rect 2276 8180 2277 8196
rect 2292 8180 2305 8340
rect 2335 8236 2348 8340
rect 2393 8318 2394 8328
rect 2409 8318 2422 8328
rect 2393 8314 2422 8318
rect 2427 8314 2457 8340
rect 2475 8326 2491 8328
rect 2563 8326 2616 8340
rect 2564 8324 2628 8326
rect 2671 8324 2686 8340
rect 2735 8337 2765 8340
rect 2735 8334 2771 8337
rect 2701 8326 2717 8328
rect 2475 8314 2490 8318
rect 2393 8312 2490 8314
rect 2518 8312 2686 8324
rect 2702 8314 2717 8318
rect 2735 8315 2774 8334
rect 2793 8328 2800 8329
rect 2799 8321 2800 8328
rect 2783 8318 2784 8321
rect 2799 8318 2812 8321
rect 2735 8314 2765 8315
rect 2774 8314 2780 8315
rect 2783 8314 2812 8318
rect 2702 8313 2812 8314
rect 2702 8312 2818 8313
rect 2377 8304 2428 8312
rect 2377 8292 2402 8304
rect 2409 8292 2428 8304
rect 2459 8304 2509 8312
rect 2459 8296 2475 8304
rect 2482 8302 2509 8304
rect 2518 8302 2739 8312
rect 2482 8292 2739 8302
rect 2768 8304 2818 8312
rect 2768 8295 2784 8304
rect 2377 8284 2428 8292
rect 2475 8284 2739 8292
rect 2765 8292 2784 8295
rect 2791 8292 2818 8304
rect 2765 8284 2818 8292
rect 2393 8276 2394 8284
rect 2409 8276 2422 8284
rect 2393 8268 2409 8276
rect 2390 8261 2409 8264
rect 2390 8252 2412 8261
rect 2363 8242 2412 8252
rect 2363 8236 2393 8242
rect 2412 8237 2417 8242
rect 2335 8220 2409 8236
rect 2427 8228 2457 8284
rect 2492 8274 2700 8284
rect 2735 8280 2780 8284
rect 2783 8283 2784 8284
rect 2799 8283 2812 8284
rect 2518 8244 2707 8274
rect 2533 8241 2707 8244
rect 2526 8238 2707 8241
rect 2335 8218 2348 8220
rect 2363 8218 2397 8220
rect 2335 8202 2409 8218
rect 2436 8214 2449 8228
rect 2464 8214 2480 8230
rect 2526 8225 2537 8238
rect 2319 8180 2320 8196
rect 2335 8180 2348 8202
rect 2363 8180 2393 8202
rect 2436 8198 2498 8214
rect 2526 8207 2537 8223
rect 2542 8218 2552 8238
rect 2562 8218 2576 8238
rect 2579 8225 2588 8238
rect 2604 8225 2613 8238
rect 2542 8207 2576 8218
rect 2579 8207 2588 8223
rect 2604 8207 2613 8223
rect 2620 8218 2630 8238
rect 2640 8218 2654 8238
rect 2655 8225 2666 8238
rect 2620 8207 2654 8218
rect 2655 8207 2666 8223
rect 2712 8214 2728 8230
rect 2735 8228 2765 8280
rect 2799 8276 2800 8283
rect 2784 8268 2800 8276
rect 2771 8236 2784 8255
rect 2799 8236 2829 8252
rect 2771 8220 2845 8236
rect 2771 8218 2784 8220
rect 2799 8218 2833 8220
rect 2436 8196 2449 8198
rect 2464 8196 2498 8198
rect 2436 8180 2498 8196
rect 2542 8191 2558 8194
rect 2620 8191 2650 8202
rect 2698 8198 2744 8214
rect 2771 8202 2845 8218
rect 2698 8196 2732 8198
rect 2697 8180 2744 8196
rect 2771 8180 2784 8202
rect 2799 8180 2829 8202
rect 2856 8180 2857 8196
rect 2872 8180 2885 8340
rect 2915 8236 2928 8340
rect 2973 8318 2974 8328
rect 2989 8318 3002 8328
rect 2973 8314 3002 8318
rect 3007 8314 3037 8340
rect 3055 8326 3071 8328
rect 3143 8326 3196 8340
rect 3144 8324 3208 8326
rect 3251 8324 3266 8340
rect 3315 8337 3345 8340
rect 3315 8334 3351 8337
rect 3281 8326 3297 8328
rect 3055 8314 3070 8318
rect 2973 8312 3070 8314
rect 3098 8312 3266 8324
rect 3282 8314 3297 8318
rect 3315 8315 3354 8334
rect 3373 8328 3380 8329
rect 3379 8321 3380 8328
rect 3363 8318 3364 8321
rect 3379 8318 3392 8321
rect 3315 8314 3345 8315
rect 3354 8314 3360 8315
rect 3363 8314 3392 8318
rect 3282 8313 3392 8314
rect 3282 8312 3398 8313
rect 2957 8304 3008 8312
rect 2957 8292 2982 8304
rect 2989 8292 3008 8304
rect 3039 8304 3089 8312
rect 3039 8296 3055 8304
rect 3062 8302 3089 8304
rect 3098 8302 3319 8312
rect 3062 8292 3319 8302
rect 3348 8304 3398 8312
rect 3348 8295 3364 8304
rect 2957 8284 3008 8292
rect 3055 8284 3319 8292
rect 3345 8292 3364 8295
rect 3371 8292 3398 8304
rect 3345 8284 3398 8292
rect 2973 8276 2974 8284
rect 2989 8276 3002 8284
rect 2973 8268 2989 8276
rect 2970 8261 2989 8264
rect 2970 8252 2992 8261
rect 2943 8242 2992 8252
rect 2943 8236 2973 8242
rect 2992 8237 2997 8242
rect 2915 8220 2989 8236
rect 3007 8228 3037 8284
rect 3072 8274 3280 8284
rect 3315 8280 3360 8284
rect 3363 8283 3364 8284
rect 3379 8283 3392 8284
rect 3098 8244 3287 8274
rect 3113 8241 3287 8244
rect 3106 8238 3287 8241
rect 2915 8218 2928 8220
rect 2943 8218 2977 8220
rect 2915 8202 2989 8218
rect 3016 8214 3029 8228
rect 3044 8214 3060 8230
rect 3106 8225 3117 8238
rect 2899 8180 2900 8196
rect 2915 8180 2928 8202
rect 2943 8180 2973 8202
rect 3016 8198 3078 8214
rect 3106 8207 3117 8223
rect 3122 8218 3132 8238
rect 3142 8218 3156 8238
rect 3159 8225 3168 8238
rect 3184 8225 3193 8238
rect 3122 8207 3156 8218
rect 3159 8207 3168 8223
rect 3184 8207 3193 8223
rect 3200 8218 3210 8238
rect 3220 8218 3234 8238
rect 3235 8225 3246 8238
rect 3200 8207 3234 8218
rect 3235 8207 3246 8223
rect 3292 8214 3308 8230
rect 3315 8228 3345 8280
rect 3379 8276 3380 8283
rect 3364 8268 3380 8276
rect 3351 8236 3364 8255
rect 3379 8236 3409 8252
rect 3351 8220 3425 8236
rect 3351 8218 3364 8220
rect 3379 8218 3413 8220
rect 3016 8196 3029 8198
rect 3044 8196 3078 8198
rect 3016 8180 3078 8196
rect 3122 8191 3138 8194
rect 3200 8191 3230 8202
rect 3278 8198 3324 8214
rect 3351 8202 3425 8218
rect 3278 8196 3312 8198
rect 3277 8180 3324 8196
rect 3351 8180 3364 8202
rect 3379 8180 3409 8202
rect 3436 8180 3437 8196
rect 3452 8180 3465 8340
rect 3495 8236 3508 8340
rect 3553 8318 3554 8328
rect 3569 8318 3582 8328
rect 3553 8314 3582 8318
rect 3587 8314 3617 8340
rect 3635 8326 3651 8328
rect 3723 8326 3776 8340
rect 3724 8324 3788 8326
rect 3831 8324 3846 8340
rect 3895 8337 3925 8340
rect 3895 8334 3931 8337
rect 3861 8326 3877 8328
rect 3635 8314 3650 8318
rect 3553 8312 3650 8314
rect 3678 8312 3846 8324
rect 3862 8314 3877 8318
rect 3895 8315 3934 8334
rect 3953 8328 3960 8329
rect 3959 8321 3960 8328
rect 3943 8318 3944 8321
rect 3959 8318 3972 8321
rect 3895 8314 3925 8315
rect 3934 8314 3940 8315
rect 3943 8314 3972 8318
rect 3862 8313 3972 8314
rect 3862 8312 3978 8313
rect 3537 8304 3588 8312
rect 3537 8292 3562 8304
rect 3569 8292 3588 8304
rect 3619 8304 3669 8312
rect 3619 8296 3635 8304
rect 3642 8302 3669 8304
rect 3678 8302 3899 8312
rect 3642 8292 3899 8302
rect 3928 8304 3978 8312
rect 3928 8295 3944 8304
rect 3537 8284 3588 8292
rect 3635 8284 3899 8292
rect 3925 8292 3944 8295
rect 3951 8292 3978 8304
rect 3925 8284 3978 8292
rect 3553 8276 3554 8284
rect 3569 8276 3582 8284
rect 3553 8268 3569 8276
rect 3550 8261 3569 8264
rect 3550 8252 3572 8261
rect 3523 8242 3572 8252
rect 3523 8236 3553 8242
rect 3572 8237 3577 8242
rect 3495 8220 3569 8236
rect 3587 8228 3617 8284
rect 3652 8274 3860 8284
rect 3895 8280 3940 8284
rect 3943 8283 3944 8284
rect 3959 8283 3972 8284
rect 3678 8244 3867 8274
rect 3693 8241 3867 8244
rect 3686 8238 3867 8241
rect 3495 8218 3508 8220
rect 3523 8218 3557 8220
rect 3495 8202 3569 8218
rect 3596 8214 3609 8228
rect 3624 8214 3640 8230
rect 3686 8225 3697 8238
rect 3479 8180 3480 8196
rect 3495 8180 3508 8202
rect 3523 8180 3553 8202
rect 3596 8198 3658 8214
rect 3686 8207 3697 8223
rect 3702 8218 3712 8238
rect 3722 8218 3736 8238
rect 3739 8225 3748 8238
rect 3764 8225 3773 8238
rect 3702 8207 3736 8218
rect 3739 8207 3748 8223
rect 3764 8207 3773 8223
rect 3780 8218 3790 8238
rect 3800 8218 3814 8238
rect 3815 8225 3826 8238
rect 3780 8207 3814 8218
rect 3815 8207 3826 8223
rect 3872 8214 3888 8230
rect 3895 8228 3925 8280
rect 3959 8276 3960 8283
rect 3944 8268 3960 8276
rect 3931 8236 3944 8255
rect 3959 8236 3989 8252
rect 3931 8220 4005 8236
rect 3931 8218 3944 8220
rect 3959 8218 3993 8220
rect 3596 8196 3609 8198
rect 3624 8196 3658 8198
rect 3596 8180 3658 8196
rect 3702 8191 3718 8194
rect 3780 8191 3810 8202
rect 3858 8198 3904 8214
rect 3931 8202 4005 8218
rect 3858 8196 3892 8198
rect 3857 8180 3904 8196
rect 3931 8180 3944 8202
rect 3959 8180 3989 8202
rect 4016 8180 4017 8196
rect 4032 8180 4045 8340
rect 4075 8236 4088 8340
rect 4133 8318 4134 8328
rect 4149 8318 4162 8328
rect 4133 8314 4162 8318
rect 4167 8314 4197 8340
rect 4215 8326 4231 8328
rect 4303 8326 4356 8340
rect 4304 8324 4368 8326
rect 4411 8324 4426 8340
rect 4475 8337 4505 8340
rect 4475 8334 4511 8337
rect 4441 8326 4457 8328
rect 4215 8314 4230 8318
rect 4133 8312 4230 8314
rect 4258 8312 4426 8324
rect 4442 8314 4457 8318
rect 4475 8315 4514 8334
rect 4533 8328 4540 8329
rect 4539 8321 4540 8328
rect 4523 8318 4524 8321
rect 4539 8318 4552 8321
rect 4475 8314 4505 8315
rect 4514 8314 4520 8315
rect 4523 8314 4552 8318
rect 4442 8313 4552 8314
rect 4442 8312 4558 8313
rect 4117 8304 4168 8312
rect 4117 8292 4142 8304
rect 4149 8292 4168 8304
rect 4199 8304 4249 8312
rect 4199 8296 4215 8304
rect 4222 8302 4249 8304
rect 4258 8302 4479 8312
rect 4222 8292 4479 8302
rect 4508 8304 4558 8312
rect 4508 8295 4524 8304
rect 4117 8284 4168 8292
rect 4215 8284 4479 8292
rect 4505 8292 4524 8295
rect 4531 8292 4558 8304
rect 4505 8284 4558 8292
rect 4133 8276 4134 8284
rect 4149 8276 4162 8284
rect 4133 8268 4149 8276
rect 4130 8261 4149 8264
rect 4130 8252 4152 8261
rect 4103 8242 4152 8252
rect 4103 8236 4133 8242
rect 4152 8237 4157 8242
rect 4075 8220 4149 8236
rect 4167 8228 4197 8284
rect 4232 8274 4440 8284
rect 4475 8280 4520 8284
rect 4523 8283 4524 8284
rect 4539 8283 4552 8284
rect 4258 8244 4447 8274
rect 4273 8241 4447 8244
rect 4266 8238 4447 8241
rect 4075 8218 4088 8220
rect 4103 8218 4137 8220
rect 4075 8202 4149 8218
rect 4176 8214 4189 8228
rect 4204 8214 4220 8230
rect 4266 8225 4277 8238
rect 4059 8180 4060 8196
rect 4075 8180 4088 8202
rect 4103 8180 4133 8202
rect 4176 8198 4238 8214
rect 4266 8207 4277 8223
rect 4282 8218 4292 8238
rect 4302 8218 4316 8238
rect 4319 8225 4328 8238
rect 4344 8225 4353 8238
rect 4282 8207 4316 8218
rect 4319 8207 4328 8223
rect 4344 8207 4353 8223
rect 4360 8218 4370 8238
rect 4380 8218 4394 8238
rect 4395 8225 4406 8238
rect 4360 8207 4394 8218
rect 4395 8207 4406 8223
rect 4452 8214 4468 8230
rect 4475 8228 4505 8280
rect 4539 8276 4540 8283
rect 4524 8268 4540 8276
rect 4511 8236 4524 8255
rect 4539 8236 4569 8252
rect 4511 8220 4585 8236
rect 4511 8218 4524 8220
rect 4539 8218 4573 8220
rect 4176 8196 4189 8198
rect 4204 8196 4238 8198
rect 4176 8180 4238 8196
rect 4282 8191 4298 8194
rect 4360 8191 4390 8202
rect 4438 8198 4484 8214
rect 4511 8202 4585 8218
rect 4438 8196 4472 8198
rect 4437 8180 4484 8196
rect 4511 8180 4524 8202
rect 4539 8180 4569 8202
rect 4596 8180 4597 8196
rect 4612 8180 4625 8340
rect -7 8172 34 8180
rect -7 8146 8 8172
rect 15 8146 34 8172
rect 98 8168 160 8180
rect 172 8168 247 8180
rect 305 8168 380 8180
rect 392 8168 423 8180
rect 429 8168 464 8180
rect 98 8166 260 8168
rect -7 8138 34 8146
rect 116 8142 129 8166
rect 144 8164 159 8166
rect -1 8128 0 8138
rect 15 8128 28 8138
rect 43 8128 73 8142
rect 116 8128 159 8142
rect 183 8139 190 8146
rect 193 8142 260 8166
rect 292 8166 464 8168
rect 262 8144 290 8148
rect 292 8144 372 8166
rect 393 8164 408 8166
rect 262 8142 372 8144
rect 193 8138 372 8142
rect 166 8128 196 8138
rect 198 8128 351 8138
rect 359 8128 389 8138
rect 393 8128 423 8142
rect 451 8128 464 8166
rect 536 8172 571 8180
rect 536 8146 537 8172
rect 544 8146 571 8172
rect 479 8128 509 8142
rect 536 8138 571 8146
rect 573 8172 614 8180
rect 573 8146 588 8172
rect 595 8146 614 8172
rect 678 8168 740 8180
rect 752 8168 827 8180
rect 885 8168 960 8180
rect 972 8168 1003 8180
rect 1009 8168 1044 8180
rect 678 8166 840 8168
rect 573 8138 614 8146
rect 696 8142 709 8166
rect 724 8164 739 8166
rect 536 8128 537 8138
rect 552 8128 565 8138
rect 579 8128 580 8138
rect 595 8128 608 8138
rect 623 8128 653 8142
rect 696 8128 739 8142
rect 763 8139 770 8146
rect 773 8142 840 8166
rect 872 8166 1044 8168
rect 842 8144 870 8148
rect 872 8144 952 8166
rect 973 8164 988 8166
rect 842 8142 952 8144
rect 773 8138 952 8142
rect 746 8128 776 8138
rect 778 8128 931 8138
rect 939 8128 969 8138
rect 973 8128 1003 8142
rect 1031 8128 1044 8166
rect 1116 8172 1151 8180
rect 1116 8146 1117 8172
rect 1124 8146 1151 8172
rect 1059 8128 1089 8142
rect 1116 8138 1151 8146
rect 1153 8172 1194 8180
rect 1153 8146 1168 8172
rect 1175 8146 1194 8172
rect 1258 8168 1320 8180
rect 1332 8168 1407 8180
rect 1465 8168 1540 8180
rect 1552 8168 1583 8180
rect 1589 8168 1624 8180
rect 1258 8166 1420 8168
rect 1153 8138 1194 8146
rect 1276 8142 1289 8166
rect 1304 8164 1319 8166
rect 1116 8128 1117 8138
rect 1132 8128 1145 8138
rect 1159 8128 1160 8138
rect 1175 8128 1188 8138
rect 1203 8128 1233 8142
rect 1276 8128 1319 8142
rect 1343 8139 1350 8146
rect 1353 8142 1420 8166
rect 1452 8166 1624 8168
rect 1422 8144 1450 8148
rect 1452 8144 1532 8166
rect 1553 8164 1568 8166
rect 1422 8142 1532 8144
rect 1353 8138 1532 8142
rect 1326 8128 1356 8138
rect 1358 8128 1511 8138
rect 1519 8128 1549 8138
rect 1553 8128 1583 8142
rect 1611 8128 1624 8166
rect 1696 8172 1731 8180
rect 1696 8146 1697 8172
rect 1704 8146 1731 8172
rect 1639 8128 1669 8142
rect 1696 8138 1731 8146
rect 1733 8172 1774 8180
rect 1733 8146 1748 8172
rect 1755 8146 1774 8172
rect 1838 8168 1900 8180
rect 1912 8168 1987 8180
rect 2045 8168 2120 8180
rect 2132 8168 2163 8180
rect 2169 8168 2204 8180
rect 1838 8166 2000 8168
rect 1733 8138 1774 8146
rect 1856 8142 1869 8166
rect 1884 8164 1899 8166
rect 1696 8128 1697 8138
rect 1712 8128 1725 8138
rect 1739 8128 1740 8138
rect 1755 8128 1768 8138
rect 1783 8128 1813 8142
rect 1856 8128 1899 8142
rect 1923 8139 1930 8146
rect 1933 8142 2000 8166
rect 2032 8166 2204 8168
rect 2002 8144 2030 8148
rect 2032 8144 2112 8166
rect 2133 8164 2148 8166
rect 2002 8142 2112 8144
rect 1933 8138 2112 8142
rect 1906 8128 1936 8138
rect 1938 8128 2091 8138
rect 2099 8128 2129 8138
rect 2133 8128 2163 8142
rect 2191 8128 2204 8166
rect 2276 8172 2311 8180
rect 2276 8146 2277 8172
rect 2284 8146 2311 8172
rect 2219 8128 2249 8142
rect 2276 8138 2311 8146
rect 2313 8172 2354 8180
rect 2313 8146 2328 8172
rect 2335 8146 2354 8172
rect 2418 8168 2480 8180
rect 2492 8168 2567 8180
rect 2625 8168 2700 8180
rect 2712 8168 2743 8180
rect 2749 8168 2784 8180
rect 2418 8166 2580 8168
rect 2313 8138 2354 8146
rect 2436 8142 2449 8166
rect 2464 8164 2479 8166
rect 2276 8128 2277 8138
rect 2292 8128 2305 8138
rect 2319 8128 2320 8138
rect 2335 8128 2348 8138
rect 2363 8128 2393 8142
rect 2436 8128 2479 8142
rect 2503 8139 2510 8146
rect 2513 8142 2580 8166
rect 2612 8166 2784 8168
rect 2582 8144 2610 8148
rect 2612 8144 2692 8166
rect 2713 8164 2728 8166
rect 2582 8142 2692 8144
rect 2513 8138 2692 8142
rect 2486 8128 2516 8138
rect 2518 8128 2671 8138
rect 2679 8128 2709 8138
rect 2713 8128 2743 8142
rect 2771 8128 2784 8166
rect 2856 8172 2891 8180
rect 2856 8146 2857 8172
rect 2864 8146 2891 8172
rect 2799 8128 2829 8142
rect 2856 8138 2891 8146
rect 2893 8172 2934 8180
rect 2893 8146 2908 8172
rect 2915 8146 2934 8172
rect 2998 8168 3060 8180
rect 3072 8168 3147 8180
rect 3205 8168 3280 8180
rect 3292 8168 3323 8180
rect 3329 8168 3364 8180
rect 2998 8166 3160 8168
rect 2893 8138 2934 8146
rect 3016 8142 3029 8166
rect 3044 8164 3059 8166
rect 2856 8128 2857 8138
rect 2872 8128 2885 8138
rect 2899 8128 2900 8138
rect 2915 8128 2928 8138
rect 2943 8128 2973 8142
rect 3016 8128 3059 8142
rect 3083 8139 3090 8146
rect 3093 8142 3160 8166
rect 3192 8166 3364 8168
rect 3162 8144 3190 8148
rect 3192 8144 3272 8166
rect 3293 8164 3308 8166
rect 3162 8142 3272 8144
rect 3093 8138 3272 8142
rect 3066 8128 3096 8138
rect 3098 8128 3251 8138
rect 3259 8128 3289 8138
rect 3293 8128 3323 8142
rect 3351 8128 3364 8166
rect 3436 8172 3471 8180
rect 3436 8146 3437 8172
rect 3444 8146 3471 8172
rect 3379 8128 3409 8142
rect 3436 8138 3471 8146
rect 3473 8172 3514 8180
rect 3473 8146 3488 8172
rect 3495 8146 3514 8172
rect 3578 8168 3640 8180
rect 3652 8168 3727 8180
rect 3785 8168 3860 8180
rect 3872 8168 3903 8180
rect 3909 8168 3944 8180
rect 3578 8166 3740 8168
rect 3473 8138 3514 8146
rect 3596 8142 3609 8166
rect 3624 8164 3639 8166
rect 3436 8128 3437 8138
rect 3452 8128 3465 8138
rect 3479 8128 3480 8138
rect 3495 8128 3508 8138
rect 3523 8128 3553 8142
rect 3596 8128 3639 8142
rect 3663 8139 3670 8146
rect 3673 8142 3740 8166
rect 3772 8166 3944 8168
rect 3742 8144 3770 8148
rect 3772 8144 3852 8166
rect 3873 8164 3888 8166
rect 3742 8142 3852 8144
rect 3673 8138 3852 8142
rect 3646 8128 3676 8138
rect 3678 8128 3831 8138
rect 3839 8128 3869 8138
rect 3873 8128 3903 8142
rect 3931 8128 3944 8166
rect 4016 8172 4051 8180
rect 4016 8146 4017 8172
rect 4024 8146 4051 8172
rect 3959 8128 3989 8142
rect 4016 8138 4051 8146
rect 4053 8172 4094 8180
rect 4053 8146 4068 8172
rect 4075 8146 4094 8172
rect 4158 8168 4220 8180
rect 4232 8168 4307 8180
rect 4365 8168 4440 8180
rect 4452 8168 4483 8180
rect 4489 8168 4524 8180
rect 4158 8166 4320 8168
rect 4053 8138 4094 8146
rect 4176 8142 4189 8166
rect 4204 8164 4219 8166
rect 4016 8128 4017 8138
rect 4032 8128 4045 8138
rect 4059 8128 4060 8138
rect 4075 8128 4088 8138
rect 4103 8128 4133 8142
rect 4176 8128 4219 8142
rect 4243 8139 4250 8146
rect 4253 8142 4320 8166
rect 4352 8166 4524 8168
rect 4322 8144 4350 8148
rect 4352 8144 4432 8166
rect 4453 8164 4468 8166
rect 4322 8142 4432 8144
rect 4253 8138 4432 8142
rect 4226 8128 4256 8138
rect 4258 8128 4411 8138
rect 4419 8128 4449 8138
rect 4453 8128 4483 8142
rect 4511 8128 4524 8166
rect 4596 8172 4631 8180
rect 4596 8146 4597 8172
rect 4604 8146 4631 8172
rect 4539 8128 4569 8142
rect 4596 8138 4631 8146
rect 4596 8128 4597 8138
rect 4612 8128 4625 8138
rect -1 8122 4625 8128
rect 0 8114 4625 8122
rect 15 8084 28 8114
rect 43 8096 73 8114
rect 116 8100 130 8114
rect 166 8100 386 8114
rect 117 8098 130 8100
rect 83 8086 98 8098
rect 80 8084 102 8086
rect 107 8084 137 8098
rect 198 8096 351 8100
rect 180 8084 372 8096
rect 415 8084 445 8098
rect 451 8084 464 8114
rect 479 8096 509 8114
rect 552 8084 565 8114
rect 595 8084 608 8114
rect 623 8096 653 8114
rect 696 8100 710 8114
rect 746 8100 966 8114
rect 697 8098 710 8100
rect 663 8086 678 8098
rect 660 8084 682 8086
rect 687 8084 717 8098
rect 778 8096 931 8100
rect 760 8084 952 8096
rect 995 8084 1025 8098
rect 1031 8084 1044 8114
rect 1059 8096 1089 8114
rect 1132 8084 1145 8114
rect 1175 8084 1188 8114
rect 1203 8096 1233 8114
rect 1276 8100 1290 8114
rect 1326 8100 1546 8114
rect 1277 8098 1290 8100
rect 1243 8086 1258 8098
rect 1240 8084 1262 8086
rect 1267 8084 1297 8098
rect 1358 8096 1511 8100
rect 1340 8084 1532 8096
rect 1575 8084 1605 8098
rect 1611 8084 1624 8114
rect 1639 8096 1669 8114
rect 1712 8084 1725 8114
rect 1755 8084 1768 8114
rect 1783 8096 1813 8114
rect 1856 8100 1870 8114
rect 1906 8100 2126 8114
rect 1857 8098 1870 8100
rect 1823 8086 1838 8098
rect 1820 8084 1842 8086
rect 1847 8084 1877 8098
rect 1938 8096 2091 8100
rect 1920 8084 2112 8096
rect 2155 8084 2185 8098
rect 2191 8084 2204 8114
rect 2219 8096 2249 8114
rect 2292 8084 2305 8114
rect 2335 8084 2348 8114
rect 2363 8096 2393 8114
rect 2436 8100 2450 8114
rect 2486 8100 2706 8114
rect 2437 8098 2450 8100
rect 2403 8086 2418 8098
rect 2400 8084 2422 8086
rect 2427 8084 2457 8098
rect 2518 8096 2671 8100
rect 2500 8084 2692 8096
rect 2735 8084 2765 8098
rect 2771 8084 2784 8114
rect 2799 8096 2829 8114
rect 2872 8084 2885 8114
rect 2915 8084 2928 8114
rect 2943 8096 2973 8114
rect 3016 8100 3030 8114
rect 3066 8100 3286 8114
rect 3017 8098 3030 8100
rect 2983 8086 2998 8098
rect 2980 8084 3002 8086
rect 3007 8084 3037 8098
rect 3098 8096 3251 8100
rect 3080 8084 3272 8096
rect 3315 8084 3345 8098
rect 3351 8084 3364 8114
rect 3379 8096 3409 8114
rect 3452 8084 3465 8114
rect 3495 8084 3508 8114
rect 3523 8096 3553 8114
rect 3596 8100 3610 8114
rect 3646 8100 3866 8114
rect 3597 8098 3610 8100
rect 3563 8086 3578 8098
rect 3560 8084 3582 8086
rect 3587 8084 3617 8098
rect 3678 8096 3831 8100
rect 3660 8084 3852 8096
rect 3895 8084 3925 8098
rect 3931 8084 3944 8114
rect 3959 8096 3989 8114
rect 4032 8084 4045 8114
rect 4075 8084 4088 8114
rect 4103 8096 4133 8114
rect 4176 8100 4190 8114
rect 4226 8100 4446 8114
rect 4177 8098 4190 8100
rect 4143 8086 4158 8098
rect 4140 8084 4162 8086
rect 4167 8084 4197 8098
rect 4258 8096 4411 8100
rect 4240 8084 4432 8096
rect 4475 8084 4505 8098
rect 4511 8084 4524 8114
rect 4539 8096 4569 8114
rect 4612 8084 4625 8114
rect 0 8070 4625 8084
rect 15 7966 28 8070
rect 73 8048 74 8058
rect 89 8048 102 8058
rect 73 8044 102 8048
rect 107 8044 137 8070
rect 155 8056 171 8058
rect 243 8056 296 8070
rect 244 8054 308 8056
rect 351 8054 366 8070
rect 415 8067 445 8070
rect 415 8064 451 8067
rect 381 8056 397 8058
rect 155 8044 170 8048
rect 73 8042 170 8044
rect 198 8042 366 8054
rect 382 8044 397 8048
rect 415 8045 454 8064
rect 473 8058 480 8059
rect 479 8051 480 8058
rect 463 8048 464 8051
rect 479 8048 492 8051
rect 415 8044 445 8045
rect 454 8044 460 8045
rect 463 8044 492 8048
rect 382 8043 492 8044
rect 382 8042 498 8043
rect 57 8034 108 8042
rect 57 8022 82 8034
rect 89 8022 108 8034
rect 139 8034 189 8042
rect 139 8026 155 8034
rect 162 8032 189 8034
rect 198 8032 419 8042
rect 162 8022 419 8032
rect 448 8034 498 8042
rect 448 8025 464 8034
rect 57 8014 108 8022
rect 155 8014 419 8022
rect 445 8022 464 8025
rect 471 8022 498 8034
rect 445 8014 498 8022
rect 73 8006 74 8014
rect 89 8006 102 8014
rect 73 7998 89 8006
rect 70 7991 89 7994
rect 70 7982 92 7991
rect 43 7972 92 7982
rect 43 7966 73 7972
rect 92 7967 97 7972
rect 15 7950 89 7966
rect 107 7958 137 8014
rect 172 8004 380 8014
rect 415 8010 460 8014
rect 463 8013 464 8014
rect 479 8013 492 8014
rect 198 7974 387 8004
rect 213 7971 387 7974
rect 206 7968 387 7971
rect 15 7948 28 7950
rect 43 7948 77 7950
rect 15 7932 89 7948
rect 116 7944 129 7958
rect 144 7944 160 7960
rect 206 7955 217 7968
rect -1 7910 0 7926
rect 15 7910 28 7932
rect 43 7910 73 7932
rect 116 7928 178 7944
rect 206 7937 217 7953
rect 222 7948 232 7968
rect 242 7948 256 7968
rect 259 7955 268 7968
rect 284 7955 293 7968
rect 222 7937 256 7948
rect 259 7937 268 7953
rect 284 7937 293 7953
rect 300 7948 310 7968
rect 320 7948 334 7968
rect 335 7955 346 7968
rect 300 7937 334 7948
rect 335 7937 346 7953
rect 392 7944 408 7960
rect 415 7958 445 8010
rect 479 8006 480 8013
rect 464 7998 480 8006
rect 451 7966 464 7985
rect 479 7966 509 7982
rect 451 7950 525 7966
rect 451 7948 464 7950
rect 479 7948 513 7950
rect 116 7926 129 7928
rect 144 7926 178 7928
rect 116 7910 178 7926
rect 222 7921 238 7924
rect 300 7921 330 7932
rect 378 7928 424 7944
rect 451 7932 525 7948
rect 378 7926 412 7928
rect 377 7910 424 7926
rect 451 7910 464 7932
rect 479 7910 509 7932
rect 536 7910 537 7926
rect 552 7910 565 8070
rect 595 7966 608 8070
rect 653 8048 654 8058
rect 669 8048 682 8058
rect 653 8044 682 8048
rect 687 8044 717 8070
rect 735 8056 751 8058
rect 823 8056 876 8070
rect 824 8054 888 8056
rect 931 8054 946 8070
rect 995 8067 1025 8070
rect 995 8064 1031 8067
rect 961 8056 977 8058
rect 735 8044 750 8048
rect 653 8042 750 8044
rect 778 8042 946 8054
rect 962 8044 977 8048
rect 995 8045 1034 8064
rect 1053 8058 1060 8059
rect 1059 8051 1060 8058
rect 1043 8048 1044 8051
rect 1059 8048 1072 8051
rect 995 8044 1025 8045
rect 1034 8044 1040 8045
rect 1043 8044 1072 8048
rect 962 8043 1072 8044
rect 962 8042 1078 8043
rect 637 8034 688 8042
rect 637 8022 662 8034
rect 669 8022 688 8034
rect 719 8034 769 8042
rect 719 8026 735 8034
rect 742 8032 769 8034
rect 778 8032 999 8042
rect 742 8022 999 8032
rect 1028 8034 1078 8042
rect 1028 8025 1044 8034
rect 637 8014 688 8022
rect 735 8014 999 8022
rect 1025 8022 1044 8025
rect 1051 8022 1078 8034
rect 1025 8014 1078 8022
rect 653 8006 654 8014
rect 669 8006 682 8014
rect 653 7998 669 8006
rect 650 7991 669 7994
rect 650 7982 672 7991
rect 623 7972 672 7982
rect 623 7966 653 7972
rect 672 7967 677 7972
rect 595 7950 669 7966
rect 687 7958 717 8014
rect 752 8004 960 8014
rect 995 8010 1040 8014
rect 1043 8013 1044 8014
rect 1059 8013 1072 8014
rect 778 7974 967 8004
rect 793 7971 967 7974
rect 786 7968 967 7971
rect 595 7948 608 7950
rect 623 7948 657 7950
rect 595 7932 669 7948
rect 696 7944 709 7958
rect 724 7944 740 7960
rect 786 7955 797 7968
rect 579 7910 580 7926
rect 595 7910 608 7932
rect 623 7910 653 7932
rect 696 7928 758 7944
rect 786 7937 797 7953
rect 802 7948 812 7968
rect 822 7948 836 7968
rect 839 7955 848 7968
rect 864 7955 873 7968
rect 802 7937 836 7948
rect 839 7937 848 7953
rect 864 7937 873 7953
rect 880 7948 890 7968
rect 900 7948 914 7968
rect 915 7955 926 7968
rect 880 7937 914 7948
rect 915 7937 926 7953
rect 972 7944 988 7960
rect 995 7958 1025 8010
rect 1059 8006 1060 8013
rect 1044 7998 1060 8006
rect 1031 7966 1044 7985
rect 1059 7966 1089 7982
rect 1031 7950 1105 7966
rect 1031 7948 1044 7950
rect 1059 7948 1093 7950
rect 696 7926 709 7928
rect 724 7926 758 7928
rect 696 7910 758 7926
rect 802 7921 818 7924
rect 880 7921 910 7932
rect 958 7928 1004 7944
rect 1031 7932 1105 7948
rect 958 7926 992 7928
rect 957 7910 1004 7926
rect 1031 7910 1044 7932
rect 1059 7910 1089 7932
rect 1116 7910 1117 7926
rect 1132 7910 1145 8070
rect 1175 7966 1188 8070
rect 1233 8048 1234 8058
rect 1249 8048 1262 8058
rect 1233 8044 1262 8048
rect 1267 8044 1297 8070
rect 1315 8056 1331 8058
rect 1403 8056 1456 8070
rect 1404 8054 1468 8056
rect 1511 8054 1526 8070
rect 1575 8067 1605 8070
rect 1575 8064 1611 8067
rect 1541 8056 1557 8058
rect 1315 8044 1330 8048
rect 1233 8042 1330 8044
rect 1358 8042 1526 8054
rect 1542 8044 1557 8048
rect 1575 8045 1614 8064
rect 1633 8058 1640 8059
rect 1639 8051 1640 8058
rect 1623 8048 1624 8051
rect 1639 8048 1652 8051
rect 1575 8044 1605 8045
rect 1614 8044 1620 8045
rect 1623 8044 1652 8048
rect 1542 8043 1652 8044
rect 1542 8042 1658 8043
rect 1217 8034 1268 8042
rect 1217 8022 1242 8034
rect 1249 8022 1268 8034
rect 1299 8034 1349 8042
rect 1299 8026 1315 8034
rect 1322 8032 1349 8034
rect 1358 8032 1579 8042
rect 1322 8022 1579 8032
rect 1608 8034 1658 8042
rect 1608 8025 1624 8034
rect 1217 8014 1268 8022
rect 1315 8014 1579 8022
rect 1605 8022 1624 8025
rect 1631 8022 1658 8034
rect 1605 8014 1658 8022
rect 1233 8006 1234 8014
rect 1249 8006 1262 8014
rect 1233 7998 1249 8006
rect 1230 7991 1249 7994
rect 1230 7982 1252 7991
rect 1203 7972 1252 7982
rect 1203 7966 1233 7972
rect 1252 7967 1257 7972
rect 1175 7950 1249 7966
rect 1267 7958 1297 8014
rect 1332 8004 1540 8014
rect 1575 8010 1620 8014
rect 1623 8013 1624 8014
rect 1639 8013 1652 8014
rect 1358 7974 1547 8004
rect 1373 7971 1547 7974
rect 1366 7968 1547 7971
rect 1175 7948 1188 7950
rect 1203 7948 1237 7950
rect 1175 7932 1249 7948
rect 1276 7944 1289 7958
rect 1304 7944 1320 7960
rect 1366 7955 1377 7968
rect 1159 7910 1160 7926
rect 1175 7910 1188 7932
rect 1203 7910 1233 7932
rect 1276 7928 1338 7944
rect 1366 7937 1377 7953
rect 1382 7948 1392 7968
rect 1402 7948 1416 7968
rect 1419 7955 1428 7968
rect 1444 7955 1453 7968
rect 1382 7937 1416 7948
rect 1419 7937 1428 7953
rect 1444 7937 1453 7953
rect 1460 7948 1470 7968
rect 1480 7948 1494 7968
rect 1495 7955 1506 7968
rect 1460 7937 1494 7948
rect 1495 7937 1506 7953
rect 1552 7944 1568 7960
rect 1575 7958 1605 8010
rect 1639 8006 1640 8013
rect 1624 7998 1640 8006
rect 1611 7966 1624 7985
rect 1639 7966 1669 7982
rect 1611 7950 1685 7966
rect 1611 7948 1624 7950
rect 1639 7948 1673 7950
rect 1276 7926 1289 7928
rect 1304 7926 1338 7928
rect 1276 7910 1338 7926
rect 1382 7921 1398 7924
rect 1460 7921 1490 7932
rect 1538 7928 1584 7944
rect 1611 7932 1685 7948
rect 1538 7926 1572 7928
rect 1537 7910 1584 7926
rect 1611 7910 1624 7932
rect 1639 7910 1669 7932
rect 1696 7910 1697 7926
rect 1712 7910 1725 8070
rect 1755 7966 1768 8070
rect 1813 8048 1814 8058
rect 1829 8048 1842 8058
rect 1813 8044 1842 8048
rect 1847 8044 1877 8070
rect 1895 8056 1911 8058
rect 1983 8056 2036 8070
rect 1984 8054 2048 8056
rect 2091 8054 2106 8070
rect 2155 8067 2185 8070
rect 2155 8064 2191 8067
rect 2121 8056 2137 8058
rect 1895 8044 1910 8048
rect 1813 8042 1910 8044
rect 1938 8042 2106 8054
rect 2122 8044 2137 8048
rect 2155 8045 2194 8064
rect 2213 8058 2220 8059
rect 2219 8051 2220 8058
rect 2203 8048 2204 8051
rect 2219 8048 2232 8051
rect 2155 8044 2185 8045
rect 2194 8044 2200 8045
rect 2203 8044 2232 8048
rect 2122 8043 2232 8044
rect 2122 8042 2238 8043
rect 1797 8034 1848 8042
rect 1797 8022 1822 8034
rect 1829 8022 1848 8034
rect 1879 8034 1929 8042
rect 1879 8026 1895 8034
rect 1902 8032 1929 8034
rect 1938 8032 2159 8042
rect 1902 8022 2159 8032
rect 2188 8034 2238 8042
rect 2188 8025 2204 8034
rect 1797 8014 1848 8022
rect 1895 8014 2159 8022
rect 2185 8022 2204 8025
rect 2211 8022 2238 8034
rect 2185 8014 2238 8022
rect 1813 8006 1814 8014
rect 1829 8006 1842 8014
rect 1813 7998 1829 8006
rect 1810 7991 1829 7994
rect 1810 7982 1832 7991
rect 1783 7972 1832 7982
rect 1783 7966 1813 7972
rect 1832 7967 1837 7972
rect 1755 7950 1829 7966
rect 1847 7958 1877 8014
rect 1912 8004 2120 8014
rect 2155 8010 2200 8014
rect 2203 8013 2204 8014
rect 2219 8013 2232 8014
rect 1938 7974 2127 8004
rect 1953 7971 2127 7974
rect 1946 7968 2127 7971
rect 1755 7948 1768 7950
rect 1783 7948 1817 7950
rect 1755 7932 1829 7948
rect 1856 7944 1869 7958
rect 1884 7944 1900 7960
rect 1946 7955 1957 7968
rect 1739 7910 1740 7926
rect 1755 7910 1768 7932
rect 1783 7910 1813 7932
rect 1856 7928 1918 7944
rect 1946 7937 1957 7953
rect 1962 7948 1972 7968
rect 1982 7948 1996 7968
rect 1999 7955 2008 7968
rect 2024 7955 2033 7968
rect 1962 7937 1996 7948
rect 1999 7937 2008 7953
rect 2024 7937 2033 7953
rect 2040 7948 2050 7968
rect 2060 7948 2074 7968
rect 2075 7955 2086 7968
rect 2040 7937 2074 7948
rect 2075 7937 2086 7953
rect 2132 7944 2148 7960
rect 2155 7958 2185 8010
rect 2219 8006 2220 8013
rect 2204 7998 2220 8006
rect 2191 7966 2204 7985
rect 2219 7966 2249 7982
rect 2191 7950 2265 7966
rect 2191 7948 2204 7950
rect 2219 7948 2253 7950
rect 1856 7926 1869 7928
rect 1884 7926 1918 7928
rect 1856 7910 1918 7926
rect 1962 7921 1978 7924
rect 2040 7921 2070 7932
rect 2118 7928 2164 7944
rect 2191 7932 2265 7948
rect 2118 7926 2152 7928
rect 2117 7910 2164 7926
rect 2191 7910 2204 7932
rect 2219 7910 2249 7932
rect 2276 7910 2277 7926
rect 2292 7910 2305 8070
rect 2335 7966 2348 8070
rect 2393 8048 2394 8058
rect 2409 8048 2422 8058
rect 2393 8044 2422 8048
rect 2427 8044 2457 8070
rect 2475 8056 2491 8058
rect 2563 8056 2616 8070
rect 2564 8054 2628 8056
rect 2671 8054 2686 8070
rect 2735 8067 2765 8070
rect 2735 8064 2771 8067
rect 2701 8056 2717 8058
rect 2475 8044 2490 8048
rect 2393 8042 2490 8044
rect 2518 8042 2686 8054
rect 2702 8044 2717 8048
rect 2735 8045 2774 8064
rect 2793 8058 2800 8059
rect 2799 8051 2800 8058
rect 2783 8048 2784 8051
rect 2799 8048 2812 8051
rect 2735 8044 2765 8045
rect 2774 8044 2780 8045
rect 2783 8044 2812 8048
rect 2702 8043 2812 8044
rect 2702 8042 2818 8043
rect 2377 8034 2428 8042
rect 2377 8022 2402 8034
rect 2409 8022 2428 8034
rect 2459 8034 2509 8042
rect 2459 8026 2475 8034
rect 2482 8032 2509 8034
rect 2518 8032 2739 8042
rect 2482 8022 2739 8032
rect 2768 8034 2818 8042
rect 2768 8025 2784 8034
rect 2377 8014 2428 8022
rect 2475 8014 2739 8022
rect 2765 8022 2784 8025
rect 2791 8022 2818 8034
rect 2765 8014 2818 8022
rect 2393 8006 2394 8014
rect 2409 8006 2422 8014
rect 2393 7998 2409 8006
rect 2390 7991 2409 7994
rect 2390 7982 2412 7991
rect 2363 7972 2412 7982
rect 2363 7966 2393 7972
rect 2412 7967 2417 7972
rect 2335 7950 2409 7966
rect 2427 7958 2457 8014
rect 2492 8004 2700 8014
rect 2735 8010 2780 8014
rect 2783 8013 2784 8014
rect 2799 8013 2812 8014
rect 2518 7974 2707 8004
rect 2533 7971 2707 7974
rect 2526 7968 2707 7971
rect 2335 7948 2348 7950
rect 2363 7948 2397 7950
rect 2335 7932 2409 7948
rect 2436 7944 2449 7958
rect 2464 7944 2480 7960
rect 2526 7955 2537 7968
rect 2319 7910 2320 7926
rect 2335 7910 2348 7932
rect 2363 7910 2393 7932
rect 2436 7928 2498 7944
rect 2526 7937 2537 7953
rect 2542 7948 2552 7968
rect 2562 7948 2576 7968
rect 2579 7955 2588 7968
rect 2604 7955 2613 7968
rect 2542 7937 2576 7948
rect 2579 7937 2588 7953
rect 2604 7937 2613 7953
rect 2620 7948 2630 7968
rect 2640 7948 2654 7968
rect 2655 7955 2666 7968
rect 2620 7937 2654 7948
rect 2655 7937 2666 7953
rect 2712 7944 2728 7960
rect 2735 7958 2765 8010
rect 2799 8006 2800 8013
rect 2784 7998 2800 8006
rect 2771 7966 2784 7985
rect 2799 7966 2829 7982
rect 2771 7950 2845 7966
rect 2771 7948 2784 7950
rect 2799 7948 2833 7950
rect 2436 7926 2449 7928
rect 2464 7926 2498 7928
rect 2436 7910 2498 7926
rect 2542 7921 2558 7924
rect 2620 7921 2650 7932
rect 2698 7928 2744 7944
rect 2771 7932 2845 7948
rect 2698 7926 2732 7928
rect 2697 7910 2744 7926
rect 2771 7910 2784 7932
rect 2799 7910 2829 7932
rect 2856 7910 2857 7926
rect 2872 7910 2885 8070
rect 2915 7966 2928 8070
rect 2973 8048 2974 8058
rect 2989 8048 3002 8058
rect 2973 8044 3002 8048
rect 3007 8044 3037 8070
rect 3055 8056 3071 8058
rect 3143 8056 3196 8070
rect 3144 8054 3208 8056
rect 3251 8054 3266 8070
rect 3315 8067 3345 8070
rect 3315 8064 3351 8067
rect 3281 8056 3297 8058
rect 3055 8044 3070 8048
rect 2973 8042 3070 8044
rect 3098 8042 3266 8054
rect 3282 8044 3297 8048
rect 3315 8045 3354 8064
rect 3373 8058 3380 8059
rect 3379 8051 3380 8058
rect 3363 8048 3364 8051
rect 3379 8048 3392 8051
rect 3315 8044 3345 8045
rect 3354 8044 3360 8045
rect 3363 8044 3392 8048
rect 3282 8043 3392 8044
rect 3282 8042 3398 8043
rect 2957 8034 3008 8042
rect 2957 8022 2982 8034
rect 2989 8022 3008 8034
rect 3039 8034 3089 8042
rect 3039 8026 3055 8034
rect 3062 8032 3089 8034
rect 3098 8032 3319 8042
rect 3062 8022 3319 8032
rect 3348 8034 3398 8042
rect 3348 8025 3364 8034
rect 2957 8014 3008 8022
rect 3055 8014 3319 8022
rect 3345 8022 3364 8025
rect 3371 8022 3398 8034
rect 3345 8014 3398 8022
rect 2973 8006 2974 8014
rect 2989 8006 3002 8014
rect 2973 7998 2989 8006
rect 2970 7991 2989 7994
rect 2970 7982 2992 7991
rect 2943 7972 2992 7982
rect 2943 7966 2973 7972
rect 2992 7967 2997 7972
rect 2915 7950 2989 7966
rect 3007 7958 3037 8014
rect 3072 8004 3280 8014
rect 3315 8010 3360 8014
rect 3363 8013 3364 8014
rect 3379 8013 3392 8014
rect 3098 7974 3287 8004
rect 3113 7971 3287 7974
rect 3106 7968 3287 7971
rect 2915 7948 2928 7950
rect 2943 7948 2977 7950
rect 2915 7932 2989 7948
rect 3016 7944 3029 7958
rect 3044 7944 3060 7960
rect 3106 7955 3117 7968
rect 2899 7910 2900 7926
rect 2915 7910 2928 7932
rect 2943 7910 2973 7932
rect 3016 7928 3078 7944
rect 3106 7937 3117 7953
rect 3122 7948 3132 7968
rect 3142 7948 3156 7968
rect 3159 7955 3168 7968
rect 3184 7955 3193 7968
rect 3122 7937 3156 7948
rect 3159 7937 3168 7953
rect 3184 7937 3193 7953
rect 3200 7948 3210 7968
rect 3220 7948 3234 7968
rect 3235 7955 3246 7968
rect 3200 7937 3234 7948
rect 3235 7937 3246 7953
rect 3292 7944 3308 7960
rect 3315 7958 3345 8010
rect 3379 8006 3380 8013
rect 3364 7998 3380 8006
rect 3351 7966 3364 7985
rect 3379 7966 3409 7982
rect 3351 7950 3425 7966
rect 3351 7948 3364 7950
rect 3379 7948 3413 7950
rect 3016 7926 3029 7928
rect 3044 7926 3078 7928
rect 3016 7910 3078 7926
rect 3122 7921 3138 7924
rect 3200 7921 3230 7932
rect 3278 7928 3324 7944
rect 3351 7932 3425 7948
rect 3278 7926 3312 7928
rect 3277 7910 3324 7926
rect 3351 7910 3364 7932
rect 3379 7910 3409 7932
rect 3436 7910 3437 7926
rect 3452 7910 3465 8070
rect 3495 7966 3508 8070
rect 3553 8048 3554 8058
rect 3569 8048 3582 8058
rect 3553 8044 3582 8048
rect 3587 8044 3617 8070
rect 3635 8056 3651 8058
rect 3723 8056 3776 8070
rect 3724 8054 3788 8056
rect 3831 8054 3846 8070
rect 3895 8067 3925 8070
rect 3895 8064 3931 8067
rect 3861 8056 3877 8058
rect 3635 8044 3650 8048
rect 3553 8042 3650 8044
rect 3678 8042 3846 8054
rect 3862 8044 3877 8048
rect 3895 8045 3934 8064
rect 3953 8058 3960 8059
rect 3959 8051 3960 8058
rect 3943 8048 3944 8051
rect 3959 8048 3972 8051
rect 3895 8044 3925 8045
rect 3934 8044 3940 8045
rect 3943 8044 3972 8048
rect 3862 8043 3972 8044
rect 3862 8042 3978 8043
rect 3537 8034 3588 8042
rect 3537 8022 3562 8034
rect 3569 8022 3588 8034
rect 3619 8034 3669 8042
rect 3619 8026 3635 8034
rect 3642 8032 3669 8034
rect 3678 8032 3899 8042
rect 3642 8022 3899 8032
rect 3928 8034 3978 8042
rect 3928 8025 3944 8034
rect 3537 8014 3588 8022
rect 3635 8014 3899 8022
rect 3925 8022 3944 8025
rect 3951 8022 3978 8034
rect 3925 8014 3978 8022
rect 3553 8006 3554 8014
rect 3569 8006 3582 8014
rect 3553 7998 3569 8006
rect 3550 7991 3569 7994
rect 3550 7982 3572 7991
rect 3523 7972 3572 7982
rect 3523 7966 3553 7972
rect 3572 7967 3577 7972
rect 3495 7950 3569 7966
rect 3587 7958 3617 8014
rect 3652 8004 3860 8014
rect 3895 8010 3940 8014
rect 3943 8013 3944 8014
rect 3959 8013 3972 8014
rect 3678 7974 3867 8004
rect 3693 7971 3867 7974
rect 3686 7968 3867 7971
rect 3495 7948 3508 7950
rect 3523 7948 3557 7950
rect 3495 7932 3569 7948
rect 3596 7944 3609 7958
rect 3624 7944 3640 7960
rect 3686 7955 3697 7968
rect 3479 7910 3480 7926
rect 3495 7910 3508 7932
rect 3523 7910 3553 7932
rect 3596 7928 3658 7944
rect 3686 7937 3697 7953
rect 3702 7948 3712 7968
rect 3722 7948 3736 7968
rect 3739 7955 3748 7968
rect 3764 7955 3773 7968
rect 3702 7937 3736 7948
rect 3739 7937 3748 7953
rect 3764 7937 3773 7953
rect 3780 7948 3790 7968
rect 3800 7948 3814 7968
rect 3815 7955 3826 7968
rect 3780 7937 3814 7948
rect 3815 7937 3826 7953
rect 3872 7944 3888 7960
rect 3895 7958 3925 8010
rect 3959 8006 3960 8013
rect 3944 7998 3960 8006
rect 3931 7966 3944 7985
rect 3959 7966 3989 7982
rect 3931 7950 4005 7966
rect 3931 7948 3944 7950
rect 3959 7948 3993 7950
rect 3596 7926 3609 7928
rect 3624 7926 3658 7928
rect 3596 7910 3658 7926
rect 3702 7921 3718 7924
rect 3780 7921 3810 7932
rect 3858 7928 3904 7944
rect 3931 7932 4005 7948
rect 3858 7926 3892 7928
rect 3857 7910 3904 7926
rect 3931 7910 3944 7932
rect 3959 7910 3989 7932
rect 4016 7910 4017 7926
rect 4032 7910 4045 8070
rect 4075 7966 4088 8070
rect 4133 8048 4134 8058
rect 4149 8048 4162 8058
rect 4133 8044 4162 8048
rect 4167 8044 4197 8070
rect 4215 8056 4231 8058
rect 4303 8056 4356 8070
rect 4304 8054 4368 8056
rect 4411 8054 4426 8070
rect 4475 8067 4505 8070
rect 4475 8064 4511 8067
rect 4441 8056 4457 8058
rect 4215 8044 4230 8048
rect 4133 8042 4230 8044
rect 4258 8042 4426 8054
rect 4442 8044 4457 8048
rect 4475 8045 4514 8064
rect 4533 8058 4540 8059
rect 4539 8051 4540 8058
rect 4523 8048 4524 8051
rect 4539 8048 4552 8051
rect 4475 8044 4505 8045
rect 4514 8044 4520 8045
rect 4523 8044 4552 8048
rect 4442 8043 4552 8044
rect 4442 8042 4558 8043
rect 4117 8034 4168 8042
rect 4117 8022 4142 8034
rect 4149 8022 4168 8034
rect 4199 8034 4249 8042
rect 4199 8026 4215 8034
rect 4222 8032 4249 8034
rect 4258 8032 4479 8042
rect 4222 8022 4479 8032
rect 4508 8034 4558 8042
rect 4508 8025 4524 8034
rect 4117 8014 4168 8022
rect 4215 8014 4479 8022
rect 4505 8022 4524 8025
rect 4531 8022 4558 8034
rect 4505 8014 4558 8022
rect 4133 8006 4134 8014
rect 4149 8006 4162 8014
rect 4133 7998 4149 8006
rect 4130 7991 4149 7994
rect 4130 7982 4152 7991
rect 4103 7972 4152 7982
rect 4103 7966 4133 7972
rect 4152 7967 4157 7972
rect 4075 7950 4149 7966
rect 4167 7958 4197 8014
rect 4232 8004 4440 8014
rect 4475 8010 4520 8014
rect 4523 8013 4524 8014
rect 4539 8013 4552 8014
rect 4258 7974 4447 8004
rect 4273 7971 4447 7974
rect 4266 7968 4447 7971
rect 4075 7948 4088 7950
rect 4103 7948 4137 7950
rect 4075 7932 4149 7948
rect 4176 7944 4189 7958
rect 4204 7944 4220 7960
rect 4266 7955 4277 7968
rect 4059 7910 4060 7926
rect 4075 7910 4088 7932
rect 4103 7910 4133 7932
rect 4176 7928 4238 7944
rect 4266 7937 4277 7953
rect 4282 7948 4292 7968
rect 4302 7948 4316 7968
rect 4319 7955 4328 7968
rect 4344 7955 4353 7968
rect 4282 7937 4316 7948
rect 4319 7937 4328 7953
rect 4344 7937 4353 7953
rect 4360 7948 4370 7968
rect 4380 7948 4394 7968
rect 4395 7955 4406 7968
rect 4360 7937 4394 7948
rect 4395 7937 4406 7953
rect 4452 7944 4468 7960
rect 4475 7958 4505 8010
rect 4539 8006 4540 8013
rect 4524 7998 4540 8006
rect 4511 7966 4524 7985
rect 4539 7966 4569 7982
rect 4511 7950 4585 7966
rect 4511 7948 4524 7950
rect 4539 7948 4573 7950
rect 4176 7926 4189 7928
rect 4204 7926 4238 7928
rect 4176 7910 4238 7926
rect 4282 7921 4298 7924
rect 4360 7921 4390 7932
rect 4438 7928 4484 7944
rect 4511 7932 4585 7948
rect 4438 7926 4472 7928
rect 4437 7910 4484 7926
rect 4511 7910 4524 7932
rect 4539 7910 4569 7932
rect 4596 7910 4597 7926
rect 4612 7910 4625 8070
rect -7 7902 34 7910
rect -7 7876 8 7902
rect 15 7876 34 7902
rect 98 7898 160 7910
rect 172 7898 247 7910
rect 305 7898 380 7910
rect 392 7898 423 7910
rect 429 7898 464 7910
rect 98 7896 260 7898
rect -7 7868 34 7876
rect 116 7872 129 7896
rect 144 7894 159 7896
rect -1 7858 0 7868
rect 15 7858 28 7868
rect 43 7858 73 7872
rect 116 7858 159 7872
rect 183 7869 190 7876
rect 193 7872 260 7896
rect 292 7896 464 7898
rect 262 7874 290 7878
rect 292 7874 372 7896
rect 393 7894 408 7896
rect 262 7872 372 7874
rect 193 7868 372 7872
rect 166 7858 196 7868
rect 198 7858 351 7868
rect 359 7858 389 7868
rect 393 7858 423 7872
rect 451 7858 464 7896
rect 536 7902 571 7910
rect 536 7876 537 7902
rect 544 7876 571 7902
rect 479 7858 509 7872
rect 536 7868 571 7876
rect 573 7902 614 7910
rect 573 7876 588 7902
rect 595 7876 614 7902
rect 678 7898 740 7910
rect 752 7898 827 7910
rect 885 7898 960 7910
rect 972 7898 1003 7910
rect 1009 7898 1044 7910
rect 678 7896 840 7898
rect 573 7868 614 7876
rect 696 7872 709 7896
rect 724 7894 739 7896
rect 536 7858 537 7868
rect 552 7858 565 7868
rect 579 7858 580 7868
rect 595 7858 608 7868
rect 623 7858 653 7872
rect 696 7858 739 7872
rect 763 7869 770 7876
rect 773 7872 840 7896
rect 872 7896 1044 7898
rect 842 7874 870 7878
rect 872 7874 952 7896
rect 973 7894 988 7896
rect 842 7872 952 7874
rect 773 7868 952 7872
rect 746 7858 776 7868
rect 778 7858 931 7868
rect 939 7858 969 7868
rect 973 7858 1003 7872
rect 1031 7858 1044 7896
rect 1116 7902 1151 7910
rect 1116 7876 1117 7902
rect 1124 7876 1151 7902
rect 1059 7858 1089 7872
rect 1116 7868 1151 7876
rect 1153 7902 1194 7910
rect 1153 7876 1168 7902
rect 1175 7876 1194 7902
rect 1258 7898 1320 7910
rect 1332 7898 1407 7910
rect 1465 7898 1540 7910
rect 1552 7898 1583 7910
rect 1589 7898 1624 7910
rect 1258 7896 1420 7898
rect 1153 7868 1194 7876
rect 1276 7872 1289 7896
rect 1304 7894 1319 7896
rect 1116 7858 1117 7868
rect 1132 7858 1145 7868
rect 1159 7858 1160 7868
rect 1175 7858 1188 7868
rect 1203 7858 1233 7872
rect 1276 7858 1319 7872
rect 1343 7869 1350 7876
rect 1353 7872 1420 7896
rect 1452 7896 1624 7898
rect 1422 7874 1450 7878
rect 1452 7874 1532 7896
rect 1553 7894 1568 7896
rect 1422 7872 1532 7874
rect 1353 7868 1532 7872
rect 1326 7858 1356 7868
rect 1358 7858 1511 7868
rect 1519 7858 1549 7868
rect 1553 7858 1583 7872
rect 1611 7858 1624 7896
rect 1696 7902 1731 7910
rect 1696 7876 1697 7902
rect 1704 7876 1731 7902
rect 1639 7858 1669 7872
rect 1696 7868 1731 7876
rect 1733 7902 1774 7910
rect 1733 7876 1748 7902
rect 1755 7876 1774 7902
rect 1838 7898 1900 7910
rect 1912 7898 1987 7910
rect 2045 7898 2120 7910
rect 2132 7898 2163 7910
rect 2169 7898 2204 7910
rect 1838 7896 2000 7898
rect 1733 7868 1774 7876
rect 1856 7872 1869 7896
rect 1884 7894 1899 7896
rect 1696 7858 1697 7868
rect 1712 7858 1725 7868
rect 1739 7858 1740 7868
rect 1755 7858 1768 7868
rect 1783 7858 1813 7872
rect 1856 7858 1899 7872
rect 1923 7869 1930 7876
rect 1933 7872 2000 7896
rect 2032 7896 2204 7898
rect 2002 7874 2030 7878
rect 2032 7874 2112 7896
rect 2133 7894 2148 7896
rect 2002 7872 2112 7874
rect 1933 7868 2112 7872
rect 1906 7858 1936 7868
rect 1938 7858 2091 7868
rect 2099 7858 2129 7868
rect 2133 7858 2163 7872
rect 2191 7858 2204 7896
rect 2276 7902 2311 7910
rect 2276 7876 2277 7902
rect 2284 7876 2311 7902
rect 2219 7858 2249 7872
rect 2276 7868 2311 7876
rect 2313 7902 2354 7910
rect 2313 7876 2328 7902
rect 2335 7876 2354 7902
rect 2418 7898 2480 7910
rect 2492 7898 2567 7910
rect 2625 7898 2700 7910
rect 2712 7898 2743 7910
rect 2749 7898 2784 7910
rect 2418 7896 2580 7898
rect 2313 7868 2354 7876
rect 2436 7872 2449 7896
rect 2464 7894 2479 7896
rect 2276 7858 2277 7868
rect 2292 7858 2305 7868
rect 2319 7858 2320 7868
rect 2335 7858 2348 7868
rect 2363 7858 2393 7872
rect 2436 7858 2479 7872
rect 2503 7869 2510 7876
rect 2513 7872 2580 7896
rect 2612 7896 2784 7898
rect 2582 7874 2610 7878
rect 2612 7874 2692 7896
rect 2713 7894 2728 7896
rect 2582 7872 2692 7874
rect 2513 7868 2692 7872
rect 2486 7858 2516 7868
rect 2518 7858 2671 7868
rect 2679 7858 2709 7868
rect 2713 7858 2743 7872
rect 2771 7858 2784 7896
rect 2856 7902 2891 7910
rect 2856 7876 2857 7902
rect 2864 7876 2891 7902
rect 2799 7858 2829 7872
rect 2856 7868 2891 7876
rect 2893 7902 2934 7910
rect 2893 7876 2908 7902
rect 2915 7876 2934 7902
rect 2998 7898 3060 7910
rect 3072 7898 3147 7910
rect 3205 7898 3280 7910
rect 3292 7898 3323 7910
rect 3329 7898 3364 7910
rect 2998 7896 3160 7898
rect 2893 7868 2934 7876
rect 3016 7872 3029 7896
rect 3044 7894 3059 7896
rect 2856 7858 2857 7868
rect 2872 7858 2885 7868
rect 2899 7858 2900 7868
rect 2915 7858 2928 7868
rect 2943 7858 2973 7872
rect 3016 7858 3059 7872
rect 3083 7869 3090 7876
rect 3093 7872 3160 7896
rect 3192 7896 3364 7898
rect 3162 7874 3190 7878
rect 3192 7874 3272 7896
rect 3293 7894 3308 7896
rect 3162 7872 3272 7874
rect 3093 7868 3272 7872
rect 3066 7858 3096 7868
rect 3098 7858 3251 7868
rect 3259 7858 3289 7868
rect 3293 7858 3323 7872
rect 3351 7858 3364 7896
rect 3436 7902 3471 7910
rect 3436 7876 3437 7902
rect 3444 7876 3471 7902
rect 3379 7858 3409 7872
rect 3436 7868 3471 7876
rect 3473 7902 3514 7910
rect 3473 7876 3488 7902
rect 3495 7876 3514 7902
rect 3578 7898 3640 7910
rect 3652 7898 3727 7910
rect 3785 7898 3860 7910
rect 3872 7898 3903 7910
rect 3909 7898 3944 7910
rect 3578 7896 3740 7898
rect 3473 7868 3514 7876
rect 3596 7872 3609 7896
rect 3624 7894 3639 7896
rect 3436 7858 3437 7868
rect 3452 7858 3465 7868
rect 3479 7858 3480 7868
rect 3495 7858 3508 7868
rect 3523 7858 3553 7872
rect 3596 7858 3639 7872
rect 3663 7869 3670 7876
rect 3673 7872 3740 7896
rect 3772 7896 3944 7898
rect 3742 7874 3770 7878
rect 3772 7874 3852 7896
rect 3873 7894 3888 7896
rect 3742 7872 3852 7874
rect 3673 7868 3852 7872
rect 3646 7858 3676 7868
rect 3678 7858 3831 7868
rect 3839 7858 3869 7868
rect 3873 7858 3903 7872
rect 3931 7858 3944 7896
rect 4016 7902 4051 7910
rect 4016 7876 4017 7902
rect 4024 7876 4051 7902
rect 3959 7858 3989 7872
rect 4016 7868 4051 7876
rect 4053 7902 4094 7910
rect 4053 7876 4068 7902
rect 4075 7876 4094 7902
rect 4158 7898 4220 7910
rect 4232 7898 4307 7910
rect 4365 7898 4440 7910
rect 4452 7898 4483 7910
rect 4489 7898 4524 7910
rect 4158 7896 4320 7898
rect 4053 7868 4094 7876
rect 4176 7872 4189 7896
rect 4204 7894 4219 7896
rect 4016 7858 4017 7868
rect 4032 7858 4045 7868
rect 4059 7858 4060 7868
rect 4075 7858 4088 7868
rect 4103 7858 4133 7872
rect 4176 7858 4219 7872
rect 4243 7869 4250 7876
rect 4253 7872 4320 7896
rect 4352 7896 4524 7898
rect 4322 7874 4350 7878
rect 4352 7874 4432 7896
rect 4453 7894 4468 7896
rect 4322 7872 4432 7874
rect 4253 7868 4432 7872
rect 4226 7858 4256 7868
rect 4258 7858 4411 7868
rect 4419 7858 4449 7868
rect 4453 7858 4483 7872
rect 4511 7858 4524 7896
rect 4596 7902 4631 7910
rect 4596 7876 4597 7902
rect 4604 7876 4631 7902
rect 4539 7858 4569 7872
rect 4596 7868 4631 7876
rect 4596 7858 4597 7868
rect 4612 7858 4625 7868
rect -1 7852 4625 7858
rect 0 7844 4625 7852
rect 15 7814 28 7844
rect 43 7826 73 7844
rect 116 7830 130 7844
rect 166 7830 386 7844
rect 117 7828 130 7830
rect 83 7816 98 7828
rect 80 7814 102 7816
rect 107 7814 137 7828
rect 198 7826 351 7830
rect 180 7814 372 7826
rect 415 7814 445 7828
rect 451 7814 464 7844
rect 479 7826 509 7844
rect 552 7814 565 7844
rect 595 7814 608 7844
rect 623 7826 653 7844
rect 696 7830 710 7844
rect 746 7830 966 7844
rect 697 7828 710 7830
rect 663 7816 678 7828
rect 660 7814 682 7816
rect 687 7814 717 7828
rect 778 7826 931 7830
rect 760 7814 952 7826
rect 995 7814 1025 7828
rect 1031 7814 1044 7844
rect 1059 7826 1089 7844
rect 1132 7814 1145 7844
rect 1175 7814 1188 7844
rect 1203 7826 1233 7844
rect 1276 7830 1290 7844
rect 1326 7830 1546 7844
rect 1277 7828 1290 7830
rect 1243 7816 1258 7828
rect 1240 7814 1262 7816
rect 1267 7814 1297 7828
rect 1358 7826 1511 7830
rect 1340 7814 1532 7826
rect 1575 7814 1605 7828
rect 1611 7814 1624 7844
rect 1639 7826 1669 7844
rect 1712 7814 1725 7844
rect 1755 7814 1768 7844
rect 1783 7826 1813 7844
rect 1856 7830 1870 7844
rect 1906 7830 2126 7844
rect 1857 7828 1870 7830
rect 1823 7816 1838 7828
rect 1820 7814 1842 7816
rect 1847 7814 1877 7828
rect 1938 7826 2091 7830
rect 1920 7814 2112 7826
rect 2155 7814 2185 7828
rect 2191 7814 2204 7844
rect 2219 7826 2249 7844
rect 2292 7814 2305 7844
rect 2335 7814 2348 7844
rect 2363 7826 2393 7844
rect 2436 7830 2450 7844
rect 2486 7830 2706 7844
rect 2437 7828 2450 7830
rect 2403 7816 2418 7828
rect 2400 7814 2422 7816
rect 2427 7814 2457 7828
rect 2518 7826 2671 7830
rect 2500 7814 2692 7826
rect 2735 7814 2765 7828
rect 2771 7814 2784 7844
rect 2799 7826 2829 7844
rect 2872 7814 2885 7844
rect 2915 7814 2928 7844
rect 2943 7826 2973 7844
rect 3016 7830 3030 7844
rect 3066 7830 3286 7844
rect 3017 7828 3030 7830
rect 2983 7816 2998 7828
rect 2980 7814 3002 7816
rect 3007 7814 3037 7828
rect 3098 7826 3251 7830
rect 3080 7814 3272 7826
rect 3315 7814 3345 7828
rect 3351 7814 3364 7844
rect 3379 7826 3409 7844
rect 3452 7814 3465 7844
rect 3495 7814 3508 7844
rect 3523 7826 3553 7844
rect 3596 7830 3610 7844
rect 3646 7830 3866 7844
rect 3597 7828 3610 7830
rect 3563 7816 3578 7828
rect 3560 7814 3582 7816
rect 3587 7814 3617 7828
rect 3678 7826 3831 7830
rect 3660 7814 3852 7826
rect 3895 7814 3925 7828
rect 3931 7814 3944 7844
rect 3959 7826 3989 7844
rect 4032 7814 4045 7844
rect 4075 7814 4088 7844
rect 4103 7826 4133 7844
rect 4176 7830 4190 7844
rect 4226 7830 4446 7844
rect 4177 7828 4190 7830
rect 4143 7816 4158 7828
rect 4140 7814 4162 7816
rect 4167 7814 4197 7828
rect 4258 7826 4411 7830
rect 4240 7814 4432 7826
rect 4475 7814 4505 7828
rect 4511 7814 4524 7844
rect 4539 7826 4569 7844
rect 4612 7814 4625 7844
rect 0 7800 4625 7814
rect 15 7696 28 7800
rect 73 7778 74 7788
rect 89 7778 102 7788
rect 73 7774 102 7778
rect 107 7774 137 7800
rect 155 7786 171 7788
rect 243 7786 296 7800
rect 244 7784 308 7786
rect 351 7784 366 7800
rect 415 7797 445 7800
rect 415 7794 451 7797
rect 381 7786 397 7788
rect 155 7774 170 7778
rect 73 7772 170 7774
rect 198 7772 366 7784
rect 382 7774 397 7778
rect 415 7775 454 7794
rect 473 7788 480 7789
rect 479 7781 480 7788
rect 463 7778 464 7781
rect 479 7778 492 7781
rect 415 7774 445 7775
rect 454 7774 460 7775
rect 463 7774 492 7778
rect 382 7773 492 7774
rect 382 7772 498 7773
rect 57 7764 108 7772
rect 57 7752 82 7764
rect 89 7752 108 7764
rect 139 7764 189 7772
rect 139 7756 155 7764
rect 162 7762 189 7764
rect 198 7762 419 7772
rect 162 7752 419 7762
rect 448 7764 498 7772
rect 448 7755 464 7764
rect 57 7744 108 7752
rect 155 7744 419 7752
rect 445 7752 464 7755
rect 471 7752 498 7764
rect 445 7744 498 7752
rect 73 7736 74 7744
rect 89 7736 102 7744
rect 73 7728 89 7736
rect 70 7721 89 7724
rect 70 7712 92 7721
rect 43 7702 92 7712
rect 43 7696 73 7702
rect 92 7697 97 7702
rect 15 7680 89 7696
rect 107 7688 137 7744
rect 172 7734 380 7744
rect 415 7740 460 7744
rect 463 7743 464 7744
rect 479 7743 492 7744
rect 198 7704 387 7734
rect 213 7701 387 7704
rect 206 7698 387 7701
rect 15 7678 28 7680
rect 43 7678 77 7680
rect 15 7662 89 7678
rect 116 7674 129 7688
rect 144 7674 160 7690
rect 206 7685 217 7698
rect -1 7640 0 7656
rect 15 7640 28 7662
rect 43 7640 73 7662
rect 116 7658 178 7674
rect 206 7667 217 7683
rect 222 7678 232 7698
rect 242 7678 256 7698
rect 259 7685 268 7698
rect 284 7685 293 7698
rect 222 7667 256 7678
rect 259 7667 268 7683
rect 284 7667 293 7683
rect 300 7678 310 7698
rect 320 7678 334 7698
rect 335 7685 346 7698
rect 300 7667 334 7678
rect 335 7667 346 7683
rect 392 7674 408 7690
rect 415 7688 445 7740
rect 479 7736 480 7743
rect 464 7728 480 7736
rect 451 7696 464 7715
rect 479 7696 509 7712
rect 451 7680 525 7696
rect 451 7678 464 7680
rect 479 7678 513 7680
rect 116 7656 129 7658
rect 144 7656 178 7658
rect 116 7640 178 7656
rect 222 7651 238 7654
rect 300 7651 330 7662
rect 378 7658 424 7674
rect 451 7662 525 7678
rect 378 7656 412 7658
rect 377 7640 424 7656
rect 451 7640 464 7662
rect 479 7640 509 7662
rect 536 7640 537 7656
rect 552 7640 565 7800
rect 595 7696 608 7800
rect 653 7778 654 7788
rect 669 7778 682 7788
rect 653 7774 682 7778
rect 687 7774 717 7800
rect 735 7786 751 7788
rect 823 7786 876 7800
rect 824 7784 888 7786
rect 931 7784 946 7800
rect 995 7797 1025 7800
rect 995 7794 1031 7797
rect 961 7786 977 7788
rect 735 7774 750 7778
rect 653 7772 750 7774
rect 778 7772 946 7784
rect 962 7774 977 7778
rect 995 7775 1034 7794
rect 1053 7788 1060 7789
rect 1059 7781 1060 7788
rect 1043 7778 1044 7781
rect 1059 7778 1072 7781
rect 995 7774 1025 7775
rect 1034 7774 1040 7775
rect 1043 7774 1072 7778
rect 962 7773 1072 7774
rect 962 7772 1078 7773
rect 637 7764 688 7772
rect 637 7752 662 7764
rect 669 7752 688 7764
rect 719 7764 769 7772
rect 719 7756 735 7764
rect 742 7762 769 7764
rect 778 7762 999 7772
rect 742 7752 999 7762
rect 1028 7764 1078 7772
rect 1028 7755 1044 7764
rect 637 7744 688 7752
rect 735 7744 999 7752
rect 1025 7752 1044 7755
rect 1051 7752 1078 7764
rect 1025 7744 1078 7752
rect 653 7736 654 7744
rect 669 7736 682 7744
rect 653 7728 669 7736
rect 650 7721 669 7724
rect 650 7712 672 7721
rect 623 7702 672 7712
rect 623 7696 653 7702
rect 672 7697 677 7702
rect 595 7680 669 7696
rect 687 7688 717 7744
rect 752 7734 960 7744
rect 995 7740 1040 7744
rect 1043 7743 1044 7744
rect 1059 7743 1072 7744
rect 778 7704 967 7734
rect 793 7701 967 7704
rect 786 7698 967 7701
rect 595 7678 608 7680
rect 623 7678 657 7680
rect 595 7662 669 7678
rect 696 7674 709 7688
rect 724 7674 740 7690
rect 786 7685 797 7698
rect 579 7640 580 7656
rect 595 7640 608 7662
rect 623 7640 653 7662
rect 696 7658 758 7674
rect 786 7667 797 7683
rect 802 7678 812 7698
rect 822 7678 836 7698
rect 839 7685 848 7698
rect 864 7685 873 7698
rect 802 7667 836 7678
rect 839 7667 848 7683
rect 864 7667 873 7683
rect 880 7678 890 7698
rect 900 7678 914 7698
rect 915 7685 926 7698
rect 880 7667 914 7678
rect 915 7667 926 7683
rect 972 7674 988 7690
rect 995 7688 1025 7740
rect 1059 7736 1060 7743
rect 1044 7728 1060 7736
rect 1031 7696 1044 7715
rect 1059 7696 1089 7712
rect 1031 7680 1105 7696
rect 1031 7678 1044 7680
rect 1059 7678 1093 7680
rect 696 7656 709 7658
rect 724 7656 758 7658
rect 696 7640 758 7656
rect 802 7651 818 7654
rect 880 7651 910 7662
rect 958 7658 1004 7674
rect 1031 7662 1105 7678
rect 958 7656 992 7658
rect 957 7640 1004 7656
rect 1031 7640 1044 7662
rect 1059 7640 1089 7662
rect 1116 7640 1117 7656
rect 1132 7640 1145 7800
rect 1175 7696 1188 7800
rect 1233 7778 1234 7788
rect 1249 7778 1262 7788
rect 1233 7774 1262 7778
rect 1267 7774 1297 7800
rect 1315 7786 1331 7788
rect 1403 7786 1456 7800
rect 1404 7784 1468 7786
rect 1511 7784 1526 7800
rect 1575 7797 1605 7800
rect 1575 7794 1611 7797
rect 1541 7786 1557 7788
rect 1315 7774 1330 7778
rect 1233 7772 1330 7774
rect 1358 7772 1526 7784
rect 1542 7774 1557 7778
rect 1575 7775 1614 7794
rect 1633 7788 1640 7789
rect 1639 7781 1640 7788
rect 1623 7778 1624 7781
rect 1639 7778 1652 7781
rect 1575 7774 1605 7775
rect 1614 7774 1620 7775
rect 1623 7774 1652 7778
rect 1542 7773 1652 7774
rect 1542 7772 1658 7773
rect 1217 7764 1268 7772
rect 1217 7752 1242 7764
rect 1249 7752 1268 7764
rect 1299 7764 1349 7772
rect 1299 7756 1315 7764
rect 1322 7762 1349 7764
rect 1358 7762 1579 7772
rect 1322 7752 1579 7762
rect 1608 7764 1658 7772
rect 1608 7755 1624 7764
rect 1217 7744 1268 7752
rect 1315 7744 1579 7752
rect 1605 7752 1624 7755
rect 1631 7752 1658 7764
rect 1605 7744 1658 7752
rect 1233 7736 1234 7744
rect 1249 7736 1262 7744
rect 1233 7728 1249 7736
rect 1230 7721 1249 7724
rect 1230 7712 1252 7721
rect 1203 7702 1252 7712
rect 1203 7696 1233 7702
rect 1252 7697 1257 7702
rect 1175 7680 1249 7696
rect 1267 7688 1297 7744
rect 1332 7734 1540 7744
rect 1575 7740 1620 7744
rect 1623 7743 1624 7744
rect 1639 7743 1652 7744
rect 1358 7704 1547 7734
rect 1373 7701 1547 7704
rect 1366 7698 1547 7701
rect 1175 7678 1188 7680
rect 1203 7678 1237 7680
rect 1175 7662 1249 7678
rect 1276 7674 1289 7688
rect 1304 7674 1320 7690
rect 1366 7685 1377 7698
rect 1159 7640 1160 7656
rect 1175 7640 1188 7662
rect 1203 7640 1233 7662
rect 1276 7658 1338 7674
rect 1366 7667 1377 7683
rect 1382 7678 1392 7698
rect 1402 7678 1416 7698
rect 1419 7685 1428 7698
rect 1444 7685 1453 7698
rect 1382 7667 1416 7678
rect 1419 7667 1428 7683
rect 1444 7667 1453 7683
rect 1460 7678 1470 7698
rect 1480 7678 1494 7698
rect 1495 7685 1506 7698
rect 1460 7667 1494 7678
rect 1495 7667 1506 7683
rect 1552 7674 1568 7690
rect 1575 7688 1605 7740
rect 1639 7736 1640 7743
rect 1624 7728 1640 7736
rect 1611 7696 1624 7715
rect 1639 7696 1669 7712
rect 1611 7680 1685 7696
rect 1611 7678 1624 7680
rect 1639 7678 1673 7680
rect 1276 7656 1289 7658
rect 1304 7656 1338 7658
rect 1276 7640 1338 7656
rect 1382 7651 1398 7654
rect 1460 7651 1490 7662
rect 1538 7658 1584 7674
rect 1611 7662 1685 7678
rect 1538 7656 1572 7658
rect 1537 7640 1584 7656
rect 1611 7640 1624 7662
rect 1639 7640 1669 7662
rect 1696 7640 1697 7656
rect 1712 7640 1725 7800
rect 1755 7696 1768 7800
rect 1813 7778 1814 7788
rect 1829 7778 1842 7788
rect 1813 7774 1842 7778
rect 1847 7774 1877 7800
rect 1895 7786 1911 7788
rect 1983 7786 2036 7800
rect 1984 7784 2048 7786
rect 2091 7784 2106 7800
rect 2155 7797 2185 7800
rect 2155 7794 2191 7797
rect 2121 7786 2137 7788
rect 1895 7774 1910 7778
rect 1813 7772 1910 7774
rect 1938 7772 2106 7784
rect 2122 7774 2137 7778
rect 2155 7775 2194 7794
rect 2213 7788 2220 7789
rect 2219 7781 2220 7788
rect 2203 7778 2204 7781
rect 2219 7778 2232 7781
rect 2155 7774 2185 7775
rect 2194 7774 2200 7775
rect 2203 7774 2232 7778
rect 2122 7773 2232 7774
rect 2122 7772 2238 7773
rect 1797 7764 1848 7772
rect 1797 7752 1822 7764
rect 1829 7752 1848 7764
rect 1879 7764 1929 7772
rect 1879 7756 1895 7764
rect 1902 7762 1929 7764
rect 1938 7762 2159 7772
rect 1902 7752 2159 7762
rect 2188 7764 2238 7772
rect 2188 7755 2204 7764
rect 1797 7744 1848 7752
rect 1895 7744 2159 7752
rect 2185 7752 2204 7755
rect 2211 7752 2238 7764
rect 2185 7744 2238 7752
rect 1813 7736 1814 7744
rect 1829 7736 1842 7744
rect 1813 7728 1829 7736
rect 1810 7721 1829 7724
rect 1810 7712 1832 7721
rect 1783 7702 1832 7712
rect 1783 7696 1813 7702
rect 1832 7697 1837 7702
rect 1755 7680 1829 7696
rect 1847 7688 1877 7744
rect 1912 7734 2120 7744
rect 2155 7740 2200 7744
rect 2203 7743 2204 7744
rect 2219 7743 2232 7744
rect 1938 7704 2127 7734
rect 1953 7701 2127 7704
rect 1946 7698 2127 7701
rect 1755 7678 1768 7680
rect 1783 7678 1817 7680
rect 1755 7662 1829 7678
rect 1856 7674 1869 7688
rect 1884 7674 1900 7690
rect 1946 7685 1957 7698
rect 1739 7640 1740 7656
rect 1755 7640 1768 7662
rect 1783 7640 1813 7662
rect 1856 7658 1918 7674
rect 1946 7667 1957 7683
rect 1962 7678 1972 7698
rect 1982 7678 1996 7698
rect 1999 7685 2008 7698
rect 2024 7685 2033 7698
rect 1962 7667 1996 7678
rect 1999 7667 2008 7683
rect 2024 7667 2033 7683
rect 2040 7678 2050 7698
rect 2060 7678 2074 7698
rect 2075 7685 2086 7698
rect 2040 7667 2074 7678
rect 2075 7667 2086 7683
rect 2132 7674 2148 7690
rect 2155 7688 2185 7740
rect 2219 7736 2220 7743
rect 2204 7728 2220 7736
rect 2191 7696 2204 7715
rect 2219 7696 2249 7712
rect 2191 7680 2265 7696
rect 2191 7678 2204 7680
rect 2219 7678 2253 7680
rect 1856 7656 1869 7658
rect 1884 7656 1918 7658
rect 1856 7640 1918 7656
rect 1962 7651 1978 7654
rect 2040 7651 2070 7662
rect 2118 7658 2164 7674
rect 2191 7662 2265 7678
rect 2118 7656 2152 7658
rect 2117 7640 2164 7656
rect 2191 7640 2204 7662
rect 2219 7640 2249 7662
rect 2276 7640 2277 7656
rect 2292 7640 2305 7800
rect 2335 7696 2348 7800
rect 2393 7778 2394 7788
rect 2409 7778 2422 7788
rect 2393 7774 2422 7778
rect 2427 7774 2457 7800
rect 2475 7786 2491 7788
rect 2563 7786 2616 7800
rect 2564 7784 2628 7786
rect 2671 7784 2686 7800
rect 2735 7797 2765 7800
rect 2735 7794 2771 7797
rect 2701 7786 2717 7788
rect 2475 7774 2490 7778
rect 2393 7772 2490 7774
rect 2518 7772 2686 7784
rect 2702 7774 2717 7778
rect 2735 7775 2774 7794
rect 2793 7788 2800 7789
rect 2799 7781 2800 7788
rect 2783 7778 2784 7781
rect 2799 7778 2812 7781
rect 2735 7774 2765 7775
rect 2774 7774 2780 7775
rect 2783 7774 2812 7778
rect 2702 7773 2812 7774
rect 2702 7772 2818 7773
rect 2377 7764 2428 7772
rect 2377 7752 2402 7764
rect 2409 7752 2428 7764
rect 2459 7764 2509 7772
rect 2459 7756 2475 7764
rect 2482 7762 2509 7764
rect 2518 7762 2739 7772
rect 2482 7752 2739 7762
rect 2768 7764 2818 7772
rect 2768 7755 2784 7764
rect 2377 7744 2428 7752
rect 2475 7744 2739 7752
rect 2765 7752 2784 7755
rect 2791 7752 2818 7764
rect 2765 7744 2818 7752
rect 2393 7736 2394 7744
rect 2409 7736 2422 7744
rect 2393 7728 2409 7736
rect 2390 7721 2409 7724
rect 2390 7712 2412 7721
rect 2363 7702 2412 7712
rect 2363 7696 2393 7702
rect 2412 7697 2417 7702
rect 2335 7680 2409 7696
rect 2427 7688 2457 7744
rect 2492 7734 2700 7744
rect 2735 7740 2780 7744
rect 2783 7743 2784 7744
rect 2799 7743 2812 7744
rect 2518 7704 2707 7734
rect 2533 7701 2707 7704
rect 2526 7698 2707 7701
rect 2335 7678 2348 7680
rect 2363 7678 2397 7680
rect 2335 7662 2409 7678
rect 2436 7674 2449 7688
rect 2464 7674 2480 7690
rect 2526 7685 2537 7698
rect 2319 7640 2320 7656
rect 2335 7640 2348 7662
rect 2363 7640 2393 7662
rect 2436 7658 2498 7674
rect 2526 7667 2537 7683
rect 2542 7678 2552 7698
rect 2562 7678 2576 7698
rect 2579 7685 2588 7698
rect 2604 7685 2613 7698
rect 2542 7667 2576 7678
rect 2579 7667 2588 7683
rect 2604 7667 2613 7683
rect 2620 7678 2630 7698
rect 2640 7678 2654 7698
rect 2655 7685 2666 7698
rect 2620 7667 2654 7678
rect 2655 7667 2666 7683
rect 2712 7674 2728 7690
rect 2735 7688 2765 7740
rect 2799 7736 2800 7743
rect 2784 7728 2800 7736
rect 2771 7696 2784 7715
rect 2799 7696 2829 7712
rect 2771 7680 2845 7696
rect 2771 7678 2784 7680
rect 2799 7678 2833 7680
rect 2436 7656 2449 7658
rect 2464 7656 2498 7658
rect 2436 7640 2498 7656
rect 2542 7651 2558 7654
rect 2620 7651 2650 7662
rect 2698 7658 2744 7674
rect 2771 7662 2845 7678
rect 2698 7656 2732 7658
rect 2697 7640 2744 7656
rect 2771 7640 2784 7662
rect 2799 7640 2829 7662
rect 2856 7640 2857 7656
rect 2872 7640 2885 7800
rect 2915 7696 2928 7800
rect 2973 7778 2974 7788
rect 2989 7778 3002 7788
rect 2973 7774 3002 7778
rect 3007 7774 3037 7800
rect 3055 7786 3071 7788
rect 3143 7786 3196 7800
rect 3144 7784 3208 7786
rect 3251 7784 3266 7800
rect 3315 7797 3345 7800
rect 3315 7794 3351 7797
rect 3281 7786 3297 7788
rect 3055 7774 3070 7778
rect 2973 7772 3070 7774
rect 3098 7772 3266 7784
rect 3282 7774 3297 7778
rect 3315 7775 3354 7794
rect 3373 7788 3380 7789
rect 3379 7781 3380 7788
rect 3363 7778 3364 7781
rect 3379 7778 3392 7781
rect 3315 7774 3345 7775
rect 3354 7774 3360 7775
rect 3363 7774 3392 7778
rect 3282 7773 3392 7774
rect 3282 7772 3398 7773
rect 2957 7764 3008 7772
rect 2957 7752 2982 7764
rect 2989 7752 3008 7764
rect 3039 7764 3089 7772
rect 3039 7756 3055 7764
rect 3062 7762 3089 7764
rect 3098 7762 3319 7772
rect 3062 7752 3319 7762
rect 3348 7764 3398 7772
rect 3348 7755 3364 7764
rect 2957 7744 3008 7752
rect 3055 7744 3319 7752
rect 3345 7752 3364 7755
rect 3371 7752 3398 7764
rect 3345 7744 3398 7752
rect 2973 7736 2974 7744
rect 2989 7736 3002 7744
rect 2973 7728 2989 7736
rect 2970 7721 2989 7724
rect 2970 7712 2992 7721
rect 2943 7702 2992 7712
rect 2943 7696 2973 7702
rect 2992 7697 2997 7702
rect 2915 7680 2989 7696
rect 3007 7688 3037 7744
rect 3072 7734 3280 7744
rect 3315 7740 3360 7744
rect 3363 7743 3364 7744
rect 3379 7743 3392 7744
rect 3098 7704 3287 7734
rect 3113 7701 3287 7704
rect 3106 7698 3287 7701
rect 2915 7678 2928 7680
rect 2943 7678 2977 7680
rect 2915 7662 2989 7678
rect 3016 7674 3029 7688
rect 3044 7674 3060 7690
rect 3106 7685 3117 7698
rect 2899 7640 2900 7656
rect 2915 7640 2928 7662
rect 2943 7640 2973 7662
rect 3016 7658 3078 7674
rect 3106 7667 3117 7683
rect 3122 7678 3132 7698
rect 3142 7678 3156 7698
rect 3159 7685 3168 7698
rect 3184 7685 3193 7698
rect 3122 7667 3156 7678
rect 3159 7667 3168 7683
rect 3184 7667 3193 7683
rect 3200 7678 3210 7698
rect 3220 7678 3234 7698
rect 3235 7685 3246 7698
rect 3200 7667 3234 7678
rect 3235 7667 3246 7683
rect 3292 7674 3308 7690
rect 3315 7688 3345 7740
rect 3379 7736 3380 7743
rect 3364 7728 3380 7736
rect 3351 7696 3364 7715
rect 3379 7696 3409 7712
rect 3351 7680 3425 7696
rect 3351 7678 3364 7680
rect 3379 7678 3413 7680
rect 3016 7656 3029 7658
rect 3044 7656 3078 7658
rect 3016 7640 3078 7656
rect 3122 7651 3138 7654
rect 3200 7651 3230 7662
rect 3278 7658 3324 7674
rect 3351 7662 3425 7678
rect 3278 7656 3312 7658
rect 3277 7640 3324 7656
rect 3351 7640 3364 7662
rect 3379 7640 3409 7662
rect 3436 7640 3437 7656
rect 3452 7640 3465 7800
rect 3495 7696 3508 7800
rect 3553 7778 3554 7788
rect 3569 7778 3582 7788
rect 3553 7774 3582 7778
rect 3587 7774 3617 7800
rect 3635 7786 3651 7788
rect 3723 7786 3776 7800
rect 3724 7784 3788 7786
rect 3831 7784 3846 7800
rect 3895 7797 3925 7800
rect 3895 7794 3931 7797
rect 3861 7786 3877 7788
rect 3635 7774 3650 7778
rect 3553 7772 3650 7774
rect 3678 7772 3846 7784
rect 3862 7774 3877 7778
rect 3895 7775 3934 7794
rect 3953 7788 3960 7789
rect 3959 7781 3960 7788
rect 3943 7778 3944 7781
rect 3959 7778 3972 7781
rect 3895 7774 3925 7775
rect 3934 7774 3940 7775
rect 3943 7774 3972 7778
rect 3862 7773 3972 7774
rect 3862 7772 3978 7773
rect 3537 7764 3588 7772
rect 3537 7752 3562 7764
rect 3569 7752 3588 7764
rect 3619 7764 3669 7772
rect 3619 7756 3635 7764
rect 3642 7762 3669 7764
rect 3678 7762 3899 7772
rect 3642 7752 3899 7762
rect 3928 7764 3978 7772
rect 3928 7755 3944 7764
rect 3537 7744 3588 7752
rect 3635 7744 3899 7752
rect 3925 7752 3944 7755
rect 3951 7752 3978 7764
rect 3925 7744 3978 7752
rect 3553 7736 3554 7744
rect 3569 7736 3582 7744
rect 3553 7728 3569 7736
rect 3550 7721 3569 7724
rect 3550 7712 3572 7721
rect 3523 7702 3572 7712
rect 3523 7696 3553 7702
rect 3572 7697 3577 7702
rect 3495 7680 3569 7696
rect 3587 7688 3617 7744
rect 3652 7734 3860 7744
rect 3895 7740 3940 7744
rect 3943 7743 3944 7744
rect 3959 7743 3972 7744
rect 3678 7704 3867 7734
rect 3693 7701 3867 7704
rect 3686 7698 3867 7701
rect 3495 7678 3508 7680
rect 3523 7678 3557 7680
rect 3495 7662 3569 7678
rect 3596 7674 3609 7688
rect 3624 7674 3640 7690
rect 3686 7685 3697 7698
rect 3479 7640 3480 7656
rect 3495 7640 3508 7662
rect 3523 7640 3553 7662
rect 3596 7658 3658 7674
rect 3686 7667 3697 7683
rect 3702 7678 3712 7698
rect 3722 7678 3736 7698
rect 3739 7685 3748 7698
rect 3764 7685 3773 7698
rect 3702 7667 3736 7678
rect 3739 7667 3748 7683
rect 3764 7667 3773 7683
rect 3780 7678 3790 7698
rect 3800 7678 3814 7698
rect 3815 7685 3826 7698
rect 3780 7667 3814 7678
rect 3815 7667 3826 7683
rect 3872 7674 3888 7690
rect 3895 7688 3925 7740
rect 3959 7736 3960 7743
rect 3944 7728 3960 7736
rect 3931 7696 3944 7715
rect 3959 7696 3989 7712
rect 3931 7680 4005 7696
rect 3931 7678 3944 7680
rect 3959 7678 3993 7680
rect 3596 7656 3609 7658
rect 3624 7656 3658 7658
rect 3596 7640 3658 7656
rect 3702 7651 3718 7654
rect 3780 7651 3810 7662
rect 3858 7658 3904 7674
rect 3931 7662 4005 7678
rect 3858 7656 3892 7658
rect 3857 7640 3904 7656
rect 3931 7640 3944 7662
rect 3959 7640 3989 7662
rect 4016 7640 4017 7656
rect 4032 7640 4045 7800
rect 4075 7696 4088 7800
rect 4133 7778 4134 7788
rect 4149 7778 4162 7788
rect 4133 7774 4162 7778
rect 4167 7774 4197 7800
rect 4215 7786 4231 7788
rect 4303 7786 4356 7800
rect 4304 7784 4368 7786
rect 4411 7784 4426 7800
rect 4475 7797 4505 7800
rect 4475 7794 4511 7797
rect 4441 7786 4457 7788
rect 4215 7774 4230 7778
rect 4133 7772 4230 7774
rect 4258 7772 4426 7784
rect 4442 7774 4457 7778
rect 4475 7775 4514 7794
rect 4533 7788 4540 7789
rect 4539 7781 4540 7788
rect 4523 7778 4524 7781
rect 4539 7778 4552 7781
rect 4475 7774 4505 7775
rect 4514 7774 4520 7775
rect 4523 7774 4552 7778
rect 4442 7773 4552 7774
rect 4442 7772 4558 7773
rect 4117 7764 4168 7772
rect 4117 7752 4142 7764
rect 4149 7752 4168 7764
rect 4199 7764 4249 7772
rect 4199 7756 4215 7764
rect 4222 7762 4249 7764
rect 4258 7762 4479 7772
rect 4222 7752 4479 7762
rect 4508 7764 4558 7772
rect 4508 7755 4524 7764
rect 4117 7744 4168 7752
rect 4215 7744 4479 7752
rect 4505 7752 4524 7755
rect 4531 7752 4558 7764
rect 4505 7744 4558 7752
rect 4133 7736 4134 7744
rect 4149 7736 4162 7744
rect 4133 7728 4149 7736
rect 4130 7721 4149 7724
rect 4130 7712 4152 7721
rect 4103 7702 4152 7712
rect 4103 7696 4133 7702
rect 4152 7697 4157 7702
rect 4075 7680 4149 7696
rect 4167 7688 4197 7744
rect 4232 7734 4440 7744
rect 4475 7740 4520 7744
rect 4523 7743 4524 7744
rect 4539 7743 4552 7744
rect 4258 7704 4447 7734
rect 4273 7701 4447 7704
rect 4266 7698 4447 7701
rect 4075 7678 4088 7680
rect 4103 7678 4137 7680
rect 4075 7662 4149 7678
rect 4176 7674 4189 7688
rect 4204 7674 4220 7690
rect 4266 7685 4277 7698
rect 4059 7640 4060 7656
rect 4075 7640 4088 7662
rect 4103 7640 4133 7662
rect 4176 7658 4238 7674
rect 4266 7667 4277 7683
rect 4282 7678 4292 7698
rect 4302 7678 4316 7698
rect 4319 7685 4328 7698
rect 4344 7685 4353 7698
rect 4282 7667 4316 7678
rect 4319 7667 4328 7683
rect 4344 7667 4353 7683
rect 4360 7678 4370 7698
rect 4380 7678 4394 7698
rect 4395 7685 4406 7698
rect 4360 7667 4394 7678
rect 4395 7667 4406 7683
rect 4452 7674 4468 7690
rect 4475 7688 4505 7740
rect 4539 7736 4540 7743
rect 4524 7728 4540 7736
rect 4511 7696 4524 7715
rect 4539 7696 4569 7712
rect 4511 7680 4585 7696
rect 4511 7678 4524 7680
rect 4539 7678 4573 7680
rect 4176 7656 4189 7658
rect 4204 7656 4238 7658
rect 4176 7640 4238 7656
rect 4282 7651 4298 7654
rect 4360 7651 4390 7662
rect 4438 7658 4484 7674
rect 4511 7662 4585 7678
rect 4438 7656 4472 7658
rect 4437 7640 4484 7656
rect 4511 7640 4524 7662
rect 4539 7640 4569 7662
rect 4596 7640 4597 7656
rect 4612 7640 4625 7800
rect -7 7632 34 7640
rect -7 7606 8 7632
rect 15 7606 34 7632
rect 98 7628 160 7640
rect 172 7628 247 7640
rect 305 7628 380 7640
rect 392 7628 423 7640
rect 429 7628 464 7640
rect 98 7626 260 7628
rect -7 7598 34 7606
rect 116 7602 129 7626
rect 144 7624 159 7626
rect -1 7588 0 7598
rect 15 7588 28 7598
rect 43 7588 73 7602
rect 116 7588 159 7602
rect 183 7599 190 7606
rect 193 7602 260 7626
rect 292 7626 464 7628
rect 262 7604 290 7608
rect 292 7604 372 7626
rect 393 7624 408 7626
rect 262 7602 372 7604
rect 193 7598 372 7602
rect 166 7588 196 7598
rect 198 7588 351 7598
rect 359 7588 389 7598
rect 393 7588 423 7602
rect 451 7588 464 7626
rect 536 7632 571 7640
rect 536 7606 537 7632
rect 544 7606 571 7632
rect 479 7588 509 7602
rect 536 7598 571 7606
rect 573 7632 614 7640
rect 573 7606 588 7632
rect 595 7606 614 7632
rect 678 7628 740 7640
rect 752 7628 827 7640
rect 885 7628 960 7640
rect 972 7628 1003 7640
rect 1009 7628 1044 7640
rect 678 7626 840 7628
rect 573 7598 614 7606
rect 696 7602 709 7626
rect 724 7624 739 7626
rect 536 7588 537 7598
rect 552 7588 565 7598
rect 579 7588 580 7598
rect 595 7588 608 7598
rect 623 7588 653 7602
rect 696 7588 739 7602
rect 763 7599 770 7606
rect 773 7602 840 7626
rect 872 7626 1044 7628
rect 842 7604 870 7608
rect 872 7604 952 7626
rect 973 7624 988 7626
rect 842 7602 952 7604
rect 773 7598 952 7602
rect 746 7588 776 7598
rect 778 7588 931 7598
rect 939 7588 969 7598
rect 973 7588 1003 7602
rect 1031 7588 1044 7626
rect 1116 7632 1151 7640
rect 1116 7606 1117 7632
rect 1124 7606 1151 7632
rect 1059 7588 1089 7602
rect 1116 7598 1151 7606
rect 1153 7632 1194 7640
rect 1153 7606 1168 7632
rect 1175 7606 1194 7632
rect 1258 7628 1320 7640
rect 1332 7628 1407 7640
rect 1465 7628 1540 7640
rect 1552 7628 1583 7640
rect 1589 7628 1624 7640
rect 1258 7626 1420 7628
rect 1153 7598 1194 7606
rect 1276 7602 1289 7626
rect 1304 7624 1319 7626
rect 1116 7588 1117 7598
rect 1132 7588 1145 7598
rect 1159 7588 1160 7598
rect 1175 7588 1188 7598
rect 1203 7588 1233 7602
rect 1276 7588 1319 7602
rect 1343 7599 1350 7606
rect 1353 7602 1420 7626
rect 1452 7626 1624 7628
rect 1422 7604 1450 7608
rect 1452 7604 1532 7626
rect 1553 7624 1568 7626
rect 1422 7602 1532 7604
rect 1353 7598 1532 7602
rect 1326 7588 1356 7598
rect 1358 7588 1511 7598
rect 1519 7588 1549 7598
rect 1553 7588 1583 7602
rect 1611 7588 1624 7626
rect 1696 7632 1731 7640
rect 1696 7606 1697 7632
rect 1704 7606 1731 7632
rect 1639 7588 1669 7602
rect 1696 7598 1731 7606
rect 1733 7632 1774 7640
rect 1733 7606 1748 7632
rect 1755 7606 1774 7632
rect 1838 7628 1900 7640
rect 1912 7628 1987 7640
rect 2045 7628 2120 7640
rect 2132 7628 2163 7640
rect 2169 7628 2204 7640
rect 1838 7626 2000 7628
rect 1733 7598 1774 7606
rect 1856 7602 1869 7626
rect 1884 7624 1899 7626
rect 1696 7588 1697 7598
rect 1712 7588 1725 7598
rect 1739 7588 1740 7598
rect 1755 7588 1768 7598
rect 1783 7588 1813 7602
rect 1856 7588 1899 7602
rect 1923 7599 1930 7606
rect 1933 7602 2000 7626
rect 2032 7626 2204 7628
rect 2002 7604 2030 7608
rect 2032 7604 2112 7626
rect 2133 7624 2148 7626
rect 2002 7602 2112 7604
rect 1933 7598 2112 7602
rect 1906 7588 1936 7598
rect 1938 7588 2091 7598
rect 2099 7588 2129 7598
rect 2133 7588 2163 7602
rect 2191 7588 2204 7626
rect 2276 7632 2311 7640
rect 2276 7606 2277 7632
rect 2284 7606 2311 7632
rect 2219 7588 2249 7602
rect 2276 7598 2311 7606
rect 2313 7632 2354 7640
rect 2313 7606 2328 7632
rect 2335 7606 2354 7632
rect 2418 7628 2480 7640
rect 2492 7628 2567 7640
rect 2625 7628 2700 7640
rect 2712 7628 2743 7640
rect 2749 7628 2784 7640
rect 2418 7626 2580 7628
rect 2313 7598 2354 7606
rect 2436 7602 2449 7626
rect 2464 7624 2479 7626
rect 2276 7588 2277 7598
rect 2292 7588 2305 7598
rect 2319 7588 2320 7598
rect 2335 7588 2348 7598
rect 2363 7588 2393 7602
rect 2436 7588 2479 7602
rect 2503 7599 2510 7606
rect 2513 7602 2580 7626
rect 2612 7626 2784 7628
rect 2582 7604 2610 7608
rect 2612 7604 2692 7626
rect 2713 7624 2728 7626
rect 2582 7602 2692 7604
rect 2513 7598 2692 7602
rect 2486 7588 2516 7598
rect 2518 7588 2671 7598
rect 2679 7588 2709 7598
rect 2713 7588 2743 7602
rect 2771 7588 2784 7626
rect 2856 7632 2891 7640
rect 2856 7606 2857 7632
rect 2864 7606 2891 7632
rect 2799 7588 2829 7602
rect 2856 7598 2891 7606
rect 2893 7632 2934 7640
rect 2893 7606 2908 7632
rect 2915 7606 2934 7632
rect 2998 7628 3060 7640
rect 3072 7628 3147 7640
rect 3205 7628 3280 7640
rect 3292 7628 3323 7640
rect 3329 7628 3364 7640
rect 2998 7626 3160 7628
rect 2893 7598 2934 7606
rect 3016 7602 3029 7626
rect 3044 7624 3059 7626
rect 2856 7588 2857 7598
rect 2872 7588 2885 7598
rect 2899 7588 2900 7598
rect 2915 7588 2928 7598
rect 2943 7588 2973 7602
rect 3016 7588 3059 7602
rect 3083 7599 3090 7606
rect 3093 7602 3160 7626
rect 3192 7626 3364 7628
rect 3162 7604 3190 7608
rect 3192 7604 3272 7626
rect 3293 7624 3308 7626
rect 3162 7602 3272 7604
rect 3093 7598 3272 7602
rect 3066 7588 3096 7598
rect 3098 7588 3251 7598
rect 3259 7588 3289 7598
rect 3293 7588 3323 7602
rect 3351 7588 3364 7626
rect 3436 7632 3471 7640
rect 3436 7606 3437 7632
rect 3444 7606 3471 7632
rect 3379 7588 3409 7602
rect 3436 7598 3471 7606
rect 3473 7632 3514 7640
rect 3473 7606 3488 7632
rect 3495 7606 3514 7632
rect 3578 7628 3640 7640
rect 3652 7628 3727 7640
rect 3785 7628 3860 7640
rect 3872 7628 3903 7640
rect 3909 7628 3944 7640
rect 3578 7626 3740 7628
rect 3473 7598 3514 7606
rect 3596 7602 3609 7626
rect 3624 7624 3639 7626
rect 3436 7588 3437 7598
rect 3452 7588 3465 7598
rect 3479 7588 3480 7598
rect 3495 7588 3508 7598
rect 3523 7588 3553 7602
rect 3596 7588 3639 7602
rect 3663 7599 3670 7606
rect 3673 7602 3740 7626
rect 3772 7626 3944 7628
rect 3742 7604 3770 7608
rect 3772 7604 3852 7626
rect 3873 7624 3888 7626
rect 3742 7602 3852 7604
rect 3673 7598 3852 7602
rect 3646 7588 3676 7598
rect 3678 7588 3831 7598
rect 3839 7588 3869 7598
rect 3873 7588 3903 7602
rect 3931 7588 3944 7626
rect 4016 7632 4051 7640
rect 4016 7606 4017 7632
rect 4024 7606 4051 7632
rect 3959 7588 3989 7602
rect 4016 7598 4051 7606
rect 4053 7632 4094 7640
rect 4053 7606 4068 7632
rect 4075 7606 4094 7632
rect 4158 7628 4220 7640
rect 4232 7628 4307 7640
rect 4365 7628 4440 7640
rect 4452 7628 4483 7640
rect 4489 7628 4524 7640
rect 4158 7626 4320 7628
rect 4053 7598 4094 7606
rect 4176 7602 4189 7626
rect 4204 7624 4219 7626
rect 4016 7588 4017 7598
rect 4032 7588 4045 7598
rect 4059 7588 4060 7598
rect 4075 7588 4088 7598
rect 4103 7588 4133 7602
rect 4176 7588 4219 7602
rect 4243 7599 4250 7606
rect 4253 7602 4320 7626
rect 4352 7626 4524 7628
rect 4322 7604 4350 7608
rect 4352 7604 4432 7626
rect 4453 7624 4468 7626
rect 4322 7602 4432 7604
rect 4253 7598 4432 7602
rect 4226 7588 4256 7598
rect 4258 7588 4411 7598
rect 4419 7588 4449 7598
rect 4453 7588 4483 7602
rect 4511 7588 4524 7626
rect 4596 7632 4631 7640
rect 4596 7606 4597 7632
rect 4604 7606 4631 7632
rect 4539 7588 4569 7602
rect 4596 7598 4631 7606
rect 4596 7588 4597 7598
rect 4612 7588 4625 7598
rect -1 7582 4625 7588
rect 0 7574 4625 7582
rect 15 7544 28 7574
rect 43 7556 73 7574
rect 116 7560 130 7574
rect 166 7560 386 7574
rect 117 7558 130 7560
rect 83 7546 98 7558
rect 80 7544 102 7546
rect 107 7544 137 7558
rect 198 7556 351 7560
rect 180 7544 372 7556
rect 415 7544 445 7558
rect 451 7544 464 7574
rect 479 7556 509 7574
rect 552 7544 565 7574
rect 595 7544 608 7574
rect 623 7556 653 7574
rect 696 7560 710 7574
rect 746 7560 966 7574
rect 697 7558 710 7560
rect 663 7546 678 7558
rect 660 7544 682 7546
rect 687 7544 717 7558
rect 778 7556 931 7560
rect 760 7544 952 7556
rect 995 7544 1025 7558
rect 1031 7544 1044 7574
rect 1059 7556 1089 7574
rect 1132 7544 1145 7574
rect 1175 7544 1188 7574
rect 1203 7556 1233 7574
rect 1276 7560 1290 7574
rect 1326 7560 1546 7574
rect 1277 7558 1290 7560
rect 1243 7546 1258 7558
rect 1240 7544 1262 7546
rect 1267 7544 1297 7558
rect 1358 7556 1511 7560
rect 1340 7544 1532 7556
rect 1575 7544 1605 7558
rect 1611 7544 1624 7574
rect 1639 7556 1669 7574
rect 1712 7544 1725 7574
rect 1755 7544 1768 7574
rect 1783 7556 1813 7574
rect 1856 7560 1870 7574
rect 1906 7560 2126 7574
rect 1857 7558 1870 7560
rect 1823 7546 1838 7558
rect 1820 7544 1842 7546
rect 1847 7544 1877 7558
rect 1938 7556 2091 7560
rect 1920 7544 2112 7556
rect 2155 7544 2185 7558
rect 2191 7544 2204 7574
rect 2219 7556 2249 7574
rect 2292 7544 2305 7574
rect 2335 7544 2348 7574
rect 2363 7556 2393 7574
rect 2436 7560 2450 7574
rect 2486 7560 2706 7574
rect 2437 7558 2450 7560
rect 2403 7546 2418 7558
rect 2400 7544 2422 7546
rect 2427 7544 2457 7558
rect 2518 7556 2671 7560
rect 2500 7544 2692 7556
rect 2735 7544 2765 7558
rect 2771 7544 2784 7574
rect 2799 7556 2829 7574
rect 2872 7544 2885 7574
rect 2915 7544 2928 7574
rect 2943 7556 2973 7574
rect 3016 7560 3030 7574
rect 3066 7560 3286 7574
rect 3017 7558 3030 7560
rect 2983 7546 2998 7558
rect 2980 7544 3002 7546
rect 3007 7544 3037 7558
rect 3098 7556 3251 7560
rect 3080 7544 3272 7556
rect 3315 7544 3345 7558
rect 3351 7544 3364 7574
rect 3379 7556 3409 7574
rect 3452 7544 3465 7574
rect 3495 7544 3508 7574
rect 3523 7556 3553 7574
rect 3596 7560 3610 7574
rect 3646 7560 3866 7574
rect 3597 7558 3610 7560
rect 3563 7546 3578 7558
rect 3560 7544 3582 7546
rect 3587 7544 3617 7558
rect 3678 7556 3831 7560
rect 3660 7544 3852 7556
rect 3895 7544 3925 7558
rect 3931 7544 3944 7574
rect 3959 7556 3989 7574
rect 4032 7544 4045 7574
rect 4075 7544 4088 7574
rect 4103 7556 4133 7574
rect 4176 7560 4190 7574
rect 4226 7560 4446 7574
rect 4177 7558 4190 7560
rect 4143 7546 4158 7558
rect 4140 7544 4162 7546
rect 4167 7544 4197 7558
rect 4258 7556 4411 7560
rect 4240 7544 4432 7556
rect 4475 7544 4505 7558
rect 4511 7544 4524 7574
rect 4539 7556 4569 7574
rect 4612 7544 4625 7574
rect 0 7530 4625 7544
rect 15 7426 28 7530
rect 73 7508 74 7518
rect 89 7508 102 7518
rect 73 7504 102 7508
rect 107 7504 137 7530
rect 155 7516 171 7518
rect 243 7516 296 7530
rect 244 7514 308 7516
rect 351 7514 366 7530
rect 415 7527 445 7530
rect 415 7524 451 7527
rect 381 7516 397 7518
rect 155 7504 170 7508
rect 73 7502 170 7504
rect 198 7502 366 7514
rect 382 7504 397 7508
rect 415 7505 454 7524
rect 473 7518 480 7519
rect 479 7511 480 7518
rect 463 7508 464 7511
rect 479 7508 492 7511
rect 415 7504 445 7505
rect 454 7504 460 7505
rect 463 7504 492 7508
rect 382 7503 492 7504
rect 382 7502 498 7503
rect 57 7494 108 7502
rect 57 7482 82 7494
rect 89 7482 108 7494
rect 139 7494 189 7502
rect 139 7486 155 7494
rect 162 7492 189 7494
rect 198 7492 419 7502
rect 162 7482 419 7492
rect 448 7494 498 7502
rect 448 7485 464 7494
rect 57 7474 108 7482
rect 155 7474 419 7482
rect 445 7482 464 7485
rect 471 7482 498 7494
rect 445 7474 498 7482
rect 73 7466 74 7474
rect 89 7466 102 7474
rect 73 7458 89 7466
rect 70 7451 89 7454
rect 70 7442 92 7451
rect 43 7432 92 7442
rect 43 7426 73 7432
rect 92 7427 97 7432
rect 15 7410 89 7426
rect 107 7418 137 7474
rect 172 7464 380 7474
rect 415 7470 460 7474
rect 463 7473 464 7474
rect 479 7473 492 7474
rect 198 7434 387 7464
rect 213 7431 387 7434
rect 206 7428 387 7431
rect 15 7408 28 7410
rect 43 7408 77 7410
rect 15 7392 89 7408
rect 116 7404 129 7418
rect 144 7404 160 7420
rect 206 7415 217 7428
rect -1 7370 0 7386
rect 15 7370 28 7392
rect 43 7370 73 7392
rect 116 7388 178 7404
rect 206 7397 217 7413
rect 222 7408 232 7428
rect 242 7408 256 7428
rect 259 7415 268 7428
rect 284 7415 293 7428
rect 222 7397 256 7408
rect 259 7397 268 7413
rect 284 7397 293 7413
rect 300 7408 310 7428
rect 320 7408 334 7428
rect 335 7415 346 7428
rect 300 7397 334 7408
rect 335 7397 346 7413
rect 392 7404 408 7420
rect 415 7418 445 7470
rect 479 7466 480 7473
rect 464 7458 480 7466
rect 451 7426 464 7445
rect 479 7426 509 7442
rect 451 7410 525 7426
rect 451 7408 464 7410
rect 479 7408 513 7410
rect 116 7386 129 7388
rect 144 7386 178 7388
rect 116 7370 178 7386
rect 222 7381 238 7384
rect 300 7381 330 7392
rect 378 7388 424 7404
rect 451 7392 525 7408
rect 378 7386 412 7388
rect 377 7370 424 7386
rect 451 7370 464 7392
rect 479 7370 509 7392
rect 536 7370 537 7386
rect 552 7370 565 7530
rect 595 7426 608 7530
rect 653 7508 654 7518
rect 669 7508 682 7518
rect 653 7504 682 7508
rect 687 7504 717 7530
rect 735 7516 751 7518
rect 823 7516 876 7530
rect 824 7514 888 7516
rect 931 7514 946 7530
rect 995 7527 1025 7530
rect 995 7524 1031 7527
rect 961 7516 977 7518
rect 735 7504 750 7508
rect 653 7502 750 7504
rect 778 7502 946 7514
rect 962 7504 977 7508
rect 995 7505 1034 7524
rect 1053 7518 1060 7519
rect 1059 7511 1060 7518
rect 1043 7508 1044 7511
rect 1059 7508 1072 7511
rect 995 7504 1025 7505
rect 1034 7504 1040 7505
rect 1043 7504 1072 7508
rect 962 7503 1072 7504
rect 962 7502 1078 7503
rect 637 7494 688 7502
rect 637 7482 662 7494
rect 669 7482 688 7494
rect 719 7494 769 7502
rect 719 7486 735 7494
rect 742 7492 769 7494
rect 778 7492 999 7502
rect 742 7482 999 7492
rect 1028 7494 1078 7502
rect 1028 7485 1044 7494
rect 637 7474 688 7482
rect 735 7474 999 7482
rect 1025 7482 1044 7485
rect 1051 7482 1078 7494
rect 1025 7474 1078 7482
rect 653 7466 654 7474
rect 669 7466 682 7474
rect 653 7458 669 7466
rect 650 7451 669 7454
rect 650 7442 672 7451
rect 623 7432 672 7442
rect 623 7426 653 7432
rect 672 7427 677 7432
rect 595 7410 669 7426
rect 687 7418 717 7474
rect 752 7464 960 7474
rect 995 7470 1040 7474
rect 1043 7473 1044 7474
rect 1059 7473 1072 7474
rect 778 7434 967 7464
rect 793 7431 967 7434
rect 786 7428 967 7431
rect 595 7408 608 7410
rect 623 7408 657 7410
rect 595 7392 669 7408
rect 696 7404 709 7418
rect 724 7404 740 7420
rect 786 7415 797 7428
rect 579 7370 580 7386
rect 595 7370 608 7392
rect 623 7370 653 7392
rect 696 7388 758 7404
rect 786 7397 797 7413
rect 802 7408 812 7428
rect 822 7408 836 7428
rect 839 7415 848 7428
rect 864 7415 873 7428
rect 802 7397 836 7408
rect 839 7397 848 7413
rect 864 7397 873 7413
rect 880 7408 890 7428
rect 900 7408 914 7428
rect 915 7415 926 7428
rect 880 7397 914 7408
rect 915 7397 926 7413
rect 972 7404 988 7420
rect 995 7418 1025 7470
rect 1059 7466 1060 7473
rect 1044 7458 1060 7466
rect 1031 7426 1044 7445
rect 1059 7426 1089 7442
rect 1031 7410 1105 7426
rect 1031 7408 1044 7410
rect 1059 7408 1093 7410
rect 696 7386 709 7388
rect 724 7386 758 7388
rect 696 7370 758 7386
rect 802 7381 818 7384
rect 880 7381 910 7392
rect 958 7388 1004 7404
rect 1031 7392 1105 7408
rect 958 7386 992 7388
rect 957 7370 1004 7386
rect 1031 7370 1044 7392
rect 1059 7370 1089 7392
rect 1116 7370 1117 7386
rect 1132 7370 1145 7530
rect 1175 7426 1188 7530
rect 1233 7508 1234 7518
rect 1249 7508 1262 7518
rect 1233 7504 1262 7508
rect 1267 7504 1297 7530
rect 1315 7516 1331 7518
rect 1403 7516 1456 7530
rect 1404 7514 1468 7516
rect 1511 7514 1526 7530
rect 1575 7527 1605 7530
rect 1575 7524 1611 7527
rect 1541 7516 1557 7518
rect 1315 7504 1330 7508
rect 1233 7502 1330 7504
rect 1358 7502 1526 7514
rect 1542 7504 1557 7508
rect 1575 7505 1614 7524
rect 1633 7518 1640 7519
rect 1639 7511 1640 7518
rect 1623 7508 1624 7511
rect 1639 7508 1652 7511
rect 1575 7504 1605 7505
rect 1614 7504 1620 7505
rect 1623 7504 1652 7508
rect 1542 7503 1652 7504
rect 1542 7502 1658 7503
rect 1217 7494 1268 7502
rect 1217 7482 1242 7494
rect 1249 7482 1268 7494
rect 1299 7494 1349 7502
rect 1299 7486 1315 7494
rect 1322 7492 1349 7494
rect 1358 7492 1579 7502
rect 1322 7482 1579 7492
rect 1608 7494 1658 7502
rect 1608 7485 1624 7494
rect 1217 7474 1268 7482
rect 1315 7474 1579 7482
rect 1605 7482 1624 7485
rect 1631 7482 1658 7494
rect 1605 7474 1658 7482
rect 1233 7466 1234 7474
rect 1249 7466 1262 7474
rect 1233 7458 1249 7466
rect 1230 7451 1249 7454
rect 1230 7442 1252 7451
rect 1203 7432 1252 7442
rect 1203 7426 1233 7432
rect 1252 7427 1257 7432
rect 1175 7410 1249 7426
rect 1267 7418 1297 7474
rect 1332 7464 1540 7474
rect 1575 7470 1620 7474
rect 1623 7473 1624 7474
rect 1639 7473 1652 7474
rect 1358 7434 1547 7464
rect 1373 7431 1547 7434
rect 1366 7428 1547 7431
rect 1175 7408 1188 7410
rect 1203 7408 1237 7410
rect 1175 7392 1249 7408
rect 1276 7404 1289 7418
rect 1304 7404 1320 7420
rect 1366 7415 1377 7428
rect 1159 7370 1160 7386
rect 1175 7370 1188 7392
rect 1203 7370 1233 7392
rect 1276 7388 1338 7404
rect 1366 7397 1377 7413
rect 1382 7408 1392 7428
rect 1402 7408 1416 7428
rect 1419 7415 1428 7428
rect 1444 7415 1453 7428
rect 1382 7397 1416 7408
rect 1419 7397 1428 7413
rect 1444 7397 1453 7413
rect 1460 7408 1470 7428
rect 1480 7408 1494 7428
rect 1495 7415 1506 7428
rect 1460 7397 1494 7408
rect 1495 7397 1506 7413
rect 1552 7404 1568 7420
rect 1575 7418 1605 7470
rect 1639 7466 1640 7473
rect 1624 7458 1640 7466
rect 1611 7426 1624 7445
rect 1639 7426 1669 7442
rect 1611 7410 1685 7426
rect 1611 7408 1624 7410
rect 1639 7408 1673 7410
rect 1276 7386 1289 7388
rect 1304 7386 1338 7388
rect 1276 7370 1338 7386
rect 1382 7381 1398 7384
rect 1460 7381 1490 7392
rect 1538 7388 1584 7404
rect 1611 7392 1685 7408
rect 1538 7386 1572 7388
rect 1537 7370 1584 7386
rect 1611 7370 1624 7392
rect 1639 7370 1669 7392
rect 1696 7370 1697 7386
rect 1712 7370 1725 7530
rect 1755 7426 1768 7530
rect 1813 7508 1814 7518
rect 1829 7508 1842 7518
rect 1813 7504 1842 7508
rect 1847 7504 1877 7530
rect 1895 7516 1911 7518
rect 1983 7516 2036 7530
rect 1984 7514 2048 7516
rect 2091 7514 2106 7530
rect 2155 7527 2185 7530
rect 2155 7524 2191 7527
rect 2121 7516 2137 7518
rect 1895 7504 1910 7508
rect 1813 7502 1910 7504
rect 1938 7502 2106 7514
rect 2122 7504 2137 7508
rect 2155 7505 2194 7524
rect 2213 7518 2220 7519
rect 2219 7511 2220 7518
rect 2203 7508 2204 7511
rect 2219 7508 2232 7511
rect 2155 7504 2185 7505
rect 2194 7504 2200 7505
rect 2203 7504 2232 7508
rect 2122 7503 2232 7504
rect 2122 7502 2238 7503
rect 1797 7494 1848 7502
rect 1797 7482 1822 7494
rect 1829 7482 1848 7494
rect 1879 7494 1929 7502
rect 1879 7486 1895 7494
rect 1902 7492 1929 7494
rect 1938 7492 2159 7502
rect 1902 7482 2159 7492
rect 2188 7494 2238 7502
rect 2188 7485 2204 7494
rect 1797 7474 1848 7482
rect 1895 7474 2159 7482
rect 2185 7482 2204 7485
rect 2211 7482 2238 7494
rect 2185 7474 2238 7482
rect 1813 7466 1814 7474
rect 1829 7466 1842 7474
rect 1813 7458 1829 7466
rect 1810 7451 1829 7454
rect 1810 7442 1832 7451
rect 1783 7432 1832 7442
rect 1783 7426 1813 7432
rect 1832 7427 1837 7432
rect 1755 7410 1829 7426
rect 1847 7418 1877 7474
rect 1912 7464 2120 7474
rect 2155 7470 2200 7474
rect 2203 7473 2204 7474
rect 2219 7473 2232 7474
rect 1938 7434 2127 7464
rect 1953 7431 2127 7434
rect 1946 7428 2127 7431
rect 1755 7408 1768 7410
rect 1783 7408 1817 7410
rect 1755 7392 1829 7408
rect 1856 7404 1869 7418
rect 1884 7404 1900 7420
rect 1946 7415 1957 7428
rect 1739 7370 1740 7386
rect 1755 7370 1768 7392
rect 1783 7370 1813 7392
rect 1856 7388 1918 7404
rect 1946 7397 1957 7413
rect 1962 7408 1972 7428
rect 1982 7408 1996 7428
rect 1999 7415 2008 7428
rect 2024 7415 2033 7428
rect 1962 7397 1996 7408
rect 1999 7397 2008 7413
rect 2024 7397 2033 7413
rect 2040 7408 2050 7428
rect 2060 7408 2074 7428
rect 2075 7415 2086 7428
rect 2040 7397 2074 7408
rect 2075 7397 2086 7413
rect 2132 7404 2148 7420
rect 2155 7418 2185 7470
rect 2219 7466 2220 7473
rect 2204 7458 2220 7466
rect 2191 7426 2204 7445
rect 2219 7426 2249 7442
rect 2191 7410 2265 7426
rect 2191 7408 2204 7410
rect 2219 7408 2253 7410
rect 1856 7386 1869 7388
rect 1884 7386 1918 7388
rect 1856 7370 1918 7386
rect 1962 7381 1978 7384
rect 2040 7381 2070 7392
rect 2118 7388 2164 7404
rect 2191 7392 2265 7408
rect 2118 7386 2152 7388
rect 2117 7370 2164 7386
rect 2191 7370 2204 7392
rect 2219 7370 2249 7392
rect 2276 7370 2277 7386
rect 2292 7370 2305 7530
rect 2335 7426 2348 7530
rect 2393 7508 2394 7518
rect 2409 7508 2422 7518
rect 2393 7504 2422 7508
rect 2427 7504 2457 7530
rect 2475 7516 2491 7518
rect 2563 7516 2616 7530
rect 2564 7514 2628 7516
rect 2671 7514 2686 7530
rect 2735 7527 2765 7530
rect 2735 7524 2771 7527
rect 2701 7516 2717 7518
rect 2475 7504 2490 7508
rect 2393 7502 2490 7504
rect 2518 7502 2686 7514
rect 2702 7504 2717 7508
rect 2735 7505 2774 7524
rect 2793 7518 2800 7519
rect 2799 7511 2800 7518
rect 2783 7508 2784 7511
rect 2799 7508 2812 7511
rect 2735 7504 2765 7505
rect 2774 7504 2780 7505
rect 2783 7504 2812 7508
rect 2702 7503 2812 7504
rect 2702 7502 2818 7503
rect 2377 7494 2428 7502
rect 2377 7482 2402 7494
rect 2409 7482 2428 7494
rect 2459 7494 2509 7502
rect 2459 7486 2475 7494
rect 2482 7492 2509 7494
rect 2518 7492 2739 7502
rect 2482 7482 2739 7492
rect 2768 7494 2818 7502
rect 2768 7485 2784 7494
rect 2377 7474 2428 7482
rect 2475 7474 2739 7482
rect 2765 7482 2784 7485
rect 2791 7482 2818 7494
rect 2765 7474 2818 7482
rect 2393 7466 2394 7474
rect 2409 7466 2422 7474
rect 2393 7458 2409 7466
rect 2390 7451 2409 7454
rect 2390 7442 2412 7451
rect 2363 7432 2412 7442
rect 2363 7426 2393 7432
rect 2412 7427 2417 7432
rect 2335 7410 2409 7426
rect 2427 7418 2457 7474
rect 2492 7464 2700 7474
rect 2735 7470 2780 7474
rect 2783 7473 2784 7474
rect 2799 7473 2812 7474
rect 2518 7434 2707 7464
rect 2533 7431 2707 7434
rect 2526 7428 2707 7431
rect 2335 7408 2348 7410
rect 2363 7408 2397 7410
rect 2335 7392 2409 7408
rect 2436 7404 2449 7418
rect 2464 7404 2480 7420
rect 2526 7415 2537 7428
rect 2319 7370 2320 7386
rect 2335 7370 2348 7392
rect 2363 7370 2393 7392
rect 2436 7388 2498 7404
rect 2526 7397 2537 7413
rect 2542 7408 2552 7428
rect 2562 7408 2576 7428
rect 2579 7415 2588 7428
rect 2604 7415 2613 7428
rect 2542 7397 2576 7408
rect 2579 7397 2588 7413
rect 2604 7397 2613 7413
rect 2620 7408 2630 7428
rect 2640 7408 2654 7428
rect 2655 7415 2666 7428
rect 2620 7397 2654 7408
rect 2655 7397 2666 7413
rect 2712 7404 2728 7420
rect 2735 7418 2765 7470
rect 2799 7466 2800 7473
rect 2784 7458 2800 7466
rect 2771 7426 2784 7445
rect 2799 7426 2829 7442
rect 2771 7410 2845 7426
rect 2771 7408 2784 7410
rect 2799 7408 2833 7410
rect 2436 7386 2449 7388
rect 2464 7386 2498 7388
rect 2436 7370 2498 7386
rect 2542 7381 2558 7384
rect 2620 7381 2650 7392
rect 2698 7388 2744 7404
rect 2771 7392 2845 7408
rect 2698 7386 2732 7388
rect 2697 7370 2744 7386
rect 2771 7370 2784 7392
rect 2799 7370 2829 7392
rect 2856 7370 2857 7386
rect 2872 7370 2885 7530
rect 2915 7426 2928 7530
rect 2973 7508 2974 7518
rect 2989 7508 3002 7518
rect 2973 7504 3002 7508
rect 3007 7504 3037 7530
rect 3055 7516 3071 7518
rect 3143 7516 3196 7530
rect 3144 7514 3208 7516
rect 3251 7514 3266 7530
rect 3315 7527 3345 7530
rect 3315 7524 3351 7527
rect 3281 7516 3297 7518
rect 3055 7504 3070 7508
rect 2973 7502 3070 7504
rect 3098 7502 3266 7514
rect 3282 7504 3297 7508
rect 3315 7505 3354 7524
rect 3373 7518 3380 7519
rect 3379 7511 3380 7518
rect 3363 7508 3364 7511
rect 3379 7508 3392 7511
rect 3315 7504 3345 7505
rect 3354 7504 3360 7505
rect 3363 7504 3392 7508
rect 3282 7503 3392 7504
rect 3282 7502 3398 7503
rect 2957 7494 3008 7502
rect 2957 7482 2982 7494
rect 2989 7482 3008 7494
rect 3039 7494 3089 7502
rect 3039 7486 3055 7494
rect 3062 7492 3089 7494
rect 3098 7492 3319 7502
rect 3062 7482 3319 7492
rect 3348 7494 3398 7502
rect 3348 7485 3364 7494
rect 2957 7474 3008 7482
rect 3055 7474 3319 7482
rect 3345 7482 3364 7485
rect 3371 7482 3398 7494
rect 3345 7474 3398 7482
rect 2973 7466 2974 7474
rect 2989 7466 3002 7474
rect 2973 7458 2989 7466
rect 2970 7451 2989 7454
rect 2970 7442 2992 7451
rect 2943 7432 2992 7442
rect 2943 7426 2973 7432
rect 2992 7427 2997 7432
rect 2915 7410 2989 7426
rect 3007 7418 3037 7474
rect 3072 7464 3280 7474
rect 3315 7470 3360 7474
rect 3363 7473 3364 7474
rect 3379 7473 3392 7474
rect 3098 7434 3287 7464
rect 3113 7431 3287 7434
rect 3106 7428 3287 7431
rect 2915 7408 2928 7410
rect 2943 7408 2977 7410
rect 2915 7392 2989 7408
rect 3016 7404 3029 7418
rect 3044 7404 3060 7420
rect 3106 7415 3117 7428
rect 2899 7370 2900 7386
rect 2915 7370 2928 7392
rect 2943 7370 2973 7392
rect 3016 7388 3078 7404
rect 3106 7397 3117 7413
rect 3122 7408 3132 7428
rect 3142 7408 3156 7428
rect 3159 7415 3168 7428
rect 3184 7415 3193 7428
rect 3122 7397 3156 7408
rect 3159 7397 3168 7413
rect 3184 7397 3193 7413
rect 3200 7408 3210 7428
rect 3220 7408 3234 7428
rect 3235 7415 3246 7428
rect 3200 7397 3234 7408
rect 3235 7397 3246 7413
rect 3292 7404 3308 7420
rect 3315 7418 3345 7470
rect 3379 7466 3380 7473
rect 3364 7458 3380 7466
rect 3351 7426 3364 7445
rect 3379 7426 3409 7442
rect 3351 7410 3425 7426
rect 3351 7408 3364 7410
rect 3379 7408 3413 7410
rect 3016 7386 3029 7388
rect 3044 7386 3078 7388
rect 3016 7370 3078 7386
rect 3122 7381 3138 7384
rect 3200 7381 3230 7392
rect 3278 7388 3324 7404
rect 3351 7392 3425 7408
rect 3278 7386 3312 7388
rect 3277 7370 3324 7386
rect 3351 7370 3364 7392
rect 3379 7370 3409 7392
rect 3436 7370 3437 7386
rect 3452 7370 3465 7530
rect 3495 7426 3508 7530
rect 3553 7508 3554 7518
rect 3569 7508 3582 7518
rect 3553 7504 3582 7508
rect 3587 7504 3617 7530
rect 3635 7516 3651 7518
rect 3723 7516 3776 7530
rect 3724 7514 3788 7516
rect 3831 7514 3846 7530
rect 3895 7527 3925 7530
rect 3895 7524 3931 7527
rect 3861 7516 3877 7518
rect 3635 7504 3650 7508
rect 3553 7502 3650 7504
rect 3678 7502 3846 7514
rect 3862 7504 3877 7508
rect 3895 7505 3934 7524
rect 3953 7518 3960 7519
rect 3959 7511 3960 7518
rect 3943 7508 3944 7511
rect 3959 7508 3972 7511
rect 3895 7504 3925 7505
rect 3934 7504 3940 7505
rect 3943 7504 3972 7508
rect 3862 7503 3972 7504
rect 3862 7502 3978 7503
rect 3537 7494 3588 7502
rect 3537 7482 3562 7494
rect 3569 7482 3588 7494
rect 3619 7494 3669 7502
rect 3619 7486 3635 7494
rect 3642 7492 3669 7494
rect 3678 7492 3899 7502
rect 3642 7482 3899 7492
rect 3928 7494 3978 7502
rect 3928 7485 3944 7494
rect 3537 7474 3588 7482
rect 3635 7474 3899 7482
rect 3925 7482 3944 7485
rect 3951 7482 3978 7494
rect 3925 7474 3978 7482
rect 3553 7466 3554 7474
rect 3569 7466 3582 7474
rect 3553 7458 3569 7466
rect 3550 7451 3569 7454
rect 3550 7442 3572 7451
rect 3523 7432 3572 7442
rect 3523 7426 3553 7432
rect 3572 7427 3577 7432
rect 3495 7410 3569 7426
rect 3587 7418 3617 7474
rect 3652 7464 3860 7474
rect 3895 7470 3940 7474
rect 3943 7473 3944 7474
rect 3959 7473 3972 7474
rect 3678 7434 3867 7464
rect 3693 7431 3867 7434
rect 3686 7428 3867 7431
rect 3495 7408 3508 7410
rect 3523 7408 3557 7410
rect 3495 7392 3569 7408
rect 3596 7404 3609 7418
rect 3624 7404 3640 7420
rect 3686 7415 3697 7428
rect 3479 7370 3480 7386
rect 3495 7370 3508 7392
rect 3523 7370 3553 7392
rect 3596 7388 3658 7404
rect 3686 7397 3697 7413
rect 3702 7408 3712 7428
rect 3722 7408 3736 7428
rect 3739 7415 3748 7428
rect 3764 7415 3773 7428
rect 3702 7397 3736 7408
rect 3739 7397 3748 7413
rect 3764 7397 3773 7413
rect 3780 7408 3790 7428
rect 3800 7408 3814 7428
rect 3815 7415 3826 7428
rect 3780 7397 3814 7408
rect 3815 7397 3826 7413
rect 3872 7404 3888 7420
rect 3895 7418 3925 7470
rect 3959 7466 3960 7473
rect 3944 7458 3960 7466
rect 3931 7426 3944 7445
rect 3959 7426 3989 7442
rect 3931 7410 4005 7426
rect 3931 7408 3944 7410
rect 3959 7408 3993 7410
rect 3596 7386 3609 7388
rect 3624 7386 3658 7388
rect 3596 7370 3658 7386
rect 3702 7381 3718 7384
rect 3780 7381 3810 7392
rect 3858 7388 3904 7404
rect 3931 7392 4005 7408
rect 3858 7386 3892 7388
rect 3857 7370 3904 7386
rect 3931 7370 3944 7392
rect 3959 7370 3989 7392
rect 4016 7370 4017 7386
rect 4032 7370 4045 7530
rect 4075 7426 4088 7530
rect 4133 7508 4134 7518
rect 4149 7508 4162 7518
rect 4133 7504 4162 7508
rect 4167 7504 4197 7530
rect 4215 7516 4231 7518
rect 4303 7516 4356 7530
rect 4304 7514 4368 7516
rect 4411 7514 4426 7530
rect 4475 7527 4505 7530
rect 4475 7524 4511 7527
rect 4441 7516 4457 7518
rect 4215 7504 4230 7508
rect 4133 7502 4230 7504
rect 4258 7502 4426 7514
rect 4442 7504 4457 7508
rect 4475 7505 4514 7524
rect 4533 7518 4540 7519
rect 4539 7511 4540 7518
rect 4523 7508 4524 7511
rect 4539 7508 4552 7511
rect 4475 7504 4505 7505
rect 4514 7504 4520 7505
rect 4523 7504 4552 7508
rect 4442 7503 4552 7504
rect 4442 7502 4558 7503
rect 4117 7494 4168 7502
rect 4117 7482 4142 7494
rect 4149 7482 4168 7494
rect 4199 7494 4249 7502
rect 4199 7486 4215 7494
rect 4222 7492 4249 7494
rect 4258 7492 4479 7502
rect 4222 7482 4479 7492
rect 4508 7494 4558 7502
rect 4508 7485 4524 7494
rect 4117 7474 4168 7482
rect 4215 7474 4479 7482
rect 4505 7482 4524 7485
rect 4531 7482 4558 7494
rect 4505 7474 4558 7482
rect 4133 7466 4134 7474
rect 4149 7466 4162 7474
rect 4133 7458 4149 7466
rect 4130 7451 4149 7454
rect 4130 7442 4152 7451
rect 4103 7432 4152 7442
rect 4103 7426 4133 7432
rect 4152 7427 4157 7432
rect 4075 7410 4149 7426
rect 4167 7418 4197 7474
rect 4232 7464 4440 7474
rect 4475 7470 4520 7474
rect 4523 7473 4524 7474
rect 4539 7473 4552 7474
rect 4258 7434 4447 7464
rect 4273 7431 4447 7434
rect 4266 7428 4447 7431
rect 4075 7408 4088 7410
rect 4103 7408 4137 7410
rect 4075 7392 4149 7408
rect 4176 7404 4189 7418
rect 4204 7404 4220 7420
rect 4266 7415 4277 7428
rect 4059 7370 4060 7386
rect 4075 7370 4088 7392
rect 4103 7370 4133 7392
rect 4176 7388 4238 7404
rect 4266 7397 4277 7413
rect 4282 7408 4292 7428
rect 4302 7408 4316 7428
rect 4319 7415 4328 7428
rect 4344 7415 4353 7428
rect 4282 7397 4316 7408
rect 4319 7397 4328 7413
rect 4344 7397 4353 7413
rect 4360 7408 4370 7428
rect 4380 7408 4394 7428
rect 4395 7415 4406 7428
rect 4360 7397 4394 7408
rect 4395 7397 4406 7413
rect 4452 7404 4468 7420
rect 4475 7418 4505 7470
rect 4539 7466 4540 7473
rect 4524 7458 4540 7466
rect 4511 7426 4524 7445
rect 4539 7426 4569 7442
rect 4511 7410 4585 7426
rect 4511 7408 4524 7410
rect 4539 7408 4573 7410
rect 4176 7386 4189 7388
rect 4204 7386 4238 7388
rect 4176 7370 4238 7386
rect 4282 7381 4298 7384
rect 4360 7381 4390 7392
rect 4438 7388 4484 7404
rect 4511 7392 4585 7408
rect 4438 7386 4472 7388
rect 4437 7370 4484 7386
rect 4511 7370 4524 7392
rect 4539 7370 4569 7392
rect 4596 7370 4597 7386
rect 4612 7370 4625 7530
rect -7 7362 34 7370
rect -7 7336 8 7362
rect 15 7336 34 7362
rect 98 7358 160 7370
rect 172 7358 247 7370
rect 305 7358 380 7370
rect 392 7358 423 7370
rect 429 7358 464 7370
rect 98 7356 260 7358
rect -7 7328 34 7336
rect 116 7332 129 7356
rect 144 7354 159 7356
rect -1 7318 0 7328
rect 15 7318 28 7328
rect 43 7318 73 7332
rect 116 7318 159 7332
rect 183 7329 190 7336
rect 193 7332 260 7356
rect 292 7356 464 7358
rect 262 7334 290 7338
rect 292 7334 372 7356
rect 393 7354 408 7356
rect 262 7332 372 7334
rect 193 7328 372 7332
rect 166 7318 196 7328
rect 198 7318 351 7328
rect 359 7318 389 7328
rect 393 7318 423 7332
rect 451 7318 464 7356
rect 536 7362 571 7370
rect 536 7336 537 7362
rect 544 7336 571 7362
rect 479 7318 509 7332
rect 536 7328 571 7336
rect 573 7362 614 7370
rect 573 7336 588 7362
rect 595 7336 614 7362
rect 678 7358 740 7370
rect 752 7358 827 7370
rect 885 7358 960 7370
rect 972 7358 1003 7370
rect 1009 7358 1044 7370
rect 678 7356 840 7358
rect 573 7328 614 7336
rect 696 7332 709 7356
rect 724 7354 739 7356
rect 536 7318 537 7328
rect 552 7318 565 7328
rect 579 7318 580 7328
rect 595 7318 608 7328
rect 623 7318 653 7332
rect 696 7318 739 7332
rect 763 7329 770 7336
rect 773 7332 840 7356
rect 872 7356 1044 7358
rect 842 7334 870 7338
rect 872 7334 952 7356
rect 973 7354 988 7356
rect 842 7332 952 7334
rect 773 7328 952 7332
rect 746 7318 776 7328
rect 778 7318 931 7328
rect 939 7318 969 7328
rect 973 7318 1003 7332
rect 1031 7318 1044 7356
rect 1116 7362 1151 7370
rect 1116 7336 1117 7362
rect 1124 7336 1151 7362
rect 1059 7318 1089 7332
rect 1116 7328 1151 7336
rect 1153 7362 1194 7370
rect 1153 7336 1168 7362
rect 1175 7336 1194 7362
rect 1258 7358 1320 7370
rect 1332 7358 1407 7370
rect 1465 7358 1540 7370
rect 1552 7358 1583 7370
rect 1589 7358 1624 7370
rect 1258 7356 1420 7358
rect 1153 7328 1194 7336
rect 1276 7332 1289 7356
rect 1304 7354 1319 7356
rect 1116 7318 1117 7328
rect 1132 7318 1145 7328
rect 1159 7318 1160 7328
rect 1175 7318 1188 7328
rect 1203 7318 1233 7332
rect 1276 7318 1319 7332
rect 1343 7329 1350 7336
rect 1353 7332 1420 7356
rect 1452 7356 1624 7358
rect 1422 7334 1450 7338
rect 1452 7334 1532 7356
rect 1553 7354 1568 7356
rect 1422 7332 1532 7334
rect 1353 7328 1532 7332
rect 1326 7318 1356 7328
rect 1358 7318 1511 7328
rect 1519 7318 1549 7328
rect 1553 7318 1583 7332
rect 1611 7318 1624 7356
rect 1696 7362 1731 7370
rect 1696 7336 1697 7362
rect 1704 7336 1731 7362
rect 1639 7318 1669 7332
rect 1696 7328 1731 7336
rect 1733 7362 1774 7370
rect 1733 7336 1748 7362
rect 1755 7336 1774 7362
rect 1838 7358 1900 7370
rect 1912 7358 1987 7370
rect 2045 7358 2120 7370
rect 2132 7358 2163 7370
rect 2169 7358 2204 7370
rect 1838 7356 2000 7358
rect 1733 7328 1774 7336
rect 1856 7332 1869 7356
rect 1884 7354 1899 7356
rect 1696 7318 1697 7328
rect 1712 7318 1725 7328
rect 1739 7318 1740 7328
rect 1755 7318 1768 7328
rect 1783 7318 1813 7332
rect 1856 7318 1899 7332
rect 1923 7329 1930 7336
rect 1933 7332 2000 7356
rect 2032 7356 2204 7358
rect 2002 7334 2030 7338
rect 2032 7334 2112 7356
rect 2133 7354 2148 7356
rect 2002 7332 2112 7334
rect 1933 7328 2112 7332
rect 1906 7318 1936 7328
rect 1938 7318 2091 7328
rect 2099 7318 2129 7328
rect 2133 7318 2163 7332
rect 2191 7318 2204 7356
rect 2276 7362 2311 7370
rect 2276 7336 2277 7362
rect 2284 7336 2311 7362
rect 2219 7318 2249 7332
rect 2276 7328 2311 7336
rect 2313 7362 2354 7370
rect 2313 7336 2328 7362
rect 2335 7336 2354 7362
rect 2418 7358 2480 7370
rect 2492 7358 2567 7370
rect 2625 7358 2700 7370
rect 2712 7358 2743 7370
rect 2749 7358 2784 7370
rect 2418 7356 2580 7358
rect 2313 7328 2354 7336
rect 2436 7332 2449 7356
rect 2464 7354 2479 7356
rect 2276 7318 2277 7328
rect 2292 7318 2305 7328
rect 2319 7318 2320 7328
rect 2335 7318 2348 7328
rect 2363 7318 2393 7332
rect 2436 7318 2479 7332
rect 2503 7329 2510 7336
rect 2513 7332 2580 7356
rect 2612 7356 2784 7358
rect 2582 7334 2610 7338
rect 2612 7334 2692 7356
rect 2713 7354 2728 7356
rect 2582 7332 2692 7334
rect 2513 7328 2692 7332
rect 2486 7318 2516 7328
rect 2518 7318 2671 7328
rect 2679 7318 2709 7328
rect 2713 7318 2743 7332
rect 2771 7318 2784 7356
rect 2856 7362 2891 7370
rect 2856 7336 2857 7362
rect 2864 7336 2891 7362
rect 2799 7318 2829 7332
rect 2856 7328 2891 7336
rect 2893 7362 2934 7370
rect 2893 7336 2908 7362
rect 2915 7336 2934 7362
rect 2998 7358 3060 7370
rect 3072 7358 3147 7370
rect 3205 7358 3280 7370
rect 3292 7358 3323 7370
rect 3329 7358 3364 7370
rect 2998 7356 3160 7358
rect 2893 7328 2934 7336
rect 3016 7332 3029 7356
rect 3044 7354 3059 7356
rect 2856 7318 2857 7328
rect 2872 7318 2885 7328
rect 2899 7318 2900 7328
rect 2915 7318 2928 7328
rect 2943 7318 2973 7332
rect 3016 7318 3059 7332
rect 3083 7329 3090 7336
rect 3093 7332 3160 7356
rect 3192 7356 3364 7358
rect 3162 7334 3190 7338
rect 3192 7334 3272 7356
rect 3293 7354 3308 7356
rect 3162 7332 3272 7334
rect 3093 7328 3272 7332
rect 3066 7318 3096 7328
rect 3098 7318 3251 7328
rect 3259 7318 3289 7328
rect 3293 7318 3323 7332
rect 3351 7318 3364 7356
rect 3436 7362 3471 7370
rect 3436 7336 3437 7362
rect 3444 7336 3471 7362
rect 3379 7318 3409 7332
rect 3436 7328 3471 7336
rect 3473 7362 3514 7370
rect 3473 7336 3488 7362
rect 3495 7336 3514 7362
rect 3578 7358 3640 7370
rect 3652 7358 3727 7370
rect 3785 7358 3860 7370
rect 3872 7358 3903 7370
rect 3909 7358 3944 7370
rect 3578 7356 3740 7358
rect 3473 7328 3514 7336
rect 3596 7332 3609 7356
rect 3624 7354 3639 7356
rect 3436 7318 3437 7328
rect 3452 7318 3465 7328
rect 3479 7318 3480 7328
rect 3495 7318 3508 7328
rect 3523 7318 3553 7332
rect 3596 7318 3639 7332
rect 3663 7329 3670 7336
rect 3673 7332 3740 7356
rect 3772 7356 3944 7358
rect 3742 7334 3770 7338
rect 3772 7334 3852 7356
rect 3873 7354 3888 7356
rect 3742 7332 3852 7334
rect 3673 7328 3852 7332
rect 3646 7318 3676 7328
rect 3678 7318 3831 7328
rect 3839 7318 3869 7328
rect 3873 7318 3903 7332
rect 3931 7318 3944 7356
rect 4016 7362 4051 7370
rect 4016 7336 4017 7362
rect 4024 7336 4051 7362
rect 3959 7318 3989 7332
rect 4016 7328 4051 7336
rect 4053 7362 4094 7370
rect 4053 7336 4068 7362
rect 4075 7336 4094 7362
rect 4158 7358 4220 7370
rect 4232 7358 4307 7370
rect 4365 7358 4440 7370
rect 4452 7358 4483 7370
rect 4489 7358 4524 7370
rect 4158 7356 4320 7358
rect 4053 7328 4094 7336
rect 4176 7332 4189 7356
rect 4204 7354 4219 7356
rect 4016 7318 4017 7328
rect 4032 7318 4045 7328
rect 4059 7318 4060 7328
rect 4075 7318 4088 7328
rect 4103 7318 4133 7332
rect 4176 7318 4219 7332
rect 4243 7329 4250 7336
rect 4253 7332 4320 7356
rect 4352 7356 4524 7358
rect 4322 7334 4350 7338
rect 4352 7334 4432 7356
rect 4453 7354 4468 7356
rect 4322 7332 4432 7334
rect 4253 7328 4432 7332
rect 4226 7318 4256 7328
rect 4258 7318 4411 7328
rect 4419 7318 4449 7328
rect 4453 7318 4483 7332
rect 4511 7318 4524 7356
rect 4596 7362 4631 7370
rect 4596 7336 4597 7362
rect 4604 7336 4631 7362
rect 4539 7318 4569 7332
rect 4596 7328 4631 7336
rect 4596 7318 4597 7328
rect 4612 7318 4625 7328
rect -1 7312 4625 7318
rect 0 7304 4625 7312
rect 15 7274 28 7304
rect 43 7286 73 7304
rect 116 7290 130 7304
rect 166 7290 386 7304
rect 117 7288 130 7290
rect 83 7276 98 7288
rect 80 7274 102 7276
rect 107 7274 137 7288
rect 198 7286 351 7290
rect 180 7274 372 7286
rect 415 7274 445 7288
rect 451 7274 464 7304
rect 479 7286 509 7304
rect 552 7274 565 7304
rect 595 7274 608 7304
rect 623 7286 653 7304
rect 696 7290 710 7304
rect 746 7290 966 7304
rect 697 7288 710 7290
rect 663 7276 678 7288
rect 660 7274 682 7276
rect 687 7274 717 7288
rect 778 7286 931 7290
rect 760 7274 952 7286
rect 995 7274 1025 7288
rect 1031 7274 1044 7304
rect 1059 7286 1089 7304
rect 1132 7274 1145 7304
rect 1175 7274 1188 7304
rect 1203 7286 1233 7304
rect 1276 7290 1290 7304
rect 1326 7290 1546 7304
rect 1277 7288 1290 7290
rect 1243 7276 1258 7288
rect 1240 7274 1262 7276
rect 1267 7274 1297 7288
rect 1358 7286 1511 7290
rect 1340 7274 1532 7286
rect 1575 7274 1605 7288
rect 1611 7274 1624 7304
rect 1639 7286 1669 7304
rect 1712 7274 1725 7304
rect 1755 7274 1768 7304
rect 1783 7286 1813 7304
rect 1856 7290 1870 7304
rect 1906 7290 2126 7304
rect 1857 7288 1870 7290
rect 1823 7276 1838 7288
rect 1820 7274 1842 7276
rect 1847 7274 1877 7288
rect 1938 7286 2091 7290
rect 1920 7274 2112 7286
rect 2155 7274 2185 7288
rect 2191 7274 2204 7304
rect 2219 7286 2249 7304
rect 2292 7274 2305 7304
rect 2335 7274 2348 7304
rect 2363 7286 2393 7304
rect 2436 7290 2450 7304
rect 2486 7290 2706 7304
rect 2437 7288 2450 7290
rect 2403 7276 2418 7288
rect 2400 7274 2422 7276
rect 2427 7274 2457 7288
rect 2518 7286 2671 7290
rect 2500 7274 2692 7286
rect 2735 7274 2765 7288
rect 2771 7274 2784 7304
rect 2799 7286 2829 7304
rect 2872 7274 2885 7304
rect 2915 7274 2928 7304
rect 2943 7286 2973 7304
rect 3016 7290 3030 7304
rect 3066 7290 3286 7304
rect 3017 7288 3030 7290
rect 2983 7276 2998 7288
rect 2980 7274 3002 7276
rect 3007 7274 3037 7288
rect 3098 7286 3251 7290
rect 3080 7274 3272 7286
rect 3315 7274 3345 7288
rect 3351 7274 3364 7304
rect 3379 7286 3409 7304
rect 3452 7274 3465 7304
rect 3495 7274 3508 7304
rect 3523 7286 3553 7304
rect 3596 7290 3610 7304
rect 3646 7290 3866 7304
rect 3597 7288 3610 7290
rect 3563 7276 3578 7288
rect 3560 7274 3582 7276
rect 3587 7274 3617 7288
rect 3678 7286 3831 7290
rect 3660 7274 3852 7286
rect 3895 7274 3925 7288
rect 3931 7274 3944 7304
rect 3959 7286 3989 7304
rect 4032 7274 4045 7304
rect 4075 7274 4088 7304
rect 4103 7286 4133 7304
rect 4176 7290 4190 7304
rect 4226 7290 4446 7304
rect 4177 7288 4190 7290
rect 4143 7276 4158 7288
rect 4140 7274 4162 7276
rect 4167 7274 4197 7288
rect 4258 7286 4411 7290
rect 4240 7274 4432 7286
rect 4475 7274 4505 7288
rect 4511 7274 4524 7304
rect 4539 7286 4569 7304
rect 4612 7274 4625 7304
rect 0 7260 4625 7274
rect 15 7156 28 7260
rect 73 7238 74 7248
rect 89 7238 102 7248
rect 73 7234 102 7238
rect 107 7234 137 7260
rect 155 7246 171 7248
rect 243 7246 296 7260
rect 244 7244 308 7246
rect 351 7244 366 7260
rect 415 7257 445 7260
rect 415 7254 451 7257
rect 381 7246 397 7248
rect 155 7234 170 7238
rect 73 7232 170 7234
rect 198 7232 366 7244
rect 382 7234 397 7238
rect 415 7235 454 7254
rect 473 7248 480 7249
rect 479 7241 480 7248
rect 463 7238 464 7241
rect 479 7238 492 7241
rect 415 7234 445 7235
rect 454 7234 460 7235
rect 463 7234 492 7238
rect 382 7233 492 7234
rect 382 7232 498 7233
rect 57 7224 108 7232
rect 57 7212 82 7224
rect 89 7212 108 7224
rect 139 7224 189 7232
rect 139 7216 155 7224
rect 162 7222 189 7224
rect 198 7222 419 7232
rect 162 7212 419 7222
rect 448 7224 498 7232
rect 448 7215 464 7224
rect 57 7204 108 7212
rect 155 7204 419 7212
rect 445 7212 464 7215
rect 471 7212 498 7224
rect 445 7204 498 7212
rect 73 7196 74 7204
rect 89 7196 102 7204
rect 73 7188 89 7196
rect 70 7181 89 7184
rect 70 7172 92 7181
rect 43 7162 92 7172
rect 43 7156 73 7162
rect 92 7157 97 7162
rect 15 7140 89 7156
rect 107 7148 137 7204
rect 172 7194 380 7204
rect 415 7200 460 7204
rect 463 7203 464 7204
rect 479 7203 492 7204
rect 198 7164 387 7194
rect 213 7161 387 7164
rect 206 7158 387 7161
rect 15 7138 28 7140
rect 43 7138 77 7140
rect 15 7122 89 7138
rect 116 7134 129 7148
rect 144 7134 160 7150
rect 206 7145 217 7158
rect -1 7100 0 7116
rect 15 7100 28 7122
rect 43 7100 73 7122
rect 116 7118 178 7134
rect 206 7127 217 7143
rect 222 7138 232 7158
rect 242 7138 256 7158
rect 259 7145 268 7158
rect 284 7145 293 7158
rect 222 7127 256 7138
rect 259 7127 268 7143
rect 284 7127 293 7143
rect 300 7138 310 7158
rect 320 7138 334 7158
rect 335 7145 346 7158
rect 300 7127 334 7138
rect 335 7127 346 7143
rect 392 7134 408 7150
rect 415 7148 445 7200
rect 479 7196 480 7203
rect 464 7188 480 7196
rect 451 7156 464 7175
rect 479 7156 509 7172
rect 451 7140 525 7156
rect 451 7138 464 7140
rect 479 7138 513 7140
rect 116 7116 129 7118
rect 144 7116 178 7118
rect 116 7100 178 7116
rect 222 7111 238 7114
rect 300 7111 330 7122
rect 378 7118 424 7134
rect 451 7122 525 7138
rect 378 7116 412 7118
rect 377 7100 424 7116
rect 451 7100 464 7122
rect 479 7100 509 7122
rect 536 7100 537 7116
rect 552 7100 565 7260
rect 595 7156 608 7260
rect 653 7238 654 7248
rect 669 7238 682 7248
rect 653 7234 682 7238
rect 687 7234 717 7260
rect 735 7246 751 7248
rect 823 7246 876 7260
rect 824 7244 888 7246
rect 931 7244 946 7260
rect 995 7257 1025 7260
rect 995 7254 1031 7257
rect 961 7246 977 7248
rect 735 7234 750 7238
rect 653 7232 750 7234
rect 778 7232 946 7244
rect 962 7234 977 7238
rect 995 7235 1034 7254
rect 1053 7248 1060 7249
rect 1059 7241 1060 7248
rect 1043 7238 1044 7241
rect 1059 7238 1072 7241
rect 995 7234 1025 7235
rect 1034 7234 1040 7235
rect 1043 7234 1072 7238
rect 962 7233 1072 7234
rect 962 7232 1078 7233
rect 637 7224 688 7232
rect 637 7212 662 7224
rect 669 7212 688 7224
rect 719 7224 769 7232
rect 719 7216 735 7224
rect 742 7222 769 7224
rect 778 7222 999 7232
rect 742 7212 999 7222
rect 1028 7224 1078 7232
rect 1028 7215 1044 7224
rect 637 7204 688 7212
rect 735 7204 999 7212
rect 1025 7212 1044 7215
rect 1051 7212 1078 7224
rect 1025 7204 1078 7212
rect 653 7196 654 7204
rect 669 7196 682 7204
rect 653 7188 669 7196
rect 650 7181 669 7184
rect 650 7172 672 7181
rect 623 7162 672 7172
rect 623 7156 653 7162
rect 672 7157 677 7162
rect 595 7140 669 7156
rect 687 7148 717 7204
rect 752 7194 960 7204
rect 995 7200 1040 7204
rect 1043 7203 1044 7204
rect 1059 7203 1072 7204
rect 778 7164 967 7194
rect 793 7161 967 7164
rect 786 7158 967 7161
rect 595 7138 608 7140
rect 623 7138 657 7140
rect 595 7122 669 7138
rect 696 7134 709 7148
rect 724 7134 740 7150
rect 786 7145 797 7158
rect 579 7100 580 7116
rect 595 7100 608 7122
rect 623 7100 653 7122
rect 696 7118 758 7134
rect 786 7127 797 7143
rect 802 7138 812 7158
rect 822 7138 836 7158
rect 839 7145 848 7158
rect 864 7145 873 7158
rect 802 7127 836 7138
rect 839 7127 848 7143
rect 864 7127 873 7143
rect 880 7138 890 7158
rect 900 7138 914 7158
rect 915 7145 926 7158
rect 880 7127 914 7138
rect 915 7127 926 7143
rect 972 7134 988 7150
rect 995 7148 1025 7200
rect 1059 7196 1060 7203
rect 1044 7188 1060 7196
rect 1031 7156 1044 7175
rect 1059 7156 1089 7172
rect 1031 7140 1105 7156
rect 1031 7138 1044 7140
rect 1059 7138 1093 7140
rect 696 7116 709 7118
rect 724 7116 758 7118
rect 696 7100 758 7116
rect 802 7111 818 7114
rect 880 7111 910 7122
rect 958 7118 1004 7134
rect 1031 7122 1105 7138
rect 958 7116 992 7118
rect 957 7100 1004 7116
rect 1031 7100 1044 7122
rect 1059 7100 1089 7122
rect 1116 7100 1117 7116
rect 1132 7100 1145 7260
rect 1175 7156 1188 7260
rect 1233 7238 1234 7248
rect 1249 7238 1262 7248
rect 1233 7234 1262 7238
rect 1267 7234 1297 7260
rect 1315 7246 1331 7248
rect 1403 7246 1456 7260
rect 1404 7244 1468 7246
rect 1511 7244 1526 7260
rect 1575 7257 1605 7260
rect 1575 7254 1611 7257
rect 1541 7246 1557 7248
rect 1315 7234 1330 7238
rect 1233 7232 1330 7234
rect 1358 7232 1526 7244
rect 1542 7234 1557 7238
rect 1575 7235 1614 7254
rect 1633 7248 1640 7249
rect 1639 7241 1640 7248
rect 1623 7238 1624 7241
rect 1639 7238 1652 7241
rect 1575 7234 1605 7235
rect 1614 7234 1620 7235
rect 1623 7234 1652 7238
rect 1542 7233 1652 7234
rect 1542 7232 1658 7233
rect 1217 7224 1268 7232
rect 1217 7212 1242 7224
rect 1249 7212 1268 7224
rect 1299 7224 1349 7232
rect 1299 7216 1315 7224
rect 1322 7222 1349 7224
rect 1358 7222 1579 7232
rect 1322 7212 1579 7222
rect 1608 7224 1658 7232
rect 1608 7215 1624 7224
rect 1217 7204 1268 7212
rect 1315 7204 1579 7212
rect 1605 7212 1624 7215
rect 1631 7212 1658 7224
rect 1605 7204 1658 7212
rect 1233 7196 1234 7204
rect 1249 7196 1262 7204
rect 1233 7188 1249 7196
rect 1230 7181 1249 7184
rect 1230 7172 1252 7181
rect 1203 7162 1252 7172
rect 1203 7156 1233 7162
rect 1252 7157 1257 7162
rect 1175 7140 1249 7156
rect 1267 7148 1297 7204
rect 1332 7194 1540 7204
rect 1575 7200 1620 7204
rect 1623 7203 1624 7204
rect 1639 7203 1652 7204
rect 1358 7164 1547 7194
rect 1373 7161 1547 7164
rect 1366 7158 1547 7161
rect 1175 7138 1188 7140
rect 1203 7138 1237 7140
rect 1175 7122 1249 7138
rect 1276 7134 1289 7148
rect 1304 7134 1320 7150
rect 1366 7145 1377 7158
rect 1159 7100 1160 7116
rect 1175 7100 1188 7122
rect 1203 7100 1233 7122
rect 1276 7118 1338 7134
rect 1366 7127 1377 7143
rect 1382 7138 1392 7158
rect 1402 7138 1416 7158
rect 1419 7145 1428 7158
rect 1444 7145 1453 7158
rect 1382 7127 1416 7138
rect 1419 7127 1428 7143
rect 1444 7127 1453 7143
rect 1460 7138 1470 7158
rect 1480 7138 1494 7158
rect 1495 7145 1506 7158
rect 1460 7127 1494 7138
rect 1495 7127 1506 7143
rect 1552 7134 1568 7150
rect 1575 7148 1605 7200
rect 1639 7196 1640 7203
rect 1624 7188 1640 7196
rect 1611 7156 1624 7175
rect 1639 7156 1669 7172
rect 1611 7140 1685 7156
rect 1611 7138 1624 7140
rect 1639 7138 1673 7140
rect 1276 7116 1289 7118
rect 1304 7116 1338 7118
rect 1276 7100 1338 7116
rect 1382 7111 1398 7114
rect 1460 7111 1490 7122
rect 1538 7118 1584 7134
rect 1611 7122 1685 7138
rect 1538 7116 1572 7118
rect 1537 7100 1584 7116
rect 1611 7100 1624 7122
rect 1639 7100 1669 7122
rect 1696 7100 1697 7116
rect 1712 7100 1725 7260
rect 1755 7156 1768 7260
rect 1813 7238 1814 7248
rect 1829 7238 1842 7248
rect 1813 7234 1842 7238
rect 1847 7234 1877 7260
rect 1895 7246 1911 7248
rect 1983 7246 2036 7260
rect 1984 7244 2048 7246
rect 2091 7244 2106 7260
rect 2155 7257 2185 7260
rect 2155 7254 2191 7257
rect 2121 7246 2137 7248
rect 1895 7234 1910 7238
rect 1813 7232 1910 7234
rect 1938 7232 2106 7244
rect 2122 7234 2137 7238
rect 2155 7235 2194 7254
rect 2213 7248 2220 7249
rect 2219 7241 2220 7248
rect 2203 7238 2204 7241
rect 2219 7238 2232 7241
rect 2155 7234 2185 7235
rect 2194 7234 2200 7235
rect 2203 7234 2232 7238
rect 2122 7233 2232 7234
rect 2122 7232 2238 7233
rect 1797 7224 1848 7232
rect 1797 7212 1822 7224
rect 1829 7212 1848 7224
rect 1879 7224 1929 7232
rect 1879 7216 1895 7224
rect 1902 7222 1929 7224
rect 1938 7222 2159 7232
rect 1902 7212 2159 7222
rect 2188 7224 2238 7232
rect 2188 7215 2204 7224
rect 1797 7204 1848 7212
rect 1895 7204 2159 7212
rect 2185 7212 2204 7215
rect 2211 7212 2238 7224
rect 2185 7204 2238 7212
rect 1813 7196 1814 7204
rect 1829 7196 1842 7204
rect 1813 7188 1829 7196
rect 1810 7181 1829 7184
rect 1810 7172 1832 7181
rect 1783 7162 1832 7172
rect 1783 7156 1813 7162
rect 1832 7157 1837 7162
rect 1755 7140 1829 7156
rect 1847 7148 1877 7204
rect 1912 7194 2120 7204
rect 2155 7200 2200 7204
rect 2203 7203 2204 7204
rect 2219 7203 2232 7204
rect 1938 7164 2127 7194
rect 1953 7161 2127 7164
rect 1946 7158 2127 7161
rect 1755 7138 1768 7140
rect 1783 7138 1817 7140
rect 1755 7122 1829 7138
rect 1856 7134 1869 7148
rect 1884 7134 1900 7150
rect 1946 7145 1957 7158
rect 1739 7100 1740 7116
rect 1755 7100 1768 7122
rect 1783 7100 1813 7122
rect 1856 7118 1918 7134
rect 1946 7127 1957 7143
rect 1962 7138 1972 7158
rect 1982 7138 1996 7158
rect 1999 7145 2008 7158
rect 2024 7145 2033 7158
rect 1962 7127 1996 7138
rect 1999 7127 2008 7143
rect 2024 7127 2033 7143
rect 2040 7138 2050 7158
rect 2060 7138 2074 7158
rect 2075 7145 2086 7158
rect 2040 7127 2074 7138
rect 2075 7127 2086 7143
rect 2132 7134 2148 7150
rect 2155 7148 2185 7200
rect 2219 7196 2220 7203
rect 2204 7188 2220 7196
rect 2191 7156 2204 7175
rect 2219 7156 2249 7172
rect 2191 7140 2265 7156
rect 2191 7138 2204 7140
rect 2219 7138 2253 7140
rect 1856 7116 1869 7118
rect 1884 7116 1918 7118
rect 1856 7100 1918 7116
rect 1962 7111 1978 7114
rect 2040 7111 2070 7122
rect 2118 7118 2164 7134
rect 2191 7122 2265 7138
rect 2118 7116 2152 7118
rect 2117 7100 2164 7116
rect 2191 7100 2204 7122
rect 2219 7100 2249 7122
rect 2276 7100 2277 7116
rect 2292 7100 2305 7260
rect 2335 7156 2348 7260
rect 2393 7238 2394 7248
rect 2409 7238 2422 7248
rect 2393 7234 2422 7238
rect 2427 7234 2457 7260
rect 2475 7246 2491 7248
rect 2563 7246 2616 7260
rect 2564 7244 2628 7246
rect 2671 7244 2686 7260
rect 2735 7257 2765 7260
rect 2735 7254 2771 7257
rect 2701 7246 2717 7248
rect 2475 7234 2490 7238
rect 2393 7232 2490 7234
rect 2518 7232 2686 7244
rect 2702 7234 2717 7238
rect 2735 7235 2774 7254
rect 2793 7248 2800 7249
rect 2799 7241 2800 7248
rect 2783 7238 2784 7241
rect 2799 7238 2812 7241
rect 2735 7234 2765 7235
rect 2774 7234 2780 7235
rect 2783 7234 2812 7238
rect 2702 7233 2812 7234
rect 2702 7232 2818 7233
rect 2377 7224 2428 7232
rect 2377 7212 2402 7224
rect 2409 7212 2428 7224
rect 2459 7224 2509 7232
rect 2459 7216 2475 7224
rect 2482 7222 2509 7224
rect 2518 7222 2739 7232
rect 2482 7212 2739 7222
rect 2768 7224 2818 7232
rect 2768 7215 2784 7224
rect 2377 7204 2428 7212
rect 2475 7204 2739 7212
rect 2765 7212 2784 7215
rect 2791 7212 2818 7224
rect 2765 7204 2818 7212
rect 2393 7196 2394 7204
rect 2409 7196 2422 7204
rect 2393 7188 2409 7196
rect 2390 7181 2409 7184
rect 2390 7172 2412 7181
rect 2363 7162 2412 7172
rect 2363 7156 2393 7162
rect 2412 7157 2417 7162
rect 2335 7140 2409 7156
rect 2427 7148 2457 7204
rect 2492 7194 2700 7204
rect 2735 7200 2780 7204
rect 2783 7203 2784 7204
rect 2799 7203 2812 7204
rect 2518 7164 2707 7194
rect 2533 7161 2707 7164
rect 2526 7158 2707 7161
rect 2335 7138 2348 7140
rect 2363 7138 2397 7140
rect 2335 7122 2409 7138
rect 2436 7134 2449 7148
rect 2464 7134 2480 7150
rect 2526 7145 2537 7158
rect 2319 7100 2320 7116
rect 2335 7100 2348 7122
rect 2363 7100 2393 7122
rect 2436 7118 2498 7134
rect 2526 7127 2537 7143
rect 2542 7138 2552 7158
rect 2562 7138 2576 7158
rect 2579 7145 2588 7158
rect 2604 7145 2613 7158
rect 2542 7127 2576 7138
rect 2579 7127 2588 7143
rect 2604 7127 2613 7143
rect 2620 7138 2630 7158
rect 2640 7138 2654 7158
rect 2655 7145 2666 7158
rect 2620 7127 2654 7138
rect 2655 7127 2666 7143
rect 2712 7134 2728 7150
rect 2735 7148 2765 7200
rect 2799 7196 2800 7203
rect 2784 7188 2800 7196
rect 2771 7156 2784 7175
rect 2799 7156 2829 7172
rect 2771 7140 2845 7156
rect 2771 7138 2784 7140
rect 2799 7138 2833 7140
rect 2436 7116 2449 7118
rect 2464 7116 2498 7118
rect 2436 7100 2498 7116
rect 2542 7111 2558 7114
rect 2620 7111 2650 7122
rect 2698 7118 2744 7134
rect 2771 7122 2845 7138
rect 2698 7116 2732 7118
rect 2697 7100 2744 7116
rect 2771 7100 2784 7122
rect 2799 7100 2829 7122
rect 2856 7100 2857 7116
rect 2872 7100 2885 7260
rect 2915 7156 2928 7260
rect 2973 7238 2974 7248
rect 2989 7238 3002 7248
rect 2973 7234 3002 7238
rect 3007 7234 3037 7260
rect 3055 7246 3071 7248
rect 3143 7246 3196 7260
rect 3144 7244 3208 7246
rect 3251 7244 3266 7260
rect 3315 7257 3345 7260
rect 3315 7254 3351 7257
rect 3281 7246 3297 7248
rect 3055 7234 3070 7238
rect 2973 7232 3070 7234
rect 3098 7232 3266 7244
rect 3282 7234 3297 7238
rect 3315 7235 3354 7254
rect 3373 7248 3380 7249
rect 3379 7241 3380 7248
rect 3363 7238 3364 7241
rect 3379 7238 3392 7241
rect 3315 7234 3345 7235
rect 3354 7234 3360 7235
rect 3363 7234 3392 7238
rect 3282 7233 3392 7234
rect 3282 7232 3398 7233
rect 2957 7224 3008 7232
rect 2957 7212 2982 7224
rect 2989 7212 3008 7224
rect 3039 7224 3089 7232
rect 3039 7216 3055 7224
rect 3062 7222 3089 7224
rect 3098 7222 3319 7232
rect 3062 7212 3319 7222
rect 3348 7224 3398 7232
rect 3348 7215 3364 7224
rect 2957 7204 3008 7212
rect 3055 7204 3319 7212
rect 3345 7212 3364 7215
rect 3371 7212 3398 7224
rect 3345 7204 3398 7212
rect 2973 7196 2974 7204
rect 2989 7196 3002 7204
rect 2973 7188 2989 7196
rect 2970 7181 2989 7184
rect 2970 7172 2992 7181
rect 2943 7162 2992 7172
rect 2943 7156 2973 7162
rect 2992 7157 2997 7162
rect 2915 7140 2989 7156
rect 3007 7148 3037 7204
rect 3072 7194 3280 7204
rect 3315 7200 3360 7204
rect 3363 7203 3364 7204
rect 3379 7203 3392 7204
rect 3098 7164 3287 7194
rect 3113 7161 3287 7164
rect 3106 7158 3287 7161
rect 2915 7138 2928 7140
rect 2943 7138 2977 7140
rect 2915 7122 2989 7138
rect 3016 7134 3029 7148
rect 3044 7134 3060 7150
rect 3106 7145 3117 7158
rect 2899 7100 2900 7116
rect 2915 7100 2928 7122
rect 2943 7100 2973 7122
rect 3016 7118 3078 7134
rect 3106 7127 3117 7143
rect 3122 7138 3132 7158
rect 3142 7138 3156 7158
rect 3159 7145 3168 7158
rect 3184 7145 3193 7158
rect 3122 7127 3156 7138
rect 3159 7127 3168 7143
rect 3184 7127 3193 7143
rect 3200 7138 3210 7158
rect 3220 7138 3234 7158
rect 3235 7145 3246 7158
rect 3200 7127 3234 7138
rect 3235 7127 3246 7143
rect 3292 7134 3308 7150
rect 3315 7148 3345 7200
rect 3379 7196 3380 7203
rect 3364 7188 3380 7196
rect 3351 7156 3364 7175
rect 3379 7156 3409 7172
rect 3351 7140 3425 7156
rect 3351 7138 3364 7140
rect 3379 7138 3413 7140
rect 3016 7116 3029 7118
rect 3044 7116 3078 7118
rect 3016 7100 3078 7116
rect 3122 7111 3138 7114
rect 3200 7111 3230 7122
rect 3278 7118 3324 7134
rect 3351 7122 3425 7138
rect 3278 7116 3312 7118
rect 3277 7100 3324 7116
rect 3351 7100 3364 7122
rect 3379 7100 3409 7122
rect 3436 7100 3437 7116
rect 3452 7100 3465 7260
rect 3495 7156 3508 7260
rect 3553 7238 3554 7248
rect 3569 7238 3582 7248
rect 3553 7234 3582 7238
rect 3587 7234 3617 7260
rect 3635 7246 3651 7248
rect 3723 7246 3776 7260
rect 3724 7244 3788 7246
rect 3831 7244 3846 7260
rect 3895 7257 3925 7260
rect 3895 7254 3931 7257
rect 3861 7246 3877 7248
rect 3635 7234 3650 7238
rect 3553 7232 3650 7234
rect 3678 7232 3846 7244
rect 3862 7234 3877 7238
rect 3895 7235 3934 7254
rect 3953 7248 3960 7249
rect 3959 7241 3960 7248
rect 3943 7238 3944 7241
rect 3959 7238 3972 7241
rect 3895 7234 3925 7235
rect 3934 7234 3940 7235
rect 3943 7234 3972 7238
rect 3862 7233 3972 7234
rect 3862 7232 3978 7233
rect 3537 7224 3588 7232
rect 3537 7212 3562 7224
rect 3569 7212 3588 7224
rect 3619 7224 3669 7232
rect 3619 7216 3635 7224
rect 3642 7222 3669 7224
rect 3678 7222 3899 7232
rect 3642 7212 3899 7222
rect 3928 7224 3978 7232
rect 3928 7215 3944 7224
rect 3537 7204 3588 7212
rect 3635 7204 3899 7212
rect 3925 7212 3944 7215
rect 3951 7212 3978 7224
rect 3925 7204 3978 7212
rect 3553 7196 3554 7204
rect 3569 7196 3582 7204
rect 3553 7188 3569 7196
rect 3550 7181 3569 7184
rect 3550 7172 3572 7181
rect 3523 7162 3572 7172
rect 3523 7156 3553 7162
rect 3572 7157 3577 7162
rect 3495 7140 3569 7156
rect 3587 7148 3617 7204
rect 3652 7194 3860 7204
rect 3895 7200 3940 7204
rect 3943 7203 3944 7204
rect 3959 7203 3972 7204
rect 3678 7164 3867 7194
rect 3693 7161 3867 7164
rect 3686 7158 3867 7161
rect 3495 7138 3508 7140
rect 3523 7138 3557 7140
rect 3495 7122 3569 7138
rect 3596 7134 3609 7148
rect 3624 7134 3640 7150
rect 3686 7145 3697 7158
rect 3479 7100 3480 7116
rect 3495 7100 3508 7122
rect 3523 7100 3553 7122
rect 3596 7118 3658 7134
rect 3686 7127 3697 7143
rect 3702 7138 3712 7158
rect 3722 7138 3736 7158
rect 3739 7145 3748 7158
rect 3764 7145 3773 7158
rect 3702 7127 3736 7138
rect 3739 7127 3748 7143
rect 3764 7127 3773 7143
rect 3780 7138 3790 7158
rect 3800 7138 3814 7158
rect 3815 7145 3826 7158
rect 3780 7127 3814 7138
rect 3815 7127 3826 7143
rect 3872 7134 3888 7150
rect 3895 7148 3925 7200
rect 3959 7196 3960 7203
rect 3944 7188 3960 7196
rect 3931 7156 3944 7175
rect 3959 7156 3989 7172
rect 3931 7140 4005 7156
rect 3931 7138 3944 7140
rect 3959 7138 3993 7140
rect 3596 7116 3609 7118
rect 3624 7116 3658 7118
rect 3596 7100 3658 7116
rect 3702 7111 3718 7114
rect 3780 7111 3810 7122
rect 3858 7118 3904 7134
rect 3931 7122 4005 7138
rect 3858 7116 3892 7118
rect 3857 7100 3904 7116
rect 3931 7100 3944 7122
rect 3959 7100 3989 7122
rect 4016 7100 4017 7116
rect 4032 7100 4045 7260
rect 4075 7156 4088 7260
rect 4133 7238 4134 7248
rect 4149 7238 4162 7248
rect 4133 7234 4162 7238
rect 4167 7234 4197 7260
rect 4215 7246 4231 7248
rect 4303 7246 4356 7260
rect 4304 7244 4368 7246
rect 4411 7244 4426 7260
rect 4475 7257 4505 7260
rect 4475 7254 4511 7257
rect 4441 7246 4457 7248
rect 4215 7234 4230 7238
rect 4133 7232 4230 7234
rect 4258 7232 4426 7244
rect 4442 7234 4457 7238
rect 4475 7235 4514 7254
rect 4533 7248 4540 7249
rect 4539 7241 4540 7248
rect 4523 7238 4524 7241
rect 4539 7238 4552 7241
rect 4475 7234 4505 7235
rect 4514 7234 4520 7235
rect 4523 7234 4552 7238
rect 4442 7233 4552 7234
rect 4442 7232 4558 7233
rect 4117 7224 4168 7232
rect 4117 7212 4142 7224
rect 4149 7212 4168 7224
rect 4199 7224 4249 7232
rect 4199 7216 4215 7224
rect 4222 7222 4249 7224
rect 4258 7222 4479 7232
rect 4222 7212 4479 7222
rect 4508 7224 4558 7232
rect 4508 7215 4524 7224
rect 4117 7204 4168 7212
rect 4215 7204 4479 7212
rect 4505 7212 4524 7215
rect 4531 7212 4558 7224
rect 4505 7204 4558 7212
rect 4133 7196 4134 7204
rect 4149 7196 4162 7204
rect 4133 7188 4149 7196
rect 4130 7181 4149 7184
rect 4130 7172 4152 7181
rect 4103 7162 4152 7172
rect 4103 7156 4133 7162
rect 4152 7157 4157 7162
rect 4075 7140 4149 7156
rect 4167 7148 4197 7204
rect 4232 7194 4440 7204
rect 4475 7200 4520 7204
rect 4523 7203 4524 7204
rect 4539 7203 4552 7204
rect 4258 7164 4447 7194
rect 4273 7161 4447 7164
rect 4266 7158 4447 7161
rect 4075 7138 4088 7140
rect 4103 7138 4137 7140
rect 4075 7122 4149 7138
rect 4176 7134 4189 7148
rect 4204 7134 4220 7150
rect 4266 7145 4277 7158
rect 4059 7100 4060 7116
rect 4075 7100 4088 7122
rect 4103 7100 4133 7122
rect 4176 7118 4238 7134
rect 4266 7127 4277 7143
rect 4282 7138 4292 7158
rect 4302 7138 4316 7158
rect 4319 7145 4328 7158
rect 4344 7145 4353 7158
rect 4282 7127 4316 7138
rect 4319 7127 4328 7143
rect 4344 7127 4353 7143
rect 4360 7138 4370 7158
rect 4380 7138 4394 7158
rect 4395 7145 4406 7158
rect 4360 7127 4394 7138
rect 4395 7127 4406 7143
rect 4452 7134 4468 7150
rect 4475 7148 4505 7200
rect 4539 7196 4540 7203
rect 4524 7188 4540 7196
rect 4511 7156 4524 7175
rect 4539 7156 4569 7172
rect 4511 7140 4585 7156
rect 4511 7138 4524 7140
rect 4539 7138 4573 7140
rect 4176 7116 4189 7118
rect 4204 7116 4238 7118
rect 4176 7100 4238 7116
rect 4282 7111 4298 7114
rect 4360 7111 4390 7122
rect 4438 7118 4484 7134
rect 4511 7122 4585 7138
rect 4438 7116 4472 7118
rect 4437 7100 4484 7116
rect 4511 7100 4524 7122
rect 4539 7100 4569 7122
rect 4596 7100 4597 7116
rect 4612 7100 4625 7260
rect -7 7092 34 7100
rect -7 7066 8 7092
rect 15 7066 34 7092
rect 98 7088 160 7100
rect 172 7088 247 7100
rect 305 7088 380 7100
rect 392 7088 423 7100
rect 429 7088 464 7100
rect 98 7086 260 7088
rect -7 7058 34 7066
rect 116 7062 129 7086
rect 144 7084 159 7086
rect -1 7048 0 7058
rect 15 7048 28 7058
rect 43 7048 73 7062
rect 116 7048 159 7062
rect 183 7059 190 7066
rect 193 7062 260 7086
rect 292 7086 464 7088
rect 262 7064 290 7068
rect 292 7064 372 7086
rect 393 7084 408 7086
rect 262 7062 372 7064
rect 193 7058 372 7062
rect 166 7048 196 7058
rect 198 7048 351 7058
rect 359 7048 389 7058
rect 393 7048 423 7062
rect 451 7048 464 7086
rect 536 7092 571 7100
rect 536 7066 537 7092
rect 544 7066 571 7092
rect 479 7048 509 7062
rect 536 7058 571 7066
rect 573 7092 614 7100
rect 573 7066 588 7092
rect 595 7066 614 7092
rect 678 7088 740 7100
rect 752 7088 827 7100
rect 885 7088 960 7100
rect 972 7088 1003 7100
rect 1009 7088 1044 7100
rect 678 7086 840 7088
rect 573 7058 614 7066
rect 696 7062 709 7086
rect 724 7084 739 7086
rect 536 7048 537 7058
rect 552 7048 565 7058
rect 579 7048 580 7058
rect 595 7048 608 7058
rect 623 7048 653 7062
rect 696 7048 739 7062
rect 763 7059 770 7066
rect 773 7062 840 7086
rect 872 7086 1044 7088
rect 842 7064 870 7068
rect 872 7064 952 7086
rect 973 7084 988 7086
rect 842 7062 952 7064
rect 773 7058 952 7062
rect 746 7048 776 7058
rect 778 7048 931 7058
rect 939 7048 969 7058
rect 973 7048 1003 7062
rect 1031 7048 1044 7086
rect 1116 7092 1151 7100
rect 1116 7066 1117 7092
rect 1124 7066 1151 7092
rect 1059 7048 1089 7062
rect 1116 7058 1151 7066
rect 1153 7092 1194 7100
rect 1153 7066 1168 7092
rect 1175 7066 1194 7092
rect 1258 7088 1320 7100
rect 1332 7088 1407 7100
rect 1465 7088 1540 7100
rect 1552 7088 1583 7100
rect 1589 7088 1624 7100
rect 1258 7086 1420 7088
rect 1153 7058 1194 7066
rect 1276 7062 1289 7086
rect 1304 7084 1319 7086
rect 1116 7048 1117 7058
rect 1132 7048 1145 7058
rect 1159 7048 1160 7058
rect 1175 7048 1188 7058
rect 1203 7048 1233 7062
rect 1276 7048 1319 7062
rect 1343 7059 1350 7066
rect 1353 7062 1420 7086
rect 1452 7086 1624 7088
rect 1422 7064 1450 7068
rect 1452 7064 1532 7086
rect 1553 7084 1568 7086
rect 1422 7062 1532 7064
rect 1353 7058 1532 7062
rect 1326 7048 1356 7058
rect 1358 7048 1511 7058
rect 1519 7048 1549 7058
rect 1553 7048 1583 7062
rect 1611 7048 1624 7086
rect 1696 7092 1731 7100
rect 1696 7066 1697 7092
rect 1704 7066 1731 7092
rect 1639 7048 1669 7062
rect 1696 7058 1731 7066
rect 1733 7092 1774 7100
rect 1733 7066 1748 7092
rect 1755 7066 1774 7092
rect 1838 7088 1900 7100
rect 1912 7088 1987 7100
rect 2045 7088 2120 7100
rect 2132 7088 2163 7100
rect 2169 7088 2204 7100
rect 1838 7086 2000 7088
rect 1733 7058 1774 7066
rect 1856 7062 1869 7086
rect 1884 7084 1899 7086
rect 1696 7048 1697 7058
rect 1712 7048 1725 7058
rect 1739 7048 1740 7058
rect 1755 7048 1768 7058
rect 1783 7048 1813 7062
rect 1856 7048 1899 7062
rect 1923 7059 1930 7066
rect 1933 7062 2000 7086
rect 2032 7086 2204 7088
rect 2002 7064 2030 7068
rect 2032 7064 2112 7086
rect 2133 7084 2148 7086
rect 2002 7062 2112 7064
rect 1933 7058 2112 7062
rect 1906 7048 1936 7058
rect 1938 7048 2091 7058
rect 2099 7048 2129 7058
rect 2133 7048 2163 7062
rect 2191 7048 2204 7086
rect 2276 7092 2311 7100
rect 2276 7066 2277 7092
rect 2284 7066 2311 7092
rect 2219 7048 2249 7062
rect 2276 7058 2311 7066
rect 2313 7092 2354 7100
rect 2313 7066 2328 7092
rect 2335 7066 2354 7092
rect 2418 7088 2480 7100
rect 2492 7088 2567 7100
rect 2625 7088 2700 7100
rect 2712 7088 2743 7100
rect 2749 7088 2784 7100
rect 2418 7086 2580 7088
rect 2313 7058 2354 7066
rect 2436 7062 2449 7086
rect 2464 7084 2479 7086
rect 2276 7048 2277 7058
rect 2292 7048 2305 7058
rect 2319 7048 2320 7058
rect 2335 7048 2348 7058
rect 2363 7048 2393 7062
rect 2436 7048 2479 7062
rect 2503 7059 2510 7066
rect 2513 7062 2580 7086
rect 2612 7086 2784 7088
rect 2582 7064 2610 7068
rect 2612 7064 2692 7086
rect 2713 7084 2728 7086
rect 2582 7062 2692 7064
rect 2513 7058 2692 7062
rect 2486 7048 2516 7058
rect 2518 7048 2671 7058
rect 2679 7048 2709 7058
rect 2713 7048 2743 7062
rect 2771 7048 2784 7086
rect 2856 7092 2891 7100
rect 2856 7066 2857 7092
rect 2864 7066 2891 7092
rect 2799 7048 2829 7062
rect 2856 7058 2891 7066
rect 2893 7092 2934 7100
rect 2893 7066 2908 7092
rect 2915 7066 2934 7092
rect 2998 7088 3060 7100
rect 3072 7088 3147 7100
rect 3205 7088 3280 7100
rect 3292 7088 3323 7100
rect 3329 7088 3364 7100
rect 2998 7086 3160 7088
rect 2893 7058 2934 7066
rect 3016 7062 3029 7086
rect 3044 7084 3059 7086
rect 2856 7048 2857 7058
rect 2872 7048 2885 7058
rect 2899 7048 2900 7058
rect 2915 7048 2928 7058
rect 2943 7048 2973 7062
rect 3016 7048 3059 7062
rect 3083 7059 3090 7066
rect 3093 7062 3160 7086
rect 3192 7086 3364 7088
rect 3162 7064 3190 7068
rect 3192 7064 3272 7086
rect 3293 7084 3308 7086
rect 3162 7062 3272 7064
rect 3093 7058 3272 7062
rect 3066 7048 3096 7058
rect 3098 7048 3251 7058
rect 3259 7048 3289 7058
rect 3293 7048 3323 7062
rect 3351 7048 3364 7086
rect 3436 7092 3471 7100
rect 3436 7066 3437 7092
rect 3444 7066 3471 7092
rect 3379 7048 3409 7062
rect 3436 7058 3471 7066
rect 3473 7092 3514 7100
rect 3473 7066 3488 7092
rect 3495 7066 3514 7092
rect 3578 7088 3640 7100
rect 3652 7088 3727 7100
rect 3785 7088 3860 7100
rect 3872 7088 3903 7100
rect 3909 7088 3944 7100
rect 3578 7086 3740 7088
rect 3473 7058 3514 7066
rect 3596 7062 3609 7086
rect 3624 7084 3639 7086
rect 3436 7048 3437 7058
rect 3452 7048 3465 7058
rect 3479 7048 3480 7058
rect 3495 7048 3508 7058
rect 3523 7048 3553 7062
rect 3596 7048 3639 7062
rect 3663 7059 3670 7066
rect 3673 7062 3740 7086
rect 3772 7086 3944 7088
rect 3742 7064 3770 7068
rect 3772 7064 3852 7086
rect 3873 7084 3888 7086
rect 3742 7062 3852 7064
rect 3673 7058 3852 7062
rect 3646 7048 3676 7058
rect 3678 7048 3831 7058
rect 3839 7048 3869 7058
rect 3873 7048 3903 7062
rect 3931 7048 3944 7086
rect 4016 7092 4051 7100
rect 4016 7066 4017 7092
rect 4024 7066 4051 7092
rect 3959 7048 3989 7062
rect 4016 7058 4051 7066
rect 4053 7092 4094 7100
rect 4053 7066 4068 7092
rect 4075 7066 4094 7092
rect 4158 7088 4220 7100
rect 4232 7088 4307 7100
rect 4365 7088 4440 7100
rect 4452 7088 4483 7100
rect 4489 7088 4524 7100
rect 4158 7086 4320 7088
rect 4053 7058 4094 7066
rect 4176 7062 4189 7086
rect 4204 7084 4219 7086
rect 4016 7048 4017 7058
rect 4032 7048 4045 7058
rect 4059 7048 4060 7058
rect 4075 7048 4088 7058
rect 4103 7048 4133 7062
rect 4176 7048 4219 7062
rect 4243 7059 4250 7066
rect 4253 7062 4320 7086
rect 4352 7086 4524 7088
rect 4322 7064 4350 7068
rect 4352 7064 4432 7086
rect 4453 7084 4468 7086
rect 4322 7062 4432 7064
rect 4253 7058 4432 7062
rect 4226 7048 4256 7058
rect 4258 7048 4411 7058
rect 4419 7048 4449 7058
rect 4453 7048 4483 7062
rect 4511 7048 4524 7086
rect 4596 7092 4631 7100
rect 4596 7066 4597 7092
rect 4604 7066 4631 7092
rect 4539 7048 4569 7062
rect 4596 7058 4631 7066
rect 4596 7048 4597 7058
rect 4612 7048 4625 7058
rect -1 7042 4625 7048
rect 0 7034 4625 7042
rect 15 7004 28 7034
rect 43 7016 73 7034
rect 116 7020 130 7034
rect 166 7020 386 7034
rect 117 7018 130 7020
rect 83 7006 98 7018
rect 80 7004 102 7006
rect 107 7004 137 7018
rect 198 7016 351 7020
rect 180 7004 372 7016
rect 415 7004 445 7018
rect 451 7004 464 7034
rect 479 7016 509 7034
rect 552 7004 565 7034
rect 595 7004 608 7034
rect 623 7016 653 7034
rect 696 7020 710 7034
rect 746 7020 966 7034
rect 697 7018 710 7020
rect 663 7006 678 7018
rect 660 7004 682 7006
rect 687 7004 717 7018
rect 778 7016 931 7020
rect 760 7004 952 7016
rect 995 7004 1025 7018
rect 1031 7004 1044 7034
rect 1059 7016 1089 7034
rect 1132 7004 1145 7034
rect 1175 7004 1188 7034
rect 1203 7016 1233 7034
rect 1276 7020 1290 7034
rect 1326 7020 1546 7034
rect 1277 7018 1290 7020
rect 1243 7006 1258 7018
rect 1240 7004 1262 7006
rect 1267 7004 1297 7018
rect 1358 7016 1511 7020
rect 1340 7004 1532 7016
rect 1575 7004 1605 7018
rect 1611 7004 1624 7034
rect 1639 7016 1669 7034
rect 1712 7004 1725 7034
rect 1755 7004 1768 7034
rect 1783 7016 1813 7034
rect 1856 7020 1870 7034
rect 1906 7020 2126 7034
rect 1857 7018 1870 7020
rect 1823 7006 1838 7018
rect 1820 7004 1842 7006
rect 1847 7004 1877 7018
rect 1938 7016 2091 7020
rect 1920 7004 2112 7016
rect 2155 7004 2185 7018
rect 2191 7004 2204 7034
rect 2219 7016 2249 7034
rect 2292 7004 2305 7034
rect 2335 7004 2348 7034
rect 2363 7016 2393 7034
rect 2436 7020 2450 7034
rect 2486 7020 2706 7034
rect 2437 7018 2450 7020
rect 2403 7006 2418 7018
rect 2400 7004 2422 7006
rect 2427 7004 2457 7018
rect 2518 7016 2671 7020
rect 2500 7004 2692 7016
rect 2735 7004 2765 7018
rect 2771 7004 2784 7034
rect 2799 7016 2829 7034
rect 2872 7004 2885 7034
rect 2915 7004 2928 7034
rect 2943 7016 2973 7034
rect 3016 7020 3030 7034
rect 3066 7020 3286 7034
rect 3017 7018 3030 7020
rect 2983 7006 2998 7018
rect 2980 7004 3002 7006
rect 3007 7004 3037 7018
rect 3098 7016 3251 7020
rect 3080 7004 3272 7016
rect 3315 7004 3345 7018
rect 3351 7004 3364 7034
rect 3379 7016 3409 7034
rect 3452 7004 3465 7034
rect 3495 7004 3508 7034
rect 3523 7016 3553 7034
rect 3596 7020 3610 7034
rect 3646 7020 3866 7034
rect 3597 7018 3610 7020
rect 3563 7006 3578 7018
rect 3560 7004 3582 7006
rect 3587 7004 3617 7018
rect 3678 7016 3831 7020
rect 3660 7004 3852 7016
rect 3895 7004 3925 7018
rect 3931 7004 3944 7034
rect 3959 7016 3989 7034
rect 4032 7004 4045 7034
rect 4075 7004 4088 7034
rect 4103 7016 4133 7034
rect 4176 7020 4190 7034
rect 4226 7020 4446 7034
rect 4177 7018 4190 7020
rect 4143 7006 4158 7018
rect 4140 7004 4162 7006
rect 4167 7004 4197 7018
rect 4258 7016 4411 7020
rect 4240 7004 4432 7016
rect 4475 7004 4505 7018
rect 4511 7004 4524 7034
rect 4539 7016 4569 7034
rect 4612 7004 4625 7034
rect 0 6990 4625 7004
rect 15 6886 28 6990
rect 73 6968 74 6978
rect 89 6968 102 6978
rect 73 6964 102 6968
rect 107 6964 137 6990
rect 155 6976 171 6978
rect 243 6976 296 6990
rect 244 6974 308 6976
rect 351 6974 366 6990
rect 415 6987 445 6990
rect 415 6984 451 6987
rect 381 6976 397 6978
rect 155 6964 170 6968
rect 73 6962 170 6964
rect 198 6962 366 6974
rect 382 6964 397 6968
rect 415 6965 454 6984
rect 473 6978 480 6979
rect 479 6971 480 6978
rect 463 6968 464 6971
rect 479 6968 492 6971
rect 415 6964 445 6965
rect 454 6964 460 6965
rect 463 6964 492 6968
rect 382 6963 492 6964
rect 382 6962 498 6963
rect 57 6954 108 6962
rect 57 6942 82 6954
rect 89 6942 108 6954
rect 139 6954 189 6962
rect 139 6946 155 6954
rect 162 6952 189 6954
rect 198 6952 419 6962
rect 162 6942 419 6952
rect 448 6954 498 6962
rect 448 6945 464 6954
rect 57 6934 108 6942
rect 155 6934 419 6942
rect 445 6942 464 6945
rect 471 6942 498 6954
rect 445 6934 498 6942
rect 73 6926 74 6934
rect 89 6926 102 6934
rect 73 6918 89 6926
rect 70 6911 89 6914
rect 70 6902 92 6911
rect 43 6892 92 6902
rect 43 6886 73 6892
rect 92 6887 97 6892
rect 15 6870 89 6886
rect 107 6878 137 6934
rect 172 6924 380 6934
rect 415 6930 460 6934
rect 463 6933 464 6934
rect 479 6933 492 6934
rect 198 6894 387 6924
rect 213 6891 387 6894
rect 206 6888 387 6891
rect 15 6868 28 6870
rect 43 6868 77 6870
rect 15 6852 89 6868
rect 116 6864 129 6878
rect 144 6864 160 6880
rect 206 6875 217 6888
rect -1 6830 0 6846
rect 15 6830 28 6852
rect 43 6830 73 6852
rect 116 6848 178 6864
rect 206 6857 217 6873
rect 222 6868 232 6888
rect 242 6868 256 6888
rect 259 6875 268 6888
rect 284 6875 293 6888
rect 222 6857 256 6868
rect 259 6857 268 6873
rect 284 6857 293 6873
rect 300 6868 310 6888
rect 320 6868 334 6888
rect 335 6875 346 6888
rect 300 6857 334 6868
rect 335 6857 346 6873
rect 392 6864 408 6880
rect 415 6878 445 6930
rect 479 6926 480 6933
rect 464 6918 480 6926
rect 451 6886 464 6905
rect 479 6886 509 6902
rect 451 6870 525 6886
rect 451 6868 464 6870
rect 479 6868 513 6870
rect 116 6846 129 6848
rect 144 6846 178 6848
rect 116 6830 178 6846
rect 222 6841 238 6844
rect 300 6841 330 6852
rect 378 6848 424 6864
rect 451 6852 525 6868
rect 378 6846 412 6848
rect 377 6830 424 6846
rect 451 6830 464 6852
rect 479 6830 509 6852
rect 536 6830 537 6846
rect 552 6830 565 6990
rect 595 6886 608 6990
rect 653 6968 654 6978
rect 669 6968 682 6978
rect 653 6964 682 6968
rect 687 6964 717 6990
rect 735 6976 751 6978
rect 823 6976 876 6990
rect 824 6974 888 6976
rect 931 6974 946 6990
rect 995 6987 1025 6990
rect 995 6984 1031 6987
rect 961 6976 977 6978
rect 735 6964 750 6968
rect 653 6962 750 6964
rect 778 6962 946 6974
rect 962 6964 977 6968
rect 995 6965 1034 6984
rect 1053 6978 1060 6979
rect 1059 6971 1060 6978
rect 1043 6968 1044 6971
rect 1059 6968 1072 6971
rect 995 6964 1025 6965
rect 1034 6964 1040 6965
rect 1043 6964 1072 6968
rect 962 6963 1072 6964
rect 962 6962 1078 6963
rect 637 6954 688 6962
rect 637 6942 662 6954
rect 669 6942 688 6954
rect 719 6954 769 6962
rect 719 6946 735 6954
rect 742 6952 769 6954
rect 778 6952 999 6962
rect 742 6942 999 6952
rect 1028 6954 1078 6962
rect 1028 6945 1044 6954
rect 637 6934 688 6942
rect 735 6934 999 6942
rect 1025 6942 1044 6945
rect 1051 6942 1078 6954
rect 1025 6934 1078 6942
rect 653 6926 654 6934
rect 669 6926 682 6934
rect 653 6918 669 6926
rect 650 6911 669 6914
rect 650 6902 672 6911
rect 623 6892 672 6902
rect 623 6886 653 6892
rect 672 6887 677 6892
rect 595 6870 669 6886
rect 687 6878 717 6934
rect 752 6924 960 6934
rect 995 6930 1040 6934
rect 1043 6933 1044 6934
rect 1059 6933 1072 6934
rect 778 6894 967 6924
rect 793 6891 967 6894
rect 786 6888 967 6891
rect 595 6868 608 6870
rect 623 6868 657 6870
rect 595 6852 669 6868
rect 696 6864 709 6878
rect 724 6864 740 6880
rect 786 6875 797 6888
rect 579 6830 580 6846
rect 595 6830 608 6852
rect 623 6830 653 6852
rect 696 6848 758 6864
rect 786 6857 797 6873
rect 802 6868 812 6888
rect 822 6868 836 6888
rect 839 6875 848 6888
rect 864 6875 873 6888
rect 802 6857 836 6868
rect 839 6857 848 6873
rect 864 6857 873 6873
rect 880 6868 890 6888
rect 900 6868 914 6888
rect 915 6875 926 6888
rect 880 6857 914 6868
rect 915 6857 926 6873
rect 972 6864 988 6880
rect 995 6878 1025 6930
rect 1059 6926 1060 6933
rect 1044 6918 1060 6926
rect 1031 6886 1044 6905
rect 1059 6886 1089 6902
rect 1031 6870 1105 6886
rect 1031 6868 1044 6870
rect 1059 6868 1093 6870
rect 696 6846 709 6848
rect 724 6846 758 6848
rect 696 6830 758 6846
rect 802 6841 818 6844
rect 880 6841 910 6852
rect 958 6848 1004 6864
rect 1031 6852 1105 6868
rect 958 6846 992 6848
rect 957 6830 1004 6846
rect 1031 6830 1044 6852
rect 1059 6830 1089 6852
rect 1116 6830 1117 6846
rect 1132 6830 1145 6990
rect 1175 6886 1188 6990
rect 1233 6968 1234 6978
rect 1249 6968 1262 6978
rect 1233 6964 1262 6968
rect 1267 6964 1297 6990
rect 1315 6976 1331 6978
rect 1403 6976 1456 6990
rect 1404 6974 1468 6976
rect 1511 6974 1526 6990
rect 1575 6987 1605 6990
rect 1575 6984 1611 6987
rect 1541 6976 1557 6978
rect 1315 6964 1330 6968
rect 1233 6962 1330 6964
rect 1358 6962 1526 6974
rect 1542 6964 1557 6968
rect 1575 6965 1614 6984
rect 1633 6978 1640 6979
rect 1639 6971 1640 6978
rect 1623 6968 1624 6971
rect 1639 6968 1652 6971
rect 1575 6964 1605 6965
rect 1614 6964 1620 6965
rect 1623 6964 1652 6968
rect 1542 6963 1652 6964
rect 1542 6962 1658 6963
rect 1217 6954 1268 6962
rect 1217 6942 1242 6954
rect 1249 6942 1268 6954
rect 1299 6954 1349 6962
rect 1299 6946 1315 6954
rect 1322 6952 1349 6954
rect 1358 6952 1579 6962
rect 1322 6942 1579 6952
rect 1608 6954 1658 6962
rect 1608 6945 1624 6954
rect 1217 6934 1268 6942
rect 1315 6934 1579 6942
rect 1605 6942 1624 6945
rect 1631 6942 1658 6954
rect 1605 6934 1658 6942
rect 1233 6926 1234 6934
rect 1249 6926 1262 6934
rect 1233 6918 1249 6926
rect 1230 6911 1249 6914
rect 1230 6902 1252 6911
rect 1203 6892 1252 6902
rect 1203 6886 1233 6892
rect 1252 6887 1257 6892
rect 1175 6870 1249 6886
rect 1267 6878 1297 6934
rect 1332 6924 1540 6934
rect 1575 6930 1620 6934
rect 1623 6933 1624 6934
rect 1639 6933 1652 6934
rect 1358 6894 1547 6924
rect 1373 6891 1547 6894
rect 1366 6888 1547 6891
rect 1175 6868 1188 6870
rect 1203 6868 1237 6870
rect 1175 6852 1249 6868
rect 1276 6864 1289 6878
rect 1304 6864 1320 6880
rect 1366 6875 1377 6888
rect 1159 6830 1160 6846
rect 1175 6830 1188 6852
rect 1203 6830 1233 6852
rect 1276 6848 1338 6864
rect 1366 6857 1377 6873
rect 1382 6868 1392 6888
rect 1402 6868 1416 6888
rect 1419 6875 1428 6888
rect 1444 6875 1453 6888
rect 1382 6857 1416 6868
rect 1419 6857 1428 6873
rect 1444 6857 1453 6873
rect 1460 6868 1470 6888
rect 1480 6868 1494 6888
rect 1495 6875 1506 6888
rect 1460 6857 1494 6868
rect 1495 6857 1506 6873
rect 1552 6864 1568 6880
rect 1575 6878 1605 6930
rect 1639 6926 1640 6933
rect 1624 6918 1640 6926
rect 1611 6886 1624 6905
rect 1639 6886 1669 6902
rect 1611 6870 1685 6886
rect 1611 6868 1624 6870
rect 1639 6868 1673 6870
rect 1276 6846 1289 6848
rect 1304 6846 1338 6848
rect 1276 6830 1338 6846
rect 1382 6841 1398 6844
rect 1460 6841 1490 6852
rect 1538 6848 1584 6864
rect 1611 6852 1685 6868
rect 1538 6846 1572 6848
rect 1537 6830 1584 6846
rect 1611 6830 1624 6852
rect 1639 6830 1669 6852
rect 1696 6830 1697 6846
rect 1712 6830 1725 6990
rect 1755 6886 1768 6990
rect 1813 6968 1814 6978
rect 1829 6968 1842 6978
rect 1813 6964 1842 6968
rect 1847 6964 1877 6990
rect 1895 6976 1911 6978
rect 1983 6976 2036 6990
rect 1984 6974 2048 6976
rect 2091 6974 2106 6990
rect 2155 6987 2185 6990
rect 2155 6984 2191 6987
rect 2121 6976 2137 6978
rect 1895 6964 1910 6968
rect 1813 6962 1910 6964
rect 1938 6962 2106 6974
rect 2122 6964 2137 6968
rect 2155 6965 2194 6984
rect 2213 6978 2220 6979
rect 2219 6971 2220 6978
rect 2203 6968 2204 6971
rect 2219 6968 2232 6971
rect 2155 6964 2185 6965
rect 2194 6964 2200 6965
rect 2203 6964 2232 6968
rect 2122 6963 2232 6964
rect 2122 6962 2238 6963
rect 1797 6954 1848 6962
rect 1797 6942 1822 6954
rect 1829 6942 1848 6954
rect 1879 6954 1929 6962
rect 1879 6946 1895 6954
rect 1902 6952 1929 6954
rect 1938 6952 2159 6962
rect 1902 6942 2159 6952
rect 2188 6954 2238 6962
rect 2188 6945 2204 6954
rect 1797 6934 1848 6942
rect 1895 6934 2159 6942
rect 2185 6942 2204 6945
rect 2211 6942 2238 6954
rect 2185 6934 2238 6942
rect 1813 6926 1814 6934
rect 1829 6926 1842 6934
rect 1813 6918 1829 6926
rect 1810 6911 1829 6914
rect 1810 6902 1832 6911
rect 1783 6892 1832 6902
rect 1783 6886 1813 6892
rect 1832 6887 1837 6892
rect 1755 6870 1829 6886
rect 1847 6878 1877 6934
rect 1912 6924 2120 6934
rect 2155 6930 2200 6934
rect 2203 6933 2204 6934
rect 2219 6933 2232 6934
rect 1938 6894 2127 6924
rect 1953 6891 2127 6894
rect 1946 6888 2127 6891
rect 1755 6868 1768 6870
rect 1783 6868 1817 6870
rect 1755 6852 1829 6868
rect 1856 6864 1869 6878
rect 1884 6864 1900 6880
rect 1946 6875 1957 6888
rect 1739 6830 1740 6846
rect 1755 6830 1768 6852
rect 1783 6830 1813 6852
rect 1856 6848 1918 6864
rect 1946 6857 1957 6873
rect 1962 6868 1972 6888
rect 1982 6868 1996 6888
rect 1999 6875 2008 6888
rect 2024 6875 2033 6888
rect 1962 6857 1996 6868
rect 1999 6857 2008 6873
rect 2024 6857 2033 6873
rect 2040 6868 2050 6888
rect 2060 6868 2074 6888
rect 2075 6875 2086 6888
rect 2040 6857 2074 6868
rect 2075 6857 2086 6873
rect 2132 6864 2148 6880
rect 2155 6878 2185 6930
rect 2219 6926 2220 6933
rect 2204 6918 2220 6926
rect 2191 6886 2204 6905
rect 2219 6886 2249 6902
rect 2191 6870 2265 6886
rect 2191 6868 2204 6870
rect 2219 6868 2253 6870
rect 1856 6846 1869 6848
rect 1884 6846 1918 6848
rect 1856 6830 1918 6846
rect 1962 6841 1978 6844
rect 2040 6841 2070 6852
rect 2118 6848 2164 6864
rect 2191 6852 2265 6868
rect 2118 6846 2152 6848
rect 2117 6830 2164 6846
rect 2191 6830 2204 6852
rect 2219 6830 2249 6852
rect 2276 6830 2277 6846
rect 2292 6830 2305 6990
rect 2335 6886 2348 6990
rect 2393 6968 2394 6978
rect 2409 6968 2422 6978
rect 2393 6964 2422 6968
rect 2427 6964 2457 6990
rect 2475 6976 2491 6978
rect 2563 6976 2616 6990
rect 2564 6974 2628 6976
rect 2671 6974 2686 6990
rect 2735 6987 2765 6990
rect 2735 6984 2771 6987
rect 2701 6976 2717 6978
rect 2475 6964 2490 6968
rect 2393 6962 2490 6964
rect 2518 6962 2686 6974
rect 2702 6964 2717 6968
rect 2735 6965 2774 6984
rect 2793 6978 2800 6979
rect 2799 6971 2800 6978
rect 2783 6968 2784 6971
rect 2799 6968 2812 6971
rect 2735 6964 2765 6965
rect 2774 6964 2780 6965
rect 2783 6964 2812 6968
rect 2702 6963 2812 6964
rect 2702 6962 2818 6963
rect 2377 6954 2428 6962
rect 2377 6942 2402 6954
rect 2409 6942 2428 6954
rect 2459 6954 2509 6962
rect 2459 6946 2475 6954
rect 2482 6952 2509 6954
rect 2518 6952 2739 6962
rect 2482 6942 2739 6952
rect 2768 6954 2818 6962
rect 2768 6945 2784 6954
rect 2377 6934 2428 6942
rect 2475 6934 2739 6942
rect 2765 6942 2784 6945
rect 2791 6942 2818 6954
rect 2765 6934 2818 6942
rect 2393 6926 2394 6934
rect 2409 6926 2422 6934
rect 2393 6918 2409 6926
rect 2390 6911 2409 6914
rect 2390 6902 2412 6911
rect 2363 6892 2412 6902
rect 2363 6886 2393 6892
rect 2412 6887 2417 6892
rect 2335 6870 2409 6886
rect 2427 6878 2457 6934
rect 2492 6924 2700 6934
rect 2735 6930 2780 6934
rect 2783 6933 2784 6934
rect 2799 6933 2812 6934
rect 2518 6894 2707 6924
rect 2533 6891 2707 6894
rect 2526 6888 2707 6891
rect 2335 6868 2348 6870
rect 2363 6868 2397 6870
rect 2335 6852 2409 6868
rect 2436 6864 2449 6878
rect 2464 6864 2480 6880
rect 2526 6875 2537 6888
rect 2319 6830 2320 6846
rect 2335 6830 2348 6852
rect 2363 6830 2393 6852
rect 2436 6848 2498 6864
rect 2526 6857 2537 6873
rect 2542 6868 2552 6888
rect 2562 6868 2576 6888
rect 2579 6875 2588 6888
rect 2604 6875 2613 6888
rect 2542 6857 2576 6868
rect 2579 6857 2588 6873
rect 2604 6857 2613 6873
rect 2620 6868 2630 6888
rect 2640 6868 2654 6888
rect 2655 6875 2666 6888
rect 2620 6857 2654 6868
rect 2655 6857 2666 6873
rect 2712 6864 2728 6880
rect 2735 6878 2765 6930
rect 2799 6926 2800 6933
rect 2784 6918 2800 6926
rect 2771 6886 2784 6905
rect 2799 6886 2829 6902
rect 2771 6870 2845 6886
rect 2771 6868 2784 6870
rect 2799 6868 2833 6870
rect 2436 6846 2449 6848
rect 2464 6846 2498 6848
rect 2436 6830 2498 6846
rect 2542 6841 2558 6844
rect 2620 6841 2650 6852
rect 2698 6848 2744 6864
rect 2771 6852 2845 6868
rect 2698 6846 2732 6848
rect 2697 6830 2744 6846
rect 2771 6830 2784 6852
rect 2799 6830 2829 6852
rect 2856 6830 2857 6846
rect 2872 6830 2885 6990
rect 2915 6886 2928 6990
rect 2973 6968 2974 6978
rect 2989 6968 3002 6978
rect 2973 6964 3002 6968
rect 3007 6964 3037 6990
rect 3055 6976 3071 6978
rect 3143 6976 3196 6990
rect 3144 6974 3208 6976
rect 3251 6974 3266 6990
rect 3315 6987 3345 6990
rect 3315 6984 3351 6987
rect 3281 6976 3297 6978
rect 3055 6964 3070 6968
rect 2973 6962 3070 6964
rect 3098 6962 3266 6974
rect 3282 6964 3297 6968
rect 3315 6965 3354 6984
rect 3373 6978 3380 6979
rect 3379 6971 3380 6978
rect 3363 6968 3364 6971
rect 3379 6968 3392 6971
rect 3315 6964 3345 6965
rect 3354 6964 3360 6965
rect 3363 6964 3392 6968
rect 3282 6963 3392 6964
rect 3282 6962 3398 6963
rect 2957 6954 3008 6962
rect 2957 6942 2982 6954
rect 2989 6942 3008 6954
rect 3039 6954 3089 6962
rect 3039 6946 3055 6954
rect 3062 6952 3089 6954
rect 3098 6952 3319 6962
rect 3062 6942 3319 6952
rect 3348 6954 3398 6962
rect 3348 6945 3364 6954
rect 2957 6934 3008 6942
rect 3055 6934 3319 6942
rect 3345 6942 3364 6945
rect 3371 6942 3398 6954
rect 3345 6934 3398 6942
rect 2973 6926 2974 6934
rect 2989 6926 3002 6934
rect 2973 6918 2989 6926
rect 2970 6911 2989 6914
rect 2970 6902 2992 6911
rect 2943 6892 2992 6902
rect 2943 6886 2973 6892
rect 2992 6887 2997 6892
rect 2915 6870 2989 6886
rect 3007 6878 3037 6934
rect 3072 6924 3280 6934
rect 3315 6930 3360 6934
rect 3363 6933 3364 6934
rect 3379 6933 3392 6934
rect 3098 6894 3287 6924
rect 3113 6891 3287 6894
rect 3106 6888 3287 6891
rect 2915 6868 2928 6870
rect 2943 6868 2977 6870
rect 2915 6852 2989 6868
rect 3016 6864 3029 6878
rect 3044 6864 3060 6880
rect 3106 6875 3117 6888
rect 2899 6830 2900 6846
rect 2915 6830 2928 6852
rect 2943 6830 2973 6852
rect 3016 6848 3078 6864
rect 3106 6857 3117 6873
rect 3122 6868 3132 6888
rect 3142 6868 3156 6888
rect 3159 6875 3168 6888
rect 3184 6875 3193 6888
rect 3122 6857 3156 6868
rect 3159 6857 3168 6873
rect 3184 6857 3193 6873
rect 3200 6868 3210 6888
rect 3220 6868 3234 6888
rect 3235 6875 3246 6888
rect 3200 6857 3234 6868
rect 3235 6857 3246 6873
rect 3292 6864 3308 6880
rect 3315 6878 3345 6930
rect 3379 6926 3380 6933
rect 3364 6918 3380 6926
rect 3351 6886 3364 6905
rect 3379 6886 3409 6902
rect 3351 6870 3425 6886
rect 3351 6868 3364 6870
rect 3379 6868 3413 6870
rect 3016 6846 3029 6848
rect 3044 6846 3078 6848
rect 3016 6830 3078 6846
rect 3122 6841 3138 6844
rect 3200 6841 3230 6852
rect 3278 6848 3324 6864
rect 3351 6852 3425 6868
rect 3278 6846 3312 6848
rect 3277 6830 3324 6846
rect 3351 6830 3364 6852
rect 3379 6830 3409 6852
rect 3436 6830 3437 6846
rect 3452 6830 3465 6990
rect 3495 6886 3508 6990
rect 3553 6968 3554 6978
rect 3569 6968 3582 6978
rect 3553 6964 3582 6968
rect 3587 6964 3617 6990
rect 3635 6976 3651 6978
rect 3723 6976 3776 6990
rect 3724 6974 3788 6976
rect 3831 6974 3846 6990
rect 3895 6987 3925 6990
rect 3895 6984 3931 6987
rect 3861 6976 3877 6978
rect 3635 6964 3650 6968
rect 3553 6962 3650 6964
rect 3678 6962 3846 6974
rect 3862 6964 3877 6968
rect 3895 6965 3934 6984
rect 3953 6978 3960 6979
rect 3959 6971 3960 6978
rect 3943 6968 3944 6971
rect 3959 6968 3972 6971
rect 3895 6964 3925 6965
rect 3934 6964 3940 6965
rect 3943 6964 3972 6968
rect 3862 6963 3972 6964
rect 3862 6962 3978 6963
rect 3537 6954 3588 6962
rect 3537 6942 3562 6954
rect 3569 6942 3588 6954
rect 3619 6954 3669 6962
rect 3619 6946 3635 6954
rect 3642 6952 3669 6954
rect 3678 6952 3899 6962
rect 3642 6942 3899 6952
rect 3928 6954 3978 6962
rect 3928 6945 3944 6954
rect 3537 6934 3588 6942
rect 3635 6934 3899 6942
rect 3925 6942 3944 6945
rect 3951 6942 3978 6954
rect 3925 6934 3978 6942
rect 3553 6926 3554 6934
rect 3569 6926 3582 6934
rect 3553 6918 3569 6926
rect 3550 6911 3569 6914
rect 3550 6902 3572 6911
rect 3523 6892 3572 6902
rect 3523 6886 3553 6892
rect 3572 6887 3577 6892
rect 3495 6870 3569 6886
rect 3587 6878 3617 6934
rect 3652 6924 3860 6934
rect 3895 6930 3940 6934
rect 3943 6933 3944 6934
rect 3959 6933 3972 6934
rect 3678 6894 3867 6924
rect 3693 6891 3867 6894
rect 3686 6888 3867 6891
rect 3495 6868 3508 6870
rect 3523 6868 3557 6870
rect 3495 6852 3569 6868
rect 3596 6864 3609 6878
rect 3624 6864 3640 6880
rect 3686 6875 3697 6888
rect 3479 6830 3480 6846
rect 3495 6830 3508 6852
rect 3523 6830 3553 6852
rect 3596 6848 3658 6864
rect 3686 6857 3697 6873
rect 3702 6868 3712 6888
rect 3722 6868 3736 6888
rect 3739 6875 3748 6888
rect 3764 6875 3773 6888
rect 3702 6857 3736 6868
rect 3739 6857 3748 6873
rect 3764 6857 3773 6873
rect 3780 6868 3790 6888
rect 3800 6868 3814 6888
rect 3815 6875 3826 6888
rect 3780 6857 3814 6868
rect 3815 6857 3826 6873
rect 3872 6864 3888 6880
rect 3895 6878 3925 6930
rect 3959 6926 3960 6933
rect 3944 6918 3960 6926
rect 3931 6886 3944 6905
rect 3959 6886 3989 6902
rect 3931 6870 4005 6886
rect 3931 6868 3944 6870
rect 3959 6868 3993 6870
rect 3596 6846 3609 6848
rect 3624 6846 3658 6848
rect 3596 6830 3658 6846
rect 3702 6841 3718 6844
rect 3780 6841 3810 6852
rect 3858 6848 3904 6864
rect 3931 6852 4005 6868
rect 3858 6846 3892 6848
rect 3857 6830 3904 6846
rect 3931 6830 3944 6852
rect 3959 6830 3989 6852
rect 4016 6830 4017 6846
rect 4032 6830 4045 6990
rect 4075 6886 4088 6990
rect 4133 6968 4134 6978
rect 4149 6968 4162 6978
rect 4133 6964 4162 6968
rect 4167 6964 4197 6990
rect 4215 6976 4231 6978
rect 4303 6976 4356 6990
rect 4304 6974 4368 6976
rect 4411 6974 4426 6990
rect 4475 6987 4505 6990
rect 4475 6984 4511 6987
rect 4441 6976 4457 6978
rect 4215 6964 4230 6968
rect 4133 6962 4230 6964
rect 4258 6962 4426 6974
rect 4442 6964 4457 6968
rect 4475 6965 4514 6984
rect 4533 6978 4540 6979
rect 4539 6971 4540 6978
rect 4523 6968 4524 6971
rect 4539 6968 4552 6971
rect 4475 6964 4505 6965
rect 4514 6964 4520 6965
rect 4523 6964 4552 6968
rect 4442 6963 4552 6964
rect 4442 6962 4558 6963
rect 4117 6954 4168 6962
rect 4117 6942 4142 6954
rect 4149 6942 4168 6954
rect 4199 6954 4249 6962
rect 4199 6946 4215 6954
rect 4222 6952 4249 6954
rect 4258 6952 4479 6962
rect 4222 6942 4479 6952
rect 4508 6954 4558 6962
rect 4508 6945 4524 6954
rect 4117 6934 4168 6942
rect 4215 6934 4479 6942
rect 4505 6942 4524 6945
rect 4531 6942 4558 6954
rect 4505 6934 4558 6942
rect 4133 6926 4134 6934
rect 4149 6926 4162 6934
rect 4133 6918 4149 6926
rect 4130 6911 4149 6914
rect 4130 6902 4152 6911
rect 4103 6892 4152 6902
rect 4103 6886 4133 6892
rect 4152 6887 4157 6892
rect 4075 6870 4149 6886
rect 4167 6878 4197 6934
rect 4232 6924 4440 6934
rect 4475 6930 4520 6934
rect 4523 6933 4524 6934
rect 4539 6933 4552 6934
rect 4258 6894 4447 6924
rect 4273 6891 4447 6894
rect 4266 6888 4447 6891
rect 4075 6868 4088 6870
rect 4103 6868 4137 6870
rect 4075 6852 4149 6868
rect 4176 6864 4189 6878
rect 4204 6864 4220 6880
rect 4266 6875 4277 6888
rect 4059 6830 4060 6846
rect 4075 6830 4088 6852
rect 4103 6830 4133 6852
rect 4176 6848 4238 6864
rect 4266 6857 4277 6873
rect 4282 6868 4292 6888
rect 4302 6868 4316 6888
rect 4319 6875 4328 6888
rect 4344 6875 4353 6888
rect 4282 6857 4316 6868
rect 4319 6857 4328 6873
rect 4344 6857 4353 6873
rect 4360 6868 4370 6888
rect 4380 6868 4394 6888
rect 4395 6875 4406 6888
rect 4360 6857 4394 6868
rect 4395 6857 4406 6873
rect 4452 6864 4468 6880
rect 4475 6878 4505 6930
rect 4539 6926 4540 6933
rect 4524 6918 4540 6926
rect 4511 6886 4524 6905
rect 4539 6886 4569 6902
rect 4511 6870 4585 6886
rect 4511 6868 4524 6870
rect 4539 6868 4573 6870
rect 4176 6846 4189 6848
rect 4204 6846 4238 6848
rect 4176 6830 4238 6846
rect 4282 6841 4298 6844
rect 4360 6841 4390 6852
rect 4438 6848 4484 6864
rect 4511 6852 4585 6868
rect 4438 6846 4472 6848
rect 4437 6830 4484 6846
rect 4511 6830 4524 6852
rect 4539 6830 4569 6852
rect 4596 6830 4597 6846
rect 4612 6830 4625 6990
rect -7 6822 34 6830
rect -7 6796 8 6822
rect 15 6796 34 6822
rect 98 6818 160 6830
rect 172 6818 247 6830
rect 305 6818 380 6830
rect 392 6818 423 6830
rect 429 6818 464 6830
rect 98 6816 260 6818
rect -7 6788 34 6796
rect 116 6792 129 6816
rect 144 6814 159 6816
rect -1 6778 0 6788
rect 15 6778 28 6788
rect 43 6778 73 6792
rect 116 6778 159 6792
rect 183 6789 190 6796
rect 193 6792 260 6816
rect 292 6816 464 6818
rect 262 6794 290 6798
rect 292 6794 372 6816
rect 393 6814 408 6816
rect 262 6792 372 6794
rect 193 6788 372 6792
rect 166 6778 196 6788
rect 198 6778 351 6788
rect 359 6778 389 6788
rect 393 6778 423 6792
rect 451 6778 464 6816
rect 536 6822 571 6830
rect 536 6796 537 6822
rect 544 6796 571 6822
rect 479 6778 509 6792
rect 536 6788 571 6796
rect 573 6822 614 6830
rect 573 6796 588 6822
rect 595 6796 614 6822
rect 678 6818 740 6830
rect 752 6818 827 6830
rect 885 6818 960 6830
rect 972 6818 1003 6830
rect 1009 6818 1044 6830
rect 678 6816 840 6818
rect 573 6788 614 6796
rect 696 6792 709 6816
rect 724 6814 739 6816
rect 536 6778 537 6788
rect 552 6778 565 6788
rect 579 6778 580 6788
rect 595 6778 608 6788
rect 623 6778 653 6792
rect 696 6778 739 6792
rect 763 6789 770 6796
rect 773 6792 840 6816
rect 872 6816 1044 6818
rect 842 6794 870 6798
rect 872 6794 952 6816
rect 973 6814 988 6816
rect 842 6792 952 6794
rect 773 6788 952 6792
rect 746 6778 776 6788
rect 778 6778 931 6788
rect 939 6778 969 6788
rect 973 6778 1003 6792
rect 1031 6778 1044 6816
rect 1116 6822 1151 6830
rect 1116 6796 1117 6822
rect 1124 6796 1151 6822
rect 1059 6778 1089 6792
rect 1116 6788 1151 6796
rect 1153 6822 1194 6830
rect 1153 6796 1168 6822
rect 1175 6796 1194 6822
rect 1258 6818 1320 6830
rect 1332 6818 1407 6830
rect 1465 6818 1540 6830
rect 1552 6818 1583 6830
rect 1589 6818 1624 6830
rect 1258 6816 1420 6818
rect 1153 6788 1194 6796
rect 1276 6792 1289 6816
rect 1304 6814 1319 6816
rect 1116 6778 1117 6788
rect 1132 6778 1145 6788
rect 1159 6778 1160 6788
rect 1175 6778 1188 6788
rect 1203 6778 1233 6792
rect 1276 6778 1319 6792
rect 1343 6789 1350 6796
rect 1353 6792 1420 6816
rect 1452 6816 1624 6818
rect 1422 6794 1450 6798
rect 1452 6794 1532 6816
rect 1553 6814 1568 6816
rect 1422 6792 1532 6794
rect 1353 6788 1532 6792
rect 1326 6778 1356 6788
rect 1358 6778 1511 6788
rect 1519 6778 1549 6788
rect 1553 6778 1583 6792
rect 1611 6778 1624 6816
rect 1696 6822 1731 6830
rect 1696 6796 1697 6822
rect 1704 6796 1731 6822
rect 1639 6778 1669 6792
rect 1696 6788 1731 6796
rect 1733 6822 1774 6830
rect 1733 6796 1748 6822
rect 1755 6796 1774 6822
rect 1838 6818 1900 6830
rect 1912 6818 1987 6830
rect 2045 6818 2120 6830
rect 2132 6818 2163 6830
rect 2169 6818 2204 6830
rect 1838 6816 2000 6818
rect 1733 6788 1774 6796
rect 1856 6792 1869 6816
rect 1884 6814 1899 6816
rect 1696 6778 1697 6788
rect 1712 6778 1725 6788
rect 1739 6778 1740 6788
rect 1755 6778 1768 6788
rect 1783 6778 1813 6792
rect 1856 6778 1899 6792
rect 1923 6789 1930 6796
rect 1933 6792 2000 6816
rect 2032 6816 2204 6818
rect 2002 6794 2030 6798
rect 2032 6794 2112 6816
rect 2133 6814 2148 6816
rect 2002 6792 2112 6794
rect 1933 6788 2112 6792
rect 1906 6778 1936 6788
rect 1938 6778 2091 6788
rect 2099 6778 2129 6788
rect 2133 6778 2163 6792
rect 2191 6778 2204 6816
rect 2276 6822 2311 6830
rect 2276 6796 2277 6822
rect 2284 6796 2311 6822
rect 2219 6778 2249 6792
rect 2276 6788 2311 6796
rect 2313 6822 2354 6830
rect 2313 6796 2328 6822
rect 2335 6796 2354 6822
rect 2418 6818 2480 6830
rect 2492 6818 2567 6830
rect 2625 6818 2700 6830
rect 2712 6818 2743 6830
rect 2749 6818 2784 6830
rect 2418 6816 2580 6818
rect 2313 6788 2354 6796
rect 2436 6792 2449 6816
rect 2464 6814 2479 6816
rect 2276 6778 2277 6788
rect 2292 6778 2305 6788
rect 2319 6778 2320 6788
rect 2335 6778 2348 6788
rect 2363 6778 2393 6792
rect 2436 6778 2479 6792
rect 2503 6789 2510 6796
rect 2513 6792 2580 6816
rect 2612 6816 2784 6818
rect 2582 6794 2610 6798
rect 2612 6794 2692 6816
rect 2713 6814 2728 6816
rect 2582 6792 2692 6794
rect 2513 6788 2692 6792
rect 2486 6778 2516 6788
rect 2518 6778 2671 6788
rect 2679 6778 2709 6788
rect 2713 6778 2743 6792
rect 2771 6778 2784 6816
rect 2856 6822 2891 6830
rect 2856 6796 2857 6822
rect 2864 6796 2891 6822
rect 2799 6778 2829 6792
rect 2856 6788 2891 6796
rect 2893 6822 2934 6830
rect 2893 6796 2908 6822
rect 2915 6796 2934 6822
rect 2998 6818 3060 6830
rect 3072 6818 3147 6830
rect 3205 6818 3280 6830
rect 3292 6818 3323 6830
rect 3329 6818 3364 6830
rect 2998 6816 3160 6818
rect 2893 6788 2934 6796
rect 3016 6792 3029 6816
rect 3044 6814 3059 6816
rect 2856 6778 2857 6788
rect 2872 6778 2885 6788
rect 2899 6778 2900 6788
rect 2915 6778 2928 6788
rect 2943 6778 2973 6792
rect 3016 6778 3059 6792
rect 3083 6789 3090 6796
rect 3093 6792 3160 6816
rect 3192 6816 3364 6818
rect 3162 6794 3190 6798
rect 3192 6794 3272 6816
rect 3293 6814 3308 6816
rect 3162 6792 3272 6794
rect 3093 6788 3272 6792
rect 3066 6778 3096 6788
rect 3098 6778 3251 6788
rect 3259 6778 3289 6788
rect 3293 6778 3323 6792
rect 3351 6778 3364 6816
rect 3436 6822 3471 6830
rect 3436 6796 3437 6822
rect 3444 6796 3471 6822
rect 3379 6778 3409 6792
rect 3436 6788 3471 6796
rect 3473 6822 3514 6830
rect 3473 6796 3488 6822
rect 3495 6796 3514 6822
rect 3578 6818 3640 6830
rect 3652 6818 3727 6830
rect 3785 6818 3860 6830
rect 3872 6818 3903 6830
rect 3909 6818 3944 6830
rect 3578 6816 3740 6818
rect 3473 6788 3514 6796
rect 3596 6792 3609 6816
rect 3624 6814 3639 6816
rect 3436 6778 3437 6788
rect 3452 6778 3465 6788
rect 3479 6778 3480 6788
rect 3495 6778 3508 6788
rect 3523 6778 3553 6792
rect 3596 6778 3639 6792
rect 3663 6789 3670 6796
rect 3673 6792 3740 6816
rect 3772 6816 3944 6818
rect 3742 6794 3770 6798
rect 3772 6794 3852 6816
rect 3873 6814 3888 6816
rect 3742 6792 3852 6794
rect 3673 6788 3852 6792
rect 3646 6778 3676 6788
rect 3678 6778 3831 6788
rect 3839 6778 3869 6788
rect 3873 6778 3903 6792
rect 3931 6778 3944 6816
rect 4016 6822 4051 6830
rect 4016 6796 4017 6822
rect 4024 6796 4051 6822
rect 3959 6778 3989 6792
rect 4016 6788 4051 6796
rect 4053 6822 4094 6830
rect 4053 6796 4068 6822
rect 4075 6796 4094 6822
rect 4158 6818 4220 6830
rect 4232 6818 4307 6830
rect 4365 6818 4440 6830
rect 4452 6818 4483 6830
rect 4489 6818 4524 6830
rect 4158 6816 4320 6818
rect 4053 6788 4094 6796
rect 4176 6792 4189 6816
rect 4204 6814 4219 6816
rect 4016 6778 4017 6788
rect 4032 6778 4045 6788
rect 4059 6778 4060 6788
rect 4075 6778 4088 6788
rect 4103 6778 4133 6792
rect 4176 6778 4219 6792
rect 4243 6789 4250 6796
rect 4253 6792 4320 6816
rect 4352 6816 4524 6818
rect 4322 6794 4350 6798
rect 4352 6794 4432 6816
rect 4453 6814 4468 6816
rect 4322 6792 4432 6794
rect 4253 6788 4432 6792
rect 4226 6778 4256 6788
rect 4258 6778 4411 6788
rect 4419 6778 4449 6788
rect 4453 6778 4483 6792
rect 4511 6778 4524 6816
rect 4596 6822 4631 6830
rect 4596 6796 4597 6822
rect 4604 6796 4631 6822
rect 4539 6778 4569 6792
rect 4596 6788 4631 6796
rect 4596 6778 4597 6788
rect 4612 6778 4625 6788
rect -1 6772 4625 6778
rect 0 6764 4625 6772
rect 15 6734 28 6764
rect 43 6746 73 6764
rect 116 6750 130 6764
rect 166 6750 386 6764
rect 117 6748 130 6750
rect 83 6736 98 6748
rect 80 6734 102 6736
rect 107 6734 137 6748
rect 198 6746 351 6750
rect 180 6734 372 6746
rect 415 6734 445 6748
rect 451 6734 464 6764
rect 479 6746 509 6764
rect 552 6734 565 6764
rect 595 6734 608 6764
rect 623 6746 653 6764
rect 696 6750 710 6764
rect 746 6750 966 6764
rect 697 6748 710 6750
rect 663 6736 678 6748
rect 660 6734 682 6736
rect 687 6734 717 6748
rect 778 6746 931 6750
rect 760 6734 952 6746
rect 995 6734 1025 6748
rect 1031 6734 1044 6764
rect 1059 6746 1089 6764
rect 1132 6734 1145 6764
rect 1175 6734 1188 6764
rect 1203 6746 1233 6764
rect 1276 6750 1290 6764
rect 1326 6750 1546 6764
rect 1277 6748 1290 6750
rect 1243 6736 1258 6748
rect 1240 6734 1262 6736
rect 1267 6734 1297 6748
rect 1358 6746 1511 6750
rect 1340 6734 1532 6746
rect 1575 6734 1605 6748
rect 1611 6734 1624 6764
rect 1639 6746 1669 6764
rect 1712 6734 1725 6764
rect 1755 6734 1768 6764
rect 1783 6746 1813 6764
rect 1856 6750 1870 6764
rect 1906 6750 2126 6764
rect 1857 6748 1870 6750
rect 1823 6736 1838 6748
rect 1820 6734 1842 6736
rect 1847 6734 1877 6748
rect 1938 6746 2091 6750
rect 1920 6734 2112 6746
rect 2155 6734 2185 6748
rect 2191 6734 2204 6764
rect 2219 6746 2249 6764
rect 2292 6734 2305 6764
rect 2335 6734 2348 6764
rect 2363 6746 2393 6764
rect 2436 6750 2450 6764
rect 2486 6750 2706 6764
rect 2437 6748 2450 6750
rect 2403 6736 2418 6748
rect 2400 6734 2422 6736
rect 2427 6734 2457 6748
rect 2518 6746 2671 6750
rect 2500 6734 2692 6746
rect 2735 6734 2765 6748
rect 2771 6734 2784 6764
rect 2799 6746 2829 6764
rect 2872 6734 2885 6764
rect 2915 6734 2928 6764
rect 2943 6746 2973 6764
rect 3016 6750 3030 6764
rect 3066 6750 3286 6764
rect 3017 6748 3030 6750
rect 2983 6736 2998 6748
rect 2980 6734 3002 6736
rect 3007 6734 3037 6748
rect 3098 6746 3251 6750
rect 3080 6734 3272 6746
rect 3315 6734 3345 6748
rect 3351 6734 3364 6764
rect 3379 6746 3409 6764
rect 3452 6734 3465 6764
rect 3495 6734 3508 6764
rect 3523 6746 3553 6764
rect 3596 6750 3610 6764
rect 3646 6750 3866 6764
rect 3597 6748 3610 6750
rect 3563 6736 3578 6748
rect 3560 6734 3582 6736
rect 3587 6734 3617 6748
rect 3678 6746 3831 6750
rect 3660 6734 3852 6746
rect 3895 6734 3925 6748
rect 3931 6734 3944 6764
rect 3959 6746 3989 6764
rect 4032 6734 4045 6764
rect 4075 6734 4088 6764
rect 4103 6746 4133 6764
rect 4176 6750 4190 6764
rect 4226 6750 4446 6764
rect 4177 6748 4190 6750
rect 4143 6736 4158 6748
rect 4140 6734 4162 6736
rect 4167 6734 4197 6748
rect 4258 6746 4411 6750
rect 4240 6734 4432 6746
rect 4475 6734 4505 6748
rect 4511 6734 4524 6764
rect 4539 6746 4569 6764
rect 4612 6734 4625 6764
rect 0 6720 4625 6734
rect 15 6616 28 6720
rect 73 6698 74 6708
rect 89 6698 102 6708
rect 73 6694 102 6698
rect 107 6694 137 6720
rect 155 6706 171 6708
rect 243 6706 296 6720
rect 244 6704 308 6706
rect 351 6704 366 6720
rect 415 6717 445 6720
rect 415 6714 451 6717
rect 381 6706 397 6708
rect 155 6694 170 6698
rect 73 6692 170 6694
rect 198 6692 366 6704
rect 382 6694 397 6698
rect 415 6695 454 6714
rect 473 6708 480 6709
rect 479 6701 480 6708
rect 463 6698 464 6701
rect 479 6698 492 6701
rect 415 6694 445 6695
rect 454 6694 460 6695
rect 463 6694 492 6698
rect 382 6693 492 6694
rect 382 6692 498 6693
rect 57 6684 108 6692
rect 57 6672 82 6684
rect 89 6672 108 6684
rect 139 6684 189 6692
rect 139 6676 155 6684
rect 162 6682 189 6684
rect 198 6682 419 6692
rect 162 6672 419 6682
rect 448 6684 498 6692
rect 448 6675 464 6684
rect 57 6664 108 6672
rect 155 6664 419 6672
rect 445 6672 464 6675
rect 471 6672 498 6684
rect 445 6664 498 6672
rect 73 6656 74 6664
rect 89 6656 102 6664
rect 73 6648 89 6656
rect 70 6641 89 6644
rect 70 6632 92 6641
rect 43 6622 92 6632
rect 43 6616 73 6622
rect 92 6617 97 6622
rect 15 6600 89 6616
rect 107 6608 137 6664
rect 172 6654 380 6664
rect 415 6660 460 6664
rect 463 6663 464 6664
rect 479 6663 492 6664
rect 198 6624 387 6654
rect 213 6621 387 6624
rect 206 6618 387 6621
rect 15 6598 28 6600
rect 43 6598 77 6600
rect 15 6582 89 6598
rect 116 6594 129 6608
rect 144 6594 160 6610
rect 206 6605 217 6618
rect -1 6560 0 6576
rect 15 6560 28 6582
rect 43 6560 73 6582
rect 116 6578 178 6594
rect 206 6587 217 6603
rect 222 6598 232 6618
rect 242 6598 256 6618
rect 259 6605 268 6618
rect 284 6605 293 6618
rect 222 6587 256 6598
rect 259 6587 268 6603
rect 284 6587 293 6603
rect 300 6598 310 6618
rect 320 6598 334 6618
rect 335 6605 346 6618
rect 300 6587 334 6598
rect 335 6587 346 6603
rect 392 6594 408 6610
rect 415 6608 445 6660
rect 479 6656 480 6663
rect 464 6648 480 6656
rect 451 6616 464 6635
rect 479 6616 509 6632
rect 451 6600 525 6616
rect 451 6598 464 6600
rect 479 6598 513 6600
rect 116 6576 129 6578
rect 144 6576 178 6578
rect 116 6560 178 6576
rect 222 6571 238 6574
rect 300 6571 330 6582
rect 378 6578 424 6594
rect 451 6582 525 6598
rect 378 6576 412 6578
rect 377 6560 424 6576
rect 451 6560 464 6582
rect 479 6560 509 6582
rect 536 6560 537 6576
rect 552 6560 565 6720
rect 595 6616 608 6720
rect 653 6698 654 6708
rect 669 6698 682 6708
rect 653 6694 682 6698
rect 687 6694 717 6720
rect 735 6706 751 6708
rect 823 6706 876 6720
rect 824 6704 888 6706
rect 931 6704 946 6720
rect 995 6717 1025 6720
rect 995 6714 1031 6717
rect 961 6706 977 6708
rect 735 6694 750 6698
rect 653 6692 750 6694
rect 778 6692 946 6704
rect 962 6694 977 6698
rect 995 6695 1034 6714
rect 1053 6708 1060 6709
rect 1059 6701 1060 6708
rect 1043 6698 1044 6701
rect 1059 6698 1072 6701
rect 995 6694 1025 6695
rect 1034 6694 1040 6695
rect 1043 6694 1072 6698
rect 962 6693 1072 6694
rect 962 6692 1078 6693
rect 637 6684 688 6692
rect 637 6672 662 6684
rect 669 6672 688 6684
rect 719 6684 769 6692
rect 719 6676 735 6684
rect 742 6682 769 6684
rect 778 6682 999 6692
rect 742 6672 999 6682
rect 1028 6684 1078 6692
rect 1028 6675 1044 6684
rect 637 6664 688 6672
rect 735 6664 999 6672
rect 1025 6672 1044 6675
rect 1051 6672 1078 6684
rect 1025 6664 1078 6672
rect 653 6656 654 6664
rect 669 6656 682 6664
rect 653 6648 669 6656
rect 650 6641 669 6644
rect 650 6632 672 6641
rect 623 6622 672 6632
rect 623 6616 653 6622
rect 672 6617 677 6622
rect 595 6600 669 6616
rect 687 6608 717 6664
rect 752 6654 960 6664
rect 995 6660 1040 6664
rect 1043 6663 1044 6664
rect 1059 6663 1072 6664
rect 778 6624 967 6654
rect 793 6621 967 6624
rect 786 6618 967 6621
rect 595 6598 608 6600
rect 623 6598 657 6600
rect 595 6582 669 6598
rect 696 6594 709 6608
rect 724 6594 740 6610
rect 786 6605 797 6618
rect 579 6560 580 6576
rect 595 6560 608 6582
rect 623 6560 653 6582
rect 696 6578 758 6594
rect 786 6587 797 6603
rect 802 6598 812 6618
rect 822 6598 836 6618
rect 839 6605 848 6618
rect 864 6605 873 6618
rect 802 6587 836 6598
rect 839 6587 848 6603
rect 864 6587 873 6603
rect 880 6598 890 6618
rect 900 6598 914 6618
rect 915 6605 926 6618
rect 880 6587 914 6598
rect 915 6587 926 6603
rect 972 6594 988 6610
rect 995 6608 1025 6660
rect 1059 6656 1060 6663
rect 1044 6648 1060 6656
rect 1031 6616 1044 6635
rect 1059 6616 1089 6632
rect 1031 6600 1105 6616
rect 1031 6598 1044 6600
rect 1059 6598 1093 6600
rect 696 6576 709 6578
rect 724 6576 758 6578
rect 696 6560 758 6576
rect 802 6571 818 6574
rect 880 6571 910 6582
rect 958 6578 1004 6594
rect 1031 6582 1105 6598
rect 958 6576 992 6578
rect 957 6560 1004 6576
rect 1031 6560 1044 6582
rect 1059 6560 1089 6582
rect 1116 6560 1117 6576
rect 1132 6560 1145 6720
rect 1175 6616 1188 6720
rect 1233 6698 1234 6708
rect 1249 6698 1262 6708
rect 1233 6694 1262 6698
rect 1267 6694 1297 6720
rect 1315 6706 1331 6708
rect 1403 6706 1456 6720
rect 1404 6704 1468 6706
rect 1511 6704 1526 6720
rect 1575 6717 1605 6720
rect 1575 6714 1611 6717
rect 1541 6706 1557 6708
rect 1315 6694 1330 6698
rect 1233 6692 1330 6694
rect 1358 6692 1526 6704
rect 1542 6694 1557 6698
rect 1575 6695 1614 6714
rect 1633 6708 1640 6709
rect 1639 6701 1640 6708
rect 1623 6698 1624 6701
rect 1639 6698 1652 6701
rect 1575 6694 1605 6695
rect 1614 6694 1620 6695
rect 1623 6694 1652 6698
rect 1542 6693 1652 6694
rect 1542 6692 1658 6693
rect 1217 6684 1268 6692
rect 1217 6672 1242 6684
rect 1249 6672 1268 6684
rect 1299 6684 1349 6692
rect 1299 6676 1315 6684
rect 1322 6682 1349 6684
rect 1358 6682 1579 6692
rect 1322 6672 1579 6682
rect 1608 6684 1658 6692
rect 1608 6675 1624 6684
rect 1217 6664 1268 6672
rect 1315 6664 1579 6672
rect 1605 6672 1624 6675
rect 1631 6672 1658 6684
rect 1605 6664 1658 6672
rect 1233 6656 1234 6664
rect 1249 6656 1262 6664
rect 1233 6648 1249 6656
rect 1230 6641 1249 6644
rect 1230 6632 1252 6641
rect 1203 6622 1252 6632
rect 1203 6616 1233 6622
rect 1252 6617 1257 6622
rect 1175 6600 1249 6616
rect 1267 6608 1297 6664
rect 1332 6654 1540 6664
rect 1575 6660 1620 6664
rect 1623 6663 1624 6664
rect 1639 6663 1652 6664
rect 1358 6624 1547 6654
rect 1373 6621 1547 6624
rect 1366 6618 1547 6621
rect 1175 6598 1188 6600
rect 1203 6598 1237 6600
rect 1175 6582 1249 6598
rect 1276 6594 1289 6608
rect 1304 6594 1320 6610
rect 1366 6605 1377 6618
rect 1159 6560 1160 6576
rect 1175 6560 1188 6582
rect 1203 6560 1233 6582
rect 1276 6578 1338 6594
rect 1366 6587 1377 6603
rect 1382 6598 1392 6618
rect 1402 6598 1416 6618
rect 1419 6605 1428 6618
rect 1444 6605 1453 6618
rect 1382 6587 1416 6598
rect 1419 6587 1428 6603
rect 1444 6587 1453 6603
rect 1460 6598 1470 6618
rect 1480 6598 1494 6618
rect 1495 6605 1506 6618
rect 1460 6587 1494 6598
rect 1495 6587 1506 6603
rect 1552 6594 1568 6610
rect 1575 6608 1605 6660
rect 1639 6656 1640 6663
rect 1624 6648 1640 6656
rect 1611 6616 1624 6635
rect 1639 6616 1669 6632
rect 1611 6600 1685 6616
rect 1611 6598 1624 6600
rect 1639 6598 1673 6600
rect 1276 6576 1289 6578
rect 1304 6576 1338 6578
rect 1276 6560 1338 6576
rect 1382 6571 1398 6574
rect 1460 6571 1490 6582
rect 1538 6578 1584 6594
rect 1611 6582 1685 6598
rect 1538 6576 1572 6578
rect 1537 6560 1584 6576
rect 1611 6560 1624 6582
rect 1639 6560 1669 6582
rect 1696 6560 1697 6576
rect 1712 6560 1725 6720
rect 1755 6616 1768 6720
rect 1813 6698 1814 6708
rect 1829 6698 1842 6708
rect 1813 6694 1842 6698
rect 1847 6694 1877 6720
rect 1895 6706 1911 6708
rect 1983 6706 2036 6720
rect 1984 6704 2048 6706
rect 2091 6704 2106 6720
rect 2155 6717 2185 6720
rect 2155 6714 2191 6717
rect 2121 6706 2137 6708
rect 1895 6694 1910 6698
rect 1813 6692 1910 6694
rect 1938 6692 2106 6704
rect 2122 6694 2137 6698
rect 2155 6695 2194 6714
rect 2213 6708 2220 6709
rect 2219 6701 2220 6708
rect 2203 6698 2204 6701
rect 2219 6698 2232 6701
rect 2155 6694 2185 6695
rect 2194 6694 2200 6695
rect 2203 6694 2232 6698
rect 2122 6693 2232 6694
rect 2122 6692 2238 6693
rect 1797 6684 1848 6692
rect 1797 6672 1822 6684
rect 1829 6672 1848 6684
rect 1879 6684 1929 6692
rect 1879 6676 1895 6684
rect 1902 6682 1929 6684
rect 1938 6682 2159 6692
rect 1902 6672 2159 6682
rect 2188 6684 2238 6692
rect 2188 6675 2204 6684
rect 1797 6664 1848 6672
rect 1895 6664 2159 6672
rect 2185 6672 2204 6675
rect 2211 6672 2238 6684
rect 2185 6664 2238 6672
rect 1813 6656 1814 6664
rect 1829 6656 1842 6664
rect 1813 6648 1829 6656
rect 1810 6641 1829 6644
rect 1810 6632 1832 6641
rect 1783 6622 1832 6632
rect 1783 6616 1813 6622
rect 1832 6617 1837 6622
rect 1755 6600 1829 6616
rect 1847 6608 1877 6664
rect 1912 6654 2120 6664
rect 2155 6660 2200 6664
rect 2203 6663 2204 6664
rect 2219 6663 2232 6664
rect 1938 6624 2127 6654
rect 1953 6621 2127 6624
rect 1946 6618 2127 6621
rect 1755 6598 1768 6600
rect 1783 6598 1817 6600
rect 1755 6582 1829 6598
rect 1856 6594 1869 6608
rect 1884 6594 1900 6610
rect 1946 6605 1957 6618
rect 1739 6560 1740 6576
rect 1755 6560 1768 6582
rect 1783 6560 1813 6582
rect 1856 6578 1918 6594
rect 1946 6587 1957 6603
rect 1962 6598 1972 6618
rect 1982 6598 1996 6618
rect 1999 6605 2008 6618
rect 2024 6605 2033 6618
rect 1962 6587 1996 6598
rect 1999 6587 2008 6603
rect 2024 6587 2033 6603
rect 2040 6598 2050 6618
rect 2060 6598 2074 6618
rect 2075 6605 2086 6618
rect 2040 6587 2074 6598
rect 2075 6587 2086 6603
rect 2132 6594 2148 6610
rect 2155 6608 2185 6660
rect 2219 6656 2220 6663
rect 2204 6648 2220 6656
rect 2191 6616 2204 6635
rect 2219 6616 2249 6632
rect 2191 6600 2265 6616
rect 2191 6598 2204 6600
rect 2219 6598 2253 6600
rect 1856 6576 1869 6578
rect 1884 6576 1918 6578
rect 1856 6560 1918 6576
rect 1962 6571 1978 6574
rect 2040 6571 2070 6582
rect 2118 6578 2164 6594
rect 2191 6582 2265 6598
rect 2118 6576 2152 6578
rect 2117 6560 2164 6576
rect 2191 6560 2204 6582
rect 2219 6560 2249 6582
rect 2276 6560 2277 6576
rect 2292 6560 2305 6720
rect 2335 6616 2348 6720
rect 2393 6698 2394 6708
rect 2409 6698 2422 6708
rect 2393 6694 2422 6698
rect 2427 6694 2457 6720
rect 2475 6706 2491 6708
rect 2563 6706 2616 6720
rect 2564 6704 2628 6706
rect 2671 6704 2686 6720
rect 2735 6717 2765 6720
rect 2735 6714 2771 6717
rect 2701 6706 2717 6708
rect 2475 6694 2490 6698
rect 2393 6692 2490 6694
rect 2518 6692 2686 6704
rect 2702 6694 2717 6698
rect 2735 6695 2774 6714
rect 2793 6708 2800 6709
rect 2799 6701 2800 6708
rect 2783 6698 2784 6701
rect 2799 6698 2812 6701
rect 2735 6694 2765 6695
rect 2774 6694 2780 6695
rect 2783 6694 2812 6698
rect 2702 6693 2812 6694
rect 2702 6692 2818 6693
rect 2377 6684 2428 6692
rect 2377 6672 2402 6684
rect 2409 6672 2428 6684
rect 2459 6684 2509 6692
rect 2459 6676 2475 6684
rect 2482 6682 2509 6684
rect 2518 6682 2739 6692
rect 2482 6672 2739 6682
rect 2768 6684 2818 6692
rect 2768 6675 2784 6684
rect 2377 6664 2428 6672
rect 2475 6664 2739 6672
rect 2765 6672 2784 6675
rect 2791 6672 2818 6684
rect 2765 6664 2818 6672
rect 2393 6656 2394 6664
rect 2409 6656 2422 6664
rect 2393 6648 2409 6656
rect 2390 6641 2409 6644
rect 2390 6632 2412 6641
rect 2363 6622 2412 6632
rect 2363 6616 2393 6622
rect 2412 6617 2417 6622
rect 2335 6600 2409 6616
rect 2427 6608 2457 6664
rect 2492 6654 2700 6664
rect 2735 6660 2780 6664
rect 2783 6663 2784 6664
rect 2799 6663 2812 6664
rect 2518 6624 2707 6654
rect 2533 6621 2707 6624
rect 2526 6618 2707 6621
rect 2335 6598 2348 6600
rect 2363 6598 2397 6600
rect 2335 6582 2409 6598
rect 2436 6594 2449 6608
rect 2464 6594 2480 6610
rect 2526 6605 2537 6618
rect 2319 6560 2320 6576
rect 2335 6560 2348 6582
rect 2363 6560 2393 6582
rect 2436 6578 2498 6594
rect 2526 6587 2537 6603
rect 2542 6598 2552 6618
rect 2562 6598 2576 6618
rect 2579 6605 2588 6618
rect 2604 6605 2613 6618
rect 2542 6587 2576 6598
rect 2579 6587 2588 6603
rect 2604 6587 2613 6603
rect 2620 6598 2630 6618
rect 2640 6598 2654 6618
rect 2655 6605 2666 6618
rect 2620 6587 2654 6598
rect 2655 6587 2666 6603
rect 2712 6594 2728 6610
rect 2735 6608 2765 6660
rect 2799 6656 2800 6663
rect 2784 6648 2800 6656
rect 2771 6616 2784 6635
rect 2799 6616 2829 6632
rect 2771 6600 2845 6616
rect 2771 6598 2784 6600
rect 2799 6598 2833 6600
rect 2436 6576 2449 6578
rect 2464 6576 2498 6578
rect 2436 6560 2498 6576
rect 2542 6571 2558 6574
rect 2620 6571 2650 6582
rect 2698 6578 2744 6594
rect 2771 6582 2845 6598
rect 2698 6576 2732 6578
rect 2697 6560 2744 6576
rect 2771 6560 2784 6582
rect 2799 6560 2829 6582
rect 2856 6560 2857 6576
rect 2872 6560 2885 6720
rect 2915 6616 2928 6720
rect 2973 6698 2974 6708
rect 2989 6698 3002 6708
rect 2973 6694 3002 6698
rect 3007 6694 3037 6720
rect 3055 6706 3071 6708
rect 3143 6706 3196 6720
rect 3144 6704 3208 6706
rect 3251 6704 3266 6720
rect 3315 6717 3345 6720
rect 3315 6714 3351 6717
rect 3281 6706 3297 6708
rect 3055 6694 3070 6698
rect 2973 6692 3070 6694
rect 3098 6692 3266 6704
rect 3282 6694 3297 6698
rect 3315 6695 3354 6714
rect 3373 6708 3380 6709
rect 3379 6701 3380 6708
rect 3363 6698 3364 6701
rect 3379 6698 3392 6701
rect 3315 6694 3345 6695
rect 3354 6694 3360 6695
rect 3363 6694 3392 6698
rect 3282 6693 3392 6694
rect 3282 6692 3398 6693
rect 2957 6684 3008 6692
rect 2957 6672 2982 6684
rect 2989 6672 3008 6684
rect 3039 6684 3089 6692
rect 3039 6676 3055 6684
rect 3062 6682 3089 6684
rect 3098 6682 3319 6692
rect 3062 6672 3319 6682
rect 3348 6684 3398 6692
rect 3348 6675 3364 6684
rect 2957 6664 3008 6672
rect 3055 6664 3319 6672
rect 3345 6672 3364 6675
rect 3371 6672 3398 6684
rect 3345 6664 3398 6672
rect 2973 6656 2974 6664
rect 2989 6656 3002 6664
rect 2973 6648 2989 6656
rect 2970 6641 2989 6644
rect 2970 6632 2992 6641
rect 2943 6622 2992 6632
rect 2943 6616 2973 6622
rect 2992 6617 2997 6622
rect 2915 6600 2989 6616
rect 3007 6608 3037 6664
rect 3072 6654 3280 6664
rect 3315 6660 3360 6664
rect 3363 6663 3364 6664
rect 3379 6663 3392 6664
rect 3098 6624 3287 6654
rect 3113 6621 3287 6624
rect 3106 6618 3287 6621
rect 2915 6598 2928 6600
rect 2943 6598 2977 6600
rect 2915 6582 2989 6598
rect 3016 6594 3029 6608
rect 3044 6594 3060 6610
rect 3106 6605 3117 6618
rect 2899 6560 2900 6576
rect 2915 6560 2928 6582
rect 2943 6560 2973 6582
rect 3016 6578 3078 6594
rect 3106 6587 3117 6603
rect 3122 6598 3132 6618
rect 3142 6598 3156 6618
rect 3159 6605 3168 6618
rect 3184 6605 3193 6618
rect 3122 6587 3156 6598
rect 3159 6587 3168 6603
rect 3184 6587 3193 6603
rect 3200 6598 3210 6618
rect 3220 6598 3234 6618
rect 3235 6605 3246 6618
rect 3200 6587 3234 6598
rect 3235 6587 3246 6603
rect 3292 6594 3308 6610
rect 3315 6608 3345 6660
rect 3379 6656 3380 6663
rect 3364 6648 3380 6656
rect 3351 6616 3364 6635
rect 3379 6616 3409 6632
rect 3351 6600 3425 6616
rect 3351 6598 3364 6600
rect 3379 6598 3413 6600
rect 3016 6576 3029 6578
rect 3044 6576 3078 6578
rect 3016 6560 3078 6576
rect 3122 6571 3138 6574
rect 3200 6571 3230 6582
rect 3278 6578 3324 6594
rect 3351 6582 3425 6598
rect 3278 6576 3312 6578
rect 3277 6560 3324 6576
rect 3351 6560 3364 6582
rect 3379 6560 3409 6582
rect 3436 6560 3437 6576
rect 3452 6560 3465 6720
rect 3495 6616 3508 6720
rect 3553 6698 3554 6708
rect 3569 6698 3582 6708
rect 3553 6694 3582 6698
rect 3587 6694 3617 6720
rect 3635 6706 3651 6708
rect 3723 6706 3776 6720
rect 3724 6704 3788 6706
rect 3831 6704 3846 6720
rect 3895 6717 3925 6720
rect 3895 6714 3931 6717
rect 3861 6706 3877 6708
rect 3635 6694 3650 6698
rect 3553 6692 3650 6694
rect 3678 6692 3846 6704
rect 3862 6694 3877 6698
rect 3895 6695 3934 6714
rect 3953 6708 3960 6709
rect 3959 6701 3960 6708
rect 3943 6698 3944 6701
rect 3959 6698 3972 6701
rect 3895 6694 3925 6695
rect 3934 6694 3940 6695
rect 3943 6694 3972 6698
rect 3862 6693 3972 6694
rect 3862 6692 3978 6693
rect 3537 6684 3588 6692
rect 3537 6672 3562 6684
rect 3569 6672 3588 6684
rect 3619 6684 3669 6692
rect 3619 6676 3635 6684
rect 3642 6682 3669 6684
rect 3678 6682 3899 6692
rect 3642 6672 3899 6682
rect 3928 6684 3978 6692
rect 3928 6675 3944 6684
rect 3537 6664 3588 6672
rect 3635 6664 3899 6672
rect 3925 6672 3944 6675
rect 3951 6672 3978 6684
rect 3925 6664 3978 6672
rect 3553 6656 3554 6664
rect 3569 6656 3582 6664
rect 3553 6648 3569 6656
rect 3550 6641 3569 6644
rect 3550 6632 3572 6641
rect 3523 6622 3572 6632
rect 3523 6616 3553 6622
rect 3572 6617 3577 6622
rect 3495 6600 3569 6616
rect 3587 6608 3617 6664
rect 3652 6654 3860 6664
rect 3895 6660 3940 6664
rect 3943 6663 3944 6664
rect 3959 6663 3972 6664
rect 3678 6624 3867 6654
rect 3693 6621 3867 6624
rect 3686 6618 3867 6621
rect 3495 6598 3508 6600
rect 3523 6598 3557 6600
rect 3495 6582 3569 6598
rect 3596 6594 3609 6608
rect 3624 6594 3640 6610
rect 3686 6605 3697 6618
rect 3479 6560 3480 6576
rect 3495 6560 3508 6582
rect 3523 6560 3553 6582
rect 3596 6578 3658 6594
rect 3686 6587 3697 6603
rect 3702 6598 3712 6618
rect 3722 6598 3736 6618
rect 3739 6605 3748 6618
rect 3764 6605 3773 6618
rect 3702 6587 3736 6598
rect 3739 6587 3748 6603
rect 3764 6587 3773 6603
rect 3780 6598 3790 6618
rect 3800 6598 3814 6618
rect 3815 6605 3826 6618
rect 3780 6587 3814 6598
rect 3815 6587 3826 6603
rect 3872 6594 3888 6610
rect 3895 6608 3925 6660
rect 3959 6656 3960 6663
rect 3944 6648 3960 6656
rect 3931 6616 3944 6635
rect 3959 6616 3989 6632
rect 3931 6600 4005 6616
rect 3931 6598 3944 6600
rect 3959 6598 3993 6600
rect 3596 6576 3609 6578
rect 3624 6576 3658 6578
rect 3596 6560 3658 6576
rect 3702 6571 3718 6574
rect 3780 6571 3810 6582
rect 3858 6578 3904 6594
rect 3931 6582 4005 6598
rect 3858 6576 3892 6578
rect 3857 6560 3904 6576
rect 3931 6560 3944 6582
rect 3959 6560 3989 6582
rect 4016 6560 4017 6576
rect 4032 6560 4045 6720
rect 4075 6616 4088 6720
rect 4133 6698 4134 6708
rect 4149 6698 4162 6708
rect 4133 6694 4162 6698
rect 4167 6694 4197 6720
rect 4215 6706 4231 6708
rect 4303 6706 4356 6720
rect 4304 6704 4368 6706
rect 4411 6704 4426 6720
rect 4475 6717 4505 6720
rect 4475 6714 4511 6717
rect 4441 6706 4457 6708
rect 4215 6694 4230 6698
rect 4133 6692 4230 6694
rect 4258 6692 4426 6704
rect 4442 6694 4457 6698
rect 4475 6695 4514 6714
rect 4533 6708 4540 6709
rect 4539 6701 4540 6708
rect 4523 6698 4524 6701
rect 4539 6698 4552 6701
rect 4475 6694 4505 6695
rect 4514 6694 4520 6695
rect 4523 6694 4552 6698
rect 4442 6693 4552 6694
rect 4442 6692 4558 6693
rect 4117 6684 4168 6692
rect 4117 6672 4142 6684
rect 4149 6672 4168 6684
rect 4199 6684 4249 6692
rect 4199 6676 4215 6684
rect 4222 6682 4249 6684
rect 4258 6682 4479 6692
rect 4222 6672 4479 6682
rect 4508 6684 4558 6692
rect 4508 6675 4524 6684
rect 4117 6664 4168 6672
rect 4215 6664 4479 6672
rect 4505 6672 4524 6675
rect 4531 6672 4558 6684
rect 4505 6664 4558 6672
rect 4133 6656 4134 6664
rect 4149 6656 4162 6664
rect 4133 6648 4149 6656
rect 4130 6641 4149 6644
rect 4130 6632 4152 6641
rect 4103 6622 4152 6632
rect 4103 6616 4133 6622
rect 4152 6617 4157 6622
rect 4075 6600 4149 6616
rect 4167 6608 4197 6664
rect 4232 6654 4440 6664
rect 4475 6660 4520 6664
rect 4523 6663 4524 6664
rect 4539 6663 4552 6664
rect 4258 6624 4447 6654
rect 4273 6621 4447 6624
rect 4266 6618 4447 6621
rect 4075 6598 4088 6600
rect 4103 6598 4137 6600
rect 4075 6582 4149 6598
rect 4176 6594 4189 6608
rect 4204 6594 4220 6610
rect 4266 6605 4277 6618
rect 4059 6560 4060 6576
rect 4075 6560 4088 6582
rect 4103 6560 4133 6582
rect 4176 6578 4238 6594
rect 4266 6587 4277 6603
rect 4282 6598 4292 6618
rect 4302 6598 4316 6618
rect 4319 6605 4328 6618
rect 4344 6605 4353 6618
rect 4282 6587 4316 6598
rect 4319 6587 4328 6603
rect 4344 6587 4353 6603
rect 4360 6598 4370 6618
rect 4380 6598 4394 6618
rect 4395 6605 4406 6618
rect 4360 6587 4394 6598
rect 4395 6587 4406 6603
rect 4452 6594 4468 6610
rect 4475 6608 4505 6660
rect 4539 6656 4540 6663
rect 4524 6648 4540 6656
rect 4511 6616 4524 6635
rect 4539 6616 4569 6632
rect 4511 6600 4585 6616
rect 4511 6598 4524 6600
rect 4539 6598 4573 6600
rect 4176 6576 4189 6578
rect 4204 6576 4238 6578
rect 4176 6560 4238 6576
rect 4282 6571 4298 6574
rect 4360 6571 4390 6582
rect 4438 6578 4484 6594
rect 4511 6582 4585 6598
rect 4438 6576 4472 6578
rect 4437 6560 4484 6576
rect 4511 6560 4524 6582
rect 4539 6560 4569 6582
rect 4596 6560 4597 6576
rect 4612 6560 4625 6720
rect -7 6552 34 6560
rect -7 6526 8 6552
rect 15 6526 34 6552
rect 98 6548 160 6560
rect 172 6548 247 6560
rect 305 6548 380 6560
rect 392 6548 423 6560
rect 429 6548 464 6560
rect 98 6546 260 6548
rect -7 6518 34 6526
rect 116 6522 129 6546
rect 144 6544 159 6546
rect -1 6508 0 6518
rect 15 6508 28 6518
rect 43 6508 73 6522
rect 116 6508 159 6522
rect 183 6519 190 6526
rect 193 6522 260 6546
rect 292 6546 464 6548
rect 262 6524 290 6528
rect 292 6524 372 6546
rect 393 6544 408 6546
rect 262 6522 372 6524
rect 193 6518 372 6522
rect 166 6508 196 6518
rect 198 6508 351 6518
rect 359 6508 389 6518
rect 393 6508 423 6522
rect 451 6508 464 6546
rect 536 6552 571 6560
rect 536 6526 537 6552
rect 544 6526 571 6552
rect 479 6508 509 6522
rect 536 6518 571 6526
rect 573 6552 614 6560
rect 573 6526 588 6552
rect 595 6526 614 6552
rect 678 6548 740 6560
rect 752 6548 827 6560
rect 885 6548 960 6560
rect 972 6548 1003 6560
rect 1009 6548 1044 6560
rect 678 6546 840 6548
rect 573 6518 614 6526
rect 696 6522 709 6546
rect 724 6544 739 6546
rect 536 6508 537 6518
rect 552 6508 565 6518
rect 579 6508 580 6518
rect 595 6508 608 6518
rect 623 6508 653 6522
rect 696 6508 739 6522
rect 763 6519 770 6526
rect 773 6522 840 6546
rect 872 6546 1044 6548
rect 842 6524 870 6528
rect 872 6524 952 6546
rect 973 6544 988 6546
rect 842 6522 952 6524
rect 773 6518 952 6522
rect 746 6508 776 6518
rect 778 6508 931 6518
rect 939 6508 969 6518
rect 973 6508 1003 6522
rect 1031 6508 1044 6546
rect 1116 6552 1151 6560
rect 1116 6526 1117 6552
rect 1124 6526 1151 6552
rect 1059 6508 1089 6522
rect 1116 6518 1151 6526
rect 1153 6552 1194 6560
rect 1153 6526 1168 6552
rect 1175 6526 1194 6552
rect 1258 6548 1320 6560
rect 1332 6548 1407 6560
rect 1465 6548 1540 6560
rect 1552 6548 1583 6560
rect 1589 6548 1624 6560
rect 1258 6546 1420 6548
rect 1153 6518 1194 6526
rect 1276 6522 1289 6546
rect 1304 6544 1319 6546
rect 1116 6508 1117 6518
rect 1132 6508 1145 6518
rect 1159 6508 1160 6518
rect 1175 6508 1188 6518
rect 1203 6508 1233 6522
rect 1276 6508 1319 6522
rect 1343 6519 1350 6526
rect 1353 6522 1420 6546
rect 1452 6546 1624 6548
rect 1422 6524 1450 6528
rect 1452 6524 1532 6546
rect 1553 6544 1568 6546
rect 1422 6522 1532 6524
rect 1353 6518 1532 6522
rect 1326 6508 1356 6518
rect 1358 6508 1511 6518
rect 1519 6508 1549 6518
rect 1553 6508 1583 6522
rect 1611 6508 1624 6546
rect 1696 6552 1731 6560
rect 1696 6526 1697 6552
rect 1704 6526 1731 6552
rect 1639 6508 1669 6522
rect 1696 6518 1731 6526
rect 1733 6552 1774 6560
rect 1733 6526 1748 6552
rect 1755 6526 1774 6552
rect 1838 6548 1900 6560
rect 1912 6548 1987 6560
rect 2045 6548 2120 6560
rect 2132 6548 2163 6560
rect 2169 6548 2204 6560
rect 1838 6546 2000 6548
rect 1733 6518 1774 6526
rect 1856 6522 1869 6546
rect 1884 6544 1899 6546
rect 1696 6508 1697 6518
rect 1712 6508 1725 6518
rect 1739 6508 1740 6518
rect 1755 6508 1768 6518
rect 1783 6508 1813 6522
rect 1856 6508 1899 6522
rect 1923 6519 1930 6526
rect 1933 6522 2000 6546
rect 2032 6546 2204 6548
rect 2002 6524 2030 6528
rect 2032 6524 2112 6546
rect 2133 6544 2148 6546
rect 2002 6522 2112 6524
rect 1933 6518 2112 6522
rect 1906 6508 1936 6518
rect 1938 6508 2091 6518
rect 2099 6508 2129 6518
rect 2133 6508 2163 6522
rect 2191 6508 2204 6546
rect 2276 6552 2311 6560
rect 2276 6526 2277 6552
rect 2284 6526 2311 6552
rect 2219 6508 2249 6522
rect 2276 6518 2311 6526
rect 2313 6552 2354 6560
rect 2313 6526 2328 6552
rect 2335 6526 2354 6552
rect 2418 6548 2480 6560
rect 2492 6548 2567 6560
rect 2625 6548 2700 6560
rect 2712 6548 2743 6560
rect 2749 6548 2784 6560
rect 2418 6546 2580 6548
rect 2313 6518 2354 6526
rect 2436 6522 2449 6546
rect 2464 6544 2479 6546
rect 2276 6508 2277 6518
rect 2292 6508 2305 6518
rect 2319 6508 2320 6518
rect 2335 6508 2348 6518
rect 2363 6508 2393 6522
rect 2436 6508 2479 6522
rect 2503 6519 2510 6526
rect 2513 6522 2580 6546
rect 2612 6546 2784 6548
rect 2582 6524 2610 6528
rect 2612 6524 2692 6546
rect 2713 6544 2728 6546
rect 2582 6522 2692 6524
rect 2513 6518 2692 6522
rect 2486 6508 2516 6518
rect 2518 6508 2671 6518
rect 2679 6508 2709 6518
rect 2713 6508 2743 6522
rect 2771 6508 2784 6546
rect 2856 6552 2891 6560
rect 2856 6526 2857 6552
rect 2864 6526 2891 6552
rect 2799 6508 2829 6522
rect 2856 6518 2891 6526
rect 2893 6552 2934 6560
rect 2893 6526 2908 6552
rect 2915 6526 2934 6552
rect 2998 6548 3060 6560
rect 3072 6548 3147 6560
rect 3205 6548 3280 6560
rect 3292 6548 3323 6560
rect 3329 6548 3364 6560
rect 2998 6546 3160 6548
rect 2893 6518 2934 6526
rect 3016 6522 3029 6546
rect 3044 6544 3059 6546
rect 2856 6508 2857 6518
rect 2872 6508 2885 6518
rect 2899 6508 2900 6518
rect 2915 6508 2928 6518
rect 2943 6508 2973 6522
rect 3016 6508 3059 6522
rect 3083 6519 3090 6526
rect 3093 6522 3160 6546
rect 3192 6546 3364 6548
rect 3162 6524 3190 6528
rect 3192 6524 3272 6546
rect 3293 6544 3308 6546
rect 3162 6522 3272 6524
rect 3093 6518 3272 6522
rect 3066 6508 3096 6518
rect 3098 6508 3251 6518
rect 3259 6508 3289 6518
rect 3293 6508 3323 6522
rect 3351 6508 3364 6546
rect 3436 6552 3471 6560
rect 3436 6526 3437 6552
rect 3444 6526 3471 6552
rect 3379 6508 3409 6522
rect 3436 6518 3471 6526
rect 3473 6552 3514 6560
rect 3473 6526 3488 6552
rect 3495 6526 3514 6552
rect 3578 6548 3640 6560
rect 3652 6548 3727 6560
rect 3785 6548 3860 6560
rect 3872 6548 3903 6560
rect 3909 6548 3944 6560
rect 3578 6546 3740 6548
rect 3473 6518 3514 6526
rect 3596 6522 3609 6546
rect 3624 6544 3639 6546
rect 3436 6508 3437 6518
rect 3452 6508 3465 6518
rect 3479 6508 3480 6518
rect 3495 6508 3508 6518
rect 3523 6508 3553 6522
rect 3596 6508 3639 6522
rect 3663 6519 3670 6526
rect 3673 6522 3740 6546
rect 3772 6546 3944 6548
rect 3742 6524 3770 6528
rect 3772 6524 3852 6546
rect 3873 6544 3888 6546
rect 3742 6522 3852 6524
rect 3673 6518 3852 6522
rect 3646 6508 3676 6518
rect 3678 6508 3831 6518
rect 3839 6508 3869 6518
rect 3873 6508 3903 6522
rect 3931 6508 3944 6546
rect 4016 6552 4051 6560
rect 4016 6526 4017 6552
rect 4024 6526 4051 6552
rect 3959 6508 3989 6522
rect 4016 6518 4051 6526
rect 4053 6552 4094 6560
rect 4053 6526 4068 6552
rect 4075 6526 4094 6552
rect 4158 6548 4220 6560
rect 4232 6548 4307 6560
rect 4365 6548 4440 6560
rect 4452 6548 4483 6560
rect 4489 6548 4524 6560
rect 4158 6546 4320 6548
rect 4053 6518 4094 6526
rect 4176 6522 4189 6546
rect 4204 6544 4219 6546
rect 4016 6508 4017 6518
rect 4032 6508 4045 6518
rect 4059 6508 4060 6518
rect 4075 6508 4088 6518
rect 4103 6508 4133 6522
rect 4176 6508 4219 6522
rect 4243 6519 4250 6526
rect 4253 6522 4320 6546
rect 4352 6546 4524 6548
rect 4322 6524 4350 6528
rect 4352 6524 4432 6546
rect 4453 6544 4468 6546
rect 4322 6522 4432 6524
rect 4253 6518 4432 6522
rect 4226 6508 4256 6518
rect 4258 6508 4411 6518
rect 4419 6508 4449 6518
rect 4453 6508 4483 6522
rect 4511 6508 4524 6546
rect 4596 6552 4631 6560
rect 4596 6526 4597 6552
rect 4604 6526 4631 6552
rect 4539 6508 4569 6522
rect 4596 6518 4631 6526
rect 4596 6508 4597 6518
rect 4612 6508 4625 6518
rect -1 6502 4625 6508
rect 0 6494 4625 6502
rect 15 6464 28 6494
rect 43 6476 73 6494
rect 116 6480 130 6494
rect 166 6480 386 6494
rect 117 6478 130 6480
rect 83 6466 98 6478
rect 80 6464 102 6466
rect 107 6464 137 6478
rect 198 6476 351 6480
rect 180 6464 372 6476
rect 415 6464 445 6478
rect 451 6464 464 6494
rect 479 6476 509 6494
rect 552 6464 565 6494
rect 595 6464 608 6494
rect 623 6476 653 6494
rect 696 6480 710 6494
rect 746 6480 966 6494
rect 697 6478 710 6480
rect 663 6466 678 6478
rect 660 6464 682 6466
rect 687 6464 717 6478
rect 778 6476 931 6480
rect 760 6464 952 6476
rect 995 6464 1025 6478
rect 1031 6464 1044 6494
rect 1059 6476 1089 6494
rect 1132 6464 1145 6494
rect 1175 6464 1188 6494
rect 1203 6476 1233 6494
rect 1276 6480 1290 6494
rect 1326 6480 1546 6494
rect 1277 6478 1290 6480
rect 1243 6466 1258 6478
rect 1240 6464 1262 6466
rect 1267 6464 1297 6478
rect 1358 6476 1511 6480
rect 1340 6464 1532 6476
rect 1575 6464 1605 6478
rect 1611 6464 1624 6494
rect 1639 6476 1669 6494
rect 1712 6464 1725 6494
rect 1755 6464 1768 6494
rect 1783 6476 1813 6494
rect 1856 6480 1870 6494
rect 1906 6480 2126 6494
rect 1857 6478 1870 6480
rect 1823 6466 1838 6478
rect 1820 6464 1842 6466
rect 1847 6464 1877 6478
rect 1938 6476 2091 6480
rect 1920 6464 2112 6476
rect 2155 6464 2185 6478
rect 2191 6464 2204 6494
rect 2219 6476 2249 6494
rect 2292 6464 2305 6494
rect 2335 6464 2348 6494
rect 2363 6476 2393 6494
rect 2436 6480 2450 6494
rect 2486 6480 2706 6494
rect 2437 6478 2450 6480
rect 2403 6466 2418 6478
rect 2400 6464 2422 6466
rect 2427 6464 2457 6478
rect 2518 6476 2671 6480
rect 2500 6464 2692 6476
rect 2735 6464 2765 6478
rect 2771 6464 2784 6494
rect 2799 6476 2829 6494
rect 2872 6464 2885 6494
rect 2915 6464 2928 6494
rect 2943 6476 2973 6494
rect 3016 6480 3030 6494
rect 3066 6480 3286 6494
rect 3017 6478 3030 6480
rect 2983 6466 2998 6478
rect 2980 6464 3002 6466
rect 3007 6464 3037 6478
rect 3098 6476 3251 6480
rect 3080 6464 3272 6476
rect 3315 6464 3345 6478
rect 3351 6464 3364 6494
rect 3379 6476 3409 6494
rect 3452 6464 3465 6494
rect 3495 6464 3508 6494
rect 3523 6476 3553 6494
rect 3596 6480 3610 6494
rect 3646 6480 3866 6494
rect 3597 6478 3610 6480
rect 3563 6466 3578 6478
rect 3560 6464 3582 6466
rect 3587 6464 3617 6478
rect 3678 6476 3831 6480
rect 3660 6464 3852 6476
rect 3895 6464 3925 6478
rect 3931 6464 3944 6494
rect 3959 6476 3989 6494
rect 4032 6464 4045 6494
rect 4075 6464 4088 6494
rect 4103 6476 4133 6494
rect 4176 6480 4190 6494
rect 4226 6480 4446 6494
rect 4177 6478 4190 6480
rect 4143 6466 4158 6478
rect 4140 6464 4162 6466
rect 4167 6464 4197 6478
rect 4258 6476 4411 6480
rect 4240 6464 4432 6476
rect 4475 6464 4505 6478
rect 4511 6464 4524 6494
rect 4539 6476 4569 6494
rect 4612 6464 4625 6494
rect 0 6450 4625 6464
rect 15 6346 28 6450
rect 73 6428 74 6438
rect 89 6428 102 6438
rect 73 6424 102 6428
rect 107 6424 137 6450
rect 155 6436 171 6438
rect 243 6436 296 6450
rect 244 6434 308 6436
rect 351 6434 366 6450
rect 415 6447 445 6450
rect 415 6444 451 6447
rect 381 6436 397 6438
rect 155 6424 170 6428
rect 73 6422 170 6424
rect 198 6422 366 6434
rect 382 6424 397 6428
rect 415 6425 454 6444
rect 473 6438 480 6439
rect 479 6431 480 6438
rect 463 6428 464 6431
rect 479 6428 492 6431
rect 415 6424 445 6425
rect 454 6424 460 6425
rect 463 6424 492 6428
rect 382 6423 492 6424
rect 382 6422 498 6423
rect 57 6414 108 6422
rect 57 6402 82 6414
rect 89 6402 108 6414
rect 139 6414 189 6422
rect 139 6406 155 6414
rect 162 6412 189 6414
rect 198 6412 419 6422
rect 162 6402 419 6412
rect 448 6414 498 6422
rect 448 6405 464 6414
rect 57 6394 108 6402
rect 155 6394 419 6402
rect 445 6402 464 6405
rect 471 6402 498 6414
rect 445 6394 498 6402
rect 73 6386 74 6394
rect 89 6386 102 6394
rect 73 6378 89 6386
rect 70 6371 89 6374
rect 70 6362 92 6371
rect 43 6352 92 6362
rect 43 6346 73 6352
rect 92 6347 97 6352
rect 15 6330 89 6346
rect 107 6338 137 6394
rect 172 6384 380 6394
rect 415 6390 460 6394
rect 463 6393 464 6394
rect 479 6393 492 6394
rect 198 6354 387 6384
rect 213 6351 387 6354
rect 206 6348 387 6351
rect 15 6328 28 6330
rect 43 6328 77 6330
rect 15 6312 89 6328
rect 116 6324 129 6338
rect 144 6324 160 6340
rect 206 6335 217 6348
rect -1 6290 0 6306
rect 15 6290 28 6312
rect 43 6290 73 6312
rect 116 6308 178 6324
rect 206 6317 217 6333
rect 222 6328 232 6348
rect 242 6328 256 6348
rect 259 6335 268 6348
rect 284 6335 293 6348
rect 222 6317 256 6328
rect 259 6317 268 6333
rect 284 6317 293 6333
rect 300 6328 310 6348
rect 320 6328 334 6348
rect 335 6335 346 6348
rect 300 6317 334 6328
rect 335 6317 346 6333
rect 392 6324 408 6340
rect 415 6338 445 6390
rect 479 6386 480 6393
rect 464 6378 480 6386
rect 451 6346 464 6365
rect 479 6346 509 6362
rect 451 6330 525 6346
rect 451 6328 464 6330
rect 479 6328 513 6330
rect 116 6306 129 6308
rect 144 6306 178 6308
rect 116 6290 178 6306
rect 222 6301 238 6304
rect 300 6301 330 6312
rect 378 6308 424 6324
rect 451 6312 525 6328
rect 378 6306 412 6308
rect 377 6290 424 6306
rect 451 6290 464 6312
rect 479 6290 509 6312
rect 536 6290 537 6306
rect 552 6290 565 6450
rect 595 6346 608 6450
rect 653 6428 654 6438
rect 669 6428 682 6438
rect 653 6424 682 6428
rect 687 6424 717 6450
rect 735 6436 751 6438
rect 823 6436 876 6450
rect 824 6434 888 6436
rect 931 6434 946 6450
rect 995 6447 1025 6450
rect 995 6444 1031 6447
rect 961 6436 977 6438
rect 735 6424 750 6428
rect 653 6422 750 6424
rect 778 6422 946 6434
rect 962 6424 977 6428
rect 995 6425 1034 6444
rect 1053 6438 1060 6439
rect 1059 6431 1060 6438
rect 1043 6428 1044 6431
rect 1059 6428 1072 6431
rect 995 6424 1025 6425
rect 1034 6424 1040 6425
rect 1043 6424 1072 6428
rect 962 6423 1072 6424
rect 962 6422 1078 6423
rect 637 6414 688 6422
rect 637 6402 662 6414
rect 669 6402 688 6414
rect 719 6414 769 6422
rect 719 6406 735 6414
rect 742 6412 769 6414
rect 778 6412 999 6422
rect 742 6402 999 6412
rect 1028 6414 1078 6422
rect 1028 6405 1044 6414
rect 637 6394 688 6402
rect 735 6394 999 6402
rect 1025 6402 1044 6405
rect 1051 6402 1078 6414
rect 1025 6394 1078 6402
rect 653 6386 654 6394
rect 669 6386 682 6394
rect 653 6378 669 6386
rect 650 6371 669 6374
rect 650 6362 672 6371
rect 623 6352 672 6362
rect 623 6346 653 6352
rect 672 6347 677 6352
rect 595 6330 669 6346
rect 687 6338 717 6394
rect 752 6384 960 6394
rect 995 6390 1040 6394
rect 1043 6393 1044 6394
rect 1059 6393 1072 6394
rect 778 6354 967 6384
rect 793 6351 967 6354
rect 786 6348 967 6351
rect 595 6328 608 6330
rect 623 6328 657 6330
rect 595 6312 669 6328
rect 696 6324 709 6338
rect 724 6324 740 6340
rect 786 6335 797 6348
rect 579 6290 580 6306
rect 595 6290 608 6312
rect 623 6290 653 6312
rect 696 6308 758 6324
rect 786 6317 797 6333
rect 802 6328 812 6348
rect 822 6328 836 6348
rect 839 6335 848 6348
rect 864 6335 873 6348
rect 802 6317 836 6328
rect 839 6317 848 6333
rect 864 6317 873 6333
rect 880 6328 890 6348
rect 900 6328 914 6348
rect 915 6335 926 6348
rect 880 6317 914 6328
rect 915 6317 926 6333
rect 972 6324 988 6340
rect 995 6338 1025 6390
rect 1059 6386 1060 6393
rect 1044 6378 1060 6386
rect 1031 6346 1044 6365
rect 1059 6346 1089 6362
rect 1031 6330 1105 6346
rect 1031 6328 1044 6330
rect 1059 6328 1093 6330
rect 696 6306 709 6308
rect 724 6306 758 6308
rect 696 6290 758 6306
rect 802 6301 818 6304
rect 880 6301 910 6312
rect 958 6308 1004 6324
rect 1031 6312 1105 6328
rect 958 6306 992 6308
rect 957 6290 1004 6306
rect 1031 6290 1044 6312
rect 1059 6290 1089 6312
rect 1116 6290 1117 6306
rect 1132 6290 1145 6450
rect 1175 6346 1188 6450
rect 1233 6428 1234 6438
rect 1249 6428 1262 6438
rect 1233 6424 1262 6428
rect 1267 6424 1297 6450
rect 1315 6436 1331 6438
rect 1403 6436 1456 6450
rect 1404 6434 1468 6436
rect 1511 6434 1526 6450
rect 1575 6447 1605 6450
rect 1575 6444 1611 6447
rect 1541 6436 1557 6438
rect 1315 6424 1330 6428
rect 1233 6422 1330 6424
rect 1358 6422 1526 6434
rect 1542 6424 1557 6428
rect 1575 6425 1614 6444
rect 1633 6438 1640 6439
rect 1639 6431 1640 6438
rect 1623 6428 1624 6431
rect 1639 6428 1652 6431
rect 1575 6424 1605 6425
rect 1614 6424 1620 6425
rect 1623 6424 1652 6428
rect 1542 6423 1652 6424
rect 1542 6422 1658 6423
rect 1217 6414 1268 6422
rect 1217 6402 1242 6414
rect 1249 6402 1268 6414
rect 1299 6414 1349 6422
rect 1299 6406 1315 6414
rect 1322 6412 1349 6414
rect 1358 6412 1579 6422
rect 1322 6402 1579 6412
rect 1608 6414 1658 6422
rect 1608 6405 1624 6414
rect 1217 6394 1268 6402
rect 1315 6394 1579 6402
rect 1605 6402 1624 6405
rect 1631 6402 1658 6414
rect 1605 6394 1658 6402
rect 1233 6386 1234 6394
rect 1249 6386 1262 6394
rect 1233 6378 1249 6386
rect 1230 6371 1249 6374
rect 1230 6362 1252 6371
rect 1203 6352 1252 6362
rect 1203 6346 1233 6352
rect 1252 6347 1257 6352
rect 1175 6330 1249 6346
rect 1267 6338 1297 6394
rect 1332 6384 1540 6394
rect 1575 6390 1620 6394
rect 1623 6393 1624 6394
rect 1639 6393 1652 6394
rect 1358 6354 1547 6384
rect 1373 6351 1547 6354
rect 1366 6348 1547 6351
rect 1175 6328 1188 6330
rect 1203 6328 1237 6330
rect 1175 6312 1249 6328
rect 1276 6324 1289 6338
rect 1304 6324 1320 6340
rect 1366 6335 1377 6348
rect 1159 6290 1160 6306
rect 1175 6290 1188 6312
rect 1203 6290 1233 6312
rect 1276 6308 1338 6324
rect 1366 6317 1377 6333
rect 1382 6328 1392 6348
rect 1402 6328 1416 6348
rect 1419 6335 1428 6348
rect 1444 6335 1453 6348
rect 1382 6317 1416 6328
rect 1419 6317 1428 6333
rect 1444 6317 1453 6333
rect 1460 6328 1470 6348
rect 1480 6328 1494 6348
rect 1495 6335 1506 6348
rect 1460 6317 1494 6328
rect 1495 6317 1506 6333
rect 1552 6324 1568 6340
rect 1575 6338 1605 6390
rect 1639 6386 1640 6393
rect 1624 6378 1640 6386
rect 1611 6346 1624 6365
rect 1639 6346 1669 6362
rect 1611 6330 1685 6346
rect 1611 6328 1624 6330
rect 1639 6328 1673 6330
rect 1276 6306 1289 6308
rect 1304 6306 1338 6308
rect 1276 6290 1338 6306
rect 1382 6301 1398 6304
rect 1460 6301 1490 6312
rect 1538 6308 1584 6324
rect 1611 6312 1685 6328
rect 1538 6306 1572 6308
rect 1537 6290 1584 6306
rect 1611 6290 1624 6312
rect 1639 6290 1669 6312
rect 1696 6290 1697 6306
rect 1712 6290 1725 6450
rect 1755 6346 1768 6450
rect 1813 6428 1814 6438
rect 1829 6428 1842 6438
rect 1813 6424 1842 6428
rect 1847 6424 1877 6450
rect 1895 6436 1911 6438
rect 1983 6436 2036 6450
rect 1984 6434 2048 6436
rect 2091 6434 2106 6450
rect 2155 6447 2185 6450
rect 2155 6444 2191 6447
rect 2121 6436 2137 6438
rect 1895 6424 1910 6428
rect 1813 6422 1910 6424
rect 1938 6422 2106 6434
rect 2122 6424 2137 6428
rect 2155 6425 2194 6444
rect 2213 6438 2220 6439
rect 2219 6431 2220 6438
rect 2203 6428 2204 6431
rect 2219 6428 2232 6431
rect 2155 6424 2185 6425
rect 2194 6424 2200 6425
rect 2203 6424 2232 6428
rect 2122 6423 2232 6424
rect 2122 6422 2238 6423
rect 1797 6414 1848 6422
rect 1797 6402 1822 6414
rect 1829 6402 1848 6414
rect 1879 6414 1929 6422
rect 1879 6406 1895 6414
rect 1902 6412 1929 6414
rect 1938 6412 2159 6422
rect 1902 6402 2159 6412
rect 2188 6414 2238 6422
rect 2188 6405 2204 6414
rect 1797 6394 1848 6402
rect 1895 6394 2159 6402
rect 2185 6402 2204 6405
rect 2211 6402 2238 6414
rect 2185 6394 2238 6402
rect 1813 6386 1814 6394
rect 1829 6386 1842 6394
rect 1813 6378 1829 6386
rect 1810 6371 1829 6374
rect 1810 6362 1832 6371
rect 1783 6352 1832 6362
rect 1783 6346 1813 6352
rect 1832 6347 1837 6352
rect 1755 6330 1829 6346
rect 1847 6338 1877 6394
rect 1912 6384 2120 6394
rect 2155 6390 2200 6394
rect 2203 6393 2204 6394
rect 2219 6393 2232 6394
rect 1938 6354 2127 6384
rect 1953 6351 2127 6354
rect 1946 6348 2127 6351
rect 1755 6328 1768 6330
rect 1783 6328 1817 6330
rect 1755 6312 1829 6328
rect 1856 6324 1869 6338
rect 1884 6324 1900 6340
rect 1946 6335 1957 6348
rect 1739 6290 1740 6306
rect 1755 6290 1768 6312
rect 1783 6290 1813 6312
rect 1856 6308 1918 6324
rect 1946 6317 1957 6333
rect 1962 6328 1972 6348
rect 1982 6328 1996 6348
rect 1999 6335 2008 6348
rect 2024 6335 2033 6348
rect 1962 6317 1996 6328
rect 1999 6317 2008 6333
rect 2024 6317 2033 6333
rect 2040 6328 2050 6348
rect 2060 6328 2074 6348
rect 2075 6335 2086 6348
rect 2040 6317 2074 6328
rect 2075 6317 2086 6333
rect 2132 6324 2148 6340
rect 2155 6338 2185 6390
rect 2219 6386 2220 6393
rect 2204 6378 2220 6386
rect 2191 6346 2204 6365
rect 2219 6346 2249 6362
rect 2191 6330 2265 6346
rect 2191 6328 2204 6330
rect 2219 6328 2253 6330
rect 1856 6306 1869 6308
rect 1884 6306 1918 6308
rect 1856 6290 1918 6306
rect 1962 6301 1978 6304
rect 2040 6301 2070 6312
rect 2118 6308 2164 6324
rect 2191 6312 2265 6328
rect 2118 6306 2152 6308
rect 2117 6290 2164 6306
rect 2191 6290 2204 6312
rect 2219 6290 2249 6312
rect 2276 6290 2277 6306
rect 2292 6290 2305 6450
rect 2335 6346 2348 6450
rect 2393 6428 2394 6438
rect 2409 6428 2422 6438
rect 2393 6424 2422 6428
rect 2427 6424 2457 6450
rect 2475 6436 2491 6438
rect 2563 6436 2616 6450
rect 2564 6434 2628 6436
rect 2671 6434 2686 6450
rect 2735 6447 2765 6450
rect 2735 6444 2771 6447
rect 2701 6436 2717 6438
rect 2475 6424 2490 6428
rect 2393 6422 2490 6424
rect 2518 6422 2686 6434
rect 2702 6424 2717 6428
rect 2735 6425 2774 6444
rect 2793 6438 2800 6439
rect 2799 6431 2800 6438
rect 2783 6428 2784 6431
rect 2799 6428 2812 6431
rect 2735 6424 2765 6425
rect 2774 6424 2780 6425
rect 2783 6424 2812 6428
rect 2702 6423 2812 6424
rect 2702 6422 2818 6423
rect 2377 6414 2428 6422
rect 2377 6402 2402 6414
rect 2409 6402 2428 6414
rect 2459 6414 2509 6422
rect 2459 6406 2475 6414
rect 2482 6412 2509 6414
rect 2518 6412 2739 6422
rect 2482 6402 2739 6412
rect 2768 6414 2818 6422
rect 2768 6405 2784 6414
rect 2377 6394 2428 6402
rect 2475 6394 2739 6402
rect 2765 6402 2784 6405
rect 2791 6402 2818 6414
rect 2765 6394 2818 6402
rect 2393 6386 2394 6394
rect 2409 6386 2422 6394
rect 2393 6378 2409 6386
rect 2390 6371 2409 6374
rect 2390 6362 2412 6371
rect 2363 6352 2412 6362
rect 2363 6346 2393 6352
rect 2412 6347 2417 6352
rect 2335 6330 2409 6346
rect 2427 6338 2457 6394
rect 2492 6384 2700 6394
rect 2735 6390 2780 6394
rect 2783 6393 2784 6394
rect 2799 6393 2812 6394
rect 2518 6354 2707 6384
rect 2533 6351 2707 6354
rect 2526 6348 2707 6351
rect 2335 6328 2348 6330
rect 2363 6328 2397 6330
rect 2335 6312 2409 6328
rect 2436 6324 2449 6338
rect 2464 6324 2480 6340
rect 2526 6335 2537 6348
rect 2319 6290 2320 6306
rect 2335 6290 2348 6312
rect 2363 6290 2393 6312
rect 2436 6308 2498 6324
rect 2526 6317 2537 6333
rect 2542 6328 2552 6348
rect 2562 6328 2576 6348
rect 2579 6335 2588 6348
rect 2604 6335 2613 6348
rect 2542 6317 2576 6328
rect 2579 6317 2588 6333
rect 2604 6317 2613 6333
rect 2620 6328 2630 6348
rect 2640 6328 2654 6348
rect 2655 6335 2666 6348
rect 2620 6317 2654 6328
rect 2655 6317 2666 6333
rect 2712 6324 2728 6340
rect 2735 6338 2765 6390
rect 2799 6386 2800 6393
rect 2784 6378 2800 6386
rect 2771 6346 2784 6365
rect 2799 6346 2829 6362
rect 2771 6330 2845 6346
rect 2771 6328 2784 6330
rect 2799 6328 2833 6330
rect 2436 6306 2449 6308
rect 2464 6306 2498 6308
rect 2436 6290 2498 6306
rect 2542 6301 2558 6304
rect 2620 6301 2650 6312
rect 2698 6308 2744 6324
rect 2771 6312 2845 6328
rect 2698 6306 2732 6308
rect 2697 6290 2744 6306
rect 2771 6290 2784 6312
rect 2799 6290 2829 6312
rect 2856 6290 2857 6306
rect 2872 6290 2885 6450
rect 2915 6346 2928 6450
rect 2973 6428 2974 6438
rect 2989 6428 3002 6438
rect 2973 6424 3002 6428
rect 3007 6424 3037 6450
rect 3055 6436 3071 6438
rect 3143 6436 3196 6450
rect 3144 6434 3208 6436
rect 3251 6434 3266 6450
rect 3315 6447 3345 6450
rect 3315 6444 3351 6447
rect 3281 6436 3297 6438
rect 3055 6424 3070 6428
rect 2973 6422 3070 6424
rect 3098 6422 3266 6434
rect 3282 6424 3297 6428
rect 3315 6425 3354 6444
rect 3373 6438 3380 6439
rect 3379 6431 3380 6438
rect 3363 6428 3364 6431
rect 3379 6428 3392 6431
rect 3315 6424 3345 6425
rect 3354 6424 3360 6425
rect 3363 6424 3392 6428
rect 3282 6423 3392 6424
rect 3282 6422 3398 6423
rect 2957 6414 3008 6422
rect 2957 6402 2982 6414
rect 2989 6402 3008 6414
rect 3039 6414 3089 6422
rect 3039 6406 3055 6414
rect 3062 6412 3089 6414
rect 3098 6412 3319 6422
rect 3062 6402 3319 6412
rect 3348 6414 3398 6422
rect 3348 6405 3364 6414
rect 2957 6394 3008 6402
rect 3055 6394 3319 6402
rect 3345 6402 3364 6405
rect 3371 6402 3398 6414
rect 3345 6394 3398 6402
rect 2973 6386 2974 6394
rect 2989 6386 3002 6394
rect 2973 6378 2989 6386
rect 2970 6371 2989 6374
rect 2970 6362 2992 6371
rect 2943 6352 2992 6362
rect 2943 6346 2973 6352
rect 2992 6347 2997 6352
rect 2915 6330 2989 6346
rect 3007 6338 3037 6394
rect 3072 6384 3280 6394
rect 3315 6390 3360 6394
rect 3363 6393 3364 6394
rect 3379 6393 3392 6394
rect 3098 6354 3287 6384
rect 3113 6351 3287 6354
rect 3106 6348 3287 6351
rect 2915 6328 2928 6330
rect 2943 6328 2977 6330
rect 2915 6312 2989 6328
rect 3016 6324 3029 6338
rect 3044 6324 3060 6340
rect 3106 6335 3117 6348
rect 2899 6290 2900 6306
rect 2915 6290 2928 6312
rect 2943 6290 2973 6312
rect 3016 6308 3078 6324
rect 3106 6317 3117 6333
rect 3122 6328 3132 6348
rect 3142 6328 3156 6348
rect 3159 6335 3168 6348
rect 3184 6335 3193 6348
rect 3122 6317 3156 6328
rect 3159 6317 3168 6333
rect 3184 6317 3193 6333
rect 3200 6328 3210 6348
rect 3220 6328 3234 6348
rect 3235 6335 3246 6348
rect 3200 6317 3234 6328
rect 3235 6317 3246 6333
rect 3292 6324 3308 6340
rect 3315 6338 3345 6390
rect 3379 6386 3380 6393
rect 3364 6378 3380 6386
rect 3351 6346 3364 6365
rect 3379 6346 3409 6362
rect 3351 6330 3425 6346
rect 3351 6328 3364 6330
rect 3379 6328 3413 6330
rect 3016 6306 3029 6308
rect 3044 6306 3078 6308
rect 3016 6290 3078 6306
rect 3122 6301 3138 6304
rect 3200 6301 3230 6312
rect 3278 6308 3324 6324
rect 3351 6312 3425 6328
rect 3278 6306 3312 6308
rect 3277 6290 3324 6306
rect 3351 6290 3364 6312
rect 3379 6290 3409 6312
rect 3436 6290 3437 6306
rect 3452 6290 3465 6450
rect 3495 6346 3508 6450
rect 3553 6428 3554 6438
rect 3569 6428 3582 6438
rect 3553 6424 3582 6428
rect 3587 6424 3617 6450
rect 3635 6436 3651 6438
rect 3723 6436 3776 6450
rect 3724 6434 3788 6436
rect 3831 6434 3846 6450
rect 3895 6447 3925 6450
rect 3895 6444 3931 6447
rect 3861 6436 3877 6438
rect 3635 6424 3650 6428
rect 3553 6422 3650 6424
rect 3678 6422 3846 6434
rect 3862 6424 3877 6428
rect 3895 6425 3934 6444
rect 3953 6438 3960 6439
rect 3959 6431 3960 6438
rect 3943 6428 3944 6431
rect 3959 6428 3972 6431
rect 3895 6424 3925 6425
rect 3934 6424 3940 6425
rect 3943 6424 3972 6428
rect 3862 6423 3972 6424
rect 3862 6422 3978 6423
rect 3537 6414 3588 6422
rect 3537 6402 3562 6414
rect 3569 6402 3588 6414
rect 3619 6414 3669 6422
rect 3619 6406 3635 6414
rect 3642 6412 3669 6414
rect 3678 6412 3899 6422
rect 3642 6402 3899 6412
rect 3928 6414 3978 6422
rect 3928 6405 3944 6414
rect 3537 6394 3588 6402
rect 3635 6394 3899 6402
rect 3925 6402 3944 6405
rect 3951 6402 3978 6414
rect 3925 6394 3978 6402
rect 3553 6386 3554 6394
rect 3569 6386 3582 6394
rect 3553 6378 3569 6386
rect 3550 6371 3569 6374
rect 3550 6362 3572 6371
rect 3523 6352 3572 6362
rect 3523 6346 3553 6352
rect 3572 6347 3577 6352
rect 3495 6330 3569 6346
rect 3587 6338 3617 6394
rect 3652 6384 3860 6394
rect 3895 6390 3940 6394
rect 3943 6393 3944 6394
rect 3959 6393 3972 6394
rect 3678 6354 3867 6384
rect 3693 6351 3867 6354
rect 3686 6348 3867 6351
rect 3495 6328 3508 6330
rect 3523 6328 3557 6330
rect 3495 6312 3569 6328
rect 3596 6324 3609 6338
rect 3624 6324 3640 6340
rect 3686 6335 3697 6348
rect 3479 6290 3480 6306
rect 3495 6290 3508 6312
rect 3523 6290 3553 6312
rect 3596 6308 3658 6324
rect 3686 6317 3697 6333
rect 3702 6328 3712 6348
rect 3722 6328 3736 6348
rect 3739 6335 3748 6348
rect 3764 6335 3773 6348
rect 3702 6317 3736 6328
rect 3739 6317 3748 6333
rect 3764 6317 3773 6333
rect 3780 6328 3790 6348
rect 3800 6328 3814 6348
rect 3815 6335 3826 6348
rect 3780 6317 3814 6328
rect 3815 6317 3826 6333
rect 3872 6324 3888 6340
rect 3895 6338 3925 6390
rect 3959 6386 3960 6393
rect 3944 6378 3960 6386
rect 3931 6346 3944 6365
rect 3959 6346 3989 6362
rect 3931 6330 4005 6346
rect 3931 6328 3944 6330
rect 3959 6328 3993 6330
rect 3596 6306 3609 6308
rect 3624 6306 3658 6308
rect 3596 6290 3658 6306
rect 3702 6301 3718 6304
rect 3780 6301 3810 6312
rect 3858 6308 3904 6324
rect 3931 6312 4005 6328
rect 3858 6306 3892 6308
rect 3857 6290 3904 6306
rect 3931 6290 3944 6312
rect 3959 6290 3989 6312
rect 4016 6290 4017 6306
rect 4032 6290 4045 6450
rect 4075 6346 4088 6450
rect 4133 6428 4134 6438
rect 4149 6428 4162 6438
rect 4133 6424 4162 6428
rect 4167 6424 4197 6450
rect 4215 6436 4231 6438
rect 4303 6436 4356 6450
rect 4304 6434 4368 6436
rect 4411 6434 4426 6450
rect 4475 6447 4505 6450
rect 4475 6444 4511 6447
rect 4441 6436 4457 6438
rect 4215 6424 4230 6428
rect 4133 6422 4230 6424
rect 4258 6422 4426 6434
rect 4442 6424 4457 6428
rect 4475 6425 4514 6444
rect 4533 6438 4540 6439
rect 4539 6431 4540 6438
rect 4523 6428 4524 6431
rect 4539 6428 4552 6431
rect 4475 6424 4505 6425
rect 4514 6424 4520 6425
rect 4523 6424 4552 6428
rect 4442 6423 4552 6424
rect 4442 6422 4558 6423
rect 4117 6414 4168 6422
rect 4117 6402 4142 6414
rect 4149 6402 4168 6414
rect 4199 6414 4249 6422
rect 4199 6406 4215 6414
rect 4222 6412 4249 6414
rect 4258 6412 4479 6422
rect 4222 6402 4479 6412
rect 4508 6414 4558 6422
rect 4508 6405 4524 6414
rect 4117 6394 4168 6402
rect 4215 6394 4479 6402
rect 4505 6402 4524 6405
rect 4531 6402 4558 6414
rect 4505 6394 4558 6402
rect 4133 6386 4134 6394
rect 4149 6386 4162 6394
rect 4133 6378 4149 6386
rect 4130 6371 4149 6374
rect 4130 6362 4152 6371
rect 4103 6352 4152 6362
rect 4103 6346 4133 6352
rect 4152 6347 4157 6352
rect 4075 6330 4149 6346
rect 4167 6338 4197 6394
rect 4232 6384 4440 6394
rect 4475 6390 4520 6394
rect 4523 6393 4524 6394
rect 4539 6393 4552 6394
rect 4258 6354 4447 6384
rect 4273 6351 4447 6354
rect 4266 6348 4447 6351
rect 4075 6328 4088 6330
rect 4103 6328 4137 6330
rect 4075 6312 4149 6328
rect 4176 6324 4189 6338
rect 4204 6324 4220 6340
rect 4266 6335 4277 6348
rect 4059 6290 4060 6306
rect 4075 6290 4088 6312
rect 4103 6290 4133 6312
rect 4176 6308 4238 6324
rect 4266 6317 4277 6333
rect 4282 6328 4292 6348
rect 4302 6328 4316 6348
rect 4319 6335 4328 6348
rect 4344 6335 4353 6348
rect 4282 6317 4316 6328
rect 4319 6317 4328 6333
rect 4344 6317 4353 6333
rect 4360 6328 4370 6348
rect 4380 6328 4394 6348
rect 4395 6335 4406 6348
rect 4360 6317 4394 6328
rect 4395 6317 4406 6333
rect 4452 6324 4468 6340
rect 4475 6338 4505 6390
rect 4539 6386 4540 6393
rect 4524 6378 4540 6386
rect 4511 6346 4524 6365
rect 4539 6346 4569 6362
rect 4511 6330 4585 6346
rect 4511 6328 4524 6330
rect 4539 6328 4573 6330
rect 4176 6306 4189 6308
rect 4204 6306 4238 6308
rect 4176 6290 4238 6306
rect 4282 6301 4298 6304
rect 4360 6301 4390 6312
rect 4438 6308 4484 6324
rect 4511 6312 4585 6328
rect 4438 6306 4472 6308
rect 4437 6290 4484 6306
rect 4511 6290 4524 6312
rect 4539 6290 4569 6312
rect 4596 6290 4597 6306
rect 4612 6290 4625 6450
rect -7 6282 34 6290
rect -7 6256 8 6282
rect 15 6256 34 6282
rect 98 6278 160 6290
rect 172 6278 247 6290
rect 305 6278 380 6290
rect 392 6278 423 6290
rect 429 6278 464 6290
rect 98 6276 260 6278
rect -7 6248 34 6256
rect 116 6252 129 6276
rect 144 6274 159 6276
rect -1 6238 0 6248
rect 15 6238 28 6248
rect 43 6238 73 6252
rect 116 6238 159 6252
rect 183 6249 190 6256
rect 193 6252 260 6276
rect 292 6276 464 6278
rect 262 6254 290 6258
rect 292 6254 372 6276
rect 393 6274 408 6276
rect 262 6252 372 6254
rect 193 6248 372 6252
rect 166 6238 196 6248
rect 198 6238 351 6248
rect 359 6238 389 6248
rect 393 6238 423 6252
rect 451 6238 464 6276
rect 536 6282 571 6290
rect 536 6256 537 6282
rect 544 6256 571 6282
rect 479 6238 509 6252
rect 536 6248 571 6256
rect 573 6282 614 6290
rect 573 6256 588 6282
rect 595 6256 614 6282
rect 678 6278 740 6290
rect 752 6278 827 6290
rect 885 6278 960 6290
rect 972 6278 1003 6290
rect 1009 6278 1044 6290
rect 678 6276 840 6278
rect 573 6248 614 6256
rect 696 6252 709 6276
rect 724 6274 739 6276
rect 536 6238 537 6248
rect 552 6238 565 6248
rect 579 6238 580 6248
rect 595 6238 608 6248
rect 623 6238 653 6252
rect 696 6238 739 6252
rect 763 6249 770 6256
rect 773 6252 840 6276
rect 872 6276 1044 6278
rect 842 6254 870 6258
rect 872 6254 952 6276
rect 973 6274 988 6276
rect 842 6252 952 6254
rect 773 6248 952 6252
rect 746 6238 776 6248
rect 778 6238 931 6248
rect 939 6238 969 6248
rect 973 6238 1003 6252
rect 1031 6238 1044 6276
rect 1116 6282 1151 6290
rect 1116 6256 1117 6282
rect 1124 6256 1151 6282
rect 1059 6238 1089 6252
rect 1116 6248 1151 6256
rect 1153 6282 1194 6290
rect 1153 6256 1168 6282
rect 1175 6256 1194 6282
rect 1258 6278 1320 6290
rect 1332 6278 1407 6290
rect 1465 6278 1540 6290
rect 1552 6278 1583 6290
rect 1589 6278 1624 6290
rect 1258 6276 1420 6278
rect 1153 6248 1194 6256
rect 1276 6252 1289 6276
rect 1304 6274 1319 6276
rect 1116 6238 1117 6248
rect 1132 6238 1145 6248
rect 1159 6238 1160 6248
rect 1175 6238 1188 6248
rect 1203 6238 1233 6252
rect 1276 6238 1319 6252
rect 1343 6249 1350 6256
rect 1353 6252 1420 6276
rect 1452 6276 1624 6278
rect 1422 6254 1450 6258
rect 1452 6254 1532 6276
rect 1553 6274 1568 6276
rect 1422 6252 1532 6254
rect 1353 6248 1532 6252
rect 1326 6238 1356 6248
rect 1358 6238 1511 6248
rect 1519 6238 1549 6248
rect 1553 6238 1583 6252
rect 1611 6238 1624 6276
rect 1696 6282 1731 6290
rect 1696 6256 1697 6282
rect 1704 6256 1731 6282
rect 1639 6238 1669 6252
rect 1696 6248 1731 6256
rect 1733 6282 1774 6290
rect 1733 6256 1748 6282
rect 1755 6256 1774 6282
rect 1838 6278 1900 6290
rect 1912 6278 1987 6290
rect 2045 6278 2120 6290
rect 2132 6278 2163 6290
rect 2169 6278 2204 6290
rect 1838 6276 2000 6278
rect 1733 6248 1774 6256
rect 1856 6252 1869 6276
rect 1884 6274 1899 6276
rect 1696 6238 1697 6248
rect 1712 6238 1725 6248
rect 1739 6238 1740 6248
rect 1755 6238 1768 6248
rect 1783 6238 1813 6252
rect 1856 6238 1899 6252
rect 1923 6249 1930 6256
rect 1933 6252 2000 6276
rect 2032 6276 2204 6278
rect 2002 6254 2030 6258
rect 2032 6254 2112 6276
rect 2133 6274 2148 6276
rect 2002 6252 2112 6254
rect 1933 6248 2112 6252
rect 1906 6238 1936 6248
rect 1938 6238 2091 6248
rect 2099 6238 2129 6248
rect 2133 6238 2163 6252
rect 2191 6238 2204 6276
rect 2276 6282 2311 6290
rect 2276 6256 2277 6282
rect 2284 6256 2311 6282
rect 2219 6238 2249 6252
rect 2276 6248 2311 6256
rect 2313 6282 2354 6290
rect 2313 6256 2328 6282
rect 2335 6256 2354 6282
rect 2418 6278 2480 6290
rect 2492 6278 2567 6290
rect 2625 6278 2700 6290
rect 2712 6278 2743 6290
rect 2749 6278 2784 6290
rect 2418 6276 2580 6278
rect 2313 6248 2354 6256
rect 2436 6252 2449 6276
rect 2464 6274 2479 6276
rect 2276 6238 2277 6248
rect 2292 6238 2305 6248
rect 2319 6238 2320 6248
rect 2335 6238 2348 6248
rect 2363 6238 2393 6252
rect 2436 6238 2479 6252
rect 2503 6249 2510 6256
rect 2513 6252 2580 6276
rect 2612 6276 2784 6278
rect 2582 6254 2610 6258
rect 2612 6254 2692 6276
rect 2713 6274 2728 6276
rect 2582 6252 2692 6254
rect 2513 6248 2692 6252
rect 2486 6238 2516 6248
rect 2518 6238 2671 6248
rect 2679 6238 2709 6248
rect 2713 6238 2743 6252
rect 2771 6238 2784 6276
rect 2856 6282 2891 6290
rect 2856 6256 2857 6282
rect 2864 6256 2891 6282
rect 2799 6238 2829 6252
rect 2856 6248 2891 6256
rect 2893 6282 2934 6290
rect 2893 6256 2908 6282
rect 2915 6256 2934 6282
rect 2998 6278 3060 6290
rect 3072 6278 3147 6290
rect 3205 6278 3280 6290
rect 3292 6278 3323 6290
rect 3329 6278 3364 6290
rect 2998 6276 3160 6278
rect 2893 6248 2934 6256
rect 3016 6252 3029 6276
rect 3044 6274 3059 6276
rect 2856 6238 2857 6248
rect 2872 6238 2885 6248
rect 2899 6238 2900 6248
rect 2915 6238 2928 6248
rect 2943 6238 2973 6252
rect 3016 6238 3059 6252
rect 3083 6249 3090 6256
rect 3093 6252 3160 6276
rect 3192 6276 3364 6278
rect 3162 6254 3190 6258
rect 3192 6254 3272 6276
rect 3293 6274 3308 6276
rect 3162 6252 3272 6254
rect 3093 6248 3272 6252
rect 3066 6238 3096 6248
rect 3098 6238 3251 6248
rect 3259 6238 3289 6248
rect 3293 6238 3323 6252
rect 3351 6238 3364 6276
rect 3436 6282 3471 6290
rect 3436 6256 3437 6282
rect 3444 6256 3471 6282
rect 3379 6238 3409 6252
rect 3436 6248 3471 6256
rect 3473 6282 3514 6290
rect 3473 6256 3488 6282
rect 3495 6256 3514 6282
rect 3578 6278 3640 6290
rect 3652 6278 3727 6290
rect 3785 6278 3860 6290
rect 3872 6278 3903 6290
rect 3909 6278 3944 6290
rect 3578 6276 3740 6278
rect 3473 6248 3514 6256
rect 3596 6252 3609 6276
rect 3624 6274 3639 6276
rect 3436 6238 3437 6248
rect 3452 6238 3465 6248
rect 3479 6238 3480 6248
rect 3495 6238 3508 6248
rect 3523 6238 3553 6252
rect 3596 6238 3639 6252
rect 3663 6249 3670 6256
rect 3673 6252 3740 6276
rect 3772 6276 3944 6278
rect 3742 6254 3770 6258
rect 3772 6254 3852 6276
rect 3873 6274 3888 6276
rect 3742 6252 3852 6254
rect 3673 6248 3852 6252
rect 3646 6238 3676 6248
rect 3678 6238 3831 6248
rect 3839 6238 3869 6248
rect 3873 6238 3903 6252
rect 3931 6238 3944 6276
rect 4016 6282 4051 6290
rect 4016 6256 4017 6282
rect 4024 6256 4051 6282
rect 3959 6238 3989 6252
rect 4016 6248 4051 6256
rect 4053 6282 4094 6290
rect 4053 6256 4068 6282
rect 4075 6256 4094 6282
rect 4158 6278 4220 6290
rect 4232 6278 4307 6290
rect 4365 6278 4440 6290
rect 4452 6278 4483 6290
rect 4489 6278 4524 6290
rect 4158 6276 4320 6278
rect 4053 6248 4094 6256
rect 4176 6252 4189 6276
rect 4204 6274 4219 6276
rect 4016 6238 4017 6248
rect 4032 6238 4045 6248
rect 4059 6238 4060 6248
rect 4075 6238 4088 6248
rect 4103 6238 4133 6252
rect 4176 6238 4219 6252
rect 4243 6249 4250 6256
rect 4253 6252 4320 6276
rect 4352 6276 4524 6278
rect 4322 6254 4350 6258
rect 4352 6254 4432 6276
rect 4453 6274 4468 6276
rect 4322 6252 4432 6254
rect 4253 6248 4432 6252
rect 4226 6238 4256 6248
rect 4258 6238 4411 6248
rect 4419 6238 4449 6248
rect 4453 6238 4483 6252
rect 4511 6238 4524 6276
rect 4596 6282 4631 6290
rect 4596 6256 4597 6282
rect 4604 6256 4631 6282
rect 4539 6238 4569 6252
rect 4596 6248 4631 6256
rect 4596 6238 4597 6248
rect 4612 6238 4625 6248
rect -1 6232 4625 6238
rect 0 6224 4625 6232
rect 15 6194 28 6224
rect 43 6206 73 6224
rect 116 6210 130 6224
rect 166 6210 386 6224
rect 117 6208 130 6210
rect 83 6196 98 6208
rect 80 6194 102 6196
rect 107 6194 137 6208
rect 198 6206 351 6210
rect 180 6194 372 6206
rect 415 6194 445 6208
rect 451 6194 464 6224
rect 479 6206 509 6224
rect 552 6194 565 6224
rect 595 6194 608 6224
rect 623 6206 653 6224
rect 696 6210 710 6224
rect 746 6210 966 6224
rect 697 6208 710 6210
rect 663 6196 678 6208
rect 660 6194 682 6196
rect 687 6194 717 6208
rect 778 6206 931 6210
rect 760 6194 952 6206
rect 995 6194 1025 6208
rect 1031 6194 1044 6224
rect 1059 6206 1089 6224
rect 1132 6194 1145 6224
rect 1175 6194 1188 6224
rect 1203 6206 1233 6224
rect 1276 6210 1290 6224
rect 1326 6210 1546 6224
rect 1277 6208 1290 6210
rect 1243 6196 1258 6208
rect 1240 6194 1262 6196
rect 1267 6194 1297 6208
rect 1358 6206 1511 6210
rect 1340 6194 1532 6206
rect 1575 6194 1605 6208
rect 1611 6194 1624 6224
rect 1639 6206 1669 6224
rect 1712 6194 1725 6224
rect 1755 6194 1768 6224
rect 1783 6206 1813 6224
rect 1856 6210 1870 6224
rect 1906 6210 2126 6224
rect 1857 6208 1870 6210
rect 1823 6196 1838 6208
rect 1820 6194 1842 6196
rect 1847 6194 1877 6208
rect 1938 6206 2091 6210
rect 1920 6194 2112 6206
rect 2155 6194 2185 6208
rect 2191 6194 2204 6224
rect 2219 6206 2249 6224
rect 2292 6194 2305 6224
rect 2335 6194 2348 6224
rect 2363 6206 2393 6224
rect 2436 6210 2450 6224
rect 2486 6210 2706 6224
rect 2437 6208 2450 6210
rect 2403 6196 2418 6208
rect 2400 6194 2422 6196
rect 2427 6194 2457 6208
rect 2518 6206 2671 6210
rect 2500 6194 2692 6206
rect 2735 6194 2765 6208
rect 2771 6194 2784 6224
rect 2799 6206 2829 6224
rect 2872 6194 2885 6224
rect 2915 6194 2928 6224
rect 2943 6206 2973 6224
rect 3016 6210 3030 6224
rect 3066 6210 3286 6224
rect 3017 6208 3030 6210
rect 2983 6196 2998 6208
rect 2980 6194 3002 6196
rect 3007 6194 3037 6208
rect 3098 6206 3251 6210
rect 3080 6194 3272 6206
rect 3315 6194 3345 6208
rect 3351 6194 3364 6224
rect 3379 6206 3409 6224
rect 3452 6194 3465 6224
rect 3495 6194 3508 6224
rect 3523 6206 3553 6224
rect 3596 6210 3610 6224
rect 3646 6210 3866 6224
rect 3597 6208 3610 6210
rect 3563 6196 3578 6208
rect 3560 6194 3582 6196
rect 3587 6194 3617 6208
rect 3678 6206 3831 6210
rect 3660 6194 3852 6206
rect 3895 6194 3925 6208
rect 3931 6194 3944 6224
rect 3959 6206 3989 6224
rect 4032 6194 4045 6224
rect 4075 6194 4088 6224
rect 4103 6206 4133 6224
rect 4176 6210 4190 6224
rect 4226 6210 4446 6224
rect 4177 6208 4190 6210
rect 4143 6196 4158 6208
rect 4140 6194 4162 6196
rect 4167 6194 4197 6208
rect 4258 6206 4411 6210
rect 4240 6194 4432 6206
rect 4475 6194 4505 6208
rect 4511 6194 4524 6224
rect 4539 6206 4569 6224
rect 4612 6194 4625 6224
rect 0 6180 4625 6194
rect 15 6076 28 6180
rect 73 6158 74 6168
rect 89 6158 102 6168
rect 73 6154 102 6158
rect 107 6154 137 6180
rect 155 6166 171 6168
rect 243 6166 296 6180
rect 244 6164 308 6166
rect 351 6164 366 6180
rect 415 6177 445 6180
rect 415 6174 451 6177
rect 381 6166 397 6168
rect 155 6154 170 6158
rect 73 6152 170 6154
rect 198 6152 366 6164
rect 382 6154 397 6158
rect 415 6155 454 6174
rect 473 6168 480 6169
rect 479 6161 480 6168
rect 463 6158 464 6161
rect 479 6158 492 6161
rect 415 6154 445 6155
rect 454 6154 460 6155
rect 463 6154 492 6158
rect 382 6153 492 6154
rect 382 6152 498 6153
rect 57 6144 108 6152
rect 57 6132 82 6144
rect 89 6132 108 6144
rect 139 6144 189 6152
rect 139 6136 155 6144
rect 162 6142 189 6144
rect 198 6142 419 6152
rect 162 6132 419 6142
rect 448 6144 498 6152
rect 448 6135 464 6144
rect 57 6124 108 6132
rect 155 6124 419 6132
rect 445 6132 464 6135
rect 471 6132 498 6144
rect 445 6124 498 6132
rect 73 6116 74 6124
rect 89 6116 102 6124
rect 73 6108 89 6116
rect 70 6101 89 6104
rect 70 6092 92 6101
rect 43 6082 92 6092
rect 43 6076 73 6082
rect 92 6077 97 6082
rect 15 6060 89 6076
rect 107 6068 137 6124
rect 172 6114 380 6124
rect 415 6120 460 6124
rect 463 6123 464 6124
rect 479 6123 492 6124
rect 198 6084 387 6114
rect 213 6081 387 6084
rect 206 6078 387 6081
rect 15 6058 28 6060
rect 43 6058 77 6060
rect 15 6042 89 6058
rect 116 6054 129 6068
rect 144 6054 160 6070
rect 206 6065 217 6078
rect -1 6020 0 6036
rect 15 6020 28 6042
rect 43 6020 73 6042
rect 116 6038 178 6054
rect 206 6047 217 6063
rect 222 6058 232 6078
rect 242 6058 256 6078
rect 259 6065 268 6078
rect 284 6065 293 6078
rect 222 6047 256 6058
rect 259 6047 268 6063
rect 284 6047 293 6063
rect 300 6058 310 6078
rect 320 6058 334 6078
rect 335 6065 346 6078
rect 300 6047 334 6058
rect 335 6047 346 6063
rect 392 6054 408 6070
rect 415 6068 445 6120
rect 479 6116 480 6123
rect 464 6108 480 6116
rect 451 6076 464 6095
rect 479 6076 509 6092
rect 451 6060 525 6076
rect 451 6058 464 6060
rect 479 6058 513 6060
rect 116 6036 129 6038
rect 144 6036 178 6038
rect 116 6020 178 6036
rect 222 6031 238 6034
rect 300 6031 330 6042
rect 378 6038 424 6054
rect 451 6042 525 6058
rect 378 6036 412 6038
rect 377 6020 424 6036
rect 451 6020 464 6042
rect 479 6020 509 6042
rect 536 6020 537 6036
rect 552 6020 565 6180
rect 595 6076 608 6180
rect 653 6158 654 6168
rect 669 6158 682 6168
rect 653 6154 682 6158
rect 687 6154 717 6180
rect 735 6166 751 6168
rect 823 6166 876 6180
rect 824 6164 888 6166
rect 931 6164 946 6180
rect 995 6177 1025 6180
rect 995 6174 1031 6177
rect 961 6166 977 6168
rect 735 6154 750 6158
rect 653 6152 750 6154
rect 778 6152 946 6164
rect 962 6154 977 6158
rect 995 6155 1034 6174
rect 1053 6168 1060 6169
rect 1059 6161 1060 6168
rect 1043 6158 1044 6161
rect 1059 6158 1072 6161
rect 995 6154 1025 6155
rect 1034 6154 1040 6155
rect 1043 6154 1072 6158
rect 962 6153 1072 6154
rect 962 6152 1078 6153
rect 637 6144 688 6152
rect 637 6132 662 6144
rect 669 6132 688 6144
rect 719 6144 769 6152
rect 719 6136 735 6144
rect 742 6142 769 6144
rect 778 6142 999 6152
rect 742 6132 999 6142
rect 1028 6144 1078 6152
rect 1028 6135 1044 6144
rect 637 6124 688 6132
rect 735 6124 999 6132
rect 1025 6132 1044 6135
rect 1051 6132 1078 6144
rect 1025 6124 1078 6132
rect 653 6116 654 6124
rect 669 6116 682 6124
rect 653 6108 669 6116
rect 650 6101 669 6104
rect 650 6092 672 6101
rect 623 6082 672 6092
rect 623 6076 653 6082
rect 672 6077 677 6082
rect 595 6060 669 6076
rect 687 6068 717 6124
rect 752 6114 960 6124
rect 995 6120 1040 6124
rect 1043 6123 1044 6124
rect 1059 6123 1072 6124
rect 778 6084 967 6114
rect 793 6081 967 6084
rect 786 6078 967 6081
rect 595 6058 608 6060
rect 623 6058 657 6060
rect 595 6042 669 6058
rect 696 6054 709 6068
rect 724 6054 740 6070
rect 786 6065 797 6078
rect 579 6020 580 6036
rect 595 6020 608 6042
rect 623 6020 653 6042
rect 696 6038 758 6054
rect 786 6047 797 6063
rect 802 6058 812 6078
rect 822 6058 836 6078
rect 839 6065 848 6078
rect 864 6065 873 6078
rect 802 6047 836 6058
rect 839 6047 848 6063
rect 864 6047 873 6063
rect 880 6058 890 6078
rect 900 6058 914 6078
rect 915 6065 926 6078
rect 880 6047 914 6058
rect 915 6047 926 6063
rect 972 6054 988 6070
rect 995 6068 1025 6120
rect 1059 6116 1060 6123
rect 1044 6108 1060 6116
rect 1031 6076 1044 6095
rect 1059 6076 1089 6092
rect 1031 6060 1105 6076
rect 1031 6058 1044 6060
rect 1059 6058 1093 6060
rect 696 6036 709 6038
rect 724 6036 758 6038
rect 696 6020 758 6036
rect 802 6031 818 6034
rect 880 6031 910 6042
rect 958 6038 1004 6054
rect 1031 6042 1105 6058
rect 958 6036 992 6038
rect 957 6020 1004 6036
rect 1031 6020 1044 6042
rect 1059 6020 1089 6042
rect 1116 6020 1117 6036
rect 1132 6020 1145 6180
rect 1175 6076 1188 6180
rect 1233 6158 1234 6168
rect 1249 6158 1262 6168
rect 1233 6154 1262 6158
rect 1267 6154 1297 6180
rect 1315 6166 1331 6168
rect 1403 6166 1456 6180
rect 1404 6164 1468 6166
rect 1511 6164 1526 6180
rect 1575 6177 1605 6180
rect 1575 6174 1611 6177
rect 1541 6166 1557 6168
rect 1315 6154 1330 6158
rect 1233 6152 1330 6154
rect 1358 6152 1526 6164
rect 1542 6154 1557 6158
rect 1575 6155 1614 6174
rect 1633 6168 1640 6169
rect 1639 6161 1640 6168
rect 1623 6158 1624 6161
rect 1639 6158 1652 6161
rect 1575 6154 1605 6155
rect 1614 6154 1620 6155
rect 1623 6154 1652 6158
rect 1542 6153 1652 6154
rect 1542 6152 1658 6153
rect 1217 6144 1268 6152
rect 1217 6132 1242 6144
rect 1249 6132 1268 6144
rect 1299 6144 1349 6152
rect 1299 6136 1315 6144
rect 1322 6142 1349 6144
rect 1358 6142 1579 6152
rect 1322 6132 1579 6142
rect 1608 6144 1658 6152
rect 1608 6135 1624 6144
rect 1217 6124 1268 6132
rect 1315 6124 1579 6132
rect 1605 6132 1624 6135
rect 1631 6132 1658 6144
rect 1605 6124 1658 6132
rect 1233 6116 1234 6124
rect 1249 6116 1262 6124
rect 1233 6108 1249 6116
rect 1230 6101 1249 6104
rect 1230 6092 1252 6101
rect 1203 6082 1252 6092
rect 1203 6076 1233 6082
rect 1252 6077 1257 6082
rect 1175 6060 1249 6076
rect 1267 6068 1297 6124
rect 1332 6114 1540 6124
rect 1575 6120 1620 6124
rect 1623 6123 1624 6124
rect 1639 6123 1652 6124
rect 1358 6084 1547 6114
rect 1373 6081 1547 6084
rect 1366 6078 1547 6081
rect 1175 6058 1188 6060
rect 1203 6058 1237 6060
rect 1175 6042 1249 6058
rect 1276 6054 1289 6068
rect 1304 6054 1320 6070
rect 1366 6065 1377 6078
rect 1159 6020 1160 6036
rect 1175 6020 1188 6042
rect 1203 6020 1233 6042
rect 1276 6038 1338 6054
rect 1366 6047 1377 6063
rect 1382 6058 1392 6078
rect 1402 6058 1416 6078
rect 1419 6065 1428 6078
rect 1444 6065 1453 6078
rect 1382 6047 1416 6058
rect 1419 6047 1428 6063
rect 1444 6047 1453 6063
rect 1460 6058 1470 6078
rect 1480 6058 1494 6078
rect 1495 6065 1506 6078
rect 1460 6047 1494 6058
rect 1495 6047 1506 6063
rect 1552 6054 1568 6070
rect 1575 6068 1605 6120
rect 1639 6116 1640 6123
rect 1624 6108 1640 6116
rect 1611 6076 1624 6095
rect 1639 6076 1669 6092
rect 1611 6060 1685 6076
rect 1611 6058 1624 6060
rect 1639 6058 1673 6060
rect 1276 6036 1289 6038
rect 1304 6036 1338 6038
rect 1276 6020 1338 6036
rect 1382 6031 1398 6034
rect 1460 6031 1490 6042
rect 1538 6038 1584 6054
rect 1611 6042 1685 6058
rect 1538 6036 1572 6038
rect 1537 6020 1584 6036
rect 1611 6020 1624 6042
rect 1639 6020 1669 6042
rect 1696 6020 1697 6036
rect 1712 6020 1725 6180
rect 1755 6076 1768 6180
rect 1813 6158 1814 6168
rect 1829 6158 1842 6168
rect 1813 6154 1842 6158
rect 1847 6154 1877 6180
rect 1895 6166 1911 6168
rect 1983 6166 2036 6180
rect 1984 6164 2048 6166
rect 2091 6164 2106 6180
rect 2155 6177 2185 6180
rect 2155 6174 2191 6177
rect 2121 6166 2137 6168
rect 1895 6154 1910 6158
rect 1813 6152 1910 6154
rect 1938 6152 2106 6164
rect 2122 6154 2137 6158
rect 2155 6155 2194 6174
rect 2213 6168 2220 6169
rect 2219 6161 2220 6168
rect 2203 6158 2204 6161
rect 2219 6158 2232 6161
rect 2155 6154 2185 6155
rect 2194 6154 2200 6155
rect 2203 6154 2232 6158
rect 2122 6153 2232 6154
rect 2122 6152 2238 6153
rect 1797 6144 1848 6152
rect 1797 6132 1822 6144
rect 1829 6132 1848 6144
rect 1879 6144 1929 6152
rect 1879 6136 1895 6144
rect 1902 6142 1929 6144
rect 1938 6142 2159 6152
rect 1902 6132 2159 6142
rect 2188 6144 2238 6152
rect 2188 6135 2204 6144
rect 1797 6124 1848 6132
rect 1895 6124 2159 6132
rect 2185 6132 2204 6135
rect 2211 6132 2238 6144
rect 2185 6124 2238 6132
rect 1813 6116 1814 6124
rect 1829 6116 1842 6124
rect 1813 6108 1829 6116
rect 1810 6101 1829 6104
rect 1810 6092 1832 6101
rect 1783 6082 1832 6092
rect 1783 6076 1813 6082
rect 1832 6077 1837 6082
rect 1755 6060 1829 6076
rect 1847 6068 1877 6124
rect 1912 6114 2120 6124
rect 2155 6120 2200 6124
rect 2203 6123 2204 6124
rect 2219 6123 2232 6124
rect 1938 6084 2127 6114
rect 1953 6081 2127 6084
rect 1946 6078 2127 6081
rect 1755 6058 1768 6060
rect 1783 6058 1817 6060
rect 1755 6042 1829 6058
rect 1856 6054 1869 6068
rect 1884 6054 1900 6070
rect 1946 6065 1957 6078
rect 1739 6020 1740 6036
rect 1755 6020 1768 6042
rect 1783 6020 1813 6042
rect 1856 6038 1918 6054
rect 1946 6047 1957 6063
rect 1962 6058 1972 6078
rect 1982 6058 1996 6078
rect 1999 6065 2008 6078
rect 2024 6065 2033 6078
rect 1962 6047 1996 6058
rect 1999 6047 2008 6063
rect 2024 6047 2033 6063
rect 2040 6058 2050 6078
rect 2060 6058 2074 6078
rect 2075 6065 2086 6078
rect 2040 6047 2074 6058
rect 2075 6047 2086 6063
rect 2132 6054 2148 6070
rect 2155 6068 2185 6120
rect 2219 6116 2220 6123
rect 2204 6108 2220 6116
rect 2191 6076 2204 6095
rect 2219 6076 2249 6092
rect 2191 6060 2265 6076
rect 2191 6058 2204 6060
rect 2219 6058 2253 6060
rect 1856 6036 1869 6038
rect 1884 6036 1918 6038
rect 1856 6020 1918 6036
rect 1962 6031 1978 6034
rect 2040 6031 2070 6042
rect 2118 6038 2164 6054
rect 2191 6042 2265 6058
rect 2118 6036 2152 6038
rect 2117 6020 2164 6036
rect 2191 6020 2204 6042
rect 2219 6020 2249 6042
rect 2276 6020 2277 6036
rect 2292 6020 2305 6180
rect 2335 6076 2348 6180
rect 2393 6158 2394 6168
rect 2409 6158 2422 6168
rect 2393 6154 2422 6158
rect 2427 6154 2457 6180
rect 2475 6166 2491 6168
rect 2563 6166 2616 6180
rect 2564 6164 2628 6166
rect 2671 6164 2686 6180
rect 2735 6177 2765 6180
rect 2735 6174 2771 6177
rect 2701 6166 2717 6168
rect 2475 6154 2490 6158
rect 2393 6152 2490 6154
rect 2518 6152 2686 6164
rect 2702 6154 2717 6158
rect 2735 6155 2774 6174
rect 2793 6168 2800 6169
rect 2799 6161 2800 6168
rect 2783 6158 2784 6161
rect 2799 6158 2812 6161
rect 2735 6154 2765 6155
rect 2774 6154 2780 6155
rect 2783 6154 2812 6158
rect 2702 6153 2812 6154
rect 2702 6152 2818 6153
rect 2377 6144 2428 6152
rect 2377 6132 2402 6144
rect 2409 6132 2428 6144
rect 2459 6144 2509 6152
rect 2459 6136 2475 6144
rect 2482 6142 2509 6144
rect 2518 6142 2739 6152
rect 2482 6132 2739 6142
rect 2768 6144 2818 6152
rect 2768 6135 2784 6144
rect 2377 6124 2428 6132
rect 2475 6124 2739 6132
rect 2765 6132 2784 6135
rect 2791 6132 2818 6144
rect 2765 6124 2818 6132
rect 2393 6116 2394 6124
rect 2409 6116 2422 6124
rect 2393 6108 2409 6116
rect 2390 6101 2409 6104
rect 2390 6092 2412 6101
rect 2363 6082 2412 6092
rect 2363 6076 2393 6082
rect 2412 6077 2417 6082
rect 2335 6060 2409 6076
rect 2427 6068 2457 6124
rect 2492 6114 2700 6124
rect 2735 6120 2780 6124
rect 2783 6123 2784 6124
rect 2799 6123 2812 6124
rect 2518 6084 2707 6114
rect 2533 6081 2707 6084
rect 2526 6078 2707 6081
rect 2335 6058 2348 6060
rect 2363 6058 2397 6060
rect 2335 6042 2409 6058
rect 2436 6054 2449 6068
rect 2464 6054 2480 6070
rect 2526 6065 2537 6078
rect 2319 6020 2320 6036
rect 2335 6020 2348 6042
rect 2363 6020 2393 6042
rect 2436 6038 2498 6054
rect 2526 6047 2537 6063
rect 2542 6058 2552 6078
rect 2562 6058 2576 6078
rect 2579 6065 2588 6078
rect 2604 6065 2613 6078
rect 2542 6047 2576 6058
rect 2579 6047 2588 6063
rect 2604 6047 2613 6063
rect 2620 6058 2630 6078
rect 2640 6058 2654 6078
rect 2655 6065 2666 6078
rect 2620 6047 2654 6058
rect 2655 6047 2666 6063
rect 2712 6054 2728 6070
rect 2735 6068 2765 6120
rect 2799 6116 2800 6123
rect 2784 6108 2800 6116
rect 2771 6076 2784 6095
rect 2799 6076 2829 6092
rect 2771 6060 2845 6076
rect 2771 6058 2784 6060
rect 2799 6058 2833 6060
rect 2436 6036 2449 6038
rect 2464 6036 2498 6038
rect 2436 6020 2498 6036
rect 2542 6031 2558 6034
rect 2620 6031 2650 6042
rect 2698 6038 2744 6054
rect 2771 6042 2845 6058
rect 2698 6036 2732 6038
rect 2697 6020 2744 6036
rect 2771 6020 2784 6042
rect 2799 6020 2829 6042
rect 2856 6020 2857 6036
rect 2872 6020 2885 6180
rect 2915 6076 2928 6180
rect 2973 6158 2974 6168
rect 2989 6158 3002 6168
rect 2973 6154 3002 6158
rect 3007 6154 3037 6180
rect 3055 6166 3071 6168
rect 3143 6166 3196 6180
rect 3144 6164 3208 6166
rect 3251 6164 3266 6180
rect 3315 6177 3345 6180
rect 3315 6174 3351 6177
rect 3281 6166 3297 6168
rect 3055 6154 3070 6158
rect 2973 6152 3070 6154
rect 3098 6152 3266 6164
rect 3282 6154 3297 6158
rect 3315 6155 3354 6174
rect 3373 6168 3380 6169
rect 3379 6161 3380 6168
rect 3363 6158 3364 6161
rect 3379 6158 3392 6161
rect 3315 6154 3345 6155
rect 3354 6154 3360 6155
rect 3363 6154 3392 6158
rect 3282 6153 3392 6154
rect 3282 6152 3398 6153
rect 2957 6144 3008 6152
rect 2957 6132 2982 6144
rect 2989 6132 3008 6144
rect 3039 6144 3089 6152
rect 3039 6136 3055 6144
rect 3062 6142 3089 6144
rect 3098 6142 3319 6152
rect 3062 6132 3319 6142
rect 3348 6144 3398 6152
rect 3348 6135 3364 6144
rect 2957 6124 3008 6132
rect 3055 6124 3319 6132
rect 3345 6132 3364 6135
rect 3371 6132 3398 6144
rect 3345 6124 3398 6132
rect 2973 6116 2974 6124
rect 2989 6116 3002 6124
rect 2973 6108 2989 6116
rect 2970 6101 2989 6104
rect 2970 6092 2992 6101
rect 2943 6082 2992 6092
rect 2943 6076 2973 6082
rect 2992 6077 2997 6082
rect 2915 6060 2989 6076
rect 3007 6068 3037 6124
rect 3072 6114 3280 6124
rect 3315 6120 3360 6124
rect 3363 6123 3364 6124
rect 3379 6123 3392 6124
rect 3098 6084 3287 6114
rect 3113 6081 3287 6084
rect 3106 6078 3287 6081
rect 2915 6058 2928 6060
rect 2943 6058 2977 6060
rect 2915 6042 2989 6058
rect 3016 6054 3029 6068
rect 3044 6054 3060 6070
rect 3106 6065 3117 6078
rect 2899 6020 2900 6036
rect 2915 6020 2928 6042
rect 2943 6020 2973 6042
rect 3016 6038 3078 6054
rect 3106 6047 3117 6063
rect 3122 6058 3132 6078
rect 3142 6058 3156 6078
rect 3159 6065 3168 6078
rect 3184 6065 3193 6078
rect 3122 6047 3156 6058
rect 3159 6047 3168 6063
rect 3184 6047 3193 6063
rect 3200 6058 3210 6078
rect 3220 6058 3234 6078
rect 3235 6065 3246 6078
rect 3200 6047 3234 6058
rect 3235 6047 3246 6063
rect 3292 6054 3308 6070
rect 3315 6068 3345 6120
rect 3379 6116 3380 6123
rect 3364 6108 3380 6116
rect 3351 6076 3364 6095
rect 3379 6076 3409 6092
rect 3351 6060 3425 6076
rect 3351 6058 3364 6060
rect 3379 6058 3413 6060
rect 3016 6036 3029 6038
rect 3044 6036 3078 6038
rect 3016 6020 3078 6036
rect 3122 6031 3138 6034
rect 3200 6031 3230 6042
rect 3278 6038 3324 6054
rect 3351 6042 3425 6058
rect 3278 6036 3312 6038
rect 3277 6020 3324 6036
rect 3351 6020 3364 6042
rect 3379 6020 3409 6042
rect 3436 6020 3437 6036
rect 3452 6020 3465 6180
rect 3495 6076 3508 6180
rect 3553 6158 3554 6168
rect 3569 6158 3582 6168
rect 3553 6154 3582 6158
rect 3587 6154 3617 6180
rect 3635 6166 3651 6168
rect 3723 6166 3776 6180
rect 3724 6164 3788 6166
rect 3831 6164 3846 6180
rect 3895 6177 3925 6180
rect 3895 6174 3931 6177
rect 3861 6166 3877 6168
rect 3635 6154 3650 6158
rect 3553 6152 3650 6154
rect 3678 6152 3846 6164
rect 3862 6154 3877 6158
rect 3895 6155 3934 6174
rect 3953 6168 3960 6169
rect 3959 6161 3960 6168
rect 3943 6158 3944 6161
rect 3959 6158 3972 6161
rect 3895 6154 3925 6155
rect 3934 6154 3940 6155
rect 3943 6154 3972 6158
rect 3862 6153 3972 6154
rect 3862 6152 3978 6153
rect 3537 6144 3588 6152
rect 3537 6132 3562 6144
rect 3569 6132 3588 6144
rect 3619 6144 3669 6152
rect 3619 6136 3635 6144
rect 3642 6142 3669 6144
rect 3678 6142 3899 6152
rect 3642 6132 3899 6142
rect 3928 6144 3978 6152
rect 3928 6135 3944 6144
rect 3537 6124 3588 6132
rect 3635 6124 3899 6132
rect 3925 6132 3944 6135
rect 3951 6132 3978 6144
rect 3925 6124 3978 6132
rect 3553 6116 3554 6124
rect 3569 6116 3582 6124
rect 3553 6108 3569 6116
rect 3550 6101 3569 6104
rect 3550 6092 3572 6101
rect 3523 6082 3572 6092
rect 3523 6076 3553 6082
rect 3572 6077 3577 6082
rect 3495 6060 3569 6076
rect 3587 6068 3617 6124
rect 3652 6114 3860 6124
rect 3895 6120 3940 6124
rect 3943 6123 3944 6124
rect 3959 6123 3972 6124
rect 3678 6084 3867 6114
rect 3693 6081 3867 6084
rect 3686 6078 3867 6081
rect 3495 6058 3508 6060
rect 3523 6058 3557 6060
rect 3495 6042 3569 6058
rect 3596 6054 3609 6068
rect 3624 6054 3640 6070
rect 3686 6065 3697 6078
rect 3479 6020 3480 6036
rect 3495 6020 3508 6042
rect 3523 6020 3553 6042
rect 3596 6038 3658 6054
rect 3686 6047 3697 6063
rect 3702 6058 3712 6078
rect 3722 6058 3736 6078
rect 3739 6065 3748 6078
rect 3764 6065 3773 6078
rect 3702 6047 3736 6058
rect 3739 6047 3748 6063
rect 3764 6047 3773 6063
rect 3780 6058 3790 6078
rect 3800 6058 3814 6078
rect 3815 6065 3826 6078
rect 3780 6047 3814 6058
rect 3815 6047 3826 6063
rect 3872 6054 3888 6070
rect 3895 6068 3925 6120
rect 3959 6116 3960 6123
rect 3944 6108 3960 6116
rect 3931 6076 3944 6095
rect 3959 6076 3989 6092
rect 3931 6060 4005 6076
rect 3931 6058 3944 6060
rect 3959 6058 3993 6060
rect 3596 6036 3609 6038
rect 3624 6036 3658 6038
rect 3596 6020 3658 6036
rect 3702 6031 3718 6034
rect 3780 6031 3810 6042
rect 3858 6038 3904 6054
rect 3931 6042 4005 6058
rect 3858 6036 3892 6038
rect 3857 6020 3904 6036
rect 3931 6020 3944 6042
rect 3959 6020 3989 6042
rect 4016 6020 4017 6036
rect 4032 6020 4045 6180
rect 4075 6076 4088 6180
rect 4133 6158 4134 6168
rect 4149 6158 4162 6168
rect 4133 6154 4162 6158
rect 4167 6154 4197 6180
rect 4215 6166 4231 6168
rect 4303 6166 4356 6180
rect 4304 6164 4368 6166
rect 4411 6164 4426 6180
rect 4475 6177 4505 6180
rect 4475 6174 4511 6177
rect 4441 6166 4457 6168
rect 4215 6154 4230 6158
rect 4133 6152 4230 6154
rect 4258 6152 4426 6164
rect 4442 6154 4457 6158
rect 4475 6155 4514 6174
rect 4533 6168 4540 6169
rect 4539 6161 4540 6168
rect 4523 6158 4524 6161
rect 4539 6158 4552 6161
rect 4475 6154 4505 6155
rect 4514 6154 4520 6155
rect 4523 6154 4552 6158
rect 4442 6153 4552 6154
rect 4442 6152 4558 6153
rect 4117 6144 4168 6152
rect 4117 6132 4142 6144
rect 4149 6132 4168 6144
rect 4199 6144 4249 6152
rect 4199 6136 4215 6144
rect 4222 6142 4249 6144
rect 4258 6142 4479 6152
rect 4222 6132 4479 6142
rect 4508 6144 4558 6152
rect 4508 6135 4524 6144
rect 4117 6124 4168 6132
rect 4215 6124 4479 6132
rect 4505 6132 4524 6135
rect 4531 6132 4558 6144
rect 4505 6124 4558 6132
rect 4133 6116 4134 6124
rect 4149 6116 4162 6124
rect 4133 6108 4149 6116
rect 4130 6101 4149 6104
rect 4130 6092 4152 6101
rect 4103 6082 4152 6092
rect 4103 6076 4133 6082
rect 4152 6077 4157 6082
rect 4075 6060 4149 6076
rect 4167 6068 4197 6124
rect 4232 6114 4440 6124
rect 4475 6120 4520 6124
rect 4523 6123 4524 6124
rect 4539 6123 4552 6124
rect 4258 6084 4447 6114
rect 4273 6081 4447 6084
rect 4266 6078 4447 6081
rect 4075 6058 4088 6060
rect 4103 6058 4137 6060
rect 4075 6042 4149 6058
rect 4176 6054 4189 6068
rect 4204 6054 4220 6070
rect 4266 6065 4277 6078
rect 4059 6020 4060 6036
rect 4075 6020 4088 6042
rect 4103 6020 4133 6042
rect 4176 6038 4238 6054
rect 4266 6047 4277 6063
rect 4282 6058 4292 6078
rect 4302 6058 4316 6078
rect 4319 6065 4328 6078
rect 4344 6065 4353 6078
rect 4282 6047 4316 6058
rect 4319 6047 4328 6063
rect 4344 6047 4353 6063
rect 4360 6058 4370 6078
rect 4380 6058 4394 6078
rect 4395 6065 4406 6078
rect 4360 6047 4394 6058
rect 4395 6047 4406 6063
rect 4452 6054 4468 6070
rect 4475 6068 4505 6120
rect 4539 6116 4540 6123
rect 4524 6108 4540 6116
rect 4511 6076 4524 6095
rect 4539 6076 4569 6092
rect 4511 6060 4585 6076
rect 4511 6058 4524 6060
rect 4539 6058 4573 6060
rect 4176 6036 4189 6038
rect 4204 6036 4238 6038
rect 4176 6020 4238 6036
rect 4282 6031 4298 6034
rect 4360 6031 4390 6042
rect 4438 6038 4484 6054
rect 4511 6042 4585 6058
rect 4438 6036 4472 6038
rect 4437 6020 4484 6036
rect 4511 6020 4524 6042
rect 4539 6020 4569 6042
rect 4596 6020 4597 6036
rect 4612 6020 4625 6180
rect -7 6012 34 6020
rect -7 5986 8 6012
rect 15 5986 34 6012
rect 98 6008 160 6020
rect 172 6008 247 6020
rect 305 6008 380 6020
rect 392 6008 423 6020
rect 429 6008 464 6020
rect 98 6006 260 6008
rect -7 5978 34 5986
rect 116 5982 129 6006
rect 144 6004 159 6006
rect -1 5968 0 5978
rect 15 5968 28 5978
rect 43 5968 73 5982
rect 116 5968 159 5982
rect 183 5979 190 5986
rect 193 5982 260 6006
rect 292 6006 464 6008
rect 262 5984 290 5988
rect 292 5984 372 6006
rect 393 6004 408 6006
rect 262 5982 372 5984
rect 193 5978 372 5982
rect 166 5968 196 5978
rect 198 5968 351 5978
rect 359 5968 389 5978
rect 393 5968 423 5982
rect 451 5968 464 6006
rect 536 6012 571 6020
rect 536 5986 537 6012
rect 544 5986 571 6012
rect 479 5968 509 5982
rect 536 5978 571 5986
rect 573 6012 614 6020
rect 573 5986 588 6012
rect 595 5986 614 6012
rect 678 6008 740 6020
rect 752 6008 827 6020
rect 885 6008 960 6020
rect 972 6008 1003 6020
rect 1009 6008 1044 6020
rect 678 6006 840 6008
rect 573 5978 614 5986
rect 696 5982 709 6006
rect 724 6004 739 6006
rect 536 5968 537 5978
rect 552 5968 565 5978
rect 579 5968 580 5978
rect 595 5968 608 5978
rect 623 5968 653 5982
rect 696 5968 739 5982
rect 763 5979 770 5986
rect 773 5982 840 6006
rect 872 6006 1044 6008
rect 842 5984 870 5988
rect 872 5984 952 6006
rect 973 6004 988 6006
rect 842 5982 952 5984
rect 773 5978 952 5982
rect 746 5968 776 5978
rect 778 5968 931 5978
rect 939 5968 969 5978
rect 973 5968 1003 5982
rect 1031 5968 1044 6006
rect 1116 6012 1151 6020
rect 1116 5986 1117 6012
rect 1124 5986 1151 6012
rect 1059 5968 1089 5982
rect 1116 5978 1151 5986
rect 1153 6012 1194 6020
rect 1153 5986 1168 6012
rect 1175 5986 1194 6012
rect 1258 6008 1320 6020
rect 1332 6008 1407 6020
rect 1465 6008 1540 6020
rect 1552 6008 1583 6020
rect 1589 6008 1624 6020
rect 1258 6006 1420 6008
rect 1153 5978 1194 5986
rect 1276 5982 1289 6006
rect 1304 6004 1319 6006
rect 1116 5968 1117 5978
rect 1132 5968 1145 5978
rect 1159 5968 1160 5978
rect 1175 5968 1188 5978
rect 1203 5968 1233 5982
rect 1276 5968 1319 5982
rect 1343 5979 1350 5986
rect 1353 5982 1420 6006
rect 1452 6006 1624 6008
rect 1422 5984 1450 5988
rect 1452 5984 1532 6006
rect 1553 6004 1568 6006
rect 1422 5982 1532 5984
rect 1353 5978 1532 5982
rect 1326 5968 1356 5978
rect 1358 5968 1511 5978
rect 1519 5968 1549 5978
rect 1553 5968 1583 5982
rect 1611 5968 1624 6006
rect 1696 6012 1731 6020
rect 1696 5986 1697 6012
rect 1704 5986 1731 6012
rect 1639 5968 1669 5982
rect 1696 5978 1731 5986
rect 1733 6012 1774 6020
rect 1733 5986 1748 6012
rect 1755 5986 1774 6012
rect 1838 6008 1900 6020
rect 1912 6008 1987 6020
rect 2045 6008 2120 6020
rect 2132 6008 2163 6020
rect 2169 6008 2204 6020
rect 1838 6006 2000 6008
rect 1733 5978 1774 5986
rect 1856 5982 1869 6006
rect 1884 6004 1899 6006
rect 1696 5968 1697 5978
rect 1712 5968 1725 5978
rect 1739 5968 1740 5978
rect 1755 5968 1768 5978
rect 1783 5968 1813 5982
rect 1856 5968 1899 5982
rect 1923 5979 1930 5986
rect 1933 5982 2000 6006
rect 2032 6006 2204 6008
rect 2002 5984 2030 5988
rect 2032 5984 2112 6006
rect 2133 6004 2148 6006
rect 2002 5982 2112 5984
rect 1933 5978 2112 5982
rect 1906 5968 1936 5978
rect 1938 5968 2091 5978
rect 2099 5968 2129 5978
rect 2133 5968 2163 5982
rect 2191 5968 2204 6006
rect 2276 6012 2311 6020
rect 2276 5986 2277 6012
rect 2284 5986 2311 6012
rect 2219 5968 2249 5982
rect 2276 5978 2311 5986
rect 2313 6012 2354 6020
rect 2313 5986 2328 6012
rect 2335 5986 2354 6012
rect 2418 6008 2480 6020
rect 2492 6008 2567 6020
rect 2625 6008 2700 6020
rect 2712 6008 2743 6020
rect 2749 6008 2784 6020
rect 2418 6006 2580 6008
rect 2313 5978 2354 5986
rect 2436 5982 2449 6006
rect 2464 6004 2479 6006
rect 2276 5968 2277 5978
rect 2292 5968 2305 5978
rect 2319 5968 2320 5978
rect 2335 5968 2348 5978
rect 2363 5968 2393 5982
rect 2436 5968 2479 5982
rect 2503 5979 2510 5986
rect 2513 5982 2580 6006
rect 2612 6006 2784 6008
rect 2582 5984 2610 5988
rect 2612 5984 2692 6006
rect 2713 6004 2728 6006
rect 2582 5982 2692 5984
rect 2513 5978 2692 5982
rect 2486 5968 2516 5978
rect 2518 5968 2671 5978
rect 2679 5968 2709 5978
rect 2713 5968 2743 5982
rect 2771 5968 2784 6006
rect 2856 6012 2891 6020
rect 2856 5986 2857 6012
rect 2864 5986 2891 6012
rect 2799 5968 2829 5982
rect 2856 5978 2891 5986
rect 2893 6012 2934 6020
rect 2893 5986 2908 6012
rect 2915 5986 2934 6012
rect 2998 6008 3060 6020
rect 3072 6008 3147 6020
rect 3205 6008 3280 6020
rect 3292 6008 3323 6020
rect 3329 6008 3364 6020
rect 2998 6006 3160 6008
rect 2893 5978 2934 5986
rect 3016 5982 3029 6006
rect 3044 6004 3059 6006
rect 2856 5968 2857 5978
rect 2872 5968 2885 5978
rect 2899 5968 2900 5978
rect 2915 5968 2928 5978
rect 2943 5968 2973 5982
rect 3016 5968 3059 5982
rect 3083 5979 3090 5986
rect 3093 5982 3160 6006
rect 3192 6006 3364 6008
rect 3162 5984 3190 5988
rect 3192 5984 3272 6006
rect 3293 6004 3308 6006
rect 3162 5982 3272 5984
rect 3093 5978 3272 5982
rect 3066 5968 3096 5978
rect 3098 5968 3251 5978
rect 3259 5968 3289 5978
rect 3293 5968 3323 5982
rect 3351 5968 3364 6006
rect 3436 6012 3471 6020
rect 3436 5986 3437 6012
rect 3444 5986 3471 6012
rect 3379 5968 3409 5982
rect 3436 5978 3471 5986
rect 3473 6012 3514 6020
rect 3473 5986 3488 6012
rect 3495 5986 3514 6012
rect 3578 6008 3640 6020
rect 3652 6008 3727 6020
rect 3785 6008 3860 6020
rect 3872 6008 3903 6020
rect 3909 6008 3944 6020
rect 3578 6006 3740 6008
rect 3473 5978 3514 5986
rect 3596 5982 3609 6006
rect 3624 6004 3639 6006
rect 3436 5968 3437 5978
rect 3452 5968 3465 5978
rect 3479 5968 3480 5978
rect 3495 5968 3508 5978
rect 3523 5968 3553 5982
rect 3596 5968 3639 5982
rect 3663 5979 3670 5986
rect 3673 5982 3740 6006
rect 3772 6006 3944 6008
rect 3742 5984 3770 5988
rect 3772 5984 3852 6006
rect 3873 6004 3888 6006
rect 3742 5982 3852 5984
rect 3673 5978 3852 5982
rect 3646 5968 3676 5978
rect 3678 5968 3831 5978
rect 3839 5968 3869 5978
rect 3873 5968 3903 5982
rect 3931 5968 3944 6006
rect 4016 6012 4051 6020
rect 4016 5986 4017 6012
rect 4024 5986 4051 6012
rect 3959 5968 3989 5982
rect 4016 5978 4051 5986
rect 4053 6012 4094 6020
rect 4053 5986 4068 6012
rect 4075 5986 4094 6012
rect 4158 6008 4220 6020
rect 4232 6008 4307 6020
rect 4365 6008 4440 6020
rect 4452 6008 4483 6020
rect 4489 6008 4524 6020
rect 4158 6006 4320 6008
rect 4053 5978 4094 5986
rect 4176 5982 4189 6006
rect 4204 6004 4219 6006
rect 4016 5968 4017 5978
rect 4032 5968 4045 5978
rect 4059 5968 4060 5978
rect 4075 5968 4088 5978
rect 4103 5968 4133 5982
rect 4176 5968 4219 5982
rect 4243 5979 4250 5986
rect 4253 5982 4320 6006
rect 4352 6006 4524 6008
rect 4322 5984 4350 5988
rect 4352 5984 4432 6006
rect 4453 6004 4468 6006
rect 4322 5982 4432 5984
rect 4253 5978 4432 5982
rect 4226 5968 4256 5978
rect 4258 5968 4411 5978
rect 4419 5968 4449 5978
rect 4453 5968 4483 5982
rect 4511 5968 4524 6006
rect 4596 6012 4631 6020
rect 4596 5986 4597 6012
rect 4604 5986 4631 6012
rect 4539 5968 4569 5982
rect 4596 5978 4631 5986
rect 4596 5968 4597 5978
rect 4612 5968 4625 5978
rect -1 5962 4625 5968
rect 0 5954 4625 5962
rect 15 5924 28 5954
rect 43 5936 73 5954
rect 116 5940 130 5954
rect 166 5940 386 5954
rect 117 5938 130 5940
rect 83 5926 98 5938
rect 80 5924 102 5926
rect 107 5924 137 5938
rect 198 5936 351 5940
rect 180 5924 372 5936
rect 415 5924 445 5938
rect 451 5924 464 5954
rect 479 5936 509 5954
rect 552 5924 565 5954
rect 595 5924 608 5954
rect 623 5936 653 5954
rect 696 5940 710 5954
rect 746 5940 966 5954
rect 697 5938 710 5940
rect 663 5926 678 5938
rect 660 5924 682 5926
rect 687 5924 717 5938
rect 778 5936 931 5940
rect 760 5924 952 5936
rect 995 5924 1025 5938
rect 1031 5924 1044 5954
rect 1059 5936 1089 5954
rect 1132 5924 1145 5954
rect 1175 5924 1188 5954
rect 1203 5936 1233 5954
rect 1276 5940 1290 5954
rect 1326 5940 1546 5954
rect 1277 5938 1290 5940
rect 1243 5926 1258 5938
rect 1240 5924 1262 5926
rect 1267 5924 1297 5938
rect 1358 5936 1511 5940
rect 1340 5924 1532 5936
rect 1575 5924 1605 5938
rect 1611 5924 1624 5954
rect 1639 5936 1669 5954
rect 1712 5924 1725 5954
rect 1755 5924 1768 5954
rect 1783 5936 1813 5954
rect 1856 5940 1870 5954
rect 1906 5940 2126 5954
rect 1857 5938 1870 5940
rect 1823 5926 1838 5938
rect 1820 5924 1842 5926
rect 1847 5924 1877 5938
rect 1938 5936 2091 5940
rect 1920 5924 2112 5936
rect 2155 5924 2185 5938
rect 2191 5924 2204 5954
rect 2219 5936 2249 5954
rect 2292 5924 2305 5954
rect 2335 5924 2348 5954
rect 2363 5936 2393 5954
rect 2436 5940 2450 5954
rect 2486 5940 2706 5954
rect 2437 5938 2450 5940
rect 2403 5926 2418 5938
rect 2400 5924 2422 5926
rect 2427 5924 2457 5938
rect 2518 5936 2671 5940
rect 2500 5924 2692 5936
rect 2735 5924 2765 5938
rect 2771 5924 2784 5954
rect 2799 5936 2829 5954
rect 2872 5924 2885 5954
rect 2915 5924 2928 5954
rect 2943 5936 2973 5954
rect 3016 5940 3030 5954
rect 3066 5940 3286 5954
rect 3017 5938 3030 5940
rect 2983 5926 2998 5938
rect 2980 5924 3002 5926
rect 3007 5924 3037 5938
rect 3098 5936 3251 5940
rect 3080 5924 3272 5936
rect 3315 5924 3345 5938
rect 3351 5924 3364 5954
rect 3379 5936 3409 5954
rect 3452 5924 3465 5954
rect 3495 5924 3508 5954
rect 3523 5936 3553 5954
rect 3596 5940 3610 5954
rect 3646 5940 3866 5954
rect 3597 5938 3610 5940
rect 3563 5926 3578 5938
rect 3560 5924 3582 5926
rect 3587 5924 3617 5938
rect 3678 5936 3831 5940
rect 3660 5924 3852 5936
rect 3895 5924 3925 5938
rect 3931 5924 3944 5954
rect 3959 5936 3989 5954
rect 4032 5924 4045 5954
rect 4075 5924 4088 5954
rect 4103 5936 4133 5954
rect 4176 5940 4190 5954
rect 4226 5940 4446 5954
rect 4177 5938 4190 5940
rect 4143 5926 4158 5938
rect 4140 5924 4162 5926
rect 4167 5924 4197 5938
rect 4258 5936 4411 5940
rect 4240 5924 4432 5936
rect 4475 5924 4505 5938
rect 4511 5924 4524 5954
rect 4539 5936 4569 5954
rect 4612 5924 4625 5954
rect 0 5910 4625 5924
rect 15 5806 28 5910
rect 73 5888 74 5898
rect 89 5888 102 5898
rect 73 5884 102 5888
rect 107 5884 137 5910
rect 155 5896 171 5898
rect 243 5896 296 5910
rect 244 5894 308 5896
rect 351 5894 366 5910
rect 415 5907 445 5910
rect 415 5904 451 5907
rect 381 5896 397 5898
rect 155 5884 170 5888
rect 73 5882 170 5884
rect 198 5882 366 5894
rect 382 5884 397 5888
rect 415 5885 454 5904
rect 473 5898 480 5899
rect 479 5891 480 5898
rect 463 5888 464 5891
rect 479 5888 492 5891
rect 415 5884 445 5885
rect 454 5884 460 5885
rect 463 5884 492 5888
rect 382 5883 492 5884
rect 382 5882 498 5883
rect 57 5874 108 5882
rect 57 5862 82 5874
rect 89 5862 108 5874
rect 139 5874 189 5882
rect 139 5866 155 5874
rect 162 5872 189 5874
rect 198 5872 419 5882
rect 162 5862 419 5872
rect 448 5874 498 5882
rect 448 5865 464 5874
rect 57 5854 108 5862
rect 155 5854 419 5862
rect 445 5862 464 5865
rect 471 5862 498 5874
rect 445 5854 498 5862
rect 73 5846 74 5854
rect 89 5846 102 5854
rect 73 5838 89 5846
rect 70 5831 89 5834
rect 70 5822 92 5831
rect 43 5812 92 5822
rect 43 5806 73 5812
rect 92 5807 97 5812
rect 15 5790 89 5806
rect 107 5798 137 5854
rect 172 5844 380 5854
rect 415 5850 460 5854
rect 463 5853 464 5854
rect 479 5853 492 5854
rect 198 5814 387 5844
rect 213 5811 387 5814
rect 206 5808 387 5811
rect 15 5788 28 5790
rect 43 5788 77 5790
rect 15 5772 89 5788
rect 116 5784 129 5798
rect 144 5784 160 5800
rect 206 5795 217 5808
rect -1 5750 0 5766
rect 15 5750 28 5772
rect 43 5750 73 5772
rect 116 5768 178 5784
rect 206 5777 217 5793
rect 222 5788 232 5808
rect 242 5788 256 5808
rect 259 5795 268 5808
rect 284 5795 293 5808
rect 222 5777 256 5788
rect 259 5777 268 5793
rect 284 5777 293 5793
rect 300 5788 310 5808
rect 320 5788 334 5808
rect 335 5795 346 5808
rect 300 5777 334 5788
rect 335 5777 346 5793
rect 392 5784 408 5800
rect 415 5798 445 5850
rect 479 5846 480 5853
rect 464 5838 480 5846
rect 451 5806 464 5825
rect 479 5806 509 5822
rect 451 5790 525 5806
rect 451 5788 464 5790
rect 479 5788 513 5790
rect 116 5766 129 5768
rect 144 5766 178 5768
rect 116 5750 178 5766
rect 222 5761 238 5764
rect 300 5761 330 5772
rect 378 5768 424 5784
rect 451 5772 525 5788
rect 378 5766 412 5768
rect 377 5750 424 5766
rect 451 5750 464 5772
rect 479 5750 509 5772
rect 536 5750 537 5766
rect 552 5750 565 5910
rect 595 5806 608 5910
rect 653 5888 654 5898
rect 669 5888 682 5898
rect 653 5884 682 5888
rect 687 5884 717 5910
rect 735 5896 751 5898
rect 823 5896 876 5910
rect 824 5894 888 5896
rect 931 5894 946 5910
rect 995 5907 1025 5910
rect 995 5904 1031 5907
rect 961 5896 977 5898
rect 735 5884 750 5888
rect 653 5882 750 5884
rect 778 5882 946 5894
rect 962 5884 977 5888
rect 995 5885 1034 5904
rect 1053 5898 1060 5899
rect 1059 5891 1060 5898
rect 1043 5888 1044 5891
rect 1059 5888 1072 5891
rect 995 5884 1025 5885
rect 1034 5884 1040 5885
rect 1043 5884 1072 5888
rect 962 5883 1072 5884
rect 962 5882 1078 5883
rect 637 5874 688 5882
rect 637 5862 662 5874
rect 669 5862 688 5874
rect 719 5874 769 5882
rect 719 5866 735 5874
rect 742 5872 769 5874
rect 778 5872 999 5882
rect 742 5862 999 5872
rect 1028 5874 1078 5882
rect 1028 5865 1044 5874
rect 637 5854 688 5862
rect 735 5854 999 5862
rect 1025 5862 1044 5865
rect 1051 5862 1078 5874
rect 1025 5854 1078 5862
rect 653 5846 654 5854
rect 669 5846 682 5854
rect 653 5838 669 5846
rect 650 5831 669 5834
rect 650 5822 672 5831
rect 623 5812 672 5822
rect 623 5806 653 5812
rect 672 5807 677 5812
rect 595 5790 669 5806
rect 687 5798 717 5854
rect 752 5844 960 5854
rect 995 5850 1040 5854
rect 1043 5853 1044 5854
rect 1059 5853 1072 5854
rect 778 5814 967 5844
rect 793 5811 967 5814
rect 786 5808 967 5811
rect 595 5788 608 5790
rect 623 5788 657 5790
rect 595 5772 669 5788
rect 696 5784 709 5798
rect 724 5784 740 5800
rect 786 5795 797 5808
rect 579 5750 580 5766
rect 595 5750 608 5772
rect 623 5750 653 5772
rect 696 5768 758 5784
rect 786 5777 797 5793
rect 802 5788 812 5808
rect 822 5788 836 5808
rect 839 5795 848 5808
rect 864 5795 873 5808
rect 802 5777 836 5788
rect 839 5777 848 5793
rect 864 5777 873 5793
rect 880 5788 890 5808
rect 900 5788 914 5808
rect 915 5795 926 5808
rect 880 5777 914 5788
rect 915 5777 926 5793
rect 972 5784 988 5800
rect 995 5798 1025 5850
rect 1059 5846 1060 5853
rect 1044 5838 1060 5846
rect 1031 5806 1044 5825
rect 1059 5806 1089 5822
rect 1031 5790 1105 5806
rect 1031 5788 1044 5790
rect 1059 5788 1093 5790
rect 696 5766 709 5768
rect 724 5766 758 5768
rect 696 5750 758 5766
rect 802 5761 818 5764
rect 880 5761 910 5772
rect 958 5768 1004 5784
rect 1031 5772 1105 5788
rect 958 5766 992 5768
rect 957 5750 1004 5766
rect 1031 5750 1044 5772
rect 1059 5750 1089 5772
rect 1116 5750 1117 5766
rect 1132 5750 1145 5910
rect 1175 5806 1188 5910
rect 1233 5888 1234 5898
rect 1249 5888 1262 5898
rect 1233 5884 1262 5888
rect 1267 5884 1297 5910
rect 1315 5896 1331 5898
rect 1403 5896 1456 5910
rect 1404 5894 1468 5896
rect 1511 5894 1526 5910
rect 1575 5907 1605 5910
rect 1575 5904 1611 5907
rect 1541 5896 1557 5898
rect 1315 5884 1330 5888
rect 1233 5882 1330 5884
rect 1358 5882 1526 5894
rect 1542 5884 1557 5888
rect 1575 5885 1614 5904
rect 1633 5898 1640 5899
rect 1639 5891 1640 5898
rect 1623 5888 1624 5891
rect 1639 5888 1652 5891
rect 1575 5884 1605 5885
rect 1614 5884 1620 5885
rect 1623 5884 1652 5888
rect 1542 5883 1652 5884
rect 1542 5882 1658 5883
rect 1217 5874 1268 5882
rect 1217 5862 1242 5874
rect 1249 5862 1268 5874
rect 1299 5874 1349 5882
rect 1299 5866 1315 5874
rect 1322 5872 1349 5874
rect 1358 5872 1579 5882
rect 1322 5862 1579 5872
rect 1608 5874 1658 5882
rect 1608 5865 1624 5874
rect 1217 5854 1268 5862
rect 1315 5854 1579 5862
rect 1605 5862 1624 5865
rect 1631 5862 1658 5874
rect 1605 5854 1658 5862
rect 1233 5846 1234 5854
rect 1249 5846 1262 5854
rect 1233 5838 1249 5846
rect 1230 5831 1249 5834
rect 1230 5822 1252 5831
rect 1203 5812 1252 5822
rect 1203 5806 1233 5812
rect 1252 5807 1257 5812
rect 1175 5790 1249 5806
rect 1267 5798 1297 5854
rect 1332 5844 1540 5854
rect 1575 5850 1620 5854
rect 1623 5853 1624 5854
rect 1639 5853 1652 5854
rect 1358 5814 1547 5844
rect 1373 5811 1547 5814
rect 1366 5808 1547 5811
rect 1175 5788 1188 5790
rect 1203 5788 1237 5790
rect 1175 5772 1249 5788
rect 1276 5784 1289 5798
rect 1304 5784 1320 5800
rect 1366 5795 1377 5808
rect 1159 5750 1160 5766
rect 1175 5750 1188 5772
rect 1203 5750 1233 5772
rect 1276 5768 1338 5784
rect 1366 5777 1377 5793
rect 1382 5788 1392 5808
rect 1402 5788 1416 5808
rect 1419 5795 1428 5808
rect 1444 5795 1453 5808
rect 1382 5777 1416 5788
rect 1419 5777 1428 5793
rect 1444 5777 1453 5793
rect 1460 5788 1470 5808
rect 1480 5788 1494 5808
rect 1495 5795 1506 5808
rect 1460 5777 1494 5788
rect 1495 5777 1506 5793
rect 1552 5784 1568 5800
rect 1575 5798 1605 5850
rect 1639 5846 1640 5853
rect 1624 5838 1640 5846
rect 1611 5806 1624 5825
rect 1639 5806 1669 5822
rect 1611 5790 1685 5806
rect 1611 5788 1624 5790
rect 1639 5788 1673 5790
rect 1276 5766 1289 5768
rect 1304 5766 1338 5768
rect 1276 5750 1338 5766
rect 1382 5761 1398 5764
rect 1460 5761 1490 5772
rect 1538 5768 1584 5784
rect 1611 5772 1685 5788
rect 1538 5766 1572 5768
rect 1537 5750 1584 5766
rect 1611 5750 1624 5772
rect 1639 5750 1669 5772
rect 1696 5750 1697 5766
rect 1712 5750 1725 5910
rect 1755 5806 1768 5910
rect 1813 5888 1814 5898
rect 1829 5888 1842 5898
rect 1813 5884 1842 5888
rect 1847 5884 1877 5910
rect 1895 5896 1911 5898
rect 1983 5896 2036 5910
rect 1984 5894 2048 5896
rect 2091 5894 2106 5910
rect 2155 5907 2185 5910
rect 2155 5904 2191 5907
rect 2121 5896 2137 5898
rect 1895 5884 1910 5888
rect 1813 5882 1910 5884
rect 1938 5882 2106 5894
rect 2122 5884 2137 5888
rect 2155 5885 2194 5904
rect 2213 5898 2220 5899
rect 2219 5891 2220 5898
rect 2203 5888 2204 5891
rect 2219 5888 2232 5891
rect 2155 5884 2185 5885
rect 2194 5884 2200 5885
rect 2203 5884 2232 5888
rect 2122 5883 2232 5884
rect 2122 5882 2238 5883
rect 1797 5874 1848 5882
rect 1797 5862 1822 5874
rect 1829 5862 1848 5874
rect 1879 5874 1929 5882
rect 1879 5866 1895 5874
rect 1902 5872 1929 5874
rect 1938 5872 2159 5882
rect 1902 5862 2159 5872
rect 2188 5874 2238 5882
rect 2188 5865 2204 5874
rect 1797 5854 1848 5862
rect 1895 5854 2159 5862
rect 2185 5862 2204 5865
rect 2211 5862 2238 5874
rect 2185 5854 2238 5862
rect 1813 5846 1814 5854
rect 1829 5846 1842 5854
rect 1813 5838 1829 5846
rect 1810 5831 1829 5834
rect 1810 5822 1832 5831
rect 1783 5812 1832 5822
rect 1783 5806 1813 5812
rect 1832 5807 1837 5812
rect 1755 5790 1829 5806
rect 1847 5798 1877 5854
rect 1912 5844 2120 5854
rect 2155 5850 2200 5854
rect 2203 5853 2204 5854
rect 2219 5853 2232 5854
rect 1938 5814 2127 5844
rect 1953 5811 2127 5814
rect 1946 5808 2127 5811
rect 1755 5788 1768 5790
rect 1783 5788 1817 5790
rect 1755 5772 1829 5788
rect 1856 5784 1869 5798
rect 1884 5784 1900 5800
rect 1946 5795 1957 5808
rect 1739 5750 1740 5766
rect 1755 5750 1768 5772
rect 1783 5750 1813 5772
rect 1856 5768 1918 5784
rect 1946 5777 1957 5793
rect 1962 5788 1972 5808
rect 1982 5788 1996 5808
rect 1999 5795 2008 5808
rect 2024 5795 2033 5808
rect 1962 5777 1996 5788
rect 1999 5777 2008 5793
rect 2024 5777 2033 5793
rect 2040 5788 2050 5808
rect 2060 5788 2074 5808
rect 2075 5795 2086 5808
rect 2040 5777 2074 5788
rect 2075 5777 2086 5793
rect 2132 5784 2148 5800
rect 2155 5798 2185 5850
rect 2219 5846 2220 5853
rect 2204 5838 2220 5846
rect 2191 5806 2204 5825
rect 2219 5806 2249 5822
rect 2191 5790 2265 5806
rect 2191 5788 2204 5790
rect 2219 5788 2253 5790
rect 1856 5766 1869 5768
rect 1884 5766 1918 5768
rect 1856 5750 1918 5766
rect 1962 5761 1978 5764
rect 2040 5761 2070 5772
rect 2118 5768 2164 5784
rect 2191 5772 2265 5788
rect 2118 5766 2152 5768
rect 2117 5750 2164 5766
rect 2191 5750 2204 5772
rect 2219 5750 2249 5772
rect 2276 5750 2277 5766
rect 2292 5750 2305 5910
rect 2335 5806 2348 5910
rect 2393 5888 2394 5898
rect 2409 5888 2422 5898
rect 2393 5884 2422 5888
rect 2427 5884 2457 5910
rect 2475 5896 2491 5898
rect 2563 5896 2616 5910
rect 2564 5894 2628 5896
rect 2671 5894 2686 5910
rect 2735 5907 2765 5910
rect 2735 5904 2771 5907
rect 2701 5896 2717 5898
rect 2475 5884 2490 5888
rect 2393 5882 2490 5884
rect 2518 5882 2686 5894
rect 2702 5884 2717 5888
rect 2735 5885 2774 5904
rect 2793 5898 2800 5899
rect 2799 5891 2800 5898
rect 2783 5888 2784 5891
rect 2799 5888 2812 5891
rect 2735 5884 2765 5885
rect 2774 5884 2780 5885
rect 2783 5884 2812 5888
rect 2702 5883 2812 5884
rect 2702 5882 2818 5883
rect 2377 5874 2428 5882
rect 2377 5862 2402 5874
rect 2409 5862 2428 5874
rect 2459 5874 2509 5882
rect 2459 5866 2475 5874
rect 2482 5872 2509 5874
rect 2518 5872 2739 5882
rect 2482 5862 2739 5872
rect 2768 5874 2818 5882
rect 2768 5865 2784 5874
rect 2377 5854 2428 5862
rect 2475 5854 2739 5862
rect 2765 5862 2784 5865
rect 2791 5862 2818 5874
rect 2765 5854 2818 5862
rect 2393 5846 2394 5854
rect 2409 5846 2422 5854
rect 2393 5838 2409 5846
rect 2390 5831 2409 5834
rect 2390 5822 2412 5831
rect 2363 5812 2412 5822
rect 2363 5806 2393 5812
rect 2412 5807 2417 5812
rect 2335 5790 2409 5806
rect 2427 5798 2457 5854
rect 2492 5844 2700 5854
rect 2735 5850 2780 5854
rect 2783 5853 2784 5854
rect 2799 5853 2812 5854
rect 2518 5814 2707 5844
rect 2533 5811 2707 5814
rect 2526 5808 2707 5811
rect 2335 5788 2348 5790
rect 2363 5788 2397 5790
rect 2335 5772 2409 5788
rect 2436 5784 2449 5798
rect 2464 5784 2480 5800
rect 2526 5795 2537 5808
rect 2319 5750 2320 5766
rect 2335 5750 2348 5772
rect 2363 5750 2393 5772
rect 2436 5768 2498 5784
rect 2526 5777 2537 5793
rect 2542 5788 2552 5808
rect 2562 5788 2576 5808
rect 2579 5795 2588 5808
rect 2604 5795 2613 5808
rect 2542 5777 2576 5788
rect 2579 5777 2588 5793
rect 2604 5777 2613 5793
rect 2620 5788 2630 5808
rect 2640 5788 2654 5808
rect 2655 5795 2666 5808
rect 2620 5777 2654 5788
rect 2655 5777 2666 5793
rect 2712 5784 2728 5800
rect 2735 5798 2765 5850
rect 2799 5846 2800 5853
rect 2784 5838 2800 5846
rect 2771 5806 2784 5825
rect 2799 5806 2829 5822
rect 2771 5790 2845 5806
rect 2771 5788 2784 5790
rect 2799 5788 2833 5790
rect 2436 5766 2449 5768
rect 2464 5766 2498 5768
rect 2436 5750 2498 5766
rect 2542 5761 2558 5764
rect 2620 5761 2650 5772
rect 2698 5768 2744 5784
rect 2771 5772 2845 5788
rect 2698 5766 2732 5768
rect 2697 5750 2744 5766
rect 2771 5750 2784 5772
rect 2799 5750 2829 5772
rect 2856 5750 2857 5766
rect 2872 5750 2885 5910
rect 2915 5806 2928 5910
rect 2973 5888 2974 5898
rect 2989 5888 3002 5898
rect 2973 5884 3002 5888
rect 3007 5884 3037 5910
rect 3055 5896 3071 5898
rect 3143 5896 3196 5910
rect 3144 5894 3208 5896
rect 3251 5894 3266 5910
rect 3315 5907 3345 5910
rect 3315 5904 3351 5907
rect 3281 5896 3297 5898
rect 3055 5884 3070 5888
rect 2973 5882 3070 5884
rect 3098 5882 3266 5894
rect 3282 5884 3297 5888
rect 3315 5885 3354 5904
rect 3373 5898 3380 5899
rect 3379 5891 3380 5898
rect 3363 5888 3364 5891
rect 3379 5888 3392 5891
rect 3315 5884 3345 5885
rect 3354 5884 3360 5885
rect 3363 5884 3392 5888
rect 3282 5883 3392 5884
rect 3282 5882 3398 5883
rect 2957 5874 3008 5882
rect 2957 5862 2982 5874
rect 2989 5862 3008 5874
rect 3039 5874 3089 5882
rect 3039 5866 3055 5874
rect 3062 5872 3089 5874
rect 3098 5872 3319 5882
rect 3062 5862 3319 5872
rect 3348 5874 3398 5882
rect 3348 5865 3364 5874
rect 2957 5854 3008 5862
rect 3055 5854 3319 5862
rect 3345 5862 3364 5865
rect 3371 5862 3398 5874
rect 3345 5854 3398 5862
rect 2973 5846 2974 5854
rect 2989 5846 3002 5854
rect 2973 5838 2989 5846
rect 2970 5831 2989 5834
rect 2970 5822 2992 5831
rect 2943 5812 2992 5822
rect 2943 5806 2973 5812
rect 2992 5807 2997 5812
rect 2915 5790 2989 5806
rect 3007 5798 3037 5854
rect 3072 5844 3280 5854
rect 3315 5850 3360 5854
rect 3363 5853 3364 5854
rect 3379 5853 3392 5854
rect 3098 5814 3287 5844
rect 3113 5811 3287 5814
rect 3106 5808 3287 5811
rect 2915 5788 2928 5790
rect 2943 5788 2977 5790
rect 2915 5772 2989 5788
rect 3016 5784 3029 5798
rect 3044 5784 3060 5800
rect 3106 5795 3117 5808
rect 2899 5750 2900 5766
rect 2915 5750 2928 5772
rect 2943 5750 2973 5772
rect 3016 5768 3078 5784
rect 3106 5777 3117 5793
rect 3122 5788 3132 5808
rect 3142 5788 3156 5808
rect 3159 5795 3168 5808
rect 3184 5795 3193 5808
rect 3122 5777 3156 5788
rect 3159 5777 3168 5793
rect 3184 5777 3193 5793
rect 3200 5788 3210 5808
rect 3220 5788 3234 5808
rect 3235 5795 3246 5808
rect 3200 5777 3234 5788
rect 3235 5777 3246 5793
rect 3292 5784 3308 5800
rect 3315 5798 3345 5850
rect 3379 5846 3380 5853
rect 3364 5838 3380 5846
rect 3351 5806 3364 5825
rect 3379 5806 3409 5822
rect 3351 5790 3425 5806
rect 3351 5788 3364 5790
rect 3379 5788 3413 5790
rect 3016 5766 3029 5768
rect 3044 5766 3078 5768
rect 3016 5750 3078 5766
rect 3122 5761 3138 5764
rect 3200 5761 3230 5772
rect 3278 5768 3324 5784
rect 3351 5772 3425 5788
rect 3278 5766 3312 5768
rect 3277 5750 3324 5766
rect 3351 5750 3364 5772
rect 3379 5750 3409 5772
rect 3436 5750 3437 5766
rect 3452 5750 3465 5910
rect 3495 5806 3508 5910
rect 3553 5888 3554 5898
rect 3569 5888 3582 5898
rect 3553 5884 3582 5888
rect 3587 5884 3617 5910
rect 3635 5896 3651 5898
rect 3723 5896 3776 5910
rect 3724 5894 3788 5896
rect 3831 5894 3846 5910
rect 3895 5907 3925 5910
rect 3895 5904 3931 5907
rect 3861 5896 3877 5898
rect 3635 5884 3650 5888
rect 3553 5882 3650 5884
rect 3678 5882 3846 5894
rect 3862 5884 3877 5888
rect 3895 5885 3934 5904
rect 3953 5898 3960 5899
rect 3959 5891 3960 5898
rect 3943 5888 3944 5891
rect 3959 5888 3972 5891
rect 3895 5884 3925 5885
rect 3934 5884 3940 5885
rect 3943 5884 3972 5888
rect 3862 5883 3972 5884
rect 3862 5882 3978 5883
rect 3537 5874 3588 5882
rect 3537 5862 3562 5874
rect 3569 5862 3588 5874
rect 3619 5874 3669 5882
rect 3619 5866 3635 5874
rect 3642 5872 3669 5874
rect 3678 5872 3899 5882
rect 3642 5862 3899 5872
rect 3928 5874 3978 5882
rect 3928 5865 3944 5874
rect 3537 5854 3588 5862
rect 3635 5854 3899 5862
rect 3925 5862 3944 5865
rect 3951 5862 3978 5874
rect 3925 5854 3978 5862
rect 3553 5846 3554 5854
rect 3569 5846 3582 5854
rect 3553 5838 3569 5846
rect 3550 5831 3569 5834
rect 3550 5822 3572 5831
rect 3523 5812 3572 5822
rect 3523 5806 3553 5812
rect 3572 5807 3577 5812
rect 3495 5790 3569 5806
rect 3587 5798 3617 5854
rect 3652 5844 3860 5854
rect 3895 5850 3940 5854
rect 3943 5853 3944 5854
rect 3959 5853 3972 5854
rect 3678 5814 3867 5844
rect 3693 5811 3867 5814
rect 3686 5808 3867 5811
rect 3495 5788 3508 5790
rect 3523 5788 3557 5790
rect 3495 5772 3569 5788
rect 3596 5784 3609 5798
rect 3624 5784 3640 5800
rect 3686 5795 3697 5808
rect 3479 5750 3480 5766
rect 3495 5750 3508 5772
rect 3523 5750 3553 5772
rect 3596 5768 3658 5784
rect 3686 5777 3697 5793
rect 3702 5788 3712 5808
rect 3722 5788 3736 5808
rect 3739 5795 3748 5808
rect 3764 5795 3773 5808
rect 3702 5777 3736 5788
rect 3739 5777 3748 5793
rect 3764 5777 3773 5793
rect 3780 5788 3790 5808
rect 3800 5788 3814 5808
rect 3815 5795 3826 5808
rect 3780 5777 3814 5788
rect 3815 5777 3826 5793
rect 3872 5784 3888 5800
rect 3895 5798 3925 5850
rect 3959 5846 3960 5853
rect 3944 5838 3960 5846
rect 3931 5806 3944 5825
rect 3959 5806 3989 5822
rect 3931 5790 4005 5806
rect 3931 5788 3944 5790
rect 3959 5788 3993 5790
rect 3596 5766 3609 5768
rect 3624 5766 3658 5768
rect 3596 5750 3658 5766
rect 3702 5761 3718 5764
rect 3780 5761 3810 5772
rect 3858 5768 3904 5784
rect 3931 5772 4005 5788
rect 3858 5766 3892 5768
rect 3857 5750 3904 5766
rect 3931 5750 3944 5772
rect 3959 5750 3989 5772
rect 4016 5750 4017 5766
rect 4032 5750 4045 5910
rect 4075 5806 4088 5910
rect 4133 5888 4134 5898
rect 4149 5888 4162 5898
rect 4133 5884 4162 5888
rect 4167 5884 4197 5910
rect 4215 5896 4231 5898
rect 4303 5896 4356 5910
rect 4304 5894 4368 5896
rect 4411 5894 4426 5910
rect 4475 5907 4505 5910
rect 4475 5904 4511 5907
rect 4441 5896 4457 5898
rect 4215 5884 4230 5888
rect 4133 5882 4230 5884
rect 4258 5882 4426 5894
rect 4442 5884 4457 5888
rect 4475 5885 4514 5904
rect 4533 5898 4540 5899
rect 4539 5891 4540 5898
rect 4523 5888 4524 5891
rect 4539 5888 4552 5891
rect 4475 5884 4505 5885
rect 4514 5884 4520 5885
rect 4523 5884 4552 5888
rect 4442 5883 4552 5884
rect 4442 5882 4558 5883
rect 4117 5874 4168 5882
rect 4117 5862 4142 5874
rect 4149 5862 4168 5874
rect 4199 5874 4249 5882
rect 4199 5866 4215 5874
rect 4222 5872 4249 5874
rect 4258 5872 4479 5882
rect 4222 5862 4479 5872
rect 4508 5874 4558 5882
rect 4508 5865 4524 5874
rect 4117 5854 4168 5862
rect 4215 5854 4479 5862
rect 4505 5862 4524 5865
rect 4531 5862 4558 5874
rect 4505 5854 4558 5862
rect 4133 5846 4134 5854
rect 4149 5846 4162 5854
rect 4133 5838 4149 5846
rect 4130 5831 4149 5834
rect 4130 5822 4152 5831
rect 4103 5812 4152 5822
rect 4103 5806 4133 5812
rect 4152 5807 4157 5812
rect 4075 5790 4149 5806
rect 4167 5798 4197 5854
rect 4232 5844 4440 5854
rect 4475 5850 4520 5854
rect 4523 5853 4524 5854
rect 4539 5853 4552 5854
rect 4258 5814 4447 5844
rect 4273 5811 4447 5814
rect 4266 5808 4447 5811
rect 4075 5788 4088 5790
rect 4103 5788 4137 5790
rect 4075 5772 4149 5788
rect 4176 5784 4189 5798
rect 4204 5784 4220 5800
rect 4266 5795 4277 5808
rect 4059 5750 4060 5766
rect 4075 5750 4088 5772
rect 4103 5750 4133 5772
rect 4176 5768 4238 5784
rect 4266 5777 4277 5793
rect 4282 5788 4292 5808
rect 4302 5788 4316 5808
rect 4319 5795 4328 5808
rect 4344 5795 4353 5808
rect 4282 5777 4316 5788
rect 4319 5777 4328 5793
rect 4344 5777 4353 5793
rect 4360 5788 4370 5808
rect 4380 5788 4394 5808
rect 4395 5795 4406 5808
rect 4360 5777 4394 5788
rect 4395 5777 4406 5793
rect 4452 5784 4468 5800
rect 4475 5798 4505 5850
rect 4539 5846 4540 5853
rect 4524 5838 4540 5846
rect 4511 5806 4524 5825
rect 4539 5806 4569 5822
rect 4511 5790 4585 5806
rect 4511 5788 4524 5790
rect 4539 5788 4573 5790
rect 4176 5766 4189 5768
rect 4204 5766 4238 5768
rect 4176 5750 4238 5766
rect 4282 5761 4298 5764
rect 4360 5761 4390 5772
rect 4438 5768 4484 5784
rect 4511 5772 4585 5788
rect 4438 5766 4472 5768
rect 4437 5750 4484 5766
rect 4511 5750 4524 5772
rect 4539 5750 4569 5772
rect 4596 5750 4597 5766
rect 4612 5750 4625 5910
rect -7 5742 34 5750
rect -7 5716 8 5742
rect 15 5716 34 5742
rect 98 5738 160 5750
rect 172 5738 247 5750
rect 305 5738 380 5750
rect 392 5738 423 5750
rect 429 5738 464 5750
rect 98 5736 260 5738
rect -7 5708 34 5716
rect 116 5712 129 5736
rect 144 5734 159 5736
rect -1 5698 0 5708
rect 15 5698 28 5708
rect 43 5698 73 5712
rect 116 5698 159 5712
rect 183 5709 190 5716
rect 193 5712 260 5736
rect 292 5736 464 5738
rect 262 5714 290 5718
rect 292 5714 372 5736
rect 393 5734 408 5736
rect 262 5712 372 5714
rect 193 5708 372 5712
rect 166 5698 196 5708
rect 198 5698 351 5708
rect 359 5698 389 5708
rect 393 5698 423 5712
rect 451 5698 464 5736
rect 536 5742 571 5750
rect 536 5716 537 5742
rect 544 5716 571 5742
rect 479 5698 509 5712
rect 536 5708 571 5716
rect 573 5742 614 5750
rect 573 5716 588 5742
rect 595 5716 614 5742
rect 678 5738 740 5750
rect 752 5738 827 5750
rect 885 5738 960 5750
rect 972 5738 1003 5750
rect 1009 5738 1044 5750
rect 678 5736 840 5738
rect 573 5708 614 5716
rect 696 5712 709 5736
rect 724 5734 739 5736
rect 536 5698 537 5708
rect 552 5698 565 5708
rect 579 5698 580 5708
rect 595 5698 608 5708
rect 623 5698 653 5712
rect 696 5698 739 5712
rect 763 5709 770 5716
rect 773 5712 840 5736
rect 872 5736 1044 5738
rect 842 5714 870 5718
rect 872 5714 952 5736
rect 973 5734 988 5736
rect 842 5712 952 5714
rect 773 5708 952 5712
rect 746 5698 776 5708
rect 778 5698 931 5708
rect 939 5698 969 5708
rect 973 5698 1003 5712
rect 1031 5698 1044 5736
rect 1116 5742 1151 5750
rect 1116 5716 1117 5742
rect 1124 5716 1151 5742
rect 1059 5698 1089 5712
rect 1116 5708 1151 5716
rect 1153 5742 1194 5750
rect 1153 5716 1168 5742
rect 1175 5716 1194 5742
rect 1258 5738 1320 5750
rect 1332 5738 1407 5750
rect 1465 5738 1540 5750
rect 1552 5738 1583 5750
rect 1589 5738 1624 5750
rect 1258 5736 1420 5738
rect 1153 5708 1194 5716
rect 1276 5712 1289 5736
rect 1304 5734 1319 5736
rect 1116 5698 1117 5708
rect 1132 5698 1145 5708
rect 1159 5698 1160 5708
rect 1175 5698 1188 5708
rect 1203 5698 1233 5712
rect 1276 5698 1319 5712
rect 1343 5709 1350 5716
rect 1353 5712 1420 5736
rect 1452 5736 1624 5738
rect 1422 5714 1450 5718
rect 1452 5714 1532 5736
rect 1553 5734 1568 5736
rect 1422 5712 1532 5714
rect 1353 5708 1532 5712
rect 1326 5698 1356 5708
rect 1358 5698 1511 5708
rect 1519 5698 1549 5708
rect 1553 5698 1583 5712
rect 1611 5698 1624 5736
rect 1696 5742 1731 5750
rect 1696 5716 1697 5742
rect 1704 5716 1731 5742
rect 1639 5698 1669 5712
rect 1696 5708 1731 5716
rect 1733 5742 1774 5750
rect 1733 5716 1748 5742
rect 1755 5716 1774 5742
rect 1838 5738 1900 5750
rect 1912 5738 1987 5750
rect 2045 5738 2120 5750
rect 2132 5738 2163 5750
rect 2169 5738 2204 5750
rect 1838 5736 2000 5738
rect 1733 5708 1774 5716
rect 1856 5712 1869 5736
rect 1884 5734 1899 5736
rect 1696 5698 1697 5708
rect 1712 5698 1725 5708
rect 1739 5698 1740 5708
rect 1755 5698 1768 5708
rect 1783 5698 1813 5712
rect 1856 5698 1899 5712
rect 1923 5709 1930 5716
rect 1933 5712 2000 5736
rect 2032 5736 2204 5738
rect 2002 5714 2030 5718
rect 2032 5714 2112 5736
rect 2133 5734 2148 5736
rect 2002 5712 2112 5714
rect 1933 5708 2112 5712
rect 1906 5698 1936 5708
rect 1938 5698 2091 5708
rect 2099 5698 2129 5708
rect 2133 5698 2163 5712
rect 2191 5698 2204 5736
rect 2276 5742 2311 5750
rect 2276 5716 2277 5742
rect 2284 5716 2311 5742
rect 2219 5698 2249 5712
rect 2276 5708 2311 5716
rect 2313 5742 2354 5750
rect 2313 5716 2328 5742
rect 2335 5716 2354 5742
rect 2418 5738 2480 5750
rect 2492 5738 2567 5750
rect 2625 5738 2700 5750
rect 2712 5738 2743 5750
rect 2749 5738 2784 5750
rect 2418 5736 2580 5738
rect 2313 5708 2354 5716
rect 2436 5712 2449 5736
rect 2464 5734 2479 5736
rect 2276 5698 2277 5708
rect 2292 5698 2305 5708
rect 2319 5698 2320 5708
rect 2335 5698 2348 5708
rect 2363 5698 2393 5712
rect 2436 5698 2479 5712
rect 2503 5709 2510 5716
rect 2513 5712 2580 5736
rect 2612 5736 2784 5738
rect 2582 5714 2610 5718
rect 2612 5714 2692 5736
rect 2713 5734 2728 5736
rect 2582 5712 2692 5714
rect 2513 5708 2692 5712
rect 2486 5698 2516 5708
rect 2518 5698 2671 5708
rect 2679 5698 2709 5708
rect 2713 5698 2743 5712
rect 2771 5698 2784 5736
rect 2856 5742 2891 5750
rect 2856 5716 2857 5742
rect 2864 5716 2891 5742
rect 2799 5698 2829 5712
rect 2856 5708 2891 5716
rect 2893 5742 2934 5750
rect 2893 5716 2908 5742
rect 2915 5716 2934 5742
rect 2998 5738 3060 5750
rect 3072 5738 3147 5750
rect 3205 5738 3280 5750
rect 3292 5738 3323 5750
rect 3329 5738 3364 5750
rect 2998 5736 3160 5738
rect 2893 5708 2934 5716
rect 3016 5712 3029 5736
rect 3044 5734 3059 5736
rect 2856 5698 2857 5708
rect 2872 5698 2885 5708
rect 2899 5698 2900 5708
rect 2915 5698 2928 5708
rect 2943 5698 2973 5712
rect 3016 5698 3059 5712
rect 3083 5709 3090 5716
rect 3093 5712 3160 5736
rect 3192 5736 3364 5738
rect 3162 5714 3190 5718
rect 3192 5714 3272 5736
rect 3293 5734 3308 5736
rect 3162 5712 3272 5714
rect 3093 5708 3272 5712
rect 3066 5698 3096 5708
rect 3098 5698 3251 5708
rect 3259 5698 3289 5708
rect 3293 5698 3323 5712
rect 3351 5698 3364 5736
rect 3436 5742 3471 5750
rect 3436 5716 3437 5742
rect 3444 5716 3471 5742
rect 3379 5698 3409 5712
rect 3436 5708 3471 5716
rect 3473 5742 3514 5750
rect 3473 5716 3488 5742
rect 3495 5716 3514 5742
rect 3578 5738 3640 5750
rect 3652 5738 3727 5750
rect 3785 5738 3860 5750
rect 3872 5738 3903 5750
rect 3909 5738 3944 5750
rect 3578 5736 3740 5738
rect 3473 5708 3514 5716
rect 3596 5712 3609 5736
rect 3624 5734 3639 5736
rect 3436 5698 3437 5708
rect 3452 5698 3465 5708
rect 3479 5698 3480 5708
rect 3495 5698 3508 5708
rect 3523 5698 3553 5712
rect 3596 5698 3639 5712
rect 3663 5709 3670 5716
rect 3673 5712 3740 5736
rect 3772 5736 3944 5738
rect 3742 5714 3770 5718
rect 3772 5714 3852 5736
rect 3873 5734 3888 5736
rect 3742 5712 3852 5714
rect 3673 5708 3852 5712
rect 3646 5698 3676 5708
rect 3678 5698 3831 5708
rect 3839 5698 3869 5708
rect 3873 5698 3903 5712
rect 3931 5698 3944 5736
rect 4016 5742 4051 5750
rect 4016 5716 4017 5742
rect 4024 5716 4051 5742
rect 3959 5698 3989 5712
rect 4016 5708 4051 5716
rect 4053 5742 4094 5750
rect 4053 5716 4068 5742
rect 4075 5716 4094 5742
rect 4158 5738 4220 5750
rect 4232 5738 4307 5750
rect 4365 5738 4440 5750
rect 4452 5738 4483 5750
rect 4489 5738 4524 5750
rect 4158 5736 4320 5738
rect 4053 5708 4094 5716
rect 4176 5712 4189 5736
rect 4204 5734 4219 5736
rect 4016 5698 4017 5708
rect 4032 5698 4045 5708
rect 4059 5698 4060 5708
rect 4075 5698 4088 5708
rect 4103 5698 4133 5712
rect 4176 5698 4219 5712
rect 4243 5709 4250 5716
rect 4253 5712 4320 5736
rect 4352 5736 4524 5738
rect 4322 5714 4350 5718
rect 4352 5714 4432 5736
rect 4453 5734 4468 5736
rect 4322 5712 4432 5714
rect 4253 5708 4432 5712
rect 4226 5698 4256 5708
rect 4258 5698 4411 5708
rect 4419 5698 4449 5708
rect 4453 5698 4483 5712
rect 4511 5698 4524 5736
rect 4596 5742 4631 5750
rect 4596 5716 4597 5742
rect 4604 5716 4631 5742
rect 4539 5698 4569 5712
rect 4596 5708 4631 5716
rect 4596 5698 4597 5708
rect 4612 5698 4625 5708
rect -1 5692 4625 5698
rect 0 5684 4625 5692
rect 15 5654 28 5684
rect 43 5666 73 5684
rect 116 5670 130 5684
rect 166 5670 386 5684
rect 117 5668 130 5670
rect 83 5656 98 5668
rect 80 5654 102 5656
rect 107 5654 137 5668
rect 198 5666 351 5670
rect 180 5654 372 5666
rect 415 5654 445 5668
rect 451 5654 464 5684
rect 479 5666 509 5684
rect 552 5654 565 5684
rect 595 5654 608 5684
rect 623 5666 653 5684
rect 696 5670 710 5684
rect 746 5670 966 5684
rect 697 5668 710 5670
rect 663 5656 678 5668
rect 660 5654 682 5656
rect 687 5654 717 5668
rect 778 5666 931 5670
rect 760 5654 952 5666
rect 995 5654 1025 5668
rect 1031 5654 1044 5684
rect 1059 5666 1089 5684
rect 1132 5654 1145 5684
rect 1175 5654 1188 5684
rect 1203 5666 1233 5684
rect 1276 5670 1290 5684
rect 1326 5670 1546 5684
rect 1277 5668 1290 5670
rect 1243 5656 1258 5668
rect 1240 5654 1262 5656
rect 1267 5654 1297 5668
rect 1358 5666 1511 5670
rect 1340 5654 1532 5666
rect 1575 5654 1605 5668
rect 1611 5654 1624 5684
rect 1639 5666 1669 5684
rect 1712 5654 1725 5684
rect 1755 5654 1768 5684
rect 1783 5666 1813 5684
rect 1856 5670 1870 5684
rect 1906 5670 2126 5684
rect 1857 5668 1870 5670
rect 1823 5656 1838 5668
rect 1820 5654 1842 5656
rect 1847 5654 1877 5668
rect 1938 5666 2091 5670
rect 1920 5654 2112 5666
rect 2155 5654 2185 5668
rect 2191 5654 2204 5684
rect 2219 5666 2249 5684
rect 2292 5654 2305 5684
rect 2335 5654 2348 5684
rect 2363 5666 2393 5684
rect 2436 5670 2450 5684
rect 2486 5670 2706 5684
rect 2437 5668 2450 5670
rect 2403 5656 2418 5668
rect 2400 5654 2422 5656
rect 2427 5654 2457 5668
rect 2518 5666 2671 5670
rect 2500 5654 2692 5666
rect 2735 5654 2765 5668
rect 2771 5654 2784 5684
rect 2799 5666 2829 5684
rect 2872 5654 2885 5684
rect 2915 5654 2928 5684
rect 2943 5666 2973 5684
rect 3016 5670 3030 5684
rect 3066 5670 3286 5684
rect 3017 5668 3030 5670
rect 2983 5656 2998 5668
rect 2980 5654 3002 5656
rect 3007 5654 3037 5668
rect 3098 5666 3251 5670
rect 3080 5654 3272 5666
rect 3315 5654 3345 5668
rect 3351 5654 3364 5684
rect 3379 5666 3409 5684
rect 3452 5654 3465 5684
rect 3495 5654 3508 5684
rect 3523 5666 3553 5684
rect 3596 5670 3610 5684
rect 3646 5670 3866 5684
rect 3597 5668 3610 5670
rect 3563 5656 3578 5668
rect 3560 5654 3582 5656
rect 3587 5654 3617 5668
rect 3678 5666 3831 5670
rect 3660 5654 3852 5666
rect 3895 5654 3925 5668
rect 3931 5654 3944 5684
rect 3959 5666 3989 5684
rect 4032 5654 4045 5684
rect 4075 5654 4088 5684
rect 4103 5666 4133 5684
rect 4176 5670 4190 5684
rect 4226 5670 4446 5684
rect 4177 5668 4190 5670
rect 4143 5656 4158 5668
rect 4140 5654 4162 5656
rect 4167 5654 4197 5668
rect 4258 5666 4411 5670
rect 4240 5654 4432 5666
rect 4475 5654 4505 5668
rect 4511 5654 4524 5684
rect 4539 5666 4569 5684
rect 4612 5654 4625 5684
rect 0 5640 4625 5654
rect 15 5536 28 5640
rect 73 5618 74 5628
rect 89 5618 102 5628
rect 73 5614 102 5618
rect 107 5614 137 5640
rect 155 5626 171 5628
rect 243 5626 296 5640
rect 244 5624 308 5626
rect 351 5624 366 5640
rect 415 5637 445 5640
rect 415 5634 451 5637
rect 381 5626 397 5628
rect 155 5614 170 5618
rect 73 5612 170 5614
rect 198 5612 366 5624
rect 382 5614 397 5618
rect 415 5615 454 5634
rect 473 5628 480 5629
rect 479 5621 480 5628
rect 463 5618 464 5621
rect 479 5618 492 5621
rect 415 5614 445 5615
rect 454 5614 460 5615
rect 463 5614 492 5618
rect 382 5613 492 5614
rect 382 5612 498 5613
rect 57 5604 108 5612
rect 57 5592 82 5604
rect 89 5592 108 5604
rect 139 5604 189 5612
rect 139 5596 155 5604
rect 162 5602 189 5604
rect 198 5602 419 5612
rect 162 5592 419 5602
rect 448 5604 498 5612
rect 448 5595 464 5604
rect 57 5584 108 5592
rect 155 5584 419 5592
rect 445 5592 464 5595
rect 471 5592 498 5604
rect 445 5584 498 5592
rect 73 5576 74 5584
rect 89 5576 102 5584
rect 73 5568 89 5576
rect 70 5561 89 5564
rect 70 5552 92 5561
rect 43 5542 92 5552
rect 43 5536 73 5542
rect 92 5537 97 5542
rect 15 5520 89 5536
rect 107 5528 137 5584
rect 172 5574 380 5584
rect 415 5580 460 5584
rect 463 5583 464 5584
rect 479 5583 492 5584
rect 198 5544 387 5574
rect 213 5541 387 5544
rect 206 5538 387 5541
rect 15 5518 28 5520
rect 43 5518 77 5520
rect 15 5502 89 5518
rect 116 5514 129 5528
rect 144 5514 160 5530
rect 206 5525 217 5538
rect -1 5480 0 5496
rect 15 5480 28 5502
rect 43 5480 73 5502
rect 116 5498 178 5514
rect 206 5507 217 5523
rect 222 5518 232 5538
rect 242 5518 256 5538
rect 259 5525 268 5538
rect 284 5525 293 5538
rect 222 5507 256 5518
rect 259 5507 268 5523
rect 284 5507 293 5523
rect 300 5518 310 5538
rect 320 5518 334 5538
rect 335 5525 346 5538
rect 300 5507 334 5518
rect 335 5507 346 5523
rect 392 5514 408 5530
rect 415 5528 445 5580
rect 479 5576 480 5583
rect 464 5568 480 5576
rect 451 5536 464 5555
rect 479 5536 509 5552
rect 451 5520 525 5536
rect 451 5518 464 5520
rect 479 5518 513 5520
rect 116 5496 129 5498
rect 144 5496 178 5498
rect 116 5480 178 5496
rect 222 5491 238 5494
rect 300 5491 330 5502
rect 378 5498 424 5514
rect 451 5502 525 5518
rect 378 5496 412 5498
rect 377 5480 424 5496
rect 451 5480 464 5502
rect 479 5480 509 5502
rect 536 5480 537 5496
rect 552 5480 565 5640
rect 595 5536 608 5640
rect 653 5618 654 5628
rect 669 5618 682 5628
rect 653 5614 682 5618
rect 687 5614 717 5640
rect 735 5626 751 5628
rect 823 5626 876 5640
rect 824 5624 888 5626
rect 931 5624 946 5640
rect 995 5637 1025 5640
rect 995 5634 1031 5637
rect 961 5626 977 5628
rect 735 5614 750 5618
rect 653 5612 750 5614
rect 778 5612 946 5624
rect 962 5614 977 5618
rect 995 5615 1034 5634
rect 1053 5628 1060 5629
rect 1059 5621 1060 5628
rect 1043 5618 1044 5621
rect 1059 5618 1072 5621
rect 995 5614 1025 5615
rect 1034 5614 1040 5615
rect 1043 5614 1072 5618
rect 962 5613 1072 5614
rect 962 5612 1078 5613
rect 637 5604 688 5612
rect 637 5592 662 5604
rect 669 5592 688 5604
rect 719 5604 769 5612
rect 719 5596 735 5604
rect 742 5602 769 5604
rect 778 5602 999 5612
rect 742 5592 999 5602
rect 1028 5604 1078 5612
rect 1028 5595 1044 5604
rect 637 5584 688 5592
rect 735 5584 999 5592
rect 1025 5592 1044 5595
rect 1051 5592 1078 5604
rect 1025 5584 1078 5592
rect 653 5576 654 5584
rect 669 5576 682 5584
rect 653 5568 669 5576
rect 650 5561 669 5564
rect 650 5552 672 5561
rect 623 5542 672 5552
rect 623 5536 653 5542
rect 672 5537 677 5542
rect 595 5520 669 5536
rect 687 5528 717 5584
rect 752 5574 960 5584
rect 995 5580 1040 5584
rect 1043 5583 1044 5584
rect 1059 5583 1072 5584
rect 778 5544 967 5574
rect 793 5541 967 5544
rect 786 5538 967 5541
rect 595 5518 608 5520
rect 623 5518 657 5520
rect 595 5502 669 5518
rect 696 5514 709 5528
rect 724 5514 740 5530
rect 786 5525 797 5538
rect 579 5480 580 5496
rect 595 5480 608 5502
rect 623 5480 653 5502
rect 696 5498 758 5514
rect 786 5507 797 5523
rect 802 5518 812 5538
rect 822 5518 836 5538
rect 839 5525 848 5538
rect 864 5525 873 5538
rect 802 5507 836 5518
rect 839 5507 848 5523
rect 864 5507 873 5523
rect 880 5518 890 5538
rect 900 5518 914 5538
rect 915 5525 926 5538
rect 880 5507 914 5518
rect 915 5507 926 5523
rect 972 5514 988 5530
rect 995 5528 1025 5580
rect 1059 5576 1060 5583
rect 1044 5568 1060 5576
rect 1031 5536 1044 5555
rect 1059 5536 1089 5552
rect 1031 5520 1105 5536
rect 1031 5518 1044 5520
rect 1059 5518 1093 5520
rect 696 5496 709 5498
rect 724 5496 758 5498
rect 696 5480 758 5496
rect 802 5491 818 5494
rect 880 5491 910 5502
rect 958 5498 1004 5514
rect 1031 5502 1105 5518
rect 958 5496 992 5498
rect 957 5480 1004 5496
rect 1031 5480 1044 5502
rect 1059 5480 1089 5502
rect 1116 5480 1117 5496
rect 1132 5480 1145 5640
rect 1175 5536 1188 5640
rect 1233 5618 1234 5628
rect 1249 5618 1262 5628
rect 1233 5614 1262 5618
rect 1267 5614 1297 5640
rect 1315 5626 1331 5628
rect 1403 5626 1456 5640
rect 1404 5624 1468 5626
rect 1511 5624 1526 5640
rect 1575 5637 1605 5640
rect 1575 5634 1611 5637
rect 1541 5626 1557 5628
rect 1315 5614 1330 5618
rect 1233 5612 1330 5614
rect 1358 5612 1526 5624
rect 1542 5614 1557 5618
rect 1575 5615 1614 5634
rect 1633 5628 1640 5629
rect 1639 5621 1640 5628
rect 1623 5618 1624 5621
rect 1639 5618 1652 5621
rect 1575 5614 1605 5615
rect 1614 5614 1620 5615
rect 1623 5614 1652 5618
rect 1542 5613 1652 5614
rect 1542 5612 1658 5613
rect 1217 5604 1268 5612
rect 1217 5592 1242 5604
rect 1249 5592 1268 5604
rect 1299 5604 1349 5612
rect 1299 5596 1315 5604
rect 1322 5602 1349 5604
rect 1358 5602 1579 5612
rect 1322 5592 1579 5602
rect 1608 5604 1658 5612
rect 1608 5595 1624 5604
rect 1217 5584 1268 5592
rect 1315 5584 1579 5592
rect 1605 5592 1624 5595
rect 1631 5592 1658 5604
rect 1605 5584 1658 5592
rect 1233 5576 1234 5584
rect 1249 5576 1262 5584
rect 1233 5568 1249 5576
rect 1230 5561 1249 5564
rect 1230 5552 1252 5561
rect 1203 5542 1252 5552
rect 1203 5536 1233 5542
rect 1252 5537 1257 5542
rect 1175 5520 1249 5536
rect 1267 5528 1297 5584
rect 1332 5574 1540 5584
rect 1575 5580 1620 5584
rect 1623 5583 1624 5584
rect 1639 5583 1652 5584
rect 1358 5544 1547 5574
rect 1373 5541 1547 5544
rect 1366 5538 1547 5541
rect 1175 5518 1188 5520
rect 1203 5518 1237 5520
rect 1175 5502 1249 5518
rect 1276 5514 1289 5528
rect 1304 5514 1320 5530
rect 1366 5525 1377 5538
rect 1159 5480 1160 5496
rect 1175 5480 1188 5502
rect 1203 5480 1233 5502
rect 1276 5498 1338 5514
rect 1366 5507 1377 5523
rect 1382 5518 1392 5538
rect 1402 5518 1416 5538
rect 1419 5525 1428 5538
rect 1444 5525 1453 5538
rect 1382 5507 1416 5518
rect 1419 5507 1428 5523
rect 1444 5507 1453 5523
rect 1460 5518 1470 5538
rect 1480 5518 1494 5538
rect 1495 5525 1506 5538
rect 1460 5507 1494 5518
rect 1495 5507 1506 5523
rect 1552 5514 1568 5530
rect 1575 5528 1605 5580
rect 1639 5576 1640 5583
rect 1624 5568 1640 5576
rect 1611 5536 1624 5555
rect 1639 5536 1669 5552
rect 1611 5520 1685 5536
rect 1611 5518 1624 5520
rect 1639 5518 1673 5520
rect 1276 5496 1289 5498
rect 1304 5496 1338 5498
rect 1276 5480 1338 5496
rect 1382 5491 1398 5494
rect 1460 5491 1490 5502
rect 1538 5498 1584 5514
rect 1611 5502 1685 5518
rect 1538 5496 1572 5498
rect 1537 5480 1584 5496
rect 1611 5480 1624 5502
rect 1639 5480 1669 5502
rect 1696 5480 1697 5496
rect 1712 5480 1725 5640
rect 1755 5536 1768 5640
rect 1813 5618 1814 5628
rect 1829 5618 1842 5628
rect 1813 5614 1842 5618
rect 1847 5614 1877 5640
rect 1895 5626 1911 5628
rect 1983 5626 2036 5640
rect 1984 5624 2048 5626
rect 2091 5624 2106 5640
rect 2155 5637 2185 5640
rect 2155 5634 2191 5637
rect 2121 5626 2137 5628
rect 1895 5614 1910 5618
rect 1813 5612 1910 5614
rect 1938 5612 2106 5624
rect 2122 5614 2137 5618
rect 2155 5615 2194 5634
rect 2213 5628 2220 5629
rect 2219 5621 2220 5628
rect 2203 5618 2204 5621
rect 2219 5618 2232 5621
rect 2155 5614 2185 5615
rect 2194 5614 2200 5615
rect 2203 5614 2232 5618
rect 2122 5613 2232 5614
rect 2122 5612 2238 5613
rect 1797 5604 1848 5612
rect 1797 5592 1822 5604
rect 1829 5592 1848 5604
rect 1879 5604 1929 5612
rect 1879 5596 1895 5604
rect 1902 5602 1929 5604
rect 1938 5602 2159 5612
rect 1902 5592 2159 5602
rect 2188 5604 2238 5612
rect 2188 5595 2204 5604
rect 1797 5584 1848 5592
rect 1895 5584 2159 5592
rect 2185 5592 2204 5595
rect 2211 5592 2238 5604
rect 2185 5584 2238 5592
rect 1813 5576 1814 5584
rect 1829 5576 1842 5584
rect 1813 5568 1829 5576
rect 1810 5561 1829 5564
rect 1810 5552 1832 5561
rect 1783 5542 1832 5552
rect 1783 5536 1813 5542
rect 1832 5537 1837 5542
rect 1755 5520 1829 5536
rect 1847 5528 1877 5584
rect 1912 5574 2120 5584
rect 2155 5580 2200 5584
rect 2203 5583 2204 5584
rect 2219 5583 2232 5584
rect 1938 5544 2127 5574
rect 1953 5541 2127 5544
rect 1946 5538 2127 5541
rect 1755 5518 1768 5520
rect 1783 5518 1817 5520
rect 1755 5502 1829 5518
rect 1856 5514 1869 5528
rect 1884 5514 1900 5530
rect 1946 5525 1957 5538
rect 1739 5480 1740 5496
rect 1755 5480 1768 5502
rect 1783 5480 1813 5502
rect 1856 5498 1918 5514
rect 1946 5507 1957 5523
rect 1962 5518 1972 5538
rect 1982 5518 1996 5538
rect 1999 5525 2008 5538
rect 2024 5525 2033 5538
rect 1962 5507 1996 5518
rect 1999 5507 2008 5523
rect 2024 5507 2033 5523
rect 2040 5518 2050 5538
rect 2060 5518 2074 5538
rect 2075 5525 2086 5538
rect 2040 5507 2074 5518
rect 2075 5507 2086 5523
rect 2132 5514 2148 5530
rect 2155 5528 2185 5580
rect 2219 5576 2220 5583
rect 2204 5568 2220 5576
rect 2191 5536 2204 5555
rect 2219 5536 2249 5552
rect 2191 5520 2265 5536
rect 2191 5518 2204 5520
rect 2219 5518 2253 5520
rect 1856 5496 1869 5498
rect 1884 5496 1918 5498
rect 1856 5480 1918 5496
rect 1962 5491 1978 5494
rect 2040 5491 2070 5502
rect 2118 5498 2164 5514
rect 2191 5502 2265 5518
rect 2118 5496 2152 5498
rect 2117 5480 2164 5496
rect 2191 5480 2204 5502
rect 2219 5480 2249 5502
rect 2276 5480 2277 5496
rect 2292 5480 2305 5640
rect 2335 5536 2348 5640
rect 2393 5618 2394 5628
rect 2409 5618 2422 5628
rect 2393 5614 2422 5618
rect 2427 5614 2457 5640
rect 2475 5626 2491 5628
rect 2563 5626 2616 5640
rect 2564 5624 2628 5626
rect 2671 5624 2686 5640
rect 2735 5637 2765 5640
rect 2735 5634 2771 5637
rect 2701 5626 2717 5628
rect 2475 5614 2490 5618
rect 2393 5612 2490 5614
rect 2518 5612 2686 5624
rect 2702 5614 2717 5618
rect 2735 5615 2774 5634
rect 2793 5628 2800 5629
rect 2799 5621 2800 5628
rect 2783 5618 2784 5621
rect 2799 5618 2812 5621
rect 2735 5614 2765 5615
rect 2774 5614 2780 5615
rect 2783 5614 2812 5618
rect 2702 5613 2812 5614
rect 2702 5612 2818 5613
rect 2377 5604 2428 5612
rect 2377 5592 2402 5604
rect 2409 5592 2428 5604
rect 2459 5604 2509 5612
rect 2459 5596 2475 5604
rect 2482 5602 2509 5604
rect 2518 5602 2739 5612
rect 2482 5592 2739 5602
rect 2768 5604 2818 5612
rect 2768 5595 2784 5604
rect 2377 5584 2428 5592
rect 2475 5584 2739 5592
rect 2765 5592 2784 5595
rect 2791 5592 2818 5604
rect 2765 5584 2818 5592
rect 2393 5576 2394 5584
rect 2409 5576 2422 5584
rect 2393 5568 2409 5576
rect 2390 5561 2409 5564
rect 2390 5552 2412 5561
rect 2363 5542 2412 5552
rect 2363 5536 2393 5542
rect 2412 5537 2417 5542
rect 2335 5520 2409 5536
rect 2427 5528 2457 5584
rect 2492 5574 2700 5584
rect 2735 5580 2780 5584
rect 2783 5583 2784 5584
rect 2799 5583 2812 5584
rect 2518 5544 2707 5574
rect 2533 5541 2707 5544
rect 2526 5538 2707 5541
rect 2335 5518 2348 5520
rect 2363 5518 2397 5520
rect 2335 5502 2409 5518
rect 2436 5514 2449 5528
rect 2464 5514 2480 5530
rect 2526 5525 2537 5538
rect 2319 5480 2320 5496
rect 2335 5480 2348 5502
rect 2363 5480 2393 5502
rect 2436 5498 2498 5514
rect 2526 5507 2537 5523
rect 2542 5518 2552 5538
rect 2562 5518 2576 5538
rect 2579 5525 2588 5538
rect 2604 5525 2613 5538
rect 2542 5507 2576 5518
rect 2579 5507 2588 5523
rect 2604 5507 2613 5523
rect 2620 5518 2630 5538
rect 2640 5518 2654 5538
rect 2655 5525 2666 5538
rect 2620 5507 2654 5518
rect 2655 5507 2666 5523
rect 2712 5514 2728 5530
rect 2735 5528 2765 5580
rect 2799 5576 2800 5583
rect 2784 5568 2800 5576
rect 2771 5536 2784 5555
rect 2799 5536 2829 5552
rect 2771 5520 2845 5536
rect 2771 5518 2784 5520
rect 2799 5518 2833 5520
rect 2436 5496 2449 5498
rect 2464 5496 2498 5498
rect 2436 5480 2498 5496
rect 2542 5491 2558 5494
rect 2620 5491 2650 5502
rect 2698 5498 2744 5514
rect 2771 5502 2845 5518
rect 2698 5496 2732 5498
rect 2697 5480 2744 5496
rect 2771 5480 2784 5502
rect 2799 5480 2829 5502
rect 2856 5480 2857 5496
rect 2872 5480 2885 5640
rect 2915 5536 2928 5640
rect 2973 5618 2974 5628
rect 2989 5618 3002 5628
rect 2973 5614 3002 5618
rect 3007 5614 3037 5640
rect 3055 5626 3071 5628
rect 3143 5626 3196 5640
rect 3144 5624 3208 5626
rect 3251 5624 3266 5640
rect 3315 5637 3345 5640
rect 3315 5634 3351 5637
rect 3281 5626 3297 5628
rect 3055 5614 3070 5618
rect 2973 5612 3070 5614
rect 3098 5612 3266 5624
rect 3282 5614 3297 5618
rect 3315 5615 3354 5634
rect 3373 5628 3380 5629
rect 3379 5621 3380 5628
rect 3363 5618 3364 5621
rect 3379 5618 3392 5621
rect 3315 5614 3345 5615
rect 3354 5614 3360 5615
rect 3363 5614 3392 5618
rect 3282 5613 3392 5614
rect 3282 5612 3398 5613
rect 2957 5604 3008 5612
rect 2957 5592 2982 5604
rect 2989 5592 3008 5604
rect 3039 5604 3089 5612
rect 3039 5596 3055 5604
rect 3062 5602 3089 5604
rect 3098 5602 3319 5612
rect 3062 5592 3319 5602
rect 3348 5604 3398 5612
rect 3348 5595 3364 5604
rect 2957 5584 3008 5592
rect 3055 5584 3319 5592
rect 3345 5592 3364 5595
rect 3371 5592 3398 5604
rect 3345 5584 3398 5592
rect 2973 5576 2974 5584
rect 2989 5576 3002 5584
rect 2973 5568 2989 5576
rect 2970 5561 2989 5564
rect 2970 5552 2992 5561
rect 2943 5542 2992 5552
rect 2943 5536 2973 5542
rect 2992 5537 2997 5542
rect 2915 5520 2989 5536
rect 3007 5528 3037 5584
rect 3072 5574 3280 5584
rect 3315 5580 3360 5584
rect 3363 5583 3364 5584
rect 3379 5583 3392 5584
rect 3098 5544 3287 5574
rect 3113 5541 3287 5544
rect 3106 5538 3287 5541
rect 2915 5518 2928 5520
rect 2943 5518 2977 5520
rect 2915 5502 2989 5518
rect 3016 5514 3029 5528
rect 3044 5514 3060 5530
rect 3106 5525 3117 5538
rect 2899 5480 2900 5496
rect 2915 5480 2928 5502
rect 2943 5480 2973 5502
rect 3016 5498 3078 5514
rect 3106 5507 3117 5523
rect 3122 5518 3132 5538
rect 3142 5518 3156 5538
rect 3159 5525 3168 5538
rect 3184 5525 3193 5538
rect 3122 5507 3156 5518
rect 3159 5507 3168 5523
rect 3184 5507 3193 5523
rect 3200 5518 3210 5538
rect 3220 5518 3234 5538
rect 3235 5525 3246 5538
rect 3200 5507 3234 5518
rect 3235 5507 3246 5523
rect 3292 5514 3308 5530
rect 3315 5528 3345 5580
rect 3379 5576 3380 5583
rect 3364 5568 3380 5576
rect 3351 5536 3364 5555
rect 3379 5536 3409 5552
rect 3351 5520 3425 5536
rect 3351 5518 3364 5520
rect 3379 5518 3413 5520
rect 3016 5496 3029 5498
rect 3044 5496 3078 5498
rect 3016 5480 3078 5496
rect 3122 5491 3138 5494
rect 3200 5491 3230 5502
rect 3278 5498 3324 5514
rect 3351 5502 3425 5518
rect 3278 5496 3312 5498
rect 3277 5480 3324 5496
rect 3351 5480 3364 5502
rect 3379 5480 3409 5502
rect 3436 5480 3437 5496
rect 3452 5480 3465 5640
rect 3495 5536 3508 5640
rect 3553 5618 3554 5628
rect 3569 5618 3582 5628
rect 3553 5614 3582 5618
rect 3587 5614 3617 5640
rect 3635 5626 3651 5628
rect 3723 5626 3776 5640
rect 3724 5624 3788 5626
rect 3831 5624 3846 5640
rect 3895 5637 3925 5640
rect 3895 5634 3931 5637
rect 3861 5626 3877 5628
rect 3635 5614 3650 5618
rect 3553 5612 3650 5614
rect 3678 5612 3846 5624
rect 3862 5614 3877 5618
rect 3895 5615 3934 5634
rect 3953 5628 3960 5629
rect 3959 5621 3960 5628
rect 3943 5618 3944 5621
rect 3959 5618 3972 5621
rect 3895 5614 3925 5615
rect 3934 5614 3940 5615
rect 3943 5614 3972 5618
rect 3862 5613 3972 5614
rect 3862 5612 3978 5613
rect 3537 5604 3588 5612
rect 3537 5592 3562 5604
rect 3569 5592 3588 5604
rect 3619 5604 3669 5612
rect 3619 5596 3635 5604
rect 3642 5602 3669 5604
rect 3678 5602 3899 5612
rect 3642 5592 3899 5602
rect 3928 5604 3978 5612
rect 3928 5595 3944 5604
rect 3537 5584 3588 5592
rect 3635 5584 3899 5592
rect 3925 5592 3944 5595
rect 3951 5592 3978 5604
rect 3925 5584 3978 5592
rect 3553 5576 3554 5584
rect 3569 5576 3582 5584
rect 3553 5568 3569 5576
rect 3550 5561 3569 5564
rect 3550 5552 3572 5561
rect 3523 5542 3572 5552
rect 3523 5536 3553 5542
rect 3572 5537 3577 5542
rect 3495 5520 3569 5536
rect 3587 5528 3617 5584
rect 3652 5574 3860 5584
rect 3895 5580 3940 5584
rect 3943 5583 3944 5584
rect 3959 5583 3972 5584
rect 3678 5544 3867 5574
rect 3693 5541 3867 5544
rect 3686 5538 3867 5541
rect 3495 5518 3508 5520
rect 3523 5518 3557 5520
rect 3495 5502 3569 5518
rect 3596 5514 3609 5528
rect 3624 5514 3640 5530
rect 3686 5525 3697 5538
rect 3479 5480 3480 5496
rect 3495 5480 3508 5502
rect 3523 5480 3553 5502
rect 3596 5498 3658 5514
rect 3686 5507 3697 5523
rect 3702 5518 3712 5538
rect 3722 5518 3736 5538
rect 3739 5525 3748 5538
rect 3764 5525 3773 5538
rect 3702 5507 3736 5518
rect 3739 5507 3748 5523
rect 3764 5507 3773 5523
rect 3780 5518 3790 5538
rect 3800 5518 3814 5538
rect 3815 5525 3826 5538
rect 3780 5507 3814 5518
rect 3815 5507 3826 5523
rect 3872 5514 3888 5530
rect 3895 5528 3925 5580
rect 3959 5576 3960 5583
rect 3944 5568 3960 5576
rect 3931 5536 3944 5555
rect 3959 5536 3989 5552
rect 3931 5520 4005 5536
rect 3931 5518 3944 5520
rect 3959 5518 3993 5520
rect 3596 5496 3609 5498
rect 3624 5496 3658 5498
rect 3596 5480 3658 5496
rect 3702 5491 3718 5494
rect 3780 5491 3810 5502
rect 3858 5498 3904 5514
rect 3931 5502 4005 5518
rect 3858 5496 3892 5498
rect 3857 5480 3904 5496
rect 3931 5480 3944 5502
rect 3959 5480 3989 5502
rect 4016 5480 4017 5496
rect 4032 5480 4045 5640
rect 4075 5536 4088 5640
rect 4133 5618 4134 5628
rect 4149 5618 4162 5628
rect 4133 5614 4162 5618
rect 4167 5614 4197 5640
rect 4215 5626 4231 5628
rect 4303 5626 4356 5640
rect 4304 5624 4368 5626
rect 4411 5624 4426 5640
rect 4475 5637 4505 5640
rect 4475 5634 4511 5637
rect 4441 5626 4457 5628
rect 4215 5614 4230 5618
rect 4133 5612 4230 5614
rect 4258 5612 4426 5624
rect 4442 5614 4457 5618
rect 4475 5615 4514 5634
rect 4533 5628 4540 5629
rect 4539 5621 4540 5628
rect 4523 5618 4524 5621
rect 4539 5618 4552 5621
rect 4475 5614 4505 5615
rect 4514 5614 4520 5615
rect 4523 5614 4552 5618
rect 4442 5613 4552 5614
rect 4442 5612 4558 5613
rect 4117 5604 4168 5612
rect 4117 5592 4142 5604
rect 4149 5592 4168 5604
rect 4199 5604 4249 5612
rect 4199 5596 4215 5604
rect 4222 5602 4249 5604
rect 4258 5602 4479 5612
rect 4222 5592 4479 5602
rect 4508 5604 4558 5612
rect 4508 5595 4524 5604
rect 4117 5584 4168 5592
rect 4215 5584 4479 5592
rect 4505 5592 4524 5595
rect 4531 5592 4558 5604
rect 4505 5584 4558 5592
rect 4133 5576 4134 5584
rect 4149 5576 4162 5584
rect 4133 5568 4149 5576
rect 4130 5561 4149 5564
rect 4130 5552 4152 5561
rect 4103 5542 4152 5552
rect 4103 5536 4133 5542
rect 4152 5537 4157 5542
rect 4075 5520 4149 5536
rect 4167 5528 4197 5584
rect 4232 5574 4440 5584
rect 4475 5580 4520 5584
rect 4523 5583 4524 5584
rect 4539 5583 4552 5584
rect 4258 5544 4447 5574
rect 4273 5541 4447 5544
rect 4266 5538 4447 5541
rect 4075 5518 4088 5520
rect 4103 5518 4137 5520
rect 4075 5502 4149 5518
rect 4176 5514 4189 5528
rect 4204 5514 4220 5530
rect 4266 5525 4277 5538
rect 4059 5480 4060 5496
rect 4075 5480 4088 5502
rect 4103 5480 4133 5502
rect 4176 5498 4238 5514
rect 4266 5507 4277 5523
rect 4282 5518 4292 5538
rect 4302 5518 4316 5538
rect 4319 5525 4328 5538
rect 4344 5525 4353 5538
rect 4282 5507 4316 5518
rect 4319 5507 4328 5523
rect 4344 5507 4353 5523
rect 4360 5518 4370 5538
rect 4380 5518 4394 5538
rect 4395 5525 4406 5538
rect 4360 5507 4394 5518
rect 4395 5507 4406 5523
rect 4452 5514 4468 5530
rect 4475 5528 4505 5580
rect 4539 5576 4540 5583
rect 4524 5568 4540 5576
rect 4511 5536 4524 5555
rect 4539 5536 4569 5552
rect 4511 5520 4585 5536
rect 4511 5518 4524 5520
rect 4539 5518 4573 5520
rect 4176 5496 4189 5498
rect 4204 5496 4238 5498
rect 4176 5480 4238 5496
rect 4282 5491 4298 5494
rect 4360 5491 4390 5502
rect 4438 5498 4484 5514
rect 4511 5502 4585 5518
rect 4438 5496 4472 5498
rect 4437 5480 4484 5496
rect 4511 5480 4524 5502
rect 4539 5480 4569 5502
rect 4596 5480 4597 5496
rect 4612 5480 4625 5640
rect -7 5472 34 5480
rect -7 5446 8 5472
rect 15 5446 34 5472
rect 98 5468 160 5480
rect 172 5468 247 5480
rect 305 5468 380 5480
rect 392 5468 423 5480
rect 429 5468 464 5480
rect 98 5466 260 5468
rect -7 5438 34 5446
rect 116 5442 129 5466
rect 144 5464 159 5466
rect -1 5428 0 5438
rect 15 5428 28 5438
rect 43 5428 73 5442
rect 116 5428 159 5442
rect 183 5439 190 5446
rect 193 5442 260 5466
rect 292 5466 464 5468
rect 262 5444 290 5448
rect 292 5444 372 5466
rect 393 5464 408 5466
rect 262 5442 372 5444
rect 193 5438 372 5442
rect 166 5428 196 5438
rect 198 5428 351 5438
rect 359 5428 389 5438
rect 393 5428 423 5442
rect 451 5428 464 5466
rect 536 5472 571 5480
rect 536 5446 537 5472
rect 544 5446 571 5472
rect 479 5428 509 5442
rect 536 5438 571 5446
rect 573 5472 614 5480
rect 573 5446 588 5472
rect 595 5446 614 5472
rect 678 5468 740 5480
rect 752 5468 827 5480
rect 885 5468 960 5480
rect 972 5468 1003 5480
rect 1009 5468 1044 5480
rect 678 5466 840 5468
rect 573 5438 614 5446
rect 696 5442 709 5466
rect 724 5464 739 5466
rect 536 5428 537 5438
rect 552 5428 565 5438
rect 579 5428 580 5438
rect 595 5428 608 5438
rect 623 5428 653 5442
rect 696 5428 739 5442
rect 763 5439 770 5446
rect 773 5442 840 5466
rect 872 5466 1044 5468
rect 842 5444 870 5448
rect 872 5444 952 5466
rect 973 5464 988 5466
rect 842 5442 952 5444
rect 773 5438 952 5442
rect 746 5428 776 5438
rect 778 5428 931 5438
rect 939 5428 969 5438
rect 973 5428 1003 5442
rect 1031 5428 1044 5466
rect 1116 5472 1151 5480
rect 1116 5446 1117 5472
rect 1124 5446 1151 5472
rect 1059 5428 1089 5442
rect 1116 5438 1151 5446
rect 1153 5472 1194 5480
rect 1153 5446 1168 5472
rect 1175 5446 1194 5472
rect 1258 5468 1320 5480
rect 1332 5468 1407 5480
rect 1465 5468 1540 5480
rect 1552 5468 1583 5480
rect 1589 5468 1624 5480
rect 1258 5466 1420 5468
rect 1153 5438 1194 5446
rect 1276 5442 1289 5466
rect 1304 5464 1319 5466
rect 1116 5428 1117 5438
rect 1132 5428 1145 5438
rect 1159 5428 1160 5438
rect 1175 5428 1188 5438
rect 1203 5428 1233 5442
rect 1276 5428 1319 5442
rect 1343 5439 1350 5446
rect 1353 5442 1420 5466
rect 1452 5466 1624 5468
rect 1422 5444 1450 5448
rect 1452 5444 1532 5466
rect 1553 5464 1568 5466
rect 1422 5442 1532 5444
rect 1353 5438 1532 5442
rect 1326 5428 1356 5438
rect 1358 5428 1511 5438
rect 1519 5428 1549 5438
rect 1553 5428 1583 5442
rect 1611 5428 1624 5466
rect 1696 5472 1731 5480
rect 1696 5446 1697 5472
rect 1704 5446 1731 5472
rect 1639 5428 1669 5442
rect 1696 5438 1731 5446
rect 1733 5472 1774 5480
rect 1733 5446 1748 5472
rect 1755 5446 1774 5472
rect 1838 5468 1900 5480
rect 1912 5468 1987 5480
rect 2045 5468 2120 5480
rect 2132 5468 2163 5480
rect 2169 5468 2204 5480
rect 1838 5466 2000 5468
rect 1733 5438 1774 5446
rect 1856 5442 1869 5466
rect 1884 5464 1899 5466
rect 1696 5428 1697 5438
rect 1712 5428 1725 5438
rect 1739 5428 1740 5438
rect 1755 5428 1768 5438
rect 1783 5428 1813 5442
rect 1856 5428 1899 5442
rect 1923 5439 1930 5446
rect 1933 5442 2000 5466
rect 2032 5466 2204 5468
rect 2002 5444 2030 5448
rect 2032 5444 2112 5466
rect 2133 5464 2148 5466
rect 2002 5442 2112 5444
rect 1933 5438 2112 5442
rect 1906 5428 1936 5438
rect 1938 5428 2091 5438
rect 2099 5428 2129 5438
rect 2133 5428 2163 5442
rect 2191 5428 2204 5466
rect 2276 5472 2311 5480
rect 2276 5446 2277 5472
rect 2284 5446 2311 5472
rect 2219 5428 2249 5442
rect 2276 5438 2311 5446
rect 2313 5472 2354 5480
rect 2313 5446 2328 5472
rect 2335 5446 2354 5472
rect 2418 5468 2480 5480
rect 2492 5468 2567 5480
rect 2625 5468 2700 5480
rect 2712 5468 2743 5480
rect 2749 5468 2784 5480
rect 2418 5466 2580 5468
rect 2313 5438 2354 5446
rect 2436 5442 2449 5466
rect 2464 5464 2479 5466
rect 2276 5428 2277 5438
rect 2292 5428 2305 5438
rect 2319 5428 2320 5438
rect 2335 5428 2348 5438
rect 2363 5428 2393 5442
rect 2436 5428 2479 5442
rect 2503 5439 2510 5446
rect 2513 5442 2580 5466
rect 2612 5466 2784 5468
rect 2582 5444 2610 5448
rect 2612 5444 2692 5466
rect 2713 5464 2728 5466
rect 2582 5442 2692 5444
rect 2513 5438 2692 5442
rect 2486 5428 2516 5438
rect 2518 5428 2671 5438
rect 2679 5428 2709 5438
rect 2713 5428 2743 5442
rect 2771 5428 2784 5466
rect 2856 5472 2891 5480
rect 2856 5446 2857 5472
rect 2864 5446 2891 5472
rect 2799 5428 2829 5442
rect 2856 5438 2891 5446
rect 2893 5472 2934 5480
rect 2893 5446 2908 5472
rect 2915 5446 2934 5472
rect 2998 5468 3060 5480
rect 3072 5468 3147 5480
rect 3205 5468 3280 5480
rect 3292 5468 3323 5480
rect 3329 5468 3364 5480
rect 2998 5466 3160 5468
rect 2893 5438 2934 5446
rect 3016 5442 3029 5466
rect 3044 5464 3059 5466
rect 2856 5428 2857 5438
rect 2872 5428 2885 5438
rect 2899 5428 2900 5438
rect 2915 5428 2928 5438
rect 2943 5428 2973 5442
rect 3016 5428 3059 5442
rect 3083 5439 3090 5446
rect 3093 5442 3160 5466
rect 3192 5466 3364 5468
rect 3162 5444 3190 5448
rect 3192 5444 3272 5466
rect 3293 5464 3308 5466
rect 3162 5442 3272 5444
rect 3093 5438 3272 5442
rect 3066 5428 3096 5438
rect 3098 5428 3251 5438
rect 3259 5428 3289 5438
rect 3293 5428 3323 5442
rect 3351 5428 3364 5466
rect 3436 5472 3471 5480
rect 3436 5446 3437 5472
rect 3444 5446 3471 5472
rect 3379 5428 3409 5442
rect 3436 5438 3471 5446
rect 3473 5472 3514 5480
rect 3473 5446 3488 5472
rect 3495 5446 3514 5472
rect 3578 5468 3640 5480
rect 3652 5468 3727 5480
rect 3785 5468 3860 5480
rect 3872 5468 3903 5480
rect 3909 5468 3944 5480
rect 3578 5466 3740 5468
rect 3473 5438 3514 5446
rect 3596 5442 3609 5466
rect 3624 5464 3639 5466
rect 3436 5428 3437 5438
rect 3452 5428 3465 5438
rect 3479 5428 3480 5438
rect 3495 5428 3508 5438
rect 3523 5428 3553 5442
rect 3596 5428 3639 5442
rect 3663 5439 3670 5446
rect 3673 5442 3740 5466
rect 3772 5466 3944 5468
rect 3742 5444 3770 5448
rect 3772 5444 3852 5466
rect 3873 5464 3888 5466
rect 3742 5442 3852 5444
rect 3673 5438 3852 5442
rect 3646 5428 3676 5438
rect 3678 5428 3831 5438
rect 3839 5428 3869 5438
rect 3873 5428 3903 5442
rect 3931 5428 3944 5466
rect 4016 5472 4051 5480
rect 4016 5446 4017 5472
rect 4024 5446 4051 5472
rect 3959 5428 3989 5442
rect 4016 5438 4051 5446
rect 4053 5472 4094 5480
rect 4053 5446 4068 5472
rect 4075 5446 4094 5472
rect 4158 5468 4220 5480
rect 4232 5468 4307 5480
rect 4365 5468 4440 5480
rect 4452 5468 4483 5480
rect 4489 5468 4524 5480
rect 4158 5466 4320 5468
rect 4053 5438 4094 5446
rect 4176 5442 4189 5466
rect 4204 5464 4219 5466
rect 4016 5428 4017 5438
rect 4032 5428 4045 5438
rect 4059 5428 4060 5438
rect 4075 5428 4088 5438
rect 4103 5428 4133 5442
rect 4176 5428 4219 5442
rect 4243 5439 4250 5446
rect 4253 5442 4320 5466
rect 4352 5466 4524 5468
rect 4322 5444 4350 5448
rect 4352 5444 4432 5466
rect 4453 5464 4468 5466
rect 4322 5442 4432 5444
rect 4253 5438 4432 5442
rect 4226 5428 4256 5438
rect 4258 5428 4411 5438
rect 4419 5428 4449 5438
rect 4453 5428 4483 5442
rect 4511 5428 4524 5466
rect 4596 5472 4631 5480
rect 4596 5446 4597 5472
rect 4604 5446 4631 5472
rect 4539 5428 4569 5442
rect 4596 5438 4631 5446
rect 4596 5428 4597 5438
rect 4612 5428 4625 5438
rect -1 5422 4625 5428
rect 0 5414 4625 5422
rect 15 5384 28 5414
rect 43 5396 73 5414
rect 116 5400 130 5414
rect 166 5400 386 5414
rect 117 5398 130 5400
rect 83 5386 98 5398
rect 80 5384 102 5386
rect 107 5384 137 5398
rect 198 5396 351 5400
rect 180 5384 372 5396
rect 415 5384 445 5398
rect 451 5384 464 5414
rect 479 5396 509 5414
rect 552 5384 565 5414
rect 595 5384 608 5414
rect 623 5396 653 5414
rect 696 5400 710 5414
rect 746 5400 966 5414
rect 697 5398 710 5400
rect 663 5386 678 5398
rect 660 5384 682 5386
rect 687 5384 717 5398
rect 778 5396 931 5400
rect 760 5384 952 5396
rect 995 5384 1025 5398
rect 1031 5384 1044 5414
rect 1059 5396 1089 5414
rect 1132 5384 1145 5414
rect 1175 5384 1188 5414
rect 1203 5396 1233 5414
rect 1276 5400 1290 5414
rect 1326 5400 1546 5414
rect 1277 5398 1290 5400
rect 1243 5386 1258 5398
rect 1240 5384 1262 5386
rect 1267 5384 1297 5398
rect 1358 5396 1511 5400
rect 1340 5384 1532 5396
rect 1575 5384 1605 5398
rect 1611 5384 1624 5414
rect 1639 5396 1669 5414
rect 1712 5384 1725 5414
rect 1755 5384 1768 5414
rect 1783 5396 1813 5414
rect 1856 5400 1870 5414
rect 1906 5400 2126 5414
rect 1857 5398 1870 5400
rect 1823 5386 1838 5398
rect 1820 5384 1842 5386
rect 1847 5384 1877 5398
rect 1938 5396 2091 5400
rect 1920 5384 2112 5396
rect 2155 5384 2185 5398
rect 2191 5384 2204 5414
rect 2219 5396 2249 5414
rect 2292 5384 2305 5414
rect 2335 5384 2348 5414
rect 2363 5396 2393 5414
rect 2436 5400 2450 5414
rect 2486 5400 2706 5414
rect 2437 5398 2450 5400
rect 2403 5386 2418 5398
rect 2400 5384 2422 5386
rect 2427 5384 2457 5398
rect 2518 5396 2671 5400
rect 2500 5384 2692 5396
rect 2735 5384 2765 5398
rect 2771 5384 2784 5414
rect 2799 5396 2829 5414
rect 2872 5384 2885 5414
rect 2915 5384 2928 5414
rect 2943 5396 2973 5414
rect 3016 5400 3030 5414
rect 3066 5400 3286 5414
rect 3017 5398 3030 5400
rect 2983 5386 2998 5398
rect 2980 5384 3002 5386
rect 3007 5384 3037 5398
rect 3098 5396 3251 5400
rect 3080 5384 3272 5396
rect 3315 5384 3345 5398
rect 3351 5384 3364 5414
rect 3379 5396 3409 5414
rect 3452 5384 3465 5414
rect 3495 5384 3508 5414
rect 3523 5396 3553 5414
rect 3596 5400 3610 5414
rect 3646 5400 3866 5414
rect 3597 5398 3610 5400
rect 3563 5386 3578 5398
rect 3560 5384 3582 5386
rect 3587 5384 3617 5398
rect 3678 5396 3831 5400
rect 3660 5384 3852 5396
rect 3895 5384 3925 5398
rect 3931 5384 3944 5414
rect 3959 5396 3989 5414
rect 4032 5384 4045 5414
rect 4075 5384 4088 5414
rect 4103 5396 4133 5414
rect 4176 5400 4190 5414
rect 4226 5400 4446 5414
rect 4177 5398 4190 5400
rect 4143 5386 4158 5398
rect 4140 5384 4162 5386
rect 4167 5384 4197 5398
rect 4258 5396 4411 5400
rect 4240 5384 4432 5396
rect 4475 5384 4505 5398
rect 4511 5384 4524 5414
rect 4539 5396 4569 5414
rect 4612 5384 4625 5414
rect 0 5370 4625 5384
rect 15 5266 28 5370
rect 73 5348 74 5358
rect 89 5348 102 5358
rect 73 5344 102 5348
rect 107 5344 137 5370
rect 155 5356 171 5358
rect 243 5356 296 5370
rect 244 5354 308 5356
rect 351 5354 366 5370
rect 415 5367 445 5370
rect 415 5364 451 5367
rect 381 5356 397 5358
rect 155 5344 170 5348
rect 73 5342 170 5344
rect 198 5342 366 5354
rect 382 5344 397 5348
rect 415 5345 454 5364
rect 473 5358 480 5359
rect 479 5351 480 5358
rect 463 5348 464 5351
rect 479 5348 492 5351
rect 415 5344 445 5345
rect 454 5344 460 5345
rect 463 5344 492 5348
rect 382 5343 492 5344
rect 382 5342 498 5343
rect 57 5334 108 5342
rect 57 5322 82 5334
rect 89 5322 108 5334
rect 139 5334 189 5342
rect 139 5326 155 5334
rect 162 5332 189 5334
rect 198 5332 419 5342
rect 162 5322 419 5332
rect 448 5334 498 5342
rect 448 5325 464 5334
rect 57 5314 108 5322
rect 155 5314 419 5322
rect 445 5322 464 5325
rect 471 5322 498 5334
rect 445 5314 498 5322
rect 73 5306 74 5314
rect 89 5306 102 5314
rect 73 5298 89 5306
rect 70 5291 89 5294
rect 70 5282 92 5291
rect 43 5272 92 5282
rect 43 5266 73 5272
rect 92 5267 97 5272
rect 15 5250 89 5266
rect 107 5258 137 5314
rect 172 5304 380 5314
rect 415 5310 460 5314
rect 463 5313 464 5314
rect 479 5313 492 5314
rect 198 5274 387 5304
rect 213 5271 387 5274
rect 206 5268 387 5271
rect 15 5248 28 5250
rect 43 5248 77 5250
rect 15 5232 89 5248
rect 116 5244 129 5258
rect 144 5244 160 5260
rect 206 5255 217 5268
rect -1 5210 0 5226
rect 15 5210 28 5232
rect 43 5210 73 5232
rect 116 5228 178 5244
rect 206 5237 217 5253
rect 222 5248 232 5268
rect 242 5248 256 5268
rect 259 5255 268 5268
rect 284 5255 293 5268
rect 222 5237 256 5248
rect 259 5237 268 5253
rect 284 5237 293 5253
rect 300 5248 310 5268
rect 320 5248 334 5268
rect 335 5255 346 5268
rect 300 5237 334 5248
rect 335 5237 346 5253
rect 392 5244 408 5260
rect 415 5258 445 5310
rect 479 5306 480 5313
rect 464 5298 480 5306
rect 451 5266 464 5285
rect 479 5266 509 5282
rect 451 5250 525 5266
rect 451 5248 464 5250
rect 479 5248 513 5250
rect 116 5226 129 5228
rect 144 5226 178 5228
rect 116 5210 178 5226
rect 222 5221 238 5224
rect 300 5221 330 5232
rect 378 5228 424 5244
rect 451 5232 525 5248
rect 378 5226 412 5228
rect 377 5210 424 5226
rect 451 5210 464 5232
rect 479 5210 509 5232
rect 536 5210 537 5226
rect 552 5210 565 5370
rect 595 5266 608 5370
rect 653 5348 654 5358
rect 669 5348 682 5358
rect 653 5344 682 5348
rect 687 5344 717 5370
rect 735 5356 751 5358
rect 823 5356 876 5370
rect 824 5354 888 5356
rect 931 5354 946 5370
rect 995 5367 1025 5370
rect 995 5364 1031 5367
rect 961 5356 977 5358
rect 735 5344 750 5348
rect 653 5342 750 5344
rect 778 5342 946 5354
rect 962 5344 977 5348
rect 995 5345 1034 5364
rect 1053 5358 1060 5359
rect 1059 5351 1060 5358
rect 1043 5348 1044 5351
rect 1059 5348 1072 5351
rect 995 5344 1025 5345
rect 1034 5344 1040 5345
rect 1043 5344 1072 5348
rect 962 5343 1072 5344
rect 962 5342 1078 5343
rect 637 5334 688 5342
rect 637 5322 662 5334
rect 669 5322 688 5334
rect 719 5334 769 5342
rect 719 5326 735 5334
rect 742 5332 769 5334
rect 778 5332 999 5342
rect 742 5322 999 5332
rect 1028 5334 1078 5342
rect 1028 5325 1044 5334
rect 637 5314 688 5322
rect 735 5314 999 5322
rect 1025 5322 1044 5325
rect 1051 5322 1078 5334
rect 1025 5314 1078 5322
rect 653 5306 654 5314
rect 669 5306 682 5314
rect 653 5298 669 5306
rect 650 5291 669 5294
rect 650 5282 672 5291
rect 623 5272 672 5282
rect 623 5266 653 5272
rect 672 5267 677 5272
rect 595 5250 669 5266
rect 687 5258 717 5314
rect 752 5304 960 5314
rect 995 5310 1040 5314
rect 1043 5313 1044 5314
rect 1059 5313 1072 5314
rect 778 5274 967 5304
rect 793 5271 967 5274
rect 786 5268 967 5271
rect 595 5248 608 5250
rect 623 5248 657 5250
rect 595 5232 669 5248
rect 696 5244 709 5258
rect 724 5244 740 5260
rect 786 5255 797 5268
rect 579 5210 580 5226
rect 595 5210 608 5232
rect 623 5210 653 5232
rect 696 5228 758 5244
rect 786 5237 797 5253
rect 802 5248 812 5268
rect 822 5248 836 5268
rect 839 5255 848 5268
rect 864 5255 873 5268
rect 802 5237 836 5248
rect 839 5237 848 5253
rect 864 5237 873 5253
rect 880 5248 890 5268
rect 900 5248 914 5268
rect 915 5255 926 5268
rect 880 5237 914 5248
rect 915 5237 926 5253
rect 972 5244 988 5260
rect 995 5258 1025 5310
rect 1059 5306 1060 5313
rect 1044 5298 1060 5306
rect 1031 5266 1044 5285
rect 1059 5266 1089 5282
rect 1031 5250 1105 5266
rect 1031 5248 1044 5250
rect 1059 5248 1093 5250
rect 696 5226 709 5228
rect 724 5226 758 5228
rect 696 5210 758 5226
rect 802 5221 818 5224
rect 880 5221 910 5232
rect 958 5228 1004 5244
rect 1031 5232 1105 5248
rect 958 5226 992 5228
rect 957 5210 1004 5226
rect 1031 5210 1044 5232
rect 1059 5210 1089 5232
rect 1116 5210 1117 5226
rect 1132 5210 1145 5370
rect 1175 5266 1188 5370
rect 1233 5348 1234 5358
rect 1249 5348 1262 5358
rect 1233 5344 1262 5348
rect 1267 5344 1297 5370
rect 1315 5356 1331 5358
rect 1403 5356 1456 5370
rect 1404 5354 1468 5356
rect 1511 5354 1526 5370
rect 1575 5367 1605 5370
rect 1575 5364 1611 5367
rect 1541 5356 1557 5358
rect 1315 5344 1330 5348
rect 1233 5342 1330 5344
rect 1358 5342 1526 5354
rect 1542 5344 1557 5348
rect 1575 5345 1614 5364
rect 1633 5358 1640 5359
rect 1639 5351 1640 5358
rect 1623 5348 1624 5351
rect 1639 5348 1652 5351
rect 1575 5344 1605 5345
rect 1614 5344 1620 5345
rect 1623 5344 1652 5348
rect 1542 5343 1652 5344
rect 1542 5342 1658 5343
rect 1217 5334 1268 5342
rect 1217 5322 1242 5334
rect 1249 5322 1268 5334
rect 1299 5334 1349 5342
rect 1299 5326 1315 5334
rect 1322 5332 1349 5334
rect 1358 5332 1579 5342
rect 1322 5322 1579 5332
rect 1608 5334 1658 5342
rect 1608 5325 1624 5334
rect 1217 5314 1268 5322
rect 1315 5314 1579 5322
rect 1605 5322 1624 5325
rect 1631 5322 1658 5334
rect 1605 5314 1658 5322
rect 1233 5306 1234 5314
rect 1249 5306 1262 5314
rect 1233 5298 1249 5306
rect 1230 5291 1249 5294
rect 1230 5282 1252 5291
rect 1203 5272 1252 5282
rect 1203 5266 1233 5272
rect 1252 5267 1257 5272
rect 1175 5250 1249 5266
rect 1267 5258 1297 5314
rect 1332 5304 1540 5314
rect 1575 5310 1620 5314
rect 1623 5313 1624 5314
rect 1639 5313 1652 5314
rect 1358 5274 1547 5304
rect 1373 5271 1547 5274
rect 1366 5268 1547 5271
rect 1175 5248 1188 5250
rect 1203 5248 1237 5250
rect 1175 5232 1249 5248
rect 1276 5244 1289 5258
rect 1304 5244 1320 5260
rect 1366 5255 1377 5268
rect 1159 5210 1160 5226
rect 1175 5210 1188 5232
rect 1203 5210 1233 5232
rect 1276 5228 1338 5244
rect 1366 5237 1377 5253
rect 1382 5248 1392 5268
rect 1402 5248 1416 5268
rect 1419 5255 1428 5268
rect 1444 5255 1453 5268
rect 1382 5237 1416 5248
rect 1419 5237 1428 5253
rect 1444 5237 1453 5253
rect 1460 5248 1470 5268
rect 1480 5248 1494 5268
rect 1495 5255 1506 5268
rect 1460 5237 1494 5248
rect 1495 5237 1506 5253
rect 1552 5244 1568 5260
rect 1575 5258 1605 5310
rect 1639 5306 1640 5313
rect 1624 5298 1640 5306
rect 1611 5266 1624 5285
rect 1639 5266 1669 5282
rect 1611 5250 1685 5266
rect 1611 5248 1624 5250
rect 1639 5248 1673 5250
rect 1276 5226 1289 5228
rect 1304 5226 1338 5228
rect 1276 5210 1338 5226
rect 1382 5221 1398 5224
rect 1460 5221 1490 5232
rect 1538 5228 1584 5244
rect 1611 5232 1685 5248
rect 1538 5226 1572 5228
rect 1537 5210 1584 5226
rect 1611 5210 1624 5232
rect 1639 5210 1669 5232
rect 1696 5210 1697 5226
rect 1712 5210 1725 5370
rect 1755 5266 1768 5370
rect 1813 5348 1814 5358
rect 1829 5348 1842 5358
rect 1813 5344 1842 5348
rect 1847 5344 1877 5370
rect 1895 5356 1911 5358
rect 1983 5356 2036 5370
rect 1984 5354 2048 5356
rect 2091 5354 2106 5370
rect 2155 5367 2185 5370
rect 2155 5364 2191 5367
rect 2121 5356 2137 5358
rect 1895 5344 1910 5348
rect 1813 5342 1910 5344
rect 1938 5342 2106 5354
rect 2122 5344 2137 5348
rect 2155 5345 2194 5364
rect 2213 5358 2220 5359
rect 2219 5351 2220 5358
rect 2203 5348 2204 5351
rect 2219 5348 2232 5351
rect 2155 5344 2185 5345
rect 2194 5344 2200 5345
rect 2203 5344 2232 5348
rect 2122 5343 2232 5344
rect 2122 5342 2238 5343
rect 1797 5334 1848 5342
rect 1797 5322 1822 5334
rect 1829 5322 1848 5334
rect 1879 5334 1929 5342
rect 1879 5326 1895 5334
rect 1902 5332 1929 5334
rect 1938 5332 2159 5342
rect 1902 5322 2159 5332
rect 2188 5334 2238 5342
rect 2188 5325 2204 5334
rect 1797 5314 1848 5322
rect 1895 5314 2159 5322
rect 2185 5322 2204 5325
rect 2211 5322 2238 5334
rect 2185 5314 2238 5322
rect 1813 5306 1814 5314
rect 1829 5306 1842 5314
rect 1813 5298 1829 5306
rect 1810 5291 1829 5294
rect 1810 5282 1832 5291
rect 1783 5272 1832 5282
rect 1783 5266 1813 5272
rect 1832 5267 1837 5272
rect 1755 5250 1829 5266
rect 1847 5258 1877 5314
rect 1912 5304 2120 5314
rect 2155 5310 2200 5314
rect 2203 5313 2204 5314
rect 2219 5313 2232 5314
rect 1938 5274 2127 5304
rect 1953 5271 2127 5274
rect 1946 5268 2127 5271
rect 1755 5248 1768 5250
rect 1783 5248 1817 5250
rect 1755 5232 1829 5248
rect 1856 5244 1869 5258
rect 1884 5244 1900 5260
rect 1946 5255 1957 5268
rect 1739 5210 1740 5226
rect 1755 5210 1768 5232
rect 1783 5210 1813 5232
rect 1856 5228 1918 5244
rect 1946 5237 1957 5253
rect 1962 5248 1972 5268
rect 1982 5248 1996 5268
rect 1999 5255 2008 5268
rect 2024 5255 2033 5268
rect 1962 5237 1996 5248
rect 1999 5237 2008 5253
rect 2024 5237 2033 5253
rect 2040 5248 2050 5268
rect 2060 5248 2074 5268
rect 2075 5255 2086 5268
rect 2040 5237 2074 5248
rect 2075 5237 2086 5253
rect 2132 5244 2148 5260
rect 2155 5258 2185 5310
rect 2219 5306 2220 5313
rect 2204 5298 2220 5306
rect 2191 5266 2204 5285
rect 2219 5266 2249 5282
rect 2191 5250 2265 5266
rect 2191 5248 2204 5250
rect 2219 5248 2253 5250
rect 1856 5226 1869 5228
rect 1884 5226 1918 5228
rect 1856 5210 1918 5226
rect 1962 5221 1978 5224
rect 2040 5221 2070 5232
rect 2118 5228 2164 5244
rect 2191 5232 2265 5248
rect 2118 5226 2152 5228
rect 2117 5210 2164 5226
rect 2191 5210 2204 5232
rect 2219 5210 2249 5232
rect 2276 5210 2277 5226
rect 2292 5210 2305 5370
rect 2335 5266 2348 5370
rect 2393 5348 2394 5358
rect 2409 5348 2422 5358
rect 2393 5344 2422 5348
rect 2427 5344 2457 5370
rect 2475 5356 2491 5358
rect 2563 5356 2616 5370
rect 2564 5354 2628 5356
rect 2671 5354 2686 5370
rect 2735 5367 2765 5370
rect 2735 5364 2771 5367
rect 2701 5356 2717 5358
rect 2475 5344 2490 5348
rect 2393 5342 2490 5344
rect 2518 5342 2686 5354
rect 2702 5344 2717 5348
rect 2735 5345 2774 5364
rect 2793 5358 2800 5359
rect 2799 5351 2800 5358
rect 2783 5348 2784 5351
rect 2799 5348 2812 5351
rect 2735 5344 2765 5345
rect 2774 5344 2780 5345
rect 2783 5344 2812 5348
rect 2702 5343 2812 5344
rect 2702 5342 2818 5343
rect 2377 5334 2428 5342
rect 2377 5322 2402 5334
rect 2409 5322 2428 5334
rect 2459 5334 2509 5342
rect 2459 5326 2475 5334
rect 2482 5332 2509 5334
rect 2518 5332 2739 5342
rect 2482 5322 2739 5332
rect 2768 5334 2818 5342
rect 2768 5325 2784 5334
rect 2377 5314 2428 5322
rect 2475 5314 2739 5322
rect 2765 5322 2784 5325
rect 2791 5322 2818 5334
rect 2765 5314 2818 5322
rect 2393 5306 2394 5314
rect 2409 5306 2422 5314
rect 2393 5298 2409 5306
rect 2390 5291 2409 5294
rect 2390 5282 2412 5291
rect 2363 5272 2412 5282
rect 2363 5266 2393 5272
rect 2412 5267 2417 5272
rect 2335 5250 2409 5266
rect 2427 5258 2457 5314
rect 2492 5304 2700 5314
rect 2735 5310 2780 5314
rect 2783 5313 2784 5314
rect 2799 5313 2812 5314
rect 2518 5274 2707 5304
rect 2533 5271 2707 5274
rect 2526 5268 2707 5271
rect 2335 5248 2348 5250
rect 2363 5248 2397 5250
rect 2335 5232 2409 5248
rect 2436 5244 2449 5258
rect 2464 5244 2480 5260
rect 2526 5255 2537 5268
rect 2319 5210 2320 5226
rect 2335 5210 2348 5232
rect 2363 5210 2393 5232
rect 2436 5228 2498 5244
rect 2526 5237 2537 5253
rect 2542 5248 2552 5268
rect 2562 5248 2576 5268
rect 2579 5255 2588 5268
rect 2604 5255 2613 5268
rect 2542 5237 2576 5248
rect 2579 5237 2588 5253
rect 2604 5237 2613 5253
rect 2620 5248 2630 5268
rect 2640 5248 2654 5268
rect 2655 5255 2666 5268
rect 2620 5237 2654 5248
rect 2655 5237 2666 5253
rect 2712 5244 2728 5260
rect 2735 5258 2765 5310
rect 2799 5306 2800 5313
rect 2784 5298 2800 5306
rect 2771 5266 2784 5285
rect 2799 5266 2829 5282
rect 2771 5250 2845 5266
rect 2771 5248 2784 5250
rect 2799 5248 2833 5250
rect 2436 5226 2449 5228
rect 2464 5226 2498 5228
rect 2436 5210 2498 5226
rect 2542 5221 2558 5224
rect 2620 5221 2650 5232
rect 2698 5228 2744 5244
rect 2771 5232 2845 5248
rect 2698 5226 2732 5228
rect 2697 5210 2744 5226
rect 2771 5210 2784 5232
rect 2799 5210 2829 5232
rect 2856 5210 2857 5226
rect 2872 5210 2885 5370
rect 2915 5266 2928 5370
rect 2973 5348 2974 5358
rect 2989 5348 3002 5358
rect 2973 5344 3002 5348
rect 3007 5344 3037 5370
rect 3055 5356 3071 5358
rect 3143 5356 3196 5370
rect 3144 5354 3208 5356
rect 3251 5354 3266 5370
rect 3315 5367 3345 5370
rect 3315 5364 3351 5367
rect 3281 5356 3297 5358
rect 3055 5344 3070 5348
rect 2973 5342 3070 5344
rect 3098 5342 3266 5354
rect 3282 5344 3297 5348
rect 3315 5345 3354 5364
rect 3373 5358 3380 5359
rect 3379 5351 3380 5358
rect 3363 5348 3364 5351
rect 3379 5348 3392 5351
rect 3315 5344 3345 5345
rect 3354 5344 3360 5345
rect 3363 5344 3392 5348
rect 3282 5343 3392 5344
rect 3282 5342 3398 5343
rect 2957 5334 3008 5342
rect 2957 5322 2982 5334
rect 2989 5322 3008 5334
rect 3039 5334 3089 5342
rect 3039 5326 3055 5334
rect 3062 5332 3089 5334
rect 3098 5332 3319 5342
rect 3062 5322 3319 5332
rect 3348 5334 3398 5342
rect 3348 5325 3364 5334
rect 2957 5314 3008 5322
rect 3055 5314 3319 5322
rect 3345 5322 3364 5325
rect 3371 5322 3398 5334
rect 3345 5314 3398 5322
rect 2973 5306 2974 5314
rect 2989 5306 3002 5314
rect 2973 5298 2989 5306
rect 2970 5291 2989 5294
rect 2970 5282 2992 5291
rect 2943 5272 2992 5282
rect 2943 5266 2973 5272
rect 2992 5267 2997 5272
rect 2915 5250 2989 5266
rect 3007 5258 3037 5314
rect 3072 5304 3280 5314
rect 3315 5310 3360 5314
rect 3363 5313 3364 5314
rect 3379 5313 3392 5314
rect 3098 5274 3287 5304
rect 3113 5271 3287 5274
rect 3106 5268 3287 5271
rect 2915 5248 2928 5250
rect 2943 5248 2977 5250
rect 2915 5232 2989 5248
rect 3016 5244 3029 5258
rect 3044 5244 3060 5260
rect 3106 5255 3117 5268
rect 2899 5210 2900 5226
rect 2915 5210 2928 5232
rect 2943 5210 2973 5232
rect 3016 5228 3078 5244
rect 3106 5237 3117 5253
rect 3122 5248 3132 5268
rect 3142 5248 3156 5268
rect 3159 5255 3168 5268
rect 3184 5255 3193 5268
rect 3122 5237 3156 5248
rect 3159 5237 3168 5253
rect 3184 5237 3193 5253
rect 3200 5248 3210 5268
rect 3220 5248 3234 5268
rect 3235 5255 3246 5268
rect 3200 5237 3234 5248
rect 3235 5237 3246 5253
rect 3292 5244 3308 5260
rect 3315 5258 3345 5310
rect 3379 5306 3380 5313
rect 3364 5298 3380 5306
rect 3351 5266 3364 5285
rect 3379 5266 3409 5282
rect 3351 5250 3425 5266
rect 3351 5248 3364 5250
rect 3379 5248 3413 5250
rect 3016 5226 3029 5228
rect 3044 5226 3078 5228
rect 3016 5210 3078 5226
rect 3122 5221 3138 5224
rect 3200 5221 3230 5232
rect 3278 5228 3324 5244
rect 3351 5232 3425 5248
rect 3278 5226 3312 5228
rect 3277 5210 3324 5226
rect 3351 5210 3364 5232
rect 3379 5210 3409 5232
rect 3436 5210 3437 5226
rect 3452 5210 3465 5370
rect 3495 5266 3508 5370
rect 3553 5348 3554 5358
rect 3569 5348 3582 5358
rect 3553 5344 3582 5348
rect 3587 5344 3617 5370
rect 3635 5356 3651 5358
rect 3723 5356 3776 5370
rect 3724 5354 3788 5356
rect 3831 5354 3846 5370
rect 3895 5367 3925 5370
rect 3895 5364 3931 5367
rect 3861 5356 3877 5358
rect 3635 5344 3650 5348
rect 3553 5342 3650 5344
rect 3678 5342 3846 5354
rect 3862 5344 3877 5348
rect 3895 5345 3934 5364
rect 3953 5358 3960 5359
rect 3959 5351 3960 5358
rect 3943 5348 3944 5351
rect 3959 5348 3972 5351
rect 3895 5344 3925 5345
rect 3934 5344 3940 5345
rect 3943 5344 3972 5348
rect 3862 5343 3972 5344
rect 3862 5342 3978 5343
rect 3537 5334 3588 5342
rect 3537 5322 3562 5334
rect 3569 5322 3588 5334
rect 3619 5334 3669 5342
rect 3619 5326 3635 5334
rect 3642 5332 3669 5334
rect 3678 5332 3899 5342
rect 3642 5322 3899 5332
rect 3928 5334 3978 5342
rect 3928 5325 3944 5334
rect 3537 5314 3588 5322
rect 3635 5314 3899 5322
rect 3925 5322 3944 5325
rect 3951 5322 3978 5334
rect 3925 5314 3978 5322
rect 3553 5306 3554 5314
rect 3569 5306 3582 5314
rect 3553 5298 3569 5306
rect 3550 5291 3569 5294
rect 3550 5282 3572 5291
rect 3523 5272 3572 5282
rect 3523 5266 3553 5272
rect 3572 5267 3577 5272
rect 3495 5250 3569 5266
rect 3587 5258 3617 5314
rect 3652 5304 3860 5314
rect 3895 5310 3940 5314
rect 3943 5313 3944 5314
rect 3959 5313 3972 5314
rect 3678 5274 3867 5304
rect 3693 5271 3867 5274
rect 3686 5268 3867 5271
rect 3495 5248 3508 5250
rect 3523 5248 3557 5250
rect 3495 5232 3569 5248
rect 3596 5244 3609 5258
rect 3624 5244 3640 5260
rect 3686 5255 3697 5268
rect 3479 5210 3480 5226
rect 3495 5210 3508 5232
rect 3523 5210 3553 5232
rect 3596 5228 3658 5244
rect 3686 5237 3697 5253
rect 3702 5248 3712 5268
rect 3722 5248 3736 5268
rect 3739 5255 3748 5268
rect 3764 5255 3773 5268
rect 3702 5237 3736 5248
rect 3739 5237 3748 5253
rect 3764 5237 3773 5253
rect 3780 5248 3790 5268
rect 3800 5248 3814 5268
rect 3815 5255 3826 5268
rect 3780 5237 3814 5248
rect 3815 5237 3826 5253
rect 3872 5244 3888 5260
rect 3895 5258 3925 5310
rect 3959 5306 3960 5313
rect 3944 5298 3960 5306
rect 3931 5266 3944 5285
rect 3959 5266 3989 5282
rect 3931 5250 4005 5266
rect 3931 5248 3944 5250
rect 3959 5248 3993 5250
rect 3596 5226 3609 5228
rect 3624 5226 3658 5228
rect 3596 5210 3658 5226
rect 3702 5221 3718 5224
rect 3780 5221 3810 5232
rect 3858 5228 3904 5244
rect 3931 5232 4005 5248
rect 3858 5226 3892 5228
rect 3857 5210 3904 5226
rect 3931 5210 3944 5232
rect 3959 5210 3989 5232
rect 4016 5210 4017 5226
rect 4032 5210 4045 5370
rect 4075 5266 4088 5370
rect 4133 5348 4134 5358
rect 4149 5348 4162 5358
rect 4133 5344 4162 5348
rect 4167 5344 4197 5370
rect 4215 5356 4231 5358
rect 4303 5356 4356 5370
rect 4304 5354 4368 5356
rect 4411 5354 4426 5370
rect 4475 5367 4505 5370
rect 4475 5364 4511 5367
rect 4441 5356 4457 5358
rect 4215 5344 4230 5348
rect 4133 5342 4230 5344
rect 4258 5342 4426 5354
rect 4442 5344 4457 5348
rect 4475 5345 4514 5364
rect 4533 5358 4540 5359
rect 4539 5351 4540 5358
rect 4523 5348 4524 5351
rect 4539 5348 4552 5351
rect 4475 5344 4505 5345
rect 4514 5344 4520 5345
rect 4523 5344 4552 5348
rect 4442 5343 4552 5344
rect 4442 5342 4558 5343
rect 4117 5334 4168 5342
rect 4117 5322 4142 5334
rect 4149 5322 4168 5334
rect 4199 5334 4249 5342
rect 4199 5326 4215 5334
rect 4222 5332 4249 5334
rect 4258 5332 4479 5342
rect 4222 5322 4479 5332
rect 4508 5334 4558 5342
rect 4508 5325 4524 5334
rect 4117 5314 4168 5322
rect 4215 5314 4479 5322
rect 4505 5322 4524 5325
rect 4531 5322 4558 5334
rect 4505 5314 4558 5322
rect 4133 5306 4134 5314
rect 4149 5306 4162 5314
rect 4133 5298 4149 5306
rect 4130 5291 4149 5294
rect 4130 5282 4152 5291
rect 4103 5272 4152 5282
rect 4103 5266 4133 5272
rect 4152 5267 4157 5272
rect 4075 5250 4149 5266
rect 4167 5258 4197 5314
rect 4232 5304 4440 5314
rect 4475 5310 4520 5314
rect 4523 5313 4524 5314
rect 4539 5313 4552 5314
rect 4258 5274 4447 5304
rect 4273 5271 4447 5274
rect 4266 5268 4447 5271
rect 4075 5248 4088 5250
rect 4103 5248 4137 5250
rect 4075 5232 4149 5248
rect 4176 5244 4189 5258
rect 4204 5244 4220 5260
rect 4266 5255 4277 5268
rect 4059 5210 4060 5226
rect 4075 5210 4088 5232
rect 4103 5210 4133 5232
rect 4176 5228 4238 5244
rect 4266 5237 4277 5253
rect 4282 5248 4292 5268
rect 4302 5248 4316 5268
rect 4319 5255 4328 5268
rect 4344 5255 4353 5268
rect 4282 5237 4316 5248
rect 4319 5237 4328 5253
rect 4344 5237 4353 5253
rect 4360 5248 4370 5268
rect 4380 5248 4394 5268
rect 4395 5255 4406 5268
rect 4360 5237 4394 5248
rect 4395 5237 4406 5253
rect 4452 5244 4468 5260
rect 4475 5258 4505 5310
rect 4539 5306 4540 5313
rect 4524 5298 4540 5306
rect 4511 5266 4524 5285
rect 4539 5266 4569 5282
rect 4511 5250 4585 5266
rect 4511 5248 4524 5250
rect 4539 5248 4573 5250
rect 4176 5226 4189 5228
rect 4204 5226 4238 5228
rect 4176 5210 4238 5226
rect 4282 5221 4298 5224
rect 4360 5221 4390 5232
rect 4438 5228 4484 5244
rect 4511 5232 4585 5248
rect 4438 5226 4472 5228
rect 4437 5210 4484 5226
rect 4511 5210 4524 5232
rect 4539 5210 4569 5232
rect 4596 5210 4597 5226
rect 4612 5210 4625 5370
rect -7 5202 34 5210
rect -7 5176 8 5202
rect 15 5176 34 5202
rect 98 5198 160 5210
rect 172 5198 247 5210
rect 305 5198 380 5210
rect 392 5198 423 5210
rect 429 5198 464 5210
rect 98 5196 260 5198
rect -7 5168 34 5176
rect 116 5172 129 5196
rect 144 5194 159 5196
rect -1 5158 0 5168
rect 15 5158 28 5168
rect 43 5158 73 5172
rect 116 5158 159 5172
rect 183 5169 190 5176
rect 193 5172 260 5196
rect 292 5196 464 5198
rect 262 5174 290 5178
rect 292 5174 372 5196
rect 393 5194 408 5196
rect 262 5172 372 5174
rect 193 5168 372 5172
rect 166 5158 196 5168
rect 198 5158 351 5168
rect 359 5158 389 5168
rect 393 5158 423 5172
rect 451 5158 464 5196
rect 536 5202 571 5210
rect 536 5176 537 5202
rect 544 5176 571 5202
rect 479 5158 509 5172
rect 536 5168 571 5176
rect 573 5202 614 5210
rect 573 5176 588 5202
rect 595 5176 614 5202
rect 678 5198 740 5210
rect 752 5198 827 5210
rect 885 5198 960 5210
rect 972 5198 1003 5210
rect 1009 5198 1044 5210
rect 678 5196 840 5198
rect 573 5168 614 5176
rect 696 5172 709 5196
rect 724 5194 739 5196
rect 536 5158 537 5168
rect 552 5158 565 5168
rect 579 5158 580 5168
rect 595 5158 608 5168
rect 623 5158 653 5172
rect 696 5158 739 5172
rect 763 5169 770 5176
rect 773 5172 840 5196
rect 872 5196 1044 5198
rect 842 5174 870 5178
rect 872 5174 952 5196
rect 973 5194 988 5196
rect 842 5172 952 5174
rect 773 5168 952 5172
rect 746 5158 776 5168
rect 778 5158 931 5168
rect 939 5158 969 5168
rect 973 5158 1003 5172
rect 1031 5158 1044 5196
rect 1116 5202 1151 5210
rect 1116 5176 1117 5202
rect 1124 5176 1151 5202
rect 1059 5158 1089 5172
rect 1116 5168 1151 5176
rect 1153 5202 1194 5210
rect 1153 5176 1168 5202
rect 1175 5176 1194 5202
rect 1258 5198 1320 5210
rect 1332 5198 1407 5210
rect 1465 5198 1540 5210
rect 1552 5198 1583 5210
rect 1589 5198 1624 5210
rect 1258 5196 1420 5198
rect 1153 5168 1194 5176
rect 1276 5172 1289 5196
rect 1304 5194 1319 5196
rect 1116 5158 1117 5168
rect 1132 5158 1145 5168
rect 1159 5158 1160 5168
rect 1175 5158 1188 5168
rect 1203 5158 1233 5172
rect 1276 5158 1319 5172
rect 1343 5169 1350 5176
rect 1353 5172 1420 5196
rect 1452 5196 1624 5198
rect 1422 5174 1450 5178
rect 1452 5174 1532 5196
rect 1553 5194 1568 5196
rect 1422 5172 1532 5174
rect 1353 5168 1532 5172
rect 1326 5158 1356 5168
rect 1358 5158 1511 5168
rect 1519 5158 1549 5168
rect 1553 5158 1583 5172
rect 1611 5158 1624 5196
rect 1696 5202 1731 5210
rect 1696 5176 1697 5202
rect 1704 5176 1731 5202
rect 1639 5158 1669 5172
rect 1696 5168 1731 5176
rect 1733 5202 1774 5210
rect 1733 5176 1748 5202
rect 1755 5176 1774 5202
rect 1838 5198 1900 5210
rect 1912 5198 1987 5210
rect 2045 5198 2120 5210
rect 2132 5198 2163 5210
rect 2169 5198 2204 5210
rect 1838 5196 2000 5198
rect 1733 5168 1774 5176
rect 1856 5172 1869 5196
rect 1884 5194 1899 5196
rect 1696 5158 1697 5168
rect 1712 5158 1725 5168
rect 1739 5158 1740 5168
rect 1755 5158 1768 5168
rect 1783 5158 1813 5172
rect 1856 5158 1899 5172
rect 1923 5169 1930 5176
rect 1933 5172 2000 5196
rect 2032 5196 2204 5198
rect 2002 5174 2030 5178
rect 2032 5174 2112 5196
rect 2133 5194 2148 5196
rect 2002 5172 2112 5174
rect 1933 5168 2112 5172
rect 1906 5158 1936 5168
rect 1938 5158 2091 5168
rect 2099 5158 2129 5168
rect 2133 5158 2163 5172
rect 2191 5158 2204 5196
rect 2276 5202 2311 5210
rect 2276 5176 2277 5202
rect 2284 5176 2311 5202
rect 2219 5158 2249 5172
rect 2276 5168 2311 5176
rect 2313 5202 2354 5210
rect 2313 5176 2328 5202
rect 2335 5176 2354 5202
rect 2418 5198 2480 5210
rect 2492 5198 2567 5210
rect 2625 5198 2700 5210
rect 2712 5198 2743 5210
rect 2749 5198 2784 5210
rect 2418 5196 2580 5198
rect 2313 5168 2354 5176
rect 2436 5172 2449 5196
rect 2464 5194 2479 5196
rect 2276 5158 2277 5168
rect 2292 5158 2305 5168
rect 2319 5158 2320 5168
rect 2335 5158 2348 5168
rect 2363 5158 2393 5172
rect 2436 5158 2479 5172
rect 2503 5169 2510 5176
rect 2513 5172 2580 5196
rect 2612 5196 2784 5198
rect 2582 5174 2610 5178
rect 2612 5174 2692 5196
rect 2713 5194 2728 5196
rect 2582 5172 2692 5174
rect 2513 5168 2692 5172
rect 2486 5158 2516 5168
rect 2518 5158 2671 5168
rect 2679 5158 2709 5168
rect 2713 5158 2743 5172
rect 2771 5158 2784 5196
rect 2856 5202 2891 5210
rect 2856 5176 2857 5202
rect 2864 5176 2891 5202
rect 2799 5158 2829 5172
rect 2856 5168 2891 5176
rect 2893 5202 2934 5210
rect 2893 5176 2908 5202
rect 2915 5176 2934 5202
rect 2998 5198 3060 5210
rect 3072 5198 3147 5210
rect 3205 5198 3280 5210
rect 3292 5198 3323 5210
rect 3329 5198 3364 5210
rect 2998 5196 3160 5198
rect 2893 5168 2934 5176
rect 3016 5172 3029 5196
rect 3044 5194 3059 5196
rect 2856 5158 2857 5168
rect 2872 5158 2885 5168
rect 2899 5158 2900 5168
rect 2915 5158 2928 5168
rect 2943 5158 2973 5172
rect 3016 5158 3059 5172
rect 3083 5169 3090 5176
rect 3093 5172 3160 5196
rect 3192 5196 3364 5198
rect 3162 5174 3190 5178
rect 3192 5174 3272 5196
rect 3293 5194 3308 5196
rect 3162 5172 3272 5174
rect 3093 5168 3272 5172
rect 3066 5158 3096 5168
rect 3098 5158 3251 5168
rect 3259 5158 3289 5168
rect 3293 5158 3323 5172
rect 3351 5158 3364 5196
rect 3436 5202 3471 5210
rect 3436 5176 3437 5202
rect 3444 5176 3471 5202
rect 3379 5158 3409 5172
rect 3436 5168 3471 5176
rect 3473 5202 3514 5210
rect 3473 5176 3488 5202
rect 3495 5176 3514 5202
rect 3578 5198 3640 5210
rect 3652 5198 3727 5210
rect 3785 5198 3860 5210
rect 3872 5198 3903 5210
rect 3909 5198 3944 5210
rect 3578 5196 3740 5198
rect 3473 5168 3514 5176
rect 3596 5172 3609 5196
rect 3624 5194 3639 5196
rect 3436 5158 3437 5168
rect 3452 5158 3465 5168
rect 3479 5158 3480 5168
rect 3495 5158 3508 5168
rect 3523 5158 3553 5172
rect 3596 5158 3639 5172
rect 3663 5169 3670 5176
rect 3673 5172 3740 5196
rect 3772 5196 3944 5198
rect 3742 5174 3770 5178
rect 3772 5174 3852 5196
rect 3873 5194 3888 5196
rect 3742 5172 3852 5174
rect 3673 5168 3852 5172
rect 3646 5158 3676 5168
rect 3678 5158 3831 5168
rect 3839 5158 3869 5168
rect 3873 5158 3903 5172
rect 3931 5158 3944 5196
rect 4016 5202 4051 5210
rect 4016 5176 4017 5202
rect 4024 5176 4051 5202
rect 3959 5158 3989 5172
rect 4016 5168 4051 5176
rect 4053 5202 4094 5210
rect 4053 5176 4068 5202
rect 4075 5176 4094 5202
rect 4158 5198 4220 5210
rect 4232 5198 4307 5210
rect 4365 5198 4440 5210
rect 4452 5198 4483 5210
rect 4489 5198 4524 5210
rect 4158 5196 4320 5198
rect 4053 5168 4094 5176
rect 4176 5172 4189 5196
rect 4204 5194 4219 5196
rect 4016 5158 4017 5168
rect 4032 5158 4045 5168
rect 4059 5158 4060 5168
rect 4075 5158 4088 5168
rect 4103 5158 4133 5172
rect 4176 5158 4219 5172
rect 4243 5169 4250 5176
rect 4253 5172 4320 5196
rect 4352 5196 4524 5198
rect 4322 5174 4350 5178
rect 4352 5174 4432 5196
rect 4453 5194 4468 5196
rect 4322 5172 4432 5174
rect 4253 5168 4432 5172
rect 4226 5158 4256 5168
rect 4258 5158 4411 5168
rect 4419 5158 4449 5168
rect 4453 5158 4483 5172
rect 4511 5158 4524 5196
rect 4596 5202 4631 5210
rect 4596 5176 4597 5202
rect 4604 5176 4631 5202
rect 4539 5158 4569 5172
rect 4596 5168 4631 5176
rect 4596 5158 4597 5168
rect 4612 5158 4625 5168
rect -1 5152 4625 5158
rect 0 5144 4625 5152
rect 15 5114 28 5144
rect 43 5126 73 5144
rect 116 5130 130 5144
rect 166 5130 386 5144
rect 117 5128 130 5130
rect 83 5116 98 5128
rect 80 5114 102 5116
rect 107 5114 137 5128
rect 198 5126 351 5130
rect 180 5114 372 5126
rect 415 5114 445 5128
rect 451 5114 464 5144
rect 479 5126 509 5144
rect 552 5114 565 5144
rect 595 5114 608 5144
rect 623 5126 653 5144
rect 696 5130 710 5144
rect 746 5130 966 5144
rect 697 5128 710 5130
rect 663 5116 678 5128
rect 660 5114 682 5116
rect 687 5114 717 5128
rect 778 5126 931 5130
rect 760 5114 952 5126
rect 995 5114 1025 5128
rect 1031 5114 1044 5144
rect 1059 5126 1089 5144
rect 1132 5114 1145 5144
rect 1175 5114 1188 5144
rect 1203 5126 1233 5144
rect 1276 5130 1290 5144
rect 1326 5130 1546 5144
rect 1277 5128 1290 5130
rect 1243 5116 1258 5128
rect 1240 5114 1262 5116
rect 1267 5114 1297 5128
rect 1358 5126 1511 5130
rect 1340 5114 1532 5126
rect 1575 5114 1605 5128
rect 1611 5114 1624 5144
rect 1639 5126 1669 5144
rect 1712 5114 1725 5144
rect 1755 5114 1768 5144
rect 1783 5126 1813 5144
rect 1856 5130 1870 5144
rect 1906 5130 2126 5144
rect 1857 5128 1870 5130
rect 1823 5116 1838 5128
rect 1820 5114 1842 5116
rect 1847 5114 1877 5128
rect 1938 5126 2091 5130
rect 1920 5114 2112 5126
rect 2155 5114 2185 5128
rect 2191 5114 2204 5144
rect 2219 5126 2249 5144
rect 2292 5114 2305 5144
rect 2335 5114 2348 5144
rect 2363 5126 2393 5144
rect 2436 5130 2450 5144
rect 2486 5130 2706 5144
rect 2437 5128 2450 5130
rect 2403 5116 2418 5128
rect 2400 5114 2422 5116
rect 2427 5114 2457 5128
rect 2518 5126 2671 5130
rect 2500 5114 2692 5126
rect 2735 5114 2765 5128
rect 2771 5114 2784 5144
rect 2799 5126 2829 5144
rect 2872 5114 2885 5144
rect 2915 5114 2928 5144
rect 2943 5126 2973 5144
rect 3016 5130 3030 5144
rect 3066 5130 3286 5144
rect 3017 5128 3030 5130
rect 2983 5116 2998 5128
rect 2980 5114 3002 5116
rect 3007 5114 3037 5128
rect 3098 5126 3251 5130
rect 3080 5114 3272 5126
rect 3315 5114 3345 5128
rect 3351 5114 3364 5144
rect 3379 5126 3409 5144
rect 3452 5114 3465 5144
rect 3495 5114 3508 5144
rect 3523 5126 3553 5144
rect 3596 5130 3610 5144
rect 3646 5130 3866 5144
rect 3597 5128 3610 5130
rect 3563 5116 3578 5128
rect 3560 5114 3582 5116
rect 3587 5114 3617 5128
rect 3678 5126 3831 5130
rect 3660 5114 3852 5126
rect 3895 5114 3925 5128
rect 3931 5114 3944 5144
rect 3959 5126 3989 5144
rect 4032 5114 4045 5144
rect 4075 5114 4088 5144
rect 4103 5126 4133 5144
rect 4176 5130 4190 5144
rect 4226 5130 4446 5144
rect 4177 5128 4190 5130
rect 4143 5116 4158 5128
rect 4140 5114 4162 5116
rect 4167 5114 4197 5128
rect 4258 5126 4411 5130
rect 4240 5114 4432 5126
rect 4475 5114 4505 5128
rect 4511 5114 4524 5144
rect 4539 5126 4569 5144
rect 4612 5114 4625 5144
rect 0 5100 4625 5114
rect 15 4996 28 5100
rect 73 5078 74 5088
rect 89 5078 102 5088
rect 73 5074 102 5078
rect 107 5074 137 5100
rect 155 5086 171 5088
rect 243 5086 296 5100
rect 244 5084 308 5086
rect 351 5084 366 5100
rect 415 5097 445 5100
rect 415 5094 451 5097
rect 381 5086 397 5088
rect 155 5074 170 5078
rect 73 5072 170 5074
rect 198 5072 366 5084
rect 382 5074 397 5078
rect 415 5075 454 5094
rect 473 5088 480 5089
rect 479 5081 480 5088
rect 463 5078 464 5081
rect 479 5078 492 5081
rect 415 5074 445 5075
rect 454 5074 460 5075
rect 463 5074 492 5078
rect 382 5073 492 5074
rect 382 5072 498 5073
rect 57 5064 108 5072
rect 57 5052 82 5064
rect 89 5052 108 5064
rect 139 5064 189 5072
rect 139 5056 155 5064
rect 162 5062 189 5064
rect 198 5062 419 5072
rect 162 5052 419 5062
rect 448 5064 498 5072
rect 448 5055 464 5064
rect 57 5044 108 5052
rect 155 5044 419 5052
rect 445 5052 464 5055
rect 471 5052 498 5064
rect 445 5044 498 5052
rect 73 5036 74 5044
rect 89 5036 102 5044
rect 73 5028 89 5036
rect 70 5021 89 5024
rect 70 5012 92 5021
rect 43 5002 92 5012
rect 43 4996 73 5002
rect 92 4997 97 5002
rect 15 4980 89 4996
rect 107 4988 137 5044
rect 172 5034 380 5044
rect 415 5040 460 5044
rect 463 5043 464 5044
rect 479 5043 492 5044
rect 198 5004 387 5034
rect 213 5001 387 5004
rect 206 4998 387 5001
rect 15 4978 28 4980
rect 43 4978 77 4980
rect 15 4962 89 4978
rect 116 4974 129 4988
rect 144 4974 160 4990
rect 206 4985 217 4998
rect -1 4940 0 4956
rect 15 4940 28 4962
rect 43 4940 73 4962
rect 116 4958 178 4974
rect 206 4967 217 4983
rect 222 4978 232 4998
rect 242 4978 256 4998
rect 259 4985 268 4998
rect 284 4985 293 4998
rect 222 4967 256 4978
rect 259 4967 268 4983
rect 284 4967 293 4983
rect 300 4978 310 4998
rect 320 4978 334 4998
rect 335 4985 346 4998
rect 300 4967 334 4978
rect 335 4967 346 4983
rect 392 4974 408 4990
rect 415 4988 445 5040
rect 479 5036 480 5043
rect 464 5028 480 5036
rect 451 4996 464 5015
rect 479 4996 509 5012
rect 451 4980 525 4996
rect 451 4978 464 4980
rect 479 4978 513 4980
rect 116 4956 129 4958
rect 144 4956 178 4958
rect 116 4940 178 4956
rect 222 4951 238 4954
rect 300 4951 330 4962
rect 378 4958 424 4974
rect 451 4962 525 4978
rect 378 4956 412 4958
rect 377 4940 424 4956
rect 451 4940 464 4962
rect 479 4940 509 4962
rect 536 4940 537 4956
rect 552 4940 565 5100
rect 595 4996 608 5100
rect 653 5078 654 5088
rect 669 5078 682 5088
rect 653 5074 682 5078
rect 687 5074 717 5100
rect 735 5086 751 5088
rect 823 5086 876 5100
rect 824 5084 888 5086
rect 931 5084 946 5100
rect 995 5097 1025 5100
rect 995 5094 1031 5097
rect 961 5086 977 5088
rect 735 5074 750 5078
rect 653 5072 750 5074
rect 778 5072 946 5084
rect 962 5074 977 5078
rect 995 5075 1034 5094
rect 1053 5088 1060 5089
rect 1059 5081 1060 5088
rect 1043 5078 1044 5081
rect 1059 5078 1072 5081
rect 995 5074 1025 5075
rect 1034 5074 1040 5075
rect 1043 5074 1072 5078
rect 962 5073 1072 5074
rect 962 5072 1078 5073
rect 637 5064 688 5072
rect 637 5052 662 5064
rect 669 5052 688 5064
rect 719 5064 769 5072
rect 719 5056 735 5064
rect 742 5062 769 5064
rect 778 5062 999 5072
rect 742 5052 999 5062
rect 1028 5064 1078 5072
rect 1028 5055 1044 5064
rect 637 5044 688 5052
rect 735 5044 999 5052
rect 1025 5052 1044 5055
rect 1051 5052 1078 5064
rect 1025 5044 1078 5052
rect 653 5036 654 5044
rect 669 5036 682 5044
rect 653 5028 669 5036
rect 650 5021 669 5024
rect 650 5012 672 5021
rect 623 5002 672 5012
rect 623 4996 653 5002
rect 672 4997 677 5002
rect 595 4980 669 4996
rect 687 4988 717 5044
rect 752 5034 960 5044
rect 995 5040 1040 5044
rect 1043 5043 1044 5044
rect 1059 5043 1072 5044
rect 778 5004 967 5034
rect 793 5001 967 5004
rect 786 4998 967 5001
rect 595 4978 608 4980
rect 623 4978 657 4980
rect 595 4962 669 4978
rect 696 4974 709 4988
rect 724 4974 740 4990
rect 786 4985 797 4998
rect 579 4940 580 4956
rect 595 4940 608 4962
rect 623 4940 653 4962
rect 696 4958 758 4974
rect 786 4967 797 4983
rect 802 4978 812 4998
rect 822 4978 836 4998
rect 839 4985 848 4998
rect 864 4985 873 4998
rect 802 4967 836 4978
rect 839 4967 848 4983
rect 864 4967 873 4983
rect 880 4978 890 4998
rect 900 4978 914 4998
rect 915 4985 926 4998
rect 880 4967 914 4978
rect 915 4967 926 4983
rect 972 4974 988 4990
rect 995 4988 1025 5040
rect 1059 5036 1060 5043
rect 1044 5028 1060 5036
rect 1031 4996 1044 5015
rect 1059 4996 1089 5012
rect 1031 4980 1105 4996
rect 1031 4978 1044 4980
rect 1059 4978 1093 4980
rect 696 4956 709 4958
rect 724 4956 758 4958
rect 696 4940 758 4956
rect 802 4951 818 4954
rect 880 4951 910 4962
rect 958 4958 1004 4974
rect 1031 4962 1105 4978
rect 958 4956 992 4958
rect 957 4940 1004 4956
rect 1031 4940 1044 4962
rect 1059 4940 1089 4962
rect 1116 4940 1117 4956
rect 1132 4940 1145 5100
rect 1175 4996 1188 5100
rect 1233 5078 1234 5088
rect 1249 5078 1262 5088
rect 1233 5074 1262 5078
rect 1267 5074 1297 5100
rect 1315 5086 1331 5088
rect 1403 5086 1456 5100
rect 1404 5084 1468 5086
rect 1511 5084 1526 5100
rect 1575 5097 1605 5100
rect 1575 5094 1611 5097
rect 1541 5086 1557 5088
rect 1315 5074 1330 5078
rect 1233 5072 1330 5074
rect 1358 5072 1526 5084
rect 1542 5074 1557 5078
rect 1575 5075 1614 5094
rect 1633 5088 1640 5089
rect 1639 5081 1640 5088
rect 1623 5078 1624 5081
rect 1639 5078 1652 5081
rect 1575 5074 1605 5075
rect 1614 5074 1620 5075
rect 1623 5074 1652 5078
rect 1542 5073 1652 5074
rect 1542 5072 1658 5073
rect 1217 5064 1268 5072
rect 1217 5052 1242 5064
rect 1249 5052 1268 5064
rect 1299 5064 1349 5072
rect 1299 5056 1315 5064
rect 1322 5062 1349 5064
rect 1358 5062 1579 5072
rect 1322 5052 1579 5062
rect 1608 5064 1658 5072
rect 1608 5055 1624 5064
rect 1217 5044 1268 5052
rect 1315 5044 1579 5052
rect 1605 5052 1624 5055
rect 1631 5052 1658 5064
rect 1605 5044 1658 5052
rect 1233 5036 1234 5044
rect 1249 5036 1262 5044
rect 1233 5028 1249 5036
rect 1230 5021 1249 5024
rect 1230 5012 1252 5021
rect 1203 5002 1252 5012
rect 1203 4996 1233 5002
rect 1252 4997 1257 5002
rect 1175 4980 1249 4996
rect 1267 4988 1297 5044
rect 1332 5034 1540 5044
rect 1575 5040 1620 5044
rect 1623 5043 1624 5044
rect 1639 5043 1652 5044
rect 1358 5004 1547 5034
rect 1373 5001 1547 5004
rect 1366 4998 1547 5001
rect 1175 4978 1188 4980
rect 1203 4978 1237 4980
rect 1175 4962 1249 4978
rect 1276 4974 1289 4988
rect 1304 4974 1320 4990
rect 1366 4985 1377 4998
rect 1159 4940 1160 4956
rect 1175 4940 1188 4962
rect 1203 4940 1233 4962
rect 1276 4958 1338 4974
rect 1366 4967 1377 4983
rect 1382 4978 1392 4998
rect 1402 4978 1416 4998
rect 1419 4985 1428 4998
rect 1444 4985 1453 4998
rect 1382 4967 1416 4978
rect 1419 4967 1428 4983
rect 1444 4967 1453 4983
rect 1460 4978 1470 4998
rect 1480 4978 1494 4998
rect 1495 4985 1506 4998
rect 1460 4967 1494 4978
rect 1495 4967 1506 4983
rect 1552 4974 1568 4990
rect 1575 4988 1605 5040
rect 1639 5036 1640 5043
rect 1624 5028 1640 5036
rect 1611 4996 1624 5015
rect 1639 4996 1669 5012
rect 1611 4980 1685 4996
rect 1611 4978 1624 4980
rect 1639 4978 1673 4980
rect 1276 4956 1289 4958
rect 1304 4956 1338 4958
rect 1276 4940 1338 4956
rect 1382 4951 1398 4954
rect 1460 4951 1490 4962
rect 1538 4958 1584 4974
rect 1611 4962 1685 4978
rect 1538 4956 1572 4958
rect 1537 4940 1584 4956
rect 1611 4940 1624 4962
rect 1639 4940 1669 4962
rect 1696 4940 1697 4956
rect 1712 4940 1725 5100
rect 1755 4996 1768 5100
rect 1813 5078 1814 5088
rect 1829 5078 1842 5088
rect 1813 5074 1842 5078
rect 1847 5074 1877 5100
rect 1895 5086 1911 5088
rect 1983 5086 2036 5100
rect 1984 5084 2048 5086
rect 2091 5084 2106 5100
rect 2155 5097 2185 5100
rect 2155 5094 2191 5097
rect 2121 5086 2137 5088
rect 1895 5074 1910 5078
rect 1813 5072 1910 5074
rect 1938 5072 2106 5084
rect 2122 5074 2137 5078
rect 2155 5075 2194 5094
rect 2213 5088 2220 5089
rect 2219 5081 2220 5088
rect 2203 5078 2204 5081
rect 2219 5078 2232 5081
rect 2155 5074 2185 5075
rect 2194 5074 2200 5075
rect 2203 5074 2232 5078
rect 2122 5073 2232 5074
rect 2122 5072 2238 5073
rect 1797 5064 1848 5072
rect 1797 5052 1822 5064
rect 1829 5052 1848 5064
rect 1879 5064 1929 5072
rect 1879 5056 1895 5064
rect 1902 5062 1929 5064
rect 1938 5062 2159 5072
rect 1902 5052 2159 5062
rect 2188 5064 2238 5072
rect 2188 5055 2204 5064
rect 1797 5044 1848 5052
rect 1895 5044 2159 5052
rect 2185 5052 2204 5055
rect 2211 5052 2238 5064
rect 2185 5044 2238 5052
rect 1813 5036 1814 5044
rect 1829 5036 1842 5044
rect 1813 5028 1829 5036
rect 1810 5021 1829 5024
rect 1810 5012 1832 5021
rect 1783 5002 1832 5012
rect 1783 4996 1813 5002
rect 1832 4997 1837 5002
rect 1755 4980 1829 4996
rect 1847 4988 1877 5044
rect 1912 5034 2120 5044
rect 2155 5040 2200 5044
rect 2203 5043 2204 5044
rect 2219 5043 2232 5044
rect 1938 5004 2127 5034
rect 1953 5001 2127 5004
rect 1946 4998 2127 5001
rect 1755 4978 1768 4980
rect 1783 4978 1817 4980
rect 1755 4962 1829 4978
rect 1856 4974 1869 4988
rect 1884 4974 1900 4990
rect 1946 4985 1957 4998
rect 1739 4940 1740 4956
rect 1755 4940 1768 4962
rect 1783 4940 1813 4962
rect 1856 4958 1918 4974
rect 1946 4967 1957 4983
rect 1962 4978 1972 4998
rect 1982 4978 1996 4998
rect 1999 4985 2008 4998
rect 2024 4985 2033 4998
rect 1962 4967 1996 4978
rect 1999 4967 2008 4983
rect 2024 4967 2033 4983
rect 2040 4978 2050 4998
rect 2060 4978 2074 4998
rect 2075 4985 2086 4998
rect 2040 4967 2074 4978
rect 2075 4967 2086 4983
rect 2132 4974 2148 4990
rect 2155 4988 2185 5040
rect 2219 5036 2220 5043
rect 2204 5028 2220 5036
rect 2191 4996 2204 5015
rect 2219 4996 2249 5012
rect 2191 4980 2265 4996
rect 2191 4978 2204 4980
rect 2219 4978 2253 4980
rect 1856 4956 1869 4958
rect 1884 4956 1918 4958
rect 1856 4940 1918 4956
rect 1962 4951 1978 4954
rect 2040 4951 2070 4962
rect 2118 4958 2164 4974
rect 2191 4962 2265 4978
rect 2118 4956 2152 4958
rect 2117 4940 2164 4956
rect 2191 4940 2204 4962
rect 2219 4940 2249 4962
rect 2276 4940 2277 4956
rect 2292 4940 2305 5100
rect 2335 4996 2348 5100
rect 2393 5078 2394 5088
rect 2409 5078 2422 5088
rect 2393 5074 2422 5078
rect 2427 5074 2457 5100
rect 2475 5086 2491 5088
rect 2563 5086 2616 5100
rect 2564 5084 2628 5086
rect 2671 5084 2686 5100
rect 2735 5097 2765 5100
rect 2735 5094 2771 5097
rect 2701 5086 2717 5088
rect 2475 5074 2490 5078
rect 2393 5072 2490 5074
rect 2518 5072 2686 5084
rect 2702 5074 2717 5078
rect 2735 5075 2774 5094
rect 2793 5088 2800 5089
rect 2799 5081 2800 5088
rect 2783 5078 2784 5081
rect 2799 5078 2812 5081
rect 2735 5074 2765 5075
rect 2774 5074 2780 5075
rect 2783 5074 2812 5078
rect 2702 5073 2812 5074
rect 2702 5072 2818 5073
rect 2377 5064 2428 5072
rect 2377 5052 2402 5064
rect 2409 5052 2428 5064
rect 2459 5064 2509 5072
rect 2459 5056 2475 5064
rect 2482 5062 2509 5064
rect 2518 5062 2739 5072
rect 2482 5052 2739 5062
rect 2768 5064 2818 5072
rect 2768 5055 2784 5064
rect 2377 5044 2428 5052
rect 2475 5044 2739 5052
rect 2765 5052 2784 5055
rect 2791 5052 2818 5064
rect 2765 5044 2818 5052
rect 2393 5036 2394 5044
rect 2409 5036 2422 5044
rect 2393 5028 2409 5036
rect 2390 5021 2409 5024
rect 2390 5012 2412 5021
rect 2363 5002 2412 5012
rect 2363 4996 2393 5002
rect 2412 4997 2417 5002
rect 2335 4980 2409 4996
rect 2427 4988 2457 5044
rect 2492 5034 2700 5044
rect 2735 5040 2780 5044
rect 2783 5043 2784 5044
rect 2799 5043 2812 5044
rect 2518 5004 2707 5034
rect 2533 5001 2707 5004
rect 2526 4998 2707 5001
rect 2335 4978 2348 4980
rect 2363 4978 2397 4980
rect 2335 4962 2409 4978
rect 2436 4974 2449 4988
rect 2464 4974 2480 4990
rect 2526 4985 2537 4998
rect 2319 4940 2320 4956
rect 2335 4940 2348 4962
rect 2363 4940 2393 4962
rect 2436 4958 2498 4974
rect 2526 4967 2537 4983
rect 2542 4978 2552 4998
rect 2562 4978 2576 4998
rect 2579 4985 2588 4998
rect 2604 4985 2613 4998
rect 2542 4967 2576 4978
rect 2579 4967 2588 4983
rect 2604 4967 2613 4983
rect 2620 4978 2630 4998
rect 2640 4978 2654 4998
rect 2655 4985 2666 4998
rect 2620 4967 2654 4978
rect 2655 4967 2666 4983
rect 2712 4974 2728 4990
rect 2735 4988 2765 5040
rect 2799 5036 2800 5043
rect 2784 5028 2800 5036
rect 2771 4996 2784 5015
rect 2799 4996 2829 5012
rect 2771 4980 2845 4996
rect 2771 4978 2784 4980
rect 2799 4978 2833 4980
rect 2436 4956 2449 4958
rect 2464 4956 2498 4958
rect 2436 4940 2498 4956
rect 2542 4951 2558 4954
rect 2620 4951 2650 4962
rect 2698 4958 2744 4974
rect 2771 4962 2845 4978
rect 2698 4956 2732 4958
rect 2697 4940 2744 4956
rect 2771 4940 2784 4962
rect 2799 4940 2829 4962
rect 2856 4940 2857 4956
rect 2872 4940 2885 5100
rect 2915 4996 2928 5100
rect 2973 5078 2974 5088
rect 2989 5078 3002 5088
rect 2973 5074 3002 5078
rect 3007 5074 3037 5100
rect 3055 5086 3071 5088
rect 3143 5086 3196 5100
rect 3144 5084 3208 5086
rect 3251 5084 3266 5100
rect 3315 5097 3345 5100
rect 3315 5094 3351 5097
rect 3281 5086 3297 5088
rect 3055 5074 3070 5078
rect 2973 5072 3070 5074
rect 3098 5072 3266 5084
rect 3282 5074 3297 5078
rect 3315 5075 3354 5094
rect 3373 5088 3380 5089
rect 3379 5081 3380 5088
rect 3363 5078 3364 5081
rect 3379 5078 3392 5081
rect 3315 5074 3345 5075
rect 3354 5074 3360 5075
rect 3363 5074 3392 5078
rect 3282 5073 3392 5074
rect 3282 5072 3398 5073
rect 2957 5064 3008 5072
rect 2957 5052 2982 5064
rect 2989 5052 3008 5064
rect 3039 5064 3089 5072
rect 3039 5056 3055 5064
rect 3062 5062 3089 5064
rect 3098 5062 3319 5072
rect 3062 5052 3319 5062
rect 3348 5064 3398 5072
rect 3348 5055 3364 5064
rect 2957 5044 3008 5052
rect 3055 5044 3319 5052
rect 3345 5052 3364 5055
rect 3371 5052 3398 5064
rect 3345 5044 3398 5052
rect 2973 5036 2974 5044
rect 2989 5036 3002 5044
rect 2973 5028 2989 5036
rect 2970 5021 2989 5024
rect 2970 5012 2992 5021
rect 2943 5002 2992 5012
rect 2943 4996 2973 5002
rect 2992 4997 2997 5002
rect 2915 4980 2989 4996
rect 3007 4988 3037 5044
rect 3072 5034 3280 5044
rect 3315 5040 3360 5044
rect 3363 5043 3364 5044
rect 3379 5043 3392 5044
rect 3098 5004 3287 5034
rect 3113 5001 3287 5004
rect 3106 4998 3287 5001
rect 2915 4978 2928 4980
rect 2943 4978 2977 4980
rect 2915 4962 2989 4978
rect 3016 4974 3029 4988
rect 3044 4974 3060 4990
rect 3106 4985 3117 4998
rect 2899 4940 2900 4956
rect 2915 4940 2928 4962
rect 2943 4940 2973 4962
rect 3016 4958 3078 4974
rect 3106 4967 3117 4983
rect 3122 4978 3132 4998
rect 3142 4978 3156 4998
rect 3159 4985 3168 4998
rect 3184 4985 3193 4998
rect 3122 4967 3156 4978
rect 3159 4967 3168 4983
rect 3184 4967 3193 4983
rect 3200 4978 3210 4998
rect 3220 4978 3234 4998
rect 3235 4985 3246 4998
rect 3200 4967 3234 4978
rect 3235 4967 3246 4983
rect 3292 4974 3308 4990
rect 3315 4988 3345 5040
rect 3379 5036 3380 5043
rect 3364 5028 3380 5036
rect 3351 4996 3364 5015
rect 3379 4996 3409 5012
rect 3351 4980 3425 4996
rect 3351 4978 3364 4980
rect 3379 4978 3413 4980
rect 3016 4956 3029 4958
rect 3044 4956 3078 4958
rect 3016 4940 3078 4956
rect 3122 4951 3138 4954
rect 3200 4951 3230 4962
rect 3278 4958 3324 4974
rect 3351 4962 3425 4978
rect 3278 4956 3312 4958
rect 3277 4940 3324 4956
rect 3351 4940 3364 4962
rect 3379 4940 3409 4962
rect 3436 4940 3437 4956
rect 3452 4940 3465 5100
rect 3495 4996 3508 5100
rect 3553 5078 3554 5088
rect 3569 5078 3582 5088
rect 3553 5074 3582 5078
rect 3587 5074 3617 5100
rect 3635 5086 3651 5088
rect 3723 5086 3776 5100
rect 3724 5084 3788 5086
rect 3831 5084 3846 5100
rect 3895 5097 3925 5100
rect 3895 5094 3931 5097
rect 3861 5086 3877 5088
rect 3635 5074 3650 5078
rect 3553 5072 3650 5074
rect 3678 5072 3846 5084
rect 3862 5074 3877 5078
rect 3895 5075 3934 5094
rect 3953 5088 3960 5089
rect 3959 5081 3960 5088
rect 3943 5078 3944 5081
rect 3959 5078 3972 5081
rect 3895 5074 3925 5075
rect 3934 5074 3940 5075
rect 3943 5074 3972 5078
rect 3862 5073 3972 5074
rect 3862 5072 3978 5073
rect 3537 5064 3588 5072
rect 3537 5052 3562 5064
rect 3569 5052 3588 5064
rect 3619 5064 3669 5072
rect 3619 5056 3635 5064
rect 3642 5062 3669 5064
rect 3678 5062 3899 5072
rect 3642 5052 3899 5062
rect 3928 5064 3978 5072
rect 3928 5055 3944 5064
rect 3537 5044 3588 5052
rect 3635 5044 3899 5052
rect 3925 5052 3944 5055
rect 3951 5052 3978 5064
rect 3925 5044 3978 5052
rect 3553 5036 3554 5044
rect 3569 5036 3582 5044
rect 3553 5028 3569 5036
rect 3550 5021 3569 5024
rect 3550 5012 3572 5021
rect 3523 5002 3572 5012
rect 3523 4996 3553 5002
rect 3572 4997 3577 5002
rect 3495 4980 3569 4996
rect 3587 4988 3617 5044
rect 3652 5034 3860 5044
rect 3895 5040 3940 5044
rect 3943 5043 3944 5044
rect 3959 5043 3972 5044
rect 3678 5004 3867 5034
rect 3693 5001 3867 5004
rect 3686 4998 3867 5001
rect 3495 4978 3508 4980
rect 3523 4978 3557 4980
rect 3495 4962 3569 4978
rect 3596 4974 3609 4988
rect 3624 4974 3640 4990
rect 3686 4985 3697 4998
rect 3479 4940 3480 4956
rect 3495 4940 3508 4962
rect 3523 4940 3553 4962
rect 3596 4958 3658 4974
rect 3686 4967 3697 4983
rect 3702 4978 3712 4998
rect 3722 4978 3736 4998
rect 3739 4985 3748 4998
rect 3764 4985 3773 4998
rect 3702 4967 3736 4978
rect 3739 4967 3748 4983
rect 3764 4967 3773 4983
rect 3780 4978 3790 4998
rect 3800 4978 3814 4998
rect 3815 4985 3826 4998
rect 3780 4967 3814 4978
rect 3815 4967 3826 4983
rect 3872 4974 3888 4990
rect 3895 4988 3925 5040
rect 3959 5036 3960 5043
rect 3944 5028 3960 5036
rect 3931 4996 3944 5015
rect 3959 4996 3989 5012
rect 3931 4980 4005 4996
rect 3931 4978 3944 4980
rect 3959 4978 3993 4980
rect 3596 4956 3609 4958
rect 3624 4956 3658 4958
rect 3596 4940 3658 4956
rect 3702 4951 3718 4954
rect 3780 4951 3810 4962
rect 3858 4958 3904 4974
rect 3931 4962 4005 4978
rect 3858 4956 3892 4958
rect 3857 4940 3904 4956
rect 3931 4940 3944 4962
rect 3959 4940 3989 4962
rect 4016 4940 4017 4956
rect 4032 4940 4045 5100
rect 4075 4996 4088 5100
rect 4133 5078 4134 5088
rect 4149 5078 4162 5088
rect 4133 5074 4162 5078
rect 4167 5074 4197 5100
rect 4215 5086 4231 5088
rect 4303 5086 4356 5100
rect 4304 5084 4368 5086
rect 4411 5084 4426 5100
rect 4475 5097 4505 5100
rect 4475 5094 4511 5097
rect 4441 5086 4457 5088
rect 4215 5074 4230 5078
rect 4133 5072 4230 5074
rect 4258 5072 4426 5084
rect 4442 5074 4457 5078
rect 4475 5075 4514 5094
rect 4533 5088 4540 5089
rect 4539 5081 4540 5088
rect 4523 5078 4524 5081
rect 4539 5078 4552 5081
rect 4475 5074 4505 5075
rect 4514 5074 4520 5075
rect 4523 5074 4552 5078
rect 4442 5073 4552 5074
rect 4442 5072 4558 5073
rect 4117 5064 4168 5072
rect 4117 5052 4142 5064
rect 4149 5052 4168 5064
rect 4199 5064 4249 5072
rect 4199 5056 4215 5064
rect 4222 5062 4249 5064
rect 4258 5062 4479 5072
rect 4222 5052 4479 5062
rect 4508 5064 4558 5072
rect 4508 5055 4524 5064
rect 4117 5044 4168 5052
rect 4215 5044 4479 5052
rect 4505 5052 4524 5055
rect 4531 5052 4558 5064
rect 4505 5044 4558 5052
rect 4133 5036 4134 5044
rect 4149 5036 4162 5044
rect 4133 5028 4149 5036
rect 4130 5021 4149 5024
rect 4130 5012 4152 5021
rect 4103 5002 4152 5012
rect 4103 4996 4133 5002
rect 4152 4997 4157 5002
rect 4075 4980 4149 4996
rect 4167 4988 4197 5044
rect 4232 5034 4440 5044
rect 4475 5040 4520 5044
rect 4523 5043 4524 5044
rect 4539 5043 4552 5044
rect 4258 5004 4447 5034
rect 4273 5001 4447 5004
rect 4266 4998 4447 5001
rect 4075 4978 4088 4980
rect 4103 4978 4137 4980
rect 4075 4962 4149 4978
rect 4176 4974 4189 4988
rect 4204 4974 4220 4990
rect 4266 4985 4277 4998
rect 4059 4940 4060 4956
rect 4075 4940 4088 4962
rect 4103 4940 4133 4962
rect 4176 4958 4238 4974
rect 4266 4967 4277 4983
rect 4282 4978 4292 4998
rect 4302 4978 4316 4998
rect 4319 4985 4328 4998
rect 4344 4985 4353 4998
rect 4282 4967 4316 4978
rect 4319 4967 4328 4983
rect 4344 4967 4353 4983
rect 4360 4978 4370 4998
rect 4380 4978 4394 4998
rect 4395 4985 4406 4998
rect 4360 4967 4394 4978
rect 4395 4967 4406 4983
rect 4452 4974 4468 4990
rect 4475 4988 4505 5040
rect 4539 5036 4540 5043
rect 4524 5028 4540 5036
rect 4511 4996 4524 5015
rect 4539 4996 4569 5012
rect 4511 4980 4585 4996
rect 4511 4978 4524 4980
rect 4539 4978 4573 4980
rect 4176 4956 4189 4958
rect 4204 4956 4238 4958
rect 4176 4940 4238 4956
rect 4282 4951 4298 4954
rect 4360 4951 4390 4962
rect 4438 4958 4484 4974
rect 4511 4962 4585 4978
rect 4438 4956 4472 4958
rect 4437 4940 4484 4956
rect 4511 4940 4524 4962
rect 4539 4940 4569 4962
rect 4596 4940 4597 4956
rect 4612 4940 4625 5100
rect -7 4932 34 4940
rect -7 4906 8 4932
rect 15 4906 34 4932
rect 98 4928 160 4940
rect 172 4928 247 4940
rect 305 4928 380 4940
rect 392 4928 423 4940
rect 429 4928 464 4940
rect 98 4926 260 4928
rect -7 4898 34 4906
rect 116 4902 129 4926
rect 144 4924 159 4926
rect -1 4888 0 4898
rect 15 4888 28 4898
rect 43 4888 73 4902
rect 116 4888 159 4902
rect 183 4899 190 4906
rect 193 4902 260 4926
rect 292 4926 464 4928
rect 262 4904 290 4908
rect 292 4904 372 4926
rect 393 4924 408 4926
rect 262 4902 372 4904
rect 193 4898 372 4902
rect 166 4888 196 4898
rect 198 4888 351 4898
rect 359 4888 389 4898
rect 393 4888 423 4902
rect 451 4888 464 4926
rect 536 4932 571 4940
rect 536 4906 537 4932
rect 544 4906 571 4932
rect 479 4888 509 4902
rect 536 4898 571 4906
rect 573 4932 614 4940
rect 573 4906 588 4932
rect 595 4906 614 4932
rect 678 4928 740 4940
rect 752 4928 827 4940
rect 885 4928 960 4940
rect 972 4928 1003 4940
rect 1009 4928 1044 4940
rect 678 4926 840 4928
rect 573 4898 614 4906
rect 696 4902 709 4926
rect 724 4924 739 4926
rect 536 4888 537 4898
rect 552 4888 565 4898
rect 579 4888 580 4898
rect 595 4888 608 4898
rect 623 4888 653 4902
rect 696 4888 739 4902
rect 763 4899 770 4906
rect 773 4902 840 4926
rect 872 4926 1044 4928
rect 842 4904 870 4908
rect 872 4904 952 4926
rect 973 4924 988 4926
rect 842 4902 952 4904
rect 773 4898 952 4902
rect 746 4888 776 4898
rect 778 4888 931 4898
rect 939 4888 969 4898
rect 973 4888 1003 4902
rect 1031 4888 1044 4926
rect 1116 4932 1151 4940
rect 1116 4906 1117 4932
rect 1124 4906 1151 4932
rect 1059 4888 1089 4902
rect 1116 4898 1151 4906
rect 1153 4932 1194 4940
rect 1153 4906 1168 4932
rect 1175 4906 1194 4932
rect 1258 4928 1320 4940
rect 1332 4928 1407 4940
rect 1465 4928 1540 4940
rect 1552 4928 1583 4940
rect 1589 4928 1624 4940
rect 1258 4926 1420 4928
rect 1153 4898 1194 4906
rect 1276 4902 1289 4926
rect 1304 4924 1319 4926
rect 1116 4888 1117 4898
rect 1132 4888 1145 4898
rect 1159 4888 1160 4898
rect 1175 4888 1188 4898
rect 1203 4888 1233 4902
rect 1276 4888 1319 4902
rect 1343 4899 1350 4906
rect 1353 4902 1420 4926
rect 1452 4926 1624 4928
rect 1422 4904 1450 4908
rect 1452 4904 1532 4926
rect 1553 4924 1568 4926
rect 1422 4902 1532 4904
rect 1353 4898 1532 4902
rect 1326 4888 1356 4898
rect 1358 4888 1511 4898
rect 1519 4888 1549 4898
rect 1553 4888 1583 4902
rect 1611 4888 1624 4926
rect 1696 4932 1731 4940
rect 1696 4906 1697 4932
rect 1704 4906 1731 4932
rect 1639 4888 1669 4902
rect 1696 4898 1731 4906
rect 1733 4932 1774 4940
rect 1733 4906 1748 4932
rect 1755 4906 1774 4932
rect 1838 4928 1900 4940
rect 1912 4928 1987 4940
rect 2045 4928 2120 4940
rect 2132 4928 2163 4940
rect 2169 4928 2204 4940
rect 1838 4926 2000 4928
rect 1733 4898 1774 4906
rect 1856 4902 1869 4926
rect 1884 4924 1899 4926
rect 1696 4888 1697 4898
rect 1712 4888 1725 4898
rect 1739 4888 1740 4898
rect 1755 4888 1768 4898
rect 1783 4888 1813 4902
rect 1856 4888 1899 4902
rect 1923 4899 1930 4906
rect 1933 4902 2000 4926
rect 2032 4926 2204 4928
rect 2002 4904 2030 4908
rect 2032 4904 2112 4926
rect 2133 4924 2148 4926
rect 2002 4902 2112 4904
rect 1933 4898 2112 4902
rect 1906 4888 1936 4898
rect 1938 4888 2091 4898
rect 2099 4888 2129 4898
rect 2133 4888 2163 4902
rect 2191 4888 2204 4926
rect 2276 4932 2311 4940
rect 2276 4906 2277 4932
rect 2284 4906 2311 4932
rect 2219 4888 2249 4902
rect 2276 4898 2311 4906
rect 2313 4932 2354 4940
rect 2313 4906 2328 4932
rect 2335 4906 2354 4932
rect 2418 4928 2480 4940
rect 2492 4928 2567 4940
rect 2625 4928 2700 4940
rect 2712 4928 2743 4940
rect 2749 4928 2784 4940
rect 2418 4926 2580 4928
rect 2313 4898 2354 4906
rect 2436 4902 2449 4926
rect 2464 4924 2479 4926
rect 2276 4888 2277 4898
rect 2292 4888 2305 4898
rect 2319 4888 2320 4898
rect 2335 4888 2348 4898
rect 2363 4888 2393 4902
rect 2436 4888 2479 4902
rect 2503 4899 2510 4906
rect 2513 4902 2580 4926
rect 2612 4926 2784 4928
rect 2582 4904 2610 4908
rect 2612 4904 2692 4926
rect 2713 4924 2728 4926
rect 2582 4902 2692 4904
rect 2513 4898 2692 4902
rect 2486 4888 2516 4898
rect 2518 4888 2671 4898
rect 2679 4888 2709 4898
rect 2713 4888 2743 4902
rect 2771 4888 2784 4926
rect 2856 4932 2891 4940
rect 2856 4906 2857 4932
rect 2864 4906 2891 4932
rect 2799 4888 2829 4902
rect 2856 4898 2891 4906
rect 2893 4932 2934 4940
rect 2893 4906 2908 4932
rect 2915 4906 2934 4932
rect 2998 4928 3060 4940
rect 3072 4928 3147 4940
rect 3205 4928 3280 4940
rect 3292 4928 3323 4940
rect 3329 4928 3364 4940
rect 2998 4926 3160 4928
rect 2893 4898 2934 4906
rect 3016 4902 3029 4926
rect 3044 4924 3059 4926
rect 2856 4888 2857 4898
rect 2872 4888 2885 4898
rect 2899 4888 2900 4898
rect 2915 4888 2928 4898
rect 2943 4888 2973 4902
rect 3016 4888 3059 4902
rect 3083 4899 3090 4906
rect 3093 4902 3160 4926
rect 3192 4926 3364 4928
rect 3162 4904 3190 4908
rect 3192 4904 3272 4926
rect 3293 4924 3308 4926
rect 3162 4902 3272 4904
rect 3093 4898 3272 4902
rect 3066 4888 3096 4898
rect 3098 4888 3251 4898
rect 3259 4888 3289 4898
rect 3293 4888 3323 4902
rect 3351 4888 3364 4926
rect 3436 4932 3471 4940
rect 3436 4906 3437 4932
rect 3444 4906 3471 4932
rect 3379 4888 3409 4902
rect 3436 4898 3471 4906
rect 3473 4932 3514 4940
rect 3473 4906 3488 4932
rect 3495 4906 3514 4932
rect 3578 4928 3640 4940
rect 3652 4928 3727 4940
rect 3785 4928 3860 4940
rect 3872 4928 3903 4940
rect 3909 4928 3944 4940
rect 3578 4926 3740 4928
rect 3473 4898 3514 4906
rect 3596 4902 3609 4926
rect 3624 4924 3639 4926
rect 3436 4888 3437 4898
rect 3452 4888 3465 4898
rect 3479 4888 3480 4898
rect 3495 4888 3508 4898
rect 3523 4888 3553 4902
rect 3596 4888 3639 4902
rect 3663 4899 3670 4906
rect 3673 4902 3740 4926
rect 3772 4926 3944 4928
rect 3742 4904 3770 4908
rect 3772 4904 3852 4926
rect 3873 4924 3888 4926
rect 3742 4902 3852 4904
rect 3673 4898 3852 4902
rect 3646 4888 3676 4898
rect 3678 4888 3831 4898
rect 3839 4888 3869 4898
rect 3873 4888 3903 4902
rect 3931 4888 3944 4926
rect 4016 4932 4051 4940
rect 4016 4906 4017 4932
rect 4024 4906 4051 4932
rect 3959 4888 3989 4902
rect 4016 4898 4051 4906
rect 4053 4932 4094 4940
rect 4053 4906 4068 4932
rect 4075 4906 4094 4932
rect 4158 4928 4220 4940
rect 4232 4928 4307 4940
rect 4365 4928 4440 4940
rect 4452 4928 4483 4940
rect 4489 4928 4524 4940
rect 4158 4926 4320 4928
rect 4053 4898 4094 4906
rect 4176 4902 4189 4926
rect 4204 4924 4219 4926
rect 4016 4888 4017 4898
rect 4032 4888 4045 4898
rect 4059 4888 4060 4898
rect 4075 4888 4088 4898
rect 4103 4888 4133 4902
rect 4176 4888 4219 4902
rect 4243 4899 4250 4906
rect 4253 4902 4320 4926
rect 4352 4926 4524 4928
rect 4322 4904 4350 4908
rect 4352 4904 4432 4926
rect 4453 4924 4468 4926
rect 4322 4902 4432 4904
rect 4253 4898 4432 4902
rect 4226 4888 4256 4898
rect 4258 4888 4411 4898
rect 4419 4888 4449 4898
rect 4453 4888 4483 4902
rect 4511 4888 4524 4926
rect 4596 4932 4631 4940
rect 4596 4906 4597 4932
rect 4604 4906 4631 4932
rect 4539 4888 4569 4902
rect 4596 4898 4631 4906
rect 4596 4888 4597 4898
rect 4612 4888 4625 4898
rect -1 4882 4625 4888
rect 0 4874 4625 4882
rect 15 4844 28 4874
rect 43 4856 73 4874
rect 116 4860 130 4874
rect 166 4860 386 4874
rect 117 4858 130 4860
rect 83 4846 98 4858
rect 80 4844 102 4846
rect 107 4844 137 4858
rect 198 4856 351 4860
rect 180 4844 372 4856
rect 415 4844 445 4858
rect 451 4844 464 4874
rect 479 4856 509 4874
rect 552 4844 565 4874
rect 595 4844 608 4874
rect 623 4856 653 4874
rect 696 4860 710 4874
rect 746 4860 966 4874
rect 697 4858 710 4860
rect 663 4846 678 4858
rect 660 4844 682 4846
rect 687 4844 717 4858
rect 778 4856 931 4860
rect 760 4844 952 4856
rect 995 4844 1025 4858
rect 1031 4844 1044 4874
rect 1059 4856 1089 4874
rect 1132 4844 1145 4874
rect 1175 4844 1188 4874
rect 1203 4856 1233 4874
rect 1276 4860 1290 4874
rect 1326 4860 1546 4874
rect 1277 4858 1290 4860
rect 1243 4846 1258 4858
rect 1240 4844 1262 4846
rect 1267 4844 1297 4858
rect 1358 4856 1511 4860
rect 1340 4844 1532 4856
rect 1575 4844 1605 4858
rect 1611 4844 1624 4874
rect 1639 4856 1669 4874
rect 1712 4844 1725 4874
rect 1755 4844 1768 4874
rect 1783 4856 1813 4874
rect 1856 4860 1870 4874
rect 1906 4860 2126 4874
rect 1857 4858 1870 4860
rect 1823 4846 1838 4858
rect 1820 4844 1842 4846
rect 1847 4844 1877 4858
rect 1938 4856 2091 4860
rect 1920 4844 2112 4856
rect 2155 4844 2185 4858
rect 2191 4844 2204 4874
rect 2219 4856 2249 4874
rect 2292 4844 2305 4874
rect 2335 4844 2348 4874
rect 2363 4856 2393 4874
rect 2436 4860 2450 4874
rect 2486 4860 2706 4874
rect 2437 4858 2450 4860
rect 2403 4846 2418 4858
rect 2400 4844 2422 4846
rect 2427 4844 2457 4858
rect 2518 4856 2671 4860
rect 2500 4844 2692 4856
rect 2735 4844 2765 4858
rect 2771 4844 2784 4874
rect 2799 4856 2829 4874
rect 2872 4844 2885 4874
rect 2915 4844 2928 4874
rect 2943 4856 2973 4874
rect 3016 4860 3030 4874
rect 3066 4860 3286 4874
rect 3017 4858 3030 4860
rect 2983 4846 2998 4858
rect 2980 4844 3002 4846
rect 3007 4844 3037 4858
rect 3098 4856 3251 4860
rect 3080 4844 3272 4856
rect 3315 4844 3345 4858
rect 3351 4844 3364 4874
rect 3379 4856 3409 4874
rect 3452 4844 3465 4874
rect 3495 4844 3508 4874
rect 3523 4856 3553 4874
rect 3596 4860 3610 4874
rect 3646 4860 3866 4874
rect 3597 4858 3610 4860
rect 3563 4846 3578 4858
rect 3560 4844 3582 4846
rect 3587 4844 3617 4858
rect 3678 4856 3831 4860
rect 3660 4844 3852 4856
rect 3895 4844 3925 4858
rect 3931 4844 3944 4874
rect 3959 4856 3989 4874
rect 4032 4844 4045 4874
rect 4075 4844 4088 4874
rect 4103 4856 4133 4874
rect 4176 4860 4190 4874
rect 4226 4860 4446 4874
rect 4177 4858 4190 4860
rect 4143 4846 4158 4858
rect 4140 4844 4162 4846
rect 4167 4844 4197 4858
rect 4258 4856 4411 4860
rect 4240 4844 4432 4856
rect 4475 4844 4505 4858
rect 4511 4844 4524 4874
rect 4539 4856 4569 4874
rect 4612 4844 4625 4874
rect 0 4830 4625 4844
rect 15 4726 28 4830
rect 73 4808 74 4818
rect 89 4808 102 4818
rect 73 4804 102 4808
rect 107 4804 137 4830
rect 155 4816 171 4818
rect 243 4816 296 4830
rect 244 4814 308 4816
rect 351 4814 366 4830
rect 415 4827 445 4830
rect 415 4824 451 4827
rect 381 4816 397 4818
rect 155 4804 170 4808
rect 73 4802 170 4804
rect 198 4802 366 4814
rect 382 4804 397 4808
rect 415 4805 454 4824
rect 473 4818 480 4819
rect 479 4811 480 4818
rect 463 4808 464 4811
rect 479 4808 492 4811
rect 415 4804 445 4805
rect 454 4804 460 4805
rect 463 4804 492 4808
rect 382 4803 492 4804
rect 382 4802 498 4803
rect 57 4794 108 4802
rect 57 4782 82 4794
rect 89 4782 108 4794
rect 139 4794 189 4802
rect 139 4786 155 4794
rect 162 4792 189 4794
rect 198 4792 419 4802
rect 162 4782 419 4792
rect 448 4794 498 4802
rect 448 4785 464 4794
rect 57 4774 108 4782
rect 155 4774 419 4782
rect 445 4782 464 4785
rect 471 4782 498 4794
rect 445 4774 498 4782
rect 73 4766 74 4774
rect 89 4766 102 4774
rect 73 4758 89 4766
rect 70 4751 89 4754
rect 70 4742 92 4751
rect 43 4732 92 4742
rect 43 4726 73 4732
rect 92 4727 97 4732
rect 15 4710 89 4726
rect 107 4718 137 4774
rect 172 4764 380 4774
rect 415 4770 460 4774
rect 463 4773 464 4774
rect 479 4773 492 4774
rect 198 4734 387 4764
rect 213 4731 387 4734
rect 206 4728 387 4731
rect 15 4708 28 4710
rect 43 4708 77 4710
rect 15 4692 89 4708
rect 116 4704 129 4718
rect 144 4704 160 4720
rect 206 4715 217 4728
rect -1 4670 0 4686
rect 15 4670 28 4692
rect 43 4670 73 4692
rect 116 4688 178 4704
rect 206 4697 217 4713
rect 222 4708 232 4728
rect 242 4708 256 4728
rect 259 4715 268 4728
rect 284 4715 293 4728
rect 222 4697 256 4708
rect 259 4697 268 4713
rect 284 4697 293 4713
rect 300 4708 310 4728
rect 320 4708 334 4728
rect 335 4715 346 4728
rect 300 4697 334 4708
rect 335 4697 346 4713
rect 392 4704 408 4720
rect 415 4718 445 4770
rect 479 4766 480 4773
rect 464 4758 480 4766
rect 451 4726 464 4745
rect 479 4726 509 4742
rect 451 4710 525 4726
rect 451 4708 464 4710
rect 479 4708 513 4710
rect 116 4686 129 4688
rect 144 4686 178 4688
rect 116 4670 178 4686
rect 222 4681 238 4684
rect 300 4681 330 4692
rect 378 4688 424 4704
rect 451 4692 525 4708
rect 378 4686 412 4688
rect 377 4670 424 4686
rect 451 4670 464 4692
rect 479 4670 509 4692
rect 536 4670 537 4686
rect 552 4670 565 4830
rect 595 4726 608 4830
rect 653 4808 654 4818
rect 669 4808 682 4818
rect 653 4804 682 4808
rect 687 4804 717 4830
rect 735 4816 751 4818
rect 823 4816 876 4830
rect 824 4814 888 4816
rect 931 4814 946 4830
rect 995 4827 1025 4830
rect 995 4824 1031 4827
rect 961 4816 977 4818
rect 735 4804 750 4808
rect 653 4802 750 4804
rect 778 4802 946 4814
rect 962 4804 977 4808
rect 995 4805 1034 4824
rect 1053 4818 1060 4819
rect 1059 4811 1060 4818
rect 1043 4808 1044 4811
rect 1059 4808 1072 4811
rect 995 4804 1025 4805
rect 1034 4804 1040 4805
rect 1043 4804 1072 4808
rect 962 4803 1072 4804
rect 962 4802 1078 4803
rect 637 4794 688 4802
rect 637 4782 662 4794
rect 669 4782 688 4794
rect 719 4794 769 4802
rect 719 4786 735 4794
rect 742 4792 769 4794
rect 778 4792 999 4802
rect 742 4782 999 4792
rect 1028 4794 1078 4802
rect 1028 4785 1044 4794
rect 637 4774 688 4782
rect 735 4774 999 4782
rect 1025 4782 1044 4785
rect 1051 4782 1078 4794
rect 1025 4774 1078 4782
rect 653 4766 654 4774
rect 669 4766 682 4774
rect 653 4758 669 4766
rect 650 4751 669 4754
rect 650 4742 672 4751
rect 623 4732 672 4742
rect 623 4726 653 4732
rect 672 4727 677 4732
rect 595 4710 669 4726
rect 687 4718 717 4774
rect 752 4764 960 4774
rect 995 4770 1040 4774
rect 1043 4773 1044 4774
rect 1059 4773 1072 4774
rect 778 4734 967 4764
rect 793 4731 967 4734
rect 786 4728 967 4731
rect 595 4708 608 4710
rect 623 4708 657 4710
rect 595 4692 669 4708
rect 696 4704 709 4718
rect 724 4704 740 4720
rect 786 4715 797 4728
rect 579 4670 580 4686
rect 595 4670 608 4692
rect 623 4670 653 4692
rect 696 4688 758 4704
rect 786 4697 797 4713
rect 802 4708 812 4728
rect 822 4708 836 4728
rect 839 4715 848 4728
rect 864 4715 873 4728
rect 802 4697 836 4708
rect 839 4697 848 4713
rect 864 4697 873 4713
rect 880 4708 890 4728
rect 900 4708 914 4728
rect 915 4715 926 4728
rect 880 4697 914 4708
rect 915 4697 926 4713
rect 972 4704 988 4720
rect 995 4718 1025 4770
rect 1059 4766 1060 4773
rect 1044 4758 1060 4766
rect 1031 4726 1044 4745
rect 1059 4726 1089 4742
rect 1031 4710 1105 4726
rect 1031 4708 1044 4710
rect 1059 4708 1093 4710
rect 696 4686 709 4688
rect 724 4686 758 4688
rect 696 4670 758 4686
rect 802 4681 818 4684
rect 880 4681 910 4692
rect 958 4688 1004 4704
rect 1031 4692 1105 4708
rect 958 4686 992 4688
rect 957 4670 1004 4686
rect 1031 4670 1044 4692
rect 1059 4670 1089 4692
rect 1116 4670 1117 4686
rect 1132 4670 1145 4830
rect 1175 4726 1188 4830
rect 1233 4808 1234 4818
rect 1249 4808 1262 4818
rect 1233 4804 1262 4808
rect 1267 4804 1297 4830
rect 1315 4816 1331 4818
rect 1403 4816 1456 4830
rect 1404 4814 1468 4816
rect 1511 4814 1526 4830
rect 1575 4827 1605 4830
rect 1575 4824 1611 4827
rect 1541 4816 1557 4818
rect 1315 4804 1330 4808
rect 1233 4802 1330 4804
rect 1358 4802 1526 4814
rect 1542 4804 1557 4808
rect 1575 4805 1614 4824
rect 1633 4818 1640 4819
rect 1639 4811 1640 4818
rect 1623 4808 1624 4811
rect 1639 4808 1652 4811
rect 1575 4804 1605 4805
rect 1614 4804 1620 4805
rect 1623 4804 1652 4808
rect 1542 4803 1652 4804
rect 1542 4802 1658 4803
rect 1217 4794 1268 4802
rect 1217 4782 1242 4794
rect 1249 4782 1268 4794
rect 1299 4794 1349 4802
rect 1299 4786 1315 4794
rect 1322 4792 1349 4794
rect 1358 4792 1579 4802
rect 1322 4782 1579 4792
rect 1608 4794 1658 4802
rect 1608 4785 1624 4794
rect 1217 4774 1268 4782
rect 1315 4774 1579 4782
rect 1605 4782 1624 4785
rect 1631 4782 1658 4794
rect 1605 4774 1658 4782
rect 1233 4766 1234 4774
rect 1249 4766 1262 4774
rect 1233 4758 1249 4766
rect 1230 4751 1249 4754
rect 1230 4742 1252 4751
rect 1203 4732 1252 4742
rect 1203 4726 1233 4732
rect 1252 4727 1257 4732
rect 1175 4710 1249 4726
rect 1267 4718 1297 4774
rect 1332 4764 1540 4774
rect 1575 4770 1620 4774
rect 1623 4773 1624 4774
rect 1639 4773 1652 4774
rect 1358 4734 1547 4764
rect 1373 4731 1547 4734
rect 1366 4728 1547 4731
rect 1175 4708 1188 4710
rect 1203 4708 1237 4710
rect 1175 4692 1249 4708
rect 1276 4704 1289 4718
rect 1304 4704 1320 4720
rect 1366 4715 1377 4728
rect 1159 4670 1160 4686
rect 1175 4670 1188 4692
rect 1203 4670 1233 4692
rect 1276 4688 1338 4704
rect 1366 4697 1377 4713
rect 1382 4708 1392 4728
rect 1402 4708 1416 4728
rect 1419 4715 1428 4728
rect 1444 4715 1453 4728
rect 1382 4697 1416 4708
rect 1419 4697 1428 4713
rect 1444 4697 1453 4713
rect 1460 4708 1470 4728
rect 1480 4708 1494 4728
rect 1495 4715 1506 4728
rect 1460 4697 1494 4708
rect 1495 4697 1506 4713
rect 1552 4704 1568 4720
rect 1575 4718 1605 4770
rect 1639 4766 1640 4773
rect 1624 4758 1640 4766
rect 1611 4726 1624 4745
rect 1639 4726 1669 4742
rect 1611 4710 1685 4726
rect 1611 4708 1624 4710
rect 1639 4708 1673 4710
rect 1276 4686 1289 4688
rect 1304 4686 1338 4688
rect 1276 4670 1338 4686
rect 1382 4681 1398 4684
rect 1460 4681 1490 4692
rect 1538 4688 1584 4704
rect 1611 4692 1685 4708
rect 1538 4686 1572 4688
rect 1537 4670 1584 4686
rect 1611 4670 1624 4692
rect 1639 4670 1669 4692
rect 1696 4670 1697 4686
rect 1712 4670 1725 4830
rect 1755 4726 1768 4830
rect 1813 4808 1814 4818
rect 1829 4808 1842 4818
rect 1813 4804 1842 4808
rect 1847 4804 1877 4830
rect 1895 4816 1911 4818
rect 1983 4816 2036 4830
rect 1984 4814 2048 4816
rect 2091 4814 2106 4830
rect 2155 4827 2185 4830
rect 2155 4824 2191 4827
rect 2121 4816 2137 4818
rect 1895 4804 1910 4808
rect 1813 4802 1910 4804
rect 1938 4802 2106 4814
rect 2122 4804 2137 4808
rect 2155 4805 2194 4824
rect 2213 4818 2220 4819
rect 2219 4811 2220 4818
rect 2203 4808 2204 4811
rect 2219 4808 2232 4811
rect 2155 4804 2185 4805
rect 2194 4804 2200 4805
rect 2203 4804 2232 4808
rect 2122 4803 2232 4804
rect 2122 4802 2238 4803
rect 1797 4794 1848 4802
rect 1797 4782 1822 4794
rect 1829 4782 1848 4794
rect 1879 4794 1929 4802
rect 1879 4786 1895 4794
rect 1902 4792 1929 4794
rect 1938 4792 2159 4802
rect 1902 4782 2159 4792
rect 2188 4794 2238 4802
rect 2188 4785 2204 4794
rect 1797 4774 1848 4782
rect 1895 4774 2159 4782
rect 2185 4782 2204 4785
rect 2211 4782 2238 4794
rect 2185 4774 2238 4782
rect 1813 4766 1814 4774
rect 1829 4766 1842 4774
rect 1813 4758 1829 4766
rect 1810 4751 1829 4754
rect 1810 4742 1832 4751
rect 1783 4732 1832 4742
rect 1783 4726 1813 4732
rect 1832 4727 1837 4732
rect 1755 4710 1829 4726
rect 1847 4718 1877 4774
rect 1912 4764 2120 4774
rect 2155 4770 2200 4774
rect 2203 4773 2204 4774
rect 2219 4773 2232 4774
rect 1938 4734 2127 4764
rect 1953 4731 2127 4734
rect 1946 4728 2127 4731
rect 1755 4708 1768 4710
rect 1783 4708 1817 4710
rect 1755 4692 1829 4708
rect 1856 4704 1869 4718
rect 1884 4704 1900 4720
rect 1946 4715 1957 4728
rect 1739 4670 1740 4686
rect 1755 4670 1768 4692
rect 1783 4670 1813 4692
rect 1856 4688 1918 4704
rect 1946 4697 1957 4713
rect 1962 4708 1972 4728
rect 1982 4708 1996 4728
rect 1999 4715 2008 4728
rect 2024 4715 2033 4728
rect 1962 4697 1996 4708
rect 1999 4697 2008 4713
rect 2024 4697 2033 4713
rect 2040 4708 2050 4728
rect 2060 4708 2074 4728
rect 2075 4715 2086 4728
rect 2040 4697 2074 4708
rect 2075 4697 2086 4713
rect 2132 4704 2148 4720
rect 2155 4718 2185 4770
rect 2219 4766 2220 4773
rect 2204 4758 2220 4766
rect 2191 4726 2204 4745
rect 2219 4726 2249 4742
rect 2191 4710 2265 4726
rect 2191 4708 2204 4710
rect 2219 4708 2253 4710
rect 1856 4686 1869 4688
rect 1884 4686 1918 4688
rect 1856 4670 1918 4686
rect 1962 4681 1978 4684
rect 2040 4681 2070 4692
rect 2118 4688 2164 4704
rect 2191 4692 2265 4708
rect 2118 4686 2152 4688
rect 2117 4670 2164 4686
rect 2191 4670 2204 4692
rect 2219 4670 2249 4692
rect 2276 4670 2277 4686
rect 2292 4670 2305 4830
rect 2335 4726 2348 4830
rect 2393 4808 2394 4818
rect 2409 4808 2422 4818
rect 2393 4804 2422 4808
rect 2427 4804 2457 4830
rect 2475 4816 2491 4818
rect 2563 4816 2616 4830
rect 2564 4814 2628 4816
rect 2671 4814 2686 4830
rect 2735 4827 2765 4830
rect 2735 4824 2771 4827
rect 2701 4816 2717 4818
rect 2475 4804 2490 4808
rect 2393 4802 2490 4804
rect 2518 4802 2686 4814
rect 2702 4804 2717 4808
rect 2735 4805 2774 4824
rect 2793 4818 2800 4819
rect 2799 4811 2800 4818
rect 2783 4808 2784 4811
rect 2799 4808 2812 4811
rect 2735 4804 2765 4805
rect 2774 4804 2780 4805
rect 2783 4804 2812 4808
rect 2702 4803 2812 4804
rect 2702 4802 2818 4803
rect 2377 4794 2428 4802
rect 2377 4782 2402 4794
rect 2409 4782 2428 4794
rect 2459 4794 2509 4802
rect 2459 4786 2475 4794
rect 2482 4792 2509 4794
rect 2518 4792 2739 4802
rect 2482 4782 2739 4792
rect 2768 4794 2818 4802
rect 2768 4785 2784 4794
rect 2377 4774 2428 4782
rect 2475 4774 2739 4782
rect 2765 4782 2784 4785
rect 2791 4782 2818 4794
rect 2765 4774 2818 4782
rect 2393 4766 2394 4774
rect 2409 4766 2422 4774
rect 2393 4758 2409 4766
rect 2390 4751 2409 4754
rect 2390 4742 2412 4751
rect 2363 4732 2412 4742
rect 2363 4726 2393 4732
rect 2412 4727 2417 4732
rect 2335 4710 2409 4726
rect 2427 4718 2457 4774
rect 2492 4764 2700 4774
rect 2735 4770 2780 4774
rect 2783 4773 2784 4774
rect 2799 4773 2812 4774
rect 2518 4734 2707 4764
rect 2533 4731 2707 4734
rect 2526 4728 2707 4731
rect 2335 4708 2348 4710
rect 2363 4708 2397 4710
rect 2335 4692 2409 4708
rect 2436 4704 2449 4718
rect 2464 4704 2480 4720
rect 2526 4715 2537 4728
rect 2319 4670 2320 4686
rect 2335 4670 2348 4692
rect 2363 4670 2393 4692
rect 2436 4688 2498 4704
rect 2526 4697 2537 4713
rect 2542 4708 2552 4728
rect 2562 4708 2576 4728
rect 2579 4715 2588 4728
rect 2604 4715 2613 4728
rect 2542 4697 2576 4708
rect 2579 4697 2588 4713
rect 2604 4697 2613 4713
rect 2620 4708 2630 4728
rect 2640 4708 2654 4728
rect 2655 4715 2666 4728
rect 2620 4697 2654 4708
rect 2655 4697 2666 4713
rect 2712 4704 2728 4720
rect 2735 4718 2765 4770
rect 2799 4766 2800 4773
rect 2784 4758 2800 4766
rect 2771 4726 2784 4745
rect 2799 4726 2829 4742
rect 2771 4710 2845 4726
rect 2771 4708 2784 4710
rect 2799 4708 2833 4710
rect 2436 4686 2449 4688
rect 2464 4686 2498 4688
rect 2436 4670 2498 4686
rect 2542 4681 2558 4684
rect 2620 4681 2650 4692
rect 2698 4688 2744 4704
rect 2771 4692 2845 4708
rect 2698 4686 2732 4688
rect 2697 4670 2744 4686
rect 2771 4670 2784 4692
rect 2799 4670 2829 4692
rect 2856 4670 2857 4686
rect 2872 4670 2885 4830
rect 2915 4726 2928 4830
rect 2973 4808 2974 4818
rect 2989 4808 3002 4818
rect 2973 4804 3002 4808
rect 3007 4804 3037 4830
rect 3055 4816 3071 4818
rect 3143 4816 3196 4830
rect 3144 4814 3208 4816
rect 3251 4814 3266 4830
rect 3315 4827 3345 4830
rect 3315 4824 3351 4827
rect 3281 4816 3297 4818
rect 3055 4804 3070 4808
rect 2973 4802 3070 4804
rect 3098 4802 3266 4814
rect 3282 4804 3297 4808
rect 3315 4805 3354 4824
rect 3373 4818 3380 4819
rect 3379 4811 3380 4818
rect 3363 4808 3364 4811
rect 3379 4808 3392 4811
rect 3315 4804 3345 4805
rect 3354 4804 3360 4805
rect 3363 4804 3392 4808
rect 3282 4803 3392 4804
rect 3282 4802 3398 4803
rect 2957 4794 3008 4802
rect 2957 4782 2982 4794
rect 2989 4782 3008 4794
rect 3039 4794 3089 4802
rect 3039 4786 3055 4794
rect 3062 4792 3089 4794
rect 3098 4792 3319 4802
rect 3062 4782 3319 4792
rect 3348 4794 3398 4802
rect 3348 4785 3364 4794
rect 2957 4774 3008 4782
rect 3055 4774 3319 4782
rect 3345 4782 3364 4785
rect 3371 4782 3398 4794
rect 3345 4774 3398 4782
rect 2973 4766 2974 4774
rect 2989 4766 3002 4774
rect 2973 4758 2989 4766
rect 2970 4751 2989 4754
rect 2970 4742 2992 4751
rect 2943 4732 2992 4742
rect 2943 4726 2973 4732
rect 2992 4727 2997 4732
rect 2915 4710 2989 4726
rect 3007 4718 3037 4774
rect 3072 4764 3280 4774
rect 3315 4770 3360 4774
rect 3363 4773 3364 4774
rect 3379 4773 3392 4774
rect 3098 4734 3287 4764
rect 3113 4731 3287 4734
rect 3106 4728 3287 4731
rect 2915 4708 2928 4710
rect 2943 4708 2977 4710
rect 2915 4692 2989 4708
rect 3016 4704 3029 4718
rect 3044 4704 3060 4720
rect 3106 4715 3117 4728
rect 2899 4670 2900 4686
rect 2915 4670 2928 4692
rect 2943 4670 2973 4692
rect 3016 4688 3078 4704
rect 3106 4697 3117 4713
rect 3122 4708 3132 4728
rect 3142 4708 3156 4728
rect 3159 4715 3168 4728
rect 3184 4715 3193 4728
rect 3122 4697 3156 4708
rect 3159 4697 3168 4713
rect 3184 4697 3193 4713
rect 3200 4708 3210 4728
rect 3220 4708 3234 4728
rect 3235 4715 3246 4728
rect 3200 4697 3234 4708
rect 3235 4697 3246 4713
rect 3292 4704 3308 4720
rect 3315 4718 3345 4770
rect 3379 4766 3380 4773
rect 3364 4758 3380 4766
rect 3351 4726 3364 4745
rect 3379 4726 3409 4742
rect 3351 4710 3425 4726
rect 3351 4708 3364 4710
rect 3379 4708 3413 4710
rect 3016 4686 3029 4688
rect 3044 4686 3078 4688
rect 3016 4670 3078 4686
rect 3122 4681 3138 4684
rect 3200 4681 3230 4692
rect 3278 4688 3324 4704
rect 3351 4692 3425 4708
rect 3278 4686 3312 4688
rect 3277 4670 3324 4686
rect 3351 4670 3364 4692
rect 3379 4670 3409 4692
rect 3436 4670 3437 4686
rect 3452 4670 3465 4830
rect 3495 4726 3508 4830
rect 3553 4808 3554 4818
rect 3569 4808 3582 4818
rect 3553 4804 3582 4808
rect 3587 4804 3617 4830
rect 3635 4816 3651 4818
rect 3723 4816 3776 4830
rect 3724 4814 3788 4816
rect 3831 4814 3846 4830
rect 3895 4827 3925 4830
rect 3895 4824 3931 4827
rect 3861 4816 3877 4818
rect 3635 4804 3650 4808
rect 3553 4802 3650 4804
rect 3678 4802 3846 4814
rect 3862 4804 3877 4808
rect 3895 4805 3934 4824
rect 3953 4818 3960 4819
rect 3959 4811 3960 4818
rect 3943 4808 3944 4811
rect 3959 4808 3972 4811
rect 3895 4804 3925 4805
rect 3934 4804 3940 4805
rect 3943 4804 3972 4808
rect 3862 4803 3972 4804
rect 3862 4802 3978 4803
rect 3537 4794 3588 4802
rect 3537 4782 3562 4794
rect 3569 4782 3588 4794
rect 3619 4794 3669 4802
rect 3619 4786 3635 4794
rect 3642 4792 3669 4794
rect 3678 4792 3899 4802
rect 3642 4782 3899 4792
rect 3928 4794 3978 4802
rect 3928 4785 3944 4794
rect 3537 4774 3588 4782
rect 3635 4774 3899 4782
rect 3925 4782 3944 4785
rect 3951 4782 3978 4794
rect 3925 4774 3978 4782
rect 3553 4766 3554 4774
rect 3569 4766 3582 4774
rect 3553 4758 3569 4766
rect 3550 4751 3569 4754
rect 3550 4742 3572 4751
rect 3523 4732 3572 4742
rect 3523 4726 3553 4732
rect 3572 4727 3577 4732
rect 3495 4710 3569 4726
rect 3587 4718 3617 4774
rect 3652 4764 3860 4774
rect 3895 4770 3940 4774
rect 3943 4773 3944 4774
rect 3959 4773 3972 4774
rect 3678 4734 3867 4764
rect 3693 4731 3867 4734
rect 3686 4728 3867 4731
rect 3495 4708 3508 4710
rect 3523 4708 3557 4710
rect 3495 4692 3569 4708
rect 3596 4704 3609 4718
rect 3624 4704 3640 4720
rect 3686 4715 3697 4728
rect 3479 4670 3480 4686
rect 3495 4670 3508 4692
rect 3523 4670 3553 4692
rect 3596 4688 3658 4704
rect 3686 4697 3697 4713
rect 3702 4708 3712 4728
rect 3722 4708 3736 4728
rect 3739 4715 3748 4728
rect 3764 4715 3773 4728
rect 3702 4697 3736 4708
rect 3739 4697 3748 4713
rect 3764 4697 3773 4713
rect 3780 4708 3790 4728
rect 3800 4708 3814 4728
rect 3815 4715 3826 4728
rect 3780 4697 3814 4708
rect 3815 4697 3826 4713
rect 3872 4704 3888 4720
rect 3895 4718 3925 4770
rect 3959 4766 3960 4773
rect 3944 4758 3960 4766
rect 3931 4726 3944 4745
rect 3959 4726 3989 4742
rect 3931 4710 4005 4726
rect 3931 4708 3944 4710
rect 3959 4708 3993 4710
rect 3596 4686 3609 4688
rect 3624 4686 3658 4688
rect 3596 4670 3658 4686
rect 3702 4681 3718 4684
rect 3780 4681 3810 4692
rect 3858 4688 3904 4704
rect 3931 4692 4005 4708
rect 3858 4686 3892 4688
rect 3857 4670 3904 4686
rect 3931 4670 3944 4692
rect 3959 4670 3989 4692
rect 4016 4670 4017 4686
rect 4032 4670 4045 4830
rect 4075 4726 4088 4830
rect 4133 4808 4134 4818
rect 4149 4808 4162 4818
rect 4133 4804 4162 4808
rect 4167 4804 4197 4830
rect 4215 4816 4231 4818
rect 4303 4816 4356 4830
rect 4304 4814 4368 4816
rect 4411 4814 4426 4830
rect 4475 4827 4505 4830
rect 4475 4824 4511 4827
rect 4441 4816 4457 4818
rect 4215 4804 4230 4808
rect 4133 4802 4230 4804
rect 4258 4802 4426 4814
rect 4442 4804 4457 4808
rect 4475 4805 4514 4824
rect 4533 4818 4540 4819
rect 4539 4811 4540 4818
rect 4523 4808 4524 4811
rect 4539 4808 4552 4811
rect 4475 4804 4505 4805
rect 4514 4804 4520 4805
rect 4523 4804 4552 4808
rect 4442 4803 4552 4804
rect 4442 4802 4558 4803
rect 4117 4794 4168 4802
rect 4117 4782 4142 4794
rect 4149 4782 4168 4794
rect 4199 4794 4249 4802
rect 4199 4786 4215 4794
rect 4222 4792 4249 4794
rect 4258 4792 4479 4802
rect 4222 4782 4479 4792
rect 4508 4794 4558 4802
rect 4508 4785 4524 4794
rect 4117 4774 4168 4782
rect 4215 4774 4479 4782
rect 4505 4782 4524 4785
rect 4531 4782 4558 4794
rect 4505 4774 4558 4782
rect 4133 4766 4134 4774
rect 4149 4766 4162 4774
rect 4133 4758 4149 4766
rect 4130 4751 4149 4754
rect 4130 4742 4152 4751
rect 4103 4732 4152 4742
rect 4103 4726 4133 4732
rect 4152 4727 4157 4732
rect 4075 4710 4149 4726
rect 4167 4718 4197 4774
rect 4232 4764 4440 4774
rect 4475 4770 4520 4774
rect 4523 4773 4524 4774
rect 4539 4773 4552 4774
rect 4258 4734 4447 4764
rect 4273 4731 4447 4734
rect 4266 4728 4447 4731
rect 4075 4708 4088 4710
rect 4103 4708 4137 4710
rect 4075 4692 4149 4708
rect 4176 4704 4189 4718
rect 4204 4704 4220 4720
rect 4266 4715 4277 4728
rect 4059 4670 4060 4686
rect 4075 4670 4088 4692
rect 4103 4670 4133 4692
rect 4176 4688 4238 4704
rect 4266 4697 4277 4713
rect 4282 4708 4292 4728
rect 4302 4708 4316 4728
rect 4319 4715 4328 4728
rect 4344 4715 4353 4728
rect 4282 4697 4316 4708
rect 4319 4697 4328 4713
rect 4344 4697 4353 4713
rect 4360 4708 4370 4728
rect 4380 4708 4394 4728
rect 4395 4715 4406 4728
rect 4360 4697 4394 4708
rect 4395 4697 4406 4713
rect 4452 4704 4468 4720
rect 4475 4718 4505 4770
rect 4539 4766 4540 4773
rect 4524 4758 4540 4766
rect 4511 4726 4524 4745
rect 4539 4726 4569 4742
rect 4511 4710 4585 4726
rect 4511 4708 4524 4710
rect 4539 4708 4573 4710
rect 4176 4686 4189 4688
rect 4204 4686 4238 4688
rect 4176 4670 4238 4686
rect 4282 4681 4298 4684
rect 4360 4681 4390 4692
rect 4438 4688 4484 4704
rect 4511 4692 4585 4708
rect 4438 4686 4472 4688
rect 4437 4670 4484 4686
rect 4511 4670 4524 4692
rect 4539 4670 4569 4692
rect 4596 4670 4597 4686
rect 4612 4670 4625 4830
rect -7 4662 34 4670
rect -7 4636 8 4662
rect 15 4636 34 4662
rect 98 4658 160 4670
rect 172 4658 247 4670
rect 305 4658 380 4670
rect 392 4658 423 4670
rect 429 4658 464 4670
rect 98 4656 260 4658
rect -7 4628 34 4636
rect 116 4632 129 4656
rect 144 4654 159 4656
rect -1 4618 0 4628
rect 15 4618 28 4628
rect 43 4618 73 4632
rect 116 4618 159 4632
rect 183 4629 190 4636
rect 193 4632 260 4656
rect 292 4656 464 4658
rect 262 4634 290 4638
rect 292 4634 372 4656
rect 393 4654 408 4656
rect 262 4632 372 4634
rect 193 4628 372 4632
rect 166 4618 196 4628
rect 198 4618 351 4628
rect 359 4618 389 4628
rect 393 4618 423 4632
rect 451 4618 464 4656
rect 536 4662 571 4670
rect 536 4636 537 4662
rect 544 4636 571 4662
rect 479 4618 509 4632
rect 536 4628 571 4636
rect 573 4662 614 4670
rect 573 4636 588 4662
rect 595 4636 614 4662
rect 678 4658 740 4670
rect 752 4658 827 4670
rect 885 4658 960 4670
rect 972 4658 1003 4670
rect 1009 4658 1044 4670
rect 678 4656 840 4658
rect 573 4628 614 4636
rect 696 4632 709 4656
rect 724 4654 739 4656
rect 536 4618 537 4628
rect 552 4618 565 4628
rect 579 4618 580 4628
rect 595 4618 608 4628
rect 623 4618 653 4632
rect 696 4618 739 4632
rect 763 4629 770 4636
rect 773 4632 840 4656
rect 872 4656 1044 4658
rect 842 4634 870 4638
rect 872 4634 952 4656
rect 973 4654 988 4656
rect 842 4632 952 4634
rect 773 4628 952 4632
rect 746 4618 776 4628
rect 778 4618 931 4628
rect 939 4618 969 4628
rect 973 4618 1003 4632
rect 1031 4618 1044 4656
rect 1116 4662 1151 4670
rect 1116 4636 1117 4662
rect 1124 4636 1151 4662
rect 1059 4618 1089 4632
rect 1116 4628 1151 4636
rect 1153 4662 1194 4670
rect 1153 4636 1168 4662
rect 1175 4636 1194 4662
rect 1258 4658 1320 4670
rect 1332 4658 1407 4670
rect 1465 4658 1540 4670
rect 1552 4658 1583 4670
rect 1589 4658 1624 4670
rect 1258 4656 1420 4658
rect 1153 4628 1194 4636
rect 1276 4632 1289 4656
rect 1304 4654 1319 4656
rect 1116 4618 1117 4628
rect 1132 4618 1145 4628
rect 1159 4618 1160 4628
rect 1175 4618 1188 4628
rect 1203 4618 1233 4632
rect 1276 4618 1319 4632
rect 1343 4629 1350 4636
rect 1353 4632 1420 4656
rect 1452 4656 1624 4658
rect 1422 4634 1450 4638
rect 1452 4634 1532 4656
rect 1553 4654 1568 4656
rect 1422 4632 1532 4634
rect 1353 4628 1532 4632
rect 1326 4618 1356 4628
rect 1358 4618 1511 4628
rect 1519 4618 1549 4628
rect 1553 4618 1583 4632
rect 1611 4618 1624 4656
rect 1696 4662 1731 4670
rect 1696 4636 1697 4662
rect 1704 4636 1731 4662
rect 1639 4618 1669 4632
rect 1696 4628 1731 4636
rect 1733 4662 1774 4670
rect 1733 4636 1748 4662
rect 1755 4636 1774 4662
rect 1838 4658 1900 4670
rect 1912 4658 1987 4670
rect 2045 4658 2120 4670
rect 2132 4658 2163 4670
rect 2169 4658 2204 4670
rect 1838 4656 2000 4658
rect 1733 4628 1774 4636
rect 1856 4632 1869 4656
rect 1884 4654 1899 4656
rect 1696 4618 1697 4628
rect 1712 4618 1725 4628
rect 1739 4618 1740 4628
rect 1755 4618 1768 4628
rect 1783 4618 1813 4632
rect 1856 4618 1899 4632
rect 1923 4629 1930 4636
rect 1933 4632 2000 4656
rect 2032 4656 2204 4658
rect 2002 4634 2030 4638
rect 2032 4634 2112 4656
rect 2133 4654 2148 4656
rect 2002 4632 2112 4634
rect 1933 4628 2112 4632
rect 1906 4618 1936 4628
rect 1938 4618 2091 4628
rect 2099 4618 2129 4628
rect 2133 4618 2163 4632
rect 2191 4618 2204 4656
rect 2276 4662 2311 4670
rect 2276 4636 2277 4662
rect 2284 4636 2311 4662
rect 2219 4618 2249 4632
rect 2276 4628 2311 4636
rect 2313 4662 2354 4670
rect 2313 4636 2328 4662
rect 2335 4636 2354 4662
rect 2418 4658 2480 4670
rect 2492 4658 2567 4670
rect 2625 4658 2700 4670
rect 2712 4658 2743 4670
rect 2749 4658 2784 4670
rect 2418 4656 2580 4658
rect 2313 4628 2354 4636
rect 2436 4632 2449 4656
rect 2464 4654 2479 4656
rect 2276 4618 2277 4628
rect 2292 4618 2305 4628
rect 2319 4618 2320 4628
rect 2335 4618 2348 4628
rect 2363 4618 2393 4632
rect 2436 4618 2479 4632
rect 2503 4629 2510 4636
rect 2513 4632 2580 4656
rect 2612 4656 2784 4658
rect 2582 4634 2610 4638
rect 2612 4634 2692 4656
rect 2713 4654 2728 4656
rect 2582 4632 2692 4634
rect 2513 4628 2692 4632
rect 2486 4618 2516 4628
rect 2518 4618 2671 4628
rect 2679 4618 2709 4628
rect 2713 4618 2743 4632
rect 2771 4618 2784 4656
rect 2856 4662 2891 4670
rect 2856 4636 2857 4662
rect 2864 4636 2891 4662
rect 2799 4618 2829 4632
rect 2856 4628 2891 4636
rect 2893 4662 2934 4670
rect 2893 4636 2908 4662
rect 2915 4636 2934 4662
rect 2998 4658 3060 4670
rect 3072 4658 3147 4670
rect 3205 4658 3280 4670
rect 3292 4658 3323 4670
rect 3329 4658 3364 4670
rect 2998 4656 3160 4658
rect 2893 4628 2934 4636
rect 3016 4632 3029 4656
rect 3044 4654 3059 4656
rect 2856 4618 2857 4628
rect 2872 4618 2885 4628
rect 2899 4618 2900 4628
rect 2915 4618 2928 4628
rect 2943 4618 2973 4632
rect 3016 4618 3059 4632
rect 3083 4629 3090 4636
rect 3093 4632 3160 4656
rect 3192 4656 3364 4658
rect 3162 4634 3190 4638
rect 3192 4634 3272 4656
rect 3293 4654 3308 4656
rect 3162 4632 3272 4634
rect 3093 4628 3272 4632
rect 3066 4618 3096 4628
rect 3098 4618 3251 4628
rect 3259 4618 3289 4628
rect 3293 4618 3323 4632
rect 3351 4618 3364 4656
rect 3436 4662 3471 4670
rect 3436 4636 3437 4662
rect 3444 4636 3471 4662
rect 3379 4618 3409 4632
rect 3436 4628 3471 4636
rect 3473 4662 3514 4670
rect 3473 4636 3488 4662
rect 3495 4636 3514 4662
rect 3578 4658 3640 4670
rect 3652 4658 3727 4670
rect 3785 4658 3860 4670
rect 3872 4658 3903 4670
rect 3909 4658 3944 4670
rect 3578 4656 3740 4658
rect 3473 4628 3514 4636
rect 3596 4632 3609 4656
rect 3624 4654 3639 4656
rect 3436 4618 3437 4628
rect 3452 4618 3465 4628
rect 3479 4618 3480 4628
rect 3495 4618 3508 4628
rect 3523 4618 3553 4632
rect 3596 4618 3639 4632
rect 3663 4629 3670 4636
rect 3673 4632 3740 4656
rect 3772 4656 3944 4658
rect 3742 4634 3770 4638
rect 3772 4634 3852 4656
rect 3873 4654 3888 4656
rect 3742 4632 3852 4634
rect 3673 4628 3852 4632
rect 3646 4618 3676 4628
rect 3678 4618 3831 4628
rect 3839 4618 3869 4628
rect 3873 4618 3903 4632
rect 3931 4618 3944 4656
rect 4016 4662 4051 4670
rect 4016 4636 4017 4662
rect 4024 4636 4051 4662
rect 3959 4618 3989 4632
rect 4016 4628 4051 4636
rect 4053 4662 4094 4670
rect 4053 4636 4068 4662
rect 4075 4636 4094 4662
rect 4158 4658 4220 4670
rect 4232 4658 4307 4670
rect 4365 4658 4440 4670
rect 4452 4658 4483 4670
rect 4489 4658 4524 4670
rect 4158 4656 4320 4658
rect 4053 4628 4094 4636
rect 4176 4632 4189 4656
rect 4204 4654 4219 4656
rect 4016 4618 4017 4628
rect 4032 4618 4045 4628
rect 4059 4618 4060 4628
rect 4075 4618 4088 4628
rect 4103 4618 4133 4632
rect 4176 4618 4219 4632
rect 4243 4629 4250 4636
rect 4253 4632 4320 4656
rect 4352 4656 4524 4658
rect 4322 4634 4350 4638
rect 4352 4634 4432 4656
rect 4453 4654 4468 4656
rect 4322 4632 4432 4634
rect 4253 4628 4432 4632
rect 4226 4618 4256 4628
rect 4258 4618 4411 4628
rect 4419 4618 4449 4628
rect 4453 4618 4483 4632
rect 4511 4618 4524 4656
rect 4596 4662 4631 4670
rect 4596 4636 4597 4662
rect 4604 4636 4631 4662
rect 4539 4618 4569 4632
rect 4596 4628 4631 4636
rect 4596 4618 4597 4628
rect 4612 4618 4625 4628
rect -1 4612 4625 4618
rect 0 4604 4625 4612
rect 15 4574 28 4604
rect 43 4586 73 4604
rect 116 4590 130 4604
rect 166 4590 386 4604
rect 117 4588 130 4590
rect 83 4576 98 4588
rect 80 4574 102 4576
rect 107 4574 137 4588
rect 198 4586 351 4590
rect 180 4574 372 4586
rect 415 4574 445 4588
rect 451 4574 464 4604
rect 479 4586 509 4604
rect 552 4574 565 4604
rect 595 4574 608 4604
rect 623 4586 653 4604
rect 696 4590 710 4604
rect 746 4590 966 4604
rect 697 4588 710 4590
rect 663 4576 678 4588
rect 660 4574 682 4576
rect 687 4574 717 4588
rect 778 4586 931 4590
rect 760 4574 952 4586
rect 995 4574 1025 4588
rect 1031 4574 1044 4604
rect 1059 4586 1089 4604
rect 1132 4574 1145 4604
rect 1175 4574 1188 4604
rect 1203 4586 1233 4604
rect 1276 4590 1290 4604
rect 1326 4590 1546 4604
rect 1277 4588 1290 4590
rect 1243 4576 1258 4588
rect 1240 4574 1262 4576
rect 1267 4574 1297 4588
rect 1358 4586 1511 4590
rect 1340 4574 1532 4586
rect 1575 4574 1605 4588
rect 1611 4574 1624 4604
rect 1639 4586 1669 4604
rect 1712 4574 1725 4604
rect 1755 4574 1768 4604
rect 1783 4586 1813 4604
rect 1856 4590 1870 4604
rect 1906 4590 2126 4604
rect 1857 4588 1870 4590
rect 1823 4576 1838 4588
rect 1820 4574 1842 4576
rect 1847 4574 1877 4588
rect 1938 4586 2091 4590
rect 1920 4574 2112 4586
rect 2155 4574 2185 4588
rect 2191 4574 2204 4604
rect 2219 4586 2249 4604
rect 2292 4574 2305 4604
rect 2335 4574 2348 4604
rect 2363 4586 2393 4604
rect 2436 4590 2450 4604
rect 2486 4590 2706 4604
rect 2437 4588 2450 4590
rect 2403 4576 2418 4588
rect 2400 4574 2422 4576
rect 2427 4574 2457 4588
rect 2518 4586 2671 4590
rect 2500 4574 2692 4586
rect 2735 4574 2765 4588
rect 2771 4574 2784 4604
rect 2799 4586 2829 4604
rect 2872 4574 2885 4604
rect 2915 4574 2928 4604
rect 2943 4586 2973 4604
rect 3016 4590 3030 4604
rect 3066 4590 3286 4604
rect 3017 4588 3030 4590
rect 2983 4576 2998 4588
rect 2980 4574 3002 4576
rect 3007 4574 3037 4588
rect 3098 4586 3251 4590
rect 3080 4574 3272 4586
rect 3315 4574 3345 4588
rect 3351 4574 3364 4604
rect 3379 4586 3409 4604
rect 3452 4574 3465 4604
rect 3495 4574 3508 4604
rect 3523 4586 3553 4604
rect 3596 4590 3610 4604
rect 3646 4590 3866 4604
rect 3597 4588 3610 4590
rect 3563 4576 3578 4588
rect 3560 4574 3582 4576
rect 3587 4574 3617 4588
rect 3678 4586 3831 4590
rect 3660 4574 3852 4586
rect 3895 4574 3925 4588
rect 3931 4574 3944 4604
rect 3959 4586 3989 4604
rect 4032 4574 4045 4604
rect 4075 4574 4088 4604
rect 4103 4586 4133 4604
rect 4176 4590 4190 4604
rect 4226 4590 4446 4604
rect 4177 4588 4190 4590
rect 4143 4576 4158 4588
rect 4140 4574 4162 4576
rect 4167 4574 4197 4588
rect 4258 4586 4411 4590
rect 4240 4574 4432 4586
rect 4475 4574 4505 4588
rect 4511 4574 4524 4604
rect 4539 4586 4569 4604
rect 4612 4574 4625 4604
rect 0 4560 4625 4574
rect 15 4456 28 4560
rect 73 4538 74 4548
rect 89 4538 102 4548
rect 73 4534 102 4538
rect 107 4534 137 4560
rect 155 4546 171 4548
rect 243 4546 296 4560
rect 244 4544 308 4546
rect 351 4544 366 4560
rect 415 4557 445 4560
rect 415 4554 451 4557
rect 381 4546 397 4548
rect 155 4534 170 4538
rect 73 4532 170 4534
rect 198 4532 366 4544
rect 382 4534 397 4538
rect 415 4535 454 4554
rect 473 4548 480 4549
rect 479 4541 480 4548
rect 463 4538 464 4541
rect 479 4538 492 4541
rect 415 4534 445 4535
rect 454 4534 460 4535
rect 463 4534 492 4538
rect 382 4533 492 4534
rect 382 4532 498 4533
rect 57 4524 108 4532
rect 57 4512 82 4524
rect 89 4512 108 4524
rect 139 4524 189 4532
rect 139 4516 155 4524
rect 162 4522 189 4524
rect 198 4522 419 4532
rect 162 4512 419 4522
rect 448 4524 498 4532
rect 448 4515 464 4524
rect 57 4504 108 4512
rect 155 4504 419 4512
rect 445 4512 464 4515
rect 471 4512 498 4524
rect 445 4504 498 4512
rect 73 4496 74 4504
rect 89 4496 102 4504
rect 73 4488 89 4496
rect 70 4481 89 4484
rect 70 4472 92 4481
rect 43 4462 92 4472
rect 43 4456 73 4462
rect 92 4457 97 4462
rect 15 4440 89 4456
rect 107 4448 137 4504
rect 172 4494 380 4504
rect 415 4500 460 4504
rect 463 4503 464 4504
rect 479 4503 492 4504
rect 198 4464 387 4494
rect 213 4461 387 4464
rect 206 4458 387 4461
rect 15 4438 28 4440
rect 43 4438 77 4440
rect 15 4422 89 4438
rect 116 4434 129 4448
rect 144 4434 160 4450
rect 206 4445 217 4458
rect -1 4400 0 4416
rect 15 4400 28 4422
rect 43 4400 73 4422
rect 116 4418 178 4434
rect 206 4427 217 4443
rect 222 4438 232 4458
rect 242 4438 256 4458
rect 259 4445 268 4458
rect 284 4445 293 4458
rect 222 4427 256 4438
rect 259 4427 268 4443
rect 284 4427 293 4443
rect 300 4438 310 4458
rect 320 4438 334 4458
rect 335 4445 346 4458
rect 300 4427 334 4438
rect 335 4427 346 4443
rect 392 4434 408 4450
rect 415 4448 445 4500
rect 479 4496 480 4503
rect 464 4488 480 4496
rect 451 4456 464 4475
rect 479 4456 509 4472
rect 451 4440 525 4456
rect 451 4438 464 4440
rect 479 4438 513 4440
rect 116 4416 129 4418
rect 144 4416 178 4418
rect 116 4400 178 4416
rect 222 4411 238 4414
rect 300 4411 330 4422
rect 378 4418 424 4434
rect 451 4422 525 4438
rect 378 4416 412 4418
rect 377 4400 424 4416
rect 451 4400 464 4422
rect 479 4400 509 4422
rect 536 4400 537 4416
rect 552 4400 565 4560
rect 595 4456 608 4560
rect 653 4538 654 4548
rect 669 4538 682 4548
rect 653 4534 682 4538
rect 687 4534 717 4560
rect 735 4546 751 4548
rect 823 4546 876 4560
rect 824 4544 888 4546
rect 931 4544 946 4560
rect 995 4557 1025 4560
rect 995 4554 1031 4557
rect 961 4546 977 4548
rect 735 4534 750 4538
rect 653 4532 750 4534
rect 778 4532 946 4544
rect 962 4534 977 4538
rect 995 4535 1034 4554
rect 1053 4548 1060 4549
rect 1059 4541 1060 4548
rect 1043 4538 1044 4541
rect 1059 4538 1072 4541
rect 995 4534 1025 4535
rect 1034 4534 1040 4535
rect 1043 4534 1072 4538
rect 962 4533 1072 4534
rect 962 4532 1078 4533
rect 637 4524 688 4532
rect 637 4512 662 4524
rect 669 4512 688 4524
rect 719 4524 769 4532
rect 719 4516 735 4524
rect 742 4522 769 4524
rect 778 4522 999 4532
rect 742 4512 999 4522
rect 1028 4524 1078 4532
rect 1028 4515 1044 4524
rect 637 4504 688 4512
rect 735 4504 999 4512
rect 1025 4512 1044 4515
rect 1051 4512 1078 4524
rect 1025 4504 1078 4512
rect 653 4496 654 4504
rect 669 4496 682 4504
rect 653 4488 669 4496
rect 650 4481 669 4484
rect 650 4472 672 4481
rect 623 4462 672 4472
rect 623 4456 653 4462
rect 672 4457 677 4462
rect 595 4440 669 4456
rect 687 4448 717 4504
rect 752 4494 960 4504
rect 995 4500 1040 4504
rect 1043 4503 1044 4504
rect 1059 4503 1072 4504
rect 778 4464 967 4494
rect 793 4461 967 4464
rect 786 4458 967 4461
rect 595 4438 608 4440
rect 623 4438 657 4440
rect 595 4422 669 4438
rect 696 4434 709 4448
rect 724 4434 740 4450
rect 786 4445 797 4458
rect 579 4400 580 4416
rect 595 4400 608 4422
rect 623 4400 653 4422
rect 696 4418 758 4434
rect 786 4427 797 4443
rect 802 4438 812 4458
rect 822 4438 836 4458
rect 839 4445 848 4458
rect 864 4445 873 4458
rect 802 4427 836 4438
rect 839 4427 848 4443
rect 864 4427 873 4443
rect 880 4438 890 4458
rect 900 4438 914 4458
rect 915 4445 926 4458
rect 880 4427 914 4438
rect 915 4427 926 4443
rect 972 4434 988 4450
rect 995 4448 1025 4500
rect 1059 4496 1060 4503
rect 1044 4488 1060 4496
rect 1031 4456 1044 4475
rect 1059 4456 1089 4472
rect 1031 4440 1105 4456
rect 1031 4438 1044 4440
rect 1059 4438 1093 4440
rect 696 4416 709 4418
rect 724 4416 758 4418
rect 696 4400 758 4416
rect 802 4411 818 4414
rect 880 4411 910 4422
rect 958 4418 1004 4434
rect 1031 4422 1105 4438
rect 958 4416 992 4418
rect 957 4400 1004 4416
rect 1031 4400 1044 4422
rect 1059 4400 1089 4422
rect 1116 4400 1117 4416
rect 1132 4400 1145 4560
rect 1175 4456 1188 4560
rect 1233 4538 1234 4548
rect 1249 4538 1262 4548
rect 1233 4534 1262 4538
rect 1267 4534 1297 4560
rect 1315 4546 1331 4548
rect 1403 4546 1456 4560
rect 1404 4544 1468 4546
rect 1511 4544 1526 4560
rect 1575 4557 1605 4560
rect 1575 4554 1611 4557
rect 1541 4546 1557 4548
rect 1315 4534 1330 4538
rect 1233 4532 1330 4534
rect 1358 4532 1526 4544
rect 1542 4534 1557 4538
rect 1575 4535 1614 4554
rect 1633 4548 1640 4549
rect 1639 4541 1640 4548
rect 1623 4538 1624 4541
rect 1639 4538 1652 4541
rect 1575 4534 1605 4535
rect 1614 4534 1620 4535
rect 1623 4534 1652 4538
rect 1542 4533 1652 4534
rect 1542 4532 1658 4533
rect 1217 4524 1268 4532
rect 1217 4512 1242 4524
rect 1249 4512 1268 4524
rect 1299 4524 1349 4532
rect 1299 4516 1315 4524
rect 1322 4522 1349 4524
rect 1358 4522 1579 4532
rect 1322 4512 1579 4522
rect 1608 4524 1658 4532
rect 1608 4515 1624 4524
rect 1217 4504 1268 4512
rect 1315 4504 1579 4512
rect 1605 4512 1624 4515
rect 1631 4512 1658 4524
rect 1605 4504 1658 4512
rect 1233 4496 1234 4504
rect 1249 4496 1262 4504
rect 1233 4488 1249 4496
rect 1230 4481 1249 4484
rect 1230 4472 1252 4481
rect 1203 4462 1252 4472
rect 1203 4456 1233 4462
rect 1252 4457 1257 4462
rect 1175 4440 1249 4456
rect 1267 4448 1297 4504
rect 1332 4494 1540 4504
rect 1575 4500 1620 4504
rect 1623 4503 1624 4504
rect 1639 4503 1652 4504
rect 1358 4464 1547 4494
rect 1373 4461 1547 4464
rect 1366 4458 1547 4461
rect 1175 4438 1188 4440
rect 1203 4438 1237 4440
rect 1175 4422 1249 4438
rect 1276 4434 1289 4448
rect 1304 4434 1320 4450
rect 1366 4445 1377 4458
rect 1159 4400 1160 4416
rect 1175 4400 1188 4422
rect 1203 4400 1233 4422
rect 1276 4418 1338 4434
rect 1366 4427 1377 4443
rect 1382 4438 1392 4458
rect 1402 4438 1416 4458
rect 1419 4445 1428 4458
rect 1444 4445 1453 4458
rect 1382 4427 1416 4438
rect 1419 4427 1428 4443
rect 1444 4427 1453 4443
rect 1460 4438 1470 4458
rect 1480 4438 1494 4458
rect 1495 4445 1506 4458
rect 1460 4427 1494 4438
rect 1495 4427 1506 4443
rect 1552 4434 1568 4450
rect 1575 4448 1605 4500
rect 1639 4496 1640 4503
rect 1624 4488 1640 4496
rect 1611 4456 1624 4475
rect 1639 4456 1669 4472
rect 1611 4440 1685 4456
rect 1611 4438 1624 4440
rect 1639 4438 1673 4440
rect 1276 4416 1289 4418
rect 1304 4416 1338 4418
rect 1276 4400 1338 4416
rect 1382 4411 1398 4414
rect 1460 4411 1490 4422
rect 1538 4418 1584 4434
rect 1611 4422 1685 4438
rect 1538 4416 1572 4418
rect 1537 4400 1584 4416
rect 1611 4400 1624 4422
rect 1639 4400 1669 4422
rect 1696 4400 1697 4416
rect 1712 4400 1725 4560
rect 1755 4456 1768 4560
rect 1813 4538 1814 4548
rect 1829 4538 1842 4548
rect 1813 4534 1842 4538
rect 1847 4534 1877 4560
rect 1895 4546 1911 4548
rect 1983 4546 2036 4560
rect 1984 4544 2048 4546
rect 2091 4544 2106 4560
rect 2155 4557 2185 4560
rect 2155 4554 2191 4557
rect 2121 4546 2137 4548
rect 1895 4534 1910 4538
rect 1813 4532 1910 4534
rect 1938 4532 2106 4544
rect 2122 4534 2137 4538
rect 2155 4535 2194 4554
rect 2213 4548 2220 4549
rect 2219 4541 2220 4548
rect 2203 4538 2204 4541
rect 2219 4538 2232 4541
rect 2155 4534 2185 4535
rect 2194 4534 2200 4535
rect 2203 4534 2232 4538
rect 2122 4533 2232 4534
rect 2122 4532 2238 4533
rect 1797 4524 1848 4532
rect 1797 4512 1822 4524
rect 1829 4512 1848 4524
rect 1879 4524 1929 4532
rect 1879 4516 1895 4524
rect 1902 4522 1929 4524
rect 1938 4522 2159 4532
rect 1902 4512 2159 4522
rect 2188 4524 2238 4532
rect 2188 4515 2204 4524
rect 1797 4504 1848 4512
rect 1895 4504 2159 4512
rect 2185 4512 2204 4515
rect 2211 4512 2238 4524
rect 2185 4504 2238 4512
rect 1813 4496 1814 4504
rect 1829 4496 1842 4504
rect 1813 4488 1829 4496
rect 1810 4481 1829 4484
rect 1810 4472 1832 4481
rect 1783 4462 1832 4472
rect 1783 4456 1813 4462
rect 1832 4457 1837 4462
rect 1755 4440 1829 4456
rect 1847 4448 1877 4504
rect 1912 4494 2120 4504
rect 2155 4500 2200 4504
rect 2203 4503 2204 4504
rect 2219 4503 2232 4504
rect 1938 4464 2127 4494
rect 1953 4461 2127 4464
rect 1946 4458 2127 4461
rect 1755 4438 1768 4440
rect 1783 4438 1817 4440
rect 1755 4422 1829 4438
rect 1856 4434 1869 4448
rect 1884 4434 1900 4450
rect 1946 4445 1957 4458
rect 1739 4400 1740 4416
rect 1755 4400 1768 4422
rect 1783 4400 1813 4422
rect 1856 4418 1918 4434
rect 1946 4427 1957 4443
rect 1962 4438 1972 4458
rect 1982 4438 1996 4458
rect 1999 4445 2008 4458
rect 2024 4445 2033 4458
rect 1962 4427 1996 4438
rect 1999 4427 2008 4443
rect 2024 4427 2033 4443
rect 2040 4438 2050 4458
rect 2060 4438 2074 4458
rect 2075 4445 2086 4458
rect 2040 4427 2074 4438
rect 2075 4427 2086 4443
rect 2132 4434 2148 4450
rect 2155 4448 2185 4500
rect 2219 4496 2220 4503
rect 2204 4488 2220 4496
rect 2191 4456 2204 4475
rect 2219 4456 2249 4472
rect 2191 4440 2265 4456
rect 2191 4438 2204 4440
rect 2219 4438 2253 4440
rect 1856 4416 1869 4418
rect 1884 4416 1918 4418
rect 1856 4400 1918 4416
rect 1962 4411 1978 4414
rect 2040 4411 2070 4422
rect 2118 4418 2164 4434
rect 2191 4422 2265 4438
rect 2118 4416 2152 4418
rect 2117 4400 2164 4416
rect 2191 4400 2204 4422
rect 2219 4400 2249 4422
rect 2276 4400 2277 4416
rect 2292 4400 2305 4560
rect 2335 4456 2348 4560
rect 2393 4538 2394 4548
rect 2409 4538 2422 4548
rect 2393 4534 2422 4538
rect 2427 4534 2457 4560
rect 2475 4546 2491 4548
rect 2563 4546 2616 4560
rect 2564 4544 2628 4546
rect 2671 4544 2686 4560
rect 2735 4557 2765 4560
rect 2735 4554 2771 4557
rect 2701 4546 2717 4548
rect 2475 4534 2490 4538
rect 2393 4532 2490 4534
rect 2518 4532 2686 4544
rect 2702 4534 2717 4538
rect 2735 4535 2774 4554
rect 2793 4548 2800 4549
rect 2799 4541 2800 4548
rect 2783 4538 2784 4541
rect 2799 4538 2812 4541
rect 2735 4534 2765 4535
rect 2774 4534 2780 4535
rect 2783 4534 2812 4538
rect 2702 4533 2812 4534
rect 2702 4532 2818 4533
rect 2377 4524 2428 4532
rect 2377 4512 2402 4524
rect 2409 4512 2428 4524
rect 2459 4524 2509 4532
rect 2459 4516 2475 4524
rect 2482 4522 2509 4524
rect 2518 4522 2739 4532
rect 2482 4512 2739 4522
rect 2768 4524 2818 4532
rect 2768 4515 2784 4524
rect 2377 4504 2428 4512
rect 2475 4504 2739 4512
rect 2765 4512 2784 4515
rect 2791 4512 2818 4524
rect 2765 4504 2818 4512
rect 2393 4496 2394 4504
rect 2409 4496 2422 4504
rect 2393 4488 2409 4496
rect 2390 4481 2409 4484
rect 2390 4472 2412 4481
rect 2363 4462 2412 4472
rect 2363 4456 2393 4462
rect 2412 4457 2417 4462
rect 2335 4440 2409 4456
rect 2427 4448 2457 4504
rect 2492 4494 2700 4504
rect 2735 4500 2780 4504
rect 2783 4503 2784 4504
rect 2799 4503 2812 4504
rect 2518 4464 2707 4494
rect 2533 4461 2707 4464
rect 2526 4458 2707 4461
rect 2335 4438 2348 4440
rect 2363 4438 2397 4440
rect 2335 4422 2409 4438
rect 2436 4434 2449 4448
rect 2464 4434 2480 4450
rect 2526 4445 2537 4458
rect 2319 4400 2320 4416
rect 2335 4400 2348 4422
rect 2363 4400 2393 4422
rect 2436 4418 2498 4434
rect 2526 4427 2537 4443
rect 2542 4438 2552 4458
rect 2562 4438 2576 4458
rect 2579 4445 2588 4458
rect 2604 4445 2613 4458
rect 2542 4427 2576 4438
rect 2579 4427 2588 4443
rect 2604 4427 2613 4443
rect 2620 4438 2630 4458
rect 2640 4438 2654 4458
rect 2655 4445 2666 4458
rect 2620 4427 2654 4438
rect 2655 4427 2666 4443
rect 2712 4434 2728 4450
rect 2735 4448 2765 4500
rect 2799 4496 2800 4503
rect 2784 4488 2800 4496
rect 2771 4456 2784 4475
rect 2799 4456 2829 4472
rect 2771 4440 2845 4456
rect 2771 4438 2784 4440
rect 2799 4438 2833 4440
rect 2436 4416 2449 4418
rect 2464 4416 2498 4418
rect 2436 4400 2498 4416
rect 2542 4411 2558 4414
rect 2620 4411 2650 4422
rect 2698 4418 2744 4434
rect 2771 4422 2845 4438
rect 2698 4416 2732 4418
rect 2697 4400 2744 4416
rect 2771 4400 2784 4422
rect 2799 4400 2829 4422
rect 2856 4400 2857 4416
rect 2872 4400 2885 4560
rect 2915 4456 2928 4560
rect 2973 4538 2974 4548
rect 2989 4538 3002 4548
rect 2973 4534 3002 4538
rect 3007 4534 3037 4560
rect 3055 4546 3071 4548
rect 3143 4546 3196 4560
rect 3144 4544 3208 4546
rect 3251 4544 3266 4560
rect 3315 4557 3345 4560
rect 3315 4554 3351 4557
rect 3281 4546 3297 4548
rect 3055 4534 3070 4538
rect 2973 4532 3070 4534
rect 3098 4532 3266 4544
rect 3282 4534 3297 4538
rect 3315 4535 3354 4554
rect 3373 4548 3380 4549
rect 3379 4541 3380 4548
rect 3363 4538 3364 4541
rect 3379 4538 3392 4541
rect 3315 4534 3345 4535
rect 3354 4534 3360 4535
rect 3363 4534 3392 4538
rect 3282 4533 3392 4534
rect 3282 4532 3398 4533
rect 2957 4524 3008 4532
rect 2957 4512 2982 4524
rect 2989 4512 3008 4524
rect 3039 4524 3089 4532
rect 3039 4516 3055 4524
rect 3062 4522 3089 4524
rect 3098 4522 3319 4532
rect 3062 4512 3319 4522
rect 3348 4524 3398 4532
rect 3348 4515 3364 4524
rect 2957 4504 3008 4512
rect 3055 4504 3319 4512
rect 3345 4512 3364 4515
rect 3371 4512 3398 4524
rect 3345 4504 3398 4512
rect 2973 4496 2974 4504
rect 2989 4496 3002 4504
rect 2973 4488 2989 4496
rect 2970 4481 2989 4484
rect 2970 4472 2992 4481
rect 2943 4462 2992 4472
rect 2943 4456 2973 4462
rect 2992 4457 2997 4462
rect 2915 4440 2989 4456
rect 3007 4448 3037 4504
rect 3072 4494 3280 4504
rect 3315 4500 3360 4504
rect 3363 4503 3364 4504
rect 3379 4503 3392 4504
rect 3098 4464 3287 4494
rect 3113 4461 3287 4464
rect 3106 4458 3287 4461
rect 2915 4438 2928 4440
rect 2943 4438 2977 4440
rect 2915 4422 2989 4438
rect 3016 4434 3029 4448
rect 3044 4434 3060 4450
rect 3106 4445 3117 4458
rect 2899 4400 2900 4416
rect 2915 4400 2928 4422
rect 2943 4400 2973 4422
rect 3016 4418 3078 4434
rect 3106 4427 3117 4443
rect 3122 4438 3132 4458
rect 3142 4438 3156 4458
rect 3159 4445 3168 4458
rect 3184 4445 3193 4458
rect 3122 4427 3156 4438
rect 3159 4427 3168 4443
rect 3184 4427 3193 4443
rect 3200 4438 3210 4458
rect 3220 4438 3234 4458
rect 3235 4445 3246 4458
rect 3200 4427 3234 4438
rect 3235 4427 3246 4443
rect 3292 4434 3308 4450
rect 3315 4448 3345 4500
rect 3379 4496 3380 4503
rect 3364 4488 3380 4496
rect 3351 4456 3364 4475
rect 3379 4456 3409 4472
rect 3351 4440 3425 4456
rect 3351 4438 3364 4440
rect 3379 4438 3413 4440
rect 3016 4416 3029 4418
rect 3044 4416 3078 4418
rect 3016 4400 3078 4416
rect 3122 4411 3138 4414
rect 3200 4411 3230 4422
rect 3278 4418 3324 4434
rect 3351 4422 3425 4438
rect 3278 4416 3312 4418
rect 3277 4400 3324 4416
rect 3351 4400 3364 4422
rect 3379 4400 3409 4422
rect 3436 4400 3437 4416
rect 3452 4400 3465 4560
rect 3495 4456 3508 4560
rect 3553 4538 3554 4548
rect 3569 4538 3582 4548
rect 3553 4534 3582 4538
rect 3587 4534 3617 4560
rect 3635 4546 3651 4548
rect 3723 4546 3776 4560
rect 3724 4544 3788 4546
rect 3831 4544 3846 4560
rect 3895 4557 3925 4560
rect 3895 4554 3931 4557
rect 3861 4546 3877 4548
rect 3635 4534 3650 4538
rect 3553 4532 3650 4534
rect 3678 4532 3846 4544
rect 3862 4534 3877 4538
rect 3895 4535 3934 4554
rect 3953 4548 3960 4549
rect 3959 4541 3960 4548
rect 3943 4538 3944 4541
rect 3959 4538 3972 4541
rect 3895 4534 3925 4535
rect 3934 4534 3940 4535
rect 3943 4534 3972 4538
rect 3862 4533 3972 4534
rect 3862 4532 3978 4533
rect 3537 4524 3588 4532
rect 3537 4512 3562 4524
rect 3569 4512 3588 4524
rect 3619 4524 3669 4532
rect 3619 4516 3635 4524
rect 3642 4522 3669 4524
rect 3678 4522 3899 4532
rect 3642 4512 3899 4522
rect 3928 4524 3978 4532
rect 3928 4515 3944 4524
rect 3537 4504 3588 4512
rect 3635 4504 3899 4512
rect 3925 4512 3944 4515
rect 3951 4512 3978 4524
rect 3925 4504 3978 4512
rect 3553 4496 3554 4504
rect 3569 4496 3582 4504
rect 3553 4488 3569 4496
rect 3550 4481 3569 4484
rect 3550 4472 3572 4481
rect 3523 4462 3572 4472
rect 3523 4456 3553 4462
rect 3572 4457 3577 4462
rect 3495 4440 3569 4456
rect 3587 4448 3617 4504
rect 3652 4494 3860 4504
rect 3895 4500 3940 4504
rect 3943 4503 3944 4504
rect 3959 4503 3972 4504
rect 3678 4464 3867 4494
rect 3693 4461 3867 4464
rect 3686 4458 3867 4461
rect 3495 4438 3508 4440
rect 3523 4438 3557 4440
rect 3495 4422 3569 4438
rect 3596 4434 3609 4448
rect 3624 4434 3640 4450
rect 3686 4445 3697 4458
rect 3479 4400 3480 4416
rect 3495 4400 3508 4422
rect 3523 4400 3553 4422
rect 3596 4418 3658 4434
rect 3686 4427 3697 4443
rect 3702 4438 3712 4458
rect 3722 4438 3736 4458
rect 3739 4445 3748 4458
rect 3764 4445 3773 4458
rect 3702 4427 3736 4438
rect 3739 4427 3748 4443
rect 3764 4427 3773 4443
rect 3780 4438 3790 4458
rect 3800 4438 3814 4458
rect 3815 4445 3826 4458
rect 3780 4427 3814 4438
rect 3815 4427 3826 4443
rect 3872 4434 3888 4450
rect 3895 4448 3925 4500
rect 3959 4496 3960 4503
rect 3944 4488 3960 4496
rect 3931 4456 3944 4475
rect 3959 4456 3989 4472
rect 3931 4440 4005 4456
rect 3931 4438 3944 4440
rect 3959 4438 3993 4440
rect 3596 4416 3609 4418
rect 3624 4416 3658 4418
rect 3596 4400 3658 4416
rect 3702 4411 3718 4414
rect 3780 4411 3810 4422
rect 3858 4418 3904 4434
rect 3931 4422 4005 4438
rect 3858 4416 3892 4418
rect 3857 4400 3904 4416
rect 3931 4400 3944 4422
rect 3959 4400 3989 4422
rect 4016 4400 4017 4416
rect 4032 4400 4045 4560
rect 4075 4456 4088 4560
rect 4133 4538 4134 4548
rect 4149 4538 4162 4548
rect 4133 4534 4162 4538
rect 4167 4534 4197 4560
rect 4215 4546 4231 4548
rect 4303 4546 4356 4560
rect 4304 4544 4368 4546
rect 4411 4544 4426 4560
rect 4475 4557 4505 4560
rect 4475 4554 4511 4557
rect 4441 4546 4457 4548
rect 4215 4534 4230 4538
rect 4133 4532 4230 4534
rect 4258 4532 4426 4544
rect 4442 4534 4457 4538
rect 4475 4535 4514 4554
rect 4533 4548 4540 4549
rect 4539 4541 4540 4548
rect 4523 4538 4524 4541
rect 4539 4538 4552 4541
rect 4475 4534 4505 4535
rect 4514 4534 4520 4535
rect 4523 4534 4552 4538
rect 4442 4533 4552 4534
rect 4442 4532 4558 4533
rect 4117 4524 4168 4532
rect 4117 4512 4142 4524
rect 4149 4512 4168 4524
rect 4199 4524 4249 4532
rect 4199 4516 4215 4524
rect 4222 4522 4249 4524
rect 4258 4522 4479 4532
rect 4222 4512 4479 4522
rect 4508 4524 4558 4532
rect 4508 4515 4524 4524
rect 4117 4504 4168 4512
rect 4215 4504 4479 4512
rect 4505 4512 4524 4515
rect 4531 4512 4558 4524
rect 4505 4504 4558 4512
rect 4133 4496 4134 4504
rect 4149 4496 4162 4504
rect 4133 4488 4149 4496
rect 4130 4481 4149 4484
rect 4130 4472 4152 4481
rect 4103 4462 4152 4472
rect 4103 4456 4133 4462
rect 4152 4457 4157 4462
rect 4075 4440 4149 4456
rect 4167 4448 4197 4504
rect 4232 4494 4440 4504
rect 4475 4500 4520 4504
rect 4523 4503 4524 4504
rect 4539 4503 4552 4504
rect 4258 4464 4447 4494
rect 4273 4461 4447 4464
rect 4266 4458 4447 4461
rect 4075 4438 4088 4440
rect 4103 4438 4137 4440
rect 4075 4422 4149 4438
rect 4176 4434 4189 4448
rect 4204 4434 4220 4450
rect 4266 4445 4277 4458
rect 4059 4400 4060 4416
rect 4075 4400 4088 4422
rect 4103 4400 4133 4422
rect 4176 4418 4238 4434
rect 4266 4427 4277 4443
rect 4282 4438 4292 4458
rect 4302 4438 4316 4458
rect 4319 4445 4328 4458
rect 4344 4445 4353 4458
rect 4282 4427 4316 4438
rect 4319 4427 4328 4443
rect 4344 4427 4353 4443
rect 4360 4438 4370 4458
rect 4380 4438 4394 4458
rect 4395 4445 4406 4458
rect 4360 4427 4394 4438
rect 4395 4427 4406 4443
rect 4452 4434 4468 4450
rect 4475 4448 4505 4500
rect 4539 4496 4540 4503
rect 4524 4488 4540 4496
rect 4511 4456 4524 4475
rect 4539 4456 4569 4472
rect 4511 4440 4585 4456
rect 4511 4438 4524 4440
rect 4539 4438 4573 4440
rect 4176 4416 4189 4418
rect 4204 4416 4238 4418
rect 4176 4400 4238 4416
rect 4282 4411 4298 4414
rect 4360 4411 4390 4422
rect 4438 4418 4484 4434
rect 4511 4422 4585 4438
rect 4438 4416 4472 4418
rect 4437 4400 4484 4416
rect 4511 4400 4524 4422
rect 4539 4400 4569 4422
rect 4596 4400 4597 4416
rect 4612 4400 4625 4560
rect -7 4392 34 4400
rect -7 4366 8 4392
rect 15 4366 34 4392
rect 98 4388 160 4400
rect 172 4388 247 4400
rect 305 4388 380 4400
rect 392 4388 423 4400
rect 429 4388 464 4400
rect 98 4386 260 4388
rect -7 4358 34 4366
rect 116 4362 129 4386
rect 144 4384 159 4386
rect -1 4348 0 4358
rect 15 4348 28 4358
rect 43 4348 73 4362
rect 116 4348 159 4362
rect 183 4359 190 4366
rect 193 4362 260 4386
rect 292 4386 464 4388
rect 262 4364 290 4368
rect 292 4364 372 4386
rect 393 4384 408 4386
rect 262 4362 372 4364
rect 193 4358 372 4362
rect 166 4348 196 4358
rect 198 4348 351 4358
rect 359 4348 389 4358
rect 393 4348 423 4362
rect 451 4348 464 4386
rect 536 4392 571 4400
rect 536 4366 537 4392
rect 544 4366 571 4392
rect 479 4348 509 4362
rect 536 4358 571 4366
rect 573 4392 614 4400
rect 573 4366 588 4392
rect 595 4366 614 4392
rect 678 4388 740 4400
rect 752 4388 827 4400
rect 885 4388 960 4400
rect 972 4388 1003 4400
rect 1009 4388 1044 4400
rect 678 4386 840 4388
rect 573 4358 614 4366
rect 696 4362 709 4386
rect 724 4384 739 4386
rect 536 4348 537 4358
rect 552 4348 565 4358
rect 579 4348 580 4358
rect 595 4348 608 4358
rect 623 4348 653 4362
rect 696 4348 739 4362
rect 763 4359 770 4366
rect 773 4362 840 4386
rect 872 4386 1044 4388
rect 842 4364 870 4368
rect 872 4364 952 4386
rect 973 4384 988 4386
rect 842 4362 952 4364
rect 773 4358 952 4362
rect 746 4348 776 4358
rect 778 4348 931 4358
rect 939 4348 969 4358
rect 973 4348 1003 4362
rect 1031 4348 1044 4386
rect 1116 4392 1151 4400
rect 1116 4366 1117 4392
rect 1124 4366 1151 4392
rect 1059 4348 1089 4362
rect 1116 4358 1151 4366
rect 1153 4392 1194 4400
rect 1153 4366 1168 4392
rect 1175 4366 1194 4392
rect 1258 4388 1320 4400
rect 1332 4388 1407 4400
rect 1465 4388 1540 4400
rect 1552 4388 1583 4400
rect 1589 4388 1624 4400
rect 1258 4386 1420 4388
rect 1153 4358 1194 4366
rect 1276 4362 1289 4386
rect 1304 4384 1319 4386
rect 1116 4348 1117 4358
rect 1132 4348 1145 4358
rect 1159 4348 1160 4358
rect 1175 4348 1188 4358
rect 1203 4348 1233 4362
rect 1276 4348 1319 4362
rect 1343 4359 1350 4366
rect 1353 4362 1420 4386
rect 1452 4386 1624 4388
rect 1422 4364 1450 4368
rect 1452 4364 1532 4386
rect 1553 4384 1568 4386
rect 1422 4362 1532 4364
rect 1353 4358 1532 4362
rect 1326 4348 1356 4358
rect 1358 4348 1511 4358
rect 1519 4348 1549 4358
rect 1553 4348 1583 4362
rect 1611 4348 1624 4386
rect 1696 4392 1731 4400
rect 1696 4366 1697 4392
rect 1704 4366 1731 4392
rect 1639 4348 1669 4362
rect 1696 4358 1731 4366
rect 1733 4392 1774 4400
rect 1733 4366 1748 4392
rect 1755 4366 1774 4392
rect 1838 4388 1900 4400
rect 1912 4388 1987 4400
rect 2045 4388 2120 4400
rect 2132 4388 2163 4400
rect 2169 4388 2204 4400
rect 1838 4386 2000 4388
rect 1733 4358 1774 4366
rect 1856 4362 1869 4386
rect 1884 4384 1899 4386
rect 1696 4348 1697 4358
rect 1712 4348 1725 4358
rect 1739 4348 1740 4358
rect 1755 4348 1768 4358
rect 1783 4348 1813 4362
rect 1856 4348 1899 4362
rect 1923 4359 1930 4366
rect 1933 4362 2000 4386
rect 2032 4386 2204 4388
rect 2002 4364 2030 4368
rect 2032 4364 2112 4386
rect 2133 4384 2148 4386
rect 2002 4362 2112 4364
rect 1933 4358 2112 4362
rect 1906 4348 1936 4358
rect 1938 4348 2091 4358
rect 2099 4348 2129 4358
rect 2133 4348 2163 4362
rect 2191 4348 2204 4386
rect 2276 4392 2311 4400
rect 2276 4366 2277 4392
rect 2284 4366 2311 4392
rect 2219 4348 2249 4362
rect 2276 4358 2311 4366
rect 2313 4392 2354 4400
rect 2313 4366 2328 4392
rect 2335 4366 2354 4392
rect 2418 4388 2480 4400
rect 2492 4388 2567 4400
rect 2625 4388 2700 4400
rect 2712 4388 2743 4400
rect 2749 4388 2784 4400
rect 2418 4386 2580 4388
rect 2313 4358 2354 4366
rect 2436 4362 2449 4386
rect 2464 4384 2479 4386
rect 2276 4348 2277 4358
rect 2292 4348 2305 4358
rect 2319 4348 2320 4358
rect 2335 4348 2348 4358
rect 2363 4348 2393 4362
rect 2436 4348 2479 4362
rect 2503 4359 2510 4366
rect 2513 4362 2580 4386
rect 2612 4386 2784 4388
rect 2582 4364 2610 4368
rect 2612 4364 2692 4386
rect 2713 4384 2728 4386
rect 2582 4362 2692 4364
rect 2513 4358 2692 4362
rect 2486 4348 2516 4358
rect 2518 4348 2671 4358
rect 2679 4348 2709 4358
rect 2713 4348 2743 4362
rect 2771 4348 2784 4386
rect 2856 4392 2891 4400
rect 2856 4366 2857 4392
rect 2864 4366 2891 4392
rect 2799 4348 2829 4362
rect 2856 4358 2891 4366
rect 2893 4392 2934 4400
rect 2893 4366 2908 4392
rect 2915 4366 2934 4392
rect 2998 4388 3060 4400
rect 3072 4388 3147 4400
rect 3205 4388 3280 4400
rect 3292 4388 3323 4400
rect 3329 4388 3364 4400
rect 2998 4386 3160 4388
rect 2893 4358 2934 4366
rect 3016 4362 3029 4386
rect 3044 4384 3059 4386
rect 2856 4348 2857 4358
rect 2872 4348 2885 4358
rect 2899 4348 2900 4358
rect 2915 4348 2928 4358
rect 2943 4348 2973 4362
rect 3016 4348 3059 4362
rect 3083 4359 3090 4366
rect 3093 4362 3160 4386
rect 3192 4386 3364 4388
rect 3162 4364 3190 4368
rect 3192 4364 3272 4386
rect 3293 4384 3308 4386
rect 3162 4362 3272 4364
rect 3093 4358 3272 4362
rect 3066 4348 3096 4358
rect 3098 4348 3251 4358
rect 3259 4348 3289 4358
rect 3293 4348 3323 4362
rect 3351 4348 3364 4386
rect 3436 4392 3471 4400
rect 3436 4366 3437 4392
rect 3444 4366 3471 4392
rect 3379 4348 3409 4362
rect 3436 4358 3471 4366
rect 3473 4392 3514 4400
rect 3473 4366 3488 4392
rect 3495 4366 3514 4392
rect 3578 4388 3640 4400
rect 3652 4388 3727 4400
rect 3785 4388 3860 4400
rect 3872 4388 3903 4400
rect 3909 4388 3944 4400
rect 3578 4386 3740 4388
rect 3473 4358 3514 4366
rect 3596 4362 3609 4386
rect 3624 4384 3639 4386
rect 3436 4348 3437 4358
rect 3452 4348 3465 4358
rect 3479 4348 3480 4358
rect 3495 4348 3508 4358
rect 3523 4348 3553 4362
rect 3596 4348 3639 4362
rect 3663 4359 3670 4366
rect 3673 4362 3740 4386
rect 3772 4386 3944 4388
rect 3742 4364 3770 4368
rect 3772 4364 3852 4386
rect 3873 4384 3888 4386
rect 3742 4362 3852 4364
rect 3673 4358 3852 4362
rect 3646 4348 3676 4358
rect 3678 4348 3831 4358
rect 3839 4348 3869 4358
rect 3873 4348 3903 4362
rect 3931 4348 3944 4386
rect 4016 4392 4051 4400
rect 4016 4366 4017 4392
rect 4024 4366 4051 4392
rect 3959 4348 3989 4362
rect 4016 4358 4051 4366
rect 4053 4392 4094 4400
rect 4053 4366 4068 4392
rect 4075 4366 4094 4392
rect 4158 4388 4220 4400
rect 4232 4388 4307 4400
rect 4365 4388 4440 4400
rect 4452 4388 4483 4400
rect 4489 4388 4524 4400
rect 4158 4386 4320 4388
rect 4053 4358 4094 4366
rect 4176 4362 4189 4386
rect 4204 4384 4219 4386
rect 4016 4348 4017 4358
rect 4032 4348 4045 4358
rect 4059 4348 4060 4358
rect 4075 4348 4088 4358
rect 4103 4348 4133 4362
rect 4176 4348 4219 4362
rect 4243 4359 4250 4366
rect 4253 4362 4320 4386
rect 4352 4386 4524 4388
rect 4322 4364 4350 4368
rect 4352 4364 4432 4386
rect 4453 4384 4468 4386
rect 4322 4362 4432 4364
rect 4253 4358 4432 4362
rect 4226 4348 4256 4358
rect 4258 4348 4411 4358
rect 4419 4348 4449 4358
rect 4453 4348 4483 4362
rect 4511 4348 4524 4386
rect 4596 4392 4631 4400
rect 4596 4366 4597 4392
rect 4604 4366 4631 4392
rect 4539 4348 4569 4362
rect 4596 4358 4631 4366
rect 4596 4348 4597 4358
rect 4612 4348 4625 4358
rect -1 4342 4625 4348
rect 0 4334 4625 4342
rect 15 4304 28 4334
rect 43 4316 73 4334
rect 116 4320 130 4334
rect 166 4320 386 4334
rect 117 4318 130 4320
rect 83 4306 98 4318
rect 80 4304 102 4306
rect 107 4304 137 4318
rect 198 4316 351 4320
rect 180 4304 372 4316
rect 415 4304 445 4318
rect 451 4304 464 4334
rect 479 4316 509 4334
rect 552 4304 565 4334
rect 595 4304 608 4334
rect 623 4316 653 4334
rect 696 4320 710 4334
rect 746 4320 966 4334
rect 697 4318 710 4320
rect 663 4306 678 4318
rect 660 4304 682 4306
rect 687 4304 717 4318
rect 778 4316 931 4320
rect 760 4304 952 4316
rect 995 4304 1025 4318
rect 1031 4304 1044 4334
rect 1059 4316 1089 4334
rect 1132 4304 1145 4334
rect 1175 4304 1188 4334
rect 1203 4316 1233 4334
rect 1276 4320 1290 4334
rect 1326 4320 1546 4334
rect 1277 4318 1290 4320
rect 1243 4306 1258 4318
rect 1240 4304 1262 4306
rect 1267 4304 1297 4318
rect 1358 4316 1511 4320
rect 1340 4304 1532 4316
rect 1575 4304 1605 4318
rect 1611 4304 1624 4334
rect 1639 4316 1669 4334
rect 1712 4304 1725 4334
rect 1755 4304 1768 4334
rect 1783 4316 1813 4334
rect 1856 4320 1870 4334
rect 1906 4320 2126 4334
rect 1857 4318 1870 4320
rect 1823 4306 1838 4318
rect 1820 4304 1842 4306
rect 1847 4304 1877 4318
rect 1938 4316 2091 4320
rect 1920 4304 2112 4316
rect 2155 4304 2185 4318
rect 2191 4304 2204 4334
rect 2219 4316 2249 4334
rect 2292 4304 2305 4334
rect 2335 4304 2348 4334
rect 2363 4316 2393 4334
rect 2436 4320 2450 4334
rect 2486 4320 2706 4334
rect 2437 4318 2450 4320
rect 2403 4306 2418 4318
rect 2400 4304 2422 4306
rect 2427 4304 2457 4318
rect 2518 4316 2671 4320
rect 2500 4304 2692 4316
rect 2735 4304 2765 4318
rect 2771 4304 2784 4334
rect 2799 4316 2829 4334
rect 2872 4304 2885 4334
rect 2915 4304 2928 4334
rect 2943 4316 2973 4334
rect 3016 4320 3030 4334
rect 3066 4320 3286 4334
rect 3017 4318 3030 4320
rect 2983 4306 2998 4318
rect 2980 4304 3002 4306
rect 3007 4304 3037 4318
rect 3098 4316 3251 4320
rect 3080 4304 3272 4316
rect 3315 4304 3345 4318
rect 3351 4304 3364 4334
rect 3379 4316 3409 4334
rect 3452 4304 3465 4334
rect 3495 4304 3508 4334
rect 3523 4316 3553 4334
rect 3596 4320 3610 4334
rect 3646 4320 3866 4334
rect 3597 4318 3610 4320
rect 3563 4306 3578 4318
rect 3560 4304 3582 4306
rect 3587 4304 3617 4318
rect 3678 4316 3831 4320
rect 3660 4304 3852 4316
rect 3895 4304 3925 4318
rect 3931 4304 3944 4334
rect 3959 4316 3989 4334
rect 4032 4304 4045 4334
rect 4075 4304 4088 4334
rect 4103 4316 4133 4334
rect 4176 4320 4190 4334
rect 4226 4320 4446 4334
rect 4177 4318 4190 4320
rect 4143 4306 4158 4318
rect 4140 4304 4162 4306
rect 4167 4304 4197 4318
rect 4258 4316 4411 4320
rect 4240 4304 4432 4316
rect 4475 4304 4505 4318
rect 4511 4304 4524 4334
rect 4539 4316 4569 4334
rect 4612 4304 4625 4334
rect 0 4290 4625 4304
rect 15 4186 28 4290
rect 73 4268 74 4278
rect 89 4268 102 4278
rect 73 4264 102 4268
rect 107 4264 137 4290
rect 155 4276 171 4278
rect 243 4276 296 4290
rect 244 4274 308 4276
rect 351 4274 366 4290
rect 415 4287 445 4290
rect 415 4284 451 4287
rect 381 4276 397 4278
rect 155 4264 170 4268
rect 73 4262 170 4264
rect 198 4262 366 4274
rect 382 4264 397 4268
rect 415 4265 454 4284
rect 473 4278 480 4279
rect 479 4271 480 4278
rect 463 4268 464 4271
rect 479 4268 492 4271
rect 415 4264 445 4265
rect 454 4264 460 4265
rect 463 4264 492 4268
rect 382 4263 492 4264
rect 382 4262 498 4263
rect 57 4254 108 4262
rect 57 4242 82 4254
rect 89 4242 108 4254
rect 139 4254 189 4262
rect 139 4246 155 4254
rect 162 4252 189 4254
rect 198 4252 419 4262
rect 162 4242 419 4252
rect 448 4254 498 4262
rect 448 4245 464 4254
rect 57 4234 108 4242
rect 155 4234 419 4242
rect 445 4242 464 4245
rect 471 4242 498 4254
rect 445 4234 498 4242
rect 73 4226 74 4234
rect 89 4226 102 4234
rect 73 4218 89 4226
rect 70 4211 89 4214
rect 70 4202 92 4211
rect 43 4192 92 4202
rect 43 4186 73 4192
rect 92 4187 97 4192
rect 15 4170 89 4186
rect 107 4178 137 4234
rect 172 4224 380 4234
rect 415 4230 460 4234
rect 463 4233 464 4234
rect 479 4233 492 4234
rect 198 4194 387 4224
rect 213 4191 387 4194
rect 206 4188 387 4191
rect 15 4168 28 4170
rect 43 4168 77 4170
rect 15 4152 89 4168
rect 116 4164 129 4178
rect 144 4164 160 4180
rect 206 4175 217 4188
rect -1 4130 0 4146
rect 15 4130 28 4152
rect 43 4130 73 4152
rect 116 4148 178 4164
rect 206 4157 217 4173
rect 222 4168 232 4188
rect 242 4168 256 4188
rect 259 4175 268 4188
rect 284 4175 293 4188
rect 222 4157 256 4168
rect 259 4157 268 4173
rect 284 4157 293 4173
rect 300 4168 310 4188
rect 320 4168 334 4188
rect 335 4175 346 4188
rect 300 4157 334 4168
rect 335 4157 346 4173
rect 392 4164 408 4180
rect 415 4178 445 4230
rect 479 4226 480 4233
rect 464 4218 480 4226
rect 451 4186 464 4205
rect 479 4186 509 4202
rect 451 4170 525 4186
rect 451 4168 464 4170
rect 479 4168 513 4170
rect 116 4146 129 4148
rect 144 4146 178 4148
rect 116 4130 178 4146
rect 222 4141 238 4144
rect 300 4141 330 4152
rect 378 4148 424 4164
rect 451 4152 525 4168
rect 378 4146 412 4148
rect 377 4130 424 4146
rect 451 4130 464 4152
rect 479 4130 509 4152
rect 536 4130 537 4146
rect 552 4130 565 4290
rect 595 4186 608 4290
rect 653 4268 654 4278
rect 669 4268 682 4278
rect 653 4264 682 4268
rect 687 4264 717 4290
rect 735 4276 751 4278
rect 823 4276 876 4290
rect 824 4274 888 4276
rect 931 4274 946 4290
rect 995 4287 1025 4290
rect 995 4284 1031 4287
rect 961 4276 977 4278
rect 735 4264 750 4268
rect 653 4262 750 4264
rect 778 4262 946 4274
rect 962 4264 977 4268
rect 995 4265 1034 4284
rect 1053 4278 1060 4279
rect 1059 4271 1060 4278
rect 1043 4268 1044 4271
rect 1059 4268 1072 4271
rect 995 4264 1025 4265
rect 1034 4264 1040 4265
rect 1043 4264 1072 4268
rect 962 4263 1072 4264
rect 962 4262 1078 4263
rect 637 4254 688 4262
rect 637 4242 662 4254
rect 669 4242 688 4254
rect 719 4254 769 4262
rect 719 4246 735 4254
rect 742 4252 769 4254
rect 778 4252 999 4262
rect 742 4242 999 4252
rect 1028 4254 1078 4262
rect 1028 4245 1044 4254
rect 637 4234 688 4242
rect 735 4234 999 4242
rect 1025 4242 1044 4245
rect 1051 4242 1078 4254
rect 1025 4234 1078 4242
rect 653 4226 654 4234
rect 669 4226 682 4234
rect 653 4218 669 4226
rect 650 4211 669 4214
rect 650 4202 672 4211
rect 623 4192 672 4202
rect 623 4186 653 4192
rect 672 4187 677 4192
rect 595 4170 669 4186
rect 687 4178 717 4234
rect 752 4224 960 4234
rect 995 4230 1040 4234
rect 1043 4233 1044 4234
rect 1059 4233 1072 4234
rect 778 4194 967 4224
rect 793 4191 967 4194
rect 786 4188 967 4191
rect 595 4168 608 4170
rect 623 4168 657 4170
rect 595 4152 669 4168
rect 696 4164 709 4178
rect 724 4164 740 4180
rect 786 4175 797 4188
rect 579 4130 580 4146
rect 595 4130 608 4152
rect 623 4130 653 4152
rect 696 4148 758 4164
rect 786 4157 797 4173
rect 802 4168 812 4188
rect 822 4168 836 4188
rect 839 4175 848 4188
rect 864 4175 873 4188
rect 802 4157 836 4168
rect 839 4157 848 4173
rect 864 4157 873 4173
rect 880 4168 890 4188
rect 900 4168 914 4188
rect 915 4175 926 4188
rect 880 4157 914 4168
rect 915 4157 926 4173
rect 972 4164 988 4180
rect 995 4178 1025 4230
rect 1059 4226 1060 4233
rect 1044 4218 1060 4226
rect 1031 4186 1044 4205
rect 1059 4186 1089 4202
rect 1031 4170 1105 4186
rect 1031 4168 1044 4170
rect 1059 4168 1093 4170
rect 696 4146 709 4148
rect 724 4146 758 4148
rect 696 4130 758 4146
rect 802 4141 818 4144
rect 880 4141 910 4152
rect 958 4148 1004 4164
rect 1031 4152 1105 4168
rect 958 4146 992 4148
rect 957 4130 1004 4146
rect 1031 4130 1044 4152
rect 1059 4130 1089 4152
rect 1116 4130 1117 4146
rect 1132 4130 1145 4290
rect 1175 4186 1188 4290
rect 1233 4268 1234 4278
rect 1249 4268 1262 4278
rect 1233 4264 1262 4268
rect 1267 4264 1297 4290
rect 1315 4276 1331 4278
rect 1403 4276 1456 4290
rect 1404 4274 1468 4276
rect 1511 4274 1526 4290
rect 1575 4287 1605 4290
rect 1575 4284 1611 4287
rect 1541 4276 1557 4278
rect 1315 4264 1330 4268
rect 1233 4262 1330 4264
rect 1358 4262 1526 4274
rect 1542 4264 1557 4268
rect 1575 4265 1614 4284
rect 1633 4278 1640 4279
rect 1639 4271 1640 4278
rect 1623 4268 1624 4271
rect 1639 4268 1652 4271
rect 1575 4264 1605 4265
rect 1614 4264 1620 4265
rect 1623 4264 1652 4268
rect 1542 4263 1652 4264
rect 1542 4262 1658 4263
rect 1217 4254 1268 4262
rect 1217 4242 1242 4254
rect 1249 4242 1268 4254
rect 1299 4254 1349 4262
rect 1299 4246 1315 4254
rect 1322 4252 1349 4254
rect 1358 4252 1579 4262
rect 1322 4242 1579 4252
rect 1608 4254 1658 4262
rect 1608 4245 1624 4254
rect 1217 4234 1268 4242
rect 1315 4234 1579 4242
rect 1605 4242 1624 4245
rect 1631 4242 1658 4254
rect 1605 4234 1658 4242
rect 1233 4226 1234 4234
rect 1249 4226 1262 4234
rect 1233 4218 1249 4226
rect 1230 4211 1249 4214
rect 1230 4202 1252 4211
rect 1203 4192 1252 4202
rect 1203 4186 1233 4192
rect 1252 4187 1257 4192
rect 1175 4170 1249 4186
rect 1267 4178 1297 4234
rect 1332 4224 1540 4234
rect 1575 4230 1620 4234
rect 1623 4233 1624 4234
rect 1639 4233 1652 4234
rect 1358 4194 1547 4224
rect 1373 4191 1547 4194
rect 1366 4188 1547 4191
rect 1175 4168 1188 4170
rect 1203 4168 1237 4170
rect 1175 4152 1249 4168
rect 1276 4164 1289 4178
rect 1304 4164 1320 4180
rect 1366 4175 1377 4188
rect 1159 4130 1160 4146
rect 1175 4130 1188 4152
rect 1203 4130 1233 4152
rect 1276 4148 1338 4164
rect 1366 4157 1377 4173
rect 1382 4168 1392 4188
rect 1402 4168 1416 4188
rect 1419 4175 1428 4188
rect 1444 4175 1453 4188
rect 1382 4157 1416 4168
rect 1419 4157 1428 4173
rect 1444 4157 1453 4173
rect 1460 4168 1470 4188
rect 1480 4168 1494 4188
rect 1495 4175 1506 4188
rect 1460 4157 1494 4168
rect 1495 4157 1506 4173
rect 1552 4164 1568 4180
rect 1575 4178 1605 4230
rect 1639 4226 1640 4233
rect 1624 4218 1640 4226
rect 1611 4186 1624 4205
rect 1639 4186 1669 4202
rect 1611 4170 1685 4186
rect 1611 4168 1624 4170
rect 1639 4168 1673 4170
rect 1276 4146 1289 4148
rect 1304 4146 1338 4148
rect 1276 4130 1338 4146
rect 1382 4141 1398 4144
rect 1460 4141 1490 4152
rect 1538 4148 1584 4164
rect 1611 4152 1685 4168
rect 1538 4146 1572 4148
rect 1537 4130 1584 4146
rect 1611 4130 1624 4152
rect 1639 4130 1669 4152
rect 1696 4130 1697 4146
rect 1712 4130 1725 4290
rect 1755 4186 1768 4290
rect 1813 4268 1814 4278
rect 1829 4268 1842 4278
rect 1813 4264 1842 4268
rect 1847 4264 1877 4290
rect 1895 4276 1911 4278
rect 1983 4276 2036 4290
rect 1984 4274 2048 4276
rect 2091 4274 2106 4290
rect 2155 4287 2185 4290
rect 2155 4284 2191 4287
rect 2121 4276 2137 4278
rect 1895 4264 1910 4268
rect 1813 4262 1910 4264
rect 1938 4262 2106 4274
rect 2122 4264 2137 4268
rect 2155 4265 2194 4284
rect 2213 4278 2220 4279
rect 2219 4271 2220 4278
rect 2203 4268 2204 4271
rect 2219 4268 2232 4271
rect 2155 4264 2185 4265
rect 2194 4264 2200 4265
rect 2203 4264 2232 4268
rect 2122 4263 2232 4264
rect 2122 4262 2238 4263
rect 1797 4254 1848 4262
rect 1797 4242 1822 4254
rect 1829 4242 1848 4254
rect 1879 4254 1929 4262
rect 1879 4246 1895 4254
rect 1902 4252 1929 4254
rect 1938 4252 2159 4262
rect 1902 4242 2159 4252
rect 2188 4254 2238 4262
rect 2188 4245 2204 4254
rect 1797 4234 1848 4242
rect 1895 4234 2159 4242
rect 2185 4242 2204 4245
rect 2211 4242 2238 4254
rect 2185 4234 2238 4242
rect 1813 4226 1814 4234
rect 1829 4226 1842 4234
rect 1813 4218 1829 4226
rect 1810 4211 1829 4214
rect 1810 4202 1832 4211
rect 1783 4192 1832 4202
rect 1783 4186 1813 4192
rect 1832 4187 1837 4192
rect 1755 4170 1829 4186
rect 1847 4178 1877 4234
rect 1912 4224 2120 4234
rect 2155 4230 2200 4234
rect 2203 4233 2204 4234
rect 2219 4233 2232 4234
rect 1938 4194 2127 4224
rect 1953 4191 2127 4194
rect 1946 4188 2127 4191
rect 1755 4168 1768 4170
rect 1783 4168 1817 4170
rect 1755 4152 1829 4168
rect 1856 4164 1869 4178
rect 1884 4164 1900 4180
rect 1946 4175 1957 4188
rect 1739 4130 1740 4146
rect 1755 4130 1768 4152
rect 1783 4130 1813 4152
rect 1856 4148 1918 4164
rect 1946 4157 1957 4173
rect 1962 4168 1972 4188
rect 1982 4168 1996 4188
rect 1999 4175 2008 4188
rect 2024 4175 2033 4188
rect 1962 4157 1996 4168
rect 1999 4157 2008 4173
rect 2024 4157 2033 4173
rect 2040 4168 2050 4188
rect 2060 4168 2074 4188
rect 2075 4175 2086 4188
rect 2040 4157 2074 4168
rect 2075 4157 2086 4173
rect 2132 4164 2148 4180
rect 2155 4178 2185 4230
rect 2219 4226 2220 4233
rect 2204 4218 2220 4226
rect 2191 4186 2204 4205
rect 2219 4186 2249 4202
rect 2191 4170 2265 4186
rect 2191 4168 2204 4170
rect 2219 4168 2253 4170
rect 1856 4146 1869 4148
rect 1884 4146 1918 4148
rect 1856 4130 1918 4146
rect 1962 4141 1978 4144
rect 2040 4141 2070 4152
rect 2118 4148 2164 4164
rect 2191 4152 2265 4168
rect 2118 4146 2152 4148
rect 2117 4130 2164 4146
rect 2191 4130 2204 4152
rect 2219 4130 2249 4152
rect 2276 4130 2277 4146
rect 2292 4130 2305 4290
rect 2335 4186 2348 4290
rect 2393 4268 2394 4278
rect 2409 4268 2422 4278
rect 2393 4264 2422 4268
rect 2427 4264 2457 4290
rect 2475 4276 2491 4278
rect 2563 4276 2616 4290
rect 2564 4274 2628 4276
rect 2671 4274 2686 4290
rect 2735 4287 2765 4290
rect 2735 4284 2771 4287
rect 2701 4276 2717 4278
rect 2475 4264 2490 4268
rect 2393 4262 2490 4264
rect 2518 4262 2686 4274
rect 2702 4264 2717 4268
rect 2735 4265 2774 4284
rect 2793 4278 2800 4279
rect 2799 4271 2800 4278
rect 2783 4268 2784 4271
rect 2799 4268 2812 4271
rect 2735 4264 2765 4265
rect 2774 4264 2780 4265
rect 2783 4264 2812 4268
rect 2702 4263 2812 4264
rect 2702 4262 2818 4263
rect 2377 4254 2428 4262
rect 2377 4242 2402 4254
rect 2409 4242 2428 4254
rect 2459 4254 2509 4262
rect 2459 4246 2475 4254
rect 2482 4252 2509 4254
rect 2518 4252 2739 4262
rect 2482 4242 2739 4252
rect 2768 4254 2818 4262
rect 2768 4245 2784 4254
rect 2377 4234 2428 4242
rect 2475 4234 2739 4242
rect 2765 4242 2784 4245
rect 2791 4242 2818 4254
rect 2765 4234 2818 4242
rect 2393 4226 2394 4234
rect 2409 4226 2422 4234
rect 2393 4218 2409 4226
rect 2390 4211 2409 4214
rect 2390 4202 2412 4211
rect 2363 4192 2412 4202
rect 2363 4186 2393 4192
rect 2412 4187 2417 4192
rect 2335 4170 2409 4186
rect 2427 4178 2457 4234
rect 2492 4224 2700 4234
rect 2735 4230 2780 4234
rect 2783 4233 2784 4234
rect 2799 4233 2812 4234
rect 2518 4194 2707 4224
rect 2533 4191 2707 4194
rect 2526 4188 2707 4191
rect 2335 4168 2348 4170
rect 2363 4168 2397 4170
rect 2335 4152 2409 4168
rect 2436 4164 2449 4178
rect 2464 4164 2480 4180
rect 2526 4175 2537 4188
rect 2319 4130 2320 4146
rect 2335 4130 2348 4152
rect 2363 4130 2393 4152
rect 2436 4148 2498 4164
rect 2526 4157 2537 4173
rect 2542 4168 2552 4188
rect 2562 4168 2576 4188
rect 2579 4175 2588 4188
rect 2604 4175 2613 4188
rect 2542 4157 2576 4168
rect 2579 4157 2588 4173
rect 2604 4157 2613 4173
rect 2620 4168 2630 4188
rect 2640 4168 2654 4188
rect 2655 4175 2666 4188
rect 2620 4157 2654 4168
rect 2655 4157 2666 4173
rect 2712 4164 2728 4180
rect 2735 4178 2765 4230
rect 2799 4226 2800 4233
rect 2784 4218 2800 4226
rect 2771 4186 2784 4205
rect 2799 4186 2829 4202
rect 2771 4170 2845 4186
rect 2771 4168 2784 4170
rect 2799 4168 2833 4170
rect 2436 4146 2449 4148
rect 2464 4146 2498 4148
rect 2436 4130 2498 4146
rect 2542 4141 2558 4144
rect 2620 4141 2650 4152
rect 2698 4148 2744 4164
rect 2771 4152 2845 4168
rect 2698 4146 2732 4148
rect 2697 4130 2744 4146
rect 2771 4130 2784 4152
rect 2799 4130 2829 4152
rect 2856 4130 2857 4146
rect 2872 4130 2885 4290
rect 2915 4186 2928 4290
rect 2973 4268 2974 4278
rect 2989 4268 3002 4278
rect 2973 4264 3002 4268
rect 3007 4264 3037 4290
rect 3055 4276 3071 4278
rect 3143 4276 3196 4290
rect 3144 4274 3208 4276
rect 3251 4274 3266 4290
rect 3315 4287 3345 4290
rect 3315 4284 3351 4287
rect 3281 4276 3297 4278
rect 3055 4264 3070 4268
rect 2973 4262 3070 4264
rect 3098 4262 3266 4274
rect 3282 4264 3297 4268
rect 3315 4265 3354 4284
rect 3373 4278 3380 4279
rect 3379 4271 3380 4278
rect 3363 4268 3364 4271
rect 3379 4268 3392 4271
rect 3315 4264 3345 4265
rect 3354 4264 3360 4265
rect 3363 4264 3392 4268
rect 3282 4263 3392 4264
rect 3282 4262 3398 4263
rect 2957 4254 3008 4262
rect 2957 4242 2982 4254
rect 2989 4242 3008 4254
rect 3039 4254 3089 4262
rect 3039 4246 3055 4254
rect 3062 4252 3089 4254
rect 3098 4252 3319 4262
rect 3062 4242 3319 4252
rect 3348 4254 3398 4262
rect 3348 4245 3364 4254
rect 2957 4234 3008 4242
rect 3055 4234 3319 4242
rect 3345 4242 3364 4245
rect 3371 4242 3398 4254
rect 3345 4234 3398 4242
rect 2973 4226 2974 4234
rect 2989 4226 3002 4234
rect 2973 4218 2989 4226
rect 2970 4211 2989 4214
rect 2970 4202 2992 4211
rect 2943 4192 2992 4202
rect 2943 4186 2973 4192
rect 2992 4187 2997 4192
rect 2915 4170 2989 4186
rect 3007 4178 3037 4234
rect 3072 4224 3280 4234
rect 3315 4230 3360 4234
rect 3363 4233 3364 4234
rect 3379 4233 3392 4234
rect 3098 4194 3287 4224
rect 3113 4191 3287 4194
rect 3106 4188 3287 4191
rect 2915 4168 2928 4170
rect 2943 4168 2977 4170
rect 2915 4152 2989 4168
rect 3016 4164 3029 4178
rect 3044 4164 3060 4180
rect 3106 4175 3117 4188
rect 2899 4130 2900 4146
rect 2915 4130 2928 4152
rect 2943 4130 2973 4152
rect 3016 4148 3078 4164
rect 3106 4157 3117 4173
rect 3122 4168 3132 4188
rect 3142 4168 3156 4188
rect 3159 4175 3168 4188
rect 3184 4175 3193 4188
rect 3122 4157 3156 4168
rect 3159 4157 3168 4173
rect 3184 4157 3193 4173
rect 3200 4168 3210 4188
rect 3220 4168 3234 4188
rect 3235 4175 3246 4188
rect 3200 4157 3234 4168
rect 3235 4157 3246 4173
rect 3292 4164 3308 4180
rect 3315 4178 3345 4230
rect 3379 4226 3380 4233
rect 3364 4218 3380 4226
rect 3351 4186 3364 4205
rect 3379 4186 3409 4202
rect 3351 4170 3425 4186
rect 3351 4168 3364 4170
rect 3379 4168 3413 4170
rect 3016 4146 3029 4148
rect 3044 4146 3078 4148
rect 3016 4130 3078 4146
rect 3122 4141 3138 4144
rect 3200 4141 3230 4152
rect 3278 4148 3324 4164
rect 3351 4152 3425 4168
rect 3278 4146 3312 4148
rect 3277 4130 3324 4146
rect 3351 4130 3364 4152
rect 3379 4130 3409 4152
rect 3436 4130 3437 4146
rect 3452 4130 3465 4290
rect 3495 4186 3508 4290
rect 3553 4268 3554 4278
rect 3569 4268 3582 4278
rect 3553 4264 3582 4268
rect 3587 4264 3617 4290
rect 3635 4276 3651 4278
rect 3723 4276 3776 4290
rect 3724 4274 3788 4276
rect 3831 4274 3846 4290
rect 3895 4287 3925 4290
rect 3895 4284 3931 4287
rect 3861 4276 3877 4278
rect 3635 4264 3650 4268
rect 3553 4262 3650 4264
rect 3678 4262 3846 4274
rect 3862 4264 3877 4268
rect 3895 4265 3934 4284
rect 3953 4278 3960 4279
rect 3959 4271 3960 4278
rect 3943 4268 3944 4271
rect 3959 4268 3972 4271
rect 3895 4264 3925 4265
rect 3934 4264 3940 4265
rect 3943 4264 3972 4268
rect 3862 4263 3972 4264
rect 3862 4262 3978 4263
rect 3537 4254 3588 4262
rect 3537 4242 3562 4254
rect 3569 4242 3588 4254
rect 3619 4254 3669 4262
rect 3619 4246 3635 4254
rect 3642 4252 3669 4254
rect 3678 4252 3899 4262
rect 3642 4242 3899 4252
rect 3928 4254 3978 4262
rect 3928 4245 3944 4254
rect 3537 4234 3588 4242
rect 3635 4234 3899 4242
rect 3925 4242 3944 4245
rect 3951 4242 3978 4254
rect 3925 4234 3978 4242
rect 3553 4226 3554 4234
rect 3569 4226 3582 4234
rect 3553 4218 3569 4226
rect 3550 4211 3569 4214
rect 3550 4202 3572 4211
rect 3523 4192 3572 4202
rect 3523 4186 3553 4192
rect 3572 4187 3577 4192
rect 3495 4170 3569 4186
rect 3587 4178 3617 4234
rect 3652 4224 3860 4234
rect 3895 4230 3940 4234
rect 3943 4233 3944 4234
rect 3959 4233 3972 4234
rect 3678 4194 3867 4224
rect 3693 4191 3867 4194
rect 3686 4188 3867 4191
rect 3495 4168 3508 4170
rect 3523 4168 3557 4170
rect 3495 4152 3569 4168
rect 3596 4164 3609 4178
rect 3624 4164 3640 4180
rect 3686 4175 3697 4188
rect 3479 4130 3480 4146
rect 3495 4130 3508 4152
rect 3523 4130 3553 4152
rect 3596 4148 3658 4164
rect 3686 4157 3697 4173
rect 3702 4168 3712 4188
rect 3722 4168 3736 4188
rect 3739 4175 3748 4188
rect 3764 4175 3773 4188
rect 3702 4157 3736 4168
rect 3739 4157 3748 4173
rect 3764 4157 3773 4173
rect 3780 4168 3790 4188
rect 3800 4168 3814 4188
rect 3815 4175 3826 4188
rect 3780 4157 3814 4168
rect 3815 4157 3826 4173
rect 3872 4164 3888 4180
rect 3895 4178 3925 4230
rect 3959 4226 3960 4233
rect 3944 4218 3960 4226
rect 3931 4186 3944 4205
rect 3959 4186 3989 4202
rect 3931 4170 4005 4186
rect 3931 4168 3944 4170
rect 3959 4168 3993 4170
rect 3596 4146 3609 4148
rect 3624 4146 3658 4148
rect 3596 4130 3658 4146
rect 3702 4141 3718 4144
rect 3780 4141 3810 4152
rect 3858 4148 3904 4164
rect 3931 4152 4005 4168
rect 3858 4146 3892 4148
rect 3857 4130 3904 4146
rect 3931 4130 3944 4152
rect 3959 4130 3989 4152
rect 4016 4130 4017 4146
rect 4032 4130 4045 4290
rect 4075 4186 4088 4290
rect 4133 4268 4134 4278
rect 4149 4268 4162 4278
rect 4133 4264 4162 4268
rect 4167 4264 4197 4290
rect 4215 4276 4231 4278
rect 4303 4276 4356 4290
rect 4304 4274 4368 4276
rect 4411 4274 4426 4290
rect 4475 4287 4505 4290
rect 4475 4284 4511 4287
rect 4441 4276 4457 4278
rect 4215 4264 4230 4268
rect 4133 4262 4230 4264
rect 4258 4262 4426 4274
rect 4442 4264 4457 4268
rect 4475 4265 4514 4284
rect 4533 4278 4540 4279
rect 4539 4271 4540 4278
rect 4523 4268 4524 4271
rect 4539 4268 4552 4271
rect 4475 4264 4505 4265
rect 4514 4264 4520 4265
rect 4523 4264 4552 4268
rect 4442 4263 4552 4264
rect 4442 4262 4558 4263
rect 4117 4254 4168 4262
rect 4117 4242 4142 4254
rect 4149 4242 4168 4254
rect 4199 4254 4249 4262
rect 4199 4246 4215 4254
rect 4222 4252 4249 4254
rect 4258 4252 4479 4262
rect 4222 4242 4479 4252
rect 4508 4254 4558 4262
rect 4508 4245 4524 4254
rect 4117 4234 4168 4242
rect 4215 4234 4479 4242
rect 4505 4242 4524 4245
rect 4531 4242 4558 4254
rect 4505 4234 4558 4242
rect 4133 4226 4134 4234
rect 4149 4226 4162 4234
rect 4133 4218 4149 4226
rect 4130 4211 4149 4214
rect 4130 4202 4152 4211
rect 4103 4192 4152 4202
rect 4103 4186 4133 4192
rect 4152 4187 4157 4192
rect 4075 4170 4149 4186
rect 4167 4178 4197 4234
rect 4232 4224 4440 4234
rect 4475 4230 4520 4234
rect 4523 4233 4524 4234
rect 4539 4233 4552 4234
rect 4258 4194 4447 4224
rect 4273 4191 4447 4194
rect 4266 4188 4447 4191
rect 4075 4168 4088 4170
rect 4103 4168 4137 4170
rect 4075 4152 4149 4168
rect 4176 4164 4189 4178
rect 4204 4164 4220 4180
rect 4266 4175 4277 4188
rect 4059 4130 4060 4146
rect 4075 4130 4088 4152
rect 4103 4130 4133 4152
rect 4176 4148 4238 4164
rect 4266 4157 4277 4173
rect 4282 4168 4292 4188
rect 4302 4168 4316 4188
rect 4319 4175 4328 4188
rect 4344 4175 4353 4188
rect 4282 4157 4316 4168
rect 4319 4157 4328 4173
rect 4344 4157 4353 4173
rect 4360 4168 4370 4188
rect 4380 4168 4394 4188
rect 4395 4175 4406 4188
rect 4360 4157 4394 4168
rect 4395 4157 4406 4173
rect 4452 4164 4468 4180
rect 4475 4178 4505 4230
rect 4539 4226 4540 4233
rect 4524 4218 4540 4226
rect 4511 4186 4524 4205
rect 4539 4186 4569 4202
rect 4511 4170 4585 4186
rect 4511 4168 4524 4170
rect 4539 4168 4573 4170
rect 4176 4146 4189 4148
rect 4204 4146 4238 4148
rect 4176 4130 4238 4146
rect 4282 4141 4298 4144
rect 4360 4141 4390 4152
rect 4438 4148 4484 4164
rect 4511 4152 4585 4168
rect 4438 4146 4472 4148
rect 4437 4130 4484 4146
rect 4511 4130 4524 4152
rect 4539 4130 4569 4152
rect 4596 4130 4597 4146
rect 4612 4130 4625 4290
rect -7 4122 34 4130
rect -7 4096 8 4122
rect 15 4096 34 4122
rect 98 4118 160 4130
rect 172 4118 247 4130
rect 305 4118 380 4130
rect 392 4118 423 4130
rect 429 4118 464 4130
rect 98 4116 260 4118
rect -7 4088 34 4096
rect 116 4092 129 4116
rect 144 4114 159 4116
rect -1 4078 0 4088
rect 15 4078 28 4088
rect 43 4078 73 4092
rect 116 4078 159 4092
rect 183 4089 190 4096
rect 193 4092 260 4116
rect 292 4116 464 4118
rect 262 4094 290 4098
rect 292 4094 372 4116
rect 393 4114 408 4116
rect 262 4092 372 4094
rect 193 4088 372 4092
rect 166 4078 196 4088
rect 198 4078 351 4088
rect 359 4078 389 4088
rect 393 4078 423 4092
rect 451 4078 464 4116
rect 536 4122 571 4130
rect 536 4096 537 4122
rect 544 4096 571 4122
rect 479 4078 509 4092
rect 536 4088 571 4096
rect 573 4122 614 4130
rect 573 4096 588 4122
rect 595 4096 614 4122
rect 678 4118 740 4130
rect 752 4118 827 4130
rect 885 4118 960 4130
rect 972 4118 1003 4130
rect 1009 4118 1044 4130
rect 678 4116 840 4118
rect 573 4088 614 4096
rect 696 4092 709 4116
rect 724 4114 739 4116
rect 536 4078 537 4088
rect 552 4078 565 4088
rect 579 4078 580 4088
rect 595 4078 608 4088
rect 623 4078 653 4092
rect 696 4078 739 4092
rect 763 4089 770 4096
rect 773 4092 840 4116
rect 872 4116 1044 4118
rect 842 4094 870 4098
rect 872 4094 952 4116
rect 973 4114 988 4116
rect 842 4092 952 4094
rect 773 4088 952 4092
rect 746 4078 776 4088
rect 778 4078 931 4088
rect 939 4078 969 4088
rect 973 4078 1003 4092
rect 1031 4078 1044 4116
rect 1116 4122 1151 4130
rect 1116 4096 1117 4122
rect 1124 4096 1151 4122
rect 1059 4078 1089 4092
rect 1116 4088 1151 4096
rect 1153 4122 1194 4130
rect 1153 4096 1168 4122
rect 1175 4096 1194 4122
rect 1258 4118 1320 4130
rect 1332 4118 1407 4130
rect 1465 4118 1540 4130
rect 1552 4118 1583 4130
rect 1589 4118 1624 4130
rect 1258 4116 1420 4118
rect 1153 4088 1194 4096
rect 1276 4092 1289 4116
rect 1304 4114 1319 4116
rect 1116 4078 1117 4088
rect 1132 4078 1145 4088
rect 1159 4078 1160 4088
rect 1175 4078 1188 4088
rect 1203 4078 1233 4092
rect 1276 4078 1319 4092
rect 1343 4089 1350 4096
rect 1353 4092 1420 4116
rect 1452 4116 1624 4118
rect 1422 4094 1450 4098
rect 1452 4094 1532 4116
rect 1553 4114 1568 4116
rect 1422 4092 1532 4094
rect 1353 4088 1532 4092
rect 1326 4078 1356 4088
rect 1358 4078 1511 4088
rect 1519 4078 1549 4088
rect 1553 4078 1583 4092
rect 1611 4078 1624 4116
rect 1696 4122 1731 4130
rect 1696 4096 1697 4122
rect 1704 4096 1731 4122
rect 1639 4078 1669 4092
rect 1696 4088 1731 4096
rect 1733 4122 1774 4130
rect 1733 4096 1748 4122
rect 1755 4096 1774 4122
rect 1838 4118 1900 4130
rect 1912 4118 1987 4130
rect 2045 4118 2120 4130
rect 2132 4118 2163 4130
rect 2169 4118 2204 4130
rect 1838 4116 2000 4118
rect 1733 4088 1774 4096
rect 1856 4092 1869 4116
rect 1884 4114 1899 4116
rect 1696 4078 1697 4088
rect 1712 4078 1725 4088
rect 1739 4078 1740 4088
rect 1755 4078 1768 4088
rect 1783 4078 1813 4092
rect 1856 4078 1899 4092
rect 1923 4089 1930 4096
rect 1933 4092 2000 4116
rect 2032 4116 2204 4118
rect 2002 4094 2030 4098
rect 2032 4094 2112 4116
rect 2133 4114 2148 4116
rect 2002 4092 2112 4094
rect 1933 4088 2112 4092
rect 1906 4078 1936 4088
rect 1938 4078 2091 4088
rect 2099 4078 2129 4088
rect 2133 4078 2163 4092
rect 2191 4078 2204 4116
rect 2276 4122 2311 4130
rect 2276 4096 2277 4122
rect 2284 4096 2311 4122
rect 2219 4078 2249 4092
rect 2276 4088 2311 4096
rect 2313 4122 2354 4130
rect 2313 4096 2328 4122
rect 2335 4096 2354 4122
rect 2418 4118 2480 4130
rect 2492 4118 2567 4130
rect 2625 4118 2700 4130
rect 2712 4118 2743 4130
rect 2749 4118 2784 4130
rect 2418 4116 2580 4118
rect 2313 4088 2354 4096
rect 2436 4092 2449 4116
rect 2464 4114 2479 4116
rect 2276 4078 2277 4088
rect 2292 4078 2305 4088
rect 2319 4078 2320 4088
rect 2335 4078 2348 4088
rect 2363 4078 2393 4092
rect 2436 4078 2479 4092
rect 2503 4089 2510 4096
rect 2513 4092 2580 4116
rect 2612 4116 2784 4118
rect 2582 4094 2610 4098
rect 2612 4094 2692 4116
rect 2713 4114 2728 4116
rect 2582 4092 2692 4094
rect 2513 4088 2692 4092
rect 2486 4078 2516 4088
rect 2518 4078 2671 4088
rect 2679 4078 2709 4088
rect 2713 4078 2743 4092
rect 2771 4078 2784 4116
rect 2856 4122 2891 4130
rect 2856 4096 2857 4122
rect 2864 4096 2891 4122
rect 2799 4078 2829 4092
rect 2856 4088 2891 4096
rect 2893 4122 2934 4130
rect 2893 4096 2908 4122
rect 2915 4096 2934 4122
rect 2998 4118 3060 4130
rect 3072 4118 3147 4130
rect 3205 4118 3280 4130
rect 3292 4118 3323 4130
rect 3329 4118 3364 4130
rect 2998 4116 3160 4118
rect 2893 4088 2934 4096
rect 3016 4092 3029 4116
rect 3044 4114 3059 4116
rect 2856 4078 2857 4088
rect 2872 4078 2885 4088
rect 2899 4078 2900 4088
rect 2915 4078 2928 4088
rect 2943 4078 2973 4092
rect 3016 4078 3059 4092
rect 3083 4089 3090 4096
rect 3093 4092 3160 4116
rect 3192 4116 3364 4118
rect 3162 4094 3190 4098
rect 3192 4094 3272 4116
rect 3293 4114 3308 4116
rect 3162 4092 3272 4094
rect 3093 4088 3272 4092
rect 3066 4078 3096 4088
rect 3098 4078 3251 4088
rect 3259 4078 3289 4088
rect 3293 4078 3323 4092
rect 3351 4078 3364 4116
rect 3436 4122 3471 4130
rect 3436 4096 3437 4122
rect 3444 4096 3471 4122
rect 3379 4078 3409 4092
rect 3436 4088 3471 4096
rect 3473 4122 3514 4130
rect 3473 4096 3488 4122
rect 3495 4096 3514 4122
rect 3578 4118 3640 4130
rect 3652 4118 3727 4130
rect 3785 4118 3860 4130
rect 3872 4118 3903 4130
rect 3909 4118 3944 4130
rect 3578 4116 3740 4118
rect 3473 4088 3514 4096
rect 3596 4092 3609 4116
rect 3624 4114 3639 4116
rect 3436 4078 3437 4088
rect 3452 4078 3465 4088
rect 3479 4078 3480 4088
rect 3495 4078 3508 4088
rect 3523 4078 3553 4092
rect 3596 4078 3639 4092
rect 3663 4089 3670 4096
rect 3673 4092 3740 4116
rect 3772 4116 3944 4118
rect 3742 4094 3770 4098
rect 3772 4094 3852 4116
rect 3873 4114 3888 4116
rect 3742 4092 3852 4094
rect 3673 4088 3852 4092
rect 3646 4078 3676 4088
rect 3678 4078 3831 4088
rect 3839 4078 3869 4088
rect 3873 4078 3903 4092
rect 3931 4078 3944 4116
rect 4016 4122 4051 4130
rect 4016 4096 4017 4122
rect 4024 4096 4051 4122
rect 3959 4078 3989 4092
rect 4016 4088 4051 4096
rect 4053 4122 4094 4130
rect 4053 4096 4068 4122
rect 4075 4096 4094 4122
rect 4158 4118 4220 4130
rect 4232 4118 4307 4130
rect 4365 4118 4440 4130
rect 4452 4118 4483 4130
rect 4489 4118 4524 4130
rect 4158 4116 4320 4118
rect 4053 4088 4094 4096
rect 4176 4092 4189 4116
rect 4204 4114 4219 4116
rect 4016 4078 4017 4088
rect 4032 4078 4045 4088
rect 4059 4078 4060 4088
rect 4075 4078 4088 4088
rect 4103 4078 4133 4092
rect 4176 4078 4219 4092
rect 4243 4089 4250 4096
rect 4253 4092 4320 4116
rect 4352 4116 4524 4118
rect 4322 4094 4350 4098
rect 4352 4094 4432 4116
rect 4453 4114 4468 4116
rect 4322 4092 4432 4094
rect 4253 4088 4432 4092
rect 4226 4078 4256 4088
rect 4258 4078 4411 4088
rect 4419 4078 4449 4088
rect 4453 4078 4483 4092
rect 4511 4078 4524 4116
rect 4596 4122 4631 4130
rect 4596 4096 4597 4122
rect 4604 4096 4631 4122
rect 4539 4078 4569 4092
rect 4596 4088 4631 4096
rect 4596 4078 4597 4088
rect 4612 4078 4625 4088
rect -1 4072 4625 4078
rect 0 4064 4625 4072
rect 15 4034 28 4064
rect 43 4046 73 4064
rect 116 4050 130 4064
rect 166 4050 386 4064
rect 117 4048 130 4050
rect 83 4036 98 4048
rect 80 4034 102 4036
rect 107 4034 137 4048
rect 198 4046 351 4050
rect 180 4034 372 4046
rect 415 4034 445 4048
rect 451 4034 464 4064
rect 479 4046 509 4064
rect 552 4034 565 4064
rect 595 4034 608 4064
rect 623 4046 653 4064
rect 696 4050 710 4064
rect 746 4050 966 4064
rect 697 4048 710 4050
rect 663 4036 678 4048
rect 660 4034 682 4036
rect 687 4034 717 4048
rect 778 4046 931 4050
rect 760 4034 952 4046
rect 995 4034 1025 4048
rect 1031 4034 1044 4064
rect 1059 4046 1089 4064
rect 1132 4034 1145 4064
rect 1175 4034 1188 4064
rect 1203 4046 1233 4064
rect 1276 4050 1290 4064
rect 1326 4050 1546 4064
rect 1277 4048 1290 4050
rect 1243 4036 1258 4048
rect 1240 4034 1262 4036
rect 1267 4034 1297 4048
rect 1358 4046 1511 4050
rect 1340 4034 1532 4046
rect 1575 4034 1605 4048
rect 1611 4034 1624 4064
rect 1639 4046 1669 4064
rect 1712 4034 1725 4064
rect 1755 4034 1768 4064
rect 1783 4046 1813 4064
rect 1856 4050 1870 4064
rect 1906 4050 2126 4064
rect 1857 4048 1870 4050
rect 1823 4036 1838 4048
rect 1820 4034 1842 4036
rect 1847 4034 1877 4048
rect 1938 4046 2091 4050
rect 1920 4034 2112 4046
rect 2155 4034 2185 4048
rect 2191 4034 2204 4064
rect 2219 4046 2249 4064
rect 2292 4034 2305 4064
rect 2335 4034 2348 4064
rect 2363 4046 2393 4064
rect 2436 4050 2450 4064
rect 2486 4050 2706 4064
rect 2437 4048 2450 4050
rect 2403 4036 2418 4048
rect 2400 4034 2422 4036
rect 2427 4034 2457 4048
rect 2518 4046 2671 4050
rect 2500 4034 2692 4046
rect 2735 4034 2765 4048
rect 2771 4034 2784 4064
rect 2799 4046 2829 4064
rect 2872 4034 2885 4064
rect 2915 4034 2928 4064
rect 2943 4046 2973 4064
rect 3016 4050 3030 4064
rect 3066 4050 3286 4064
rect 3017 4048 3030 4050
rect 2983 4036 2998 4048
rect 2980 4034 3002 4036
rect 3007 4034 3037 4048
rect 3098 4046 3251 4050
rect 3080 4034 3272 4046
rect 3315 4034 3345 4048
rect 3351 4034 3364 4064
rect 3379 4046 3409 4064
rect 3452 4034 3465 4064
rect 3495 4034 3508 4064
rect 3523 4046 3553 4064
rect 3596 4050 3610 4064
rect 3646 4050 3866 4064
rect 3597 4048 3610 4050
rect 3563 4036 3578 4048
rect 3560 4034 3582 4036
rect 3587 4034 3617 4048
rect 3678 4046 3831 4050
rect 3660 4034 3852 4046
rect 3895 4034 3925 4048
rect 3931 4034 3944 4064
rect 3959 4046 3989 4064
rect 4032 4034 4045 4064
rect 4075 4034 4088 4064
rect 4103 4046 4133 4064
rect 4176 4050 4190 4064
rect 4226 4050 4446 4064
rect 4177 4048 4190 4050
rect 4143 4036 4158 4048
rect 4140 4034 4162 4036
rect 4167 4034 4197 4048
rect 4258 4046 4411 4050
rect 4240 4034 4432 4046
rect 4475 4034 4505 4048
rect 4511 4034 4524 4064
rect 4539 4046 4569 4064
rect 4612 4034 4625 4064
rect 0 4020 4625 4034
rect 15 3916 28 4020
rect 73 3998 74 4008
rect 89 3998 102 4008
rect 73 3994 102 3998
rect 107 3994 137 4020
rect 155 4006 171 4008
rect 243 4006 296 4020
rect 244 4004 308 4006
rect 351 4004 366 4020
rect 415 4017 445 4020
rect 415 4014 451 4017
rect 381 4006 397 4008
rect 155 3994 170 3998
rect 73 3992 170 3994
rect 198 3992 366 4004
rect 382 3994 397 3998
rect 415 3995 454 4014
rect 473 4008 480 4009
rect 479 4001 480 4008
rect 463 3998 464 4001
rect 479 3998 492 4001
rect 415 3994 445 3995
rect 454 3994 460 3995
rect 463 3994 492 3998
rect 382 3993 492 3994
rect 382 3992 498 3993
rect 57 3984 108 3992
rect 57 3972 82 3984
rect 89 3972 108 3984
rect 139 3984 189 3992
rect 139 3976 155 3984
rect 162 3982 189 3984
rect 198 3982 419 3992
rect 162 3972 419 3982
rect 448 3984 498 3992
rect 448 3975 464 3984
rect 57 3964 108 3972
rect 155 3964 419 3972
rect 445 3972 464 3975
rect 471 3972 498 3984
rect 445 3964 498 3972
rect 73 3956 74 3964
rect 89 3956 102 3964
rect 73 3948 89 3956
rect 70 3941 89 3944
rect 70 3932 92 3941
rect 43 3922 92 3932
rect 43 3916 73 3922
rect 92 3917 97 3922
rect 15 3900 89 3916
rect 107 3908 137 3964
rect 172 3954 380 3964
rect 415 3960 460 3964
rect 463 3963 464 3964
rect 479 3963 492 3964
rect 198 3924 387 3954
rect 213 3921 387 3924
rect 206 3918 387 3921
rect 15 3898 28 3900
rect 43 3898 77 3900
rect 15 3882 89 3898
rect 116 3894 129 3908
rect 144 3894 160 3910
rect 206 3905 217 3918
rect -1 3860 0 3876
rect 15 3860 28 3882
rect 43 3860 73 3882
rect 116 3878 178 3894
rect 206 3887 217 3903
rect 222 3898 232 3918
rect 242 3898 256 3918
rect 259 3905 268 3918
rect 284 3905 293 3918
rect 222 3887 256 3898
rect 259 3887 268 3903
rect 284 3887 293 3903
rect 300 3898 310 3918
rect 320 3898 334 3918
rect 335 3905 346 3918
rect 300 3887 334 3898
rect 335 3887 346 3903
rect 392 3894 408 3910
rect 415 3908 445 3960
rect 479 3956 480 3963
rect 464 3948 480 3956
rect 451 3916 464 3935
rect 479 3916 509 3932
rect 451 3900 525 3916
rect 451 3898 464 3900
rect 479 3898 513 3900
rect 116 3876 129 3878
rect 144 3876 178 3878
rect 116 3860 178 3876
rect 222 3871 238 3874
rect 300 3871 330 3882
rect 378 3878 424 3894
rect 451 3882 525 3898
rect 378 3876 412 3878
rect 377 3860 424 3876
rect 451 3860 464 3882
rect 479 3860 509 3882
rect 536 3860 537 3876
rect 552 3860 565 4020
rect 595 3916 608 4020
rect 653 3998 654 4008
rect 669 3998 682 4008
rect 653 3994 682 3998
rect 687 3994 717 4020
rect 735 4006 751 4008
rect 823 4006 876 4020
rect 824 4004 888 4006
rect 931 4004 946 4020
rect 995 4017 1025 4020
rect 995 4014 1031 4017
rect 961 4006 977 4008
rect 735 3994 750 3998
rect 653 3992 750 3994
rect 778 3992 946 4004
rect 962 3994 977 3998
rect 995 3995 1034 4014
rect 1053 4008 1060 4009
rect 1059 4001 1060 4008
rect 1043 3998 1044 4001
rect 1059 3998 1072 4001
rect 995 3994 1025 3995
rect 1034 3994 1040 3995
rect 1043 3994 1072 3998
rect 962 3993 1072 3994
rect 962 3992 1078 3993
rect 637 3984 688 3992
rect 637 3972 662 3984
rect 669 3972 688 3984
rect 719 3984 769 3992
rect 719 3976 735 3984
rect 742 3982 769 3984
rect 778 3982 999 3992
rect 742 3972 999 3982
rect 1028 3984 1078 3992
rect 1028 3975 1044 3984
rect 637 3964 688 3972
rect 735 3964 999 3972
rect 1025 3972 1044 3975
rect 1051 3972 1078 3984
rect 1025 3964 1078 3972
rect 653 3956 654 3964
rect 669 3956 682 3964
rect 653 3948 669 3956
rect 650 3941 669 3944
rect 650 3932 672 3941
rect 623 3922 672 3932
rect 623 3916 653 3922
rect 672 3917 677 3922
rect 595 3900 669 3916
rect 687 3908 717 3964
rect 752 3954 960 3964
rect 995 3960 1040 3964
rect 1043 3963 1044 3964
rect 1059 3963 1072 3964
rect 778 3924 967 3954
rect 793 3921 967 3924
rect 786 3918 967 3921
rect 595 3898 608 3900
rect 623 3898 657 3900
rect 595 3882 669 3898
rect 696 3894 709 3908
rect 724 3894 740 3910
rect 786 3905 797 3918
rect 579 3860 580 3876
rect 595 3860 608 3882
rect 623 3860 653 3882
rect 696 3878 758 3894
rect 786 3887 797 3903
rect 802 3898 812 3918
rect 822 3898 836 3918
rect 839 3905 848 3918
rect 864 3905 873 3918
rect 802 3887 836 3898
rect 839 3887 848 3903
rect 864 3887 873 3903
rect 880 3898 890 3918
rect 900 3898 914 3918
rect 915 3905 926 3918
rect 880 3887 914 3898
rect 915 3887 926 3903
rect 972 3894 988 3910
rect 995 3908 1025 3960
rect 1059 3956 1060 3963
rect 1044 3948 1060 3956
rect 1031 3916 1044 3935
rect 1059 3916 1089 3932
rect 1031 3900 1105 3916
rect 1031 3898 1044 3900
rect 1059 3898 1093 3900
rect 696 3876 709 3878
rect 724 3876 758 3878
rect 696 3860 758 3876
rect 802 3871 818 3874
rect 880 3871 910 3882
rect 958 3878 1004 3894
rect 1031 3882 1105 3898
rect 958 3876 992 3878
rect 957 3860 1004 3876
rect 1031 3860 1044 3882
rect 1059 3860 1089 3882
rect 1116 3860 1117 3876
rect 1132 3860 1145 4020
rect 1175 3916 1188 4020
rect 1233 3998 1234 4008
rect 1249 3998 1262 4008
rect 1233 3994 1262 3998
rect 1267 3994 1297 4020
rect 1315 4006 1331 4008
rect 1403 4006 1456 4020
rect 1404 4004 1468 4006
rect 1511 4004 1526 4020
rect 1575 4017 1605 4020
rect 1575 4014 1611 4017
rect 1541 4006 1557 4008
rect 1315 3994 1330 3998
rect 1233 3992 1330 3994
rect 1358 3992 1526 4004
rect 1542 3994 1557 3998
rect 1575 3995 1614 4014
rect 1633 4008 1640 4009
rect 1639 4001 1640 4008
rect 1623 3998 1624 4001
rect 1639 3998 1652 4001
rect 1575 3994 1605 3995
rect 1614 3994 1620 3995
rect 1623 3994 1652 3998
rect 1542 3993 1652 3994
rect 1542 3992 1658 3993
rect 1217 3984 1268 3992
rect 1217 3972 1242 3984
rect 1249 3972 1268 3984
rect 1299 3984 1349 3992
rect 1299 3976 1315 3984
rect 1322 3982 1349 3984
rect 1358 3982 1579 3992
rect 1322 3972 1579 3982
rect 1608 3984 1658 3992
rect 1608 3975 1624 3984
rect 1217 3964 1268 3972
rect 1315 3964 1579 3972
rect 1605 3972 1624 3975
rect 1631 3972 1658 3984
rect 1605 3964 1658 3972
rect 1233 3956 1234 3964
rect 1249 3956 1262 3964
rect 1233 3948 1249 3956
rect 1230 3941 1249 3944
rect 1230 3932 1252 3941
rect 1203 3922 1252 3932
rect 1203 3916 1233 3922
rect 1252 3917 1257 3922
rect 1175 3900 1249 3916
rect 1267 3908 1297 3964
rect 1332 3954 1540 3964
rect 1575 3960 1620 3964
rect 1623 3963 1624 3964
rect 1639 3963 1652 3964
rect 1358 3924 1547 3954
rect 1373 3921 1547 3924
rect 1366 3918 1547 3921
rect 1175 3898 1188 3900
rect 1203 3898 1237 3900
rect 1175 3882 1249 3898
rect 1276 3894 1289 3908
rect 1304 3894 1320 3910
rect 1366 3905 1377 3918
rect 1159 3860 1160 3876
rect 1175 3860 1188 3882
rect 1203 3860 1233 3882
rect 1276 3878 1338 3894
rect 1366 3887 1377 3903
rect 1382 3898 1392 3918
rect 1402 3898 1416 3918
rect 1419 3905 1428 3918
rect 1444 3905 1453 3918
rect 1382 3887 1416 3898
rect 1419 3887 1428 3903
rect 1444 3887 1453 3903
rect 1460 3898 1470 3918
rect 1480 3898 1494 3918
rect 1495 3905 1506 3918
rect 1460 3887 1494 3898
rect 1495 3887 1506 3903
rect 1552 3894 1568 3910
rect 1575 3908 1605 3960
rect 1639 3956 1640 3963
rect 1624 3948 1640 3956
rect 1611 3916 1624 3935
rect 1639 3916 1669 3932
rect 1611 3900 1685 3916
rect 1611 3898 1624 3900
rect 1639 3898 1673 3900
rect 1276 3876 1289 3878
rect 1304 3876 1338 3878
rect 1276 3860 1338 3876
rect 1382 3871 1398 3874
rect 1460 3871 1490 3882
rect 1538 3878 1584 3894
rect 1611 3882 1685 3898
rect 1538 3876 1572 3878
rect 1537 3860 1584 3876
rect 1611 3860 1624 3882
rect 1639 3860 1669 3882
rect 1696 3860 1697 3876
rect 1712 3860 1725 4020
rect 1755 3916 1768 4020
rect 1813 3998 1814 4008
rect 1829 3998 1842 4008
rect 1813 3994 1842 3998
rect 1847 3994 1877 4020
rect 1895 4006 1911 4008
rect 1983 4006 2036 4020
rect 1984 4004 2048 4006
rect 2091 4004 2106 4020
rect 2155 4017 2185 4020
rect 2155 4014 2191 4017
rect 2121 4006 2137 4008
rect 1895 3994 1910 3998
rect 1813 3992 1910 3994
rect 1938 3992 2106 4004
rect 2122 3994 2137 3998
rect 2155 3995 2194 4014
rect 2213 4008 2220 4009
rect 2219 4001 2220 4008
rect 2203 3998 2204 4001
rect 2219 3998 2232 4001
rect 2155 3994 2185 3995
rect 2194 3994 2200 3995
rect 2203 3994 2232 3998
rect 2122 3993 2232 3994
rect 2122 3992 2238 3993
rect 1797 3984 1848 3992
rect 1797 3972 1822 3984
rect 1829 3972 1848 3984
rect 1879 3984 1929 3992
rect 1879 3976 1895 3984
rect 1902 3982 1929 3984
rect 1938 3982 2159 3992
rect 1902 3972 2159 3982
rect 2188 3984 2238 3992
rect 2188 3975 2204 3984
rect 1797 3964 1848 3972
rect 1895 3964 2159 3972
rect 2185 3972 2204 3975
rect 2211 3972 2238 3984
rect 2185 3964 2238 3972
rect 1813 3956 1814 3964
rect 1829 3956 1842 3964
rect 1813 3948 1829 3956
rect 1810 3941 1829 3944
rect 1810 3932 1832 3941
rect 1783 3922 1832 3932
rect 1783 3916 1813 3922
rect 1832 3917 1837 3922
rect 1755 3900 1829 3916
rect 1847 3908 1877 3964
rect 1912 3954 2120 3964
rect 2155 3960 2200 3964
rect 2203 3963 2204 3964
rect 2219 3963 2232 3964
rect 1938 3924 2127 3954
rect 1953 3921 2127 3924
rect 1946 3918 2127 3921
rect 1755 3898 1768 3900
rect 1783 3898 1817 3900
rect 1755 3882 1829 3898
rect 1856 3894 1869 3908
rect 1884 3894 1900 3910
rect 1946 3905 1957 3918
rect 1739 3860 1740 3876
rect 1755 3860 1768 3882
rect 1783 3860 1813 3882
rect 1856 3878 1918 3894
rect 1946 3887 1957 3903
rect 1962 3898 1972 3918
rect 1982 3898 1996 3918
rect 1999 3905 2008 3918
rect 2024 3905 2033 3918
rect 1962 3887 1996 3898
rect 1999 3887 2008 3903
rect 2024 3887 2033 3903
rect 2040 3898 2050 3918
rect 2060 3898 2074 3918
rect 2075 3905 2086 3918
rect 2040 3887 2074 3898
rect 2075 3887 2086 3903
rect 2132 3894 2148 3910
rect 2155 3908 2185 3960
rect 2219 3956 2220 3963
rect 2204 3948 2220 3956
rect 2191 3916 2204 3935
rect 2219 3916 2249 3932
rect 2191 3900 2265 3916
rect 2191 3898 2204 3900
rect 2219 3898 2253 3900
rect 1856 3876 1869 3878
rect 1884 3876 1918 3878
rect 1856 3860 1918 3876
rect 1962 3871 1978 3874
rect 2040 3871 2070 3882
rect 2118 3878 2164 3894
rect 2191 3882 2265 3898
rect 2118 3876 2152 3878
rect 2117 3860 2164 3876
rect 2191 3860 2204 3882
rect 2219 3860 2249 3882
rect 2276 3860 2277 3876
rect 2292 3860 2305 4020
rect 2335 3916 2348 4020
rect 2393 3998 2394 4008
rect 2409 3998 2422 4008
rect 2393 3994 2422 3998
rect 2427 3994 2457 4020
rect 2475 4006 2491 4008
rect 2563 4006 2616 4020
rect 2564 4004 2628 4006
rect 2671 4004 2686 4020
rect 2735 4017 2765 4020
rect 2735 4014 2771 4017
rect 2701 4006 2717 4008
rect 2475 3994 2490 3998
rect 2393 3992 2490 3994
rect 2518 3992 2686 4004
rect 2702 3994 2717 3998
rect 2735 3995 2774 4014
rect 2793 4008 2800 4009
rect 2799 4001 2800 4008
rect 2783 3998 2784 4001
rect 2799 3998 2812 4001
rect 2735 3994 2765 3995
rect 2774 3994 2780 3995
rect 2783 3994 2812 3998
rect 2702 3993 2812 3994
rect 2702 3992 2818 3993
rect 2377 3984 2428 3992
rect 2377 3972 2402 3984
rect 2409 3972 2428 3984
rect 2459 3984 2509 3992
rect 2459 3976 2475 3984
rect 2482 3982 2509 3984
rect 2518 3982 2739 3992
rect 2482 3972 2739 3982
rect 2768 3984 2818 3992
rect 2768 3975 2784 3984
rect 2377 3964 2428 3972
rect 2475 3964 2739 3972
rect 2765 3972 2784 3975
rect 2791 3972 2818 3984
rect 2765 3964 2818 3972
rect 2393 3956 2394 3964
rect 2409 3956 2422 3964
rect 2393 3948 2409 3956
rect 2390 3941 2409 3944
rect 2390 3932 2412 3941
rect 2363 3922 2412 3932
rect 2363 3916 2393 3922
rect 2412 3917 2417 3922
rect 2335 3900 2409 3916
rect 2427 3908 2457 3964
rect 2492 3954 2700 3964
rect 2735 3960 2780 3964
rect 2783 3963 2784 3964
rect 2799 3963 2812 3964
rect 2518 3924 2707 3954
rect 2533 3921 2707 3924
rect 2526 3918 2707 3921
rect 2335 3898 2348 3900
rect 2363 3898 2397 3900
rect 2335 3882 2409 3898
rect 2436 3894 2449 3908
rect 2464 3894 2480 3910
rect 2526 3905 2537 3918
rect 2319 3860 2320 3876
rect 2335 3860 2348 3882
rect 2363 3860 2393 3882
rect 2436 3878 2498 3894
rect 2526 3887 2537 3903
rect 2542 3898 2552 3918
rect 2562 3898 2576 3918
rect 2579 3905 2588 3918
rect 2604 3905 2613 3918
rect 2542 3887 2576 3898
rect 2579 3887 2588 3903
rect 2604 3887 2613 3903
rect 2620 3898 2630 3918
rect 2640 3898 2654 3918
rect 2655 3905 2666 3918
rect 2620 3887 2654 3898
rect 2655 3887 2666 3903
rect 2712 3894 2728 3910
rect 2735 3908 2765 3960
rect 2799 3956 2800 3963
rect 2784 3948 2800 3956
rect 2771 3916 2784 3935
rect 2799 3916 2829 3932
rect 2771 3900 2845 3916
rect 2771 3898 2784 3900
rect 2799 3898 2833 3900
rect 2436 3876 2449 3878
rect 2464 3876 2498 3878
rect 2436 3860 2498 3876
rect 2542 3871 2558 3874
rect 2620 3871 2650 3882
rect 2698 3878 2744 3894
rect 2771 3882 2845 3898
rect 2698 3876 2732 3878
rect 2697 3860 2744 3876
rect 2771 3860 2784 3882
rect 2799 3860 2829 3882
rect 2856 3860 2857 3876
rect 2872 3860 2885 4020
rect 2915 3916 2928 4020
rect 2973 3998 2974 4008
rect 2989 3998 3002 4008
rect 2973 3994 3002 3998
rect 3007 3994 3037 4020
rect 3055 4006 3071 4008
rect 3143 4006 3196 4020
rect 3144 4004 3208 4006
rect 3251 4004 3266 4020
rect 3315 4017 3345 4020
rect 3315 4014 3351 4017
rect 3281 4006 3297 4008
rect 3055 3994 3070 3998
rect 2973 3992 3070 3994
rect 3098 3992 3266 4004
rect 3282 3994 3297 3998
rect 3315 3995 3354 4014
rect 3373 4008 3380 4009
rect 3379 4001 3380 4008
rect 3363 3998 3364 4001
rect 3379 3998 3392 4001
rect 3315 3994 3345 3995
rect 3354 3994 3360 3995
rect 3363 3994 3392 3998
rect 3282 3993 3392 3994
rect 3282 3992 3398 3993
rect 2957 3984 3008 3992
rect 2957 3972 2982 3984
rect 2989 3972 3008 3984
rect 3039 3984 3089 3992
rect 3039 3976 3055 3984
rect 3062 3982 3089 3984
rect 3098 3982 3319 3992
rect 3062 3972 3319 3982
rect 3348 3984 3398 3992
rect 3348 3975 3364 3984
rect 2957 3964 3008 3972
rect 3055 3964 3319 3972
rect 3345 3972 3364 3975
rect 3371 3972 3398 3984
rect 3345 3964 3398 3972
rect 2973 3956 2974 3964
rect 2989 3956 3002 3964
rect 2973 3948 2989 3956
rect 2970 3941 2989 3944
rect 2970 3932 2992 3941
rect 2943 3922 2992 3932
rect 2943 3916 2973 3922
rect 2992 3917 2997 3922
rect 2915 3900 2989 3916
rect 3007 3908 3037 3964
rect 3072 3954 3280 3964
rect 3315 3960 3360 3964
rect 3363 3963 3364 3964
rect 3379 3963 3392 3964
rect 3098 3924 3287 3954
rect 3113 3921 3287 3924
rect 3106 3918 3287 3921
rect 2915 3898 2928 3900
rect 2943 3898 2977 3900
rect 2915 3882 2989 3898
rect 3016 3894 3029 3908
rect 3044 3894 3060 3910
rect 3106 3905 3117 3918
rect 2899 3860 2900 3876
rect 2915 3860 2928 3882
rect 2943 3860 2973 3882
rect 3016 3878 3078 3894
rect 3106 3887 3117 3903
rect 3122 3898 3132 3918
rect 3142 3898 3156 3918
rect 3159 3905 3168 3918
rect 3184 3905 3193 3918
rect 3122 3887 3156 3898
rect 3159 3887 3168 3903
rect 3184 3887 3193 3903
rect 3200 3898 3210 3918
rect 3220 3898 3234 3918
rect 3235 3905 3246 3918
rect 3200 3887 3234 3898
rect 3235 3887 3246 3903
rect 3292 3894 3308 3910
rect 3315 3908 3345 3960
rect 3379 3956 3380 3963
rect 3364 3948 3380 3956
rect 3351 3916 3364 3935
rect 3379 3916 3409 3932
rect 3351 3900 3425 3916
rect 3351 3898 3364 3900
rect 3379 3898 3413 3900
rect 3016 3876 3029 3878
rect 3044 3876 3078 3878
rect 3016 3860 3078 3876
rect 3122 3871 3138 3874
rect 3200 3871 3230 3882
rect 3278 3878 3324 3894
rect 3351 3882 3425 3898
rect 3278 3876 3312 3878
rect 3277 3860 3324 3876
rect 3351 3860 3364 3882
rect 3379 3860 3409 3882
rect 3436 3860 3437 3876
rect 3452 3860 3465 4020
rect 3495 3916 3508 4020
rect 3553 3998 3554 4008
rect 3569 3998 3582 4008
rect 3553 3994 3582 3998
rect 3587 3994 3617 4020
rect 3635 4006 3651 4008
rect 3723 4006 3776 4020
rect 3724 4004 3788 4006
rect 3831 4004 3846 4020
rect 3895 4017 3925 4020
rect 3895 4014 3931 4017
rect 3861 4006 3877 4008
rect 3635 3994 3650 3998
rect 3553 3992 3650 3994
rect 3678 3992 3846 4004
rect 3862 3994 3877 3998
rect 3895 3995 3934 4014
rect 3953 4008 3960 4009
rect 3959 4001 3960 4008
rect 3943 3998 3944 4001
rect 3959 3998 3972 4001
rect 3895 3994 3925 3995
rect 3934 3994 3940 3995
rect 3943 3994 3972 3998
rect 3862 3993 3972 3994
rect 3862 3992 3978 3993
rect 3537 3984 3588 3992
rect 3537 3972 3562 3984
rect 3569 3972 3588 3984
rect 3619 3984 3669 3992
rect 3619 3976 3635 3984
rect 3642 3982 3669 3984
rect 3678 3982 3899 3992
rect 3642 3972 3899 3982
rect 3928 3984 3978 3992
rect 3928 3975 3944 3984
rect 3537 3964 3588 3972
rect 3635 3964 3899 3972
rect 3925 3972 3944 3975
rect 3951 3972 3978 3984
rect 3925 3964 3978 3972
rect 3553 3956 3554 3964
rect 3569 3956 3582 3964
rect 3553 3948 3569 3956
rect 3550 3941 3569 3944
rect 3550 3932 3572 3941
rect 3523 3922 3572 3932
rect 3523 3916 3553 3922
rect 3572 3917 3577 3922
rect 3495 3900 3569 3916
rect 3587 3908 3617 3964
rect 3652 3954 3860 3964
rect 3895 3960 3940 3964
rect 3943 3963 3944 3964
rect 3959 3963 3972 3964
rect 3678 3924 3867 3954
rect 3693 3921 3867 3924
rect 3686 3918 3867 3921
rect 3495 3898 3508 3900
rect 3523 3898 3557 3900
rect 3495 3882 3569 3898
rect 3596 3894 3609 3908
rect 3624 3894 3640 3910
rect 3686 3905 3697 3918
rect 3479 3860 3480 3876
rect 3495 3860 3508 3882
rect 3523 3860 3553 3882
rect 3596 3878 3658 3894
rect 3686 3887 3697 3903
rect 3702 3898 3712 3918
rect 3722 3898 3736 3918
rect 3739 3905 3748 3918
rect 3764 3905 3773 3918
rect 3702 3887 3736 3898
rect 3739 3887 3748 3903
rect 3764 3887 3773 3903
rect 3780 3898 3790 3918
rect 3800 3898 3814 3918
rect 3815 3905 3826 3918
rect 3780 3887 3814 3898
rect 3815 3887 3826 3903
rect 3872 3894 3888 3910
rect 3895 3908 3925 3960
rect 3959 3956 3960 3963
rect 3944 3948 3960 3956
rect 3931 3916 3944 3935
rect 3959 3916 3989 3932
rect 3931 3900 4005 3916
rect 3931 3898 3944 3900
rect 3959 3898 3993 3900
rect 3596 3876 3609 3878
rect 3624 3876 3658 3878
rect 3596 3860 3658 3876
rect 3702 3871 3718 3874
rect 3780 3871 3810 3882
rect 3858 3878 3904 3894
rect 3931 3882 4005 3898
rect 3858 3876 3892 3878
rect 3857 3860 3904 3876
rect 3931 3860 3944 3882
rect 3959 3860 3989 3882
rect 4016 3860 4017 3876
rect 4032 3860 4045 4020
rect 4075 3916 4088 4020
rect 4133 3998 4134 4008
rect 4149 3998 4162 4008
rect 4133 3994 4162 3998
rect 4167 3994 4197 4020
rect 4215 4006 4231 4008
rect 4303 4006 4356 4020
rect 4304 4004 4368 4006
rect 4411 4004 4426 4020
rect 4475 4017 4505 4020
rect 4475 4014 4511 4017
rect 4441 4006 4457 4008
rect 4215 3994 4230 3998
rect 4133 3992 4230 3994
rect 4258 3992 4426 4004
rect 4442 3994 4457 3998
rect 4475 3995 4514 4014
rect 4533 4008 4540 4009
rect 4539 4001 4540 4008
rect 4523 3998 4524 4001
rect 4539 3998 4552 4001
rect 4475 3994 4505 3995
rect 4514 3994 4520 3995
rect 4523 3994 4552 3998
rect 4442 3993 4552 3994
rect 4442 3992 4558 3993
rect 4117 3984 4168 3992
rect 4117 3972 4142 3984
rect 4149 3972 4168 3984
rect 4199 3984 4249 3992
rect 4199 3976 4215 3984
rect 4222 3982 4249 3984
rect 4258 3982 4479 3992
rect 4222 3972 4479 3982
rect 4508 3984 4558 3992
rect 4508 3975 4524 3984
rect 4117 3964 4168 3972
rect 4215 3964 4479 3972
rect 4505 3972 4524 3975
rect 4531 3972 4558 3984
rect 4505 3964 4558 3972
rect 4133 3956 4134 3964
rect 4149 3956 4162 3964
rect 4133 3948 4149 3956
rect 4130 3941 4149 3944
rect 4130 3932 4152 3941
rect 4103 3922 4152 3932
rect 4103 3916 4133 3922
rect 4152 3917 4157 3922
rect 4075 3900 4149 3916
rect 4167 3908 4197 3964
rect 4232 3954 4440 3964
rect 4475 3960 4520 3964
rect 4523 3963 4524 3964
rect 4539 3963 4552 3964
rect 4258 3924 4447 3954
rect 4273 3921 4447 3924
rect 4266 3918 4447 3921
rect 4075 3898 4088 3900
rect 4103 3898 4137 3900
rect 4075 3882 4149 3898
rect 4176 3894 4189 3908
rect 4204 3894 4220 3910
rect 4266 3905 4277 3918
rect 4059 3860 4060 3876
rect 4075 3860 4088 3882
rect 4103 3860 4133 3882
rect 4176 3878 4238 3894
rect 4266 3887 4277 3903
rect 4282 3898 4292 3918
rect 4302 3898 4316 3918
rect 4319 3905 4328 3918
rect 4344 3905 4353 3918
rect 4282 3887 4316 3898
rect 4319 3887 4328 3903
rect 4344 3887 4353 3903
rect 4360 3898 4370 3918
rect 4380 3898 4394 3918
rect 4395 3905 4406 3918
rect 4360 3887 4394 3898
rect 4395 3887 4406 3903
rect 4452 3894 4468 3910
rect 4475 3908 4505 3960
rect 4539 3956 4540 3963
rect 4524 3948 4540 3956
rect 4511 3916 4524 3935
rect 4539 3916 4569 3932
rect 4511 3900 4585 3916
rect 4511 3898 4524 3900
rect 4539 3898 4573 3900
rect 4176 3876 4189 3878
rect 4204 3876 4238 3878
rect 4176 3860 4238 3876
rect 4282 3871 4298 3874
rect 4360 3871 4390 3882
rect 4438 3878 4484 3894
rect 4511 3882 4585 3898
rect 4438 3876 4472 3878
rect 4437 3860 4484 3876
rect 4511 3860 4524 3882
rect 4539 3860 4569 3882
rect 4596 3860 4597 3876
rect 4612 3860 4625 4020
rect -7 3852 34 3860
rect -7 3826 8 3852
rect 15 3826 34 3852
rect 98 3848 160 3860
rect 172 3848 247 3860
rect 305 3848 380 3860
rect 392 3848 423 3860
rect 429 3848 464 3860
rect 98 3846 260 3848
rect -7 3818 34 3826
rect 116 3822 129 3846
rect 144 3844 159 3846
rect -1 3808 0 3818
rect 15 3808 28 3818
rect 43 3808 73 3822
rect 116 3808 159 3822
rect 183 3819 190 3826
rect 193 3822 260 3846
rect 292 3846 464 3848
rect 262 3824 290 3828
rect 292 3824 372 3846
rect 393 3844 408 3846
rect 262 3822 372 3824
rect 193 3818 372 3822
rect 166 3808 196 3818
rect 198 3808 351 3818
rect 359 3808 389 3818
rect 393 3808 423 3822
rect 451 3808 464 3846
rect 536 3852 571 3860
rect 536 3826 537 3852
rect 544 3826 571 3852
rect 479 3808 509 3822
rect 536 3818 571 3826
rect 573 3852 614 3860
rect 573 3826 588 3852
rect 595 3826 614 3852
rect 678 3848 740 3860
rect 752 3848 827 3860
rect 885 3848 960 3860
rect 972 3848 1003 3860
rect 1009 3848 1044 3860
rect 678 3846 840 3848
rect 573 3818 614 3826
rect 696 3822 709 3846
rect 724 3844 739 3846
rect 536 3808 537 3818
rect 552 3808 565 3818
rect 579 3808 580 3818
rect 595 3808 608 3818
rect 623 3808 653 3822
rect 696 3808 739 3822
rect 763 3819 770 3826
rect 773 3822 840 3846
rect 872 3846 1044 3848
rect 842 3824 870 3828
rect 872 3824 952 3846
rect 973 3844 988 3846
rect 842 3822 952 3824
rect 773 3818 952 3822
rect 746 3808 776 3818
rect 778 3808 931 3818
rect 939 3808 969 3818
rect 973 3808 1003 3822
rect 1031 3808 1044 3846
rect 1116 3852 1151 3860
rect 1116 3826 1117 3852
rect 1124 3826 1151 3852
rect 1059 3808 1089 3822
rect 1116 3818 1151 3826
rect 1153 3852 1194 3860
rect 1153 3826 1168 3852
rect 1175 3826 1194 3852
rect 1258 3848 1320 3860
rect 1332 3848 1407 3860
rect 1465 3848 1540 3860
rect 1552 3848 1583 3860
rect 1589 3848 1624 3860
rect 1258 3846 1420 3848
rect 1153 3818 1194 3826
rect 1276 3822 1289 3846
rect 1304 3844 1319 3846
rect 1116 3808 1117 3818
rect 1132 3808 1145 3818
rect 1159 3808 1160 3818
rect 1175 3808 1188 3818
rect 1203 3808 1233 3822
rect 1276 3808 1319 3822
rect 1343 3819 1350 3826
rect 1353 3822 1420 3846
rect 1452 3846 1624 3848
rect 1422 3824 1450 3828
rect 1452 3824 1532 3846
rect 1553 3844 1568 3846
rect 1422 3822 1532 3824
rect 1353 3818 1532 3822
rect 1326 3808 1356 3818
rect 1358 3808 1511 3818
rect 1519 3808 1549 3818
rect 1553 3808 1583 3822
rect 1611 3808 1624 3846
rect 1696 3852 1731 3860
rect 1696 3826 1697 3852
rect 1704 3826 1731 3852
rect 1639 3808 1669 3822
rect 1696 3818 1731 3826
rect 1733 3852 1774 3860
rect 1733 3826 1748 3852
rect 1755 3826 1774 3852
rect 1838 3848 1900 3860
rect 1912 3848 1987 3860
rect 2045 3848 2120 3860
rect 2132 3848 2163 3860
rect 2169 3848 2204 3860
rect 1838 3846 2000 3848
rect 1733 3818 1774 3826
rect 1856 3822 1869 3846
rect 1884 3844 1899 3846
rect 1696 3808 1697 3818
rect 1712 3808 1725 3818
rect 1739 3808 1740 3818
rect 1755 3808 1768 3818
rect 1783 3808 1813 3822
rect 1856 3808 1899 3822
rect 1923 3819 1930 3826
rect 1933 3822 2000 3846
rect 2032 3846 2204 3848
rect 2002 3824 2030 3828
rect 2032 3824 2112 3846
rect 2133 3844 2148 3846
rect 2002 3822 2112 3824
rect 1933 3818 2112 3822
rect 1906 3808 1936 3818
rect 1938 3808 2091 3818
rect 2099 3808 2129 3818
rect 2133 3808 2163 3822
rect 2191 3808 2204 3846
rect 2276 3852 2311 3860
rect 2276 3826 2277 3852
rect 2284 3826 2311 3852
rect 2219 3808 2249 3822
rect 2276 3818 2311 3826
rect 2313 3852 2354 3860
rect 2313 3826 2328 3852
rect 2335 3826 2354 3852
rect 2418 3848 2480 3860
rect 2492 3848 2567 3860
rect 2625 3848 2700 3860
rect 2712 3848 2743 3860
rect 2749 3848 2784 3860
rect 2418 3846 2580 3848
rect 2313 3818 2354 3826
rect 2436 3822 2449 3846
rect 2464 3844 2479 3846
rect 2276 3808 2277 3818
rect 2292 3808 2305 3818
rect 2319 3808 2320 3818
rect 2335 3808 2348 3818
rect 2363 3808 2393 3822
rect 2436 3808 2479 3822
rect 2503 3819 2510 3826
rect 2513 3822 2580 3846
rect 2612 3846 2784 3848
rect 2582 3824 2610 3828
rect 2612 3824 2692 3846
rect 2713 3844 2728 3846
rect 2582 3822 2692 3824
rect 2513 3818 2692 3822
rect 2486 3808 2516 3818
rect 2518 3808 2671 3818
rect 2679 3808 2709 3818
rect 2713 3808 2743 3822
rect 2771 3808 2784 3846
rect 2856 3852 2891 3860
rect 2856 3826 2857 3852
rect 2864 3826 2891 3852
rect 2799 3808 2829 3822
rect 2856 3818 2891 3826
rect 2893 3852 2934 3860
rect 2893 3826 2908 3852
rect 2915 3826 2934 3852
rect 2998 3848 3060 3860
rect 3072 3848 3147 3860
rect 3205 3848 3280 3860
rect 3292 3848 3323 3860
rect 3329 3848 3364 3860
rect 2998 3846 3160 3848
rect 2893 3818 2934 3826
rect 3016 3822 3029 3846
rect 3044 3844 3059 3846
rect 2856 3808 2857 3818
rect 2872 3808 2885 3818
rect 2899 3808 2900 3818
rect 2915 3808 2928 3818
rect 2943 3808 2973 3822
rect 3016 3808 3059 3822
rect 3083 3819 3090 3826
rect 3093 3822 3160 3846
rect 3192 3846 3364 3848
rect 3162 3824 3190 3828
rect 3192 3824 3272 3846
rect 3293 3844 3308 3846
rect 3162 3822 3272 3824
rect 3093 3818 3272 3822
rect 3066 3808 3096 3818
rect 3098 3808 3251 3818
rect 3259 3808 3289 3818
rect 3293 3808 3323 3822
rect 3351 3808 3364 3846
rect 3436 3852 3471 3860
rect 3436 3826 3437 3852
rect 3444 3826 3471 3852
rect 3379 3808 3409 3822
rect 3436 3818 3471 3826
rect 3473 3852 3514 3860
rect 3473 3826 3488 3852
rect 3495 3826 3514 3852
rect 3578 3848 3640 3860
rect 3652 3848 3727 3860
rect 3785 3848 3860 3860
rect 3872 3848 3903 3860
rect 3909 3848 3944 3860
rect 3578 3846 3740 3848
rect 3473 3818 3514 3826
rect 3596 3822 3609 3846
rect 3624 3844 3639 3846
rect 3436 3808 3437 3818
rect 3452 3808 3465 3818
rect 3479 3808 3480 3818
rect 3495 3808 3508 3818
rect 3523 3808 3553 3822
rect 3596 3808 3639 3822
rect 3663 3819 3670 3826
rect 3673 3822 3740 3846
rect 3772 3846 3944 3848
rect 3742 3824 3770 3828
rect 3772 3824 3852 3846
rect 3873 3844 3888 3846
rect 3742 3822 3852 3824
rect 3673 3818 3852 3822
rect 3646 3808 3676 3818
rect 3678 3808 3831 3818
rect 3839 3808 3869 3818
rect 3873 3808 3903 3822
rect 3931 3808 3944 3846
rect 4016 3852 4051 3860
rect 4016 3826 4017 3852
rect 4024 3826 4051 3852
rect 3959 3808 3989 3822
rect 4016 3818 4051 3826
rect 4053 3852 4094 3860
rect 4053 3826 4068 3852
rect 4075 3826 4094 3852
rect 4158 3848 4220 3860
rect 4232 3848 4307 3860
rect 4365 3848 4440 3860
rect 4452 3848 4483 3860
rect 4489 3848 4524 3860
rect 4158 3846 4320 3848
rect 4053 3818 4094 3826
rect 4176 3822 4189 3846
rect 4204 3844 4219 3846
rect 4016 3808 4017 3818
rect 4032 3808 4045 3818
rect 4059 3808 4060 3818
rect 4075 3808 4088 3818
rect 4103 3808 4133 3822
rect 4176 3808 4219 3822
rect 4243 3819 4250 3826
rect 4253 3822 4320 3846
rect 4352 3846 4524 3848
rect 4322 3824 4350 3828
rect 4352 3824 4432 3846
rect 4453 3844 4468 3846
rect 4322 3822 4432 3824
rect 4253 3818 4432 3822
rect 4226 3808 4256 3818
rect 4258 3808 4411 3818
rect 4419 3808 4449 3818
rect 4453 3808 4483 3822
rect 4511 3808 4524 3846
rect 4596 3852 4631 3860
rect 4596 3826 4597 3852
rect 4604 3826 4631 3852
rect 4539 3808 4569 3822
rect 4596 3818 4631 3826
rect 4596 3808 4597 3818
rect 4612 3808 4625 3818
rect -1 3802 4625 3808
rect 0 3794 4625 3802
rect 15 3764 28 3794
rect 43 3776 73 3794
rect 116 3780 130 3794
rect 166 3780 386 3794
rect 117 3778 130 3780
rect 83 3766 98 3778
rect 80 3764 102 3766
rect 107 3764 137 3778
rect 198 3776 351 3780
rect 180 3764 372 3776
rect 415 3764 445 3778
rect 451 3764 464 3794
rect 479 3776 509 3794
rect 552 3764 565 3794
rect 595 3764 608 3794
rect 623 3776 653 3794
rect 696 3780 710 3794
rect 746 3780 966 3794
rect 697 3778 710 3780
rect 663 3766 678 3778
rect 660 3764 682 3766
rect 687 3764 717 3778
rect 778 3776 931 3780
rect 760 3764 952 3776
rect 995 3764 1025 3778
rect 1031 3764 1044 3794
rect 1059 3776 1089 3794
rect 1132 3764 1145 3794
rect 1175 3764 1188 3794
rect 1203 3776 1233 3794
rect 1276 3780 1290 3794
rect 1326 3780 1546 3794
rect 1277 3778 1290 3780
rect 1243 3766 1258 3778
rect 1240 3764 1262 3766
rect 1267 3764 1297 3778
rect 1358 3776 1511 3780
rect 1340 3764 1532 3776
rect 1575 3764 1605 3778
rect 1611 3764 1624 3794
rect 1639 3776 1669 3794
rect 1712 3764 1725 3794
rect 1755 3764 1768 3794
rect 1783 3776 1813 3794
rect 1856 3780 1870 3794
rect 1906 3780 2126 3794
rect 1857 3778 1870 3780
rect 1823 3766 1838 3778
rect 1820 3764 1842 3766
rect 1847 3764 1877 3778
rect 1938 3776 2091 3780
rect 1920 3764 2112 3776
rect 2155 3764 2185 3778
rect 2191 3764 2204 3794
rect 2219 3776 2249 3794
rect 2292 3764 2305 3794
rect 2335 3764 2348 3794
rect 2363 3776 2393 3794
rect 2436 3780 2450 3794
rect 2486 3780 2706 3794
rect 2437 3778 2450 3780
rect 2403 3766 2418 3778
rect 2400 3764 2422 3766
rect 2427 3764 2457 3778
rect 2518 3776 2671 3780
rect 2500 3764 2692 3776
rect 2735 3764 2765 3778
rect 2771 3764 2784 3794
rect 2799 3776 2829 3794
rect 2872 3764 2885 3794
rect 2915 3764 2928 3794
rect 2943 3776 2973 3794
rect 3016 3780 3030 3794
rect 3066 3780 3286 3794
rect 3017 3778 3030 3780
rect 2983 3766 2998 3778
rect 2980 3764 3002 3766
rect 3007 3764 3037 3778
rect 3098 3776 3251 3780
rect 3080 3764 3272 3776
rect 3315 3764 3345 3778
rect 3351 3764 3364 3794
rect 3379 3776 3409 3794
rect 3452 3764 3465 3794
rect 3495 3764 3508 3794
rect 3523 3776 3553 3794
rect 3596 3780 3610 3794
rect 3646 3780 3866 3794
rect 3597 3778 3610 3780
rect 3563 3766 3578 3778
rect 3560 3764 3582 3766
rect 3587 3764 3617 3778
rect 3678 3776 3831 3780
rect 3660 3764 3852 3776
rect 3895 3764 3925 3778
rect 3931 3764 3944 3794
rect 3959 3776 3989 3794
rect 4032 3764 4045 3794
rect 4075 3764 4088 3794
rect 4103 3776 4133 3794
rect 4176 3780 4190 3794
rect 4226 3780 4446 3794
rect 4177 3778 4190 3780
rect 4143 3766 4158 3778
rect 4140 3764 4162 3766
rect 4167 3764 4197 3778
rect 4258 3776 4411 3780
rect 4240 3764 4432 3776
rect 4475 3764 4505 3778
rect 4511 3764 4524 3794
rect 4539 3776 4569 3794
rect 4612 3764 4625 3794
rect 0 3750 4625 3764
rect 15 3646 28 3750
rect 73 3728 74 3738
rect 89 3728 102 3738
rect 73 3724 102 3728
rect 107 3724 137 3750
rect 155 3736 171 3738
rect 243 3736 296 3750
rect 244 3734 308 3736
rect 351 3734 366 3750
rect 415 3747 445 3750
rect 415 3744 451 3747
rect 381 3736 397 3738
rect 155 3724 170 3728
rect 73 3722 170 3724
rect 198 3722 366 3734
rect 382 3724 397 3728
rect 415 3725 454 3744
rect 473 3738 480 3739
rect 479 3731 480 3738
rect 463 3728 464 3731
rect 479 3728 492 3731
rect 415 3724 445 3725
rect 454 3724 460 3725
rect 463 3724 492 3728
rect 382 3723 492 3724
rect 382 3722 498 3723
rect 57 3714 108 3722
rect 57 3702 82 3714
rect 89 3702 108 3714
rect 139 3714 189 3722
rect 139 3706 155 3714
rect 162 3712 189 3714
rect 198 3712 419 3722
rect 162 3702 419 3712
rect 448 3714 498 3722
rect 448 3705 464 3714
rect 57 3694 108 3702
rect 155 3694 419 3702
rect 445 3702 464 3705
rect 471 3702 498 3714
rect 445 3694 498 3702
rect 73 3686 74 3694
rect 89 3686 102 3694
rect 73 3678 89 3686
rect 70 3671 89 3674
rect 70 3662 92 3671
rect 43 3652 92 3662
rect 43 3646 73 3652
rect 92 3647 97 3652
rect 15 3630 89 3646
rect 107 3638 137 3694
rect 172 3684 380 3694
rect 415 3690 460 3694
rect 463 3693 464 3694
rect 479 3693 492 3694
rect 198 3654 387 3684
rect 213 3651 387 3654
rect 206 3648 387 3651
rect 15 3628 28 3630
rect 43 3628 77 3630
rect 15 3612 89 3628
rect 116 3624 129 3638
rect 144 3624 160 3640
rect 206 3635 217 3648
rect -1 3590 0 3606
rect 15 3590 28 3612
rect 43 3590 73 3612
rect 116 3608 178 3624
rect 206 3617 217 3633
rect 222 3628 232 3648
rect 242 3628 256 3648
rect 259 3635 268 3648
rect 284 3635 293 3648
rect 222 3617 256 3628
rect 259 3617 268 3633
rect 284 3617 293 3633
rect 300 3628 310 3648
rect 320 3628 334 3648
rect 335 3635 346 3648
rect 300 3617 334 3628
rect 335 3617 346 3633
rect 392 3624 408 3640
rect 415 3638 445 3690
rect 479 3686 480 3693
rect 464 3678 480 3686
rect 451 3646 464 3665
rect 479 3646 509 3662
rect 451 3630 525 3646
rect 451 3628 464 3630
rect 479 3628 513 3630
rect 116 3606 129 3608
rect 144 3606 178 3608
rect 116 3590 178 3606
rect 222 3601 238 3604
rect 300 3601 330 3612
rect 378 3608 424 3624
rect 451 3612 525 3628
rect 378 3606 412 3608
rect 377 3590 424 3606
rect 451 3590 464 3612
rect 479 3590 509 3612
rect 536 3590 537 3606
rect 552 3590 565 3750
rect 595 3646 608 3750
rect 653 3728 654 3738
rect 669 3728 682 3738
rect 653 3724 682 3728
rect 687 3724 717 3750
rect 735 3736 751 3738
rect 823 3736 876 3750
rect 824 3734 888 3736
rect 931 3734 946 3750
rect 995 3747 1025 3750
rect 995 3744 1031 3747
rect 961 3736 977 3738
rect 735 3724 750 3728
rect 653 3722 750 3724
rect 778 3722 946 3734
rect 962 3724 977 3728
rect 995 3725 1034 3744
rect 1053 3738 1060 3739
rect 1059 3731 1060 3738
rect 1043 3728 1044 3731
rect 1059 3728 1072 3731
rect 995 3724 1025 3725
rect 1034 3724 1040 3725
rect 1043 3724 1072 3728
rect 962 3723 1072 3724
rect 962 3722 1078 3723
rect 637 3714 688 3722
rect 637 3702 662 3714
rect 669 3702 688 3714
rect 719 3714 769 3722
rect 719 3706 735 3714
rect 742 3712 769 3714
rect 778 3712 999 3722
rect 742 3702 999 3712
rect 1028 3714 1078 3722
rect 1028 3705 1044 3714
rect 637 3694 688 3702
rect 735 3694 999 3702
rect 1025 3702 1044 3705
rect 1051 3702 1078 3714
rect 1025 3694 1078 3702
rect 653 3686 654 3694
rect 669 3686 682 3694
rect 653 3678 669 3686
rect 650 3671 669 3674
rect 650 3662 672 3671
rect 623 3652 672 3662
rect 623 3646 653 3652
rect 672 3647 677 3652
rect 595 3630 669 3646
rect 687 3638 717 3694
rect 752 3684 960 3694
rect 995 3690 1040 3694
rect 1043 3693 1044 3694
rect 1059 3693 1072 3694
rect 778 3654 967 3684
rect 793 3651 967 3654
rect 786 3648 967 3651
rect 595 3628 608 3630
rect 623 3628 657 3630
rect 595 3612 669 3628
rect 696 3624 709 3638
rect 724 3624 740 3640
rect 786 3635 797 3648
rect 579 3590 580 3606
rect 595 3590 608 3612
rect 623 3590 653 3612
rect 696 3608 758 3624
rect 786 3617 797 3633
rect 802 3628 812 3648
rect 822 3628 836 3648
rect 839 3635 848 3648
rect 864 3635 873 3648
rect 802 3617 836 3628
rect 839 3617 848 3633
rect 864 3617 873 3633
rect 880 3628 890 3648
rect 900 3628 914 3648
rect 915 3635 926 3648
rect 880 3617 914 3628
rect 915 3617 926 3633
rect 972 3624 988 3640
rect 995 3638 1025 3690
rect 1059 3686 1060 3693
rect 1044 3678 1060 3686
rect 1031 3646 1044 3665
rect 1059 3646 1089 3662
rect 1031 3630 1105 3646
rect 1031 3628 1044 3630
rect 1059 3628 1093 3630
rect 696 3606 709 3608
rect 724 3606 758 3608
rect 696 3590 758 3606
rect 802 3601 818 3604
rect 880 3601 910 3612
rect 958 3608 1004 3624
rect 1031 3612 1105 3628
rect 958 3606 992 3608
rect 957 3590 1004 3606
rect 1031 3590 1044 3612
rect 1059 3590 1089 3612
rect 1116 3590 1117 3606
rect 1132 3590 1145 3750
rect 1175 3646 1188 3750
rect 1233 3728 1234 3738
rect 1249 3728 1262 3738
rect 1233 3724 1262 3728
rect 1267 3724 1297 3750
rect 1315 3736 1331 3738
rect 1403 3736 1456 3750
rect 1404 3734 1468 3736
rect 1511 3734 1526 3750
rect 1575 3747 1605 3750
rect 1575 3744 1611 3747
rect 1541 3736 1557 3738
rect 1315 3724 1330 3728
rect 1233 3722 1330 3724
rect 1358 3722 1526 3734
rect 1542 3724 1557 3728
rect 1575 3725 1614 3744
rect 1633 3738 1640 3739
rect 1639 3731 1640 3738
rect 1623 3728 1624 3731
rect 1639 3728 1652 3731
rect 1575 3724 1605 3725
rect 1614 3724 1620 3725
rect 1623 3724 1652 3728
rect 1542 3723 1652 3724
rect 1542 3722 1658 3723
rect 1217 3714 1268 3722
rect 1217 3702 1242 3714
rect 1249 3702 1268 3714
rect 1299 3714 1349 3722
rect 1299 3706 1315 3714
rect 1322 3712 1349 3714
rect 1358 3712 1579 3722
rect 1322 3702 1579 3712
rect 1608 3714 1658 3722
rect 1608 3705 1624 3714
rect 1217 3694 1268 3702
rect 1315 3694 1579 3702
rect 1605 3702 1624 3705
rect 1631 3702 1658 3714
rect 1605 3694 1658 3702
rect 1233 3686 1234 3694
rect 1249 3686 1262 3694
rect 1233 3678 1249 3686
rect 1230 3671 1249 3674
rect 1230 3662 1252 3671
rect 1203 3652 1252 3662
rect 1203 3646 1233 3652
rect 1252 3647 1257 3652
rect 1175 3630 1249 3646
rect 1267 3638 1297 3694
rect 1332 3684 1540 3694
rect 1575 3690 1620 3694
rect 1623 3693 1624 3694
rect 1639 3693 1652 3694
rect 1358 3654 1547 3684
rect 1373 3651 1547 3654
rect 1366 3648 1547 3651
rect 1175 3628 1188 3630
rect 1203 3628 1237 3630
rect 1175 3612 1249 3628
rect 1276 3624 1289 3638
rect 1304 3624 1320 3640
rect 1366 3635 1377 3648
rect 1159 3590 1160 3606
rect 1175 3590 1188 3612
rect 1203 3590 1233 3612
rect 1276 3608 1338 3624
rect 1366 3617 1377 3633
rect 1382 3628 1392 3648
rect 1402 3628 1416 3648
rect 1419 3635 1428 3648
rect 1444 3635 1453 3648
rect 1382 3617 1416 3628
rect 1419 3617 1428 3633
rect 1444 3617 1453 3633
rect 1460 3628 1470 3648
rect 1480 3628 1494 3648
rect 1495 3635 1506 3648
rect 1460 3617 1494 3628
rect 1495 3617 1506 3633
rect 1552 3624 1568 3640
rect 1575 3638 1605 3690
rect 1639 3686 1640 3693
rect 1624 3678 1640 3686
rect 1611 3646 1624 3665
rect 1639 3646 1669 3662
rect 1611 3630 1685 3646
rect 1611 3628 1624 3630
rect 1639 3628 1673 3630
rect 1276 3606 1289 3608
rect 1304 3606 1338 3608
rect 1276 3590 1338 3606
rect 1382 3601 1398 3604
rect 1460 3601 1490 3612
rect 1538 3608 1584 3624
rect 1611 3612 1685 3628
rect 1538 3606 1572 3608
rect 1537 3590 1584 3606
rect 1611 3590 1624 3612
rect 1639 3590 1669 3612
rect 1696 3590 1697 3606
rect 1712 3590 1725 3750
rect 1755 3646 1768 3750
rect 1813 3728 1814 3738
rect 1829 3728 1842 3738
rect 1813 3724 1842 3728
rect 1847 3724 1877 3750
rect 1895 3736 1911 3738
rect 1983 3736 2036 3750
rect 1984 3734 2048 3736
rect 2091 3734 2106 3750
rect 2155 3747 2185 3750
rect 2155 3744 2191 3747
rect 2121 3736 2137 3738
rect 1895 3724 1910 3728
rect 1813 3722 1910 3724
rect 1938 3722 2106 3734
rect 2122 3724 2137 3728
rect 2155 3725 2194 3744
rect 2213 3738 2220 3739
rect 2219 3731 2220 3738
rect 2203 3728 2204 3731
rect 2219 3728 2232 3731
rect 2155 3724 2185 3725
rect 2194 3724 2200 3725
rect 2203 3724 2232 3728
rect 2122 3723 2232 3724
rect 2122 3722 2238 3723
rect 1797 3714 1848 3722
rect 1797 3702 1822 3714
rect 1829 3702 1848 3714
rect 1879 3714 1929 3722
rect 1879 3706 1895 3714
rect 1902 3712 1929 3714
rect 1938 3712 2159 3722
rect 1902 3702 2159 3712
rect 2188 3714 2238 3722
rect 2188 3705 2204 3714
rect 1797 3694 1848 3702
rect 1895 3694 2159 3702
rect 2185 3702 2204 3705
rect 2211 3702 2238 3714
rect 2185 3694 2238 3702
rect 1813 3686 1814 3694
rect 1829 3686 1842 3694
rect 1813 3678 1829 3686
rect 1810 3671 1829 3674
rect 1810 3662 1832 3671
rect 1783 3652 1832 3662
rect 1783 3646 1813 3652
rect 1832 3647 1837 3652
rect 1755 3630 1829 3646
rect 1847 3638 1877 3694
rect 1912 3684 2120 3694
rect 2155 3690 2200 3694
rect 2203 3693 2204 3694
rect 2219 3693 2232 3694
rect 1938 3654 2127 3684
rect 1953 3651 2127 3654
rect 1946 3648 2127 3651
rect 1755 3628 1768 3630
rect 1783 3628 1817 3630
rect 1755 3612 1829 3628
rect 1856 3624 1869 3638
rect 1884 3624 1900 3640
rect 1946 3635 1957 3648
rect 1739 3590 1740 3606
rect 1755 3590 1768 3612
rect 1783 3590 1813 3612
rect 1856 3608 1918 3624
rect 1946 3617 1957 3633
rect 1962 3628 1972 3648
rect 1982 3628 1996 3648
rect 1999 3635 2008 3648
rect 2024 3635 2033 3648
rect 1962 3617 1996 3628
rect 1999 3617 2008 3633
rect 2024 3617 2033 3633
rect 2040 3628 2050 3648
rect 2060 3628 2074 3648
rect 2075 3635 2086 3648
rect 2040 3617 2074 3628
rect 2075 3617 2086 3633
rect 2132 3624 2148 3640
rect 2155 3638 2185 3690
rect 2219 3686 2220 3693
rect 2204 3678 2220 3686
rect 2191 3646 2204 3665
rect 2219 3646 2249 3662
rect 2191 3630 2265 3646
rect 2191 3628 2204 3630
rect 2219 3628 2253 3630
rect 1856 3606 1869 3608
rect 1884 3606 1918 3608
rect 1856 3590 1918 3606
rect 1962 3601 1978 3604
rect 2040 3601 2070 3612
rect 2118 3608 2164 3624
rect 2191 3612 2265 3628
rect 2118 3606 2152 3608
rect 2117 3590 2164 3606
rect 2191 3590 2204 3612
rect 2219 3590 2249 3612
rect 2276 3590 2277 3606
rect 2292 3590 2305 3750
rect 2335 3646 2348 3750
rect 2393 3728 2394 3738
rect 2409 3728 2422 3738
rect 2393 3724 2422 3728
rect 2427 3724 2457 3750
rect 2475 3736 2491 3738
rect 2563 3736 2616 3750
rect 2564 3734 2628 3736
rect 2671 3734 2686 3750
rect 2735 3747 2765 3750
rect 2735 3744 2771 3747
rect 2701 3736 2717 3738
rect 2475 3724 2490 3728
rect 2393 3722 2490 3724
rect 2518 3722 2686 3734
rect 2702 3724 2717 3728
rect 2735 3725 2774 3744
rect 2793 3738 2800 3739
rect 2799 3731 2800 3738
rect 2783 3728 2784 3731
rect 2799 3728 2812 3731
rect 2735 3724 2765 3725
rect 2774 3724 2780 3725
rect 2783 3724 2812 3728
rect 2702 3723 2812 3724
rect 2702 3722 2818 3723
rect 2377 3714 2428 3722
rect 2377 3702 2402 3714
rect 2409 3702 2428 3714
rect 2459 3714 2509 3722
rect 2459 3706 2475 3714
rect 2482 3712 2509 3714
rect 2518 3712 2739 3722
rect 2482 3702 2739 3712
rect 2768 3714 2818 3722
rect 2768 3705 2784 3714
rect 2377 3694 2428 3702
rect 2475 3694 2739 3702
rect 2765 3702 2784 3705
rect 2791 3702 2818 3714
rect 2765 3694 2818 3702
rect 2393 3686 2394 3694
rect 2409 3686 2422 3694
rect 2393 3678 2409 3686
rect 2390 3671 2409 3674
rect 2390 3662 2412 3671
rect 2363 3652 2412 3662
rect 2363 3646 2393 3652
rect 2412 3647 2417 3652
rect 2335 3630 2409 3646
rect 2427 3638 2457 3694
rect 2492 3684 2700 3694
rect 2735 3690 2780 3694
rect 2783 3693 2784 3694
rect 2799 3693 2812 3694
rect 2518 3654 2707 3684
rect 2533 3651 2707 3654
rect 2526 3648 2707 3651
rect 2335 3628 2348 3630
rect 2363 3628 2397 3630
rect 2335 3612 2409 3628
rect 2436 3624 2449 3638
rect 2464 3624 2480 3640
rect 2526 3635 2537 3648
rect 2319 3590 2320 3606
rect 2335 3590 2348 3612
rect 2363 3590 2393 3612
rect 2436 3608 2498 3624
rect 2526 3617 2537 3633
rect 2542 3628 2552 3648
rect 2562 3628 2576 3648
rect 2579 3635 2588 3648
rect 2604 3635 2613 3648
rect 2542 3617 2576 3628
rect 2579 3617 2588 3633
rect 2604 3617 2613 3633
rect 2620 3628 2630 3648
rect 2640 3628 2654 3648
rect 2655 3635 2666 3648
rect 2620 3617 2654 3628
rect 2655 3617 2666 3633
rect 2712 3624 2728 3640
rect 2735 3638 2765 3690
rect 2799 3686 2800 3693
rect 2784 3678 2800 3686
rect 2771 3646 2784 3665
rect 2799 3646 2829 3662
rect 2771 3630 2845 3646
rect 2771 3628 2784 3630
rect 2799 3628 2833 3630
rect 2436 3606 2449 3608
rect 2464 3606 2498 3608
rect 2436 3590 2498 3606
rect 2542 3601 2558 3604
rect 2620 3601 2650 3612
rect 2698 3608 2744 3624
rect 2771 3612 2845 3628
rect 2698 3606 2732 3608
rect 2697 3590 2744 3606
rect 2771 3590 2784 3612
rect 2799 3590 2829 3612
rect 2856 3590 2857 3606
rect 2872 3590 2885 3750
rect 2915 3646 2928 3750
rect 2973 3728 2974 3738
rect 2989 3728 3002 3738
rect 2973 3724 3002 3728
rect 3007 3724 3037 3750
rect 3055 3736 3071 3738
rect 3143 3736 3196 3750
rect 3144 3734 3208 3736
rect 3251 3734 3266 3750
rect 3315 3747 3345 3750
rect 3315 3744 3351 3747
rect 3281 3736 3297 3738
rect 3055 3724 3070 3728
rect 2973 3722 3070 3724
rect 3098 3722 3266 3734
rect 3282 3724 3297 3728
rect 3315 3725 3354 3744
rect 3373 3738 3380 3739
rect 3379 3731 3380 3738
rect 3363 3728 3364 3731
rect 3379 3728 3392 3731
rect 3315 3724 3345 3725
rect 3354 3724 3360 3725
rect 3363 3724 3392 3728
rect 3282 3723 3392 3724
rect 3282 3722 3398 3723
rect 2957 3714 3008 3722
rect 2957 3702 2982 3714
rect 2989 3702 3008 3714
rect 3039 3714 3089 3722
rect 3039 3706 3055 3714
rect 3062 3712 3089 3714
rect 3098 3712 3319 3722
rect 3062 3702 3319 3712
rect 3348 3714 3398 3722
rect 3348 3705 3364 3714
rect 2957 3694 3008 3702
rect 3055 3694 3319 3702
rect 3345 3702 3364 3705
rect 3371 3702 3398 3714
rect 3345 3694 3398 3702
rect 2973 3686 2974 3694
rect 2989 3686 3002 3694
rect 2973 3678 2989 3686
rect 2970 3671 2989 3674
rect 2970 3662 2992 3671
rect 2943 3652 2992 3662
rect 2943 3646 2973 3652
rect 2992 3647 2997 3652
rect 2915 3630 2989 3646
rect 3007 3638 3037 3694
rect 3072 3684 3280 3694
rect 3315 3690 3360 3694
rect 3363 3693 3364 3694
rect 3379 3693 3392 3694
rect 3098 3654 3287 3684
rect 3113 3651 3287 3654
rect 3106 3648 3287 3651
rect 2915 3628 2928 3630
rect 2943 3628 2977 3630
rect 2915 3612 2989 3628
rect 3016 3624 3029 3638
rect 3044 3624 3060 3640
rect 3106 3635 3117 3648
rect 2899 3590 2900 3606
rect 2915 3590 2928 3612
rect 2943 3590 2973 3612
rect 3016 3608 3078 3624
rect 3106 3617 3117 3633
rect 3122 3628 3132 3648
rect 3142 3628 3156 3648
rect 3159 3635 3168 3648
rect 3184 3635 3193 3648
rect 3122 3617 3156 3628
rect 3159 3617 3168 3633
rect 3184 3617 3193 3633
rect 3200 3628 3210 3648
rect 3220 3628 3234 3648
rect 3235 3635 3246 3648
rect 3200 3617 3234 3628
rect 3235 3617 3246 3633
rect 3292 3624 3308 3640
rect 3315 3638 3345 3690
rect 3379 3686 3380 3693
rect 3364 3678 3380 3686
rect 3351 3646 3364 3665
rect 3379 3646 3409 3662
rect 3351 3630 3425 3646
rect 3351 3628 3364 3630
rect 3379 3628 3413 3630
rect 3016 3606 3029 3608
rect 3044 3606 3078 3608
rect 3016 3590 3078 3606
rect 3122 3601 3138 3604
rect 3200 3601 3230 3612
rect 3278 3608 3324 3624
rect 3351 3612 3425 3628
rect 3278 3606 3312 3608
rect 3277 3590 3324 3606
rect 3351 3590 3364 3612
rect 3379 3590 3409 3612
rect 3436 3590 3437 3606
rect 3452 3590 3465 3750
rect 3495 3646 3508 3750
rect 3553 3728 3554 3738
rect 3569 3728 3582 3738
rect 3553 3724 3582 3728
rect 3587 3724 3617 3750
rect 3635 3736 3651 3738
rect 3723 3736 3776 3750
rect 3724 3734 3788 3736
rect 3831 3734 3846 3750
rect 3895 3747 3925 3750
rect 3895 3744 3931 3747
rect 3861 3736 3877 3738
rect 3635 3724 3650 3728
rect 3553 3722 3650 3724
rect 3678 3722 3846 3734
rect 3862 3724 3877 3728
rect 3895 3725 3934 3744
rect 3953 3738 3960 3739
rect 3959 3731 3960 3738
rect 3943 3728 3944 3731
rect 3959 3728 3972 3731
rect 3895 3724 3925 3725
rect 3934 3724 3940 3725
rect 3943 3724 3972 3728
rect 3862 3723 3972 3724
rect 3862 3722 3978 3723
rect 3537 3714 3588 3722
rect 3537 3702 3562 3714
rect 3569 3702 3588 3714
rect 3619 3714 3669 3722
rect 3619 3706 3635 3714
rect 3642 3712 3669 3714
rect 3678 3712 3899 3722
rect 3642 3702 3899 3712
rect 3928 3714 3978 3722
rect 3928 3705 3944 3714
rect 3537 3694 3588 3702
rect 3635 3694 3899 3702
rect 3925 3702 3944 3705
rect 3951 3702 3978 3714
rect 3925 3694 3978 3702
rect 3553 3686 3554 3694
rect 3569 3686 3582 3694
rect 3553 3678 3569 3686
rect 3550 3671 3569 3674
rect 3550 3662 3572 3671
rect 3523 3652 3572 3662
rect 3523 3646 3553 3652
rect 3572 3647 3577 3652
rect 3495 3630 3569 3646
rect 3587 3638 3617 3694
rect 3652 3684 3860 3694
rect 3895 3690 3940 3694
rect 3943 3693 3944 3694
rect 3959 3693 3972 3694
rect 3678 3654 3867 3684
rect 3693 3651 3867 3654
rect 3686 3648 3867 3651
rect 3495 3628 3508 3630
rect 3523 3628 3557 3630
rect 3495 3612 3569 3628
rect 3596 3624 3609 3638
rect 3624 3624 3640 3640
rect 3686 3635 3697 3648
rect 3479 3590 3480 3606
rect 3495 3590 3508 3612
rect 3523 3590 3553 3612
rect 3596 3608 3658 3624
rect 3686 3617 3697 3633
rect 3702 3628 3712 3648
rect 3722 3628 3736 3648
rect 3739 3635 3748 3648
rect 3764 3635 3773 3648
rect 3702 3617 3736 3628
rect 3739 3617 3748 3633
rect 3764 3617 3773 3633
rect 3780 3628 3790 3648
rect 3800 3628 3814 3648
rect 3815 3635 3826 3648
rect 3780 3617 3814 3628
rect 3815 3617 3826 3633
rect 3872 3624 3888 3640
rect 3895 3638 3925 3690
rect 3959 3686 3960 3693
rect 3944 3678 3960 3686
rect 3931 3646 3944 3665
rect 3959 3646 3989 3662
rect 3931 3630 4005 3646
rect 3931 3628 3944 3630
rect 3959 3628 3993 3630
rect 3596 3606 3609 3608
rect 3624 3606 3658 3608
rect 3596 3590 3658 3606
rect 3702 3601 3718 3604
rect 3780 3601 3810 3612
rect 3858 3608 3904 3624
rect 3931 3612 4005 3628
rect 3858 3606 3892 3608
rect 3857 3590 3904 3606
rect 3931 3590 3944 3612
rect 3959 3590 3989 3612
rect 4016 3590 4017 3606
rect 4032 3590 4045 3750
rect 4075 3646 4088 3750
rect 4133 3728 4134 3738
rect 4149 3728 4162 3738
rect 4133 3724 4162 3728
rect 4167 3724 4197 3750
rect 4215 3736 4231 3738
rect 4303 3736 4356 3750
rect 4304 3734 4368 3736
rect 4411 3734 4426 3750
rect 4475 3747 4505 3750
rect 4475 3744 4511 3747
rect 4441 3736 4457 3738
rect 4215 3724 4230 3728
rect 4133 3722 4230 3724
rect 4258 3722 4426 3734
rect 4442 3724 4457 3728
rect 4475 3725 4514 3744
rect 4533 3738 4540 3739
rect 4539 3731 4540 3738
rect 4523 3728 4524 3731
rect 4539 3728 4552 3731
rect 4475 3724 4505 3725
rect 4514 3724 4520 3725
rect 4523 3724 4552 3728
rect 4442 3723 4552 3724
rect 4442 3722 4558 3723
rect 4117 3714 4168 3722
rect 4117 3702 4142 3714
rect 4149 3702 4168 3714
rect 4199 3714 4249 3722
rect 4199 3706 4215 3714
rect 4222 3712 4249 3714
rect 4258 3712 4479 3722
rect 4222 3702 4479 3712
rect 4508 3714 4558 3722
rect 4508 3705 4524 3714
rect 4117 3694 4168 3702
rect 4215 3694 4479 3702
rect 4505 3702 4524 3705
rect 4531 3702 4558 3714
rect 4505 3694 4558 3702
rect 4133 3686 4134 3694
rect 4149 3686 4162 3694
rect 4133 3678 4149 3686
rect 4130 3671 4149 3674
rect 4130 3662 4152 3671
rect 4103 3652 4152 3662
rect 4103 3646 4133 3652
rect 4152 3647 4157 3652
rect 4075 3630 4149 3646
rect 4167 3638 4197 3694
rect 4232 3684 4440 3694
rect 4475 3690 4520 3694
rect 4523 3693 4524 3694
rect 4539 3693 4552 3694
rect 4258 3654 4447 3684
rect 4273 3651 4447 3654
rect 4266 3648 4447 3651
rect 4075 3628 4088 3630
rect 4103 3628 4137 3630
rect 4075 3612 4149 3628
rect 4176 3624 4189 3638
rect 4204 3624 4220 3640
rect 4266 3635 4277 3648
rect 4059 3590 4060 3606
rect 4075 3590 4088 3612
rect 4103 3590 4133 3612
rect 4176 3608 4238 3624
rect 4266 3617 4277 3633
rect 4282 3628 4292 3648
rect 4302 3628 4316 3648
rect 4319 3635 4328 3648
rect 4344 3635 4353 3648
rect 4282 3617 4316 3628
rect 4319 3617 4328 3633
rect 4344 3617 4353 3633
rect 4360 3628 4370 3648
rect 4380 3628 4394 3648
rect 4395 3635 4406 3648
rect 4360 3617 4394 3628
rect 4395 3617 4406 3633
rect 4452 3624 4468 3640
rect 4475 3638 4505 3690
rect 4539 3686 4540 3693
rect 4524 3678 4540 3686
rect 4511 3646 4524 3665
rect 4539 3646 4569 3662
rect 4511 3630 4585 3646
rect 4511 3628 4524 3630
rect 4539 3628 4573 3630
rect 4176 3606 4189 3608
rect 4204 3606 4238 3608
rect 4176 3590 4238 3606
rect 4282 3601 4298 3604
rect 4360 3601 4390 3612
rect 4438 3608 4484 3624
rect 4511 3612 4585 3628
rect 4438 3606 4472 3608
rect 4437 3590 4484 3606
rect 4511 3590 4524 3612
rect 4539 3590 4569 3612
rect 4596 3590 4597 3606
rect 4612 3590 4625 3750
rect -7 3582 34 3590
rect -7 3556 8 3582
rect 15 3556 34 3582
rect 98 3578 160 3590
rect 172 3578 247 3590
rect 305 3578 380 3590
rect 392 3578 423 3590
rect 429 3578 464 3590
rect 98 3576 260 3578
rect -7 3548 34 3556
rect 116 3552 129 3576
rect 144 3574 159 3576
rect -1 3538 0 3548
rect 15 3538 28 3548
rect 43 3538 73 3552
rect 116 3538 159 3552
rect 183 3549 190 3556
rect 193 3552 260 3576
rect 292 3576 464 3578
rect 262 3554 290 3558
rect 292 3554 372 3576
rect 393 3574 408 3576
rect 262 3552 372 3554
rect 193 3548 372 3552
rect 166 3538 196 3548
rect 198 3538 351 3548
rect 359 3538 389 3548
rect 393 3538 423 3552
rect 451 3538 464 3576
rect 536 3582 571 3590
rect 536 3556 537 3582
rect 544 3556 571 3582
rect 479 3538 509 3552
rect 536 3548 571 3556
rect 573 3582 614 3590
rect 573 3556 588 3582
rect 595 3556 614 3582
rect 678 3578 740 3590
rect 752 3578 827 3590
rect 885 3578 960 3590
rect 972 3578 1003 3590
rect 1009 3578 1044 3590
rect 678 3576 840 3578
rect 573 3548 614 3556
rect 696 3552 709 3576
rect 724 3574 739 3576
rect 536 3538 537 3548
rect 552 3538 565 3548
rect 579 3538 580 3548
rect 595 3538 608 3548
rect 623 3538 653 3552
rect 696 3538 739 3552
rect 763 3549 770 3556
rect 773 3552 840 3576
rect 872 3576 1044 3578
rect 842 3554 870 3558
rect 872 3554 952 3576
rect 973 3574 988 3576
rect 842 3552 952 3554
rect 773 3548 952 3552
rect 746 3538 776 3548
rect 778 3538 931 3548
rect 939 3538 969 3548
rect 973 3538 1003 3552
rect 1031 3538 1044 3576
rect 1116 3582 1151 3590
rect 1116 3556 1117 3582
rect 1124 3556 1151 3582
rect 1059 3538 1089 3552
rect 1116 3548 1151 3556
rect 1153 3582 1194 3590
rect 1153 3556 1168 3582
rect 1175 3556 1194 3582
rect 1258 3578 1320 3590
rect 1332 3578 1407 3590
rect 1465 3578 1540 3590
rect 1552 3578 1583 3590
rect 1589 3578 1624 3590
rect 1258 3576 1420 3578
rect 1153 3548 1194 3556
rect 1276 3552 1289 3576
rect 1304 3574 1319 3576
rect 1116 3538 1117 3548
rect 1132 3538 1145 3548
rect 1159 3538 1160 3548
rect 1175 3538 1188 3548
rect 1203 3538 1233 3552
rect 1276 3538 1319 3552
rect 1343 3549 1350 3556
rect 1353 3552 1420 3576
rect 1452 3576 1624 3578
rect 1422 3554 1450 3558
rect 1452 3554 1532 3576
rect 1553 3574 1568 3576
rect 1422 3552 1532 3554
rect 1353 3548 1532 3552
rect 1326 3538 1356 3548
rect 1358 3538 1511 3548
rect 1519 3538 1549 3548
rect 1553 3538 1583 3552
rect 1611 3538 1624 3576
rect 1696 3582 1731 3590
rect 1696 3556 1697 3582
rect 1704 3556 1731 3582
rect 1639 3538 1669 3552
rect 1696 3548 1731 3556
rect 1733 3582 1774 3590
rect 1733 3556 1748 3582
rect 1755 3556 1774 3582
rect 1838 3578 1900 3590
rect 1912 3578 1987 3590
rect 2045 3578 2120 3590
rect 2132 3578 2163 3590
rect 2169 3578 2204 3590
rect 1838 3576 2000 3578
rect 1733 3548 1774 3556
rect 1856 3552 1869 3576
rect 1884 3574 1899 3576
rect 1696 3538 1697 3548
rect 1712 3538 1725 3548
rect 1739 3538 1740 3548
rect 1755 3538 1768 3548
rect 1783 3538 1813 3552
rect 1856 3538 1899 3552
rect 1923 3549 1930 3556
rect 1933 3552 2000 3576
rect 2032 3576 2204 3578
rect 2002 3554 2030 3558
rect 2032 3554 2112 3576
rect 2133 3574 2148 3576
rect 2002 3552 2112 3554
rect 1933 3548 2112 3552
rect 1906 3538 1936 3548
rect 1938 3538 2091 3548
rect 2099 3538 2129 3548
rect 2133 3538 2163 3552
rect 2191 3538 2204 3576
rect 2276 3582 2311 3590
rect 2276 3556 2277 3582
rect 2284 3556 2311 3582
rect 2219 3538 2249 3552
rect 2276 3548 2311 3556
rect 2313 3582 2354 3590
rect 2313 3556 2328 3582
rect 2335 3556 2354 3582
rect 2418 3578 2480 3590
rect 2492 3578 2567 3590
rect 2625 3578 2700 3590
rect 2712 3578 2743 3590
rect 2749 3578 2784 3590
rect 2418 3576 2580 3578
rect 2313 3548 2354 3556
rect 2436 3552 2449 3576
rect 2464 3574 2479 3576
rect 2276 3538 2277 3548
rect 2292 3538 2305 3548
rect 2319 3538 2320 3548
rect 2335 3538 2348 3548
rect 2363 3538 2393 3552
rect 2436 3538 2479 3552
rect 2503 3549 2510 3556
rect 2513 3552 2580 3576
rect 2612 3576 2784 3578
rect 2582 3554 2610 3558
rect 2612 3554 2692 3576
rect 2713 3574 2728 3576
rect 2582 3552 2692 3554
rect 2513 3548 2692 3552
rect 2486 3538 2516 3548
rect 2518 3538 2671 3548
rect 2679 3538 2709 3548
rect 2713 3538 2743 3552
rect 2771 3538 2784 3576
rect 2856 3582 2891 3590
rect 2856 3556 2857 3582
rect 2864 3556 2891 3582
rect 2799 3538 2829 3552
rect 2856 3548 2891 3556
rect 2893 3582 2934 3590
rect 2893 3556 2908 3582
rect 2915 3556 2934 3582
rect 2998 3578 3060 3590
rect 3072 3578 3147 3590
rect 3205 3578 3280 3590
rect 3292 3578 3323 3590
rect 3329 3578 3364 3590
rect 2998 3576 3160 3578
rect 2893 3548 2934 3556
rect 3016 3552 3029 3576
rect 3044 3574 3059 3576
rect 2856 3538 2857 3548
rect 2872 3538 2885 3548
rect 2899 3538 2900 3548
rect 2915 3538 2928 3548
rect 2943 3538 2973 3552
rect 3016 3538 3059 3552
rect 3083 3549 3090 3556
rect 3093 3552 3160 3576
rect 3192 3576 3364 3578
rect 3162 3554 3190 3558
rect 3192 3554 3272 3576
rect 3293 3574 3308 3576
rect 3162 3552 3272 3554
rect 3093 3548 3272 3552
rect 3066 3538 3096 3548
rect 3098 3538 3251 3548
rect 3259 3538 3289 3548
rect 3293 3538 3323 3552
rect 3351 3538 3364 3576
rect 3436 3582 3471 3590
rect 3436 3556 3437 3582
rect 3444 3556 3471 3582
rect 3379 3538 3409 3552
rect 3436 3548 3471 3556
rect 3473 3582 3514 3590
rect 3473 3556 3488 3582
rect 3495 3556 3514 3582
rect 3578 3578 3640 3590
rect 3652 3578 3727 3590
rect 3785 3578 3860 3590
rect 3872 3578 3903 3590
rect 3909 3578 3944 3590
rect 3578 3576 3740 3578
rect 3473 3548 3514 3556
rect 3596 3552 3609 3576
rect 3624 3574 3639 3576
rect 3436 3538 3437 3548
rect 3452 3538 3465 3548
rect 3479 3538 3480 3548
rect 3495 3538 3508 3548
rect 3523 3538 3553 3552
rect 3596 3538 3639 3552
rect 3663 3549 3670 3556
rect 3673 3552 3740 3576
rect 3772 3576 3944 3578
rect 3742 3554 3770 3558
rect 3772 3554 3852 3576
rect 3873 3574 3888 3576
rect 3742 3552 3852 3554
rect 3673 3548 3852 3552
rect 3646 3538 3676 3548
rect 3678 3538 3831 3548
rect 3839 3538 3869 3548
rect 3873 3538 3903 3552
rect 3931 3538 3944 3576
rect 4016 3582 4051 3590
rect 4016 3556 4017 3582
rect 4024 3556 4051 3582
rect 3959 3538 3989 3552
rect 4016 3548 4051 3556
rect 4053 3582 4094 3590
rect 4053 3556 4068 3582
rect 4075 3556 4094 3582
rect 4158 3578 4220 3590
rect 4232 3578 4307 3590
rect 4365 3578 4440 3590
rect 4452 3578 4483 3590
rect 4489 3578 4524 3590
rect 4158 3576 4320 3578
rect 4053 3548 4094 3556
rect 4176 3552 4189 3576
rect 4204 3574 4219 3576
rect 4016 3538 4017 3548
rect 4032 3538 4045 3548
rect 4059 3538 4060 3548
rect 4075 3538 4088 3548
rect 4103 3538 4133 3552
rect 4176 3538 4219 3552
rect 4243 3549 4250 3556
rect 4253 3552 4320 3576
rect 4352 3576 4524 3578
rect 4322 3554 4350 3558
rect 4352 3554 4432 3576
rect 4453 3574 4468 3576
rect 4322 3552 4432 3554
rect 4253 3548 4432 3552
rect 4226 3538 4256 3548
rect 4258 3538 4411 3548
rect 4419 3538 4449 3548
rect 4453 3538 4483 3552
rect 4511 3538 4524 3576
rect 4596 3582 4631 3590
rect 4596 3556 4597 3582
rect 4604 3556 4631 3582
rect 4539 3538 4569 3552
rect 4596 3548 4631 3556
rect 4596 3538 4597 3548
rect 4612 3538 4625 3548
rect -1 3532 4625 3538
rect 0 3524 4625 3532
rect 15 3494 28 3524
rect 43 3506 73 3524
rect 116 3510 130 3524
rect 166 3510 386 3524
rect 117 3508 130 3510
rect 83 3496 98 3508
rect 80 3494 102 3496
rect 107 3494 137 3508
rect 198 3506 351 3510
rect 180 3494 372 3506
rect 415 3494 445 3508
rect 451 3494 464 3524
rect 479 3506 509 3524
rect 552 3494 565 3524
rect 595 3494 608 3524
rect 623 3506 653 3524
rect 696 3510 710 3524
rect 746 3510 966 3524
rect 697 3508 710 3510
rect 663 3496 678 3508
rect 660 3494 682 3496
rect 687 3494 717 3508
rect 778 3506 931 3510
rect 760 3494 952 3506
rect 995 3494 1025 3508
rect 1031 3494 1044 3524
rect 1059 3506 1089 3524
rect 1132 3494 1145 3524
rect 1175 3494 1188 3524
rect 1203 3506 1233 3524
rect 1276 3510 1290 3524
rect 1326 3510 1546 3524
rect 1277 3508 1290 3510
rect 1243 3496 1258 3508
rect 1240 3494 1262 3496
rect 1267 3494 1297 3508
rect 1358 3506 1511 3510
rect 1340 3494 1532 3506
rect 1575 3494 1605 3508
rect 1611 3494 1624 3524
rect 1639 3506 1669 3524
rect 1712 3494 1725 3524
rect 1755 3494 1768 3524
rect 1783 3506 1813 3524
rect 1856 3510 1870 3524
rect 1906 3510 2126 3524
rect 1857 3508 1870 3510
rect 1823 3496 1838 3508
rect 1820 3494 1842 3496
rect 1847 3494 1877 3508
rect 1938 3506 2091 3510
rect 1920 3494 2112 3506
rect 2155 3494 2185 3508
rect 2191 3494 2204 3524
rect 2219 3506 2249 3524
rect 2292 3494 2305 3524
rect 2335 3494 2348 3524
rect 2363 3506 2393 3524
rect 2436 3510 2450 3524
rect 2486 3510 2706 3524
rect 2437 3508 2450 3510
rect 2403 3496 2418 3508
rect 2400 3494 2422 3496
rect 2427 3494 2457 3508
rect 2518 3506 2671 3510
rect 2500 3494 2692 3506
rect 2735 3494 2765 3508
rect 2771 3494 2784 3524
rect 2799 3506 2829 3524
rect 2872 3494 2885 3524
rect 2915 3494 2928 3524
rect 2943 3506 2973 3524
rect 3016 3510 3030 3524
rect 3066 3510 3286 3524
rect 3017 3508 3030 3510
rect 2983 3496 2998 3508
rect 2980 3494 3002 3496
rect 3007 3494 3037 3508
rect 3098 3506 3251 3510
rect 3080 3494 3272 3506
rect 3315 3494 3345 3508
rect 3351 3494 3364 3524
rect 3379 3506 3409 3524
rect 3452 3494 3465 3524
rect 3495 3494 3508 3524
rect 3523 3506 3553 3524
rect 3596 3510 3610 3524
rect 3646 3510 3866 3524
rect 3597 3508 3610 3510
rect 3563 3496 3578 3508
rect 3560 3494 3582 3496
rect 3587 3494 3617 3508
rect 3678 3506 3831 3510
rect 3660 3494 3852 3506
rect 3895 3494 3925 3508
rect 3931 3494 3944 3524
rect 3959 3506 3989 3524
rect 4032 3494 4045 3524
rect 4075 3494 4088 3524
rect 4103 3506 4133 3524
rect 4176 3510 4190 3524
rect 4226 3510 4446 3524
rect 4177 3508 4190 3510
rect 4143 3496 4158 3508
rect 4140 3494 4162 3496
rect 4167 3494 4197 3508
rect 4258 3506 4411 3510
rect 4240 3494 4432 3506
rect 4475 3494 4505 3508
rect 4511 3494 4524 3524
rect 4539 3506 4569 3524
rect 4612 3494 4625 3524
rect 0 3480 4625 3494
rect 15 3376 28 3480
rect 73 3458 74 3468
rect 89 3458 102 3468
rect 73 3454 102 3458
rect 107 3454 137 3480
rect 155 3466 171 3468
rect 243 3466 296 3480
rect 244 3464 308 3466
rect 351 3464 366 3480
rect 415 3477 445 3480
rect 415 3474 451 3477
rect 381 3466 397 3468
rect 155 3454 170 3458
rect 73 3452 170 3454
rect 198 3452 366 3464
rect 382 3454 397 3458
rect 415 3455 454 3474
rect 473 3468 480 3469
rect 479 3461 480 3468
rect 463 3458 464 3461
rect 479 3458 492 3461
rect 415 3454 445 3455
rect 454 3454 460 3455
rect 463 3454 492 3458
rect 382 3453 492 3454
rect 382 3452 498 3453
rect 57 3444 108 3452
rect 57 3432 82 3444
rect 89 3432 108 3444
rect 139 3444 189 3452
rect 139 3436 155 3444
rect 162 3442 189 3444
rect 198 3442 419 3452
rect 162 3432 419 3442
rect 448 3444 498 3452
rect 448 3435 464 3444
rect 57 3424 108 3432
rect 155 3424 419 3432
rect 445 3432 464 3435
rect 471 3432 498 3444
rect 445 3424 498 3432
rect 73 3416 74 3424
rect 89 3416 102 3424
rect 73 3408 89 3416
rect 70 3401 89 3404
rect 70 3392 92 3401
rect 43 3382 92 3392
rect 43 3376 73 3382
rect 92 3377 97 3382
rect 15 3360 89 3376
rect 107 3368 137 3424
rect 172 3414 380 3424
rect 415 3420 460 3424
rect 463 3423 464 3424
rect 479 3423 492 3424
rect 198 3384 387 3414
rect 213 3381 387 3384
rect 206 3378 387 3381
rect 15 3358 28 3360
rect 43 3358 77 3360
rect 15 3342 89 3358
rect 116 3354 129 3368
rect 144 3354 160 3370
rect 206 3365 217 3378
rect -1 3320 0 3336
rect 15 3320 28 3342
rect 43 3320 73 3342
rect 116 3338 178 3354
rect 206 3347 217 3363
rect 222 3358 232 3378
rect 242 3358 256 3378
rect 259 3365 268 3378
rect 284 3365 293 3378
rect 222 3347 256 3358
rect 259 3347 268 3363
rect 284 3347 293 3363
rect 300 3358 310 3378
rect 320 3358 334 3378
rect 335 3365 346 3378
rect 300 3347 334 3358
rect 335 3347 346 3363
rect 392 3354 408 3370
rect 415 3368 445 3420
rect 479 3416 480 3423
rect 464 3408 480 3416
rect 451 3376 464 3395
rect 479 3376 509 3392
rect 451 3360 525 3376
rect 451 3358 464 3360
rect 479 3358 513 3360
rect 116 3336 129 3338
rect 144 3336 178 3338
rect 116 3320 178 3336
rect 222 3331 238 3334
rect 300 3331 330 3342
rect 378 3338 424 3354
rect 451 3342 525 3358
rect 378 3336 412 3338
rect 377 3320 424 3336
rect 451 3320 464 3342
rect 479 3320 509 3342
rect 536 3320 537 3336
rect 552 3320 565 3480
rect 595 3376 608 3480
rect 653 3458 654 3468
rect 669 3458 682 3468
rect 653 3454 682 3458
rect 687 3454 717 3480
rect 735 3466 751 3468
rect 823 3466 876 3480
rect 824 3464 888 3466
rect 931 3464 946 3480
rect 995 3477 1025 3480
rect 995 3474 1031 3477
rect 961 3466 977 3468
rect 735 3454 750 3458
rect 653 3452 750 3454
rect 778 3452 946 3464
rect 962 3454 977 3458
rect 995 3455 1034 3474
rect 1053 3468 1060 3469
rect 1059 3461 1060 3468
rect 1043 3458 1044 3461
rect 1059 3458 1072 3461
rect 995 3454 1025 3455
rect 1034 3454 1040 3455
rect 1043 3454 1072 3458
rect 962 3453 1072 3454
rect 962 3452 1078 3453
rect 637 3444 688 3452
rect 637 3432 662 3444
rect 669 3432 688 3444
rect 719 3444 769 3452
rect 719 3436 735 3444
rect 742 3442 769 3444
rect 778 3442 999 3452
rect 742 3432 999 3442
rect 1028 3444 1078 3452
rect 1028 3435 1044 3444
rect 637 3424 688 3432
rect 735 3424 999 3432
rect 1025 3432 1044 3435
rect 1051 3432 1078 3444
rect 1025 3424 1078 3432
rect 653 3416 654 3424
rect 669 3416 682 3424
rect 653 3408 669 3416
rect 650 3401 669 3404
rect 650 3392 672 3401
rect 623 3382 672 3392
rect 623 3376 653 3382
rect 672 3377 677 3382
rect 595 3360 669 3376
rect 687 3368 717 3424
rect 752 3414 960 3424
rect 995 3420 1040 3424
rect 1043 3423 1044 3424
rect 1059 3423 1072 3424
rect 778 3384 967 3414
rect 793 3381 967 3384
rect 786 3378 967 3381
rect 595 3358 608 3360
rect 623 3358 657 3360
rect 595 3342 669 3358
rect 696 3354 709 3368
rect 724 3354 740 3370
rect 786 3365 797 3378
rect 579 3320 580 3336
rect 595 3320 608 3342
rect 623 3320 653 3342
rect 696 3338 758 3354
rect 786 3347 797 3363
rect 802 3358 812 3378
rect 822 3358 836 3378
rect 839 3365 848 3378
rect 864 3365 873 3378
rect 802 3347 836 3358
rect 839 3347 848 3363
rect 864 3347 873 3363
rect 880 3358 890 3378
rect 900 3358 914 3378
rect 915 3365 926 3378
rect 880 3347 914 3358
rect 915 3347 926 3363
rect 972 3354 988 3370
rect 995 3368 1025 3420
rect 1059 3416 1060 3423
rect 1044 3408 1060 3416
rect 1031 3376 1044 3395
rect 1059 3376 1089 3392
rect 1031 3360 1105 3376
rect 1031 3358 1044 3360
rect 1059 3358 1093 3360
rect 696 3336 709 3338
rect 724 3336 758 3338
rect 696 3320 758 3336
rect 802 3331 818 3334
rect 880 3331 910 3342
rect 958 3338 1004 3354
rect 1031 3342 1105 3358
rect 958 3336 992 3338
rect 957 3320 1004 3336
rect 1031 3320 1044 3342
rect 1059 3320 1089 3342
rect 1116 3320 1117 3336
rect 1132 3320 1145 3480
rect 1175 3376 1188 3480
rect 1233 3458 1234 3468
rect 1249 3458 1262 3468
rect 1233 3454 1262 3458
rect 1267 3454 1297 3480
rect 1315 3466 1331 3468
rect 1403 3466 1456 3480
rect 1404 3464 1468 3466
rect 1511 3464 1526 3480
rect 1575 3477 1605 3480
rect 1575 3474 1611 3477
rect 1541 3466 1557 3468
rect 1315 3454 1330 3458
rect 1233 3452 1330 3454
rect 1358 3452 1526 3464
rect 1542 3454 1557 3458
rect 1575 3455 1614 3474
rect 1633 3468 1640 3469
rect 1639 3461 1640 3468
rect 1623 3458 1624 3461
rect 1639 3458 1652 3461
rect 1575 3454 1605 3455
rect 1614 3454 1620 3455
rect 1623 3454 1652 3458
rect 1542 3453 1652 3454
rect 1542 3452 1658 3453
rect 1217 3444 1268 3452
rect 1217 3432 1242 3444
rect 1249 3432 1268 3444
rect 1299 3444 1349 3452
rect 1299 3436 1315 3444
rect 1322 3442 1349 3444
rect 1358 3442 1579 3452
rect 1322 3432 1579 3442
rect 1608 3444 1658 3452
rect 1608 3435 1624 3444
rect 1217 3424 1268 3432
rect 1315 3424 1579 3432
rect 1605 3432 1624 3435
rect 1631 3432 1658 3444
rect 1605 3424 1658 3432
rect 1233 3416 1234 3424
rect 1249 3416 1262 3424
rect 1233 3408 1249 3416
rect 1230 3401 1249 3404
rect 1230 3392 1252 3401
rect 1203 3382 1252 3392
rect 1203 3376 1233 3382
rect 1252 3377 1257 3382
rect 1175 3360 1249 3376
rect 1267 3368 1297 3424
rect 1332 3414 1540 3424
rect 1575 3420 1620 3424
rect 1623 3423 1624 3424
rect 1639 3423 1652 3424
rect 1358 3384 1547 3414
rect 1373 3381 1547 3384
rect 1366 3378 1547 3381
rect 1175 3358 1188 3360
rect 1203 3358 1237 3360
rect 1175 3342 1249 3358
rect 1276 3354 1289 3368
rect 1304 3354 1320 3370
rect 1366 3365 1377 3378
rect 1159 3320 1160 3336
rect 1175 3320 1188 3342
rect 1203 3320 1233 3342
rect 1276 3338 1338 3354
rect 1366 3347 1377 3363
rect 1382 3358 1392 3378
rect 1402 3358 1416 3378
rect 1419 3365 1428 3378
rect 1444 3365 1453 3378
rect 1382 3347 1416 3358
rect 1419 3347 1428 3363
rect 1444 3347 1453 3363
rect 1460 3358 1470 3378
rect 1480 3358 1494 3378
rect 1495 3365 1506 3378
rect 1460 3347 1494 3358
rect 1495 3347 1506 3363
rect 1552 3354 1568 3370
rect 1575 3368 1605 3420
rect 1639 3416 1640 3423
rect 1624 3408 1640 3416
rect 1611 3376 1624 3395
rect 1639 3376 1669 3392
rect 1611 3360 1685 3376
rect 1611 3358 1624 3360
rect 1639 3358 1673 3360
rect 1276 3336 1289 3338
rect 1304 3336 1338 3338
rect 1276 3320 1338 3336
rect 1382 3331 1398 3334
rect 1460 3331 1490 3342
rect 1538 3338 1584 3354
rect 1611 3342 1685 3358
rect 1538 3336 1572 3338
rect 1537 3320 1584 3336
rect 1611 3320 1624 3342
rect 1639 3320 1669 3342
rect 1696 3320 1697 3336
rect 1712 3320 1725 3480
rect 1755 3376 1768 3480
rect 1813 3458 1814 3468
rect 1829 3458 1842 3468
rect 1813 3454 1842 3458
rect 1847 3454 1877 3480
rect 1895 3466 1911 3468
rect 1983 3466 2036 3480
rect 1984 3464 2048 3466
rect 2091 3464 2106 3480
rect 2155 3477 2185 3480
rect 2155 3474 2191 3477
rect 2121 3466 2137 3468
rect 1895 3454 1910 3458
rect 1813 3452 1910 3454
rect 1938 3452 2106 3464
rect 2122 3454 2137 3458
rect 2155 3455 2194 3474
rect 2213 3468 2220 3469
rect 2219 3461 2220 3468
rect 2203 3458 2204 3461
rect 2219 3458 2232 3461
rect 2155 3454 2185 3455
rect 2194 3454 2200 3455
rect 2203 3454 2232 3458
rect 2122 3453 2232 3454
rect 2122 3452 2238 3453
rect 1797 3444 1848 3452
rect 1797 3432 1822 3444
rect 1829 3432 1848 3444
rect 1879 3444 1929 3452
rect 1879 3436 1895 3444
rect 1902 3442 1929 3444
rect 1938 3442 2159 3452
rect 1902 3432 2159 3442
rect 2188 3444 2238 3452
rect 2188 3435 2204 3444
rect 1797 3424 1848 3432
rect 1895 3424 2159 3432
rect 2185 3432 2204 3435
rect 2211 3432 2238 3444
rect 2185 3424 2238 3432
rect 1813 3416 1814 3424
rect 1829 3416 1842 3424
rect 1813 3408 1829 3416
rect 1810 3401 1829 3404
rect 1810 3392 1832 3401
rect 1783 3382 1832 3392
rect 1783 3376 1813 3382
rect 1832 3377 1837 3382
rect 1755 3360 1829 3376
rect 1847 3368 1877 3424
rect 1912 3414 2120 3424
rect 2155 3420 2200 3424
rect 2203 3423 2204 3424
rect 2219 3423 2232 3424
rect 1938 3384 2127 3414
rect 1953 3381 2127 3384
rect 1946 3378 2127 3381
rect 1755 3358 1768 3360
rect 1783 3358 1817 3360
rect 1755 3342 1829 3358
rect 1856 3354 1869 3368
rect 1884 3354 1900 3370
rect 1946 3365 1957 3378
rect 1739 3320 1740 3336
rect 1755 3320 1768 3342
rect 1783 3320 1813 3342
rect 1856 3338 1918 3354
rect 1946 3347 1957 3363
rect 1962 3358 1972 3378
rect 1982 3358 1996 3378
rect 1999 3365 2008 3378
rect 2024 3365 2033 3378
rect 1962 3347 1996 3358
rect 1999 3347 2008 3363
rect 2024 3347 2033 3363
rect 2040 3358 2050 3378
rect 2060 3358 2074 3378
rect 2075 3365 2086 3378
rect 2040 3347 2074 3358
rect 2075 3347 2086 3363
rect 2132 3354 2148 3370
rect 2155 3368 2185 3420
rect 2219 3416 2220 3423
rect 2204 3408 2220 3416
rect 2191 3376 2204 3395
rect 2219 3376 2249 3392
rect 2191 3360 2265 3376
rect 2191 3358 2204 3360
rect 2219 3358 2253 3360
rect 1856 3336 1869 3338
rect 1884 3336 1918 3338
rect 1856 3320 1918 3336
rect 1962 3331 1978 3334
rect 2040 3331 2070 3342
rect 2118 3338 2164 3354
rect 2191 3342 2265 3358
rect 2118 3336 2152 3338
rect 2117 3320 2164 3336
rect 2191 3320 2204 3342
rect 2219 3320 2249 3342
rect 2276 3320 2277 3336
rect 2292 3320 2305 3480
rect 2335 3376 2348 3480
rect 2393 3458 2394 3468
rect 2409 3458 2422 3468
rect 2393 3454 2422 3458
rect 2427 3454 2457 3480
rect 2475 3466 2491 3468
rect 2563 3466 2616 3480
rect 2564 3464 2628 3466
rect 2671 3464 2686 3480
rect 2735 3477 2765 3480
rect 2735 3474 2771 3477
rect 2701 3466 2717 3468
rect 2475 3454 2490 3458
rect 2393 3452 2490 3454
rect 2518 3452 2686 3464
rect 2702 3454 2717 3458
rect 2735 3455 2774 3474
rect 2793 3468 2800 3469
rect 2799 3461 2800 3468
rect 2783 3458 2784 3461
rect 2799 3458 2812 3461
rect 2735 3454 2765 3455
rect 2774 3454 2780 3455
rect 2783 3454 2812 3458
rect 2702 3453 2812 3454
rect 2702 3452 2818 3453
rect 2377 3444 2428 3452
rect 2377 3432 2402 3444
rect 2409 3432 2428 3444
rect 2459 3444 2509 3452
rect 2459 3436 2475 3444
rect 2482 3442 2509 3444
rect 2518 3442 2739 3452
rect 2482 3432 2739 3442
rect 2768 3444 2818 3452
rect 2768 3435 2784 3444
rect 2377 3424 2428 3432
rect 2475 3424 2739 3432
rect 2765 3432 2784 3435
rect 2791 3432 2818 3444
rect 2765 3424 2818 3432
rect 2393 3416 2394 3424
rect 2409 3416 2422 3424
rect 2393 3408 2409 3416
rect 2390 3401 2409 3404
rect 2390 3392 2412 3401
rect 2363 3382 2412 3392
rect 2363 3376 2393 3382
rect 2412 3377 2417 3382
rect 2335 3360 2409 3376
rect 2427 3368 2457 3424
rect 2492 3414 2700 3424
rect 2735 3420 2780 3424
rect 2783 3423 2784 3424
rect 2799 3423 2812 3424
rect 2518 3384 2707 3414
rect 2533 3381 2707 3384
rect 2526 3378 2707 3381
rect 2335 3358 2348 3360
rect 2363 3358 2397 3360
rect 2335 3342 2409 3358
rect 2436 3354 2449 3368
rect 2464 3354 2480 3370
rect 2526 3365 2537 3378
rect 2319 3320 2320 3336
rect 2335 3320 2348 3342
rect 2363 3320 2393 3342
rect 2436 3338 2498 3354
rect 2526 3347 2537 3363
rect 2542 3358 2552 3378
rect 2562 3358 2576 3378
rect 2579 3365 2588 3378
rect 2604 3365 2613 3378
rect 2542 3347 2576 3358
rect 2579 3347 2588 3363
rect 2604 3347 2613 3363
rect 2620 3358 2630 3378
rect 2640 3358 2654 3378
rect 2655 3365 2666 3378
rect 2620 3347 2654 3358
rect 2655 3347 2666 3363
rect 2712 3354 2728 3370
rect 2735 3368 2765 3420
rect 2799 3416 2800 3423
rect 2784 3408 2800 3416
rect 2771 3376 2784 3395
rect 2799 3376 2829 3392
rect 2771 3360 2845 3376
rect 2771 3358 2784 3360
rect 2799 3358 2833 3360
rect 2436 3336 2449 3338
rect 2464 3336 2498 3338
rect 2436 3320 2498 3336
rect 2542 3331 2558 3334
rect 2620 3331 2650 3342
rect 2698 3338 2744 3354
rect 2771 3342 2845 3358
rect 2698 3336 2732 3338
rect 2697 3320 2744 3336
rect 2771 3320 2784 3342
rect 2799 3320 2829 3342
rect 2856 3320 2857 3336
rect 2872 3320 2885 3480
rect 2915 3376 2928 3480
rect 2973 3458 2974 3468
rect 2989 3458 3002 3468
rect 2973 3454 3002 3458
rect 3007 3454 3037 3480
rect 3055 3466 3071 3468
rect 3143 3466 3196 3480
rect 3144 3464 3208 3466
rect 3251 3464 3266 3480
rect 3315 3477 3345 3480
rect 3315 3474 3351 3477
rect 3281 3466 3297 3468
rect 3055 3454 3070 3458
rect 2973 3452 3070 3454
rect 3098 3452 3266 3464
rect 3282 3454 3297 3458
rect 3315 3455 3354 3474
rect 3373 3468 3380 3469
rect 3379 3461 3380 3468
rect 3363 3458 3364 3461
rect 3379 3458 3392 3461
rect 3315 3454 3345 3455
rect 3354 3454 3360 3455
rect 3363 3454 3392 3458
rect 3282 3453 3392 3454
rect 3282 3452 3398 3453
rect 2957 3444 3008 3452
rect 2957 3432 2982 3444
rect 2989 3432 3008 3444
rect 3039 3444 3089 3452
rect 3039 3436 3055 3444
rect 3062 3442 3089 3444
rect 3098 3442 3319 3452
rect 3062 3432 3319 3442
rect 3348 3444 3398 3452
rect 3348 3435 3364 3444
rect 2957 3424 3008 3432
rect 3055 3424 3319 3432
rect 3345 3432 3364 3435
rect 3371 3432 3398 3444
rect 3345 3424 3398 3432
rect 2973 3416 2974 3424
rect 2989 3416 3002 3424
rect 2973 3408 2989 3416
rect 2970 3401 2989 3404
rect 2970 3392 2992 3401
rect 2943 3382 2992 3392
rect 2943 3376 2973 3382
rect 2992 3377 2997 3382
rect 2915 3360 2989 3376
rect 3007 3368 3037 3424
rect 3072 3414 3280 3424
rect 3315 3420 3360 3424
rect 3363 3423 3364 3424
rect 3379 3423 3392 3424
rect 3098 3384 3287 3414
rect 3113 3381 3287 3384
rect 3106 3378 3287 3381
rect 2915 3358 2928 3360
rect 2943 3358 2977 3360
rect 2915 3342 2989 3358
rect 3016 3354 3029 3368
rect 3044 3354 3060 3370
rect 3106 3365 3117 3378
rect 2899 3320 2900 3336
rect 2915 3320 2928 3342
rect 2943 3320 2973 3342
rect 3016 3338 3078 3354
rect 3106 3347 3117 3363
rect 3122 3358 3132 3378
rect 3142 3358 3156 3378
rect 3159 3365 3168 3378
rect 3184 3365 3193 3378
rect 3122 3347 3156 3358
rect 3159 3347 3168 3363
rect 3184 3347 3193 3363
rect 3200 3358 3210 3378
rect 3220 3358 3234 3378
rect 3235 3365 3246 3378
rect 3200 3347 3234 3358
rect 3235 3347 3246 3363
rect 3292 3354 3308 3370
rect 3315 3368 3345 3420
rect 3379 3416 3380 3423
rect 3364 3408 3380 3416
rect 3351 3376 3364 3395
rect 3379 3376 3409 3392
rect 3351 3360 3425 3376
rect 3351 3358 3364 3360
rect 3379 3358 3413 3360
rect 3016 3336 3029 3338
rect 3044 3336 3078 3338
rect 3016 3320 3078 3336
rect 3122 3331 3138 3334
rect 3200 3331 3230 3342
rect 3278 3338 3324 3354
rect 3351 3342 3425 3358
rect 3278 3336 3312 3338
rect 3277 3320 3324 3336
rect 3351 3320 3364 3342
rect 3379 3320 3409 3342
rect 3436 3320 3437 3336
rect 3452 3320 3465 3480
rect 3495 3376 3508 3480
rect 3553 3458 3554 3468
rect 3569 3458 3582 3468
rect 3553 3454 3582 3458
rect 3587 3454 3617 3480
rect 3635 3466 3651 3468
rect 3723 3466 3776 3480
rect 3724 3464 3788 3466
rect 3831 3464 3846 3480
rect 3895 3477 3925 3480
rect 3895 3474 3931 3477
rect 3861 3466 3877 3468
rect 3635 3454 3650 3458
rect 3553 3452 3650 3454
rect 3678 3452 3846 3464
rect 3862 3454 3877 3458
rect 3895 3455 3934 3474
rect 3953 3468 3960 3469
rect 3959 3461 3960 3468
rect 3943 3458 3944 3461
rect 3959 3458 3972 3461
rect 3895 3454 3925 3455
rect 3934 3454 3940 3455
rect 3943 3454 3972 3458
rect 3862 3453 3972 3454
rect 3862 3452 3978 3453
rect 3537 3444 3588 3452
rect 3537 3432 3562 3444
rect 3569 3432 3588 3444
rect 3619 3444 3669 3452
rect 3619 3436 3635 3444
rect 3642 3442 3669 3444
rect 3678 3442 3899 3452
rect 3642 3432 3899 3442
rect 3928 3444 3978 3452
rect 3928 3435 3944 3444
rect 3537 3424 3588 3432
rect 3635 3424 3899 3432
rect 3925 3432 3944 3435
rect 3951 3432 3978 3444
rect 3925 3424 3978 3432
rect 3553 3416 3554 3424
rect 3569 3416 3582 3424
rect 3553 3408 3569 3416
rect 3550 3401 3569 3404
rect 3550 3392 3572 3401
rect 3523 3382 3572 3392
rect 3523 3376 3553 3382
rect 3572 3377 3577 3382
rect 3495 3360 3569 3376
rect 3587 3368 3617 3424
rect 3652 3414 3860 3424
rect 3895 3420 3940 3424
rect 3943 3423 3944 3424
rect 3959 3423 3972 3424
rect 3678 3384 3867 3414
rect 3693 3381 3867 3384
rect 3686 3378 3867 3381
rect 3495 3358 3508 3360
rect 3523 3358 3557 3360
rect 3495 3342 3569 3358
rect 3596 3354 3609 3368
rect 3624 3354 3640 3370
rect 3686 3365 3697 3378
rect 3479 3320 3480 3336
rect 3495 3320 3508 3342
rect 3523 3320 3553 3342
rect 3596 3338 3658 3354
rect 3686 3347 3697 3363
rect 3702 3358 3712 3378
rect 3722 3358 3736 3378
rect 3739 3365 3748 3378
rect 3764 3365 3773 3378
rect 3702 3347 3736 3358
rect 3739 3347 3748 3363
rect 3764 3347 3773 3363
rect 3780 3358 3790 3378
rect 3800 3358 3814 3378
rect 3815 3365 3826 3378
rect 3780 3347 3814 3358
rect 3815 3347 3826 3363
rect 3872 3354 3888 3370
rect 3895 3368 3925 3420
rect 3959 3416 3960 3423
rect 3944 3408 3960 3416
rect 3931 3376 3944 3395
rect 3959 3376 3989 3392
rect 3931 3360 4005 3376
rect 3931 3358 3944 3360
rect 3959 3358 3993 3360
rect 3596 3336 3609 3338
rect 3624 3336 3658 3338
rect 3596 3320 3658 3336
rect 3702 3331 3718 3334
rect 3780 3331 3810 3342
rect 3858 3338 3904 3354
rect 3931 3342 4005 3358
rect 3858 3336 3892 3338
rect 3857 3320 3904 3336
rect 3931 3320 3944 3342
rect 3959 3320 3989 3342
rect 4016 3320 4017 3336
rect 4032 3320 4045 3480
rect 4075 3376 4088 3480
rect 4133 3458 4134 3468
rect 4149 3458 4162 3468
rect 4133 3454 4162 3458
rect 4167 3454 4197 3480
rect 4215 3466 4231 3468
rect 4303 3466 4356 3480
rect 4304 3464 4368 3466
rect 4411 3464 4426 3480
rect 4475 3477 4505 3480
rect 4475 3474 4511 3477
rect 4441 3466 4457 3468
rect 4215 3454 4230 3458
rect 4133 3452 4230 3454
rect 4258 3452 4426 3464
rect 4442 3454 4457 3458
rect 4475 3455 4514 3474
rect 4533 3468 4540 3469
rect 4539 3461 4540 3468
rect 4523 3458 4524 3461
rect 4539 3458 4552 3461
rect 4475 3454 4505 3455
rect 4514 3454 4520 3455
rect 4523 3454 4552 3458
rect 4442 3453 4552 3454
rect 4442 3452 4558 3453
rect 4117 3444 4168 3452
rect 4117 3432 4142 3444
rect 4149 3432 4168 3444
rect 4199 3444 4249 3452
rect 4199 3436 4215 3444
rect 4222 3442 4249 3444
rect 4258 3442 4479 3452
rect 4222 3432 4479 3442
rect 4508 3444 4558 3452
rect 4508 3435 4524 3444
rect 4117 3424 4168 3432
rect 4215 3424 4479 3432
rect 4505 3432 4524 3435
rect 4531 3432 4558 3444
rect 4505 3424 4558 3432
rect 4133 3416 4134 3424
rect 4149 3416 4162 3424
rect 4133 3408 4149 3416
rect 4130 3401 4149 3404
rect 4130 3392 4152 3401
rect 4103 3382 4152 3392
rect 4103 3376 4133 3382
rect 4152 3377 4157 3382
rect 4075 3360 4149 3376
rect 4167 3368 4197 3424
rect 4232 3414 4440 3424
rect 4475 3420 4520 3424
rect 4523 3423 4524 3424
rect 4539 3423 4552 3424
rect 4258 3384 4447 3414
rect 4273 3381 4447 3384
rect 4266 3378 4447 3381
rect 4075 3358 4088 3360
rect 4103 3358 4137 3360
rect 4075 3342 4149 3358
rect 4176 3354 4189 3368
rect 4204 3354 4220 3370
rect 4266 3365 4277 3378
rect 4059 3320 4060 3336
rect 4075 3320 4088 3342
rect 4103 3320 4133 3342
rect 4176 3338 4238 3354
rect 4266 3347 4277 3363
rect 4282 3358 4292 3378
rect 4302 3358 4316 3378
rect 4319 3365 4328 3378
rect 4344 3365 4353 3378
rect 4282 3347 4316 3358
rect 4319 3347 4328 3363
rect 4344 3347 4353 3363
rect 4360 3358 4370 3378
rect 4380 3358 4394 3378
rect 4395 3365 4406 3378
rect 4360 3347 4394 3358
rect 4395 3347 4406 3363
rect 4452 3354 4468 3370
rect 4475 3368 4505 3420
rect 4539 3416 4540 3423
rect 4524 3408 4540 3416
rect 4511 3376 4524 3395
rect 4539 3376 4569 3392
rect 4511 3360 4585 3376
rect 4511 3358 4524 3360
rect 4539 3358 4573 3360
rect 4176 3336 4189 3338
rect 4204 3336 4238 3338
rect 4176 3320 4238 3336
rect 4282 3331 4298 3334
rect 4360 3331 4390 3342
rect 4438 3338 4484 3354
rect 4511 3342 4585 3358
rect 4438 3336 4472 3338
rect 4437 3320 4484 3336
rect 4511 3320 4524 3342
rect 4539 3320 4569 3342
rect 4596 3320 4597 3336
rect 4612 3320 4625 3480
rect -7 3312 34 3320
rect -7 3286 8 3312
rect 15 3286 34 3312
rect 98 3308 160 3320
rect 172 3308 247 3320
rect 305 3308 380 3320
rect 392 3308 423 3320
rect 429 3308 464 3320
rect 98 3306 260 3308
rect -7 3278 34 3286
rect 116 3282 129 3306
rect 144 3304 159 3306
rect -1 3268 0 3278
rect 15 3268 28 3278
rect 43 3268 73 3282
rect 116 3268 159 3282
rect 183 3279 190 3286
rect 193 3282 260 3306
rect 292 3306 464 3308
rect 262 3284 290 3288
rect 292 3284 372 3306
rect 393 3304 408 3306
rect 262 3282 372 3284
rect 193 3278 372 3282
rect 166 3268 196 3278
rect 198 3268 351 3278
rect 359 3268 389 3278
rect 393 3268 423 3282
rect 451 3268 464 3306
rect 536 3312 571 3320
rect 536 3286 537 3312
rect 544 3286 571 3312
rect 479 3268 509 3282
rect 536 3278 571 3286
rect 573 3312 614 3320
rect 573 3286 588 3312
rect 595 3286 614 3312
rect 678 3308 740 3320
rect 752 3308 827 3320
rect 885 3308 960 3320
rect 972 3308 1003 3320
rect 1009 3308 1044 3320
rect 678 3306 840 3308
rect 573 3278 614 3286
rect 696 3282 709 3306
rect 724 3304 739 3306
rect 536 3268 537 3278
rect 552 3268 565 3278
rect 579 3268 580 3278
rect 595 3268 608 3278
rect 623 3268 653 3282
rect 696 3268 739 3282
rect 763 3279 770 3286
rect 773 3282 840 3306
rect 872 3306 1044 3308
rect 842 3284 870 3288
rect 872 3284 952 3306
rect 973 3304 988 3306
rect 842 3282 952 3284
rect 773 3278 952 3282
rect 746 3268 776 3278
rect 778 3268 931 3278
rect 939 3268 969 3278
rect 973 3268 1003 3282
rect 1031 3268 1044 3306
rect 1116 3312 1151 3320
rect 1116 3286 1117 3312
rect 1124 3286 1151 3312
rect 1059 3268 1089 3282
rect 1116 3278 1151 3286
rect 1153 3312 1194 3320
rect 1153 3286 1168 3312
rect 1175 3286 1194 3312
rect 1258 3308 1320 3320
rect 1332 3308 1407 3320
rect 1465 3308 1540 3320
rect 1552 3308 1583 3320
rect 1589 3308 1624 3320
rect 1258 3306 1420 3308
rect 1153 3278 1194 3286
rect 1276 3282 1289 3306
rect 1304 3304 1319 3306
rect 1116 3268 1117 3278
rect 1132 3268 1145 3278
rect 1159 3268 1160 3278
rect 1175 3268 1188 3278
rect 1203 3268 1233 3282
rect 1276 3268 1319 3282
rect 1343 3279 1350 3286
rect 1353 3282 1420 3306
rect 1452 3306 1624 3308
rect 1422 3284 1450 3288
rect 1452 3284 1532 3306
rect 1553 3304 1568 3306
rect 1422 3282 1532 3284
rect 1353 3278 1532 3282
rect 1326 3268 1356 3278
rect 1358 3268 1511 3278
rect 1519 3268 1549 3278
rect 1553 3268 1583 3282
rect 1611 3268 1624 3306
rect 1696 3312 1731 3320
rect 1696 3286 1697 3312
rect 1704 3286 1731 3312
rect 1639 3268 1669 3282
rect 1696 3278 1731 3286
rect 1733 3312 1774 3320
rect 1733 3286 1748 3312
rect 1755 3286 1774 3312
rect 1838 3308 1900 3320
rect 1912 3308 1987 3320
rect 2045 3308 2120 3320
rect 2132 3308 2163 3320
rect 2169 3308 2204 3320
rect 1838 3306 2000 3308
rect 1733 3278 1774 3286
rect 1856 3282 1869 3306
rect 1884 3304 1899 3306
rect 1696 3268 1697 3278
rect 1712 3268 1725 3278
rect 1739 3268 1740 3278
rect 1755 3268 1768 3278
rect 1783 3268 1813 3282
rect 1856 3268 1899 3282
rect 1923 3279 1930 3286
rect 1933 3282 2000 3306
rect 2032 3306 2204 3308
rect 2002 3284 2030 3288
rect 2032 3284 2112 3306
rect 2133 3304 2148 3306
rect 2002 3282 2112 3284
rect 1933 3278 2112 3282
rect 1906 3268 1936 3278
rect 1938 3268 2091 3278
rect 2099 3268 2129 3278
rect 2133 3268 2163 3282
rect 2191 3268 2204 3306
rect 2276 3312 2311 3320
rect 2276 3286 2277 3312
rect 2284 3286 2311 3312
rect 2219 3268 2249 3282
rect 2276 3278 2311 3286
rect 2313 3312 2354 3320
rect 2313 3286 2328 3312
rect 2335 3286 2354 3312
rect 2418 3308 2480 3320
rect 2492 3308 2567 3320
rect 2625 3308 2700 3320
rect 2712 3308 2743 3320
rect 2749 3308 2784 3320
rect 2418 3306 2580 3308
rect 2313 3278 2354 3286
rect 2436 3282 2449 3306
rect 2464 3304 2479 3306
rect 2276 3268 2277 3278
rect 2292 3268 2305 3278
rect 2319 3268 2320 3278
rect 2335 3268 2348 3278
rect 2363 3268 2393 3282
rect 2436 3268 2479 3282
rect 2503 3279 2510 3286
rect 2513 3282 2580 3306
rect 2612 3306 2784 3308
rect 2582 3284 2610 3288
rect 2612 3284 2692 3306
rect 2713 3304 2728 3306
rect 2582 3282 2692 3284
rect 2513 3278 2692 3282
rect 2486 3268 2516 3278
rect 2518 3268 2671 3278
rect 2679 3268 2709 3278
rect 2713 3268 2743 3282
rect 2771 3268 2784 3306
rect 2856 3312 2891 3320
rect 2856 3286 2857 3312
rect 2864 3286 2891 3312
rect 2799 3268 2829 3282
rect 2856 3278 2891 3286
rect 2893 3312 2934 3320
rect 2893 3286 2908 3312
rect 2915 3286 2934 3312
rect 2998 3308 3060 3320
rect 3072 3308 3147 3320
rect 3205 3308 3280 3320
rect 3292 3308 3323 3320
rect 3329 3308 3364 3320
rect 2998 3306 3160 3308
rect 2893 3278 2934 3286
rect 3016 3282 3029 3306
rect 3044 3304 3059 3306
rect 2856 3268 2857 3278
rect 2872 3268 2885 3278
rect 2899 3268 2900 3278
rect 2915 3268 2928 3278
rect 2943 3268 2973 3282
rect 3016 3268 3059 3282
rect 3083 3279 3090 3286
rect 3093 3282 3160 3306
rect 3192 3306 3364 3308
rect 3162 3284 3190 3288
rect 3192 3284 3272 3306
rect 3293 3304 3308 3306
rect 3162 3282 3272 3284
rect 3093 3278 3272 3282
rect 3066 3268 3096 3278
rect 3098 3268 3251 3278
rect 3259 3268 3289 3278
rect 3293 3268 3323 3282
rect 3351 3268 3364 3306
rect 3436 3312 3471 3320
rect 3436 3286 3437 3312
rect 3444 3286 3471 3312
rect 3379 3268 3409 3282
rect 3436 3278 3471 3286
rect 3473 3312 3514 3320
rect 3473 3286 3488 3312
rect 3495 3286 3514 3312
rect 3578 3308 3640 3320
rect 3652 3308 3727 3320
rect 3785 3308 3860 3320
rect 3872 3308 3903 3320
rect 3909 3308 3944 3320
rect 3578 3306 3740 3308
rect 3473 3278 3514 3286
rect 3596 3282 3609 3306
rect 3624 3304 3639 3306
rect 3436 3268 3437 3278
rect 3452 3268 3465 3278
rect 3479 3268 3480 3278
rect 3495 3268 3508 3278
rect 3523 3268 3553 3282
rect 3596 3268 3639 3282
rect 3663 3279 3670 3286
rect 3673 3282 3740 3306
rect 3772 3306 3944 3308
rect 3742 3284 3770 3288
rect 3772 3284 3852 3306
rect 3873 3304 3888 3306
rect 3742 3282 3852 3284
rect 3673 3278 3852 3282
rect 3646 3268 3676 3278
rect 3678 3268 3831 3278
rect 3839 3268 3869 3278
rect 3873 3268 3903 3282
rect 3931 3268 3944 3306
rect 4016 3312 4051 3320
rect 4016 3286 4017 3312
rect 4024 3286 4051 3312
rect 3959 3268 3989 3282
rect 4016 3278 4051 3286
rect 4053 3312 4094 3320
rect 4053 3286 4068 3312
rect 4075 3286 4094 3312
rect 4158 3308 4220 3320
rect 4232 3308 4307 3320
rect 4365 3308 4440 3320
rect 4452 3308 4483 3320
rect 4489 3308 4524 3320
rect 4158 3306 4320 3308
rect 4053 3278 4094 3286
rect 4176 3282 4189 3306
rect 4204 3304 4219 3306
rect 4016 3268 4017 3278
rect 4032 3268 4045 3278
rect 4059 3268 4060 3278
rect 4075 3268 4088 3278
rect 4103 3268 4133 3282
rect 4176 3268 4219 3282
rect 4243 3279 4250 3286
rect 4253 3282 4320 3306
rect 4352 3306 4524 3308
rect 4322 3284 4350 3288
rect 4352 3284 4432 3306
rect 4453 3304 4468 3306
rect 4322 3282 4432 3284
rect 4253 3278 4432 3282
rect 4226 3268 4256 3278
rect 4258 3268 4411 3278
rect 4419 3268 4449 3278
rect 4453 3268 4483 3282
rect 4511 3268 4524 3306
rect 4596 3312 4631 3320
rect 4596 3286 4597 3312
rect 4604 3286 4631 3312
rect 4539 3268 4569 3282
rect 4596 3278 4631 3286
rect 4596 3268 4597 3278
rect 4612 3268 4625 3278
rect -1 3262 4625 3268
rect 0 3254 4625 3262
rect 15 3224 28 3254
rect 43 3236 73 3254
rect 116 3240 130 3254
rect 166 3240 386 3254
rect 117 3238 130 3240
rect 83 3226 98 3238
rect 80 3224 102 3226
rect 107 3224 137 3238
rect 198 3236 351 3240
rect 180 3224 372 3236
rect 415 3224 445 3238
rect 451 3224 464 3254
rect 479 3236 509 3254
rect 552 3224 565 3254
rect 595 3224 608 3254
rect 623 3236 653 3254
rect 696 3240 710 3254
rect 746 3240 966 3254
rect 697 3238 710 3240
rect 663 3226 678 3238
rect 660 3224 682 3226
rect 687 3224 717 3238
rect 778 3236 931 3240
rect 760 3224 952 3236
rect 995 3224 1025 3238
rect 1031 3224 1044 3254
rect 1059 3236 1089 3254
rect 1132 3224 1145 3254
rect 1175 3224 1188 3254
rect 1203 3236 1233 3254
rect 1276 3240 1290 3254
rect 1326 3240 1546 3254
rect 1277 3238 1290 3240
rect 1243 3226 1258 3238
rect 1240 3224 1262 3226
rect 1267 3224 1297 3238
rect 1358 3236 1511 3240
rect 1340 3224 1532 3236
rect 1575 3224 1605 3238
rect 1611 3224 1624 3254
rect 1639 3236 1669 3254
rect 1712 3224 1725 3254
rect 1755 3224 1768 3254
rect 1783 3236 1813 3254
rect 1856 3240 1870 3254
rect 1906 3240 2126 3254
rect 1857 3238 1870 3240
rect 1823 3226 1838 3238
rect 1820 3224 1842 3226
rect 1847 3224 1877 3238
rect 1938 3236 2091 3240
rect 1920 3224 2112 3236
rect 2155 3224 2185 3238
rect 2191 3224 2204 3254
rect 2219 3236 2249 3254
rect 2292 3224 2305 3254
rect 2335 3224 2348 3254
rect 2363 3236 2393 3254
rect 2436 3240 2450 3254
rect 2486 3240 2706 3254
rect 2437 3238 2450 3240
rect 2403 3226 2418 3238
rect 2400 3224 2422 3226
rect 2427 3224 2457 3238
rect 2518 3236 2671 3240
rect 2500 3224 2692 3236
rect 2735 3224 2765 3238
rect 2771 3224 2784 3254
rect 2799 3236 2829 3254
rect 2872 3224 2885 3254
rect 2915 3224 2928 3254
rect 2943 3236 2973 3254
rect 3016 3240 3030 3254
rect 3066 3240 3286 3254
rect 3017 3238 3030 3240
rect 2983 3226 2998 3238
rect 2980 3224 3002 3226
rect 3007 3224 3037 3238
rect 3098 3236 3251 3240
rect 3080 3224 3272 3236
rect 3315 3224 3345 3238
rect 3351 3224 3364 3254
rect 3379 3236 3409 3254
rect 3452 3224 3465 3254
rect 3495 3224 3508 3254
rect 3523 3236 3553 3254
rect 3596 3240 3610 3254
rect 3646 3240 3866 3254
rect 3597 3238 3610 3240
rect 3563 3226 3578 3238
rect 3560 3224 3582 3226
rect 3587 3224 3617 3238
rect 3678 3236 3831 3240
rect 3660 3224 3852 3236
rect 3895 3224 3925 3238
rect 3931 3224 3944 3254
rect 3959 3236 3989 3254
rect 4032 3224 4045 3254
rect 4075 3224 4088 3254
rect 4103 3236 4133 3254
rect 4176 3240 4190 3254
rect 4226 3240 4446 3254
rect 4177 3238 4190 3240
rect 4143 3226 4158 3238
rect 4140 3224 4162 3226
rect 4167 3224 4197 3238
rect 4258 3236 4411 3240
rect 4240 3224 4432 3236
rect 4475 3224 4505 3238
rect 4511 3224 4524 3254
rect 4539 3236 4569 3254
rect 4612 3224 4625 3254
rect 0 3210 4625 3224
rect 15 3106 28 3210
rect 73 3188 74 3198
rect 89 3188 102 3198
rect 73 3184 102 3188
rect 107 3184 137 3210
rect 155 3196 171 3198
rect 243 3196 296 3210
rect 244 3194 308 3196
rect 351 3194 366 3210
rect 415 3207 445 3210
rect 415 3204 451 3207
rect 381 3196 397 3198
rect 155 3184 170 3188
rect 73 3182 170 3184
rect 198 3182 366 3194
rect 382 3184 397 3188
rect 415 3185 454 3204
rect 473 3198 480 3199
rect 479 3191 480 3198
rect 463 3188 464 3191
rect 479 3188 492 3191
rect 415 3184 445 3185
rect 454 3184 460 3185
rect 463 3184 492 3188
rect 382 3183 492 3184
rect 382 3182 498 3183
rect 57 3174 108 3182
rect 57 3162 82 3174
rect 89 3162 108 3174
rect 139 3174 189 3182
rect 139 3166 155 3174
rect 162 3172 189 3174
rect 198 3172 419 3182
rect 162 3162 419 3172
rect 448 3174 498 3182
rect 448 3165 464 3174
rect 57 3154 108 3162
rect 155 3154 419 3162
rect 445 3162 464 3165
rect 471 3162 498 3174
rect 445 3154 498 3162
rect 73 3146 74 3154
rect 89 3146 102 3154
rect 73 3138 89 3146
rect 70 3131 89 3134
rect 70 3122 92 3131
rect 43 3112 92 3122
rect 43 3106 73 3112
rect 92 3107 97 3112
rect 15 3090 89 3106
rect 107 3098 137 3154
rect 172 3144 380 3154
rect 415 3150 460 3154
rect 463 3153 464 3154
rect 479 3153 492 3154
rect 198 3114 387 3144
rect 213 3111 387 3114
rect 206 3108 387 3111
rect 15 3088 28 3090
rect 43 3088 77 3090
rect 15 3072 89 3088
rect 116 3084 129 3098
rect 144 3084 160 3100
rect 206 3095 217 3108
rect -1 3050 0 3066
rect 15 3050 28 3072
rect 43 3050 73 3072
rect 116 3068 178 3084
rect 206 3077 217 3093
rect 222 3088 232 3108
rect 242 3088 256 3108
rect 259 3095 268 3108
rect 284 3095 293 3108
rect 222 3077 256 3088
rect 259 3077 268 3093
rect 284 3077 293 3093
rect 300 3088 310 3108
rect 320 3088 334 3108
rect 335 3095 346 3108
rect 300 3077 334 3088
rect 335 3077 346 3093
rect 392 3084 408 3100
rect 415 3098 445 3150
rect 479 3146 480 3153
rect 464 3138 480 3146
rect 451 3106 464 3125
rect 479 3106 509 3122
rect 451 3090 525 3106
rect 451 3088 464 3090
rect 479 3088 513 3090
rect 116 3066 129 3068
rect 144 3066 178 3068
rect 116 3050 178 3066
rect 222 3061 238 3064
rect 300 3061 330 3072
rect 378 3068 424 3084
rect 451 3072 525 3088
rect 378 3066 412 3068
rect 377 3050 424 3066
rect 451 3050 464 3072
rect 479 3050 509 3072
rect 536 3050 537 3066
rect 552 3050 565 3210
rect 595 3106 608 3210
rect 653 3188 654 3198
rect 669 3188 682 3198
rect 653 3184 682 3188
rect 687 3184 717 3210
rect 735 3196 751 3198
rect 823 3196 876 3210
rect 824 3194 888 3196
rect 931 3194 946 3210
rect 995 3207 1025 3210
rect 995 3204 1031 3207
rect 961 3196 977 3198
rect 735 3184 750 3188
rect 653 3182 750 3184
rect 778 3182 946 3194
rect 962 3184 977 3188
rect 995 3185 1034 3204
rect 1053 3198 1060 3199
rect 1059 3191 1060 3198
rect 1043 3188 1044 3191
rect 1059 3188 1072 3191
rect 995 3184 1025 3185
rect 1034 3184 1040 3185
rect 1043 3184 1072 3188
rect 962 3183 1072 3184
rect 962 3182 1078 3183
rect 637 3174 688 3182
rect 637 3162 662 3174
rect 669 3162 688 3174
rect 719 3174 769 3182
rect 719 3166 735 3174
rect 742 3172 769 3174
rect 778 3172 999 3182
rect 742 3162 999 3172
rect 1028 3174 1078 3182
rect 1028 3165 1044 3174
rect 637 3154 688 3162
rect 735 3154 999 3162
rect 1025 3162 1044 3165
rect 1051 3162 1078 3174
rect 1025 3154 1078 3162
rect 653 3146 654 3154
rect 669 3146 682 3154
rect 653 3138 669 3146
rect 650 3131 669 3134
rect 650 3122 672 3131
rect 623 3112 672 3122
rect 623 3106 653 3112
rect 672 3107 677 3112
rect 595 3090 669 3106
rect 687 3098 717 3154
rect 752 3144 960 3154
rect 995 3150 1040 3154
rect 1043 3153 1044 3154
rect 1059 3153 1072 3154
rect 778 3114 967 3144
rect 793 3111 967 3114
rect 786 3108 967 3111
rect 595 3088 608 3090
rect 623 3088 657 3090
rect 595 3072 669 3088
rect 696 3084 709 3098
rect 724 3084 740 3100
rect 786 3095 797 3108
rect 579 3050 580 3066
rect 595 3050 608 3072
rect 623 3050 653 3072
rect 696 3068 758 3084
rect 786 3077 797 3093
rect 802 3088 812 3108
rect 822 3088 836 3108
rect 839 3095 848 3108
rect 864 3095 873 3108
rect 802 3077 836 3088
rect 839 3077 848 3093
rect 864 3077 873 3093
rect 880 3088 890 3108
rect 900 3088 914 3108
rect 915 3095 926 3108
rect 880 3077 914 3088
rect 915 3077 926 3093
rect 972 3084 988 3100
rect 995 3098 1025 3150
rect 1059 3146 1060 3153
rect 1044 3138 1060 3146
rect 1031 3106 1044 3125
rect 1059 3106 1089 3122
rect 1031 3090 1105 3106
rect 1031 3088 1044 3090
rect 1059 3088 1093 3090
rect 696 3066 709 3068
rect 724 3066 758 3068
rect 696 3050 758 3066
rect 802 3061 818 3064
rect 880 3061 910 3072
rect 958 3068 1004 3084
rect 1031 3072 1105 3088
rect 958 3066 992 3068
rect 957 3050 1004 3066
rect 1031 3050 1044 3072
rect 1059 3050 1089 3072
rect 1116 3050 1117 3066
rect 1132 3050 1145 3210
rect 1175 3106 1188 3210
rect 1233 3188 1234 3198
rect 1249 3188 1262 3198
rect 1233 3184 1262 3188
rect 1267 3184 1297 3210
rect 1315 3196 1331 3198
rect 1403 3196 1456 3210
rect 1404 3194 1468 3196
rect 1511 3194 1526 3210
rect 1575 3207 1605 3210
rect 1575 3204 1611 3207
rect 1541 3196 1557 3198
rect 1315 3184 1330 3188
rect 1233 3182 1330 3184
rect 1358 3182 1526 3194
rect 1542 3184 1557 3188
rect 1575 3185 1614 3204
rect 1633 3198 1640 3199
rect 1639 3191 1640 3198
rect 1623 3188 1624 3191
rect 1639 3188 1652 3191
rect 1575 3184 1605 3185
rect 1614 3184 1620 3185
rect 1623 3184 1652 3188
rect 1542 3183 1652 3184
rect 1542 3182 1658 3183
rect 1217 3174 1268 3182
rect 1217 3162 1242 3174
rect 1249 3162 1268 3174
rect 1299 3174 1349 3182
rect 1299 3166 1315 3174
rect 1322 3172 1349 3174
rect 1358 3172 1579 3182
rect 1322 3162 1579 3172
rect 1608 3174 1658 3182
rect 1608 3165 1624 3174
rect 1217 3154 1268 3162
rect 1315 3154 1579 3162
rect 1605 3162 1624 3165
rect 1631 3162 1658 3174
rect 1605 3154 1658 3162
rect 1233 3146 1234 3154
rect 1249 3146 1262 3154
rect 1233 3138 1249 3146
rect 1230 3131 1249 3134
rect 1230 3122 1252 3131
rect 1203 3112 1252 3122
rect 1203 3106 1233 3112
rect 1252 3107 1257 3112
rect 1175 3090 1249 3106
rect 1267 3098 1297 3154
rect 1332 3144 1540 3154
rect 1575 3150 1620 3154
rect 1623 3153 1624 3154
rect 1639 3153 1652 3154
rect 1358 3114 1547 3144
rect 1373 3111 1547 3114
rect 1366 3108 1547 3111
rect 1175 3088 1188 3090
rect 1203 3088 1237 3090
rect 1175 3072 1249 3088
rect 1276 3084 1289 3098
rect 1304 3084 1320 3100
rect 1366 3095 1377 3108
rect 1159 3050 1160 3066
rect 1175 3050 1188 3072
rect 1203 3050 1233 3072
rect 1276 3068 1338 3084
rect 1366 3077 1377 3093
rect 1382 3088 1392 3108
rect 1402 3088 1416 3108
rect 1419 3095 1428 3108
rect 1444 3095 1453 3108
rect 1382 3077 1416 3088
rect 1419 3077 1428 3093
rect 1444 3077 1453 3093
rect 1460 3088 1470 3108
rect 1480 3088 1494 3108
rect 1495 3095 1506 3108
rect 1460 3077 1494 3088
rect 1495 3077 1506 3093
rect 1552 3084 1568 3100
rect 1575 3098 1605 3150
rect 1639 3146 1640 3153
rect 1624 3138 1640 3146
rect 1611 3106 1624 3125
rect 1639 3106 1669 3122
rect 1611 3090 1685 3106
rect 1611 3088 1624 3090
rect 1639 3088 1673 3090
rect 1276 3066 1289 3068
rect 1304 3066 1338 3068
rect 1276 3050 1338 3066
rect 1382 3061 1398 3064
rect 1460 3061 1490 3072
rect 1538 3068 1584 3084
rect 1611 3072 1685 3088
rect 1538 3066 1572 3068
rect 1537 3050 1584 3066
rect 1611 3050 1624 3072
rect 1639 3050 1669 3072
rect 1696 3050 1697 3066
rect 1712 3050 1725 3210
rect 1755 3106 1768 3210
rect 1813 3188 1814 3198
rect 1829 3188 1842 3198
rect 1813 3184 1842 3188
rect 1847 3184 1877 3210
rect 1895 3196 1911 3198
rect 1983 3196 2036 3210
rect 1984 3194 2048 3196
rect 2091 3194 2106 3210
rect 2155 3207 2185 3210
rect 2155 3204 2191 3207
rect 2121 3196 2137 3198
rect 1895 3184 1910 3188
rect 1813 3182 1910 3184
rect 1938 3182 2106 3194
rect 2122 3184 2137 3188
rect 2155 3185 2194 3204
rect 2213 3198 2220 3199
rect 2219 3191 2220 3198
rect 2203 3188 2204 3191
rect 2219 3188 2232 3191
rect 2155 3184 2185 3185
rect 2194 3184 2200 3185
rect 2203 3184 2232 3188
rect 2122 3183 2232 3184
rect 2122 3182 2238 3183
rect 1797 3174 1848 3182
rect 1797 3162 1822 3174
rect 1829 3162 1848 3174
rect 1879 3174 1929 3182
rect 1879 3166 1895 3174
rect 1902 3172 1929 3174
rect 1938 3172 2159 3182
rect 1902 3162 2159 3172
rect 2188 3174 2238 3182
rect 2188 3165 2204 3174
rect 1797 3154 1848 3162
rect 1895 3154 2159 3162
rect 2185 3162 2204 3165
rect 2211 3162 2238 3174
rect 2185 3154 2238 3162
rect 1813 3146 1814 3154
rect 1829 3146 1842 3154
rect 1813 3138 1829 3146
rect 1810 3131 1829 3134
rect 1810 3122 1832 3131
rect 1783 3112 1832 3122
rect 1783 3106 1813 3112
rect 1832 3107 1837 3112
rect 1755 3090 1829 3106
rect 1847 3098 1877 3154
rect 1912 3144 2120 3154
rect 2155 3150 2200 3154
rect 2203 3153 2204 3154
rect 2219 3153 2232 3154
rect 1938 3114 2127 3144
rect 1953 3111 2127 3114
rect 1946 3108 2127 3111
rect 1755 3088 1768 3090
rect 1783 3088 1817 3090
rect 1755 3072 1829 3088
rect 1856 3084 1869 3098
rect 1884 3084 1900 3100
rect 1946 3095 1957 3108
rect 1739 3050 1740 3066
rect 1755 3050 1768 3072
rect 1783 3050 1813 3072
rect 1856 3068 1918 3084
rect 1946 3077 1957 3093
rect 1962 3088 1972 3108
rect 1982 3088 1996 3108
rect 1999 3095 2008 3108
rect 2024 3095 2033 3108
rect 1962 3077 1996 3088
rect 1999 3077 2008 3093
rect 2024 3077 2033 3093
rect 2040 3088 2050 3108
rect 2060 3088 2074 3108
rect 2075 3095 2086 3108
rect 2040 3077 2074 3088
rect 2075 3077 2086 3093
rect 2132 3084 2148 3100
rect 2155 3098 2185 3150
rect 2219 3146 2220 3153
rect 2204 3138 2220 3146
rect 2191 3106 2204 3125
rect 2219 3106 2249 3122
rect 2191 3090 2265 3106
rect 2191 3088 2204 3090
rect 2219 3088 2253 3090
rect 1856 3066 1869 3068
rect 1884 3066 1918 3068
rect 1856 3050 1918 3066
rect 1962 3061 1978 3064
rect 2040 3061 2070 3072
rect 2118 3068 2164 3084
rect 2191 3072 2265 3088
rect 2118 3066 2152 3068
rect 2117 3050 2164 3066
rect 2191 3050 2204 3072
rect 2219 3050 2249 3072
rect 2276 3050 2277 3066
rect 2292 3050 2305 3210
rect 2335 3106 2348 3210
rect 2393 3188 2394 3198
rect 2409 3188 2422 3198
rect 2393 3184 2422 3188
rect 2427 3184 2457 3210
rect 2475 3196 2491 3198
rect 2563 3196 2616 3210
rect 2564 3194 2628 3196
rect 2671 3194 2686 3210
rect 2735 3207 2765 3210
rect 2735 3204 2771 3207
rect 2701 3196 2717 3198
rect 2475 3184 2490 3188
rect 2393 3182 2490 3184
rect 2518 3182 2686 3194
rect 2702 3184 2717 3188
rect 2735 3185 2774 3204
rect 2793 3198 2800 3199
rect 2799 3191 2800 3198
rect 2783 3188 2784 3191
rect 2799 3188 2812 3191
rect 2735 3184 2765 3185
rect 2774 3184 2780 3185
rect 2783 3184 2812 3188
rect 2702 3183 2812 3184
rect 2702 3182 2818 3183
rect 2377 3174 2428 3182
rect 2377 3162 2402 3174
rect 2409 3162 2428 3174
rect 2459 3174 2509 3182
rect 2459 3166 2475 3174
rect 2482 3172 2509 3174
rect 2518 3172 2739 3182
rect 2482 3162 2739 3172
rect 2768 3174 2818 3182
rect 2768 3165 2784 3174
rect 2377 3154 2428 3162
rect 2475 3154 2739 3162
rect 2765 3162 2784 3165
rect 2791 3162 2818 3174
rect 2765 3154 2818 3162
rect 2393 3146 2394 3154
rect 2409 3146 2422 3154
rect 2393 3138 2409 3146
rect 2390 3131 2409 3134
rect 2390 3122 2412 3131
rect 2363 3112 2412 3122
rect 2363 3106 2393 3112
rect 2412 3107 2417 3112
rect 2335 3090 2409 3106
rect 2427 3098 2457 3154
rect 2492 3144 2700 3154
rect 2735 3150 2780 3154
rect 2783 3153 2784 3154
rect 2799 3153 2812 3154
rect 2518 3114 2707 3144
rect 2533 3111 2707 3114
rect 2526 3108 2707 3111
rect 2335 3088 2348 3090
rect 2363 3088 2397 3090
rect 2335 3072 2409 3088
rect 2436 3084 2449 3098
rect 2464 3084 2480 3100
rect 2526 3095 2537 3108
rect 2319 3050 2320 3066
rect 2335 3050 2348 3072
rect 2363 3050 2393 3072
rect 2436 3068 2498 3084
rect 2526 3077 2537 3093
rect 2542 3088 2552 3108
rect 2562 3088 2576 3108
rect 2579 3095 2588 3108
rect 2604 3095 2613 3108
rect 2542 3077 2576 3088
rect 2579 3077 2588 3093
rect 2604 3077 2613 3093
rect 2620 3088 2630 3108
rect 2640 3088 2654 3108
rect 2655 3095 2666 3108
rect 2620 3077 2654 3088
rect 2655 3077 2666 3093
rect 2712 3084 2728 3100
rect 2735 3098 2765 3150
rect 2799 3146 2800 3153
rect 2784 3138 2800 3146
rect 2771 3106 2784 3125
rect 2799 3106 2829 3122
rect 2771 3090 2845 3106
rect 2771 3088 2784 3090
rect 2799 3088 2833 3090
rect 2436 3066 2449 3068
rect 2464 3066 2498 3068
rect 2436 3050 2498 3066
rect 2542 3061 2558 3064
rect 2620 3061 2650 3072
rect 2698 3068 2744 3084
rect 2771 3072 2845 3088
rect 2698 3066 2732 3068
rect 2697 3050 2744 3066
rect 2771 3050 2784 3072
rect 2799 3050 2829 3072
rect 2856 3050 2857 3066
rect 2872 3050 2885 3210
rect 2915 3106 2928 3210
rect 2973 3188 2974 3198
rect 2989 3188 3002 3198
rect 2973 3184 3002 3188
rect 3007 3184 3037 3210
rect 3055 3196 3071 3198
rect 3143 3196 3196 3210
rect 3144 3194 3208 3196
rect 3251 3194 3266 3210
rect 3315 3207 3345 3210
rect 3315 3204 3351 3207
rect 3281 3196 3297 3198
rect 3055 3184 3070 3188
rect 2973 3182 3070 3184
rect 3098 3182 3266 3194
rect 3282 3184 3297 3188
rect 3315 3185 3354 3204
rect 3373 3198 3380 3199
rect 3379 3191 3380 3198
rect 3363 3188 3364 3191
rect 3379 3188 3392 3191
rect 3315 3184 3345 3185
rect 3354 3184 3360 3185
rect 3363 3184 3392 3188
rect 3282 3183 3392 3184
rect 3282 3182 3398 3183
rect 2957 3174 3008 3182
rect 2957 3162 2982 3174
rect 2989 3162 3008 3174
rect 3039 3174 3089 3182
rect 3039 3166 3055 3174
rect 3062 3172 3089 3174
rect 3098 3172 3319 3182
rect 3062 3162 3319 3172
rect 3348 3174 3398 3182
rect 3348 3165 3364 3174
rect 2957 3154 3008 3162
rect 3055 3154 3319 3162
rect 3345 3162 3364 3165
rect 3371 3162 3398 3174
rect 3345 3154 3398 3162
rect 2973 3146 2974 3154
rect 2989 3146 3002 3154
rect 2973 3138 2989 3146
rect 2970 3131 2989 3134
rect 2970 3122 2992 3131
rect 2943 3112 2992 3122
rect 2943 3106 2973 3112
rect 2992 3107 2997 3112
rect 2915 3090 2989 3106
rect 3007 3098 3037 3154
rect 3072 3144 3280 3154
rect 3315 3150 3360 3154
rect 3363 3153 3364 3154
rect 3379 3153 3392 3154
rect 3098 3114 3287 3144
rect 3113 3111 3287 3114
rect 3106 3108 3287 3111
rect 2915 3088 2928 3090
rect 2943 3088 2977 3090
rect 2915 3072 2989 3088
rect 3016 3084 3029 3098
rect 3044 3084 3060 3100
rect 3106 3095 3117 3108
rect 2899 3050 2900 3066
rect 2915 3050 2928 3072
rect 2943 3050 2973 3072
rect 3016 3068 3078 3084
rect 3106 3077 3117 3093
rect 3122 3088 3132 3108
rect 3142 3088 3156 3108
rect 3159 3095 3168 3108
rect 3184 3095 3193 3108
rect 3122 3077 3156 3088
rect 3159 3077 3168 3093
rect 3184 3077 3193 3093
rect 3200 3088 3210 3108
rect 3220 3088 3234 3108
rect 3235 3095 3246 3108
rect 3200 3077 3234 3088
rect 3235 3077 3246 3093
rect 3292 3084 3308 3100
rect 3315 3098 3345 3150
rect 3379 3146 3380 3153
rect 3364 3138 3380 3146
rect 3351 3106 3364 3125
rect 3379 3106 3409 3122
rect 3351 3090 3425 3106
rect 3351 3088 3364 3090
rect 3379 3088 3413 3090
rect 3016 3066 3029 3068
rect 3044 3066 3078 3068
rect 3016 3050 3078 3066
rect 3122 3061 3138 3064
rect 3200 3061 3230 3072
rect 3278 3068 3324 3084
rect 3351 3072 3425 3088
rect 3278 3066 3312 3068
rect 3277 3050 3324 3066
rect 3351 3050 3364 3072
rect 3379 3050 3409 3072
rect 3436 3050 3437 3066
rect 3452 3050 3465 3210
rect 3495 3106 3508 3210
rect 3553 3188 3554 3198
rect 3569 3188 3582 3198
rect 3553 3184 3582 3188
rect 3587 3184 3617 3210
rect 3635 3196 3651 3198
rect 3723 3196 3776 3210
rect 3724 3194 3788 3196
rect 3831 3194 3846 3210
rect 3895 3207 3925 3210
rect 3895 3204 3931 3207
rect 3861 3196 3877 3198
rect 3635 3184 3650 3188
rect 3553 3182 3650 3184
rect 3678 3182 3846 3194
rect 3862 3184 3877 3188
rect 3895 3185 3934 3204
rect 3953 3198 3960 3199
rect 3959 3191 3960 3198
rect 3943 3188 3944 3191
rect 3959 3188 3972 3191
rect 3895 3184 3925 3185
rect 3934 3184 3940 3185
rect 3943 3184 3972 3188
rect 3862 3183 3972 3184
rect 3862 3182 3978 3183
rect 3537 3174 3588 3182
rect 3537 3162 3562 3174
rect 3569 3162 3588 3174
rect 3619 3174 3669 3182
rect 3619 3166 3635 3174
rect 3642 3172 3669 3174
rect 3678 3172 3899 3182
rect 3642 3162 3899 3172
rect 3928 3174 3978 3182
rect 3928 3165 3944 3174
rect 3537 3154 3588 3162
rect 3635 3154 3899 3162
rect 3925 3162 3944 3165
rect 3951 3162 3978 3174
rect 3925 3154 3978 3162
rect 3553 3146 3554 3154
rect 3569 3146 3582 3154
rect 3553 3138 3569 3146
rect 3550 3131 3569 3134
rect 3550 3122 3572 3131
rect 3523 3112 3572 3122
rect 3523 3106 3553 3112
rect 3572 3107 3577 3112
rect 3495 3090 3569 3106
rect 3587 3098 3617 3154
rect 3652 3144 3860 3154
rect 3895 3150 3940 3154
rect 3943 3153 3944 3154
rect 3959 3153 3972 3154
rect 3678 3114 3867 3144
rect 3693 3111 3867 3114
rect 3686 3108 3867 3111
rect 3495 3088 3508 3090
rect 3523 3088 3557 3090
rect 3495 3072 3569 3088
rect 3596 3084 3609 3098
rect 3624 3084 3640 3100
rect 3686 3095 3697 3108
rect 3479 3050 3480 3066
rect 3495 3050 3508 3072
rect 3523 3050 3553 3072
rect 3596 3068 3658 3084
rect 3686 3077 3697 3093
rect 3702 3088 3712 3108
rect 3722 3088 3736 3108
rect 3739 3095 3748 3108
rect 3764 3095 3773 3108
rect 3702 3077 3736 3088
rect 3739 3077 3748 3093
rect 3764 3077 3773 3093
rect 3780 3088 3790 3108
rect 3800 3088 3814 3108
rect 3815 3095 3826 3108
rect 3780 3077 3814 3088
rect 3815 3077 3826 3093
rect 3872 3084 3888 3100
rect 3895 3098 3925 3150
rect 3959 3146 3960 3153
rect 3944 3138 3960 3146
rect 3931 3106 3944 3125
rect 3959 3106 3989 3122
rect 3931 3090 4005 3106
rect 3931 3088 3944 3090
rect 3959 3088 3993 3090
rect 3596 3066 3609 3068
rect 3624 3066 3658 3068
rect 3596 3050 3658 3066
rect 3702 3061 3718 3064
rect 3780 3061 3810 3072
rect 3858 3068 3904 3084
rect 3931 3072 4005 3088
rect 3858 3066 3892 3068
rect 3857 3050 3904 3066
rect 3931 3050 3944 3072
rect 3959 3050 3989 3072
rect 4016 3050 4017 3066
rect 4032 3050 4045 3210
rect 4075 3106 4088 3210
rect 4133 3188 4134 3198
rect 4149 3188 4162 3198
rect 4133 3184 4162 3188
rect 4167 3184 4197 3210
rect 4215 3196 4231 3198
rect 4303 3196 4356 3210
rect 4304 3194 4368 3196
rect 4411 3194 4426 3210
rect 4475 3207 4505 3210
rect 4475 3204 4511 3207
rect 4441 3196 4457 3198
rect 4215 3184 4230 3188
rect 4133 3182 4230 3184
rect 4258 3182 4426 3194
rect 4442 3184 4457 3188
rect 4475 3185 4514 3204
rect 4533 3198 4540 3199
rect 4539 3191 4540 3198
rect 4523 3188 4524 3191
rect 4539 3188 4552 3191
rect 4475 3184 4505 3185
rect 4514 3184 4520 3185
rect 4523 3184 4552 3188
rect 4442 3183 4552 3184
rect 4442 3182 4558 3183
rect 4117 3174 4168 3182
rect 4117 3162 4142 3174
rect 4149 3162 4168 3174
rect 4199 3174 4249 3182
rect 4199 3166 4215 3174
rect 4222 3172 4249 3174
rect 4258 3172 4479 3182
rect 4222 3162 4479 3172
rect 4508 3174 4558 3182
rect 4508 3165 4524 3174
rect 4117 3154 4168 3162
rect 4215 3154 4479 3162
rect 4505 3162 4524 3165
rect 4531 3162 4558 3174
rect 4505 3154 4558 3162
rect 4133 3146 4134 3154
rect 4149 3146 4162 3154
rect 4133 3138 4149 3146
rect 4130 3131 4149 3134
rect 4130 3122 4152 3131
rect 4103 3112 4152 3122
rect 4103 3106 4133 3112
rect 4152 3107 4157 3112
rect 4075 3090 4149 3106
rect 4167 3098 4197 3154
rect 4232 3144 4440 3154
rect 4475 3150 4520 3154
rect 4523 3153 4524 3154
rect 4539 3153 4552 3154
rect 4258 3114 4447 3144
rect 4273 3111 4447 3114
rect 4266 3108 4447 3111
rect 4075 3088 4088 3090
rect 4103 3088 4137 3090
rect 4075 3072 4149 3088
rect 4176 3084 4189 3098
rect 4204 3084 4220 3100
rect 4266 3095 4277 3108
rect 4059 3050 4060 3066
rect 4075 3050 4088 3072
rect 4103 3050 4133 3072
rect 4176 3068 4238 3084
rect 4266 3077 4277 3093
rect 4282 3088 4292 3108
rect 4302 3088 4316 3108
rect 4319 3095 4328 3108
rect 4344 3095 4353 3108
rect 4282 3077 4316 3088
rect 4319 3077 4328 3093
rect 4344 3077 4353 3093
rect 4360 3088 4370 3108
rect 4380 3088 4394 3108
rect 4395 3095 4406 3108
rect 4360 3077 4394 3088
rect 4395 3077 4406 3093
rect 4452 3084 4468 3100
rect 4475 3098 4505 3150
rect 4539 3146 4540 3153
rect 4524 3138 4540 3146
rect 4511 3106 4524 3125
rect 4539 3106 4569 3122
rect 4511 3090 4585 3106
rect 4511 3088 4524 3090
rect 4539 3088 4573 3090
rect 4176 3066 4189 3068
rect 4204 3066 4238 3068
rect 4176 3050 4238 3066
rect 4282 3061 4298 3064
rect 4360 3061 4390 3072
rect 4438 3068 4484 3084
rect 4511 3072 4585 3088
rect 4438 3066 4472 3068
rect 4437 3050 4484 3066
rect 4511 3050 4524 3072
rect 4539 3050 4569 3072
rect 4596 3050 4597 3066
rect 4612 3050 4625 3210
rect -7 3042 34 3050
rect -7 3016 8 3042
rect 15 3016 34 3042
rect 98 3038 160 3050
rect 172 3038 247 3050
rect 305 3038 380 3050
rect 392 3038 423 3050
rect 429 3038 464 3050
rect 98 3036 260 3038
rect -7 3008 34 3016
rect 116 3012 129 3036
rect 144 3034 159 3036
rect -1 2998 0 3008
rect 15 2998 28 3008
rect 43 2998 73 3012
rect 116 2998 159 3012
rect 183 3009 190 3016
rect 193 3012 260 3036
rect 292 3036 464 3038
rect 262 3014 290 3018
rect 292 3014 372 3036
rect 393 3034 408 3036
rect 262 3012 372 3014
rect 193 3008 372 3012
rect 166 2998 196 3008
rect 198 2998 351 3008
rect 359 2998 389 3008
rect 393 2998 423 3012
rect 451 2998 464 3036
rect 536 3042 571 3050
rect 536 3016 537 3042
rect 544 3016 571 3042
rect 479 2998 509 3012
rect 536 3008 571 3016
rect 573 3042 614 3050
rect 573 3016 588 3042
rect 595 3016 614 3042
rect 678 3038 740 3050
rect 752 3038 827 3050
rect 885 3038 960 3050
rect 972 3038 1003 3050
rect 1009 3038 1044 3050
rect 678 3036 840 3038
rect 573 3008 614 3016
rect 696 3012 709 3036
rect 724 3034 739 3036
rect 536 2998 537 3008
rect 552 2998 565 3008
rect 579 2998 580 3008
rect 595 2998 608 3008
rect 623 2998 653 3012
rect 696 2998 739 3012
rect 763 3009 770 3016
rect 773 3012 840 3036
rect 872 3036 1044 3038
rect 842 3014 870 3018
rect 872 3014 952 3036
rect 973 3034 988 3036
rect 842 3012 952 3014
rect 773 3008 952 3012
rect 746 2998 776 3008
rect 778 2998 931 3008
rect 939 2998 969 3008
rect 973 2998 1003 3012
rect 1031 2998 1044 3036
rect 1116 3042 1151 3050
rect 1116 3016 1117 3042
rect 1124 3016 1151 3042
rect 1059 2998 1089 3012
rect 1116 3008 1151 3016
rect 1153 3042 1194 3050
rect 1153 3016 1168 3042
rect 1175 3016 1194 3042
rect 1258 3038 1320 3050
rect 1332 3038 1407 3050
rect 1465 3038 1540 3050
rect 1552 3038 1583 3050
rect 1589 3038 1624 3050
rect 1258 3036 1420 3038
rect 1153 3008 1194 3016
rect 1276 3012 1289 3036
rect 1304 3034 1319 3036
rect 1116 2998 1117 3008
rect 1132 2998 1145 3008
rect 1159 2998 1160 3008
rect 1175 2998 1188 3008
rect 1203 2998 1233 3012
rect 1276 2998 1319 3012
rect 1343 3009 1350 3016
rect 1353 3012 1420 3036
rect 1452 3036 1624 3038
rect 1422 3014 1450 3018
rect 1452 3014 1532 3036
rect 1553 3034 1568 3036
rect 1422 3012 1532 3014
rect 1353 3008 1532 3012
rect 1326 2998 1356 3008
rect 1358 2998 1511 3008
rect 1519 2998 1549 3008
rect 1553 2998 1583 3012
rect 1611 2998 1624 3036
rect 1696 3042 1731 3050
rect 1696 3016 1697 3042
rect 1704 3016 1731 3042
rect 1639 2998 1669 3012
rect 1696 3008 1731 3016
rect 1733 3042 1774 3050
rect 1733 3016 1748 3042
rect 1755 3016 1774 3042
rect 1838 3038 1900 3050
rect 1912 3038 1987 3050
rect 2045 3038 2120 3050
rect 2132 3038 2163 3050
rect 2169 3038 2204 3050
rect 1838 3036 2000 3038
rect 1733 3008 1774 3016
rect 1856 3012 1869 3036
rect 1884 3034 1899 3036
rect 1696 2998 1697 3008
rect 1712 2998 1725 3008
rect 1739 2998 1740 3008
rect 1755 2998 1768 3008
rect 1783 2998 1813 3012
rect 1856 2998 1899 3012
rect 1923 3009 1930 3016
rect 1933 3012 2000 3036
rect 2032 3036 2204 3038
rect 2002 3014 2030 3018
rect 2032 3014 2112 3036
rect 2133 3034 2148 3036
rect 2002 3012 2112 3014
rect 1933 3008 2112 3012
rect 1906 2998 1936 3008
rect 1938 2998 2091 3008
rect 2099 2998 2129 3008
rect 2133 2998 2163 3012
rect 2191 2998 2204 3036
rect 2276 3042 2311 3050
rect 2276 3016 2277 3042
rect 2284 3016 2311 3042
rect 2219 2998 2249 3012
rect 2276 3008 2311 3016
rect 2313 3042 2354 3050
rect 2313 3016 2328 3042
rect 2335 3016 2354 3042
rect 2418 3038 2480 3050
rect 2492 3038 2567 3050
rect 2625 3038 2700 3050
rect 2712 3038 2743 3050
rect 2749 3038 2784 3050
rect 2418 3036 2580 3038
rect 2313 3008 2354 3016
rect 2436 3012 2449 3036
rect 2464 3034 2479 3036
rect 2276 2998 2277 3008
rect 2292 2998 2305 3008
rect 2319 2998 2320 3008
rect 2335 2998 2348 3008
rect 2363 2998 2393 3012
rect 2436 2998 2479 3012
rect 2503 3009 2510 3016
rect 2513 3012 2580 3036
rect 2612 3036 2784 3038
rect 2582 3014 2610 3018
rect 2612 3014 2692 3036
rect 2713 3034 2728 3036
rect 2582 3012 2692 3014
rect 2513 3008 2692 3012
rect 2486 2998 2516 3008
rect 2518 2998 2671 3008
rect 2679 2998 2709 3008
rect 2713 2998 2743 3012
rect 2771 2998 2784 3036
rect 2856 3042 2891 3050
rect 2856 3016 2857 3042
rect 2864 3016 2891 3042
rect 2799 2998 2829 3012
rect 2856 3008 2891 3016
rect 2893 3042 2934 3050
rect 2893 3016 2908 3042
rect 2915 3016 2934 3042
rect 2998 3038 3060 3050
rect 3072 3038 3147 3050
rect 3205 3038 3280 3050
rect 3292 3038 3323 3050
rect 3329 3038 3364 3050
rect 2998 3036 3160 3038
rect 2893 3008 2934 3016
rect 3016 3012 3029 3036
rect 3044 3034 3059 3036
rect 2856 2998 2857 3008
rect 2872 2998 2885 3008
rect 2899 2998 2900 3008
rect 2915 2998 2928 3008
rect 2943 2998 2973 3012
rect 3016 2998 3059 3012
rect 3083 3009 3090 3016
rect 3093 3012 3160 3036
rect 3192 3036 3364 3038
rect 3162 3014 3190 3018
rect 3192 3014 3272 3036
rect 3293 3034 3308 3036
rect 3162 3012 3272 3014
rect 3093 3008 3272 3012
rect 3066 2998 3096 3008
rect 3098 2998 3251 3008
rect 3259 2998 3289 3008
rect 3293 2998 3323 3012
rect 3351 2998 3364 3036
rect 3436 3042 3471 3050
rect 3436 3016 3437 3042
rect 3444 3016 3471 3042
rect 3379 2998 3409 3012
rect 3436 3008 3471 3016
rect 3473 3042 3514 3050
rect 3473 3016 3488 3042
rect 3495 3016 3514 3042
rect 3578 3038 3640 3050
rect 3652 3038 3727 3050
rect 3785 3038 3860 3050
rect 3872 3038 3903 3050
rect 3909 3038 3944 3050
rect 3578 3036 3740 3038
rect 3473 3008 3514 3016
rect 3596 3012 3609 3036
rect 3624 3034 3639 3036
rect 3436 2998 3437 3008
rect 3452 2998 3465 3008
rect 3479 2998 3480 3008
rect 3495 2998 3508 3008
rect 3523 2998 3553 3012
rect 3596 2998 3639 3012
rect 3663 3009 3670 3016
rect 3673 3012 3740 3036
rect 3772 3036 3944 3038
rect 3742 3014 3770 3018
rect 3772 3014 3852 3036
rect 3873 3034 3888 3036
rect 3742 3012 3852 3014
rect 3673 3008 3852 3012
rect 3646 2998 3676 3008
rect 3678 2998 3831 3008
rect 3839 2998 3869 3008
rect 3873 2998 3903 3012
rect 3931 2998 3944 3036
rect 4016 3042 4051 3050
rect 4016 3016 4017 3042
rect 4024 3016 4051 3042
rect 3959 2998 3989 3012
rect 4016 3008 4051 3016
rect 4053 3042 4094 3050
rect 4053 3016 4068 3042
rect 4075 3016 4094 3042
rect 4158 3038 4220 3050
rect 4232 3038 4307 3050
rect 4365 3038 4440 3050
rect 4452 3038 4483 3050
rect 4489 3038 4524 3050
rect 4158 3036 4320 3038
rect 4053 3008 4094 3016
rect 4176 3012 4189 3036
rect 4204 3034 4219 3036
rect 4016 2998 4017 3008
rect 4032 2998 4045 3008
rect 4059 2998 4060 3008
rect 4075 2998 4088 3008
rect 4103 2998 4133 3012
rect 4176 2998 4219 3012
rect 4243 3009 4250 3016
rect 4253 3012 4320 3036
rect 4352 3036 4524 3038
rect 4322 3014 4350 3018
rect 4352 3014 4432 3036
rect 4453 3034 4468 3036
rect 4322 3012 4432 3014
rect 4253 3008 4432 3012
rect 4226 2998 4256 3008
rect 4258 2998 4411 3008
rect 4419 2998 4449 3008
rect 4453 2998 4483 3012
rect 4511 2998 4524 3036
rect 4596 3042 4631 3050
rect 4596 3016 4597 3042
rect 4604 3016 4631 3042
rect 4539 2998 4569 3012
rect 4596 3008 4631 3016
rect 4596 2998 4597 3008
rect 4612 2998 4625 3008
rect -1 2992 4625 2998
rect 0 2984 4625 2992
rect 15 2954 28 2984
rect 43 2966 73 2984
rect 116 2970 130 2984
rect 166 2970 386 2984
rect 117 2968 130 2970
rect 83 2956 98 2968
rect 80 2954 102 2956
rect 107 2954 137 2968
rect 198 2966 351 2970
rect 180 2954 372 2966
rect 415 2954 445 2968
rect 451 2954 464 2984
rect 479 2966 509 2984
rect 552 2954 565 2984
rect 595 2954 608 2984
rect 623 2966 653 2984
rect 696 2970 710 2984
rect 746 2970 966 2984
rect 697 2968 710 2970
rect 663 2956 678 2968
rect 660 2954 682 2956
rect 687 2954 717 2968
rect 778 2966 931 2970
rect 760 2954 952 2966
rect 995 2954 1025 2968
rect 1031 2954 1044 2984
rect 1059 2966 1089 2984
rect 1132 2954 1145 2984
rect 1175 2954 1188 2984
rect 1203 2966 1233 2984
rect 1276 2970 1290 2984
rect 1326 2970 1546 2984
rect 1277 2968 1290 2970
rect 1243 2956 1258 2968
rect 1240 2954 1262 2956
rect 1267 2954 1297 2968
rect 1358 2966 1511 2970
rect 1340 2954 1532 2966
rect 1575 2954 1605 2968
rect 1611 2954 1624 2984
rect 1639 2966 1669 2984
rect 1712 2954 1725 2984
rect 1755 2954 1768 2984
rect 1783 2966 1813 2984
rect 1856 2970 1870 2984
rect 1906 2970 2126 2984
rect 1857 2968 1870 2970
rect 1823 2956 1838 2968
rect 1820 2954 1842 2956
rect 1847 2954 1877 2968
rect 1938 2966 2091 2970
rect 1920 2954 2112 2966
rect 2155 2954 2185 2968
rect 2191 2954 2204 2984
rect 2219 2966 2249 2984
rect 2292 2954 2305 2984
rect 2335 2954 2348 2984
rect 2363 2966 2393 2984
rect 2436 2970 2450 2984
rect 2486 2970 2706 2984
rect 2437 2968 2450 2970
rect 2403 2956 2418 2968
rect 2400 2954 2422 2956
rect 2427 2954 2457 2968
rect 2518 2966 2671 2970
rect 2500 2954 2692 2966
rect 2735 2954 2765 2968
rect 2771 2954 2784 2984
rect 2799 2966 2829 2984
rect 2872 2954 2885 2984
rect 2915 2954 2928 2984
rect 2943 2966 2973 2984
rect 3016 2970 3030 2984
rect 3066 2970 3286 2984
rect 3017 2968 3030 2970
rect 2983 2956 2998 2968
rect 2980 2954 3002 2956
rect 3007 2954 3037 2968
rect 3098 2966 3251 2970
rect 3080 2954 3272 2966
rect 3315 2954 3345 2968
rect 3351 2954 3364 2984
rect 3379 2966 3409 2984
rect 3452 2954 3465 2984
rect 3495 2954 3508 2984
rect 3523 2966 3553 2984
rect 3596 2970 3610 2984
rect 3646 2970 3866 2984
rect 3597 2968 3610 2970
rect 3563 2956 3578 2968
rect 3560 2954 3582 2956
rect 3587 2954 3617 2968
rect 3678 2966 3831 2970
rect 3660 2954 3852 2966
rect 3895 2954 3925 2968
rect 3931 2954 3944 2984
rect 3959 2966 3989 2984
rect 4032 2954 4045 2984
rect 4075 2954 4088 2984
rect 4103 2966 4133 2984
rect 4176 2970 4190 2984
rect 4226 2970 4446 2984
rect 4177 2968 4190 2970
rect 4143 2956 4158 2968
rect 4140 2954 4162 2956
rect 4167 2954 4197 2968
rect 4258 2966 4411 2970
rect 4240 2954 4432 2966
rect 4475 2954 4505 2968
rect 4511 2954 4524 2984
rect 4539 2966 4569 2984
rect 4612 2954 4625 2984
rect 0 2940 4625 2954
rect 15 2836 28 2940
rect 73 2918 74 2928
rect 89 2918 102 2928
rect 73 2914 102 2918
rect 107 2914 137 2940
rect 155 2926 171 2928
rect 243 2926 296 2940
rect 244 2924 308 2926
rect 351 2924 366 2940
rect 415 2937 445 2940
rect 415 2934 451 2937
rect 381 2926 397 2928
rect 155 2914 170 2918
rect 73 2912 170 2914
rect 198 2912 366 2924
rect 382 2914 397 2918
rect 415 2915 454 2934
rect 473 2928 480 2929
rect 479 2921 480 2928
rect 463 2918 464 2921
rect 479 2918 492 2921
rect 415 2914 445 2915
rect 454 2914 460 2915
rect 463 2914 492 2918
rect 382 2913 492 2914
rect 382 2912 498 2913
rect 57 2904 108 2912
rect 57 2892 82 2904
rect 89 2892 108 2904
rect 139 2904 189 2912
rect 139 2896 155 2904
rect 162 2902 189 2904
rect 198 2902 419 2912
rect 162 2892 419 2902
rect 448 2904 498 2912
rect 448 2895 464 2904
rect 57 2884 108 2892
rect 155 2884 419 2892
rect 445 2892 464 2895
rect 471 2892 498 2904
rect 445 2884 498 2892
rect 73 2876 74 2884
rect 89 2876 102 2884
rect 73 2868 89 2876
rect 70 2861 89 2864
rect 70 2852 92 2861
rect 43 2842 92 2852
rect 43 2836 73 2842
rect 92 2837 97 2842
rect 15 2820 89 2836
rect 107 2828 137 2884
rect 172 2874 380 2884
rect 415 2880 460 2884
rect 463 2883 464 2884
rect 479 2883 492 2884
rect 198 2844 387 2874
rect 213 2841 387 2844
rect 206 2838 387 2841
rect 15 2818 28 2820
rect 43 2818 77 2820
rect 15 2802 89 2818
rect 116 2814 129 2828
rect 144 2814 160 2830
rect 206 2825 217 2838
rect -1 2780 0 2796
rect 15 2780 28 2802
rect 43 2780 73 2802
rect 116 2798 178 2814
rect 206 2807 217 2823
rect 222 2818 232 2838
rect 242 2818 256 2838
rect 259 2825 268 2838
rect 284 2825 293 2838
rect 222 2807 256 2818
rect 259 2807 268 2823
rect 284 2807 293 2823
rect 300 2818 310 2838
rect 320 2818 334 2838
rect 335 2825 346 2838
rect 300 2807 334 2818
rect 335 2807 346 2823
rect 392 2814 408 2830
rect 415 2828 445 2880
rect 479 2876 480 2883
rect 464 2868 480 2876
rect 451 2836 464 2855
rect 479 2836 509 2852
rect 451 2820 525 2836
rect 451 2818 464 2820
rect 479 2818 513 2820
rect 116 2796 129 2798
rect 144 2796 178 2798
rect 116 2780 178 2796
rect 222 2791 238 2794
rect 300 2791 330 2802
rect 378 2798 424 2814
rect 451 2802 525 2818
rect 378 2796 412 2798
rect 377 2780 424 2796
rect 451 2780 464 2802
rect 479 2780 509 2802
rect 536 2780 537 2796
rect 552 2780 565 2940
rect 595 2836 608 2940
rect 653 2918 654 2928
rect 669 2918 682 2928
rect 653 2914 682 2918
rect 687 2914 717 2940
rect 735 2926 751 2928
rect 823 2926 876 2940
rect 824 2924 888 2926
rect 931 2924 946 2940
rect 995 2937 1025 2940
rect 995 2934 1031 2937
rect 961 2926 977 2928
rect 735 2914 750 2918
rect 653 2912 750 2914
rect 778 2912 946 2924
rect 962 2914 977 2918
rect 995 2915 1034 2934
rect 1053 2928 1060 2929
rect 1059 2921 1060 2928
rect 1043 2918 1044 2921
rect 1059 2918 1072 2921
rect 995 2914 1025 2915
rect 1034 2914 1040 2915
rect 1043 2914 1072 2918
rect 962 2913 1072 2914
rect 962 2912 1078 2913
rect 637 2904 688 2912
rect 637 2892 662 2904
rect 669 2892 688 2904
rect 719 2904 769 2912
rect 719 2896 735 2904
rect 742 2902 769 2904
rect 778 2902 999 2912
rect 742 2892 999 2902
rect 1028 2904 1078 2912
rect 1028 2895 1044 2904
rect 637 2884 688 2892
rect 735 2884 999 2892
rect 1025 2892 1044 2895
rect 1051 2892 1078 2904
rect 1025 2884 1078 2892
rect 653 2876 654 2884
rect 669 2876 682 2884
rect 653 2868 669 2876
rect 650 2861 669 2864
rect 650 2852 672 2861
rect 623 2842 672 2852
rect 623 2836 653 2842
rect 672 2837 677 2842
rect 595 2820 669 2836
rect 687 2828 717 2884
rect 752 2874 960 2884
rect 995 2880 1040 2884
rect 1043 2883 1044 2884
rect 1059 2883 1072 2884
rect 778 2844 967 2874
rect 793 2841 967 2844
rect 786 2838 967 2841
rect 595 2818 608 2820
rect 623 2818 657 2820
rect 595 2802 669 2818
rect 696 2814 709 2828
rect 724 2814 740 2830
rect 786 2825 797 2838
rect 579 2780 580 2796
rect 595 2780 608 2802
rect 623 2780 653 2802
rect 696 2798 758 2814
rect 786 2807 797 2823
rect 802 2818 812 2838
rect 822 2818 836 2838
rect 839 2825 848 2838
rect 864 2825 873 2838
rect 802 2807 836 2818
rect 839 2807 848 2823
rect 864 2807 873 2823
rect 880 2818 890 2838
rect 900 2818 914 2838
rect 915 2825 926 2838
rect 880 2807 914 2818
rect 915 2807 926 2823
rect 972 2814 988 2830
rect 995 2828 1025 2880
rect 1059 2876 1060 2883
rect 1044 2868 1060 2876
rect 1031 2836 1044 2855
rect 1059 2836 1089 2852
rect 1031 2820 1105 2836
rect 1031 2818 1044 2820
rect 1059 2818 1093 2820
rect 696 2796 709 2798
rect 724 2796 758 2798
rect 696 2780 758 2796
rect 802 2791 818 2794
rect 880 2791 910 2802
rect 958 2798 1004 2814
rect 1031 2802 1105 2818
rect 958 2796 992 2798
rect 957 2780 1004 2796
rect 1031 2780 1044 2802
rect 1059 2780 1089 2802
rect 1116 2780 1117 2796
rect 1132 2780 1145 2940
rect 1175 2836 1188 2940
rect 1233 2918 1234 2928
rect 1249 2918 1262 2928
rect 1233 2914 1262 2918
rect 1267 2914 1297 2940
rect 1315 2926 1331 2928
rect 1403 2926 1456 2940
rect 1404 2924 1468 2926
rect 1511 2924 1526 2940
rect 1575 2937 1605 2940
rect 1575 2934 1611 2937
rect 1541 2926 1557 2928
rect 1315 2914 1330 2918
rect 1233 2912 1330 2914
rect 1358 2912 1526 2924
rect 1542 2914 1557 2918
rect 1575 2915 1614 2934
rect 1633 2928 1640 2929
rect 1639 2921 1640 2928
rect 1623 2918 1624 2921
rect 1639 2918 1652 2921
rect 1575 2914 1605 2915
rect 1614 2914 1620 2915
rect 1623 2914 1652 2918
rect 1542 2913 1652 2914
rect 1542 2912 1658 2913
rect 1217 2904 1268 2912
rect 1217 2892 1242 2904
rect 1249 2892 1268 2904
rect 1299 2904 1349 2912
rect 1299 2896 1315 2904
rect 1322 2902 1349 2904
rect 1358 2902 1579 2912
rect 1322 2892 1579 2902
rect 1608 2904 1658 2912
rect 1608 2895 1624 2904
rect 1217 2884 1268 2892
rect 1315 2884 1579 2892
rect 1605 2892 1624 2895
rect 1631 2892 1658 2904
rect 1605 2884 1658 2892
rect 1233 2876 1234 2884
rect 1249 2876 1262 2884
rect 1233 2868 1249 2876
rect 1230 2861 1249 2864
rect 1230 2852 1252 2861
rect 1203 2842 1252 2852
rect 1203 2836 1233 2842
rect 1252 2837 1257 2842
rect 1175 2820 1249 2836
rect 1267 2828 1297 2884
rect 1332 2874 1540 2884
rect 1575 2880 1620 2884
rect 1623 2883 1624 2884
rect 1639 2883 1652 2884
rect 1358 2844 1547 2874
rect 1373 2841 1547 2844
rect 1366 2838 1547 2841
rect 1175 2818 1188 2820
rect 1203 2818 1237 2820
rect 1175 2802 1249 2818
rect 1276 2814 1289 2828
rect 1304 2814 1320 2830
rect 1366 2825 1377 2838
rect 1159 2780 1160 2796
rect 1175 2780 1188 2802
rect 1203 2780 1233 2802
rect 1276 2798 1338 2814
rect 1366 2807 1377 2823
rect 1382 2818 1392 2838
rect 1402 2818 1416 2838
rect 1419 2825 1428 2838
rect 1444 2825 1453 2838
rect 1382 2807 1416 2818
rect 1419 2807 1428 2823
rect 1444 2807 1453 2823
rect 1460 2818 1470 2838
rect 1480 2818 1494 2838
rect 1495 2825 1506 2838
rect 1460 2807 1494 2818
rect 1495 2807 1506 2823
rect 1552 2814 1568 2830
rect 1575 2828 1605 2880
rect 1639 2876 1640 2883
rect 1624 2868 1640 2876
rect 1611 2836 1624 2855
rect 1639 2836 1669 2852
rect 1611 2820 1685 2836
rect 1611 2818 1624 2820
rect 1639 2818 1673 2820
rect 1276 2796 1289 2798
rect 1304 2796 1338 2798
rect 1276 2780 1338 2796
rect 1382 2791 1398 2794
rect 1460 2791 1490 2802
rect 1538 2798 1584 2814
rect 1611 2802 1685 2818
rect 1538 2796 1572 2798
rect 1537 2780 1584 2796
rect 1611 2780 1624 2802
rect 1639 2780 1669 2802
rect 1696 2780 1697 2796
rect 1712 2780 1725 2940
rect 1755 2836 1768 2940
rect 1813 2918 1814 2928
rect 1829 2918 1842 2928
rect 1813 2914 1842 2918
rect 1847 2914 1877 2940
rect 1895 2926 1911 2928
rect 1983 2926 2036 2940
rect 1984 2924 2048 2926
rect 2091 2924 2106 2940
rect 2155 2937 2185 2940
rect 2155 2934 2191 2937
rect 2121 2926 2137 2928
rect 1895 2914 1910 2918
rect 1813 2912 1910 2914
rect 1938 2912 2106 2924
rect 2122 2914 2137 2918
rect 2155 2915 2194 2934
rect 2213 2928 2220 2929
rect 2219 2921 2220 2928
rect 2203 2918 2204 2921
rect 2219 2918 2232 2921
rect 2155 2914 2185 2915
rect 2194 2914 2200 2915
rect 2203 2914 2232 2918
rect 2122 2913 2232 2914
rect 2122 2912 2238 2913
rect 1797 2904 1848 2912
rect 1797 2892 1822 2904
rect 1829 2892 1848 2904
rect 1879 2904 1929 2912
rect 1879 2896 1895 2904
rect 1902 2902 1929 2904
rect 1938 2902 2159 2912
rect 1902 2892 2159 2902
rect 2188 2904 2238 2912
rect 2188 2895 2204 2904
rect 1797 2884 1848 2892
rect 1895 2884 2159 2892
rect 2185 2892 2204 2895
rect 2211 2892 2238 2904
rect 2185 2884 2238 2892
rect 1813 2876 1814 2884
rect 1829 2876 1842 2884
rect 1813 2868 1829 2876
rect 1810 2861 1829 2864
rect 1810 2852 1832 2861
rect 1783 2842 1832 2852
rect 1783 2836 1813 2842
rect 1832 2837 1837 2842
rect 1755 2820 1829 2836
rect 1847 2828 1877 2884
rect 1912 2874 2120 2884
rect 2155 2880 2200 2884
rect 2203 2883 2204 2884
rect 2219 2883 2232 2884
rect 1938 2844 2127 2874
rect 1953 2841 2127 2844
rect 1946 2838 2127 2841
rect 1755 2818 1768 2820
rect 1783 2818 1817 2820
rect 1755 2802 1829 2818
rect 1856 2814 1869 2828
rect 1884 2814 1900 2830
rect 1946 2825 1957 2838
rect 1739 2780 1740 2796
rect 1755 2780 1768 2802
rect 1783 2780 1813 2802
rect 1856 2798 1918 2814
rect 1946 2807 1957 2823
rect 1962 2818 1972 2838
rect 1982 2818 1996 2838
rect 1999 2825 2008 2838
rect 2024 2825 2033 2838
rect 1962 2807 1996 2818
rect 1999 2807 2008 2823
rect 2024 2807 2033 2823
rect 2040 2818 2050 2838
rect 2060 2818 2074 2838
rect 2075 2825 2086 2838
rect 2040 2807 2074 2818
rect 2075 2807 2086 2823
rect 2132 2814 2148 2830
rect 2155 2828 2185 2880
rect 2219 2876 2220 2883
rect 2204 2868 2220 2876
rect 2191 2836 2204 2855
rect 2219 2836 2249 2852
rect 2191 2820 2265 2836
rect 2191 2818 2204 2820
rect 2219 2818 2253 2820
rect 1856 2796 1869 2798
rect 1884 2796 1918 2798
rect 1856 2780 1918 2796
rect 1962 2791 1978 2794
rect 2040 2791 2070 2802
rect 2118 2798 2164 2814
rect 2191 2802 2265 2818
rect 2118 2796 2152 2798
rect 2117 2780 2164 2796
rect 2191 2780 2204 2802
rect 2219 2780 2249 2802
rect 2276 2780 2277 2796
rect 2292 2780 2305 2940
rect 2335 2836 2348 2940
rect 2393 2918 2394 2928
rect 2409 2918 2422 2928
rect 2393 2914 2422 2918
rect 2427 2914 2457 2940
rect 2475 2926 2491 2928
rect 2563 2926 2616 2940
rect 2564 2924 2628 2926
rect 2671 2924 2686 2940
rect 2735 2937 2765 2940
rect 2735 2934 2771 2937
rect 2701 2926 2717 2928
rect 2475 2914 2490 2918
rect 2393 2912 2490 2914
rect 2518 2912 2686 2924
rect 2702 2914 2717 2918
rect 2735 2915 2774 2934
rect 2793 2928 2800 2929
rect 2799 2921 2800 2928
rect 2783 2918 2784 2921
rect 2799 2918 2812 2921
rect 2735 2914 2765 2915
rect 2774 2914 2780 2915
rect 2783 2914 2812 2918
rect 2702 2913 2812 2914
rect 2702 2912 2818 2913
rect 2377 2904 2428 2912
rect 2377 2892 2402 2904
rect 2409 2892 2428 2904
rect 2459 2904 2509 2912
rect 2459 2896 2475 2904
rect 2482 2902 2509 2904
rect 2518 2902 2739 2912
rect 2482 2892 2739 2902
rect 2768 2904 2818 2912
rect 2768 2895 2784 2904
rect 2377 2884 2428 2892
rect 2475 2884 2739 2892
rect 2765 2892 2784 2895
rect 2791 2892 2818 2904
rect 2765 2884 2818 2892
rect 2393 2876 2394 2884
rect 2409 2876 2422 2884
rect 2393 2868 2409 2876
rect 2390 2861 2409 2864
rect 2390 2852 2412 2861
rect 2363 2842 2412 2852
rect 2363 2836 2393 2842
rect 2412 2837 2417 2842
rect 2335 2820 2409 2836
rect 2427 2828 2457 2884
rect 2492 2874 2700 2884
rect 2735 2880 2780 2884
rect 2783 2883 2784 2884
rect 2799 2883 2812 2884
rect 2518 2844 2707 2874
rect 2533 2841 2707 2844
rect 2526 2838 2707 2841
rect 2335 2818 2348 2820
rect 2363 2818 2397 2820
rect 2335 2802 2409 2818
rect 2436 2814 2449 2828
rect 2464 2814 2480 2830
rect 2526 2825 2537 2838
rect 2319 2780 2320 2796
rect 2335 2780 2348 2802
rect 2363 2780 2393 2802
rect 2436 2798 2498 2814
rect 2526 2807 2537 2823
rect 2542 2818 2552 2838
rect 2562 2818 2576 2838
rect 2579 2825 2588 2838
rect 2604 2825 2613 2838
rect 2542 2807 2576 2818
rect 2579 2807 2588 2823
rect 2604 2807 2613 2823
rect 2620 2818 2630 2838
rect 2640 2818 2654 2838
rect 2655 2825 2666 2838
rect 2620 2807 2654 2818
rect 2655 2807 2666 2823
rect 2712 2814 2728 2830
rect 2735 2828 2765 2880
rect 2799 2876 2800 2883
rect 2784 2868 2800 2876
rect 2771 2836 2784 2855
rect 2799 2836 2829 2852
rect 2771 2820 2845 2836
rect 2771 2818 2784 2820
rect 2799 2818 2833 2820
rect 2436 2796 2449 2798
rect 2464 2796 2498 2798
rect 2436 2780 2498 2796
rect 2542 2791 2558 2794
rect 2620 2791 2650 2802
rect 2698 2798 2744 2814
rect 2771 2802 2845 2818
rect 2698 2796 2732 2798
rect 2697 2780 2744 2796
rect 2771 2780 2784 2802
rect 2799 2780 2829 2802
rect 2856 2780 2857 2796
rect 2872 2780 2885 2940
rect 2915 2836 2928 2940
rect 2973 2918 2974 2928
rect 2989 2918 3002 2928
rect 2973 2914 3002 2918
rect 3007 2914 3037 2940
rect 3055 2926 3071 2928
rect 3143 2926 3196 2940
rect 3144 2924 3208 2926
rect 3251 2924 3266 2940
rect 3315 2937 3345 2940
rect 3315 2934 3351 2937
rect 3281 2926 3297 2928
rect 3055 2914 3070 2918
rect 2973 2912 3070 2914
rect 3098 2912 3266 2924
rect 3282 2914 3297 2918
rect 3315 2915 3354 2934
rect 3373 2928 3380 2929
rect 3379 2921 3380 2928
rect 3363 2918 3364 2921
rect 3379 2918 3392 2921
rect 3315 2914 3345 2915
rect 3354 2914 3360 2915
rect 3363 2914 3392 2918
rect 3282 2913 3392 2914
rect 3282 2912 3398 2913
rect 2957 2904 3008 2912
rect 2957 2892 2982 2904
rect 2989 2892 3008 2904
rect 3039 2904 3089 2912
rect 3039 2896 3055 2904
rect 3062 2902 3089 2904
rect 3098 2902 3319 2912
rect 3062 2892 3319 2902
rect 3348 2904 3398 2912
rect 3348 2895 3364 2904
rect 2957 2884 3008 2892
rect 3055 2884 3319 2892
rect 3345 2892 3364 2895
rect 3371 2892 3398 2904
rect 3345 2884 3398 2892
rect 2973 2876 2974 2884
rect 2989 2876 3002 2884
rect 2973 2868 2989 2876
rect 2970 2861 2989 2864
rect 2970 2852 2992 2861
rect 2943 2842 2992 2852
rect 2943 2836 2973 2842
rect 2992 2837 2997 2842
rect 2915 2820 2989 2836
rect 3007 2828 3037 2884
rect 3072 2874 3280 2884
rect 3315 2880 3360 2884
rect 3363 2883 3364 2884
rect 3379 2883 3392 2884
rect 3098 2844 3287 2874
rect 3113 2841 3287 2844
rect 3106 2838 3287 2841
rect 2915 2818 2928 2820
rect 2943 2818 2977 2820
rect 2915 2802 2989 2818
rect 3016 2814 3029 2828
rect 3044 2814 3060 2830
rect 3106 2825 3117 2838
rect 2899 2780 2900 2796
rect 2915 2780 2928 2802
rect 2943 2780 2973 2802
rect 3016 2798 3078 2814
rect 3106 2807 3117 2823
rect 3122 2818 3132 2838
rect 3142 2818 3156 2838
rect 3159 2825 3168 2838
rect 3184 2825 3193 2838
rect 3122 2807 3156 2818
rect 3159 2807 3168 2823
rect 3184 2807 3193 2823
rect 3200 2818 3210 2838
rect 3220 2818 3234 2838
rect 3235 2825 3246 2838
rect 3200 2807 3234 2818
rect 3235 2807 3246 2823
rect 3292 2814 3308 2830
rect 3315 2828 3345 2880
rect 3379 2876 3380 2883
rect 3364 2868 3380 2876
rect 3351 2836 3364 2855
rect 3379 2836 3409 2852
rect 3351 2820 3425 2836
rect 3351 2818 3364 2820
rect 3379 2818 3413 2820
rect 3016 2796 3029 2798
rect 3044 2796 3078 2798
rect 3016 2780 3078 2796
rect 3122 2791 3138 2794
rect 3200 2791 3230 2802
rect 3278 2798 3324 2814
rect 3351 2802 3425 2818
rect 3278 2796 3312 2798
rect 3277 2780 3324 2796
rect 3351 2780 3364 2802
rect 3379 2780 3409 2802
rect 3436 2780 3437 2796
rect 3452 2780 3465 2940
rect 3495 2836 3508 2940
rect 3553 2918 3554 2928
rect 3569 2918 3582 2928
rect 3553 2914 3582 2918
rect 3587 2914 3617 2940
rect 3635 2926 3651 2928
rect 3723 2926 3776 2940
rect 3724 2924 3788 2926
rect 3831 2924 3846 2940
rect 3895 2937 3925 2940
rect 3895 2934 3931 2937
rect 3861 2926 3877 2928
rect 3635 2914 3650 2918
rect 3553 2912 3650 2914
rect 3678 2912 3846 2924
rect 3862 2914 3877 2918
rect 3895 2915 3934 2934
rect 3953 2928 3960 2929
rect 3959 2921 3960 2928
rect 3943 2918 3944 2921
rect 3959 2918 3972 2921
rect 3895 2914 3925 2915
rect 3934 2914 3940 2915
rect 3943 2914 3972 2918
rect 3862 2913 3972 2914
rect 3862 2912 3978 2913
rect 3537 2904 3588 2912
rect 3537 2892 3562 2904
rect 3569 2892 3588 2904
rect 3619 2904 3669 2912
rect 3619 2896 3635 2904
rect 3642 2902 3669 2904
rect 3678 2902 3899 2912
rect 3642 2892 3899 2902
rect 3928 2904 3978 2912
rect 3928 2895 3944 2904
rect 3537 2884 3588 2892
rect 3635 2884 3899 2892
rect 3925 2892 3944 2895
rect 3951 2892 3978 2904
rect 3925 2884 3978 2892
rect 3553 2876 3554 2884
rect 3569 2876 3582 2884
rect 3553 2868 3569 2876
rect 3550 2861 3569 2864
rect 3550 2852 3572 2861
rect 3523 2842 3572 2852
rect 3523 2836 3553 2842
rect 3572 2837 3577 2842
rect 3495 2820 3569 2836
rect 3587 2828 3617 2884
rect 3652 2874 3860 2884
rect 3895 2880 3940 2884
rect 3943 2883 3944 2884
rect 3959 2883 3972 2884
rect 3678 2844 3867 2874
rect 3693 2841 3867 2844
rect 3686 2838 3867 2841
rect 3495 2818 3508 2820
rect 3523 2818 3557 2820
rect 3495 2802 3569 2818
rect 3596 2814 3609 2828
rect 3624 2814 3640 2830
rect 3686 2825 3697 2838
rect 3479 2780 3480 2796
rect 3495 2780 3508 2802
rect 3523 2780 3553 2802
rect 3596 2798 3658 2814
rect 3686 2807 3697 2823
rect 3702 2818 3712 2838
rect 3722 2818 3736 2838
rect 3739 2825 3748 2838
rect 3764 2825 3773 2838
rect 3702 2807 3736 2818
rect 3739 2807 3748 2823
rect 3764 2807 3773 2823
rect 3780 2818 3790 2838
rect 3800 2818 3814 2838
rect 3815 2825 3826 2838
rect 3780 2807 3814 2818
rect 3815 2807 3826 2823
rect 3872 2814 3888 2830
rect 3895 2828 3925 2880
rect 3959 2876 3960 2883
rect 3944 2868 3960 2876
rect 3931 2836 3944 2855
rect 3959 2836 3989 2852
rect 3931 2820 4005 2836
rect 3931 2818 3944 2820
rect 3959 2818 3993 2820
rect 3596 2796 3609 2798
rect 3624 2796 3658 2798
rect 3596 2780 3658 2796
rect 3702 2791 3718 2794
rect 3780 2791 3810 2802
rect 3858 2798 3904 2814
rect 3931 2802 4005 2818
rect 3858 2796 3892 2798
rect 3857 2780 3904 2796
rect 3931 2780 3944 2802
rect 3959 2780 3989 2802
rect 4016 2780 4017 2796
rect 4032 2780 4045 2940
rect 4075 2836 4088 2940
rect 4133 2918 4134 2928
rect 4149 2918 4162 2928
rect 4133 2914 4162 2918
rect 4167 2914 4197 2940
rect 4215 2926 4231 2928
rect 4303 2926 4356 2940
rect 4304 2924 4368 2926
rect 4411 2924 4426 2940
rect 4475 2937 4505 2940
rect 4475 2934 4511 2937
rect 4441 2926 4457 2928
rect 4215 2914 4230 2918
rect 4133 2912 4230 2914
rect 4258 2912 4426 2924
rect 4442 2914 4457 2918
rect 4475 2915 4514 2934
rect 4533 2928 4540 2929
rect 4539 2921 4540 2928
rect 4523 2918 4524 2921
rect 4539 2918 4552 2921
rect 4475 2914 4505 2915
rect 4514 2914 4520 2915
rect 4523 2914 4552 2918
rect 4442 2913 4552 2914
rect 4442 2912 4558 2913
rect 4117 2904 4168 2912
rect 4117 2892 4142 2904
rect 4149 2892 4168 2904
rect 4199 2904 4249 2912
rect 4199 2896 4215 2904
rect 4222 2902 4249 2904
rect 4258 2902 4479 2912
rect 4222 2892 4479 2902
rect 4508 2904 4558 2912
rect 4508 2895 4524 2904
rect 4117 2884 4168 2892
rect 4215 2884 4479 2892
rect 4505 2892 4524 2895
rect 4531 2892 4558 2904
rect 4505 2884 4558 2892
rect 4133 2876 4134 2884
rect 4149 2876 4162 2884
rect 4133 2868 4149 2876
rect 4130 2861 4149 2864
rect 4130 2852 4152 2861
rect 4103 2842 4152 2852
rect 4103 2836 4133 2842
rect 4152 2837 4157 2842
rect 4075 2820 4149 2836
rect 4167 2828 4197 2884
rect 4232 2874 4440 2884
rect 4475 2880 4520 2884
rect 4523 2883 4524 2884
rect 4539 2883 4552 2884
rect 4258 2844 4447 2874
rect 4273 2841 4447 2844
rect 4266 2838 4447 2841
rect 4075 2818 4088 2820
rect 4103 2818 4137 2820
rect 4075 2802 4149 2818
rect 4176 2814 4189 2828
rect 4204 2814 4220 2830
rect 4266 2825 4277 2838
rect 4059 2780 4060 2796
rect 4075 2780 4088 2802
rect 4103 2780 4133 2802
rect 4176 2798 4238 2814
rect 4266 2807 4277 2823
rect 4282 2818 4292 2838
rect 4302 2818 4316 2838
rect 4319 2825 4328 2838
rect 4344 2825 4353 2838
rect 4282 2807 4316 2818
rect 4319 2807 4328 2823
rect 4344 2807 4353 2823
rect 4360 2818 4370 2838
rect 4380 2818 4394 2838
rect 4395 2825 4406 2838
rect 4360 2807 4394 2818
rect 4395 2807 4406 2823
rect 4452 2814 4468 2830
rect 4475 2828 4505 2880
rect 4539 2876 4540 2883
rect 4524 2868 4540 2876
rect 4511 2836 4524 2855
rect 4539 2836 4569 2852
rect 4511 2820 4585 2836
rect 4511 2818 4524 2820
rect 4539 2818 4573 2820
rect 4176 2796 4189 2798
rect 4204 2796 4238 2798
rect 4176 2780 4238 2796
rect 4282 2791 4298 2794
rect 4360 2791 4390 2802
rect 4438 2798 4484 2814
rect 4511 2802 4585 2818
rect 4438 2796 4472 2798
rect 4437 2780 4484 2796
rect 4511 2780 4524 2802
rect 4539 2780 4569 2802
rect 4596 2780 4597 2796
rect 4612 2780 4625 2940
rect -7 2772 34 2780
rect -7 2746 8 2772
rect 15 2746 34 2772
rect 98 2768 160 2780
rect 172 2768 247 2780
rect 305 2768 380 2780
rect 392 2768 423 2780
rect 429 2768 464 2780
rect 98 2766 260 2768
rect -7 2738 34 2746
rect 116 2742 129 2766
rect 144 2764 159 2766
rect -1 2728 0 2738
rect 15 2728 28 2738
rect 43 2728 73 2742
rect 116 2728 159 2742
rect 183 2739 190 2746
rect 193 2742 260 2766
rect 292 2766 464 2768
rect 262 2744 290 2748
rect 292 2744 372 2766
rect 393 2764 408 2766
rect 262 2742 372 2744
rect 193 2738 372 2742
rect 166 2728 196 2738
rect 198 2728 351 2738
rect 359 2728 389 2738
rect 393 2728 423 2742
rect 451 2728 464 2766
rect 536 2772 571 2780
rect 536 2746 537 2772
rect 544 2746 571 2772
rect 479 2728 509 2742
rect 536 2738 571 2746
rect 573 2772 614 2780
rect 573 2746 588 2772
rect 595 2746 614 2772
rect 678 2768 740 2780
rect 752 2768 827 2780
rect 885 2768 960 2780
rect 972 2768 1003 2780
rect 1009 2768 1044 2780
rect 678 2766 840 2768
rect 573 2738 614 2746
rect 696 2742 709 2766
rect 724 2764 739 2766
rect 536 2728 537 2738
rect 552 2728 565 2738
rect 579 2728 580 2738
rect 595 2728 608 2738
rect 623 2728 653 2742
rect 696 2728 739 2742
rect 763 2739 770 2746
rect 773 2742 840 2766
rect 872 2766 1044 2768
rect 842 2744 870 2748
rect 872 2744 952 2766
rect 973 2764 988 2766
rect 842 2742 952 2744
rect 773 2738 952 2742
rect 746 2728 776 2738
rect 778 2728 931 2738
rect 939 2728 969 2738
rect 973 2728 1003 2742
rect 1031 2728 1044 2766
rect 1116 2772 1151 2780
rect 1116 2746 1117 2772
rect 1124 2746 1151 2772
rect 1059 2728 1089 2742
rect 1116 2738 1151 2746
rect 1153 2772 1194 2780
rect 1153 2746 1168 2772
rect 1175 2746 1194 2772
rect 1258 2768 1320 2780
rect 1332 2768 1407 2780
rect 1465 2768 1540 2780
rect 1552 2768 1583 2780
rect 1589 2768 1624 2780
rect 1258 2766 1420 2768
rect 1153 2738 1194 2746
rect 1276 2742 1289 2766
rect 1304 2764 1319 2766
rect 1116 2728 1117 2738
rect 1132 2728 1145 2738
rect 1159 2728 1160 2738
rect 1175 2728 1188 2738
rect 1203 2728 1233 2742
rect 1276 2728 1319 2742
rect 1343 2739 1350 2746
rect 1353 2742 1420 2766
rect 1452 2766 1624 2768
rect 1422 2744 1450 2748
rect 1452 2744 1532 2766
rect 1553 2764 1568 2766
rect 1422 2742 1532 2744
rect 1353 2738 1532 2742
rect 1326 2728 1356 2738
rect 1358 2728 1511 2738
rect 1519 2728 1549 2738
rect 1553 2728 1583 2742
rect 1611 2728 1624 2766
rect 1696 2772 1731 2780
rect 1696 2746 1697 2772
rect 1704 2746 1731 2772
rect 1639 2728 1669 2742
rect 1696 2738 1731 2746
rect 1733 2772 1774 2780
rect 1733 2746 1748 2772
rect 1755 2746 1774 2772
rect 1838 2768 1900 2780
rect 1912 2768 1987 2780
rect 2045 2768 2120 2780
rect 2132 2768 2163 2780
rect 2169 2768 2204 2780
rect 1838 2766 2000 2768
rect 1733 2738 1774 2746
rect 1856 2742 1869 2766
rect 1884 2764 1899 2766
rect 1696 2728 1697 2738
rect 1712 2728 1725 2738
rect 1739 2728 1740 2738
rect 1755 2728 1768 2738
rect 1783 2728 1813 2742
rect 1856 2728 1899 2742
rect 1923 2739 1930 2746
rect 1933 2742 2000 2766
rect 2032 2766 2204 2768
rect 2002 2744 2030 2748
rect 2032 2744 2112 2766
rect 2133 2764 2148 2766
rect 2002 2742 2112 2744
rect 1933 2738 2112 2742
rect 1906 2728 1936 2738
rect 1938 2728 2091 2738
rect 2099 2728 2129 2738
rect 2133 2728 2163 2742
rect 2191 2728 2204 2766
rect 2276 2772 2311 2780
rect 2276 2746 2277 2772
rect 2284 2746 2311 2772
rect 2219 2728 2249 2742
rect 2276 2738 2311 2746
rect 2313 2772 2354 2780
rect 2313 2746 2328 2772
rect 2335 2746 2354 2772
rect 2418 2768 2480 2780
rect 2492 2768 2567 2780
rect 2625 2768 2700 2780
rect 2712 2768 2743 2780
rect 2749 2768 2784 2780
rect 2418 2766 2580 2768
rect 2313 2738 2354 2746
rect 2436 2742 2449 2766
rect 2464 2764 2479 2766
rect 2276 2728 2277 2738
rect 2292 2728 2305 2738
rect 2319 2728 2320 2738
rect 2335 2728 2348 2738
rect 2363 2728 2393 2742
rect 2436 2728 2479 2742
rect 2503 2739 2510 2746
rect 2513 2742 2580 2766
rect 2612 2766 2784 2768
rect 2582 2744 2610 2748
rect 2612 2744 2692 2766
rect 2713 2764 2728 2766
rect 2582 2742 2692 2744
rect 2513 2738 2692 2742
rect 2486 2728 2516 2738
rect 2518 2728 2671 2738
rect 2679 2728 2709 2738
rect 2713 2728 2743 2742
rect 2771 2728 2784 2766
rect 2856 2772 2891 2780
rect 2856 2746 2857 2772
rect 2864 2746 2891 2772
rect 2799 2728 2829 2742
rect 2856 2738 2891 2746
rect 2893 2772 2934 2780
rect 2893 2746 2908 2772
rect 2915 2746 2934 2772
rect 2998 2768 3060 2780
rect 3072 2768 3147 2780
rect 3205 2768 3280 2780
rect 3292 2768 3323 2780
rect 3329 2768 3364 2780
rect 2998 2766 3160 2768
rect 2893 2738 2934 2746
rect 3016 2742 3029 2766
rect 3044 2764 3059 2766
rect 2856 2728 2857 2738
rect 2872 2728 2885 2738
rect 2899 2728 2900 2738
rect 2915 2728 2928 2738
rect 2943 2728 2973 2742
rect 3016 2728 3059 2742
rect 3083 2739 3090 2746
rect 3093 2742 3160 2766
rect 3192 2766 3364 2768
rect 3162 2744 3190 2748
rect 3192 2744 3272 2766
rect 3293 2764 3308 2766
rect 3162 2742 3272 2744
rect 3093 2738 3272 2742
rect 3066 2728 3096 2738
rect 3098 2728 3251 2738
rect 3259 2728 3289 2738
rect 3293 2728 3323 2742
rect 3351 2728 3364 2766
rect 3436 2772 3471 2780
rect 3436 2746 3437 2772
rect 3444 2746 3471 2772
rect 3379 2728 3409 2742
rect 3436 2738 3471 2746
rect 3473 2772 3514 2780
rect 3473 2746 3488 2772
rect 3495 2746 3514 2772
rect 3578 2768 3640 2780
rect 3652 2768 3727 2780
rect 3785 2768 3860 2780
rect 3872 2768 3903 2780
rect 3909 2768 3944 2780
rect 3578 2766 3740 2768
rect 3473 2738 3514 2746
rect 3596 2742 3609 2766
rect 3624 2764 3639 2766
rect 3436 2728 3437 2738
rect 3452 2728 3465 2738
rect 3479 2728 3480 2738
rect 3495 2728 3508 2738
rect 3523 2728 3553 2742
rect 3596 2728 3639 2742
rect 3663 2739 3670 2746
rect 3673 2742 3740 2766
rect 3772 2766 3944 2768
rect 3742 2744 3770 2748
rect 3772 2744 3852 2766
rect 3873 2764 3888 2766
rect 3742 2742 3852 2744
rect 3673 2738 3852 2742
rect 3646 2728 3676 2738
rect 3678 2728 3831 2738
rect 3839 2728 3869 2738
rect 3873 2728 3903 2742
rect 3931 2728 3944 2766
rect 4016 2772 4051 2780
rect 4016 2746 4017 2772
rect 4024 2746 4051 2772
rect 3959 2728 3989 2742
rect 4016 2738 4051 2746
rect 4053 2772 4094 2780
rect 4053 2746 4068 2772
rect 4075 2746 4094 2772
rect 4158 2768 4220 2780
rect 4232 2768 4307 2780
rect 4365 2768 4440 2780
rect 4452 2768 4483 2780
rect 4489 2768 4524 2780
rect 4158 2766 4320 2768
rect 4053 2738 4094 2746
rect 4176 2742 4189 2766
rect 4204 2764 4219 2766
rect 4016 2728 4017 2738
rect 4032 2728 4045 2738
rect 4059 2728 4060 2738
rect 4075 2728 4088 2738
rect 4103 2728 4133 2742
rect 4176 2728 4219 2742
rect 4243 2739 4250 2746
rect 4253 2742 4320 2766
rect 4352 2766 4524 2768
rect 4322 2744 4350 2748
rect 4352 2744 4432 2766
rect 4453 2764 4468 2766
rect 4322 2742 4432 2744
rect 4253 2738 4432 2742
rect 4226 2728 4256 2738
rect 4258 2728 4411 2738
rect 4419 2728 4449 2738
rect 4453 2728 4483 2742
rect 4511 2728 4524 2766
rect 4596 2772 4631 2780
rect 4596 2746 4597 2772
rect 4604 2746 4631 2772
rect 4539 2728 4569 2742
rect 4596 2738 4631 2746
rect 4596 2728 4597 2738
rect 4612 2728 4625 2738
rect -1 2722 4625 2728
rect 0 2714 4625 2722
rect 15 2684 28 2714
rect 43 2696 73 2714
rect 116 2700 130 2714
rect 166 2700 386 2714
rect 117 2698 130 2700
rect 83 2686 98 2698
rect 80 2684 102 2686
rect 107 2684 137 2698
rect 198 2696 351 2700
rect 180 2684 372 2696
rect 415 2684 445 2698
rect 451 2684 464 2714
rect 479 2696 509 2714
rect 552 2684 565 2714
rect 595 2684 608 2714
rect 623 2696 653 2714
rect 696 2700 710 2714
rect 746 2700 966 2714
rect 697 2698 710 2700
rect 663 2686 678 2698
rect 660 2684 682 2686
rect 687 2684 717 2698
rect 778 2696 931 2700
rect 760 2684 952 2696
rect 995 2684 1025 2698
rect 1031 2684 1044 2714
rect 1059 2696 1089 2714
rect 1132 2684 1145 2714
rect 1175 2684 1188 2714
rect 1203 2696 1233 2714
rect 1276 2700 1290 2714
rect 1326 2700 1546 2714
rect 1277 2698 1290 2700
rect 1243 2686 1258 2698
rect 1240 2684 1262 2686
rect 1267 2684 1297 2698
rect 1358 2696 1511 2700
rect 1340 2684 1532 2696
rect 1575 2684 1605 2698
rect 1611 2684 1624 2714
rect 1639 2696 1669 2714
rect 1712 2684 1725 2714
rect 1755 2684 1768 2714
rect 1783 2696 1813 2714
rect 1856 2700 1870 2714
rect 1906 2700 2126 2714
rect 1857 2698 1870 2700
rect 1823 2686 1838 2698
rect 1820 2684 1842 2686
rect 1847 2684 1877 2698
rect 1938 2696 2091 2700
rect 1920 2684 2112 2696
rect 2155 2684 2185 2698
rect 2191 2684 2204 2714
rect 2219 2696 2249 2714
rect 2292 2684 2305 2714
rect 2335 2684 2348 2714
rect 2363 2696 2393 2714
rect 2436 2700 2450 2714
rect 2486 2700 2706 2714
rect 2437 2698 2450 2700
rect 2403 2686 2418 2698
rect 2400 2684 2422 2686
rect 2427 2684 2457 2698
rect 2518 2696 2671 2700
rect 2500 2684 2692 2696
rect 2735 2684 2765 2698
rect 2771 2684 2784 2714
rect 2799 2696 2829 2714
rect 2872 2684 2885 2714
rect 2915 2684 2928 2714
rect 2943 2696 2973 2714
rect 3016 2700 3030 2714
rect 3066 2700 3286 2714
rect 3017 2698 3030 2700
rect 2983 2686 2998 2698
rect 2980 2684 3002 2686
rect 3007 2684 3037 2698
rect 3098 2696 3251 2700
rect 3080 2684 3272 2696
rect 3315 2684 3345 2698
rect 3351 2684 3364 2714
rect 3379 2696 3409 2714
rect 3452 2684 3465 2714
rect 3495 2684 3508 2714
rect 3523 2696 3553 2714
rect 3596 2700 3610 2714
rect 3646 2700 3866 2714
rect 3597 2698 3610 2700
rect 3563 2686 3578 2698
rect 3560 2684 3582 2686
rect 3587 2684 3617 2698
rect 3678 2696 3831 2700
rect 3660 2684 3852 2696
rect 3895 2684 3925 2698
rect 3931 2684 3944 2714
rect 3959 2696 3989 2714
rect 4032 2684 4045 2714
rect 4075 2684 4088 2714
rect 4103 2696 4133 2714
rect 4176 2700 4190 2714
rect 4226 2700 4446 2714
rect 4177 2698 4190 2700
rect 4143 2686 4158 2698
rect 4140 2684 4162 2686
rect 4167 2684 4197 2698
rect 4258 2696 4411 2700
rect 4240 2684 4432 2696
rect 4475 2684 4505 2698
rect 4511 2684 4524 2714
rect 4539 2696 4569 2714
rect 4612 2684 4625 2714
rect 0 2670 4625 2684
rect 15 2566 28 2670
rect 73 2648 74 2658
rect 89 2648 102 2658
rect 73 2644 102 2648
rect 107 2644 137 2670
rect 155 2656 171 2658
rect 243 2656 296 2670
rect 244 2654 308 2656
rect 351 2654 366 2670
rect 415 2667 445 2670
rect 415 2664 451 2667
rect 381 2656 397 2658
rect 155 2644 170 2648
rect 73 2642 170 2644
rect 198 2642 366 2654
rect 382 2644 397 2648
rect 415 2645 454 2664
rect 473 2658 480 2659
rect 479 2651 480 2658
rect 463 2648 464 2651
rect 479 2648 492 2651
rect 415 2644 445 2645
rect 454 2644 460 2645
rect 463 2644 492 2648
rect 382 2643 492 2644
rect 382 2642 498 2643
rect 57 2634 108 2642
rect 57 2622 82 2634
rect 89 2622 108 2634
rect 139 2634 189 2642
rect 139 2626 155 2634
rect 162 2632 189 2634
rect 198 2632 419 2642
rect 162 2622 419 2632
rect 448 2634 498 2642
rect 448 2625 464 2634
rect 57 2614 108 2622
rect 155 2614 419 2622
rect 445 2622 464 2625
rect 471 2622 498 2634
rect 445 2614 498 2622
rect 73 2606 74 2614
rect 89 2606 102 2614
rect 73 2598 89 2606
rect 70 2591 89 2594
rect 70 2582 92 2591
rect 43 2572 92 2582
rect 43 2566 73 2572
rect 92 2567 97 2572
rect 15 2550 89 2566
rect 107 2558 137 2614
rect 172 2604 380 2614
rect 415 2610 460 2614
rect 463 2613 464 2614
rect 479 2613 492 2614
rect 198 2574 387 2604
rect 213 2571 387 2574
rect 206 2568 387 2571
rect 15 2548 28 2550
rect 43 2548 77 2550
rect 15 2532 89 2548
rect 116 2544 129 2558
rect 144 2544 160 2560
rect 206 2555 217 2568
rect -1 2510 0 2526
rect 15 2510 28 2532
rect 43 2510 73 2532
rect 116 2528 178 2544
rect 206 2537 217 2553
rect 222 2548 232 2568
rect 242 2548 256 2568
rect 259 2555 268 2568
rect 284 2555 293 2568
rect 222 2537 256 2548
rect 259 2537 268 2553
rect 284 2537 293 2553
rect 300 2548 310 2568
rect 320 2548 334 2568
rect 335 2555 346 2568
rect 300 2537 334 2548
rect 335 2537 346 2553
rect 392 2544 408 2560
rect 415 2558 445 2610
rect 479 2606 480 2613
rect 464 2598 480 2606
rect 451 2566 464 2585
rect 479 2566 509 2582
rect 451 2550 525 2566
rect 451 2548 464 2550
rect 479 2548 513 2550
rect 116 2526 129 2528
rect 144 2526 178 2528
rect 116 2510 178 2526
rect 222 2521 238 2524
rect 300 2521 330 2532
rect 378 2528 424 2544
rect 451 2532 525 2548
rect 378 2526 412 2528
rect 377 2510 424 2526
rect 451 2510 464 2532
rect 479 2510 509 2532
rect 536 2510 537 2526
rect 552 2510 565 2670
rect 595 2566 608 2670
rect 653 2648 654 2658
rect 669 2648 682 2658
rect 653 2644 682 2648
rect 687 2644 717 2670
rect 735 2656 751 2658
rect 823 2656 876 2670
rect 824 2654 888 2656
rect 931 2654 946 2670
rect 995 2667 1025 2670
rect 995 2664 1031 2667
rect 961 2656 977 2658
rect 735 2644 750 2648
rect 653 2642 750 2644
rect 778 2642 946 2654
rect 962 2644 977 2648
rect 995 2645 1034 2664
rect 1053 2658 1060 2659
rect 1059 2651 1060 2658
rect 1043 2648 1044 2651
rect 1059 2648 1072 2651
rect 995 2644 1025 2645
rect 1034 2644 1040 2645
rect 1043 2644 1072 2648
rect 962 2643 1072 2644
rect 962 2642 1078 2643
rect 637 2634 688 2642
rect 637 2622 662 2634
rect 669 2622 688 2634
rect 719 2634 769 2642
rect 719 2626 735 2634
rect 742 2632 769 2634
rect 778 2632 999 2642
rect 742 2622 999 2632
rect 1028 2634 1078 2642
rect 1028 2625 1044 2634
rect 637 2614 688 2622
rect 735 2614 999 2622
rect 1025 2622 1044 2625
rect 1051 2622 1078 2634
rect 1025 2614 1078 2622
rect 653 2606 654 2614
rect 669 2606 682 2614
rect 653 2598 669 2606
rect 650 2591 669 2594
rect 650 2582 672 2591
rect 623 2572 672 2582
rect 623 2566 653 2572
rect 672 2567 677 2572
rect 595 2550 669 2566
rect 687 2558 717 2614
rect 752 2604 960 2614
rect 995 2610 1040 2614
rect 1043 2613 1044 2614
rect 1059 2613 1072 2614
rect 778 2574 967 2604
rect 793 2571 967 2574
rect 786 2568 967 2571
rect 595 2548 608 2550
rect 623 2548 657 2550
rect 595 2532 669 2548
rect 696 2544 709 2558
rect 724 2544 740 2560
rect 786 2555 797 2568
rect 579 2510 580 2526
rect 595 2510 608 2532
rect 623 2510 653 2532
rect 696 2528 758 2544
rect 786 2537 797 2553
rect 802 2548 812 2568
rect 822 2548 836 2568
rect 839 2555 848 2568
rect 864 2555 873 2568
rect 802 2537 836 2548
rect 839 2537 848 2553
rect 864 2537 873 2553
rect 880 2548 890 2568
rect 900 2548 914 2568
rect 915 2555 926 2568
rect 880 2537 914 2548
rect 915 2537 926 2553
rect 972 2544 988 2560
rect 995 2558 1025 2610
rect 1059 2606 1060 2613
rect 1044 2598 1060 2606
rect 1031 2566 1044 2585
rect 1059 2566 1089 2582
rect 1031 2550 1105 2566
rect 1031 2548 1044 2550
rect 1059 2548 1093 2550
rect 696 2526 709 2528
rect 724 2526 758 2528
rect 696 2510 758 2526
rect 802 2521 818 2524
rect 880 2521 910 2532
rect 958 2528 1004 2544
rect 1031 2532 1105 2548
rect 958 2526 992 2528
rect 957 2510 1004 2526
rect 1031 2510 1044 2532
rect 1059 2510 1089 2532
rect 1116 2510 1117 2526
rect 1132 2510 1145 2670
rect 1175 2566 1188 2670
rect 1233 2648 1234 2658
rect 1249 2648 1262 2658
rect 1233 2644 1262 2648
rect 1267 2644 1297 2670
rect 1315 2656 1331 2658
rect 1403 2656 1456 2670
rect 1404 2654 1468 2656
rect 1511 2654 1526 2670
rect 1575 2667 1605 2670
rect 1575 2664 1611 2667
rect 1541 2656 1557 2658
rect 1315 2644 1330 2648
rect 1233 2642 1330 2644
rect 1358 2642 1526 2654
rect 1542 2644 1557 2648
rect 1575 2645 1614 2664
rect 1633 2658 1640 2659
rect 1639 2651 1640 2658
rect 1623 2648 1624 2651
rect 1639 2648 1652 2651
rect 1575 2644 1605 2645
rect 1614 2644 1620 2645
rect 1623 2644 1652 2648
rect 1542 2643 1652 2644
rect 1542 2642 1658 2643
rect 1217 2634 1268 2642
rect 1217 2622 1242 2634
rect 1249 2622 1268 2634
rect 1299 2634 1349 2642
rect 1299 2626 1315 2634
rect 1322 2632 1349 2634
rect 1358 2632 1579 2642
rect 1322 2622 1579 2632
rect 1608 2634 1658 2642
rect 1608 2625 1624 2634
rect 1217 2614 1268 2622
rect 1315 2614 1579 2622
rect 1605 2622 1624 2625
rect 1631 2622 1658 2634
rect 1605 2614 1658 2622
rect 1233 2606 1234 2614
rect 1249 2606 1262 2614
rect 1233 2598 1249 2606
rect 1230 2591 1249 2594
rect 1230 2582 1252 2591
rect 1203 2572 1252 2582
rect 1203 2566 1233 2572
rect 1252 2567 1257 2572
rect 1175 2550 1249 2566
rect 1267 2558 1297 2614
rect 1332 2604 1540 2614
rect 1575 2610 1620 2614
rect 1623 2613 1624 2614
rect 1639 2613 1652 2614
rect 1358 2574 1547 2604
rect 1373 2571 1547 2574
rect 1366 2568 1547 2571
rect 1175 2548 1188 2550
rect 1203 2548 1237 2550
rect 1175 2532 1249 2548
rect 1276 2544 1289 2558
rect 1304 2544 1320 2560
rect 1366 2555 1377 2568
rect 1159 2510 1160 2526
rect 1175 2510 1188 2532
rect 1203 2510 1233 2532
rect 1276 2528 1338 2544
rect 1366 2537 1377 2553
rect 1382 2548 1392 2568
rect 1402 2548 1416 2568
rect 1419 2555 1428 2568
rect 1444 2555 1453 2568
rect 1382 2537 1416 2548
rect 1419 2537 1428 2553
rect 1444 2537 1453 2553
rect 1460 2548 1470 2568
rect 1480 2548 1494 2568
rect 1495 2555 1506 2568
rect 1460 2537 1494 2548
rect 1495 2537 1506 2553
rect 1552 2544 1568 2560
rect 1575 2558 1605 2610
rect 1639 2606 1640 2613
rect 1624 2598 1640 2606
rect 1611 2566 1624 2585
rect 1639 2566 1669 2582
rect 1611 2550 1685 2566
rect 1611 2548 1624 2550
rect 1639 2548 1673 2550
rect 1276 2526 1289 2528
rect 1304 2526 1338 2528
rect 1276 2510 1338 2526
rect 1382 2521 1398 2524
rect 1460 2521 1490 2532
rect 1538 2528 1584 2544
rect 1611 2532 1685 2548
rect 1538 2526 1572 2528
rect 1537 2510 1584 2526
rect 1611 2510 1624 2532
rect 1639 2510 1669 2532
rect 1696 2510 1697 2526
rect 1712 2510 1725 2670
rect 1755 2566 1768 2670
rect 1813 2648 1814 2658
rect 1829 2648 1842 2658
rect 1813 2644 1842 2648
rect 1847 2644 1877 2670
rect 1895 2656 1911 2658
rect 1983 2656 2036 2670
rect 1984 2654 2048 2656
rect 2091 2654 2106 2670
rect 2155 2667 2185 2670
rect 2155 2664 2191 2667
rect 2121 2656 2137 2658
rect 1895 2644 1910 2648
rect 1813 2642 1910 2644
rect 1938 2642 2106 2654
rect 2122 2644 2137 2648
rect 2155 2645 2194 2664
rect 2213 2658 2220 2659
rect 2219 2651 2220 2658
rect 2203 2648 2204 2651
rect 2219 2648 2232 2651
rect 2155 2644 2185 2645
rect 2194 2644 2200 2645
rect 2203 2644 2232 2648
rect 2122 2643 2232 2644
rect 2122 2642 2238 2643
rect 1797 2634 1848 2642
rect 1797 2622 1822 2634
rect 1829 2622 1848 2634
rect 1879 2634 1929 2642
rect 1879 2626 1895 2634
rect 1902 2632 1929 2634
rect 1938 2632 2159 2642
rect 1902 2622 2159 2632
rect 2188 2634 2238 2642
rect 2188 2625 2204 2634
rect 1797 2614 1848 2622
rect 1895 2614 2159 2622
rect 2185 2622 2204 2625
rect 2211 2622 2238 2634
rect 2185 2614 2238 2622
rect 1813 2606 1814 2614
rect 1829 2606 1842 2614
rect 1813 2598 1829 2606
rect 1810 2591 1829 2594
rect 1810 2582 1832 2591
rect 1783 2572 1832 2582
rect 1783 2566 1813 2572
rect 1832 2567 1837 2572
rect 1755 2550 1829 2566
rect 1847 2558 1877 2614
rect 1912 2604 2120 2614
rect 2155 2610 2200 2614
rect 2203 2613 2204 2614
rect 2219 2613 2232 2614
rect 1938 2574 2127 2604
rect 1953 2571 2127 2574
rect 1946 2568 2127 2571
rect 1755 2548 1768 2550
rect 1783 2548 1817 2550
rect 1755 2532 1829 2548
rect 1856 2544 1869 2558
rect 1884 2544 1900 2560
rect 1946 2555 1957 2568
rect 1739 2510 1740 2526
rect 1755 2510 1768 2532
rect 1783 2510 1813 2532
rect 1856 2528 1918 2544
rect 1946 2537 1957 2553
rect 1962 2548 1972 2568
rect 1982 2548 1996 2568
rect 1999 2555 2008 2568
rect 2024 2555 2033 2568
rect 1962 2537 1996 2548
rect 1999 2537 2008 2553
rect 2024 2537 2033 2553
rect 2040 2548 2050 2568
rect 2060 2548 2074 2568
rect 2075 2555 2086 2568
rect 2040 2537 2074 2548
rect 2075 2537 2086 2553
rect 2132 2544 2148 2560
rect 2155 2558 2185 2610
rect 2219 2606 2220 2613
rect 2204 2598 2220 2606
rect 2191 2566 2204 2585
rect 2219 2566 2249 2582
rect 2191 2550 2265 2566
rect 2191 2548 2204 2550
rect 2219 2548 2253 2550
rect 1856 2526 1869 2528
rect 1884 2526 1918 2528
rect 1856 2510 1918 2526
rect 1962 2521 1978 2524
rect 2040 2521 2070 2532
rect 2118 2528 2164 2544
rect 2191 2532 2265 2548
rect 2118 2526 2152 2528
rect 2117 2510 2164 2526
rect 2191 2510 2204 2532
rect 2219 2510 2249 2532
rect 2276 2510 2277 2526
rect 2292 2510 2305 2670
rect 2335 2566 2348 2670
rect 2393 2648 2394 2658
rect 2409 2648 2422 2658
rect 2393 2644 2422 2648
rect 2427 2644 2457 2670
rect 2475 2656 2491 2658
rect 2563 2656 2616 2670
rect 2564 2654 2628 2656
rect 2671 2654 2686 2670
rect 2735 2667 2765 2670
rect 2735 2664 2771 2667
rect 2701 2656 2717 2658
rect 2475 2644 2490 2648
rect 2393 2642 2490 2644
rect 2518 2642 2686 2654
rect 2702 2644 2717 2648
rect 2735 2645 2774 2664
rect 2793 2658 2800 2659
rect 2799 2651 2800 2658
rect 2783 2648 2784 2651
rect 2799 2648 2812 2651
rect 2735 2644 2765 2645
rect 2774 2644 2780 2645
rect 2783 2644 2812 2648
rect 2702 2643 2812 2644
rect 2702 2642 2818 2643
rect 2377 2634 2428 2642
rect 2377 2622 2402 2634
rect 2409 2622 2428 2634
rect 2459 2634 2509 2642
rect 2459 2626 2475 2634
rect 2482 2632 2509 2634
rect 2518 2632 2739 2642
rect 2482 2622 2739 2632
rect 2768 2634 2818 2642
rect 2768 2625 2784 2634
rect 2377 2614 2428 2622
rect 2475 2614 2739 2622
rect 2765 2622 2784 2625
rect 2791 2622 2818 2634
rect 2765 2614 2818 2622
rect 2393 2606 2394 2614
rect 2409 2606 2422 2614
rect 2393 2598 2409 2606
rect 2390 2591 2409 2594
rect 2390 2582 2412 2591
rect 2363 2572 2412 2582
rect 2363 2566 2393 2572
rect 2412 2567 2417 2572
rect 2335 2550 2409 2566
rect 2427 2558 2457 2614
rect 2492 2604 2700 2614
rect 2735 2610 2780 2614
rect 2783 2613 2784 2614
rect 2799 2613 2812 2614
rect 2518 2574 2707 2604
rect 2533 2571 2707 2574
rect 2526 2568 2707 2571
rect 2335 2548 2348 2550
rect 2363 2548 2397 2550
rect 2335 2532 2409 2548
rect 2436 2544 2449 2558
rect 2464 2544 2480 2560
rect 2526 2555 2537 2568
rect 2319 2510 2320 2526
rect 2335 2510 2348 2532
rect 2363 2510 2393 2532
rect 2436 2528 2498 2544
rect 2526 2537 2537 2553
rect 2542 2548 2552 2568
rect 2562 2548 2576 2568
rect 2579 2555 2588 2568
rect 2604 2555 2613 2568
rect 2542 2537 2576 2548
rect 2579 2537 2588 2553
rect 2604 2537 2613 2553
rect 2620 2548 2630 2568
rect 2640 2548 2654 2568
rect 2655 2555 2666 2568
rect 2620 2537 2654 2548
rect 2655 2537 2666 2553
rect 2712 2544 2728 2560
rect 2735 2558 2765 2610
rect 2799 2606 2800 2613
rect 2784 2598 2800 2606
rect 2771 2566 2784 2585
rect 2799 2566 2829 2582
rect 2771 2550 2845 2566
rect 2771 2548 2784 2550
rect 2799 2548 2833 2550
rect 2436 2526 2449 2528
rect 2464 2526 2498 2528
rect 2436 2510 2498 2526
rect 2542 2521 2558 2524
rect 2620 2521 2650 2532
rect 2698 2528 2744 2544
rect 2771 2532 2845 2548
rect 2698 2526 2732 2528
rect 2697 2510 2744 2526
rect 2771 2510 2784 2532
rect 2799 2510 2829 2532
rect 2856 2510 2857 2526
rect 2872 2510 2885 2670
rect 2915 2566 2928 2670
rect 2973 2648 2974 2658
rect 2989 2648 3002 2658
rect 2973 2644 3002 2648
rect 3007 2644 3037 2670
rect 3055 2656 3071 2658
rect 3143 2656 3196 2670
rect 3144 2654 3208 2656
rect 3251 2654 3266 2670
rect 3315 2667 3345 2670
rect 3315 2664 3351 2667
rect 3281 2656 3297 2658
rect 3055 2644 3070 2648
rect 2973 2642 3070 2644
rect 3098 2642 3266 2654
rect 3282 2644 3297 2648
rect 3315 2645 3354 2664
rect 3373 2658 3380 2659
rect 3379 2651 3380 2658
rect 3363 2648 3364 2651
rect 3379 2648 3392 2651
rect 3315 2644 3345 2645
rect 3354 2644 3360 2645
rect 3363 2644 3392 2648
rect 3282 2643 3392 2644
rect 3282 2642 3398 2643
rect 2957 2634 3008 2642
rect 2957 2622 2982 2634
rect 2989 2622 3008 2634
rect 3039 2634 3089 2642
rect 3039 2626 3055 2634
rect 3062 2632 3089 2634
rect 3098 2632 3319 2642
rect 3062 2622 3319 2632
rect 3348 2634 3398 2642
rect 3348 2625 3364 2634
rect 2957 2614 3008 2622
rect 3055 2614 3319 2622
rect 3345 2622 3364 2625
rect 3371 2622 3398 2634
rect 3345 2614 3398 2622
rect 2973 2606 2974 2614
rect 2989 2606 3002 2614
rect 2973 2598 2989 2606
rect 2970 2591 2989 2594
rect 2970 2582 2992 2591
rect 2943 2572 2992 2582
rect 2943 2566 2973 2572
rect 2992 2567 2997 2572
rect 2915 2550 2989 2566
rect 3007 2558 3037 2614
rect 3072 2604 3280 2614
rect 3315 2610 3360 2614
rect 3363 2613 3364 2614
rect 3379 2613 3392 2614
rect 3098 2574 3287 2604
rect 3113 2571 3287 2574
rect 3106 2568 3287 2571
rect 2915 2548 2928 2550
rect 2943 2548 2977 2550
rect 2915 2532 2989 2548
rect 3016 2544 3029 2558
rect 3044 2544 3060 2560
rect 3106 2555 3117 2568
rect 2899 2510 2900 2526
rect 2915 2510 2928 2532
rect 2943 2510 2973 2532
rect 3016 2528 3078 2544
rect 3106 2537 3117 2553
rect 3122 2548 3132 2568
rect 3142 2548 3156 2568
rect 3159 2555 3168 2568
rect 3184 2555 3193 2568
rect 3122 2537 3156 2548
rect 3159 2537 3168 2553
rect 3184 2537 3193 2553
rect 3200 2548 3210 2568
rect 3220 2548 3234 2568
rect 3235 2555 3246 2568
rect 3200 2537 3234 2548
rect 3235 2537 3246 2553
rect 3292 2544 3308 2560
rect 3315 2558 3345 2610
rect 3379 2606 3380 2613
rect 3364 2598 3380 2606
rect 3351 2566 3364 2585
rect 3379 2566 3409 2582
rect 3351 2550 3425 2566
rect 3351 2548 3364 2550
rect 3379 2548 3413 2550
rect 3016 2526 3029 2528
rect 3044 2526 3078 2528
rect 3016 2510 3078 2526
rect 3122 2521 3138 2524
rect 3200 2521 3230 2532
rect 3278 2528 3324 2544
rect 3351 2532 3425 2548
rect 3278 2526 3312 2528
rect 3277 2510 3324 2526
rect 3351 2510 3364 2532
rect 3379 2510 3409 2532
rect 3436 2510 3437 2526
rect 3452 2510 3465 2670
rect 3495 2566 3508 2670
rect 3553 2648 3554 2658
rect 3569 2648 3582 2658
rect 3553 2644 3582 2648
rect 3587 2644 3617 2670
rect 3635 2656 3651 2658
rect 3723 2656 3776 2670
rect 3724 2654 3788 2656
rect 3831 2654 3846 2670
rect 3895 2667 3925 2670
rect 3895 2664 3931 2667
rect 3861 2656 3877 2658
rect 3635 2644 3650 2648
rect 3553 2642 3650 2644
rect 3678 2642 3846 2654
rect 3862 2644 3877 2648
rect 3895 2645 3934 2664
rect 3953 2658 3960 2659
rect 3959 2651 3960 2658
rect 3943 2648 3944 2651
rect 3959 2648 3972 2651
rect 3895 2644 3925 2645
rect 3934 2644 3940 2645
rect 3943 2644 3972 2648
rect 3862 2643 3972 2644
rect 3862 2642 3978 2643
rect 3537 2634 3588 2642
rect 3537 2622 3562 2634
rect 3569 2622 3588 2634
rect 3619 2634 3669 2642
rect 3619 2626 3635 2634
rect 3642 2632 3669 2634
rect 3678 2632 3899 2642
rect 3642 2622 3899 2632
rect 3928 2634 3978 2642
rect 3928 2625 3944 2634
rect 3537 2614 3588 2622
rect 3635 2614 3899 2622
rect 3925 2622 3944 2625
rect 3951 2622 3978 2634
rect 3925 2614 3978 2622
rect 3553 2606 3554 2614
rect 3569 2606 3582 2614
rect 3553 2598 3569 2606
rect 3550 2591 3569 2594
rect 3550 2582 3572 2591
rect 3523 2572 3572 2582
rect 3523 2566 3553 2572
rect 3572 2567 3577 2572
rect 3495 2550 3569 2566
rect 3587 2558 3617 2614
rect 3652 2604 3860 2614
rect 3895 2610 3940 2614
rect 3943 2613 3944 2614
rect 3959 2613 3972 2614
rect 3678 2574 3867 2604
rect 3693 2571 3867 2574
rect 3686 2568 3867 2571
rect 3495 2548 3508 2550
rect 3523 2548 3557 2550
rect 3495 2532 3569 2548
rect 3596 2544 3609 2558
rect 3624 2544 3640 2560
rect 3686 2555 3697 2568
rect 3479 2510 3480 2526
rect 3495 2510 3508 2532
rect 3523 2510 3553 2532
rect 3596 2528 3658 2544
rect 3686 2537 3697 2553
rect 3702 2548 3712 2568
rect 3722 2548 3736 2568
rect 3739 2555 3748 2568
rect 3764 2555 3773 2568
rect 3702 2537 3736 2548
rect 3739 2537 3748 2553
rect 3764 2537 3773 2553
rect 3780 2548 3790 2568
rect 3800 2548 3814 2568
rect 3815 2555 3826 2568
rect 3780 2537 3814 2548
rect 3815 2537 3826 2553
rect 3872 2544 3888 2560
rect 3895 2558 3925 2610
rect 3959 2606 3960 2613
rect 3944 2598 3960 2606
rect 3931 2566 3944 2585
rect 3959 2566 3989 2582
rect 3931 2550 4005 2566
rect 3931 2548 3944 2550
rect 3959 2548 3993 2550
rect 3596 2526 3609 2528
rect 3624 2526 3658 2528
rect 3596 2510 3658 2526
rect 3702 2521 3718 2524
rect 3780 2521 3810 2532
rect 3858 2528 3904 2544
rect 3931 2532 4005 2548
rect 3858 2526 3892 2528
rect 3857 2510 3904 2526
rect 3931 2510 3944 2532
rect 3959 2510 3989 2532
rect 4016 2510 4017 2526
rect 4032 2510 4045 2670
rect 4075 2566 4088 2670
rect 4133 2648 4134 2658
rect 4149 2648 4162 2658
rect 4133 2644 4162 2648
rect 4167 2644 4197 2670
rect 4215 2656 4231 2658
rect 4303 2656 4356 2670
rect 4304 2654 4368 2656
rect 4411 2654 4426 2670
rect 4475 2667 4505 2670
rect 4475 2664 4511 2667
rect 4441 2656 4457 2658
rect 4215 2644 4230 2648
rect 4133 2642 4230 2644
rect 4258 2642 4426 2654
rect 4442 2644 4457 2648
rect 4475 2645 4514 2664
rect 4533 2658 4540 2659
rect 4539 2651 4540 2658
rect 4523 2648 4524 2651
rect 4539 2648 4552 2651
rect 4475 2644 4505 2645
rect 4514 2644 4520 2645
rect 4523 2644 4552 2648
rect 4442 2643 4552 2644
rect 4442 2642 4558 2643
rect 4117 2634 4168 2642
rect 4117 2622 4142 2634
rect 4149 2622 4168 2634
rect 4199 2634 4249 2642
rect 4199 2626 4215 2634
rect 4222 2632 4249 2634
rect 4258 2632 4479 2642
rect 4222 2622 4479 2632
rect 4508 2634 4558 2642
rect 4508 2625 4524 2634
rect 4117 2614 4168 2622
rect 4215 2614 4479 2622
rect 4505 2622 4524 2625
rect 4531 2622 4558 2634
rect 4505 2614 4558 2622
rect 4133 2606 4134 2614
rect 4149 2606 4162 2614
rect 4133 2598 4149 2606
rect 4130 2591 4149 2594
rect 4130 2582 4152 2591
rect 4103 2572 4152 2582
rect 4103 2566 4133 2572
rect 4152 2567 4157 2572
rect 4075 2550 4149 2566
rect 4167 2558 4197 2614
rect 4232 2604 4440 2614
rect 4475 2610 4520 2614
rect 4523 2613 4524 2614
rect 4539 2613 4552 2614
rect 4258 2574 4447 2604
rect 4273 2571 4447 2574
rect 4266 2568 4447 2571
rect 4075 2548 4088 2550
rect 4103 2548 4137 2550
rect 4075 2532 4149 2548
rect 4176 2544 4189 2558
rect 4204 2544 4220 2560
rect 4266 2555 4277 2568
rect 4059 2510 4060 2526
rect 4075 2510 4088 2532
rect 4103 2510 4133 2532
rect 4176 2528 4238 2544
rect 4266 2537 4277 2553
rect 4282 2548 4292 2568
rect 4302 2548 4316 2568
rect 4319 2555 4328 2568
rect 4344 2555 4353 2568
rect 4282 2537 4316 2548
rect 4319 2537 4328 2553
rect 4344 2537 4353 2553
rect 4360 2548 4370 2568
rect 4380 2548 4394 2568
rect 4395 2555 4406 2568
rect 4360 2537 4394 2548
rect 4395 2537 4406 2553
rect 4452 2544 4468 2560
rect 4475 2558 4505 2610
rect 4539 2606 4540 2613
rect 4524 2598 4540 2606
rect 4511 2566 4524 2585
rect 4539 2566 4569 2582
rect 4511 2550 4585 2566
rect 4511 2548 4524 2550
rect 4539 2548 4573 2550
rect 4176 2526 4189 2528
rect 4204 2526 4238 2528
rect 4176 2510 4238 2526
rect 4282 2521 4298 2524
rect 4360 2521 4390 2532
rect 4438 2528 4484 2544
rect 4511 2532 4585 2548
rect 4438 2526 4472 2528
rect 4437 2510 4484 2526
rect 4511 2510 4524 2532
rect 4539 2510 4569 2532
rect 4596 2510 4597 2526
rect 4612 2510 4625 2670
rect -7 2502 34 2510
rect -7 2476 8 2502
rect 15 2476 34 2502
rect 98 2498 160 2510
rect 172 2498 247 2510
rect 305 2498 380 2510
rect 392 2498 423 2510
rect 429 2498 464 2510
rect 98 2496 260 2498
rect -7 2468 34 2476
rect 116 2472 129 2496
rect 144 2494 159 2496
rect -1 2458 0 2468
rect 15 2458 28 2468
rect 43 2458 73 2472
rect 116 2458 159 2472
rect 183 2469 190 2476
rect 193 2472 260 2496
rect 292 2496 464 2498
rect 262 2474 290 2478
rect 292 2474 372 2496
rect 393 2494 408 2496
rect 262 2472 372 2474
rect 193 2468 372 2472
rect 166 2458 196 2468
rect 198 2458 351 2468
rect 359 2458 389 2468
rect 393 2458 423 2472
rect 451 2458 464 2496
rect 536 2502 571 2510
rect 536 2476 537 2502
rect 544 2476 571 2502
rect 479 2458 509 2472
rect 536 2468 571 2476
rect 573 2502 614 2510
rect 573 2476 588 2502
rect 595 2476 614 2502
rect 678 2498 740 2510
rect 752 2498 827 2510
rect 885 2498 960 2510
rect 972 2498 1003 2510
rect 1009 2498 1044 2510
rect 678 2496 840 2498
rect 573 2468 614 2476
rect 696 2472 709 2496
rect 724 2494 739 2496
rect 536 2458 537 2468
rect 552 2458 565 2468
rect 579 2458 580 2468
rect 595 2458 608 2468
rect 623 2458 653 2472
rect 696 2458 739 2472
rect 763 2469 770 2476
rect 773 2472 840 2496
rect 872 2496 1044 2498
rect 842 2474 870 2478
rect 872 2474 952 2496
rect 973 2494 988 2496
rect 842 2472 952 2474
rect 773 2468 952 2472
rect 746 2458 776 2468
rect 778 2458 931 2468
rect 939 2458 969 2468
rect 973 2458 1003 2472
rect 1031 2458 1044 2496
rect 1116 2502 1151 2510
rect 1116 2476 1117 2502
rect 1124 2476 1151 2502
rect 1059 2458 1089 2472
rect 1116 2468 1151 2476
rect 1153 2502 1194 2510
rect 1153 2476 1168 2502
rect 1175 2476 1194 2502
rect 1258 2498 1320 2510
rect 1332 2498 1407 2510
rect 1465 2498 1540 2510
rect 1552 2498 1583 2510
rect 1589 2498 1624 2510
rect 1258 2496 1420 2498
rect 1153 2468 1194 2476
rect 1276 2472 1289 2496
rect 1304 2494 1319 2496
rect 1116 2458 1117 2468
rect 1132 2458 1145 2468
rect 1159 2458 1160 2468
rect 1175 2458 1188 2468
rect 1203 2458 1233 2472
rect 1276 2458 1319 2472
rect 1343 2469 1350 2476
rect 1353 2472 1420 2496
rect 1452 2496 1624 2498
rect 1422 2474 1450 2478
rect 1452 2474 1532 2496
rect 1553 2494 1568 2496
rect 1422 2472 1532 2474
rect 1353 2468 1532 2472
rect 1326 2458 1356 2468
rect 1358 2458 1511 2468
rect 1519 2458 1549 2468
rect 1553 2458 1583 2472
rect 1611 2458 1624 2496
rect 1696 2502 1731 2510
rect 1696 2476 1697 2502
rect 1704 2476 1731 2502
rect 1639 2458 1669 2472
rect 1696 2468 1731 2476
rect 1733 2502 1774 2510
rect 1733 2476 1748 2502
rect 1755 2476 1774 2502
rect 1838 2498 1900 2510
rect 1912 2498 1987 2510
rect 2045 2498 2120 2510
rect 2132 2498 2163 2510
rect 2169 2498 2204 2510
rect 1838 2496 2000 2498
rect 1733 2468 1774 2476
rect 1856 2472 1869 2496
rect 1884 2494 1899 2496
rect 1696 2458 1697 2468
rect 1712 2458 1725 2468
rect 1739 2458 1740 2468
rect 1755 2458 1768 2468
rect 1783 2458 1813 2472
rect 1856 2458 1899 2472
rect 1923 2469 1930 2476
rect 1933 2472 2000 2496
rect 2032 2496 2204 2498
rect 2002 2474 2030 2478
rect 2032 2474 2112 2496
rect 2133 2494 2148 2496
rect 2002 2472 2112 2474
rect 1933 2468 2112 2472
rect 1906 2458 1936 2468
rect 1938 2458 2091 2468
rect 2099 2458 2129 2468
rect 2133 2458 2163 2472
rect 2191 2458 2204 2496
rect 2276 2502 2311 2510
rect 2276 2476 2277 2502
rect 2284 2476 2311 2502
rect 2219 2458 2249 2472
rect 2276 2468 2311 2476
rect 2313 2502 2354 2510
rect 2313 2476 2328 2502
rect 2335 2476 2354 2502
rect 2418 2498 2480 2510
rect 2492 2498 2567 2510
rect 2625 2498 2700 2510
rect 2712 2498 2743 2510
rect 2749 2498 2784 2510
rect 2418 2496 2580 2498
rect 2313 2468 2354 2476
rect 2436 2472 2449 2496
rect 2464 2494 2479 2496
rect 2276 2458 2277 2468
rect 2292 2458 2305 2468
rect 2319 2458 2320 2468
rect 2335 2458 2348 2468
rect 2363 2458 2393 2472
rect 2436 2458 2479 2472
rect 2503 2469 2510 2476
rect 2513 2472 2580 2496
rect 2612 2496 2784 2498
rect 2582 2474 2610 2478
rect 2612 2474 2692 2496
rect 2713 2494 2728 2496
rect 2582 2472 2692 2474
rect 2513 2468 2692 2472
rect 2486 2458 2516 2468
rect 2518 2458 2671 2468
rect 2679 2458 2709 2468
rect 2713 2458 2743 2472
rect 2771 2458 2784 2496
rect 2856 2502 2891 2510
rect 2856 2476 2857 2502
rect 2864 2476 2891 2502
rect 2799 2458 2829 2472
rect 2856 2468 2891 2476
rect 2893 2502 2934 2510
rect 2893 2476 2908 2502
rect 2915 2476 2934 2502
rect 2998 2498 3060 2510
rect 3072 2498 3147 2510
rect 3205 2498 3280 2510
rect 3292 2498 3323 2510
rect 3329 2498 3364 2510
rect 2998 2496 3160 2498
rect 2893 2468 2934 2476
rect 3016 2472 3029 2496
rect 3044 2494 3059 2496
rect 2856 2458 2857 2468
rect 2872 2458 2885 2468
rect 2899 2458 2900 2468
rect 2915 2458 2928 2468
rect 2943 2458 2973 2472
rect 3016 2458 3059 2472
rect 3083 2469 3090 2476
rect 3093 2472 3160 2496
rect 3192 2496 3364 2498
rect 3162 2474 3190 2478
rect 3192 2474 3272 2496
rect 3293 2494 3308 2496
rect 3162 2472 3272 2474
rect 3093 2468 3272 2472
rect 3066 2458 3096 2468
rect 3098 2458 3251 2468
rect 3259 2458 3289 2468
rect 3293 2458 3323 2472
rect 3351 2458 3364 2496
rect 3436 2502 3471 2510
rect 3436 2476 3437 2502
rect 3444 2476 3471 2502
rect 3379 2458 3409 2472
rect 3436 2468 3471 2476
rect 3473 2502 3514 2510
rect 3473 2476 3488 2502
rect 3495 2476 3514 2502
rect 3578 2498 3640 2510
rect 3652 2498 3727 2510
rect 3785 2498 3860 2510
rect 3872 2498 3903 2510
rect 3909 2498 3944 2510
rect 3578 2496 3740 2498
rect 3473 2468 3514 2476
rect 3596 2472 3609 2496
rect 3624 2494 3639 2496
rect 3436 2458 3437 2468
rect 3452 2458 3465 2468
rect 3479 2458 3480 2468
rect 3495 2458 3508 2468
rect 3523 2458 3553 2472
rect 3596 2458 3639 2472
rect 3663 2469 3670 2476
rect 3673 2472 3740 2496
rect 3772 2496 3944 2498
rect 3742 2474 3770 2478
rect 3772 2474 3852 2496
rect 3873 2494 3888 2496
rect 3742 2472 3852 2474
rect 3673 2468 3852 2472
rect 3646 2458 3676 2468
rect 3678 2458 3831 2468
rect 3839 2458 3869 2468
rect 3873 2458 3903 2472
rect 3931 2458 3944 2496
rect 4016 2502 4051 2510
rect 4016 2476 4017 2502
rect 4024 2476 4051 2502
rect 3959 2458 3989 2472
rect 4016 2468 4051 2476
rect 4053 2502 4094 2510
rect 4053 2476 4068 2502
rect 4075 2476 4094 2502
rect 4158 2498 4220 2510
rect 4232 2498 4307 2510
rect 4365 2498 4440 2510
rect 4452 2498 4483 2510
rect 4489 2498 4524 2510
rect 4158 2496 4320 2498
rect 4053 2468 4094 2476
rect 4176 2472 4189 2496
rect 4204 2494 4219 2496
rect 4016 2458 4017 2468
rect 4032 2458 4045 2468
rect 4059 2458 4060 2468
rect 4075 2458 4088 2468
rect 4103 2458 4133 2472
rect 4176 2458 4219 2472
rect 4243 2469 4250 2476
rect 4253 2472 4320 2496
rect 4352 2496 4524 2498
rect 4322 2474 4350 2478
rect 4352 2474 4432 2496
rect 4453 2494 4468 2496
rect 4322 2472 4432 2474
rect 4253 2468 4432 2472
rect 4226 2458 4256 2468
rect 4258 2458 4411 2468
rect 4419 2458 4449 2468
rect 4453 2458 4483 2472
rect 4511 2458 4524 2496
rect 4596 2502 4631 2510
rect 4596 2476 4597 2502
rect 4604 2476 4631 2502
rect 4539 2458 4569 2472
rect 4596 2468 4631 2476
rect 4596 2458 4597 2468
rect 4612 2458 4625 2468
rect -1 2452 4625 2458
rect 0 2444 4625 2452
rect 15 2414 28 2444
rect 43 2426 73 2444
rect 116 2430 130 2444
rect 166 2430 386 2444
rect 117 2428 130 2430
rect 83 2416 98 2428
rect 80 2414 102 2416
rect 107 2414 137 2428
rect 198 2426 351 2430
rect 180 2414 372 2426
rect 415 2414 445 2428
rect 451 2414 464 2444
rect 479 2426 509 2444
rect 552 2414 565 2444
rect 595 2414 608 2444
rect 623 2426 653 2444
rect 696 2430 710 2444
rect 746 2430 966 2444
rect 697 2428 710 2430
rect 663 2416 678 2428
rect 660 2414 682 2416
rect 687 2414 717 2428
rect 778 2426 931 2430
rect 760 2414 952 2426
rect 995 2414 1025 2428
rect 1031 2414 1044 2444
rect 1059 2426 1089 2444
rect 1132 2414 1145 2444
rect 1175 2414 1188 2444
rect 1203 2426 1233 2444
rect 1276 2430 1290 2444
rect 1326 2430 1546 2444
rect 1277 2428 1290 2430
rect 1243 2416 1258 2428
rect 1240 2414 1262 2416
rect 1267 2414 1297 2428
rect 1358 2426 1511 2430
rect 1340 2414 1532 2426
rect 1575 2414 1605 2428
rect 1611 2414 1624 2444
rect 1639 2426 1669 2444
rect 1712 2414 1725 2444
rect 1755 2414 1768 2444
rect 1783 2426 1813 2444
rect 1856 2430 1870 2444
rect 1906 2430 2126 2444
rect 1857 2428 1870 2430
rect 1823 2416 1838 2428
rect 1820 2414 1842 2416
rect 1847 2414 1877 2428
rect 1938 2426 2091 2430
rect 1920 2414 2112 2426
rect 2155 2414 2185 2428
rect 2191 2414 2204 2444
rect 2219 2426 2249 2444
rect 2292 2414 2305 2444
rect 2335 2414 2348 2444
rect 2363 2426 2393 2444
rect 2436 2430 2450 2444
rect 2486 2430 2706 2444
rect 2437 2428 2450 2430
rect 2403 2416 2418 2428
rect 2400 2414 2422 2416
rect 2427 2414 2457 2428
rect 2518 2426 2671 2430
rect 2500 2414 2692 2426
rect 2735 2414 2765 2428
rect 2771 2414 2784 2444
rect 2799 2426 2829 2444
rect 2872 2414 2885 2444
rect 2915 2414 2928 2444
rect 2943 2426 2973 2444
rect 3016 2430 3030 2444
rect 3066 2430 3286 2444
rect 3017 2428 3030 2430
rect 2983 2416 2998 2428
rect 2980 2414 3002 2416
rect 3007 2414 3037 2428
rect 3098 2426 3251 2430
rect 3080 2414 3272 2426
rect 3315 2414 3345 2428
rect 3351 2414 3364 2444
rect 3379 2426 3409 2444
rect 3452 2414 3465 2444
rect 3495 2414 3508 2444
rect 3523 2426 3553 2444
rect 3596 2430 3610 2444
rect 3646 2430 3866 2444
rect 3597 2428 3610 2430
rect 3563 2416 3578 2428
rect 3560 2414 3582 2416
rect 3587 2414 3617 2428
rect 3678 2426 3831 2430
rect 3660 2414 3852 2426
rect 3895 2414 3925 2428
rect 3931 2414 3944 2444
rect 3959 2426 3989 2444
rect 4032 2414 4045 2444
rect 4075 2414 4088 2444
rect 4103 2426 4133 2444
rect 4176 2430 4190 2444
rect 4226 2430 4446 2444
rect 4177 2428 4190 2430
rect 4143 2416 4158 2428
rect 4140 2414 4162 2416
rect 4167 2414 4197 2428
rect 4258 2426 4411 2430
rect 4240 2414 4432 2426
rect 4475 2414 4505 2428
rect 4511 2414 4524 2444
rect 4539 2426 4569 2444
rect 4612 2414 4625 2444
rect 0 2400 4625 2414
rect 15 2296 28 2400
rect 73 2378 74 2388
rect 89 2378 102 2388
rect 73 2374 102 2378
rect 107 2374 137 2400
rect 155 2386 171 2388
rect 243 2386 296 2400
rect 244 2384 308 2386
rect 351 2384 366 2400
rect 415 2397 445 2400
rect 415 2394 451 2397
rect 381 2386 397 2388
rect 155 2374 170 2378
rect 73 2372 170 2374
rect 198 2372 366 2384
rect 382 2374 397 2378
rect 415 2375 454 2394
rect 473 2388 480 2389
rect 479 2381 480 2388
rect 463 2378 464 2381
rect 479 2378 492 2381
rect 415 2374 445 2375
rect 454 2374 460 2375
rect 463 2374 492 2378
rect 382 2373 492 2374
rect 382 2372 498 2373
rect 57 2364 108 2372
rect 57 2352 82 2364
rect 89 2352 108 2364
rect 139 2364 189 2372
rect 139 2356 155 2364
rect 162 2362 189 2364
rect 198 2362 419 2372
rect 162 2352 419 2362
rect 448 2364 498 2372
rect 448 2355 464 2364
rect 57 2344 108 2352
rect 155 2344 419 2352
rect 445 2352 464 2355
rect 471 2352 498 2364
rect 445 2344 498 2352
rect 73 2336 74 2344
rect 89 2336 102 2344
rect 73 2328 89 2336
rect 70 2321 89 2324
rect 70 2312 92 2321
rect 43 2302 92 2312
rect 43 2296 73 2302
rect 92 2297 97 2302
rect 15 2280 89 2296
rect 107 2288 137 2344
rect 172 2334 380 2344
rect 415 2340 460 2344
rect 463 2343 464 2344
rect 479 2343 492 2344
rect 198 2304 387 2334
rect 213 2301 387 2304
rect 206 2298 387 2301
rect 15 2278 28 2280
rect 43 2278 77 2280
rect 15 2262 89 2278
rect 116 2274 129 2288
rect 144 2274 160 2290
rect 206 2285 217 2298
rect -1 2240 0 2256
rect 15 2240 28 2262
rect 43 2240 73 2262
rect 116 2258 178 2274
rect 206 2267 217 2283
rect 222 2278 232 2298
rect 242 2278 256 2298
rect 259 2285 268 2298
rect 284 2285 293 2298
rect 222 2267 256 2278
rect 259 2267 268 2283
rect 284 2267 293 2283
rect 300 2278 310 2298
rect 320 2278 334 2298
rect 335 2285 346 2298
rect 300 2267 334 2278
rect 335 2267 346 2283
rect 392 2274 408 2290
rect 415 2288 445 2340
rect 479 2336 480 2343
rect 464 2328 480 2336
rect 451 2296 464 2315
rect 479 2296 509 2312
rect 451 2280 525 2296
rect 451 2278 464 2280
rect 479 2278 513 2280
rect 116 2256 129 2258
rect 144 2256 178 2258
rect 116 2240 178 2256
rect 222 2251 238 2254
rect 300 2251 330 2262
rect 378 2258 424 2274
rect 451 2262 525 2278
rect 378 2256 412 2258
rect 377 2240 424 2256
rect 451 2240 464 2262
rect 479 2240 509 2262
rect 536 2240 537 2256
rect 552 2240 565 2400
rect 595 2296 608 2400
rect 653 2378 654 2388
rect 669 2378 682 2388
rect 653 2374 682 2378
rect 687 2374 717 2400
rect 735 2386 751 2388
rect 823 2386 876 2400
rect 824 2384 888 2386
rect 931 2384 946 2400
rect 995 2397 1025 2400
rect 995 2394 1031 2397
rect 961 2386 977 2388
rect 735 2374 750 2378
rect 653 2372 750 2374
rect 778 2372 946 2384
rect 962 2374 977 2378
rect 995 2375 1034 2394
rect 1053 2388 1060 2389
rect 1059 2381 1060 2388
rect 1043 2378 1044 2381
rect 1059 2378 1072 2381
rect 995 2374 1025 2375
rect 1034 2374 1040 2375
rect 1043 2374 1072 2378
rect 962 2373 1072 2374
rect 962 2372 1078 2373
rect 637 2364 688 2372
rect 637 2352 662 2364
rect 669 2352 688 2364
rect 719 2364 769 2372
rect 719 2356 735 2364
rect 742 2362 769 2364
rect 778 2362 999 2372
rect 742 2352 999 2362
rect 1028 2364 1078 2372
rect 1028 2355 1044 2364
rect 637 2344 688 2352
rect 735 2344 999 2352
rect 1025 2352 1044 2355
rect 1051 2352 1078 2364
rect 1025 2344 1078 2352
rect 653 2336 654 2344
rect 669 2336 682 2344
rect 653 2328 669 2336
rect 650 2321 669 2324
rect 650 2312 672 2321
rect 623 2302 672 2312
rect 623 2296 653 2302
rect 672 2297 677 2302
rect 595 2280 669 2296
rect 687 2288 717 2344
rect 752 2334 960 2344
rect 995 2340 1040 2344
rect 1043 2343 1044 2344
rect 1059 2343 1072 2344
rect 778 2304 967 2334
rect 793 2301 967 2304
rect 786 2298 967 2301
rect 595 2278 608 2280
rect 623 2278 657 2280
rect 595 2262 669 2278
rect 696 2274 709 2288
rect 724 2274 740 2290
rect 786 2285 797 2298
rect 579 2240 580 2256
rect 595 2240 608 2262
rect 623 2240 653 2262
rect 696 2258 758 2274
rect 786 2267 797 2283
rect 802 2278 812 2298
rect 822 2278 836 2298
rect 839 2285 848 2298
rect 864 2285 873 2298
rect 802 2267 836 2278
rect 839 2267 848 2283
rect 864 2267 873 2283
rect 880 2278 890 2298
rect 900 2278 914 2298
rect 915 2285 926 2298
rect 880 2267 914 2278
rect 915 2267 926 2283
rect 972 2274 988 2290
rect 995 2288 1025 2340
rect 1059 2336 1060 2343
rect 1044 2328 1060 2336
rect 1031 2296 1044 2315
rect 1059 2296 1089 2312
rect 1031 2280 1105 2296
rect 1031 2278 1044 2280
rect 1059 2278 1093 2280
rect 696 2256 709 2258
rect 724 2256 758 2258
rect 696 2240 758 2256
rect 802 2251 818 2254
rect 880 2251 910 2262
rect 958 2258 1004 2274
rect 1031 2262 1105 2278
rect 958 2256 992 2258
rect 957 2240 1004 2256
rect 1031 2240 1044 2262
rect 1059 2240 1089 2262
rect 1116 2240 1117 2256
rect 1132 2240 1145 2400
rect 1175 2296 1188 2400
rect 1233 2378 1234 2388
rect 1249 2378 1262 2388
rect 1233 2374 1262 2378
rect 1267 2374 1297 2400
rect 1315 2386 1331 2388
rect 1403 2386 1456 2400
rect 1404 2384 1468 2386
rect 1511 2384 1526 2400
rect 1575 2397 1605 2400
rect 1575 2394 1611 2397
rect 1541 2386 1557 2388
rect 1315 2374 1330 2378
rect 1233 2372 1330 2374
rect 1358 2372 1526 2384
rect 1542 2374 1557 2378
rect 1575 2375 1614 2394
rect 1633 2388 1640 2389
rect 1639 2381 1640 2388
rect 1623 2378 1624 2381
rect 1639 2378 1652 2381
rect 1575 2374 1605 2375
rect 1614 2374 1620 2375
rect 1623 2374 1652 2378
rect 1542 2373 1652 2374
rect 1542 2372 1658 2373
rect 1217 2364 1268 2372
rect 1217 2352 1242 2364
rect 1249 2352 1268 2364
rect 1299 2364 1349 2372
rect 1299 2356 1315 2364
rect 1322 2362 1349 2364
rect 1358 2362 1579 2372
rect 1322 2352 1579 2362
rect 1608 2364 1658 2372
rect 1608 2355 1624 2364
rect 1217 2344 1268 2352
rect 1315 2344 1579 2352
rect 1605 2352 1624 2355
rect 1631 2352 1658 2364
rect 1605 2344 1658 2352
rect 1233 2336 1234 2344
rect 1249 2336 1262 2344
rect 1233 2328 1249 2336
rect 1230 2321 1249 2324
rect 1230 2312 1252 2321
rect 1203 2302 1252 2312
rect 1203 2296 1233 2302
rect 1252 2297 1257 2302
rect 1175 2280 1249 2296
rect 1267 2288 1297 2344
rect 1332 2334 1540 2344
rect 1575 2340 1620 2344
rect 1623 2343 1624 2344
rect 1639 2343 1652 2344
rect 1358 2304 1547 2334
rect 1373 2301 1547 2304
rect 1366 2298 1547 2301
rect 1175 2278 1188 2280
rect 1203 2278 1237 2280
rect 1175 2262 1249 2278
rect 1276 2274 1289 2288
rect 1304 2274 1320 2290
rect 1366 2285 1377 2298
rect 1159 2240 1160 2256
rect 1175 2240 1188 2262
rect 1203 2240 1233 2262
rect 1276 2258 1338 2274
rect 1366 2267 1377 2283
rect 1382 2278 1392 2298
rect 1402 2278 1416 2298
rect 1419 2285 1428 2298
rect 1444 2285 1453 2298
rect 1382 2267 1416 2278
rect 1419 2267 1428 2283
rect 1444 2267 1453 2283
rect 1460 2278 1470 2298
rect 1480 2278 1494 2298
rect 1495 2285 1506 2298
rect 1460 2267 1494 2278
rect 1495 2267 1506 2283
rect 1552 2274 1568 2290
rect 1575 2288 1605 2340
rect 1639 2336 1640 2343
rect 1624 2328 1640 2336
rect 1611 2296 1624 2315
rect 1639 2296 1669 2312
rect 1611 2280 1685 2296
rect 1611 2278 1624 2280
rect 1639 2278 1673 2280
rect 1276 2256 1289 2258
rect 1304 2256 1338 2258
rect 1276 2240 1338 2256
rect 1382 2251 1398 2254
rect 1460 2251 1490 2262
rect 1538 2258 1584 2274
rect 1611 2262 1685 2278
rect 1538 2256 1572 2258
rect 1537 2240 1584 2256
rect 1611 2240 1624 2262
rect 1639 2240 1669 2262
rect 1696 2240 1697 2256
rect 1712 2240 1725 2400
rect 1755 2296 1768 2400
rect 1813 2378 1814 2388
rect 1829 2378 1842 2388
rect 1813 2374 1842 2378
rect 1847 2374 1877 2400
rect 1895 2386 1911 2388
rect 1983 2386 2036 2400
rect 1984 2384 2048 2386
rect 2091 2384 2106 2400
rect 2155 2397 2185 2400
rect 2155 2394 2191 2397
rect 2121 2386 2137 2388
rect 1895 2374 1910 2378
rect 1813 2372 1910 2374
rect 1938 2372 2106 2384
rect 2122 2374 2137 2378
rect 2155 2375 2194 2394
rect 2213 2388 2220 2389
rect 2219 2381 2220 2388
rect 2203 2378 2204 2381
rect 2219 2378 2232 2381
rect 2155 2374 2185 2375
rect 2194 2374 2200 2375
rect 2203 2374 2232 2378
rect 2122 2373 2232 2374
rect 2122 2372 2238 2373
rect 1797 2364 1848 2372
rect 1797 2352 1822 2364
rect 1829 2352 1848 2364
rect 1879 2364 1929 2372
rect 1879 2356 1895 2364
rect 1902 2362 1929 2364
rect 1938 2362 2159 2372
rect 1902 2352 2159 2362
rect 2188 2364 2238 2372
rect 2188 2355 2204 2364
rect 1797 2344 1848 2352
rect 1895 2344 2159 2352
rect 2185 2352 2204 2355
rect 2211 2352 2238 2364
rect 2185 2344 2238 2352
rect 1813 2336 1814 2344
rect 1829 2336 1842 2344
rect 1813 2328 1829 2336
rect 1810 2321 1829 2324
rect 1810 2312 1832 2321
rect 1783 2302 1832 2312
rect 1783 2296 1813 2302
rect 1832 2297 1837 2302
rect 1755 2280 1829 2296
rect 1847 2288 1877 2344
rect 1912 2334 2120 2344
rect 2155 2340 2200 2344
rect 2203 2343 2204 2344
rect 2219 2343 2232 2344
rect 1938 2304 2127 2334
rect 1953 2301 2127 2304
rect 1946 2298 2127 2301
rect 1755 2278 1768 2280
rect 1783 2278 1817 2280
rect 1755 2262 1829 2278
rect 1856 2274 1869 2288
rect 1884 2274 1900 2290
rect 1946 2285 1957 2298
rect 1739 2240 1740 2256
rect 1755 2240 1768 2262
rect 1783 2240 1813 2262
rect 1856 2258 1918 2274
rect 1946 2267 1957 2283
rect 1962 2278 1972 2298
rect 1982 2278 1996 2298
rect 1999 2285 2008 2298
rect 2024 2285 2033 2298
rect 1962 2267 1996 2278
rect 1999 2267 2008 2283
rect 2024 2267 2033 2283
rect 2040 2278 2050 2298
rect 2060 2278 2074 2298
rect 2075 2285 2086 2298
rect 2040 2267 2074 2278
rect 2075 2267 2086 2283
rect 2132 2274 2148 2290
rect 2155 2288 2185 2340
rect 2219 2336 2220 2343
rect 2204 2328 2220 2336
rect 2191 2296 2204 2315
rect 2219 2296 2249 2312
rect 2191 2280 2265 2296
rect 2191 2278 2204 2280
rect 2219 2278 2253 2280
rect 1856 2256 1869 2258
rect 1884 2256 1918 2258
rect 1856 2240 1918 2256
rect 1962 2251 1978 2254
rect 2040 2251 2070 2262
rect 2118 2258 2164 2274
rect 2191 2262 2265 2278
rect 2118 2256 2152 2258
rect 2117 2240 2164 2256
rect 2191 2240 2204 2262
rect 2219 2240 2249 2262
rect 2276 2240 2277 2256
rect 2292 2240 2305 2400
rect 2335 2296 2348 2400
rect 2393 2378 2394 2388
rect 2409 2378 2422 2388
rect 2393 2374 2422 2378
rect 2427 2374 2457 2400
rect 2475 2386 2491 2388
rect 2563 2386 2616 2400
rect 2564 2384 2628 2386
rect 2671 2384 2686 2400
rect 2735 2397 2765 2400
rect 2735 2394 2771 2397
rect 2701 2386 2717 2388
rect 2475 2374 2490 2378
rect 2393 2372 2490 2374
rect 2518 2372 2686 2384
rect 2702 2374 2717 2378
rect 2735 2375 2774 2394
rect 2793 2388 2800 2389
rect 2799 2381 2800 2388
rect 2783 2378 2784 2381
rect 2799 2378 2812 2381
rect 2735 2374 2765 2375
rect 2774 2374 2780 2375
rect 2783 2374 2812 2378
rect 2702 2373 2812 2374
rect 2702 2372 2818 2373
rect 2377 2364 2428 2372
rect 2377 2352 2402 2364
rect 2409 2352 2428 2364
rect 2459 2364 2509 2372
rect 2459 2356 2475 2364
rect 2482 2362 2509 2364
rect 2518 2362 2739 2372
rect 2482 2352 2739 2362
rect 2768 2364 2818 2372
rect 2768 2355 2784 2364
rect 2377 2344 2428 2352
rect 2475 2344 2739 2352
rect 2765 2352 2784 2355
rect 2791 2352 2818 2364
rect 2765 2344 2818 2352
rect 2393 2336 2394 2344
rect 2409 2336 2422 2344
rect 2393 2328 2409 2336
rect 2390 2321 2409 2324
rect 2390 2312 2412 2321
rect 2363 2302 2412 2312
rect 2363 2296 2393 2302
rect 2412 2297 2417 2302
rect 2335 2280 2409 2296
rect 2427 2288 2457 2344
rect 2492 2334 2700 2344
rect 2735 2340 2780 2344
rect 2783 2343 2784 2344
rect 2799 2343 2812 2344
rect 2518 2304 2707 2334
rect 2533 2301 2707 2304
rect 2526 2298 2707 2301
rect 2335 2278 2348 2280
rect 2363 2278 2397 2280
rect 2335 2262 2409 2278
rect 2436 2274 2449 2288
rect 2464 2274 2480 2290
rect 2526 2285 2537 2298
rect 2319 2240 2320 2256
rect 2335 2240 2348 2262
rect 2363 2240 2393 2262
rect 2436 2258 2498 2274
rect 2526 2267 2537 2283
rect 2542 2278 2552 2298
rect 2562 2278 2576 2298
rect 2579 2285 2588 2298
rect 2604 2285 2613 2298
rect 2542 2267 2576 2278
rect 2579 2267 2588 2283
rect 2604 2267 2613 2283
rect 2620 2278 2630 2298
rect 2640 2278 2654 2298
rect 2655 2285 2666 2298
rect 2620 2267 2654 2278
rect 2655 2267 2666 2283
rect 2712 2274 2728 2290
rect 2735 2288 2765 2340
rect 2799 2336 2800 2343
rect 2784 2328 2800 2336
rect 2771 2296 2784 2315
rect 2799 2296 2829 2312
rect 2771 2280 2845 2296
rect 2771 2278 2784 2280
rect 2799 2278 2833 2280
rect 2436 2256 2449 2258
rect 2464 2256 2498 2258
rect 2436 2240 2498 2256
rect 2542 2251 2558 2254
rect 2620 2251 2650 2262
rect 2698 2258 2744 2274
rect 2771 2262 2845 2278
rect 2698 2256 2732 2258
rect 2697 2240 2744 2256
rect 2771 2240 2784 2262
rect 2799 2240 2829 2262
rect 2856 2240 2857 2256
rect 2872 2240 2885 2400
rect 2915 2296 2928 2400
rect 2973 2378 2974 2388
rect 2989 2378 3002 2388
rect 2973 2374 3002 2378
rect 3007 2374 3037 2400
rect 3055 2386 3071 2388
rect 3143 2386 3196 2400
rect 3144 2384 3208 2386
rect 3251 2384 3266 2400
rect 3315 2397 3345 2400
rect 3315 2394 3351 2397
rect 3281 2386 3297 2388
rect 3055 2374 3070 2378
rect 2973 2372 3070 2374
rect 3098 2372 3266 2384
rect 3282 2374 3297 2378
rect 3315 2375 3354 2394
rect 3373 2388 3380 2389
rect 3379 2381 3380 2388
rect 3363 2378 3364 2381
rect 3379 2378 3392 2381
rect 3315 2374 3345 2375
rect 3354 2374 3360 2375
rect 3363 2374 3392 2378
rect 3282 2373 3392 2374
rect 3282 2372 3398 2373
rect 2957 2364 3008 2372
rect 2957 2352 2982 2364
rect 2989 2352 3008 2364
rect 3039 2364 3089 2372
rect 3039 2356 3055 2364
rect 3062 2362 3089 2364
rect 3098 2362 3319 2372
rect 3062 2352 3319 2362
rect 3348 2364 3398 2372
rect 3348 2355 3364 2364
rect 2957 2344 3008 2352
rect 3055 2344 3319 2352
rect 3345 2352 3364 2355
rect 3371 2352 3398 2364
rect 3345 2344 3398 2352
rect 2973 2336 2974 2344
rect 2989 2336 3002 2344
rect 2973 2328 2989 2336
rect 2970 2321 2989 2324
rect 2970 2312 2992 2321
rect 2943 2302 2992 2312
rect 2943 2296 2973 2302
rect 2992 2297 2997 2302
rect 2915 2280 2989 2296
rect 3007 2288 3037 2344
rect 3072 2334 3280 2344
rect 3315 2340 3360 2344
rect 3363 2343 3364 2344
rect 3379 2343 3392 2344
rect 3098 2304 3287 2334
rect 3113 2301 3287 2304
rect 3106 2298 3287 2301
rect 2915 2278 2928 2280
rect 2943 2278 2977 2280
rect 2915 2262 2989 2278
rect 3016 2274 3029 2288
rect 3044 2274 3060 2290
rect 3106 2285 3117 2298
rect 2899 2240 2900 2256
rect 2915 2240 2928 2262
rect 2943 2240 2973 2262
rect 3016 2258 3078 2274
rect 3106 2267 3117 2283
rect 3122 2278 3132 2298
rect 3142 2278 3156 2298
rect 3159 2285 3168 2298
rect 3184 2285 3193 2298
rect 3122 2267 3156 2278
rect 3159 2267 3168 2283
rect 3184 2267 3193 2283
rect 3200 2278 3210 2298
rect 3220 2278 3234 2298
rect 3235 2285 3246 2298
rect 3200 2267 3234 2278
rect 3235 2267 3246 2283
rect 3292 2274 3308 2290
rect 3315 2288 3345 2340
rect 3379 2336 3380 2343
rect 3364 2328 3380 2336
rect 3351 2296 3364 2315
rect 3379 2296 3409 2312
rect 3351 2280 3425 2296
rect 3351 2278 3364 2280
rect 3379 2278 3413 2280
rect 3016 2256 3029 2258
rect 3044 2256 3078 2258
rect 3016 2240 3078 2256
rect 3122 2251 3138 2254
rect 3200 2251 3230 2262
rect 3278 2258 3324 2274
rect 3351 2262 3425 2278
rect 3278 2256 3312 2258
rect 3277 2240 3324 2256
rect 3351 2240 3364 2262
rect 3379 2240 3409 2262
rect 3436 2240 3437 2256
rect 3452 2240 3465 2400
rect 3495 2296 3508 2400
rect 3553 2378 3554 2388
rect 3569 2378 3582 2388
rect 3553 2374 3582 2378
rect 3587 2374 3617 2400
rect 3635 2386 3651 2388
rect 3723 2386 3776 2400
rect 3724 2384 3788 2386
rect 3831 2384 3846 2400
rect 3895 2397 3925 2400
rect 3895 2394 3931 2397
rect 3861 2386 3877 2388
rect 3635 2374 3650 2378
rect 3553 2372 3650 2374
rect 3678 2372 3846 2384
rect 3862 2374 3877 2378
rect 3895 2375 3934 2394
rect 3953 2388 3960 2389
rect 3959 2381 3960 2388
rect 3943 2378 3944 2381
rect 3959 2378 3972 2381
rect 3895 2374 3925 2375
rect 3934 2374 3940 2375
rect 3943 2374 3972 2378
rect 3862 2373 3972 2374
rect 3862 2372 3978 2373
rect 3537 2364 3588 2372
rect 3537 2352 3562 2364
rect 3569 2352 3588 2364
rect 3619 2364 3669 2372
rect 3619 2356 3635 2364
rect 3642 2362 3669 2364
rect 3678 2362 3899 2372
rect 3642 2352 3899 2362
rect 3928 2364 3978 2372
rect 3928 2355 3944 2364
rect 3537 2344 3588 2352
rect 3635 2344 3899 2352
rect 3925 2352 3944 2355
rect 3951 2352 3978 2364
rect 3925 2344 3978 2352
rect 3553 2336 3554 2344
rect 3569 2336 3582 2344
rect 3553 2328 3569 2336
rect 3550 2321 3569 2324
rect 3550 2312 3572 2321
rect 3523 2302 3572 2312
rect 3523 2296 3553 2302
rect 3572 2297 3577 2302
rect 3495 2280 3569 2296
rect 3587 2288 3617 2344
rect 3652 2334 3860 2344
rect 3895 2340 3940 2344
rect 3943 2343 3944 2344
rect 3959 2343 3972 2344
rect 3678 2304 3867 2334
rect 3693 2301 3867 2304
rect 3686 2298 3867 2301
rect 3495 2278 3508 2280
rect 3523 2278 3557 2280
rect 3495 2262 3569 2278
rect 3596 2274 3609 2288
rect 3624 2274 3640 2290
rect 3686 2285 3697 2298
rect 3479 2240 3480 2256
rect 3495 2240 3508 2262
rect 3523 2240 3553 2262
rect 3596 2258 3658 2274
rect 3686 2267 3697 2283
rect 3702 2278 3712 2298
rect 3722 2278 3736 2298
rect 3739 2285 3748 2298
rect 3764 2285 3773 2298
rect 3702 2267 3736 2278
rect 3739 2267 3748 2283
rect 3764 2267 3773 2283
rect 3780 2278 3790 2298
rect 3800 2278 3814 2298
rect 3815 2285 3826 2298
rect 3780 2267 3814 2278
rect 3815 2267 3826 2283
rect 3872 2274 3888 2290
rect 3895 2288 3925 2340
rect 3959 2336 3960 2343
rect 3944 2328 3960 2336
rect 3931 2296 3944 2315
rect 3959 2296 3989 2312
rect 3931 2280 4005 2296
rect 3931 2278 3944 2280
rect 3959 2278 3993 2280
rect 3596 2256 3609 2258
rect 3624 2256 3658 2258
rect 3596 2240 3658 2256
rect 3702 2251 3718 2254
rect 3780 2251 3810 2262
rect 3858 2258 3904 2274
rect 3931 2262 4005 2278
rect 3858 2256 3892 2258
rect 3857 2240 3904 2256
rect 3931 2240 3944 2262
rect 3959 2240 3989 2262
rect 4016 2240 4017 2256
rect 4032 2240 4045 2400
rect 4075 2296 4088 2400
rect 4133 2378 4134 2388
rect 4149 2378 4162 2388
rect 4133 2374 4162 2378
rect 4167 2374 4197 2400
rect 4215 2386 4231 2388
rect 4303 2386 4356 2400
rect 4304 2384 4368 2386
rect 4411 2384 4426 2400
rect 4475 2397 4505 2400
rect 4475 2394 4511 2397
rect 4441 2386 4457 2388
rect 4215 2374 4230 2378
rect 4133 2372 4230 2374
rect 4258 2372 4426 2384
rect 4442 2374 4457 2378
rect 4475 2375 4514 2394
rect 4533 2388 4540 2389
rect 4539 2381 4540 2388
rect 4523 2378 4524 2381
rect 4539 2378 4552 2381
rect 4475 2374 4505 2375
rect 4514 2374 4520 2375
rect 4523 2374 4552 2378
rect 4442 2373 4552 2374
rect 4442 2372 4558 2373
rect 4117 2364 4168 2372
rect 4117 2352 4142 2364
rect 4149 2352 4168 2364
rect 4199 2364 4249 2372
rect 4199 2356 4215 2364
rect 4222 2362 4249 2364
rect 4258 2362 4479 2372
rect 4222 2352 4479 2362
rect 4508 2364 4558 2372
rect 4508 2355 4524 2364
rect 4117 2344 4168 2352
rect 4215 2344 4479 2352
rect 4505 2352 4524 2355
rect 4531 2352 4558 2364
rect 4505 2344 4558 2352
rect 4133 2336 4134 2344
rect 4149 2336 4162 2344
rect 4133 2328 4149 2336
rect 4130 2321 4149 2324
rect 4130 2312 4152 2321
rect 4103 2302 4152 2312
rect 4103 2296 4133 2302
rect 4152 2297 4157 2302
rect 4075 2280 4149 2296
rect 4167 2288 4197 2344
rect 4232 2334 4440 2344
rect 4475 2340 4520 2344
rect 4523 2343 4524 2344
rect 4539 2343 4552 2344
rect 4258 2304 4447 2334
rect 4273 2301 4447 2304
rect 4266 2298 4447 2301
rect 4075 2278 4088 2280
rect 4103 2278 4137 2280
rect 4075 2262 4149 2278
rect 4176 2274 4189 2288
rect 4204 2274 4220 2290
rect 4266 2285 4277 2298
rect 4059 2240 4060 2256
rect 4075 2240 4088 2262
rect 4103 2240 4133 2262
rect 4176 2258 4238 2274
rect 4266 2267 4277 2283
rect 4282 2278 4292 2298
rect 4302 2278 4316 2298
rect 4319 2285 4328 2298
rect 4344 2285 4353 2298
rect 4282 2267 4316 2278
rect 4319 2267 4328 2283
rect 4344 2267 4353 2283
rect 4360 2278 4370 2298
rect 4380 2278 4394 2298
rect 4395 2285 4406 2298
rect 4360 2267 4394 2278
rect 4395 2267 4406 2283
rect 4452 2274 4468 2290
rect 4475 2288 4505 2340
rect 4539 2336 4540 2343
rect 4524 2328 4540 2336
rect 4511 2296 4524 2315
rect 4539 2296 4569 2312
rect 4511 2280 4585 2296
rect 4511 2278 4524 2280
rect 4539 2278 4573 2280
rect 4176 2256 4189 2258
rect 4204 2256 4238 2258
rect 4176 2240 4238 2256
rect 4282 2251 4298 2254
rect 4360 2251 4390 2262
rect 4438 2258 4484 2274
rect 4511 2262 4585 2278
rect 4438 2256 4472 2258
rect 4437 2240 4484 2256
rect 4511 2240 4524 2262
rect 4539 2240 4569 2262
rect 4596 2240 4597 2256
rect 4612 2240 4625 2400
rect -7 2232 34 2240
rect -7 2206 8 2232
rect 15 2206 34 2232
rect 98 2228 160 2240
rect 172 2228 247 2240
rect 305 2228 380 2240
rect 392 2228 423 2240
rect 429 2228 464 2240
rect 98 2226 260 2228
rect -7 2198 34 2206
rect 116 2202 129 2226
rect 144 2224 159 2226
rect -1 2188 0 2198
rect 15 2188 28 2198
rect 43 2188 73 2202
rect 116 2188 159 2202
rect 183 2199 190 2206
rect 193 2202 260 2226
rect 292 2226 464 2228
rect 262 2204 290 2208
rect 292 2204 372 2226
rect 393 2224 408 2226
rect 262 2202 372 2204
rect 193 2198 372 2202
rect 166 2188 196 2198
rect 198 2188 351 2198
rect 359 2188 389 2198
rect 393 2188 423 2202
rect 451 2188 464 2226
rect 536 2232 571 2240
rect 536 2206 537 2232
rect 544 2206 571 2232
rect 479 2188 509 2202
rect 536 2198 571 2206
rect 573 2232 614 2240
rect 573 2206 588 2232
rect 595 2206 614 2232
rect 678 2228 740 2240
rect 752 2228 827 2240
rect 885 2228 960 2240
rect 972 2228 1003 2240
rect 1009 2228 1044 2240
rect 678 2226 840 2228
rect 573 2198 614 2206
rect 696 2202 709 2226
rect 724 2224 739 2226
rect 536 2188 537 2198
rect 552 2188 565 2198
rect 579 2188 580 2198
rect 595 2188 608 2198
rect 623 2188 653 2202
rect 696 2188 739 2202
rect 763 2199 770 2206
rect 773 2202 840 2226
rect 872 2226 1044 2228
rect 842 2204 870 2208
rect 872 2204 952 2226
rect 973 2224 988 2226
rect 842 2202 952 2204
rect 773 2198 952 2202
rect 746 2188 776 2198
rect 778 2188 931 2198
rect 939 2188 969 2198
rect 973 2188 1003 2202
rect 1031 2188 1044 2226
rect 1116 2232 1151 2240
rect 1116 2206 1117 2232
rect 1124 2206 1151 2232
rect 1059 2188 1089 2202
rect 1116 2198 1151 2206
rect 1153 2232 1194 2240
rect 1153 2206 1168 2232
rect 1175 2206 1194 2232
rect 1258 2228 1320 2240
rect 1332 2228 1407 2240
rect 1465 2228 1540 2240
rect 1552 2228 1583 2240
rect 1589 2228 1624 2240
rect 1258 2226 1420 2228
rect 1153 2198 1194 2206
rect 1276 2202 1289 2226
rect 1304 2224 1319 2226
rect 1116 2188 1117 2198
rect 1132 2188 1145 2198
rect 1159 2188 1160 2198
rect 1175 2188 1188 2198
rect 1203 2188 1233 2202
rect 1276 2188 1319 2202
rect 1343 2199 1350 2206
rect 1353 2202 1420 2226
rect 1452 2226 1624 2228
rect 1422 2204 1450 2208
rect 1452 2204 1532 2226
rect 1553 2224 1568 2226
rect 1422 2202 1532 2204
rect 1353 2198 1532 2202
rect 1326 2188 1356 2198
rect 1358 2188 1511 2198
rect 1519 2188 1549 2198
rect 1553 2188 1583 2202
rect 1611 2188 1624 2226
rect 1696 2232 1731 2240
rect 1696 2206 1697 2232
rect 1704 2206 1731 2232
rect 1639 2188 1669 2202
rect 1696 2198 1731 2206
rect 1733 2232 1774 2240
rect 1733 2206 1748 2232
rect 1755 2206 1774 2232
rect 1838 2228 1900 2240
rect 1912 2228 1987 2240
rect 2045 2228 2120 2240
rect 2132 2228 2163 2240
rect 2169 2228 2204 2240
rect 1838 2226 2000 2228
rect 1733 2198 1774 2206
rect 1856 2202 1869 2226
rect 1884 2224 1899 2226
rect 1696 2188 1697 2198
rect 1712 2188 1725 2198
rect 1739 2188 1740 2198
rect 1755 2188 1768 2198
rect 1783 2188 1813 2202
rect 1856 2188 1899 2202
rect 1923 2199 1930 2206
rect 1933 2202 2000 2226
rect 2032 2226 2204 2228
rect 2002 2204 2030 2208
rect 2032 2204 2112 2226
rect 2133 2224 2148 2226
rect 2002 2202 2112 2204
rect 1933 2198 2112 2202
rect 1906 2188 1936 2198
rect 1938 2188 2091 2198
rect 2099 2188 2129 2198
rect 2133 2188 2163 2202
rect 2191 2188 2204 2226
rect 2276 2232 2311 2240
rect 2276 2206 2277 2232
rect 2284 2206 2311 2232
rect 2219 2188 2249 2202
rect 2276 2198 2311 2206
rect 2313 2232 2354 2240
rect 2313 2206 2328 2232
rect 2335 2206 2354 2232
rect 2418 2228 2480 2240
rect 2492 2228 2567 2240
rect 2625 2228 2700 2240
rect 2712 2228 2743 2240
rect 2749 2228 2784 2240
rect 2418 2226 2580 2228
rect 2313 2198 2354 2206
rect 2436 2202 2449 2226
rect 2464 2224 2479 2226
rect 2276 2188 2277 2198
rect 2292 2188 2305 2198
rect 2319 2188 2320 2198
rect 2335 2188 2348 2198
rect 2363 2188 2393 2202
rect 2436 2188 2479 2202
rect 2503 2199 2510 2206
rect 2513 2202 2580 2226
rect 2612 2226 2784 2228
rect 2582 2204 2610 2208
rect 2612 2204 2692 2226
rect 2713 2224 2728 2226
rect 2582 2202 2692 2204
rect 2513 2198 2692 2202
rect 2486 2188 2516 2198
rect 2518 2188 2671 2198
rect 2679 2188 2709 2198
rect 2713 2188 2743 2202
rect 2771 2188 2784 2226
rect 2856 2232 2891 2240
rect 2856 2206 2857 2232
rect 2864 2206 2891 2232
rect 2799 2188 2829 2202
rect 2856 2198 2891 2206
rect 2893 2232 2934 2240
rect 2893 2206 2908 2232
rect 2915 2206 2934 2232
rect 2998 2228 3060 2240
rect 3072 2228 3147 2240
rect 3205 2228 3280 2240
rect 3292 2228 3323 2240
rect 3329 2228 3364 2240
rect 2998 2226 3160 2228
rect 2893 2198 2934 2206
rect 3016 2202 3029 2226
rect 3044 2224 3059 2226
rect 2856 2188 2857 2198
rect 2872 2188 2885 2198
rect 2899 2188 2900 2198
rect 2915 2188 2928 2198
rect 2943 2188 2973 2202
rect 3016 2188 3059 2202
rect 3083 2199 3090 2206
rect 3093 2202 3160 2226
rect 3192 2226 3364 2228
rect 3162 2204 3190 2208
rect 3192 2204 3272 2226
rect 3293 2224 3308 2226
rect 3162 2202 3272 2204
rect 3093 2198 3272 2202
rect 3066 2188 3096 2198
rect 3098 2188 3251 2198
rect 3259 2188 3289 2198
rect 3293 2188 3323 2202
rect 3351 2188 3364 2226
rect 3436 2232 3471 2240
rect 3436 2206 3437 2232
rect 3444 2206 3471 2232
rect 3379 2188 3409 2202
rect 3436 2198 3471 2206
rect 3473 2232 3514 2240
rect 3473 2206 3488 2232
rect 3495 2206 3514 2232
rect 3578 2228 3640 2240
rect 3652 2228 3727 2240
rect 3785 2228 3860 2240
rect 3872 2228 3903 2240
rect 3909 2228 3944 2240
rect 3578 2226 3740 2228
rect 3473 2198 3514 2206
rect 3596 2202 3609 2226
rect 3624 2224 3639 2226
rect 3436 2188 3437 2198
rect 3452 2188 3465 2198
rect 3479 2188 3480 2198
rect 3495 2188 3508 2198
rect 3523 2188 3553 2202
rect 3596 2188 3639 2202
rect 3663 2199 3670 2206
rect 3673 2202 3740 2226
rect 3772 2226 3944 2228
rect 3742 2204 3770 2208
rect 3772 2204 3852 2226
rect 3873 2224 3888 2226
rect 3742 2202 3852 2204
rect 3673 2198 3852 2202
rect 3646 2188 3676 2198
rect 3678 2188 3831 2198
rect 3839 2188 3869 2198
rect 3873 2188 3903 2202
rect 3931 2188 3944 2226
rect 4016 2232 4051 2240
rect 4016 2206 4017 2232
rect 4024 2206 4051 2232
rect 3959 2188 3989 2202
rect 4016 2198 4051 2206
rect 4053 2232 4094 2240
rect 4053 2206 4068 2232
rect 4075 2206 4094 2232
rect 4158 2228 4220 2240
rect 4232 2228 4307 2240
rect 4365 2228 4440 2240
rect 4452 2228 4483 2240
rect 4489 2228 4524 2240
rect 4158 2226 4320 2228
rect 4053 2198 4094 2206
rect 4176 2202 4189 2226
rect 4204 2224 4219 2226
rect 4016 2188 4017 2198
rect 4032 2188 4045 2198
rect 4059 2188 4060 2198
rect 4075 2188 4088 2198
rect 4103 2188 4133 2202
rect 4176 2188 4219 2202
rect 4243 2199 4250 2206
rect 4253 2202 4320 2226
rect 4352 2226 4524 2228
rect 4322 2204 4350 2208
rect 4352 2204 4432 2226
rect 4453 2224 4468 2226
rect 4322 2202 4432 2204
rect 4253 2198 4432 2202
rect 4226 2188 4256 2198
rect 4258 2188 4411 2198
rect 4419 2188 4449 2198
rect 4453 2188 4483 2202
rect 4511 2188 4524 2226
rect 4596 2232 4631 2240
rect 4596 2206 4597 2232
rect 4604 2206 4631 2232
rect 4539 2188 4569 2202
rect 4596 2198 4631 2206
rect 4596 2188 4597 2198
rect 4612 2188 4625 2198
rect -1 2182 4625 2188
rect 0 2174 4625 2182
rect 15 2144 28 2174
rect 43 2156 73 2174
rect 116 2160 130 2174
rect 166 2160 386 2174
rect 117 2158 130 2160
rect 83 2146 98 2158
rect 80 2144 102 2146
rect 107 2144 137 2158
rect 198 2156 351 2160
rect 180 2144 372 2156
rect 415 2144 445 2158
rect 451 2144 464 2174
rect 479 2156 509 2174
rect 552 2144 565 2174
rect 595 2144 608 2174
rect 623 2156 653 2174
rect 696 2160 710 2174
rect 746 2160 966 2174
rect 697 2158 710 2160
rect 663 2146 678 2158
rect 660 2144 682 2146
rect 687 2144 717 2158
rect 778 2156 931 2160
rect 760 2144 952 2156
rect 995 2144 1025 2158
rect 1031 2144 1044 2174
rect 1059 2156 1089 2174
rect 1132 2144 1145 2174
rect 1175 2144 1188 2174
rect 1203 2156 1233 2174
rect 1276 2160 1290 2174
rect 1326 2160 1546 2174
rect 1277 2158 1290 2160
rect 1243 2146 1258 2158
rect 1240 2144 1262 2146
rect 1267 2144 1297 2158
rect 1358 2156 1511 2160
rect 1340 2144 1532 2156
rect 1575 2144 1605 2158
rect 1611 2144 1624 2174
rect 1639 2156 1669 2174
rect 1712 2144 1725 2174
rect 1755 2144 1768 2174
rect 1783 2156 1813 2174
rect 1856 2160 1870 2174
rect 1906 2160 2126 2174
rect 1857 2158 1870 2160
rect 1823 2146 1838 2158
rect 1820 2144 1842 2146
rect 1847 2144 1877 2158
rect 1938 2156 2091 2160
rect 1920 2144 2112 2156
rect 2155 2144 2185 2158
rect 2191 2144 2204 2174
rect 2219 2156 2249 2174
rect 2292 2144 2305 2174
rect 2335 2144 2348 2174
rect 2363 2156 2393 2174
rect 2436 2160 2450 2174
rect 2486 2160 2706 2174
rect 2437 2158 2450 2160
rect 2403 2146 2418 2158
rect 2400 2144 2422 2146
rect 2427 2144 2457 2158
rect 2518 2156 2671 2160
rect 2500 2144 2692 2156
rect 2735 2144 2765 2158
rect 2771 2144 2784 2174
rect 2799 2156 2829 2174
rect 2872 2144 2885 2174
rect 2915 2144 2928 2174
rect 2943 2156 2973 2174
rect 3016 2160 3030 2174
rect 3066 2160 3286 2174
rect 3017 2158 3030 2160
rect 2983 2146 2998 2158
rect 2980 2144 3002 2146
rect 3007 2144 3037 2158
rect 3098 2156 3251 2160
rect 3080 2144 3272 2156
rect 3315 2144 3345 2158
rect 3351 2144 3364 2174
rect 3379 2156 3409 2174
rect 3452 2144 3465 2174
rect 3495 2144 3508 2174
rect 3523 2156 3553 2174
rect 3596 2160 3610 2174
rect 3646 2160 3866 2174
rect 3597 2158 3610 2160
rect 3563 2146 3578 2158
rect 3560 2144 3582 2146
rect 3587 2144 3617 2158
rect 3678 2156 3831 2160
rect 3660 2144 3852 2156
rect 3895 2144 3925 2158
rect 3931 2144 3944 2174
rect 3959 2156 3989 2174
rect 4032 2144 4045 2174
rect 4075 2144 4088 2174
rect 4103 2156 4133 2174
rect 4176 2160 4190 2174
rect 4226 2160 4446 2174
rect 4177 2158 4190 2160
rect 4143 2146 4158 2158
rect 4140 2144 4162 2146
rect 4167 2144 4197 2158
rect 4258 2156 4411 2160
rect 4240 2144 4432 2156
rect 4475 2144 4505 2158
rect 4511 2144 4524 2174
rect 4539 2156 4569 2174
rect 4612 2144 4625 2174
rect 0 2130 4625 2144
rect 15 2026 28 2130
rect 73 2108 74 2118
rect 89 2108 102 2118
rect 73 2104 102 2108
rect 107 2104 137 2130
rect 155 2116 171 2118
rect 243 2116 296 2130
rect 244 2114 308 2116
rect 351 2114 366 2130
rect 415 2127 445 2130
rect 415 2124 451 2127
rect 381 2116 397 2118
rect 155 2104 170 2108
rect 73 2102 170 2104
rect 198 2102 366 2114
rect 382 2104 397 2108
rect 415 2105 454 2124
rect 473 2118 480 2119
rect 479 2111 480 2118
rect 463 2108 464 2111
rect 479 2108 492 2111
rect 415 2104 445 2105
rect 454 2104 460 2105
rect 463 2104 492 2108
rect 382 2103 492 2104
rect 382 2102 498 2103
rect 57 2094 108 2102
rect 57 2082 82 2094
rect 89 2082 108 2094
rect 139 2094 189 2102
rect 139 2086 155 2094
rect 162 2092 189 2094
rect 198 2092 419 2102
rect 162 2082 419 2092
rect 448 2094 498 2102
rect 448 2085 464 2094
rect 57 2074 108 2082
rect 155 2074 419 2082
rect 445 2082 464 2085
rect 471 2082 498 2094
rect 445 2074 498 2082
rect 73 2066 74 2074
rect 89 2066 102 2074
rect 73 2058 89 2066
rect 70 2051 89 2054
rect 70 2042 92 2051
rect 43 2032 92 2042
rect 43 2026 73 2032
rect 92 2027 97 2032
rect 15 2010 89 2026
rect 107 2018 137 2074
rect 172 2064 380 2074
rect 415 2070 460 2074
rect 463 2073 464 2074
rect 479 2073 492 2074
rect 198 2034 387 2064
rect 213 2031 387 2034
rect 206 2028 387 2031
rect 15 2008 28 2010
rect 43 2008 77 2010
rect 15 1992 89 2008
rect 116 2004 129 2018
rect 144 2004 160 2020
rect 206 2015 217 2028
rect -1 1970 0 1986
rect 15 1970 28 1992
rect 43 1970 73 1992
rect 116 1988 178 2004
rect 206 1997 217 2013
rect 222 2008 232 2028
rect 242 2008 256 2028
rect 259 2015 268 2028
rect 284 2015 293 2028
rect 222 1997 256 2008
rect 259 1997 268 2013
rect 284 1997 293 2013
rect 300 2008 310 2028
rect 320 2008 334 2028
rect 335 2015 346 2028
rect 300 1997 334 2008
rect 335 1997 346 2013
rect 392 2004 408 2020
rect 415 2018 445 2070
rect 479 2066 480 2073
rect 464 2058 480 2066
rect 451 2026 464 2045
rect 479 2026 509 2042
rect 451 2010 525 2026
rect 451 2008 464 2010
rect 479 2008 513 2010
rect 116 1986 129 1988
rect 144 1986 178 1988
rect 116 1970 178 1986
rect 222 1981 238 1984
rect 300 1981 330 1992
rect 378 1988 424 2004
rect 451 1992 525 2008
rect 378 1986 412 1988
rect 377 1970 424 1986
rect 451 1970 464 1992
rect 479 1970 509 1992
rect 536 1970 537 1986
rect 552 1970 565 2130
rect 595 2026 608 2130
rect 653 2108 654 2118
rect 669 2108 682 2118
rect 653 2104 682 2108
rect 687 2104 717 2130
rect 735 2116 751 2118
rect 823 2116 876 2130
rect 824 2114 888 2116
rect 931 2114 946 2130
rect 995 2127 1025 2130
rect 995 2124 1031 2127
rect 961 2116 977 2118
rect 735 2104 750 2108
rect 653 2102 750 2104
rect 778 2102 946 2114
rect 962 2104 977 2108
rect 995 2105 1034 2124
rect 1053 2118 1060 2119
rect 1059 2111 1060 2118
rect 1043 2108 1044 2111
rect 1059 2108 1072 2111
rect 995 2104 1025 2105
rect 1034 2104 1040 2105
rect 1043 2104 1072 2108
rect 962 2103 1072 2104
rect 962 2102 1078 2103
rect 637 2094 688 2102
rect 637 2082 662 2094
rect 669 2082 688 2094
rect 719 2094 769 2102
rect 719 2086 735 2094
rect 742 2092 769 2094
rect 778 2092 999 2102
rect 742 2082 999 2092
rect 1028 2094 1078 2102
rect 1028 2085 1044 2094
rect 637 2074 688 2082
rect 735 2074 999 2082
rect 1025 2082 1044 2085
rect 1051 2082 1078 2094
rect 1025 2074 1078 2082
rect 653 2066 654 2074
rect 669 2066 682 2074
rect 653 2058 669 2066
rect 650 2051 669 2054
rect 650 2042 672 2051
rect 623 2032 672 2042
rect 623 2026 653 2032
rect 672 2027 677 2032
rect 595 2010 669 2026
rect 687 2018 717 2074
rect 752 2064 960 2074
rect 995 2070 1040 2074
rect 1043 2073 1044 2074
rect 1059 2073 1072 2074
rect 778 2034 967 2064
rect 793 2031 967 2034
rect 786 2028 967 2031
rect 595 2008 608 2010
rect 623 2008 657 2010
rect 595 1992 669 2008
rect 696 2004 709 2018
rect 724 2004 740 2020
rect 786 2015 797 2028
rect 579 1970 580 1986
rect 595 1970 608 1992
rect 623 1970 653 1992
rect 696 1988 758 2004
rect 786 1997 797 2013
rect 802 2008 812 2028
rect 822 2008 836 2028
rect 839 2015 848 2028
rect 864 2015 873 2028
rect 802 1997 836 2008
rect 839 1997 848 2013
rect 864 1997 873 2013
rect 880 2008 890 2028
rect 900 2008 914 2028
rect 915 2015 926 2028
rect 880 1997 914 2008
rect 915 1997 926 2013
rect 972 2004 988 2020
rect 995 2018 1025 2070
rect 1059 2066 1060 2073
rect 1044 2058 1060 2066
rect 1031 2026 1044 2045
rect 1059 2026 1089 2042
rect 1031 2010 1105 2026
rect 1031 2008 1044 2010
rect 1059 2008 1093 2010
rect 696 1986 709 1988
rect 724 1986 758 1988
rect 696 1970 758 1986
rect 802 1981 818 1984
rect 880 1981 910 1992
rect 958 1988 1004 2004
rect 1031 1992 1105 2008
rect 958 1986 992 1988
rect 957 1970 1004 1986
rect 1031 1970 1044 1992
rect 1059 1970 1089 1992
rect 1116 1970 1117 1986
rect 1132 1970 1145 2130
rect 1175 2026 1188 2130
rect 1233 2108 1234 2118
rect 1249 2108 1262 2118
rect 1233 2104 1262 2108
rect 1267 2104 1297 2130
rect 1315 2116 1331 2118
rect 1403 2116 1456 2130
rect 1404 2114 1468 2116
rect 1511 2114 1526 2130
rect 1575 2127 1605 2130
rect 1575 2124 1611 2127
rect 1541 2116 1557 2118
rect 1315 2104 1330 2108
rect 1233 2102 1330 2104
rect 1358 2102 1526 2114
rect 1542 2104 1557 2108
rect 1575 2105 1614 2124
rect 1633 2118 1640 2119
rect 1639 2111 1640 2118
rect 1623 2108 1624 2111
rect 1639 2108 1652 2111
rect 1575 2104 1605 2105
rect 1614 2104 1620 2105
rect 1623 2104 1652 2108
rect 1542 2103 1652 2104
rect 1542 2102 1658 2103
rect 1217 2094 1268 2102
rect 1217 2082 1242 2094
rect 1249 2082 1268 2094
rect 1299 2094 1349 2102
rect 1299 2086 1315 2094
rect 1322 2092 1349 2094
rect 1358 2092 1579 2102
rect 1322 2082 1579 2092
rect 1608 2094 1658 2102
rect 1608 2085 1624 2094
rect 1217 2074 1268 2082
rect 1315 2074 1579 2082
rect 1605 2082 1624 2085
rect 1631 2082 1658 2094
rect 1605 2074 1658 2082
rect 1233 2066 1234 2074
rect 1249 2066 1262 2074
rect 1233 2058 1249 2066
rect 1230 2051 1249 2054
rect 1230 2042 1252 2051
rect 1203 2032 1252 2042
rect 1203 2026 1233 2032
rect 1252 2027 1257 2032
rect 1175 2010 1249 2026
rect 1267 2018 1297 2074
rect 1332 2064 1540 2074
rect 1575 2070 1620 2074
rect 1623 2073 1624 2074
rect 1639 2073 1652 2074
rect 1358 2034 1547 2064
rect 1373 2031 1547 2034
rect 1366 2028 1547 2031
rect 1175 2008 1188 2010
rect 1203 2008 1237 2010
rect 1175 1992 1249 2008
rect 1276 2004 1289 2018
rect 1304 2004 1320 2020
rect 1366 2015 1377 2028
rect 1159 1970 1160 1986
rect 1175 1970 1188 1992
rect 1203 1970 1233 1992
rect 1276 1988 1338 2004
rect 1366 1997 1377 2013
rect 1382 2008 1392 2028
rect 1402 2008 1416 2028
rect 1419 2015 1428 2028
rect 1444 2015 1453 2028
rect 1382 1997 1416 2008
rect 1419 1997 1428 2013
rect 1444 1997 1453 2013
rect 1460 2008 1470 2028
rect 1480 2008 1494 2028
rect 1495 2015 1506 2028
rect 1460 1997 1494 2008
rect 1495 1997 1506 2013
rect 1552 2004 1568 2020
rect 1575 2018 1605 2070
rect 1639 2066 1640 2073
rect 1624 2058 1640 2066
rect 1611 2026 1624 2045
rect 1639 2026 1669 2042
rect 1611 2010 1685 2026
rect 1611 2008 1624 2010
rect 1639 2008 1673 2010
rect 1276 1986 1289 1988
rect 1304 1986 1338 1988
rect 1276 1970 1338 1986
rect 1382 1981 1398 1984
rect 1460 1981 1490 1992
rect 1538 1988 1584 2004
rect 1611 1992 1685 2008
rect 1538 1986 1572 1988
rect 1537 1970 1584 1986
rect 1611 1970 1624 1992
rect 1639 1970 1669 1992
rect 1696 1970 1697 1986
rect 1712 1970 1725 2130
rect 1755 2026 1768 2130
rect 1813 2108 1814 2118
rect 1829 2108 1842 2118
rect 1813 2104 1842 2108
rect 1847 2104 1877 2130
rect 1895 2116 1911 2118
rect 1983 2116 2036 2130
rect 1984 2114 2048 2116
rect 2091 2114 2106 2130
rect 2155 2127 2185 2130
rect 2155 2124 2191 2127
rect 2121 2116 2137 2118
rect 1895 2104 1910 2108
rect 1813 2102 1910 2104
rect 1938 2102 2106 2114
rect 2122 2104 2137 2108
rect 2155 2105 2194 2124
rect 2213 2118 2220 2119
rect 2219 2111 2220 2118
rect 2203 2108 2204 2111
rect 2219 2108 2232 2111
rect 2155 2104 2185 2105
rect 2194 2104 2200 2105
rect 2203 2104 2232 2108
rect 2122 2103 2232 2104
rect 2122 2102 2238 2103
rect 1797 2094 1848 2102
rect 1797 2082 1822 2094
rect 1829 2082 1848 2094
rect 1879 2094 1929 2102
rect 1879 2086 1895 2094
rect 1902 2092 1929 2094
rect 1938 2092 2159 2102
rect 1902 2082 2159 2092
rect 2188 2094 2238 2102
rect 2188 2085 2204 2094
rect 1797 2074 1848 2082
rect 1895 2074 2159 2082
rect 2185 2082 2204 2085
rect 2211 2082 2238 2094
rect 2185 2074 2238 2082
rect 1813 2066 1814 2074
rect 1829 2066 1842 2074
rect 1813 2058 1829 2066
rect 1810 2051 1829 2054
rect 1810 2042 1832 2051
rect 1783 2032 1832 2042
rect 1783 2026 1813 2032
rect 1832 2027 1837 2032
rect 1755 2010 1829 2026
rect 1847 2018 1877 2074
rect 1912 2064 2120 2074
rect 2155 2070 2200 2074
rect 2203 2073 2204 2074
rect 2219 2073 2232 2074
rect 1938 2034 2127 2064
rect 1953 2031 2127 2034
rect 1946 2028 2127 2031
rect 1755 2008 1768 2010
rect 1783 2008 1817 2010
rect 1755 1992 1829 2008
rect 1856 2004 1869 2018
rect 1884 2004 1900 2020
rect 1946 2015 1957 2028
rect 1739 1970 1740 1986
rect 1755 1970 1768 1992
rect 1783 1970 1813 1992
rect 1856 1988 1918 2004
rect 1946 1997 1957 2013
rect 1962 2008 1972 2028
rect 1982 2008 1996 2028
rect 1999 2015 2008 2028
rect 2024 2015 2033 2028
rect 1962 1997 1996 2008
rect 1999 1997 2008 2013
rect 2024 1997 2033 2013
rect 2040 2008 2050 2028
rect 2060 2008 2074 2028
rect 2075 2015 2086 2028
rect 2040 1997 2074 2008
rect 2075 1997 2086 2013
rect 2132 2004 2148 2020
rect 2155 2018 2185 2070
rect 2219 2066 2220 2073
rect 2204 2058 2220 2066
rect 2191 2026 2204 2045
rect 2219 2026 2249 2042
rect 2191 2010 2265 2026
rect 2191 2008 2204 2010
rect 2219 2008 2253 2010
rect 1856 1986 1869 1988
rect 1884 1986 1918 1988
rect 1856 1970 1918 1986
rect 1962 1981 1978 1984
rect 2040 1981 2070 1992
rect 2118 1988 2164 2004
rect 2191 1992 2265 2008
rect 2118 1986 2152 1988
rect 2117 1970 2164 1986
rect 2191 1970 2204 1992
rect 2219 1970 2249 1992
rect 2276 1970 2277 1986
rect 2292 1970 2305 2130
rect 2335 2026 2348 2130
rect 2393 2108 2394 2118
rect 2409 2108 2422 2118
rect 2393 2104 2422 2108
rect 2427 2104 2457 2130
rect 2475 2116 2491 2118
rect 2563 2116 2616 2130
rect 2564 2114 2628 2116
rect 2671 2114 2686 2130
rect 2735 2127 2765 2130
rect 2735 2124 2771 2127
rect 2701 2116 2717 2118
rect 2475 2104 2490 2108
rect 2393 2102 2490 2104
rect 2518 2102 2686 2114
rect 2702 2104 2717 2108
rect 2735 2105 2774 2124
rect 2793 2118 2800 2119
rect 2799 2111 2800 2118
rect 2783 2108 2784 2111
rect 2799 2108 2812 2111
rect 2735 2104 2765 2105
rect 2774 2104 2780 2105
rect 2783 2104 2812 2108
rect 2702 2103 2812 2104
rect 2702 2102 2818 2103
rect 2377 2094 2428 2102
rect 2377 2082 2402 2094
rect 2409 2082 2428 2094
rect 2459 2094 2509 2102
rect 2459 2086 2475 2094
rect 2482 2092 2509 2094
rect 2518 2092 2739 2102
rect 2482 2082 2739 2092
rect 2768 2094 2818 2102
rect 2768 2085 2784 2094
rect 2377 2074 2428 2082
rect 2475 2074 2739 2082
rect 2765 2082 2784 2085
rect 2791 2082 2818 2094
rect 2765 2074 2818 2082
rect 2393 2066 2394 2074
rect 2409 2066 2422 2074
rect 2393 2058 2409 2066
rect 2390 2051 2409 2054
rect 2390 2042 2412 2051
rect 2363 2032 2412 2042
rect 2363 2026 2393 2032
rect 2412 2027 2417 2032
rect 2335 2010 2409 2026
rect 2427 2018 2457 2074
rect 2492 2064 2700 2074
rect 2735 2070 2780 2074
rect 2783 2073 2784 2074
rect 2799 2073 2812 2074
rect 2518 2034 2707 2064
rect 2533 2031 2707 2034
rect 2526 2028 2707 2031
rect 2335 2008 2348 2010
rect 2363 2008 2397 2010
rect 2335 1992 2409 2008
rect 2436 2004 2449 2018
rect 2464 2004 2480 2020
rect 2526 2015 2537 2028
rect 2319 1970 2320 1986
rect 2335 1970 2348 1992
rect 2363 1970 2393 1992
rect 2436 1988 2498 2004
rect 2526 1997 2537 2013
rect 2542 2008 2552 2028
rect 2562 2008 2576 2028
rect 2579 2015 2588 2028
rect 2604 2015 2613 2028
rect 2542 1997 2576 2008
rect 2579 1997 2588 2013
rect 2604 1997 2613 2013
rect 2620 2008 2630 2028
rect 2640 2008 2654 2028
rect 2655 2015 2666 2028
rect 2620 1997 2654 2008
rect 2655 1997 2666 2013
rect 2712 2004 2728 2020
rect 2735 2018 2765 2070
rect 2799 2066 2800 2073
rect 2784 2058 2800 2066
rect 2771 2026 2784 2045
rect 2799 2026 2829 2042
rect 2771 2010 2845 2026
rect 2771 2008 2784 2010
rect 2799 2008 2833 2010
rect 2436 1986 2449 1988
rect 2464 1986 2498 1988
rect 2436 1970 2498 1986
rect 2542 1981 2558 1984
rect 2620 1981 2650 1992
rect 2698 1988 2744 2004
rect 2771 1992 2845 2008
rect 2698 1986 2732 1988
rect 2697 1970 2744 1986
rect 2771 1970 2784 1992
rect 2799 1970 2829 1992
rect 2856 1970 2857 1986
rect 2872 1970 2885 2130
rect 2915 2026 2928 2130
rect 2973 2108 2974 2118
rect 2989 2108 3002 2118
rect 2973 2104 3002 2108
rect 3007 2104 3037 2130
rect 3055 2116 3071 2118
rect 3143 2116 3196 2130
rect 3144 2114 3208 2116
rect 3251 2114 3266 2130
rect 3315 2127 3345 2130
rect 3315 2124 3351 2127
rect 3281 2116 3297 2118
rect 3055 2104 3070 2108
rect 2973 2102 3070 2104
rect 3098 2102 3266 2114
rect 3282 2104 3297 2108
rect 3315 2105 3354 2124
rect 3373 2118 3380 2119
rect 3379 2111 3380 2118
rect 3363 2108 3364 2111
rect 3379 2108 3392 2111
rect 3315 2104 3345 2105
rect 3354 2104 3360 2105
rect 3363 2104 3392 2108
rect 3282 2103 3392 2104
rect 3282 2102 3398 2103
rect 2957 2094 3008 2102
rect 2957 2082 2982 2094
rect 2989 2082 3008 2094
rect 3039 2094 3089 2102
rect 3039 2086 3055 2094
rect 3062 2092 3089 2094
rect 3098 2092 3319 2102
rect 3062 2082 3319 2092
rect 3348 2094 3398 2102
rect 3348 2085 3364 2094
rect 2957 2074 3008 2082
rect 3055 2074 3319 2082
rect 3345 2082 3364 2085
rect 3371 2082 3398 2094
rect 3345 2074 3398 2082
rect 2973 2066 2974 2074
rect 2989 2066 3002 2074
rect 2973 2058 2989 2066
rect 2970 2051 2989 2054
rect 2970 2042 2992 2051
rect 2943 2032 2992 2042
rect 2943 2026 2973 2032
rect 2992 2027 2997 2032
rect 2915 2010 2989 2026
rect 3007 2018 3037 2074
rect 3072 2064 3280 2074
rect 3315 2070 3360 2074
rect 3363 2073 3364 2074
rect 3379 2073 3392 2074
rect 3098 2034 3287 2064
rect 3113 2031 3287 2034
rect 3106 2028 3287 2031
rect 2915 2008 2928 2010
rect 2943 2008 2977 2010
rect 2915 1992 2989 2008
rect 3016 2004 3029 2018
rect 3044 2004 3060 2020
rect 3106 2015 3117 2028
rect 2899 1970 2900 1986
rect 2915 1970 2928 1992
rect 2943 1970 2973 1992
rect 3016 1988 3078 2004
rect 3106 1997 3117 2013
rect 3122 2008 3132 2028
rect 3142 2008 3156 2028
rect 3159 2015 3168 2028
rect 3184 2015 3193 2028
rect 3122 1997 3156 2008
rect 3159 1997 3168 2013
rect 3184 1997 3193 2013
rect 3200 2008 3210 2028
rect 3220 2008 3234 2028
rect 3235 2015 3246 2028
rect 3200 1997 3234 2008
rect 3235 1997 3246 2013
rect 3292 2004 3308 2020
rect 3315 2018 3345 2070
rect 3379 2066 3380 2073
rect 3364 2058 3380 2066
rect 3351 2026 3364 2045
rect 3379 2026 3409 2042
rect 3351 2010 3425 2026
rect 3351 2008 3364 2010
rect 3379 2008 3413 2010
rect 3016 1986 3029 1988
rect 3044 1986 3078 1988
rect 3016 1970 3078 1986
rect 3122 1981 3138 1984
rect 3200 1981 3230 1992
rect 3278 1988 3324 2004
rect 3351 1992 3425 2008
rect 3278 1986 3312 1988
rect 3277 1970 3324 1986
rect 3351 1970 3364 1992
rect 3379 1970 3409 1992
rect 3436 1970 3437 1986
rect 3452 1970 3465 2130
rect 3495 2026 3508 2130
rect 3553 2108 3554 2118
rect 3569 2108 3582 2118
rect 3553 2104 3582 2108
rect 3587 2104 3617 2130
rect 3635 2116 3651 2118
rect 3723 2116 3776 2130
rect 3724 2114 3788 2116
rect 3831 2114 3846 2130
rect 3895 2127 3925 2130
rect 3895 2124 3931 2127
rect 3861 2116 3877 2118
rect 3635 2104 3650 2108
rect 3553 2102 3650 2104
rect 3678 2102 3846 2114
rect 3862 2104 3877 2108
rect 3895 2105 3934 2124
rect 3953 2118 3960 2119
rect 3959 2111 3960 2118
rect 3943 2108 3944 2111
rect 3959 2108 3972 2111
rect 3895 2104 3925 2105
rect 3934 2104 3940 2105
rect 3943 2104 3972 2108
rect 3862 2103 3972 2104
rect 3862 2102 3978 2103
rect 3537 2094 3588 2102
rect 3537 2082 3562 2094
rect 3569 2082 3588 2094
rect 3619 2094 3669 2102
rect 3619 2086 3635 2094
rect 3642 2092 3669 2094
rect 3678 2092 3899 2102
rect 3642 2082 3899 2092
rect 3928 2094 3978 2102
rect 3928 2085 3944 2094
rect 3537 2074 3588 2082
rect 3635 2074 3899 2082
rect 3925 2082 3944 2085
rect 3951 2082 3978 2094
rect 3925 2074 3978 2082
rect 3553 2066 3554 2074
rect 3569 2066 3582 2074
rect 3553 2058 3569 2066
rect 3550 2051 3569 2054
rect 3550 2042 3572 2051
rect 3523 2032 3572 2042
rect 3523 2026 3553 2032
rect 3572 2027 3577 2032
rect 3495 2010 3569 2026
rect 3587 2018 3617 2074
rect 3652 2064 3860 2074
rect 3895 2070 3940 2074
rect 3943 2073 3944 2074
rect 3959 2073 3972 2074
rect 3678 2034 3867 2064
rect 3693 2031 3867 2034
rect 3686 2028 3867 2031
rect 3495 2008 3508 2010
rect 3523 2008 3557 2010
rect 3495 1992 3569 2008
rect 3596 2004 3609 2018
rect 3624 2004 3640 2020
rect 3686 2015 3697 2028
rect 3479 1970 3480 1986
rect 3495 1970 3508 1992
rect 3523 1970 3553 1992
rect 3596 1988 3658 2004
rect 3686 1997 3697 2013
rect 3702 2008 3712 2028
rect 3722 2008 3736 2028
rect 3739 2015 3748 2028
rect 3764 2015 3773 2028
rect 3702 1997 3736 2008
rect 3739 1997 3748 2013
rect 3764 1997 3773 2013
rect 3780 2008 3790 2028
rect 3800 2008 3814 2028
rect 3815 2015 3826 2028
rect 3780 1997 3814 2008
rect 3815 1997 3826 2013
rect 3872 2004 3888 2020
rect 3895 2018 3925 2070
rect 3959 2066 3960 2073
rect 3944 2058 3960 2066
rect 3931 2026 3944 2045
rect 3959 2026 3989 2042
rect 3931 2010 4005 2026
rect 3931 2008 3944 2010
rect 3959 2008 3993 2010
rect 3596 1986 3609 1988
rect 3624 1986 3658 1988
rect 3596 1970 3658 1986
rect 3702 1981 3718 1984
rect 3780 1981 3810 1992
rect 3858 1988 3904 2004
rect 3931 1992 4005 2008
rect 3858 1986 3892 1988
rect 3857 1970 3904 1986
rect 3931 1970 3944 1992
rect 3959 1970 3989 1992
rect 4016 1970 4017 1986
rect 4032 1970 4045 2130
rect 4075 2026 4088 2130
rect 4133 2108 4134 2118
rect 4149 2108 4162 2118
rect 4133 2104 4162 2108
rect 4167 2104 4197 2130
rect 4215 2116 4231 2118
rect 4303 2116 4356 2130
rect 4304 2114 4368 2116
rect 4411 2114 4426 2130
rect 4475 2127 4505 2130
rect 4475 2124 4511 2127
rect 4441 2116 4457 2118
rect 4215 2104 4230 2108
rect 4133 2102 4230 2104
rect 4258 2102 4426 2114
rect 4442 2104 4457 2108
rect 4475 2105 4514 2124
rect 4533 2118 4540 2119
rect 4539 2111 4540 2118
rect 4523 2108 4524 2111
rect 4539 2108 4552 2111
rect 4475 2104 4505 2105
rect 4514 2104 4520 2105
rect 4523 2104 4552 2108
rect 4442 2103 4552 2104
rect 4442 2102 4558 2103
rect 4117 2094 4168 2102
rect 4117 2082 4142 2094
rect 4149 2082 4168 2094
rect 4199 2094 4249 2102
rect 4199 2086 4215 2094
rect 4222 2092 4249 2094
rect 4258 2092 4479 2102
rect 4222 2082 4479 2092
rect 4508 2094 4558 2102
rect 4508 2085 4524 2094
rect 4117 2074 4168 2082
rect 4215 2074 4479 2082
rect 4505 2082 4524 2085
rect 4531 2082 4558 2094
rect 4505 2074 4558 2082
rect 4133 2066 4134 2074
rect 4149 2066 4162 2074
rect 4133 2058 4149 2066
rect 4130 2051 4149 2054
rect 4130 2042 4152 2051
rect 4103 2032 4152 2042
rect 4103 2026 4133 2032
rect 4152 2027 4157 2032
rect 4075 2010 4149 2026
rect 4167 2018 4197 2074
rect 4232 2064 4440 2074
rect 4475 2070 4520 2074
rect 4523 2073 4524 2074
rect 4539 2073 4552 2074
rect 4258 2034 4447 2064
rect 4273 2031 4447 2034
rect 4266 2028 4447 2031
rect 4075 2008 4088 2010
rect 4103 2008 4137 2010
rect 4075 1992 4149 2008
rect 4176 2004 4189 2018
rect 4204 2004 4220 2020
rect 4266 2015 4277 2028
rect 4059 1970 4060 1986
rect 4075 1970 4088 1992
rect 4103 1970 4133 1992
rect 4176 1988 4238 2004
rect 4266 1997 4277 2013
rect 4282 2008 4292 2028
rect 4302 2008 4316 2028
rect 4319 2015 4328 2028
rect 4344 2015 4353 2028
rect 4282 1997 4316 2008
rect 4319 1997 4328 2013
rect 4344 1997 4353 2013
rect 4360 2008 4370 2028
rect 4380 2008 4394 2028
rect 4395 2015 4406 2028
rect 4360 1997 4394 2008
rect 4395 1997 4406 2013
rect 4452 2004 4468 2020
rect 4475 2018 4505 2070
rect 4539 2066 4540 2073
rect 4524 2058 4540 2066
rect 4511 2026 4524 2045
rect 4539 2026 4569 2042
rect 4511 2010 4585 2026
rect 4511 2008 4524 2010
rect 4539 2008 4573 2010
rect 4176 1986 4189 1988
rect 4204 1986 4238 1988
rect 4176 1970 4238 1986
rect 4282 1981 4298 1984
rect 4360 1981 4390 1992
rect 4438 1988 4484 2004
rect 4511 1992 4585 2008
rect 4438 1986 4472 1988
rect 4437 1970 4484 1986
rect 4511 1970 4524 1992
rect 4539 1970 4569 1992
rect 4596 1970 4597 1986
rect 4612 1970 4625 2130
rect -7 1962 34 1970
rect -7 1936 8 1962
rect 15 1936 34 1962
rect 98 1958 160 1970
rect 172 1958 247 1970
rect 305 1958 380 1970
rect 392 1958 423 1970
rect 429 1958 464 1970
rect 98 1956 260 1958
rect -7 1928 34 1936
rect 116 1932 129 1956
rect 144 1954 159 1956
rect -1 1918 0 1928
rect 15 1918 28 1928
rect 43 1918 73 1932
rect 116 1918 159 1932
rect 183 1929 190 1936
rect 193 1932 260 1956
rect 292 1956 464 1958
rect 262 1934 290 1938
rect 292 1934 372 1956
rect 393 1954 408 1956
rect 262 1932 372 1934
rect 193 1928 372 1932
rect 166 1918 196 1928
rect 198 1918 351 1928
rect 359 1918 389 1928
rect 393 1918 423 1932
rect 451 1918 464 1956
rect 536 1962 571 1970
rect 536 1936 537 1962
rect 544 1936 571 1962
rect 479 1918 509 1932
rect 536 1928 571 1936
rect 573 1962 614 1970
rect 573 1936 588 1962
rect 595 1936 614 1962
rect 678 1958 740 1970
rect 752 1958 827 1970
rect 885 1958 960 1970
rect 972 1958 1003 1970
rect 1009 1958 1044 1970
rect 678 1956 840 1958
rect 573 1928 614 1936
rect 696 1932 709 1956
rect 724 1954 739 1956
rect 536 1918 537 1928
rect 552 1918 565 1928
rect 579 1918 580 1928
rect 595 1918 608 1928
rect 623 1918 653 1932
rect 696 1918 739 1932
rect 763 1929 770 1936
rect 773 1932 840 1956
rect 872 1956 1044 1958
rect 842 1934 870 1938
rect 872 1934 952 1956
rect 973 1954 988 1956
rect 842 1932 952 1934
rect 773 1928 952 1932
rect 746 1918 776 1928
rect 778 1918 931 1928
rect 939 1918 969 1928
rect 973 1918 1003 1932
rect 1031 1918 1044 1956
rect 1116 1962 1151 1970
rect 1116 1936 1117 1962
rect 1124 1936 1151 1962
rect 1059 1918 1089 1932
rect 1116 1928 1151 1936
rect 1153 1962 1194 1970
rect 1153 1936 1168 1962
rect 1175 1936 1194 1962
rect 1258 1958 1320 1970
rect 1332 1958 1407 1970
rect 1465 1958 1540 1970
rect 1552 1958 1583 1970
rect 1589 1958 1624 1970
rect 1258 1956 1420 1958
rect 1153 1928 1194 1936
rect 1276 1932 1289 1956
rect 1304 1954 1319 1956
rect 1116 1918 1117 1928
rect 1132 1918 1145 1928
rect 1159 1918 1160 1928
rect 1175 1918 1188 1928
rect 1203 1918 1233 1932
rect 1276 1918 1319 1932
rect 1343 1929 1350 1936
rect 1353 1932 1420 1956
rect 1452 1956 1624 1958
rect 1422 1934 1450 1938
rect 1452 1934 1532 1956
rect 1553 1954 1568 1956
rect 1422 1932 1532 1934
rect 1353 1928 1532 1932
rect 1326 1918 1356 1928
rect 1358 1918 1511 1928
rect 1519 1918 1549 1928
rect 1553 1918 1583 1932
rect 1611 1918 1624 1956
rect 1696 1962 1731 1970
rect 1696 1936 1697 1962
rect 1704 1936 1731 1962
rect 1639 1918 1669 1932
rect 1696 1928 1731 1936
rect 1733 1962 1774 1970
rect 1733 1936 1748 1962
rect 1755 1936 1774 1962
rect 1838 1958 1900 1970
rect 1912 1958 1987 1970
rect 2045 1958 2120 1970
rect 2132 1958 2163 1970
rect 2169 1958 2204 1970
rect 1838 1956 2000 1958
rect 1733 1928 1774 1936
rect 1856 1932 1869 1956
rect 1884 1954 1899 1956
rect 1696 1918 1697 1928
rect 1712 1918 1725 1928
rect 1739 1918 1740 1928
rect 1755 1918 1768 1928
rect 1783 1918 1813 1932
rect 1856 1918 1899 1932
rect 1923 1929 1930 1936
rect 1933 1932 2000 1956
rect 2032 1956 2204 1958
rect 2002 1934 2030 1938
rect 2032 1934 2112 1956
rect 2133 1954 2148 1956
rect 2002 1932 2112 1934
rect 1933 1928 2112 1932
rect 1906 1918 1936 1928
rect 1938 1918 2091 1928
rect 2099 1918 2129 1928
rect 2133 1918 2163 1932
rect 2191 1918 2204 1956
rect 2276 1962 2311 1970
rect 2276 1936 2277 1962
rect 2284 1936 2311 1962
rect 2219 1918 2249 1932
rect 2276 1928 2311 1936
rect 2313 1962 2354 1970
rect 2313 1936 2328 1962
rect 2335 1936 2354 1962
rect 2418 1958 2480 1970
rect 2492 1958 2567 1970
rect 2625 1958 2700 1970
rect 2712 1958 2743 1970
rect 2749 1958 2784 1970
rect 2418 1956 2580 1958
rect 2313 1928 2354 1936
rect 2436 1932 2449 1956
rect 2464 1954 2479 1956
rect 2276 1918 2277 1928
rect 2292 1918 2305 1928
rect 2319 1918 2320 1928
rect 2335 1918 2348 1928
rect 2363 1918 2393 1932
rect 2436 1918 2479 1932
rect 2503 1929 2510 1936
rect 2513 1932 2580 1956
rect 2612 1956 2784 1958
rect 2582 1934 2610 1938
rect 2612 1934 2692 1956
rect 2713 1954 2728 1956
rect 2582 1932 2692 1934
rect 2513 1928 2692 1932
rect 2486 1918 2516 1928
rect 2518 1918 2671 1928
rect 2679 1918 2709 1928
rect 2713 1918 2743 1932
rect 2771 1918 2784 1956
rect 2856 1962 2891 1970
rect 2856 1936 2857 1962
rect 2864 1936 2891 1962
rect 2799 1918 2829 1932
rect 2856 1928 2891 1936
rect 2893 1962 2934 1970
rect 2893 1936 2908 1962
rect 2915 1936 2934 1962
rect 2998 1958 3060 1970
rect 3072 1958 3147 1970
rect 3205 1958 3280 1970
rect 3292 1958 3323 1970
rect 3329 1958 3364 1970
rect 2998 1956 3160 1958
rect 2893 1928 2934 1936
rect 3016 1932 3029 1956
rect 3044 1954 3059 1956
rect 2856 1918 2857 1928
rect 2872 1918 2885 1928
rect 2899 1918 2900 1928
rect 2915 1918 2928 1928
rect 2943 1918 2973 1932
rect 3016 1918 3059 1932
rect 3083 1929 3090 1936
rect 3093 1932 3160 1956
rect 3192 1956 3364 1958
rect 3162 1934 3190 1938
rect 3192 1934 3272 1956
rect 3293 1954 3308 1956
rect 3162 1932 3272 1934
rect 3093 1928 3272 1932
rect 3066 1918 3096 1928
rect 3098 1918 3251 1928
rect 3259 1918 3289 1928
rect 3293 1918 3323 1932
rect 3351 1918 3364 1956
rect 3436 1962 3471 1970
rect 3436 1936 3437 1962
rect 3444 1936 3471 1962
rect 3379 1918 3409 1932
rect 3436 1928 3471 1936
rect 3473 1962 3514 1970
rect 3473 1936 3488 1962
rect 3495 1936 3514 1962
rect 3578 1958 3640 1970
rect 3652 1958 3727 1970
rect 3785 1958 3860 1970
rect 3872 1958 3903 1970
rect 3909 1958 3944 1970
rect 3578 1956 3740 1958
rect 3473 1928 3514 1936
rect 3596 1932 3609 1956
rect 3624 1954 3639 1956
rect 3436 1918 3437 1928
rect 3452 1918 3465 1928
rect 3479 1918 3480 1928
rect 3495 1918 3508 1928
rect 3523 1918 3553 1932
rect 3596 1918 3639 1932
rect 3663 1929 3670 1936
rect 3673 1932 3740 1956
rect 3772 1956 3944 1958
rect 3742 1934 3770 1938
rect 3772 1934 3852 1956
rect 3873 1954 3888 1956
rect 3742 1932 3852 1934
rect 3673 1928 3852 1932
rect 3646 1918 3676 1928
rect 3678 1918 3831 1928
rect 3839 1918 3869 1928
rect 3873 1918 3903 1932
rect 3931 1918 3944 1956
rect 4016 1962 4051 1970
rect 4016 1936 4017 1962
rect 4024 1936 4051 1962
rect 3959 1918 3989 1932
rect 4016 1928 4051 1936
rect 4053 1962 4094 1970
rect 4053 1936 4068 1962
rect 4075 1936 4094 1962
rect 4158 1958 4220 1970
rect 4232 1958 4307 1970
rect 4365 1958 4440 1970
rect 4452 1958 4483 1970
rect 4489 1958 4524 1970
rect 4158 1956 4320 1958
rect 4053 1928 4094 1936
rect 4176 1932 4189 1956
rect 4204 1954 4219 1956
rect 4016 1918 4017 1928
rect 4032 1918 4045 1928
rect 4059 1918 4060 1928
rect 4075 1918 4088 1928
rect 4103 1918 4133 1932
rect 4176 1918 4219 1932
rect 4243 1929 4250 1936
rect 4253 1932 4320 1956
rect 4352 1956 4524 1958
rect 4322 1934 4350 1938
rect 4352 1934 4432 1956
rect 4453 1954 4468 1956
rect 4322 1932 4432 1934
rect 4253 1928 4432 1932
rect 4226 1918 4256 1928
rect 4258 1918 4411 1928
rect 4419 1918 4449 1928
rect 4453 1918 4483 1932
rect 4511 1918 4524 1956
rect 4596 1962 4631 1970
rect 4596 1936 4597 1962
rect 4604 1936 4631 1962
rect 4539 1918 4569 1932
rect 4596 1928 4631 1936
rect 4596 1918 4597 1928
rect 4612 1918 4625 1928
rect -1 1912 4625 1918
rect 0 1904 4625 1912
rect 15 1874 28 1904
rect 43 1886 73 1904
rect 116 1890 130 1904
rect 166 1890 386 1904
rect 117 1888 130 1890
rect 83 1876 98 1888
rect 80 1874 102 1876
rect 107 1874 137 1888
rect 198 1886 351 1890
rect 180 1874 372 1886
rect 415 1874 445 1888
rect 451 1874 464 1904
rect 479 1886 509 1904
rect 552 1874 565 1904
rect 595 1874 608 1904
rect 623 1886 653 1904
rect 696 1890 710 1904
rect 746 1890 966 1904
rect 697 1888 710 1890
rect 663 1876 678 1888
rect 660 1874 682 1876
rect 687 1874 717 1888
rect 778 1886 931 1890
rect 760 1874 952 1886
rect 995 1874 1025 1888
rect 1031 1874 1044 1904
rect 1059 1886 1089 1904
rect 1132 1874 1145 1904
rect 1175 1874 1188 1904
rect 1203 1886 1233 1904
rect 1276 1890 1290 1904
rect 1326 1890 1546 1904
rect 1277 1888 1290 1890
rect 1243 1876 1258 1888
rect 1240 1874 1262 1876
rect 1267 1874 1297 1888
rect 1358 1886 1511 1890
rect 1340 1874 1532 1886
rect 1575 1874 1605 1888
rect 1611 1874 1624 1904
rect 1639 1886 1669 1904
rect 1712 1874 1725 1904
rect 1755 1874 1768 1904
rect 1783 1886 1813 1904
rect 1856 1890 1870 1904
rect 1906 1890 2126 1904
rect 1857 1888 1870 1890
rect 1823 1876 1838 1888
rect 1820 1874 1842 1876
rect 1847 1874 1877 1888
rect 1938 1886 2091 1890
rect 1920 1874 2112 1886
rect 2155 1874 2185 1888
rect 2191 1874 2204 1904
rect 2219 1886 2249 1904
rect 2292 1874 2305 1904
rect 2335 1874 2348 1904
rect 2363 1886 2393 1904
rect 2436 1890 2450 1904
rect 2486 1890 2706 1904
rect 2437 1888 2450 1890
rect 2403 1876 2418 1888
rect 2400 1874 2422 1876
rect 2427 1874 2457 1888
rect 2518 1886 2671 1890
rect 2500 1874 2692 1886
rect 2735 1874 2765 1888
rect 2771 1874 2784 1904
rect 2799 1886 2829 1904
rect 2872 1874 2885 1904
rect 2915 1874 2928 1904
rect 2943 1886 2973 1904
rect 3016 1890 3030 1904
rect 3066 1890 3286 1904
rect 3017 1888 3030 1890
rect 2983 1876 2998 1888
rect 2980 1874 3002 1876
rect 3007 1874 3037 1888
rect 3098 1886 3251 1890
rect 3080 1874 3272 1886
rect 3315 1874 3345 1888
rect 3351 1874 3364 1904
rect 3379 1886 3409 1904
rect 3452 1874 3465 1904
rect 3495 1874 3508 1904
rect 3523 1886 3553 1904
rect 3596 1890 3610 1904
rect 3646 1890 3866 1904
rect 3597 1888 3610 1890
rect 3563 1876 3578 1888
rect 3560 1874 3582 1876
rect 3587 1874 3617 1888
rect 3678 1886 3831 1890
rect 3660 1874 3852 1886
rect 3895 1874 3925 1888
rect 3931 1874 3944 1904
rect 3959 1886 3989 1904
rect 4032 1874 4045 1904
rect 4075 1874 4088 1904
rect 4103 1886 4133 1904
rect 4176 1890 4190 1904
rect 4226 1890 4446 1904
rect 4177 1888 4190 1890
rect 4143 1876 4158 1888
rect 4140 1874 4162 1876
rect 4167 1874 4197 1888
rect 4258 1886 4411 1890
rect 4240 1874 4432 1886
rect 4475 1874 4505 1888
rect 4511 1874 4524 1904
rect 4539 1886 4569 1904
rect 4612 1874 4625 1904
rect 0 1860 4625 1874
rect 15 1756 28 1860
rect 73 1838 74 1848
rect 89 1838 102 1848
rect 73 1834 102 1838
rect 107 1834 137 1860
rect 155 1846 171 1848
rect 243 1846 296 1860
rect 244 1844 308 1846
rect 351 1844 366 1860
rect 415 1857 445 1860
rect 415 1854 451 1857
rect 381 1846 397 1848
rect 155 1834 170 1838
rect 73 1832 170 1834
rect 198 1832 366 1844
rect 382 1834 397 1838
rect 415 1835 454 1854
rect 473 1848 480 1849
rect 479 1841 480 1848
rect 463 1838 464 1841
rect 479 1838 492 1841
rect 415 1834 445 1835
rect 454 1834 460 1835
rect 463 1834 492 1838
rect 382 1833 492 1834
rect 382 1832 498 1833
rect 57 1824 108 1832
rect 57 1812 82 1824
rect 89 1812 108 1824
rect 139 1824 189 1832
rect 139 1816 155 1824
rect 162 1822 189 1824
rect 198 1822 419 1832
rect 162 1812 419 1822
rect 448 1824 498 1832
rect 448 1815 464 1824
rect 57 1804 108 1812
rect 155 1804 419 1812
rect 445 1812 464 1815
rect 471 1812 498 1824
rect 445 1804 498 1812
rect 73 1796 74 1804
rect 89 1796 102 1804
rect 73 1788 89 1796
rect 70 1781 89 1784
rect 70 1772 92 1781
rect 43 1762 92 1772
rect 43 1756 73 1762
rect 92 1757 97 1762
rect 15 1740 89 1756
rect 107 1748 137 1804
rect 172 1794 380 1804
rect 415 1800 460 1804
rect 463 1803 464 1804
rect 479 1803 492 1804
rect 198 1764 387 1794
rect 213 1761 387 1764
rect 206 1758 387 1761
rect 15 1738 28 1740
rect 43 1738 77 1740
rect 15 1722 89 1738
rect 116 1734 129 1748
rect 144 1734 160 1750
rect 206 1745 217 1758
rect -1 1700 0 1716
rect 15 1700 28 1722
rect 43 1700 73 1722
rect 116 1718 178 1734
rect 206 1727 217 1743
rect 222 1738 232 1758
rect 242 1738 256 1758
rect 259 1745 268 1758
rect 284 1745 293 1758
rect 222 1727 256 1738
rect 259 1727 268 1743
rect 284 1727 293 1743
rect 300 1738 310 1758
rect 320 1738 334 1758
rect 335 1745 346 1758
rect 300 1727 334 1738
rect 335 1727 346 1743
rect 392 1734 408 1750
rect 415 1748 445 1800
rect 479 1796 480 1803
rect 464 1788 480 1796
rect 451 1756 464 1775
rect 479 1756 509 1772
rect 451 1740 525 1756
rect 451 1738 464 1740
rect 479 1738 513 1740
rect 116 1716 129 1718
rect 144 1716 178 1718
rect 116 1700 178 1716
rect 222 1711 238 1714
rect 300 1711 330 1722
rect 378 1718 424 1734
rect 451 1722 525 1738
rect 378 1716 412 1718
rect 377 1700 424 1716
rect 451 1700 464 1722
rect 479 1700 509 1722
rect 536 1700 537 1716
rect 552 1700 565 1860
rect 595 1756 608 1860
rect 653 1838 654 1848
rect 669 1838 682 1848
rect 653 1834 682 1838
rect 687 1834 717 1860
rect 735 1846 751 1848
rect 823 1846 876 1860
rect 824 1844 888 1846
rect 931 1844 946 1860
rect 995 1857 1025 1860
rect 995 1854 1031 1857
rect 961 1846 977 1848
rect 735 1834 750 1838
rect 653 1832 750 1834
rect 778 1832 946 1844
rect 962 1834 977 1838
rect 995 1835 1034 1854
rect 1053 1848 1060 1849
rect 1059 1841 1060 1848
rect 1043 1838 1044 1841
rect 1059 1838 1072 1841
rect 995 1834 1025 1835
rect 1034 1834 1040 1835
rect 1043 1834 1072 1838
rect 962 1833 1072 1834
rect 962 1832 1078 1833
rect 637 1824 688 1832
rect 637 1812 662 1824
rect 669 1812 688 1824
rect 719 1824 769 1832
rect 719 1816 735 1824
rect 742 1822 769 1824
rect 778 1822 999 1832
rect 742 1812 999 1822
rect 1028 1824 1078 1832
rect 1028 1815 1044 1824
rect 637 1804 688 1812
rect 735 1804 999 1812
rect 1025 1812 1044 1815
rect 1051 1812 1078 1824
rect 1025 1804 1078 1812
rect 653 1796 654 1804
rect 669 1796 682 1804
rect 653 1788 669 1796
rect 650 1781 669 1784
rect 650 1772 672 1781
rect 623 1762 672 1772
rect 623 1756 653 1762
rect 672 1757 677 1762
rect 595 1740 669 1756
rect 687 1748 717 1804
rect 752 1794 960 1804
rect 995 1800 1040 1804
rect 1043 1803 1044 1804
rect 1059 1803 1072 1804
rect 778 1764 967 1794
rect 793 1761 967 1764
rect 786 1758 967 1761
rect 595 1738 608 1740
rect 623 1738 657 1740
rect 595 1722 669 1738
rect 696 1734 709 1748
rect 724 1734 740 1750
rect 786 1745 797 1758
rect 579 1700 580 1716
rect 595 1700 608 1722
rect 623 1700 653 1722
rect 696 1718 758 1734
rect 786 1727 797 1743
rect 802 1738 812 1758
rect 822 1738 836 1758
rect 839 1745 848 1758
rect 864 1745 873 1758
rect 802 1727 836 1738
rect 839 1727 848 1743
rect 864 1727 873 1743
rect 880 1738 890 1758
rect 900 1738 914 1758
rect 915 1745 926 1758
rect 880 1727 914 1738
rect 915 1727 926 1743
rect 972 1734 988 1750
rect 995 1748 1025 1800
rect 1059 1796 1060 1803
rect 1044 1788 1060 1796
rect 1031 1756 1044 1775
rect 1059 1756 1089 1772
rect 1031 1740 1105 1756
rect 1031 1738 1044 1740
rect 1059 1738 1093 1740
rect 696 1716 709 1718
rect 724 1716 758 1718
rect 696 1700 758 1716
rect 802 1711 818 1714
rect 880 1711 910 1722
rect 958 1718 1004 1734
rect 1031 1722 1105 1738
rect 958 1716 992 1718
rect 957 1700 1004 1716
rect 1031 1700 1044 1722
rect 1059 1700 1089 1722
rect 1116 1700 1117 1716
rect 1132 1700 1145 1860
rect 1175 1756 1188 1860
rect 1233 1838 1234 1848
rect 1249 1838 1262 1848
rect 1233 1834 1262 1838
rect 1267 1834 1297 1860
rect 1315 1846 1331 1848
rect 1403 1846 1456 1860
rect 1404 1844 1468 1846
rect 1511 1844 1526 1860
rect 1575 1857 1605 1860
rect 1575 1854 1611 1857
rect 1541 1846 1557 1848
rect 1315 1834 1330 1838
rect 1233 1832 1330 1834
rect 1358 1832 1526 1844
rect 1542 1834 1557 1838
rect 1575 1835 1614 1854
rect 1633 1848 1640 1849
rect 1639 1841 1640 1848
rect 1623 1838 1624 1841
rect 1639 1838 1652 1841
rect 1575 1834 1605 1835
rect 1614 1834 1620 1835
rect 1623 1834 1652 1838
rect 1542 1833 1652 1834
rect 1542 1832 1658 1833
rect 1217 1824 1268 1832
rect 1217 1812 1242 1824
rect 1249 1812 1268 1824
rect 1299 1824 1349 1832
rect 1299 1816 1315 1824
rect 1322 1822 1349 1824
rect 1358 1822 1579 1832
rect 1322 1812 1579 1822
rect 1608 1824 1658 1832
rect 1608 1815 1624 1824
rect 1217 1804 1268 1812
rect 1315 1804 1579 1812
rect 1605 1812 1624 1815
rect 1631 1812 1658 1824
rect 1605 1804 1658 1812
rect 1233 1796 1234 1804
rect 1249 1796 1262 1804
rect 1233 1788 1249 1796
rect 1230 1781 1249 1784
rect 1230 1772 1252 1781
rect 1203 1762 1252 1772
rect 1203 1756 1233 1762
rect 1252 1757 1257 1762
rect 1175 1740 1249 1756
rect 1267 1748 1297 1804
rect 1332 1794 1540 1804
rect 1575 1800 1620 1804
rect 1623 1803 1624 1804
rect 1639 1803 1652 1804
rect 1358 1764 1547 1794
rect 1373 1761 1547 1764
rect 1366 1758 1547 1761
rect 1175 1738 1188 1740
rect 1203 1738 1237 1740
rect 1175 1722 1249 1738
rect 1276 1734 1289 1748
rect 1304 1734 1320 1750
rect 1366 1745 1377 1758
rect 1159 1700 1160 1716
rect 1175 1700 1188 1722
rect 1203 1700 1233 1722
rect 1276 1718 1338 1734
rect 1366 1727 1377 1743
rect 1382 1738 1392 1758
rect 1402 1738 1416 1758
rect 1419 1745 1428 1758
rect 1444 1745 1453 1758
rect 1382 1727 1416 1738
rect 1419 1727 1428 1743
rect 1444 1727 1453 1743
rect 1460 1738 1470 1758
rect 1480 1738 1494 1758
rect 1495 1745 1506 1758
rect 1460 1727 1494 1738
rect 1495 1727 1506 1743
rect 1552 1734 1568 1750
rect 1575 1748 1605 1800
rect 1639 1796 1640 1803
rect 1624 1788 1640 1796
rect 1611 1756 1624 1775
rect 1639 1756 1669 1772
rect 1611 1740 1685 1756
rect 1611 1738 1624 1740
rect 1639 1738 1673 1740
rect 1276 1716 1289 1718
rect 1304 1716 1338 1718
rect 1276 1700 1338 1716
rect 1382 1711 1398 1714
rect 1460 1711 1490 1722
rect 1538 1718 1584 1734
rect 1611 1722 1685 1738
rect 1538 1716 1572 1718
rect 1537 1700 1584 1716
rect 1611 1700 1624 1722
rect 1639 1700 1669 1722
rect 1696 1700 1697 1716
rect 1712 1700 1725 1860
rect 1755 1756 1768 1860
rect 1813 1838 1814 1848
rect 1829 1838 1842 1848
rect 1813 1834 1842 1838
rect 1847 1834 1877 1860
rect 1895 1846 1911 1848
rect 1983 1846 2036 1860
rect 1984 1844 2048 1846
rect 2091 1844 2106 1860
rect 2155 1857 2185 1860
rect 2155 1854 2191 1857
rect 2121 1846 2137 1848
rect 1895 1834 1910 1838
rect 1813 1832 1910 1834
rect 1938 1832 2106 1844
rect 2122 1834 2137 1838
rect 2155 1835 2194 1854
rect 2213 1848 2220 1849
rect 2219 1841 2220 1848
rect 2203 1838 2204 1841
rect 2219 1838 2232 1841
rect 2155 1834 2185 1835
rect 2194 1834 2200 1835
rect 2203 1834 2232 1838
rect 2122 1833 2232 1834
rect 2122 1832 2238 1833
rect 1797 1824 1848 1832
rect 1797 1812 1822 1824
rect 1829 1812 1848 1824
rect 1879 1824 1929 1832
rect 1879 1816 1895 1824
rect 1902 1822 1929 1824
rect 1938 1822 2159 1832
rect 1902 1812 2159 1822
rect 2188 1824 2238 1832
rect 2188 1815 2204 1824
rect 1797 1804 1848 1812
rect 1895 1804 2159 1812
rect 2185 1812 2204 1815
rect 2211 1812 2238 1824
rect 2185 1804 2238 1812
rect 1813 1796 1814 1804
rect 1829 1796 1842 1804
rect 1813 1788 1829 1796
rect 1810 1781 1829 1784
rect 1810 1772 1832 1781
rect 1783 1762 1832 1772
rect 1783 1756 1813 1762
rect 1832 1757 1837 1762
rect 1755 1740 1829 1756
rect 1847 1748 1877 1804
rect 1912 1794 2120 1804
rect 2155 1800 2200 1804
rect 2203 1803 2204 1804
rect 2219 1803 2232 1804
rect 1938 1764 2127 1794
rect 1953 1761 2127 1764
rect 1946 1758 2127 1761
rect 1755 1738 1768 1740
rect 1783 1738 1817 1740
rect 1755 1722 1829 1738
rect 1856 1734 1869 1748
rect 1884 1734 1900 1750
rect 1946 1745 1957 1758
rect 1739 1700 1740 1716
rect 1755 1700 1768 1722
rect 1783 1700 1813 1722
rect 1856 1718 1918 1734
rect 1946 1727 1957 1743
rect 1962 1738 1972 1758
rect 1982 1738 1996 1758
rect 1999 1745 2008 1758
rect 2024 1745 2033 1758
rect 1962 1727 1996 1738
rect 1999 1727 2008 1743
rect 2024 1727 2033 1743
rect 2040 1738 2050 1758
rect 2060 1738 2074 1758
rect 2075 1745 2086 1758
rect 2040 1727 2074 1738
rect 2075 1727 2086 1743
rect 2132 1734 2148 1750
rect 2155 1748 2185 1800
rect 2219 1796 2220 1803
rect 2204 1788 2220 1796
rect 2191 1756 2204 1775
rect 2219 1756 2249 1772
rect 2191 1740 2265 1756
rect 2191 1738 2204 1740
rect 2219 1738 2253 1740
rect 1856 1716 1869 1718
rect 1884 1716 1918 1718
rect 1856 1700 1918 1716
rect 1962 1711 1978 1714
rect 2040 1711 2070 1722
rect 2118 1718 2164 1734
rect 2191 1722 2265 1738
rect 2118 1716 2152 1718
rect 2117 1700 2164 1716
rect 2191 1700 2204 1722
rect 2219 1700 2249 1722
rect 2276 1700 2277 1716
rect 2292 1700 2305 1860
rect 2335 1756 2348 1860
rect 2393 1838 2394 1848
rect 2409 1838 2422 1848
rect 2393 1834 2422 1838
rect 2427 1834 2457 1860
rect 2475 1846 2491 1848
rect 2563 1846 2616 1860
rect 2564 1844 2628 1846
rect 2671 1844 2686 1860
rect 2735 1857 2765 1860
rect 2735 1854 2771 1857
rect 2701 1846 2717 1848
rect 2475 1834 2490 1838
rect 2393 1832 2490 1834
rect 2518 1832 2686 1844
rect 2702 1834 2717 1838
rect 2735 1835 2774 1854
rect 2793 1848 2800 1849
rect 2799 1841 2800 1848
rect 2783 1838 2784 1841
rect 2799 1838 2812 1841
rect 2735 1834 2765 1835
rect 2774 1834 2780 1835
rect 2783 1834 2812 1838
rect 2702 1833 2812 1834
rect 2702 1832 2818 1833
rect 2377 1824 2428 1832
rect 2377 1812 2402 1824
rect 2409 1812 2428 1824
rect 2459 1824 2509 1832
rect 2459 1816 2475 1824
rect 2482 1822 2509 1824
rect 2518 1822 2739 1832
rect 2482 1812 2739 1822
rect 2768 1824 2818 1832
rect 2768 1815 2784 1824
rect 2377 1804 2428 1812
rect 2475 1804 2739 1812
rect 2765 1812 2784 1815
rect 2791 1812 2818 1824
rect 2765 1804 2818 1812
rect 2393 1796 2394 1804
rect 2409 1796 2422 1804
rect 2393 1788 2409 1796
rect 2390 1781 2409 1784
rect 2390 1772 2412 1781
rect 2363 1762 2412 1772
rect 2363 1756 2393 1762
rect 2412 1757 2417 1762
rect 2335 1740 2409 1756
rect 2427 1748 2457 1804
rect 2492 1794 2700 1804
rect 2735 1800 2780 1804
rect 2783 1803 2784 1804
rect 2799 1803 2812 1804
rect 2518 1764 2707 1794
rect 2533 1761 2707 1764
rect 2526 1758 2707 1761
rect 2335 1738 2348 1740
rect 2363 1738 2397 1740
rect 2335 1722 2409 1738
rect 2436 1734 2449 1748
rect 2464 1734 2480 1750
rect 2526 1745 2537 1758
rect 2319 1700 2320 1716
rect 2335 1700 2348 1722
rect 2363 1700 2393 1722
rect 2436 1718 2498 1734
rect 2526 1727 2537 1743
rect 2542 1738 2552 1758
rect 2562 1738 2576 1758
rect 2579 1745 2588 1758
rect 2604 1745 2613 1758
rect 2542 1727 2576 1738
rect 2579 1727 2588 1743
rect 2604 1727 2613 1743
rect 2620 1738 2630 1758
rect 2640 1738 2654 1758
rect 2655 1745 2666 1758
rect 2620 1727 2654 1738
rect 2655 1727 2666 1743
rect 2712 1734 2728 1750
rect 2735 1748 2765 1800
rect 2799 1796 2800 1803
rect 2784 1788 2800 1796
rect 2771 1756 2784 1775
rect 2799 1756 2829 1772
rect 2771 1740 2845 1756
rect 2771 1738 2784 1740
rect 2799 1738 2833 1740
rect 2436 1716 2449 1718
rect 2464 1716 2498 1718
rect 2436 1700 2498 1716
rect 2542 1711 2558 1714
rect 2620 1711 2650 1722
rect 2698 1718 2744 1734
rect 2771 1722 2845 1738
rect 2698 1716 2732 1718
rect 2697 1700 2744 1716
rect 2771 1700 2784 1722
rect 2799 1700 2829 1722
rect 2856 1700 2857 1716
rect 2872 1700 2885 1860
rect 2915 1756 2928 1860
rect 2973 1838 2974 1848
rect 2989 1838 3002 1848
rect 2973 1834 3002 1838
rect 3007 1834 3037 1860
rect 3055 1846 3071 1848
rect 3143 1846 3196 1860
rect 3144 1844 3208 1846
rect 3251 1844 3266 1860
rect 3315 1857 3345 1860
rect 3315 1854 3351 1857
rect 3281 1846 3297 1848
rect 3055 1834 3070 1838
rect 2973 1832 3070 1834
rect 3098 1832 3266 1844
rect 3282 1834 3297 1838
rect 3315 1835 3354 1854
rect 3373 1848 3380 1849
rect 3379 1841 3380 1848
rect 3363 1838 3364 1841
rect 3379 1838 3392 1841
rect 3315 1834 3345 1835
rect 3354 1834 3360 1835
rect 3363 1834 3392 1838
rect 3282 1833 3392 1834
rect 3282 1832 3398 1833
rect 2957 1824 3008 1832
rect 2957 1812 2982 1824
rect 2989 1812 3008 1824
rect 3039 1824 3089 1832
rect 3039 1816 3055 1824
rect 3062 1822 3089 1824
rect 3098 1822 3319 1832
rect 3062 1812 3319 1822
rect 3348 1824 3398 1832
rect 3348 1815 3364 1824
rect 2957 1804 3008 1812
rect 3055 1804 3319 1812
rect 3345 1812 3364 1815
rect 3371 1812 3398 1824
rect 3345 1804 3398 1812
rect 2973 1796 2974 1804
rect 2989 1796 3002 1804
rect 2973 1788 2989 1796
rect 2970 1781 2989 1784
rect 2970 1772 2992 1781
rect 2943 1762 2992 1772
rect 2943 1756 2973 1762
rect 2992 1757 2997 1762
rect 2915 1740 2989 1756
rect 3007 1748 3037 1804
rect 3072 1794 3280 1804
rect 3315 1800 3360 1804
rect 3363 1803 3364 1804
rect 3379 1803 3392 1804
rect 3098 1764 3287 1794
rect 3113 1761 3287 1764
rect 3106 1758 3287 1761
rect 2915 1738 2928 1740
rect 2943 1738 2977 1740
rect 2915 1722 2989 1738
rect 3016 1734 3029 1748
rect 3044 1734 3060 1750
rect 3106 1745 3117 1758
rect 2899 1700 2900 1716
rect 2915 1700 2928 1722
rect 2943 1700 2973 1722
rect 3016 1718 3078 1734
rect 3106 1727 3117 1743
rect 3122 1738 3132 1758
rect 3142 1738 3156 1758
rect 3159 1745 3168 1758
rect 3184 1745 3193 1758
rect 3122 1727 3156 1738
rect 3159 1727 3168 1743
rect 3184 1727 3193 1743
rect 3200 1738 3210 1758
rect 3220 1738 3234 1758
rect 3235 1745 3246 1758
rect 3200 1727 3234 1738
rect 3235 1727 3246 1743
rect 3292 1734 3308 1750
rect 3315 1748 3345 1800
rect 3379 1796 3380 1803
rect 3364 1788 3380 1796
rect 3351 1756 3364 1775
rect 3379 1756 3409 1772
rect 3351 1740 3425 1756
rect 3351 1738 3364 1740
rect 3379 1738 3413 1740
rect 3016 1716 3029 1718
rect 3044 1716 3078 1718
rect 3016 1700 3078 1716
rect 3122 1711 3138 1714
rect 3200 1711 3230 1722
rect 3278 1718 3324 1734
rect 3351 1722 3425 1738
rect 3278 1716 3312 1718
rect 3277 1700 3324 1716
rect 3351 1700 3364 1722
rect 3379 1700 3409 1722
rect 3436 1700 3437 1716
rect 3452 1700 3465 1860
rect 3495 1756 3508 1860
rect 3553 1838 3554 1848
rect 3569 1838 3582 1848
rect 3553 1834 3582 1838
rect 3587 1834 3617 1860
rect 3635 1846 3651 1848
rect 3723 1846 3776 1860
rect 3724 1844 3788 1846
rect 3831 1844 3846 1860
rect 3895 1857 3925 1860
rect 3895 1854 3931 1857
rect 3861 1846 3877 1848
rect 3635 1834 3650 1838
rect 3553 1832 3650 1834
rect 3678 1832 3846 1844
rect 3862 1834 3877 1838
rect 3895 1835 3934 1854
rect 3953 1848 3960 1849
rect 3959 1841 3960 1848
rect 3943 1838 3944 1841
rect 3959 1838 3972 1841
rect 3895 1834 3925 1835
rect 3934 1834 3940 1835
rect 3943 1834 3972 1838
rect 3862 1833 3972 1834
rect 3862 1832 3978 1833
rect 3537 1824 3588 1832
rect 3537 1812 3562 1824
rect 3569 1812 3588 1824
rect 3619 1824 3669 1832
rect 3619 1816 3635 1824
rect 3642 1822 3669 1824
rect 3678 1822 3899 1832
rect 3642 1812 3899 1822
rect 3928 1824 3978 1832
rect 3928 1815 3944 1824
rect 3537 1804 3588 1812
rect 3635 1804 3899 1812
rect 3925 1812 3944 1815
rect 3951 1812 3978 1824
rect 3925 1804 3978 1812
rect 3553 1796 3554 1804
rect 3569 1796 3582 1804
rect 3553 1788 3569 1796
rect 3550 1781 3569 1784
rect 3550 1772 3572 1781
rect 3523 1762 3572 1772
rect 3523 1756 3553 1762
rect 3572 1757 3577 1762
rect 3495 1740 3569 1756
rect 3587 1748 3617 1804
rect 3652 1794 3860 1804
rect 3895 1800 3940 1804
rect 3943 1803 3944 1804
rect 3959 1803 3972 1804
rect 3678 1764 3867 1794
rect 3693 1761 3867 1764
rect 3686 1758 3867 1761
rect 3495 1738 3508 1740
rect 3523 1738 3557 1740
rect 3495 1722 3569 1738
rect 3596 1734 3609 1748
rect 3624 1734 3640 1750
rect 3686 1745 3697 1758
rect 3479 1700 3480 1716
rect 3495 1700 3508 1722
rect 3523 1700 3553 1722
rect 3596 1718 3658 1734
rect 3686 1727 3697 1743
rect 3702 1738 3712 1758
rect 3722 1738 3736 1758
rect 3739 1745 3748 1758
rect 3764 1745 3773 1758
rect 3702 1727 3736 1738
rect 3739 1727 3748 1743
rect 3764 1727 3773 1743
rect 3780 1738 3790 1758
rect 3800 1738 3814 1758
rect 3815 1745 3826 1758
rect 3780 1727 3814 1738
rect 3815 1727 3826 1743
rect 3872 1734 3888 1750
rect 3895 1748 3925 1800
rect 3959 1796 3960 1803
rect 3944 1788 3960 1796
rect 3931 1756 3944 1775
rect 3959 1756 3989 1772
rect 3931 1740 4005 1756
rect 3931 1738 3944 1740
rect 3959 1738 3993 1740
rect 3596 1716 3609 1718
rect 3624 1716 3658 1718
rect 3596 1700 3658 1716
rect 3702 1711 3718 1714
rect 3780 1711 3810 1722
rect 3858 1718 3904 1734
rect 3931 1722 4005 1738
rect 3858 1716 3892 1718
rect 3857 1700 3904 1716
rect 3931 1700 3944 1722
rect 3959 1700 3989 1722
rect 4016 1700 4017 1716
rect 4032 1700 4045 1860
rect 4075 1756 4088 1860
rect 4133 1838 4134 1848
rect 4149 1838 4162 1848
rect 4133 1834 4162 1838
rect 4167 1834 4197 1860
rect 4215 1846 4231 1848
rect 4303 1846 4356 1860
rect 4304 1844 4368 1846
rect 4411 1844 4426 1860
rect 4475 1857 4505 1860
rect 4475 1854 4511 1857
rect 4441 1846 4457 1848
rect 4215 1834 4230 1838
rect 4133 1832 4230 1834
rect 4258 1832 4426 1844
rect 4442 1834 4457 1838
rect 4475 1835 4514 1854
rect 4533 1848 4540 1849
rect 4539 1841 4540 1848
rect 4523 1838 4524 1841
rect 4539 1838 4552 1841
rect 4475 1834 4505 1835
rect 4514 1834 4520 1835
rect 4523 1834 4552 1838
rect 4442 1833 4552 1834
rect 4442 1832 4558 1833
rect 4117 1824 4168 1832
rect 4117 1812 4142 1824
rect 4149 1812 4168 1824
rect 4199 1824 4249 1832
rect 4199 1816 4215 1824
rect 4222 1822 4249 1824
rect 4258 1822 4479 1832
rect 4222 1812 4479 1822
rect 4508 1824 4558 1832
rect 4508 1815 4524 1824
rect 4117 1804 4168 1812
rect 4215 1804 4479 1812
rect 4505 1812 4524 1815
rect 4531 1812 4558 1824
rect 4505 1804 4558 1812
rect 4133 1796 4134 1804
rect 4149 1796 4162 1804
rect 4133 1788 4149 1796
rect 4130 1781 4149 1784
rect 4130 1772 4152 1781
rect 4103 1762 4152 1772
rect 4103 1756 4133 1762
rect 4152 1757 4157 1762
rect 4075 1740 4149 1756
rect 4167 1748 4197 1804
rect 4232 1794 4440 1804
rect 4475 1800 4520 1804
rect 4523 1803 4524 1804
rect 4539 1803 4552 1804
rect 4258 1764 4447 1794
rect 4273 1761 4447 1764
rect 4266 1758 4447 1761
rect 4075 1738 4088 1740
rect 4103 1738 4137 1740
rect 4075 1722 4149 1738
rect 4176 1734 4189 1748
rect 4204 1734 4220 1750
rect 4266 1745 4277 1758
rect 4059 1700 4060 1716
rect 4075 1700 4088 1722
rect 4103 1700 4133 1722
rect 4176 1718 4238 1734
rect 4266 1727 4277 1743
rect 4282 1738 4292 1758
rect 4302 1738 4316 1758
rect 4319 1745 4328 1758
rect 4344 1745 4353 1758
rect 4282 1727 4316 1738
rect 4319 1727 4328 1743
rect 4344 1727 4353 1743
rect 4360 1738 4370 1758
rect 4380 1738 4394 1758
rect 4395 1745 4406 1758
rect 4360 1727 4394 1738
rect 4395 1727 4406 1743
rect 4452 1734 4468 1750
rect 4475 1748 4505 1800
rect 4539 1796 4540 1803
rect 4524 1788 4540 1796
rect 4511 1756 4524 1775
rect 4539 1756 4569 1772
rect 4511 1740 4585 1756
rect 4511 1738 4524 1740
rect 4539 1738 4573 1740
rect 4176 1716 4189 1718
rect 4204 1716 4238 1718
rect 4176 1700 4238 1716
rect 4282 1711 4298 1714
rect 4360 1711 4390 1722
rect 4438 1718 4484 1734
rect 4511 1722 4585 1738
rect 4438 1716 4472 1718
rect 4437 1700 4484 1716
rect 4511 1700 4524 1722
rect 4539 1700 4569 1722
rect 4596 1700 4597 1716
rect 4612 1700 4625 1860
rect -7 1692 34 1700
rect -7 1666 8 1692
rect 15 1666 34 1692
rect 98 1688 160 1700
rect 172 1688 247 1700
rect 305 1688 380 1700
rect 392 1688 423 1700
rect 429 1688 464 1700
rect 98 1686 260 1688
rect -7 1658 34 1666
rect 116 1662 129 1686
rect 144 1684 159 1686
rect -1 1648 0 1658
rect 15 1648 28 1658
rect 43 1648 73 1662
rect 116 1648 159 1662
rect 183 1659 190 1666
rect 193 1662 260 1686
rect 292 1686 464 1688
rect 262 1664 290 1668
rect 292 1664 372 1686
rect 393 1684 408 1686
rect 262 1662 372 1664
rect 193 1658 372 1662
rect 166 1648 196 1658
rect 198 1648 351 1658
rect 359 1648 389 1658
rect 393 1648 423 1662
rect 451 1648 464 1686
rect 536 1692 571 1700
rect 536 1666 537 1692
rect 544 1666 571 1692
rect 479 1648 509 1662
rect 536 1658 571 1666
rect 573 1692 614 1700
rect 573 1666 588 1692
rect 595 1666 614 1692
rect 678 1688 740 1700
rect 752 1688 827 1700
rect 885 1688 960 1700
rect 972 1688 1003 1700
rect 1009 1688 1044 1700
rect 678 1686 840 1688
rect 573 1658 614 1666
rect 696 1662 709 1686
rect 724 1684 739 1686
rect 536 1648 537 1658
rect 552 1648 565 1658
rect 579 1648 580 1658
rect 595 1648 608 1658
rect 623 1648 653 1662
rect 696 1648 739 1662
rect 763 1659 770 1666
rect 773 1662 840 1686
rect 872 1686 1044 1688
rect 842 1664 870 1668
rect 872 1664 952 1686
rect 973 1684 988 1686
rect 842 1662 952 1664
rect 773 1658 952 1662
rect 746 1648 776 1658
rect 778 1648 931 1658
rect 939 1648 969 1658
rect 973 1648 1003 1662
rect 1031 1648 1044 1686
rect 1116 1692 1151 1700
rect 1116 1666 1117 1692
rect 1124 1666 1151 1692
rect 1059 1648 1089 1662
rect 1116 1658 1151 1666
rect 1153 1692 1194 1700
rect 1153 1666 1168 1692
rect 1175 1666 1194 1692
rect 1258 1688 1320 1700
rect 1332 1688 1407 1700
rect 1465 1688 1540 1700
rect 1552 1688 1583 1700
rect 1589 1688 1624 1700
rect 1258 1686 1420 1688
rect 1153 1658 1194 1666
rect 1276 1662 1289 1686
rect 1304 1684 1319 1686
rect 1116 1648 1117 1658
rect 1132 1648 1145 1658
rect 1159 1648 1160 1658
rect 1175 1648 1188 1658
rect 1203 1648 1233 1662
rect 1276 1648 1319 1662
rect 1343 1659 1350 1666
rect 1353 1662 1420 1686
rect 1452 1686 1624 1688
rect 1422 1664 1450 1668
rect 1452 1664 1532 1686
rect 1553 1684 1568 1686
rect 1422 1662 1532 1664
rect 1353 1658 1532 1662
rect 1326 1648 1356 1658
rect 1358 1648 1511 1658
rect 1519 1648 1549 1658
rect 1553 1648 1583 1662
rect 1611 1648 1624 1686
rect 1696 1692 1731 1700
rect 1696 1666 1697 1692
rect 1704 1666 1731 1692
rect 1639 1648 1669 1662
rect 1696 1658 1731 1666
rect 1733 1692 1774 1700
rect 1733 1666 1748 1692
rect 1755 1666 1774 1692
rect 1838 1688 1900 1700
rect 1912 1688 1987 1700
rect 2045 1688 2120 1700
rect 2132 1688 2163 1700
rect 2169 1688 2204 1700
rect 1838 1686 2000 1688
rect 1733 1658 1774 1666
rect 1856 1662 1869 1686
rect 1884 1684 1899 1686
rect 1696 1648 1697 1658
rect 1712 1648 1725 1658
rect 1739 1648 1740 1658
rect 1755 1648 1768 1658
rect 1783 1648 1813 1662
rect 1856 1648 1899 1662
rect 1923 1659 1930 1666
rect 1933 1662 2000 1686
rect 2032 1686 2204 1688
rect 2002 1664 2030 1668
rect 2032 1664 2112 1686
rect 2133 1684 2148 1686
rect 2002 1662 2112 1664
rect 1933 1658 2112 1662
rect 1906 1648 1936 1658
rect 1938 1648 2091 1658
rect 2099 1648 2129 1658
rect 2133 1648 2163 1662
rect 2191 1648 2204 1686
rect 2276 1692 2311 1700
rect 2276 1666 2277 1692
rect 2284 1666 2311 1692
rect 2219 1648 2249 1662
rect 2276 1658 2311 1666
rect 2313 1692 2354 1700
rect 2313 1666 2328 1692
rect 2335 1666 2354 1692
rect 2418 1688 2480 1700
rect 2492 1688 2567 1700
rect 2625 1688 2700 1700
rect 2712 1688 2743 1700
rect 2749 1688 2784 1700
rect 2418 1686 2580 1688
rect 2313 1658 2354 1666
rect 2436 1662 2449 1686
rect 2464 1684 2479 1686
rect 2276 1648 2277 1658
rect 2292 1648 2305 1658
rect 2319 1648 2320 1658
rect 2335 1648 2348 1658
rect 2363 1648 2393 1662
rect 2436 1648 2479 1662
rect 2503 1659 2510 1666
rect 2513 1662 2580 1686
rect 2612 1686 2784 1688
rect 2582 1664 2610 1668
rect 2612 1664 2692 1686
rect 2713 1684 2728 1686
rect 2582 1662 2692 1664
rect 2513 1658 2692 1662
rect 2486 1648 2516 1658
rect 2518 1648 2671 1658
rect 2679 1648 2709 1658
rect 2713 1648 2743 1662
rect 2771 1648 2784 1686
rect 2856 1692 2891 1700
rect 2856 1666 2857 1692
rect 2864 1666 2891 1692
rect 2799 1648 2829 1662
rect 2856 1658 2891 1666
rect 2893 1692 2934 1700
rect 2893 1666 2908 1692
rect 2915 1666 2934 1692
rect 2998 1688 3060 1700
rect 3072 1688 3147 1700
rect 3205 1688 3280 1700
rect 3292 1688 3323 1700
rect 3329 1688 3364 1700
rect 2998 1686 3160 1688
rect 2893 1658 2934 1666
rect 3016 1662 3029 1686
rect 3044 1684 3059 1686
rect 2856 1648 2857 1658
rect 2872 1648 2885 1658
rect 2899 1648 2900 1658
rect 2915 1648 2928 1658
rect 2943 1648 2973 1662
rect 3016 1648 3059 1662
rect 3083 1659 3090 1666
rect 3093 1662 3160 1686
rect 3192 1686 3364 1688
rect 3162 1664 3190 1668
rect 3192 1664 3272 1686
rect 3293 1684 3308 1686
rect 3162 1662 3272 1664
rect 3093 1658 3272 1662
rect 3066 1648 3096 1658
rect 3098 1648 3251 1658
rect 3259 1648 3289 1658
rect 3293 1648 3323 1662
rect 3351 1648 3364 1686
rect 3436 1692 3471 1700
rect 3436 1666 3437 1692
rect 3444 1666 3471 1692
rect 3379 1648 3409 1662
rect 3436 1658 3471 1666
rect 3473 1692 3514 1700
rect 3473 1666 3488 1692
rect 3495 1666 3514 1692
rect 3578 1688 3640 1700
rect 3652 1688 3727 1700
rect 3785 1688 3860 1700
rect 3872 1688 3903 1700
rect 3909 1688 3944 1700
rect 3578 1686 3740 1688
rect 3473 1658 3514 1666
rect 3596 1662 3609 1686
rect 3624 1684 3639 1686
rect 3436 1648 3437 1658
rect 3452 1648 3465 1658
rect 3479 1648 3480 1658
rect 3495 1648 3508 1658
rect 3523 1648 3553 1662
rect 3596 1648 3639 1662
rect 3663 1659 3670 1666
rect 3673 1662 3740 1686
rect 3772 1686 3944 1688
rect 3742 1664 3770 1668
rect 3772 1664 3852 1686
rect 3873 1684 3888 1686
rect 3742 1662 3852 1664
rect 3673 1658 3852 1662
rect 3646 1648 3676 1658
rect 3678 1648 3831 1658
rect 3839 1648 3869 1658
rect 3873 1648 3903 1662
rect 3931 1648 3944 1686
rect 4016 1692 4051 1700
rect 4016 1666 4017 1692
rect 4024 1666 4051 1692
rect 3959 1648 3989 1662
rect 4016 1658 4051 1666
rect 4053 1692 4094 1700
rect 4053 1666 4068 1692
rect 4075 1666 4094 1692
rect 4158 1688 4220 1700
rect 4232 1688 4307 1700
rect 4365 1688 4440 1700
rect 4452 1688 4483 1700
rect 4489 1688 4524 1700
rect 4158 1686 4320 1688
rect 4053 1658 4094 1666
rect 4176 1662 4189 1686
rect 4204 1684 4219 1686
rect 4016 1648 4017 1658
rect 4032 1648 4045 1658
rect 4059 1648 4060 1658
rect 4075 1648 4088 1658
rect 4103 1648 4133 1662
rect 4176 1648 4219 1662
rect 4243 1659 4250 1666
rect 4253 1662 4320 1686
rect 4352 1686 4524 1688
rect 4322 1664 4350 1668
rect 4352 1664 4432 1686
rect 4453 1684 4468 1686
rect 4322 1662 4432 1664
rect 4253 1658 4432 1662
rect 4226 1648 4256 1658
rect 4258 1648 4411 1658
rect 4419 1648 4449 1658
rect 4453 1648 4483 1662
rect 4511 1648 4524 1686
rect 4596 1692 4631 1700
rect 4596 1666 4597 1692
rect 4604 1666 4631 1692
rect 4539 1648 4569 1662
rect 4596 1658 4631 1666
rect 4596 1648 4597 1658
rect 4612 1648 4625 1658
rect -1 1642 4625 1648
rect 0 1634 4625 1642
rect 15 1604 28 1634
rect 43 1616 73 1634
rect 116 1620 130 1634
rect 166 1620 386 1634
rect 117 1618 130 1620
rect 83 1606 98 1618
rect 80 1604 102 1606
rect 107 1604 137 1618
rect 198 1616 351 1620
rect 180 1604 372 1616
rect 415 1604 445 1618
rect 451 1604 464 1634
rect 479 1616 509 1634
rect 552 1604 565 1634
rect 595 1604 608 1634
rect 623 1616 653 1634
rect 696 1620 710 1634
rect 746 1620 966 1634
rect 697 1618 710 1620
rect 663 1606 678 1618
rect 660 1604 682 1606
rect 687 1604 717 1618
rect 778 1616 931 1620
rect 760 1604 952 1616
rect 995 1604 1025 1618
rect 1031 1604 1044 1634
rect 1059 1616 1089 1634
rect 1132 1604 1145 1634
rect 1175 1604 1188 1634
rect 1203 1616 1233 1634
rect 1276 1620 1290 1634
rect 1326 1620 1546 1634
rect 1277 1618 1290 1620
rect 1243 1606 1258 1618
rect 1240 1604 1262 1606
rect 1267 1604 1297 1618
rect 1358 1616 1511 1620
rect 1340 1604 1532 1616
rect 1575 1604 1605 1618
rect 1611 1604 1624 1634
rect 1639 1616 1669 1634
rect 1712 1604 1725 1634
rect 1755 1604 1768 1634
rect 1783 1616 1813 1634
rect 1856 1620 1870 1634
rect 1906 1620 2126 1634
rect 1857 1618 1870 1620
rect 1823 1606 1838 1618
rect 1820 1604 1842 1606
rect 1847 1604 1877 1618
rect 1938 1616 2091 1620
rect 1920 1604 2112 1616
rect 2155 1604 2185 1618
rect 2191 1604 2204 1634
rect 2219 1616 2249 1634
rect 2292 1604 2305 1634
rect 2335 1604 2348 1634
rect 2363 1616 2393 1634
rect 2436 1620 2450 1634
rect 2486 1620 2706 1634
rect 2437 1618 2450 1620
rect 2403 1606 2418 1618
rect 2400 1604 2422 1606
rect 2427 1604 2457 1618
rect 2518 1616 2671 1620
rect 2500 1604 2692 1616
rect 2735 1604 2765 1618
rect 2771 1604 2784 1634
rect 2799 1616 2829 1634
rect 2872 1604 2885 1634
rect 2915 1604 2928 1634
rect 2943 1616 2973 1634
rect 3016 1620 3030 1634
rect 3066 1620 3286 1634
rect 3017 1618 3030 1620
rect 2983 1606 2998 1618
rect 2980 1604 3002 1606
rect 3007 1604 3037 1618
rect 3098 1616 3251 1620
rect 3080 1604 3272 1616
rect 3315 1604 3345 1618
rect 3351 1604 3364 1634
rect 3379 1616 3409 1634
rect 3452 1604 3465 1634
rect 3495 1604 3508 1634
rect 3523 1616 3553 1634
rect 3596 1620 3610 1634
rect 3646 1620 3866 1634
rect 3597 1618 3610 1620
rect 3563 1606 3578 1618
rect 3560 1604 3582 1606
rect 3587 1604 3617 1618
rect 3678 1616 3831 1620
rect 3660 1604 3852 1616
rect 3895 1604 3925 1618
rect 3931 1604 3944 1634
rect 3959 1616 3989 1634
rect 4032 1604 4045 1634
rect 4075 1604 4088 1634
rect 4103 1616 4133 1634
rect 4176 1620 4190 1634
rect 4226 1620 4446 1634
rect 4177 1618 4190 1620
rect 4143 1606 4158 1618
rect 4140 1604 4162 1606
rect 4167 1604 4197 1618
rect 4258 1616 4411 1620
rect 4240 1604 4432 1616
rect 4475 1604 4505 1618
rect 4511 1604 4524 1634
rect 4539 1616 4569 1634
rect 4612 1604 4625 1634
rect 0 1590 4625 1604
rect 15 1486 28 1590
rect 73 1568 74 1578
rect 89 1568 102 1578
rect 73 1564 102 1568
rect 107 1564 137 1590
rect 155 1576 171 1578
rect 243 1576 296 1590
rect 244 1574 308 1576
rect 351 1574 366 1590
rect 415 1587 445 1590
rect 415 1584 451 1587
rect 381 1576 397 1578
rect 155 1564 170 1568
rect 73 1562 170 1564
rect 198 1562 366 1574
rect 382 1564 397 1568
rect 415 1565 454 1584
rect 473 1578 480 1579
rect 479 1571 480 1578
rect 463 1568 464 1571
rect 479 1568 492 1571
rect 415 1564 445 1565
rect 454 1564 460 1565
rect 463 1564 492 1568
rect 382 1563 492 1564
rect 382 1562 498 1563
rect 57 1554 108 1562
rect 57 1542 82 1554
rect 89 1542 108 1554
rect 139 1554 189 1562
rect 139 1546 155 1554
rect 162 1552 189 1554
rect 198 1552 419 1562
rect 162 1542 419 1552
rect 448 1554 498 1562
rect 448 1545 464 1554
rect 57 1534 108 1542
rect 155 1534 419 1542
rect 445 1542 464 1545
rect 471 1542 498 1554
rect 445 1534 498 1542
rect 73 1526 74 1534
rect 89 1526 102 1534
rect 73 1518 89 1526
rect 70 1511 89 1514
rect 70 1502 92 1511
rect 43 1492 92 1502
rect 43 1486 73 1492
rect 92 1487 97 1492
rect 15 1470 89 1486
rect 107 1478 137 1534
rect 172 1524 380 1534
rect 415 1530 460 1534
rect 463 1533 464 1534
rect 479 1533 492 1534
rect 198 1494 387 1524
rect 213 1491 387 1494
rect 206 1488 387 1491
rect 15 1468 28 1470
rect 43 1468 77 1470
rect 15 1452 89 1468
rect 116 1464 129 1478
rect 144 1464 160 1480
rect 206 1475 217 1488
rect -1 1430 0 1446
rect 15 1430 28 1452
rect 43 1430 73 1452
rect 116 1448 178 1464
rect 206 1457 217 1473
rect 222 1468 232 1488
rect 242 1468 256 1488
rect 259 1475 268 1488
rect 284 1475 293 1488
rect 222 1457 256 1468
rect 259 1457 268 1473
rect 284 1457 293 1473
rect 300 1468 310 1488
rect 320 1468 334 1488
rect 335 1475 346 1488
rect 300 1457 334 1468
rect 335 1457 346 1473
rect 392 1464 408 1480
rect 415 1478 445 1530
rect 479 1526 480 1533
rect 464 1518 480 1526
rect 451 1486 464 1505
rect 479 1486 509 1502
rect 451 1470 525 1486
rect 451 1468 464 1470
rect 479 1468 513 1470
rect 116 1446 129 1448
rect 144 1446 178 1448
rect 116 1430 178 1446
rect 222 1441 238 1444
rect 300 1441 330 1452
rect 378 1448 424 1464
rect 451 1452 525 1468
rect 378 1446 412 1448
rect 377 1430 424 1446
rect 451 1430 464 1452
rect 479 1430 509 1452
rect 536 1430 537 1446
rect 552 1430 565 1590
rect 595 1486 608 1590
rect 653 1568 654 1578
rect 669 1568 682 1578
rect 653 1564 682 1568
rect 687 1564 717 1590
rect 735 1576 751 1578
rect 823 1576 876 1590
rect 824 1574 888 1576
rect 931 1574 946 1590
rect 995 1587 1025 1590
rect 995 1584 1031 1587
rect 961 1576 977 1578
rect 735 1564 750 1568
rect 653 1562 750 1564
rect 778 1562 946 1574
rect 962 1564 977 1568
rect 995 1565 1034 1584
rect 1053 1578 1060 1579
rect 1059 1571 1060 1578
rect 1043 1568 1044 1571
rect 1059 1568 1072 1571
rect 995 1564 1025 1565
rect 1034 1564 1040 1565
rect 1043 1564 1072 1568
rect 962 1563 1072 1564
rect 962 1562 1078 1563
rect 637 1554 688 1562
rect 637 1542 662 1554
rect 669 1542 688 1554
rect 719 1554 769 1562
rect 719 1546 735 1554
rect 742 1552 769 1554
rect 778 1552 999 1562
rect 742 1542 999 1552
rect 1028 1554 1078 1562
rect 1028 1545 1044 1554
rect 637 1534 688 1542
rect 735 1534 999 1542
rect 1025 1542 1044 1545
rect 1051 1542 1078 1554
rect 1025 1534 1078 1542
rect 653 1526 654 1534
rect 669 1526 682 1534
rect 653 1518 669 1526
rect 650 1511 669 1514
rect 650 1502 672 1511
rect 623 1492 672 1502
rect 623 1486 653 1492
rect 672 1487 677 1492
rect 595 1470 669 1486
rect 687 1478 717 1534
rect 752 1524 960 1534
rect 995 1530 1040 1534
rect 1043 1533 1044 1534
rect 1059 1533 1072 1534
rect 778 1494 967 1524
rect 793 1491 967 1494
rect 786 1488 967 1491
rect 595 1468 608 1470
rect 623 1468 657 1470
rect 595 1452 669 1468
rect 696 1464 709 1478
rect 724 1464 740 1480
rect 786 1475 797 1488
rect 579 1430 580 1446
rect 595 1430 608 1452
rect 623 1430 653 1452
rect 696 1448 758 1464
rect 786 1457 797 1473
rect 802 1468 812 1488
rect 822 1468 836 1488
rect 839 1475 848 1488
rect 864 1475 873 1488
rect 802 1457 836 1468
rect 839 1457 848 1473
rect 864 1457 873 1473
rect 880 1468 890 1488
rect 900 1468 914 1488
rect 915 1475 926 1488
rect 880 1457 914 1468
rect 915 1457 926 1473
rect 972 1464 988 1480
rect 995 1478 1025 1530
rect 1059 1526 1060 1533
rect 1044 1518 1060 1526
rect 1031 1486 1044 1505
rect 1059 1486 1089 1502
rect 1031 1470 1105 1486
rect 1031 1468 1044 1470
rect 1059 1468 1093 1470
rect 696 1446 709 1448
rect 724 1446 758 1448
rect 696 1430 758 1446
rect 802 1441 818 1444
rect 880 1441 910 1452
rect 958 1448 1004 1464
rect 1031 1452 1105 1468
rect 958 1446 992 1448
rect 957 1430 1004 1446
rect 1031 1430 1044 1452
rect 1059 1430 1089 1452
rect 1116 1430 1117 1446
rect 1132 1430 1145 1590
rect 1175 1486 1188 1590
rect 1233 1568 1234 1578
rect 1249 1568 1262 1578
rect 1233 1564 1262 1568
rect 1267 1564 1297 1590
rect 1315 1576 1331 1578
rect 1403 1576 1456 1590
rect 1404 1574 1468 1576
rect 1511 1574 1526 1590
rect 1575 1587 1605 1590
rect 1575 1584 1611 1587
rect 1541 1576 1557 1578
rect 1315 1564 1330 1568
rect 1233 1562 1330 1564
rect 1358 1562 1526 1574
rect 1542 1564 1557 1568
rect 1575 1565 1614 1584
rect 1633 1578 1640 1579
rect 1639 1571 1640 1578
rect 1623 1568 1624 1571
rect 1639 1568 1652 1571
rect 1575 1564 1605 1565
rect 1614 1564 1620 1565
rect 1623 1564 1652 1568
rect 1542 1563 1652 1564
rect 1542 1562 1658 1563
rect 1217 1554 1268 1562
rect 1217 1542 1242 1554
rect 1249 1542 1268 1554
rect 1299 1554 1349 1562
rect 1299 1546 1315 1554
rect 1322 1552 1349 1554
rect 1358 1552 1579 1562
rect 1322 1542 1579 1552
rect 1608 1554 1658 1562
rect 1608 1545 1624 1554
rect 1217 1534 1268 1542
rect 1315 1534 1579 1542
rect 1605 1542 1624 1545
rect 1631 1542 1658 1554
rect 1605 1534 1658 1542
rect 1233 1526 1234 1534
rect 1249 1526 1262 1534
rect 1233 1518 1249 1526
rect 1230 1511 1249 1514
rect 1230 1502 1252 1511
rect 1203 1492 1252 1502
rect 1203 1486 1233 1492
rect 1252 1487 1257 1492
rect 1175 1470 1249 1486
rect 1267 1478 1297 1534
rect 1332 1524 1540 1534
rect 1575 1530 1620 1534
rect 1623 1533 1624 1534
rect 1639 1533 1652 1534
rect 1358 1494 1547 1524
rect 1373 1491 1547 1494
rect 1366 1488 1547 1491
rect 1175 1468 1188 1470
rect 1203 1468 1237 1470
rect 1175 1452 1249 1468
rect 1276 1464 1289 1478
rect 1304 1464 1320 1480
rect 1366 1475 1377 1488
rect 1159 1430 1160 1446
rect 1175 1430 1188 1452
rect 1203 1430 1233 1452
rect 1276 1448 1338 1464
rect 1366 1457 1377 1473
rect 1382 1468 1392 1488
rect 1402 1468 1416 1488
rect 1419 1475 1428 1488
rect 1444 1475 1453 1488
rect 1382 1457 1416 1468
rect 1419 1457 1428 1473
rect 1444 1457 1453 1473
rect 1460 1468 1470 1488
rect 1480 1468 1494 1488
rect 1495 1475 1506 1488
rect 1460 1457 1494 1468
rect 1495 1457 1506 1473
rect 1552 1464 1568 1480
rect 1575 1478 1605 1530
rect 1639 1526 1640 1533
rect 1624 1518 1640 1526
rect 1611 1486 1624 1505
rect 1639 1486 1669 1502
rect 1611 1470 1685 1486
rect 1611 1468 1624 1470
rect 1639 1468 1673 1470
rect 1276 1446 1289 1448
rect 1304 1446 1338 1448
rect 1276 1430 1338 1446
rect 1382 1441 1398 1444
rect 1460 1441 1490 1452
rect 1538 1448 1584 1464
rect 1611 1452 1685 1468
rect 1538 1446 1572 1448
rect 1537 1430 1584 1446
rect 1611 1430 1624 1452
rect 1639 1430 1669 1452
rect 1696 1430 1697 1446
rect 1712 1430 1725 1590
rect 1755 1486 1768 1590
rect 1813 1568 1814 1578
rect 1829 1568 1842 1578
rect 1813 1564 1842 1568
rect 1847 1564 1877 1590
rect 1895 1576 1911 1578
rect 1983 1576 2036 1590
rect 1984 1574 2048 1576
rect 2091 1574 2106 1590
rect 2155 1587 2185 1590
rect 2155 1584 2191 1587
rect 2121 1576 2137 1578
rect 1895 1564 1910 1568
rect 1813 1562 1910 1564
rect 1938 1562 2106 1574
rect 2122 1564 2137 1568
rect 2155 1565 2194 1584
rect 2213 1578 2220 1579
rect 2219 1571 2220 1578
rect 2203 1568 2204 1571
rect 2219 1568 2232 1571
rect 2155 1564 2185 1565
rect 2194 1564 2200 1565
rect 2203 1564 2232 1568
rect 2122 1563 2232 1564
rect 2122 1562 2238 1563
rect 1797 1554 1848 1562
rect 1797 1542 1822 1554
rect 1829 1542 1848 1554
rect 1879 1554 1929 1562
rect 1879 1546 1895 1554
rect 1902 1552 1929 1554
rect 1938 1552 2159 1562
rect 1902 1542 2159 1552
rect 2188 1554 2238 1562
rect 2188 1545 2204 1554
rect 1797 1534 1848 1542
rect 1895 1534 2159 1542
rect 2185 1542 2204 1545
rect 2211 1542 2238 1554
rect 2185 1534 2238 1542
rect 1813 1526 1814 1534
rect 1829 1526 1842 1534
rect 1813 1518 1829 1526
rect 1810 1511 1829 1514
rect 1810 1502 1832 1511
rect 1783 1492 1832 1502
rect 1783 1486 1813 1492
rect 1832 1487 1837 1492
rect 1755 1470 1829 1486
rect 1847 1478 1877 1534
rect 1912 1524 2120 1534
rect 2155 1530 2200 1534
rect 2203 1533 2204 1534
rect 2219 1533 2232 1534
rect 1938 1494 2127 1524
rect 1953 1491 2127 1494
rect 1946 1488 2127 1491
rect 1755 1468 1768 1470
rect 1783 1468 1817 1470
rect 1755 1452 1829 1468
rect 1856 1464 1869 1478
rect 1884 1464 1900 1480
rect 1946 1475 1957 1488
rect 1739 1430 1740 1446
rect 1755 1430 1768 1452
rect 1783 1430 1813 1452
rect 1856 1448 1918 1464
rect 1946 1457 1957 1473
rect 1962 1468 1972 1488
rect 1982 1468 1996 1488
rect 1999 1475 2008 1488
rect 2024 1475 2033 1488
rect 1962 1457 1996 1468
rect 1999 1457 2008 1473
rect 2024 1457 2033 1473
rect 2040 1468 2050 1488
rect 2060 1468 2074 1488
rect 2075 1475 2086 1488
rect 2040 1457 2074 1468
rect 2075 1457 2086 1473
rect 2132 1464 2148 1480
rect 2155 1478 2185 1530
rect 2219 1526 2220 1533
rect 2204 1518 2220 1526
rect 2191 1486 2204 1505
rect 2219 1486 2249 1502
rect 2191 1470 2265 1486
rect 2191 1468 2204 1470
rect 2219 1468 2253 1470
rect 1856 1446 1869 1448
rect 1884 1446 1918 1448
rect 1856 1430 1918 1446
rect 1962 1441 1978 1444
rect 2040 1441 2070 1452
rect 2118 1448 2164 1464
rect 2191 1452 2265 1468
rect 2118 1446 2152 1448
rect 2117 1430 2164 1446
rect 2191 1430 2204 1452
rect 2219 1430 2249 1452
rect 2276 1430 2277 1446
rect 2292 1430 2305 1590
rect 2335 1486 2348 1590
rect 2393 1568 2394 1578
rect 2409 1568 2422 1578
rect 2393 1564 2422 1568
rect 2427 1564 2457 1590
rect 2475 1576 2491 1578
rect 2563 1576 2616 1590
rect 2564 1574 2628 1576
rect 2671 1574 2686 1590
rect 2735 1587 2765 1590
rect 2735 1584 2771 1587
rect 2701 1576 2717 1578
rect 2475 1564 2490 1568
rect 2393 1562 2490 1564
rect 2518 1562 2686 1574
rect 2702 1564 2717 1568
rect 2735 1565 2774 1584
rect 2793 1578 2800 1579
rect 2799 1571 2800 1578
rect 2783 1568 2784 1571
rect 2799 1568 2812 1571
rect 2735 1564 2765 1565
rect 2774 1564 2780 1565
rect 2783 1564 2812 1568
rect 2702 1563 2812 1564
rect 2702 1562 2818 1563
rect 2377 1554 2428 1562
rect 2377 1542 2402 1554
rect 2409 1542 2428 1554
rect 2459 1554 2509 1562
rect 2459 1546 2475 1554
rect 2482 1552 2509 1554
rect 2518 1552 2739 1562
rect 2482 1542 2739 1552
rect 2768 1554 2818 1562
rect 2768 1545 2784 1554
rect 2377 1534 2428 1542
rect 2475 1534 2739 1542
rect 2765 1542 2784 1545
rect 2791 1542 2818 1554
rect 2765 1534 2818 1542
rect 2393 1526 2394 1534
rect 2409 1526 2422 1534
rect 2393 1518 2409 1526
rect 2390 1511 2409 1514
rect 2390 1502 2412 1511
rect 2363 1492 2412 1502
rect 2363 1486 2393 1492
rect 2412 1487 2417 1492
rect 2335 1470 2409 1486
rect 2427 1478 2457 1534
rect 2492 1524 2700 1534
rect 2735 1530 2780 1534
rect 2783 1533 2784 1534
rect 2799 1533 2812 1534
rect 2518 1494 2707 1524
rect 2533 1491 2707 1494
rect 2526 1488 2707 1491
rect 2335 1468 2348 1470
rect 2363 1468 2397 1470
rect 2335 1452 2409 1468
rect 2436 1464 2449 1478
rect 2464 1464 2480 1480
rect 2526 1475 2537 1488
rect 2319 1430 2320 1446
rect 2335 1430 2348 1452
rect 2363 1430 2393 1452
rect 2436 1448 2498 1464
rect 2526 1457 2537 1473
rect 2542 1468 2552 1488
rect 2562 1468 2576 1488
rect 2579 1475 2588 1488
rect 2604 1475 2613 1488
rect 2542 1457 2576 1468
rect 2579 1457 2588 1473
rect 2604 1457 2613 1473
rect 2620 1468 2630 1488
rect 2640 1468 2654 1488
rect 2655 1475 2666 1488
rect 2620 1457 2654 1468
rect 2655 1457 2666 1473
rect 2712 1464 2728 1480
rect 2735 1478 2765 1530
rect 2799 1526 2800 1533
rect 2784 1518 2800 1526
rect 2771 1486 2784 1505
rect 2799 1486 2829 1502
rect 2771 1470 2845 1486
rect 2771 1468 2784 1470
rect 2799 1468 2833 1470
rect 2436 1446 2449 1448
rect 2464 1446 2498 1448
rect 2436 1430 2498 1446
rect 2542 1441 2558 1444
rect 2620 1441 2650 1452
rect 2698 1448 2744 1464
rect 2771 1452 2845 1468
rect 2698 1446 2732 1448
rect 2697 1430 2744 1446
rect 2771 1430 2784 1452
rect 2799 1430 2829 1452
rect 2856 1430 2857 1446
rect 2872 1430 2885 1590
rect 2915 1486 2928 1590
rect 2973 1568 2974 1578
rect 2989 1568 3002 1578
rect 2973 1564 3002 1568
rect 3007 1564 3037 1590
rect 3055 1576 3071 1578
rect 3143 1576 3196 1590
rect 3144 1574 3208 1576
rect 3251 1574 3266 1590
rect 3315 1587 3345 1590
rect 3315 1584 3351 1587
rect 3281 1576 3297 1578
rect 3055 1564 3070 1568
rect 2973 1562 3070 1564
rect 3098 1562 3266 1574
rect 3282 1564 3297 1568
rect 3315 1565 3354 1584
rect 3373 1578 3380 1579
rect 3379 1571 3380 1578
rect 3363 1568 3364 1571
rect 3379 1568 3392 1571
rect 3315 1564 3345 1565
rect 3354 1564 3360 1565
rect 3363 1564 3392 1568
rect 3282 1563 3392 1564
rect 3282 1562 3398 1563
rect 2957 1554 3008 1562
rect 2957 1542 2982 1554
rect 2989 1542 3008 1554
rect 3039 1554 3089 1562
rect 3039 1546 3055 1554
rect 3062 1552 3089 1554
rect 3098 1552 3319 1562
rect 3062 1542 3319 1552
rect 3348 1554 3398 1562
rect 3348 1545 3364 1554
rect 2957 1534 3008 1542
rect 3055 1534 3319 1542
rect 3345 1542 3364 1545
rect 3371 1542 3398 1554
rect 3345 1534 3398 1542
rect 2973 1526 2974 1534
rect 2989 1526 3002 1534
rect 2973 1518 2989 1526
rect 2970 1511 2989 1514
rect 2970 1502 2992 1511
rect 2943 1492 2992 1502
rect 2943 1486 2973 1492
rect 2992 1487 2997 1492
rect 2915 1470 2989 1486
rect 3007 1478 3037 1534
rect 3072 1524 3280 1534
rect 3315 1530 3360 1534
rect 3363 1533 3364 1534
rect 3379 1533 3392 1534
rect 3098 1494 3287 1524
rect 3113 1491 3287 1494
rect 3106 1488 3287 1491
rect 2915 1468 2928 1470
rect 2943 1468 2977 1470
rect 2915 1452 2989 1468
rect 3016 1464 3029 1478
rect 3044 1464 3060 1480
rect 3106 1475 3117 1488
rect 2899 1430 2900 1446
rect 2915 1430 2928 1452
rect 2943 1430 2973 1452
rect 3016 1448 3078 1464
rect 3106 1457 3117 1473
rect 3122 1468 3132 1488
rect 3142 1468 3156 1488
rect 3159 1475 3168 1488
rect 3184 1475 3193 1488
rect 3122 1457 3156 1468
rect 3159 1457 3168 1473
rect 3184 1457 3193 1473
rect 3200 1468 3210 1488
rect 3220 1468 3234 1488
rect 3235 1475 3246 1488
rect 3200 1457 3234 1468
rect 3235 1457 3246 1473
rect 3292 1464 3308 1480
rect 3315 1478 3345 1530
rect 3379 1526 3380 1533
rect 3364 1518 3380 1526
rect 3351 1486 3364 1505
rect 3379 1486 3409 1502
rect 3351 1470 3425 1486
rect 3351 1468 3364 1470
rect 3379 1468 3413 1470
rect 3016 1446 3029 1448
rect 3044 1446 3078 1448
rect 3016 1430 3078 1446
rect 3122 1441 3138 1444
rect 3200 1441 3230 1452
rect 3278 1448 3324 1464
rect 3351 1452 3425 1468
rect 3278 1446 3312 1448
rect 3277 1430 3324 1446
rect 3351 1430 3364 1452
rect 3379 1430 3409 1452
rect 3436 1430 3437 1446
rect 3452 1430 3465 1590
rect 3495 1486 3508 1590
rect 3553 1568 3554 1578
rect 3569 1568 3582 1578
rect 3553 1564 3582 1568
rect 3587 1564 3617 1590
rect 3635 1576 3651 1578
rect 3723 1576 3776 1590
rect 3724 1574 3788 1576
rect 3831 1574 3846 1590
rect 3895 1587 3925 1590
rect 3895 1584 3931 1587
rect 3861 1576 3877 1578
rect 3635 1564 3650 1568
rect 3553 1562 3650 1564
rect 3678 1562 3846 1574
rect 3862 1564 3877 1568
rect 3895 1565 3934 1584
rect 3953 1578 3960 1579
rect 3959 1571 3960 1578
rect 3943 1568 3944 1571
rect 3959 1568 3972 1571
rect 3895 1564 3925 1565
rect 3934 1564 3940 1565
rect 3943 1564 3972 1568
rect 3862 1563 3972 1564
rect 3862 1562 3978 1563
rect 3537 1554 3588 1562
rect 3537 1542 3562 1554
rect 3569 1542 3588 1554
rect 3619 1554 3669 1562
rect 3619 1546 3635 1554
rect 3642 1552 3669 1554
rect 3678 1552 3899 1562
rect 3642 1542 3899 1552
rect 3928 1554 3978 1562
rect 3928 1545 3944 1554
rect 3537 1534 3588 1542
rect 3635 1534 3899 1542
rect 3925 1542 3944 1545
rect 3951 1542 3978 1554
rect 3925 1534 3978 1542
rect 3553 1526 3554 1534
rect 3569 1526 3582 1534
rect 3553 1518 3569 1526
rect 3550 1511 3569 1514
rect 3550 1502 3572 1511
rect 3523 1492 3572 1502
rect 3523 1486 3553 1492
rect 3572 1487 3577 1492
rect 3495 1470 3569 1486
rect 3587 1478 3617 1534
rect 3652 1524 3860 1534
rect 3895 1530 3940 1534
rect 3943 1533 3944 1534
rect 3959 1533 3972 1534
rect 3678 1494 3867 1524
rect 3693 1491 3867 1494
rect 3686 1488 3867 1491
rect 3495 1468 3508 1470
rect 3523 1468 3557 1470
rect 3495 1452 3569 1468
rect 3596 1464 3609 1478
rect 3624 1464 3640 1480
rect 3686 1475 3697 1488
rect 3479 1430 3480 1446
rect 3495 1430 3508 1452
rect 3523 1430 3553 1452
rect 3596 1448 3658 1464
rect 3686 1457 3697 1473
rect 3702 1468 3712 1488
rect 3722 1468 3736 1488
rect 3739 1475 3748 1488
rect 3764 1475 3773 1488
rect 3702 1457 3736 1468
rect 3739 1457 3748 1473
rect 3764 1457 3773 1473
rect 3780 1468 3790 1488
rect 3800 1468 3814 1488
rect 3815 1475 3826 1488
rect 3780 1457 3814 1468
rect 3815 1457 3826 1473
rect 3872 1464 3888 1480
rect 3895 1478 3925 1530
rect 3959 1526 3960 1533
rect 3944 1518 3960 1526
rect 3931 1486 3944 1505
rect 3959 1486 3989 1502
rect 3931 1470 4005 1486
rect 3931 1468 3944 1470
rect 3959 1468 3993 1470
rect 3596 1446 3609 1448
rect 3624 1446 3658 1448
rect 3596 1430 3658 1446
rect 3702 1441 3718 1444
rect 3780 1441 3810 1452
rect 3858 1448 3904 1464
rect 3931 1452 4005 1468
rect 3858 1446 3892 1448
rect 3857 1430 3904 1446
rect 3931 1430 3944 1452
rect 3959 1430 3989 1452
rect 4016 1430 4017 1446
rect 4032 1430 4045 1590
rect 4075 1486 4088 1590
rect 4133 1568 4134 1578
rect 4149 1568 4162 1578
rect 4133 1564 4162 1568
rect 4167 1564 4197 1590
rect 4215 1576 4231 1578
rect 4303 1576 4356 1590
rect 4304 1574 4368 1576
rect 4411 1574 4426 1590
rect 4475 1587 4505 1590
rect 4475 1584 4511 1587
rect 4441 1576 4457 1578
rect 4215 1564 4230 1568
rect 4133 1562 4230 1564
rect 4258 1562 4426 1574
rect 4442 1564 4457 1568
rect 4475 1565 4514 1584
rect 4533 1578 4540 1579
rect 4539 1571 4540 1578
rect 4523 1568 4524 1571
rect 4539 1568 4552 1571
rect 4475 1564 4505 1565
rect 4514 1564 4520 1565
rect 4523 1564 4552 1568
rect 4442 1563 4552 1564
rect 4442 1562 4558 1563
rect 4117 1554 4168 1562
rect 4117 1542 4142 1554
rect 4149 1542 4168 1554
rect 4199 1554 4249 1562
rect 4199 1546 4215 1554
rect 4222 1552 4249 1554
rect 4258 1552 4479 1562
rect 4222 1542 4479 1552
rect 4508 1554 4558 1562
rect 4508 1545 4524 1554
rect 4117 1534 4168 1542
rect 4215 1534 4479 1542
rect 4505 1542 4524 1545
rect 4531 1542 4558 1554
rect 4505 1534 4558 1542
rect 4133 1526 4134 1534
rect 4149 1526 4162 1534
rect 4133 1518 4149 1526
rect 4130 1511 4149 1514
rect 4130 1502 4152 1511
rect 4103 1492 4152 1502
rect 4103 1486 4133 1492
rect 4152 1487 4157 1492
rect 4075 1470 4149 1486
rect 4167 1478 4197 1534
rect 4232 1524 4440 1534
rect 4475 1530 4520 1534
rect 4523 1533 4524 1534
rect 4539 1533 4552 1534
rect 4258 1494 4447 1524
rect 4273 1491 4447 1494
rect 4266 1488 4447 1491
rect 4075 1468 4088 1470
rect 4103 1468 4137 1470
rect 4075 1452 4149 1468
rect 4176 1464 4189 1478
rect 4204 1464 4220 1480
rect 4266 1475 4277 1488
rect 4059 1430 4060 1446
rect 4075 1430 4088 1452
rect 4103 1430 4133 1452
rect 4176 1448 4238 1464
rect 4266 1457 4277 1473
rect 4282 1468 4292 1488
rect 4302 1468 4316 1488
rect 4319 1475 4328 1488
rect 4344 1475 4353 1488
rect 4282 1457 4316 1468
rect 4319 1457 4328 1473
rect 4344 1457 4353 1473
rect 4360 1468 4370 1488
rect 4380 1468 4394 1488
rect 4395 1475 4406 1488
rect 4360 1457 4394 1468
rect 4395 1457 4406 1473
rect 4452 1464 4468 1480
rect 4475 1478 4505 1530
rect 4539 1526 4540 1533
rect 4524 1518 4540 1526
rect 4511 1486 4524 1505
rect 4539 1486 4569 1502
rect 4511 1470 4585 1486
rect 4511 1468 4524 1470
rect 4539 1468 4573 1470
rect 4176 1446 4189 1448
rect 4204 1446 4238 1448
rect 4176 1430 4238 1446
rect 4282 1441 4298 1444
rect 4360 1441 4390 1452
rect 4438 1448 4484 1464
rect 4511 1452 4585 1468
rect 4438 1446 4472 1448
rect 4437 1430 4484 1446
rect 4511 1430 4524 1452
rect 4539 1430 4569 1452
rect 4596 1430 4597 1446
rect 4612 1430 4625 1590
rect -7 1422 34 1430
rect -7 1396 8 1422
rect 15 1396 34 1422
rect 98 1418 160 1430
rect 172 1418 247 1430
rect 305 1418 380 1430
rect 392 1418 423 1430
rect 429 1418 464 1430
rect 98 1416 260 1418
rect -7 1388 34 1396
rect 116 1392 129 1416
rect 144 1414 159 1416
rect -1 1378 0 1388
rect 15 1378 28 1388
rect 43 1378 73 1392
rect 116 1378 159 1392
rect 183 1389 190 1396
rect 193 1392 260 1416
rect 292 1416 464 1418
rect 262 1394 290 1398
rect 292 1394 372 1416
rect 393 1414 408 1416
rect 262 1392 372 1394
rect 193 1388 372 1392
rect 166 1378 196 1388
rect 198 1378 351 1388
rect 359 1378 389 1388
rect 393 1378 423 1392
rect 451 1378 464 1416
rect 536 1422 571 1430
rect 536 1396 537 1422
rect 544 1396 571 1422
rect 479 1378 509 1392
rect 536 1388 571 1396
rect 573 1422 614 1430
rect 573 1396 588 1422
rect 595 1396 614 1422
rect 678 1418 740 1430
rect 752 1418 827 1430
rect 885 1418 960 1430
rect 972 1418 1003 1430
rect 1009 1418 1044 1430
rect 678 1416 840 1418
rect 573 1388 614 1396
rect 696 1392 709 1416
rect 724 1414 739 1416
rect 536 1378 537 1388
rect 552 1378 565 1388
rect 579 1378 580 1388
rect 595 1378 608 1388
rect 623 1378 653 1392
rect 696 1378 739 1392
rect 763 1389 770 1396
rect 773 1392 840 1416
rect 872 1416 1044 1418
rect 842 1394 870 1398
rect 872 1394 952 1416
rect 973 1414 988 1416
rect 842 1392 952 1394
rect 773 1388 952 1392
rect 746 1378 776 1388
rect 778 1378 931 1388
rect 939 1378 969 1388
rect 973 1378 1003 1392
rect 1031 1378 1044 1416
rect 1116 1422 1151 1430
rect 1116 1396 1117 1422
rect 1124 1396 1151 1422
rect 1059 1378 1089 1392
rect 1116 1388 1151 1396
rect 1153 1422 1194 1430
rect 1153 1396 1168 1422
rect 1175 1396 1194 1422
rect 1258 1418 1320 1430
rect 1332 1418 1407 1430
rect 1465 1418 1540 1430
rect 1552 1418 1583 1430
rect 1589 1418 1624 1430
rect 1258 1416 1420 1418
rect 1153 1388 1194 1396
rect 1276 1392 1289 1416
rect 1304 1414 1319 1416
rect 1116 1378 1117 1388
rect 1132 1378 1145 1388
rect 1159 1378 1160 1388
rect 1175 1378 1188 1388
rect 1203 1378 1233 1392
rect 1276 1378 1319 1392
rect 1343 1389 1350 1396
rect 1353 1392 1420 1416
rect 1452 1416 1624 1418
rect 1422 1394 1450 1398
rect 1452 1394 1532 1416
rect 1553 1414 1568 1416
rect 1422 1392 1532 1394
rect 1353 1388 1532 1392
rect 1326 1378 1356 1388
rect 1358 1378 1511 1388
rect 1519 1378 1549 1388
rect 1553 1378 1583 1392
rect 1611 1378 1624 1416
rect 1696 1422 1731 1430
rect 1696 1396 1697 1422
rect 1704 1396 1731 1422
rect 1639 1378 1669 1392
rect 1696 1388 1731 1396
rect 1733 1422 1774 1430
rect 1733 1396 1748 1422
rect 1755 1396 1774 1422
rect 1838 1418 1900 1430
rect 1912 1418 1987 1430
rect 2045 1418 2120 1430
rect 2132 1418 2163 1430
rect 2169 1418 2204 1430
rect 1838 1416 2000 1418
rect 1733 1388 1774 1396
rect 1856 1392 1869 1416
rect 1884 1414 1899 1416
rect 1696 1378 1697 1388
rect 1712 1378 1725 1388
rect 1739 1378 1740 1388
rect 1755 1378 1768 1388
rect 1783 1378 1813 1392
rect 1856 1378 1899 1392
rect 1923 1389 1930 1396
rect 1933 1392 2000 1416
rect 2032 1416 2204 1418
rect 2002 1394 2030 1398
rect 2032 1394 2112 1416
rect 2133 1414 2148 1416
rect 2002 1392 2112 1394
rect 1933 1388 2112 1392
rect 1906 1378 1936 1388
rect 1938 1378 2091 1388
rect 2099 1378 2129 1388
rect 2133 1378 2163 1392
rect 2191 1378 2204 1416
rect 2276 1422 2311 1430
rect 2276 1396 2277 1422
rect 2284 1396 2311 1422
rect 2219 1378 2249 1392
rect 2276 1388 2311 1396
rect 2313 1422 2354 1430
rect 2313 1396 2328 1422
rect 2335 1396 2354 1422
rect 2418 1418 2480 1430
rect 2492 1418 2567 1430
rect 2625 1418 2700 1430
rect 2712 1418 2743 1430
rect 2749 1418 2784 1430
rect 2418 1416 2580 1418
rect 2313 1388 2354 1396
rect 2436 1392 2449 1416
rect 2464 1414 2479 1416
rect 2276 1378 2277 1388
rect 2292 1378 2305 1388
rect 2319 1378 2320 1388
rect 2335 1378 2348 1388
rect 2363 1378 2393 1392
rect 2436 1378 2479 1392
rect 2503 1389 2510 1396
rect 2513 1392 2580 1416
rect 2612 1416 2784 1418
rect 2582 1394 2610 1398
rect 2612 1394 2692 1416
rect 2713 1414 2728 1416
rect 2582 1392 2692 1394
rect 2513 1388 2692 1392
rect 2486 1378 2516 1388
rect 2518 1378 2671 1388
rect 2679 1378 2709 1388
rect 2713 1378 2743 1392
rect 2771 1378 2784 1416
rect 2856 1422 2891 1430
rect 2856 1396 2857 1422
rect 2864 1396 2891 1422
rect 2799 1378 2829 1392
rect 2856 1388 2891 1396
rect 2893 1422 2934 1430
rect 2893 1396 2908 1422
rect 2915 1396 2934 1422
rect 2998 1418 3060 1430
rect 3072 1418 3147 1430
rect 3205 1418 3280 1430
rect 3292 1418 3323 1430
rect 3329 1418 3364 1430
rect 2998 1416 3160 1418
rect 2893 1388 2934 1396
rect 3016 1392 3029 1416
rect 3044 1414 3059 1416
rect 2856 1378 2857 1388
rect 2872 1378 2885 1388
rect 2899 1378 2900 1388
rect 2915 1378 2928 1388
rect 2943 1378 2973 1392
rect 3016 1378 3059 1392
rect 3083 1389 3090 1396
rect 3093 1392 3160 1416
rect 3192 1416 3364 1418
rect 3162 1394 3190 1398
rect 3192 1394 3272 1416
rect 3293 1414 3308 1416
rect 3162 1392 3272 1394
rect 3093 1388 3272 1392
rect 3066 1378 3096 1388
rect 3098 1378 3251 1388
rect 3259 1378 3289 1388
rect 3293 1378 3323 1392
rect 3351 1378 3364 1416
rect 3436 1422 3471 1430
rect 3436 1396 3437 1422
rect 3444 1396 3471 1422
rect 3379 1378 3409 1392
rect 3436 1388 3471 1396
rect 3473 1422 3514 1430
rect 3473 1396 3488 1422
rect 3495 1396 3514 1422
rect 3578 1418 3640 1430
rect 3652 1418 3727 1430
rect 3785 1418 3860 1430
rect 3872 1418 3903 1430
rect 3909 1418 3944 1430
rect 3578 1416 3740 1418
rect 3473 1388 3514 1396
rect 3596 1392 3609 1416
rect 3624 1414 3639 1416
rect 3436 1378 3437 1388
rect 3452 1378 3465 1388
rect 3479 1378 3480 1388
rect 3495 1378 3508 1388
rect 3523 1378 3553 1392
rect 3596 1378 3639 1392
rect 3663 1389 3670 1396
rect 3673 1392 3740 1416
rect 3772 1416 3944 1418
rect 3742 1394 3770 1398
rect 3772 1394 3852 1416
rect 3873 1414 3888 1416
rect 3742 1392 3852 1394
rect 3673 1388 3852 1392
rect 3646 1378 3676 1388
rect 3678 1378 3831 1388
rect 3839 1378 3869 1388
rect 3873 1378 3903 1392
rect 3931 1378 3944 1416
rect 4016 1422 4051 1430
rect 4016 1396 4017 1422
rect 4024 1396 4051 1422
rect 3959 1378 3989 1392
rect 4016 1388 4051 1396
rect 4053 1422 4094 1430
rect 4053 1396 4068 1422
rect 4075 1396 4094 1422
rect 4158 1418 4220 1430
rect 4232 1418 4307 1430
rect 4365 1418 4440 1430
rect 4452 1418 4483 1430
rect 4489 1418 4524 1430
rect 4158 1416 4320 1418
rect 4053 1388 4094 1396
rect 4176 1392 4189 1416
rect 4204 1414 4219 1416
rect 4016 1378 4017 1388
rect 4032 1378 4045 1388
rect 4059 1378 4060 1388
rect 4075 1378 4088 1388
rect 4103 1378 4133 1392
rect 4176 1378 4219 1392
rect 4243 1389 4250 1396
rect 4253 1392 4320 1416
rect 4352 1416 4524 1418
rect 4322 1394 4350 1398
rect 4352 1394 4432 1416
rect 4453 1414 4468 1416
rect 4322 1392 4432 1394
rect 4253 1388 4432 1392
rect 4226 1378 4256 1388
rect 4258 1378 4411 1388
rect 4419 1378 4449 1388
rect 4453 1378 4483 1392
rect 4511 1378 4524 1416
rect 4596 1422 4631 1430
rect 4596 1396 4597 1422
rect 4604 1396 4631 1422
rect 4539 1378 4569 1392
rect 4596 1388 4631 1396
rect 4596 1378 4597 1388
rect 4612 1378 4625 1388
rect -1 1372 4625 1378
rect 0 1364 4625 1372
rect 15 1334 28 1364
rect 43 1346 73 1364
rect 116 1350 130 1364
rect 166 1350 386 1364
rect 117 1348 130 1350
rect 83 1336 98 1348
rect 80 1334 102 1336
rect 107 1334 137 1348
rect 198 1346 351 1350
rect 180 1334 372 1346
rect 415 1334 445 1348
rect 451 1334 464 1364
rect 479 1346 509 1364
rect 552 1334 565 1364
rect 595 1334 608 1364
rect 623 1346 653 1364
rect 696 1350 710 1364
rect 746 1350 966 1364
rect 697 1348 710 1350
rect 663 1336 678 1348
rect 660 1334 682 1336
rect 687 1334 717 1348
rect 778 1346 931 1350
rect 760 1334 952 1346
rect 995 1334 1025 1348
rect 1031 1334 1044 1364
rect 1059 1346 1089 1364
rect 1132 1334 1145 1364
rect 1175 1334 1188 1364
rect 1203 1346 1233 1364
rect 1276 1350 1290 1364
rect 1326 1350 1546 1364
rect 1277 1348 1290 1350
rect 1243 1336 1258 1348
rect 1240 1334 1262 1336
rect 1267 1334 1297 1348
rect 1358 1346 1511 1350
rect 1340 1334 1532 1346
rect 1575 1334 1605 1348
rect 1611 1334 1624 1364
rect 1639 1346 1669 1364
rect 1712 1334 1725 1364
rect 1755 1334 1768 1364
rect 1783 1346 1813 1364
rect 1856 1350 1870 1364
rect 1906 1350 2126 1364
rect 1857 1348 1870 1350
rect 1823 1336 1838 1348
rect 1820 1334 1842 1336
rect 1847 1334 1877 1348
rect 1938 1346 2091 1350
rect 1920 1334 2112 1346
rect 2155 1334 2185 1348
rect 2191 1334 2204 1364
rect 2219 1346 2249 1364
rect 2292 1334 2305 1364
rect 2335 1334 2348 1364
rect 2363 1346 2393 1364
rect 2436 1350 2450 1364
rect 2486 1350 2706 1364
rect 2437 1348 2450 1350
rect 2403 1336 2418 1348
rect 2400 1334 2422 1336
rect 2427 1334 2457 1348
rect 2518 1346 2671 1350
rect 2500 1334 2692 1346
rect 2735 1334 2765 1348
rect 2771 1334 2784 1364
rect 2799 1346 2829 1364
rect 2872 1334 2885 1364
rect 2915 1334 2928 1364
rect 2943 1346 2973 1364
rect 3016 1350 3030 1364
rect 3066 1350 3286 1364
rect 3017 1348 3030 1350
rect 2983 1336 2998 1348
rect 2980 1334 3002 1336
rect 3007 1334 3037 1348
rect 3098 1346 3251 1350
rect 3080 1334 3272 1346
rect 3315 1334 3345 1348
rect 3351 1334 3364 1364
rect 3379 1346 3409 1364
rect 3452 1334 3465 1364
rect 3495 1334 3508 1364
rect 3523 1346 3553 1364
rect 3596 1350 3610 1364
rect 3646 1350 3866 1364
rect 3597 1348 3610 1350
rect 3563 1336 3578 1348
rect 3560 1334 3582 1336
rect 3587 1334 3617 1348
rect 3678 1346 3831 1350
rect 3660 1334 3852 1346
rect 3895 1334 3925 1348
rect 3931 1334 3944 1364
rect 3959 1346 3989 1364
rect 4032 1334 4045 1364
rect 4075 1334 4088 1364
rect 4103 1346 4133 1364
rect 4176 1350 4190 1364
rect 4226 1350 4446 1364
rect 4177 1348 4190 1350
rect 4143 1336 4158 1348
rect 4140 1334 4162 1336
rect 4167 1334 4197 1348
rect 4258 1346 4411 1350
rect 4240 1334 4432 1346
rect 4475 1334 4505 1348
rect 4511 1334 4524 1364
rect 4539 1346 4569 1364
rect 4612 1334 4625 1364
rect 0 1320 4625 1334
rect 15 1216 28 1320
rect 73 1298 74 1308
rect 89 1298 102 1308
rect 73 1294 102 1298
rect 107 1294 137 1320
rect 155 1306 171 1308
rect 243 1306 296 1320
rect 244 1304 308 1306
rect 351 1304 366 1320
rect 415 1317 445 1320
rect 415 1314 451 1317
rect 381 1306 397 1308
rect 155 1294 170 1298
rect 73 1292 170 1294
rect 198 1292 366 1304
rect 382 1294 397 1298
rect 415 1295 454 1314
rect 473 1308 480 1309
rect 479 1301 480 1308
rect 463 1298 464 1301
rect 479 1298 492 1301
rect 415 1294 445 1295
rect 454 1294 460 1295
rect 463 1294 492 1298
rect 382 1293 492 1294
rect 382 1292 498 1293
rect 57 1284 108 1292
rect 57 1272 82 1284
rect 89 1272 108 1284
rect 139 1284 189 1292
rect 139 1276 155 1284
rect 162 1282 189 1284
rect 198 1282 419 1292
rect 162 1272 419 1282
rect 448 1284 498 1292
rect 448 1275 464 1284
rect 57 1264 108 1272
rect 155 1264 419 1272
rect 445 1272 464 1275
rect 471 1272 498 1284
rect 445 1264 498 1272
rect 73 1256 74 1264
rect 89 1256 102 1264
rect 73 1248 89 1256
rect 70 1241 89 1244
rect 70 1232 92 1241
rect 43 1222 92 1232
rect 43 1216 73 1222
rect 92 1217 97 1222
rect 15 1200 89 1216
rect 107 1208 137 1264
rect 172 1254 380 1264
rect 415 1260 460 1264
rect 463 1263 464 1264
rect 479 1263 492 1264
rect 198 1224 387 1254
rect 213 1221 387 1224
rect 206 1218 387 1221
rect 15 1198 28 1200
rect 43 1198 77 1200
rect 15 1182 89 1198
rect 116 1194 129 1208
rect 144 1194 160 1210
rect 206 1205 217 1218
rect -1 1160 0 1176
rect 15 1160 28 1182
rect 43 1160 73 1182
rect 116 1178 178 1194
rect 206 1187 217 1203
rect 222 1198 232 1218
rect 242 1198 256 1218
rect 259 1205 268 1218
rect 284 1205 293 1218
rect 222 1187 256 1198
rect 259 1187 268 1203
rect 284 1187 293 1203
rect 300 1198 310 1218
rect 320 1198 334 1218
rect 335 1205 346 1218
rect 300 1187 334 1198
rect 335 1187 346 1203
rect 392 1194 408 1210
rect 415 1208 445 1260
rect 479 1256 480 1263
rect 464 1248 480 1256
rect 451 1216 464 1235
rect 479 1216 509 1232
rect 451 1200 525 1216
rect 451 1198 464 1200
rect 479 1198 513 1200
rect 116 1176 129 1178
rect 144 1176 178 1178
rect 116 1160 178 1176
rect 222 1171 238 1174
rect 300 1171 330 1182
rect 378 1178 424 1194
rect 451 1182 525 1198
rect 378 1176 412 1178
rect 377 1160 424 1176
rect 451 1160 464 1182
rect 479 1160 509 1182
rect 536 1160 537 1176
rect 552 1160 565 1320
rect 595 1216 608 1320
rect 653 1298 654 1308
rect 669 1298 682 1308
rect 653 1294 682 1298
rect 687 1294 717 1320
rect 735 1306 751 1308
rect 823 1306 876 1320
rect 824 1304 888 1306
rect 931 1304 946 1320
rect 995 1317 1025 1320
rect 995 1314 1031 1317
rect 961 1306 977 1308
rect 735 1294 750 1298
rect 653 1292 750 1294
rect 778 1292 946 1304
rect 962 1294 977 1298
rect 995 1295 1034 1314
rect 1053 1308 1060 1309
rect 1059 1301 1060 1308
rect 1043 1298 1044 1301
rect 1059 1298 1072 1301
rect 995 1294 1025 1295
rect 1034 1294 1040 1295
rect 1043 1294 1072 1298
rect 962 1293 1072 1294
rect 962 1292 1078 1293
rect 637 1284 688 1292
rect 637 1272 662 1284
rect 669 1272 688 1284
rect 719 1284 769 1292
rect 719 1276 735 1284
rect 742 1282 769 1284
rect 778 1282 999 1292
rect 742 1272 999 1282
rect 1028 1284 1078 1292
rect 1028 1275 1044 1284
rect 637 1264 688 1272
rect 735 1264 999 1272
rect 1025 1272 1044 1275
rect 1051 1272 1078 1284
rect 1025 1264 1078 1272
rect 653 1256 654 1264
rect 669 1256 682 1264
rect 653 1248 669 1256
rect 650 1241 669 1244
rect 650 1232 672 1241
rect 623 1222 672 1232
rect 623 1216 653 1222
rect 672 1217 677 1222
rect 595 1200 669 1216
rect 687 1208 717 1264
rect 752 1254 960 1264
rect 995 1260 1040 1264
rect 1043 1263 1044 1264
rect 1059 1263 1072 1264
rect 778 1224 967 1254
rect 793 1221 967 1224
rect 786 1218 967 1221
rect 595 1198 608 1200
rect 623 1198 657 1200
rect 595 1182 669 1198
rect 696 1194 709 1208
rect 724 1194 740 1210
rect 786 1205 797 1218
rect 579 1160 580 1176
rect 595 1160 608 1182
rect 623 1160 653 1182
rect 696 1178 758 1194
rect 786 1187 797 1203
rect 802 1198 812 1218
rect 822 1198 836 1218
rect 839 1205 848 1218
rect 864 1205 873 1218
rect 802 1187 836 1198
rect 839 1187 848 1203
rect 864 1187 873 1203
rect 880 1198 890 1218
rect 900 1198 914 1218
rect 915 1205 926 1218
rect 880 1187 914 1198
rect 915 1187 926 1203
rect 972 1194 988 1210
rect 995 1208 1025 1260
rect 1059 1256 1060 1263
rect 1044 1248 1060 1256
rect 1031 1216 1044 1235
rect 1059 1216 1089 1232
rect 1031 1200 1105 1216
rect 1031 1198 1044 1200
rect 1059 1198 1093 1200
rect 696 1176 709 1178
rect 724 1176 758 1178
rect 696 1160 758 1176
rect 802 1171 818 1174
rect 880 1171 910 1182
rect 958 1178 1004 1194
rect 1031 1182 1105 1198
rect 958 1176 992 1178
rect 957 1160 1004 1176
rect 1031 1160 1044 1182
rect 1059 1160 1089 1182
rect 1116 1160 1117 1176
rect 1132 1160 1145 1320
rect 1175 1216 1188 1320
rect 1233 1298 1234 1308
rect 1249 1298 1262 1308
rect 1233 1294 1262 1298
rect 1267 1294 1297 1320
rect 1315 1306 1331 1308
rect 1403 1306 1456 1320
rect 1404 1304 1468 1306
rect 1511 1304 1526 1320
rect 1575 1317 1605 1320
rect 1575 1314 1611 1317
rect 1541 1306 1557 1308
rect 1315 1294 1330 1298
rect 1233 1292 1330 1294
rect 1358 1292 1526 1304
rect 1542 1294 1557 1298
rect 1575 1295 1614 1314
rect 1633 1308 1640 1309
rect 1639 1301 1640 1308
rect 1623 1298 1624 1301
rect 1639 1298 1652 1301
rect 1575 1294 1605 1295
rect 1614 1294 1620 1295
rect 1623 1294 1652 1298
rect 1542 1293 1652 1294
rect 1542 1292 1658 1293
rect 1217 1284 1268 1292
rect 1217 1272 1242 1284
rect 1249 1272 1268 1284
rect 1299 1284 1349 1292
rect 1299 1276 1315 1284
rect 1322 1282 1349 1284
rect 1358 1282 1579 1292
rect 1322 1272 1579 1282
rect 1608 1284 1658 1292
rect 1608 1275 1624 1284
rect 1217 1264 1268 1272
rect 1315 1264 1579 1272
rect 1605 1272 1624 1275
rect 1631 1272 1658 1284
rect 1605 1264 1658 1272
rect 1233 1256 1234 1264
rect 1249 1256 1262 1264
rect 1233 1248 1249 1256
rect 1230 1241 1249 1244
rect 1230 1232 1252 1241
rect 1203 1222 1252 1232
rect 1203 1216 1233 1222
rect 1252 1217 1257 1222
rect 1175 1200 1249 1216
rect 1267 1208 1297 1264
rect 1332 1254 1540 1264
rect 1575 1260 1620 1264
rect 1623 1263 1624 1264
rect 1639 1263 1652 1264
rect 1358 1224 1547 1254
rect 1373 1221 1547 1224
rect 1366 1218 1547 1221
rect 1175 1198 1188 1200
rect 1203 1198 1237 1200
rect 1175 1182 1249 1198
rect 1276 1194 1289 1208
rect 1304 1194 1320 1210
rect 1366 1205 1377 1218
rect 1159 1160 1160 1176
rect 1175 1160 1188 1182
rect 1203 1160 1233 1182
rect 1276 1178 1338 1194
rect 1366 1187 1377 1203
rect 1382 1198 1392 1218
rect 1402 1198 1416 1218
rect 1419 1205 1428 1218
rect 1444 1205 1453 1218
rect 1382 1187 1416 1198
rect 1419 1187 1428 1203
rect 1444 1187 1453 1203
rect 1460 1198 1470 1218
rect 1480 1198 1494 1218
rect 1495 1205 1506 1218
rect 1460 1187 1494 1198
rect 1495 1187 1506 1203
rect 1552 1194 1568 1210
rect 1575 1208 1605 1260
rect 1639 1256 1640 1263
rect 1624 1248 1640 1256
rect 1611 1216 1624 1235
rect 1639 1216 1669 1232
rect 1611 1200 1685 1216
rect 1611 1198 1624 1200
rect 1639 1198 1673 1200
rect 1276 1176 1289 1178
rect 1304 1176 1338 1178
rect 1276 1160 1338 1176
rect 1382 1171 1398 1174
rect 1460 1171 1490 1182
rect 1538 1178 1584 1194
rect 1611 1182 1685 1198
rect 1538 1176 1572 1178
rect 1537 1160 1584 1176
rect 1611 1160 1624 1182
rect 1639 1160 1669 1182
rect 1696 1160 1697 1176
rect 1712 1160 1725 1320
rect 1755 1216 1768 1320
rect 1813 1298 1814 1308
rect 1829 1298 1842 1308
rect 1813 1294 1842 1298
rect 1847 1294 1877 1320
rect 1895 1306 1911 1308
rect 1983 1306 2036 1320
rect 1984 1304 2048 1306
rect 2091 1304 2106 1320
rect 2155 1317 2185 1320
rect 2155 1314 2191 1317
rect 2121 1306 2137 1308
rect 1895 1294 1910 1298
rect 1813 1292 1910 1294
rect 1938 1292 2106 1304
rect 2122 1294 2137 1298
rect 2155 1295 2194 1314
rect 2213 1308 2220 1309
rect 2219 1301 2220 1308
rect 2203 1298 2204 1301
rect 2219 1298 2232 1301
rect 2155 1294 2185 1295
rect 2194 1294 2200 1295
rect 2203 1294 2232 1298
rect 2122 1293 2232 1294
rect 2122 1292 2238 1293
rect 1797 1284 1848 1292
rect 1797 1272 1822 1284
rect 1829 1272 1848 1284
rect 1879 1284 1929 1292
rect 1879 1276 1895 1284
rect 1902 1282 1929 1284
rect 1938 1282 2159 1292
rect 1902 1272 2159 1282
rect 2188 1284 2238 1292
rect 2188 1275 2204 1284
rect 1797 1264 1848 1272
rect 1895 1264 2159 1272
rect 2185 1272 2204 1275
rect 2211 1272 2238 1284
rect 2185 1264 2238 1272
rect 1813 1256 1814 1264
rect 1829 1256 1842 1264
rect 1813 1248 1829 1256
rect 1810 1241 1829 1244
rect 1810 1232 1832 1241
rect 1783 1222 1832 1232
rect 1783 1216 1813 1222
rect 1832 1217 1837 1222
rect 1755 1200 1829 1216
rect 1847 1208 1877 1264
rect 1912 1254 2120 1264
rect 2155 1260 2200 1264
rect 2203 1263 2204 1264
rect 2219 1263 2232 1264
rect 1938 1224 2127 1254
rect 1953 1221 2127 1224
rect 1946 1218 2127 1221
rect 1755 1198 1768 1200
rect 1783 1198 1817 1200
rect 1755 1182 1829 1198
rect 1856 1194 1869 1208
rect 1884 1194 1900 1210
rect 1946 1205 1957 1218
rect 1739 1160 1740 1176
rect 1755 1160 1768 1182
rect 1783 1160 1813 1182
rect 1856 1178 1918 1194
rect 1946 1187 1957 1203
rect 1962 1198 1972 1218
rect 1982 1198 1996 1218
rect 1999 1205 2008 1218
rect 2024 1205 2033 1218
rect 1962 1187 1996 1198
rect 1999 1187 2008 1203
rect 2024 1187 2033 1203
rect 2040 1198 2050 1218
rect 2060 1198 2074 1218
rect 2075 1205 2086 1218
rect 2040 1187 2074 1198
rect 2075 1187 2086 1203
rect 2132 1194 2148 1210
rect 2155 1208 2185 1260
rect 2219 1256 2220 1263
rect 2204 1248 2220 1256
rect 2191 1216 2204 1235
rect 2219 1216 2249 1232
rect 2191 1200 2265 1216
rect 2191 1198 2204 1200
rect 2219 1198 2253 1200
rect 1856 1176 1869 1178
rect 1884 1176 1918 1178
rect 1856 1160 1918 1176
rect 1962 1171 1978 1174
rect 2040 1171 2070 1182
rect 2118 1178 2164 1194
rect 2191 1182 2265 1198
rect 2118 1176 2152 1178
rect 2117 1160 2164 1176
rect 2191 1160 2204 1182
rect 2219 1160 2249 1182
rect 2276 1160 2277 1176
rect 2292 1160 2305 1320
rect 2335 1216 2348 1320
rect 2393 1298 2394 1308
rect 2409 1298 2422 1308
rect 2393 1294 2422 1298
rect 2427 1294 2457 1320
rect 2475 1306 2491 1308
rect 2563 1306 2616 1320
rect 2564 1304 2628 1306
rect 2671 1304 2686 1320
rect 2735 1317 2765 1320
rect 2735 1314 2771 1317
rect 2701 1306 2717 1308
rect 2475 1294 2490 1298
rect 2393 1292 2490 1294
rect 2518 1292 2686 1304
rect 2702 1294 2717 1298
rect 2735 1295 2774 1314
rect 2793 1308 2800 1309
rect 2799 1301 2800 1308
rect 2783 1298 2784 1301
rect 2799 1298 2812 1301
rect 2735 1294 2765 1295
rect 2774 1294 2780 1295
rect 2783 1294 2812 1298
rect 2702 1293 2812 1294
rect 2702 1292 2818 1293
rect 2377 1284 2428 1292
rect 2377 1272 2402 1284
rect 2409 1272 2428 1284
rect 2459 1284 2509 1292
rect 2459 1276 2475 1284
rect 2482 1282 2509 1284
rect 2518 1282 2739 1292
rect 2482 1272 2739 1282
rect 2768 1284 2818 1292
rect 2768 1275 2784 1284
rect 2377 1264 2428 1272
rect 2475 1264 2739 1272
rect 2765 1272 2784 1275
rect 2791 1272 2818 1284
rect 2765 1264 2818 1272
rect 2393 1256 2394 1264
rect 2409 1256 2422 1264
rect 2393 1248 2409 1256
rect 2390 1241 2409 1244
rect 2390 1232 2412 1241
rect 2363 1222 2412 1232
rect 2363 1216 2393 1222
rect 2412 1217 2417 1222
rect 2335 1200 2409 1216
rect 2427 1208 2457 1264
rect 2492 1254 2700 1264
rect 2735 1260 2780 1264
rect 2783 1263 2784 1264
rect 2799 1263 2812 1264
rect 2518 1224 2707 1254
rect 2533 1221 2707 1224
rect 2526 1218 2707 1221
rect 2335 1198 2348 1200
rect 2363 1198 2397 1200
rect 2335 1182 2409 1198
rect 2436 1194 2449 1208
rect 2464 1194 2480 1210
rect 2526 1205 2537 1218
rect 2319 1160 2320 1176
rect 2335 1160 2348 1182
rect 2363 1160 2393 1182
rect 2436 1178 2498 1194
rect 2526 1187 2537 1203
rect 2542 1198 2552 1218
rect 2562 1198 2576 1218
rect 2579 1205 2588 1218
rect 2604 1205 2613 1218
rect 2542 1187 2576 1198
rect 2579 1187 2588 1203
rect 2604 1187 2613 1203
rect 2620 1198 2630 1218
rect 2640 1198 2654 1218
rect 2655 1205 2666 1218
rect 2620 1187 2654 1198
rect 2655 1187 2666 1203
rect 2712 1194 2728 1210
rect 2735 1208 2765 1260
rect 2799 1256 2800 1263
rect 2784 1248 2800 1256
rect 2771 1216 2784 1235
rect 2799 1216 2829 1232
rect 2771 1200 2845 1216
rect 2771 1198 2784 1200
rect 2799 1198 2833 1200
rect 2436 1176 2449 1178
rect 2464 1176 2498 1178
rect 2436 1160 2498 1176
rect 2542 1171 2558 1174
rect 2620 1171 2650 1182
rect 2698 1178 2744 1194
rect 2771 1182 2845 1198
rect 2698 1176 2732 1178
rect 2697 1160 2744 1176
rect 2771 1160 2784 1182
rect 2799 1160 2829 1182
rect 2856 1160 2857 1176
rect 2872 1160 2885 1320
rect 2915 1216 2928 1320
rect 2973 1298 2974 1308
rect 2989 1298 3002 1308
rect 2973 1294 3002 1298
rect 3007 1294 3037 1320
rect 3055 1306 3071 1308
rect 3143 1306 3196 1320
rect 3144 1304 3208 1306
rect 3251 1304 3266 1320
rect 3315 1317 3345 1320
rect 3315 1314 3351 1317
rect 3281 1306 3297 1308
rect 3055 1294 3070 1298
rect 2973 1292 3070 1294
rect 3098 1292 3266 1304
rect 3282 1294 3297 1298
rect 3315 1295 3354 1314
rect 3373 1308 3380 1309
rect 3379 1301 3380 1308
rect 3363 1298 3364 1301
rect 3379 1298 3392 1301
rect 3315 1294 3345 1295
rect 3354 1294 3360 1295
rect 3363 1294 3392 1298
rect 3282 1293 3392 1294
rect 3282 1292 3398 1293
rect 2957 1284 3008 1292
rect 2957 1272 2982 1284
rect 2989 1272 3008 1284
rect 3039 1284 3089 1292
rect 3039 1276 3055 1284
rect 3062 1282 3089 1284
rect 3098 1282 3319 1292
rect 3062 1272 3319 1282
rect 3348 1284 3398 1292
rect 3348 1275 3364 1284
rect 2957 1264 3008 1272
rect 3055 1264 3319 1272
rect 3345 1272 3364 1275
rect 3371 1272 3398 1284
rect 3345 1264 3398 1272
rect 2973 1256 2974 1264
rect 2989 1256 3002 1264
rect 2973 1248 2989 1256
rect 2970 1241 2989 1244
rect 2970 1232 2992 1241
rect 2943 1222 2992 1232
rect 2943 1216 2973 1222
rect 2992 1217 2997 1222
rect 2915 1200 2989 1216
rect 3007 1208 3037 1264
rect 3072 1254 3280 1264
rect 3315 1260 3360 1264
rect 3363 1263 3364 1264
rect 3379 1263 3392 1264
rect 3098 1224 3287 1254
rect 3113 1221 3287 1224
rect 3106 1218 3287 1221
rect 2915 1198 2928 1200
rect 2943 1198 2977 1200
rect 2915 1182 2989 1198
rect 3016 1194 3029 1208
rect 3044 1194 3060 1210
rect 3106 1205 3117 1218
rect 2899 1160 2900 1176
rect 2915 1160 2928 1182
rect 2943 1160 2973 1182
rect 3016 1178 3078 1194
rect 3106 1187 3117 1203
rect 3122 1198 3132 1218
rect 3142 1198 3156 1218
rect 3159 1205 3168 1218
rect 3184 1205 3193 1218
rect 3122 1187 3156 1198
rect 3159 1187 3168 1203
rect 3184 1187 3193 1203
rect 3200 1198 3210 1218
rect 3220 1198 3234 1218
rect 3235 1205 3246 1218
rect 3200 1187 3234 1198
rect 3235 1187 3246 1203
rect 3292 1194 3308 1210
rect 3315 1208 3345 1260
rect 3379 1256 3380 1263
rect 3364 1248 3380 1256
rect 3351 1216 3364 1235
rect 3379 1216 3409 1232
rect 3351 1200 3425 1216
rect 3351 1198 3364 1200
rect 3379 1198 3413 1200
rect 3016 1176 3029 1178
rect 3044 1176 3078 1178
rect 3016 1160 3078 1176
rect 3122 1171 3138 1174
rect 3200 1171 3230 1182
rect 3278 1178 3324 1194
rect 3351 1182 3425 1198
rect 3278 1176 3312 1178
rect 3277 1160 3324 1176
rect 3351 1160 3364 1182
rect 3379 1160 3409 1182
rect 3436 1160 3437 1176
rect 3452 1160 3465 1320
rect 3495 1216 3508 1320
rect 3553 1298 3554 1308
rect 3569 1298 3582 1308
rect 3553 1294 3582 1298
rect 3587 1294 3617 1320
rect 3635 1306 3651 1308
rect 3723 1306 3776 1320
rect 3724 1304 3788 1306
rect 3831 1304 3846 1320
rect 3895 1317 3925 1320
rect 3895 1314 3931 1317
rect 3861 1306 3877 1308
rect 3635 1294 3650 1298
rect 3553 1292 3650 1294
rect 3678 1292 3846 1304
rect 3862 1294 3877 1298
rect 3895 1295 3934 1314
rect 3953 1308 3960 1309
rect 3959 1301 3960 1308
rect 3943 1298 3944 1301
rect 3959 1298 3972 1301
rect 3895 1294 3925 1295
rect 3934 1294 3940 1295
rect 3943 1294 3972 1298
rect 3862 1293 3972 1294
rect 3862 1292 3978 1293
rect 3537 1284 3588 1292
rect 3537 1272 3562 1284
rect 3569 1272 3588 1284
rect 3619 1284 3669 1292
rect 3619 1276 3635 1284
rect 3642 1282 3669 1284
rect 3678 1282 3899 1292
rect 3642 1272 3899 1282
rect 3928 1284 3978 1292
rect 3928 1275 3944 1284
rect 3537 1264 3588 1272
rect 3635 1264 3899 1272
rect 3925 1272 3944 1275
rect 3951 1272 3978 1284
rect 3925 1264 3978 1272
rect 3553 1256 3554 1264
rect 3569 1256 3582 1264
rect 3553 1248 3569 1256
rect 3550 1241 3569 1244
rect 3550 1232 3572 1241
rect 3523 1222 3572 1232
rect 3523 1216 3553 1222
rect 3572 1217 3577 1222
rect 3495 1200 3569 1216
rect 3587 1208 3617 1264
rect 3652 1254 3860 1264
rect 3895 1260 3940 1264
rect 3943 1263 3944 1264
rect 3959 1263 3972 1264
rect 3678 1224 3867 1254
rect 3693 1221 3867 1224
rect 3686 1218 3867 1221
rect 3495 1198 3508 1200
rect 3523 1198 3557 1200
rect 3495 1182 3569 1198
rect 3596 1194 3609 1208
rect 3624 1194 3640 1210
rect 3686 1205 3697 1218
rect 3479 1160 3480 1176
rect 3495 1160 3508 1182
rect 3523 1160 3553 1182
rect 3596 1178 3658 1194
rect 3686 1187 3697 1203
rect 3702 1198 3712 1218
rect 3722 1198 3736 1218
rect 3739 1205 3748 1218
rect 3764 1205 3773 1218
rect 3702 1187 3736 1198
rect 3739 1187 3748 1203
rect 3764 1187 3773 1203
rect 3780 1198 3790 1218
rect 3800 1198 3814 1218
rect 3815 1205 3826 1218
rect 3780 1187 3814 1198
rect 3815 1187 3826 1203
rect 3872 1194 3888 1210
rect 3895 1208 3925 1260
rect 3959 1256 3960 1263
rect 3944 1248 3960 1256
rect 3931 1216 3944 1235
rect 3959 1216 3989 1232
rect 3931 1200 4005 1216
rect 3931 1198 3944 1200
rect 3959 1198 3993 1200
rect 3596 1176 3609 1178
rect 3624 1176 3658 1178
rect 3596 1160 3658 1176
rect 3702 1171 3718 1174
rect 3780 1171 3810 1182
rect 3858 1178 3904 1194
rect 3931 1182 4005 1198
rect 3858 1176 3892 1178
rect 3857 1160 3904 1176
rect 3931 1160 3944 1182
rect 3959 1160 3989 1182
rect 4016 1160 4017 1176
rect 4032 1160 4045 1320
rect 4075 1216 4088 1320
rect 4133 1298 4134 1308
rect 4149 1298 4162 1308
rect 4133 1294 4162 1298
rect 4167 1294 4197 1320
rect 4215 1306 4231 1308
rect 4303 1306 4356 1320
rect 4304 1304 4368 1306
rect 4411 1304 4426 1320
rect 4475 1317 4505 1320
rect 4475 1314 4511 1317
rect 4441 1306 4457 1308
rect 4215 1294 4230 1298
rect 4133 1292 4230 1294
rect 4258 1292 4426 1304
rect 4442 1294 4457 1298
rect 4475 1295 4514 1314
rect 4533 1308 4540 1309
rect 4539 1301 4540 1308
rect 4523 1298 4524 1301
rect 4539 1298 4552 1301
rect 4475 1294 4505 1295
rect 4514 1294 4520 1295
rect 4523 1294 4552 1298
rect 4442 1293 4552 1294
rect 4442 1292 4558 1293
rect 4117 1284 4168 1292
rect 4117 1272 4142 1284
rect 4149 1272 4168 1284
rect 4199 1284 4249 1292
rect 4199 1276 4215 1284
rect 4222 1282 4249 1284
rect 4258 1282 4479 1292
rect 4222 1272 4479 1282
rect 4508 1284 4558 1292
rect 4508 1275 4524 1284
rect 4117 1264 4168 1272
rect 4215 1264 4479 1272
rect 4505 1272 4524 1275
rect 4531 1272 4558 1284
rect 4505 1264 4558 1272
rect 4133 1256 4134 1264
rect 4149 1256 4162 1264
rect 4133 1248 4149 1256
rect 4130 1241 4149 1244
rect 4130 1232 4152 1241
rect 4103 1222 4152 1232
rect 4103 1216 4133 1222
rect 4152 1217 4157 1222
rect 4075 1200 4149 1216
rect 4167 1208 4197 1264
rect 4232 1254 4440 1264
rect 4475 1260 4520 1264
rect 4523 1263 4524 1264
rect 4539 1263 4552 1264
rect 4258 1224 4447 1254
rect 4273 1221 4447 1224
rect 4266 1218 4447 1221
rect 4075 1198 4088 1200
rect 4103 1198 4137 1200
rect 4075 1182 4149 1198
rect 4176 1194 4189 1208
rect 4204 1194 4220 1210
rect 4266 1205 4277 1218
rect 4059 1160 4060 1176
rect 4075 1160 4088 1182
rect 4103 1160 4133 1182
rect 4176 1178 4238 1194
rect 4266 1187 4277 1203
rect 4282 1198 4292 1218
rect 4302 1198 4316 1218
rect 4319 1205 4328 1218
rect 4344 1205 4353 1218
rect 4282 1187 4316 1198
rect 4319 1187 4328 1203
rect 4344 1187 4353 1203
rect 4360 1198 4370 1218
rect 4380 1198 4394 1218
rect 4395 1205 4406 1218
rect 4360 1187 4394 1198
rect 4395 1187 4406 1203
rect 4452 1194 4468 1210
rect 4475 1208 4505 1260
rect 4539 1256 4540 1263
rect 4524 1248 4540 1256
rect 4511 1216 4524 1235
rect 4539 1216 4569 1232
rect 4511 1200 4585 1216
rect 4511 1198 4524 1200
rect 4539 1198 4573 1200
rect 4176 1176 4189 1178
rect 4204 1176 4238 1178
rect 4176 1160 4238 1176
rect 4282 1171 4298 1174
rect 4360 1171 4390 1182
rect 4438 1178 4484 1194
rect 4511 1182 4585 1198
rect 4438 1176 4472 1178
rect 4437 1160 4484 1176
rect 4511 1160 4524 1182
rect 4539 1160 4569 1182
rect 4596 1160 4597 1176
rect 4612 1160 4625 1320
rect -7 1152 34 1160
rect -7 1126 8 1152
rect 15 1126 34 1152
rect 98 1148 160 1160
rect 172 1148 247 1160
rect 305 1148 380 1160
rect 392 1148 423 1160
rect 429 1148 464 1160
rect 98 1146 260 1148
rect -7 1118 34 1126
rect 116 1122 129 1146
rect 144 1144 159 1146
rect -1 1108 0 1118
rect 15 1108 28 1118
rect 43 1108 73 1122
rect 116 1108 159 1122
rect 183 1119 190 1126
rect 193 1122 260 1146
rect 292 1146 464 1148
rect 262 1124 290 1128
rect 292 1124 372 1146
rect 393 1144 408 1146
rect 262 1122 372 1124
rect 193 1118 372 1122
rect 166 1108 196 1118
rect 198 1108 351 1118
rect 359 1108 389 1118
rect 393 1108 423 1122
rect 451 1108 464 1146
rect 536 1152 571 1160
rect 536 1126 537 1152
rect 544 1126 571 1152
rect 479 1108 509 1122
rect 536 1118 571 1126
rect 573 1152 614 1160
rect 573 1126 588 1152
rect 595 1126 614 1152
rect 678 1148 740 1160
rect 752 1148 827 1160
rect 885 1148 960 1160
rect 972 1148 1003 1160
rect 1009 1148 1044 1160
rect 678 1146 840 1148
rect 573 1118 614 1126
rect 696 1122 709 1146
rect 724 1144 739 1146
rect 536 1108 537 1118
rect 552 1108 565 1118
rect 579 1108 580 1118
rect 595 1108 608 1118
rect 623 1108 653 1122
rect 696 1108 739 1122
rect 763 1119 770 1126
rect 773 1122 840 1146
rect 872 1146 1044 1148
rect 842 1124 870 1128
rect 872 1124 952 1146
rect 973 1144 988 1146
rect 842 1122 952 1124
rect 773 1118 952 1122
rect 746 1108 776 1118
rect 778 1108 931 1118
rect 939 1108 969 1118
rect 973 1108 1003 1122
rect 1031 1108 1044 1146
rect 1116 1152 1151 1160
rect 1116 1126 1117 1152
rect 1124 1126 1151 1152
rect 1059 1108 1089 1122
rect 1116 1118 1151 1126
rect 1153 1152 1194 1160
rect 1153 1126 1168 1152
rect 1175 1126 1194 1152
rect 1258 1148 1320 1160
rect 1332 1148 1407 1160
rect 1465 1148 1540 1160
rect 1552 1148 1583 1160
rect 1589 1148 1624 1160
rect 1258 1146 1420 1148
rect 1153 1118 1194 1126
rect 1276 1122 1289 1146
rect 1304 1144 1319 1146
rect 1116 1108 1117 1118
rect 1132 1108 1145 1118
rect 1159 1108 1160 1118
rect 1175 1108 1188 1118
rect 1203 1108 1233 1122
rect 1276 1108 1319 1122
rect 1343 1119 1350 1126
rect 1353 1122 1420 1146
rect 1452 1146 1624 1148
rect 1422 1124 1450 1128
rect 1452 1124 1532 1146
rect 1553 1144 1568 1146
rect 1422 1122 1532 1124
rect 1353 1118 1532 1122
rect 1326 1108 1356 1118
rect 1358 1108 1511 1118
rect 1519 1108 1549 1118
rect 1553 1108 1583 1122
rect 1611 1108 1624 1146
rect 1696 1152 1731 1160
rect 1696 1126 1697 1152
rect 1704 1126 1731 1152
rect 1639 1108 1669 1122
rect 1696 1118 1731 1126
rect 1733 1152 1774 1160
rect 1733 1126 1748 1152
rect 1755 1126 1774 1152
rect 1838 1148 1900 1160
rect 1912 1148 1987 1160
rect 2045 1148 2120 1160
rect 2132 1148 2163 1160
rect 2169 1148 2204 1160
rect 1838 1146 2000 1148
rect 1733 1118 1774 1126
rect 1856 1122 1869 1146
rect 1884 1144 1899 1146
rect 1696 1108 1697 1118
rect 1712 1108 1725 1118
rect 1739 1108 1740 1118
rect 1755 1108 1768 1118
rect 1783 1108 1813 1122
rect 1856 1108 1899 1122
rect 1923 1119 1930 1126
rect 1933 1122 2000 1146
rect 2032 1146 2204 1148
rect 2002 1124 2030 1128
rect 2032 1124 2112 1146
rect 2133 1144 2148 1146
rect 2002 1122 2112 1124
rect 1933 1118 2112 1122
rect 1906 1108 1936 1118
rect 1938 1108 2091 1118
rect 2099 1108 2129 1118
rect 2133 1108 2163 1122
rect 2191 1108 2204 1146
rect 2276 1152 2311 1160
rect 2276 1126 2277 1152
rect 2284 1126 2311 1152
rect 2219 1108 2249 1122
rect 2276 1118 2311 1126
rect 2313 1152 2354 1160
rect 2313 1126 2328 1152
rect 2335 1126 2354 1152
rect 2418 1148 2480 1160
rect 2492 1148 2567 1160
rect 2625 1148 2700 1160
rect 2712 1148 2743 1160
rect 2749 1148 2784 1160
rect 2418 1146 2580 1148
rect 2313 1118 2354 1126
rect 2436 1122 2449 1146
rect 2464 1144 2479 1146
rect 2276 1108 2277 1118
rect 2292 1108 2305 1118
rect 2319 1108 2320 1118
rect 2335 1108 2348 1118
rect 2363 1108 2393 1122
rect 2436 1108 2479 1122
rect 2503 1119 2510 1126
rect 2513 1122 2580 1146
rect 2612 1146 2784 1148
rect 2582 1124 2610 1128
rect 2612 1124 2692 1146
rect 2713 1144 2728 1146
rect 2582 1122 2692 1124
rect 2513 1118 2692 1122
rect 2486 1108 2516 1118
rect 2518 1108 2671 1118
rect 2679 1108 2709 1118
rect 2713 1108 2743 1122
rect 2771 1108 2784 1146
rect 2856 1152 2891 1160
rect 2856 1126 2857 1152
rect 2864 1126 2891 1152
rect 2799 1108 2829 1122
rect 2856 1118 2891 1126
rect 2893 1152 2934 1160
rect 2893 1126 2908 1152
rect 2915 1126 2934 1152
rect 2998 1148 3060 1160
rect 3072 1148 3147 1160
rect 3205 1148 3280 1160
rect 3292 1148 3323 1160
rect 3329 1148 3364 1160
rect 2998 1146 3160 1148
rect 2893 1118 2934 1126
rect 3016 1122 3029 1146
rect 3044 1144 3059 1146
rect 2856 1108 2857 1118
rect 2872 1108 2885 1118
rect 2899 1108 2900 1118
rect 2915 1108 2928 1118
rect 2943 1108 2973 1122
rect 3016 1108 3059 1122
rect 3083 1119 3090 1126
rect 3093 1122 3160 1146
rect 3192 1146 3364 1148
rect 3162 1124 3190 1128
rect 3192 1124 3272 1146
rect 3293 1144 3308 1146
rect 3162 1122 3272 1124
rect 3093 1118 3272 1122
rect 3066 1108 3096 1118
rect 3098 1108 3251 1118
rect 3259 1108 3289 1118
rect 3293 1108 3323 1122
rect 3351 1108 3364 1146
rect 3436 1152 3471 1160
rect 3436 1126 3437 1152
rect 3444 1126 3471 1152
rect 3379 1108 3409 1122
rect 3436 1118 3471 1126
rect 3473 1152 3514 1160
rect 3473 1126 3488 1152
rect 3495 1126 3514 1152
rect 3578 1148 3640 1160
rect 3652 1148 3727 1160
rect 3785 1148 3860 1160
rect 3872 1148 3903 1160
rect 3909 1148 3944 1160
rect 3578 1146 3740 1148
rect 3473 1118 3514 1126
rect 3596 1122 3609 1146
rect 3624 1144 3639 1146
rect 3436 1108 3437 1118
rect 3452 1108 3465 1118
rect 3479 1108 3480 1118
rect 3495 1108 3508 1118
rect 3523 1108 3553 1122
rect 3596 1108 3639 1122
rect 3663 1119 3670 1126
rect 3673 1122 3740 1146
rect 3772 1146 3944 1148
rect 3742 1124 3770 1128
rect 3772 1124 3852 1146
rect 3873 1144 3888 1146
rect 3742 1122 3852 1124
rect 3673 1118 3852 1122
rect 3646 1108 3676 1118
rect 3678 1108 3831 1118
rect 3839 1108 3869 1118
rect 3873 1108 3903 1122
rect 3931 1108 3944 1146
rect 4016 1152 4051 1160
rect 4016 1126 4017 1152
rect 4024 1126 4051 1152
rect 3959 1108 3989 1122
rect 4016 1118 4051 1126
rect 4053 1152 4094 1160
rect 4053 1126 4068 1152
rect 4075 1126 4094 1152
rect 4158 1148 4220 1160
rect 4232 1148 4307 1160
rect 4365 1148 4440 1160
rect 4452 1148 4483 1160
rect 4489 1148 4524 1160
rect 4158 1146 4320 1148
rect 4053 1118 4094 1126
rect 4176 1122 4189 1146
rect 4204 1144 4219 1146
rect 4016 1108 4017 1118
rect 4032 1108 4045 1118
rect 4059 1108 4060 1118
rect 4075 1108 4088 1118
rect 4103 1108 4133 1122
rect 4176 1108 4219 1122
rect 4243 1119 4250 1126
rect 4253 1122 4320 1146
rect 4352 1146 4524 1148
rect 4322 1124 4350 1128
rect 4352 1124 4432 1146
rect 4453 1144 4468 1146
rect 4322 1122 4432 1124
rect 4253 1118 4432 1122
rect 4226 1108 4256 1118
rect 4258 1108 4411 1118
rect 4419 1108 4449 1118
rect 4453 1108 4483 1122
rect 4511 1108 4524 1146
rect 4596 1152 4631 1160
rect 4596 1126 4597 1152
rect 4604 1126 4631 1152
rect 4539 1108 4569 1122
rect 4596 1118 4631 1126
rect 4596 1108 4597 1118
rect 4612 1108 4625 1118
rect -1 1102 4625 1108
rect 0 1094 4625 1102
rect 15 1064 28 1094
rect 43 1076 73 1094
rect 116 1080 130 1094
rect 166 1080 386 1094
rect 117 1078 130 1080
rect 83 1066 98 1078
rect 80 1064 102 1066
rect 107 1064 137 1078
rect 198 1076 351 1080
rect 180 1064 372 1076
rect 415 1064 445 1078
rect 451 1064 464 1094
rect 479 1076 509 1094
rect 552 1064 565 1094
rect 595 1064 608 1094
rect 623 1076 653 1094
rect 696 1080 710 1094
rect 746 1080 966 1094
rect 697 1078 710 1080
rect 663 1066 678 1078
rect 660 1064 682 1066
rect 687 1064 717 1078
rect 778 1076 931 1080
rect 760 1064 952 1076
rect 995 1064 1025 1078
rect 1031 1064 1044 1094
rect 1059 1076 1089 1094
rect 1132 1064 1145 1094
rect 1175 1064 1188 1094
rect 1203 1076 1233 1094
rect 1276 1080 1290 1094
rect 1326 1080 1546 1094
rect 1277 1078 1290 1080
rect 1243 1066 1258 1078
rect 1240 1064 1262 1066
rect 1267 1064 1297 1078
rect 1358 1076 1511 1080
rect 1340 1064 1532 1076
rect 1575 1064 1605 1078
rect 1611 1064 1624 1094
rect 1639 1076 1669 1094
rect 1712 1064 1725 1094
rect 1755 1064 1768 1094
rect 1783 1076 1813 1094
rect 1856 1080 1870 1094
rect 1906 1080 2126 1094
rect 1857 1078 1870 1080
rect 1823 1066 1838 1078
rect 1820 1064 1842 1066
rect 1847 1064 1877 1078
rect 1938 1076 2091 1080
rect 1920 1064 2112 1076
rect 2155 1064 2185 1078
rect 2191 1064 2204 1094
rect 2219 1076 2249 1094
rect 2292 1064 2305 1094
rect 2335 1064 2348 1094
rect 2363 1076 2393 1094
rect 2436 1080 2450 1094
rect 2486 1080 2706 1094
rect 2437 1078 2450 1080
rect 2403 1066 2418 1078
rect 2400 1064 2422 1066
rect 2427 1064 2457 1078
rect 2518 1076 2671 1080
rect 2500 1064 2692 1076
rect 2735 1064 2765 1078
rect 2771 1064 2784 1094
rect 2799 1076 2829 1094
rect 2872 1064 2885 1094
rect 2915 1064 2928 1094
rect 2943 1076 2973 1094
rect 3016 1080 3030 1094
rect 3066 1080 3286 1094
rect 3017 1078 3030 1080
rect 2983 1066 2998 1078
rect 2980 1064 3002 1066
rect 3007 1064 3037 1078
rect 3098 1076 3251 1080
rect 3080 1064 3272 1076
rect 3315 1064 3345 1078
rect 3351 1064 3364 1094
rect 3379 1076 3409 1094
rect 3452 1064 3465 1094
rect 3495 1064 3508 1094
rect 3523 1076 3553 1094
rect 3596 1080 3610 1094
rect 3646 1080 3866 1094
rect 3597 1078 3610 1080
rect 3563 1066 3578 1078
rect 3560 1064 3582 1066
rect 3587 1064 3617 1078
rect 3678 1076 3831 1080
rect 3660 1064 3852 1076
rect 3895 1064 3925 1078
rect 3931 1064 3944 1094
rect 3959 1076 3989 1094
rect 4032 1064 4045 1094
rect 4075 1064 4088 1094
rect 4103 1076 4133 1094
rect 4176 1080 4190 1094
rect 4226 1080 4446 1094
rect 4177 1078 4190 1080
rect 4143 1066 4158 1078
rect 4140 1064 4162 1066
rect 4167 1064 4197 1078
rect 4258 1076 4411 1080
rect 4240 1064 4432 1076
rect 4475 1064 4505 1078
rect 4511 1064 4524 1094
rect 4539 1076 4569 1094
rect 4612 1064 4625 1094
rect 0 1050 4625 1064
rect 15 946 28 1050
rect 73 1028 74 1038
rect 89 1028 102 1038
rect 73 1024 102 1028
rect 107 1024 137 1050
rect 155 1036 171 1038
rect 243 1036 296 1050
rect 244 1034 308 1036
rect 351 1034 366 1050
rect 415 1047 445 1050
rect 415 1044 451 1047
rect 381 1036 397 1038
rect 155 1024 170 1028
rect 73 1022 170 1024
rect 198 1022 366 1034
rect 382 1024 397 1028
rect 415 1025 454 1044
rect 473 1038 480 1039
rect 479 1031 480 1038
rect 463 1028 464 1031
rect 479 1028 492 1031
rect 415 1024 445 1025
rect 454 1024 460 1025
rect 463 1024 492 1028
rect 382 1023 492 1024
rect 382 1022 498 1023
rect 57 1014 108 1022
rect 57 1002 82 1014
rect 89 1002 108 1014
rect 139 1014 189 1022
rect 139 1006 155 1014
rect 162 1012 189 1014
rect 198 1012 419 1022
rect 162 1002 419 1012
rect 448 1014 498 1022
rect 448 1005 464 1014
rect 57 994 108 1002
rect 155 994 419 1002
rect 445 1002 464 1005
rect 471 1002 498 1014
rect 445 994 498 1002
rect 73 986 74 994
rect 89 986 102 994
rect 73 978 89 986
rect 70 971 89 974
rect 70 962 92 971
rect 43 952 92 962
rect 43 946 73 952
rect 92 947 97 952
rect 15 930 89 946
rect 107 938 137 994
rect 172 984 380 994
rect 415 990 460 994
rect 463 993 464 994
rect 479 993 492 994
rect 198 954 387 984
rect 213 951 387 954
rect 206 948 387 951
rect 15 928 28 930
rect 43 928 77 930
rect 15 912 89 928
rect 116 924 129 938
rect 144 924 160 940
rect 206 935 217 948
rect -1 890 0 906
rect 15 890 28 912
rect 43 890 73 912
rect 116 908 178 924
rect 206 917 217 933
rect 222 928 232 948
rect 242 928 256 948
rect 259 935 268 948
rect 284 935 293 948
rect 222 917 256 928
rect 259 917 268 933
rect 284 917 293 933
rect 300 928 310 948
rect 320 928 334 948
rect 335 935 346 948
rect 300 917 334 928
rect 335 917 346 933
rect 392 924 408 940
rect 415 938 445 990
rect 479 986 480 993
rect 464 978 480 986
rect 451 946 464 965
rect 479 946 509 962
rect 451 930 525 946
rect 451 928 464 930
rect 479 928 513 930
rect 116 906 129 908
rect 144 906 178 908
rect 116 890 178 906
rect 222 901 238 904
rect 300 901 330 912
rect 378 908 424 924
rect 451 912 525 928
rect 378 906 412 908
rect 377 890 424 906
rect 451 890 464 912
rect 479 890 509 912
rect 536 890 537 906
rect 552 890 565 1050
rect 595 946 608 1050
rect 653 1028 654 1038
rect 669 1028 682 1038
rect 653 1024 682 1028
rect 687 1024 717 1050
rect 735 1036 751 1038
rect 823 1036 876 1050
rect 824 1034 888 1036
rect 931 1034 946 1050
rect 995 1047 1025 1050
rect 995 1044 1031 1047
rect 961 1036 977 1038
rect 735 1024 750 1028
rect 653 1022 750 1024
rect 778 1022 946 1034
rect 962 1024 977 1028
rect 995 1025 1034 1044
rect 1053 1038 1060 1039
rect 1059 1031 1060 1038
rect 1043 1028 1044 1031
rect 1059 1028 1072 1031
rect 995 1024 1025 1025
rect 1034 1024 1040 1025
rect 1043 1024 1072 1028
rect 962 1023 1072 1024
rect 962 1022 1078 1023
rect 637 1014 688 1022
rect 637 1002 662 1014
rect 669 1002 688 1014
rect 719 1014 769 1022
rect 719 1006 735 1014
rect 742 1012 769 1014
rect 778 1012 999 1022
rect 742 1002 999 1012
rect 1028 1014 1078 1022
rect 1028 1005 1044 1014
rect 637 994 688 1002
rect 735 994 999 1002
rect 1025 1002 1044 1005
rect 1051 1002 1078 1014
rect 1025 994 1078 1002
rect 653 986 654 994
rect 669 986 682 994
rect 653 978 669 986
rect 650 971 669 974
rect 650 962 672 971
rect 623 952 672 962
rect 623 946 653 952
rect 672 947 677 952
rect 595 930 669 946
rect 687 938 717 994
rect 752 984 960 994
rect 995 990 1040 994
rect 1043 993 1044 994
rect 1059 993 1072 994
rect 778 954 967 984
rect 793 951 967 954
rect 786 948 967 951
rect 595 928 608 930
rect 623 928 657 930
rect 595 912 669 928
rect 696 924 709 938
rect 724 924 740 940
rect 786 935 797 948
rect 579 890 580 906
rect 595 890 608 912
rect 623 890 653 912
rect 696 908 758 924
rect 786 917 797 933
rect 802 928 812 948
rect 822 928 836 948
rect 839 935 848 948
rect 864 935 873 948
rect 802 917 836 928
rect 839 917 848 933
rect 864 917 873 933
rect 880 928 890 948
rect 900 928 914 948
rect 915 935 926 948
rect 880 917 914 928
rect 915 917 926 933
rect 972 924 988 940
rect 995 938 1025 990
rect 1059 986 1060 993
rect 1044 978 1060 986
rect 1031 946 1044 965
rect 1059 946 1089 962
rect 1031 930 1105 946
rect 1031 928 1044 930
rect 1059 928 1093 930
rect 696 906 709 908
rect 724 906 758 908
rect 696 890 758 906
rect 802 901 818 904
rect 880 901 910 912
rect 958 908 1004 924
rect 1031 912 1105 928
rect 958 906 992 908
rect 957 890 1004 906
rect 1031 890 1044 912
rect 1059 890 1089 912
rect 1116 890 1117 906
rect 1132 890 1145 1050
rect 1175 946 1188 1050
rect 1233 1028 1234 1038
rect 1249 1028 1262 1038
rect 1233 1024 1262 1028
rect 1267 1024 1297 1050
rect 1315 1036 1331 1038
rect 1403 1036 1456 1050
rect 1404 1034 1468 1036
rect 1511 1034 1526 1050
rect 1575 1047 1605 1050
rect 1575 1044 1611 1047
rect 1541 1036 1557 1038
rect 1315 1024 1330 1028
rect 1233 1022 1330 1024
rect 1358 1022 1526 1034
rect 1542 1024 1557 1028
rect 1575 1025 1614 1044
rect 1633 1038 1640 1039
rect 1639 1031 1640 1038
rect 1623 1028 1624 1031
rect 1639 1028 1652 1031
rect 1575 1024 1605 1025
rect 1614 1024 1620 1025
rect 1623 1024 1652 1028
rect 1542 1023 1652 1024
rect 1542 1022 1658 1023
rect 1217 1014 1268 1022
rect 1217 1002 1242 1014
rect 1249 1002 1268 1014
rect 1299 1014 1349 1022
rect 1299 1006 1315 1014
rect 1322 1012 1349 1014
rect 1358 1012 1579 1022
rect 1322 1002 1579 1012
rect 1608 1014 1658 1022
rect 1608 1005 1624 1014
rect 1217 994 1268 1002
rect 1315 994 1579 1002
rect 1605 1002 1624 1005
rect 1631 1002 1658 1014
rect 1605 994 1658 1002
rect 1233 986 1234 994
rect 1249 986 1262 994
rect 1233 978 1249 986
rect 1230 971 1249 974
rect 1230 962 1252 971
rect 1203 952 1252 962
rect 1203 946 1233 952
rect 1252 947 1257 952
rect 1175 930 1249 946
rect 1267 938 1297 994
rect 1332 984 1540 994
rect 1575 990 1620 994
rect 1623 993 1624 994
rect 1639 993 1652 994
rect 1358 954 1547 984
rect 1373 951 1547 954
rect 1366 948 1547 951
rect 1175 928 1188 930
rect 1203 928 1237 930
rect 1175 912 1249 928
rect 1276 924 1289 938
rect 1304 924 1320 940
rect 1366 935 1377 948
rect 1159 890 1160 906
rect 1175 890 1188 912
rect 1203 890 1233 912
rect 1276 908 1338 924
rect 1366 917 1377 933
rect 1382 928 1392 948
rect 1402 928 1416 948
rect 1419 935 1428 948
rect 1444 935 1453 948
rect 1382 917 1416 928
rect 1419 917 1428 933
rect 1444 917 1453 933
rect 1460 928 1470 948
rect 1480 928 1494 948
rect 1495 935 1506 948
rect 1460 917 1494 928
rect 1495 917 1506 933
rect 1552 924 1568 940
rect 1575 938 1605 990
rect 1639 986 1640 993
rect 1624 978 1640 986
rect 1611 946 1624 965
rect 1639 946 1669 962
rect 1611 930 1685 946
rect 1611 928 1624 930
rect 1639 928 1673 930
rect 1276 906 1289 908
rect 1304 906 1338 908
rect 1276 890 1338 906
rect 1382 901 1398 904
rect 1460 901 1490 912
rect 1538 908 1584 924
rect 1611 912 1685 928
rect 1538 906 1572 908
rect 1537 890 1584 906
rect 1611 890 1624 912
rect 1639 890 1669 912
rect 1696 890 1697 906
rect 1712 890 1725 1050
rect 1755 946 1768 1050
rect 1813 1028 1814 1038
rect 1829 1028 1842 1038
rect 1813 1024 1842 1028
rect 1847 1024 1877 1050
rect 1895 1036 1911 1038
rect 1983 1036 2036 1050
rect 1984 1034 2048 1036
rect 2091 1034 2106 1050
rect 2155 1047 2185 1050
rect 2155 1044 2191 1047
rect 2121 1036 2137 1038
rect 1895 1024 1910 1028
rect 1813 1022 1910 1024
rect 1938 1022 2106 1034
rect 2122 1024 2137 1028
rect 2155 1025 2194 1044
rect 2213 1038 2220 1039
rect 2219 1031 2220 1038
rect 2203 1028 2204 1031
rect 2219 1028 2232 1031
rect 2155 1024 2185 1025
rect 2194 1024 2200 1025
rect 2203 1024 2232 1028
rect 2122 1023 2232 1024
rect 2122 1022 2238 1023
rect 1797 1014 1848 1022
rect 1797 1002 1822 1014
rect 1829 1002 1848 1014
rect 1879 1014 1929 1022
rect 1879 1006 1895 1014
rect 1902 1012 1929 1014
rect 1938 1012 2159 1022
rect 1902 1002 2159 1012
rect 2188 1014 2238 1022
rect 2188 1005 2204 1014
rect 1797 994 1848 1002
rect 1895 994 2159 1002
rect 2185 1002 2204 1005
rect 2211 1002 2238 1014
rect 2185 994 2238 1002
rect 1813 986 1814 994
rect 1829 986 1842 994
rect 1813 978 1829 986
rect 1810 971 1829 974
rect 1810 962 1832 971
rect 1783 952 1832 962
rect 1783 946 1813 952
rect 1832 947 1837 952
rect 1755 930 1829 946
rect 1847 938 1877 994
rect 1912 984 2120 994
rect 2155 990 2200 994
rect 2203 993 2204 994
rect 2219 993 2232 994
rect 1938 954 2127 984
rect 1953 951 2127 954
rect 1946 948 2127 951
rect 1755 928 1768 930
rect 1783 928 1817 930
rect 1755 912 1829 928
rect 1856 924 1869 938
rect 1884 924 1900 940
rect 1946 935 1957 948
rect 1739 890 1740 906
rect 1755 890 1768 912
rect 1783 890 1813 912
rect 1856 908 1918 924
rect 1946 917 1957 933
rect 1962 928 1972 948
rect 1982 928 1996 948
rect 1999 935 2008 948
rect 2024 935 2033 948
rect 1962 917 1996 928
rect 1999 917 2008 933
rect 2024 917 2033 933
rect 2040 928 2050 948
rect 2060 928 2074 948
rect 2075 935 2086 948
rect 2040 917 2074 928
rect 2075 917 2086 933
rect 2132 924 2148 940
rect 2155 938 2185 990
rect 2219 986 2220 993
rect 2204 978 2220 986
rect 2191 946 2204 965
rect 2219 946 2249 962
rect 2191 930 2265 946
rect 2191 928 2204 930
rect 2219 928 2253 930
rect 1856 906 1869 908
rect 1884 906 1918 908
rect 1856 890 1918 906
rect 1962 901 1978 904
rect 2040 901 2070 912
rect 2118 908 2164 924
rect 2191 912 2265 928
rect 2118 906 2152 908
rect 2117 890 2164 906
rect 2191 890 2204 912
rect 2219 890 2249 912
rect 2276 890 2277 906
rect 2292 890 2305 1050
rect 2335 946 2348 1050
rect 2393 1028 2394 1038
rect 2409 1028 2422 1038
rect 2393 1024 2422 1028
rect 2427 1024 2457 1050
rect 2475 1036 2491 1038
rect 2563 1036 2616 1050
rect 2564 1034 2628 1036
rect 2671 1034 2686 1050
rect 2735 1047 2765 1050
rect 2735 1044 2771 1047
rect 2701 1036 2717 1038
rect 2475 1024 2490 1028
rect 2393 1022 2490 1024
rect 2518 1022 2686 1034
rect 2702 1024 2717 1028
rect 2735 1025 2774 1044
rect 2793 1038 2800 1039
rect 2799 1031 2800 1038
rect 2783 1028 2784 1031
rect 2799 1028 2812 1031
rect 2735 1024 2765 1025
rect 2774 1024 2780 1025
rect 2783 1024 2812 1028
rect 2702 1023 2812 1024
rect 2702 1022 2818 1023
rect 2377 1014 2428 1022
rect 2377 1002 2402 1014
rect 2409 1002 2428 1014
rect 2459 1014 2509 1022
rect 2459 1006 2475 1014
rect 2482 1012 2509 1014
rect 2518 1012 2739 1022
rect 2482 1002 2739 1012
rect 2768 1014 2818 1022
rect 2768 1005 2784 1014
rect 2377 994 2428 1002
rect 2475 994 2739 1002
rect 2765 1002 2784 1005
rect 2791 1002 2818 1014
rect 2765 994 2818 1002
rect 2393 986 2394 994
rect 2409 986 2422 994
rect 2393 978 2409 986
rect 2390 971 2409 974
rect 2390 962 2412 971
rect 2363 952 2412 962
rect 2363 946 2393 952
rect 2412 947 2417 952
rect 2335 930 2409 946
rect 2427 938 2457 994
rect 2492 984 2700 994
rect 2735 990 2780 994
rect 2783 993 2784 994
rect 2799 993 2812 994
rect 2518 954 2707 984
rect 2533 951 2707 954
rect 2526 948 2707 951
rect 2335 928 2348 930
rect 2363 928 2397 930
rect 2335 912 2409 928
rect 2436 924 2449 938
rect 2464 924 2480 940
rect 2526 935 2537 948
rect 2319 890 2320 906
rect 2335 890 2348 912
rect 2363 890 2393 912
rect 2436 908 2498 924
rect 2526 917 2537 933
rect 2542 928 2552 948
rect 2562 928 2576 948
rect 2579 935 2588 948
rect 2604 935 2613 948
rect 2542 917 2576 928
rect 2579 917 2588 933
rect 2604 917 2613 933
rect 2620 928 2630 948
rect 2640 928 2654 948
rect 2655 935 2666 948
rect 2620 917 2654 928
rect 2655 917 2666 933
rect 2712 924 2728 940
rect 2735 938 2765 990
rect 2799 986 2800 993
rect 2784 978 2800 986
rect 2771 946 2784 965
rect 2799 946 2829 962
rect 2771 930 2845 946
rect 2771 928 2784 930
rect 2799 928 2833 930
rect 2436 906 2449 908
rect 2464 906 2498 908
rect 2436 890 2498 906
rect 2542 901 2558 904
rect 2620 901 2650 912
rect 2698 908 2744 924
rect 2771 912 2845 928
rect 2698 906 2732 908
rect 2697 890 2744 906
rect 2771 890 2784 912
rect 2799 890 2829 912
rect 2856 890 2857 906
rect 2872 890 2885 1050
rect 2915 946 2928 1050
rect 2973 1028 2974 1038
rect 2989 1028 3002 1038
rect 2973 1024 3002 1028
rect 3007 1024 3037 1050
rect 3055 1036 3071 1038
rect 3143 1036 3196 1050
rect 3144 1034 3208 1036
rect 3251 1034 3266 1050
rect 3315 1047 3345 1050
rect 3315 1044 3351 1047
rect 3281 1036 3297 1038
rect 3055 1024 3070 1028
rect 2973 1022 3070 1024
rect 3098 1022 3266 1034
rect 3282 1024 3297 1028
rect 3315 1025 3354 1044
rect 3373 1038 3380 1039
rect 3379 1031 3380 1038
rect 3363 1028 3364 1031
rect 3379 1028 3392 1031
rect 3315 1024 3345 1025
rect 3354 1024 3360 1025
rect 3363 1024 3392 1028
rect 3282 1023 3392 1024
rect 3282 1022 3398 1023
rect 2957 1014 3008 1022
rect 2957 1002 2982 1014
rect 2989 1002 3008 1014
rect 3039 1014 3089 1022
rect 3039 1006 3055 1014
rect 3062 1012 3089 1014
rect 3098 1012 3319 1022
rect 3062 1002 3319 1012
rect 3348 1014 3398 1022
rect 3348 1005 3364 1014
rect 2957 994 3008 1002
rect 3055 994 3319 1002
rect 3345 1002 3364 1005
rect 3371 1002 3398 1014
rect 3345 994 3398 1002
rect 2973 986 2974 994
rect 2989 986 3002 994
rect 2973 978 2989 986
rect 2970 971 2989 974
rect 2970 962 2992 971
rect 2943 952 2992 962
rect 2943 946 2973 952
rect 2992 947 2997 952
rect 2915 930 2989 946
rect 3007 938 3037 994
rect 3072 984 3280 994
rect 3315 990 3360 994
rect 3363 993 3364 994
rect 3379 993 3392 994
rect 3098 954 3287 984
rect 3113 951 3287 954
rect 3106 948 3287 951
rect 2915 928 2928 930
rect 2943 928 2977 930
rect 2915 912 2989 928
rect 3016 924 3029 938
rect 3044 924 3060 940
rect 3106 935 3117 948
rect 2899 890 2900 906
rect 2915 890 2928 912
rect 2943 890 2973 912
rect 3016 908 3078 924
rect 3106 917 3117 933
rect 3122 928 3132 948
rect 3142 928 3156 948
rect 3159 935 3168 948
rect 3184 935 3193 948
rect 3122 917 3156 928
rect 3159 917 3168 933
rect 3184 917 3193 933
rect 3200 928 3210 948
rect 3220 928 3234 948
rect 3235 935 3246 948
rect 3200 917 3234 928
rect 3235 917 3246 933
rect 3292 924 3308 940
rect 3315 938 3345 990
rect 3379 986 3380 993
rect 3364 978 3380 986
rect 3351 946 3364 965
rect 3379 946 3409 962
rect 3351 930 3425 946
rect 3351 928 3364 930
rect 3379 928 3413 930
rect 3016 906 3029 908
rect 3044 906 3078 908
rect 3016 890 3078 906
rect 3122 901 3138 904
rect 3200 901 3230 912
rect 3278 908 3324 924
rect 3351 912 3425 928
rect 3278 906 3312 908
rect 3277 890 3324 906
rect 3351 890 3364 912
rect 3379 890 3409 912
rect 3436 890 3437 906
rect 3452 890 3465 1050
rect 3495 946 3508 1050
rect 3553 1028 3554 1038
rect 3569 1028 3582 1038
rect 3553 1024 3582 1028
rect 3587 1024 3617 1050
rect 3635 1036 3651 1038
rect 3723 1036 3776 1050
rect 3724 1034 3788 1036
rect 3831 1034 3846 1050
rect 3895 1047 3925 1050
rect 3895 1044 3931 1047
rect 3861 1036 3877 1038
rect 3635 1024 3650 1028
rect 3553 1022 3650 1024
rect 3678 1022 3846 1034
rect 3862 1024 3877 1028
rect 3895 1025 3934 1044
rect 3953 1038 3960 1039
rect 3959 1031 3960 1038
rect 3943 1028 3944 1031
rect 3959 1028 3972 1031
rect 3895 1024 3925 1025
rect 3934 1024 3940 1025
rect 3943 1024 3972 1028
rect 3862 1023 3972 1024
rect 3862 1022 3978 1023
rect 3537 1014 3588 1022
rect 3537 1002 3562 1014
rect 3569 1002 3588 1014
rect 3619 1014 3669 1022
rect 3619 1006 3635 1014
rect 3642 1012 3669 1014
rect 3678 1012 3899 1022
rect 3642 1002 3899 1012
rect 3928 1014 3978 1022
rect 3928 1005 3944 1014
rect 3537 994 3588 1002
rect 3635 994 3899 1002
rect 3925 1002 3944 1005
rect 3951 1002 3978 1014
rect 3925 994 3978 1002
rect 3553 986 3554 994
rect 3569 986 3582 994
rect 3553 978 3569 986
rect 3550 971 3569 974
rect 3550 962 3572 971
rect 3523 952 3572 962
rect 3523 946 3553 952
rect 3572 947 3577 952
rect 3495 930 3569 946
rect 3587 938 3617 994
rect 3652 984 3860 994
rect 3895 990 3940 994
rect 3943 993 3944 994
rect 3959 993 3972 994
rect 3678 954 3867 984
rect 3693 951 3867 954
rect 3686 948 3867 951
rect 3495 928 3508 930
rect 3523 928 3557 930
rect 3495 912 3569 928
rect 3596 924 3609 938
rect 3624 924 3640 940
rect 3686 935 3697 948
rect 3479 890 3480 906
rect 3495 890 3508 912
rect 3523 890 3553 912
rect 3596 908 3658 924
rect 3686 917 3697 933
rect 3702 928 3712 948
rect 3722 928 3736 948
rect 3739 935 3748 948
rect 3764 935 3773 948
rect 3702 917 3736 928
rect 3739 917 3748 933
rect 3764 917 3773 933
rect 3780 928 3790 948
rect 3800 928 3814 948
rect 3815 935 3826 948
rect 3780 917 3814 928
rect 3815 917 3826 933
rect 3872 924 3888 940
rect 3895 938 3925 990
rect 3959 986 3960 993
rect 3944 978 3960 986
rect 3931 946 3944 965
rect 3959 946 3989 962
rect 3931 930 4005 946
rect 3931 928 3944 930
rect 3959 928 3993 930
rect 3596 906 3609 908
rect 3624 906 3658 908
rect 3596 890 3658 906
rect 3702 901 3718 904
rect 3780 901 3810 912
rect 3858 908 3904 924
rect 3931 912 4005 928
rect 3858 906 3892 908
rect 3857 890 3904 906
rect 3931 890 3944 912
rect 3959 890 3989 912
rect 4016 890 4017 906
rect 4032 890 4045 1050
rect 4075 946 4088 1050
rect 4133 1028 4134 1038
rect 4149 1028 4162 1038
rect 4133 1024 4162 1028
rect 4167 1024 4197 1050
rect 4215 1036 4231 1038
rect 4303 1036 4356 1050
rect 4304 1034 4368 1036
rect 4411 1034 4426 1050
rect 4475 1047 4505 1050
rect 4475 1044 4511 1047
rect 4441 1036 4457 1038
rect 4215 1024 4230 1028
rect 4133 1022 4230 1024
rect 4258 1022 4426 1034
rect 4442 1024 4457 1028
rect 4475 1025 4514 1044
rect 4533 1038 4540 1039
rect 4539 1031 4540 1038
rect 4523 1028 4524 1031
rect 4539 1028 4552 1031
rect 4475 1024 4505 1025
rect 4514 1024 4520 1025
rect 4523 1024 4552 1028
rect 4442 1023 4552 1024
rect 4442 1022 4558 1023
rect 4117 1014 4168 1022
rect 4117 1002 4142 1014
rect 4149 1002 4168 1014
rect 4199 1014 4249 1022
rect 4199 1006 4215 1014
rect 4222 1012 4249 1014
rect 4258 1012 4479 1022
rect 4222 1002 4479 1012
rect 4508 1014 4558 1022
rect 4508 1005 4524 1014
rect 4117 994 4168 1002
rect 4215 994 4479 1002
rect 4505 1002 4524 1005
rect 4531 1002 4558 1014
rect 4505 994 4558 1002
rect 4133 986 4134 994
rect 4149 986 4162 994
rect 4133 978 4149 986
rect 4130 971 4149 974
rect 4130 962 4152 971
rect 4103 952 4152 962
rect 4103 946 4133 952
rect 4152 947 4157 952
rect 4075 930 4149 946
rect 4167 938 4197 994
rect 4232 984 4440 994
rect 4475 990 4520 994
rect 4523 993 4524 994
rect 4539 993 4552 994
rect 4258 954 4447 984
rect 4273 951 4447 954
rect 4266 948 4447 951
rect 4075 928 4088 930
rect 4103 928 4137 930
rect 4075 912 4149 928
rect 4176 924 4189 938
rect 4204 924 4220 940
rect 4266 935 4277 948
rect 4059 890 4060 906
rect 4075 890 4088 912
rect 4103 890 4133 912
rect 4176 908 4238 924
rect 4266 917 4277 933
rect 4282 928 4292 948
rect 4302 928 4316 948
rect 4319 935 4328 948
rect 4344 935 4353 948
rect 4282 917 4316 928
rect 4319 917 4328 933
rect 4344 917 4353 933
rect 4360 928 4370 948
rect 4380 928 4394 948
rect 4395 935 4406 948
rect 4360 917 4394 928
rect 4395 917 4406 933
rect 4452 924 4468 940
rect 4475 938 4505 990
rect 4539 986 4540 993
rect 4524 978 4540 986
rect 4511 946 4524 965
rect 4539 946 4569 962
rect 4511 930 4585 946
rect 4511 928 4524 930
rect 4539 928 4573 930
rect 4176 906 4189 908
rect 4204 906 4238 908
rect 4176 890 4238 906
rect 4282 901 4298 904
rect 4360 901 4390 912
rect 4438 908 4484 924
rect 4511 912 4585 928
rect 4438 906 4472 908
rect 4437 890 4484 906
rect 4511 890 4524 912
rect 4539 890 4569 912
rect 4596 890 4597 906
rect 4612 890 4625 1050
rect -7 882 34 890
rect -7 856 8 882
rect 15 856 34 882
rect 98 878 160 890
rect 172 878 247 890
rect 305 878 380 890
rect 392 878 423 890
rect 429 878 464 890
rect 98 876 260 878
rect -7 848 34 856
rect 116 852 129 876
rect 144 874 159 876
rect -1 838 0 848
rect 15 838 28 848
rect 43 838 73 852
rect 116 838 159 852
rect 183 849 190 856
rect 193 852 260 876
rect 292 876 464 878
rect 262 854 290 858
rect 292 854 372 876
rect 393 874 408 876
rect 262 852 372 854
rect 193 848 372 852
rect 166 838 196 848
rect 198 838 351 848
rect 359 838 389 848
rect 393 838 423 852
rect 451 838 464 876
rect 536 882 571 890
rect 536 856 537 882
rect 544 856 571 882
rect 479 838 509 852
rect 536 848 571 856
rect 573 882 614 890
rect 573 856 588 882
rect 595 856 614 882
rect 678 878 740 890
rect 752 878 827 890
rect 885 878 960 890
rect 972 878 1003 890
rect 1009 878 1044 890
rect 678 876 840 878
rect 573 848 614 856
rect 696 852 709 876
rect 724 874 739 876
rect 536 838 537 848
rect 552 838 565 848
rect 579 838 580 848
rect 595 838 608 848
rect 623 838 653 852
rect 696 838 739 852
rect 763 849 770 856
rect 773 852 840 876
rect 872 876 1044 878
rect 842 854 870 858
rect 872 854 952 876
rect 973 874 988 876
rect 842 852 952 854
rect 773 848 952 852
rect 746 838 776 848
rect 778 838 931 848
rect 939 838 969 848
rect 973 838 1003 852
rect 1031 838 1044 876
rect 1116 882 1151 890
rect 1116 856 1117 882
rect 1124 856 1151 882
rect 1059 838 1089 852
rect 1116 848 1151 856
rect 1153 882 1194 890
rect 1153 856 1168 882
rect 1175 856 1194 882
rect 1258 878 1320 890
rect 1332 878 1407 890
rect 1465 878 1540 890
rect 1552 878 1583 890
rect 1589 878 1624 890
rect 1258 876 1420 878
rect 1153 848 1194 856
rect 1276 852 1289 876
rect 1304 874 1319 876
rect 1116 838 1117 848
rect 1132 838 1145 848
rect 1159 838 1160 848
rect 1175 838 1188 848
rect 1203 838 1233 852
rect 1276 838 1319 852
rect 1343 849 1350 856
rect 1353 852 1420 876
rect 1452 876 1624 878
rect 1422 854 1450 858
rect 1452 854 1532 876
rect 1553 874 1568 876
rect 1422 852 1532 854
rect 1353 848 1532 852
rect 1326 838 1356 848
rect 1358 838 1511 848
rect 1519 838 1549 848
rect 1553 838 1583 852
rect 1611 838 1624 876
rect 1696 882 1731 890
rect 1696 856 1697 882
rect 1704 856 1731 882
rect 1639 838 1669 852
rect 1696 848 1731 856
rect 1733 882 1774 890
rect 1733 856 1748 882
rect 1755 856 1774 882
rect 1838 878 1900 890
rect 1912 878 1987 890
rect 2045 878 2120 890
rect 2132 878 2163 890
rect 2169 878 2204 890
rect 1838 876 2000 878
rect 1733 848 1774 856
rect 1856 852 1869 876
rect 1884 874 1899 876
rect 1696 838 1697 848
rect 1712 838 1725 848
rect 1739 838 1740 848
rect 1755 838 1768 848
rect 1783 838 1813 852
rect 1856 838 1899 852
rect 1923 849 1930 856
rect 1933 852 2000 876
rect 2032 876 2204 878
rect 2002 854 2030 858
rect 2032 854 2112 876
rect 2133 874 2148 876
rect 2002 852 2112 854
rect 1933 848 2112 852
rect 1906 838 1936 848
rect 1938 838 2091 848
rect 2099 838 2129 848
rect 2133 838 2163 852
rect 2191 838 2204 876
rect 2276 882 2311 890
rect 2276 856 2277 882
rect 2284 856 2311 882
rect 2219 838 2249 852
rect 2276 848 2311 856
rect 2313 882 2354 890
rect 2313 856 2328 882
rect 2335 856 2354 882
rect 2418 878 2480 890
rect 2492 878 2567 890
rect 2625 878 2700 890
rect 2712 878 2743 890
rect 2749 878 2784 890
rect 2418 876 2580 878
rect 2313 848 2354 856
rect 2436 852 2449 876
rect 2464 874 2479 876
rect 2276 838 2277 848
rect 2292 838 2305 848
rect 2319 838 2320 848
rect 2335 838 2348 848
rect 2363 838 2393 852
rect 2436 838 2479 852
rect 2503 849 2510 856
rect 2513 852 2580 876
rect 2612 876 2784 878
rect 2582 854 2610 858
rect 2612 854 2692 876
rect 2713 874 2728 876
rect 2582 852 2692 854
rect 2513 848 2692 852
rect 2486 838 2516 848
rect 2518 838 2671 848
rect 2679 838 2709 848
rect 2713 838 2743 852
rect 2771 838 2784 876
rect 2856 882 2891 890
rect 2856 856 2857 882
rect 2864 856 2891 882
rect 2799 838 2829 852
rect 2856 848 2891 856
rect 2893 882 2934 890
rect 2893 856 2908 882
rect 2915 856 2934 882
rect 2998 878 3060 890
rect 3072 878 3147 890
rect 3205 878 3280 890
rect 3292 878 3323 890
rect 3329 878 3364 890
rect 2998 876 3160 878
rect 2893 848 2934 856
rect 3016 852 3029 876
rect 3044 874 3059 876
rect 2856 838 2857 848
rect 2872 838 2885 848
rect 2899 838 2900 848
rect 2915 838 2928 848
rect 2943 838 2973 852
rect 3016 838 3059 852
rect 3083 849 3090 856
rect 3093 852 3160 876
rect 3192 876 3364 878
rect 3162 854 3190 858
rect 3192 854 3272 876
rect 3293 874 3308 876
rect 3162 852 3272 854
rect 3093 848 3272 852
rect 3066 838 3096 848
rect 3098 838 3251 848
rect 3259 838 3289 848
rect 3293 838 3323 852
rect 3351 838 3364 876
rect 3436 882 3471 890
rect 3436 856 3437 882
rect 3444 856 3471 882
rect 3379 838 3409 852
rect 3436 848 3471 856
rect 3473 882 3514 890
rect 3473 856 3488 882
rect 3495 856 3514 882
rect 3578 878 3640 890
rect 3652 878 3727 890
rect 3785 878 3860 890
rect 3872 878 3903 890
rect 3909 878 3944 890
rect 3578 876 3740 878
rect 3473 848 3514 856
rect 3596 852 3609 876
rect 3624 874 3639 876
rect 3436 838 3437 848
rect 3452 838 3465 848
rect 3479 838 3480 848
rect 3495 838 3508 848
rect 3523 838 3553 852
rect 3596 838 3639 852
rect 3663 849 3670 856
rect 3673 852 3740 876
rect 3772 876 3944 878
rect 3742 854 3770 858
rect 3772 854 3852 876
rect 3873 874 3888 876
rect 3742 852 3852 854
rect 3673 848 3852 852
rect 3646 838 3676 848
rect 3678 838 3831 848
rect 3839 838 3869 848
rect 3873 838 3903 852
rect 3931 838 3944 876
rect 4016 882 4051 890
rect 4016 856 4017 882
rect 4024 856 4051 882
rect 3959 838 3989 852
rect 4016 848 4051 856
rect 4053 882 4094 890
rect 4053 856 4068 882
rect 4075 856 4094 882
rect 4158 878 4220 890
rect 4232 878 4307 890
rect 4365 878 4440 890
rect 4452 878 4483 890
rect 4489 878 4524 890
rect 4158 876 4320 878
rect 4053 848 4094 856
rect 4176 852 4189 876
rect 4204 874 4219 876
rect 4016 838 4017 848
rect 4032 838 4045 848
rect 4059 838 4060 848
rect 4075 838 4088 848
rect 4103 838 4133 852
rect 4176 838 4219 852
rect 4243 849 4250 856
rect 4253 852 4320 876
rect 4352 876 4524 878
rect 4322 854 4350 858
rect 4352 854 4432 876
rect 4453 874 4468 876
rect 4322 852 4432 854
rect 4253 848 4432 852
rect 4226 838 4256 848
rect 4258 838 4411 848
rect 4419 838 4449 848
rect 4453 838 4483 852
rect 4511 838 4524 876
rect 4596 882 4631 890
rect 4596 856 4597 882
rect 4604 856 4631 882
rect 4539 838 4569 852
rect 4596 848 4631 856
rect 4596 838 4597 848
rect 4612 838 4625 848
rect -1 832 4625 838
rect 0 824 4625 832
rect 15 794 28 824
rect 43 806 73 824
rect 116 810 130 824
rect 166 810 386 824
rect 117 808 130 810
rect 83 796 98 808
rect 80 794 102 796
rect 107 794 137 808
rect 198 806 351 810
rect 180 794 372 806
rect 415 794 445 808
rect 451 794 464 824
rect 479 806 509 824
rect 552 794 565 824
rect 595 794 608 824
rect 623 806 653 824
rect 696 810 710 824
rect 746 810 966 824
rect 697 808 710 810
rect 663 796 678 808
rect 660 794 682 796
rect 687 794 717 808
rect 778 806 931 810
rect 760 794 952 806
rect 995 794 1025 808
rect 1031 794 1044 824
rect 1059 806 1089 824
rect 1132 794 1145 824
rect 1175 794 1188 824
rect 1203 806 1233 824
rect 1276 810 1290 824
rect 1326 810 1546 824
rect 1277 808 1290 810
rect 1243 796 1258 808
rect 1240 794 1262 796
rect 1267 794 1297 808
rect 1358 806 1511 810
rect 1340 794 1532 806
rect 1575 794 1605 808
rect 1611 794 1624 824
rect 1639 806 1669 824
rect 1712 794 1725 824
rect 1755 794 1768 824
rect 1783 806 1813 824
rect 1856 810 1870 824
rect 1906 810 2126 824
rect 1857 808 1870 810
rect 1823 796 1838 808
rect 1820 794 1842 796
rect 1847 794 1877 808
rect 1938 806 2091 810
rect 1920 794 2112 806
rect 2155 794 2185 808
rect 2191 794 2204 824
rect 2219 806 2249 824
rect 2292 794 2305 824
rect 2335 794 2348 824
rect 2363 806 2393 824
rect 2436 810 2450 824
rect 2486 810 2706 824
rect 2437 808 2450 810
rect 2403 796 2418 808
rect 2400 794 2422 796
rect 2427 794 2457 808
rect 2518 806 2671 810
rect 2500 794 2692 806
rect 2735 794 2765 808
rect 2771 794 2784 824
rect 2799 806 2829 824
rect 2872 794 2885 824
rect 2915 794 2928 824
rect 2943 806 2973 824
rect 3016 810 3030 824
rect 3066 810 3286 824
rect 3017 808 3030 810
rect 2983 796 2998 808
rect 2980 794 3002 796
rect 3007 794 3037 808
rect 3098 806 3251 810
rect 3080 794 3272 806
rect 3315 794 3345 808
rect 3351 794 3364 824
rect 3379 806 3409 824
rect 3452 794 3465 824
rect 3495 794 3508 824
rect 3523 806 3553 824
rect 3596 810 3610 824
rect 3646 810 3866 824
rect 3597 808 3610 810
rect 3563 796 3578 808
rect 3560 794 3582 796
rect 3587 794 3617 808
rect 3678 806 3831 810
rect 3660 794 3852 806
rect 3895 794 3925 808
rect 3931 794 3944 824
rect 3959 806 3989 824
rect 4032 794 4045 824
rect 4075 794 4088 824
rect 4103 806 4133 824
rect 4176 810 4190 824
rect 4226 810 4446 824
rect 4177 808 4190 810
rect 4143 796 4158 808
rect 4140 794 4162 796
rect 4167 794 4197 808
rect 4258 806 4411 810
rect 4240 794 4432 806
rect 4475 794 4505 808
rect 4511 794 4524 824
rect 4539 806 4569 824
rect 4612 794 4625 824
rect 0 780 4625 794
rect 15 676 28 780
rect 73 758 74 768
rect 89 758 102 768
rect 73 754 102 758
rect 107 754 137 780
rect 155 766 171 768
rect 243 766 296 780
rect 244 764 308 766
rect 351 764 366 780
rect 415 777 445 780
rect 415 774 451 777
rect 381 766 397 768
rect 155 754 170 758
rect 73 752 170 754
rect 198 752 366 764
rect 382 754 397 758
rect 415 755 454 774
rect 473 768 480 769
rect 479 761 480 768
rect 463 758 464 761
rect 479 758 492 761
rect 415 754 445 755
rect 454 754 460 755
rect 463 754 492 758
rect 382 753 492 754
rect 382 752 498 753
rect 57 744 108 752
rect 57 732 82 744
rect 89 732 108 744
rect 139 744 189 752
rect 139 736 155 744
rect 162 742 189 744
rect 198 742 419 752
rect 162 732 419 742
rect 448 744 498 752
rect 448 735 464 744
rect 57 724 108 732
rect 155 724 419 732
rect 445 732 464 735
rect 471 732 498 744
rect 445 724 498 732
rect 73 716 74 724
rect 89 716 102 724
rect 73 708 89 716
rect 70 701 89 704
rect 70 692 92 701
rect 43 682 92 692
rect 43 676 73 682
rect 92 677 97 682
rect 15 660 89 676
rect 107 668 137 724
rect 172 714 380 724
rect 415 720 460 724
rect 463 723 464 724
rect 479 723 492 724
rect 198 684 387 714
rect 213 681 387 684
rect 206 678 387 681
rect 15 658 28 660
rect 43 658 77 660
rect 15 642 89 658
rect 116 654 129 668
rect 144 654 160 670
rect 206 665 217 678
rect -1 620 0 636
rect 15 620 28 642
rect 43 620 73 642
rect 116 638 178 654
rect 206 647 217 663
rect 222 658 232 678
rect 242 658 256 678
rect 259 665 268 678
rect 284 665 293 678
rect 222 647 256 658
rect 259 647 268 663
rect 284 647 293 663
rect 300 658 310 678
rect 320 658 334 678
rect 335 665 346 678
rect 300 647 334 658
rect 335 647 346 663
rect 392 654 408 670
rect 415 668 445 720
rect 479 716 480 723
rect 464 708 480 716
rect 451 676 464 695
rect 479 676 509 692
rect 451 660 525 676
rect 451 658 464 660
rect 479 658 513 660
rect 116 636 129 638
rect 144 636 178 638
rect 116 620 178 636
rect 222 631 238 634
rect 300 631 330 642
rect 378 638 424 654
rect 451 642 525 658
rect 378 636 412 638
rect 377 620 424 636
rect 451 620 464 642
rect 479 620 509 642
rect 536 620 537 636
rect 552 620 565 780
rect 595 676 608 780
rect 653 758 654 768
rect 669 758 682 768
rect 653 754 682 758
rect 687 754 717 780
rect 735 766 751 768
rect 823 766 876 780
rect 824 764 888 766
rect 931 764 946 780
rect 995 777 1025 780
rect 995 774 1031 777
rect 961 766 977 768
rect 735 754 750 758
rect 653 752 750 754
rect 778 752 946 764
rect 962 754 977 758
rect 995 755 1034 774
rect 1053 768 1060 769
rect 1059 761 1060 768
rect 1043 758 1044 761
rect 1059 758 1072 761
rect 995 754 1025 755
rect 1034 754 1040 755
rect 1043 754 1072 758
rect 962 753 1072 754
rect 962 752 1078 753
rect 637 744 688 752
rect 637 732 662 744
rect 669 732 688 744
rect 719 744 769 752
rect 719 736 735 744
rect 742 742 769 744
rect 778 742 999 752
rect 742 732 999 742
rect 1028 744 1078 752
rect 1028 735 1044 744
rect 637 724 688 732
rect 735 724 999 732
rect 1025 732 1044 735
rect 1051 732 1078 744
rect 1025 724 1078 732
rect 653 716 654 724
rect 669 716 682 724
rect 653 708 669 716
rect 650 701 669 704
rect 650 692 672 701
rect 623 682 672 692
rect 623 676 653 682
rect 672 677 677 682
rect 595 660 669 676
rect 687 668 717 724
rect 752 714 960 724
rect 995 720 1040 724
rect 1043 723 1044 724
rect 1059 723 1072 724
rect 778 684 967 714
rect 793 681 967 684
rect 786 678 967 681
rect 595 658 608 660
rect 623 658 657 660
rect 595 642 669 658
rect 696 654 709 668
rect 724 654 740 670
rect 786 665 797 678
rect 579 620 580 636
rect 595 620 608 642
rect 623 620 653 642
rect 696 638 758 654
rect 786 647 797 663
rect 802 658 812 678
rect 822 658 836 678
rect 839 665 848 678
rect 864 665 873 678
rect 802 647 836 658
rect 839 647 848 663
rect 864 647 873 663
rect 880 658 890 678
rect 900 658 914 678
rect 915 665 926 678
rect 880 647 914 658
rect 915 647 926 663
rect 972 654 988 670
rect 995 668 1025 720
rect 1059 716 1060 723
rect 1044 708 1060 716
rect 1031 676 1044 695
rect 1059 676 1089 692
rect 1031 660 1105 676
rect 1031 658 1044 660
rect 1059 658 1093 660
rect 696 636 709 638
rect 724 636 758 638
rect 696 620 758 636
rect 802 631 818 634
rect 880 631 910 642
rect 958 638 1004 654
rect 1031 642 1105 658
rect 958 636 992 638
rect 957 620 1004 636
rect 1031 620 1044 642
rect 1059 620 1089 642
rect 1116 620 1117 636
rect 1132 620 1145 780
rect 1175 676 1188 780
rect 1233 758 1234 768
rect 1249 758 1262 768
rect 1233 754 1262 758
rect 1267 754 1297 780
rect 1315 766 1331 768
rect 1403 766 1456 780
rect 1404 764 1468 766
rect 1511 764 1526 780
rect 1575 777 1605 780
rect 1575 774 1611 777
rect 1541 766 1557 768
rect 1315 754 1330 758
rect 1233 752 1330 754
rect 1358 752 1526 764
rect 1542 754 1557 758
rect 1575 755 1614 774
rect 1633 768 1640 769
rect 1639 761 1640 768
rect 1623 758 1624 761
rect 1639 758 1652 761
rect 1575 754 1605 755
rect 1614 754 1620 755
rect 1623 754 1652 758
rect 1542 753 1652 754
rect 1542 752 1658 753
rect 1217 744 1268 752
rect 1217 732 1242 744
rect 1249 732 1268 744
rect 1299 744 1349 752
rect 1299 736 1315 744
rect 1322 742 1349 744
rect 1358 742 1579 752
rect 1322 732 1579 742
rect 1608 744 1658 752
rect 1608 735 1624 744
rect 1217 724 1268 732
rect 1315 724 1579 732
rect 1605 732 1624 735
rect 1631 732 1658 744
rect 1605 724 1658 732
rect 1233 716 1234 724
rect 1249 716 1262 724
rect 1233 708 1249 716
rect 1230 701 1249 704
rect 1230 692 1252 701
rect 1203 682 1252 692
rect 1203 676 1233 682
rect 1252 677 1257 682
rect 1175 660 1249 676
rect 1267 668 1297 724
rect 1332 714 1540 724
rect 1575 720 1620 724
rect 1623 723 1624 724
rect 1639 723 1652 724
rect 1358 684 1547 714
rect 1373 681 1547 684
rect 1366 678 1547 681
rect 1175 658 1188 660
rect 1203 658 1237 660
rect 1175 642 1249 658
rect 1276 654 1289 668
rect 1304 654 1320 670
rect 1366 665 1377 678
rect 1159 620 1160 636
rect 1175 620 1188 642
rect 1203 620 1233 642
rect 1276 638 1338 654
rect 1366 647 1377 663
rect 1382 658 1392 678
rect 1402 658 1416 678
rect 1419 665 1428 678
rect 1444 665 1453 678
rect 1382 647 1416 658
rect 1419 647 1428 663
rect 1444 647 1453 663
rect 1460 658 1470 678
rect 1480 658 1494 678
rect 1495 665 1506 678
rect 1460 647 1494 658
rect 1495 647 1506 663
rect 1552 654 1568 670
rect 1575 668 1605 720
rect 1639 716 1640 723
rect 1624 708 1640 716
rect 1611 676 1624 695
rect 1639 676 1669 692
rect 1611 660 1685 676
rect 1611 658 1624 660
rect 1639 658 1673 660
rect 1276 636 1289 638
rect 1304 636 1338 638
rect 1276 620 1338 636
rect 1382 631 1398 634
rect 1460 631 1490 642
rect 1538 638 1584 654
rect 1611 642 1685 658
rect 1538 636 1572 638
rect 1537 620 1584 636
rect 1611 620 1624 642
rect 1639 620 1669 642
rect 1696 620 1697 636
rect 1712 620 1725 780
rect 1755 676 1768 780
rect 1813 758 1814 768
rect 1829 758 1842 768
rect 1813 754 1842 758
rect 1847 754 1877 780
rect 1895 766 1911 768
rect 1983 766 2036 780
rect 1984 764 2048 766
rect 2091 764 2106 780
rect 2155 777 2185 780
rect 2155 774 2191 777
rect 2121 766 2137 768
rect 1895 754 1910 758
rect 1813 752 1910 754
rect 1938 752 2106 764
rect 2122 754 2137 758
rect 2155 755 2194 774
rect 2213 768 2220 769
rect 2219 761 2220 768
rect 2203 758 2204 761
rect 2219 758 2232 761
rect 2155 754 2185 755
rect 2194 754 2200 755
rect 2203 754 2232 758
rect 2122 753 2232 754
rect 2122 752 2238 753
rect 1797 744 1848 752
rect 1797 732 1822 744
rect 1829 732 1848 744
rect 1879 744 1929 752
rect 1879 736 1895 744
rect 1902 742 1929 744
rect 1938 742 2159 752
rect 1902 732 2159 742
rect 2188 744 2238 752
rect 2188 735 2204 744
rect 1797 724 1848 732
rect 1895 724 2159 732
rect 2185 732 2204 735
rect 2211 732 2238 744
rect 2185 724 2238 732
rect 1813 716 1814 724
rect 1829 716 1842 724
rect 1813 708 1829 716
rect 1810 701 1829 704
rect 1810 692 1832 701
rect 1783 682 1832 692
rect 1783 676 1813 682
rect 1832 677 1837 682
rect 1755 660 1829 676
rect 1847 668 1877 724
rect 1912 714 2120 724
rect 2155 720 2200 724
rect 2203 723 2204 724
rect 2219 723 2232 724
rect 1938 684 2127 714
rect 1953 681 2127 684
rect 1946 678 2127 681
rect 1755 658 1768 660
rect 1783 658 1817 660
rect 1755 642 1829 658
rect 1856 654 1869 668
rect 1884 654 1900 670
rect 1946 665 1957 678
rect 1739 620 1740 636
rect 1755 620 1768 642
rect 1783 620 1813 642
rect 1856 638 1918 654
rect 1946 647 1957 663
rect 1962 658 1972 678
rect 1982 658 1996 678
rect 1999 665 2008 678
rect 2024 665 2033 678
rect 1962 647 1996 658
rect 1999 647 2008 663
rect 2024 647 2033 663
rect 2040 658 2050 678
rect 2060 658 2074 678
rect 2075 665 2086 678
rect 2040 647 2074 658
rect 2075 647 2086 663
rect 2132 654 2148 670
rect 2155 668 2185 720
rect 2219 716 2220 723
rect 2204 708 2220 716
rect 2191 676 2204 695
rect 2219 676 2249 692
rect 2191 660 2265 676
rect 2191 658 2204 660
rect 2219 658 2253 660
rect 1856 636 1869 638
rect 1884 636 1918 638
rect 1856 620 1918 636
rect 1962 631 1978 634
rect 2040 631 2070 642
rect 2118 638 2164 654
rect 2191 642 2265 658
rect 2118 636 2152 638
rect 2117 620 2164 636
rect 2191 620 2204 642
rect 2219 620 2249 642
rect 2276 620 2277 636
rect 2292 620 2305 780
rect 2335 676 2348 780
rect 2393 758 2394 768
rect 2409 758 2422 768
rect 2393 754 2422 758
rect 2427 754 2457 780
rect 2475 766 2491 768
rect 2563 766 2616 780
rect 2564 764 2628 766
rect 2671 764 2686 780
rect 2735 777 2765 780
rect 2735 774 2771 777
rect 2701 766 2717 768
rect 2475 754 2490 758
rect 2393 752 2490 754
rect 2518 752 2686 764
rect 2702 754 2717 758
rect 2735 755 2774 774
rect 2793 768 2800 769
rect 2799 761 2800 768
rect 2783 758 2784 761
rect 2799 758 2812 761
rect 2735 754 2765 755
rect 2774 754 2780 755
rect 2783 754 2812 758
rect 2702 753 2812 754
rect 2702 752 2818 753
rect 2377 744 2428 752
rect 2377 732 2402 744
rect 2409 732 2428 744
rect 2459 744 2509 752
rect 2459 736 2475 744
rect 2482 742 2509 744
rect 2518 742 2739 752
rect 2482 732 2739 742
rect 2768 744 2818 752
rect 2768 735 2784 744
rect 2377 724 2428 732
rect 2475 724 2739 732
rect 2765 732 2784 735
rect 2791 732 2818 744
rect 2765 724 2818 732
rect 2393 716 2394 724
rect 2409 716 2422 724
rect 2393 708 2409 716
rect 2390 701 2409 704
rect 2390 692 2412 701
rect 2363 682 2412 692
rect 2363 676 2393 682
rect 2412 677 2417 682
rect 2335 660 2409 676
rect 2427 668 2457 724
rect 2492 714 2700 724
rect 2735 720 2780 724
rect 2783 723 2784 724
rect 2799 723 2812 724
rect 2518 684 2707 714
rect 2533 681 2707 684
rect 2526 678 2707 681
rect 2335 658 2348 660
rect 2363 658 2397 660
rect 2335 642 2409 658
rect 2436 654 2449 668
rect 2464 654 2480 670
rect 2526 665 2537 678
rect 2319 620 2320 636
rect 2335 620 2348 642
rect 2363 620 2393 642
rect 2436 638 2498 654
rect 2526 647 2537 663
rect 2542 658 2552 678
rect 2562 658 2576 678
rect 2579 665 2588 678
rect 2604 665 2613 678
rect 2542 647 2576 658
rect 2579 647 2588 663
rect 2604 647 2613 663
rect 2620 658 2630 678
rect 2640 658 2654 678
rect 2655 665 2666 678
rect 2620 647 2654 658
rect 2655 647 2666 663
rect 2712 654 2728 670
rect 2735 668 2765 720
rect 2799 716 2800 723
rect 2784 708 2800 716
rect 2771 676 2784 695
rect 2799 676 2829 692
rect 2771 660 2845 676
rect 2771 658 2784 660
rect 2799 658 2833 660
rect 2436 636 2449 638
rect 2464 636 2498 638
rect 2436 620 2498 636
rect 2542 631 2558 634
rect 2620 631 2650 642
rect 2698 638 2744 654
rect 2771 642 2845 658
rect 2698 636 2732 638
rect 2697 620 2744 636
rect 2771 620 2784 642
rect 2799 620 2829 642
rect 2856 620 2857 636
rect 2872 620 2885 780
rect 2915 676 2928 780
rect 2973 758 2974 768
rect 2989 758 3002 768
rect 2973 754 3002 758
rect 3007 754 3037 780
rect 3055 766 3071 768
rect 3143 766 3196 780
rect 3144 764 3208 766
rect 3251 764 3266 780
rect 3315 777 3345 780
rect 3315 774 3351 777
rect 3281 766 3297 768
rect 3055 754 3070 758
rect 2973 752 3070 754
rect 3098 752 3266 764
rect 3282 754 3297 758
rect 3315 755 3354 774
rect 3373 768 3380 769
rect 3379 761 3380 768
rect 3363 758 3364 761
rect 3379 758 3392 761
rect 3315 754 3345 755
rect 3354 754 3360 755
rect 3363 754 3392 758
rect 3282 753 3392 754
rect 3282 752 3398 753
rect 2957 744 3008 752
rect 2957 732 2982 744
rect 2989 732 3008 744
rect 3039 744 3089 752
rect 3039 736 3055 744
rect 3062 742 3089 744
rect 3098 742 3319 752
rect 3062 732 3319 742
rect 3348 744 3398 752
rect 3348 735 3364 744
rect 2957 724 3008 732
rect 3055 724 3319 732
rect 3345 732 3364 735
rect 3371 732 3398 744
rect 3345 724 3398 732
rect 2973 716 2974 724
rect 2989 716 3002 724
rect 2973 708 2989 716
rect 2970 701 2989 704
rect 2970 692 2992 701
rect 2943 682 2992 692
rect 2943 676 2973 682
rect 2992 677 2997 682
rect 2915 660 2989 676
rect 3007 668 3037 724
rect 3072 714 3280 724
rect 3315 720 3360 724
rect 3363 723 3364 724
rect 3379 723 3392 724
rect 3098 684 3287 714
rect 3113 681 3287 684
rect 3106 678 3287 681
rect 2915 658 2928 660
rect 2943 658 2977 660
rect 2915 642 2989 658
rect 3016 654 3029 668
rect 3044 654 3060 670
rect 3106 665 3117 678
rect 2899 620 2900 636
rect 2915 620 2928 642
rect 2943 620 2973 642
rect 3016 638 3078 654
rect 3106 647 3117 663
rect 3122 658 3132 678
rect 3142 658 3156 678
rect 3159 665 3168 678
rect 3184 665 3193 678
rect 3122 647 3156 658
rect 3159 647 3168 663
rect 3184 647 3193 663
rect 3200 658 3210 678
rect 3220 658 3234 678
rect 3235 665 3246 678
rect 3200 647 3234 658
rect 3235 647 3246 663
rect 3292 654 3308 670
rect 3315 668 3345 720
rect 3379 716 3380 723
rect 3364 708 3380 716
rect 3351 676 3364 695
rect 3379 676 3409 692
rect 3351 660 3425 676
rect 3351 658 3364 660
rect 3379 658 3413 660
rect 3016 636 3029 638
rect 3044 636 3078 638
rect 3016 620 3078 636
rect 3122 631 3138 634
rect 3200 631 3230 642
rect 3278 638 3324 654
rect 3351 642 3425 658
rect 3278 636 3312 638
rect 3277 620 3324 636
rect 3351 620 3364 642
rect 3379 620 3409 642
rect 3436 620 3437 636
rect 3452 620 3465 780
rect 3495 676 3508 780
rect 3553 758 3554 768
rect 3569 758 3582 768
rect 3553 754 3582 758
rect 3587 754 3617 780
rect 3635 766 3651 768
rect 3723 766 3776 780
rect 3724 764 3788 766
rect 3831 764 3846 780
rect 3895 777 3925 780
rect 3895 774 3931 777
rect 3861 766 3877 768
rect 3635 754 3650 758
rect 3553 752 3650 754
rect 3678 752 3846 764
rect 3862 754 3877 758
rect 3895 755 3934 774
rect 3953 768 3960 769
rect 3959 761 3960 768
rect 3943 758 3944 761
rect 3959 758 3972 761
rect 3895 754 3925 755
rect 3934 754 3940 755
rect 3943 754 3972 758
rect 3862 753 3972 754
rect 3862 752 3978 753
rect 3537 744 3588 752
rect 3537 732 3562 744
rect 3569 732 3588 744
rect 3619 744 3669 752
rect 3619 736 3635 744
rect 3642 742 3669 744
rect 3678 742 3899 752
rect 3642 732 3899 742
rect 3928 744 3978 752
rect 3928 735 3944 744
rect 3537 724 3588 732
rect 3635 724 3899 732
rect 3925 732 3944 735
rect 3951 732 3978 744
rect 3925 724 3978 732
rect 3553 716 3554 724
rect 3569 716 3582 724
rect 3553 708 3569 716
rect 3550 701 3569 704
rect 3550 692 3572 701
rect 3523 682 3572 692
rect 3523 676 3553 682
rect 3572 677 3577 682
rect 3495 660 3569 676
rect 3587 668 3617 724
rect 3652 714 3860 724
rect 3895 720 3940 724
rect 3943 723 3944 724
rect 3959 723 3972 724
rect 3678 684 3867 714
rect 3693 681 3867 684
rect 3686 678 3867 681
rect 3495 658 3508 660
rect 3523 658 3557 660
rect 3495 642 3569 658
rect 3596 654 3609 668
rect 3624 654 3640 670
rect 3686 665 3697 678
rect 3479 620 3480 636
rect 3495 620 3508 642
rect 3523 620 3553 642
rect 3596 638 3658 654
rect 3686 647 3697 663
rect 3702 658 3712 678
rect 3722 658 3736 678
rect 3739 665 3748 678
rect 3764 665 3773 678
rect 3702 647 3736 658
rect 3739 647 3748 663
rect 3764 647 3773 663
rect 3780 658 3790 678
rect 3800 658 3814 678
rect 3815 665 3826 678
rect 3780 647 3814 658
rect 3815 647 3826 663
rect 3872 654 3888 670
rect 3895 668 3925 720
rect 3959 716 3960 723
rect 3944 708 3960 716
rect 3931 676 3944 695
rect 3959 676 3989 692
rect 3931 660 4005 676
rect 3931 658 3944 660
rect 3959 658 3993 660
rect 3596 636 3609 638
rect 3624 636 3658 638
rect 3596 620 3658 636
rect 3702 631 3718 634
rect 3780 631 3810 642
rect 3858 638 3904 654
rect 3931 642 4005 658
rect 3858 636 3892 638
rect 3857 620 3904 636
rect 3931 620 3944 642
rect 3959 620 3989 642
rect 4016 620 4017 636
rect 4032 620 4045 780
rect 4075 676 4088 780
rect 4133 758 4134 768
rect 4149 758 4162 768
rect 4133 754 4162 758
rect 4167 754 4197 780
rect 4215 766 4231 768
rect 4303 766 4356 780
rect 4304 764 4368 766
rect 4411 764 4426 780
rect 4475 777 4505 780
rect 4475 774 4511 777
rect 4441 766 4457 768
rect 4215 754 4230 758
rect 4133 752 4230 754
rect 4258 752 4426 764
rect 4442 754 4457 758
rect 4475 755 4514 774
rect 4533 768 4540 769
rect 4539 761 4540 768
rect 4523 758 4524 761
rect 4539 758 4552 761
rect 4475 754 4505 755
rect 4514 754 4520 755
rect 4523 754 4552 758
rect 4442 753 4552 754
rect 4442 752 4558 753
rect 4117 744 4168 752
rect 4117 732 4142 744
rect 4149 732 4168 744
rect 4199 744 4249 752
rect 4199 736 4215 744
rect 4222 742 4249 744
rect 4258 742 4479 752
rect 4222 732 4479 742
rect 4508 744 4558 752
rect 4508 735 4524 744
rect 4117 724 4168 732
rect 4215 724 4479 732
rect 4505 732 4524 735
rect 4531 732 4558 744
rect 4505 724 4558 732
rect 4133 716 4134 724
rect 4149 716 4162 724
rect 4133 708 4149 716
rect 4130 701 4149 704
rect 4130 692 4152 701
rect 4103 682 4152 692
rect 4103 676 4133 682
rect 4152 677 4157 682
rect 4075 660 4149 676
rect 4167 668 4197 724
rect 4232 714 4440 724
rect 4475 720 4520 724
rect 4523 723 4524 724
rect 4539 723 4552 724
rect 4258 684 4447 714
rect 4273 681 4447 684
rect 4266 678 4447 681
rect 4075 658 4088 660
rect 4103 658 4137 660
rect 4075 642 4149 658
rect 4176 654 4189 668
rect 4204 654 4220 670
rect 4266 665 4277 678
rect 4059 620 4060 636
rect 4075 620 4088 642
rect 4103 620 4133 642
rect 4176 638 4238 654
rect 4266 647 4277 663
rect 4282 658 4292 678
rect 4302 658 4316 678
rect 4319 665 4328 678
rect 4344 665 4353 678
rect 4282 647 4316 658
rect 4319 647 4328 663
rect 4344 647 4353 663
rect 4360 658 4370 678
rect 4380 658 4394 678
rect 4395 665 4406 678
rect 4360 647 4394 658
rect 4395 647 4406 663
rect 4452 654 4468 670
rect 4475 668 4505 720
rect 4539 716 4540 723
rect 4524 708 4540 716
rect 4511 676 4524 695
rect 4539 676 4569 692
rect 4511 660 4585 676
rect 4511 658 4524 660
rect 4539 658 4573 660
rect 4176 636 4189 638
rect 4204 636 4238 638
rect 4176 620 4238 636
rect 4282 631 4298 634
rect 4360 631 4390 642
rect 4438 638 4484 654
rect 4511 642 4585 658
rect 4438 636 4472 638
rect 4437 620 4484 636
rect 4511 620 4524 642
rect 4539 620 4569 642
rect 4596 620 4597 636
rect 4612 620 4625 780
rect -7 612 34 620
rect -7 586 8 612
rect 15 586 34 612
rect 98 608 160 620
rect 172 608 247 620
rect 305 608 380 620
rect 392 608 423 620
rect 429 608 464 620
rect 98 606 260 608
rect -7 578 34 586
rect 116 582 129 606
rect 144 604 159 606
rect -1 568 0 578
rect 15 568 28 578
rect 43 568 73 582
rect 116 568 159 582
rect 183 579 190 586
rect 193 582 260 606
rect 292 606 464 608
rect 262 584 290 588
rect 292 584 372 606
rect 393 604 408 606
rect 262 582 372 584
rect 193 578 372 582
rect 166 568 196 578
rect 198 568 351 578
rect 359 568 389 578
rect 393 568 423 582
rect 451 568 464 606
rect 536 612 571 620
rect 536 586 537 612
rect 544 586 571 612
rect 479 568 509 582
rect 536 578 571 586
rect 573 612 614 620
rect 573 586 588 612
rect 595 586 614 612
rect 678 608 740 620
rect 752 608 827 620
rect 885 608 960 620
rect 972 608 1003 620
rect 1009 608 1044 620
rect 678 606 840 608
rect 573 578 614 586
rect 696 582 709 606
rect 724 604 739 606
rect 536 568 537 578
rect 552 568 565 578
rect 579 568 580 578
rect 595 568 608 578
rect 623 568 653 582
rect 696 568 739 582
rect 763 579 770 586
rect 773 582 840 606
rect 872 606 1044 608
rect 842 584 870 588
rect 872 584 952 606
rect 973 604 988 606
rect 842 582 952 584
rect 773 578 952 582
rect 746 568 776 578
rect 778 568 931 578
rect 939 568 969 578
rect 973 568 1003 582
rect 1031 568 1044 606
rect 1116 612 1151 620
rect 1116 586 1117 612
rect 1124 586 1151 612
rect 1059 568 1089 582
rect 1116 578 1151 586
rect 1153 612 1194 620
rect 1153 586 1168 612
rect 1175 586 1194 612
rect 1258 608 1320 620
rect 1332 608 1407 620
rect 1465 608 1540 620
rect 1552 608 1583 620
rect 1589 608 1624 620
rect 1258 606 1420 608
rect 1153 578 1194 586
rect 1276 582 1289 606
rect 1304 604 1319 606
rect 1116 568 1117 578
rect 1132 568 1145 578
rect 1159 568 1160 578
rect 1175 568 1188 578
rect 1203 568 1233 582
rect 1276 568 1319 582
rect 1343 579 1350 586
rect 1353 582 1420 606
rect 1452 606 1624 608
rect 1422 584 1450 588
rect 1452 584 1532 606
rect 1553 604 1568 606
rect 1422 582 1532 584
rect 1353 578 1532 582
rect 1326 568 1356 578
rect 1358 568 1511 578
rect 1519 568 1549 578
rect 1553 568 1583 582
rect 1611 568 1624 606
rect 1696 612 1731 620
rect 1696 586 1697 612
rect 1704 586 1731 612
rect 1639 568 1669 582
rect 1696 578 1731 586
rect 1733 612 1774 620
rect 1733 586 1748 612
rect 1755 586 1774 612
rect 1838 608 1900 620
rect 1912 608 1987 620
rect 2045 608 2120 620
rect 2132 608 2163 620
rect 2169 608 2204 620
rect 1838 606 2000 608
rect 1733 578 1774 586
rect 1856 582 1869 606
rect 1884 604 1899 606
rect 1696 568 1697 578
rect 1712 568 1725 578
rect 1739 568 1740 578
rect 1755 568 1768 578
rect 1783 568 1813 582
rect 1856 568 1899 582
rect 1923 579 1930 586
rect 1933 582 2000 606
rect 2032 606 2204 608
rect 2002 584 2030 588
rect 2032 584 2112 606
rect 2133 604 2148 606
rect 2002 582 2112 584
rect 1933 578 2112 582
rect 1906 568 1936 578
rect 1938 568 2091 578
rect 2099 568 2129 578
rect 2133 568 2163 582
rect 2191 568 2204 606
rect 2276 612 2311 620
rect 2276 586 2277 612
rect 2284 586 2311 612
rect 2219 568 2249 582
rect 2276 578 2311 586
rect 2313 612 2354 620
rect 2313 586 2328 612
rect 2335 586 2354 612
rect 2418 608 2480 620
rect 2492 608 2567 620
rect 2625 608 2700 620
rect 2712 608 2743 620
rect 2749 608 2784 620
rect 2418 606 2580 608
rect 2313 578 2354 586
rect 2436 582 2449 606
rect 2464 604 2479 606
rect 2276 568 2277 578
rect 2292 568 2305 578
rect 2319 568 2320 578
rect 2335 568 2348 578
rect 2363 568 2393 582
rect 2436 568 2479 582
rect 2503 579 2510 586
rect 2513 582 2580 606
rect 2612 606 2784 608
rect 2582 584 2610 588
rect 2612 584 2692 606
rect 2713 604 2728 606
rect 2582 582 2692 584
rect 2513 578 2692 582
rect 2486 568 2516 578
rect 2518 568 2671 578
rect 2679 568 2709 578
rect 2713 568 2743 582
rect 2771 568 2784 606
rect 2856 612 2891 620
rect 2856 586 2857 612
rect 2864 586 2891 612
rect 2799 568 2829 582
rect 2856 578 2891 586
rect 2893 612 2934 620
rect 2893 586 2908 612
rect 2915 586 2934 612
rect 2998 608 3060 620
rect 3072 608 3147 620
rect 3205 608 3280 620
rect 3292 608 3323 620
rect 3329 608 3364 620
rect 2998 606 3160 608
rect 2893 578 2934 586
rect 3016 582 3029 606
rect 3044 604 3059 606
rect 2856 568 2857 578
rect 2872 568 2885 578
rect 2899 568 2900 578
rect 2915 568 2928 578
rect 2943 568 2973 582
rect 3016 568 3059 582
rect 3083 579 3090 586
rect 3093 582 3160 606
rect 3192 606 3364 608
rect 3162 584 3190 588
rect 3192 584 3272 606
rect 3293 604 3308 606
rect 3162 582 3272 584
rect 3093 578 3272 582
rect 3066 568 3096 578
rect 3098 568 3251 578
rect 3259 568 3289 578
rect 3293 568 3323 582
rect 3351 568 3364 606
rect 3436 612 3471 620
rect 3436 586 3437 612
rect 3444 586 3471 612
rect 3379 568 3409 582
rect 3436 578 3471 586
rect 3473 612 3514 620
rect 3473 586 3488 612
rect 3495 586 3514 612
rect 3578 608 3640 620
rect 3652 608 3727 620
rect 3785 608 3860 620
rect 3872 608 3903 620
rect 3909 608 3944 620
rect 3578 606 3740 608
rect 3473 578 3514 586
rect 3596 582 3609 606
rect 3624 604 3639 606
rect 3436 568 3437 578
rect 3452 568 3465 578
rect 3479 568 3480 578
rect 3495 568 3508 578
rect 3523 568 3553 582
rect 3596 568 3639 582
rect 3663 579 3670 586
rect 3673 582 3740 606
rect 3772 606 3944 608
rect 3742 584 3770 588
rect 3772 584 3852 606
rect 3873 604 3888 606
rect 3742 582 3852 584
rect 3673 578 3852 582
rect 3646 568 3676 578
rect 3678 568 3831 578
rect 3839 568 3869 578
rect 3873 568 3903 582
rect 3931 568 3944 606
rect 4016 612 4051 620
rect 4016 586 4017 612
rect 4024 586 4051 612
rect 3959 568 3989 582
rect 4016 578 4051 586
rect 4053 612 4094 620
rect 4053 586 4068 612
rect 4075 586 4094 612
rect 4158 608 4220 620
rect 4232 608 4307 620
rect 4365 608 4440 620
rect 4452 608 4483 620
rect 4489 608 4524 620
rect 4158 606 4320 608
rect 4053 578 4094 586
rect 4176 582 4189 606
rect 4204 604 4219 606
rect 4016 568 4017 578
rect 4032 568 4045 578
rect 4059 568 4060 578
rect 4075 568 4088 578
rect 4103 568 4133 582
rect 4176 568 4219 582
rect 4243 579 4250 586
rect 4253 582 4320 606
rect 4352 606 4524 608
rect 4322 584 4350 588
rect 4352 584 4432 606
rect 4453 604 4468 606
rect 4322 582 4432 584
rect 4253 578 4432 582
rect 4226 568 4256 578
rect 4258 568 4411 578
rect 4419 568 4449 578
rect 4453 568 4483 582
rect 4511 568 4524 606
rect 4596 612 4631 620
rect 4596 586 4597 612
rect 4604 586 4631 612
rect 4539 568 4569 582
rect 4596 578 4631 586
rect 4596 568 4597 578
rect 4612 568 4625 578
rect -1 562 4625 568
rect 0 554 4625 562
rect 15 524 28 554
rect 43 536 73 554
rect 116 540 130 554
rect 166 540 386 554
rect 117 538 130 540
rect 83 526 98 538
rect 80 524 102 526
rect 107 524 137 538
rect 198 536 351 540
rect 180 524 372 536
rect 415 524 445 538
rect 451 524 464 554
rect 479 536 509 554
rect 552 524 565 554
rect 595 524 608 554
rect 623 536 653 554
rect 696 540 710 554
rect 746 540 966 554
rect 697 538 710 540
rect 663 526 678 538
rect 660 524 682 526
rect 687 524 717 538
rect 778 536 931 540
rect 760 524 952 536
rect 995 524 1025 538
rect 1031 524 1044 554
rect 1059 536 1089 554
rect 1132 524 1145 554
rect 1175 524 1188 554
rect 1203 536 1233 554
rect 1276 540 1290 554
rect 1326 540 1546 554
rect 1277 538 1290 540
rect 1243 526 1258 538
rect 1240 524 1262 526
rect 1267 524 1297 538
rect 1358 536 1511 540
rect 1340 524 1532 536
rect 1575 524 1605 538
rect 1611 524 1624 554
rect 1639 536 1669 554
rect 1712 524 1725 554
rect 1755 524 1768 554
rect 1783 536 1813 554
rect 1856 540 1870 554
rect 1906 540 2126 554
rect 1857 538 1870 540
rect 1823 526 1838 538
rect 1820 524 1842 526
rect 1847 524 1877 538
rect 1938 536 2091 540
rect 1920 524 2112 536
rect 2155 524 2185 538
rect 2191 524 2204 554
rect 2219 536 2249 554
rect 2292 524 2305 554
rect 2335 524 2348 554
rect 2363 536 2393 554
rect 2436 540 2450 554
rect 2486 540 2706 554
rect 2437 538 2450 540
rect 2403 526 2418 538
rect 2400 524 2422 526
rect 2427 524 2457 538
rect 2518 536 2671 540
rect 2500 524 2692 536
rect 2735 524 2765 538
rect 2771 524 2784 554
rect 2799 536 2829 554
rect 2872 524 2885 554
rect 2915 524 2928 554
rect 2943 536 2973 554
rect 3016 540 3030 554
rect 3066 540 3286 554
rect 3017 538 3030 540
rect 2983 526 2998 538
rect 2980 524 3002 526
rect 3007 524 3037 538
rect 3098 536 3251 540
rect 3080 524 3272 536
rect 3315 524 3345 538
rect 3351 524 3364 554
rect 3379 536 3409 554
rect 3452 524 3465 554
rect 3495 524 3508 554
rect 3523 536 3553 554
rect 3596 540 3610 554
rect 3646 540 3866 554
rect 3597 538 3610 540
rect 3563 526 3578 538
rect 3560 524 3582 526
rect 3587 524 3617 538
rect 3678 536 3831 540
rect 3660 524 3852 536
rect 3895 524 3925 538
rect 3931 524 3944 554
rect 3959 536 3989 554
rect 4032 524 4045 554
rect 4075 524 4088 554
rect 4103 536 4133 554
rect 4176 540 4190 554
rect 4226 540 4446 554
rect 4177 538 4190 540
rect 4143 526 4158 538
rect 4140 524 4162 526
rect 4167 524 4197 538
rect 4258 536 4411 540
rect 4240 524 4432 536
rect 4475 524 4505 538
rect 4511 524 4524 554
rect 4539 536 4569 554
rect 4612 524 4625 554
rect 0 510 4625 524
rect 15 406 28 510
rect 73 488 74 498
rect 89 488 102 498
rect 73 484 102 488
rect 107 484 137 510
rect 155 496 171 498
rect 243 496 296 510
rect 244 494 308 496
rect 351 494 366 510
rect 415 507 445 510
rect 415 504 451 507
rect 381 496 397 498
rect 155 484 170 488
rect 73 482 170 484
rect 198 482 366 494
rect 382 484 397 488
rect 415 485 454 504
rect 473 498 480 499
rect 479 491 480 498
rect 463 488 464 491
rect 479 488 492 491
rect 415 484 445 485
rect 454 484 460 485
rect 463 484 492 488
rect 382 483 492 484
rect 382 482 498 483
rect 57 474 108 482
rect 57 462 82 474
rect 89 462 108 474
rect 139 474 189 482
rect 139 466 155 474
rect 162 472 189 474
rect 198 472 419 482
rect 162 462 419 472
rect 448 474 498 482
rect 448 465 464 474
rect 57 454 108 462
rect 155 454 419 462
rect 445 462 464 465
rect 471 462 498 474
rect 445 454 498 462
rect 73 446 74 454
rect 89 446 102 454
rect 73 438 89 446
rect 70 431 89 434
rect 70 422 92 431
rect 43 412 92 422
rect 43 406 73 412
rect 92 407 97 412
rect 15 390 89 406
rect 107 398 137 454
rect 172 444 380 454
rect 415 450 460 454
rect 463 453 464 454
rect 479 453 492 454
rect 198 414 387 444
rect 213 411 387 414
rect 206 408 387 411
rect 15 388 28 390
rect 43 388 77 390
rect 15 372 89 388
rect 116 384 129 398
rect 144 384 160 400
rect 206 395 217 408
rect -1 350 0 366
rect 15 350 28 372
rect 43 350 73 372
rect 116 368 178 384
rect 206 377 217 393
rect 222 388 232 408
rect 242 388 256 408
rect 259 395 268 408
rect 284 395 293 408
rect 222 377 256 388
rect 259 377 268 393
rect 284 377 293 393
rect 300 388 310 408
rect 320 388 334 408
rect 335 395 346 408
rect 300 377 334 388
rect 335 377 346 393
rect 392 384 408 400
rect 415 398 445 450
rect 479 446 480 453
rect 464 438 480 446
rect 451 406 464 425
rect 479 406 509 422
rect 451 390 525 406
rect 451 388 464 390
rect 479 388 513 390
rect 116 366 129 368
rect 144 366 178 368
rect 116 350 178 366
rect 222 361 238 364
rect 300 361 330 372
rect 378 368 424 384
rect 451 372 525 388
rect 378 366 412 368
rect 377 350 424 366
rect 451 350 464 372
rect 479 350 509 372
rect 536 350 537 366
rect 552 350 565 510
rect 595 406 608 510
rect 653 488 654 498
rect 669 488 682 498
rect 653 484 682 488
rect 687 484 717 510
rect 735 496 751 498
rect 823 496 876 510
rect 824 494 888 496
rect 931 494 946 510
rect 995 507 1025 510
rect 995 504 1031 507
rect 961 496 977 498
rect 735 484 750 488
rect 653 482 750 484
rect 778 482 946 494
rect 962 484 977 488
rect 995 485 1034 504
rect 1053 498 1060 499
rect 1059 491 1060 498
rect 1043 488 1044 491
rect 1059 488 1072 491
rect 995 484 1025 485
rect 1034 484 1040 485
rect 1043 484 1072 488
rect 962 483 1072 484
rect 962 482 1078 483
rect 637 474 688 482
rect 637 462 662 474
rect 669 462 688 474
rect 719 474 769 482
rect 719 466 735 474
rect 742 472 769 474
rect 778 472 999 482
rect 742 462 999 472
rect 1028 474 1078 482
rect 1028 465 1044 474
rect 637 454 688 462
rect 735 454 999 462
rect 1025 462 1044 465
rect 1051 462 1078 474
rect 1025 454 1078 462
rect 653 446 654 454
rect 669 446 682 454
rect 653 438 669 446
rect 650 431 669 434
rect 650 422 672 431
rect 623 412 672 422
rect 623 406 653 412
rect 672 407 677 412
rect 595 390 669 406
rect 687 398 717 454
rect 752 444 960 454
rect 995 450 1040 454
rect 1043 453 1044 454
rect 1059 453 1072 454
rect 778 414 967 444
rect 793 411 967 414
rect 786 408 967 411
rect 595 388 608 390
rect 623 388 657 390
rect 595 372 669 388
rect 696 384 709 398
rect 724 384 740 400
rect 786 395 797 408
rect 579 350 580 366
rect 595 350 608 372
rect 623 350 653 372
rect 696 368 758 384
rect 786 377 797 393
rect 802 388 812 408
rect 822 388 836 408
rect 839 395 848 408
rect 864 395 873 408
rect 802 377 836 388
rect 839 377 848 393
rect 864 377 873 393
rect 880 388 890 408
rect 900 388 914 408
rect 915 395 926 408
rect 880 377 914 388
rect 915 377 926 393
rect 972 384 988 400
rect 995 398 1025 450
rect 1059 446 1060 453
rect 1044 438 1060 446
rect 1031 406 1044 425
rect 1059 406 1089 422
rect 1031 390 1105 406
rect 1031 388 1044 390
rect 1059 388 1093 390
rect 696 366 709 368
rect 724 366 758 368
rect 696 350 758 366
rect 802 361 818 364
rect 880 361 910 372
rect 958 368 1004 384
rect 1031 372 1105 388
rect 958 366 992 368
rect 957 350 1004 366
rect 1031 350 1044 372
rect 1059 350 1089 372
rect 1116 350 1117 366
rect 1132 350 1145 510
rect 1175 406 1188 510
rect 1233 488 1234 498
rect 1249 488 1262 498
rect 1233 484 1262 488
rect 1267 484 1297 510
rect 1315 496 1331 498
rect 1403 496 1456 510
rect 1404 494 1468 496
rect 1511 494 1526 510
rect 1575 507 1605 510
rect 1575 504 1611 507
rect 1541 496 1557 498
rect 1315 484 1330 488
rect 1233 482 1330 484
rect 1358 482 1526 494
rect 1542 484 1557 488
rect 1575 485 1614 504
rect 1633 498 1640 499
rect 1639 491 1640 498
rect 1623 488 1624 491
rect 1639 488 1652 491
rect 1575 484 1605 485
rect 1614 484 1620 485
rect 1623 484 1652 488
rect 1542 483 1652 484
rect 1542 482 1658 483
rect 1217 474 1268 482
rect 1217 462 1242 474
rect 1249 462 1268 474
rect 1299 474 1349 482
rect 1299 466 1315 474
rect 1322 472 1349 474
rect 1358 472 1579 482
rect 1322 462 1579 472
rect 1608 474 1658 482
rect 1608 465 1624 474
rect 1217 454 1268 462
rect 1315 454 1579 462
rect 1605 462 1624 465
rect 1631 462 1658 474
rect 1605 454 1658 462
rect 1233 446 1234 454
rect 1249 446 1262 454
rect 1233 438 1249 446
rect 1230 431 1249 434
rect 1230 422 1252 431
rect 1203 412 1252 422
rect 1203 406 1233 412
rect 1252 407 1257 412
rect 1175 390 1249 406
rect 1267 398 1297 454
rect 1332 444 1540 454
rect 1575 450 1620 454
rect 1623 453 1624 454
rect 1639 453 1652 454
rect 1358 414 1547 444
rect 1373 411 1547 414
rect 1366 408 1547 411
rect 1175 388 1188 390
rect 1203 388 1237 390
rect 1175 372 1249 388
rect 1276 384 1289 398
rect 1304 384 1320 400
rect 1366 395 1377 408
rect 1159 350 1160 366
rect 1175 350 1188 372
rect 1203 350 1233 372
rect 1276 368 1338 384
rect 1366 377 1377 393
rect 1382 388 1392 408
rect 1402 388 1416 408
rect 1419 395 1428 408
rect 1444 395 1453 408
rect 1382 377 1416 388
rect 1419 377 1428 393
rect 1444 377 1453 393
rect 1460 388 1470 408
rect 1480 388 1494 408
rect 1495 395 1506 408
rect 1460 377 1494 388
rect 1495 377 1506 393
rect 1552 384 1568 400
rect 1575 398 1605 450
rect 1639 446 1640 453
rect 1624 438 1640 446
rect 1611 406 1624 425
rect 1639 406 1669 422
rect 1611 390 1685 406
rect 1611 388 1624 390
rect 1639 388 1673 390
rect 1276 366 1289 368
rect 1304 366 1338 368
rect 1276 350 1338 366
rect 1382 361 1398 364
rect 1460 361 1490 372
rect 1538 368 1584 384
rect 1611 372 1685 388
rect 1538 366 1572 368
rect 1537 350 1584 366
rect 1611 350 1624 372
rect 1639 350 1669 372
rect 1696 350 1697 366
rect 1712 350 1725 510
rect 1755 406 1768 510
rect 1813 488 1814 498
rect 1829 488 1842 498
rect 1813 484 1842 488
rect 1847 484 1877 510
rect 1895 496 1911 498
rect 1983 496 2036 510
rect 1984 494 2048 496
rect 2091 494 2106 510
rect 2155 507 2185 510
rect 2155 504 2191 507
rect 2121 496 2137 498
rect 1895 484 1910 488
rect 1813 482 1910 484
rect 1938 482 2106 494
rect 2122 484 2137 488
rect 2155 485 2194 504
rect 2213 498 2220 499
rect 2219 491 2220 498
rect 2203 488 2204 491
rect 2219 488 2232 491
rect 2155 484 2185 485
rect 2194 484 2200 485
rect 2203 484 2232 488
rect 2122 483 2232 484
rect 2122 482 2238 483
rect 1797 474 1848 482
rect 1797 462 1822 474
rect 1829 462 1848 474
rect 1879 474 1929 482
rect 1879 466 1895 474
rect 1902 472 1929 474
rect 1938 472 2159 482
rect 1902 462 2159 472
rect 2188 474 2238 482
rect 2188 465 2204 474
rect 1797 454 1848 462
rect 1895 454 2159 462
rect 2185 462 2204 465
rect 2211 462 2238 474
rect 2185 454 2238 462
rect 1813 446 1814 454
rect 1829 446 1842 454
rect 1813 438 1829 446
rect 1810 431 1829 434
rect 1810 422 1832 431
rect 1783 412 1832 422
rect 1783 406 1813 412
rect 1832 407 1837 412
rect 1755 390 1829 406
rect 1847 398 1877 454
rect 1912 444 2120 454
rect 2155 450 2200 454
rect 2203 453 2204 454
rect 2219 453 2232 454
rect 1938 414 2127 444
rect 1953 411 2127 414
rect 1946 408 2127 411
rect 1755 388 1768 390
rect 1783 388 1817 390
rect 1755 372 1829 388
rect 1856 384 1869 398
rect 1884 384 1900 400
rect 1946 395 1957 408
rect 1739 350 1740 366
rect 1755 350 1768 372
rect 1783 350 1813 372
rect 1856 368 1918 384
rect 1946 377 1957 393
rect 1962 388 1972 408
rect 1982 388 1996 408
rect 1999 395 2008 408
rect 2024 395 2033 408
rect 1962 377 1996 388
rect 1999 377 2008 393
rect 2024 377 2033 393
rect 2040 388 2050 408
rect 2060 388 2074 408
rect 2075 395 2086 408
rect 2040 377 2074 388
rect 2075 377 2086 393
rect 2132 384 2148 400
rect 2155 398 2185 450
rect 2219 446 2220 453
rect 2204 438 2220 446
rect 2191 406 2204 425
rect 2219 406 2249 422
rect 2191 390 2265 406
rect 2191 388 2204 390
rect 2219 388 2253 390
rect 1856 366 1869 368
rect 1884 366 1918 368
rect 1856 350 1918 366
rect 1962 361 1978 364
rect 2040 361 2070 372
rect 2118 368 2164 384
rect 2191 372 2265 388
rect 2118 366 2152 368
rect 2117 350 2164 366
rect 2191 350 2204 372
rect 2219 350 2249 372
rect 2276 350 2277 366
rect 2292 350 2305 510
rect 2335 406 2348 510
rect 2393 488 2394 498
rect 2409 488 2422 498
rect 2393 484 2422 488
rect 2427 484 2457 510
rect 2475 496 2491 498
rect 2563 496 2616 510
rect 2564 494 2628 496
rect 2671 494 2686 510
rect 2735 507 2765 510
rect 2735 504 2771 507
rect 2701 496 2717 498
rect 2475 484 2490 488
rect 2393 482 2490 484
rect 2518 482 2686 494
rect 2702 484 2717 488
rect 2735 485 2774 504
rect 2793 498 2800 499
rect 2799 491 2800 498
rect 2783 488 2784 491
rect 2799 488 2812 491
rect 2735 484 2765 485
rect 2774 484 2780 485
rect 2783 484 2812 488
rect 2702 483 2812 484
rect 2702 482 2818 483
rect 2377 474 2428 482
rect 2377 462 2402 474
rect 2409 462 2428 474
rect 2459 474 2509 482
rect 2459 466 2475 474
rect 2482 472 2509 474
rect 2518 472 2739 482
rect 2482 462 2739 472
rect 2768 474 2818 482
rect 2768 465 2784 474
rect 2377 454 2428 462
rect 2475 454 2739 462
rect 2765 462 2784 465
rect 2791 462 2818 474
rect 2765 454 2818 462
rect 2393 446 2394 454
rect 2409 446 2422 454
rect 2393 438 2409 446
rect 2390 431 2409 434
rect 2390 422 2412 431
rect 2363 412 2412 422
rect 2363 406 2393 412
rect 2412 407 2417 412
rect 2335 390 2409 406
rect 2427 398 2457 454
rect 2492 444 2700 454
rect 2735 450 2780 454
rect 2783 453 2784 454
rect 2799 453 2812 454
rect 2518 414 2707 444
rect 2533 411 2707 414
rect 2526 408 2707 411
rect 2335 388 2348 390
rect 2363 388 2397 390
rect 2335 372 2409 388
rect 2436 384 2449 398
rect 2464 384 2480 400
rect 2526 395 2537 408
rect 2319 350 2320 366
rect 2335 350 2348 372
rect 2363 350 2393 372
rect 2436 368 2498 384
rect 2526 377 2537 393
rect 2542 388 2552 408
rect 2562 388 2576 408
rect 2579 395 2588 408
rect 2604 395 2613 408
rect 2542 377 2576 388
rect 2579 377 2588 393
rect 2604 377 2613 393
rect 2620 388 2630 408
rect 2640 388 2654 408
rect 2655 395 2666 408
rect 2620 377 2654 388
rect 2655 377 2666 393
rect 2712 384 2728 400
rect 2735 398 2765 450
rect 2799 446 2800 453
rect 2784 438 2800 446
rect 2771 406 2784 425
rect 2799 406 2829 422
rect 2771 390 2845 406
rect 2771 388 2784 390
rect 2799 388 2833 390
rect 2436 366 2449 368
rect 2464 366 2498 368
rect 2436 350 2498 366
rect 2542 361 2558 364
rect 2620 361 2650 372
rect 2698 368 2744 384
rect 2771 372 2845 388
rect 2698 366 2732 368
rect 2697 350 2744 366
rect 2771 350 2784 372
rect 2799 350 2829 372
rect 2856 350 2857 366
rect 2872 350 2885 510
rect 2915 406 2928 510
rect 2973 488 2974 498
rect 2989 488 3002 498
rect 2973 484 3002 488
rect 3007 484 3037 510
rect 3055 496 3071 498
rect 3143 496 3196 510
rect 3144 494 3208 496
rect 3251 494 3266 510
rect 3315 507 3345 510
rect 3315 504 3351 507
rect 3281 496 3297 498
rect 3055 484 3070 488
rect 2973 482 3070 484
rect 3098 482 3266 494
rect 3282 484 3297 488
rect 3315 485 3354 504
rect 3373 498 3380 499
rect 3379 491 3380 498
rect 3363 488 3364 491
rect 3379 488 3392 491
rect 3315 484 3345 485
rect 3354 484 3360 485
rect 3363 484 3392 488
rect 3282 483 3392 484
rect 3282 482 3398 483
rect 2957 474 3008 482
rect 2957 462 2982 474
rect 2989 462 3008 474
rect 3039 474 3089 482
rect 3039 466 3055 474
rect 3062 472 3089 474
rect 3098 472 3319 482
rect 3062 462 3319 472
rect 3348 474 3398 482
rect 3348 465 3364 474
rect 2957 454 3008 462
rect 3055 454 3319 462
rect 3345 462 3364 465
rect 3371 462 3398 474
rect 3345 454 3398 462
rect 2973 446 2974 454
rect 2989 446 3002 454
rect 2973 438 2989 446
rect 2970 431 2989 434
rect 2970 422 2992 431
rect 2943 412 2992 422
rect 2943 406 2973 412
rect 2992 407 2997 412
rect 2915 390 2989 406
rect 3007 398 3037 454
rect 3072 444 3280 454
rect 3315 450 3360 454
rect 3363 453 3364 454
rect 3379 453 3392 454
rect 3098 414 3287 444
rect 3113 411 3287 414
rect 3106 408 3287 411
rect 2915 388 2928 390
rect 2943 388 2977 390
rect 2915 372 2989 388
rect 3016 384 3029 398
rect 3044 384 3060 400
rect 3106 395 3117 408
rect 2899 350 2900 366
rect 2915 350 2928 372
rect 2943 350 2973 372
rect 3016 368 3078 384
rect 3106 377 3117 393
rect 3122 388 3132 408
rect 3142 388 3156 408
rect 3159 395 3168 408
rect 3184 395 3193 408
rect 3122 377 3156 388
rect 3159 377 3168 393
rect 3184 377 3193 393
rect 3200 388 3210 408
rect 3220 388 3234 408
rect 3235 395 3246 408
rect 3200 377 3234 388
rect 3235 377 3246 393
rect 3292 384 3308 400
rect 3315 398 3345 450
rect 3379 446 3380 453
rect 3364 438 3380 446
rect 3351 406 3364 425
rect 3379 406 3409 422
rect 3351 390 3425 406
rect 3351 388 3364 390
rect 3379 388 3413 390
rect 3016 366 3029 368
rect 3044 366 3078 368
rect 3016 350 3078 366
rect 3122 361 3138 364
rect 3200 361 3230 372
rect 3278 368 3324 384
rect 3351 372 3425 388
rect 3278 366 3312 368
rect 3277 350 3324 366
rect 3351 350 3364 372
rect 3379 350 3409 372
rect 3436 350 3437 366
rect 3452 350 3465 510
rect 3495 406 3508 510
rect 3553 488 3554 498
rect 3569 488 3582 498
rect 3553 484 3582 488
rect 3587 484 3617 510
rect 3635 496 3651 498
rect 3723 496 3776 510
rect 3724 494 3788 496
rect 3831 494 3846 510
rect 3895 507 3925 510
rect 3895 504 3931 507
rect 3861 496 3877 498
rect 3635 484 3650 488
rect 3553 482 3650 484
rect 3678 482 3846 494
rect 3862 484 3877 488
rect 3895 485 3934 504
rect 3953 498 3960 499
rect 3959 491 3960 498
rect 3943 488 3944 491
rect 3959 488 3972 491
rect 3895 484 3925 485
rect 3934 484 3940 485
rect 3943 484 3972 488
rect 3862 483 3972 484
rect 3862 482 3978 483
rect 3537 474 3588 482
rect 3537 462 3562 474
rect 3569 462 3588 474
rect 3619 474 3669 482
rect 3619 466 3635 474
rect 3642 472 3669 474
rect 3678 472 3899 482
rect 3642 462 3899 472
rect 3928 474 3978 482
rect 3928 465 3944 474
rect 3537 454 3588 462
rect 3635 454 3899 462
rect 3925 462 3944 465
rect 3951 462 3978 474
rect 3925 454 3978 462
rect 3553 446 3554 454
rect 3569 446 3582 454
rect 3553 438 3569 446
rect 3550 431 3569 434
rect 3550 422 3572 431
rect 3523 412 3572 422
rect 3523 406 3553 412
rect 3572 407 3577 412
rect 3495 390 3569 406
rect 3587 398 3617 454
rect 3652 444 3860 454
rect 3895 450 3940 454
rect 3943 453 3944 454
rect 3959 453 3972 454
rect 3678 414 3867 444
rect 3693 411 3867 414
rect 3686 408 3867 411
rect 3495 388 3508 390
rect 3523 388 3557 390
rect 3495 372 3569 388
rect 3596 384 3609 398
rect 3624 384 3640 400
rect 3686 395 3697 408
rect 3479 350 3480 366
rect 3495 350 3508 372
rect 3523 350 3553 372
rect 3596 368 3658 384
rect 3686 377 3697 393
rect 3702 388 3712 408
rect 3722 388 3736 408
rect 3739 395 3748 408
rect 3764 395 3773 408
rect 3702 377 3736 388
rect 3739 377 3748 393
rect 3764 377 3773 393
rect 3780 388 3790 408
rect 3800 388 3814 408
rect 3815 395 3826 408
rect 3780 377 3814 388
rect 3815 377 3826 393
rect 3872 384 3888 400
rect 3895 398 3925 450
rect 3959 446 3960 453
rect 3944 438 3960 446
rect 3931 406 3944 425
rect 3959 406 3989 422
rect 3931 390 4005 406
rect 3931 388 3944 390
rect 3959 388 3993 390
rect 3596 366 3609 368
rect 3624 366 3658 368
rect 3596 350 3658 366
rect 3702 361 3718 364
rect 3780 361 3810 372
rect 3858 368 3904 384
rect 3931 372 4005 388
rect 3858 366 3892 368
rect 3857 350 3904 366
rect 3931 350 3944 372
rect 3959 350 3989 372
rect 4016 350 4017 366
rect 4032 350 4045 510
rect 4075 406 4088 510
rect 4133 488 4134 498
rect 4149 488 4162 498
rect 4133 484 4162 488
rect 4167 484 4197 510
rect 4215 496 4231 498
rect 4303 496 4356 510
rect 4304 494 4368 496
rect 4411 494 4426 510
rect 4475 507 4505 510
rect 4475 504 4511 507
rect 4441 496 4457 498
rect 4215 484 4230 488
rect 4133 482 4230 484
rect 4258 482 4426 494
rect 4442 484 4457 488
rect 4475 485 4514 504
rect 4533 498 4540 499
rect 4539 491 4540 498
rect 4523 488 4524 491
rect 4539 488 4552 491
rect 4475 484 4505 485
rect 4514 484 4520 485
rect 4523 484 4552 488
rect 4442 483 4552 484
rect 4442 482 4558 483
rect 4117 474 4168 482
rect 4117 462 4142 474
rect 4149 462 4168 474
rect 4199 474 4249 482
rect 4199 466 4215 474
rect 4222 472 4249 474
rect 4258 472 4479 482
rect 4222 462 4479 472
rect 4508 474 4558 482
rect 4508 465 4524 474
rect 4117 454 4168 462
rect 4215 454 4479 462
rect 4505 462 4524 465
rect 4531 462 4558 474
rect 4505 454 4558 462
rect 4133 446 4134 454
rect 4149 446 4162 454
rect 4133 438 4149 446
rect 4130 431 4149 434
rect 4130 422 4152 431
rect 4103 412 4152 422
rect 4103 406 4133 412
rect 4152 407 4157 412
rect 4075 390 4149 406
rect 4167 398 4197 454
rect 4232 444 4440 454
rect 4475 450 4520 454
rect 4523 453 4524 454
rect 4539 453 4552 454
rect 4258 414 4447 444
rect 4273 411 4447 414
rect 4266 408 4447 411
rect 4075 388 4088 390
rect 4103 388 4137 390
rect 4075 372 4149 388
rect 4176 384 4189 398
rect 4204 384 4220 400
rect 4266 395 4277 408
rect 4059 350 4060 366
rect 4075 350 4088 372
rect 4103 350 4133 372
rect 4176 368 4238 384
rect 4266 377 4277 393
rect 4282 388 4292 408
rect 4302 388 4316 408
rect 4319 395 4328 408
rect 4344 395 4353 408
rect 4282 377 4316 388
rect 4319 377 4328 393
rect 4344 377 4353 393
rect 4360 388 4370 408
rect 4380 388 4394 408
rect 4395 395 4406 408
rect 4360 377 4394 388
rect 4395 377 4406 393
rect 4452 384 4468 400
rect 4475 398 4505 450
rect 4539 446 4540 453
rect 4524 438 4540 446
rect 4511 406 4524 425
rect 4539 406 4569 422
rect 4511 390 4585 406
rect 4511 388 4524 390
rect 4539 388 4573 390
rect 4176 366 4189 368
rect 4204 366 4238 368
rect 4176 350 4238 366
rect 4282 361 4298 364
rect 4360 361 4390 372
rect 4438 368 4484 384
rect 4511 372 4585 388
rect 4438 366 4472 368
rect 4437 350 4484 366
rect 4511 350 4524 372
rect 4539 350 4569 372
rect 4596 350 4597 366
rect 4612 350 4625 510
rect -7 342 34 350
rect -7 316 8 342
rect 15 316 34 342
rect 98 338 160 350
rect 172 338 247 350
rect 305 338 380 350
rect 392 338 423 350
rect 429 338 464 350
rect 98 336 260 338
rect -7 308 34 316
rect 116 312 129 336
rect 144 334 159 336
rect -1 298 0 308
rect 15 298 28 308
rect 43 298 73 312
rect 116 298 159 312
rect 183 309 190 316
rect 193 312 260 336
rect 292 336 464 338
rect 262 314 290 318
rect 292 314 372 336
rect 393 334 408 336
rect 262 312 372 314
rect 193 308 372 312
rect 166 298 196 308
rect 198 298 351 308
rect 359 298 389 308
rect 393 298 423 312
rect 451 298 464 336
rect 536 342 571 350
rect 536 316 537 342
rect 544 316 571 342
rect 479 298 509 312
rect 536 308 571 316
rect 573 342 614 350
rect 573 316 588 342
rect 595 316 614 342
rect 678 338 740 350
rect 752 338 827 350
rect 885 338 960 350
rect 972 338 1003 350
rect 1009 338 1044 350
rect 678 336 840 338
rect 573 308 614 316
rect 696 312 709 336
rect 724 334 739 336
rect 536 298 537 308
rect 552 298 565 308
rect 579 298 580 308
rect 595 298 608 308
rect 623 298 653 312
rect 696 298 739 312
rect 763 309 770 316
rect 773 312 840 336
rect 872 336 1044 338
rect 842 314 870 318
rect 872 314 952 336
rect 973 334 988 336
rect 842 312 952 314
rect 773 308 952 312
rect 746 298 776 308
rect 778 298 931 308
rect 939 298 969 308
rect 973 298 1003 312
rect 1031 298 1044 336
rect 1116 342 1151 350
rect 1116 316 1117 342
rect 1124 316 1151 342
rect 1059 298 1089 312
rect 1116 308 1151 316
rect 1153 342 1194 350
rect 1153 316 1168 342
rect 1175 316 1194 342
rect 1258 338 1320 350
rect 1332 338 1407 350
rect 1465 338 1540 350
rect 1552 338 1583 350
rect 1589 338 1624 350
rect 1258 336 1420 338
rect 1153 308 1194 316
rect 1276 312 1289 336
rect 1304 334 1319 336
rect 1116 298 1117 308
rect 1132 298 1145 308
rect 1159 298 1160 308
rect 1175 298 1188 308
rect 1203 298 1233 312
rect 1276 298 1319 312
rect 1343 309 1350 316
rect 1353 312 1420 336
rect 1452 336 1624 338
rect 1422 314 1450 318
rect 1452 314 1532 336
rect 1553 334 1568 336
rect 1422 312 1532 314
rect 1353 308 1532 312
rect 1326 298 1356 308
rect 1358 298 1511 308
rect 1519 298 1549 308
rect 1553 298 1583 312
rect 1611 298 1624 336
rect 1696 342 1731 350
rect 1696 316 1697 342
rect 1704 316 1731 342
rect 1639 298 1669 312
rect 1696 308 1731 316
rect 1733 342 1774 350
rect 1733 316 1748 342
rect 1755 316 1774 342
rect 1838 338 1900 350
rect 1912 338 1987 350
rect 2045 338 2120 350
rect 2132 338 2163 350
rect 2169 338 2204 350
rect 1838 336 2000 338
rect 1733 308 1774 316
rect 1856 312 1869 336
rect 1884 334 1899 336
rect 1696 298 1697 308
rect 1712 298 1725 308
rect 1739 298 1740 308
rect 1755 298 1768 308
rect 1783 298 1813 312
rect 1856 298 1899 312
rect 1923 309 1930 316
rect 1933 312 2000 336
rect 2032 336 2204 338
rect 2002 314 2030 318
rect 2032 314 2112 336
rect 2133 334 2148 336
rect 2002 312 2112 314
rect 1933 308 2112 312
rect 1906 298 1936 308
rect 1938 298 2091 308
rect 2099 298 2129 308
rect 2133 298 2163 312
rect 2191 298 2204 336
rect 2276 342 2311 350
rect 2276 316 2277 342
rect 2284 316 2311 342
rect 2219 298 2249 312
rect 2276 308 2311 316
rect 2313 342 2354 350
rect 2313 316 2328 342
rect 2335 316 2354 342
rect 2418 338 2480 350
rect 2492 338 2567 350
rect 2625 338 2700 350
rect 2712 338 2743 350
rect 2749 338 2784 350
rect 2418 336 2580 338
rect 2313 308 2354 316
rect 2436 312 2449 336
rect 2464 334 2479 336
rect 2276 298 2277 308
rect 2292 298 2305 308
rect 2319 298 2320 308
rect 2335 298 2348 308
rect 2363 298 2393 312
rect 2436 298 2479 312
rect 2503 309 2510 316
rect 2513 312 2580 336
rect 2612 336 2784 338
rect 2582 314 2610 318
rect 2612 314 2692 336
rect 2713 334 2728 336
rect 2582 312 2692 314
rect 2513 308 2692 312
rect 2486 298 2516 308
rect 2518 298 2671 308
rect 2679 298 2709 308
rect 2713 298 2743 312
rect 2771 298 2784 336
rect 2856 342 2891 350
rect 2856 316 2857 342
rect 2864 316 2891 342
rect 2799 298 2829 312
rect 2856 308 2891 316
rect 2893 342 2934 350
rect 2893 316 2908 342
rect 2915 316 2934 342
rect 2998 338 3060 350
rect 3072 338 3147 350
rect 3205 338 3280 350
rect 3292 338 3323 350
rect 3329 338 3364 350
rect 2998 336 3160 338
rect 2893 308 2934 316
rect 3016 312 3029 336
rect 3044 334 3059 336
rect 2856 298 2857 308
rect 2872 298 2885 308
rect 2899 298 2900 308
rect 2915 298 2928 308
rect 2943 298 2973 312
rect 3016 298 3059 312
rect 3083 309 3090 316
rect 3093 312 3160 336
rect 3192 336 3364 338
rect 3162 314 3190 318
rect 3192 314 3272 336
rect 3293 334 3308 336
rect 3162 312 3272 314
rect 3093 308 3272 312
rect 3066 298 3096 308
rect 3098 298 3251 308
rect 3259 298 3289 308
rect 3293 298 3323 312
rect 3351 298 3364 336
rect 3436 342 3471 350
rect 3436 316 3437 342
rect 3444 316 3471 342
rect 3379 298 3409 312
rect 3436 308 3471 316
rect 3473 342 3514 350
rect 3473 316 3488 342
rect 3495 316 3514 342
rect 3578 338 3640 350
rect 3652 338 3727 350
rect 3785 338 3860 350
rect 3872 338 3903 350
rect 3909 338 3944 350
rect 3578 336 3740 338
rect 3473 308 3514 316
rect 3596 312 3609 336
rect 3624 334 3639 336
rect 3436 298 3437 308
rect 3452 298 3465 308
rect 3479 298 3480 308
rect 3495 298 3508 308
rect 3523 298 3553 312
rect 3596 298 3639 312
rect 3663 309 3670 316
rect 3673 312 3740 336
rect 3772 336 3944 338
rect 3742 314 3770 318
rect 3772 314 3852 336
rect 3873 334 3888 336
rect 3742 312 3852 314
rect 3673 308 3852 312
rect 3646 298 3676 308
rect 3678 298 3831 308
rect 3839 298 3869 308
rect 3873 298 3903 312
rect 3931 298 3944 336
rect 4016 342 4051 350
rect 4016 316 4017 342
rect 4024 316 4051 342
rect 3959 298 3989 312
rect 4016 308 4051 316
rect 4053 342 4094 350
rect 4053 316 4068 342
rect 4075 316 4094 342
rect 4158 338 4220 350
rect 4232 338 4307 350
rect 4365 338 4440 350
rect 4452 338 4483 350
rect 4489 338 4524 350
rect 4158 336 4320 338
rect 4053 308 4094 316
rect 4176 312 4189 336
rect 4204 334 4219 336
rect 4016 298 4017 308
rect 4032 298 4045 308
rect 4059 298 4060 308
rect 4075 298 4088 308
rect 4103 298 4133 312
rect 4176 298 4219 312
rect 4243 309 4250 316
rect 4253 312 4320 336
rect 4352 336 4524 338
rect 4322 314 4350 318
rect 4352 314 4432 336
rect 4453 334 4468 336
rect 4322 312 4432 314
rect 4253 308 4432 312
rect 4226 298 4256 308
rect 4258 298 4411 308
rect 4419 298 4449 308
rect 4453 298 4483 312
rect 4511 298 4524 336
rect 4596 342 4631 350
rect 4596 316 4597 342
rect 4604 316 4631 342
rect 4539 298 4569 312
rect 4596 308 4631 316
rect 4596 298 4597 308
rect 4612 298 4625 308
rect -1 292 4625 298
rect 0 284 4625 292
rect 15 254 28 284
rect 43 266 73 284
rect 116 270 130 284
rect 166 270 386 284
rect 117 268 130 270
rect 83 256 98 268
rect 80 254 102 256
rect 107 254 137 268
rect 198 266 351 270
rect 180 254 372 266
rect 415 254 445 268
rect 451 254 464 284
rect 479 266 509 284
rect 552 254 565 284
rect 595 254 608 284
rect 623 266 653 284
rect 696 270 710 284
rect 746 270 966 284
rect 697 268 710 270
rect 663 256 678 268
rect 660 254 682 256
rect 687 254 717 268
rect 778 266 931 270
rect 760 254 952 266
rect 995 254 1025 268
rect 1031 254 1044 284
rect 1059 266 1089 284
rect 1132 254 1145 284
rect 1175 254 1188 284
rect 1203 266 1233 284
rect 1276 270 1290 284
rect 1326 270 1546 284
rect 1277 268 1290 270
rect 1243 256 1258 268
rect 1240 254 1262 256
rect 1267 254 1297 268
rect 1358 266 1511 270
rect 1340 254 1532 266
rect 1575 254 1605 268
rect 1611 254 1624 284
rect 1639 266 1669 284
rect 1712 254 1725 284
rect 1755 254 1768 284
rect 1783 266 1813 284
rect 1856 270 1870 284
rect 1906 270 2126 284
rect 1857 268 1870 270
rect 1823 256 1838 268
rect 1820 254 1842 256
rect 1847 254 1877 268
rect 1938 266 2091 270
rect 1920 254 2112 266
rect 2155 254 2185 268
rect 2191 254 2204 284
rect 2219 266 2249 284
rect 2292 254 2305 284
rect 2335 254 2348 284
rect 2363 266 2393 284
rect 2436 270 2450 284
rect 2486 270 2706 284
rect 2437 268 2450 270
rect 2403 256 2418 268
rect 2400 254 2422 256
rect 2427 254 2457 268
rect 2518 266 2671 270
rect 2500 254 2692 266
rect 2735 254 2765 268
rect 2771 254 2784 284
rect 2799 266 2829 284
rect 2872 254 2885 284
rect 2915 254 2928 284
rect 2943 266 2973 284
rect 3016 270 3030 284
rect 3066 270 3286 284
rect 3017 268 3030 270
rect 2983 256 2998 268
rect 2980 254 3002 256
rect 3007 254 3037 268
rect 3098 266 3251 270
rect 3080 254 3272 266
rect 3315 254 3345 268
rect 3351 254 3364 284
rect 3379 266 3409 284
rect 3452 254 3465 284
rect 3495 254 3508 284
rect 3523 266 3553 284
rect 3596 270 3610 284
rect 3646 270 3866 284
rect 3597 268 3610 270
rect 3563 256 3578 268
rect 3560 254 3582 256
rect 3587 254 3617 268
rect 3678 266 3831 270
rect 3660 254 3852 266
rect 3895 254 3925 268
rect 3931 254 3944 284
rect 3959 266 3989 284
rect 4032 254 4045 284
rect 4075 254 4088 284
rect 4103 266 4133 284
rect 4176 270 4190 284
rect 4226 270 4446 284
rect 4177 268 4190 270
rect 4143 256 4158 268
rect 4140 254 4162 256
rect 4167 254 4197 268
rect 4258 266 4411 270
rect 4240 254 4432 266
rect 4475 254 4505 268
rect 4511 254 4524 284
rect 4539 266 4569 284
rect 4612 254 4625 284
rect 0 240 4625 254
rect 15 136 28 240
rect 73 218 74 228
rect 89 218 102 228
rect 73 214 102 218
rect 107 214 137 240
rect 155 226 171 228
rect 243 226 296 240
rect 244 224 308 226
rect 155 214 170 218
rect 73 212 170 214
rect 57 204 108 212
rect 57 192 82 204
rect 89 192 108 204
rect 139 204 189 212
rect 139 196 155 204
rect 162 202 189 204
rect 198 204 213 208
rect 260 204 292 224
rect 351 212 366 240
rect 415 237 445 240
rect 415 234 451 237
rect 381 226 397 228
rect 382 214 397 218
rect 415 215 454 234
rect 473 228 480 229
rect 479 221 480 228
rect 463 218 464 221
rect 479 218 492 221
rect 415 214 445 215
rect 454 214 460 215
rect 463 214 492 218
rect 382 213 492 214
rect 382 212 498 213
rect 351 204 419 212
rect 198 202 267 204
rect 285 202 419 204
rect 162 198 234 202
rect 162 196 287 198
rect 162 192 234 196
rect 57 184 108 192
rect 155 188 234 192
rect 315 188 419 202
rect 448 204 498 212
rect 448 195 464 204
rect 155 184 419 188
rect 445 192 464 195
rect 471 192 498 204
rect 445 184 498 192
rect 73 176 74 184
rect 89 176 102 184
rect 73 168 89 176
rect 70 161 89 164
rect 70 152 92 161
rect 43 142 92 152
rect 43 136 73 142
rect 92 137 97 142
rect 15 120 89 136
rect 107 128 137 184
rect 172 174 380 184
rect 415 180 460 184
rect 463 183 464 184
rect 479 183 492 184
rect 339 170 387 174
rect 222 148 252 157
rect 315 150 330 157
rect 351 148 387 170
rect 198 144 387 148
rect 213 141 387 144
rect 206 138 387 141
rect 15 118 28 120
rect 43 118 77 120
rect 15 102 89 118
rect 116 114 129 128
rect 144 114 160 130
rect 206 125 217 138
rect -1 80 0 96
rect 15 80 28 102
rect 43 80 73 102
rect 116 98 178 114
rect 206 107 217 123
rect 222 118 232 138
rect 242 118 256 138
rect 259 125 268 138
rect 284 125 293 138
rect 222 107 256 118
rect 259 107 267 123
rect 284 107 293 123
rect 300 118 310 138
rect 320 118 334 138
rect 335 125 346 138
rect 300 107 334 118
rect 335 107 346 123
rect 392 114 408 130
rect 415 128 445 180
rect 479 176 480 183
rect 464 168 480 176
rect 451 136 464 155
rect 479 136 509 152
rect 451 120 525 136
rect 451 118 464 120
rect 479 118 513 120
rect 116 96 129 98
rect 144 96 178 98
rect 116 80 178 96
rect 222 91 235 94
rect 300 91 330 102
rect 378 98 424 114
rect 451 102 525 118
rect 378 96 412 98
rect 377 80 424 96
rect 451 80 464 102
rect 479 80 509 102
rect 536 80 537 96
rect 552 80 565 240
rect 595 136 608 240
rect 653 218 654 228
rect 669 218 682 228
rect 653 214 682 218
rect 687 214 717 240
rect 735 226 751 228
rect 823 226 876 240
rect 824 224 888 226
rect 735 214 750 218
rect 653 212 750 214
rect 637 204 688 212
rect 637 192 662 204
rect 669 192 688 204
rect 719 204 769 212
rect 719 196 735 204
rect 742 202 769 204
rect 778 204 793 208
rect 840 204 872 224
rect 931 212 946 240
rect 995 237 1025 240
rect 995 234 1031 237
rect 961 226 977 228
rect 962 214 977 218
rect 995 215 1034 234
rect 1053 228 1060 229
rect 1059 221 1060 228
rect 1043 218 1044 221
rect 1059 218 1072 221
rect 995 214 1025 215
rect 1034 214 1040 215
rect 1043 214 1072 218
rect 962 213 1072 214
rect 962 212 1078 213
rect 931 204 999 212
rect 778 202 847 204
rect 865 202 999 204
rect 742 198 814 202
rect 742 196 867 198
rect 742 192 814 196
rect 637 184 688 192
rect 735 188 814 192
rect 895 188 999 202
rect 1028 204 1078 212
rect 1028 195 1044 204
rect 735 184 999 188
rect 1025 192 1044 195
rect 1051 192 1078 204
rect 1025 184 1078 192
rect 653 176 654 184
rect 669 176 682 184
rect 653 168 669 176
rect 650 161 669 164
rect 650 152 672 161
rect 623 142 672 152
rect 623 136 653 142
rect 672 137 677 142
rect 595 120 669 136
rect 687 128 717 184
rect 752 174 960 184
rect 995 180 1040 184
rect 1043 183 1044 184
rect 1059 183 1072 184
rect 919 170 967 174
rect 802 148 832 157
rect 895 150 910 157
rect 931 148 967 170
rect 778 144 967 148
rect 793 141 967 144
rect 786 138 967 141
rect 595 118 608 120
rect 623 118 657 120
rect 595 102 669 118
rect 696 114 709 128
rect 724 114 740 130
rect 786 125 797 138
rect 579 80 580 96
rect 595 80 608 102
rect 623 80 653 102
rect 696 98 758 114
rect 786 107 797 123
rect 802 118 812 138
rect 822 118 836 138
rect 839 125 848 138
rect 864 125 873 138
rect 802 107 836 118
rect 839 107 847 123
rect 864 107 873 123
rect 880 118 890 138
rect 900 118 914 138
rect 915 125 926 138
rect 880 107 914 118
rect 915 107 926 123
rect 972 114 988 130
rect 995 128 1025 180
rect 1059 176 1060 183
rect 1044 168 1060 176
rect 1031 136 1044 155
rect 1059 136 1089 152
rect 1031 120 1105 136
rect 1031 118 1044 120
rect 1059 118 1093 120
rect 696 96 709 98
rect 724 96 758 98
rect 696 80 758 96
rect 802 91 815 94
rect 880 91 910 102
rect 958 98 1004 114
rect 1031 102 1105 118
rect 958 96 992 98
rect 957 80 1004 96
rect 1031 80 1044 102
rect 1059 80 1089 102
rect 1116 80 1117 96
rect 1132 80 1145 240
rect 1175 136 1188 240
rect 1233 218 1234 228
rect 1249 218 1262 228
rect 1233 214 1262 218
rect 1267 214 1297 240
rect 1315 226 1331 228
rect 1403 226 1456 240
rect 1404 224 1468 226
rect 1315 214 1330 218
rect 1233 212 1330 214
rect 1217 204 1268 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1299 204 1349 212
rect 1299 196 1315 204
rect 1322 202 1349 204
rect 1358 204 1373 208
rect 1420 204 1452 224
rect 1511 212 1526 240
rect 1575 237 1605 240
rect 1575 234 1611 237
rect 1541 226 1557 228
rect 1542 214 1557 218
rect 1575 215 1614 234
rect 1633 228 1640 229
rect 1639 221 1640 228
rect 1623 218 1624 221
rect 1639 218 1652 221
rect 1575 214 1605 215
rect 1614 214 1620 215
rect 1623 214 1652 218
rect 1542 213 1652 214
rect 1542 212 1658 213
rect 1511 204 1579 212
rect 1358 202 1427 204
rect 1445 202 1579 204
rect 1322 198 1394 202
rect 1322 196 1447 198
rect 1322 192 1394 196
rect 1217 184 1268 192
rect 1315 188 1394 192
rect 1475 188 1579 202
rect 1608 204 1658 212
rect 1608 195 1624 204
rect 1315 184 1579 188
rect 1605 192 1624 195
rect 1631 192 1658 204
rect 1605 184 1658 192
rect 1233 176 1234 184
rect 1249 176 1262 184
rect 1233 168 1249 176
rect 1230 161 1249 164
rect 1230 152 1252 161
rect 1203 142 1252 152
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1175 120 1249 136
rect 1267 128 1297 184
rect 1332 174 1540 184
rect 1575 180 1620 184
rect 1623 183 1624 184
rect 1639 183 1652 184
rect 1499 170 1547 174
rect 1382 148 1412 157
rect 1475 150 1490 157
rect 1511 148 1547 170
rect 1358 144 1547 148
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1175 118 1188 120
rect 1203 118 1237 120
rect 1175 102 1249 118
rect 1276 114 1289 128
rect 1304 114 1320 130
rect 1366 125 1377 138
rect 1159 80 1160 96
rect 1175 80 1188 102
rect 1203 80 1233 102
rect 1276 98 1338 114
rect 1366 107 1377 123
rect 1382 118 1392 138
rect 1402 118 1416 138
rect 1419 125 1428 138
rect 1444 125 1453 138
rect 1382 107 1416 118
rect 1419 107 1427 123
rect 1444 107 1453 123
rect 1460 118 1470 138
rect 1480 118 1494 138
rect 1495 125 1506 138
rect 1460 107 1494 118
rect 1495 107 1506 123
rect 1552 114 1568 130
rect 1575 128 1605 180
rect 1639 176 1640 183
rect 1624 168 1640 176
rect 1611 136 1624 155
rect 1639 136 1669 152
rect 1611 120 1685 136
rect 1611 118 1624 120
rect 1639 118 1673 120
rect 1276 96 1289 98
rect 1304 96 1338 98
rect 1276 80 1338 96
rect 1382 91 1395 94
rect 1460 91 1490 102
rect 1538 98 1584 114
rect 1611 102 1685 118
rect 1538 96 1572 98
rect 1537 80 1584 96
rect 1611 80 1624 102
rect 1639 80 1669 102
rect 1696 80 1697 96
rect 1712 80 1725 240
rect 1755 136 1768 240
rect 1813 218 1814 228
rect 1829 218 1842 228
rect 1813 214 1842 218
rect 1847 214 1877 240
rect 1895 226 1911 228
rect 1983 226 2036 240
rect 1984 224 2048 226
rect 1895 214 1910 218
rect 1813 212 1910 214
rect 1797 204 1848 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1879 204 1929 212
rect 1879 196 1895 204
rect 1902 202 1929 204
rect 1938 204 1953 208
rect 2000 204 2032 224
rect 2091 212 2106 240
rect 2155 237 2185 240
rect 2155 234 2191 237
rect 2121 226 2137 228
rect 2122 214 2137 218
rect 2155 215 2194 234
rect 2213 228 2220 229
rect 2219 221 2220 228
rect 2203 218 2204 221
rect 2219 218 2232 221
rect 2155 214 2185 215
rect 2194 214 2200 215
rect 2203 214 2232 218
rect 2122 213 2232 214
rect 2122 212 2238 213
rect 2091 204 2159 212
rect 1938 202 2007 204
rect 2025 202 2159 204
rect 1902 198 1974 202
rect 1902 196 2027 198
rect 1902 192 1974 196
rect 1797 184 1848 192
rect 1895 188 1974 192
rect 2055 188 2159 202
rect 2188 204 2238 212
rect 2188 195 2204 204
rect 1895 184 2159 188
rect 2185 192 2204 195
rect 2211 192 2238 204
rect 2185 184 2238 192
rect 1813 176 1814 184
rect 1829 176 1842 184
rect 1813 168 1829 176
rect 1810 161 1829 164
rect 1810 152 1832 161
rect 1783 142 1832 152
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1755 120 1829 136
rect 1847 128 1877 184
rect 1912 174 2120 184
rect 2155 180 2200 184
rect 2203 183 2204 184
rect 2219 183 2232 184
rect 2079 170 2127 174
rect 1962 148 1992 157
rect 2055 150 2070 157
rect 2091 148 2127 170
rect 1938 144 2127 148
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 1755 118 1768 120
rect 1783 118 1817 120
rect 1755 102 1829 118
rect 1856 114 1869 128
rect 1884 114 1900 130
rect 1946 125 1957 138
rect 1739 80 1740 96
rect 1755 80 1768 102
rect 1783 80 1813 102
rect 1856 98 1918 114
rect 1946 107 1957 123
rect 1962 118 1972 138
rect 1982 118 1996 138
rect 1999 125 2008 138
rect 2024 125 2033 138
rect 1962 107 1996 118
rect 1999 107 2007 123
rect 2024 107 2033 123
rect 2040 118 2050 138
rect 2060 118 2074 138
rect 2075 125 2086 138
rect 2040 107 2074 118
rect 2075 107 2086 123
rect 2132 114 2148 130
rect 2155 128 2185 180
rect 2219 176 2220 183
rect 2204 168 2220 176
rect 2191 136 2204 155
rect 2219 136 2249 152
rect 2191 120 2265 136
rect 2191 118 2204 120
rect 2219 118 2253 120
rect 1856 96 1869 98
rect 1884 96 1918 98
rect 1856 80 1918 96
rect 1962 91 1975 94
rect 2040 91 2070 102
rect 2118 98 2164 114
rect 2191 102 2265 118
rect 2118 96 2152 98
rect 2117 80 2164 96
rect 2191 80 2204 102
rect 2219 80 2249 102
rect 2276 80 2277 96
rect 2292 80 2305 240
rect 2335 136 2348 240
rect 2393 218 2394 228
rect 2409 218 2422 228
rect 2393 214 2422 218
rect 2427 214 2457 240
rect 2475 226 2491 228
rect 2563 226 2616 240
rect 2564 224 2628 226
rect 2475 214 2490 218
rect 2393 212 2490 214
rect 2377 204 2428 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2459 204 2509 212
rect 2459 196 2475 204
rect 2482 202 2509 204
rect 2518 204 2533 208
rect 2580 204 2612 224
rect 2671 212 2686 240
rect 2735 237 2765 240
rect 2735 234 2771 237
rect 2701 226 2717 228
rect 2702 214 2717 218
rect 2735 215 2774 234
rect 2793 228 2800 229
rect 2799 221 2800 228
rect 2783 218 2784 221
rect 2799 218 2812 221
rect 2735 214 2765 215
rect 2774 214 2780 215
rect 2783 214 2812 218
rect 2702 213 2812 214
rect 2702 212 2818 213
rect 2671 204 2739 212
rect 2518 202 2587 204
rect 2605 202 2739 204
rect 2482 198 2554 202
rect 2482 196 2607 198
rect 2482 192 2554 196
rect 2377 184 2428 192
rect 2475 188 2554 192
rect 2635 188 2739 202
rect 2768 204 2818 212
rect 2768 195 2784 204
rect 2475 184 2739 188
rect 2765 192 2784 195
rect 2791 192 2818 204
rect 2765 184 2818 192
rect 2393 176 2394 184
rect 2409 176 2422 184
rect 2393 168 2409 176
rect 2390 161 2409 164
rect 2390 152 2412 161
rect 2363 142 2412 152
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2335 120 2409 136
rect 2427 128 2457 184
rect 2492 174 2700 184
rect 2735 180 2780 184
rect 2783 183 2784 184
rect 2799 183 2812 184
rect 2659 170 2707 174
rect 2542 148 2572 157
rect 2635 150 2650 157
rect 2671 148 2707 170
rect 2518 144 2707 148
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2335 118 2348 120
rect 2363 118 2397 120
rect 2335 102 2409 118
rect 2436 114 2449 128
rect 2464 114 2480 130
rect 2526 125 2537 138
rect 2319 80 2320 96
rect 2335 80 2348 102
rect 2363 80 2393 102
rect 2436 98 2498 114
rect 2526 107 2537 123
rect 2542 118 2552 138
rect 2562 118 2576 138
rect 2579 125 2588 138
rect 2604 125 2613 138
rect 2542 107 2576 118
rect 2579 107 2587 123
rect 2604 107 2613 123
rect 2620 118 2630 138
rect 2640 118 2654 138
rect 2655 125 2666 138
rect 2620 107 2654 118
rect 2655 107 2666 123
rect 2712 114 2728 130
rect 2735 128 2765 180
rect 2799 176 2800 183
rect 2784 168 2800 176
rect 2771 136 2784 155
rect 2799 136 2829 152
rect 2771 120 2845 136
rect 2771 118 2784 120
rect 2799 118 2833 120
rect 2436 96 2449 98
rect 2464 96 2498 98
rect 2436 80 2498 96
rect 2542 91 2555 94
rect 2620 91 2650 102
rect 2698 98 2744 114
rect 2771 102 2845 118
rect 2698 96 2732 98
rect 2697 80 2744 96
rect 2771 80 2784 102
rect 2799 80 2829 102
rect 2856 80 2857 96
rect 2872 80 2885 240
rect 2915 136 2928 240
rect 2973 218 2974 228
rect 2989 218 3002 228
rect 2973 214 3002 218
rect 3007 214 3037 240
rect 3055 226 3071 228
rect 3143 226 3196 240
rect 3144 224 3208 226
rect 3055 214 3070 218
rect 2973 212 3070 214
rect 2957 204 3008 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3039 204 3089 212
rect 3039 196 3055 204
rect 3062 202 3089 204
rect 3098 204 3113 208
rect 3160 204 3192 224
rect 3251 212 3266 240
rect 3315 237 3345 240
rect 3315 234 3351 237
rect 3281 226 3297 228
rect 3282 214 3297 218
rect 3315 215 3354 234
rect 3373 228 3380 229
rect 3379 221 3380 228
rect 3363 218 3364 221
rect 3379 218 3392 221
rect 3315 214 3345 215
rect 3354 214 3360 215
rect 3363 214 3392 218
rect 3282 213 3392 214
rect 3282 212 3398 213
rect 3251 204 3319 212
rect 3098 202 3167 204
rect 3185 202 3319 204
rect 3062 198 3134 202
rect 3062 196 3187 198
rect 3062 192 3134 196
rect 2957 184 3008 192
rect 3055 188 3134 192
rect 3215 188 3319 202
rect 3348 204 3398 212
rect 3348 195 3364 204
rect 3055 184 3319 188
rect 3345 192 3364 195
rect 3371 192 3398 204
rect 3345 184 3398 192
rect 2973 176 2974 184
rect 2989 176 3002 184
rect 2973 168 2989 176
rect 2970 161 2989 164
rect 2970 152 2992 161
rect 2943 142 2992 152
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2915 120 2989 136
rect 3007 128 3037 184
rect 3072 174 3280 184
rect 3315 180 3360 184
rect 3363 183 3364 184
rect 3379 183 3392 184
rect 3239 170 3287 174
rect 3122 148 3152 157
rect 3215 150 3230 157
rect 3251 148 3287 170
rect 3098 144 3287 148
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 2915 118 2928 120
rect 2943 118 2977 120
rect 2915 102 2989 118
rect 3016 114 3029 128
rect 3044 114 3060 130
rect 3106 125 3117 138
rect 2899 80 2900 96
rect 2915 80 2928 102
rect 2943 80 2973 102
rect 3016 98 3078 114
rect 3106 107 3117 123
rect 3122 118 3132 138
rect 3142 118 3156 138
rect 3159 125 3168 138
rect 3184 125 3193 138
rect 3122 107 3156 118
rect 3159 107 3167 123
rect 3184 107 3193 123
rect 3200 118 3210 138
rect 3220 118 3234 138
rect 3235 125 3246 138
rect 3200 107 3234 118
rect 3235 107 3246 123
rect 3292 114 3308 130
rect 3315 128 3345 180
rect 3379 176 3380 183
rect 3364 168 3380 176
rect 3351 136 3364 155
rect 3379 136 3409 152
rect 3351 120 3425 136
rect 3351 118 3364 120
rect 3379 118 3413 120
rect 3016 96 3029 98
rect 3044 96 3078 98
rect 3016 80 3078 96
rect 3122 91 3135 94
rect 3200 91 3230 102
rect 3278 98 3324 114
rect 3351 102 3425 118
rect 3278 96 3312 98
rect 3277 80 3324 96
rect 3351 80 3364 102
rect 3379 80 3409 102
rect 3436 80 3437 96
rect 3452 80 3465 240
rect 3495 136 3508 240
rect 3553 218 3554 228
rect 3569 218 3582 228
rect 3553 214 3582 218
rect 3587 214 3617 240
rect 3635 226 3651 228
rect 3723 226 3776 240
rect 3724 224 3788 226
rect 3635 214 3650 218
rect 3553 212 3650 214
rect 3537 204 3588 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3619 204 3669 212
rect 3619 196 3635 204
rect 3642 202 3669 204
rect 3678 204 3693 208
rect 3740 204 3772 224
rect 3831 212 3846 240
rect 3895 237 3925 240
rect 3895 234 3931 237
rect 3861 226 3877 228
rect 3862 214 3877 218
rect 3895 215 3934 234
rect 3953 228 3960 229
rect 3959 221 3960 228
rect 3943 218 3944 221
rect 3959 218 3972 221
rect 3895 214 3925 215
rect 3934 214 3940 215
rect 3943 214 3972 218
rect 3862 213 3972 214
rect 3862 212 3978 213
rect 3831 204 3899 212
rect 3678 202 3747 204
rect 3765 202 3899 204
rect 3642 198 3714 202
rect 3642 196 3767 198
rect 3642 192 3714 196
rect 3537 184 3588 192
rect 3635 188 3714 192
rect 3795 188 3899 202
rect 3928 204 3978 212
rect 3928 195 3944 204
rect 3635 184 3899 188
rect 3925 192 3944 195
rect 3951 192 3978 204
rect 3925 184 3978 192
rect 3553 176 3554 184
rect 3569 176 3582 184
rect 3553 168 3569 176
rect 3550 161 3569 164
rect 3550 152 3572 161
rect 3523 142 3572 152
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3495 120 3569 136
rect 3587 128 3617 184
rect 3652 174 3860 184
rect 3895 180 3940 184
rect 3943 183 3944 184
rect 3959 183 3972 184
rect 3819 170 3867 174
rect 3702 148 3732 157
rect 3795 150 3810 157
rect 3831 148 3867 170
rect 3678 144 3867 148
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3495 118 3508 120
rect 3523 118 3557 120
rect 3495 102 3569 118
rect 3596 114 3609 128
rect 3624 114 3640 130
rect 3686 125 3697 138
rect 3479 80 3480 96
rect 3495 80 3508 102
rect 3523 80 3553 102
rect 3596 98 3658 114
rect 3686 107 3697 123
rect 3702 118 3712 138
rect 3722 118 3736 138
rect 3739 125 3748 138
rect 3764 125 3773 138
rect 3702 107 3736 118
rect 3739 107 3747 123
rect 3764 107 3773 123
rect 3780 118 3790 138
rect 3800 118 3814 138
rect 3815 125 3826 138
rect 3780 107 3814 118
rect 3815 107 3826 123
rect 3872 114 3888 130
rect 3895 128 3925 180
rect 3959 176 3960 183
rect 3944 168 3960 176
rect 3931 136 3944 155
rect 3959 136 3989 152
rect 3931 120 4005 136
rect 3931 118 3944 120
rect 3959 118 3993 120
rect 3596 96 3609 98
rect 3624 96 3658 98
rect 3596 80 3658 96
rect 3702 91 3715 94
rect 3780 91 3810 102
rect 3858 98 3904 114
rect 3931 102 4005 118
rect 3858 96 3892 98
rect 3857 80 3904 96
rect 3931 80 3944 102
rect 3959 80 3989 102
rect 4016 80 4017 96
rect 4032 80 4045 240
rect 4075 136 4088 240
rect 4133 218 4134 228
rect 4149 218 4162 228
rect 4133 214 4162 218
rect 4167 214 4197 240
rect 4215 226 4231 228
rect 4303 226 4356 240
rect 4304 224 4368 226
rect 4215 214 4230 218
rect 4133 212 4230 214
rect 4117 204 4168 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4199 204 4249 212
rect 4199 196 4215 204
rect 4222 202 4249 204
rect 4258 204 4273 208
rect 4320 204 4352 224
rect 4411 212 4426 240
rect 4475 237 4505 240
rect 4475 234 4511 237
rect 4441 226 4457 228
rect 4442 214 4457 218
rect 4475 215 4514 234
rect 4533 228 4540 229
rect 4539 221 4540 228
rect 4523 218 4524 221
rect 4539 218 4552 221
rect 4475 214 4505 215
rect 4514 214 4520 215
rect 4523 214 4552 218
rect 4442 213 4552 214
rect 4442 212 4558 213
rect 4411 204 4479 212
rect 4258 202 4327 204
rect 4345 202 4479 204
rect 4222 198 4294 202
rect 4222 196 4347 198
rect 4222 192 4294 196
rect 4117 184 4168 192
rect 4215 188 4294 192
rect 4375 188 4479 202
rect 4508 204 4558 212
rect 4508 195 4524 204
rect 4215 184 4479 188
rect 4505 192 4524 195
rect 4531 192 4558 204
rect 4505 184 4558 192
rect 4133 176 4134 184
rect 4149 176 4162 184
rect 4133 168 4149 176
rect 4130 161 4149 164
rect 4130 152 4152 161
rect 4103 142 4152 152
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4075 120 4149 136
rect 4167 128 4197 184
rect 4232 174 4440 184
rect 4475 180 4520 184
rect 4523 183 4524 184
rect 4539 183 4552 184
rect 4399 170 4447 174
rect 4282 148 4312 157
rect 4375 150 4390 157
rect 4411 148 4447 170
rect 4258 144 4447 148
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4075 118 4088 120
rect 4103 118 4137 120
rect 4075 102 4149 118
rect 4176 114 4189 128
rect 4204 114 4220 130
rect 4266 125 4277 138
rect 4059 80 4060 96
rect 4075 80 4088 102
rect 4103 80 4133 102
rect 4176 98 4238 114
rect 4266 107 4277 123
rect 4282 118 4292 138
rect 4302 118 4316 138
rect 4319 125 4328 138
rect 4344 125 4353 138
rect 4282 107 4316 118
rect 4319 107 4327 123
rect 4344 107 4353 123
rect 4360 118 4370 138
rect 4380 118 4394 138
rect 4395 125 4406 138
rect 4360 107 4394 118
rect 4395 107 4406 123
rect 4452 114 4468 130
rect 4475 128 4505 180
rect 4539 176 4540 183
rect 4524 168 4540 176
rect 4511 136 4524 155
rect 4539 136 4569 152
rect 4511 120 4585 136
rect 4511 118 4524 120
rect 4539 118 4573 120
rect 4176 96 4189 98
rect 4204 96 4238 98
rect 4176 80 4238 96
rect 4282 91 4295 94
rect 4360 91 4390 102
rect 4438 98 4484 114
rect 4511 102 4585 118
rect 4438 96 4472 98
rect 4437 80 4484 96
rect 4511 80 4524 102
rect 4539 80 4569 102
rect 4596 80 4597 96
rect 4612 80 4625 240
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 160 80
rect 172 68 247 80
rect 305 68 380 80
rect 392 68 423 80
rect 429 68 464 80
rect 98 66 260 68
rect -7 38 34 46
rect 116 38 129 66
rect 144 64 159 66
rect 183 39 190 46
rect 193 38 260 66
rect 292 66 464 68
rect 262 44 290 48
rect 292 44 372 66
rect 393 64 408 66
rect 262 42 372 44
rect 262 38 290 42
rect 292 38 372 42
rect -1 28 0 38
rect 15 28 28 38
rect 43 28 73 38
rect 116 28 159 38
rect 166 28 174 38
rect 193 30 196 38
rect 260 30 292 38
rect 193 28 359 30
rect 378 28 389 38
rect 393 28 423 38
rect 451 28 464 66
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 740 80
rect 752 68 827 80
rect 885 68 960 80
rect 972 68 1003 80
rect 1009 68 1044 80
rect 678 66 840 68
rect 573 38 614 46
rect 696 38 709 66
rect 724 64 739 66
rect 763 39 770 46
rect 773 38 840 66
rect 872 66 1044 68
rect 842 44 870 48
rect 872 44 952 66
rect 973 64 988 66
rect 842 42 952 44
rect 842 38 870 42
rect 872 38 952 42
rect 479 28 509 38
rect 536 28 537 38
rect 552 28 565 38
rect 579 28 580 38
rect 595 28 608 38
rect 623 28 653 38
rect 696 28 739 38
rect 746 28 754 38
rect 773 30 776 38
rect 840 30 872 38
rect 773 28 939 30
rect 958 28 969 38
rect 973 28 1003 38
rect 1031 28 1044 66
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1320 80
rect 1332 68 1407 80
rect 1465 68 1540 80
rect 1552 68 1583 80
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1153 38 1194 46
rect 1276 38 1289 66
rect 1304 64 1319 66
rect 1343 39 1350 46
rect 1353 38 1420 66
rect 1452 66 1624 68
rect 1422 44 1450 48
rect 1452 44 1532 66
rect 1553 64 1568 66
rect 1422 42 1532 44
rect 1422 38 1450 42
rect 1452 38 1532 42
rect 1059 28 1089 38
rect 1116 28 1117 38
rect 1132 28 1145 38
rect 1159 28 1160 38
rect 1175 28 1188 38
rect 1203 28 1233 38
rect 1276 28 1319 38
rect 1326 28 1334 38
rect 1353 30 1356 38
rect 1420 30 1452 38
rect 1353 28 1519 30
rect 1538 28 1549 38
rect 1553 28 1583 38
rect 1611 28 1624 66
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1900 80
rect 1912 68 1987 80
rect 2045 68 2120 80
rect 2132 68 2163 80
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1733 38 1774 46
rect 1856 38 1869 66
rect 1884 64 1899 66
rect 1923 39 1930 46
rect 1933 38 2000 66
rect 2032 66 2204 68
rect 2002 44 2030 48
rect 2032 44 2112 66
rect 2133 64 2148 66
rect 2002 42 2112 44
rect 2002 38 2030 42
rect 2032 38 2112 42
rect 1639 28 1669 38
rect 1696 28 1697 38
rect 1712 28 1725 38
rect 1739 28 1740 38
rect 1755 28 1768 38
rect 1783 28 1813 38
rect 1856 28 1899 38
rect 1906 28 1914 38
rect 1933 30 1936 38
rect 2000 30 2032 38
rect 1933 28 2099 30
rect 2118 28 2129 38
rect 2133 28 2163 38
rect 2191 28 2204 66
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2480 80
rect 2492 68 2567 80
rect 2625 68 2700 80
rect 2712 68 2743 80
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2313 38 2354 46
rect 2436 38 2449 66
rect 2464 64 2479 66
rect 2503 39 2510 46
rect 2513 38 2580 66
rect 2612 66 2784 68
rect 2582 44 2610 48
rect 2612 44 2692 66
rect 2713 64 2728 66
rect 2582 42 2692 44
rect 2582 38 2610 42
rect 2612 38 2692 42
rect 2219 28 2249 38
rect 2276 28 2277 38
rect 2292 28 2305 38
rect 2319 28 2320 38
rect 2335 28 2348 38
rect 2363 28 2393 38
rect 2436 28 2479 38
rect 2486 28 2494 38
rect 2513 30 2516 38
rect 2580 30 2612 38
rect 2513 28 2679 30
rect 2698 28 2709 38
rect 2713 28 2743 38
rect 2771 28 2784 66
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3060 80
rect 3072 68 3147 80
rect 3205 68 3280 80
rect 3292 68 3323 80
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 2893 38 2934 46
rect 3016 38 3029 66
rect 3044 64 3059 66
rect 3083 39 3090 46
rect 3093 38 3160 66
rect 3192 66 3364 68
rect 3162 44 3190 48
rect 3192 44 3272 66
rect 3293 64 3308 66
rect 3162 42 3272 44
rect 3162 38 3190 42
rect 3192 38 3272 42
rect 2799 28 2829 38
rect 2856 28 2857 38
rect 2872 28 2885 38
rect 2899 28 2900 38
rect 2915 28 2928 38
rect 2943 28 2973 38
rect 3016 28 3059 38
rect 3066 28 3074 38
rect 3093 30 3096 38
rect 3160 30 3192 38
rect 3093 28 3259 30
rect 3278 28 3289 38
rect 3293 28 3323 38
rect 3351 28 3364 66
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3640 80
rect 3652 68 3727 80
rect 3785 68 3860 80
rect 3872 68 3903 80
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3473 38 3514 46
rect 3596 38 3609 66
rect 3624 64 3639 66
rect 3663 39 3670 46
rect 3673 38 3740 66
rect 3772 66 3944 68
rect 3742 44 3770 48
rect 3772 44 3852 66
rect 3873 64 3888 66
rect 3742 42 3852 44
rect 3742 38 3770 42
rect 3772 38 3852 42
rect 3379 28 3409 38
rect 3436 28 3437 38
rect 3452 28 3465 38
rect 3479 28 3480 38
rect 3495 28 3508 38
rect 3523 28 3553 38
rect 3596 28 3639 38
rect 3646 28 3654 38
rect 3673 30 3676 38
rect 3740 30 3772 38
rect 3673 28 3839 30
rect 3858 28 3869 38
rect 3873 28 3903 38
rect 3931 28 3944 66
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4220 80
rect 4232 68 4307 80
rect 4365 68 4440 80
rect 4452 68 4483 80
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4053 38 4094 46
rect 4176 38 4189 66
rect 4204 64 4219 66
rect 4243 39 4250 46
rect 4253 38 4320 66
rect 4352 66 4524 68
rect 4322 44 4350 48
rect 4352 44 4432 66
rect 4453 64 4468 66
rect 4322 42 4432 44
rect 4322 38 4350 42
rect 4352 38 4432 42
rect 3959 28 3989 38
rect 4016 28 4017 38
rect 4032 28 4045 38
rect 4059 28 4060 38
rect 4075 28 4088 38
rect 4103 28 4133 38
rect 4176 28 4219 38
rect 4226 28 4234 38
rect 4253 30 4256 38
rect 4320 30 4352 38
rect 4253 28 4419 30
rect 4438 28 4449 38
rect 4453 28 4483 38
rect 4511 28 4524 66
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4596 38 4631 46
rect 4539 28 4569 38
rect 4596 28 4597 38
rect 4612 28 4625 38
rect -1 22 4625 28
rect 0 14 4625 22
rect 15 0 28 14
rect 43 -4 73 14
rect 116 0 129 14
rect 166 1 174 14
rect 207 1 345 14
rect 378 1 386 14
rect 243 0 294 1
rect 451 0 464 14
rect 244 -2 308 0
rect 479 -4 509 14
rect 552 0 565 14
rect 595 0 608 14
rect 623 -4 653 14
rect 696 0 709 14
rect 746 1 754 14
rect 787 1 925 14
rect 958 1 966 14
rect 823 0 874 1
rect 1031 0 1044 14
rect 824 -2 888 0
rect 1059 -4 1089 14
rect 1132 0 1145 14
rect 1175 0 1188 14
rect 1203 -4 1233 14
rect 1276 0 1289 14
rect 1326 1 1334 14
rect 1367 1 1505 14
rect 1538 1 1546 14
rect 1403 0 1454 1
rect 1611 0 1624 14
rect 1404 -2 1468 0
rect 1639 -4 1669 14
rect 1712 0 1725 14
rect 1755 0 1768 14
rect 1783 -4 1813 14
rect 1856 0 1869 14
rect 1906 1 1914 14
rect 1947 1 2085 14
rect 2118 1 2126 14
rect 1983 0 2034 1
rect 2191 0 2204 14
rect 1984 -2 2048 0
rect 2219 -4 2249 14
rect 2292 0 2305 14
rect 2335 0 2348 14
rect 2363 -4 2393 14
rect 2436 0 2449 14
rect 2486 1 2494 14
rect 2527 1 2665 14
rect 2698 1 2706 14
rect 2563 0 2614 1
rect 2771 0 2784 14
rect 2564 -2 2628 0
rect 2799 -4 2829 14
rect 2872 0 2885 14
rect 2915 0 2928 14
rect 2943 -4 2973 14
rect 3016 0 3029 14
rect 3066 1 3074 14
rect 3107 1 3245 14
rect 3278 1 3286 14
rect 3143 0 3194 1
rect 3351 0 3364 14
rect 3144 -2 3208 0
rect 3379 -4 3409 14
rect 3452 0 3465 14
rect 3495 0 3508 14
rect 3523 -4 3553 14
rect 3596 0 3609 14
rect 3646 1 3654 14
rect 3687 1 3825 14
rect 3858 1 3866 14
rect 3723 0 3774 1
rect 3931 0 3944 14
rect 3724 -2 3788 0
rect 3959 -4 3989 14
rect 4032 0 4045 14
rect 4075 0 4088 14
rect 4103 -4 4133 14
rect 4176 0 4189 14
rect 4226 1 4234 14
rect 4267 1 4405 14
rect 4438 1 4446 14
rect 4303 0 4354 1
rect 4511 0 4524 14
rect 4304 -2 4368 0
rect 4539 -4 4569 14
rect 4612 0 4625 14
<< pwell >>
rect 74 184 89 212
rect 464 184 479 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
<< ndiffc >>
rect 74 184 89 212
rect 464 184 479 213
rect 654 184 669 212
rect 1044 184 1059 213
rect 1234 184 1249 212
rect 1624 184 1639 213
rect 1814 184 1829 212
rect 2204 184 2219 213
rect 2394 184 2409 212
rect 2784 184 2799 213
rect 2974 184 2989 212
rect 3364 184 3379 213
rect 3554 184 3569 212
rect 3944 184 3959 213
rect 4134 184 4149 212
rect 4524 184 4539 213
rect 0 38 15 80
rect 537 38 552 80
rect 580 38 595 80
rect 1117 38 1132 80
rect 1160 38 1175 80
rect 1697 38 1712 80
rect 1740 38 1755 80
rect 2277 38 2292 80
rect 2320 38 2335 80
rect 2857 38 2872 80
rect 2900 38 2915 80
rect 3437 38 3452 80
rect 3480 38 3495 80
rect 4017 38 4032 80
rect 4060 38 4075 80
rect 4597 38 4612 80
<< poly >>
rect 0 8610 30 8640
rect 0 8340 30 8370
rect 0 8070 30 8100
rect 0 7800 30 7830
rect 0 7530 30 7560
rect 0 7260 30 7290
rect 0 6990 30 7020
rect 0 6720 30 6750
rect 0 6450 30 6480
rect 0 6180 30 6210
rect 0 5910 30 5940
rect 0 5640 30 5670
rect 0 5370 30 5400
rect 0 5100 30 5130
rect 0 4830 30 4860
rect 0 4560 30 4590
rect 0 4290 30 4320
rect 0 4020 30 4050
rect 0 3750 30 3780
rect 0 3480 30 3510
rect 0 3210 30 3240
rect 0 2940 30 2970
rect 0 2670 30 2700
rect 0 2400 30 2430
rect 0 2130 30 2160
rect 0 1860 30 1890
rect 0 1590 30 1620
rect 0 1320 30 1350
rect 0 1050 30 1080
rect 0 780 30 810
rect 0 510 30 540
rect 0 240 30 270
<< metal1 >>
rect 0 8596 15 8610
rect 0 8472 15 8506
rect 0 8370 15 8384
rect 0 8326 15 8340
rect 0 8202 15 8236
rect 0 8100 15 8114
rect 0 8056 15 8070
rect 0 7932 15 7966
rect 0 7830 15 7844
rect 0 7786 15 7800
rect 0 7662 15 7696
rect 0 7560 15 7574
rect 0 7516 15 7530
rect 0 7392 15 7426
rect 0 7290 15 7304
rect 0 7246 15 7260
rect 0 7122 15 7156
rect 0 7020 15 7034
rect 0 6976 15 6990
rect 0 6852 15 6886
rect 0 6750 15 6764
rect 0 6706 15 6720
rect 0 6582 15 6616
rect 0 6480 15 6494
rect 0 6436 15 6450
rect 0 6312 15 6346
rect 0 6210 15 6224
rect 0 6166 15 6180
rect 0 6042 15 6076
rect 0 5940 15 5954
rect 0 5896 15 5910
rect 0 5772 15 5806
rect 0 5670 15 5684
rect 0 5626 15 5640
rect 0 5502 15 5536
rect 0 5400 15 5414
rect 0 5356 15 5370
rect 0 5232 15 5266
rect 0 5130 15 5144
rect 0 5086 15 5100
rect 0 4962 15 4996
rect 0 4860 15 4874
rect 0 4816 15 4830
rect 0 4692 15 4726
rect 0 4590 15 4604
rect 0 4546 15 4560
rect 0 4422 15 4456
rect 0 4320 15 4334
rect 0 4276 15 4290
rect 0 4152 15 4186
rect 0 4050 15 4064
rect 0 4006 15 4020
rect 0 3882 15 3916
rect 0 3780 15 3794
rect 0 3736 15 3750
rect 0 3612 15 3646
rect 0 3510 15 3524
rect 0 3466 15 3480
rect 0 3342 15 3376
rect 0 3240 15 3254
rect 0 3196 15 3210
rect 0 3072 15 3106
rect 0 2970 15 2984
rect 0 2926 15 2940
rect 0 2802 15 2836
rect 0 2700 15 2714
rect 0 2656 15 2670
rect 0 2532 15 2566
rect 0 2430 15 2444
rect 0 2386 15 2400
rect 0 2262 15 2296
rect 0 2160 15 2174
rect 0 2116 15 2130
rect 0 1992 15 2026
rect 0 1890 15 1904
rect 0 1846 15 1860
rect 0 1722 15 1756
rect 0 1620 15 1634
rect 0 1576 15 1590
rect 0 1452 15 1486
rect 0 1350 15 1364
rect 0 1306 15 1320
rect 0 1182 15 1216
rect 0 1080 15 1094
rect 0 1036 15 1050
rect 0 912 15 946
rect 0 810 15 824
rect 0 766 15 780
rect 0 642 15 676
rect 0 540 15 554
rect 0 496 15 510
rect 0 372 15 406
rect 0 270 15 284
rect 0 226 15 240
rect 0 102 15 136
rect 0 0 15 14
use 10T_1x8_magic  10T_1x8_magic_16
timestamp 1656019537
transform 1 0 0 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_18
timestamp 1656019537
transform 1 0 0 0 1 270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_19
timestamp 1656019537
transform 1 0 0 0 1 1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_22
timestamp 1656019537
transform 1 0 0 0 1 1350
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_17
timestamp 1656019537
transform 1 0 0 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_20
timestamp 1656019537
transform 1 0 0 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_23
timestamp 1656019537
transform 1 0 0 0 1 2160
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_21
timestamp 1656019537
transform 1 0 0 0 1 1620
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_24
timestamp 1656019537
transform 1 0 0 0 1 1890
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_27
timestamp 1656019537
transform 1 0 0 0 1 3240
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_25
timestamp 1656019537
transform 1 0 0 0 1 2700
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_28
timestamp 1656019537
transform 1 0 0 0 1 2970
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_26
timestamp 1656019537
transform 1 0 0 0 1 2430
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_9
timestamp 1656019537
transform 1 0 0 0 1 4320
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_29
timestamp 1656019537
transform 1 0 0 0 1 3780
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_31
timestamp 1656019537
transform 1 0 0 0 1 4050
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_30
timestamp 1656019537
transform 1 0 0 0 1 3510
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_10
timestamp 1656019537
transform 1 0 0 0 1 4860
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_11
timestamp 1656019537
transform 1 0 0 0 1 5130
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_8
timestamp 1656019537
transform 1 0 0 0 1 4590
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_15
timestamp 1656019537
transform 1 0 0 0 1 5940
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_14
timestamp 1656019537
transform 1 0 0 0 1 6210
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_12
timestamp 1656019537
transform 1 0 0 0 1 5400
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_13
timestamp 1656019537
transform 1 0 0 0 1 5670
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1656019537
transform 1 0 0 0 1 7020
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1656019537
transform 1 0 0 0 1 7290
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1656019537
transform 1 0 0 0 1 6480
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1656019537
transform 1 0 0 0 1 6750
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1656019537
transform 1 0 0 0 1 7560
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1656019537
transform 1 0 0 0 1 7830
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1656019537
transform 1 0 0 0 1 8100
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1656019537
transform 1 0 0 0 1 8370
box -7 -4 4631 312
<< labels >>
rlabel metal1 0 4422 15 4456 1 RWL_15
port 64 ew signal input
rlabel poly 0 4560 30 4590 1 WWL_15
port 63 ew signal input
rlabel metal1 0 4692 15 4726 1 RWL_14
port 62 ew signal input
rlabel poly 0 4830 30 4860 1 WWL_14
port 61 ew signal input
rlabel metal1 0 4962 15 4996 1 RWL_13
port 60 ew signal input
rlabel poly 0 5100 30 5130 1 WWL_13
port 59 ew signal input
rlabel metal1 0 5232 15 5266 1 RWL_12
port 58 ew signal input
rlabel poly 0 5370 30 5400 1 WWL_12
port 57 ew signal input
rlabel metal1 0 5502 15 5536 1 RWL_11
port 56 ew signal input
rlabel poly 0 5640 30 5670 1 WWL_11
port 55 ew signal input
rlabel metal1 0 5772 15 5806 1 RWL_10
port 54 ew signal input
rlabel poly 0 5910 30 5940 1 WWL_10
port 53 ew signal input
rlabel metal1 0 6042 15 6076 1 RWL_9
port 52 ew signal input
rlabel poly 0 6180 30 6210 1 WWL_9
port 51 ew signal input
rlabel metal1 0 6312 15 6346 1 RWL_8
port 50 ew signal input
rlabel poly 0 6450 30 6480 1 WWL_8
port 49 ew signal input
rlabel metal1 0 6436 15 6450 1 VDD
rlabel metal1 0 6210 15 6224 1 GND
rlabel metal1 0 5896 15 5910 1 VDD
rlabel metal1 0 5626 15 5640 1 VDD
rlabel metal1 0 6166 15 6180 1 VDD
rlabel metal1 0 5356 15 5370 1 VDD
rlabel metal1 0 4816 15 4830 1 VDD
rlabel metal1 0 4546 15 4560 1 VDD
rlabel metal1 0 5086 15 5100 1 VDD
rlabel metal1 0 5400 15 5414 1 GND
rlabel metal1 0 5670 15 5684 1 GND
rlabel metal1 0 5940 15 5954 1 GND
rlabel metal1 0 5130 15 5144 1 GND
rlabel metal1 0 4320 15 4334 1 GND
rlabel metal1 0 4590 15 4604 1 GND
rlabel metal1 0 4860 15 4874 1 GND
rlabel poly 0 8610 30 8640 1 WWL_0
port 33 ew signal input
rlabel metal1 0 7020 15 7034 1 GND
rlabel metal1 0 6750 15 6764 1 GND
rlabel metal1 0 6480 15 6494 1 GND
rlabel metal1 0 7290 15 7304 1 GND
rlabel metal1 0 8100 15 8114 1 GND
rlabel metal1 0 7830 15 7844 1 GND
rlabel metal1 0 7560 15 7574 1 GND
rlabel metal1 0 7246 15 7260 1 VDD
rlabel metal1 0 6706 15 6720 1 VDD
rlabel metal1 0 6976 15 6990 1 VDD
rlabel metal1 0 7516 15 7530 1 VDD
rlabel metal1 0 8326 15 8340 1 VDD
rlabel metal1 0 7786 15 7800 1 VDD
rlabel metal1 0 8056 15 8070 1 VDD
rlabel metal1 0 8370 15 8384 1 GND
port 98 ew ground bidirectional abutment
rlabel metal1 0 8596 15 8610 1 VDD
port 97 ew power bidirectional abutment
rlabel metal1 0 6582 15 6616 1 RWL_7
port 48 ew signal input
rlabel poly 0 6720 30 6750 1 WWL_7
port 47 ew signal input
rlabel metal1 0 6852 15 6886 1 RWL_6
port 46 ew signal input
rlabel poly 0 6990 30 7020 1 WWL_6
port 45 ew signal input
rlabel metal1 0 7122 15 7156 1 RWL_5
port 44 ew signal input
rlabel poly 0 7260 30 7290 1 WWL_5
port 43 ew signal input
rlabel metal1 0 7392 15 7426 1 RWL_4
port 42 ew signal input
rlabel poly 0 7530 30 7560 1 WWL_4
port 41 ew signal input
rlabel metal1 0 7662 15 7696 1 RWL_3
port 40 ew signal input
rlabel poly 0 7800 30 7830 1 WWL_3
port 39 ew signal input
rlabel metal1 0 7932 15 7966 1 RWL_2
port 38 ew signal input
rlabel poly 0 8070 30 8100 1 WWL_2
port 37 ew signal input
rlabel metal1 0 8202 15 8236 1 RWL_1
port 36 ew signal input
rlabel poly 0 8340 30 8370 1 WWL_1
port 35 ew signal input
rlabel metal1 0 8472 15 8506 1 RWL_0
port 34 ew signal input
rlabel locali 0 38 15 80 1 RBL1_0
port 1 ns signal output
rlabel locali 537 38 552 80 1 RBL0_0
port 2 ns signal output
rlabel locali 580 38 595 80 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 38 1132 80 1 RBL0_1
port 4 ns signal output
rlabel locali 1160 38 1175 80 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 38 1712 80 1 RBL0_2
port 6 ns signal output
rlabel locali 1740 38 1755 80 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 38 2292 80 1 RBL0_3
port 8 ns signal output
rlabel locali 2320 38 2335 80 1 RBL1_4
port 9 ns signal output
rlabel locali 2857 38 2872 80 1 RBL0_4
port 10 ns signal output
rlabel locali 2900 38 2915 80 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 38 3452 80 1 RBL0_5
port 12 ns signal output
rlabel locali 3480 38 3495 80 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 38 4032 80 1 RBL0_6
port 14 ns signal output
rlabel locali 4060 38 4075 80 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 38 4612 80 1 RBL0_7
port 16 ns signal output
rlabel locali 464 184 479 213 1 WBL_0
port 17 ns signal input
rlabel locali 74 184 89 212 1 WBLb_0
port 18 ns signal input
rlabel locali 1044 184 1059 213 1 WBL_1
port 19 ns signal input
rlabel locali 654 184 669 212 1 WBLb_1
port 20 ns signal input
rlabel locali 1624 184 1639 213 1 WBL_2
port 21 ns signal input
rlabel locali 1234 184 1249 212 1 WBLb_2
port 22 ns signal input
rlabel locali 2204 184 2219 213 1 WBL_3
port 23 ns signal input
rlabel locali 1814 184 1829 212 1 WBLb_3
port 24 ns signal input
rlabel locali 2784 184 2799 213 1 WBL_4
port 25 ns signal input
rlabel locali 2394 184 2409 212 1 WBLb_4
port 26 ns signal input
rlabel locali 3364 184 3379 213 1 WBL_5
port 27 ns signal input
rlabel locali 2974 184 2989 212 1 WBLb_5
port 28 ns signal input
rlabel locali 3944 184 3959 213 1 WBL_6
port 29 ns signal input
rlabel locali 3554 184 3569 212 1 WBLb_6
port 30 ns signal input
rlabel locali 4524 184 4539 213 1 WBL_7
port 31 ns signal input
rlabel locali 4134 184 4149 212 1 WBLb_7
port 32 ns signal input
rlabel metal1 0 2116 15 2130 1 VDD
rlabel metal1 0 1890 15 1904 1 GND
rlabel metal1 0 1576 15 1590 1 VDD
rlabel metal1 0 1306 15 1320 1 VDD
rlabel metal1 0 1846 15 1860 1 VDD
rlabel metal1 0 1036 15 1050 1 VDD
rlabel metal1 0 496 15 510 1 VDD
rlabel metal1 0 226 15 240 1 VDD
rlabel metal1 0 766 15 780 1 VDD
rlabel metal1 0 1080 15 1094 1 GND
rlabel metal1 0 1350 15 1364 1 GND
rlabel metal1 0 1620 15 1634 1 GND
rlabel metal1 0 810 15 824 1 GND
rlabel metal1 0 0 15 14 1 GND
rlabel metal1 0 270 15 284 1 GND
rlabel metal1 0 540 15 554 1 GND
rlabel metal1 0 2700 15 2714 1 GND
rlabel metal1 0 2430 15 2444 1 GND
rlabel metal1 0 2160 15 2174 1 GND
rlabel metal1 0 2970 15 2984 1 GND
rlabel metal1 0 3780 15 3794 1 GND
rlabel metal1 0 3510 15 3524 1 GND
rlabel metal1 0 3240 15 3254 1 GND
rlabel metal1 0 2926 15 2940 1 VDD
rlabel metal1 0 2386 15 2400 1 VDD
rlabel metal1 0 2656 15 2670 1 VDD
rlabel metal1 0 3196 15 3210 1 VDD
rlabel metal1 0 4006 15 4020 1 VDD
rlabel metal1 0 3466 15 3480 1 VDD
rlabel metal1 0 3736 15 3750 1 VDD
rlabel metal1 0 4050 15 4064 1 GND
port 98 ew ground bidirectional abutment
rlabel metal1 0 4276 15 4290 1 VDD
port 97 ew power bidirectional abutment
rlabel poly 0 4290 30 4320 1 WWL_16
port 65 ew signal input
rlabel metal1 0 4152 15 4186 1 RWL_16
port 66 ew signal input
rlabel poly 0 4020 30 4050 1 WWL_17
port 67 ew signal input
rlabel metal1 0 3882 15 3916 1 RWL_17
port 68 ew signal input
rlabel poly 0 3750 30 3780 1 WWL_18
port 69 ew signal input
rlabel metal1 0 3612 15 3646 1 RWL_18
port 70 ew signal input
rlabel poly 0 3480 30 3510 1 WWL_19
port 71 ew signal input
rlabel metal1 0 3342 15 3376 1 RWL_19
port 72 ew signal input
rlabel poly 0 3210 30 3240 1 WWL_20
port 73 ew signal input
rlabel metal1 0 3072 15 3106 1 RWL_20
port 74 ew signal input
rlabel poly 0 2940 30 2970 1 WWL_21
port 75 ew signal input
rlabel metal1 0 2802 15 2836 1 RWL_21
port 76 ew signal input
rlabel poly 0 2670 30 2700 1 WWL_22
port 77 ew signal input
rlabel metal1 0 2532 15 2566 1 RWL_22
port 78 ew signal input
rlabel poly 0 2400 30 2430 1 WWL_23
port 79 ew signal input
rlabel metal1 0 2262 15 2296 1 RWL_23
port 80 ew signal input
rlabel poly 0 2130 30 2160 1 WWL_24
port 81 ew signal input
rlabel metal1 0 1992 15 2026 1 RWL_24
port 82 ew signal input
rlabel poly 0 1860 30 1890 1 WWL_25
port 83 ew signal input
rlabel metal1 0 1722 15 1756 1 RWL_25
port 84 ew signal input
rlabel poly 0 1590 30 1620 1 WWL_26
port 85 ew signal input
rlabel metal1 0 1452 15 1486 1 RWL_26
port 86 ew signal input
rlabel poly 0 1320 30 1350 1 WWL_27
port 87 ew signal input
rlabel metal1 0 1182 15 1216 1 RWL_27
port 88 ew signal input
rlabel poly 0 1050 30 1080 1 WWL_28
port 89 ew signal input
rlabel metal1 0 912 15 946 1 RWL_28
port 90 ew signal input
rlabel poly 0 780 30 810 1 WWL_29
port 91 ew signal input
rlabel metal1 0 642 15 676 1 RWL_29
port 92 ew signal input
rlabel poly 0 510 30 540 1 WWL_30
port 93 ew signal input
rlabel metal1 0 372 15 406 1 RWL_30
port 94 ew signal input
rlabel poly 0 240 30 270 1 WWL_31
port 95 ew signal input
rlabel metal1 0 102 15 136 1 RWL_31
port 96 ew signal input
<< end >>
