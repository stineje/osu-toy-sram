magic
tech sky130
magscale 1 2
timestamp 1668460924
<< error_p >>
rect 14 2158 27 2174
rect 116 2172 129 2174
rect 82 2158 97 2172
rect 106 2158 136 2172
rect 197 2170 350 2216
rect 179 2158 371 2170
rect 414 2158 444 2172
rect 450 2158 463 2174
rect 551 2158 564 2174
rect 594 2158 607 2174
rect 696 2172 709 2174
rect 662 2158 677 2172
rect 686 2158 716 2172
rect 777 2170 930 2216
rect 759 2158 951 2170
rect 994 2158 1024 2172
rect 1030 2158 1043 2174
rect 1131 2158 1144 2174
rect 1174 2158 1187 2174
rect 1276 2172 1281 2174
rect 1242 2158 1257 2172
rect 1266 2158 1281 2172
rect 3494 2158 3507 2174
rect 3596 2172 3609 2174
rect 3562 2158 3577 2172
rect 3586 2158 3616 2172
rect 3677 2170 3830 2216
rect 3659 2158 3851 2170
rect 3894 2158 3924 2172
rect 3930 2158 3943 2174
rect 4031 2158 4044 2174
rect 4074 2158 4087 2174
rect 4176 2172 4189 2174
rect 4142 2158 4157 2172
rect 4166 2158 4196 2172
rect 4257 2170 4410 2216
rect 4239 2158 4431 2170
rect 4474 2158 4504 2172
rect 4510 2158 4523 2174
rect 4611 2158 4624 2174
rect 4654 2158 4667 2174
rect 4756 2172 4769 2174
rect 4722 2158 4737 2172
rect 4746 2158 4776 2172
rect 4837 2170 4990 2216
rect 4819 2158 5011 2170
rect 5054 2158 5084 2172
rect 5090 2158 5103 2174
rect 5191 2158 5204 2174
rect 5234 2158 5247 2174
rect 5336 2172 5349 2174
rect 5302 2158 5317 2172
rect 5326 2158 5356 2172
rect 5417 2170 5570 2216
rect 5399 2158 5591 2170
rect 5634 2158 5664 2172
rect 5670 2158 5683 2174
rect 5771 2158 5784 2174
rect 5814 2158 5827 2174
rect 5916 2172 5929 2174
rect 5882 2158 5897 2172
rect 5906 2158 5936 2172
rect 5997 2170 6150 2216
rect 5979 2158 6171 2170
rect 6214 2158 6244 2172
rect 6250 2158 6263 2174
rect 6351 2158 6364 2174
rect 6394 2158 6407 2174
rect 6496 2172 6509 2174
rect 6462 2158 6477 2172
rect 6486 2158 6516 2172
rect 6577 2170 6730 2216
rect 6559 2158 6751 2170
rect 6794 2158 6824 2172
rect 6830 2158 6843 2174
rect 6931 2158 6944 2174
rect -1 2144 1281 2158
rect 3481 2144 6944 2158
rect 14 2040 27 2144
rect 72 2122 73 2132
rect 88 2122 101 2132
rect 72 2118 101 2122
rect 106 2118 136 2144
rect 154 2130 170 2132
rect 242 2130 295 2144
rect 243 2128 307 2130
rect 350 2128 365 2144
rect 414 2141 444 2144
rect 414 2138 450 2141
rect 380 2130 396 2132
rect 154 2118 169 2122
rect 72 2116 169 2118
rect 197 2116 365 2128
rect 381 2118 396 2122
rect 414 2119 453 2138
rect 472 2132 479 2133
rect 478 2125 479 2132
rect 462 2122 463 2125
rect 478 2122 491 2125
rect 414 2118 444 2119
rect 453 2118 459 2119
rect 462 2118 491 2122
rect 381 2117 491 2118
rect 381 2116 497 2117
rect 56 2108 107 2116
rect 56 2096 81 2108
rect 88 2096 107 2108
rect 138 2108 188 2116
rect 138 2100 154 2108
rect 161 2106 188 2108
rect 197 2106 418 2116
rect 161 2096 418 2106
rect 447 2108 497 2116
rect 447 2099 463 2108
rect 56 2088 107 2096
rect 154 2088 418 2096
rect 444 2096 463 2099
rect 470 2096 497 2108
rect 444 2088 497 2096
rect 72 2080 73 2088
rect 88 2080 101 2088
rect 72 2072 88 2080
rect 69 2065 88 2068
rect 69 2056 91 2065
rect 42 2046 91 2056
rect 42 2040 72 2046
rect 91 2041 96 2046
rect 14 2024 88 2040
rect 106 2032 136 2088
rect 171 2078 379 2088
rect 414 2084 459 2088
rect 462 2087 463 2088
rect 478 2087 491 2088
rect 197 2048 386 2078
rect 212 2045 386 2048
rect 205 2042 386 2045
rect 14 2022 27 2024
rect 42 2022 76 2024
rect 14 2006 88 2022
rect 115 2018 128 2032
rect 143 2018 159 2034
rect 205 2029 216 2042
rect -2 1984 -1 2000
rect 14 1984 27 2006
rect 42 1984 72 2006
rect 115 2002 177 2018
rect 205 2011 216 2027
rect 221 2022 231 2042
rect 241 2022 255 2042
rect 258 2029 267 2042
rect 283 2029 292 2042
rect 221 2011 255 2022
rect 258 2011 267 2027
rect 283 2011 292 2027
rect 299 2022 309 2042
rect 319 2022 333 2042
rect 334 2029 345 2042
rect 299 2011 333 2022
rect 334 2011 345 2027
rect 391 2018 407 2034
rect 414 2032 444 2084
rect 478 2080 479 2087
rect 463 2072 479 2080
rect 450 2040 463 2059
rect 478 2040 508 2056
rect 450 2024 524 2040
rect 450 2022 463 2024
rect 478 2022 512 2024
rect 115 2000 128 2002
rect 143 2000 177 2002
rect 115 1984 177 2000
rect 221 1995 237 2002
rect 299 1995 329 2006
rect 377 2002 423 2018
rect 450 2006 524 2022
rect 377 2000 411 2002
rect 376 1984 423 2000
rect 450 1984 463 2006
rect 478 1984 508 2006
rect 535 1984 536 2000
rect 551 1984 564 2144
rect 594 2040 607 2144
rect 652 2122 653 2132
rect 668 2122 681 2132
rect 652 2118 681 2122
rect 686 2118 716 2144
rect 734 2130 750 2132
rect 822 2130 875 2144
rect 823 2128 887 2130
rect 930 2128 945 2144
rect 994 2141 1024 2144
rect 994 2138 1030 2141
rect 960 2130 976 2132
rect 734 2118 749 2122
rect 652 2116 749 2118
rect 777 2116 945 2128
rect 961 2118 976 2122
rect 994 2119 1033 2138
rect 1052 2132 1059 2133
rect 1058 2125 1059 2132
rect 1042 2122 1043 2125
rect 1058 2122 1071 2125
rect 994 2118 1024 2119
rect 1033 2118 1039 2119
rect 1042 2118 1071 2122
rect 961 2117 1071 2118
rect 961 2116 1077 2117
rect 636 2108 687 2116
rect 636 2096 661 2108
rect 668 2096 687 2108
rect 718 2108 768 2116
rect 718 2100 734 2108
rect 741 2106 768 2108
rect 777 2106 998 2116
rect 741 2096 998 2106
rect 1027 2108 1077 2116
rect 1027 2099 1043 2108
rect 636 2088 687 2096
rect 734 2088 998 2096
rect 1024 2096 1043 2099
rect 1050 2096 1077 2108
rect 1024 2088 1077 2096
rect 652 2080 653 2088
rect 668 2080 681 2088
rect 652 2072 668 2080
rect 649 2065 668 2068
rect 649 2056 671 2065
rect 622 2046 671 2056
rect 622 2040 652 2046
rect 671 2041 676 2046
rect 594 2024 668 2040
rect 686 2032 716 2088
rect 751 2078 959 2088
rect 994 2084 1039 2088
rect 1042 2087 1043 2088
rect 1058 2087 1071 2088
rect 777 2048 966 2078
rect 792 2045 966 2048
rect 785 2042 966 2045
rect 594 2022 607 2024
rect 622 2022 656 2024
rect 594 2006 668 2022
rect 695 2018 708 2032
rect 723 2018 739 2034
rect 785 2029 796 2042
rect 578 1984 579 2000
rect 594 1984 607 2006
rect 622 1984 652 2006
rect 695 2002 757 2018
rect 785 2011 796 2027
rect 801 2022 811 2042
rect 821 2022 835 2042
rect 838 2029 847 2042
rect 863 2029 872 2042
rect 801 2011 835 2022
rect 838 2011 847 2027
rect 863 2011 872 2027
rect 879 2022 889 2042
rect 899 2022 913 2042
rect 914 2029 925 2042
rect 879 2011 913 2022
rect 914 2011 925 2027
rect 971 2018 987 2034
rect 994 2032 1024 2084
rect 1058 2080 1059 2087
rect 1043 2072 1059 2080
rect 1030 2040 1043 2059
rect 1058 2040 1088 2056
rect 1030 2024 1104 2040
rect 1030 2022 1043 2024
rect 1058 2022 1092 2024
rect 695 2000 708 2002
rect 723 2000 757 2002
rect 695 1984 757 2000
rect 801 1995 817 2002
rect 879 1995 909 2006
rect 957 2002 1003 2018
rect 1030 2006 1104 2022
rect 957 2000 991 2002
rect 956 1984 1003 2000
rect 1030 1984 1043 2006
rect 1058 1984 1088 2006
rect 1115 1984 1116 2000
rect 1131 1984 1144 2144
rect 1174 2040 1187 2144
rect 1232 2122 1233 2132
rect 1248 2122 1261 2132
rect 1232 2118 1261 2122
rect 1266 2118 1281 2144
rect 1232 2116 1281 2118
rect 1216 2108 1267 2116
rect 1216 2096 1241 2108
rect 1248 2096 1267 2108
rect 1216 2088 1267 2096
rect 1232 2080 1233 2088
rect 1248 2080 1261 2088
rect 1232 2072 1248 2080
rect 1229 2065 1248 2068
rect 1229 2056 1251 2065
rect 1202 2046 1251 2056
rect 1202 2040 1232 2046
rect 1251 2041 1256 2046
rect 1174 2024 1248 2040
rect 1266 2032 1281 2088
rect 1174 2022 1187 2024
rect 1202 2022 1236 2024
rect 1174 2006 1248 2022
rect 1158 1984 1159 2000
rect 1174 1984 1187 2006
rect 1202 1984 1232 2006
rect 1275 1984 1281 2032
rect 3494 2040 3507 2144
rect 3552 2122 3553 2132
rect 3568 2122 3581 2132
rect 3552 2118 3581 2122
rect 3586 2118 3616 2144
rect 3634 2130 3650 2132
rect 3722 2130 3775 2144
rect 3723 2128 3787 2130
rect 3830 2128 3845 2144
rect 3894 2141 3924 2144
rect 3894 2138 3930 2141
rect 3860 2130 3876 2132
rect 3634 2118 3649 2122
rect 3552 2116 3649 2118
rect 3677 2116 3845 2128
rect 3861 2118 3876 2122
rect 3894 2119 3933 2138
rect 3952 2132 3959 2133
rect 3958 2125 3959 2132
rect 3942 2122 3943 2125
rect 3958 2122 3971 2125
rect 3894 2118 3924 2119
rect 3933 2118 3939 2119
rect 3942 2118 3971 2122
rect 3861 2117 3971 2118
rect 3861 2116 3977 2117
rect 3536 2108 3587 2116
rect 3536 2096 3561 2108
rect 3568 2096 3587 2108
rect 3618 2108 3668 2116
rect 3618 2100 3634 2108
rect 3641 2106 3668 2108
rect 3677 2106 3898 2116
rect 3641 2096 3898 2106
rect 3927 2108 3977 2116
rect 3927 2099 3943 2108
rect 3536 2088 3587 2096
rect 3634 2088 3898 2096
rect 3924 2096 3943 2099
rect 3950 2096 3977 2108
rect 3924 2088 3977 2096
rect 3552 2080 3553 2088
rect 3568 2080 3581 2088
rect 3552 2072 3568 2080
rect 3549 2065 3568 2068
rect 3549 2056 3571 2065
rect 3522 2046 3571 2056
rect 3522 2040 3552 2046
rect 3571 2041 3576 2046
rect 3494 2024 3568 2040
rect 3586 2032 3616 2088
rect 3651 2078 3859 2088
rect 3894 2084 3939 2088
rect 3942 2087 3943 2088
rect 3958 2087 3971 2088
rect 3677 2048 3866 2078
rect 3692 2045 3866 2048
rect 3685 2042 3866 2045
rect 3494 2022 3507 2024
rect 3522 2022 3556 2024
rect 3494 2006 3568 2022
rect 3595 2018 3608 2032
rect 3623 2018 3639 2034
rect 3685 2029 3696 2042
rect 3494 1984 3507 2006
rect 3522 1984 3552 2006
rect 3595 2002 3657 2018
rect 3685 2011 3696 2027
rect 3701 2022 3711 2042
rect 3721 2022 3735 2042
rect 3738 2029 3747 2042
rect 3763 2029 3772 2042
rect 3701 2011 3735 2022
rect 3738 2011 3747 2027
rect 3763 2011 3772 2027
rect 3779 2022 3789 2042
rect 3799 2022 3813 2042
rect 3814 2029 3825 2042
rect 3779 2011 3813 2022
rect 3814 2011 3825 2027
rect 3871 2018 3887 2034
rect 3894 2032 3924 2084
rect 3958 2080 3959 2087
rect 3943 2072 3959 2080
rect 3930 2040 3943 2059
rect 3958 2040 3988 2056
rect 3930 2024 4004 2040
rect 3930 2022 3943 2024
rect 3958 2022 3992 2024
rect 3595 2000 3608 2002
rect 3623 2000 3657 2002
rect 3595 1984 3657 2000
rect 3701 1995 3717 2002
rect 3779 1995 3809 2006
rect 3857 2002 3903 2018
rect 3930 2006 4004 2022
rect 3857 2000 3891 2002
rect 3856 1984 3903 2000
rect 3930 1984 3943 2006
rect 3958 1984 3988 2006
rect 4015 1984 4016 2000
rect 4031 1984 4044 2144
rect 4074 2040 4087 2144
rect 4132 2122 4133 2132
rect 4148 2122 4161 2132
rect 4132 2118 4161 2122
rect 4166 2118 4196 2144
rect 4214 2130 4230 2132
rect 4302 2130 4355 2144
rect 4303 2128 4367 2130
rect 4410 2128 4425 2144
rect 4474 2141 4504 2144
rect 4474 2138 4510 2141
rect 4440 2130 4456 2132
rect 4214 2118 4229 2122
rect 4132 2116 4229 2118
rect 4257 2116 4425 2128
rect 4441 2118 4456 2122
rect 4474 2119 4513 2138
rect 4532 2132 4539 2133
rect 4538 2125 4539 2132
rect 4522 2122 4523 2125
rect 4538 2122 4551 2125
rect 4474 2118 4504 2119
rect 4513 2118 4519 2119
rect 4522 2118 4551 2122
rect 4441 2117 4551 2118
rect 4441 2116 4557 2117
rect 4116 2108 4167 2116
rect 4116 2096 4141 2108
rect 4148 2096 4167 2108
rect 4198 2108 4248 2116
rect 4198 2100 4214 2108
rect 4221 2106 4248 2108
rect 4257 2106 4478 2116
rect 4221 2096 4478 2106
rect 4507 2108 4557 2116
rect 4507 2099 4523 2108
rect 4116 2088 4167 2096
rect 4214 2088 4478 2096
rect 4504 2096 4523 2099
rect 4530 2096 4557 2108
rect 4504 2088 4557 2096
rect 4132 2080 4133 2088
rect 4148 2080 4161 2088
rect 4132 2072 4148 2080
rect 4129 2065 4148 2068
rect 4129 2056 4151 2065
rect 4102 2046 4151 2056
rect 4102 2040 4132 2046
rect 4151 2041 4156 2046
rect 4074 2024 4148 2040
rect 4166 2032 4196 2088
rect 4231 2078 4439 2088
rect 4474 2084 4519 2088
rect 4522 2087 4523 2088
rect 4538 2087 4551 2088
rect 4257 2048 4446 2078
rect 4272 2045 4446 2048
rect 4265 2042 4446 2045
rect 4074 2022 4087 2024
rect 4102 2022 4136 2024
rect 4074 2006 4148 2022
rect 4175 2018 4188 2032
rect 4203 2018 4219 2034
rect 4265 2029 4276 2042
rect 4058 1984 4059 2000
rect 4074 1984 4087 2006
rect 4102 1984 4132 2006
rect 4175 2002 4237 2018
rect 4265 2011 4276 2027
rect 4281 2022 4291 2042
rect 4301 2022 4315 2042
rect 4318 2029 4327 2042
rect 4343 2029 4352 2042
rect 4281 2011 4315 2022
rect 4318 2011 4327 2027
rect 4343 2011 4352 2027
rect 4359 2022 4369 2042
rect 4379 2022 4393 2042
rect 4394 2029 4405 2042
rect 4359 2011 4393 2022
rect 4394 2011 4405 2027
rect 4451 2018 4467 2034
rect 4474 2032 4504 2084
rect 4538 2080 4539 2087
rect 4523 2072 4539 2080
rect 4510 2040 4523 2059
rect 4538 2040 4568 2056
rect 4510 2024 4584 2040
rect 4510 2022 4523 2024
rect 4538 2022 4572 2024
rect 4175 2000 4188 2002
rect 4203 2000 4237 2002
rect 4175 1984 4237 2000
rect 4281 1995 4297 2002
rect 4359 1995 4389 2006
rect 4437 2002 4483 2018
rect 4510 2006 4584 2022
rect 4437 2000 4471 2002
rect 4436 1984 4483 2000
rect 4510 1984 4523 2006
rect 4538 1984 4568 2006
rect 4595 1984 4596 2000
rect 4611 1984 4624 2144
rect 4654 2040 4667 2144
rect 4712 2122 4713 2132
rect 4728 2122 4741 2132
rect 4712 2118 4741 2122
rect 4746 2118 4776 2144
rect 4794 2130 4810 2132
rect 4882 2130 4933 2144
rect 4883 2128 4947 2130
rect 4990 2128 5005 2144
rect 5054 2141 5084 2144
rect 5054 2138 5090 2141
rect 5020 2130 5036 2132
rect 4794 2118 4809 2122
rect 4712 2116 4809 2118
rect 4837 2116 5005 2128
rect 5021 2118 5036 2122
rect 5054 2119 5093 2138
rect 5112 2132 5119 2133
rect 5118 2125 5119 2132
rect 5102 2122 5103 2125
rect 5118 2122 5131 2125
rect 5054 2118 5084 2119
rect 5093 2118 5099 2119
rect 5102 2118 5131 2122
rect 5021 2117 5131 2118
rect 5021 2116 5137 2117
rect 4696 2108 4747 2116
rect 4696 2096 4721 2108
rect 4728 2096 4747 2108
rect 4778 2108 4828 2116
rect 4778 2100 4794 2108
rect 4801 2106 4828 2108
rect 4837 2106 5058 2116
rect 4801 2096 5058 2106
rect 5087 2108 5137 2116
rect 5087 2099 5103 2108
rect 4696 2088 4747 2096
rect 4794 2088 5058 2096
rect 5084 2096 5103 2099
rect 5110 2096 5137 2108
rect 5084 2088 5137 2096
rect 4712 2080 4713 2088
rect 4728 2080 4741 2088
rect 4712 2072 4728 2080
rect 4709 2065 4728 2068
rect 4709 2056 4731 2065
rect 4682 2046 4731 2056
rect 4682 2040 4712 2046
rect 4731 2041 4736 2046
rect 4654 2024 4728 2040
rect 4746 2032 4776 2088
rect 4811 2078 5019 2088
rect 5054 2084 5099 2088
rect 5102 2087 5103 2088
rect 5118 2087 5131 2088
rect 4837 2048 5026 2078
rect 4852 2045 5026 2048
rect 4845 2042 5026 2045
rect 4654 2022 4667 2024
rect 4682 2022 4716 2024
rect 4654 2006 4728 2022
rect 4755 2018 4768 2032
rect 4783 2018 4799 2034
rect 4845 2029 4856 2042
rect 4638 1984 4639 2000
rect 4654 1984 4667 2006
rect 4682 1984 4712 2006
rect 4755 2002 4817 2018
rect 4845 2011 4856 2027
rect 4861 2022 4871 2042
rect 4881 2022 4895 2042
rect 4898 2029 4907 2042
rect 4923 2029 4932 2042
rect 4861 2011 4895 2022
rect 4898 2011 4907 2027
rect 4923 2011 4932 2027
rect 4939 2022 4949 2042
rect 4959 2022 4973 2042
rect 4974 2029 4985 2042
rect 4939 2011 4973 2022
rect 4974 2011 4985 2027
rect 5031 2018 5047 2034
rect 5054 2032 5084 2084
rect 5118 2080 5119 2087
rect 5103 2072 5119 2080
rect 5090 2040 5103 2059
rect 5118 2040 5148 2056
rect 5090 2024 5164 2040
rect 5090 2022 5103 2024
rect 5118 2022 5152 2024
rect 4755 2000 4768 2002
rect 4783 2000 4817 2002
rect 4755 1984 4817 2000
rect 4861 1995 4877 2002
rect 4939 1995 4969 2006
rect 5017 2002 5063 2018
rect 5090 2006 5164 2022
rect 5017 2000 5051 2002
rect 5016 1984 5063 2000
rect 5090 1984 5103 2006
rect 5118 1984 5148 2006
rect 5175 1984 5176 2000
rect 5191 1984 5204 2144
rect 5234 2040 5247 2144
rect 5292 2122 5293 2132
rect 5308 2122 5321 2132
rect 5292 2118 5321 2122
rect 5326 2118 5356 2144
rect 5374 2130 5390 2132
rect 5462 2130 5513 2144
rect 5463 2128 5527 2130
rect 5570 2128 5585 2144
rect 5634 2141 5664 2144
rect 5634 2138 5670 2141
rect 5600 2130 5616 2132
rect 5374 2118 5389 2122
rect 5292 2116 5389 2118
rect 5417 2116 5585 2128
rect 5601 2118 5616 2122
rect 5634 2119 5673 2138
rect 5692 2132 5699 2133
rect 5698 2125 5699 2132
rect 5682 2122 5683 2125
rect 5698 2122 5711 2125
rect 5634 2118 5664 2119
rect 5673 2118 5679 2119
rect 5682 2118 5711 2122
rect 5601 2117 5711 2118
rect 5601 2116 5717 2117
rect 5276 2108 5327 2116
rect 5276 2096 5301 2108
rect 5308 2096 5327 2108
rect 5358 2108 5408 2116
rect 5358 2100 5374 2108
rect 5381 2106 5408 2108
rect 5417 2106 5638 2116
rect 5381 2096 5638 2106
rect 5667 2108 5717 2116
rect 5667 2099 5683 2108
rect 5276 2088 5327 2096
rect 5374 2088 5638 2096
rect 5664 2096 5683 2099
rect 5690 2096 5717 2108
rect 5664 2088 5717 2096
rect 5292 2080 5293 2088
rect 5308 2080 5321 2088
rect 5292 2072 5308 2080
rect 5289 2065 5308 2068
rect 5289 2056 5311 2065
rect 5262 2046 5311 2056
rect 5262 2040 5292 2046
rect 5311 2041 5316 2046
rect 5234 2024 5308 2040
rect 5326 2032 5356 2088
rect 5391 2078 5599 2088
rect 5634 2084 5679 2088
rect 5682 2087 5683 2088
rect 5698 2087 5711 2088
rect 5417 2048 5606 2078
rect 5432 2045 5606 2048
rect 5425 2042 5606 2045
rect 5234 2022 5247 2024
rect 5262 2022 5296 2024
rect 5234 2006 5308 2022
rect 5335 2018 5348 2032
rect 5363 2018 5379 2034
rect 5425 2029 5436 2042
rect 5218 1984 5219 2000
rect 5234 1984 5247 2006
rect 5262 1984 5292 2006
rect 5335 2002 5397 2018
rect 5425 2011 5436 2027
rect 5441 2022 5451 2042
rect 5461 2022 5475 2042
rect 5478 2029 5487 2042
rect 5503 2029 5512 2042
rect 5441 2011 5475 2022
rect 5478 2011 5487 2027
rect 5503 2011 5512 2027
rect 5519 2022 5529 2042
rect 5539 2022 5553 2042
rect 5554 2029 5565 2042
rect 5519 2011 5553 2022
rect 5554 2011 5565 2027
rect 5611 2018 5627 2034
rect 5634 2032 5664 2084
rect 5698 2080 5699 2087
rect 5683 2072 5699 2080
rect 5670 2040 5683 2059
rect 5698 2040 5728 2056
rect 5670 2024 5744 2040
rect 5670 2022 5683 2024
rect 5698 2022 5732 2024
rect 5335 2000 5348 2002
rect 5363 2000 5397 2002
rect 5335 1984 5397 2000
rect 5441 1995 5457 2002
rect 5519 1995 5549 2006
rect 5597 2002 5643 2018
rect 5670 2006 5744 2022
rect 5597 2000 5631 2002
rect 5596 1984 5643 2000
rect 5670 1984 5683 2006
rect 5698 1984 5728 2006
rect 5755 1984 5756 2000
rect 5771 1984 5784 2144
rect 5814 2040 5827 2144
rect 5872 2122 5873 2132
rect 5888 2122 5901 2132
rect 5872 2118 5901 2122
rect 5906 2118 5936 2144
rect 5954 2130 5970 2132
rect 6042 2130 6093 2144
rect 6043 2128 6107 2130
rect 6150 2128 6165 2144
rect 6214 2141 6244 2144
rect 6214 2138 6250 2141
rect 6180 2130 6196 2132
rect 5954 2118 5969 2122
rect 5872 2116 5969 2118
rect 5997 2116 6165 2128
rect 6181 2118 6196 2122
rect 6214 2119 6253 2138
rect 6272 2132 6279 2133
rect 6278 2125 6279 2132
rect 6262 2122 6263 2125
rect 6278 2122 6291 2125
rect 6214 2118 6244 2119
rect 6253 2118 6259 2119
rect 6262 2118 6291 2122
rect 6181 2117 6291 2118
rect 6181 2116 6297 2117
rect 5856 2108 5907 2116
rect 5856 2096 5881 2108
rect 5888 2096 5907 2108
rect 5938 2108 5988 2116
rect 5938 2100 5954 2108
rect 5961 2106 5988 2108
rect 5997 2106 6218 2116
rect 5961 2096 6218 2106
rect 6247 2108 6297 2116
rect 6247 2099 6263 2108
rect 5856 2088 5907 2096
rect 5954 2088 6218 2096
rect 6244 2096 6263 2099
rect 6270 2096 6297 2108
rect 6244 2088 6297 2096
rect 5872 2080 5873 2088
rect 5888 2080 5901 2088
rect 5872 2072 5888 2080
rect 5869 2065 5888 2068
rect 5869 2056 5891 2065
rect 5842 2046 5891 2056
rect 5842 2040 5872 2046
rect 5891 2041 5896 2046
rect 5814 2024 5888 2040
rect 5906 2032 5936 2088
rect 5971 2078 6179 2088
rect 6214 2084 6259 2088
rect 6262 2087 6263 2088
rect 6278 2087 6291 2088
rect 5997 2048 6186 2078
rect 6012 2045 6186 2048
rect 6005 2042 6186 2045
rect 5814 2022 5827 2024
rect 5842 2022 5876 2024
rect 5814 2006 5888 2022
rect 5915 2018 5928 2032
rect 5943 2018 5959 2034
rect 6005 2029 6016 2042
rect 5798 1984 5799 2000
rect 5814 1984 5827 2006
rect 5842 1984 5872 2006
rect 5915 2002 5977 2018
rect 6005 2011 6016 2027
rect 6021 2022 6031 2042
rect 6041 2022 6055 2042
rect 6058 2029 6067 2042
rect 6083 2029 6092 2042
rect 6021 2011 6055 2022
rect 6058 2011 6067 2027
rect 6083 2011 6092 2027
rect 6099 2022 6109 2042
rect 6119 2022 6133 2042
rect 6134 2029 6145 2042
rect 6099 2011 6133 2022
rect 6134 2011 6145 2027
rect 6191 2018 6207 2034
rect 6214 2032 6244 2084
rect 6278 2080 6279 2087
rect 6263 2072 6279 2080
rect 6250 2040 6263 2059
rect 6278 2040 6308 2056
rect 6250 2024 6324 2040
rect 6250 2022 6263 2024
rect 6278 2022 6312 2024
rect 5915 2000 5928 2002
rect 5943 2000 5977 2002
rect 5915 1984 5977 2000
rect 6021 1995 6037 2002
rect 6099 1995 6129 2006
rect 6177 2002 6223 2018
rect 6250 2006 6324 2022
rect 6177 2000 6211 2002
rect 6176 1984 6223 2000
rect 6250 1984 6263 2006
rect 6278 1984 6308 2006
rect 6335 1984 6336 2000
rect 6351 1984 6364 2144
rect 6394 2040 6407 2144
rect 6452 2122 6453 2132
rect 6468 2122 6481 2132
rect 6452 2118 6481 2122
rect 6486 2118 6516 2144
rect 6534 2130 6550 2132
rect 6622 2130 6673 2144
rect 6623 2128 6687 2130
rect 6730 2128 6745 2144
rect 6794 2141 6824 2144
rect 6794 2138 6830 2141
rect 6760 2130 6776 2132
rect 6534 2118 6549 2122
rect 6452 2116 6549 2118
rect 6577 2116 6745 2128
rect 6761 2118 6776 2122
rect 6794 2119 6833 2138
rect 6852 2132 6859 2133
rect 6858 2125 6859 2132
rect 6842 2122 6843 2125
rect 6858 2122 6871 2125
rect 6794 2118 6824 2119
rect 6833 2118 6839 2119
rect 6842 2118 6871 2122
rect 6761 2117 6871 2118
rect 6761 2116 6877 2117
rect 6436 2108 6487 2116
rect 6436 2096 6461 2108
rect 6468 2096 6487 2108
rect 6518 2108 6568 2116
rect 6518 2100 6534 2108
rect 6541 2106 6568 2108
rect 6577 2106 6798 2116
rect 6541 2096 6798 2106
rect 6827 2108 6877 2116
rect 6827 2099 6843 2108
rect 6436 2088 6487 2096
rect 6534 2088 6798 2096
rect 6824 2096 6843 2099
rect 6850 2096 6877 2108
rect 6824 2088 6877 2096
rect 6452 2080 6453 2088
rect 6468 2080 6481 2088
rect 6452 2072 6468 2080
rect 6449 2065 6468 2068
rect 6449 2056 6471 2065
rect 6422 2046 6471 2056
rect 6422 2040 6452 2046
rect 6471 2041 6476 2046
rect 6394 2024 6468 2040
rect 6486 2032 6516 2088
rect 6551 2078 6759 2088
rect 6794 2084 6839 2088
rect 6842 2087 6843 2088
rect 6858 2087 6871 2088
rect 6577 2048 6766 2078
rect 6592 2045 6766 2048
rect 6585 2042 6766 2045
rect 6394 2022 6407 2024
rect 6422 2022 6456 2024
rect 6394 2006 6468 2022
rect 6495 2018 6508 2032
rect 6523 2018 6539 2034
rect 6585 2029 6596 2042
rect 6378 1984 6379 2000
rect 6394 1984 6407 2006
rect 6422 1984 6452 2006
rect 6495 2002 6557 2018
rect 6585 2011 6596 2027
rect 6601 2022 6611 2042
rect 6621 2022 6635 2042
rect 6638 2029 6647 2042
rect 6663 2029 6672 2042
rect 6601 2011 6635 2022
rect 6638 2011 6647 2027
rect 6663 2011 6672 2027
rect 6679 2022 6689 2042
rect 6699 2022 6713 2042
rect 6714 2029 6725 2042
rect 6679 2011 6713 2022
rect 6714 2011 6725 2027
rect 6771 2018 6787 2034
rect 6794 2032 6824 2084
rect 6858 2080 6859 2087
rect 6843 2072 6859 2080
rect 6830 2040 6843 2059
rect 6858 2040 6888 2056
rect 6830 2024 6904 2040
rect 6830 2022 6843 2024
rect 6858 2022 6892 2024
rect 6495 2000 6508 2002
rect 6523 2000 6557 2002
rect 6495 1984 6557 2000
rect 6601 1995 6617 2002
rect 6679 1995 6709 2006
rect 6757 2002 6803 2018
rect 6830 2006 6904 2022
rect 6757 2000 6791 2002
rect 6756 1984 6803 2000
rect 6830 1984 6843 2006
rect 6858 1984 6888 2006
rect 6915 1984 6916 2000
rect 6931 1984 6944 2144
rect -8 1976 33 1984
rect -8 1950 7 1976
rect 14 1950 33 1976
rect 97 1972 159 1984
rect 171 1972 246 1984
rect 304 1972 379 1984
rect 391 1972 422 1984
rect 428 1972 463 1984
rect 97 1970 259 1972
rect -8 1942 33 1950
rect 115 1946 128 1970
rect 143 1968 158 1970
rect -2 1932 -1 1942
rect 14 1932 27 1942
rect 42 1932 72 1946
rect 115 1932 158 1946
rect 182 1943 189 1950
rect 192 1946 259 1970
rect 291 1970 463 1972
rect 261 1948 289 1952
rect 291 1948 371 1970
rect 392 1968 407 1970
rect 261 1946 371 1948
rect 192 1942 371 1946
rect 165 1932 195 1942
rect 197 1932 350 1942
rect 358 1932 388 1942
rect 392 1932 422 1946
rect 450 1932 463 1970
rect 535 1976 570 1984
rect 535 1950 536 1976
rect 543 1950 570 1976
rect 478 1932 508 1946
rect 535 1942 570 1950
rect 572 1976 613 1984
rect 572 1950 587 1976
rect 594 1950 613 1976
rect 677 1972 739 1984
rect 751 1972 826 1984
rect 884 1972 959 1984
rect 971 1972 1002 1984
rect 1008 1972 1043 1984
rect 677 1970 839 1972
rect 572 1942 613 1950
rect 695 1946 708 1970
rect 723 1968 738 1970
rect 535 1932 536 1942
rect 551 1932 564 1942
rect 578 1932 579 1942
rect 594 1932 607 1942
rect 622 1932 652 1946
rect 695 1932 738 1946
rect 762 1943 769 1950
rect 772 1946 839 1970
rect 871 1970 1043 1972
rect 841 1948 869 1952
rect 871 1948 951 1970
rect 972 1968 987 1970
rect 841 1946 951 1948
rect 772 1942 951 1946
rect 745 1932 775 1942
rect 777 1932 930 1942
rect 938 1932 968 1942
rect 972 1932 1002 1946
rect 1030 1932 1043 1970
rect 1115 1976 1150 1984
rect 1115 1950 1116 1976
rect 1123 1950 1150 1976
rect 1058 1932 1088 1946
rect 1115 1942 1150 1950
rect 1152 1976 1193 1984
rect 1152 1950 1167 1976
rect 1174 1950 1193 1976
rect 1257 1970 1281 1984
rect 1152 1942 1193 1950
rect 1115 1932 1116 1942
rect 1131 1932 1144 1942
rect 1158 1932 1159 1942
rect 1174 1932 1187 1942
rect 1202 1932 1232 1946
rect 1275 1932 1281 1970
rect 3481 1976 3513 1984
rect 3481 1950 3487 1976
rect 3494 1950 3513 1976
rect 3577 1972 3639 1984
rect 3651 1972 3726 1984
rect 3784 1972 3859 1984
rect 3871 1972 3902 1984
rect 3908 1972 3943 1984
rect 3577 1970 3739 1972
rect 3481 1942 3513 1950
rect 3595 1946 3608 1970
rect 3623 1968 3638 1970
rect 3494 1932 3507 1942
rect 3522 1932 3552 1946
rect 3595 1932 3638 1946
rect 3662 1943 3669 1950
rect 3672 1946 3739 1970
rect 3771 1970 3943 1972
rect 3741 1948 3769 1952
rect 3771 1948 3851 1970
rect 3872 1968 3887 1970
rect 3741 1946 3851 1948
rect 3672 1942 3851 1946
rect 3645 1932 3675 1942
rect 3677 1932 3830 1942
rect 3838 1932 3868 1942
rect 3872 1932 3902 1946
rect 3930 1932 3943 1970
rect 4015 1976 4050 1984
rect 4015 1950 4016 1976
rect 4023 1950 4050 1976
rect 3958 1932 3988 1946
rect 4015 1942 4050 1950
rect 4052 1976 4093 1984
rect 4052 1950 4067 1976
rect 4074 1950 4093 1976
rect 4157 1972 4219 1984
rect 4231 1972 4306 1984
rect 4364 1972 4439 1984
rect 4451 1972 4482 1984
rect 4488 1972 4523 1984
rect 4157 1970 4319 1972
rect 4052 1942 4093 1950
rect 4175 1946 4188 1970
rect 4203 1968 4218 1970
rect 4015 1932 4016 1942
rect 4031 1932 4044 1942
rect 4058 1932 4059 1942
rect 4074 1932 4087 1942
rect 4102 1932 4132 1946
rect 4175 1932 4218 1946
rect 4242 1943 4249 1950
rect 4252 1946 4319 1970
rect 4351 1970 4523 1972
rect 4321 1948 4349 1952
rect 4351 1948 4431 1970
rect 4452 1968 4467 1970
rect 4321 1946 4431 1948
rect 4252 1942 4431 1946
rect 4225 1932 4255 1942
rect 4257 1932 4410 1942
rect 4418 1932 4448 1942
rect 4452 1932 4482 1946
rect 4510 1932 4523 1970
rect 4595 1976 4630 1984
rect 4595 1950 4596 1976
rect 4603 1950 4630 1976
rect 4538 1932 4568 1946
rect 4595 1942 4630 1950
rect 4632 1976 4673 1984
rect 4632 1950 4647 1976
rect 4654 1950 4673 1976
rect 4737 1972 4799 1984
rect 4811 1972 4886 1984
rect 4944 1972 5019 1984
rect 5031 1972 5062 1984
rect 5068 1972 5103 1984
rect 4737 1970 4899 1972
rect 4632 1942 4673 1950
rect 4755 1946 4768 1970
rect 4783 1968 4798 1970
rect 4832 1952 4899 1970
rect 4931 1970 5103 1972
rect 4931 1952 5011 1970
rect 5032 1968 5047 1970
rect 4595 1932 4596 1942
rect 4611 1932 4624 1942
rect 4638 1932 4639 1942
rect 4654 1932 4667 1942
rect 4682 1932 4712 1946
rect 4755 1932 4798 1946
rect 4822 1943 4829 1950
rect 4832 1942 5011 1952
rect 4805 1932 4835 1942
rect 4837 1932 4990 1942
rect 4998 1932 5028 1942
rect 5032 1932 5062 1946
rect 5090 1932 5103 1970
rect 5175 1976 5210 1984
rect 5175 1950 5176 1976
rect 5183 1950 5210 1976
rect 5118 1932 5148 1946
rect 5175 1942 5210 1950
rect 5212 1976 5253 1984
rect 5212 1950 5227 1976
rect 5234 1950 5253 1976
rect 5317 1972 5379 1984
rect 5391 1972 5466 1984
rect 5524 1972 5599 1984
rect 5611 1972 5642 1984
rect 5648 1972 5683 1984
rect 5317 1970 5479 1972
rect 5212 1942 5253 1950
rect 5335 1946 5348 1970
rect 5363 1968 5378 1970
rect 5412 1952 5479 1970
rect 5511 1970 5683 1972
rect 5511 1952 5591 1970
rect 5612 1968 5627 1970
rect 5175 1932 5176 1942
rect 5191 1932 5204 1942
rect 5218 1932 5219 1942
rect 5234 1932 5247 1942
rect 5262 1932 5292 1946
rect 5335 1932 5378 1946
rect 5402 1943 5409 1950
rect 5412 1942 5591 1952
rect 5385 1932 5415 1942
rect 5417 1932 5570 1942
rect 5578 1932 5608 1942
rect 5612 1932 5642 1946
rect 5670 1932 5683 1970
rect 5755 1976 5790 1984
rect 5755 1950 5756 1976
rect 5763 1950 5790 1976
rect 5698 1932 5728 1946
rect 5755 1942 5790 1950
rect 5792 1976 5833 1984
rect 5792 1950 5807 1976
rect 5814 1950 5833 1976
rect 5897 1972 5959 1984
rect 5971 1972 6046 1984
rect 6104 1972 6179 1984
rect 6191 1972 6222 1984
rect 6228 1972 6263 1984
rect 5897 1970 6059 1972
rect 5792 1942 5833 1950
rect 5915 1946 5928 1970
rect 5943 1968 5958 1970
rect 5992 1952 6059 1970
rect 6091 1970 6263 1972
rect 6091 1952 6171 1970
rect 6192 1968 6207 1970
rect 5755 1932 5756 1942
rect 5771 1932 5784 1942
rect 5798 1932 5799 1942
rect 5814 1932 5827 1942
rect 5842 1932 5872 1946
rect 5915 1932 5958 1946
rect 5982 1943 5989 1950
rect 5992 1942 6171 1952
rect 5965 1932 5995 1942
rect 5997 1932 6150 1942
rect 6158 1932 6188 1942
rect 6192 1932 6222 1946
rect 6250 1932 6263 1970
rect 6335 1976 6370 1984
rect 6335 1950 6336 1976
rect 6343 1950 6370 1976
rect 6278 1932 6308 1946
rect 6335 1942 6370 1950
rect 6372 1976 6413 1984
rect 6372 1950 6387 1976
rect 6394 1950 6413 1976
rect 6477 1972 6539 1984
rect 6551 1972 6626 1984
rect 6684 1972 6759 1984
rect 6771 1972 6802 1984
rect 6808 1972 6843 1984
rect 6477 1970 6639 1972
rect 6372 1942 6413 1950
rect 6495 1946 6508 1970
rect 6523 1968 6538 1970
rect 6572 1952 6639 1970
rect 6671 1970 6843 1972
rect 6671 1952 6751 1970
rect 6772 1968 6787 1970
rect 6335 1932 6336 1942
rect 6351 1932 6364 1942
rect 6378 1932 6379 1942
rect 6394 1932 6407 1942
rect 6422 1932 6452 1946
rect 6495 1932 6538 1946
rect 6562 1943 6569 1950
rect 6572 1942 6751 1952
rect 6545 1932 6575 1942
rect 6577 1932 6730 1942
rect 6738 1932 6768 1942
rect 6772 1932 6802 1946
rect 6830 1932 6843 1970
rect 6915 1976 6950 1984
rect 6915 1950 6916 1976
rect 6923 1950 6950 1976
rect 6858 1932 6888 1946
rect 6915 1942 6950 1950
rect 6915 1932 6916 1942
rect 6931 1932 6944 1942
rect -2 1926 1281 1932
rect -1 1918 1281 1926
rect 3481 1918 6944 1932
rect 14 1888 27 1918
rect 42 1900 72 1918
rect 115 1904 129 1918
rect 165 1904 385 1918
rect 116 1902 129 1904
rect 82 1890 97 1902
rect 79 1888 101 1890
rect 106 1888 136 1902
rect 197 1900 350 1904
rect 179 1888 371 1900
rect 414 1888 444 1902
rect 450 1888 463 1918
rect 478 1900 508 1918
rect 551 1888 564 1918
rect 594 1888 607 1918
rect 622 1900 652 1918
rect 695 1904 709 1918
rect 745 1904 965 1918
rect 696 1902 709 1904
rect 662 1890 677 1902
rect 659 1888 681 1890
rect 686 1888 716 1902
rect 777 1900 930 1904
rect 759 1888 951 1900
rect 994 1888 1024 1902
rect 1030 1888 1043 1918
rect 1058 1900 1088 1918
rect 1131 1888 1144 1918
rect 1174 1888 1187 1918
rect 1202 1900 1232 1918
rect 1275 1904 1281 1918
rect 1276 1902 1281 1904
rect 1242 1890 1257 1902
rect 1239 1888 1261 1890
rect 1266 1888 1281 1902
rect 3494 1888 3507 1918
rect 3522 1900 3552 1918
rect 3595 1904 3609 1918
rect 3645 1904 3865 1918
rect 3596 1902 3609 1904
rect 3562 1890 3577 1902
rect 3559 1888 3581 1890
rect 3586 1888 3616 1902
rect 3677 1900 3830 1904
rect 3659 1888 3851 1900
rect 3894 1888 3924 1902
rect 3930 1888 3943 1918
rect 3958 1900 3988 1918
rect 4031 1888 4044 1918
rect 4074 1888 4087 1918
rect 4102 1900 4132 1918
rect 4175 1904 4189 1918
rect 4225 1904 4445 1918
rect 4176 1902 4189 1904
rect 4142 1890 4157 1902
rect 4139 1888 4161 1890
rect 4166 1888 4196 1902
rect 4257 1900 4410 1904
rect 4239 1888 4431 1900
rect 4474 1888 4504 1902
rect 4510 1888 4523 1918
rect 4538 1900 4568 1918
rect 4611 1888 4624 1918
rect 4654 1888 4667 1918
rect 4682 1900 4712 1918
rect 4755 1904 4769 1918
rect 4805 1904 5025 1918
rect 4756 1902 4769 1904
rect 4722 1890 4737 1902
rect 4719 1888 4741 1890
rect 4746 1888 4776 1902
rect 4837 1900 4990 1904
rect 4819 1888 5011 1900
rect 5054 1888 5084 1902
rect 5090 1888 5103 1918
rect 5118 1900 5148 1918
rect 5191 1888 5204 1918
rect 5234 1888 5247 1918
rect 5262 1900 5292 1918
rect 5335 1904 5349 1918
rect 5385 1904 5605 1918
rect 5336 1902 5349 1904
rect 5302 1890 5317 1902
rect 5299 1888 5321 1890
rect 5326 1888 5356 1902
rect 5417 1900 5570 1904
rect 5399 1888 5591 1900
rect 5634 1888 5664 1902
rect 5670 1888 5683 1918
rect 5698 1900 5728 1918
rect 5771 1888 5784 1918
rect 5814 1888 5827 1918
rect 5842 1900 5872 1918
rect 5915 1904 5929 1918
rect 5965 1904 6185 1918
rect 5916 1902 5929 1904
rect 5882 1890 5897 1902
rect 5879 1888 5901 1890
rect 5906 1888 5936 1902
rect 5997 1900 6150 1904
rect 5979 1888 6171 1900
rect 6214 1888 6244 1902
rect 6250 1888 6263 1918
rect 6278 1900 6308 1918
rect 6351 1888 6364 1918
rect 6394 1888 6407 1918
rect 6422 1900 6452 1918
rect 6495 1904 6509 1918
rect 6545 1904 6765 1918
rect 6496 1902 6509 1904
rect 6462 1890 6477 1902
rect 6459 1888 6481 1890
rect 6486 1888 6516 1902
rect 6577 1900 6730 1904
rect 6559 1888 6751 1900
rect 6794 1888 6824 1902
rect 6830 1888 6843 1918
rect 6858 1900 6888 1918
rect 6931 1888 6944 1918
rect -1 1874 1281 1888
rect 3481 1874 6944 1888
rect 14 1770 27 1874
rect 72 1852 73 1862
rect 88 1852 101 1862
rect 72 1848 101 1852
rect 106 1848 136 1874
rect 154 1860 170 1862
rect 242 1860 295 1874
rect 243 1858 307 1860
rect 350 1858 365 1874
rect 414 1871 444 1874
rect 414 1868 450 1871
rect 380 1860 396 1862
rect 154 1848 169 1852
rect 72 1846 169 1848
rect 197 1846 365 1858
rect 381 1848 396 1852
rect 414 1849 453 1868
rect 472 1862 479 1863
rect 478 1855 479 1862
rect 462 1852 463 1855
rect 478 1852 491 1855
rect 414 1848 444 1849
rect 453 1848 459 1849
rect 462 1848 491 1852
rect 381 1847 491 1848
rect 381 1846 497 1847
rect 56 1838 107 1846
rect 56 1826 81 1838
rect 88 1826 107 1838
rect 138 1838 188 1846
rect 138 1830 154 1838
rect 161 1836 188 1838
rect 197 1836 418 1846
rect 161 1826 418 1836
rect 447 1838 497 1846
rect 447 1829 463 1838
rect 56 1818 107 1826
rect 154 1818 418 1826
rect 444 1826 463 1829
rect 470 1826 497 1838
rect 444 1818 497 1826
rect 72 1810 73 1818
rect 88 1810 101 1818
rect 72 1802 88 1810
rect 69 1795 88 1798
rect 69 1786 91 1795
rect 42 1776 91 1786
rect 42 1770 72 1776
rect 91 1771 96 1776
rect 14 1754 88 1770
rect 106 1762 136 1818
rect 171 1808 379 1818
rect 414 1814 459 1818
rect 462 1817 463 1818
rect 478 1817 491 1818
rect 197 1778 386 1808
rect 212 1775 386 1778
rect 205 1772 386 1775
rect 14 1752 27 1754
rect 42 1752 76 1754
rect 14 1736 88 1752
rect 115 1748 128 1762
rect 143 1748 159 1764
rect 205 1759 216 1772
rect -2 1714 -1 1730
rect 14 1714 27 1736
rect 42 1714 72 1736
rect 115 1732 177 1748
rect 205 1741 216 1757
rect 221 1752 231 1772
rect 241 1752 255 1772
rect 258 1759 267 1772
rect 283 1759 292 1772
rect 221 1741 255 1752
rect 258 1741 267 1757
rect 283 1741 292 1757
rect 299 1752 309 1772
rect 319 1752 333 1772
rect 334 1759 345 1772
rect 299 1741 333 1752
rect 334 1741 345 1757
rect 391 1748 407 1764
rect 414 1762 444 1814
rect 478 1810 479 1817
rect 463 1802 479 1810
rect 450 1770 463 1789
rect 478 1770 508 1786
rect 450 1754 524 1770
rect 450 1752 463 1754
rect 478 1752 512 1754
rect 115 1730 128 1732
rect 143 1730 177 1732
rect 115 1714 177 1730
rect 221 1725 237 1732
rect 299 1725 329 1736
rect 377 1732 423 1748
rect 450 1736 524 1752
rect 377 1730 411 1732
rect 376 1714 423 1730
rect 450 1714 463 1736
rect 478 1714 508 1736
rect 535 1714 536 1730
rect 551 1714 564 1874
rect 594 1770 607 1874
rect 652 1852 653 1862
rect 668 1852 681 1862
rect 652 1848 681 1852
rect 686 1848 716 1874
rect 734 1860 750 1862
rect 822 1860 875 1874
rect 823 1858 887 1860
rect 930 1858 945 1874
rect 994 1871 1024 1874
rect 994 1868 1030 1871
rect 960 1860 976 1862
rect 734 1848 749 1852
rect 652 1846 749 1848
rect 777 1846 945 1858
rect 961 1848 976 1852
rect 994 1849 1033 1868
rect 1052 1862 1059 1863
rect 1058 1855 1059 1862
rect 1042 1852 1043 1855
rect 1058 1852 1071 1855
rect 994 1848 1024 1849
rect 1033 1848 1039 1849
rect 1042 1848 1071 1852
rect 961 1847 1071 1848
rect 961 1846 1077 1847
rect 636 1838 687 1846
rect 636 1826 661 1838
rect 668 1826 687 1838
rect 718 1838 768 1846
rect 718 1830 734 1838
rect 741 1836 768 1838
rect 777 1836 998 1846
rect 741 1826 998 1836
rect 1027 1838 1077 1846
rect 1027 1829 1043 1838
rect 636 1818 687 1826
rect 734 1818 998 1826
rect 1024 1826 1043 1829
rect 1050 1826 1077 1838
rect 1024 1818 1077 1826
rect 652 1810 653 1818
rect 668 1810 681 1818
rect 652 1802 668 1810
rect 649 1795 668 1798
rect 649 1786 671 1795
rect 622 1776 671 1786
rect 622 1770 652 1776
rect 671 1771 676 1776
rect 594 1754 668 1770
rect 686 1762 716 1818
rect 751 1808 959 1818
rect 994 1814 1039 1818
rect 1042 1817 1043 1818
rect 1058 1817 1071 1818
rect 777 1778 966 1808
rect 792 1775 966 1778
rect 785 1772 966 1775
rect 594 1752 607 1754
rect 622 1752 656 1754
rect 594 1736 668 1752
rect 695 1748 708 1762
rect 723 1748 739 1764
rect 785 1759 796 1772
rect 578 1714 579 1730
rect 594 1714 607 1736
rect 622 1714 652 1736
rect 695 1732 757 1748
rect 785 1741 796 1757
rect 801 1752 811 1772
rect 821 1752 835 1772
rect 838 1759 847 1772
rect 863 1759 872 1772
rect 801 1741 835 1752
rect 838 1741 847 1757
rect 863 1741 872 1757
rect 879 1752 889 1772
rect 899 1752 913 1772
rect 914 1759 925 1772
rect 879 1741 913 1752
rect 914 1741 925 1757
rect 971 1748 987 1764
rect 994 1762 1024 1814
rect 1058 1810 1059 1817
rect 1043 1802 1059 1810
rect 1030 1770 1043 1789
rect 1058 1770 1088 1786
rect 1030 1754 1104 1770
rect 1030 1752 1043 1754
rect 1058 1752 1092 1754
rect 695 1730 708 1732
rect 723 1730 757 1732
rect 695 1714 757 1730
rect 801 1725 817 1732
rect 879 1725 909 1736
rect 957 1732 1003 1748
rect 1030 1736 1104 1752
rect 957 1730 991 1732
rect 956 1714 1003 1730
rect 1030 1714 1043 1736
rect 1058 1714 1088 1736
rect 1115 1714 1116 1730
rect 1131 1714 1144 1874
rect 1174 1770 1187 1874
rect 1232 1852 1233 1862
rect 1248 1852 1261 1862
rect 1232 1848 1261 1852
rect 1266 1848 1281 1874
rect 1232 1846 1281 1848
rect 1216 1838 1267 1846
rect 1216 1826 1241 1838
rect 1248 1826 1267 1838
rect 1216 1818 1267 1826
rect 1232 1810 1233 1818
rect 1248 1810 1261 1818
rect 1232 1802 1248 1810
rect 1229 1795 1248 1798
rect 1229 1786 1251 1795
rect 1202 1776 1251 1786
rect 1202 1770 1232 1776
rect 1251 1771 1256 1776
rect 1174 1754 1248 1770
rect 1266 1762 1281 1818
rect 1174 1752 1187 1754
rect 1202 1752 1236 1754
rect 1174 1736 1248 1752
rect 1158 1714 1159 1730
rect 1174 1714 1187 1736
rect 1202 1714 1232 1736
rect 1275 1714 1281 1762
rect 3494 1770 3507 1874
rect 3552 1852 3553 1862
rect 3568 1852 3581 1862
rect 3552 1848 3581 1852
rect 3586 1848 3616 1874
rect 3634 1860 3650 1862
rect 3722 1860 3775 1874
rect 3723 1858 3787 1860
rect 3830 1858 3845 1874
rect 3894 1871 3924 1874
rect 3894 1868 3930 1871
rect 3860 1860 3876 1862
rect 3634 1848 3649 1852
rect 3552 1846 3649 1848
rect 3677 1846 3845 1858
rect 3861 1848 3876 1852
rect 3894 1849 3933 1868
rect 3952 1862 3959 1863
rect 3958 1855 3959 1862
rect 3942 1852 3943 1855
rect 3958 1852 3971 1855
rect 3894 1848 3924 1849
rect 3933 1848 3939 1849
rect 3942 1848 3971 1852
rect 3861 1847 3971 1848
rect 3861 1846 3977 1847
rect 3536 1838 3587 1846
rect 3536 1826 3561 1838
rect 3568 1826 3587 1838
rect 3618 1838 3668 1846
rect 3618 1830 3634 1838
rect 3641 1836 3668 1838
rect 3677 1836 3898 1846
rect 3641 1826 3898 1836
rect 3927 1838 3977 1846
rect 3927 1829 3943 1838
rect 3536 1818 3587 1826
rect 3634 1818 3898 1826
rect 3924 1826 3943 1829
rect 3950 1826 3977 1838
rect 3924 1818 3977 1826
rect 3552 1810 3553 1818
rect 3568 1810 3581 1818
rect 3552 1802 3568 1810
rect 3549 1795 3568 1798
rect 3549 1786 3571 1795
rect 3522 1776 3571 1786
rect 3522 1770 3552 1776
rect 3571 1771 3576 1776
rect 3494 1754 3568 1770
rect 3586 1762 3616 1818
rect 3651 1808 3859 1818
rect 3894 1814 3939 1818
rect 3942 1817 3943 1818
rect 3958 1817 3971 1818
rect 3677 1778 3866 1808
rect 3692 1775 3866 1778
rect 3685 1772 3866 1775
rect 3494 1752 3507 1754
rect 3522 1752 3556 1754
rect 3494 1736 3568 1752
rect 3595 1748 3608 1762
rect 3623 1748 3639 1764
rect 3685 1759 3696 1772
rect 3494 1714 3507 1736
rect 3522 1714 3552 1736
rect 3595 1732 3657 1748
rect 3685 1741 3696 1757
rect 3701 1752 3711 1772
rect 3721 1752 3735 1772
rect 3738 1759 3747 1772
rect 3763 1759 3772 1772
rect 3701 1741 3735 1752
rect 3738 1741 3747 1757
rect 3763 1741 3772 1757
rect 3779 1752 3789 1772
rect 3799 1752 3813 1772
rect 3814 1759 3825 1772
rect 3779 1741 3813 1752
rect 3814 1741 3825 1757
rect 3871 1748 3887 1764
rect 3894 1762 3924 1814
rect 3958 1810 3959 1817
rect 3943 1802 3959 1810
rect 3930 1770 3943 1789
rect 3958 1770 3988 1786
rect 3930 1754 4004 1770
rect 3930 1752 3943 1754
rect 3958 1752 3992 1754
rect 3595 1730 3608 1732
rect 3623 1730 3657 1732
rect 3595 1714 3657 1730
rect 3701 1725 3717 1732
rect 3779 1725 3809 1736
rect 3857 1732 3903 1748
rect 3930 1736 4004 1752
rect 3857 1730 3891 1732
rect 3856 1714 3903 1730
rect 3930 1714 3943 1736
rect 3958 1714 3988 1736
rect 4015 1714 4016 1730
rect 4031 1714 4044 1874
rect 4074 1770 4087 1874
rect 4132 1852 4133 1862
rect 4148 1852 4161 1862
rect 4132 1848 4161 1852
rect 4166 1848 4196 1874
rect 4214 1860 4230 1862
rect 4302 1860 4355 1874
rect 4303 1858 4367 1860
rect 4410 1858 4425 1874
rect 4474 1871 4504 1874
rect 4474 1868 4510 1871
rect 4440 1860 4456 1862
rect 4214 1848 4229 1852
rect 4132 1846 4229 1848
rect 4257 1846 4425 1858
rect 4441 1848 4456 1852
rect 4474 1849 4513 1868
rect 4532 1862 4539 1863
rect 4538 1855 4539 1862
rect 4522 1852 4523 1855
rect 4538 1852 4551 1855
rect 4474 1848 4504 1849
rect 4513 1848 4519 1849
rect 4522 1848 4551 1852
rect 4441 1847 4551 1848
rect 4441 1846 4557 1847
rect 4116 1838 4167 1846
rect 4116 1826 4141 1838
rect 4148 1826 4167 1838
rect 4198 1838 4248 1846
rect 4198 1830 4214 1838
rect 4221 1836 4248 1838
rect 4257 1836 4478 1846
rect 4221 1826 4478 1836
rect 4507 1838 4557 1846
rect 4507 1829 4523 1838
rect 4116 1818 4167 1826
rect 4214 1818 4478 1826
rect 4504 1826 4523 1829
rect 4530 1826 4557 1838
rect 4504 1818 4557 1826
rect 4132 1810 4133 1818
rect 4148 1810 4161 1818
rect 4132 1802 4148 1810
rect 4129 1795 4148 1798
rect 4129 1786 4151 1795
rect 4102 1776 4151 1786
rect 4102 1770 4132 1776
rect 4151 1771 4156 1776
rect 4074 1754 4148 1770
rect 4166 1762 4196 1818
rect 4231 1808 4439 1818
rect 4474 1814 4519 1818
rect 4522 1817 4523 1818
rect 4538 1817 4551 1818
rect 4257 1778 4446 1808
rect 4272 1775 4446 1778
rect 4265 1772 4446 1775
rect 4074 1752 4087 1754
rect 4102 1752 4136 1754
rect 4074 1736 4148 1752
rect 4175 1748 4188 1762
rect 4203 1748 4219 1764
rect 4265 1759 4276 1772
rect 4058 1714 4059 1730
rect 4074 1714 4087 1736
rect 4102 1714 4132 1736
rect 4175 1732 4237 1748
rect 4265 1741 4276 1757
rect 4281 1752 4291 1772
rect 4301 1752 4315 1772
rect 4318 1759 4327 1772
rect 4343 1759 4352 1772
rect 4281 1741 4315 1752
rect 4318 1741 4327 1757
rect 4343 1741 4352 1757
rect 4359 1752 4369 1772
rect 4379 1752 4393 1772
rect 4394 1759 4405 1772
rect 4359 1741 4393 1752
rect 4394 1741 4405 1757
rect 4451 1748 4467 1764
rect 4474 1762 4504 1814
rect 4538 1810 4539 1817
rect 4523 1802 4539 1810
rect 4510 1770 4523 1789
rect 4538 1770 4568 1786
rect 4510 1754 4584 1770
rect 4510 1752 4523 1754
rect 4538 1752 4572 1754
rect 4175 1730 4188 1732
rect 4203 1730 4237 1732
rect 4175 1714 4237 1730
rect 4281 1725 4297 1732
rect 4359 1725 4389 1736
rect 4437 1732 4483 1748
rect 4510 1736 4584 1752
rect 4437 1730 4471 1732
rect 4436 1714 4483 1730
rect 4510 1714 4523 1736
rect 4538 1714 4568 1736
rect 4595 1714 4596 1730
rect 4611 1714 4624 1874
rect 4654 1770 4667 1874
rect 4712 1852 4713 1862
rect 4728 1852 4741 1862
rect 4712 1848 4741 1852
rect 4746 1848 4776 1874
rect 4794 1860 4810 1862
rect 4882 1860 4933 1874
rect 4883 1858 4947 1860
rect 4990 1858 5005 1874
rect 5054 1871 5084 1874
rect 5054 1868 5090 1871
rect 5020 1860 5036 1862
rect 4794 1848 4809 1852
rect 4712 1846 4809 1848
rect 4837 1846 5005 1858
rect 5021 1848 5036 1852
rect 5054 1849 5093 1868
rect 5112 1862 5119 1863
rect 5118 1855 5119 1862
rect 5102 1852 5103 1855
rect 5118 1852 5131 1855
rect 5054 1848 5084 1849
rect 5093 1848 5099 1849
rect 5102 1848 5131 1852
rect 5021 1847 5131 1848
rect 5021 1846 5137 1847
rect 4696 1838 4747 1846
rect 4696 1826 4721 1838
rect 4728 1826 4747 1838
rect 4778 1838 4828 1846
rect 4778 1830 4794 1838
rect 4801 1836 4828 1838
rect 4837 1836 5058 1846
rect 4801 1826 5058 1836
rect 5087 1838 5137 1846
rect 5087 1829 5103 1838
rect 4696 1818 4747 1826
rect 4794 1818 5058 1826
rect 5084 1826 5103 1829
rect 5110 1826 5137 1838
rect 5084 1818 5137 1826
rect 4712 1810 4713 1818
rect 4728 1810 4741 1818
rect 4712 1802 4728 1810
rect 4709 1795 4728 1798
rect 4709 1786 4731 1795
rect 4682 1776 4731 1786
rect 4682 1770 4712 1776
rect 4731 1771 4736 1776
rect 4654 1754 4728 1770
rect 4746 1762 4776 1818
rect 4811 1808 5019 1818
rect 5054 1814 5099 1818
rect 5102 1817 5103 1818
rect 5118 1817 5131 1818
rect 4837 1778 5026 1808
rect 4852 1775 5026 1778
rect 4845 1772 5026 1775
rect 4654 1752 4667 1754
rect 4682 1752 4716 1754
rect 4654 1736 4728 1752
rect 4755 1748 4768 1762
rect 4783 1748 4799 1764
rect 4845 1759 4856 1772
rect 4638 1714 4639 1730
rect 4654 1714 4667 1736
rect 4682 1714 4712 1736
rect 4755 1732 4817 1748
rect 4845 1741 4856 1757
rect 4861 1752 4871 1772
rect 4881 1752 4895 1772
rect 4898 1759 4907 1772
rect 4923 1759 4932 1772
rect 4861 1741 4895 1752
rect 4898 1741 4907 1757
rect 4923 1741 4932 1757
rect 4939 1752 4949 1772
rect 4959 1752 4973 1772
rect 4974 1759 4985 1772
rect 4939 1741 4973 1752
rect 4974 1741 4985 1757
rect 5031 1748 5047 1764
rect 5054 1762 5084 1814
rect 5118 1810 5119 1817
rect 5103 1802 5119 1810
rect 5090 1770 5103 1789
rect 5118 1770 5148 1786
rect 5090 1754 5164 1770
rect 5090 1752 5103 1754
rect 5118 1752 5152 1754
rect 4755 1730 4768 1732
rect 4783 1730 4817 1732
rect 4755 1714 4817 1730
rect 4861 1725 4877 1732
rect 4939 1725 4969 1736
rect 5017 1732 5063 1748
rect 5090 1736 5164 1752
rect 5017 1730 5051 1732
rect 5016 1714 5063 1730
rect 5090 1714 5103 1736
rect 5118 1714 5148 1736
rect 5175 1714 5176 1730
rect 5191 1714 5204 1874
rect 5234 1770 5247 1874
rect 5292 1852 5293 1862
rect 5308 1852 5321 1862
rect 5292 1848 5321 1852
rect 5326 1848 5356 1874
rect 5374 1860 5390 1862
rect 5462 1860 5513 1874
rect 5463 1858 5527 1860
rect 5570 1858 5585 1874
rect 5634 1871 5664 1874
rect 5634 1868 5670 1871
rect 5600 1860 5616 1862
rect 5374 1848 5389 1852
rect 5292 1846 5389 1848
rect 5417 1846 5585 1858
rect 5601 1848 5616 1852
rect 5634 1849 5673 1868
rect 5692 1862 5699 1863
rect 5698 1855 5699 1862
rect 5682 1852 5683 1855
rect 5698 1852 5711 1855
rect 5634 1848 5664 1849
rect 5673 1848 5679 1849
rect 5682 1848 5711 1852
rect 5601 1847 5711 1848
rect 5601 1846 5717 1847
rect 5276 1838 5327 1846
rect 5276 1826 5301 1838
rect 5308 1826 5327 1838
rect 5358 1838 5408 1846
rect 5358 1830 5374 1838
rect 5381 1836 5408 1838
rect 5417 1836 5638 1846
rect 5381 1826 5638 1836
rect 5667 1838 5717 1846
rect 5667 1829 5683 1838
rect 5276 1818 5327 1826
rect 5374 1818 5638 1826
rect 5664 1826 5683 1829
rect 5690 1826 5717 1838
rect 5664 1818 5717 1826
rect 5292 1810 5293 1818
rect 5308 1810 5321 1818
rect 5292 1802 5308 1810
rect 5289 1795 5308 1798
rect 5289 1786 5311 1795
rect 5262 1776 5311 1786
rect 5262 1770 5292 1776
rect 5311 1771 5316 1776
rect 5234 1754 5308 1770
rect 5326 1762 5356 1818
rect 5391 1808 5599 1818
rect 5634 1814 5679 1818
rect 5682 1817 5683 1818
rect 5698 1817 5711 1818
rect 5417 1778 5606 1808
rect 5432 1775 5606 1778
rect 5425 1772 5606 1775
rect 5234 1752 5247 1754
rect 5262 1752 5296 1754
rect 5234 1736 5308 1752
rect 5335 1748 5348 1762
rect 5363 1748 5379 1764
rect 5425 1759 5436 1772
rect 5218 1714 5219 1730
rect 5234 1714 5247 1736
rect 5262 1714 5292 1736
rect 5335 1732 5397 1748
rect 5425 1741 5436 1757
rect 5441 1752 5451 1772
rect 5461 1752 5475 1772
rect 5478 1759 5487 1772
rect 5503 1759 5512 1772
rect 5441 1741 5475 1752
rect 5478 1741 5487 1757
rect 5503 1741 5512 1757
rect 5519 1752 5529 1772
rect 5539 1752 5553 1772
rect 5554 1759 5565 1772
rect 5519 1741 5553 1752
rect 5554 1741 5565 1757
rect 5611 1748 5627 1764
rect 5634 1762 5664 1814
rect 5698 1810 5699 1817
rect 5683 1802 5699 1810
rect 5670 1770 5683 1789
rect 5698 1770 5728 1786
rect 5670 1754 5744 1770
rect 5670 1752 5683 1754
rect 5698 1752 5732 1754
rect 5335 1730 5348 1732
rect 5363 1730 5397 1732
rect 5335 1714 5397 1730
rect 5441 1725 5457 1732
rect 5519 1725 5549 1736
rect 5597 1732 5643 1748
rect 5670 1736 5744 1752
rect 5597 1730 5631 1732
rect 5596 1714 5643 1730
rect 5670 1714 5683 1736
rect 5698 1714 5728 1736
rect 5755 1714 5756 1730
rect 5771 1714 5784 1874
rect 5814 1770 5827 1874
rect 5872 1852 5873 1862
rect 5888 1852 5901 1862
rect 5872 1848 5901 1852
rect 5906 1848 5936 1874
rect 5954 1860 5970 1862
rect 6042 1860 6093 1874
rect 6043 1858 6107 1860
rect 6150 1858 6165 1874
rect 6214 1871 6244 1874
rect 6214 1868 6250 1871
rect 6180 1860 6196 1862
rect 5954 1848 5969 1852
rect 5872 1846 5969 1848
rect 5997 1846 6165 1858
rect 6181 1848 6196 1852
rect 6214 1849 6253 1868
rect 6272 1862 6279 1863
rect 6278 1855 6279 1862
rect 6262 1852 6263 1855
rect 6278 1852 6291 1855
rect 6214 1848 6244 1849
rect 6253 1848 6259 1849
rect 6262 1848 6291 1852
rect 6181 1847 6291 1848
rect 6181 1846 6297 1847
rect 5856 1838 5907 1846
rect 5856 1826 5881 1838
rect 5888 1826 5907 1838
rect 5938 1838 5988 1846
rect 5938 1830 5954 1838
rect 5961 1836 5988 1838
rect 5997 1836 6218 1846
rect 5961 1826 6218 1836
rect 6247 1838 6297 1846
rect 6247 1829 6263 1838
rect 5856 1818 5907 1826
rect 5954 1818 6218 1826
rect 6244 1826 6263 1829
rect 6270 1826 6297 1838
rect 6244 1818 6297 1826
rect 5872 1810 5873 1818
rect 5888 1810 5901 1818
rect 5872 1802 5888 1810
rect 5869 1795 5888 1798
rect 5869 1786 5891 1795
rect 5842 1776 5891 1786
rect 5842 1770 5872 1776
rect 5891 1771 5896 1776
rect 5814 1754 5888 1770
rect 5906 1762 5936 1818
rect 5971 1808 6179 1818
rect 6214 1814 6259 1818
rect 6262 1817 6263 1818
rect 6278 1817 6291 1818
rect 5997 1778 6186 1808
rect 6012 1775 6186 1778
rect 6005 1772 6186 1775
rect 5814 1752 5827 1754
rect 5842 1752 5876 1754
rect 5814 1736 5888 1752
rect 5915 1748 5928 1762
rect 5943 1748 5959 1764
rect 6005 1759 6016 1772
rect 5798 1714 5799 1730
rect 5814 1714 5827 1736
rect 5842 1714 5872 1736
rect 5915 1732 5977 1748
rect 6005 1741 6016 1757
rect 6021 1752 6031 1772
rect 6041 1752 6055 1772
rect 6058 1759 6067 1772
rect 6083 1759 6092 1772
rect 6021 1741 6055 1752
rect 6058 1741 6067 1757
rect 6083 1741 6092 1757
rect 6099 1752 6109 1772
rect 6119 1752 6133 1772
rect 6134 1759 6145 1772
rect 6099 1741 6133 1752
rect 6134 1741 6145 1757
rect 6191 1748 6207 1764
rect 6214 1762 6244 1814
rect 6278 1810 6279 1817
rect 6263 1802 6279 1810
rect 6250 1770 6263 1789
rect 6278 1770 6308 1786
rect 6250 1754 6324 1770
rect 6250 1752 6263 1754
rect 6278 1752 6312 1754
rect 5915 1730 5928 1732
rect 5943 1730 5977 1732
rect 5915 1714 5977 1730
rect 6021 1725 6037 1732
rect 6099 1725 6129 1736
rect 6177 1732 6223 1748
rect 6250 1736 6324 1752
rect 6177 1730 6211 1732
rect 6176 1714 6223 1730
rect 6250 1714 6263 1736
rect 6278 1714 6308 1736
rect 6335 1714 6336 1730
rect 6351 1714 6364 1874
rect 6394 1770 6407 1874
rect 6452 1852 6453 1862
rect 6468 1852 6481 1862
rect 6452 1848 6481 1852
rect 6486 1848 6516 1874
rect 6534 1860 6550 1862
rect 6622 1860 6673 1874
rect 6623 1858 6687 1860
rect 6730 1858 6745 1874
rect 6794 1871 6824 1874
rect 6794 1868 6830 1871
rect 6760 1860 6776 1862
rect 6534 1848 6549 1852
rect 6452 1846 6549 1848
rect 6577 1846 6745 1858
rect 6761 1848 6776 1852
rect 6794 1849 6833 1868
rect 6852 1862 6859 1863
rect 6858 1855 6859 1862
rect 6842 1852 6843 1855
rect 6858 1852 6871 1855
rect 6794 1848 6824 1849
rect 6833 1848 6839 1849
rect 6842 1848 6871 1852
rect 6761 1847 6871 1848
rect 6761 1846 6877 1847
rect 6436 1838 6487 1846
rect 6436 1826 6461 1838
rect 6468 1826 6487 1838
rect 6518 1838 6568 1846
rect 6518 1830 6534 1838
rect 6541 1836 6568 1838
rect 6577 1836 6798 1846
rect 6541 1826 6798 1836
rect 6827 1838 6877 1846
rect 6827 1829 6843 1838
rect 6436 1818 6487 1826
rect 6534 1818 6798 1826
rect 6824 1826 6843 1829
rect 6850 1826 6877 1838
rect 6824 1818 6877 1826
rect 6452 1810 6453 1818
rect 6468 1810 6481 1818
rect 6452 1802 6468 1810
rect 6449 1795 6468 1798
rect 6449 1786 6471 1795
rect 6422 1776 6471 1786
rect 6422 1770 6452 1776
rect 6471 1771 6476 1776
rect 6394 1754 6468 1770
rect 6486 1762 6516 1818
rect 6551 1808 6759 1818
rect 6794 1814 6839 1818
rect 6842 1817 6843 1818
rect 6858 1817 6871 1818
rect 6577 1778 6766 1808
rect 6592 1775 6766 1778
rect 6585 1772 6766 1775
rect 6394 1752 6407 1754
rect 6422 1752 6456 1754
rect 6394 1736 6468 1752
rect 6495 1748 6508 1762
rect 6523 1748 6539 1764
rect 6585 1759 6596 1772
rect 6378 1714 6379 1730
rect 6394 1714 6407 1736
rect 6422 1714 6452 1736
rect 6495 1732 6557 1748
rect 6585 1741 6596 1757
rect 6601 1752 6611 1772
rect 6621 1752 6635 1772
rect 6638 1759 6647 1772
rect 6663 1759 6672 1772
rect 6601 1741 6635 1752
rect 6638 1741 6647 1757
rect 6663 1741 6672 1757
rect 6679 1752 6689 1772
rect 6699 1752 6713 1772
rect 6714 1759 6725 1772
rect 6679 1741 6713 1752
rect 6714 1741 6725 1757
rect 6771 1748 6787 1764
rect 6794 1762 6824 1814
rect 6858 1810 6859 1817
rect 6843 1802 6859 1810
rect 6830 1770 6843 1789
rect 6858 1770 6888 1786
rect 6830 1754 6904 1770
rect 6830 1752 6843 1754
rect 6858 1752 6892 1754
rect 6495 1730 6508 1732
rect 6523 1730 6557 1732
rect 6495 1714 6557 1730
rect 6601 1725 6617 1732
rect 6679 1725 6709 1736
rect 6757 1732 6803 1748
rect 6830 1736 6904 1752
rect 6757 1730 6791 1732
rect 6756 1714 6803 1730
rect 6830 1714 6843 1736
rect 6858 1714 6888 1736
rect 6915 1714 6916 1730
rect 6931 1714 6944 1874
rect -8 1706 33 1714
rect -8 1680 7 1706
rect 14 1680 33 1706
rect 97 1702 159 1714
rect 171 1702 246 1714
rect 304 1702 379 1714
rect 391 1702 422 1714
rect 428 1702 463 1714
rect 97 1700 259 1702
rect -8 1672 33 1680
rect 115 1676 128 1700
rect 143 1698 158 1700
rect -2 1662 -1 1672
rect 14 1662 27 1672
rect 42 1662 72 1676
rect 115 1662 158 1676
rect 182 1673 189 1680
rect 192 1676 259 1700
rect 291 1700 463 1702
rect 261 1678 289 1682
rect 291 1678 371 1700
rect 392 1698 407 1700
rect 261 1676 371 1678
rect 192 1672 371 1676
rect 165 1662 195 1672
rect 197 1662 350 1672
rect 358 1662 388 1672
rect 392 1662 422 1676
rect 450 1662 463 1700
rect 535 1706 570 1714
rect 535 1680 536 1706
rect 543 1680 570 1706
rect 478 1662 508 1676
rect 535 1672 570 1680
rect 572 1706 613 1714
rect 572 1680 587 1706
rect 594 1680 613 1706
rect 677 1702 739 1714
rect 751 1702 826 1714
rect 884 1702 959 1714
rect 971 1702 1002 1714
rect 1008 1702 1043 1714
rect 677 1700 839 1702
rect 572 1672 613 1680
rect 695 1676 708 1700
rect 723 1698 738 1700
rect 535 1662 536 1672
rect 551 1662 564 1672
rect 578 1662 579 1672
rect 594 1662 607 1672
rect 622 1662 652 1676
rect 695 1662 738 1676
rect 762 1673 769 1680
rect 772 1676 839 1700
rect 871 1700 1043 1702
rect 841 1678 869 1682
rect 871 1678 951 1700
rect 972 1698 987 1700
rect 841 1676 951 1678
rect 772 1672 951 1676
rect 745 1662 775 1672
rect 777 1662 930 1672
rect 938 1662 968 1672
rect 972 1662 1002 1676
rect 1030 1662 1043 1700
rect 1115 1706 1150 1714
rect 1115 1680 1116 1706
rect 1123 1680 1150 1706
rect 1058 1662 1088 1676
rect 1115 1672 1150 1680
rect 1152 1706 1193 1714
rect 1152 1680 1167 1706
rect 1174 1680 1193 1706
rect 1257 1700 1281 1714
rect 1152 1672 1193 1680
rect 1115 1662 1116 1672
rect 1131 1662 1144 1672
rect 1158 1662 1159 1672
rect 1174 1662 1187 1672
rect 1202 1662 1232 1676
rect 1275 1662 1281 1700
rect 3481 1706 3513 1714
rect 3481 1680 3487 1706
rect 3494 1680 3513 1706
rect 3577 1702 3639 1714
rect 3651 1702 3726 1714
rect 3784 1702 3859 1714
rect 3871 1702 3902 1714
rect 3908 1702 3943 1714
rect 3577 1700 3739 1702
rect 3481 1672 3513 1680
rect 3595 1676 3608 1700
rect 3623 1698 3638 1700
rect 3494 1662 3507 1672
rect 3522 1662 3552 1676
rect 3595 1662 3638 1676
rect 3662 1673 3669 1680
rect 3672 1676 3739 1700
rect 3771 1700 3943 1702
rect 3741 1678 3769 1682
rect 3771 1678 3851 1700
rect 3872 1698 3887 1700
rect 3741 1676 3851 1678
rect 3672 1672 3851 1676
rect 3645 1662 3675 1672
rect 3677 1662 3830 1672
rect 3838 1662 3868 1672
rect 3872 1662 3902 1676
rect 3930 1662 3943 1700
rect 4015 1706 4050 1714
rect 4015 1680 4016 1706
rect 4023 1680 4050 1706
rect 3958 1662 3988 1676
rect 4015 1672 4050 1680
rect 4052 1706 4093 1714
rect 4052 1680 4067 1706
rect 4074 1680 4093 1706
rect 4157 1702 4219 1714
rect 4231 1702 4306 1714
rect 4364 1702 4439 1714
rect 4451 1702 4482 1714
rect 4488 1702 4523 1714
rect 4157 1700 4319 1702
rect 4052 1672 4093 1680
rect 4175 1676 4188 1700
rect 4203 1698 4218 1700
rect 4015 1662 4016 1672
rect 4031 1662 4044 1672
rect 4058 1662 4059 1672
rect 4074 1662 4087 1672
rect 4102 1662 4132 1676
rect 4175 1662 4218 1676
rect 4242 1673 4249 1680
rect 4252 1676 4319 1700
rect 4351 1700 4523 1702
rect 4321 1678 4349 1682
rect 4351 1678 4431 1700
rect 4452 1698 4467 1700
rect 4321 1676 4431 1678
rect 4252 1672 4431 1676
rect 4225 1662 4255 1672
rect 4257 1662 4410 1672
rect 4418 1662 4448 1672
rect 4452 1662 4482 1676
rect 4510 1662 4523 1700
rect 4595 1706 4630 1714
rect 4595 1680 4596 1706
rect 4603 1680 4630 1706
rect 4538 1662 4568 1676
rect 4595 1672 4630 1680
rect 4632 1706 4673 1714
rect 4632 1680 4647 1706
rect 4654 1680 4673 1706
rect 4737 1702 4799 1714
rect 4811 1702 4886 1714
rect 4944 1702 5019 1714
rect 5031 1702 5062 1714
rect 5068 1702 5103 1714
rect 4737 1700 4899 1702
rect 4755 1682 4768 1700
rect 4783 1698 4798 1700
rect 4632 1672 4673 1680
rect 4756 1676 4768 1682
rect 4832 1682 4899 1700
rect 4931 1700 5103 1702
rect 4931 1682 5011 1700
rect 5032 1698 5047 1700
rect 4595 1662 4596 1672
rect 4611 1662 4624 1672
rect 4638 1662 4639 1672
rect 4654 1662 4667 1672
rect 4682 1662 4712 1676
rect 4756 1662 4798 1676
rect 4822 1673 4829 1680
rect 4832 1672 5011 1682
rect 4805 1662 4835 1672
rect 4837 1662 4990 1672
rect 4998 1662 5028 1672
rect 5032 1662 5062 1676
rect 5090 1662 5103 1700
rect 5175 1706 5210 1714
rect 5175 1680 5176 1706
rect 5183 1680 5210 1706
rect 5118 1662 5148 1676
rect 5175 1672 5210 1680
rect 5212 1706 5253 1714
rect 5212 1680 5227 1706
rect 5234 1680 5253 1706
rect 5317 1702 5379 1714
rect 5391 1702 5466 1714
rect 5524 1702 5599 1714
rect 5611 1702 5642 1714
rect 5648 1702 5683 1714
rect 5317 1700 5479 1702
rect 5335 1682 5348 1700
rect 5363 1698 5378 1700
rect 5212 1672 5253 1680
rect 5336 1676 5348 1682
rect 5412 1682 5479 1700
rect 5511 1700 5683 1702
rect 5511 1682 5591 1700
rect 5612 1698 5627 1700
rect 5175 1662 5176 1672
rect 5191 1662 5204 1672
rect 5218 1662 5219 1672
rect 5234 1662 5247 1672
rect 5262 1662 5292 1676
rect 5336 1662 5378 1676
rect 5402 1673 5409 1680
rect 5412 1672 5591 1682
rect 5385 1662 5415 1672
rect 5417 1662 5570 1672
rect 5578 1662 5608 1672
rect 5612 1662 5642 1676
rect 5670 1662 5683 1700
rect 5755 1706 5790 1714
rect 5755 1680 5756 1706
rect 5763 1680 5790 1706
rect 5698 1662 5728 1676
rect 5755 1672 5790 1680
rect 5792 1706 5833 1714
rect 5792 1680 5807 1706
rect 5814 1680 5833 1706
rect 5897 1702 5959 1714
rect 5971 1702 6046 1714
rect 6104 1702 6179 1714
rect 6191 1702 6222 1714
rect 6228 1702 6263 1714
rect 5897 1700 6059 1702
rect 5915 1682 5928 1700
rect 5943 1698 5958 1700
rect 5792 1672 5833 1680
rect 5916 1676 5928 1682
rect 5992 1682 6059 1700
rect 6091 1700 6263 1702
rect 6091 1682 6171 1700
rect 6192 1698 6207 1700
rect 5755 1662 5756 1672
rect 5771 1662 5784 1672
rect 5798 1662 5799 1672
rect 5814 1662 5827 1672
rect 5842 1662 5872 1676
rect 5916 1662 5958 1676
rect 5982 1673 5989 1680
rect 5992 1672 6171 1682
rect 5965 1662 5995 1672
rect 5997 1662 6150 1672
rect 6158 1662 6188 1672
rect 6192 1662 6222 1676
rect 6250 1662 6263 1700
rect 6335 1706 6370 1714
rect 6335 1680 6336 1706
rect 6343 1680 6370 1706
rect 6278 1662 6308 1676
rect 6335 1672 6370 1680
rect 6372 1706 6413 1714
rect 6372 1680 6387 1706
rect 6394 1680 6413 1706
rect 6477 1702 6539 1714
rect 6551 1702 6626 1714
rect 6684 1702 6759 1714
rect 6771 1702 6802 1714
rect 6808 1702 6843 1714
rect 6477 1700 6639 1702
rect 6495 1682 6508 1700
rect 6523 1698 6538 1700
rect 6372 1672 6413 1680
rect 6496 1676 6508 1682
rect 6572 1682 6639 1700
rect 6671 1700 6843 1702
rect 6671 1682 6751 1700
rect 6772 1698 6787 1700
rect 6335 1662 6336 1672
rect 6351 1662 6364 1672
rect 6378 1662 6379 1672
rect 6394 1662 6407 1672
rect 6422 1662 6452 1676
rect 6496 1662 6538 1676
rect 6562 1673 6569 1680
rect 6572 1672 6751 1682
rect 6545 1662 6575 1672
rect 6577 1662 6730 1672
rect 6738 1662 6768 1672
rect 6772 1662 6802 1676
rect 6830 1662 6843 1700
rect 6915 1706 6950 1714
rect 6915 1680 6916 1706
rect 6923 1680 6950 1706
rect 6858 1662 6888 1676
rect 6915 1672 6950 1680
rect 6915 1662 6916 1672
rect 6931 1662 6944 1672
rect -2 1656 1281 1662
rect -1 1648 1281 1656
rect 3481 1648 6944 1662
rect 14 1618 27 1648
rect 42 1630 72 1648
rect 115 1634 129 1648
rect 165 1634 385 1648
rect 116 1632 129 1634
rect 82 1620 97 1632
rect 79 1618 101 1620
rect 106 1618 136 1632
rect 197 1630 350 1634
rect 179 1618 371 1630
rect 414 1618 444 1632
rect 450 1618 463 1648
rect 478 1630 508 1648
rect 551 1618 564 1648
rect 594 1618 607 1648
rect 622 1630 652 1648
rect 695 1634 709 1648
rect 745 1634 965 1648
rect 696 1632 709 1634
rect 662 1620 677 1632
rect 659 1618 681 1620
rect 686 1618 716 1632
rect 777 1630 930 1634
rect 759 1618 951 1630
rect 994 1618 1024 1632
rect 1030 1618 1043 1648
rect 1058 1630 1088 1648
rect 1131 1618 1144 1648
rect 1174 1618 1187 1648
rect 1202 1630 1232 1648
rect 1275 1634 1281 1648
rect 1276 1632 1281 1634
rect 1242 1620 1257 1632
rect 1239 1618 1261 1620
rect 1266 1618 1281 1632
rect 3494 1618 3507 1648
rect 3522 1630 3552 1648
rect 3595 1634 3609 1648
rect 3645 1634 3865 1648
rect 3596 1632 3609 1634
rect 3562 1620 3577 1632
rect 3559 1618 3581 1620
rect 3586 1618 3616 1632
rect 3677 1630 3830 1634
rect 3659 1618 3851 1630
rect 3894 1618 3924 1632
rect 3930 1618 3943 1648
rect 3958 1630 3988 1648
rect 4031 1618 4044 1648
rect 4074 1618 4087 1648
rect 4102 1630 4132 1648
rect 4175 1634 4189 1648
rect 4225 1634 4445 1648
rect 4176 1632 4189 1634
rect 4142 1620 4157 1632
rect 4139 1618 4161 1620
rect 4166 1618 4196 1632
rect 4257 1630 4410 1634
rect 4239 1618 4431 1630
rect 4474 1618 4504 1632
rect 4510 1618 4523 1648
rect 4538 1630 4568 1648
rect 4611 1618 4624 1648
rect 4654 1618 4667 1648
rect 4682 1630 4712 1648
rect 4756 1632 4769 1648
rect 4805 1634 5025 1648
rect 4722 1620 4737 1632
rect 4719 1618 4741 1620
rect 4746 1618 4776 1632
rect 4837 1630 4990 1634
rect 4819 1618 5011 1630
rect 5054 1618 5084 1632
rect 5090 1618 5103 1648
rect 5118 1630 5148 1648
rect 5191 1618 5204 1648
rect 5234 1618 5247 1648
rect 5262 1630 5292 1648
rect 5336 1632 5349 1648
rect 5385 1634 5605 1648
rect 5302 1620 5317 1632
rect 5299 1618 5321 1620
rect 5326 1618 5356 1632
rect 5417 1630 5570 1634
rect 5399 1618 5591 1630
rect 5634 1618 5664 1632
rect 5670 1618 5683 1648
rect 5698 1630 5728 1648
rect 5771 1618 5784 1648
rect 5814 1618 5827 1648
rect 5842 1630 5872 1648
rect 5916 1632 5929 1648
rect 5965 1634 6185 1648
rect 5882 1620 5897 1632
rect 5879 1618 5901 1620
rect 5906 1618 5936 1632
rect 5997 1630 6150 1634
rect 5979 1618 6171 1630
rect 6214 1618 6244 1632
rect 6250 1618 6263 1648
rect 6278 1630 6308 1648
rect 6351 1618 6364 1648
rect 6394 1618 6407 1648
rect 6422 1630 6452 1648
rect 6496 1632 6509 1648
rect 6545 1634 6765 1648
rect 6462 1620 6477 1632
rect 6459 1618 6481 1620
rect 6486 1618 6516 1632
rect 6577 1630 6730 1634
rect 6559 1618 6751 1630
rect 6794 1618 6824 1632
rect 6830 1618 6843 1648
rect 6858 1630 6888 1648
rect 6931 1618 6944 1648
rect -1 1604 1281 1618
rect 3481 1604 6944 1618
rect 14 1500 27 1604
rect 72 1582 73 1592
rect 88 1582 101 1592
rect 72 1578 101 1582
rect 106 1578 136 1604
rect 154 1590 170 1592
rect 242 1590 295 1604
rect 243 1588 307 1590
rect 350 1588 365 1604
rect 414 1601 444 1604
rect 414 1598 450 1601
rect 380 1590 396 1592
rect 154 1578 169 1582
rect 72 1576 169 1578
rect 197 1576 365 1588
rect 381 1578 396 1582
rect 414 1579 453 1598
rect 472 1592 479 1593
rect 478 1585 479 1592
rect 462 1582 463 1585
rect 478 1582 491 1585
rect 414 1578 444 1579
rect 453 1578 459 1579
rect 462 1578 491 1582
rect 381 1577 491 1578
rect 381 1576 497 1577
rect 56 1568 107 1576
rect 56 1556 81 1568
rect 88 1556 107 1568
rect 138 1568 188 1576
rect 138 1560 154 1568
rect 161 1566 188 1568
rect 197 1566 418 1576
rect 161 1556 418 1566
rect 447 1568 497 1576
rect 447 1559 463 1568
rect 56 1548 107 1556
rect 154 1548 418 1556
rect 444 1556 463 1559
rect 470 1556 497 1568
rect 444 1548 497 1556
rect 72 1540 73 1548
rect 88 1540 101 1548
rect 72 1532 88 1540
rect 69 1525 88 1528
rect 69 1516 91 1525
rect 42 1506 91 1516
rect 42 1500 72 1506
rect 91 1501 96 1506
rect 14 1484 88 1500
rect 106 1492 136 1548
rect 171 1538 379 1548
rect 414 1544 459 1548
rect 462 1547 463 1548
rect 478 1547 491 1548
rect 197 1508 386 1538
rect 212 1505 386 1508
rect 205 1502 386 1505
rect 14 1482 27 1484
rect 42 1482 76 1484
rect 14 1466 88 1482
rect 115 1478 128 1492
rect 143 1478 159 1494
rect 205 1489 216 1502
rect -2 1444 -1 1460
rect 14 1444 27 1466
rect 42 1444 72 1466
rect 115 1462 177 1478
rect 205 1471 216 1487
rect 221 1482 231 1502
rect 241 1482 255 1502
rect 258 1489 267 1502
rect 283 1489 292 1502
rect 221 1471 255 1482
rect 258 1471 267 1487
rect 283 1471 292 1487
rect 299 1482 309 1502
rect 319 1482 333 1502
rect 334 1489 345 1502
rect 299 1471 333 1482
rect 334 1471 345 1487
rect 391 1478 407 1494
rect 414 1492 444 1544
rect 478 1540 479 1547
rect 463 1532 479 1540
rect 450 1500 463 1519
rect 478 1500 508 1516
rect 450 1484 524 1500
rect 450 1482 463 1484
rect 478 1482 512 1484
rect 115 1460 128 1462
rect 143 1460 177 1462
rect 115 1444 177 1460
rect 221 1455 237 1462
rect 299 1455 329 1466
rect 377 1462 423 1478
rect 450 1466 524 1482
rect 377 1460 411 1462
rect 376 1444 423 1460
rect 450 1444 463 1466
rect 478 1444 508 1466
rect 535 1444 536 1460
rect 551 1444 564 1604
rect 594 1500 607 1604
rect 652 1582 653 1592
rect 668 1582 681 1592
rect 652 1578 681 1582
rect 686 1578 716 1604
rect 734 1590 750 1592
rect 822 1590 875 1604
rect 823 1588 887 1590
rect 930 1588 945 1604
rect 994 1601 1024 1604
rect 994 1598 1030 1601
rect 960 1590 976 1592
rect 734 1578 749 1582
rect 652 1576 749 1578
rect 777 1576 945 1588
rect 961 1578 976 1582
rect 994 1579 1033 1598
rect 1052 1592 1059 1593
rect 1058 1585 1059 1592
rect 1042 1582 1043 1585
rect 1058 1582 1071 1585
rect 994 1578 1024 1579
rect 1033 1578 1039 1579
rect 1042 1578 1071 1582
rect 961 1577 1071 1578
rect 961 1576 1077 1577
rect 636 1568 687 1576
rect 636 1556 661 1568
rect 668 1556 687 1568
rect 718 1568 768 1576
rect 718 1560 734 1568
rect 741 1566 768 1568
rect 777 1566 998 1576
rect 741 1556 998 1566
rect 1027 1568 1077 1576
rect 1027 1559 1043 1568
rect 636 1548 687 1556
rect 734 1548 998 1556
rect 1024 1556 1043 1559
rect 1050 1556 1077 1568
rect 1024 1548 1077 1556
rect 652 1540 653 1548
rect 668 1540 681 1548
rect 652 1532 668 1540
rect 649 1525 668 1528
rect 649 1516 671 1525
rect 622 1506 671 1516
rect 622 1500 652 1506
rect 671 1501 676 1506
rect 594 1484 668 1500
rect 686 1492 716 1548
rect 751 1538 959 1548
rect 994 1544 1039 1548
rect 1042 1547 1043 1548
rect 1058 1547 1071 1548
rect 777 1508 966 1538
rect 792 1505 966 1508
rect 785 1502 966 1505
rect 594 1482 607 1484
rect 622 1482 656 1484
rect 594 1466 668 1482
rect 695 1478 708 1492
rect 723 1478 739 1494
rect 785 1489 796 1502
rect 578 1444 579 1460
rect 594 1444 607 1466
rect 622 1444 652 1466
rect 695 1462 757 1478
rect 785 1471 796 1487
rect 801 1482 811 1502
rect 821 1482 835 1502
rect 838 1489 847 1502
rect 863 1489 872 1502
rect 801 1471 835 1482
rect 838 1471 847 1487
rect 863 1471 872 1487
rect 879 1482 889 1502
rect 899 1482 913 1502
rect 914 1489 925 1502
rect 879 1471 913 1482
rect 914 1471 925 1487
rect 971 1478 987 1494
rect 994 1492 1024 1544
rect 1058 1540 1059 1547
rect 1043 1532 1059 1540
rect 1030 1500 1043 1519
rect 1058 1500 1088 1516
rect 1030 1484 1104 1500
rect 1030 1482 1043 1484
rect 1058 1482 1092 1484
rect 695 1460 708 1462
rect 723 1460 757 1462
rect 695 1444 757 1460
rect 801 1455 817 1462
rect 879 1455 909 1466
rect 957 1462 1003 1478
rect 1030 1466 1104 1482
rect 957 1460 991 1462
rect 956 1444 1003 1460
rect 1030 1444 1043 1466
rect 1058 1444 1088 1466
rect 1115 1444 1116 1460
rect 1131 1444 1144 1604
rect 1174 1500 1187 1604
rect 1232 1582 1233 1592
rect 1248 1582 1261 1592
rect 1232 1578 1261 1582
rect 1266 1578 1281 1604
rect 1232 1576 1281 1578
rect 1216 1568 1267 1576
rect 1216 1556 1241 1568
rect 1248 1556 1267 1568
rect 1216 1548 1267 1556
rect 1232 1540 1233 1548
rect 1248 1540 1261 1548
rect 1232 1532 1248 1540
rect 1229 1525 1248 1528
rect 1229 1516 1251 1525
rect 1202 1506 1251 1516
rect 1202 1500 1232 1506
rect 1251 1501 1256 1506
rect 1174 1484 1248 1500
rect 1266 1492 1281 1548
rect 1174 1482 1187 1484
rect 1202 1482 1236 1484
rect 1174 1466 1248 1482
rect 1158 1444 1159 1460
rect 1174 1444 1187 1466
rect 1202 1444 1232 1466
rect 1275 1444 1281 1492
rect 3494 1500 3507 1604
rect 3552 1582 3553 1592
rect 3568 1582 3581 1592
rect 3552 1578 3581 1582
rect 3586 1578 3616 1604
rect 3634 1590 3650 1592
rect 3722 1590 3775 1604
rect 3723 1588 3787 1590
rect 3830 1588 3845 1604
rect 3894 1601 3924 1604
rect 3894 1598 3930 1601
rect 3860 1590 3876 1592
rect 3634 1578 3649 1582
rect 3552 1576 3649 1578
rect 3677 1576 3845 1588
rect 3861 1578 3876 1582
rect 3894 1579 3933 1598
rect 3952 1592 3959 1593
rect 3958 1585 3959 1592
rect 3942 1582 3943 1585
rect 3958 1582 3971 1585
rect 3894 1578 3924 1579
rect 3933 1578 3939 1579
rect 3942 1578 3971 1582
rect 3861 1577 3971 1578
rect 3861 1576 3977 1577
rect 3536 1568 3587 1576
rect 3536 1556 3561 1568
rect 3568 1556 3587 1568
rect 3618 1568 3668 1576
rect 3618 1560 3634 1568
rect 3641 1566 3668 1568
rect 3677 1566 3898 1576
rect 3641 1556 3898 1566
rect 3927 1568 3977 1576
rect 3927 1559 3943 1568
rect 3536 1548 3587 1556
rect 3634 1548 3898 1556
rect 3924 1556 3943 1559
rect 3950 1556 3977 1568
rect 3924 1548 3977 1556
rect 3552 1540 3553 1548
rect 3568 1540 3581 1548
rect 3552 1532 3568 1540
rect 3549 1525 3568 1528
rect 3549 1516 3571 1525
rect 3522 1506 3571 1516
rect 3522 1500 3552 1506
rect 3571 1501 3576 1506
rect 3494 1484 3568 1500
rect 3586 1492 3616 1548
rect 3651 1538 3859 1548
rect 3894 1544 3939 1548
rect 3942 1547 3943 1548
rect 3958 1547 3971 1548
rect 3677 1508 3866 1538
rect 3692 1505 3866 1508
rect 3685 1502 3866 1505
rect 3494 1482 3507 1484
rect 3522 1482 3556 1484
rect 3494 1466 3568 1482
rect 3595 1478 3608 1492
rect 3623 1478 3639 1494
rect 3685 1489 3696 1502
rect 3494 1444 3507 1466
rect 3522 1444 3552 1466
rect 3595 1462 3657 1478
rect 3685 1471 3696 1487
rect 3701 1482 3711 1502
rect 3721 1482 3735 1502
rect 3738 1489 3747 1502
rect 3763 1489 3772 1502
rect 3701 1471 3735 1482
rect 3738 1471 3747 1487
rect 3763 1471 3772 1487
rect 3779 1482 3789 1502
rect 3799 1482 3813 1502
rect 3814 1489 3825 1502
rect 3779 1471 3813 1482
rect 3814 1471 3825 1487
rect 3871 1478 3887 1494
rect 3894 1492 3924 1544
rect 3958 1540 3959 1547
rect 3943 1532 3959 1540
rect 3930 1500 3943 1519
rect 3958 1500 3988 1516
rect 3930 1484 4004 1500
rect 3930 1482 3943 1484
rect 3958 1482 3992 1484
rect 3595 1460 3608 1462
rect 3623 1460 3657 1462
rect 3595 1444 3657 1460
rect 3701 1455 3717 1462
rect 3779 1455 3809 1466
rect 3857 1462 3903 1478
rect 3930 1466 4004 1482
rect 3857 1460 3891 1462
rect 3856 1444 3903 1460
rect 3930 1444 3943 1466
rect 3958 1444 3988 1466
rect 4015 1444 4016 1460
rect 4031 1444 4044 1604
rect 4074 1500 4087 1604
rect 4132 1582 4133 1592
rect 4148 1582 4161 1592
rect 4132 1578 4161 1582
rect 4166 1578 4196 1604
rect 4214 1590 4230 1592
rect 4302 1590 4355 1604
rect 4303 1588 4367 1590
rect 4410 1588 4425 1604
rect 4474 1601 4504 1604
rect 4474 1598 4510 1601
rect 4440 1590 4456 1592
rect 4214 1578 4229 1582
rect 4132 1576 4229 1578
rect 4257 1576 4425 1588
rect 4441 1578 4456 1582
rect 4474 1579 4513 1598
rect 4532 1592 4539 1593
rect 4538 1585 4539 1592
rect 4522 1582 4523 1585
rect 4538 1582 4551 1585
rect 4474 1578 4504 1579
rect 4513 1578 4519 1579
rect 4522 1578 4551 1582
rect 4441 1577 4551 1578
rect 4441 1576 4557 1577
rect 4116 1568 4167 1576
rect 4116 1556 4141 1568
rect 4148 1556 4167 1568
rect 4198 1568 4248 1576
rect 4198 1560 4214 1568
rect 4221 1566 4248 1568
rect 4257 1566 4478 1576
rect 4221 1556 4478 1566
rect 4507 1568 4557 1576
rect 4507 1559 4523 1568
rect 4116 1548 4167 1556
rect 4214 1548 4478 1556
rect 4504 1556 4523 1559
rect 4530 1556 4557 1568
rect 4504 1548 4557 1556
rect 4132 1540 4133 1548
rect 4148 1540 4161 1548
rect 4132 1532 4148 1540
rect 4129 1525 4148 1528
rect 4129 1516 4151 1525
rect 4102 1506 4151 1516
rect 4102 1500 4132 1506
rect 4151 1501 4156 1506
rect 4074 1484 4148 1500
rect 4166 1492 4196 1548
rect 4231 1538 4439 1548
rect 4474 1544 4519 1548
rect 4522 1547 4523 1548
rect 4538 1547 4551 1548
rect 4257 1508 4446 1538
rect 4272 1505 4446 1508
rect 4265 1502 4446 1505
rect 4074 1482 4087 1484
rect 4102 1482 4136 1484
rect 4074 1466 4148 1482
rect 4175 1478 4188 1492
rect 4203 1478 4219 1494
rect 4265 1489 4276 1502
rect 4058 1444 4059 1460
rect 4074 1444 4087 1466
rect 4102 1444 4132 1466
rect 4175 1462 4237 1478
rect 4265 1471 4276 1487
rect 4281 1482 4291 1502
rect 4301 1482 4315 1502
rect 4318 1489 4327 1502
rect 4343 1489 4352 1502
rect 4281 1471 4315 1482
rect 4318 1471 4327 1487
rect 4343 1471 4352 1487
rect 4359 1482 4369 1502
rect 4379 1482 4393 1502
rect 4394 1489 4405 1502
rect 4359 1471 4393 1482
rect 4394 1471 4405 1487
rect 4451 1478 4467 1494
rect 4474 1492 4504 1544
rect 4538 1540 4539 1547
rect 4523 1532 4539 1540
rect 4510 1500 4523 1519
rect 4538 1500 4568 1516
rect 4510 1484 4584 1500
rect 4510 1482 4523 1484
rect 4538 1482 4572 1484
rect 4175 1460 4188 1462
rect 4203 1460 4237 1462
rect 4175 1444 4237 1460
rect 4281 1455 4297 1462
rect 4359 1455 4389 1466
rect 4437 1462 4483 1478
rect 4510 1466 4584 1482
rect 4437 1460 4471 1462
rect 4436 1444 4483 1460
rect 4510 1444 4523 1466
rect 4538 1444 4568 1466
rect 4595 1444 4596 1460
rect 4611 1444 4624 1604
rect 4654 1500 4667 1604
rect 4712 1582 4713 1592
rect 4728 1582 4741 1592
rect 4712 1578 4741 1582
rect 4746 1578 4776 1604
rect 4794 1590 4810 1592
rect 4882 1590 4933 1604
rect 4883 1588 4947 1590
rect 4990 1588 5005 1604
rect 5054 1601 5084 1604
rect 5054 1598 5090 1601
rect 5020 1590 5036 1592
rect 4794 1578 4809 1582
rect 4712 1576 4809 1578
rect 4837 1576 5005 1588
rect 5021 1578 5036 1582
rect 5054 1579 5093 1598
rect 5112 1592 5119 1593
rect 5118 1585 5119 1592
rect 5102 1582 5103 1585
rect 5118 1582 5131 1585
rect 5054 1578 5084 1579
rect 5093 1578 5099 1579
rect 5102 1578 5131 1582
rect 5021 1577 5131 1578
rect 5021 1576 5137 1577
rect 4696 1568 4747 1576
rect 4696 1556 4721 1568
rect 4728 1556 4747 1568
rect 4778 1568 4828 1576
rect 4778 1560 4794 1568
rect 4801 1566 4828 1568
rect 4837 1566 5058 1576
rect 4801 1556 5058 1566
rect 5087 1568 5137 1576
rect 5087 1559 5103 1568
rect 4696 1548 4747 1556
rect 4794 1548 5058 1556
rect 5084 1556 5103 1559
rect 5110 1556 5137 1568
rect 5084 1548 5137 1556
rect 4712 1540 4713 1548
rect 4728 1540 4741 1548
rect 4712 1532 4728 1540
rect 4709 1525 4728 1528
rect 4709 1516 4731 1525
rect 4682 1506 4731 1516
rect 4682 1500 4712 1506
rect 4731 1501 4736 1506
rect 4654 1484 4728 1500
rect 4746 1492 4776 1548
rect 4811 1538 5019 1548
rect 5054 1544 5099 1548
rect 5102 1547 5103 1548
rect 5118 1547 5131 1548
rect 4837 1508 5026 1538
rect 4852 1505 5026 1508
rect 4845 1502 5026 1505
rect 4654 1482 4667 1484
rect 4682 1482 4716 1484
rect 4654 1466 4728 1482
rect 4755 1478 4768 1492
rect 4783 1478 4799 1494
rect 4845 1489 4856 1502
rect 4638 1444 4639 1460
rect 4654 1444 4667 1466
rect 4682 1444 4712 1466
rect 4755 1462 4817 1478
rect 4845 1471 4856 1487
rect 4861 1482 4871 1502
rect 4881 1482 4895 1502
rect 4898 1489 4907 1502
rect 4923 1489 4932 1502
rect 4861 1471 4895 1482
rect 4898 1471 4907 1487
rect 4923 1471 4932 1487
rect 4939 1482 4949 1502
rect 4959 1482 4973 1502
rect 4974 1489 4985 1502
rect 4939 1471 4973 1482
rect 4974 1471 4985 1487
rect 5031 1478 5047 1494
rect 5054 1492 5084 1544
rect 5118 1540 5119 1547
rect 5103 1532 5119 1540
rect 5090 1500 5103 1519
rect 5118 1500 5148 1516
rect 5090 1484 5164 1500
rect 5090 1482 5103 1484
rect 5118 1482 5152 1484
rect 4755 1460 4768 1462
rect 4783 1460 4817 1462
rect 4755 1444 4817 1460
rect 4861 1455 4877 1462
rect 4939 1455 4969 1466
rect 5017 1462 5063 1478
rect 5090 1466 5164 1482
rect 5017 1460 5051 1462
rect 5016 1444 5063 1460
rect 5090 1444 5103 1466
rect 5118 1444 5148 1466
rect 5175 1444 5176 1460
rect 5191 1444 5204 1604
rect 5234 1500 5247 1604
rect 5292 1582 5293 1592
rect 5308 1582 5321 1592
rect 5292 1578 5321 1582
rect 5326 1578 5356 1604
rect 5374 1590 5390 1592
rect 5462 1590 5513 1604
rect 5463 1588 5527 1590
rect 5570 1588 5585 1604
rect 5634 1601 5664 1604
rect 5634 1598 5670 1601
rect 5600 1590 5616 1592
rect 5374 1578 5389 1582
rect 5292 1576 5389 1578
rect 5417 1576 5585 1588
rect 5601 1578 5616 1582
rect 5634 1579 5673 1598
rect 5692 1592 5699 1593
rect 5698 1585 5699 1592
rect 5682 1582 5683 1585
rect 5698 1582 5711 1585
rect 5634 1578 5664 1579
rect 5673 1578 5679 1579
rect 5682 1578 5711 1582
rect 5601 1577 5711 1578
rect 5601 1576 5717 1577
rect 5276 1568 5327 1576
rect 5276 1556 5301 1568
rect 5308 1556 5327 1568
rect 5358 1568 5408 1576
rect 5358 1560 5374 1568
rect 5381 1566 5408 1568
rect 5417 1566 5638 1576
rect 5381 1556 5638 1566
rect 5667 1568 5717 1576
rect 5667 1559 5683 1568
rect 5276 1548 5327 1556
rect 5374 1548 5638 1556
rect 5664 1556 5683 1559
rect 5690 1556 5717 1568
rect 5664 1548 5717 1556
rect 5292 1540 5293 1548
rect 5308 1540 5321 1548
rect 5292 1532 5308 1540
rect 5289 1525 5308 1528
rect 5289 1516 5311 1525
rect 5262 1506 5311 1516
rect 5262 1500 5292 1506
rect 5311 1501 5316 1506
rect 5234 1484 5308 1500
rect 5326 1492 5356 1548
rect 5391 1538 5599 1548
rect 5634 1544 5679 1548
rect 5682 1547 5683 1548
rect 5698 1547 5711 1548
rect 5417 1508 5606 1538
rect 5432 1505 5606 1508
rect 5425 1502 5606 1505
rect 5234 1482 5247 1484
rect 5262 1482 5296 1484
rect 5234 1466 5308 1482
rect 5335 1478 5348 1492
rect 5363 1478 5379 1494
rect 5425 1489 5436 1502
rect 5218 1444 5219 1460
rect 5234 1444 5247 1466
rect 5262 1444 5292 1466
rect 5335 1462 5397 1478
rect 5425 1471 5436 1487
rect 5441 1482 5451 1502
rect 5461 1482 5475 1502
rect 5478 1489 5487 1502
rect 5503 1489 5512 1502
rect 5441 1471 5475 1482
rect 5478 1471 5487 1487
rect 5503 1471 5512 1487
rect 5519 1482 5529 1502
rect 5539 1482 5553 1502
rect 5554 1489 5565 1502
rect 5519 1471 5553 1482
rect 5554 1471 5565 1487
rect 5611 1478 5627 1494
rect 5634 1492 5664 1544
rect 5698 1540 5699 1547
rect 5683 1532 5699 1540
rect 5670 1500 5683 1519
rect 5698 1500 5728 1516
rect 5670 1484 5744 1500
rect 5670 1482 5683 1484
rect 5698 1482 5732 1484
rect 5335 1460 5348 1462
rect 5363 1460 5397 1462
rect 5335 1444 5397 1460
rect 5441 1455 5457 1462
rect 5519 1455 5549 1466
rect 5597 1462 5643 1478
rect 5670 1466 5744 1482
rect 5597 1460 5631 1462
rect 5596 1444 5643 1460
rect 5670 1444 5683 1466
rect 5698 1444 5728 1466
rect 5755 1444 5756 1460
rect 5771 1444 5784 1604
rect 5814 1500 5827 1604
rect 5872 1582 5873 1592
rect 5888 1582 5901 1592
rect 5872 1578 5901 1582
rect 5906 1578 5936 1604
rect 5954 1590 5970 1592
rect 6042 1590 6093 1604
rect 6043 1588 6107 1590
rect 6150 1588 6165 1604
rect 6214 1601 6244 1604
rect 6214 1598 6250 1601
rect 6180 1590 6196 1592
rect 5954 1578 5969 1582
rect 5872 1576 5969 1578
rect 5997 1576 6165 1588
rect 6181 1578 6196 1582
rect 6214 1579 6253 1598
rect 6272 1592 6279 1593
rect 6278 1585 6279 1592
rect 6262 1582 6263 1585
rect 6278 1582 6291 1585
rect 6214 1578 6244 1579
rect 6253 1578 6259 1579
rect 6262 1578 6291 1582
rect 6181 1577 6291 1578
rect 6181 1576 6297 1577
rect 5856 1568 5907 1576
rect 5856 1556 5881 1568
rect 5888 1556 5907 1568
rect 5938 1568 5988 1576
rect 5938 1560 5954 1568
rect 5961 1566 5988 1568
rect 5997 1566 6218 1576
rect 5961 1556 6218 1566
rect 6247 1568 6297 1576
rect 6247 1559 6263 1568
rect 5856 1548 5907 1556
rect 5954 1548 6218 1556
rect 6244 1556 6263 1559
rect 6270 1556 6297 1568
rect 6244 1548 6297 1556
rect 5872 1540 5873 1548
rect 5888 1540 5901 1548
rect 5872 1532 5888 1540
rect 5869 1525 5888 1528
rect 5869 1516 5891 1525
rect 5842 1506 5891 1516
rect 5842 1500 5872 1506
rect 5891 1501 5896 1506
rect 5814 1484 5888 1500
rect 5906 1492 5936 1548
rect 5971 1538 6179 1548
rect 6214 1544 6259 1548
rect 6262 1547 6263 1548
rect 6278 1547 6291 1548
rect 5997 1508 6186 1538
rect 6012 1505 6186 1508
rect 6005 1502 6186 1505
rect 5814 1482 5827 1484
rect 5842 1482 5876 1484
rect 5814 1466 5888 1482
rect 5915 1478 5928 1492
rect 5943 1478 5959 1494
rect 6005 1489 6016 1502
rect 5798 1444 5799 1460
rect 5814 1444 5827 1466
rect 5842 1444 5872 1466
rect 5915 1462 5977 1478
rect 6005 1471 6016 1487
rect 6021 1482 6031 1502
rect 6041 1482 6055 1502
rect 6058 1489 6067 1502
rect 6083 1489 6092 1502
rect 6021 1471 6055 1482
rect 6058 1471 6067 1487
rect 6083 1471 6092 1487
rect 6099 1482 6109 1502
rect 6119 1482 6133 1502
rect 6134 1489 6145 1502
rect 6099 1471 6133 1482
rect 6134 1471 6145 1487
rect 6191 1478 6207 1494
rect 6214 1492 6244 1544
rect 6278 1540 6279 1547
rect 6263 1532 6279 1540
rect 6250 1500 6263 1519
rect 6278 1500 6308 1516
rect 6250 1484 6324 1500
rect 6250 1482 6263 1484
rect 6278 1482 6312 1484
rect 5915 1460 5928 1462
rect 5943 1460 5977 1462
rect 5915 1444 5977 1460
rect 6021 1455 6037 1462
rect 6099 1455 6129 1466
rect 6177 1462 6223 1478
rect 6250 1466 6324 1482
rect 6177 1460 6211 1462
rect 6176 1444 6223 1460
rect 6250 1444 6263 1466
rect 6278 1444 6308 1466
rect 6335 1444 6336 1460
rect 6351 1444 6364 1604
rect 6394 1500 6407 1604
rect 6452 1582 6453 1592
rect 6468 1582 6481 1592
rect 6452 1578 6481 1582
rect 6486 1578 6516 1604
rect 6534 1590 6550 1592
rect 6622 1590 6673 1604
rect 6623 1588 6687 1590
rect 6730 1588 6745 1604
rect 6794 1601 6824 1604
rect 6794 1598 6830 1601
rect 6760 1590 6776 1592
rect 6534 1578 6549 1582
rect 6452 1576 6549 1578
rect 6577 1576 6745 1588
rect 6761 1578 6776 1582
rect 6794 1579 6833 1598
rect 6852 1592 6859 1593
rect 6858 1585 6859 1592
rect 6842 1582 6843 1585
rect 6858 1582 6871 1585
rect 6794 1578 6824 1579
rect 6833 1578 6839 1579
rect 6842 1578 6871 1582
rect 6761 1577 6871 1578
rect 6761 1576 6877 1577
rect 6436 1568 6487 1576
rect 6436 1556 6461 1568
rect 6468 1556 6487 1568
rect 6518 1568 6568 1576
rect 6518 1560 6534 1568
rect 6541 1566 6568 1568
rect 6577 1566 6798 1576
rect 6541 1556 6798 1566
rect 6827 1568 6877 1576
rect 6827 1559 6843 1568
rect 6436 1548 6487 1556
rect 6534 1548 6798 1556
rect 6824 1556 6843 1559
rect 6850 1556 6877 1568
rect 6824 1548 6877 1556
rect 6452 1540 6453 1548
rect 6468 1540 6481 1548
rect 6452 1532 6468 1540
rect 6449 1525 6468 1528
rect 6449 1516 6471 1525
rect 6422 1506 6471 1516
rect 6422 1500 6452 1506
rect 6471 1501 6476 1506
rect 6394 1484 6468 1500
rect 6486 1492 6516 1548
rect 6551 1538 6759 1548
rect 6794 1544 6839 1548
rect 6842 1547 6843 1548
rect 6858 1547 6871 1548
rect 6577 1508 6766 1538
rect 6592 1505 6766 1508
rect 6585 1502 6766 1505
rect 6394 1482 6407 1484
rect 6422 1482 6456 1484
rect 6394 1466 6468 1482
rect 6495 1478 6508 1492
rect 6523 1478 6539 1494
rect 6585 1489 6596 1502
rect 6378 1444 6379 1460
rect 6394 1444 6407 1466
rect 6422 1444 6452 1466
rect 6495 1462 6557 1478
rect 6585 1471 6596 1487
rect 6601 1482 6611 1502
rect 6621 1482 6635 1502
rect 6638 1489 6647 1502
rect 6663 1489 6672 1502
rect 6601 1471 6635 1482
rect 6638 1471 6647 1487
rect 6663 1471 6672 1487
rect 6679 1482 6689 1502
rect 6699 1482 6713 1502
rect 6714 1489 6725 1502
rect 6679 1471 6713 1482
rect 6714 1471 6725 1487
rect 6771 1478 6787 1494
rect 6794 1492 6824 1544
rect 6858 1540 6859 1547
rect 6843 1532 6859 1540
rect 6830 1500 6843 1519
rect 6858 1500 6888 1516
rect 6830 1484 6904 1500
rect 6830 1482 6843 1484
rect 6858 1482 6892 1484
rect 6495 1460 6508 1462
rect 6523 1460 6557 1462
rect 6495 1444 6557 1460
rect 6601 1455 6617 1462
rect 6679 1455 6709 1466
rect 6757 1462 6803 1478
rect 6830 1466 6904 1482
rect 6757 1460 6791 1462
rect 6756 1444 6803 1460
rect 6830 1444 6843 1466
rect 6858 1444 6888 1466
rect 6915 1444 6916 1460
rect 6931 1444 6944 1604
rect -8 1436 33 1444
rect -8 1410 7 1436
rect 14 1410 33 1436
rect 97 1432 159 1444
rect 171 1432 246 1444
rect 304 1432 379 1444
rect 391 1432 422 1444
rect 428 1432 463 1444
rect 97 1430 259 1432
rect -8 1402 33 1410
rect 115 1406 128 1430
rect 143 1428 158 1430
rect -2 1392 -1 1402
rect 14 1392 27 1402
rect 42 1392 72 1406
rect 115 1392 158 1406
rect 182 1403 189 1410
rect 192 1406 259 1430
rect 291 1430 463 1432
rect 261 1408 289 1412
rect 291 1408 371 1430
rect 392 1428 407 1430
rect 261 1406 371 1408
rect 192 1402 371 1406
rect 165 1392 195 1402
rect 197 1392 350 1402
rect 358 1392 388 1402
rect 392 1392 422 1406
rect 450 1392 463 1430
rect 535 1436 570 1444
rect 535 1410 536 1436
rect 543 1410 570 1436
rect 478 1392 508 1406
rect 535 1402 570 1410
rect 572 1436 613 1444
rect 572 1410 587 1436
rect 594 1410 613 1436
rect 677 1432 739 1444
rect 751 1432 826 1444
rect 884 1432 959 1444
rect 971 1432 1002 1444
rect 1008 1432 1043 1444
rect 677 1430 839 1432
rect 572 1402 613 1410
rect 695 1406 708 1430
rect 723 1428 738 1430
rect 535 1392 536 1402
rect 551 1392 564 1402
rect 578 1392 579 1402
rect 594 1392 607 1402
rect 622 1392 652 1406
rect 695 1392 738 1406
rect 762 1403 769 1410
rect 772 1406 839 1430
rect 871 1430 1043 1432
rect 841 1408 869 1412
rect 871 1408 951 1430
rect 972 1428 987 1430
rect 841 1406 951 1408
rect 772 1402 951 1406
rect 745 1392 775 1402
rect 777 1392 930 1402
rect 938 1392 968 1402
rect 972 1392 1002 1406
rect 1030 1392 1043 1430
rect 1115 1436 1150 1444
rect 1115 1410 1116 1436
rect 1123 1410 1150 1436
rect 1058 1392 1088 1406
rect 1115 1402 1150 1410
rect 1152 1436 1193 1444
rect 1152 1410 1167 1436
rect 1174 1410 1193 1436
rect 1257 1430 1281 1444
rect 1152 1402 1193 1410
rect 1115 1392 1116 1402
rect 1131 1392 1144 1402
rect 1158 1392 1159 1402
rect 1174 1392 1187 1402
rect 1202 1392 1232 1406
rect 1275 1392 1281 1430
rect 3481 1436 3513 1444
rect 3481 1410 3487 1436
rect 3494 1410 3513 1436
rect 3577 1432 3639 1444
rect 3651 1432 3726 1444
rect 3784 1432 3859 1444
rect 3871 1432 3902 1444
rect 3908 1432 3943 1444
rect 3577 1430 3739 1432
rect 3481 1402 3513 1410
rect 3595 1406 3608 1430
rect 3623 1428 3638 1430
rect 3494 1392 3507 1402
rect 3522 1392 3552 1406
rect 3595 1392 3638 1406
rect 3662 1403 3669 1410
rect 3672 1406 3739 1430
rect 3771 1430 3943 1432
rect 3741 1408 3769 1412
rect 3771 1408 3851 1430
rect 3872 1428 3887 1430
rect 3741 1406 3851 1408
rect 3672 1402 3851 1406
rect 3645 1392 3675 1402
rect 3677 1392 3830 1402
rect 3838 1392 3868 1402
rect 3872 1392 3902 1406
rect 3930 1392 3943 1430
rect 4015 1436 4050 1444
rect 4015 1410 4016 1436
rect 4023 1410 4050 1436
rect 3958 1392 3988 1406
rect 4015 1402 4050 1410
rect 4052 1436 4093 1444
rect 4052 1410 4067 1436
rect 4074 1410 4093 1436
rect 4157 1432 4219 1444
rect 4231 1432 4306 1444
rect 4364 1432 4439 1444
rect 4451 1432 4482 1444
rect 4488 1432 4523 1444
rect 4157 1430 4319 1432
rect 4052 1402 4093 1410
rect 4175 1406 4188 1430
rect 4203 1428 4218 1430
rect 4015 1392 4016 1402
rect 4031 1392 4044 1402
rect 4058 1392 4059 1402
rect 4074 1392 4087 1402
rect 4102 1392 4132 1406
rect 4175 1392 4218 1406
rect 4242 1403 4249 1410
rect 4252 1406 4319 1430
rect 4351 1430 4523 1432
rect 4321 1408 4349 1412
rect 4351 1408 4431 1430
rect 4452 1428 4467 1430
rect 4321 1406 4431 1408
rect 4252 1402 4431 1406
rect 4225 1392 4255 1402
rect 4257 1392 4410 1402
rect 4418 1392 4448 1402
rect 4452 1392 4482 1406
rect 4510 1392 4523 1430
rect 4595 1436 4630 1444
rect 4595 1410 4596 1436
rect 4603 1410 4630 1436
rect 4538 1392 4568 1406
rect 4595 1402 4630 1410
rect 4632 1436 4673 1444
rect 4632 1410 4647 1436
rect 4654 1410 4673 1436
rect 4737 1432 4799 1444
rect 4811 1432 4886 1444
rect 4944 1432 5019 1444
rect 5031 1432 5062 1444
rect 5068 1432 5103 1444
rect 4737 1430 4899 1432
rect 4632 1402 4673 1410
rect 4755 1406 4768 1430
rect 4783 1428 4798 1430
rect 4832 1412 4899 1430
rect 4931 1430 5103 1432
rect 4931 1412 5011 1430
rect 5032 1428 5047 1430
rect 4595 1392 4596 1402
rect 4611 1392 4624 1402
rect 4638 1392 4639 1402
rect 4654 1392 4667 1402
rect 4682 1392 4712 1406
rect 4755 1392 4798 1406
rect 4822 1403 4829 1410
rect 4832 1402 5011 1412
rect 4805 1392 4835 1402
rect 4837 1392 4990 1402
rect 4998 1392 5028 1402
rect 5032 1392 5062 1406
rect 5090 1392 5103 1430
rect 5175 1436 5210 1444
rect 5175 1410 5176 1436
rect 5183 1410 5210 1436
rect 5118 1392 5148 1406
rect 5175 1402 5210 1410
rect 5212 1436 5253 1444
rect 5212 1410 5227 1436
rect 5234 1410 5253 1436
rect 5317 1432 5379 1444
rect 5391 1432 5466 1444
rect 5524 1432 5599 1444
rect 5611 1432 5642 1444
rect 5648 1432 5683 1444
rect 5317 1430 5479 1432
rect 5212 1402 5253 1410
rect 5335 1406 5348 1430
rect 5363 1428 5378 1430
rect 5412 1412 5479 1430
rect 5511 1430 5683 1432
rect 5511 1412 5591 1430
rect 5612 1428 5627 1430
rect 5175 1392 5176 1402
rect 5191 1392 5204 1402
rect 5218 1392 5219 1402
rect 5234 1392 5247 1402
rect 5262 1392 5292 1406
rect 5335 1392 5378 1406
rect 5402 1403 5409 1410
rect 5412 1402 5591 1412
rect 5385 1392 5415 1402
rect 5417 1392 5570 1402
rect 5578 1392 5608 1402
rect 5612 1392 5642 1406
rect 5670 1392 5683 1430
rect 5755 1436 5790 1444
rect 5755 1410 5756 1436
rect 5763 1410 5790 1436
rect 5698 1392 5728 1406
rect 5755 1402 5790 1410
rect 5792 1436 5833 1444
rect 5792 1410 5807 1436
rect 5814 1410 5833 1436
rect 5897 1432 5959 1444
rect 5971 1432 6046 1444
rect 6104 1432 6179 1444
rect 6191 1432 6222 1444
rect 6228 1432 6263 1444
rect 5897 1430 6059 1432
rect 5792 1402 5833 1410
rect 5915 1406 5928 1430
rect 5943 1428 5958 1430
rect 5992 1412 6059 1430
rect 6091 1430 6263 1432
rect 6091 1412 6171 1430
rect 6192 1428 6207 1430
rect 5755 1392 5756 1402
rect 5771 1392 5784 1402
rect 5798 1392 5799 1402
rect 5814 1392 5827 1402
rect 5842 1392 5872 1406
rect 5915 1392 5958 1406
rect 5982 1403 5989 1410
rect 5992 1402 6171 1412
rect 5965 1392 5995 1402
rect 5997 1392 6150 1402
rect 6158 1392 6188 1402
rect 6192 1392 6222 1406
rect 6250 1392 6263 1430
rect 6335 1436 6370 1444
rect 6335 1410 6336 1436
rect 6343 1410 6370 1436
rect 6278 1392 6308 1406
rect 6335 1402 6370 1410
rect 6372 1436 6413 1444
rect 6372 1410 6387 1436
rect 6394 1410 6413 1436
rect 6477 1432 6539 1444
rect 6551 1432 6626 1444
rect 6684 1432 6759 1444
rect 6771 1432 6802 1444
rect 6808 1432 6843 1444
rect 6477 1430 6639 1432
rect 6372 1402 6413 1410
rect 6495 1406 6508 1430
rect 6523 1428 6538 1430
rect 6572 1412 6639 1430
rect 6671 1430 6843 1432
rect 6671 1412 6751 1430
rect 6772 1428 6787 1430
rect 6335 1392 6336 1402
rect 6351 1392 6364 1402
rect 6378 1392 6379 1402
rect 6394 1392 6407 1402
rect 6422 1392 6452 1406
rect 6495 1392 6538 1406
rect 6562 1403 6569 1410
rect 6572 1402 6751 1412
rect 6545 1392 6575 1402
rect 6577 1392 6730 1402
rect 6738 1392 6768 1402
rect 6772 1392 6802 1406
rect 6830 1392 6843 1430
rect 6915 1436 6950 1444
rect 6915 1410 6916 1436
rect 6923 1410 6950 1436
rect 6858 1392 6888 1406
rect 6915 1402 6950 1410
rect 6915 1392 6916 1402
rect 6931 1392 6944 1402
rect -2 1386 1281 1392
rect -1 1378 1281 1386
rect 3481 1378 6944 1392
rect 14 1348 27 1378
rect 42 1360 72 1378
rect 115 1364 129 1378
rect 165 1364 385 1378
rect 116 1362 129 1364
rect 82 1350 97 1362
rect 79 1348 101 1350
rect 106 1348 136 1362
rect 197 1360 350 1364
rect 179 1348 371 1360
rect 414 1348 444 1362
rect 450 1348 463 1378
rect 478 1360 508 1378
rect 551 1348 564 1378
rect 594 1348 607 1378
rect 622 1360 652 1378
rect 695 1364 709 1378
rect 745 1364 965 1378
rect 696 1362 709 1364
rect 662 1350 677 1362
rect 659 1348 681 1350
rect 686 1348 716 1362
rect 777 1360 930 1364
rect 759 1348 951 1360
rect 994 1348 1024 1362
rect 1030 1348 1043 1378
rect 1058 1360 1088 1378
rect 1131 1348 1144 1378
rect 1174 1348 1187 1378
rect 1202 1360 1232 1378
rect 1275 1364 1281 1378
rect 1276 1362 1281 1364
rect 1242 1350 1257 1362
rect 1239 1348 1261 1350
rect 1266 1348 1281 1362
rect 3494 1348 3507 1378
rect 3522 1360 3552 1378
rect 3595 1364 3609 1378
rect 3645 1364 3865 1378
rect 3596 1362 3609 1364
rect 3562 1350 3577 1362
rect 3559 1348 3581 1350
rect 3586 1348 3616 1362
rect 3677 1360 3830 1364
rect 3659 1348 3851 1360
rect 3894 1348 3924 1362
rect 3930 1348 3943 1378
rect 3958 1360 3988 1378
rect 4031 1348 4044 1378
rect 4074 1348 4087 1378
rect 4102 1360 4132 1378
rect 4175 1364 4189 1378
rect 4225 1364 4445 1378
rect 4176 1362 4189 1364
rect 4142 1350 4157 1362
rect 4139 1348 4161 1350
rect 4166 1348 4196 1362
rect 4257 1360 4410 1364
rect 4239 1348 4431 1360
rect 4474 1348 4504 1362
rect 4510 1348 4523 1378
rect 4538 1360 4568 1378
rect 4611 1348 4624 1378
rect 4654 1348 4667 1378
rect 4682 1360 4712 1378
rect 4755 1364 4769 1378
rect 4805 1364 5025 1378
rect 4756 1362 4769 1364
rect 4722 1350 4737 1362
rect 4719 1348 4741 1350
rect 4746 1348 4776 1362
rect 4837 1360 4990 1364
rect 4819 1348 5011 1360
rect 5054 1348 5084 1362
rect 5090 1348 5103 1378
rect 5118 1360 5148 1378
rect 5191 1348 5204 1378
rect 5234 1348 5247 1378
rect 5262 1360 5292 1378
rect 5335 1364 5349 1378
rect 5385 1364 5605 1378
rect 5336 1362 5349 1364
rect 5302 1350 5317 1362
rect 5299 1348 5321 1350
rect 5326 1348 5356 1362
rect 5417 1360 5570 1364
rect 5399 1348 5591 1360
rect 5634 1348 5664 1362
rect 5670 1348 5683 1378
rect 5698 1360 5728 1378
rect 5771 1348 5784 1378
rect 5814 1348 5827 1378
rect 5842 1360 5872 1378
rect 5915 1364 5929 1378
rect 5965 1364 6185 1378
rect 5916 1362 5929 1364
rect 5882 1350 5897 1362
rect 5879 1348 5901 1350
rect 5906 1348 5936 1362
rect 5997 1360 6150 1364
rect 5979 1348 6171 1360
rect 6214 1348 6244 1362
rect 6250 1348 6263 1378
rect 6278 1360 6308 1378
rect 6351 1348 6364 1378
rect 6394 1348 6407 1378
rect 6422 1360 6452 1378
rect 6495 1364 6509 1378
rect 6545 1364 6765 1378
rect 6496 1362 6509 1364
rect 6462 1350 6477 1362
rect 6459 1348 6481 1350
rect 6486 1348 6516 1362
rect 6577 1360 6730 1364
rect 6559 1348 6751 1360
rect 6794 1348 6824 1362
rect 6830 1348 6843 1378
rect 6858 1360 6888 1378
rect 6931 1348 6944 1378
rect -1 1334 1281 1348
rect 3481 1334 6944 1348
rect 14 1230 27 1334
rect 72 1312 73 1322
rect 88 1312 101 1322
rect 72 1308 101 1312
rect 106 1308 136 1334
rect 154 1320 170 1322
rect 242 1320 295 1334
rect 243 1318 307 1320
rect 350 1318 365 1334
rect 414 1331 444 1334
rect 414 1328 450 1331
rect 380 1320 396 1322
rect 154 1308 169 1312
rect 72 1306 169 1308
rect 197 1306 365 1318
rect 381 1308 396 1312
rect 414 1309 453 1328
rect 472 1322 479 1323
rect 478 1315 479 1322
rect 462 1312 463 1315
rect 478 1312 491 1315
rect 414 1308 444 1309
rect 453 1308 459 1309
rect 462 1308 491 1312
rect 381 1307 491 1308
rect 381 1306 497 1307
rect 56 1298 107 1306
rect 56 1286 81 1298
rect 88 1286 107 1298
rect 138 1298 188 1306
rect 138 1290 154 1298
rect 161 1296 188 1298
rect 197 1296 418 1306
rect 161 1286 418 1296
rect 447 1298 497 1306
rect 447 1289 463 1298
rect 56 1278 107 1286
rect 154 1278 418 1286
rect 444 1286 463 1289
rect 470 1286 497 1298
rect 444 1278 497 1286
rect 72 1270 73 1278
rect 88 1270 101 1278
rect 72 1262 88 1270
rect 69 1255 88 1258
rect 69 1246 91 1255
rect 42 1236 91 1246
rect 42 1230 72 1236
rect 91 1231 96 1236
rect 14 1214 88 1230
rect 106 1222 136 1278
rect 171 1268 379 1278
rect 414 1274 459 1278
rect 462 1277 463 1278
rect 478 1277 491 1278
rect 197 1238 386 1268
rect 212 1235 386 1238
rect 205 1232 386 1235
rect 14 1212 27 1214
rect 42 1212 76 1214
rect 14 1196 88 1212
rect 115 1208 128 1222
rect 143 1208 159 1224
rect 205 1219 216 1232
rect -2 1174 -1 1190
rect 14 1174 27 1196
rect 42 1174 72 1196
rect 115 1192 177 1208
rect 205 1201 216 1217
rect 221 1212 231 1232
rect 241 1212 255 1232
rect 258 1219 267 1232
rect 283 1219 292 1232
rect 221 1201 255 1212
rect 258 1201 267 1217
rect 283 1201 292 1217
rect 299 1212 309 1232
rect 319 1212 333 1232
rect 334 1219 345 1232
rect 299 1201 333 1212
rect 334 1201 345 1217
rect 391 1208 407 1224
rect 414 1222 444 1274
rect 478 1270 479 1277
rect 463 1262 479 1270
rect 450 1230 463 1249
rect 478 1230 508 1246
rect 450 1214 524 1230
rect 450 1212 463 1214
rect 478 1212 512 1214
rect 115 1190 128 1192
rect 143 1190 177 1192
rect 115 1174 177 1190
rect 221 1185 237 1192
rect 299 1185 329 1196
rect 377 1192 423 1208
rect 450 1196 524 1212
rect 377 1190 411 1192
rect 376 1174 423 1190
rect 450 1174 463 1196
rect 478 1174 508 1196
rect 535 1174 536 1190
rect 551 1174 564 1334
rect 594 1230 607 1334
rect 652 1312 653 1322
rect 668 1312 681 1322
rect 652 1308 681 1312
rect 686 1308 716 1334
rect 734 1320 750 1322
rect 822 1320 875 1334
rect 823 1318 887 1320
rect 930 1318 945 1334
rect 994 1331 1024 1334
rect 994 1328 1030 1331
rect 960 1320 976 1322
rect 734 1308 749 1312
rect 652 1306 749 1308
rect 777 1306 945 1318
rect 961 1308 976 1312
rect 994 1309 1033 1328
rect 1052 1322 1059 1323
rect 1058 1315 1059 1322
rect 1042 1312 1043 1315
rect 1058 1312 1071 1315
rect 994 1308 1024 1309
rect 1033 1308 1039 1309
rect 1042 1308 1071 1312
rect 961 1307 1071 1308
rect 961 1306 1077 1307
rect 636 1298 687 1306
rect 636 1286 661 1298
rect 668 1286 687 1298
rect 718 1298 768 1306
rect 718 1290 734 1298
rect 741 1296 768 1298
rect 777 1296 998 1306
rect 741 1286 998 1296
rect 1027 1298 1077 1306
rect 1027 1289 1043 1298
rect 636 1278 687 1286
rect 734 1278 998 1286
rect 1024 1286 1043 1289
rect 1050 1286 1077 1298
rect 1024 1278 1077 1286
rect 652 1270 653 1278
rect 668 1270 681 1278
rect 652 1262 668 1270
rect 649 1255 668 1258
rect 649 1246 671 1255
rect 622 1236 671 1246
rect 622 1230 652 1236
rect 671 1231 676 1236
rect 594 1214 668 1230
rect 686 1222 716 1278
rect 751 1268 959 1278
rect 994 1274 1039 1278
rect 1042 1277 1043 1278
rect 1058 1277 1071 1278
rect 777 1238 966 1268
rect 792 1235 966 1238
rect 785 1232 966 1235
rect 594 1212 607 1214
rect 622 1212 656 1214
rect 594 1196 668 1212
rect 695 1208 708 1222
rect 723 1208 739 1224
rect 785 1219 796 1232
rect 578 1174 579 1190
rect 594 1174 607 1196
rect 622 1174 652 1196
rect 695 1192 757 1208
rect 785 1201 796 1217
rect 801 1212 811 1232
rect 821 1212 835 1232
rect 838 1219 847 1232
rect 863 1219 872 1232
rect 801 1201 835 1212
rect 838 1201 847 1217
rect 863 1201 872 1217
rect 879 1212 889 1232
rect 899 1212 913 1232
rect 914 1219 925 1232
rect 879 1201 913 1212
rect 914 1201 925 1217
rect 971 1208 987 1224
rect 994 1222 1024 1274
rect 1058 1270 1059 1277
rect 1043 1262 1059 1270
rect 1030 1230 1043 1249
rect 1058 1230 1088 1246
rect 1030 1214 1104 1230
rect 1030 1212 1043 1214
rect 1058 1212 1092 1214
rect 695 1190 708 1192
rect 723 1190 757 1192
rect 695 1174 757 1190
rect 801 1185 817 1192
rect 879 1185 909 1196
rect 957 1192 1003 1208
rect 1030 1196 1104 1212
rect 957 1190 991 1192
rect 956 1174 1003 1190
rect 1030 1174 1043 1196
rect 1058 1174 1088 1196
rect 1115 1174 1116 1190
rect 1131 1174 1144 1334
rect 1174 1230 1187 1334
rect 1232 1312 1233 1322
rect 1248 1312 1261 1322
rect 1232 1308 1261 1312
rect 1266 1308 1281 1334
rect 1232 1306 1281 1308
rect 1216 1298 1267 1306
rect 1216 1286 1241 1298
rect 1248 1286 1267 1298
rect 1216 1278 1267 1286
rect 1232 1270 1233 1278
rect 1248 1270 1261 1278
rect 1232 1262 1248 1270
rect 1229 1255 1248 1258
rect 1229 1246 1251 1255
rect 1202 1236 1251 1246
rect 1202 1230 1232 1236
rect 1251 1231 1256 1236
rect 1174 1214 1248 1230
rect 1266 1222 1281 1278
rect 1174 1212 1187 1214
rect 1202 1212 1236 1214
rect 1174 1196 1248 1212
rect 1158 1174 1159 1190
rect 1174 1174 1187 1196
rect 1202 1174 1232 1196
rect 1275 1174 1281 1222
rect 3494 1230 3507 1334
rect 3552 1312 3553 1322
rect 3568 1312 3581 1322
rect 3552 1308 3581 1312
rect 3586 1308 3616 1334
rect 3634 1320 3650 1322
rect 3722 1320 3775 1334
rect 3723 1318 3787 1320
rect 3830 1318 3845 1334
rect 3894 1331 3924 1334
rect 3894 1328 3930 1331
rect 3860 1320 3876 1322
rect 3634 1308 3649 1312
rect 3552 1306 3649 1308
rect 3677 1306 3845 1318
rect 3861 1308 3876 1312
rect 3894 1309 3933 1328
rect 3952 1322 3959 1323
rect 3958 1315 3959 1322
rect 3942 1312 3943 1315
rect 3958 1312 3971 1315
rect 3894 1308 3924 1309
rect 3933 1308 3939 1309
rect 3942 1308 3971 1312
rect 3861 1307 3971 1308
rect 3861 1306 3977 1307
rect 3536 1298 3587 1306
rect 3536 1286 3561 1298
rect 3568 1286 3587 1298
rect 3618 1298 3668 1306
rect 3618 1290 3634 1298
rect 3641 1296 3668 1298
rect 3677 1296 3898 1306
rect 3641 1286 3898 1296
rect 3927 1298 3977 1306
rect 3927 1289 3943 1298
rect 3536 1278 3587 1286
rect 3634 1278 3898 1286
rect 3924 1286 3943 1289
rect 3950 1286 3977 1298
rect 3924 1278 3977 1286
rect 3552 1270 3553 1278
rect 3568 1270 3581 1278
rect 3552 1262 3568 1270
rect 3549 1255 3568 1258
rect 3549 1246 3571 1255
rect 3522 1236 3571 1246
rect 3522 1230 3552 1236
rect 3571 1231 3576 1236
rect 3494 1214 3568 1230
rect 3586 1222 3616 1278
rect 3651 1268 3859 1278
rect 3894 1274 3939 1278
rect 3942 1277 3943 1278
rect 3958 1277 3971 1278
rect 3677 1238 3866 1268
rect 3692 1235 3866 1238
rect 3685 1232 3866 1235
rect 3494 1212 3507 1214
rect 3522 1212 3556 1214
rect 3494 1196 3568 1212
rect 3595 1208 3608 1222
rect 3623 1208 3639 1224
rect 3685 1219 3696 1232
rect 3494 1174 3507 1196
rect 3522 1174 3552 1196
rect 3595 1192 3657 1208
rect 3685 1201 3696 1217
rect 3701 1212 3711 1232
rect 3721 1212 3735 1232
rect 3738 1219 3747 1232
rect 3763 1219 3772 1232
rect 3701 1201 3735 1212
rect 3738 1201 3747 1217
rect 3763 1201 3772 1217
rect 3779 1212 3789 1232
rect 3799 1212 3813 1232
rect 3814 1219 3825 1232
rect 3779 1201 3813 1212
rect 3814 1201 3825 1217
rect 3871 1208 3887 1224
rect 3894 1222 3924 1274
rect 3958 1270 3959 1277
rect 3943 1262 3959 1270
rect 3930 1230 3943 1249
rect 3958 1230 3988 1246
rect 3930 1214 4004 1230
rect 3930 1212 3943 1214
rect 3958 1212 3992 1214
rect 3595 1190 3608 1192
rect 3623 1190 3657 1192
rect 3595 1174 3657 1190
rect 3701 1185 3717 1192
rect 3779 1185 3809 1196
rect 3857 1192 3903 1208
rect 3930 1196 4004 1212
rect 3857 1190 3891 1192
rect 3856 1174 3903 1190
rect 3930 1174 3943 1196
rect 3958 1174 3988 1196
rect 4015 1174 4016 1190
rect 4031 1174 4044 1334
rect 4074 1230 4087 1334
rect 4132 1312 4133 1322
rect 4148 1312 4161 1322
rect 4132 1308 4161 1312
rect 4166 1308 4196 1334
rect 4214 1320 4230 1322
rect 4302 1320 4355 1334
rect 4303 1318 4367 1320
rect 4410 1318 4425 1334
rect 4474 1331 4504 1334
rect 4474 1328 4510 1331
rect 4440 1320 4456 1322
rect 4214 1308 4229 1312
rect 4132 1306 4229 1308
rect 4257 1306 4425 1318
rect 4441 1308 4456 1312
rect 4474 1309 4513 1328
rect 4532 1322 4539 1323
rect 4538 1315 4539 1322
rect 4522 1312 4523 1315
rect 4538 1312 4551 1315
rect 4474 1308 4504 1309
rect 4513 1308 4519 1309
rect 4522 1308 4551 1312
rect 4441 1307 4551 1308
rect 4441 1306 4557 1307
rect 4116 1298 4167 1306
rect 4116 1286 4141 1298
rect 4148 1286 4167 1298
rect 4198 1298 4248 1306
rect 4198 1290 4214 1298
rect 4221 1296 4248 1298
rect 4257 1296 4478 1306
rect 4221 1286 4478 1296
rect 4507 1298 4557 1306
rect 4507 1289 4523 1298
rect 4116 1278 4167 1286
rect 4214 1278 4478 1286
rect 4504 1286 4523 1289
rect 4530 1286 4557 1298
rect 4504 1278 4557 1286
rect 4132 1270 4133 1278
rect 4148 1270 4161 1278
rect 4132 1262 4148 1270
rect 4129 1255 4148 1258
rect 4129 1246 4151 1255
rect 4102 1236 4151 1246
rect 4102 1230 4132 1236
rect 4151 1231 4156 1236
rect 4074 1214 4148 1230
rect 4166 1222 4196 1278
rect 4231 1268 4439 1278
rect 4474 1274 4519 1278
rect 4522 1277 4523 1278
rect 4538 1277 4551 1278
rect 4257 1238 4446 1268
rect 4272 1235 4446 1238
rect 4265 1232 4446 1235
rect 4074 1212 4087 1214
rect 4102 1212 4136 1214
rect 4074 1196 4148 1212
rect 4175 1208 4188 1222
rect 4203 1208 4219 1224
rect 4265 1219 4276 1232
rect 4058 1174 4059 1190
rect 4074 1174 4087 1196
rect 4102 1174 4132 1196
rect 4175 1192 4237 1208
rect 4265 1201 4276 1217
rect 4281 1212 4291 1232
rect 4301 1212 4315 1232
rect 4318 1219 4327 1232
rect 4343 1219 4352 1232
rect 4281 1201 4315 1212
rect 4318 1201 4327 1217
rect 4343 1201 4352 1217
rect 4359 1212 4369 1232
rect 4379 1212 4393 1232
rect 4394 1219 4405 1232
rect 4359 1201 4393 1212
rect 4394 1201 4405 1217
rect 4451 1208 4467 1224
rect 4474 1222 4504 1274
rect 4538 1270 4539 1277
rect 4523 1262 4539 1270
rect 4510 1230 4523 1249
rect 4538 1230 4568 1246
rect 4510 1214 4584 1230
rect 4510 1212 4523 1214
rect 4538 1212 4572 1214
rect 4175 1190 4188 1192
rect 4203 1190 4237 1192
rect 4175 1174 4237 1190
rect 4281 1185 4297 1192
rect 4359 1185 4389 1196
rect 4437 1192 4483 1208
rect 4510 1196 4584 1212
rect 4437 1190 4471 1192
rect 4436 1174 4483 1190
rect 4510 1174 4523 1196
rect 4538 1174 4568 1196
rect 4595 1174 4596 1190
rect 4611 1174 4624 1334
rect 4654 1230 4667 1334
rect 4712 1312 4713 1322
rect 4728 1312 4741 1322
rect 4712 1308 4741 1312
rect 4746 1308 4776 1334
rect 4794 1320 4810 1322
rect 4882 1320 4933 1334
rect 4883 1318 4947 1320
rect 4990 1318 5005 1334
rect 5054 1331 5084 1334
rect 5054 1328 5090 1331
rect 5020 1320 5036 1322
rect 4794 1308 4809 1312
rect 4712 1306 4809 1308
rect 4837 1306 5005 1318
rect 5021 1308 5036 1312
rect 5054 1309 5093 1328
rect 5112 1322 5119 1323
rect 5118 1315 5119 1322
rect 5102 1312 5103 1315
rect 5118 1312 5131 1315
rect 5054 1308 5084 1309
rect 5093 1308 5099 1309
rect 5102 1308 5131 1312
rect 5021 1307 5131 1308
rect 5021 1306 5137 1307
rect 4696 1298 4747 1306
rect 4696 1286 4721 1298
rect 4728 1286 4747 1298
rect 4778 1298 4828 1306
rect 4778 1290 4794 1298
rect 4801 1296 4828 1298
rect 4837 1296 5058 1306
rect 4801 1286 5058 1296
rect 5087 1298 5137 1306
rect 5087 1289 5103 1298
rect 4696 1278 4747 1286
rect 4794 1278 5058 1286
rect 5084 1286 5103 1289
rect 5110 1286 5137 1298
rect 5084 1278 5137 1286
rect 4712 1270 4713 1278
rect 4728 1270 4741 1278
rect 4712 1262 4728 1270
rect 4709 1255 4728 1258
rect 4709 1246 4731 1255
rect 4682 1236 4731 1246
rect 4682 1230 4712 1236
rect 4731 1231 4736 1236
rect 4654 1214 4728 1230
rect 4746 1222 4776 1278
rect 4811 1268 5019 1278
rect 5054 1274 5099 1278
rect 5102 1277 5103 1278
rect 5118 1277 5131 1278
rect 4837 1238 5026 1268
rect 4852 1235 5026 1238
rect 4845 1232 5026 1235
rect 4654 1212 4667 1214
rect 4682 1212 4716 1214
rect 4654 1196 4728 1212
rect 4755 1208 4768 1222
rect 4783 1208 4799 1224
rect 4845 1219 4856 1232
rect 4638 1174 4639 1190
rect 4654 1174 4667 1196
rect 4682 1174 4712 1196
rect 4755 1192 4817 1208
rect 4845 1201 4856 1217
rect 4861 1212 4871 1232
rect 4881 1212 4895 1232
rect 4898 1219 4907 1232
rect 4923 1219 4932 1232
rect 4861 1201 4895 1212
rect 4898 1201 4907 1217
rect 4923 1201 4932 1217
rect 4939 1212 4949 1232
rect 4959 1212 4973 1232
rect 4974 1219 4985 1232
rect 4939 1201 4973 1212
rect 4974 1201 4985 1217
rect 5031 1208 5047 1224
rect 5054 1222 5084 1274
rect 5118 1270 5119 1277
rect 5103 1262 5119 1270
rect 5090 1230 5103 1249
rect 5118 1230 5148 1246
rect 5090 1214 5164 1230
rect 5090 1212 5103 1214
rect 5118 1212 5152 1214
rect 4755 1190 4768 1192
rect 4783 1190 4817 1192
rect 4755 1174 4817 1190
rect 4861 1185 4877 1192
rect 4939 1185 4969 1196
rect 5017 1192 5063 1208
rect 5090 1196 5164 1212
rect 5017 1190 5051 1192
rect 5016 1174 5063 1190
rect 5090 1174 5103 1196
rect 5118 1174 5148 1196
rect 5175 1174 5176 1190
rect 5191 1174 5204 1334
rect 5234 1230 5247 1334
rect 5292 1312 5293 1322
rect 5308 1312 5321 1322
rect 5292 1308 5321 1312
rect 5326 1308 5356 1334
rect 5374 1320 5390 1322
rect 5462 1320 5513 1334
rect 5463 1318 5527 1320
rect 5570 1318 5585 1334
rect 5634 1331 5664 1334
rect 5634 1328 5670 1331
rect 5600 1320 5616 1322
rect 5374 1308 5389 1312
rect 5292 1306 5389 1308
rect 5417 1306 5585 1318
rect 5601 1308 5616 1312
rect 5634 1309 5673 1328
rect 5692 1322 5699 1323
rect 5698 1315 5699 1322
rect 5682 1312 5683 1315
rect 5698 1312 5711 1315
rect 5634 1308 5664 1309
rect 5673 1308 5679 1309
rect 5682 1308 5711 1312
rect 5601 1307 5711 1308
rect 5601 1306 5717 1307
rect 5276 1298 5327 1306
rect 5276 1286 5301 1298
rect 5308 1286 5327 1298
rect 5358 1298 5408 1306
rect 5358 1290 5374 1298
rect 5381 1296 5408 1298
rect 5417 1296 5638 1306
rect 5381 1286 5638 1296
rect 5667 1298 5717 1306
rect 5667 1289 5683 1298
rect 5276 1278 5327 1286
rect 5374 1278 5638 1286
rect 5664 1286 5683 1289
rect 5690 1286 5717 1298
rect 5664 1278 5717 1286
rect 5292 1270 5293 1278
rect 5308 1270 5321 1278
rect 5292 1262 5308 1270
rect 5289 1255 5308 1258
rect 5289 1246 5311 1255
rect 5262 1236 5311 1246
rect 5262 1230 5292 1236
rect 5311 1231 5316 1236
rect 5234 1214 5308 1230
rect 5326 1222 5356 1278
rect 5391 1268 5599 1278
rect 5634 1274 5679 1278
rect 5682 1277 5683 1278
rect 5698 1277 5711 1278
rect 5417 1238 5606 1268
rect 5432 1235 5606 1238
rect 5425 1232 5606 1235
rect 5234 1212 5247 1214
rect 5262 1212 5296 1214
rect 5234 1196 5308 1212
rect 5335 1208 5348 1222
rect 5363 1208 5379 1224
rect 5425 1219 5436 1232
rect 5218 1174 5219 1190
rect 5234 1174 5247 1196
rect 5262 1174 5292 1196
rect 5335 1192 5397 1208
rect 5425 1201 5436 1217
rect 5441 1212 5451 1232
rect 5461 1212 5475 1232
rect 5478 1219 5487 1232
rect 5503 1219 5512 1232
rect 5441 1201 5475 1212
rect 5478 1201 5487 1217
rect 5503 1201 5512 1217
rect 5519 1212 5529 1232
rect 5539 1212 5553 1232
rect 5554 1219 5565 1232
rect 5519 1201 5553 1212
rect 5554 1201 5565 1217
rect 5611 1208 5627 1224
rect 5634 1222 5664 1274
rect 5698 1270 5699 1277
rect 5683 1262 5699 1270
rect 5670 1230 5683 1249
rect 5698 1230 5728 1246
rect 5670 1214 5744 1230
rect 5670 1212 5683 1214
rect 5698 1212 5732 1214
rect 5335 1190 5348 1192
rect 5363 1190 5397 1192
rect 5335 1174 5397 1190
rect 5441 1185 5457 1192
rect 5519 1185 5549 1196
rect 5597 1192 5643 1208
rect 5670 1196 5744 1212
rect 5597 1190 5631 1192
rect 5596 1174 5643 1190
rect 5670 1174 5683 1196
rect 5698 1174 5728 1196
rect 5755 1174 5756 1190
rect 5771 1174 5784 1334
rect 5814 1230 5827 1334
rect 5872 1312 5873 1322
rect 5888 1312 5901 1322
rect 5872 1308 5901 1312
rect 5906 1308 5936 1334
rect 5954 1320 5970 1322
rect 6042 1320 6093 1334
rect 6043 1318 6107 1320
rect 6150 1318 6165 1334
rect 6214 1331 6244 1334
rect 6214 1328 6250 1331
rect 6180 1320 6196 1322
rect 5954 1308 5969 1312
rect 5872 1306 5969 1308
rect 5997 1306 6165 1318
rect 6181 1308 6196 1312
rect 6214 1309 6253 1328
rect 6272 1322 6279 1323
rect 6278 1315 6279 1322
rect 6262 1312 6263 1315
rect 6278 1312 6291 1315
rect 6214 1308 6244 1309
rect 6253 1308 6259 1309
rect 6262 1308 6291 1312
rect 6181 1307 6291 1308
rect 6181 1306 6297 1307
rect 5856 1298 5907 1306
rect 5856 1286 5881 1298
rect 5888 1286 5907 1298
rect 5938 1298 5988 1306
rect 5938 1290 5954 1298
rect 5961 1296 5988 1298
rect 5997 1296 6218 1306
rect 5961 1286 6218 1296
rect 6247 1298 6297 1306
rect 6247 1289 6263 1298
rect 5856 1278 5907 1286
rect 5954 1278 6218 1286
rect 6244 1286 6263 1289
rect 6270 1286 6297 1298
rect 6244 1278 6297 1286
rect 5872 1270 5873 1278
rect 5888 1270 5901 1278
rect 5872 1262 5888 1270
rect 5869 1255 5888 1258
rect 5869 1246 5891 1255
rect 5842 1236 5891 1246
rect 5842 1230 5872 1236
rect 5891 1231 5896 1236
rect 5814 1214 5888 1230
rect 5906 1222 5936 1278
rect 5971 1268 6179 1278
rect 6214 1274 6259 1278
rect 6262 1277 6263 1278
rect 6278 1277 6291 1278
rect 5997 1238 6186 1268
rect 6012 1235 6186 1238
rect 6005 1232 6186 1235
rect 5814 1212 5827 1214
rect 5842 1212 5876 1214
rect 5814 1196 5888 1212
rect 5915 1208 5928 1222
rect 5943 1208 5959 1224
rect 6005 1219 6016 1232
rect 5798 1174 5799 1190
rect 5814 1174 5827 1196
rect 5842 1174 5872 1196
rect 5915 1192 5977 1208
rect 6005 1201 6016 1217
rect 6021 1212 6031 1232
rect 6041 1212 6055 1232
rect 6058 1219 6067 1232
rect 6083 1219 6092 1232
rect 6021 1201 6055 1212
rect 6058 1201 6067 1217
rect 6083 1201 6092 1217
rect 6099 1212 6109 1232
rect 6119 1212 6133 1232
rect 6134 1219 6145 1232
rect 6099 1201 6133 1212
rect 6134 1201 6145 1217
rect 6191 1208 6207 1224
rect 6214 1222 6244 1274
rect 6278 1270 6279 1277
rect 6263 1262 6279 1270
rect 6250 1230 6263 1249
rect 6278 1230 6308 1246
rect 6250 1214 6324 1230
rect 6250 1212 6263 1214
rect 6278 1212 6312 1214
rect 5915 1190 5928 1192
rect 5943 1190 5977 1192
rect 5915 1174 5977 1190
rect 6021 1185 6037 1192
rect 6099 1185 6129 1196
rect 6177 1192 6223 1208
rect 6250 1196 6324 1212
rect 6177 1190 6211 1192
rect 6176 1174 6223 1190
rect 6250 1174 6263 1196
rect 6278 1174 6308 1196
rect 6335 1174 6336 1190
rect 6351 1174 6364 1334
rect 6394 1230 6407 1334
rect 6452 1312 6453 1322
rect 6468 1312 6481 1322
rect 6452 1308 6481 1312
rect 6486 1308 6516 1334
rect 6534 1320 6550 1322
rect 6622 1320 6673 1334
rect 6623 1318 6687 1320
rect 6730 1318 6745 1334
rect 6794 1331 6824 1334
rect 6794 1328 6830 1331
rect 6760 1320 6776 1322
rect 6534 1308 6549 1312
rect 6452 1306 6549 1308
rect 6577 1306 6745 1318
rect 6761 1308 6776 1312
rect 6794 1309 6833 1328
rect 6852 1322 6859 1323
rect 6858 1315 6859 1322
rect 6842 1312 6843 1315
rect 6858 1312 6871 1315
rect 6794 1308 6824 1309
rect 6833 1308 6839 1309
rect 6842 1308 6871 1312
rect 6761 1307 6871 1308
rect 6761 1306 6877 1307
rect 6436 1298 6487 1306
rect 6436 1286 6461 1298
rect 6468 1286 6487 1298
rect 6518 1298 6568 1306
rect 6518 1290 6534 1298
rect 6541 1296 6568 1298
rect 6577 1296 6798 1306
rect 6541 1286 6798 1296
rect 6827 1298 6877 1306
rect 6827 1289 6843 1298
rect 6436 1278 6487 1286
rect 6534 1278 6798 1286
rect 6824 1286 6843 1289
rect 6850 1286 6877 1298
rect 6824 1278 6877 1286
rect 6452 1270 6453 1278
rect 6468 1270 6481 1278
rect 6452 1262 6468 1270
rect 6449 1255 6468 1258
rect 6449 1246 6471 1255
rect 6422 1236 6471 1246
rect 6422 1230 6452 1236
rect 6471 1231 6476 1236
rect 6394 1214 6468 1230
rect 6486 1222 6516 1278
rect 6551 1268 6759 1278
rect 6794 1274 6839 1278
rect 6842 1277 6843 1278
rect 6858 1277 6871 1278
rect 6577 1238 6766 1268
rect 6592 1235 6766 1238
rect 6585 1232 6766 1235
rect 6394 1212 6407 1214
rect 6422 1212 6456 1214
rect 6394 1196 6468 1212
rect 6495 1208 6508 1222
rect 6523 1208 6539 1224
rect 6585 1219 6596 1232
rect 6378 1174 6379 1190
rect 6394 1174 6407 1196
rect 6422 1174 6452 1196
rect 6495 1192 6557 1208
rect 6585 1201 6596 1217
rect 6601 1212 6611 1232
rect 6621 1212 6635 1232
rect 6638 1219 6647 1232
rect 6663 1219 6672 1232
rect 6601 1201 6635 1212
rect 6638 1201 6647 1217
rect 6663 1201 6672 1217
rect 6679 1212 6689 1232
rect 6699 1212 6713 1232
rect 6714 1219 6725 1232
rect 6679 1201 6713 1212
rect 6714 1201 6725 1217
rect 6771 1208 6787 1224
rect 6794 1222 6824 1274
rect 6858 1270 6859 1277
rect 6843 1262 6859 1270
rect 6830 1230 6843 1249
rect 6858 1230 6888 1246
rect 6830 1214 6904 1230
rect 6830 1212 6843 1214
rect 6858 1212 6892 1214
rect 6495 1190 6508 1192
rect 6523 1190 6557 1192
rect 6495 1174 6557 1190
rect 6601 1185 6617 1192
rect 6679 1185 6709 1196
rect 6757 1192 6803 1208
rect 6830 1196 6904 1212
rect 6757 1190 6791 1192
rect 6756 1174 6803 1190
rect 6830 1174 6843 1196
rect 6858 1174 6888 1196
rect 6915 1174 6916 1190
rect 6931 1174 6944 1334
rect -8 1166 33 1174
rect -8 1140 7 1166
rect 14 1140 33 1166
rect 97 1162 159 1174
rect 171 1162 246 1174
rect 304 1162 379 1174
rect 391 1162 422 1174
rect 428 1162 463 1174
rect 97 1160 259 1162
rect -8 1132 33 1140
rect 115 1136 128 1160
rect 143 1158 158 1160
rect -2 1122 -1 1132
rect 14 1122 27 1132
rect 42 1122 72 1136
rect 115 1122 158 1136
rect 182 1133 189 1140
rect 192 1136 259 1160
rect 291 1160 463 1162
rect 261 1138 289 1142
rect 291 1138 371 1160
rect 392 1158 407 1160
rect 261 1136 371 1138
rect 192 1132 371 1136
rect 165 1122 195 1132
rect 197 1122 350 1132
rect 358 1122 388 1132
rect 392 1122 422 1136
rect 450 1122 463 1160
rect 535 1166 570 1174
rect 535 1140 536 1166
rect 543 1140 570 1166
rect 478 1122 508 1136
rect 535 1132 570 1140
rect 572 1166 613 1174
rect 572 1140 587 1166
rect 594 1140 613 1166
rect 677 1162 739 1174
rect 751 1162 826 1174
rect 884 1162 959 1174
rect 971 1162 1002 1174
rect 1008 1162 1043 1174
rect 677 1160 839 1162
rect 572 1132 613 1140
rect 695 1136 708 1160
rect 723 1158 738 1160
rect 535 1122 536 1132
rect 551 1122 564 1132
rect 578 1122 579 1132
rect 594 1122 607 1132
rect 622 1122 652 1136
rect 695 1122 738 1136
rect 762 1133 769 1140
rect 772 1136 839 1160
rect 871 1160 1043 1162
rect 841 1138 869 1142
rect 871 1138 951 1160
rect 972 1158 987 1160
rect 841 1136 951 1138
rect 772 1132 951 1136
rect 745 1122 775 1132
rect 777 1122 930 1132
rect 938 1122 968 1132
rect 972 1122 1002 1136
rect 1030 1122 1043 1160
rect 1115 1166 1150 1174
rect 1115 1140 1116 1166
rect 1123 1140 1150 1166
rect 1058 1122 1088 1136
rect 1115 1132 1150 1140
rect 1152 1166 1193 1174
rect 1152 1140 1167 1166
rect 1174 1140 1193 1166
rect 1257 1160 1281 1174
rect 1152 1132 1193 1140
rect 1115 1122 1116 1132
rect 1131 1122 1144 1132
rect 1158 1122 1159 1132
rect 1174 1122 1187 1132
rect 1202 1122 1232 1136
rect 1275 1122 1281 1160
rect 3481 1166 3513 1174
rect 3481 1140 3487 1166
rect 3494 1140 3513 1166
rect 3577 1162 3639 1174
rect 3651 1162 3726 1174
rect 3784 1162 3859 1174
rect 3871 1162 3902 1174
rect 3908 1162 3943 1174
rect 3577 1160 3739 1162
rect 3481 1132 3513 1140
rect 3595 1136 3608 1160
rect 3623 1158 3638 1160
rect 3494 1122 3507 1132
rect 3522 1122 3552 1136
rect 3595 1122 3638 1136
rect 3662 1133 3669 1140
rect 3672 1136 3739 1160
rect 3771 1160 3943 1162
rect 3741 1138 3769 1142
rect 3771 1138 3851 1160
rect 3872 1158 3887 1160
rect 3741 1136 3851 1138
rect 3672 1132 3851 1136
rect 3645 1122 3675 1132
rect 3677 1122 3830 1132
rect 3838 1122 3868 1132
rect 3872 1122 3902 1136
rect 3930 1122 3943 1160
rect 4015 1166 4050 1174
rect 4015 1140 4016 1166
rect 4023 1140 4050 1166
rect 3958 1122 3988 1136
rect 4015 1132 4050 1140
rect 4052 1166 4093 1174
rect 4052 1140 4067 1166
rect 4074 1140 4093 1166
rect 4157 1162 4219 1174
rect 4231 1162 4306 1174
rect 4364 1162 4439 1174
rect 4451 1162 4482 1174
rect 4488 1162 4523 1174
rect 4157 1160 4319 1162
rect 4052 1132 4093 1140
rect 4175 1136 4188 1160
rect 4203 1158 4218 1160
rect 4015 1122 4016 1132
rect 4031 1122 4044 1132
rect 4058 1122 4059 1132
rect 4074 1122 4087 1132
rect 4102 1122 4132 1136
rect 4175 1122 4218 1136
rect 4242 1133 4249 1140
rect 4252 1136 4319 1160
rect 4351 1160 4523 1162
rect 4321 1138 4349 1142
rect 4351 1138 4431 1160
rect 4452 1158 4467 1160
rect 4321 1136 4431 1138
rect 4252 1132 4431 1136
rect 4225 1122 4255 1132
rect 4257 1122 4410 1132
rect 4418 1122 4448 1132
rect 4452 1122 4482 1136
rect 4510 1122 4523 1160
rect 4595 1166 4630 1174
rect 4595 1140 4596 1166
rect 4603 1140 4630 1166
rect 4538 1122 4568 1136
rect 4595 1132 4630 1140
rect 4632 1166 4673 1174
rect 4632 1140 4647 1166
rect 4654 1140 4673 1166
rect 4737 1162 4799 1174
rect 4811 1162 4886 1174
rect 4944 1162 5019 1174
rect 5031 1162 5062 1174
rect 5068 1162 5103 1174
rect 4737 1160 4899 1162
rect 4755 1142 4768 1160
rect 4783 1158 4798 1160
rect 4632 1132 4673 1140
rect 4756 1136 4768 1142
rect 4832 1142 4899 1160
rect 4931 1160 5103 1162
rect 4931 1142 5011 1160
rect 5032 1158 5047 1160
rect 4595 1122 4596 1132
rect 4611 1122 4624 1132
rect 4638 1122 4639 1132
rect 4654 1122 4667 1132
rect 4682 1122 4712 1136
rect 4756 1122 4798 1136
rect 4822 1133 4829 1140
rect 4832 1132 5011 1142
rect 4805 1122 4835 1132
rect 4837 1122 4990 1132
rect 4998 1122 5028 1132
rect 5032 1122 5062 1136
rect 5090 1122 5103 1160
rect 5175 1166 5210 1174
rect 5175 1140 5176 1166
rect 5183 1140 5210 1166
rect 5118 1122 5148 1136
rect 5175 1132 5210 1140
rect 5212 1166 5253 1174
rect 5212 1140 5227 1166
rect 5234 1140 5253 1166
rect 5317 1162 5379 1174
rect 5391 1162 5466 1174
rect 5524 1162 5599 1174
rect 5611 1162 5642 1174
rect 5648 1162 5683 1174
rect 5317 1160 5479 1162
rect 5335 1142 5348 1160
rect 5363 1158 5378 1160
rect 5212 1132 5253 1140
rect 5336 1136 5348 1142
rect 5412 1142 5479 1160
rect 5511 1160 5683 1162
rect 5511 1142 5591 1160
rect 5612 1158 5627 1160
rect 5175 1122 5176 1132
rect 5191 1122 5204 1132
rect 5218 1122 5219 1132
rect 5234 1122 5247 1132
rect 5262 1122 5292 1136
rect 5336 1122 5378 1136
rect 5402 1133 5409 1140
rect 5412 1132 5591 1142
rect 5385 1122 5415 1132
rect 5417 1122 5570 1132
rect 5578 1122 5608 1132
rect 5612 1122 5642 1136
rect 5670 1122 5683 1160
rect 5755 1166 5790 1174
rect 5755 1140 5756 1166
rect 5763 1140 5790 1166
rect 5698 1122 5728 1136
rect 5755 1132 5790 1140
rect 5792 1166 5833 1174
rect 5792 1140 5807 1166
rect 5814 1140 5833 1166
rect 5897 1162 5959 1174
rect 5971 1162 6046 1174
rect 6104 1162 6179 1174
rect 6191 1162 6222 1174
rect 6228 1162 6263 1174
rect 5897 1160 6059 1162
rect 5915 1142 5928 1160
rect 5943 1158 5958 1160
rect 5792 1132 5833 1140
rect 5916 1136 5928 1142
rect 5992 1142 6059 1160
rect 6091 1160 6263 1162
rect 6091 1142 6171 1160
rect 6192 1158 6207 1160
rect 5755 1122 5756 1132
rect 5771 1122 5784 1132
rect 5798 1122 5799 1132
rect 5814 1122 5827 1132
rect 5842 1122 5872 1136
rect 5916 1122 5958 1136
rect 5982 1133 5989 1140
rect 5992 1132 6171 1142
rect 5965 1122 5995 1132
rect 5997 1122 6150 1132
rect 6158 1122 6188 1132
rect 6192 1122 6222 1136
rect 6250 1122 6263 1160
rect 6335 1166 6370 1174
rect 6335 1140 6336 1166
rect 6343 1140 6370 1166
rect 6278 1122 6308 1136
rect 6335 1132 6370 1140
rect 6372 1166 6413 1174
rect 6372 1140 6387 1166
rect 6394 1140 6413 1166
rect 6477 1162 6539 1174
rect 6551 1162 6626 1174
rect 6684 1162 6759 1174
rect 6771 1162 6802 1174
rect 6808 1162 6843 1174
rect 6477 1160 6639 1162
rect 6495 1142 6508 1160
rect 6523 1158 6538 1160
rect 6372 1132 6413 1140
rect 6496 1136 6508 1142
rect 6572 1142 6639 1160
rect 6671 1160 6843 1162
rect 6671 1142 6751 1160
rect 6772 1158 6787 1160
rect 6335 1122 6336 1132
rect 6351 1122 6364 1132
rect 6378 1122 6379 1132
rect 6394 1122 6407 1132
rect 6422 1122 6452 1136
rect 6496 1122 6538 1136
rect 6562 1133 6569 1140
rect 6572 1132 6751 1142
rect 6545 1122 6575 1132
rect 6577 1122 6730 1132
rect 6738 1122 6768 1132
rect 6772 1122 6802 1136
rect 6830 1122 6843 1160
rect 6915 1166 6950 1174
rect 6915 1140 6916 1166
rect 6923 1140 6950 1166
rect 6858 1122 6888 1136
rect 6915 1132 6950 1140
rect 6915 1122 6916 1132
rect 6931 1122 6944 1132
rect -2 1116 1281 1122
rect -1 1108 1281 1116
rect 3481 1108 6944 1122
rect 14 1078 27 1108
rect 42 1090 72 1108
rect 115 1094 129 1108
rect 165 1094 385 1108
rect 116 1092 129 1094
rect 82 1080 97 1092
rect 79 1078 101 1080
rect 106 1078 136 1092
rect 197 1090 350 1094
rect 179 1078 371 1090
rect 414 1078 444 1092
rect 450 1078 463 1108
rect 478 1090 508 1108
rect 551 1078 564 1108
rect 594 1078 607 1108
rect 622 1090 652 1108
rect 695 1094 709 1108
rect 745 1094 965 1108
rect 696 1092 709 1094
rect 662 1080 677 1092
rect 659 1078 681 1080
rect 686 1078 716 1092
rect 777 1090 930 1094
rect 759 1078 951 1090
rect 994 1078 1024 1092
rect 1030 1078 1043 1108
rect 1058 1090 1088 1108
rect 1131 1078 1144 1108
rect 1174 1078 1187 1108
rect 1202 1090 1232 1108
rect 1275 1094 1281 1108
rect 1276 1092 1281 1094
rect 1242 1080 1257 1092
rect 1239 1078 1261 1080
rect 1266 1078 1281 1092
rect 3494 1078 3507 1108
rect 3522 1090 3552 1108
rect 3595 1094 3609 1108
rect 3645 1094 3865 1108
rect 3596 1092 3609 1094
rect 3562 1080 3577 1092
rect 3559 1078 3581 1080
rect 3586 1078 3616 1092
rect 3677 1090 3830 1094
rect 3659 1078 3851 1090
rect 3894 1078 3924 1092
rect 3930 1078 3943 1108
rect 3958 1090 3988 1108
rect 4031 1078 4044 1108
rect 4074 1078 4087 1108
rect 4102 1090 4132 1108
rect 4175 1094 4189 1108
rect 4225 1094 4445 1108
rect 4176 1092 4189 1094
rect 4142 1080 4157 1092
rect 4139 1078 4161 1080
rect 4166 1078 4196 1092
rect 4257 1090 4410 1094
rect 4239 1078 4431 1090
rect 4474 1078 4504 1092
rect 4510 1078 4523 1108
rect 4538 1090 4568 1108
rect 4611 1078 4624 1108
rect 4654 1078 4667 1108
rect 4682 1090 4712 1108
rect 4756 1092 4769 1108
rect 4805 1094 5025 1108
rect 4722 1080 4737 1092
rect 4719 1078 4741 1080
rect 4746 1078 4776 1092
rect 4837 1090 4990 1094
rect 4819 1078 5011 1090
rect 5054 1078 5084 1092
rect 5090 1078 5103 1108
rect 5118 1090 5148 1108
rect 5191 1078 5204 1108
rect 5234 1078 5247 1108
rect 5262 1090 5292 1108
rect 5336 1092 5349 1108
rect 5385 1094 5605 1108
rect 5302 1080 5317 1092
rect 5299 1078 5321 1080
rect 5326 1078 5356 1092
rect 5417 1090 5570 1094
rect 5399 1078 5591 1090
rect 5634 1078 5664 1092
rect 5670 1078 5683 1108
rect 5698 1090 5728 1108
rect 5771 1078 5784 1108
rect 5814 1078 5827 1108
rect 5842 1090 5872 1108
rect 5916 1092 5929 1108
rect 5965 1094 6185 1108
rect 5882 1080 5897 1092
rect 5879 1078 5901 1080
rect 5906 1078 5936 1092
rect 5997 1090 6150 1094
rect 5979 1078 6171 1090
rect 6214 1078 6244 1092
rect 6250 1078 6263 1108
rect 6278 1090 6308 1108
rect 6351 1078 6364 1108
rect 6394 1078 6407 1108
rect 6422 1090 6452 1108
rect 6496 1092 6509 1108
rect 6545 1094 6765 1108
rect 6462 1080 6477 1092
rect 6459 1078 6481 1080
rect 6486 1078 6516 1092
rect 6577 1090 6730 1094
rect 6559 1078 6751 1090
rect 6794 1078 6824 1092
rect 6830 1078 6843 1108
rect 6858 1090 6888 1108
rect 6931 1078 6944 1108
rect -1 1064 1281 1078
rect 3481 1064 6944 1078
rect 14 960 27 1064
rect 72 1042 73 1052
rect 88 1042 101 1052
rect 72 1038 101 1042
rect 106 1038 136 1064
rect 154 1050 170 1052
rect 242 1050 295 1064
rect 243 1048 307 1050
rect 350 1048 365 1064
rect 414 1061 444 1064
rect 414 1058 450 1061
rect 380 1050 396 1052
rect 154 1038 169 1042
rect 72 1036 169 1038
rect 197 1036 365 1048
rect 381 1038 396 1042
rect 414 1039 453 1058
rect 472 1052 479 1053
rect 478 1045 479 1052
rect 462 1042 463 1045
rect 478 1042 491 1045
rect 414 1038 444 1039
rect 453 1038 459 1039
rect 462 1038 491 1042
rect 381 1037 491 1038
rect 381 1036 497 1037
rect 56 1028 107 1036
rect 56 1016 81 1028
rect 88 1016 107 1028
rect 138 1028 188 1036
rect 138 1020 154 1028
rect 161 1026 188 1028
rect 197 1026 418 1036
rect 161 1016 418 1026
rect 447 1028 497 1036
rect 447 1019 463 1028
rect 56 1008 107 1016
rect 154 1008 418 1016
rect 444 1016 463 1019
rect 470 1016 497 1028
rect 444 1008 497 1016
rect 72 1000 73 1008
rect 88 1000 101 1008
rect 72 992 88 1000
rect 69 985 88 988
rect 69 976 91 985
rect 42 966 91 976
rect 42 960 72 966
rect 91 961 96 966
rect 14 944 88 960
rect 106 952 136 1008
rect 171 998 379 1008
rect 414 1004 459 1008
rect 462 1007 463 1008
rect 478 1007 491 1008
rect 197 968 386 998
rect 212 965 386 968
rect 205 962 386 965
rect 14 942 27 944
rect 42 942 76 944
rect 14 926 88 942
rect 115 938 128 952
rect 143 938 159 954
rect 205 949 216 962
rect -2 904 -1 920
rect 14 904 27 926
rect 42 904 72 926
rect 115 922 177 938
rect 205 931 216 947
rect 221 942 231 962
rect 241 942 255 962
rect 258 949 267 962
rect 283 949 292 962
rect 221 931 255 942
rect 258 931 267 947
rect 283 931 292 947
rect 299 942 309 962
rect 319 942 333 962
rect 334 949 345 962
rect 299 931 333 942
rect 334 931 345 947
rect 391 938 407 954
rect 414 952 444 1004
rect 478 1000 479 1007
rect 463 992 479 1000
rect 450 960 463 979
rect 478 960 508 976
rect 450 944 524 960
rect 450 942 463 944
rect 478 942 512 944
rect 115 920 128 922
rect 143 920 177 922
rect 115 904 177 920
rect 221 915 237 922
rect 299 915 329 926
rect 377 922 423 938
rect 450 926 524 942
rect 377 920 411 922
rect 376 904 423 920
rect 450 904 463 926
rect 478 904 508 926
rect 535 904 536 920
rect 551 904 564 1064
rect 594 960 607 1064
rect 652 1042 653 1052
rect 668 1042 681 1052
rect 652 1038 681 1042
rect 686 1038 716 1064
rect 734 1050 750 1052
rect 822 1050 875 1064
rect 823 1048 887 1050
rect 930 1048 945 1064
rect 994 1061 1024 1064
rect 994 1058 1030 1061
rect 960 1050 976 1052
rect 734 1038 749 1042
rect 652 1036 749 1038
rect 777 1036 945 1048
rect 961 1038 976 1042
rect 994 1039 1033 1058
rect 1052 1052 1059 1053
rect 1058 1045 1059 1052
rect 1042 1042 1043 1045
rect 1058 1042 1071 1045
rect 994 1038 1024 1039
rect 1033 1038 1039 1039
rect 1042 1038 1071 1042
rect 961 1037 1071 1038
rect 961 1036 1077 1037
rect 636 1028 687 1036
rect 636 1016 661 1028
rect 668 1016 687 1028
rect 718 1028 768 1036
rect 718 1020 734 1028
rect 741 1026 768 1028
rect 777 1026 998 1036
rect 741 1016 998 1026
rect 1027 1028 1077 1036
rect 1027 1019 1043 1028
rect 636 1008 687 1016
rect 734 1008 998 1016
rect 1024 1016 1043 1019
rect 1050 1016 1077 1028
rect 1024 1008 1077 1016
rect 652 1000 653 1008
rect 668 1000 681 1008
rect 652 992 668 1000
rect 649 985 668 988
rect 649 976 671 985
rect 622 966 671 976
rect 622 960 652 966
rect 671 961 676 966
rect 594 944 668 960
rect 686 952 716 1008
rect 751 998 959 1008
rect 994 1004 1039 1008
rect 1042 1007 1043 1008
rect 1058 1007 1071 1008
rect 777 968 966 998
rect 792 965 966 968
rect 785 962 966 965
rect 594 942 607 944
rect 622 942 656 944
rect 594 926 668 942
rect 695 938 708 952
rect 723 938 739 954
rect 785 949 796 962
rect 578 904 579 920
rect 594 904 607 926
rect 622 904 652 926
rect 695 922 757 938
rect 785 931 796 947
rect 801 942 811 962
rect 821 942 835 962
rect 838 949 847 962
rect 863 949 872 962
rect 801 931 835 942
rect 838 931 847 947
rect 863 931 872 947
rect 879 942 889 962
rect 899 942 913 962
rect 914 949 925 962
rect 879 931 913 942
rect 914 931 925 947
rect 971 938 987 954
rect 994 952 1024 1004
rect 1058 1000 1059 1007
rect 1043 992 1059 1000
rect 1030 960 1043 979
rect 1058 960 1088 976
rect 1030 944 1104 960
rect 1030 942 1043 944
rect 1058 942 1092 944
rect 695 920 708 922
rect 723 920 757 922
rect 695 904 757 920
rect 801 915 817 922
rect 879 915 909 926
rect 957 922 1003 938
rect 1030 926 1104 942
rect 957 920 991 922
rect 956 904 1003 920
rect 1030 904 1043 926
rect 1058 904 1088 926
rect 1115 904 1116 920
rect 1131 904 1144 1064
rect 1174 960 1187 1064
rect 1232 1042 1233 1052
rect 1248 1042 1261 1052
rect 1232 1038 1261 1042
rect 1266 1038 1281 1064
rect 1232 1036 1281 1038
rect 1216 1028 1267 1036
rect 1216 1016 1241 1028
rect 1248 1016 1267 1028
rect 1216 1008 1267 1016
rect 1232 1000 1233 1008
rect 1248 1000 1261 1008
rect 1232 992 1248 1000
rect 1229 985 1248 988
rect 1229 976 1251 985
rect 1202 966 1251 976
rect 1202 960 1232 966
rect 1251 961 1256 966
rect 1174 944 1248 960
rect 1266 952 1281 1008
rect 1174 942 1187 944
rect 1202 942 1236 944
rect 1174 926 1248 942
rect 1158 904 1159 920
rect 1174 904 1187 926
rect 1202 904 1232 926
rect 1275 904 1281 952
rect 3494 960 3507 1064
rect 3552 1042 3553 1052
rect 3568 1042 3581 1052
rect 3552 1038 3581 1042
rect 3586 1038 3616 1064
rect 3634 1050 3650 1052
rect 3722 1050 3775 1064
rect 3723 1048 3787 1050
rect 3830 1048 3845 1064
rect 3894 1061 3924 1064
rect 3894 1058 3930 1061
rect 3860 1050 3876 1052
rect 3634 1038 3649 1042
rect 3552 1036 3649 1038
rect 3677 1036 3845 1048
rect 3861 1038 3876 1042
rect 3894 1039 3933 1058
rect 3952 1052 3959 1053
rect 3958 1045 3959 1052
rect 3942 1042 3943 1045
rect 3958 1042 3971 1045
rect 3894 1038 3924 1039
rect 3933 1038 3939 1039
rect 3942 1038 3971 1042
rect 3861 1037 3971 1038
rect 3861 1036 3977 1037
rect 3536 1028 3587 1036
rect 3536 1016 3561 1028
rect 3568 1016 3587 1028
rect 3618 1028 3668 1036
rect 3618 1020 3634 1028
rect 3641 1026 3668 1028
rect 3677 1026 3898 1036
rect 3641 1016 3898 1026
rect 3927 1028 3977 1036
rect 3927 1019 3943 1028
rect 3536 1008 3587 1016
rect 3634 1008 3898 1016
rect 3924 1016 3943 1019
rect 3950 1016 3977 1028
rect 3924 1008 3977 1016
rect 3552 1000 3553 1008
rect 3568 1000 3581 1008
rect 3552 992 3568 1000
rect 3549 985 3568 988
rect 3549 976 3571 985
rect 3522 966 3571 976
rect 3522 960 3552 966
rect 3571 961 3576 966
rect 3494 944 3568 960
rect 3586 952 3616 1008
rect 3651 998 3859 1008
rect 3894 1004 3939 1008
rect 3942 1007 3943 1008
rect 3958 1007 3971 1008
rect 3677 968 3866 998
rect 3692 965 3866 968
rect 3685 962 3866 965
rect 3494 942 3507 944
rect 3522 942 3556 944
rect 3494 926 3568 942
rect 3595 938 3608 952
rect 3623 938 3639 954
rect 3685 949 3696 962
rect 3494 914 3507 926
rect 3522 914 3552 926
rect 3595 922 3657 938
rect 3685 931 3696 947
rect 3701 942 3711 962
rect 3721 942 3735 962
rect 3738 949 3747 962
rect 3763 949 3772 962
rect 3701 931 3735 942
rect 3738 931 3747 947
rect 3763 931 3772 947
rect 3779 942 3789 962
rect 3799 942 3813 962
rect 3814 949 3825 962
rect 3779 931 3813 942
rect 3814 931 3825 947
rect 3871 938 3887 954
rect 3894 952 3924 1004
rect 3958 1000 3959 1007
rect 3943 992 3959 1000
rect 3930 960 3943 979
rect 3958 960 3988 976
rect 3930 944 4004 960
rect 3930 942 3943 944
rect 3958 942 3992 944
rect 3595 920 3608 922
rect 3623 920 3657 922
rect 3595 914 3657 920
rect 3701 915 3717 922
rect 3779 915 3809 926
rect 3857 922 3903 938
rect 3930 926 4004 942
rect 3857 920 3891 922
rect 3857 914 3903 920
rect 3930 914 3943 926
rect 3958 914 3988 926
rect 4031 914 4044 1064
rect 4074 960 4087 1064
rect 4132 1042 4133 1052
rect 4148 1042 4161 1052
rect 4132 1038 4161 1042
rect 4166 1038 4196 1064
rect 4214 1050 4230 1052
rect 4302 1050 4355 1064
rect 4303 1048 4367 1050
rect 4410 1048 4425 1064
rect 4474 1061 4504 1064
rect 4474 1058 4510 1061
rect 4440 1050 4456 1052
rect 4214 1038 4229 1042
rect 4132 1036 4229 1038
rect 4257 1036 4425 1048
rect 4441 1038 4456 1042
rect 4474 1039 4513 1058
rect 4532 1052 4539 1053
rect 4538 1045 4539 1052
rect 4522 1042 4523 1045
rect 4538 1042 4551 1045
rect 4474 1038 4504 1039
rect 4513 1038 4519 1039
rect 4522 1038 4551 1042
rect 4441 1037 4551 1038
rect 4441 1036 4557 1037
rect 4116 1028 4167 1036
rect 4116 1016 4141 1028
rect 4148 1016 4167 1028
rect 4198 1028 4248 1036
rect 4198 1020 4214 1028
rect 4221 1026 4248 1028
rect 4257 1026 4478 1036
rect 4221 1016 4478 1026
rect 4507 1028 4557 1036
rect 4507 1019 4523 1028
rect 4116 1008 4167 1016
rect 4214 1008 4478 1016
rect 4504 1016 4523 1019
rect 4530 1016 4557 1028
rect 4504 1008 4557 1016
rect 4132 1000 4133 1008
rect 4148 1000 4161 1008
rect 4132 992 4148 1000
rect 4129 985 4148 988
rect 4129 976 4151 985
rect 4102 966 4151 976
rect 4102 960 4132 966
rect 4151 961 4156 966
rect 4074 944 4148 960
rect 4166 952 4196 1008
rect 4231 998 4439 1008
rect 4474 1004 4519 1008
rect 4522 1007 4523 1008
rect 4538 1007 4551 1008
rect 4257 968 4446 998
rect 4272 965 4446 968
rect 4265 962 4446 965
rect 4074 942 4087 944
rect 4102 942 4136 944
rect 4074 926 4148 942
rect 4175 938 4188 952
rect 4203 938 4219 954
rect 4265 949 4276 962
rect 4074 914 4087 926
rect 4102 914 4132 926
rect 4175 922 4237 938
rect 4265 931 4276 947
rect 4281 942 4291 962
rect 4301 942 4315 962
rect 4318 949 4327 962
rect 4343 949 4352 962
rect 4281 931 4315 942
rect 4318 931 4327 947
rect 4343 931 4352 947
rect 4359 942 4369 962
rect 4379 942 4393 962
rect 4394 949 4405 962
rect 4359 931 4393 942
rect 4394 931 4405 947
rect 4451 938 4467 954
rect 4474 952 4504 1004
rect 4538 1000 4539 1007
rect 4523 992 4539 1000
rect 4510 960 4523 979
rect 4538 960 4568 976
rect 4510 944 4584 960
rect 4510 942 4523 944
rect 4538 942 4572 944
rect 4175 920 4188 922
rect 4203 920 4237 922
rect 4175 914 4237 920
rect 4281 915 4297 922
rect 4359 915 4389 926
rect 4437 922 4483 938
rect 4510 926 4584 942
rect 4437 920 4471 922
rect 4437 914 4483 920
rect 4510 914 4523 926
rect 4538 914 4568 926
rect 4611 914 4624 1064
rect 4654 960 4667 1064
rect 4712 1042 4713 1052
rect 4728 1042 4741 1052
rect 4712 1038 4741 1042
rect 4746 1038 4776 1064
rect 4794 1050 4810 1052
rect 4882 1050 4933 1064
rect 4883 1048 4947 1050
rect 4990 1048 5005 1064
rect 5054 1061 5084 1064
rect 5054 1058 5090 1061
rect 5020 1050 5036 1052
rect 4794 1038 4809 1042
rect 4712 1036 4809 1038
rect 4837 1036 5005 1048
rect 5021 1038 5036 1042
rect 5054 1039 5093 1058
rect 5112 1052 5119 1053
rect 5118 1045 5119 1052
rect 5102 1042 5103 1045
rect 5118 1042 5131 1045
rect 5054 1038 5084 1039
rect 5093 1038 5099 1039
rect 5102 1038 5131 1042
rect 5021 1037 5131 1038
rect 5021 1036 5137 1037
rect 4696 1028 4747 1036
rect 4696 1016 4721 1028
rect 4728 1016 4747 1028
rect 4778 1028 4828 1036
rect 4778 1020 4794 1028
rect 4801 1026 4828 1028
rect 4837 1026 5058 1036
rect 4801 1016 5058 1026
rect 5087 1028 5137 1036
rect 5087 1019 5103 1028
rect 4696 1008 4747 1016
rect 4794 1008 5058 1016
rect 5084 1016 5103 1019
rect 5110 1016 5137 1028
rect 5084 1008 5137 1016
rect 4712 1000 4713 1008
rect 4728 1000 4741 1008
rect 4712 992 4728 1000
rect 4709 985 4728 988
rect 4709 976 4731 985
rect 4682 966 4731 976
rect 4682 960 4712 966
rect 4731 961 4736 966
rect 4654 944 4728 960
rect 4746 952 4776 1008
rect 4811 998 5019 1008
rect 5054 1004 5099 1008
rect 5102 1007 5103 1008
rect 5118 1007 5131 1008
rect 4837 968 5026 998
rect 4852 965 5026 968
rect 4845 962 5026 965
rect 4654 942 4667 944
rect 4682 942 4716 944
rect 4654 926 4728 942
rect 4755 938 4768 952
rect 4783 938 4799 954
rect 4845 949 4856 962
rect 4654 914 4667 926
rect 4682 914 4712 926
rect 4755 922 4817 938
rect 4845 931 4856 947
rect 4861 942 4871 962
rect 4881 942 4895 962
rect 4898 949 4907 962
rect 4923 949 4932 962
rect 4861 931 4895 942
rect 4898 931 4907 947
rect 4923 931 4932 947
rect 4939 942 4949 962
rect 4959 942 4973 962
rect 4974 949 4985 962
rect 4939 931 4973 942
rect 4974 931 4985 947
rect 5031 938 5047 954
rect 5054 952 5084 1004
rect 5118 1000 5119 1007
rect 5103 992 5119 1000
rect 5090 960 5103 979
rect 5118 960 5148 976
rect 5090 944 5164 960
rect 5090 942 5103 944
rect 5118 942 5152 944
rect 4755 920 4768 922
rect 4783 920 4817 922
rect 4755 914 4817 920
rect 4861 915 4877 922
rect 4939 915 4969 926
rect 5017 922 5063 938
rect 5090 926 5164 942
rect 5017 920 5051 922
rect 5017 914 5063 920
rect 5090 914 5103 926
rect 5118 914 5148 926
rect 5191 914 5204 1064
rect 5234 960 5247 1064
rect 5292 1042 5293 1052
rect 5308 1042 5321 1052
rect 5292 1038 5321 1042
rect 5326 1038 5356 1064
rect 5374 1050 5390 1052
rect 5462 1050 5513 1064
rect 5463 1048 5527 1050
rect 5570 1048 5585 1064
rect 5634 1061 5664 1064
rect 5634 1058 5670 1061
rect 5600 1050 5616 1052
rect 5374 1038 5389 1042
rect 5292 1036 5389 1038
rect 5417 1036 5585 1048
rect 5601 1038 5616 1042
rect 5634 1039 5673 1058
rect 5692 1052 5699 1053
rect 5698 1045 5699 1052
rect 5682 1042 5683 1045
rect 5698 1042 5711 1045
rect 5634 1038 5664 1039
rect 5673 1038 5679 1039
rect 5682 1038 5711 1042
rect 5601 1037 5711 1038
rect 5601 1036 5717 1037
rect 5276 1028 5327 1036
rect 5276 1016 5301 1028
rect 5308 1016 5327 1028
rect 5358 1028 5408 1036
rect 5358 1020 5374 1028
rect 5381 1026 5408 1028
rect 5417 1026 5638 1036
rect 5381 1016 5638 1026
rect 5667 1028 5717 1036
rect 5667 1019 5683 1028
rect 5276 1008 5327 1016
rect 5374 1008 5638 1016
rect 5664 1016 5683 1019
rect 5690 1016 5717 1028
rect 5664 1008 5717 1016
rect 5292 1000 5293 1008
rect 5308 1000 5321 1008
rect 5292 992 5308 1000
rect 5289 985 5308 988
rect 5289 976 5311 985
rect 5262 966 5311 976
rect 5262 960 5292 966
rect 5311 961 5316 966
rect 5234 944 5308 960
rect 5326 952 5356 1008
rect 5391 998 5599 1008
rect 5634 1004 5679 1008
rect 5682 1007 5683 1008
rect 5698 1007 5711 1008
rect 5417 968 5606 998
rect 5432 965 5606 968
rect 5425 962 5606 965
rect 5234 942 5247 944
rect 5262 942 5296 944
rect 5234 926 5308 942
rect 5335 938 5348 952
rect 5363 938 5379 954
rect 5425 949 5436 962
rect 5234 914 5247 926
rect 5262 914 5292 926
rect 5335 922 5397 938
rect 5425 931 5436 947
rect 5441 942 5451 962
rect 5461 942 5475 962
rect 5478 949 5487 962
rect 5503 949 5512 962
rect 5441 931 5475 942
rect 5478 931 5487 947
rect 5503 931 5512 947
rect 5519 942 5529 962
rect 5539 942 5553 962
rect 5554 949 5565 962
rect 5519 931 5553 942
rect 5554 931 5565 947
rect 5611 938 5627 954
rect 5634 952 5664 1004
rect 5698 1000 5699 1007
rect 5683 992 5699 1000
rect 5670 960 5683 979
rect 5698 960 5728 976
rect 5670 944 5744 960
rect 5670 942 5683 944
rect 5698 942 5732 944
rect 5335 920 5348 922
rect 5363 920 5397 922
rect 5335 914 5397 920
rect 5441 915 5457 922
rect 5519 915 5549 926
rect 5597 922 5643 938
rect 5670 926 5744 942
rect 5597 920 5631 922
rect 5597 914 5643 920
rect 5670 914 5683 926
rect 5698 914 5728 926
rect 5771 914 5784 1064
rect 5814 960 5827 1064
rect 5872 1042 5873 1052
rect 5888 1042 5901 1052
rect 5872 1038 5901 1042
rect 5906 1038 5936 1064
rect 5954 1050 5970 1052
rect 6042 1050 6093 1064
rect 6043 1048 6107 1050
rect 6150 1048 6165 1064
rect 6214 1061 6244 1064
rect 6214 1058 6250 1061
rect 6180 1050 6196 1052
rect 5954 1038 5969 1042
rect 5872 1036 5969 1038
rect 5997 1036 6165 1048
rect 6181 1038 6196 1042
rect 6214 1039 6253 1058
rect 6272 1052 6279 1053
rect 6278 1045 6279 1052
rect 6262 1042 6263 1045
rect 6278 1042 6291 1045
rect 6214 1038 6244 1039
rect 6253 1038 6259 1039
rect 6262 1038 6291 1042
rect 6181 1037 6291 1038
rect 6181 1036 6297 1037
rect 5856 1028 5907 1036
rect 5856 1016 5881 1028
rect 5888 1016 5907 1028
rect 5938 1028 5988 1036
rect 5938 1020 5954 1028
rect 5961 1026 5988 1028
rect 5997 1026 6218 1036
rect 5961 1016 6218 1026
rect 6247 1028 6297 1036
rect 6247 1019 6263 1028
rect 5856 1008 5907 1016
rect 5954 1008 6218 1016
rect 6244 1016 6263 1019
rect 6270 1016 6297 1028
rect 6244 1008 6297 1016
rect 5872 1000 5873 1008
rect 5888 1000 5901 1008
rect 5872 992 5888 1000
rect 5869 985 5888 988
rect 5869 976 5891 985
rect 5842 966 5891 976
rect 5842 960 5872 966
rect 5891 961 5896 966
rect 5814 944 5888 960
rect 5906 952 5936 1008
rect 5971 998 6179 1008
rect 6214 1004 6259 1008
rect 6262 1007 6263 1008
rect 6278 1007 6291 1008
rect 5997 968 6186 998
rect 6012 965 6186 968
rect 6005 962 6186 965
rect 5814 942 5827 944
rect 5842 942 5876 944
rect 5814 926 5888 942
rect 5915 938 5928 952
rect 5943 938 5959 954
rect 6005 949 6016 962
rect 5814 914 5827 926
rect 5842 914 5872 926
rect 5915 922 5977 938
rect 6005 931 6016 947
rect 6021 942 6031 962
rect 6041 942 6055 962
rect 6058 949 6067 962
rect 6083 949 6092 962
rect 6021 931 6055 942
rect 6058 931 6067 947
rect 6083 931 6092 947
rect 6099 942 6109 962
rect 6119 942 6133 962
rect 6134 949 6145 962
rect 6099 931 6133 942
rect 6134 931 6145 947
rect 6191 938 6207 954
rect 6214 952 6244 1004
rect 6278 1000 6279 1007
rect 6263 992 6279 1000
rect 6250 960 6263 979
rect 6278 960 6308 976
rect 6250 944 6324 960
rect 6250 942 6263 944
rect 6278 942 6312 944
rect 5915 920 5928 922
rect 5943 920 5977 922
rect 5915 914 5977 920
rect 6021 915 6037 922
rect 6099 915 6129 926
rect 6177 922 6223 938
rect 6250 926 6324 942
rect 6177 920 6211 922
rect 6177 914 6223 920
rect 6250 914 6263 926
rect 6278 914 6308 926
rect 6351 914 6364 1064
rect 6394 960 6407 1064
rect 6452 1042 6453 1052
rect 6468 1042 6481 1052
rect 6452 1038 6481 1042
rect 6486 1038 6516 1064
rect 6534 1050 6550 1052
rect 6622 1050 6673 1064
rect 6623 1048 6687 1050
rect 6730 1048 6745 1064
rect 6794 1061 6824 1064
rect 6794 1058 6830 1061
rect 6760 1050 6776 1052
rect 6534 1038 6549 1042
rect 6452 1036 6549 1038
rect 6577 1036 6745 1048
rect 6761 1038 6776 1042
rect 6794 1039 6833 1058
rect 6852 1052 6859 1053
rect 6858 1045 6859 1052
rect 6842 1042 6843 1045
rect 6858 1042 6871 1045
rect 6794 1038 6824 1039
rect 6833 1038 6839 1039
rect 6842 1038 6871 1042
rect 6761 1037 6871 1038
rect 6761 1036 6877 1037
rect 6436 1028 6487 1036
rect 6436 1016 6461 1028
rect 6468 1016 6487 1028
rect 6518 1028 6568 1036
rect 6518 1020 6534 1028
rect 6541 1026 6568 1028
rect 6577 1026 6798 1036
rect 6541 1016 6798 1026
rect 6827 1028 6877 1036
rect 6827 1019 6843 1028
rect 6436 1008 6487 1016
rect 6534 1008 6798 1016
rect 6824 1016 6843 1019
rect 6850 1016 6877 1028
rect 6824 1008 6877 1016
rect 6452 1000 6453 1008
rect 6468 1000 6481 1008
rect 6452 992 6468 1000
rect 6449 985 6468 988
rect 6449 976 6471 985
rect 6422 966 6471 976
rect 6422 960 6452 966
rect 6471 961 6476 966
rect 6394 944 6468 960
rect 6486 952 6516 1008
rect 6551 998 6759 1008
rect 6794 1004 6839 1008
rect 6842 1007 6843 1008
rect 6858 1007 6871 1008
rect 6577 968 6766 998
rect 6592 965 6766 968
rect 6585 962 6766 965
rect 6394 942 6407 944
rect 6422 942 6456 944
rect 6394 926 6468 942
rect 6495 938 6508 952
rect 6523 938 6539 954
rect 6585 949 6596 962
rect 6394 914 6407 926
rect 6422 914 6452 926
rect 6495 922 6557 938
rect 6585 931 6596 947
rect 6601 942 6611 962
rect 6621 942 6635 962
rect 6638 949 6647 962
rect 6663 949 6672 962
rect 6601 931 6635 942
rect 6638 931 6647 947
rect 6663 931 6672 947
rect 6679 942 6689 962
rect 6699 942 6713 962
rect 6714 949 6725 962
rect 6679 931 6713 942
rect 6714 931 6725 947
rect 6771 938 6787 954
rect 6794 952 6824 1004
rect 6858 1000 6859 1007
rect 6843 992 6859 1000
rect 6830 960 6843 979
rect 6858 960 6888 976
rect 6830 944 6904 960
rect 6830 942 6843 944
rect 6858 942 6892 944
rect 6495 920 6508 922
rect 6523 920 6557 922
rect 6495 914 6557 920
rect 6601 915 6617 922
rect 6679 915 6709 926
rect 6757 922 6803 938
rect 6830 926 6904 942
rect 6757 920 6791 922
rect 6757 914 6803 920
rect 6830 914 6843 926
rect 6858 914 6888 926
rect 6931 914 6944 1064
rect -8 896 33 904
rect -8 870 7 896
rect 14 870 33 896
rect 97 892 159 904
rect 171 892 246 904
rect 304 892 379 904
rect 391 892 422 904
rect 428 892 463 904
rect 97 890 259 892
rect -8 862 33 870
rect 115 866 128 890
rect 143 888 158 890
rect -2 852 -1 862
rect 14 852 27 862
rect 42 852 72 866
rect 115 852 158 866
rect 182 863 189 870
rect 192 866 259 890
rect 291 890 463 892
rect 261 868 289 872
rect 291 868 371 890
rect 392 888 407 890
rect 261 866 371 868
rect 192 862 371 866
rect 165 852 195 862
rect 197 852 350 862
rect 358 852 388 862
rect 392 852 422 866
rect 450 852 463 890
rect 535 896 570 904
rect 535 870 536 896
rect 543 870 570 896
rect 478 852 508 866
rect 535 862 570 870
rect 572 896 613 904
rect 572 870 587 896
rect 594 870 613 896
rect 677 892 739 904
rect 751 892 826 904
rect 884 892 959 904
rect 971 892 1002 904
rect 1008 892 1043 904
rect 677 890 839 892
rect 572 862 613 870
rect 695 866 708 890
rect 723 888 738 890
rect 535 852 536 862
rect 551 852 564 862
rect 578 852 579 862
rect 594 852 607 862
rect 622 852 652 866
rect 695 852 738 866
rect 762 863 769 870
rect 772 866 839 890
rect 871 890 1043 892
rect 841 868 869 872
rect 871 868 951 890
rect 972 888 987 890
rect 841 866 951 868
rect 772 862 951 866
rect 745 852 775 862
rect 777 852 930 862
rect 938 852 968 862
rect 972 852 1002 866
rect 1030 852 1043 890
rect 1115 896 1150 904
rect 1115 870 1116 896
rect 1123 870 1150 896
rect 1058 852 1088 866
rect 1115 862 1150 870
rect 1152 896 1193 904
rect 1152 870 1167 896
rect 1174 870 1193 896
rect 1257 890 1281 904
rect 1152 862 1193 870
rect 1115 852 1116 862
rect 1131 852 1144 862
rect 1158 852 1159 862
rect 1174 852 1187 862
rect 1202 852 1232 866
rect 1275 852 1281 890
rect -2 846 1281 852
rect -1 838 1281 846
rect 14 808 27 838
rect 42 820 72 838
rect 115 824 129 838
rect 165 824 385 838
rect 116 822 129 824
rect 82 810 97 822
rect 79 808 101 810
rect 106 808 136 822
rect 197 820 350 824
rect 179 808 371 820
rect 414 808 444 822
rect 450 808 463 838
rect 478 820 508 838
rect 551 808 564 838
rect 594 808 607 838
rect 622 820 652 838
rect 695 824 709 838
rect 745 824 965 838
rect 696 822 709 824
rect 662 810 677 822
rect 659 808 681 810
rect 686 808 716 822
rect 777 820 930 824
rect 759 808 951 820
rect 994 808 1024 822
rect 1030 808 1043 838
rect 1058 820 1088 838
rect 1131 808 1144 838
rect 1174 808 1187 838
rect 1202 820 1232 838
rect 1275 824 1281 838
rect 1276 822 1281 824
rect 1242 810 1257 822
rect 1239 808 1261 810
rect 1266 808 1281 822
rect -1 794 1281 808
rect 14 690 27 794
rect 72 772 73 782
rect 88 772 101 782
rect 72 768 101 772
rect 106 768 136 794
rect 154 780 170 782
rect 242 780 295 794
rect 243 778 307 780
rect 350 778 365 794
rect 414 791 444 794
rect 414 788 450 791
rect 380 780 396 782
rect 154 768 169 772
rect 72 766 169 768
rect 197 766 365 778
rect 381 768 396 772
rect 414 769 453 788
rect 472 782 479 783
rect 478 775 479 782
rect 462 772 463 775
rect 478 772 491 775
rect 414 768 444 769
rect 453 768 459 769
rect 462 768 491 772
rect 381 767 491 768
rect 381 766 497 767
rect 56 758 107 766
rect 56 746 81 758
rect 88 746 107 758
rect 138 758 188 766
rect 138 750 154 758
rect 161 756 188 758
rect 197 756 418 766
rect 161 746 418 756
rect 447 758 497 766
rect 447 749 463 758
rect 56 738 107 746
rect 154 738 418 746
rect 444 746 463 749
rect 470 746 497 758
rect 444 738 497 746
rect 72 730 73 738
rect 88 730 101 738
rect 72 722 88 730
rect 69 715 88 718
rect 69 706 91 715
rect 42 696 91 706
rect 42 690 72 696
rect 91 691 96 696
rect 14 674 88 690
rect 106 682 136 738
rect 171 728 379 738
rect 414 734 459 738
rect 462 737 463 738
rect 478 737 491 738
rect 197 698 386 728
rect 212 695 386 698
rect 205 692 386 695
rect 14 672 27 674
rect 42 672 76 674
rect 14 656 88 672
rect 115 668 128 682
rect 143 668 159 684
rect 205 679 216 692
rect -2 634 -1 650
rect 14 634 27 656
rect 42 634 72 656
rect 115 652 177 668
rect 205 661 216 677
rect 221 672 231 692
rect 241 672 255 692
rect 258 679 267 692
rect 283 679 292 692
rect 221 661 255 672
rect 258 661 267 677
rect 283 661 292 677
rect 299 672 309 692
rect 319 672 333 692
rect 334 679 345 692
rect 299 661 333 672
rect 334 661 345 677
rect 391 668 407 684
rect 414 682 444 734
rect 478 730 479 737
rect 463 722 479 730
rect 450 690 463 709
rect 478 690 508 706
rect 450 674 524 690
rect 450 672 463 674
rect 478 672 512 674
rect 115 650 128 652
rect 143 650 177 652
rect 115 634 177 650
rect 221 645 237 652
rect 299 645 329 656
rect 377 652 423 668
rect 450 656 524 672
rect 377 650 411 652
rect 376 634 423 650
rect 450 634 463 656
rect 478 634 508 656
rect 535 634 536 650
rect 551 634 564 794
rect 594 690 607 794
rect 652 772 653 782
rect 668 772 681 782
rect 652 768 681 772
rect 686 768 716 794
rect 734 780 750 782
rect 822 780 875 794
rect 823 778 887 780
rect 930 778 945 794
rect 994 791 1024 794
rect 994 788 1030 791
rect 960 780 976 782
rect 734 768 749 772
rect 652 766 749 768
rect 777 766 945 778
rect 961 768 976 772
rect 994 769 1033 788
rect 1052 782 1059 783
rect 1058 775 1059 782
rect 1042 772 1043 775
rect 1058 772 1071 775
rect 994 768 1024 769
rect 1033 768 1039 769
rect 1042 768 1071 772
rect 961 767 1071 768
rect 961 766 1077 767
rect 636 758 687 766
rect 636 746 661 758
rect 668 746 687 758
rect 718 758 768 766
rect 718 750 734 758
rect 741 756 768 758
rect 777 756 998 766
rect 741 746 998 756
rect 1027 758 1077 766
rect 1027 749 1043 758
rect 636 738 687 746
rect 734 738 998 746
rect 1024 746 1043 749
rect 1050 746 1077 758
rect 1024 738 1077 746
rect 652 730 653 738
rect 668 730 681 738
rect 652 722 668 730
rect 649 715 668 718
rect 649 706 671 715
rect 622 696 671 706
rect 622 690 652 696
rect 671 691 676 696
rect 594 674 668 690
rect 686 682 716 738
rect 751 728 959 738
rect 994 734 1039 738
rect 1042 737 1043 738
rect 1058 737 1071 738
rect 777 698 966 728
rect 792 695 966 698
rect 785 692 966 695
rect 594 672 607 674
rect 622 672 656 674
rect 594 656 668 672
rect 695 668 708 682
rect 723 668 739 684
rect 785 679 796 692
rect 578 634 579 650
rect 594 634 607 656
rect 622 634 652 656
rect 695 652 757 668
rect 785 661 796 677
rect 801 672 811 692
rect 821 672 835 692
rect 838 679 847 692
rect 863 679 872 692
rect 801 661 835 672
rect 838 661 847 677
rect 863 661 872 677
rect 879 672 889 692
rect 899 672 913 692
rect 914 679 925 692
rect 879 661 913 672
rect 914 661 925 677
rect 971 668 987 684
rect 994 682 1024 734
rect 1058 730 1059 737
rect 1043 722 1059 730
rect 1030 690 1043 709
rect 1058 690 1088 706
rect 1030 674 1104 690
rect 1030 672 1043 674
rect 1058 672 1092 674
rect 695 650 708 652
rect 723 650 757 652
rect 695 634 757 650
rect 801 645 817 652
rect 879 645 909 656
rect 957 652 1003 668
rect 1030 656 1104 672
rect 957 650 991 652
rect 956 634 1003 650
rect 1030 634 1043 656
rect 1058 634 1088 656
rect 1115 634 1116 650
rect 1131 634 1144 794
rect 1174 690 1187 794
rect 1232 772 1233 782
rect 1248 772 1261 782
rect 1232 768 1261 772
rect 1266 768 1281 794
rect 1232 766 1281 768
rect 1216 758 1267 766
rect 1216 746 1241 758
rect 1248 746 1267 758
rect 1216 738 1267 746
rect 1232 730 1233 738
rect 1248 730 1261 738
rect 1232 722 1248 730
rect 1229 715 1248 718
rect 1229 706 1251 715
rect 1202 696 1251 706
rect 1202 690 1232 696
rect 1251 691 1256 696
rect 1174 674 1248 690
rect 1266 682 1281 738
rect 1174 672 1187 674
rect 1202 672 1236 674
rect 1174 656 1248 672
rect 1158 634 1159 650
rect 1174 634 1187 656
rect 1202 634 1232 656
rect 1275 634 1281 682
rect -8 626 33 634
rect -8 600 7 626
rect 14 600 33 626
rect 97 622 159 634
rect 171 622 246 634
rect 304 622 379 634
rect 391 622 422 634
rect 428 622 463 634
rect 97 620 259 622
rect -8 592 33 600
rect 115 596 128 620
rect 143 618 158 620
rect -2 582 -1 592
rect 14 582 27 592
rect 42 582 72 596
rect 115 582 158 596
rect 182 593 189 600
rect 192 596 259 620
rect 291 620 463 622
rect 261 598 289 602
rect 291 598 371 620
rect 392 618 407 620
rect 261 596 371 598
rect 192 592 371 596
rect 165 582 195 592
rect 197 582 350 592
rect 358 582 388 592
rect 392 582 422 596
rect 450 582 463 620
rect 535 626 570 634
rect 535 600 536 626
rect 543 600 570 626
rect 478 582 508 596
rect 535 592 570 600
rect 572 626 613 634
rect 572 600 587 626
rect 594 600 613 626
rect 677 622 739 634
rect 751 622 826 634
rect 884 622 959 634
rect 971 622 1002 634
rect 1008 622 1043 634
rect 677 620 839 622
rect 572 592 613 600
rect 695 596 708 620
rect 723 618 738 620
rect 535 582 536 592
rect 551 582 564 592
rect 578 582 579 592
rect 594 582 607 592
rect 622 582 652 596
rect 695 582 738 596
rect 762 593 769 600
rect 772 596 839 620
rect 871 620 1043 622
rect 841 598 869 602
rect 871 598 951 620
rect 972 618 987 620
rect 841 596 951 598
rect 772 592 951 596
rect 745 582 775 592
rect 777 582 930 592
rect 938 582 968 592
rect 972 582 1002 596
rect 1030 582 1043 620
rect 1115 626 1150 634
rect 1115 600 1116 626
rect 1123 600 1150 626
rect 1058 582 1088 596
rect 1115 592 1150 600
rect 1152 626 1193 634
rect 1152 600 1167 626
rect 1174 600 1193 626
rect 1257 620 1281 634
rect 1152 592 1193 600
rect 1115 582 1116 592
rect 1131 582 1144 592
rect 1158 582 1159 592
rect 1174 582 1187 592
rect 1202 582 1232 596
rect 1275 582 1281 620
rect -2 576 1281 582
rect -1 568 1281 576
rect 14 538 27 568
rect 42 550 72 568
rect 115 554 129 568
rect 165 554 385 568
rect 116 552 129 554
rect 82 540 97 552
rect 79 538 101 540
rect 106 538 136 552
rect 197 550 350 554
rect 179 538 371 550
rect 414 538 444 552
rect 450 538 463 568
rect 478 550 508 568
rect 551 538 564 568
rect 594 538 607 568
rect 622 550 652 568
rect 695 554 709 568
rect 745 554 965 568
rect 696 552 709 554
rect 662 540 677 552
rect 659 538 681 540
rect 686 538 716 552
rect 777 550 930 554
rect 759 538 951 550
rect 994 538 1024 552
rect 1030 538 1043 568
rect 1058 550 1088 568
rect 1131 538 1144 568
rect 1174 538 1187 568
rect 1202 550 1232 568
rect 1275 554 1281 568
rect 1276 552 1281 554
rect 1242 540 1257 552
rect 1239 538 1261 540
rect 1266 538 1281 552
rect -1 524 1281 538
rect 14 420 27 524
rect 72 502 73 512
rect 88 502 101 512
rect 72 498 101 502
rect 106 498 136 524
rect 154 510 170 512
rect 242 510 295 524
rect 243 508 307 510
rect 350 508 365 524
rect 414 521 444 524
rect 414 518 450 521
rect 380 510 396 512
rect 154 498 169 502
rect 72 496 169 498
rect 197 496 365 508
rect 381 498 396 502
rect 414 499 453 518
rect 472 512 479 513
rect 478 505 479 512
rect 462 502 463 505
rect 478 502 491 505
rect 414 498 444 499
rect 453 498 459 499
rect 462 498 491 502
rect 381 497 491 498
rect 381 496 497 497
rect 56 488 107 496
rect 56 476 81 488
rect 88 476 107 488
rect 138 488 188 496
rect 138 480 154 488
rect 161 486 188 488
rect 197 486 418 496
rect 161 476 418 486
rect 447 488 497 496
rect 447 479 463 488
rect 56 468 107 476
rect 154 468 418 476
rect 444 476 463 479
rect 470 476 497 488
rect 444 468 497 476
rect 72 460 73 468
rect 88 460 101 468
rect 72 452 88 460
rect 69 445 88 448
rect 69 436 91 445
rect 42 426 91 436
rect 42 420 72 426
rect 91 421 96 426
rect 14 404 88 420
rect 106 412 136 468
rect 171 458 379 468
rect 414 464 459 468
rect 462 467 463 468
rect 478 467 491 468
rect 197 428 386 458
rect 212 425 386 428
rect 205 422 386 425
rect 14 402 27 404
rect 42 402 76 404
rect 14 386 88 402
rect 115 398 128 412
rect 143 398 159 414
rect 205 409 216 422
rect -2 364 -1 380
rect 14 364 27 386
rect 42 364 72 386
rect 115 382 177 398
rect 205 391 216 407
rect 221 402 231 422
rect 241 402 255 422
rect 258 409 267 422
rect 283 409 292 422
rect 221 391 255 402
rect 258 391 267 407
rect 283 391 292 407
rect 299 402 309 422
rect 319 402 333 422
rect 334 409 345 422
rect 299 391 333 402
rect 334 391 345 407
rect 391 398 407 414
rect 414 412 444 464
rect 478 460 479 467
rect 463 452 479 460
rect 450 420 463 439
rect 478 420 508 436
rect 450 404 524 420
rect 450 402 463 404
rect 478 402 512 404
rect 115 380 128 382
rect 143 380 177 382
rect 115 364 177 380
rect 221 375 237 382
rect 299 375 329 386
rect 377 382 423 398
rect 450 386 524 402
rect 377 380 411 382
rect 376 364 423 380
rect 450 364 463 386
rect 478 364 508 386
rect 535 364 536 380
rect 551 364 564 524
rect 594 420 607 524
rect 652 502 653 512
rect 668 502 681 512
rect 652 498 681 502
rect 686 498 716 524
rect 734 510 750 512
rect 822 510 875 524
rect 823 508 887 510
rect 930 508 945 524
rect 994 521 1024 524
rect 994 518 1030 521
rect 960 510 976 512
rect 734 498 749 502
rect 652 496 749 498
rect 777 496 945 508
rect 961 498 976 502
rect 994 499 1033 518
rect 1052 512 1059 513
rect 1058 505 1059 512
rect 1042 502 1043 505
rect 1058 502 1071 505
rect 994 498 1024 499
rect 1033 498 1039 499
rect 1042 498 1071 502
rect 961 497 1071 498
rect 961 496 1077 497
rect 636 488 687 496
rect 636 476 661 488
rect 668 476 687 488
rect 718 488 768 496
rect 718 480 734 488
rect 741 486 768 488
rect 777 486 998 496
rect 741 476 998 486
rect 1027 488 1077 496
rect 1027 479 1043 488
rect 636 468 687 476
rect 734 468 998 476
rect 1024 476 1043 479
rect 1050 476 1077 488
rect 1024 468 1077 476
rect 652 460 653 468
rect 668 460 681 468
rect 652 452 668 460
rect 649 445 668 448
rect 649 436 671 445
rect 622 426 671 436
rect 622 420 652 426
rect 671 421 676 426
rect 594 404 668 420
rect 686 412 716 468
rect 751 458 959 468
rect 994 464 1039 468
rect 1042 467 1043 468
rect 1058 467 1071 468
rect 777 428 966 458
rect 792 425 966 428
rect 785 422 966 425
rect 594 402 607 404
rect 622 402 656 404
rect 594 386 668 402
rect 695 398 708 412
rect 723 398 739 414
rect 785 409 796 422
rect 578 364 579 380
rect 594 364 607 386
rect 622 364 652 386
rect 695 382 757 398
rect 785 391 796 407
rect 801 402 811 422
rect 821 402 835 422
rect 838 409 847 422
rect 863 409 872 422
rect 801 391 835 402
rect 838 391 847 407
rect 863 391 872 407
rect 879 402 889 422
rect 899 402 913 422
rect 914 409 925 422
rect 879 391 913 402
rect 914 391 925 407
rect 971 398 987 414
rect 994 412 1024 464
rect 1058 460 1059 467
rect 1043 452 1059 460
rect 1030 420 1043 439
rect 1058 420 1088 436
rect 1030 404 1104 420
rect 1030 402 1043 404
rect 1058 402 1092 404
rect 695 380 708 382
rect 723 380 757 382
rect 695 364 757 380
rect 801 375 817 382
rect 879 375 909 386
rect 957 382 1003 398
rect 1030 386 1104 402
rect 957 380 991 382
rect 956 364 1003 380
rect 1030 364 1043 386
rect 1058 364 1088 386
rect 1115 364 1116 380
rect 1131 364 1144 524
rect 1174 420 1187 524
rect 1232 502 1233 512
rect 1248 502 1261 512
rect 1232 498 1261 502
rect 1266 498 1281 524
rect 1232 496 1281 498
rect 1216 488 1267 496
rect 1216 476 1241 488
rect 1248 476 1267 488
rect 1216 468 1267 476
rect 1232 460 1233 468
rect 1248 460 1261 468
rect 1232 452 1248 460
rect 1229 445 1248 448
rect 1229 436 1251 445
rect 1202 426 1251 436
rect 1202 420 1232 426
rect 1251 421 1256 426
rect 1174 404 1248 420
rect 1266 412 1281 468
rect 1174 402 1187 404
rect 1202 402 1236 404
rect 1174 386 1248 402
rect 1158 364 1159 380
rect 1174 364 1187 386
rect 1202 364 1232 386
rect 1275 364 1281 412
rect -8 356 33 364
rect -8 330 7 356
rect 14 330 33 356
rect 97 352 159 364
rect 171 352 246 364
rect 304 352 379 364
rect 391 352 422 364
rect 428 352 463 364
rect 97 350 259 352
rect -8 322 33 330
rect 115 326 128 350
rect 143 348 158 350
rect -2 312 -1 322
rect 14 312 27 322
rect 42 312 72 326
rect 115 312 158 326
rect 182 323 189 330
rect 192 326 259 350
rect 291 350 463 352
rect 261 328 289 332
rect 291 328 371 350
rect 392 348 407 350
rect 261 326 371 328
rect 192 322 371 326
rect 165 312 195 322
rect 197 312 350 322
rect 358 312 388 322
rect 392 312 422 326
rect 450 312 463 350
rect 535 356 570 364
rect 535 330 536 356
rect 543 330 570 356
rect 478 312 508 326
rect 535 322 570 330
rect 572 356 613 364
rect 572 330 587 356
rect 594 330 613 356
rect 677 352 739 364
rect 751 352 826 364
rect 884 352 959 364
rect 971 352 1002 364
rect 1008 352 1043 364
rect 677 350 839 352
rect 572 322 613 330
rect 695 326 708 350
rect 723 348 738 350
rect 535 312 536 322
rect 551 312 564 322
rect 578 312 579 322
rect 594 312 607 322
rect 622 312 652 326
rect 695 312 738 326
rect 762 323 769 330
rect 772 326 839 350
rect 871 350 1043 352
rect 841 328 869 332
rect 871 328 951 350
rect 972 348 987 350
rect 841 326 951 328
rect 772 322 951 326
rect 745 312 775 322
rect 777 312 930 322
rect 938 312 968 322
rect 972 312 1002 326
rect 1030 312 1043 350
rect 1115 356 1150 364
rect 1115 330 1116 356
rect 1123 330 1150 356
rect 1058 312 1088 326
rect 1115 322 1150 330
rect 1152 356 1193 364
rect 1152 330 1167 356
rect 1174 330 1193 356
rect 1257 350 1281 364
rect 1152 322 1193 330
rect 1115 312 1116 322
rect 1131 312 1144 322
rect 1158 312 1159 322
rect 1174 312 1187 322
rect 1202 312 1232 326
rect 1275 312 1281 350
rect -2 306 1281 312
rect -1 298 1281 306
rect 14 268 27 298
rect 42 280 72 298
rect 115 284 129 298
rect 165 284 385 298
rect 116 282 129 284
rect 82 270 97 282
rect 79 268 101 270
rect 106 268 136 282
rect 197 280 350 284
rect 179 268 371 280
rect 414 268 444 282
rect 450 268 463 298
rect 478 280 508 298
rect 551 268 564 298
rect 594 268 607 298
rect 622 280 652 298
rect 695 284 709 298
rect 745 284 965 298
rect 696 282 709 284
rect 662 270 677 282
rect 659 268 681 270
rect 686 268 716 282
rect 777 280 930 284
rect 759 268 951 280
rect 994 268 1024 282
rect 1030 268 1043 298
rect 1058 280 1088 298
rect 1131 268 1144 298
rect 1174 268 1187 298
rect 1202 280 1232 298
rect 1275 284 1281 298
rect 1276 282 1281 284
rect 1242 270 1257 282
rect 1239 268 1261 270
rect 1266 268 1281 282
rect -1 254 1281 268
rect 14 150 27 254
rect 72 232 73 242
rect 88 232 101 242
rect 72 228 101 232
rect 106 228 136 254
rect 154 240 170 242
rect 242 240 295 254
rect 243 238 307 240
rect 350 238 365 254
rect 414 251 444 254
rect 414 248 450 251
rect 380 240 396 242
rect 154 228 169 232
rect 72 226 169 228
rect 197 226 365 238
rect 381 228 396 232
rect 414 229 453 248
rect 472 242 479 243
rect 478 235 479 242
rect 462 232 463 235
rect 478 232 491 235
rect 414 228 444 229
rect 453 228 459 229
rect 462 228 491 232
rect 381 227 491 228
rect 381 226 497 227
rect 56 218 107 226
rect 56 206 81 218
rect 88 206 107 218
rect 138 218 188 226
rect 138 210 154 218
rect 161 216 188 218
rect 197 216 418 226
rect 161 206 418 216
rect 447 218 497 226
rect 447 209 463 218
rect 56 198 107 206
rect 154 198 418 206
rect 444 206 463 209
rect 470 206 497 218
rect 444 198 497 206
rect 72 190 73 198
rect 88 190 101 198
rect 72 182 88 190
rect 69 175 88 178
rect 69 166 91 175
rect 42 156 91 166
rect 42 150 72 156
rect 91 151 96 156
rect 14 134 88 150
rect 106 142 136 198
rect 171 188 379 198
rect 414 194 459 198
rect 462 197 463 198
rect 478 197 491 198
rect 197 158 386 188
rect 212 155 386 158
rect 205 152 386 155
rect 14 132 27 134
rect 42 132 76 134
rect 14 116 88 132
rect 115 128 128 142
rect 143 128 159 144
rect 205 139 216 152
rect -2 94 -1 110
rect 14 94 27 116
rect 42 94 72 116
rect 115 112 177 128
rect 205 121 216 137
rect 221 132 231 152
rect 241 132 255 152
rect 258 139 267 152
rect 283 139 292 152
rect 221 121 255 132
rect 258 121 267 137
rect 283 121 292 137
rect 299 132 309 152
rect 319 132 333 152
rect 334 139 345 152
rect 299 121 333 132
rect 334 121 345 137
rect 391 128 407 144
rect 414 142 444 194
rect 478 190 479 197
rect 463 182 479 190
rect 450 150 463 169
rect 478 150 508 166
rect 450 134 524 150
rect 450 132 463 134
rect 478 132 512 134
rect 115 110 128 112
rect 143 110 177 112
rect 115 94 177 110
rect 221 105 237 112
rect 299 105 329 116
rect 377 112 423 128
rect 450 116 524 132
rect 377 110 411 112
rect 376 94 423 110
rect 450 94 463 116
rect 478 94 508 116
rect 535 94 536 110
rect 551 94 564 254
rect 594 150 607 254
rect 652 232 653 242
rect 668 232 681 242
rect 652 228 681 232
rect 686 228 716 254
rect 734 240 750 242
rect 822 240 875 254
rect 823 238 887 240
rect 930 238 945 254
rect 994 251 1024 254
rect 994 248 1030 251
rect 960 240 976 242
rect 734 228 749 232
rect 652 226 749 228
rect 777 226 945 238
rect 961 228 976 232
rect 994 229 1033 248
rect 1052 242 1059 243
rect 1058 235 1059 242
rect 1042 232 1043 235
rect 1058 232 1071 235
rect 994 228 1024 229
rect 1033 228 1039 229
rect 1042 228 1071 232
rect 961 227 1071 228
rect 961 226 1077 227
rect 636 218 687 226
rect 636 206 661 218
rect 668 206 687 218
rect 718 218 768 226
rect 718 210 734 218
rect 741 216 768 218
rect 777 216 998 226
rect 741 206 998 216
rect 1027 218 1077 226
rect 1027 209 1043 218
rect 636 198 687 206
rect 734 198 998 206
rect 1024 206 1043 209
rect 1050 206 1077 218
rect 1024 198 1077 206
rect 652 190 653 198
rect 668 190 681 198
rect 652 182 668 190
rect 649 175 668 178
rect 649 166 671 175
rect 622 156 671 166
rect 622 150 652 156
rect 671 151 676 156
rect 594 134 668 150
rect 686 142 716 198
rect 751 188 959 198
rect 994 194 1039 198
rect 1042 197 1043 198
rect 1058 197 1071 198
rect 777 158 966 188
rect 792 155 966 158
rect 785 152 966 155
rect 594 132 607 134
rect 622 132 656 134
rect 594 116 668 132
rect 695 128 708 142
rect 723 128 739 144
rect 785 139 796 152
rect 578 94 579 110
rect 594 94 607 116
rect 622 94 652 116
rect 695 112 757 128
rect 785 121 796 137
rect 801 132 811 152
rect 821 132 835 152
rect 838 139 847 152
rect 863 139 872 152
rect 801 121 835 132
rect 838 121 847 137
rect 863 121 872 137
rect 879 132 889 152
rect 899 132 913 152
rect 914 139 925 152
rect 879 121 913 132
rect 914 121 925 137
rect 971 128 987 144
rect 994 142 1024 194
rect 1058 190 1059 197
rect 1043 182 1059 190
rect 1030 150 1043 169
rect 1058 150 1088 166
rect 1030 134 1104 150
rect 1030 132 1043 134
rect 1058 132 1092 134
rect 695 110 708 112
rect 723 110 757 112
rect 695 94 757 110
rect 801 105 817 112
rect 879 105 909 116
rect 957 112 1003 128
rect 1030 116 1104 132
rect 957 110 991 112
rect 956 94 1003 110
rect 1030 94 1043 116
rect 1058 94 1088 116
rect 1115 94 1116 110
rect 1131 94 1144 254
rect 1174 150 1187 254
rect 1232 232 1233 242
rect 1248 232 1261 242
rect 1232 228 1261 232
rect 1266 228 1281 254
rect 1232 226 1281 228
rect 1216 218 1267 226
rect 1216 206 1241 218
rect 1248 206 1267 218
rect 1216 198 1267 206
rect 1232 190 1233 198
rect 1248 190 1261 198
rect 1232 182 1248 190
rect 1229 175 1248 178
rect 1229 166 1251 175
rect 1202 156 1251 166
rect 1202 150 1232 156
rect 1251 151 1256 156
rect 1174 134 1248 150
rect 1266 142 1281 198
rect 1174 132 1187 134
rect 1202 132 1236 134
rect 1174 116 1248 132
rect 1158 94 1159 110
rect 1174 94 1187 116
rect 1202 94 1232 116
rect 1275 94 1281 142
rect -8 86 33 94
rect -8 60 7 86
rect 14 60 33 86
rect 97 82 159 94
rect 171 82 246 94
rect 304 82 379 94
rect 391 82 422 94
rect 428 82 463 94
rect 97 80 259 82
rect -8 52 33 60
rect 115 56 128 80
rect 143 78 158 80
rect -2 42 -1 52
rect 14 42 27 52
rect 42 42 72 56
rect 115 42 158 56
rect 182 53 189 60
rect 192 56 259 80
rect 291 80 463 82
rect 261 58 289 62
rect 291 58 371 80
rect 392 78 407 80
rect 261 56 371 58
rect 192 52 371 56
rect 165 42 195 52
rect 197 42 350 52
rect 358 42 388 52
rect 392 42 422 56
rect 450 42 463 80
rect 535 86 570 94
rect 535 60 536 86
rect 543 60 570 86
rect 478 42 508 56
rect 535 52 570 60
rect 572 86 613 94
rect 572 60 587 86
rect 594 60 613 86
rect 677 82 739 94
rect 751 82 826 94
rect 884 82 959 94
rect 971 82 1002 94
rect 1008 82 1043 94
rect 677 80 839 82
rect 572 52 613 60
rect 695 56 708 80
rect 723 78 738 80
rect 535 42 536 52
rect 551 42 564 52
rect 578 42 579 52
rect 594 42 607 52
rect 622 42 652 56
rect 695 42 738 56
rect 762 53 769 60
rect 772 56 839 80
rect 871 80 1043 82
rect 841 58 869 62
rect 871 58 951 80
rect 972 78 987 80
rect 841 56 951 58
rect 772 52 951 56
rect 745 42 775 52
rect 777 42 930 52
rect 938 42 968 52
rect 972 42 1002 56
rect 1030 42 1043 80
rect 1115 86 1150 94
rect 1115 60 1116 86
rect 1123 60 1150 86
rect 1058 42 1088 56
rect 1115 52 1150 60
rect 1152 86 1193 94
rect 1152 60 1167 86
rect 1174 60 1193 86
rect 1257 80 1281 94
rect 1152 52 1193 60
rect 1115 42 1116 52
rect 1131 42 1144 52
rect 1158 42 1159 52
rect 1174 42 1187 52
rect 1202 42 1232 56
rect 1275 42 1281 80
rect -2 36 1281 42
rect -1 28 1281 36
rect 14 -2 27 28
rect 42 10 72 28
rect 115 14 129 28
rect 165 14 385 28
rect 116 12 129 14
rect 82 0 97 12
rect 79 -2 101 0
rect 106 -2 136 12
rect 197 10 350 14
rect 179 -2 371 10
rect 414 -2 444 12
rect 450 -2 463 28
rect 478 10 508 28
rect 551 -2 564 28
rect 594 -2 607 28
rect 622 10 652 28
rect 695 14 709 28
rect 745 14 965 28
rect 696 12 709 14
rect 662 0 677 12
rect 659 -2 681 0
rect 686 -2 716 12
rect 777 10 930 14
rect 759 -2 951 10
rect 994 -2 1024 12
rect 1030 -2 1043 28
rect 1058 10 1088 28
rect 1131 -2 1144 28
rect 1174 -2 1187 28
rect 1202 10 1232 28
rect 1275 14 1281 28
rect 1276 12 1281 14
rect 1242 0 1257 12
rect 1239 -2 1261 0
rect 1266 -2 1281 12
rect -1 -16 1281 -2
rect 14 -120 27 -16
rect 72 -38 73 -28
rect 88 -38 101 -28
rect 72 -42 101 -38
rect 106 -42 136 -16
rect 154 -30 170 -28
rect 242 -30 295 -16
rect 243 -32 307 -30
rect 350 -32 365 -16
rect 414 -19 444 -16
rect 414 -22 450 -19
rect 380 -30 396 -28
rect 154 -42 169 -38
rect 72 -44 169 -42
rect 197 -44 365 -32
rect 381 -42 396 -38
rect 414 -41 453 -22
rect 472 -28 479 -27
rect 478 -35 479 -28
rect 462 -38 463 -35
rect 478 -38 491 -35
rect 414 -42 444 -41
rect 453 -42 459 -41
rect 462 -42 491 -38
rect 381 -43 491 -42
rect 381 -44 497 -43
rect 56 -52 107 -44
rect 56 -64 81 -52
rect 88 -64 107 -52
rect 138 -52 188 -44
rect 138 -60 154 -52
rect 161 -54 188 -52
rect 197 -54 418 -44
rect 161 -64 418 -54
rect 447 -52 497 -44
rect 447 -61 463 -52
rect 56 -72 107 -64
rect 154 -72 418 -64
rect 444 -64 463 -61
rect 470 -64 497 -52
rect 444 -72 497 -64
rect 72 -80 73 -72
rect 88 -80 101 -72
rect 72 -88 88 -80
rect 69 -95 88 -92
rect 69 -104 91 -95
rect 42 -114 91 -104
rect 42 -120 72 -114
rect 91 -119 96 -114
rect 14 -136 88 -120
rect 106 -128 136 -72
rect 171 -82 379 -72
rect 414 -76 459 -72
rect 462 -73 463 -72
rect 478 -73 491 -72
rect 197 -112 386 -82
rect 212 -115 386 -112
rect 205 -118 386 -115
rect 14 -138 27 -136
rect 42 -138 76 -136
rect 14 -154 88 -138
rect 115 -142 128 -128
rect 143 -142 159 -126
rect 205 -131 216 -118
rect -2 -176 -1 -160
rect 14 -176 27 -154
rect 42 -176 72 -154
rect 115 -158 177 -142
rect 205 -149 216 -133
rect 221 -138 231 -118
rect 241 -138 255 -118
rect 258 -131 267 -118
rect 283 -131 292 -118
rect 221 -149 255 -138
rect 258 -149 267 -133
rect 283 -149 292 -133
rect 299 -138 309 -118
rect 319 -138 333 -118
rect 334 -131 345 -118
rect 299 -149 333 -138
rect 334 -149 345 -133
rect 391 -142 407 -126
rect 414 -128 444 -76
rect 478 -80 479 -73
rect 463 -88 479 -80
rect 450 -120 463 -101
rect 478 -120 508 -104
rect 450 -136 524 -120
rect 450 -138 463 -136
rect 478 -138 512 -136
rect 115 -160 128 -158
rect 143 -160 177 -158
rect 115 -176 177 -160
rect 221 -165 237 -158
rect 299 -165 329 -154
rect 377 -158 423 -142
rect 450 -154 524 -138
rect 377 -160 411 -158
rect 376 -176 423 -160
rect 450 -176 463 -154
rect 478 -176 508 -154
rect 535 -176 536 -160
rect 551 -176 564 -16
rect 594 -120 607 -16
rect 652 -38 653 -28
rect 668 -38 681 -28
rect 652 -42 681 -38
rect 686 -42 716 -16
rect 734 -30 750 -28
rect 822 -30 875 -16
rect 823 -32 887 -30
rect 930 -32 945 -16
rect 994 -19 1024 -16
rect 994 -22 1030 -19
rect 960 -30 976 -28
rect 734 -42 749 -38
rect 652 -44 749 -42
rect 777 -44 945 -32
rect 961 -42 976 -38
rect 994 -41 1033 -22
rect 1052 -28 1059 -27
rect 1058 -35 1059 -28
rect 1042 -38 1043 -35
rect 1058 -38 1071 -35
rect 994 -42 1024 -41
rect 1033 -42 1039 -41
rect 1042 -42 1071 -38
rect 961 -43 1071 -42
rect 961 -44 1077 -43
rect 636 -52 687 -44
rect 636 -64 661 -52
rect 668 -64 687 -52
rect 718 -52 768 -44
rect 718 -60 734 -52
rect 741 -54 768 -52
rect 777 -54 998 -44
rect 741 -64 998 -54
rect 1027 -52 1077 -44
rect 1027 -61 1043 -52
rect 636 -72 687 -64
rect 734 -72 998 -64
rect 1024 -64 1043 -61
rect 1050 -64 1077 -52
rect 1024 -72 1077 -64
rect 652 -80 653 -72
rect 668 -80 681 -72
rect 652 -88 668 -80
rect 649 -95 668 -92
rect 649 -104 671 -95
rect 622 -114 671 -104
rect 622 -120 652 -114
rect 671 -119 676 -114
rect 594 -136 668 -120
rect 686 -128 716 -72
rect 751 -82 959 -72
rect 994 -76 1039 -72
rect 1042 -73 1043 -72
rect 1058 -73 1071 -72
rect 777 -112 966 -82
rect 792 -115 966 -112
rect 785 -118 966 -115
rect 594 -138 607 -136
rect 622 -138 656 -136
rect 594 -154 668 -138
rect 695 -142 708 -128
rect 723 -142 739 -126
rect 785 -131 796 -118
rect 578 -176 579 -160
rect 594 -176 607 -154
rect 622 -176 652 -154
rect 695 -158 757 -142
rect 785 -149 796 -133
rect 801 -138 811 -118
rect 821 -138 835 -118
rect 838 -131 847 -118
rect 863 -131 872 -118
rect 801 -149 835 -138
rect 838 -149 847 -133
rect 863 -149 872 -133
rect 879 -138 889 -118
rect 899 -138 913 -118
rect 914 -131 925 -118
rect 879 -149 913 -138
rect 914 -149 925 -133
rect 971 -142 987 -126
rect 994 -128 1024 -76
rect 1058 -80 1059 -73
rect 1043 -88 1059 -80
rect 1030 -120 1043 -101
rect 1058 -120 1088 -104
rect 1030 -136 1104 -120
rect 1030 -138 1043 -136
rect 1058 -138 1092 -136
rect 695 -160 708 -158
rect 723 -160 757 -158
rect 695 -176 757 -160
rect 801 -165 817 -158
rect 879 -165 909 -154
rect 957 -158 1003 -142
rect 1030 -154 1104 -138
rect 957 -160 991 -158
rect 956 -176 1003 -160
rect 1030 -176 1043 -154
rect 1058 -176 1088 -154
rect 1115 -176 1116 -160
rect 1131 -176 1144 -16
rect 1174 -120 1187 -16
rect 1232 -38 1233 -28
rect 1248 -38 1261 -28
rect 1232 -42 1261 -38
rect 1266 -42 1281 -16
rect 1232 -44 1281 -42
rect 1216 -52 1267 -44
rect 1216 -64 1241 -52
rect 1248 -64 1267 -52
rect 1321 -64 1551 -62
rect 1216 -72 1267 -64
rect 1314 -72 1551 -64
rect 1232 -80 1233 -72
rect 1248 -80 1261 -72
rect 1232 -88 1248 -80
rect 1229 -95 1248 -92
rect 1229 -104 1251 -95
rect 1202 -114 1251 -104
rect 1202 -120 1232 -114
rect 1251 -119 1256 -114
rect 1174 -136 1248 -120
rect 1266 -128 1296 -72
rect 1331 -82 1539 -72
rect 1357 -112 1546 -82
rect 1372 -115 1546 -112
rect 1365 -118 1546 -115
rect 1174 -138 1187 -136
rect 1202 -138 1236 -136
rect 1174 -154 1248 -138
rect 1275 -142 1288 -128
rect 1303 -142 1319 -126
rect 1365 -131 1376 -118
rect 1158 -176 1159 -160
rect 1174 -176 1187 -154
rect 1202 -176 1232 -154
rect 1275 -158 1337 -142
rect 1365 -149 1376 -133
rect 1381 -138 1391 -118
rect 1401 -138 1415 -118
rect 1418 -131 1427 -118
rect 1443 -131 1452 -118
rect 1381 -149 1415 -138
rect 1418 -149 1427 -133
rect 1443 -149 1452 -133
rect 1459 -138 1469 -118
rect 1479 -138 1493 -118
rect 1494 -131 1505 -118
rect 1459 -149 1493 -138
rect 1494 -149 1505 -133
rect 1275 -160 1288 -158
rect 1303 -160 1337 -158
rect 1275 -176 1337 -160
rect 1381 -165 1397 -158
rect 1459 -165 1489 -154
rect 1537 -160 1551 -142
rect 1536 -176 1551 -160
rect -8 -184 33 -176
rect -8 -210 7 -184
rect 14 -210 33 -184
rect 97 -188 159 -176
rect 171 -188 246 -176
rect 304 -188 379 -176
rect 391 -188 422 -176
rect 428 -188 463 -176
rect 97 -190 259 -188
rect -8 -218 33 -210
rect 115 -214 128 -190
rect 143 -192 158 -190
rect -2 -228 -1 -218
rect 14 -228 27 -218
rect 42 -228 72 -214
rect 115 -228 158 -214
rect 182 -217 189 -210
rect 192 -214 259 -190
rect 291 -190 463 -188
rect 261 -212 289 -208
rect 291 -212 371 -190
rect 392 -192 407 -190
rect 261 -214 371 -212
rect 192 -218 371 -214
rect 165 -228 195 -218
rect 197 -228 350 -218
rect 358 -228 388 -218
rect 392 -228 422 -214
rect 450 -228 463 -190
rect 535 -184 570 -176
rect 535 -210 536 -184
rect 543 -210 570 -184
rect 478 -228 508 -214
rect 535 -218 570 -210
rect 572 -184 613 -176
rect 572 -210 587 -184
rect 594 -210 613 -184
rect 677 -188 739 -176
rect 751 -188 826 -176
rect 884 -188 959 -176
rect 971 -188 1002 -176
rect 1008 -188 1043 -176
rect 677 -190 839 -188
rect 572 -218 613 -210
rect 695 -214 708 -190
rect 723 -192 738 -190
rect 535 -228 536 -218
rect 551 -228 564 -218
rect 578 -228 579 -218
rect 594 -228 607 -218
rect 622 -228 652 -214
rect 695 -228 738 -214
rect 762 -217 769 -210
rect 772 -214 839 -190
rect 871 -190 1043 -188
rect 841 -212 869 -208
rect 871 -212 951 -190
rect 972 -192 987 -190
rect 841 -214 951 -212
rect 772 -218 951 -214
rect 745 -228 775 -218
rect 777 -228 930 -218
rect 938 -228 968 -218
rect 972 -228 1002 -214
rect 1030 -228 1043 -190
rect 1115 -184 1150 -176
rect 1115 -210 1116 -184
rect 1123 -210 1150 -184
rect 1058 -228 1088 -214
rect 1115 -218 1150 -210
rect 1152 -184 1193 -176
rect 1152 -210 1167 -184
rect 1174 -210 1193 -184
rect 1257 -188 1319 -176
rect 1331 -188 1406 -176
rect 1464 -188 1539 -176
rect 1257 -190 1419 -188
rect 1152 -218 1193 -210
rect 1275 -214 1288 -190
rect 1303 -192 1318 -190
rect 1115 -228 1116 -218
rect 1131 -228 1144 -218
rect 1158 -228 1159 -218
rect 1174 -228 1187 -218
rect 1202 -228 1232 -214
rect 1275 -228 1318 -214
rect 1342 -217 1349 -210
rect 1352 -214 1419 -190
rect 1451 -190 1551 -188
rect 1421 -212 1449 -208
rect 1451 -212 1531 -190
rect 1421 -214 1531 -212
rect 1352 -218 1531 -214
rect 1325 -228 1355 -218
rect 1357 -228 1510 -218
rect 1518 -228 1548 -218
rect -2 -234 1551 -228
rect -1 -242 1551 -234
rect 14 -272 27 -242
rect 42 -260 72 -242
rect 115 -256 129 -242
rect 165 -256 385 -242
rect 116 -258 129 -256
rect 82 -270 97 -258
rect 79 -272 101 -270
rect 106 -272 136 -258
rect 197 -260 350 -256
rect 179 -272 371 -260
rect 414 -272 444 -258
rect 450 -272 463 -242
rect 478 -260 508 -242
rect 551 -272 564 -242
rect 594 -272 607 -242
rect 622 -260 652 -242
rect 695 -256 709 -242
rect 745 -256 965 -242
rect 696 -258 709 -256
rect 662 -270 677 -258
rect 659 -272 681 -270
rect 686 -272 716 -258
rect 777 -260 930 -256
rect 759 -272 951 -260
rect 994 -272 1024 -258
rect 1030 -272 1043 -242
rect 1058 -260 1088 -242
rect 1131 -272 1144 -242
rect 1174 -272 1187 -242
rect 1202 -260 1232 -242
rect 1275 -256 1289 -242
rect 1325 -256 1545 -242
rect 1276 -258 1289 -256
rect 1242 -270 1257 -258
rect 1239 -272 1261 -270
rect 1266 -272 1296 -258
rect 1357 -260 1510 -256
rect 1339 -272 1531 -260
rect -1 -286 1551 -272
rect 14 -390 27 -286
rect 72 -308 73 -298
rect 88 -308 101 -298
rect 72 -312 101 -308
rect 106 -312 136 -286
rect 154 -300 170 -298
rect 242 -300 295 -286
rect 243 -302 307 -300
rect 350 -302 365 -286
rect 414 -289 444 -286
rect 414 -292 450 -289
rect 380 -300 396 -298
rect 154 -312 169 -308
rect 72 -314 169 -312
rect 197 -314 365 -302
rect 381 -312 396 -308
rect 414 -311 453 -292
rect 472 -298 479 -297
rect 478 -305 479 -298
rect 462 -308 463 -305
rect 478 -308 491 -305
rect 414 -312 444 -311
rect 453 -312 459 -311
rect 462 -312 491 -308
rect 381 -313 491 -312
rect 381 -314 497 -313
rect 56 -322 107 -314
rect 56 -334 81 -322
rect 88 -334 107 -322
rect 138 -322 188 -314
rect 138 -330 154 -322
rect 161 -324 188 -322
rect 197 -324 418 -314
rect 161 -334 418 -324
rect 447 -322 497 -314
rect 447 -331 463 -322
rect 56 -342 107 -334
rect 154 -342 418 -334
rect 444 -334 463 -331
rect 470 -334 497 -322
rect 444 -342 497 -334
rect 72 -350 73 -342
rect 88 -350 101 -342
rect 72 -358 88 -350
rect 69 -365 88 -362
rect 69 -374 91 -365
rect 42 -384 91 -374
rect 42 -390 72 -384
rect 91 -389 96 -384
rect 14 -406 88 -390
rect 106 -398 136 -342
rect 171 -352 379 -342
rect 414 -346 459 -342
rect 462 -343 463 -342
rect 478 -343 491 -342
rect 197 -382 386 -352
rect 212 -385 386 -382
rect 205 -388 386 -385
rect 14 -408 27 -406
rect 42 -408 76 -406
rect 14 -424 88 -408
rect 115 -412 128 -398
rect 143 -412 159 -396
rect 205 -401 216 -388
rect -2 -446 -1 -430
rect 14 -446 27 -424
rect 42 -446 72 -424
rect 115 -428 177 -412
rect 205 -419 216 -403
rect 221 -408 231 -388
rect 241 -408 255 -388
rect 258 -401 267 -388
rect 283 -401 292 -388
rect 221 -419 255 -408
rect 258 -419 267 -403
rect 283 -419 292 -403
rect 299 -408 309 -388
rect 319 -408 333 -388
rect 334 -401 345 -388
rect 299 -419 333 -408
rect 334 -419 345 -403
rect 391 -412 407 -396
rect 414 -398 444 -346
rect 478 -350 479 -343
rect 463 -358 479 -350
rect 450 -390 463 -371
rect 478 -390 508 -374
rect 450 -406 524 -390
rect 450 -408 463 -406
rect 478 -408 512 -406
rect 115 -430 128 -428
rect 143 -430 177 -428
rect 115 -446 177 -430
rect 221 -435 237 -428
rect 299 -435 329 -424
rect 377 -428 423 -412
rect 450 -424 524 -408
rect 377 -430 411 -428
rect 376 -446 423 -430
rect 450 -446 463 -424
rect 478 -446 508 -424
rect 535 -446 536 -430
rect 551 -446 564 -286
rect 594 -390 607 -286
rect 652 -308 653 -298
rect 668 -308 681 -298
rect 652 -312 681 -308
rect 686 -312 716 -286
rect 734 -300 750 -298
rect 822 -300 875 -286
rect 823 -302 887 -300
rect 930 -302 945 -286
rect 994 -289 1024 -286
rect 994 -292 1030 -289
rect 960 -300 976 -298
rect 734 -312 749 -308
rect 652 -314 749 -312
rect 777 -314 945 -302
rect 961 -312 976 -308
rect 994 -311 1033 -292
rect 1052 -298 1059 -297
rect 1058 -305 1059 -298
rect 1042 -308 1043 -305
rect 1058 -308 1071 -305
rect 994 -312 1024 -311
rect 1033 -312 1039 -311
rect 1042 -312 1071 -308
rect 961 -313 1071 -312
rect 961 -314 1077 -313
rect 636 -322 687 -314
rect 636 -334 661 -322
rect 668 -334 687 -322
rect 718 -322 768 -314
rect 718 -330 734 -322
rect 741 -324 768 -322
rect 777 -324 998 -314
rect 741 -334 998 -324
rect 1027 -322 1077 -314
rect 1027 -331 1043 -322
rect 636 -342 687 -334
rect 734 -342 998 -334
rect 1024 -334 1043 -331
rect 1050 -334 1077 -322
rect 1024 -342 1077 -334
rect 652 -350 653 -342
rect 668 -350 681 -342
rect 652 -358 668 -350
rect 649 -365 668 -362
rect 649 -374 671 -365
rect 622 -384 671 -374
rect 622 -390 652 -384
rect 671 -389 676 -384
rect 594 -406 668 -390
rect 686 -398 716 -342
rect 751 -352 959 -342
rect 994 -346 1039 -342
rect 1042 -343 1043 -342
rect 1058 -343 1071 -342
rect 777 -382 966 -352
rect 792 -385 966 -382
rect 785 -388 966 -385
rect 594 -408 607 -406
rect 622 -408 656 -406
rect 594 -424 668 -408
rect 695 -412 708 -398
rect 723 -412 739 -396
rect 785 -401 796 -388
rect 578 -446 579 -430
rect 594 -446 607 -424
rect 622 -446 652 -424
rect 695 -428 757 -412
rect 785 -419 796 -403
rect 801 -408 811 -388
rect 821 -408 835 -388
rect 838 -401 847 -388
rect 863 -401 872 -388
rect 801 -419 835 -408
rect 838 -419 847 -403
rect 863 -419 872 -403
rect 879 -408 889 -388
rect 899 -408 913 -388
rect 914 -401 925 -388
rect 879 -419 913 -408
rect 914 -419 925 -403
rect 971 -412 987 -396
rect 994 -398 1024 -346
rect 1058 -350 1059 -343
rect 1043 -358 1059 -350
rect 1030 -390 1043 -371
rect 1058 -390 1088 -374
rect 1030 -406 1104 -390
rect 1030 -408 1043 -406
rect 1058 -408 1092 -406
rect 695 -430 708 -428
rect 723 -430 757 -428
rect 695 -446 757 -430
rect 801 -435 817 -428
rect 879 -435 909 -424
rect 957 -428 1003 -412
rect 1030 -424 1104 -408
rect 957 -430 991 -428
rect 956 -446 1003 -430
rect 1030 -446 1043 -424
rect 1058 -446 1088 -424
rect 1115 -446 1116 -430
rect 1131 -446 1144 -286
rect 1174 -390 1187 -286
rect 1232 -308 1233 -298
rect 1248 -308 1261 -298
rect 1232 -312 1261 -308
rect 1266 -312 1296 -286
rect 1314 -300 1330 -298
rect 1402 -300 1455 -286
rect 1403 -302 1467 -300
rect 1510 -302 1525 -286
rect 1540 -300 1551 -298
rect 1314 -312 1329 -308
rect 1232 -314 1329 -312
rect 1357 -314 1525 -302
rect 1541 -314 1551 -308
rect 1216 -322 1267 -314
rect 1216 -334 1241 -322
rect 1248 -334 1267 -322
rect 1298 -322 1348 -314
rect 1298 -330 1314 -322
rect 1321 -324 1348 -322
rect 1357 -324 1551 -314
rect 1321 -334 1551 -324
rect 1216 -342 1267 -334
rect 1314 -342 1551 -334
rect 1232 -350 1233 -342
rect 1248 -350 1261 -342
rect 1232 -358 1248 -350
rect 1229 -365 1248 -362
rect 1229 -374 1251 -365
rect 1202 -384 1251 -374
rect 1202 -390 1232 -384
rect 1251 -389 1256 -384
rect 1174 -406 1248 -390
rect 1266 -398 1296 -342
rect 1331 -352 1539 -342
rect 1357 -382 1546 -352
rect 1372 -385 1546 -382
rect 1365 -388 1546 -385
rect 1174 -408 1187 -406
rect 1202 -408 1236 -406
rect 1174 -424 1248 -408
rect 1275 -412 1288 -398
rect 1303 -412 1319 -396
rect 1365 -401 1376 -388
rect 1158 -446 1159 -430
rect 1174 -446 1187 -424
rect 1202 -446 1232 -424
rect 1275 -428 1337 -412
rect 1365 -419 1376 -403
rect 1381 -408 1391 -388
rect 1401 -408 1415 -388
rect 1418 -401 1427 -388
rect 1443 -401 1452 -388
rect 1381 -419 1415 -408
rect 1418 -419 1427 -403
rect 1443 -419 1452 -403
rect 1459 -408 1469 -388
rect 1479 -408 1493 -388
rect 1494 -401 1505 -388
rect 1459 -419 1493 -408
rect 1494 -419 1505 -403
rect 1275 -430 1288 -428
rect 1303 -430 1337 -428
rect 1275 -446 1337 -430
rect 1381 -435 1397 -428
rect 1459 -435 1489 -424
rect 1537 -430 1551 -412
rect 1536 -446 1551 -430
rect -8 -454 33 -446
rect -8 -480 7 -454
rect 14 -480 33 -454
rect 97 -458 159 -446
rect 171 -458 246 -446
rect 304 -458 379 -446
rect 391 -458 422 -446
rect 428 -458 463 -446
rect 97 -460 259 -458
rect -8 -488 33 -480
rect 115 -484 128 -460
rect 143 -462 158 -460
rect -2 -498 -1 -488
rect 14 -498 27 -488
rect 42 -498 72 -484
rect 115 -498 158 -484
rect 182 -487 189 -480
rect 192 -484 259 -460
rect 291 -460 463 -458
rect 261 -482 289 -478
rect 291 -482 371 -460
rect 392 -462 407 -460
rect 261 -484 371 -482
rect 192 -488 371 -484
rect 165 -498 195 -488
rect 197 -498 350 -488
rect 358 -498 388 -488
rect 392 -498 422 -484
rect 450 -498 463 -460
rect 535 -454 570 -446
rect 535 -480 536 -454
rect 543 -480 570 -454
rect 478 -498 508 -484
rect 535 -488 570 -480
rect 572 -454 613 -446
rect 572 -480 587 -454
rect 594 -480 613 -454
rect 677 -458 739 -446
rect 751 -458 826 -446
rect 884 -458 959 -446
rect 971 -458 1002 -446
rect 1008 -458 1043 -446
rect 677 -460 839 -458
rect 572 -488 613 -480
rect 695 -484 708 -460
rect 723 -462 738 -460
rect 535 -498 536 -488
rect 551 -498 564 -488
rect 578 -498 579 -488
rect 594 -498 607 -488
rect 622 -498 652 -484
rect 695 -498 738 -484
rect 762 -487 769 -480
rect 772 -484 839 -460
rect 871 -460 1043 -458
rect 841 -482 869 -478
rect 871 -482 951 -460
rect 972 -462 987 -460
rect 841 -484 951 -482
rect 772 -488 951 -484
rect 745 -498 775 -488
rect 777 -498 930 -488
rect 938 -498 968 -488
rect 972 -498 1002 -484
rect 1030 -498 1043 -460
rect 1115 -454 1150 -446
rect 1115 -480 1116 -454
rect 1123 -480 1150 -454
rect 1058 -498 1088 -484
rect 1115 -488 1150 -480
rect 1152 -454 1193 -446
rect 1152 -480 1167 -454
rect 1174 -480 1193 -454
rect 1257 -458 1319 -446
rect 1331 -458 1406 -446
rect 1464 -458 1539 -446
rect 1257 -460 1419 -458
rect 1152 -488 1193 -480
rect 1275 -484 1288 -460
rect 1303 -462 1318 -460
rect 1115 -498 1116 -488
rect 1131 -498 1144 -488
rect 1158 -498 1159 -488
rect 1174 -498 1187 -488
rect 1202 -498 1232 -484
rect 1275 -498 1318 -484
rect 1342 -487 1349 -480
rect 1352 -484 1419 -460
rect 1451 -460 1551 -458
rect 1421 -482 1449 -478
rect 1451 -482 1531 -460
rect 1421 -484 1531 -482
rect 1352 -488 1531 -484
rect 1325 -498 1355 -488
rect 1357 -498 1510 -488
rect 1518 -498 1548 -488
rect -2 -504 1551 -498
rect -1 -512 1551 -504
rect 14 -542 27 -512
rect 42 -530 72 -512
rect 115 -526 129 -512
rect 165 -526 385 -512
rect 116 -528 129 -526
rect 82 -540 97 -528
rect 79 -542 101 -540
rect 106 -542 136 -528
rect 197 -530 350 -526
rect 179 -542 371 -530
rect 414 -542 444 -528
rect 450 -542 463 -512
rect 478 -530 508 -512
rect 551 -542 564 -512
rect 594 -542 607 -512
rect 622 -530 652 -512
rect 695 -526 709 -512
rect 745 -526 965 -512
rect 696 -528 709 -526
rect 662 -540 677 -528
rect 659 -542 681 -540
rect 686 -542 716 -528
rect 777 -530 930 -526
rect 759 -542 951 -530
rect 994 -542 1024 -528
rect 1030 -542 1043 -512
rect 1058 -530 1088 -512
rect 1131 -542 1144 -512
rect 1174 -542 1187 -512
rect 1202 -530 1232 -512
rect 1275 -526 1289 -512
rect 1325 -526 1545 -512
rect 1276 -528 1289 -526
rect 1242 -540 1257 -528
rect 1239 -542 1261 -540
rect 1266 -542 1296 -528
rect 1357 -530 1510 -526
rect 1339 -542 1531 -530
rect -1 -556 1551 -542
rect 14 -660 27 -556
rect 72 -578 73 -568
rect 88 -578 101 -568
rect 72 -582 101 -578
rect 106 -582 136 -556
rect 154 -570 170 -568
rect 242 -570 295 -556
rect 243 -572 307 -570
rect 350 -572 365 -556
rect 414 -559 444 -556
rect 414 -562 450 -559
rect 380 -570 396 -568
rect 154 -582 169 -578
rect 72 -584 169 -582
rect 197 -584 365 -572
rect 381 -582 396 -578
rect 414 -581 453 -562
rect 472 -568 479 -567
rect 478 -575 479 -568
rect 462 -578 463 -575
rect 478 -578 491 -575
rect 414 -582 444 -581
rect 453 -582 459 -581
rect 462 -582 491 -578
rect 381 -583 491 -582
rect 381 -584 497 -583
rect 56 -592 107 -584
rect 56 -604 81 -592
rect 88 -604 107 -592
rect 138 -592 188 -584
rect 138 -600 154 -592
rect 161 -594 188 -592
rect 197 -594 418 -584
rect 161 -604 418 -594
rect 447 -592 497 -584
rect 447 -601 463 -592
rect 56 -612 107 -604
rect 154 -612 418 -604
rect 444 -604 463 -601
rect 470 -604 497 -592
rect 444 -612 497 -604
rect 72 -620 73 -612
rect 88 -620 101 -612
rect 72 -628 88 -620
rect 69 -635 88 -632
rect 69 -644 91 -635
rect 42 -654 91 -644
rect 42 -660 72 -654
rect 91 -659 96 -654
rect 14 -676 88 -660
rect 106 -668 136 -612
rect 171 -622 379 -612
rect 414 -616 459 -612
rect 462 -613 463 -612
rect 478 -613 491 -612
rect 197 -652 386 -622
rect 212 -655 386 -652
rect 205 -658 386 -655
rect 14 -678 27 -676
rect 42 -678 76 -676
rect 14 -694 88 -678
rect 115 -682 128 -668
rect 143 -682 159 -666
rect 205 -671 216 -658
rect -2 -716 -1 -700
rect 14 -716 27 -694
rect 42 -716 72 -694
rect 115 -698 177 -682
rect 205 -689 216 -673
rect 221 -678 231 -658
rect 241 -678 255 -658
rect 258 -671 267 -658
rect 283 -671 292 -658
rect 221 -689 255 -678
rect 258 -689 267 -673
rect 283 -689 292 -673
rect 299 -678 309 -658
rect 319 -678 333 -658
rect 334 -671 345 -658
rect 299 -689 333 -678
rect 334 -689 345 -673
rect 391 -682 407 -666
rect 414 -668 444 -616
rect 478 -620 479 -613
rect 463 -628 479 -620
rect 450 -660 463 -641
rect 478 -660 508 -644
rect 450 -676 524 -660
rect 450 -678 463 -676
rect 478 -678 512 -676
rect 115 -700 128 -698
rect 143 -700 177 -698
rect 115 -716 177 -700
rect 221 -705 237 -698
rect 299 -705 329 -694
rect 377 -698 423 -682
rect 450 -694 524 -678
rect 377 -700 411 -698
rect 376 -716 423 -700
rect 450 -716 463 -694
rect 478 -716 508 -694
rect 535 -716 536 -700
rect 551 -716 564 -556
rect 594 -660 607 -556
rect 652 -578 653 -568
rect 668 -578 681 -568
rect 652 -582 681 -578
rect 686 -582 716 -556
rect 734 -570 750 -568
rect 822 -570 875 -556
rect 823 -572 887 -570
rect 930 -572 945 -556
rect 994 -559 1024 -556
rect 994 -562 1030 -559
rect 960 -570 976 -568
rect 734 -582 749 -578
rect 652 -584 749 -582
rect 777 -584 945 -572
rect 961 -582 976 -578
rect 994 -581 1033 -562
rect 1052 -568 1059 -567
rect 1058 -575 1059 -568
rect 1042 -578 1043 -575
rect 1058 -578 1071 -575
rect 994 -582 1024 -581
rect 1033 -582 1039 -581
rect 1042 -582 1071 -578
rect 961 -583 1071 -582
rect 961 -584 1077 -583
rect 636 -592 687 -584
rect 636 -604 661 -592
rect 668 -604 687 -592
rect 718 -592 768 -584
rect 718 -600 734 -592
rect 741 -594 768 -592
rect 777 -594 998 -584
rect 741 -604 998 -594
rect 1027 -592 1077 -584
rect 1027 -601 1043 -592
rect 636 -612 687 -604
rect 734 -612 998 -604
rect 1024 -604 1043 -601
rect 1050 -604 1077 -592
rect 1024 -612 1077 -604
rect 652 -620 653 -612
rect 668 -620 681 -612
rect 652 -628 668 -620
rect 649 -635 668 -632
rect 649 -644 671 -635
rect 622 -654 671 -644
rect 622 -660 652 -654
rect 671 -659 676 -654
rect 594 -676 668 -660
rect 686 -668 716 -612
rect 751 -622 959 -612
rect 994 -616 1039 -612
rect 1042 -613 1043 -612
rect 1058 -613 1071 -612
rect 777 -652 966 -622
rect 792 -655 966 -652
rect 785 -658 966 -655
rect 594 -678 607 -676
rect 622 -678 656 -676
rect 594 -694 668 -678
rect 695 -682 708 -668
rect 723 -682 739 -666
rect 785 -671 796 -658
rect 578 -716 579 -700
rect 594 -716 607 -694
rect 622 -716 652 -694
rect 695 -698 757 -682
rect 785 -689 796 -673
rect 801 -678 811 -658
rect 821 -678 835 -658
rect 838 -671 847 -658
rect 863 -671 872 -658
rect 801 -689 835 -678
rect 838 -689 847 -673
rect 863 -689 872 -673
rect 879 -678 889 -658
rect 899 -678 913 -658
rect 914 -671 925 -658
rect 879 -689 913 -678
rect 914 -689 925 -673
rect 971 -682 987 -666
rect 994 -668 1024 -616
rect 1058 -620 1059 -613
rect 1043 -628 1059 -620
rect 1030 -660 1043 -641
rect 1058 -660 1088 -644
rect 1030 -676 1104 -660
rect 1030 -678 1043 -676
rect 1058 -678 1092 -676
rect 695 -700 708 -698
rect 723 -700 757 -698
rect 695 -716 757 -700
rect 801 -705 817 -698
rect 879 -705 909 -694
rect 957 -698 1003 -682
rect 1030 -694 1104 -678
rect 957 -700 991 -698
rect 956 -716 1003 -700
rect 1030 -716 1043 -694
rect 1058 -716 1088 -694
rect 1115 -716 1116 -700
rect 1131 -716 1144 -556
rect 1174 -660 1187 -556
rect 1232 -578 1233 -568
rect 1248 -578 1261 -568
rect 1232 -582 1261 -578
rect 1266 -582 1296 -556
rect 1314 -570 1330 -568
rect 1402 -570 1455 -556
rect 1403 -572 1467 -570
rect 1510 -572 1525 -556
rect 1540 -570 1551 -568
rect 1314 -582 1329 -578
rect 1232 -584 1329 -582
rect 1357 -584 1525 -572
rect 1541 -584 1551 -578
rect 1216 -592 1267 -584
rect 1216 -604 1241 -592
rect 1248 -604 1267 -592
rect 1298 -592 1348 -584
rect 1298 -600 1314 -592
rect 1321 -594 1348 -592
rect 1357 -594 1551 -584
rect 1321 -604 1551 -594
rect 1216 -612 1267 -604
rect 1314 -612 1551 -604
rect 1232 -620 1233 -612
rect 1248 -620 1261 -612
rect 1232 -628 1248 -620
rect 1229 -635 1248 -632
rect 1229 -644 1251 -635
rect 1202 -654 1251 -644
rect 1202 -660 1232 -654
rect 1251 -659 1256 -654
rect 1174 -676 1248 -660
rect 1266 -668 1296 -612
rect 1331 -622 1539 -612
rect 1357 -652 1546 -622
rect 1372 -655 1546 -652
rect 1365 -658 1546 -655
rect 1174 -678 1187 -676
rect 1202 -678 1236 -676
rect 1174 -694 1248 -678
rect 1275 -682 1288 -668
rect 1303 -682 1319 -666
rect 1365 -671 1376 -658
rect 1158 -716 1159 -700
rect 1174 -716 1187 -694
rect 1202 -716 1232 -694
rect 1275 -698 1337 -682
rect 1365 -689 1376 -673
rect 1381 -678 1391 -658
rect 1401 -678 1415 -658
rect 1418 -671 1427 -658
rect 1443 -671 1452 -658
rect 1381 -689 1415 -678
rect 1418 -689 1427 -673
rect 1443 -689 1452 -673
rect 1459 -678 1469 -658
rect 1479 -678 1493 -658
rect 1494 -671 1505 -658
rect 1459 -689 1493 -678
rect 1494 -689 1505 -673
rect 1275 -700 1288 -698
rect 1303 -700 1337 -698
rect 1275 -716 1337 -700
rect 1381 -705 1397 -698
rect 1459 -705 1489 -694
rect 1537 -700 1551 -682
rect 1536 -716 1551 -700
rect -8 -724 33 -716
rect -8 -750 7 -724
rect 14 -750 33 -724
rect 97 -728 159 -716
rect 171 -728 246 -716
rect 304 -728 379 -716
rect 391 -728 422 -716
rect 428 -728 463 -716
rect 97 -730 259 -728
rect -8 -758 33 -750
rect 115 -754 128 -730
rect 143 -732 158 -730
rect -2 -768 -1 -758
rect 14 -768 27 -758
rect 42 -768 72 -754
rect 115 -768 158 -754
rect 182 -757 189 -750
rect 192 -754 259 -730
rect 291 -730 463 -728
rect 261 -752 289 -748
rect 291 -752 371 -730
rect 392 -732 407 -730
rect 261 -754 371 -752
rect 192 -758 371 -754
rect 165 -768 195 -758
rect 197 -768 350 -758
rect 358 -768 388 -758
rect 392 -768 422 -754
rect 450 -768 463 -730
rect 535 -724 570 -716
rect 535 -750 536 -724
rect 543 -750 570 -724
rect 478 -768 508 -754
rect 535 -758 570 -750
rect 572 -724 613 -716
rect 572 -750 587 -724
rect 594 -750 613 -724
rect 677 -728 739 -716
rect 751 -728 826 -716
rect 884 -728 959 -716
rect 971 -728 1002 -716
rect 1008 -728 1043 -716
rect 677 -730 839 -728
rect 572 -758 613 -750
rect 695 -754 708 -730
rect 723 -732 738 -730
rect 535 -768 536 -758
rect 551 -768 564 -758
rect 578 -768 579 -758
rect 594 -768 607 -758
rect 622 -768 652 -754
rect 695 -768 738 -754
rect 762 -757 769 -750
rect 772 -754 839 -730
rect 871 -730 1043 -728
rect 841 -752 869 -748
rect 871 -752 951 -730
rect 972 -732 987 -730
rect 841 -754 951 -752
rect 772 -758 951 -754
rect 745 -768 775 -758
rect 777 -768 930 -758
rect 938 -768 968 -758
rect 972 -768 1002 -754
rect 1030 -768 1043 -730
rect 1115 -724 1150 -716
rect 1115 -750 1116 -724
rect 1123 -750 1150 -724
rect 1058 -768 1088 -754
rect 1115 -758 1150 -750
rect 1152 -724 1193 -716
rect 1152 -750 1167 -724
rect 1174 -750 1193 -724
rect 1257 -728 1319 -716
rect 1331 -728 1406 -716
rect 1464 -728 1539 -716
rect 1257 -730 1419 -728
rect 1152 -758 1193 -750
rect 1275 -754 1288 -730
rect 1303 -732 1318 -730
rect 1115 -768 1116 -758
rect 1131 -768 1144 -758
rect 1158 -768 1159 -758
rect 1174 -768 1187 -758
rect 1202 -768 1232 -754
rect 1275 -768 1318 -754
rect 1342 -757 1349 -750
rect 1352 -754 1419 -730
rect 1451 -730 1551 -728
rect 1421 -752 1449 -748
rect 1451 -752 1531 -730
rect 1421 -754 1531 -752
rect 1352 -758 1531 -754
rect 1325 -768 1355 -758
rect 1357 -768 1510 -758
rect 1518 -768 1548 -758
rect -2 -774 1551 -768
rect -1 -782 1551 -774
rect 14 -812 27 -782
rect 42 -800 72 -782
rect 115 -796 129 -782
rect 165 -796 385 -782
rect 116 -798 129 -796
rect 82 -810 97 -798
rect 79 -812 101 -810
rect 106 -812 136 -798
rect 197 -800 350 -796
rect 179 -812 371 -800
rect 414 -812 444 -798
rect 450 -812 463 -782
rect 478 -800 508 -782
rect 551 -812 564 -782
rect 594 -812 607 -782
rect 622 -800 652 -782
rect 695 -796 709 -782
rect 745 -796 965 -782
rect 696 -798 709 -796
rect 662 -810 677 -798
rect 659 -812 681 -810
rect 686 -812 716 -798
rect 777 -800 930 -796
rect 759 -812 951 -800
rect 994 -812 1024 -798
rect 1030 -812 1043 -782
rect 1058 -800 1088 -782
rect 1131 -812 1144 -782
rect 1174 -812 1187 -782
rect 1202 -800 1232 -782
rect 1275 -796 1289 -782
rect 1325 -796 1545 -782
rect 1276 -798 1289 -796
rect 1242 -810 1257 -798
rect 1239 -812 1261 -810
rect 1266 -812 1296 -798
rect 1357 -800 1510 -796
rect 1339 -812 1531 -800
rect -1 -826 1551 -812
rect 14 -930 27 -826
rect 72 -848 73 -838
rect 88 -848 101 -838
rect 72 -852 101 -848
rect 106 -852 136 -826
rect 154 -840 170 -838
rect 242 -840 295 -826
rect 243 -842 307 -840
rect 350 -842 365 -826
rect 414 -829 444 -826
rect 414 -832 450 -829
rect 380 -840 396 -838
rect 154 -852 169 -848
rect 72 -854 169 -852
rect 197 -854 365 -842
rect 381 -852 396 -848
rect 414 -851 453 -832
rect 472 -838 479 -837
rect 478 -845 479 -838
rect 462 -848 463 -845
rect 478 -848 491 -845
rect 414 -852 444 -851
rect 453 -852 459 -851
rect 462 -852 491 -848
rect 381 -853 491 -852
rect 381 -854 497 -853
rect 56 -862 107 -854
rect 56 -874 81 -862
rect 88 -874 107 -862
rect 138 -862 188 -854
rect 138 -870 154 -862
rect 161 -864 188 -862
rect 197 -864 418 -854
rect 161 -874 418 -864
rect 447 -862 497 -854
rect 447 -871 463 -862
rect 56 -882 107 -874
rect 154 -882 418 -874
rect 444 -874 463 -871
rect 470 -874 497 -862
rect 444 -882 497 -874
rect 72 -890 73 -882
rect 88 -890 101 -882
rect 72 -898 88 -890
rect 69 -905 88 -902
rect 69 -914 91 -905
rect 42 -924 91 -914
rect 42 -930 72 -924
rect 91 -929 96 -924
rect 14 -946 88 -930
rect 106 -938 136 -882
rect 171 -892 379 -882
rect 414 -886 459 -882
rect 462 -883 463 -882
rect 478 -883 491 -882
rect 197 -922 386 -892
rect 212 -925 386 -922
rect 205 -928 386 -925
rect 14 -948 27 -946
rect 42 -948 76 -946
rect 14 -964 88 -948
rect 115 -952 128 -938
rect 143 -952 159 -936
rect 205 -941 216 -928
rect -2 -986 -1 -970
rect 14 -986 27 -964
rect 42 -986 72 -964
rect 115 -968 177 -952
rect 205 -959 216 -943
rect 221 -948 231 -928
rect 241 -948 255 -928
rect 258 -941 267 -928
rect 283 -941 292 -928
rect 221 -959 255 -948
rect 258 -959 267 -943
rect 283 -959 292 -943
rect 299 -948 309 -928
rect 319 -948 333 -928
rect 334 -941 345 -928
rect 299 -959 333 -948
rect 334 -959 345 -943
rect 391 -952 407 -936
rect 414 -938 444 -886
rect 478 -890 479 -883
rect 463 -898 479 -890
rect 450 -930 463 -911
rect 478 -930 508 -914
rect 450 -946 524 -930
rect 450 -948 463 -946
rect 478 -948 512 -946
rect 115 -970 128 -968
rect 143 -970 177 -968
rect 115 -986 177 -970
rect 221 -975 237 -968
rect 299 -975 329 -964
rect 377 -968 423 -952
rect 450 -964 524 -948
rect 377 -970 411 -968
rect 376 -986 423 -970
rect 450 -986 463 -964
rect 478 -986 508 -964
rect 535 -986 536 -970
rect 551 -986 564 -826
rect 594 -930 607 -826
rect 652 -848 653 -838
rect 668 -848 681 -838
rect 652 -852 681 -848
rect 686 -852 716 -826
rect 734 -840 750 -838
rect 822 -840 875 -826
rect 823 -842 887 -840
rect 930 -842 945 -826
rect 994 -829 1024 -826
rect 994 -832 1030 -829
rect 960 -840 976 -838
rect 734 -852 749 -848
rect 652 -854 749 -852
rect 777 -854 945 -842
rect 961 -852 976 -848
rect 994 -851 1033 -832
rect 1052 -838 1059 -837
rect 1058 -845 1059 -838
rect 1042 -848 1043 -845
rect 1058 -848 1071 -845
rect 994 -852 1024 -851
rect 1033 -852 1039 -851
rect 1042 -852 1071 -848
rect 961 -853 1071 -852
rect 961 -854 1077 -853
rect 636 -862 687 -854
rect 636 -874 661 -862
rect 668 -874 687 -862
rect 718 -862 768 -854
rect 718 -870 734 -862
rect 741 -864 768 -862
rect 777 -864 998 -854
rect 741 -874 998 -864
rect 1027 -862 1077 -854
rect 1027 -871 1043 -862
rect 636 -882 687 -874
rect 734 -882 998 -874
rect 1024 -874 1043 -871
rect 1050 -874 1077 -862
rect 1024 -882 1077 -874
rect 652 -890 653 -882
rect 668 -890 681 -882
rect 652 -898 668 -890
rect 649 -905 668 -902
rect 649 -914 671 -905
rect 622 -924 671 -914
rect 622 -930 652 -924
rect 671 -929 676 -924
rect 594 -946 668 -930
rect 686 -938 716 -882
rect 751 -892 959 -882
rect 994 -886 1039 -882
rect 1042 -883 1043 -882
rect 1058 -883 1071 -882
rect 777 -922 966 -892
rect 792 -925 966 -922
rect 785 -928 966 -925
rect 594 -948 607 -946
rect 622 -948 656 -946
rect 594 -964 668 -948
rect 695 -952 708 -938
rect 723 -952 739 -936
rect 785 -941 796 -928
rect 578 -986 579 -970
rect 594 -986 607 -964
rect 622 -986 652 -964
rect 695 -968 757 -952
rect 785 -959 796 -943
rect 801 -948 811 -928
rect 821 -948 835 -928
rect 838 -941 847 -928
rect 863 -941 872 -928
rect 801 -959 835 -948
rect 838 -959 847 -943
rect 863 -959 872 -943
rect 879 -948 889 -928
rect 899 -948 913 -928
rect 914 -941 925 -928
rect 879 -959 913 -948
rect 914 -959 925 -943
rect 971 -952 987 -936
rect 994 -938 1024 -886
rect 1058 -890 1059 -883
rect 1043 -898 1059 -890
rect 1030 -930 1043 -911
rect 1058 -930 1088 -914
rect 1030 -946 1104 -930
rect 1030 -948 1043 -946
rect 1058 -948 1092 -946
rect 695 -970 708 -968
rect 723 -970 757 -968
rect 695 -986 757 -970
rect 801 -975 817 -968
rect 879 -975 909 -964
rect 957 -968 1003 -952
rect 1030 -964 1104 -948
rect 957 -970 991 -968
rect 956 -986 1003 -970
rect 1030 -986 1043 -964
rect 1058 -986 1088 -964
rect 1115 -986 1116 -970
rect 1131 -986 1144 -826
rect 1174 -930 1187 -826
rect 1232 -848 1233 -838
rect 1248 -848 1261 -838
rect 1232 -852 1261 -848
rect 1266 -852 1296 -826
rect 1314 -840 1330 -838
rect 1402 -840 1455 -826
rect 1403 -842 1467 -840
rect 1510 -842 1525 -826
rect 1540 -840 1551 -838
rect 1314 -852 1329 -848
rect 1232 -854 1329 -852
rect 1357 -854 1525 -842
rect 1541 -854 1551 -848
rect 1216 -862 1267 -854
rect 1216 -874 1241 -862
rect 1248 -874 1267 -862
rect 1298 -862 1348 -854
rect 1298 -870 1314 -862
rect 1321 -864 1348 -862
rect 1357 -864 1551 -854
rect 1321 -874 1551 -864
rect 1216 -882 1267 -874
rect 1314 -882 1551 -874
rect 1232 -890 1233 -882
rect 1248 -890 1261 -882
rect 1232 -898 1248 -890
rect 1229 -905 1248 -902
rect 1229 -914 1251 -905
rect 1202 -924 1251 -914
rect 1202 -930 1232 -924
rect 1251 -929 1256 -924
rect 1174 -946 1248 -930
rect 1266 -938 1296 -882
rect 1331 -892 1539 -882
rect 1357 -922 1546 -892
rect 1372 -925 1546 -922
rect 1365 -928 1546 -925
rect 1174 -948 1187 -946
rect 1202 -948 1236 -946
rect 1174 -964 1248 -948
rect 1275 -952 1288 -938
rect 1303 -952 1319 -936
rect 1365 -941 1376 -928
rect 1158 -986 1159 -970
rect 1174 -986 1187 -964
rect 1202 -986 1232 -964
rect 1275 -968 1337 -952
rect 1365 -959 1376 -943
rect 1381 -948 1391 -928
rect 1401 -948 1415 -928
rect 1418 -941 1427 -928
rect 1443 -941 1452 -928
rect 1381 -959 1415 -948
rect 1418 -959 1427 -943
rect 1443 -959 1452 -943
rect 1459 -948 1469 -928
rect 1479 -948 1493 -928
rect 1494 -941 1505 -928
rect 3379 -930 3408 -914
rect 1459 -959 1493 -948
rect 1494 -959 1505 -943
rect 3379 -946 3424 -930
rect 3379 -948 3412 -946
rect 1275 -970 1288 -968
rect 1303 -970 1337 -968
rect 1275 -986 1337 -970
rect 1381 -975 1397 -968
rect 1459 -975 1489 -964
rect 1537 -970 1551 -952
rect 1536 -986 1551 -970
rect 3379 -964 3424 -948
rect 3379 -986 3408 -964
rect 3435 -986 3436 -970
rect 3451 -986 3464 -886
rect 3494 -930 3507 -886
rect 3552 -890 3553 -886
rect 3568 -890 3581 -886
rect 3552 -898 3568 -890
rect 3549 -905 3568 -902
rect 3549 -914 3571 -905
rect 3522 -924 3571 -914
rect 3522 -930 3552 -924
rect 3571 -929 3576 -924
rect 3494 -946 3568 -930
rect 3586 -938 3616 -886
rect 3651 -892 3859 -886
rect 3677 -922 3866 -892
rect 3692 -925 3866 -922
rect 3685 -928 3866 -925
rect 3494 -948 3507 -946
rect 3522 -948 3556 -946
rect 3494 -964 3568 -948
rect 3595 -952 3608 -938
rect 3623 -952 3639 -936
rect 3685 -941 3696 -928
rect 3478 -986 3479 -970
rect 3494 -986 3507 -964
rect 3522 -986 3552 -964
rect 3595 -968 3657 -952
rect 3685 -959 3696 -943
rect 3701 -948 3711 -928
rect 3721 -948 3735 -928
rect 3738 -941 3747 -928
rect 3763 -941 3772 -928
rect 3701 -959 3735 -948
rect 3738 -959 3747 -943
rect 3763 -959 3772 -943
rect 3779 -948 3789 -928
rect 3799 -948 3813 -928
rect 3814 -941 3825 -928
rect 3779 -959 3813 -948
rect 3814 -959 3825 -943
rect 3871 -952 3887 -936
rect 3894 -938 3924 -886
rect 3958 -890 3959 -886
rect 3943 -898 3959 -890
rect 3930 -930 3943 -911
rect 3958 -930 3988 -914
rect 3930 -946 4004 -930
rect 3930 -948 3943 -946
rect 3958 -948 3992 -946
rect 3595 -970 3608 -968
rect 3623 -970 3657 -968
rect 3595 -986 3657 -970
rect 3701 -975 3717 -968
rect 3779 -975 3809 -964
rect 3857 -968 3903 -952
rect 3930 -964 4004 -948
rect 3857 -970 3891 -968
rect 3856 -986 3903 -970
rect 3930 -986 3943 -964
rect 3958 -986 3988 -964
rect 4015 -986 4016 -970
rect 4031 -986 4044 -886
rect 4074 -930 4087 -886
rect 4132 -890 4133 -886
rect 4148 -890 4161 -886
rect 4132 -898 4148 -890
rect 4129 -905 4148 -902
rect 4129 -914 4151 -905
rect 4102 -924 4151 -914
rect 4102 -930 4132 -924
rect 4151 -929 4156 -924
rect 4074 -946 4148 -930
rect 4166 -938 4196 -886
rect 4231 -892 4439 -886
rect 4257 -922 4446 -892
rect 4272 -925 4446 -922
rect 4265 -928 4446 -925
rect 4074 -948 4087 -946
rect 4102 -948 4136 -946
rect 4074 -964 4148 -948
rect 4175 -952 4188 -938
rect 4203 -952 4219 -936
rect 4265 -941 4276 -928
rect 4058 -986 4059 -970
rect 4074 -986 4087 -964
rect 4102 -986 4132 -964
rect 4175 -968 4237 -952
rect 4265 -959 4276 -943
rect 4281 -948 4291 -928
rect 4301 -948 4315 -928
rect 4318 -941 4327 -928
rect 4343 -941 4352 -928
rect 4281 -959 4315 -948
rect 4318 -959 4327 -943
rect 4343 -959 4352 -943
rect 4359 -948 4369 -928
rect 4379 -948 4393 -928
rect 4394 -941 4405 -928
rect 4359 -959 4393 -948
rect 4394 -959 4405 -943
rect 4451 -952 4467 -936
rect 4474 -938 4504 -886
rect 4538 -890 4539 -886
rect 4523 -898 4539 -890
rect 4510 -930 4523 -911
rect 4538 -930 4568 -914
rect 4510 -946 4584 -930
rect 4510 -948 4523 -946
rect 4538 -948 4572 -946
rect 4175 -970 4188 -968
rect 4203 -970 4237 -968
rect 4175 -986 4237 -970
rect 4281 -975 4297 -968
rect 4359 -975 4389 -964
rect 4437 -968 4483 -952
rect 4510 -964 4584 -948
rect 4437 -970 4471 -968
rect 4436 -986 4483 -970
rect 4510 -986 4523 -964
rect 4538 -986 4568 -964
rect 4595 -986 4596 -970
rect 4611 -986 4624 -886
rect 4654 -930 4667 -886
rect 4712 -890 4713 -886
rect 4728 -890 4741 -886
rect 4712 -898 4728 -890
rect 4709 -905 4728 -902
rect 4709 -914 4731 -905
rect 4682 -924 4731 -914
rect 4682 -930 4712 -924
rect 4731 -929 4736 -924
rect 4654 -946 4728 -930
rect 4746 -938 4776 -886
rect 4811 -892 5019 -886
rect 4837 -922 5026 -892
rect 4852 -925 5026 -922
rect 4845 -928 5026 -925
rect 4654 -948 4667 -946
rect 4682 -948 4716 -946
rect 4654 -964 4728 -948
rect 4755 -952 4768 -938
rect 4783 -952 4799 -936
rect 4845 -941 4856 -928
rect 4638 -986 4639 -970
rect 4654 -986 4667 -964
rect 4682 -986 4712 -964
rect 4755 -968 4817 -952
rect 4845 -959 4856 -943
rect 4861 -948 4871 -928
rect 4881 -948 4895 -928
rect 4898 -941 4907 -928
rect 4923 -941 4932 -928
rect 4861 -959 4895 -948
rect 4898 -959 4907 -943
rect 4923 -959 4932 -943
rect 4939 -948 4949 -928
rect 4959 -948 4973 -928
rect 4974 -941 4985 -928
rect 4939 -959 4973 -948
rect 4974 -959 4985 -943
rect 5031 -952 5047 -936
rect 5054 -938 5084 -886
rect 5118 -890 5119 -886
rect 5103 -898 5119 -890
rect 5090 -930 5103 -911
rect 5118 -930 5148 -914
rect 5090 -946 5164 -930
rect 5090 -948 5103 -946
rect 5118 -948 5152 -946
rect 4755 -970 4768 -968
rect 4783 -970 4817 -968
rect 4755 -986 4817 -970
rect 4861 -975 4877 -968
rect 4939 -975 4969 -964
rect 5017 -968 5063 -952
rect 5090 -964 5164 -948
rect 5017 -970 5051 -968
rect 5016 -986 5063 -970
rect 5090 -986 5103 -964
rect 5118 -986 5148 -964
rect 5175 -986 5176 -970
rect 5191 -986 5204 -886
rect 5234 -930 5247 -886
rect 5292 -890 5293 -886
rect 5308 -890 5321 -886
rect 5292 -898 5308 -890
rect 5289 -905 5308 -902
rect 5289 -914 5311 -905
rect 5262 -924 5311 -914
rect 5262 -930 5292 -924
rect 5311 -929 5316 -924
rect 5234 -946 5308 -930
rect 5326 -938 5356 -886
rect 5391 -892 5599 -886
rect 5417 -922 5606 -892
rect 5432 -925 5606 -922
rect 5425 -928 5606 -925
rect 5234 -948 5247 -946
rect 5262 -948 5296 -946
rect 5234 -964 5308 -948
rect 5335 -952 5348 -938
rect 5363 -952 5379 -936
rect 5425 -941 5436 -928
rect 5218 -986 5219 -970
rect 5234 -986 5247 -964
rect 5262 -986 5292 -964
rect 5335 -968 5397 -952
rect 5425 -959 5436 -943
rect 5441 -948 5451 -928
rect 5461 -948 5475 -928
rect 5478 -941 5487 -928
rect 5503 -941 5512 -928
rect 5441 -959 5475 -948
rect 5478 -959 5487 -943
rect 5503 -959 5512 -943
rect 5519 -948 5529 -928
rect 5539 -948 5553 -928
rect 5554 -941 5565 -928
rect 5519 -959 5553 -948
rect 5554 -959 5565 -943
rect 5611 -952 5627 -936
rect 5634 -938 5664 -886
rect 5698 -890 5699 -886
rect 5683 -898 5699 -890
rect 5670 -930 5683 -911
rect 5698 -930 5728 -914
rect 5670 -946 5744 -930
rect 5670 -948 5683 -946
rect 5698 -948 5732 -946
rect 5335 -970 5348 -968
rect 5363 -970 5397 -968
rect 5335 -986 5397 -970
rect 5441 -975 5457 -968
rect 5519 -975 5549 -964
rect 5597 -968 5643 -952
rect 5670 -964 5744 -948
rect 5597 -970 5631 -968
rect 5596 -986 5643 -970
rect 5670 -986 5683 -964
rect 5698 -986 5728 -964
rect 5755 -986 5756 -970
rect 5771 -986 5784 -886
rect 5814 -930 5827 -886
rect 5872 -890 5873 -886
rect 5888 -890 5901 -886
rect 5872 -898 5888 -890
rect 5869 -905 5888 -902
rect 5869 -914 5891 -905
rect 5842 -924 5891 -914
rect 5842 -930 5872 -924
rect 5891 -929 5896 -924
rect 5814 -946 5888 -930
rect 5906 -938 5936 -886
rect 5971 -892 6179 -886
rect 5997 -922 6186 -892
rect 6012 -925 6186 -922
rect 6005 -928 6186 -925
rect 5814 -948 5827 -946
rect 5842 -948 5876 -946
rect 5814 -964 5888 -948
rect 5915 -952 5928 -938
rect 5943 -952 5959 -936
rect 6005 -941 6016 -928
rect 5798 -986 5799 -970
rect 5814 -986 5827 -964
rect 5842 -986 5872 -964
rect 5915 -968 5977 -952
rect 6005 -959 6016 -943
rect 6021 -948 6031 -928
rect 6041 -948 6055 -928
rect 6058 -941 6067 -928
rect 6083 -941 6092 -928
rect 6021 -959 6055 -948
rect 6058 -959 6067 -943
rect 6083 -959 6092 -943
rect 6099 -948 6109 -928
rect 6119 -948 6133 -928
rect 6134 -941 6145 -928
rect 6099 -959 6133 -948
rect 6134 -959 6145 -943
rect 6191 -952 6207 -936
rect 6214 -938 6244 -886
rect 6278 -890 6279 -886
rect 6263 -898 6279 -890
rect 6250 -930 6263 -911
rect 6278 -930 6308 -914
rect 6250 -946 6324 -930
rect 6250 -948 6263 -946
rect 6278 -948 6312 -946
rect 5915 -970 5928 -968
rect 5943 -970 5977 -968
rect 5915 -986 5977 -970
rect 6021 -975 6037 -968
rect 6099 -975 6129 -964
rect 6177 -968 6223 -952
rect 6250 -964 6324 -948
rect 6177 -970 6211 -968
rect 6176 -986 6223 -970
rect 6250 -986 6263 -964
rect 6278 -986 6308 -964
rect 6335 -986 6336 -970
rect 6351 -986 6364 -886
rect 6394 -930 6407 -886
rect 6452 -890 6453 -886
rect 6468 -890 6481 -886
rect 6452 -898 6468 -890
rect 6449 -905 6468 -902
rect 6449 -914 6471 -905
rect 6422 -924 6471 -914
rect 6422 -930 6452 -924
rect 6471 -929 6476 -924
rect 6394 -946 6468 -930
rect 6486 -938 6516 -886
rect 6551 -892 6759 -886
rect 6577 -922 6766 -892
rect 6592 -925 6766 -922
rect 6585 -928 6766 -925
rect 6394 -948 6407 -946
rect 6422 -948 6456 -946
rect 6394 -964 6468 -948
rect 6495 -952 6508 -938
rect 6523 -952 6539 -936
rect 6585 -941 6596 -928
rect 6378 -986 6379 -970
rect 6394 -986 6407 -964
rect 6422 -986 6452 -964
rect 6495 -968 6557 -952
rect 6585 -959 6596 -943
rect 6601 -948 6611 -928
rect 6621 -948 6635 -928
rect 6638 -941 6647 -928
rect 6663 -941 6672 -928
rect 6601 -959 6635 -948
rect 6638 -959 6647 -943
rect 6663 -959 6672 -943
rect 6679 -948 6689 -928
rect 6699 -948 6713 -928
rect 6714 -941 6725 -928
rect 6679 -959 6713 -948
rect 6714 -959 6725 -943
rect 6771 -952 6787 -936
rect 6794 -938 6824 -886
rect 6858 -890 6859 -886
rect 6843 -898 6859 -890
rect 6830 -930 6843 -911
rect 6858 -930 6888 -914
rect 6830 -946 6904 -930
rect 6830 -948 6843 -946
rect 6858 -948 6892 -946
rect 6495 -970 6508 -968
rect 6523 -970 6557 -968
rect 6495 -986 6557 -970
rect 6601 -975 6617 -968
rect 6679 -975 6709 -964
rect 6757 -968 6803 -952
rect 6830 -964 6904 -948
rect 6757 -970 6791 -968
rect 6756 -986 6803 -970
rect 6830 -986 6843 -964
rect 6858 -986 6888 -964
rect 6915 -986 6916 -970
rect 6931 -986 6944 -886
rect -8 -994 33 -986
rect -8 -1020 7 -994
rect 14 -1020 33 -994
rect 97 -998 159 -986
rect 171 -998 246 -986
rect 304 -998 379 -986
rect 391 -998 422 -986
rect 428 -998 463 -986
rect 97 -1000 259 -998
rect -8 -1028 33 -1020
rect 115 -1024 128 -1000
rect 143 -1002 158 -1000
rect -2 -1038 -1 -1028
rect 14 -1038 27 -1028
rect 42 -1038 72 -1024
rect 115 -1038 158 -1024
rect 182 -1027 189 -1020
rect 192 -1024 259 -1000
rect 291 -1000 463 -998
rect 261 -1022 289 -1018
rect 291 -1022 371 -1000
rect 392 -1002 407 -1000
rect 261 -1024 371 -1022
rect 192 -1028 371 -1024
rect 165 -1038 195 -1028
rect 197 -1038 350 -1028
rect 358 -1038 388 -1028
rect 392 -1038 422 -1024
rect 450 -1038 463 -1000
rect 535 -994 570 -986
rect 535 -1020 536 -994
rect 543 -1020 570 -994
rect 478 -1038 508 -1024
rect 535 -1028 570 -1020
rect 572 -994 613 -986
rect 572 -1020 587 -994
rect 594 -1020 613 -994
rect 677 -998 739 -986
rect 751 -998 826 -986
rect 884 -998 959 -986
rect 971 -998 1002 -986
rect 1008 -998 1043 -986
rect 677 -1000 839 -998
rect 572 -1028 613 -1020
rect 695 -1024 708 -1000
rect 723 -1002 738 -1000
rect 535 -1038 536 -1028
rect 551 -1038 564 -1028
rect 578 -1038 579 -1028
rect 594 -1038 607 -1028
rect 622 -1038 652 -1024
rect 695 -1038 738 -1024
rect 762 -1027 769 -1020
rect 772 -1024 839 -1000
rect 871 -1000 1043 -998
rect 841 -1022 869 -1018
rect 871 -1022 951 -1000
rect 972 -1002 987 -1000
rect 841 -1024 951 -1022
rect 772 -1028 951 -1024
rect 745 -1038 775 -1028
rect 777 -1038 930 -1028
rect 938 -1038 968 -1028
rect 972 -1038 1002 -1024
rect 1030 -1038 1043 -1000
rect 1115 -994 1150 -986
rect 1115 -1020 1116 -994
rect 1123 -1020 1150 -994
rect 1058 -1038 1088 -1024
rect 1115 -1028 1150 -1020
rect 1152 -994 1193 -986
rect 1152 -1020 1167 -994
rect 1174 -1020 1193 -994
rect 1257 -998 1319 -986
rect 1331 -998 1406 -986
rect 1464 -998 1539 -986
rect 3435 -994 3470 -986
rect 1257 -1000 1419 -998
rect 1152 -1028 1193 -1020
rect 1275 -1024 1288 -1000
rect 1303 -1002 1318 -1000
rect 1115 -1038 1116 -1028
rect 1131 -1038 1144 -1028
rect 1158 -1038 1159 -1028
rect 1174 -1038 1187 -1028
rect 1202 -1038 1232 -1024
rect 1275 -1038 1318 -1024
rect 1342 -1027 1349 -1020
rect 1352 -1024 1419 -1000
rect 1451 -1000 1551 -998
rect 1421 -1022 1449 -1018
rect 1451 -1022 1531 -1000
rect 1421 -1024 1531 -1022
rect 3435 -1020 3436 -994
rect 3443 -1020 3470 -994
rect 1352 -1028 1531 -1024
rect 1325 -1038 1355 -1028
rect 1357 -1038 1510 -1028
rect 1518 -1038 1548 -1028
rect 3379 -1038 3408 -1024
rect 3435 -1028 3470 -1020
rect 3472 -994 3513 -986
rect 3472 -1020 3487 -994
rect 3494 -1020 3513 -994
rect 3577 -998 3639 -986
rect 3651 -998 3726 -986
rect 3784 -998 3859 -986
rect 3871 -998 3902 -986
rect 3908 -998 3943 -986
rect 3577 -1000 3739 -998
rect 3472 -1028 3513 -1020
rect 3595 -1024 3608 -1000
rect 3623 -1002 3638 -1000
rect 3435 -1038 3436 -1028
rect 3451 -1038 3464 -1028
rect 3478 -1038 3479 -1028
rect 3494 -1038 3507 -1028
rect 3522 -1038 3552 -1024
rect 3595 -1038 3638 -1024
rect 3662 -1027 3669 -1020
rect 3672 -1024 3739 -1000
rect 3771 -1000 3943 -998
rect 3741 -1022 3769 -1018
rect 3771 -1022 3851 -1000
rect 3872 -1002 3887 -1000
rect 3741 -1024 3851 -1022
rect 3672 -1028 3851 -1024
rect 3645 -1038 3675 -1028
rect 3677 -1038 3830 -1028
rect 3838 -1038 3868 -1028
rect 3872 -1038 3902 -1024
rect 3930 -1038 3943 -1000
rect 4015 -994 4050 -986
rect 4015 -1020 4016 -994
rect 4023 -1020 4050 -994
rect 3958 -1038 3988 -1024
rect 4015 -1028 4050 -1020
rect 4052 -994 4093 -986
rect 4052 -1020 4067 -994
rect 4074 -1020 4093 -994
rect 4157 -998 4219 -986
rect 4231 -998 4306 -986
rect 4364 -998 4439 -986
rect 4451 -998 4482 -986
rect 4488 -998 4523 -986
rect 4157 -1000 4319 -998
rect 4052 -1028 4093 -1020
rect 4175 -1024 4188 -1000
rect 4203 -1002 4218 -1000
rect 4015 -1038 4016 -1028
rect 4031 -1038 4044 -1028
rect 4058 -1038 4059 -1028
rect 4074 -1038 4087 -1028
rect 4102 -1038 4132 -1024
rect 4175 -1038 4218 -1024
rect 4242 -1027 4249 -1020
rect 4252 -1024 4319 -1000
rect 4351 -1000 4523 -998
rect 4321 -1022 4349 -1018
rect 4351 -1022 4431 -1000
rect 4452 -1002 4467 -1000
rect 4321 -1024 4431 -1022
rect 4252 -1028 4431 -1024
rect 4225 -1038 4255 -1028
rect 4257 -1038 4410 -1028
rect 4418 -1038 4448 -1028
rect 4452 -1038 4482 -1024
rect 4510 -1038 4523 -1000
rect 4595 -994 4630 -986
rect 4595 -1020 4596 -994
rect 4603 -1020 4630 -994
rect 4538 -1038 4568 -1024
rect 4595 -1028 4630 -1020
rect 4632 -994 4673 -986
rect 4632 -1020 4647 -994
rect 4654 -1020 4673 -994
rect 4737 -998 4799 -986
rect 4811 -998 4886 -986
rect 4944 -998 5019 -986
rect 5031 -998 5062 -986
rect 5068 -998 5103 -986
rect 4737 -1000 4899 -998
rect 4755 -1018 4768 -1000
rect 4783 -1002 4798 -1000
rect 4632 -1028 4673 -1020
rect 4756 -1024 4768 -1018
rect 4832 -1018 4899 -1000
rect 4931 -1000 5103 -998
rect 4931 -1018 5011 -1000
rect 5032 -1002 5047 -1000
rect 4595 -1038 4596 -1028
rect 4611 -1038 4624 -1028
rect 4638 -1038 4639 -1028
rect 4654 -1038 4667 -1028
rect 4682 -1038 4712 -1024
rect 4756 -1038 4798 -1024
rect 4822 -1027 4829 -1020
rect 4832 -1028 5011 -1018
rect 4805 -1038 4835 -1028
rect 4837 -1038 4990 -1028
rect 4998 -1038 5028 -1028
rect 5032 -1038 5062 -1024
rect 5090 -1038 5103 -1000
rect 5175 -994 5210 -986
rect 5175 -1020 5176 -994
rect 5183 -1020 5210 -994
rect 5118 -1038 5148 -1024
rect 5175 -1028 5210 -1020
rect 5212 -994 5253 -986
rect 5212 -1020 5227 -994
rect 5234 -1020 5253 -994
rect 5317 -998 5379 -986
rect 5391 -998 5466 -986
rect 5524 -998 5599 -986
rect 5611 -998 5642 -986
rect 5648 -998 5683 -986
rect 5317 -1000 5479 -998
rect 5335 -1018 5348 -1000
rect 5363 -1002 5378 -1000
rect 5212 -1028 5253 -1020
rect 5336 -1024 5348 -1018
rect 5412 -1018 5479 -1000
rect 5511 -1000 5683 -998
rect 5511 -1018 5591 -1000
rect 5612 -1002 5627 -1000
rect 5175 -1038 5176 -1028
rect 5191 -1038 5204 -1028
rect 5218 -1038 5219 -1028
rect 5234 -1038 5247 -1028
rect 5262 -1038 5292 -1024
rect 5336 -1038 5378 -1024
rect 5402 -1027 5409 -1020
rect 5412 -1028 5591 -1018
rect 5385 -1038 5415 -1028
rect 5417 -1038 5570 -1028
rect 5578 -1038 5608 -1028
rect 5612 -1038 5642 -1024
rect 5670 -1038 5683 -1000
rect 5755 -994 5790 -986
rect 5755 -1020 5756 -994
rect 5763 -1020 5790 -994
rect 5698 -1038 5728 -1024
rect 5755 -1028 5790 -1020
rect 5792 -994 5833 -986
rect 5792 -1020 5807 -994
rect 5814 -1020 5833 -994
rect 5897 -998 5959 -986
rect 5971 -998 6046 -986
rect 6104 -998 6179 -986
rect 6191 -998 6222 -986
rect 6228 -998 6263 -986
rect 5897 -1000 6059 -998
rect 5915 -1018 5928 -1000
rect 5943 -1002 5958 -1000
rect 5792 -1028 5833 -1020
rect 5916 -1024 5928 -1018
rect 5992 -1018 6059 -1000
rect 6091 -1000 6263 -998
rect 6091 -1018 6171 -1000
rect 6192 -1002 6207 -1000
rect 5755 -1038 5756 -1028
rect 5771 -1038 5784 -1028
rect 5798 -1038 5799 -1028
rect 5814 -1038 5827 -1028
rect 5842 -1038 5872 -1024
rect 5916 -1038 5958 -1024
rect 5982 -1027 5989 -1020
rect 5992 -1028 6171 -1018
rect 5965 -1038 5995 -1028
rect 5997 -1038 6150 -1028
rect 6158 -1038 6188 -1028
rect 6192 -1038 6222 -1024
rect 6250 -1038 6263 -1000
rect 6335 -994 6370 -986
rect 6335 -1020 6336 -994
rect 6343 -1020 6370 -994
rect 6278 -1038 6308 -1024
rect 6335 -1028 6370 -1020
rect 6372 -994 6413 -986
rect 6372 -1020 6387 -994
rect 6394 -1020 6413 -994
rect 6477 -998 6539 -986
rect 6551 -998 6626 -986
rect 6684 -998 6759 -986
rect 6771 -998 6802 -986
rect 6808 -998 6843 -986
rect 6477 -1000 6639 -998
rect 6495 -1018 6508 -1000
rect 6523 -1002 6538 -1000
rect 6372 -1028 6413 -1020
rect 6496 -1024 6508 -1018
rect 6572 -1018 6639 -1000
rect 6671 -1000 6843 -998
rect 6671 -1018 6751 -1000
rect 6772 -1002 6787 -1000
rect 6335 -1038 6336 -1028
rect 6351 -1038 6364 -1028
rect 6378 -1038 6379 -1028
rect 6394 -1038 6407 -1028
rect 6422 -1038 6452 -1024
rect 6496 -1038 6538 -1024
rect 6562 -1027 6569 -1020
rect 6572 -1028 6751 -1018
rect 6545 -1038 6575 -1028
rect 6577 -1038 6730 -1028
rect 6738 -1038 6768 -1028
rect 6772 -1038 6802 -1024
rect 6830 -1038 6843 -1000
rect 6915 -994 6950 -986
rect 6915 -1020 6916 -994
rect 6923 -1020 6950 -994
rect 6858 -1038 6888 -1024
rect 6915 -1028 6950 -1020
rect 6915 -1038 6916 -1028
rect 6931 -1038 6944 -1028
rect -2 -1044 1551 -1038
rect -1 -1052 1551 -1044
rect 3379 -1052 6944 -1038
rect 14 -1082 27 -1052
rect 42 -1070 72 -1052
rect 115 -1066 129 -1052
rect 165 -1066 385 -1052
rect 116 -1068 129 -1066
rect 82 -1080 97 -1068
rect 79 -1082 101 -1080
rect 106 -1082 136 -1068
rect 197 -1070 350 -1066
rect 179 -1082 371 -1070
rect 414 -1082 444 -1068
rect 450 -1082 463 -1052
rect 478 -1070 508 -1052
rect 551 -1082 564 -1052
rect 594 -1082 607 -1052
rect 622 -1070 652 -1052
rect 695 -1066 709 -1052
rect 745 -1066 965 -1052
rect 696 -1068 709 -1066
rect 662 -1080 677 -1068
rect 659 -1082 681 -1080
rect 686 -1082 716 -1068
rect 777 -1070 930 -1066
rect 759 -1082 951 -1070
rect 994 -1082 1024 -1068
rect 1030 -1082 1043 -1052
rect 1058 -1070 1088 -1052
rect 1131 -1082 1144 -1052
rect 1174 -1082 1187 -1052
rect 1202 -1070 1232 -1052
rect 1275 -1066 1289 -1052
rect 1325 -1066 1545 -1052
rect 1276 -1068 1289 -1066
rect 1242 -1080 1257 -1068
rect 1239 -1082 1261 -1080
rect 1266 -1082 1296 -1068
rect 1357 -1070 1510 -1066
rect 3379 -1070 3408 -1052
rect 1339 -1082 1531 -1070
rect 3451 -1082 3464 -1052
rect 3494 -1082 3507 -1052
rect 3522 -1070 3552 -1052
rect 3595 -1066 3609 -1052
rect 3645 -1066 3865 -1052
rect 3596 -1068 3609 -1066
rect 3562 -1080 3577 -1068
rect 3559 -1082 3581 -1080
rect 3586 -1082 3616 -1068
rect 3677 -1070 3830 -1066
rect 3659 -1082 3851 -1070
rect 3894 -1082 3924 -1068
rect 3930 -1082 3943 -1052
rect 3958 -1070 3988 -1052
rect 4031 -1082 4044 -1052
rect 4074 -1082 4087 -1052
rect 4102 -1070 4132 -1052
rect 4175 -1066 4189 -1052
rect 4225 -1066 4445 -1052
rect 4176 -1068 4189 -1066
rect 4142 -1080 4157 -1068
rect 4139 -1082 4161 -1080
rect 4166 -1082 4196 -1068
rect 4257 -1070 4410 -1066
rect 4239 -1082 4431 -1070
rect 4474 -1082 4504 -1068
rect 4510 -1082 4523 -1052
rect 4538 -1070 4568 -1052
rect 4611 -1082 4624 -1052
rect 4654 -1082 4667 -1052
rect 4682 -1070 4712 -1052
rect 4756 -1068 4769 -1052
rect 4805 -1066 5025 -1052
rect 4722 -1080 4737 -1068
rect 4719 -1082 4741 -1080
rect 4746 -1082 4776 -1068
rect 4837 -1070 4990 -1066
rect 4819 -1082 5011 -1070
rect 5054 -1082 5084 -1068
rect 5090 -1082 5103 -1052
rect 5118 -1070 5148 -1052
rect 5191 -1082 5204 -1052
rect 5234 -1082 5247 -1052
rect 5262 -1070 5292 -1052
rect 5336 -1068 5349 -1052
rect 5385 -1066 5605 -1052
rect 5302 -1080 5317 -1068
rect 5299 -1082 5321 -1080
rect 5326 -1082 5356 -1068
rect 5417 -1070 5570 -1066
rect 5399 -1082 5591 -1070
rect 5634 -1082 5664 -1068
rect 5670 -1082 5683 -1052
rect 5698 -1070 5728 -1052
rect 5771 -1082 5784 -1052
rect 5814 -1082 5827 -1052
rect 5842 -1070 5872 -1052
rect 5916 -1068 5929 -1052
rect 5965 -1066 6185 -1052
rect 5882 -1080 5897 -1068
rect 5879 -1082 5901 -1080
rect 5906 -1082 5936 -1068
rect 5997 -1070 6150 -1066
rect 5979 -1082 6171 -1070
rect 6214 -1082 6244 -1068
rect 6250 -1082 6263 -1052
rect 6278 -1070 6308 -1052
rect 6351 -1082 6364 -1052
rect 6394 -1082 6407 -1052
rect 6422 -1070 6452 -1052
rect 6496 -1068 6509 -1052
rect 6545 -1066 6765 -1052
rect 6462 -1080 6477 -1068
rect 6459 -1082 6481 -1080
rect 6486 -1082 6516 -1068
rect 6577 -1070 6730 -1066
rect 6559 -1082 6751 -1070
rect 6794 -1082 6824 -1068
rect 6830 -1082 6843 -1052
rect 6858 -1070 6888 -1052
rect 6931 -1082 6944 -1052
rect -1 -1096 1551 -1082
rect 3379 -1096 6944 -1082
rect 14 -1200 27 -1096
rect 72 -1118 73 -1108
rect 88 -1118 101 -1108
rect 72 -1122 101 -1118
rect 106 -1122 136 -1096
rect 154 -1110 170 -1108
rect 242 -1110 295 -1096
rect 243 -1112 307 -1110
rect 350 -1112 365 -1096
rect 414 -1099 444 -1096
rect 414 -1102 450 -1099
rect 380 -1110 396 -1108
rect 154 -1122 169 -1118
rect 72 -1124 169 -1122
rect 197 -1124 365 -1112
rect 381 -1122 396 -1118
rect 414 -1121 453 -1102
rect 472 -1108 479 -1107
rect 478 -1115 479 -1108
rect 462 -1118 463 -1115
rect 478 -1118 491 -1115
rect 414 -1122 444 -1121
rect 453 -1122 459 -1121
rect 462 -1122 491 -1118
rect 381 -1123 491 -1122
rect 381 -1124 497 -1123
rect 56 -1132 107 -1124
rect 56 -1144 81 -1132
rect 88 -1144 107 -1132
rect 138 -1132 188 -1124
rect 138 -1140 154 -1132
rect 161 -1134 188 -1132
rect 197 -1134 418 -1124
rect 161 -1144 418 -1134
rect 447 -1132 497 -1124
rect 447 -1141 463 -1132
rect 56 -1152 107 -1144
rect 154 -1152 418 -1144
rect 444 -1144 463 -1141
rect 470 -1144 497 -1132
rect 444 -1152 497 -1144
rect 72 -1160 73 -1152
rect 88 -1160 101 -1152
rect 72 -1168 88 -1160
rect 69 -1175 88 -1172
rect 69 -1184 91 -1175
rect 42 -1194 91 -1184
rect 42 -1200 72 -1194
rect 91 -1199 96 -1194
rect 14 -1216 88 -1200
rect 106 -1208 136 -1152
rect 171 -1162 379 -1152
rect 414 -1156 459 -1152
rect 462 -1153 463 -1152
rect 478 -1153 491 -1152
rect 197 -1192 386 -1162
rect 212 -1195 386 -1192
rect 205 -1198 386 -1195
rect 14 -1218 27 -1216
rect 42 -1218 76 -1216
rect 14 -1234 88 -1218
rect 115 -1222 128 -1208
rect 143 -1222 159 -1206
rect 205 -1211 216 -1198
rect -2 -1256 -1 -1240
rect 14 -1256 27 -1234
rect 42 -1256 72 -1234
rect 115 -1238 177 -1222
rect 205 -1229 216 -1213
rect 221 -1218 231 -1198
rect 241 -1218 255 -1198
rect 258 -1211 267 -1198
rect 283 -1211 292 -1198
rect 221 -1229 255 -1218
rect 258 -1229 267 -1213
rect 283 -1229 292 -1213
rect 299 -1218 309 -1198
rect 319 -1218 333 -1198
rect 334 -1211 345 -1198
rect 299 -1229 333 -1218
rect 334 -1229 345 -1213
rect 391 -1222 407 -1206
rect 414 -1208 444 -1156
rect 478 -1160 479 -1153
rect 463 -1168 479 -1160
rect 450 -1200 463 -1181
rect 478 -1200 508 -1184
rect 450 -1216 524 -1200
rect 450 -1218 463 -1216
rect 478 -1218 512 -1216
rect 115 -1240 128 -1238
rect 143 -1240 177 -1238
rect 115 -1256 177 -1240
rect 221 -1245 237 -1238
rect 299 -1245 329 -1234
rect 377 -1238 423 -1222
rect 450 -1234 524 -1218
rect 377 -1240 411 -1238
rect 376 -1256 423 -1240
rect 450 -1256 463 -1234
rect 478 -1256 508 -1234
rect 535 -1256 536 -1240
rect 551 -1256 564 -1096
rect 594 -1200 607 -1096
rect 652 -1118 653 -1108
rect 668 -1118 681 -1108
rect 652 -1122 681 -1118
rect 686 -1122 716 -1096
rect 734 -1110 750 -1108
rect 822 -1110 875 -1096
rect 823 -1112 887 -1110
rect 930 -1112 945 -1096
rect 994 -1099 1024 -1096
rect 994 -1102 1030 -1099
rect 960 -1110 976 -1108
rect 734 -1122 749 -1118
rect 652 -1124 749 -1122
rect 777 -1124 945 -1112
rect 961 -1122 976 -1118
rect 994 -1121 1033 -1102
rect 1052 -1108 1059 -1107
rect 1058 -1115 1059 -1108
rect 1042 -1118 1043 -1115
rect 1058 -1118 1071 -1115
rect 994 -1122 1024 -1121
rect 1033 -1122 1039 -1121
rect 1042 -1122 1071 -1118
rect 961 -1123 1071 -1122
rect 961 -1124 1077 -1123
rect 636 -1132 687 -1124
rect 636 -1144 661 -1132
rect 668 -1144 687 -1132
rect 718 -1132 768 -1124
rect 718 -1140 734 -1132
rect 741 -1134 768 -1132
rect 777 -1134 998 -1124
rect 741 -1144 998 -1134
rect 1027 -1132 1077 -1124
rect 1027 -1141 1043 -1132
rect 636 -1152 687 -1144
rect 734 -1152 998 -1144
rect 1024 -1144 1043 -1141
rect 1050 -1144 1077 -1132
rect 1024 -1152 1077 -1144
rect 652 -1160 653 -1152
rect 668 -1160 681 -1152
rect 652 -1168 668 -1160
rect 649 -1175 668 -1172
rect 649 -1184 671 -1175
rect 622 -1194 671 -1184
rect 622 -1200 652 -1194
rect 671 -1199 676 -1194
rect 594 -1216 668 -1200
rect 686 -1208 716 -1152
rect 751 -1162 959 -1152
rect 994 -1156 1039 -1152
rect 1042 -1153 1043 -1152
rect 1058 -1153 1071 -1152
rect 777 -1192 966 -1162
rect 792 -1195 966 -1192
rect 785 -1198 966 -1195
rect 594 -1218 607 -1216
rect 622 -1218 656 -1216
rect 594 -1234 668 -1218
rect 695 -1222 708 -1208
rect 723 -1222 739 -1206
rect 785 -1211 796 -1198
rect 578 -1256 579 -1240
rect 594 -1256 607 -1234
rect 622 -1256 652 -1234
rect 695 -1238 757 -1222
rect 785 -1229 796 -1213
rect 801 -1218 811 -1198
rect 821 -1218 835 -1198
rect 838 -1211 847 -1198
rect 863 -1211 872 -1198
rect 801 -1229 835 -1218
rect 838 -1229 847 -1213
rect 863 -1229 872 -1213
rect 879 -1218 889 -1198
rect 899 -1218 913 -1198
rect 914 -1211 925 -1198
rect 879 -1229 913 -1218
rect 914 -1229 925 -1213
rect 971 -1222 987 -1206
rect 994 -1208 1024 -1156
rect 1058 -1160 1059 -1153
rect 1043 -1168 1059 -1160
rect 1030 -1200 1043 -1181
rect 1058 -1200 1088 -1184
rect 1030 -1216 1104 -1200
rect 1030 -1218 1043 -1216
rect 1058 -1218 1092 -1216
rect 695 -1240 708 -1238
rect 723 -1240 757 -1238
rect 695 -1256 757 -1240
rect 801 -1245 817 -1238
rect 879 -1245 909 -1234
rect 957 -1238 1003 -1222
rect 1030 -1234 1104 -1218
rect 957 -1240 991 -1238
rect 956 -1256 1003 -1240
rect 1030 -1256 1043 -1234
rect 1058 -1256 1088 -1234
rect 1115 -1256 1116 -1240
rect 1131 -1256 1144 -1096
rect 1174 -1200 1187 -1096
rect 1232 -1118 1233 -1108
rect 1248 -1118 1261 -1108
rect 1232 -1122 1261 -1118
rect 1266 -1122 1296 -1096
rect 1314 -1110 1330 -1108
rect 1402 -1110 1455 -1096
rect 1403 -1112 1467 -1110
rect 1510 -1112 1525 -1096
rect 1540 -1110 1551 -1108
rect 1314 -1122 1329 -1118
rect 1232 -1124 1329 -1122
rect 1357 -1124 1525 -1112
rect 1541 -1124 1551 -1118
rect 1216 -1132 1267 -1124
rect 1216 -1144 1241 -1132
rect 1248 -1144 1267 -1132
rect 1298 -1132 1348 -1124
rect 1298 -1140 1314 -1132
rect 1321 -1134 1348 -1132
rect 1357 -1134 1551 -1124
rect 1321 -1144 1551 -1134
rect 1216 -1152 1267 -1144
rect 1314 -1152 1551 -1144
rect 3379 -1123 3391 -1115
rect 3379 -1152 3397 -1123
rect 1232 -1160 1233 -1152
rect 1248 -1160 1261 -1152
rect 1232 -1168 1248 -1160
rect 1229 -1175 1248 -1172
rect 1229 -1184 1251 -1175
rect 1202 -1194 1251 -1184
rect 1202 -1200 1232 -1194
rect 1251 -1199 1256 -1194
rect 1174 -1216 1248 -1200
rect 1266 -1208 1296 -1152
rect 1331 -1162 1539 -1152
rect 3379 -1153 3391 -1152
rect 1357 -1192 1546 -1162
rect 1372 -1195 1546 -1192
rect 1365 -1198 1546 -1195
rect 1174 -1218 1187 -1216
rect 1202 -1218 1236 -1216
rect 1174 -1234 1248 -1218
rect 1275 -1222 1288 -1208
rect 1303 -1222 1319 -1206
rect 1365 -1211 1376 -1198
rect 1158 -1256 1159 -1240
rect 1174 -1256 1187 -1234
rect 1202 -1256 1232 -1234
rect 1275 -1238 1337 -1222
rect 1365 -1229 1376 -1213
rect 1381 -1218 1391 -1198
rect 1401 -1218 1415 -1198
rect 1418 -1211 1427 -1198
rect 1443 -1211 1452 -1198
rect 1381 -1229 1415 -1218
rect 1418 -1229 1427 -1213
rect 1443 -1229 1452 -1213
rect 1459 -1218 1469 -1198
rect 1479 -1218 1493 -1198
rect 1494 -1211 1505 -1198
rect 3379 -1200 3408 -1184
rect 1459 -1229 1493 -1218
rect 1494 -1229 1505 -1213
rect 3379 -1216 3424 -1200
rect 3379 -1218 3412 -1216
rect 1275 -1240 1288 -1238
rect 1303 -1240 1337 -1238
rect 1275 -1256 1337 -1240
rect 1381 -1245 1397 -1238
rect 1459 -1245 1489 -1234
rect 1537 -1240 1551 -1222
rect 1536 -1256 1551 -1240
rect 3379 -1234 3424 -1218
rect 3379 -1256 3408 -1234
rect 3435 -1256 3436 -1240
rect 3451 -1256 3464 -1096
rect 3494 -1200 3507 -1096
rect 3552 -1118 3553 -1108
rect 3568 -1118 3581 -1108
rect 3552 -1122 3581 -1118
rect 3586 -1122 3616 -1096
rect 3634 -1110 3650 -1108
rect 3722 -1110 3775 -1096
rect 3723 -1112 3787 -1110
rect 3830 -1112 3845 -1096
rect 3894 -1099 3924 -1096
rect 3894 -1102 3930 -1099
rect 3860 -1110 3876 -1108
rect 3634 -1122 3649 -1118
rect 3552 -1124 3649 -1122
rect 3677 -1124 3845 -1112
rect 3861 -1122 3876 -1118
rect 3894 -1121 3933 -1102
rect 3952 -1108 3959 -1107
rect 3958 -1115 3959 -1108
rect 3942 -1118 3943 -1115
rect 3958 -1118 3971 -1115
rect 3894 -1122 3924 -1121
rect 3933 -1122 3939 -1121
rect 3942 -1122 3971 -1118
rect 3861 -1123 3971 -1122
rect 3861 -1124 3977 -1123
rect 3536 -1132 3587 -1124
rect 3536 -1144 3561 -1132
rect 3568 -1144 3587 -1132
rect 3618 -1132 3668 -1124
rect 3618 -1140 3634 -1132
rect 3641 -1134 3668 -1132
rect 3677 -1134 3898 -1124
rect 3641 -1144 3898 -1134
rect 3927 -1132 3977 -1124
rect 3927 -1141 3943 -1132
rect 3536 -1152 3587 -1144
rect 3634 -1152 3898 -1144
rect 3924 -1144 3943 -1141
rect 3950 -1144 3977 -1132
rect 3924 -1152 3977 -1144
rect 3552 -1160 3553 -1152
rect 3568 -1160 3581 -1152
rect 3552 -1168 3568 -1160
rect 3549 -1175 3568 -1172
rect 3549 -1184 3571 -1175
rect 3522 -1194 3571 -1184
rect 3522 -1200 3552 -1194
rect 3571 -1199 3576 -1194
rect 3494 -1216 3568 -1200
rect 3586 -1208 3616 -1152
rect 3651 -1162 3859 -1152
rect 3894 -1156 3939 -1152
rect 3942 -1153 3943 -1152
rect 3958 -1153 3971 -1152
rect 3677 -1192 3866 -1162
rect 3692 -1195 3866 -1192
rect 3685 -1198 3866 -1195
rect 3494 -1218 3507 -1216
rect 3522 -1218 3556 -1216
rect 3494 -1234 3568 -1218
rect 3595 -1222 3608 -1208
rect 3623 -1222 3639 -1206
rect 3685 -1211 3696 -1198
rect 3478 -1256 3479 -1240
rect 3494 -1256 3507 -1234
rect 3522 -1256 3552 -1234
rect 3595 -1238 3657 -1222
rect 3685 -1229 3696 -1213
rect 3701 -1218 3711 -1198
rect 3721 -1218 3735 -1198
rect 3738 -1211 3747 -1198
rect 3763 -1211 3772 -1198
rect 3701 -1229 3735 -1218
rect 3738 -1229 3747 -1213
rect 3763 -1229 3772 -1213
rect 3779 -1218 3789 -1198
rect 3799 -1218 3813 -1198
rect 3814 -1211 3825 -1198
rect 3779 -1229 3813 -1218
rect 3814 -1229 3825 -1213
rect 3871 -1222 3887 -1206
rect 3894 -1208 3924 -1156
rect 3958 -1160 3959 -1153
rect 3943 -1168 3959 -1160
rect 3930 -1200 3943 -1181
rect 3958 -1200 3988 -1184
rect 3930 -1216 4004 -1200
rect 3930 -1218 3943 -1216
rect 3958 -1218 3992 -1216
rect 3595 -1240 3608 -1238
rect 3623 -1240 3657 -1238
rect 3595 -1256 3657 -1240
rect 3701 -1245 3717 -1238
rect 3779 -1245 3809 -1234
rect 3857 -1238 3903 -1222
rect 3930 -1234 4004 -1218
rect 3857 -1240 3891 -1238
rect 3856 -1256 3903 -1240
rect 3930 -1256 3943 -1234
rect 3958 -1256 3988 -1234
rect 4015 -1256 4016 -1240
rect 4031 -1256 4044 -1096
rect 4074 -1200 4087 -1096
rect 4132 -1118 4133 -1108
rect 4148 -1118 4161 -1108
rect 4132 -1122 4161 -1118
rect 4166 -1122 4196 -1096
rect 4214 -1110 4230 -1108
rect 4302 -1110 4355 -1096
rect 4303 -1112 4367 -1110
rect 4410 -1112 4425 -1096
rect 4474 -1099 4504 -1096
rect 4474 -1102 4510 -1099
rect 4440 -1110 4456 -1108
rect 4214 -1122 4229 -1118
rect 4132 -1124 4229 -1122
rect 4257 -1124 4425 -1112
rect 4441 -1122 4456 -1118
rect 4474 -1121 4513 -1102
rect 4532 -1108 4539 -1107
rect 4538 -1115 4539 -1108
rect 4522 -1118 4523 -1115
rect 4538 -1118 4551 -1115
rect 4474 -1122 4504 -1121
rect 4513 -1122 4519 -1121
rect 4522 -1122 4551 -1118
rect 4441 -1123 4551 -1122
rect 4441 -1124 4557 -1123
rect 4116 -1132 4167 -1124
rect 4116 -1144 4141 -1132
rect 4148 -1144 4167 -1132
rect 4198 -1132 4248 -1124
rect 4198 -1140 4214 -1132
rect 4221 -1134 4248 -1132
rect 4257 -1134 4478 -1124
rect 4221 -1144 4478 -1134
rect 4507 -1132 4557 -1124
rect 4507 -1141 4523 -1132
rect 4116 -1152 4167 -1144
rect 4214 -1152 4478 -1144
rect 4504 -1144 4523 -1141
rect 4530 -1144 4557 -1132
rect 4504 -1152 4557 -1144
rect 4132 -1160 4133 -1152
rect 4148 -1160 4161 -1152
rect 4132 -1168 4148 -1160
rect 4129 -1175 4148 -1172
rect 4129 -1184 4151 -1175
rect 4102 -1194 4151 -1184
rect 4102 -1200 4132 -1194
rect 4151 -1199 4156 -1194
rect 4074 -1216 4148 -1200
rect 4166 -1208 4196 -1152
rect 4231 -1162 4439 -1152
rect 4474 -1156 4519 -1152
rect 4522 -1153 4523 -1152
rect 4538 -1153 4551 -1152
rect 4257 -1192 4446 -1162
rect 4272 -1195 4446 -1192
rect 4265 -1198 4446 -1195
rect 4074 -1218 4087 -1216
rect 4102 -1218 4136 -1216
rect 4074 -1234 4148 -1218
rect 4175 -1222 4188 -1208
rect 4203 -1222 4219 -1206
rect 4265 -1211 4276 -1198
rect 4058 -1256 4059 -1240
rect 4074 -1256 4087 -1234
rect 4102 -1256 4132 -1234
rect 4175 -1238 4237 -1222
rect 4265 -1229 4276 -1213
rect 4281 -1218 4291 -1198
rect 4301 -1218 4315 -1198
rect 4318 -1211 4327 -1198
rect 4343 -1211 4352 -1198
rect 4281 -1229 4315 -1218
rect 4318 -1229 4327 -1213
rect 4343 -1229 4352 -1213
rect 4359 -1218 4369 -1198
rect 4379 -1218 4393 -1198
rect 4394 -1211 4405 -1198
rect 4359 -1229 4393 -1218
rect 4394 -1229 4405 -1213
rect 4451 -1222 4467 -1206
rect 4474 -1208 4504 -1156
rect 4538 -1160 4539 -1153
rect 4523 -1168 4539 -1160
rect 4510 -1200 4523 -1181
rect 4538 -1200 4568 -1184
rect 4510 -1216 4584 -1200
rect 4510 -1218 4523 -1216
rect 4538 -1218 4572 -1216
rect 4175 -1240 4188 -1238
rect 4203 -1240 4237 -1238
rect 4175 -1256 4237 -1240
rect 4281 -1245 4297 -1238
rect 4359 -1245 4389 -1234
rect 4437 -1238 4483 -1222
rect 4510 -1234 4584 -1218
rect 4437 -1240 4471 -1238
rect 4436 -1256 4483 -1240
rect 4510 -1256 4523 -1234
rect 4538 -1256 4568 -1234
rect 4595 -1256 4596 -1240
rect 4611 -1256 4624 -1096
rect 4654 -1200 4667 -1096
rect 4712 -1118 4713 -1108
rect 4728 -1118 4741 -1108
rect 4712 -1122 4741 -1118
rect 4746 -1122 4776 -1096
rect 4794 -1110 4810 -1108
rect 4882 -1110 4933 -1096
rect 4883 -1112 4947 -1110
rect 4990 -1112 5005 -1096
rect 5054 -1099 5084 -1096
rect 5054 -1102 5090 -1099
rect 5020 -1110 5036 -1108
rect 4794 -1122 4809 -1118
rect 4712 -1124 4809 -1122
rect 4837 -1124 5005 -1112
rect 5021 -1122 5036 -1118
rect 5054 -1121 5093 -1102
rect 5112 -1108 5119 -1107
rect 5118 -1115 5119 -1108
rect 5102 -1118 5103 -1115
rect 5118 -1118 5131 -1115
rect 5054 -1122 5084 -1121
rect 5093 -1122 5099 -1121
rect 5102 -1122 5131 -1118
rect 5021 -1123 5131 -1122
rect 5021 -1124 5137 -1123
rect 4696 -1132 4747 -1124
rect 4696 -1144 4721 -1132
rect 4728 -1144 4747 -1132
rect 4778 -1132 4828 -1124
rect 4778 -1140 4794 -1132
rect 4801 -1134 4828 -1132
rect 4837 -1134 5058 -1124
rect 4801 -1144 5058 -1134
rect 5087 -1132 5137 -1124
rect 5087 -1141 5103 -1132
rect 4696 -1152 4747 -1144
rect 4794 -1152 5058 -1144
rect 5084 -1144 5103 -1141
rect 5110 -1144 5137 -1132
rect 5084 -1152 5137 -1144
rect 4712 -1160 4713 -1152
rect 4728 -1160 4741 -1152
rect 4712 -1168 4728 -1160
rect 4709 -1175 4728 -1172
rect 4709 -1184 4731 -1175
rect 4682 -1194 4731 -1184
rect 4682 -1200 4712 -1194
rect 4731 -1199 4736 -1194
rect 4654 -1216 4728 -1200
rect 4746 -1208 4776 -1152
rect 4811 -1162 5019 -1152
rect 5054 -1156 5099 -1152
rect 5102 -1153 5103 -1152
rect 5118 -1153 5131 -1152
rect 4837 -1192 5026 -1162
rect 4852 -1195 5026 -1192
rect 4845 -1198 5026 -1195
rect 4654 -1218 4667 -1216
rect 4682 -1218 4716 -1216
rect 4654 -1234 4728 -1218
rect 4755 -1222 4768 -1208
rect 4783 -1222 4799 -1206
rect 4845 -1211 4856 -1198
rect 4638 -1256 4639 -1240
rect 4654 -1256 4667 -1234
rect 4682 -1256 4712 -1234
rect 4755 -1238 4817 -1222
rect 4845 -1229 4856 -1213
rect 4861 -1218 4871 -1198
rect 4881 -1218 4895 -1198
rect 4898 -1211 4907 -1198
rect 4923 -1211 4932 -1198
rect 4861 -1229 4895 -1218
rect 4898 -1229 4907 -1213
rect 4923 -1229 4932 -1213
rect 4939 -1218 4949 -1198
rect 4959 -1218 4973 -1198
rect 4974 -1211 4985 -1198
rect 4939 -1229 4973 -1218
rect 4974 -1229 4985 -1213
rect 5031 -1222 5047 -1206
rect 5054 -1208 5084 -1156
rect 5118 -1160 5119 -1153
rect 5103 -1168 5119 -1160
rect 5090 -1200 5103 -1181
rect 5118 -1200 5148 -1184
rect 5090 -1216 5164 -1200
rect 5090 -1218 5103 -1216
rect 5118 -1218 5152 -1216
rect 4755 -1240 4768 -1238
rect 4783 -1240 4817 -1238
rect 4755 -1256 4817 -1240
rect 4861 -1245 4877 -1238
rect 4939 -1245 4969 -1234
rect 5017 -1238 5063 -1222
rect 5090 -1234 5164 -1218
rect 5017 -1240 5051 -1238
rect 5016 -1256 5063 -1240
rect 5090 -1256 5103 -1234
rect 5118 -1256 5148 -1234
rect 5175 -1256 5176 -1240
rect 5191 -1256 5204 -1096
rect 5234 -1200 5247 -1096
rect 5292 -1118 5293 -1108
rect 5308 -1118 5321 -1108
rect 5292 -1122 5321 -1118
rect 5326 -1122 5356 -1096
rect 5374 -1110 5390 -1108
rect 5462 -1110 5513 -1096
rect 5463 -1112 5527 -1110
rect 5570 -1112 5585 -1096
rect 5634 -1099 5664 -1096
rect 5634 -1102 5670 -1099
rect 5600 -1110 5616 -1108
rect 5374 -1122 5389 -1118
rect 5292 -1124 5389 -1122
rect 5417 -1124 5585 -1112
rect 5601 -1122 5616 -1118
rect 5634 -1121 5673 -1102
rect 5692 -1108 5699 -1107
rect 5698 -1115 5699 -1108
rect 5682 -1118 5683 -1115
rect 5698 -1118 5711 -1115
rect 5634 -1122 5664 -1121
rect 5673 -1122 5679 -1121
rect 5682 -1122 5711 -1118
rect 5601 -1123 5711 -1122
rect 5601 -1124 5717 -1123
rect 5276 -1132 5327 -1124
rect 5276 -1144 5301 -1132
rect 5308 -1144 5327 -1132
rect 5358 -1132 5408 -1124
rect 5358 -1140 5374 -1132
rect 5381 -1134 5408 -1132
rect 5417 -1134 5638 -1124
rect 5381 -1144 5638 -1134
rect 5667 -1132 5717 -1124
rect 5667 -1141 5683 -1132
rect 5276 -1152 5327 -1144
rect 5374 -1152 5638 -1144
rect 5664 -1144 5683 -1141
rect 5690 -1144 5717 -1132
rect 5664 -1152 5717 -1144
rect 5292 -1160 5293 -1152
rect 5308 -1160 5321 -1152
rect 5292 -1168 5308 -1160
rect 5289 -1175 5308 -1172
rect 5289 -1184 5311 -1175
rect 5262 -1194 5311 -1184
rect 5262 -1200 5292 -1194
rect 5311 -1199 5316 -1194
rect 5234 -1216 5308 -1200
rect 5326 -1208 5356 -1152
rect 5391 -1162 5599 -1152
rect 5634 -1156 5679 -1152
rect 5682 -1153 5683 -1152
rect 5698 -1153 5711 -1152
rect 5417 -1192 5606 -1162
rect 5432 -1195 5606 -1192
rect 5425 -1198 5606 -1195
rect 5234 -1218 5247 -1216
rect 5262 -1218 5296 -1216
rect 5234 -1234 5308 -1218
rect 5335 -1222 5348 -1208
rect 5363 -1222 5379 -1206
rect 5425 -1211 5436 -1198
rect 5218 -1256 5219 -1240
rect 5234 -1256 5247 -1234
rect 5262 -1256 5292 -1234
rect 5335 -1238 5397 -1222
rect 5425 -1229 5436 -1213
rect 5441 -1218 5451 -1198
rect 5461 -1218 5475 -1198
rect 5478 -1211 5487 -1198
rect 5503 -1211 5512 -1198
rect 5441 -1229 5475 -1218
rect 5478 -1229 5487 -1213
rect 5503 -1229 5512 -1213
rect 5519 -1218 5529 -1198
rect 5539 -1218 5553 -1198
rect 5554 -1211 5565 -1198
rect 5519 -1229 5553 -1218
rect 5554 -1229 5565 -1213
rect 5611 -1222 5627 -1206
rect 5634 -1208 5664 -1156
rect 5698 -1160 5699 -1153
rect 5683 -1168 5699 -1160
rect 5670 -1200 5683 -1181
rect 5698 -1200 5728 -1184
rect 5670 -1216 5744 -1200
rect 5670 -1218 5683 -1216
rect 5698 -1218 5732 -1216
rect 5335 -1240 5348 -1238
rect 5363 -1240 5397 -1238
rect 5335 -1256 5397 -1240
rect 5441 -1245 5457 -1238
rect 5519 -1245 5549 -1234
rect 5597 -1238 5643 -1222
rect 5670 -1234 5744 -1218
rect 5597 -1240 5631 -1238
rect 5596 -1256 5643 -1240
rect 5670 -1256 5683 -1234
rect 5698 -1256 5728 -1234
rect 5755 -1256 5756 -1240
rect 5771 -1256 5784 -1096
rect 5814 -1200 5827 -1096
rect 5872 -1118 5873 -1108
rect 5888 -1118 5901 -1108
rect 5872 -1122 5901 -1118
rect 5906 -1122 5936 -1096
rect 5954 -1110 5970 -1108
rect 6042 -1110 6093 -1096
rect 6043 -1112 6107 -1110
rect 6150 -1112 6165 -1096
rect 6214 -1099 6244 -1096
rect 6214 -1102 6250 -1099
rect 6180 -1110 6196 -1108
rect 5954 -1122 5969 -1118
rect 5872 -1124 5969 -1122
rect 5997 -1124 6165 -1112
rect 6181 -1122 6196 -1118
rect 6214 -1121 6253 -1102
rect 6272 -1108 6279 -1107
rect 6278 -1115 6279 -1108
rect 6262 -1118 6263 -1115
rect 6278 -1118 6291 -1115
rect 6214 -1122 6244 -1121
rect 6253 -1122 6259 -1121
rect 6262 -1122 6291 -1118
rect 6181 -1123 6291 -1122
rect 6181 -1124 6297 -1123
rect 5856 -1132 5907 -1124
rect 5856 -1144 5881 -1132
rect 5888 -1144 5907 -1132
rect 5938 -1132 5988 -1124
rect 5938 -1140 5954 -1132
rect 5961 -1134 5988 -1132
rect 5997 -1134 6218 -1124
rect 5961 -1144 6218 -1134
rect 6247 -1132 6297 -1124
rect 6247 -1141 6263 -1132
rect 5856 -1152 5907 -1144
rect 5954 -1152 6218 -1144
rect 6244 -1144 6263 -1141
rect 6270 -1144 6297 -1132
rect 6244 -1152 6297 -1144
rect 5872 -1160 5873 -1152
rect 5888 -1160 5901 -1152
rect 5872 -1168 5888 -1160
rect 5869 -1175 5888 -1172
rect 5869 -1184 5891 -1175
rect 5842 -1194 5891 -1184
rect 5842 -1200 5872 -1194
rect 5891 -1199 5896 -1194
rect 5814 -1216 5888 -1200
rect 5906 -1208 5936 -1152
rect 5971 -1162 6179 -1152
rect 6214 -1156 6259 -1152
rect 6262 -1153 6263 -1152
rect 6278 -1153 6291 -1152
rect 5997 -1192 6186 -1162
rect 6012 -1195 6186 -1192
rect 6005 -1198 6186 -1195
rect 5814 -1218 5827 -1216
rect 5842 -1218 5876 -1216
rect 5814 -1234 5888 -1218
rect 5915 -1222 5928 -1208
rect 5943 -1222 5959 -1206
rect 6005 -1211 6016 -1198
rect 5798 -1256 5799 -1240
rect 5814 -1256 5827 -1234
rect 5842 -1256 5872 -1234
rect 5915 -1238 5977 -1222
rect 6005 -1229 6016 -1213
rect 6021 -1218 6031 -1198
rect 6041 -1218 6055 -1198
rect 6058 -1211 6067 -1198
rect 6083 -1211 6092 -1198
rect 6021 -1229 6055 -1218
rect 6058 -1229 6067 -1213
rect 6083 -1229 6092 -1213
rect 6099 -1218 6109 -1198
rect 6119 -1218 6133 -1198
rect 6134 -1211 6145 -1198
rect 6099 -1229 6133 -1218
rect 6134 -1229 6145 -1213
rect 6191 -1222 6207 -1206
rect 6214 -1208 6244 -1156
rect 6278 -1160 6279 -1153
rect 6263 -1168 6279 -1160
rect 6250 -1200 6263 -1181
rect 6278 -1200 6308 -1184
rect 6250 -1216 6324 -1200
rect 6250 -1218 6263 -1216
rect 6278 -1218 6312 -1216
rect 5915 -1240 5928 -1238
rect 5943 -1240 5977 -1238
rect 5915 -1256 5977 -1240
rect 6021 -1245 6037 -1238
rect 6099 -1245 6129 -1234
rect 6177 -1238 6223 -1222
rect 6250 -1234 6324 -1218
rect 6177 -1240 6211 -1238
rect 6176 -1256 6223 -1240
rect 6250 -1256 6263 -1234
rect 6278 -1256 6308 -1234
rect 6335 -1256 6336 -1240
rect 6351 -1256 6364 -1096
rect 6394 -1200 6407 -1096
rect 6452 -1118 6453 -1108
rect 6468 -1118 6481 -1108
rect 6452 -1122 6481 -1118
rect 6486 -1122 6516 -1096
rect 6534 -1110 6550 -1108
rect 6622 -1110 6673 -1096
rect 6623 -1112 6687 -1110
rect 6730 -1112 6745 -1096
rect 6794 -1099 6824 -1096
rect 6794 -1102 6830 -1099
rect 6760 -1110 6776 -1108
rect 6534 -1122 6549 -1118
rect 6452 -1124 6549 -1122
rect 6577 -1124 6745 -1112
rect 6761 -1122 6776 -1118
rect 6794 -1121 6833 -1102
rect 6852 -1108 6859 -1107
rect 6858 -1115 6859 -1108
rect 6842 -1118 6843 -1115
rect 6858 -1118 6871 -1115
rect 6794 -1122 6824 -1121
rect 6833 -1122 6839 -1121
rect 6842 -1122 6871 -1118
rect 6761 -1123 6871 -1122
rect 6761 -1124 6877 -1123
rect 6436 -1132 6487 -1124
rect 6436 -1144 6461 -1132
rect 6468 -1144 6487 -1132
rect 6518 -1132 6568 -1124
rect 6518 -1140 6534 -1132
rect 6541 -1134 6568 -1132
rect 6577 -1134 6798 -1124
rect 6541 -1144 6798 -1134
rect 6827 -1132 6877 -1124
rect 6827 -1141 6843 -1132
rect 6436 -1152 6487 -1144
rect 6534 -1152 6798 -1144
rect 6824 -1144 6843 -1141
rect 6850 -1144 6877 -1132
rect 6824 -1152 6877 -1144
rect 6452 -1160 6453 -1152
rect 6468 -1160 6481 -1152
rect 6452 -1168 6468 -1160
rect 6449 -1175 6468 -1172
rect 6449 -1184 6471 -1175
rect 6422 -1194 6471 -1184
rect 6422 -1200 6452 -1194
rect 6471 -1199 6476 -1194
rect 6394 -1216 6468 -1200
rect 6486 -1208 6516 -1152
rect 6551 -1162 6759 -1152
rect 6794 -1156 6839 -1152
rect 6842 -1153 6843 -1152
rect 6858 -1153 6871 -1152
rect 6577 -1192 6766 -1162
rect 6592 -1195 6766 -1192
rect 6585 -1198 6766 -1195
rect 6394 -1218 6407 -1216
rect 6422 -1218 6456 -1216
rect 6394 -1234 6468 -1218
rect 6495 -1222 6508 -1208
rect 6523 -1222 6539 -1206
rect 6585 -1211 6596 -1198
rect 6378 -1256 6379 -1240
rect 6394 -1256 6407 -1234
rect 6422 -1256 6452 -1234
rect 6495 -1238 6557 -1222
rect 6585 -1229 6596 -1213
rect 6601 -1218 6611 -1198
rect 6621 -1218 6635 -1198
rect 6638 -1211 6647 -1198
rect 6663 -1211 6672 -1198
rect 6601 -1229 6635 -1218
rect 6638 -1229 6647 -1213
rect 6663 -1229 6672 -1213
rect 6679 -1218 6689 -1198
rect 6699 -1218 6713 -1198
rect 6714 -1211 6725 -1198
rect 6679 -1229 6713 -1218
rect 6714 -1229 6725 -1213
rect 6771 -1222 6787 -1206
rect 6794 -1208 6824 -1156
rect 6858 -1160 6859 -1153
rect 6843 -1168 6859 -1160
rect 6830 -1200 6843 -1181
rect 6858 -1200 6888 -1184
rect 6830 -1216 6904 -1200
rect 6830 -1218 6843 -1216
rect 6858 -1218 6892 -1216
rect 6495 -1240 6508 -1238
rect 6523 -1240 6557 -1238
rect 6495 -1256 6557 -1240
rect 6601 -1245 6617 -1238
rect 6679 -1245 6709 -1234
rect 6757 -1238 6803 -1222
rect 6830 -1234 6904 -1218
rect 6757 -1240 6791 -1238
rect 6756 -1256 6803 -1240
rect 6830 -1256 6843 -1234
rect 6858 -1256 6888 -1234
rect 6915 -1256 6916 -1240
rect 6931 -1256 6944 -1096
rect -8 -1264 33 -1256
rect -8 -1290 7 -1264
rect 14 -1290 33 -1264
rect 97 -1268 159 -1256
rect 171 -1268 246 -1256
rect 304 -1268 379 -1256
rect 391 -1268 422 -1256
rect 428 -1268 463 -1256
rect 97 -1270 259 -1268
rect -8 -1298 33 -1290
rect 115 -1294 128 -1270
rect 143 -1272 158 -1270
rect -2 -1308 -1 -1298
rect 14 -1308 27 -1298
rect 42 -1308 72 -1294
rect 115 -1308 158 -1294
rect 182 -1297 189 -1290
rect 192 -1294 259 -1270
rect 291 -1270 463 -1268
rect 261 -1292 289 -1288
rect 291 -1292 371 -1270
rect 392 -1272 407 -1270
rect 261 -1294 371 -1292
rect 192 -1298 371 -1294
rect 165 -1308 195 -1298
rect 197 -1308 350 -1298
rect 358 -1308 388 -1298
rect 392 -1308 422 -1294
rect 450 -1308 463 -1270
rect 535 -1264 570 -1256
rect 535 -1290 536 -1264
rect 543 -1290 570 -1264
rect 478 -1308 508 -1294
rect 535 -1298 570 -1290
rect 572 -1264 613 -1256
rect 572 -1290 587 -1264
rect 594 -1290 613 -1264
rect 677 -1268 739 -1256
rect 751 -1268 826 -1256
rect 884 -1268 959 -1256
rect 971 -1268 1002 -1256
rect 1008 -1268 1043 -1256
rect 677 -1270 839 -1268
rect 572 -1298 613 -1290
rect 695 -1294 708 -1270
rect 723 -1272 738 -1270
rect 535 -1308 536 -1298
rect 551 -1308 564 -1298
rect 578 -1308 579 -1298
rect 594 -1308 607 -1298
rect 622 -1308 652 -1294
rect 695 -1308 738 -1294
rect 762 -1297 769 -1290
rect 772 -1294 839 -1270
rect 871 -1270 1043 -1268
rect 841 -1292 869 -1288
rect 871 -1292 951 -1270
rect 972 -1272 987 -1270
rect 841 -1294 951 -1292
rect 772 -1298 951 -1294
rect 745 -1308 775 -1298
rect 777 -1308 930 -1298
rect 938 -1308 968 -1298
rect 972 -1308 1002 -1294
rect 1030 -1308 1043 -1270
rect 1115 -1264 1150 -1256
rect 1115 -1290 1116 -1264
rect 1123 -1290 1150 -1264
rect 1058 -1308 1088 -1294
rect 1115 -1298 1150 -1290
rect 1152 -1264 1193 -1256
rect 1152 -1290 1167 -1264
rect 1174 -1290 1193 -1264
rect 1257 -1268 1319 -1256
rect 1331 -1268 1406 -1256
rect 1464 -1268 1539 -1256
rect 3435 -1264 3470 -1256
rect 1257 -1270 1419 -1268
rect 1152 -1298 1193 -1290
rect 1275 -1294 1288 -1270
rect 1303 -1272 1318 -1270
rect 1115 -1308 1116 -1298
rect 1131 -1308 1144 -1298
rect 1158 -1308 1159 -1298
rect 1174 -1308 1187 -1298
rect 1202 -1308 1232 -1294
rect 1275 -1308 1318 -1294
rect 1342 -1297 1349 -1290
rect 1352 -1294 1419 -1270
rect 1451 -1270 1551 -1268
rect 1421 -1292 1449 -1288
rect 1451 -1292 1531 -1270
rect 1421 -1294 1531 -1292
rect 3435 -1290 3436 -1264
rect 3443 -1290 3470 -1264
rect 1352 -1298 1531 -1294
rect 1325 -1308 1355 -1298
rect 1357 -1308 1510 -1298
rect 1518 -1308 1548 -1298
rect 3379 -1308 3408 -1294
rect 3435 -1298 3470 -1290
rect 3472 -1264 3513 -1256
rect 3472 -1290 3487 -1264
rect 3494 -1290 3513 -1264
rect 3577 -1268 3639 -1256
rect 3651 -1268 3726 -1256
rect 3784 -1268 3859 -1256
rect 3871 -1268 3902 -1256
rect 3908 -1268 3943 -1256
rect 3577 -1270 3739 -1268
rect 3472 -1298 3513 -1290
rect 3595 -1294 3608 -1270
rect 3623 -1272 3638 -1270
rect 3435 -1308 3436 -1298
rect 3451 -1308 3464 -1298
rect 3478 -1308 3479 -1298
rect 3494 -1308 3507 -1298
rect 3522 -1308 3552 -1294
rect 3595 -1308 3638 -1294
rect 3662 -1297 3669 -1290
rect 3672 -1294 3739 -1270
rect 3771 -1270 3943 -1268
rect 3741 -1292 3769 -1288
rect 3771 -1292 3851 -1270
rect 3872 -1272 3887 -1270
rect 3741 -1294 3851 -1292
rect 3672 -1298 3851 -1294
rect 3645 -1308 3675 -1298
rect 3677 -1308 3830 -1298
rect 3838 -1308 3868 -1298
rect 3872 -1308 3902 -1294
rect 3930 -1308 3943 -1270
rect 4015 -1264 4050 -1256
rect 4015 -1290 4016 -1264
rect 4023 -1290 4050 -1264
rect 3958 -1308 3988 -1294
rect 4015 -1298 4050 -1290
rect 4052 -1264 4093 -1256
rect 4052 -1290 4067 -1264
rect 4074 -1290 4093 -1264
rect 4157 -1268 4219 -1256
rect 4231 -1268 4306 -1256
rect 4364 -1268 4439 -1256
rect 4451 -1268 4482 -1256
rect 4488 -1268 4523 -1256
rect 4157 -1270 4319 -1268
rect 4052 -1298 4093 -1290
rect 4175 -1294 4188 -1270
rect 4203 -1272 4218 -1270
rect 4015 -1308 4016 -1298
rect 4031 -1308 4044 -1298
rect 4058 -1308 4059 -1298
rect 4074 -1308 4087 -1298
rect 4102 -1308 4132 -1294
rect 4175 -1308 4218 -1294
rect 4242 -1297 4249 -1290
rect 4252 -1294 4319 -1270
rect 4351 -1270 4523 -1268
rect 4321 -1292 4349 -1288
rect 4351 -1292 4431 -1270
rect 4452 -1272 4467 -1270
rect 4321 -1294 4431 -1292
rect 4252 -1298 4431 -1294
rect 4225 -1308 4255 -1298
rect 4257 -1308 4410 -1298
rect 4418 -1308 4448 -1298
rect 4452 -1308 4482 -1294
rect 4510 -1308 4523 -1270
rect 4595 -1264 4630 -1256
rect 4595 -1290 4596 -1264
rect 4603 -1290 4630 -1264
rect 4538 -1308 4568 -1294
rect 4595 -1298 4630 -1290
rect 4632 -1264 4673 -1256
rect 4632 -1290 4647 -1264
rect 4654 -1290 4673 -1264
rect 4737 -1268 4799 -1256
rect 4811 -1268 4886 -1256
rect 4944 -1268 5019 -1256
rect 5031 -1268 5062 -1256
rect 5068 -1268 5103 -1256
rect 4737 -1270 4899 -1268
rect 4632 -1298 4673 -1290
rect 4755 -1294 4768 -1270
rect 4783 -1272 4798 -1270
rect 4832 -1288 4899 -1270
rect 4931 -1270 5103 -1268
rect 4931 -1288 5011 -1270
rect 5032 -1272 5047 -1270
rect 4595 -1308 4596 -1298
rect 4611 -1308 4624 -1298
rect 4638 -1308 4639 -1298
rect 4654 -1308 4667 -1298
rect 4682 -1308 4712 -1294
rect 4755 -1308 4798 -1294
rect 4822 -1297 4829 -1290
rect 4832 -1298 5011 -1288
rect 4805 -1308 4835 -1298
rect 4837 -1308 4990 -1298
rect 4998 -1308 5028 -1298
rect 5032 -1308 5062 -1294
rect 5090 -1308 5103 -1270
rect 5175 -1264 5210 -1256
rect 5175 -1290 5176 -1264
rect 5183 -1290 5210 -1264
rect 5118 -1308 5148 -1294
rect 5175 -1298 5210 -1290
rect 5212 -1264 5253 -1256
rect 5212 -1290 5227 -1264
rect 5234 -1290 5253 -1264
rect 5317 -1268 5379 -1256
rect 5391 -1268 5466 -1256
rect 5524 -1268 5599 -1256
rect 5611 -1268 5642 -1256
rect 5648 -1268 5683 -1256
rect 5317 -1270 5479 -1268
rect 5212 -1298 5253 -1290
rect 5335 -1294 5348 -1270
rect 5363 -1272 5378 -1270
rect 5412 -1288 5479 -1270
rect 5511 -1270 5683 -1268
rect 5511 -1288 5591 -1270
rect 5612 -1272 5627 -1270
rect 5175 -1308 5176 -1298
rect 5191 -1308 5204 -1298
rect 5218 -1308 5219 -1298
rect 5234 -1308 5247 -1298
rect 5262 -1308 5292 -1294
rect 5335 -1308 5378 -1294
rect 5402 -1297 5409 -1290
rect 5412 -1298 5591 -1288
rect 5385 -1308 5415 -1298
rect 5417 -1308 5570 -1298
rect 5578 -1308 5608 -1298
rect 5612 -1308 5642 -1294
rect 5670 -1308 5683 -1270
rect 5755 -1264 5790 -1256
rect 5755 -1290 5756 -1264
rect 5763 -1290 5790 -1264
rect 5698 -1308 5728 -1294
rect 5755 -1298 5790 -1290
rect 5792 -1264 5833 -1256
rect 5792 -1290 5807 -1264
rect 5814 -1290 5833 -1264
rect 5897 -1268 5959 -1256
rect 5971 -1268 6046 -1256
rect 6104 -1268 6179 -1256
rect 6191 -1268 6222 -1256
rect 6228 -1268 6263 -1256
rect 5897 -1270 6059 -1268
rect 5792 -1298 5833 -1290
rect 5915 -1294 5928 -1270
rect 5943 -1272 5958 -1270
rect 5992 -1288 6059 -1270
rect 6091 -1270 6263 -1268
rect 6091 -1288 6171 -1270
rect 6192 -1272 6207 -1270
rect 5755 -1308 5756 -1298
rect 5771 -1308 5784 -1298
rect 5798 -1308 5799 -1298
rect 5814 -1308 5827 -1298
rect 5842 -1308 5872 -1294
rect 5915 -1308 5958 -1294
rect 5982 -1297 5989 -1290
rect 5992 -1298 6171 -1288
rect 5965 -1308 5995 -1298
rect 5997 -1308 6150 -1298
rect 6158 -1308 6188 -1298
rect 6192 -1308 6222 -1294
rect 6250 -1308 6263 -1270
rect 6335 -1264 6370 -1256
rect 6335 -1290 6336 -1264
rect 6343 -1290 6370 -1264
rect 6278 -1308 6308 -1294
rect 6335 -1298 6370 -1290
rect 6372 -1264 6413 -1256
rect 6372 -1290 6387 -1264
rect 6394 -1290 6413 -1264
rect 6477 -1268 6539 -1256
rect 6551 -1268 6626 -1256
rect 6684 -1268 6759 -1256
rect 6771 -1268 6802 -1256
rect 6808 -1268 6843 -1256
rect 6477 -1270 6639 -1268
rect 6372 -1298 6413 -1290
rect 6495 -1294 6508 -1270
rect 6523 -1272 6538 -1270
rect 6572 -1288 6639 -1270
rect 6671 -1270 6843 -1268
rect 6671 -1288 6751 -1270
rect 6772 -1272 6787 -1270
rect 6335 -1308 6336 -1298
rect 6351 -1308 6364 -1298
rect 6378 -1308 6379 -1298
rect 6394 -1308 6407 -1298
rect 6422 -1308 6452 -1294
rect 6495 -1308 6538 -1294
rect 6562 -1297 6569 -1290
rect 6572 -1298 6751 -1288
rect 6545 -1308 6575 -1298
rect 6577 -1308 6730 -1298
rect 6738 -1308 6768 -1298
rect 6772 -1308 6802 -1294
rect 6830 -1308 6843 -1270
rect 6915 -1264 6950 -1256
rect 6915 -1290 6916 -1264
rect 6923 -1290 6950 -1264
rect 6858 -1308 6888 -1294
rect 6915 -1298 6950 -1290
rect 6915 -1308 6916 -1298
rect 6931 -1308 6944 -1298
rect -2 -1314 1551 -1308
rect -1 -1322 1551 -1314
rect 3379 -1322 6944 -1308
rect 14 -1352 27 -1322
rect 42 -1340 72 -1322
rect 115 -1336 129 -1322
rect 165 -1336 385 -1322
rect 116 -1338 129 -1336
rect 82 -1350 97 -1338
rect 79 -1352 101 -1350
rect 106 -1352 136 -1338
rect 197 -1340 350 -1336
rect 179 -1352 371 -1340
rect 414 -1352 444 -1338
rect 450 -1352 463 -1322
rect 478 -1340 508 -1322
rect 551 -1352 564 -1322
rect 594 -1352 607 -1322
rect 622 -1340 652 -1322
rect 695 -1336 709 -1322
rect 745 -1336 965 -1322
rect 696 -1338 709 -1336
rect 662 -1350 677 -1338
rect 659 -1352 681 -1350
rect 686 -1352 716 -1338
rect 777 -1340 930 -1336
rect 759 -1352 951 -1340
rect 994 -1352 1024 -1338
rect 1030 -1352 1043 -1322
rect 1058 -1340 1088 -1322
rect 1131 -1352 1144 -1322
rect 1174 -1352 1187 -1322
rect 1202 -1340 1232 -1322
rect 1275 -1336 1289 -1322
rect 1325 -1336 1545 -1322
rect 1276 -1338 1289 -1336
rect 1242 -1350 1257 -1338
rect 1239 -1352 1261 -1350
rect 1266 -1352 1296 -1338
rect 1357 -1340 1510 -1336
rect 3379 -1340 3408 -1322
rect 1339 -1352 1531 -1340
rect 3451 -1352 3464 -1322
rect 3494 -1352 3507 -1322
rect 3522 -1340 3552 -1322
rect 3595 -1336 3609 -1322
rect 3645 -1336 3865 -1322
rect 3596 -1338 3609 -1336
rect 3562 -1350 3577 -1338
rect 3559 -1352 3581 -1350
rect 3586 -1352 3616 -1338
rect 3677 -1340 3830 -1336
rect 3659 -1352 3851 -1340
rect 3894 -1352 3924 -1338
rect 3930 -1352 3943 -1322
rect 3958 -1340 3988 -1322
rect 4031 -1352 4044 -1322
rect 4074 -1352 4087 -1322
rect 4102 -1340 4132 -1322
rect 4175 -1336 4189 -1322
rect 4225 -1336 4445 -1322
rect 4176 -1338 4189 -1336
rect 4142 -1350 4157 -1338
rect 4139 -1352 4161 -1350
rect 4166 -1352 4196 -1338
rect 4257 -1340 4410 -1336
rect 4239 -1352 4431 -1340
rect 4474 -1352 4504 -1338
rect 4510 -1352 4523 -1322
rect 4538 -1340 4568 -1322
rect 4611 -1352 4624 -1322
rect 4654 -1352 4667 -1322
rect 4682 -1340 4712 -1322
rect 4755 -1336 4769 -1322
rect 4805 -1336 5025 -1322
rect 4756 -1338 4769 -1336
rect 4722 -1350 4737 -1338
rect 4719 -1352 4741 -1350
rect 4746 -1352 4776 -1338
rect 4837 -1340 4990 -1336
rect 4819 -1352 5011 -1340
rect 5054 -1352 5084 -1338
rect 5090 -1352 5103 -1322
rect 5118 -1340 5148 -1322
rect 5191 -1352 5204 -1322
rect 5234 -1352 5247 -1322
rect 5262 -1340 5292 -1322
rect 5335 -1336 5349 -1322
rect 5385 -1336 5605 -1322
rect 5336 -1338 5349 -1336
rect 5302 -1350 5317 -1338
rect 5299 -1352 5321 -1350
rect 5326 -1352 5356 -1338
rect 5417 -1340 5570 -1336
rect 5399 -1352 5591 -1340
rect 5634 -1352 5664 -1338
rect 5670 -1352 5683 -1322
rect 5698 -1340 5728 -1322
rect 5771 -1352 5784 -1322
rect 5814 -1352 5827 -1322
rect 5842 -1340 5872 -1322
rect 5915 -1336 5929 -1322
rect 5965 -1336 6185 -1322
rect 5916 -1338 5929 -1336
rect 5882 -1350 5897 -1338
rect 5879 -1352 5901 -1350
rect 5906 -1352 5936 -1338
rect 5997 -1340 6150 -1336
rect 5979 -1352 6171 -1340
rect 6214 -1352 6244 -1338
rect 6250 -1352 6263 -1322
rect 6278 -1340 6308 -1322
rect 6351 -1352 6364 -1322
rect 6394 -1352 6407 -1322
rect 6422 -1340 6452 -1322
rect 6495 -1336 6509 -1322
rect 6545 -1336 6765 -1322
rect 6496 -1338 6509 -1336
rect 6462 -1350 6477 -1338
rect 6459 -1352 6481 -1350
rect 6486 -1352 6516 -1338
rect 6577 -1340 6730 -1336
rect 6559 -1352 6751 -1340
rect 6794 -1352 6824 -1338
rect 6830 -1352 6843 -1322
rect 6858 -1340 6888 -1322
rect 6931 -1352 6944 -1322
rect -1 -1366 1551 -1352
rect 3379 -1366 6944 -1352
rect 14 -1470 27 -1366
rect 72 -1388 73 -1378
rect 88 -1388 101 -1378
rect 72 -1392 101 -1388
rect 106 -1392 136 -1366
rect 154 -1380 170 -1378
rect 242 -1380 295 -1366
rect 243 -1382 307 -1380
rect 350 -1382 365 -1366
rect 414 -1369 444 -1366
rect 414 -1372 450 -1369
rect 380 -1380 396 -1378
rect 154 -1392 169 -1388
rect 72 -1394 169 -1392
rect 197 -1394 365 -1382
rect 381 -1392 396 -1388
rect 414 -1391 453 -1372
rect 472 -1378 479 -1377
rect 478 -1385 479 -1378
rect 462 -1388 463 -1385
rect 478 -1388 491 -1385
rect 414 -1392 444 -1391
rect 453 -1392 459 -1391
rect 462 -1392 491 -1388
rect 381 -1393 491 -1392
rect 381 -1394 497 -1393
rect 56 -1402 107 -1394
rect 56 -1414 81 -1402
rect 88 -1414 107 -1402
rect 138 -1402 188 -1394
rect 138 -1410 154 -1402
rect 161 -1404 188 -1402
rect 197 -1404 418 -1394
rect 161 -1414 418 -1404
rect 447 -1402 497 -1394
rect 447 -1411 463 -1402
rect 56 -1422 107 -1414
rect 154 -1422 418 -1414
rect 444 -1414 463 -1411
rect 470 -1414 497 -1402
rect 444 -1422 497 -1414
rect 72 -1430 73 -1422
rect 88 -1430 101 -1422
rect 72 -1438 88 -1430
rect 69 -1445 88 -1442
rect 69 -1454 91 -1445
rect 42 -1464 91 -1454
rect 42 -1470 72 -1464
rect 91 -1469 96 -1464
rect 14 -1486 88 -1470
rect 106 -1478 136 -1422
rect 171 -1432 379 -1422
rect 414 -1426 459 -1422
rect 462 -1423 463 -1422
rect 478 -1423 491 -1422
rect 197 -1462 386 -1432
rect 212 -1465 386 -1462
rect 205 -1468 386 -1465
rect 14 -1488 27 -1486
rect 42 -1488 76 -1486
rect 14 -1504 88 -1488
rect 115 -1492 128 -1478
rect 143 -1492 159 -1476
rect 205 -1481 216 -1468
rect -2 -1526 -1 -1510
rect 14 -1526 27 -1504
rect 42 -1526 72 -1504
rect 115 -1508 177 -1492
rect 205 -1499 216 -1483
rect 221 -1488 231 -1468
rect 241 -1488 255 -1468
rect 258 -1481 267 -1468
rect 283 -1481 292 -1468
rect 221 -1499 255 -1488
rect 258 -1499 267 -1483
rect 283 -1499 292 -1483
rect 299 -1488 309 -1468
rect 319 -1488 333 -1468
rect 334 -1481 345 -1468
rect 299 -1499 333 -1488
rect 334 -1499 345 -1483
rect 391 -1492 407 -1476
rect 414 -1478 444 -1426
rect 478 -1430 479 -1423
rect 463 -1438 479 -1430
rect 450 -1470 463 -1451
rect 478 -1470 508 -1454
rect 450 -1486 524 -1470
rect 450 -1488 463 -1486
rect 478 -1488 512 -1486
rect 115 -1510 128 -1508
rect 143 -1510 177 -1508
rect 115 -1526 177 -1510
rect 221 -1515 237 -1508
rect 299 -1515 329 -1504
rect 377 -1508 423 -1492
rect 450 -1504 524 -1488
rect 377 -1510 411 -1508
rect 376 -1526 423 -1510
rect 450 -1526 463 -1504
rect 478 -1526 508 -1504
rect 535 -1526 536 -1510
rect 551 -1526 564 -1366
rect 594 -1470 607 -1366
rect 652 -1388 653 -1378
rect 668 -1388 681 -1378
rect 652 -1392 681 -1388
rect 686 -1392 716 -1366
rect 734 -1380 750 -1378
rect 822 -1380 875 -1366
rect 823 -1382 887 -1380
rect 930 -1382 945 -1366
rect 994 -1369 1024 -1366
rect 994 -1372 1030 -1369
rect 960 -1380 976 -1378
rect 734 -1392 749 -1388
rect 652 -1394 749 -1392
rect 777 -1394 945 -1382
rect 961 -1392 976 -1388
rect 994 -1391 1033 -1372
rect 1052 -1378 1059 -1377
rect 1058 -1385 1059 -1378
rect 1042 -1388 1043 -1385
rect 1058 -1388 1071 -1385
rect 994 -1392 1024 -1391
rect 1033 -1392 1039 -1391
rect 1042 -1392 1071 -1388
rect 961 -1393 1071 -1392
rect 961 -1394 1077 -1393
rect 636 -1402 687 -1394
rect 636 -1414 661 -1402
rect 668 -1414 687 -1402
rect 718 -1402 768 -1394
rect 718 -1410 734 -1402
rect 741 -1404 768 -1402
rect 777 -1404 998 -1394
rect 741 -1414 998 -1404
rect 1027 -1402 1077 -1394
rect 1027 -1411 1043 -1402
rect 636 -1422 687 -1414
rect 734 -1422 998 -1414
rect 1024 -1414 1043 -1411
rect 1050 -1414 1077 -1402
rect 1024 -1422 1077 -1414
rect 652 -1430 653 -1422
rect 668 -1430 681 -1422
rect 652 -1438 668 -1430
rect 649 -1445 668 -1442
rect 649 -1454 671 -1445
rect 622 -1464 671 -1454
rect 622 -1470 652 -1464
rect 671 -1469 676 -1464
rect 594 -1486 668 -1470
rect 686 -1478 716 -1422
rect 751 -1432 959 -1422
rect 994 -1426 1039 -1422
rect 1042 -1423 1043 -1422
rect 1058 -1423 1071 -1422
rect 777 -1462 966 -1432
rect 792 -1465 966 -1462
rect 785 -1468 966 -1465
rect 594 -1488 607 -1486
rect 622 -1488 656 -1486
rect 594 -1504 668 -1488
rect 695 -1492 708 -1478
rect 723 -1492 739 -1476
rect 785 -1481 796 -1468
rect 578 -1526 579 -1510
rect 594 -1526 607 -1504
rect 622 -1526 652 -1504
rect 695 -1508 757 -1492
rect 785 -1499 796 -1483
rect 801 -1488 811 -1468
rect 821 -1488 835 -1468
rect 838 -1481 847 -1468
rect 863 -1481 872 -1468
rect 801 -1499 835 -1488
rect 838 -1499 847 -1483
rect 863 -1499 872 -1483
rect 879 -1488 889 -1468
rect 899 -1488 913 -1468
rect 914 -1481 925 -1468
rect 879 -1499 913 -1488
rect 914 -1499 925 -1483
rect 971 -1492 987 -1476
rect 994 -1478 1024 -1426
rect 1058 -1430 1059 -1423
rect 1043 -1438 1059 -1430
rect 1030 -1470 1043 -1451
rect 1058 -1470 1088 -1454
rect 1030 -1486 1104 -1470
rect 1030 -1488 1043 -1486
rect 1058 -1488 1092 -1486
rect 695 -1510 708 -1508
rect 723 -1510 757 -1508
rect 695 -1526 757 -1510
rect 801 -1515 817 -1508
rect 879 -1515 909 -1504
rect 957 -1508 1003 -1492
rect 1030 -1504 1104 -1488
rect 957 -1510 991 -1508
rect 956 -1526 1003 -1510
rect 1030 -1526 1043 -1504
rect 1058 -1526 1088 -1504
rect 1115 -1526 1116 -1510
rect 1131 -1526 1144 -1366
rect 1174 -1470 1187 -1366
rect 1232 -1388 1233 -1378
rect 1248 -1388 1261 -1378
rect 1232 -1392 1261 -1388
rect 1266 -1392 1296 -1366
rect 1314 -1380 1330 -1378
rect 1402 -1380 1455 -1366
rect 1403 -1382 1467 -1380
rect 1510 -1382 1525 -1366
rect 1540 -1380 1551 -1378
rect 1314 -1392 1329 -1388
rect 1232 -1394 1329 -1392
rect 1357 -1394 1525 -1382
rect 1541 -1394 1551 -1388
rect 1216 -1402 1267 -1394
rect 1216 -1414 1241 -1402
rect 1248 -1414 1267 -1402
rect 1298 -1402 1348 -1394
rect 1298 -1410 1314 -1402
rect 1321 -1404 1348 -1402
rect 1357 -1404 1551 -1394
rect 1321 -1414 1551 -1404
rect 1216 -1422 1267 -1414
rect 1314 -1422 1551 -1414
rect 3379 -1393 3391 -1385
rect 3379 -1422 3397 -1393
rect 1232 -1430 1233 -1422
rect 1248 -1430 1261 -1422
rect 1232 -1438 1248 -1430
rect 1229 -1445 1248 -1442
rect 1229 -1454 1251 -1445
rect 1202 -1464 1251 -1454
rect 1202 -1470 1232 -1464
rect 1251 -1469 1256 -1464
rect 1174 -1486 1248 -1470
rect 1266 -1478 1296 -1422
rect 1331 -1432 1539 -1422
rect 3379 -1423 3391 -1422
rect 1357 -1462 1546 -1432
rect 1372 -1465 1546 -1462
rect 1365 -1468 1546 -1465
rect 1174 -1488 1187 -1486
rect 1202 -1488 1236 -1486
rect 1174 -1504 1248 -1488
rect 1275 -1492 1288 -1478
rect 1303 -1492 1319 -1476
rect 1365 -1481 1376 -1468
rect 1158 -1526 1159 -1510
rect 1174 -1526 1187 -1504
rect 1202 -1526 1232 -1504
rect 1275 -1508 1337 -1492
rect 1365 -1499 1376 -1483
rect 1381 -1488 1391 -1468
rect 1401 -1488 1415 -1468
rect 1418 -1481 1427 -1468
rect 1443 -1481 1452 -1468
rect 1381 -1499 1415 -1488
rect 1418 -1499 1427 -1483
rect 1443 -1499 1452 -1483
rect 1459 -1488 1469 -1468
rect 1479 -1488 1493 -1468
rect 1494 -1481 1505 -1468
rect 3379 -1470 3408 -1454
rect 1459 -1499 1493 -1488
rect 1494 -1499 1505 -1483
rect 3379 -1486 3424 -1470
rect 3379 -1488 3412 -1486
rect 1275 -1510 1288 -1508
rect 1303 -1510 1337 -1508
rect 1275 -1526 1337 -1510
rect 1381 -1515 1397 -1508
rect 1459 -1515 1489 -1504
rect 1537 -1510 1551 -1492
rect 1536 -1526 1551 -1510
rect 3379 -1504 3424 -1488
rect 3379 -1526 3408 -1504
rect 3435 -1526 3436 -1510
rect 3451 -1526 3464 -1366
rect 3494 -1470 3507 -1366
rect 3552 -1388 3553 -1378
rect 3568 -1388 3581 -1378
rect 3552 -1392 3581 -1388
rect 3586 -1392 3616 -1366
rect 3634 -1380 3650 -1378
rect 3722 -1380 3775 -1366
rect 3723 -1382 3787 -1380
rect 3830 -1382 3845 -1366
rect 3894 -1369 3924 -1366
rect 3894 -1372 3930 -1369
rect 3860 -1380 3876 -1378
rect 3634 -1392 3649 -1388
rect 3552 -1394 3649 -1392
rect 3677 -1394 3845 -1382
rect 3861 -1392 3876 -1388
rect 3894 -1391 3933 -1372
rect 3952 -1378 3959 -1377
rect 3958 -1385 3959 -1378
rect 3942 -1388 3943 -1385
rect 3958 -1388 3971 -1385
rect 3894 -1392 3924 -1391
rect 3933 -1392 3939 -1391
rect 3942 -1392 3971 -1388
rect 3861 -1393 3971 -1392
rect 3861 -1394 3977 -1393
rect 3536 -1402 3587 -1394
rect 3536 -1414 3561 -1402
rect 3568 -1414 3587 -1402
rect 3618 -1402 3668 -1394
rect 3618 -1410 3634 -1402
rect 3641 -1404 3668 -1402
rect 3677 -1404 3898 -1394
rect 3641 -1414 3898 -1404
rect 3927 -1402 3977 -1394
rect 3927 -1411 3943 -1402
rect 3536 -1422 3587 -1414
rect 3634 -1422 3898 -1414
rect 3924 -1414 3943 -1411
rect 3950 -1414 3977 -1402
rect 3924 -1422 3977 -1414
rect 3552 -1430 3553 -1422
rect 3568 -1430 3581 -1422
rect 3552 -1438 3568 -1430
rect 3549 -1445 3568 -1442
rect 3549 -1454 3571 -1445
rect 3522 -1464 3571 -1454
rect 3522 -1470 3552 -1464
rect 3571 -1469 3576 -1464
rect 3494 -1486 3568 -1470
rect 3586 -1478 3616 -1422
rect 3651 -1432 3859 -1422
rect 3894 -1426 3939 -1422
rect 3942 -1423 3943 -1422
rect 3958 -1423 3971 -1422
rect 3677 -1462 3866 -1432
rect 3692 -1465 3866 -1462
rect 3685 -1468 3866 -1465
rect 3494 -1488 3507 -1486
rect 3522 -1488 3556 -1486
rect 3494 -1504 3568 -1488
rect 3595 -1492 3608 -1478
rect 3623 -1492 3639 -1476
rect 3685 -1481 3696 -1468
rect 3478 -1526 3479 -1510
rect 3494 -1526 3507 -1504
rect 3522 -1526 3552 -1504
rect 3595 -1508 3657 -1492
rect 3685 -1499 3696 -1483
rect 3701 -1488 3711 -1468
rect 3721 -1488 3735 -1468
rect 3738 -1481 3747 -1468
rect 3763 -1481 3772 -1468
rect 3701 -1499 3735 -1488
rect 3738 -1499 3747 -1483
rect 3763 -1499 3772 -1483
rect 3779 -1488 3789 -1468
rect 3799 -1488 3813 -1468
rect 3814 -1481 3825 -1468
rect 3779 -1499 3813 -1488
rect 3814 -1499 3825 -1483
rect 3871 -1492 3887 -1476
rect 3894 -1478 3924 -1426
rect 3958 -1430 3959 -1423
rect 3943 -1438 3959 -1430
rect 3930 -1470 3943 -1451
rect 3958 -1470 3988 -1454
rect 3930 -1486 4004 -1470
rect 3930 -1488 3943 -1486
rect 3958 -1488 3992 -1486
rect 3595 -1510 3608 -1508
rect 3623 -1510 3657 -1508
rect 3595 -1526 3657 -1510
rect 3701 -1515 3717 -1508
rect 3779 -1515 3809 -1504
rect 3857 -1508 3903 -1492
rect 3930 -1504 4004 -1488
rect 3857 -1510 3891 -1508
rect 3856 -1526 3903 -1510
rect 3930 -1526 3943 -1504
rect 3958 -1526 3988 -1504
rect 4015 -1526 4016 -1510
rect 4031 -1526 4044 -1366
rect 4074 -1470 4087 -1366
rect 4132 -1388 4133 -1378
rect 4148 -1388 4161 -1378
rect 4132 -1392 4161 -1388
rect 4166 -1392 4196 -1366
rect 4214 -1380 4230 -1378
rect 4302 -1380 4355 -1366
rect 4303 -1382 4367 -1380
rect 4410 -1382 4425 -1366
rect 4474 -1369 4504 -1366
rect 4474 -1372 4510 -1369
rect 4440 -1380 4456 -1378
rect 4214 -1392 4229 -1388
rect 4132 -1394 4229 -1392
rect 4257 -1394 4425 -1382
rect 4441 -1392 4456 -1388
rect 4474 -1391 4513 -1372
rect 4532 -1378 4539 -1377
rect 4538 -1385 4539 -1378
rect 4522 -1388 4523 -1385
rect 4538 -1388 4551 -1385
rect 4474 -1392 4504 -1391
rect 4513 -1392 4519 -1391
rect 4522 -1392 4551 -1388
rect 4441 -1393 4551 -1392
rect 4441 -1394 4557 -1393
rect 4116 -1402 4167 -1394
rect 4116 -1414 4141 -1402
rect 4148 -1414 4167 -1402
rect 4198 -1402 4248 -1394
rect 4198 -1410 4214 -1402
rect 4221 -1404 4248 -1402
rect 4257 -1404 4478 -1394
rect 4221 -1414 4478 -1404
rect 4507 -1402 4557 -1394
rect 4507 -1411 4523 -1402
rect 4116 -1422 4167 -1414
rect 4214 -1422 4478 -1414
rect 4504 -1414 4523 -1411
rect 4530 -1414 4557 -1402
rect 4504 -1422 4557 -1414
rect 4132 -1430 4133 -1422
rect 4148 -1430 4161 -1422
rect 4132 -1438 4148 -1430
rect 4129 -1445 4148 -1442
rect 4129 -1454 4151 -1445
rect 4102 -1464 4151 -1454
rect 4102 -1470 4132 -1464
rect 4151 -1469 4156 -1464
rect 4074 -1486 4148 -1470
rect 4166 -1478 4196 -1422
rect 4231 -1432 4439 -1422
rect 4474 -1426 4519 -1422
rect 4522 -1423 4523 -1422
rect 4538 -1423 4551 -1422
rect 4257 -1462 4446 -1432
rect 4272 -1465 4446 -1462
rect 4265 -1468 4446 -1465
rect 4074 -1488 4087 -1486
rect 4102 -1488 4136 -1486
rect 4074 -1504 4148 -1488
rect 4175 -1492 4188 -1478
rect 4203 -1492 4219 -1476
rect 4265 -1481 4276 -1468
rect 4058 -1526 4059 -1510
rect 4074 -1526 4087 -1504
rect 4102 -1526 4132 -1504
rect 4175 -1508 4237 -1492
rect 4265 -1499 4276 -1483
rect 4281 -1488 4291 -1468
rect 4301 -1488 4315 -1468
rect 4318 -1481 4327 -1468
rect 4343 -1481 4352 -1468
rect 4281 -1499 4315 -1488
rect 4318 -1499 4327 -1483
rect 4343 -1499 4352 -1483
rect 4359 -1488 4369 -1468
rect 4379 -1488 4393 -1468
rect 4394 -1481 4405 -1468
rect 4359 -1499 4393 -1488
rect 4394 -1499 4405 -1483
rect 4451 -1492 4467 -1476
rect 4474 -1478 4504 -1426
rect 4538 -1430 4539 -1423
rect 4523 -1438 4539 -1430
rect 4510 -1470 4523 -1451
rect 4538 -1470 4568 -1454
rect 4510 -1486 4584 -1470
rect 4510 -1488 4523 -1486
rect 4538 -1488 4572 -1486
rect 4175 -1510 4188 -1508
rect 4203 -1510 4237 -1508
rect 4175 -1526 4237 -1510
rect 4281 -1515 4297 -1508
rect 4359 -1515 4389 -1504
rect 4437 -1508 4483 -1492
rect 4510 -1504 4584 -1488
rect 4437 -1510 4471 -1508
rect 4436 -1526 4483 -1510
rect 4510 -1526 4523 -1504
rect 4538 -1526 4568 -1504
rect 4595 -1526 4596 -1510
rect 4611 -1526 4624 -1366
rect 4654 -1470 4667 -1366
rect 4712 -1388 4713 -1378
rect 4728 -1388 4741 -1378
rect 4712 -1392 4741 -1388
rect 4746 -1392 4776 -1366
rect 4794 -1380 4810 -1378
rect 4882 -1380 4933 -1366
rect 4883 -1382 4947 -1380
rect 4990 -1382 5005 -1366
rect 5054 -1369 5084 -1366
rect 5054 -1372 5090 -1369
rect 5020 -1380 5036 -1378
rect 4794 -1392 4809 -1388
rect 4712 -1394 4809 -1392
rect 4837 -1394 5005 -1382
rect 5021 -1392 5036 -1388
rect 5054 -1391 5093 -1372
rect 5112 -1378 5119 -1377
rect 5118 -1385 5119 -1378
rect 5102 -1388 5103 -1385
rect 5118 -1388 5131 -1385
rect 5054 -1392 5084 -1391
rect 5093 -1392 5099 -1391
rect 5102 -1392 5131 -1388
rect 5021 -1393 5131 -1392
rect 5021 -1394 5137 -1393
rect 4696 -1402 4747 -1394
rect 4696 -1414 4721 -1402
rect 4728 -1414 4747 -1402
rect 4778 -1402 4828 -1394
rect 4778 -1410 4794 -1402
rect 4801 -1404 4828 -1402
rect 4837 -1404 5058 -1394
rect 4801 -1414 5058 -1404
rect 5087 -1402 5137 -1394
rect 5087 -1411 5103 -1402
rect 4696 -1422 4747 -1414
rect 4794 -1422 5058 -1414
rect 5084 -1414 5103 -1411
rect 5110 -1414 5137 -1402
rect 5084 -1422 5137 -1414
rect 4712 -1430 4713 -1422
rect 4728 -1430 4741 -1422
rect 4712 -1438 4728 -1430
rect 4709 -1445 4728 -1442
rect 4709 -1454 4731 -1445
rect 4682 -1464 4731 -1454
rect 4682 -1470 4712 -1464
rect 4731 -1469 4736 -1464
rect 4654 -1486 4728 -1470
rect 4746 -1478 4776 -1422
rect 4811 -1432 5019 -1422
rect 5054 -1426 5099 -1422
rect 5102 -1423 5103 -1422
rect 5118 -1423 5131 -1422
rect 4837 -1462 5026 -1432
rect 4852 -1465 5026 -1462
rect 4845 -1468 5026 -1465
rect 4654 -1488 4667 -1486
rect 4682 -1488 4716 -1486
rect 4654 -1504 4728 -1488
rect 4755 -1492 4768 -1478
rect 4783 -1492 4799 -1476
rect 4845 -1481 4856 -1468
rect 4638 -1526 4639 -1510
rect 4654 -1526 4667 -1504
rect 4682 -1526 4712 -1504
rect 4755 -1508 4817 -1492
rect 4845 -1499 4856 -1483
rect 4861 -1488 4871 -1468
rect 4881 -1488 4895 -1468
rect 4898 -1481 4907 -1468
rect 4923 -1481 4932 -1468
rect 4861 -1499 4895 -1488
rect 4898 -1499 4907 -1483
rect 4923 -1499 4932 -1483
rect 4939 -1488 4949 -1468
rect 4959 -1488 4973 -1468
rect 4974 -1481 4985 -1468
rect 4939 -1499 4973 -1488
rect 4974 -1499 4985 -1483
rect 5031 -1492 5047 -1476
rect 5054 -1478 5084 -1426
rect 5118 -1430 5119 -1423
rect 5103 -1438 5119 -1430
rect 5090 -1470 5103 -1451
rect 5118 -1470 5148 -1454
rect 5090 -1486 5164 -1470
rect 5090 -1488 5103 -1486
rect 5118 -1488 5152 -1486
rect 4755 -1510 4768 -1508
rect 4783 -1510 4817 -1508
rect 4755 -1526 4817 -1510
rect 4861 -1515 4877 -1508
rect 4939 -1515 4969 -1504
rect 5017 -1508 5063 -1492
rect 5090 -1504 5164 -1488
rect 5017 -1510 5051 -1508
rect 5016 -1526 5063 -1510
rect 5090 -1526 5103 -1504
rect 5118 -1526 5148 -1504
rect 5175 -1526 5176 -1510
rect 5191 -1526 5204 -1366
rect 5234 -1470 5247 -1366
rect 5292 -1388 5293 -1378
rect 5308 -1388 5321 -1378
rect 5292 -1392 5321 -1388
rect 5326 -1392 5356 -1366
rect 5374 -1380 5390 -1378
rect 5462 -1380 5513 -1366
rect 5463 -1382 5527 -1380
rect 5570 -1382 5585 -1366
rect 5634 -1369 5664 -1366
rect 5634 -1372 5670 -1369
rect 5600 -1380 5616 -1378
rect 5374 -1392 5389 -1388
rect 5292 -1394 5389 -1392
rect 5417 -1394 5585 -1382
rect 5601 -1392 5616 -1388
rect 5634 -1391 5673 -1372
rect 5692 -1378 5699 -1377
rect 5698 -1385 5699 -1378
rect 5682 -1388 5683 -1385
rect 5698 -1388 5711 -1385
rect 5634 -1392 5664 -1391
rect 5673 -1392 5679 -1391
rect 5682 -1392 5711 -1388
rect 5601 -1393 5711 -1392
rect 5601 -1394 5717 -1393
rect 5276 -1402 5327 -1394
rect 5276 -1414 5301 -1402
rect 5308 -1414 5327 -1402
rect 5358 -1402 5408 -1394
rect 5358 -1410 5374 -1402
rect 5381 -1404 5408 -1402
rect 5417 -1404 5638 -1394
rect 5381 -1414 5638 -1404
rect 5667 -1402 5717 -1394
rect 5667 -1411 5683 -1402
rect 5276 -1422 5327 -1414
rect 5374 -1422 5638 -1414
rect 5664 -1414 5683 -1411
rect 5690 -1414 5717 -1402
rect 5664 -1422 5717 -1414
rect 5292 -1430 5293 -1422
rect 5308 -1430 5321 -1422
rect 5292 -1438 5308 -1430
rect 5289 -1445 5308 -1442
rect 5289 -1454 5311 -1445
rect 5262 -1464 5311 -1454
rect 5262 -1470 5292 -1464
rect 5311 -1469 5316 -1464
rect 5234 -1486 5308 -1470
rect 5326 -1478 5356 -1422
rect 5391 -1432 5599 -1422
rect 5634 -1426 5679 -1422
rect 5682 -1423 5683 -1422
rect 5698 -1423 5711 -1422
rect 5417 -1462 5606 -1432
rect 5432 -1465 5606 -1462
rect 5425 -1468 5606 -1465
rect 5234 -1488 5247 -1486
rect 5262 -1488 5296 -1486
rect 5234 -1504 5308 -1488
rect 5335 -1492 5348 -1478
rect 5363 -1492 5379 -1476
rect 5425 -1481 5436 -1468
rect 5218 -1526 5219 -1510
rect 5234 -1526 5247 -1504
rect 5262 -1526 5292 -1504
rect 5335 -1508 5397 -1492
rect 5425 -1499 5436 -1483
rect 5441 -1488 5451 -1468
rect 5461 -1488 5475 -1468
rect 5478 -1481 5487 -1468
rect 5503 -1481 5512 -1468
rect 5441 -1499 5475 -1488
rect 5478 -1499 5487 -1483
rect 5503 -1499 5512 -1483
rect 5519 -1488 5529 -1468
rect 5539 -1488 5553 -1468
rect 5554 -1481 5565 -1468
rect 5519 -1499 5553 -1488
rect 5554 -1499 5565 -1483
rect 5611 -1492 5627 -1476
rect 5634 -1478 5664 -1426
rect 5698 -1430 5699 -1423
rect 5683 -1438 5699 -1430
rect 5670 -1470 5683 -1451
rect 5698 -1470 5728 -1454
rect 5670 -1486 5744 -1470
rect 5670 -1488 5683 -1486
rect 5698 -1488 5732 -1486
rect 5335 -1510 5348 -1508
rect 5363 -1510 5397 -1508
rect 5335 -1526 5397 -1510
rect 5441 -1515 5457 -1508
rect 5519 -1515 5549 -1504
rect 5597 -1508 5643 -1492
rect 5670 -1504 5744 -1488
rect 5597 -1510 5631 -1508
rect 5596 -1526 5643 -1510
rect 5670 -1526 5683 -1504
rect 5698 -1526 5728 -1504
rect 5755 -1526 5756 -1510
rect 5771 -1526 5784 -1366
rect 5814 -1470 5827 -1366
rect 5872 -1388 5873 -1378
rect 5888 -1388 5901 -1378
rect 5872 -1392 5901 -1388
rect 5906 -1392 5936 -1366
rect 5954 -1380 5970 -1378
rect 6042 -1380 6093 -1366
rect 6043 -1382 6107 -1380
rect 6150 -1382 6165 -1366
rect 6214 -1369 6244 -1366
rect 6214 -1372 6250 -1369
rect 6180 -1380 6196 -1378
rect 5954 -1392 5969 -1388
rect 5872 -1394 5969 -1392
rect 5997 -1394 6165 -1382
rect 6181 -1392 6196 -1388
rect 6214 -1391 6253 -1372
rect 6272 -1378 6279 -1377
rect 6278 -1385 6279 -1378
rect 6262 -1388 6263 -1385
rect 6278 -1388 6291 -1385
rect 6214 -1392 6244 -1391
rect 6253 -1392 6259 -1391
rect 6262 -1392 6291 -1388
rect 6181 -1393 6291 -1392
rect 6181 -1394 6297 -1393
rect 5856 -1402 5907 -1394
rect 5856 -1414 5881 -1402
rect 5888 -1414 5907 -1402
rect 5938 -1402 5988 -1394
rect 5938 -1410 5954 -1402
rect 5961 -1404 5988 -1402
rect 5997 -1404 6218 -1394
rect 5961 -1414 6218 -1404
rect 6247 -1402 6297 -1394
rect 6247 -1411 6263 -1402
rect 5856 -1422 5907 -1414
rect 5954 -1422 6218 -1414
rect 6244 -1414 6263 -1411
rect 6270 -1414 6297 -1402
rect 6244 -1422 6297 -1414
rect 5872 -1430 5873 -1422
rect 5888 -1430 5901 -1422
rect 5872 -1438 5888 -1430
rect 5869 -1445 5888 -1442
rect 5869 -1454 5891 -1445
rect 5842 -1464 5891 -1454
rect 5842 -1470 5872 -1464
rect 5891 -1469 5896 -1464
rect 5814 -1486 5888 -1470
rect 5906 -1478 5936 -1422
rect 5971 -1432 6179 -1422
rect 6214 -1426 6259 -1422
rect 6262 -1423 6263 -1422
rect 6278 -1423 6291 -1422
rect 5997 -1462 6186 -1432
rect 6012 -1465 6186 -1462
rect 6005 -1468 6186 -1465
rect 5814 -1488 5827 -1486
rect 5842 -1488 5876 -1486
rect 5814 -1504 5888 -1488
rect 5915 -1492 5928 -1478
rect 5943 -1492 5959 -1476
rect 6005 -1481 6016 -1468
rect 5798 -1526 5799 -1510
rect 5814 -1526 5827 -1504
rect 5842 -1526 5872 -1504
rect 5915 -1508 5977 -1492
rect 6005 -1499 6016 -1483
rect 6021 -1488 6031 -1468
rect 6041 -1488 6055 -1468
rect 6058 -1481 6067 -1468
rect 6083 -1481 6092 -1468
rect 6021 -1499 6055 -1488
rect 6058 -1499 6067 -1483
rect 6083 -1499 6092 -1483
rect 6099 -1488 6109 -1468
rect 6119 -1488 6133 -1468
rect 6134 -1481 6145 -1468
rect 6099 -1499 6133 -1488
rect 6134 -1499 6145 -1483
rect 6191 -1492 6207 -1476
rect 6214 -1478 6244 -1426
rect 6278 -1430 6279 -1423
rect 6263 -1438 6279 -1430
rect 6250 -1470 6263 -1451
rect 6278 -1470 6308 -1454
rect 6250 -1486 6324 -1470
rect 6250 -1488 6263 -1486
rect 6278 -1488 6312 -1486
rect 5915 -1510 5928 -1508
rect 5943 -1510 5977 -1508
rect 5915 -1526 5977 -1510
rect 6021 -1515 6037 -1508
rect 6099 -1515 6129 -1504
rect 6177 -1508 6223 -1492
rect 6250 -1504 6324 -1488
rect 6177 -1510 6211 -1508
rect 6176 -1526 6223 -1510
rect 6250 -1526 6263 -1504
rect 6278 -1526 6308 -1504
rect 6335 -1526 6336 -1510
rect 6351 -1526 6364 -1366
rect 6394 -1470 6407 -1366
rect 6452 -1388 6453 -1378
rect 6468 -1388 6481 -1378
rect 6452 -1392 6481 -1388
rect 6486 -1392 6516 -1366
rect 6534 -1380 6550 -1378
rect 6622 -1380 6673 -1366
rect 6623 -1382 6687 -1380
rect 6730 -1382 6745 -1366
rect 6794 -1369 6824 -1366
rect 6794 -1372 6830 -1369
rect 6760 -1380 6776 -1378
rect 6534 -1392 6549 -1388
rect 6452 -1394 6549 -1392
rect 6577 -1394 6745 -1382
rect 6761 -1392 6776 -1388
rect 6794 -1391 6833 -1372
rect 6852 -1378 6859 -1377
rect 6858 -1385 6859 -1378
rect 6842 -1388 6843 -1385
rect 6858 -1388 6871 -1385
rect 6794 -1392 6824 -1391
rect 6833 -1392 6839 -1391
rect 6842 -1392 6871 -1388
rect 6761 -1393 6871 -1392
rect 6761 -1394 6877 -1393
rect 6436 -1402 6487 -1394
rect 6436 -1414 6461 -1402
rect 6468 -1414 6487 -1402
rect 6518 -1402 6568 -1394
rect 6518 -1410 6534 -1402
rect 6541 -1404 6568 -1402
rect 6577 -1404 6798 -1394
rect 6541 -1414 6798 -1404
rect 6827 -1402 6877 -1394
rect 6827 -1411 6843 -1402
rect 6436 -1422 6487 -1414
rect 6534 -1422 6798 -1414
rect 6824 -1414 6843 -1411
rect 6850 -1414 6877 -1402
rect 6824 -1422 6877 -1414
rect 6452 -1430 6453 -1422
rect 6468 -1430 6481 -1422
rect 6452 -1438 6468 -1430
rect 6449 -1445 6468 -1442
rect 6449 -1454 6471 -1445
rect 6422 -1464 6471 -1454
rect 6422 -1470 6452 -1464
rect 6471 -1469 6476 -1464
rect 6394 -1486 6468 -1470
rect 6486 -1478 6516 -1422
rect 6551 -1432 6759 -1422
rect 6794 -1426 6839 -1422
rect 6842 -1423 6843 -1422
rect 6858 -1423 6871 -1422
rect 6577 -1462 6766 -1432
rect 6592 -1465 6766 -1462
rect 6585 -1468 6766 -1465
rect 6394 -1488 6407 -1486
rect 6422 -1488 6456 -1486
rect 6394 -1504 6468 -1488
rect 6495 -1492 6508 -1478
rect 6523 -1492 6539 -1476
rect 6585 -1481 6596 -1468
rect 6378 -1526 6379 -1510
rect 6394 -1526 6407 -1504
rect 6422 -1526 6452 -1504
rect 6495 -1508 6557 -1492
rect 6585 -1499 6596 -1483
rect 6601 -1488 6611 -1468
rect 6621 -1488 6635 -1468
rect 6638 -1481 6647 -1468
rect 6663 -1481 6672 -1468
rect 6601 -1499 6635 -1488
rect 6638 -1499 6647 -1483
rect 6663 -1499 6672 -1483
rect 6679 -1488 6689 -1468
rect 6699 -1488 6713 -1468
rect 6714 -1481 6725 -1468
rect 6679 -1499 6713 -1488
rect 6714 -1499 6725 -1483
rect 6771 -1492 6787 -1476
rect 6794 -1478 6824 -1426
rect 6858 -1430 6859 -1423
rect 6843 -1438 6859 -1430
rect 6830 -1470 6843 -1451
rect 6858 -1470 6888 -1454
rect 6830 -1486 6904 -1470
rect 6830 -1488 6843 -1486
rect 6858 -1488 6892 -1486
rect 6495 -1510 6508 -1508
rect 6523 -1510 6557 -1508
rect 6495 -1526 6557 -1510
rect 6601 -1515 6617 -1508
rect 6679 -1515 6709 -1504
rect 6757 -1508 6803 -1492
rect 6830 -1504 6904 -1488
rect 6757 -1510 6791 -1508
rect 6756 -1526 6803 -1510
rect 6830 -1526 6843 -1504
rect 6858 -1526 6888 -1504
rect 6915 -1526 6916 -1510
rect 6931 -1526 6944 -1366
rect -8 -1534 33 -1526
rect -8 -1560 7 -1534
rect 14 -1560 33 -1534
rect 97 -1538 159 -1526
rect 171 -1538 246 -1526
rect 304 -1538 379 -1526
rect 391 -1538 422 -1526
rect 428 -1538 463 -1526
rect 97 -1540 259 -1538
rect -8 -1568 33 -1560
rect 115 -1564 128 -1540
rect 143 -1542 158 -1540
rect -2 -1578 -1 -1568
rect 14 -1578 27 -1568
rect 42 -1578 72 -1564
rect 115 -1578 158 -1564
rect 182 -1567 189 -1560
rect 192 -1564 259 -1540
rect 291 -1540 463 -1538
rect 261 -1562 289 -1558
rect 291 -1562 371 -1540
rect 392 -1542 407 -1540
rect 261 -1564 371 -1562
rect 192 -1568 371 -1564
rect 165 -1578 195 -1568
rect 197 -1578 350 -1568
rect 358 -1578 388 -1568
rect 392 -1578 422 -1564
rect 450 -1578 463 -1540
rect 535 -1534 570 -1526
rect 535 -1560 536 -1534
rect 543 -1560 570 -1534
rect 478 -1578 508 -1564
rect 535 -1568 570 -1560
rect 572 -1534 613 -1526
rect 572 -1560 587 -1534
rect 594 -1560 613 -1534
rect 677 -1538 739 -1526
rect 751 -1538 826 -1526
rect 884 -1538 959 -1526
rect 971 -1538 1002 -1526
rect 1008 -1538 1043 -1526
rect 677 -1540 839 -1538
rect 572 -1568 613 -1560
rect 695 -1564 708 -1540
rect 723 -1542 738 -1540
rect 535 -1578 536 -1568
rect 551 -1578 564 -1568
rect 578 -1578 579 -1568
rect 594 -1578 607 -1568
rect 622 -1578 652 -1564
rect 695 -1578 738 -1564
rect 762 -1567 769 -1560
rect 772 -1564 839 -1540
rect 871 -1540 1043 -1538
rect 841 -1562 869 -1558
rect 871 -1562 951 -1540
rect 972 -1542 987 -1540
rect 841 -1564 951 -1562
rect 772 -1568 951 -1564
rect 745 -1578 775 -1568
rect 777 -1578 930 -1568
rect 938 -1578 968 -1568
rect 972 -1578 1002 -1564
rect 1030 -1578 1043 -1540
rect 1115 -1534 1150 -1526
rect 1115 -1560 1116 -1534
rect 1123 -1560 1150 -1534
rect 1058 -1578 1088 -1564
rect 1115 -1568 1150 -1560
rect 1152 -1534 1193 -1526
rect 1152 -1560 1167 -1534
rect 1174 -1560 1193 -1534
rect 1257 -1538 1319 -1526
rect 1331 -1538 1406 -1526
rect 1464 -1538 1539 -1526
rect 3435 -1534 3470 -1526
rect 1257 -1540 1419 -1538
rect 1152 -1568 1193 -1560
rect 1275 -1564 1288 -1540
rect 1303 -1542 1318 -1540
rect 1115 -1578 1116 -1568
rect 1131 -1578 1144 -1568
rect 1158 -1578 1159 -1568
rect 1174 -1578 1187 -1568
rect 1202 -1578 1232 -1564
rect 1275 -1578 1318 -1564
rect 1342 -1567 1349 -1560
rect 1352 -1564 1419 -1540
rect 1451 -1540 1551 -1538
rect 1421 -1562 1449 -1558
rect 1451 -1562 1531 -1540
rect 1421 -1564 1531 -1562
rect 3435 -1560 3436 -1534
rect 3443 -1560 3470 -1534
rect 1352 -1568 1531 -1564
rect 1325 -1578 1355 -1568
rect 1357 -1578 1510 -1568
rect 1518 -1578 1548 -1568
rect 3379 -1578 3408 -1564
rect 3435 -1568 3470 -1560
rect 3472 -1534 3513 -1526
rect 3472 -1560 3487 -1534
rect 3494 -1560 3513 -1534
rect 3577 -1538 3639 -1526
rect 3651 -1538 3726 -1526
rect 3784 -1538 3859 -1526
rect 3871 -1538 3902 -1526
rect 3908 -1538 3943 -1526
rect 3577 -1540 3739 -1538
rect 3472 -1568 3513 -1560
rect 3595 -1564 3608 -1540
rect 3623 -1542 3638 -1540
rect 3435 -1578 3436 -1568
rect 3451 -1578 3464 -1568
rect 3478 -1578 3479 -1568
rect 3494 -1578 3507 -1568
rect 3522 -1578 3552 -1564
rect 3595 -1578 3638 -1564
rect 3662 -1567 3669 -1560
rect 3672 -1564 3739 -1540
rect 3771 -1540 3943 -1538
rect 3741 -1562 3769 -1558
rect 3771 -1562 3851 -1540
rect 3872 -1542 3887 -1540
rect 3741 -1564 3851 -1562
rect 3672 -1568 3851 -1564
rect 3645 -1578 3675 -1568
rect 3677 -1578 3830 -1568
rect 3838 -1578 3868 -1568
rect 3872 -1578 3902 -1564
rect 3930 -1578 3943 -1540
rect 4015 -1534 4050 -1526
rect 4015 -1560 4016 -1534
rect 4023 -1560 4050 -1534
rect 3958 -1578 3988 -1564
rect 4015 -1568 4050 -1560
rect 4052 -1534 4093 -1526
rect 4052 -1560 4067 -1534
rect 4074 -1560 4093 -1534
rect 4157 -1538 4219 -1526
rect 4231 -1538 4306 -1526
rect 4364 -1538 4439 -1526
rect 4451 -1538 4482 -1526
rect 4488 -1538 4523 -1526
rect 4157 -1540 4319 -1538
rect 4052 -1568 4093 -1560
rect 4175 -1564 4188 -1540
rect 4203 -1542 4218 -1540
rect 4015 -1578 4016 -1568
rect 4031 -1578 4044 -1568
rect 4058 -1578 4059 -1568
rect 4074 -1578 4087 -1568
rect 4102 -1578 4132 -1564
rect 4175 -1578 4218 -1564
rect 4242 -1567 4249 -1560
rect 4252 -1564 4319 -1540
rect 4351 -1540 4523 -1538
rect 4321 -1562 4349 -1558
rect 4351 -1562 4431 -1540
rect 4452 -1542 4467 -1540
rect 4321 -1564 4431 -1562
rect 4252 -1568 4431 -1564
rect 4225 -1578 4255 -1568
rect 4257 -1578 4410 -1568
rect 4418 -1578 4448 -1568
rect 4452 -1578 4482 -1564
rect 4510 -1578 4523 -1540
rect 4595 -1534 4630 -1526
rect 4595 -1560 4596 -1534
rect 4603 -1560 4630 -1534
rect 4538 -1578 4568 -1564
rect 4595 -1568 4630 -1560
rect 4632 -1534 4673 -1526
rect 4632 -1560 4647 -1534
rect 4654 -1560 4673 -1534
rect 4737 -1538 4799 -1526
rect 4811 -1538 4886 -1526
rect 4944 -1538 5019 -1526
rect 5031 -1538 5062 -1526
rect 5068 -1538 5103 -1526
rect 4737 -1540 4899 -1538
rect 4755 -1558 4768 -1540
rect 4783 -1542 4798 -1540
rect 4632 -1568 4673 -1560
rect 4756 -1564 4768 -1558
rect 4832 -1558 4899 -1540
rect 4931 -1540 5103 -1538
rect 4931 -1558 5011 -1540
rect 5032 -1542 5047 -1540
rect 4595 -1578 4596 -1568
rect 4611 -1578 4624 -1568
rect 4638 -1578 4639 -1568
rect 4654 -1578 4667 -1568
rect 4682 -1578 4712 -1564
rect 4756 -1578 4798 -1564
rect 4822 -1567 4829 -1560
rect 4832 -1568 5011 -1558
rect 4805 -1578 4835 -1568
rect 4837 -1578 4990 -1568
rect 4998 -1578 5028 -1568
rect 5032 -1578 5062 -1564
rect 5090 -1578 5103 -1540
rect 5175 -1534 5210 -1526
rect 5175 -1560 5176 -1534
rect 5183 -1560 5210 -1534
rect 5118 -1578 5148 -1564
rect 5175 -1568 5210 -1560
rect 5212 -1534 5253 -1526
rect 5212 -1560 5227 -1534
rect 5234 -1560 5253 -1534
rect 5317 -1538 5379 -1526
rect 5391 -1538 5466 -1526
rect 5524 -1538 5599 -1526
rect 5611 -1538 5642 -1526
rect 5648 -1538 5683 -1526
rect 5317 -1540 5479 -1538
rect 5335 -1558 5348 -1540
rect 5363 -1542 5378 -1540
rect 5212 -1568 5253 -1560
rect 5336 -1564 5348 -1558
rect 5412 -1558 5479 -1540
rect 5511 -1540 5683 -1538
rect 5511 -1558 5591 -1540
rect 5612 -1542 5627 -1540
rect 5175 -1578 5176 -1568
rect 5191 -1578 5204 -1568
rect 5218 -1578 5219 -1568
rect 5234 -1578 5247 -1568
rect 5262 -1578 5292 -1564
rect 5336 -1578 5378 -1564
rect 5402 -1567 5409 -1560
rect 5412 -1568 5591 -1558
rect 5385 -1578 5415 -1568
rect 5417 -1578 5570 -1568
rect 5578 -1578 5608 -1568
rect 5612 -1578 5642 -1564
rect 5670 -1578 5683 -1540
rect 5755 -1534 5790 -1526
rect 5755 -1560 5756 -1534
rect 5763 -1560 5790 -1534
rect 5698 -1578 5728 -1564
rect 5755 -1568 5790 -1560
rect 5792 -1534 5833 -1526
rect 5792 -1560 5807 -1534
rect 5814 -1560 5833 -1534
rect 5897 -1538 5959 -1526
rect 5971 -1538 6046 -1526
rect 6104 -1538 6179 -1526
rect 6191 -1538 6222 -1526
rect 6228 -1538 6263 -1526
rect 5897 -1540 6059 -1538
rect 5915 -1558 5928 -1540
rect 5943 -1542 5958 -1540
rect 5792 -1568 5833 -1560
rect 5916 -1564 5928 -1558
rect 5992 -1558 6059 -1540
rect 6091 -1540 6263 -1538
rect 6091 -1558 6171 -1540
rect 6192 -1542 6207 -1540
rect 5755 -1578 5756 -1568
rect 5771 -1578 5784 -1568
rect 5798 -1578 5799 -1568
rect 5814 -1578 5827 -1568
rect 5842 -1578 5872 -1564
rect 5916 -1578 5958 -1564
rect 5982 -1567 5989 -1560
rect 5992 -1568 6171 -1558
rect 5965 -1578 5995 -1568
rect 5997 -1578 6150 -1568
rect 6158 -1578 6188 -1568
rect 6192 -1578 6222 -1564
rect 6250 -1578 6263 -1540
rect 6335 -1534 6370 -1526
rect 6335 -1560 6336 -1534
rect 6343 -1560 6370 -1534
rect 6278 -1578 6308 -1564
rect 6335 -1568 6370 -1560
rect 6372 -1534 6413 -1526
rect 6372 -1560 6387 -1534
rect 6394 -1560 6413 -1534
rect 6477 -1538 6539 -1526
rect 6551 -1538 6626 -1526
rect 6684 -1538 6759 -1526
rect 6771 -1538 6802 -1526
rect 6808 -1538 6843 -1526
rect 6477 -1540 6639 -1538
rect 6495 -1558 6508 -1540
rect 6523 -1542 6538 -1540
rect 6372 -1568 6413 -1560
rect 6496 -1564 6508 -1558
rect 6572 -1558 6639 -1540
rect 6671 -1540 6843 -1538
rect 6671 -1558 6751 -1540
rect 6772 -1542 6787 -1540
rect 6335 -1578 6336 -1568
rect 6351 -1578 6364 -1568
rect 6378 -1578 6379 -1568
rect 6394 -1578 6407 -1568
rect 6422 -1578 6452 -1564
rect 6496 -1578 6538 -1564
rect 6562 -1567 6569 -1560
rect 6572 -1568 6751 -1558
rect 6545 -1578 6575 -1568
rect 6577 -1578 6730 -1568
rect 6738 -1578 6768 -1568
rect 6772 -1578 6802 -1564
rect 6830 -1578 6843 -1540
rect 6915 -1534 6950 -1526
rect 6915 -1560 6916 -1534
rect 6923 -1560 6950 -1534
rect 6858 -1578 6888 -1564
rect 6915 -1568 6950 -1560
rect 6915 -1578 6916 -1568
rect 6931 -1578 6944 -1568
rect -2 -1584 1551 -1578
rect -1 -1592 1551 -1584
rect 3379 -1592 6944 -1578
rect 14 -1622 27 -1592
rect 42 -1610 72 -1592
rect 115 -1606 129 -1592
rect 165 -1606 385 -1592
rect 116 -1608 129 -1606
rect 82 -1620 97 -1608
rect 79 -1622 101 -1620
rect 106 -1622 136 -1608
rect 197 -1610 350 -1606
rect 179 -1622 371 -1610
rect 414 -1622 444 -1608
rect 450 -1622 463 -1592
rect 478 -1610 508 -1592
rect 551 -1622 564 -1592
rect 594 -1622 607 -1592
rect 622 -1610 652 -1592
rect 695 -1606 709 -1592
rect 745 -1606 965 -1592
rect 696 -1608 709 -1606
rect 662 -1620 677 -1608
rect 659 -1622 681 -1620
rect 686 -1622 716 -1608
rect 777 -1610 930 -1606
rect 759 -1622 951 -1610
rect 994 -1622 1024 -1608
rect 1030 -1622 1043 -1592
rect 1058 -1610 1088 -1592
rect 1131 -1622 1144 -1592
rect 1174 -1622 1187 -1592
rect 1202 -1610 1232 -1592
rect 1275 -1606 1289 -1592
rect 1325 -1606 1545 -1592
rect 1276 -1608 1289 -1606
rect 1242 -1620 1257 -1608
rect 1239 -1622 1261 -1620
rect 1266 -1622 1296 -1608
rect 1357 -1610 1510 -1606
rect 3379 -1610 3408 -1592
rect 1339 -1622 1531 -1610
rect 3451 -1622 3464 -1592
rect 3494 -1622 3507 -1592
rect 3522 -1610 3552 -1592
rect 3595 -1606 3609 -1592
rect 3645 -1606 3865 -1592
rect 3596 -1608 3609 -1606
rect 3562 -1620 3577 -1608
rect 3559 -1622 3581 -1620
rect 3586 -1622 3616 -1608
rect 3677 -1610 3830 -1606
rect 3659 -1622 3851 -1610
rect 3894 -1622 3924 -1608
rect 3930 -1622 3943 -1592
rect 3958 -1610 3988 -1592
rect 4031 -1622 4044 -1592
rect 4074 -1622 4087 -1592
rect 4102 -1610 4132 -1592
rect 4175 -1606 4189 -1592
rect 4225 -1606 4445 -1592
rect 4176 -1608 4189 -1606
rect 4142 -1620 4157 -1608
rect 4139 -1622 4161 -1620
rect 4166 -1622 4196 -1608
rect 4257 -1610 4410 -1606
rect 4239 -1622 4431 -1610
rect 4474 -1622 4504 -1608
rect 4510 -1622 4523 -1592
rect 4538 -1610 4568 -1592
rect 4611 -1622 4624 -1592
rect 4654 -1622 4667 -1592
rect 4682 -1610 4712 -1592
rect 4756 -1608 4769 -1592
rect 4805 -1606 5025 -1592
rect 4722 -1620 4737 -1608
rect 4719 -1622 4741 -1620
rect 4746 -1622 4776 -1608
rect 4837 -1610 4990 -1606
rect 4819 -1622 5011 -1610
rect 5054 -1622 5084 -1608
rect 5090 -1622 5103 -1592
rect 5118 -1610 5148 -1592
rect 5191 -1622 5204 -1592
rect 5234 -1622 5247 -1592
rect 5262 -1610 5292 -1592
rect 5336 -1608 5349 -1592
rect 5385 -1606 5605 -1592
rect 5302 -1620 5317 -1608
rect 5299 -1622 5321 -1620
rect 5326 -1622 5356 -1608
rect 5417 -1610 5570 -1606
rect 5399 -1622 5591 -1610
rect 5634 -1622 5664 -1608
rect 5670 -1622 5683 -1592
rect 5698 -1610 5728 -1592
rect 5771 -1622 5784 -1592
rect 5814 -1622 5827 -1592
rect 5842 -1610 5872 -1592
rect 5916 -1608 5929 -1592
rect 5965 -1606 6185 -1592
rect 5882 -1620 5897 -1608
rect 5879 -1622 5901 -1620
rect 5906 -1622 5936 -1608
rect 5997 -1610 6150 -1606
rect 5979 -1622 6171 -1610
rect 6214 -1622 6244 -1608
rect 6250 -1622 6263 -1592
rect 6278 -1610 6308 -1592
rect 6351 -1622 6364 -1592
rect 6394 -1622 6407 -1592
rect 6422 -1610 6452 -1592
rect 6496 -1608 6509 -1592
rect 6545 -1606 6765 -1592
rect 6462 -1620 6477 -1608
rect 6459 -1622 6481 -1620
rect 6486 -1622 6516 -1608
rect 6577 -1610 6730 -1606
rect 6559 -1622 6751 -1610
rect 6794 -1622 6824 -1608
rect 6830 -1622 6843 -1592
rect 6858 -1610 6888 -1592
rect 6931 -1622 6944 -1592
rect -1 -1636 1551 -1622
rect 3379 -1636 6944 -1622
rect 14 -1740 27 -1636
rect 72 -1658 73 -1648
rect 88 -1658 101 -1648
rect 72 -1662 101 -1658
rect 106 -1662 136 -1636
rect 154 -1650 170 -1648
rect 242 -1650 295 -1636
rect 243 -1652 307 -1650
rect 350 -1652 365 -1636
rect 414 -1639 444 -1636
rect 414 -1642 450 -1639
rect 380 -1650 396 -1648
rect 154 -1662 169 -1658
rect 72 -1664 169 -1662
rect 197 -1664 365 -1652
rect 381 -1662 396 -1658
rect 414 -1661 453 -1642
rect 472 -1648 479 -1647
rect 478 -1655 479 -1648
rect 462 -1658 463 -1655
rect 478 -1658 491 -1655
rect 414 -1662 444 -1661
rect 453 -1662 459 -1661
rect 462 -1662 491 -1658
rect 381 -1663 491 -1662
rect 381 -1664 497 -1663
rect 56 -1672 107 -1664
rect 56 -1684 81 -1672
rect 88 -1684 107 -1672
rect 138 -1672 188 -1664
rect 138 -1680 154 -1672
rect 161 -1674 188 -1672
rect 197 -1674 418 -1664
rect 161 -1684 418 -1674
rect 447 -1672 497 -1664
rect 447 -1681 463 -1672
rect 56 -1692 107 -1684
rect 154 -1692 418 -1684
rect 444 -1684 463 -1681
rect 470 -1684 497 -1672
rect 444 -1692 497 -1684
rect 72 -1700 73 -1692
rect 88 -1700 101 -1692
rect 72 -1708 88 -1700
rect 69 -1715 88 -1712
rect 69 -1724 91 -1715
rect 42 -1734 91 -1724
rect 42 -1740 72 -1734
rect 91 -1739 96 -1734
rect 14 -1756 88 -1740
rect 106 -1748 136 -1692
rect 171 -1702 379 -1692
rect 414 -1696 459 -1692
rect 462 -1693 463 -1692
rect 478 -1693 491 -1692
rect 197 -1732 386 -1702
rect 212 -1735 386 -1732
rect 205 -1738 386 -1735
rect 14 -1758 27 -1756
rect 42 -1758 76 -1756
rect 14 -1774 88 -1758
rect 115 -1762 128 -1748
rect 143 -1762 159 -1746
rect 205 -1751 216 -1738
rect -2 -1796 -1 -1780
rect 14 -1796 27 -1774
rect 42 -1796 72 -1774
rect 115 -1778 177 -1762
rect 205 -1769 216 -1753
rect 221 -1758 231 -1738
rect 241 -1758 255 -1738
rect 258 -1751 267 -1738
rect 283 -1751 292 -1738
rect 221 -1769 255 -1758
rect 258 -1769 267 -1753
rect 283 -1769 292 -1753
rect 299 -1758 309 -1738
rect 319 -1758 333 -1738
rect 334 -1751 345 -1738
rect 299 -1769 333 -1758
rect 334 -1769 345 -1753
rect 391 -1762 407 -1746
rect 414 -1748 444 -1696
rect 478 -1700 479 -1693
rect 463 -1708 479 -1700
rect 450 -1740 463 -1721
rect 478 -1740 508 -1724
rect 450 -1756 524 -1740
rect 450 -1758 463 -1756
rect 478 -1758 512 -1756
rect 115 -1780 128 -1778
rect 143 -1780 177 -1778
rect 115 -1796 177 -1780
rect 221 -1785 237 -1778
rect 299 -1785 329 -1774
rect 377 -1778 423 -1762
rect 450 -1774 524 -1758
rect 377 -1780 411 -1778
rect 376 -1796 423 -1780
rect 450 -1796 463 -1774
rect 478 -1796 508 -1774
rect 535 -1796 536 -1780
rect 551 -1796 564 -1636
rect 594 -1740 607 -1636
rect 652 -1658 653 -1648
rect 668 -1658 681 -1648
rect 652 -1662 681 -1658
rect 686 -1662 716 -1636
rect 734 -1650 750 -1648
rect 822 -1650 875 -1636
rect 823 -1652 887 -1650
rect 930 -1652 945 -1636
rect 994 -1639 1024 -1636
rect 994 -1642 1030 -1639
rect 960 -1650 976 -1648
rect 734 -1662 749 -1658
rect 652 -1664 749 -1662
rect 777 -1664 945 -1652
rect 961 -1662 976 -1658
rect 994 -1661 1033 -1642
rect 1052 -1648 1059 -1647
rect 1058 -1655 1059 -1648
rect 1042 -1658 1043 -1655
rect 1058 -1658 1071 -1655
rect 994 -1662 1024 -1661
rect 1033 -1662 1039 -1661
rect 1042 -1662 1071 -1658
rect 961 -1663 1071 -1662
rect 961 -1664 1077 -1663
rect 636 -1672 687 -1664
rect 636 -1684 661 -1672
rect 668 -1684 687 -1672
rect 718 -1672 768 -1664
rect 718 -1680 734 -1672
rect 741 -1674 768 -1672
rect 777 -1674 998 -1664
rect 741 -1684 998 -1674
rect 1027 -1672 1077 -1664
rect 1027 -1681 1043 -1672
rect 636 -1692 687 -1684
rect 734 -1692 998 -1684
rect 1024 -1684 1043 -1681
rect 1050 -1684 1077 -1672
rect 1024 -1692 1077 -1684
rect 652 -1700 653 -1692
rect 668 -1700 681 -1692
rect 652 -1708 668 -1700
rect 649 -1715 668 -1712
rect 649 -1724 671 -1715
rect 622 -1734 671 -1724
rect 622 -1740 652 -1734
rect 671 -1739 676 -1734
rect 594 -1756 668 -1740
rect 686 -1748 716 -1692
rect 751 -1702 959 -1692
rect 994 -1696 1039 -1692
rect 1042 -1693 1043 -1692
rect 1058 -1693 1071 -1692
rect 777 -1732 966 -1702
rect 792 -1735 966 -1732
rect 785 -1738 966 -1735
rect 594 -1758 607 -1756
rect 622 -1758 656 -1756
rect 594 -1774 668 -1758
rect 695 -1762 708 -1748
rect 723 -1762 739 -1746
rect 785 -1751 796 -1738
rect 578 -1796 579 -1780
rect 594 -1796 607 -1774
rect 622 -1796 652 -1774
rect 695 -1778 757 -1762
rect 785 -1769 796 -1753
rect 801 -1758 811 -1738
rect 821 -1758 835 -1738
rect 838 -1751 847 -1738
rect 863 -1751 872 -1738
rect 801 -1769 835 -1758
rect 838 -1769 847 -1753
rect 863 -1769 872 -1753
rect 879 -1758 889 -1738
rect 899 -1758 913 -1738
rect 914 -1751 925 -1738
rect 879 -1769 913 -1758
rect 914 -1769 925 -1753
rect 971 -1762 987 -1746
rect 994 -1748 1024 -1696
rect 1058 -1700 1059 -1693
rect 1043 -1708 1059 -1700
rect 1030 -1740 1043 -1721
rect 1058 -1740 1088 -1724
rect 1030 -1756 1104 -1740
rect 1030 -1758 1043 -1756
rect 1058 -1758 1092 -1756
rect 695 -1780 708 -1778
rect 723 -1780 757 -1778
rect 695 -1796 757 -1780
rect 801 -1785 817 -1778
rect 879 -1785 909 -1774
rect 957 -1778 1003 -1762
rect 1030 -1774 1104 -1758
rect 957 -1780 991 -1778
rect 956 -1796 1003 -1780
rect 1030 -1796 1043 -1774
rect 1058 -1796 1088 -1774
rect 1115 -1796 1116 -1780
rect 1131 -1796 1144 -1636
rect 1174 -1740 1187 -1636
rect 1232 -1658 1233 -1648
rect 1248 -1658 1261 -1648
rect 1232 -1662 1261 -1658
rect 1266 -1662 1296 -1636
rect 1314 -1650 1330 -1648
rect 1402 -1650 1455 -1636
rect 1403 -1652 1467 -1650
rect 1510 -1652 1525 -1636
rect 1540 -1650 1551 -1648
rect 1314 -1662 1329 -1658
rect 1232 -1664 1329 -1662
rect 1357 -1664 1525 -1652
rect 1541 -1664 1551 -1658
rect 1216 -1672 1267 -1664
rect 1216 -1684 1241 -1672
rect 1248 -1684 1267 -1672
rect 1298 -1672 1348 -1664
rect 1298 -1680 1314 -1672
rect 1321 -1674 1348 -1672
rect 1357 -1674 1551 -1664
rect 1321 -1684 1551 -1674
rect 1216 -1692 1267 -1684
rect 1314 -1692 1551 -1684
rect 3379 -1663 3391 -1655
rect 3379 -1692 3397 -1663
rect 1232 -1700 1233 -1692
rect 1248 -1700 1261 -1692
rect 1232 -1708 1248 -1700
rect 1229 -1715 1248 -1712
rect 1229 -1724 1251 -1715
rect 1202 -1734 1251 -1724
rect 1202 -1740 1232 -1734
rect 1251 -1739 1256 -1734
rect 1174 -1756 1248 -1740
rect 1266 -1748 1296 -1692
rect 1331 -1702 1539 -1692
rect 3379 -1693 3391 -1692
rect 1357 -1732 1546 -1702
rect 1372 -1735 1546 -1732
rect 1365 -1738 1546 -1735
rect 1174 -1758 1187 -1756
rect 1202 -1758 1236 -1756
rect 1174 -1774 1248 -1758
rect 1275 -1762 1288 -1748
rect 1303 -1762 1319 -1746
rect 1365 -1751 1376 -1738
rect 1158 -1796 1159 -1780
rect 1174 -1796 1187 -1774
rect 1202 -1796 1232 -1774
rect 1275 -1778 1337 -1762
rect 1365 -1769 1376 -1753
rect 1381 -1758 1391 -1738
rect 1401 -1758 1415 -1738
rect 1418 -1751 1427 -1738
rect 1443 -1751 1452 -1738
rect 1381 -1769 1415 -1758
rect 1418 -1769 1427 -1753
rect 1443 -1769 1452 -1753
rect 1459 -1758 1469 -1738
rect 1479 -1758 1493 -1738
rect 1494 -1751 1505 -1738
rect 3379 -1740 3408 -1724
rect 1459 -1769 1493 -1758
rect 1494 -1769 1505 -1753
rect 3379 -1756 3424 -1740
rect 3379 -1758 3412 -1756
rect 1275 -1780 1288 -1778
rect 1303 -1780 1337 -1778
rect 1275 -1796 1337 -1780
rect 1381 -1785 1397 -1778
rect 1459 -1785 1489 -1774
rect 1537 -1780 1551 -1762
rect 1536 -1796 1551 -1780
rect 3379 -1774 3424 -1758
rect 3379 -1796 3408 -1774
rect 3435 -1796 3436 -1780
rect 3451 -1796 3464 -1636
rect 3494 -1740 3507 -1636
rect 3552 -1658 3553 -1648
rect 3568 -1658 3581 -1648
rect 3552 -1662 3581 -1658
rect 3586 -1662 3616 -1636
rect 3634 -1650 3650 -1648
rect 3722 -1650 3775 -1636
rect 3723 -1652 3787 -1650
rect 3830 -1652 3845 -1636
rect 3894 -1639 3924 -1636
rect 3894 -1642 3930 -1639
rect 3860 -1650 3876 -1648
rect 3634 -1662 3649 -1658
rect 3552 -1664 3649 -1662
rect 3677 -1664 3845 -1652
rect 3861 -1662 3876 -1658
rect 3894 -1661 3933 -1642
rect 3952 -1648 3959 -1647
rect 3958 -1655 3959 -1648
rect 3942 -1658 3943 -1655
rect 3958 -1658 3971 -1655
rect 3894 -1662 3924 -1661
rect 3933 -1662 3939 -1661
rect 3942 -1662 3971 -1658
rect 3861 -1663 3971 -1662
rect 3861 -1664 3977 -1663
rect 3536 -1672 3587 -1664
rect 3536 -1684 3561 -1672
rect 3568 -1684 3587 -1672
rect 3618 -1672 3668 -1664
rect 3618 -1680 3634 -1672
rect 3641 -1674 3668 -1672
rect 3677 -1674 3898 -1664
rect 3641 -1684 3898 -1674
rect 3927 -1672 3977 -1664
rect 3927 -1681 3943 -1672
rect 3536 -1692 3587 -1684
rect 3634 -1692 3898 -1684
rect 3924 -1684 3943 -1681
rect 3950 -1684 3977 -1672
rect 3924 -1692 3977 -1684
rect 3552 -1700 3553 -1692
rect 3568 -1700 3581 -1692
rect 3552 -1708 3568 -1700
rect 3549 -1715 3568 -1712
rect 3549 -1724 3571 -1715
rect 3522 -1734 3571 -1724
rect 3522 -1740 3552 -1734
rect 3571 -1739 3576 -1734
rect 3494 -1756 3568 -1740
rect 3586 -1748 3616 -1692
rect 3651 -1702 3859 -1692
rect 3894 -1696 3939 -1692
rect 3942 -1693 3943 -1692
rect 3958 -1693 3971 -1692
rect 3677 -1732 3866 -1702
rect 3692 -1735 3866 -1732
rect 3685 -1738 3866 -1735
rect 3494 -1758 3507 -1756
rect 3522 -1758 3556 -1756
rect 3494 -1774 3568 -1758
rect 3595 -1762 3608 -1748
rect 3623 -1762 3639 -1746
rect 3685 -1751 3696 -1738
rect 3478 -1796 3479 -1780
rect 3494 -1796 3507 -1774
rect 3522 -1796 3552 -1774
rect 3595 -1778 3657 -1762
rect 3685 -1769 3696 -1753
rect 3701 -1758 3711 -1738
rect 3721 -1758 3735 -1738
rect 3738 -1751 3747 -1738
rect 3763 -1751 3772 -1738
rect 3701 -1769 3735 -1758
rect 3738 -1769 3747 -1753
rect 3763 -1769 3772 -1753
rect 3779 -1758 3789 -1738
rect 3799 -1758 3813 -1738
rect 3814 -1751 3825 -1738
rect 3779 -1769 3813 -1758
rect 3814 -1769 3825 -1753
rect 3871 -1762 3887 -1746
rect 3894 -1748 3924 -1696
rect 3958 -1700 3959 -1693
rect 3943 -1708 3959 -1700
rect 3930 -1740 3943 -1721
rect 3958 -1740 3988 -1724
rect 3930 -1756 4004 -1740
rect 3930 -1758 3943 -1756
rect 3958 -1758 3992 -1756
rect 3595 -1780 3608 -1778
rect 3623 -1780 3657 -1778
rect 3595 -1796 3657 -1780
rect 3701 -1785 3717 -1778
rect 3779 -1785 3809 -1774
rect 3857 -1778 3903 -1762
rect 3930 -1774 4004 -1758
rect 3857 -1780 3891 -1778
rect 3856 -1796 3903 -1780
rect 3930 -1796 3943 -1774
rect 3958 -1796 3988 -1774
rect 4015 -1796 4016 -1780
rect 4031 -1796 4044 -1636
rect 4074 -1740 4087 -1636
rect 4132 -1658 4133 -1648
rect 4148 -1658 4161 -1648
rect 4132 -1662 4161 -1658
rect 4166 -1662 4196 -1636
rect 4214 -1650 4230 -1648
rect 4302 -1650 4355 -1636
rect 4303 -1652 4367 -1650
rect 4410 -1652 4425 -1636
rect 4474 -1639 4504 -1636
rect 4474 -1642 4510 -1639
rect 4440 -1650 4456 -1648
rect 4214 -1662 4229 -1658
rect 4132 -1664 4229 -1662
rect 4257 -1664 4425 -1652
rect 4441 -1662 4456 -1658
rect 4474 -1661 4513 -1642
rect 4532 -1648 4539 -1647
rect 4538 -1655 4539 -1648
rect 4522 -1658 4523 -1655
rect 4538 -1658 4551 -1655
rect 4474 -1662 4504 -1661
rect 4513 -1662 4519 -1661
rect 4522 -1662 4551 -1658
rect 4441 -1663 4551 -1662
rect 4441 -1664 4557 -1663
rect 4116 -1672 4167 -1664
rect 4116 -1684 4141 -1672
rect 4148 -1684 4167 -1672
rect 4198 -1672 4248 -1664
rect 4198 -1680 4214 -1672
rect 4221 -1674 4248 -1672
rect 4257 -1674 4478 -1664
rect 4221 -1684 4478 -1674
rect 4507 -1672 4557 -1664
rect 4507 -1681 4523 -1672
rect 4116 -1692 4167 -1684
rect 4214 -1692 4478 -1684
rect 4504 -1684 4523 -1681
rect 4530 -1684 4557 -1672
rect 4504 -1692 4557 -1684
rect 4132 -1700 4133 -1692
rect 4148 -1700 4161 -1692
rect 4132 -1708 4148 -1700
rect 4129 -1715 4148 -1712
rect 4129 -1724 4151 -1715
rect 4102 -1734 4151 -1724
rect 4102 -1740 4132 -1734
rect 4151 -1739 4156 -1734
rect 4074 -1756 4148 -1740
rect 4166 -1748 4196 -1692
rect 4231 -1702 4439 -1692
rect 4474 -1696 4519 -1692
rect 4522 -1693 4523 -1692
rect 4538 -1693 4551 -1692
rect 4257 -1732 4446 -1702
rect 4272 -1735 4446 -1732
rect 4265 -1738 4446 -1735
rect 4074 -1758 4087 -1756
rect 4102 -1758 4136 -1756
rect 4074 -1774 4148 -1758
rect 4175 -1762 4188 -1748
rect 4203 -1762 4219 -1746
rect 4265 -1751 4276 -1738
rect 4058 -1796 4059 -1780
rect 4074 -1796 4087 -1774
rect 4102 -1796 4132 -1774
rect 4175 -1778 4237 -1762
rect 4265 -1769 4276 -1753
rect 4281 -1758 4291 -1738
rect 4301 -1758 4315 -1738
rect 4318 -1751 4327 -1738
rect 4343 -1751 4352 -1738
rect 4281 -1769 4315 -1758
rect 4318 -1769 4327 -1753
rect 4343 -1769 4352 -1753
rect 4359 -1758 4369 -1738
rect 4379 -1758 4393 -1738
rect 4394 -1751 4405 -1738
rect 4359 -1769 4393 -1758
rect 4394 -1769 4405 -1753
rect 4451 -1762 4467 -1746
rect 4474 -1748 4504 -1696
rect 4538 -1700 4539 -1693
rect 4523 -1708 4539 -1700
rect 4510 -1740 4523 -1721
rect 4538 -1740 4568 -1724
rect 4510 -1756 4584 -1740
rect 4510 -1758 4523 -1756
rect 4538 -1758 4572 -1756
rect 4175 -1780 4188 -1778
rect 4203 -1780 4237 -1778
rect 4175 -1796 4237 -1780
rect 4281 -1785 4297 -1778
rect 4359 -1785 4389 -1774
rect 4437 -1778 4483 -1762
rect 4510 -1774 4584 -1758
rect 4437 -1780 4471 -1778
rect 4436 -1796 4483 -1780
rect 4510 -1796 4523 -1774
rect 4538 -1796 4568 -1774
rect 4595 -1796 4596 -1780
rect 4611 -1796 4624 -1636
rect 4654 -1740 4667 -1636
rect 4712 -1658 4713 -1648
rect 4728 -1658 4741 -1648
rect 4712 -1662 4741 -1658
rect 4746 -1662 4776 -1636
rect 4794 -1650 4810 -1648
rect 4882 -1650 4933 -1636
rect 4883 -1652 4947 -1650
rect 4990 -1652 5005 -1636
rect 5054 -1639 5084 -1636
rect 5054 -1642 5090 -1639
rect 5020 -1650 5036 -1648
rect 4794 -1662 4809 -1658
rect 4712 -1664 4809 -1662
rect 4837 -1664 5005 -1652
rect 5021 -1662 5036 -1658
rect 5054 -1661 5093 -1642
rect 5112 -1648 5119 -1647
rect 5118 -1655 5119 -1648
rect 5102 -1658 5103 -1655
rect 5118 -1658 5131 -1655
rect 5054 -1662 5084 -1661
rect 5093 -1662 5099 -1661
rect 5102 -1662 5131 -1658
rect 5021 -1663 5131 -1662
rect 5021 -1664 5137 -1663
rect 4696 -1672 4747 -1664
rect 4696 -1684 4721 -1672
rect 4728 -1684 4747 -1672
rect 4778 -1672 4828 -1664
rect 4778 -1680 4794 -1672
rect 4801 -1674 4828 -1672
rect 4837 -1674 5058 -1664
rect 4801 -1684 5058 -1674
rect 5087 -1672 5137 -1664
rect 5087 -1681 5103 -1672
rect 4696 -1692 4747 -1684
rect 4794 -1692 5058 -1684
rect 5084 -1684 5103 -1681
rect 5110 -1684 5137 -1672
rect 5084 -1692 5137 -1684
rect 4712 -1700 4713 -1692
rect 4728 -1700 4741 -1692
rect 4712 -1708 4728 -1700
rect 4709 -1715 4728 -1712
rect 4709 -1724 4731 -1715
rect 4682 -1734 4731 -1724
rect 4682 -1740 4712 -1734
rect 4731 -1739 4736 -1734
rect 4654 -1756 4728 -1740
rect 4746 -1748 4776 -1692
rect 4811 -1702 5019 -1692
rect 5054 -1696 5099 -1692
rect 5102 -1693 5103 -1692
rect 5118 -1693 5131 -1692
rect 4837 -1732 5026 -1702
rect 4852 -1735 5026 -1732
rect 4845 -1738 5026 -1735
rect 4654 -1758 4667 -1756
rect 4682 -1758 4716 -1756
rect 4654 -1774 4728 -1758
rect 4755 -1762 4768 -1748
rect 4783 -1762 4799 -1746
rect 4845 -1751 4856 -1738
rect 4638 -1796 4639 -1780
rect 4654 -1796 4667 -1774
rect 4682 -1796 4712 -1774
rect 4755 -1778 4817 -1762
rect 4845 -1769 4856 -1753
rect 4861 -1758 4871 -1738
rect 4881 -1758 4895 -1738
rect 4898 -1751 4907 -1738
rect 4923 -1751 4932 -1738
rect 4861 -1769 4895 -1758
rect 4898 -1769 4907 -1753
rect 4923 -1769 4932 -1753
rect 4939 -1758 4949 -1738
rect 4959 -1758 4973 -1738
rect 4974 -1751 4985 -1738
rect 4939 -1769 4973 -1758
rect 4974 -1769 4985 -1753
rect 5031 -1762 5047 -1746
rect 5054 -1748 5084 -1696
rect 5118 -1700 5119 -1693
rect 5103 -1708 5119 -1700
rect 5090 -1740 5103 -1721
rect 5118 -1740 5148 -1724
rect 5090 -1756 5164 -1740
rect 5090 -1758 5103 -1756
rect 5118 -1758 5152 -1756
rect 4755 -1780 4768 -1778
rect 4783 -1780 4817 -1778
rect 4755 -1796 4817 -1780
rect 4861 -1785 4877 -1778
rect 4939 -1785 4969 -1774
rect 5017 -1778 5063 -1762
rect 5090 -1774 5164 -1758
rect 5017 -1780 5051 -1778
rect 5016 -1796 5063 -1780
rect 5090 -1796 5103 -1774
rect 5118 -1796 5148 -1774
rect 5175 -1796 5176 -1780
rect 5191 -1796 5204 -1636
rect 5234 -1740 5247 -1636
rect 5292 -1658 5293 -1648
rect 5308 -1658 5321 -1648
rect 5292 -1662 5321 -1658
rect 5326 -1662 5356 -1636
rect 5374 -1650 5390 -1648
rect 5462 -1650 5513 -1636
rect 5463 -1652 5527 -1650
rect 5570 -1652 5585 -1636
rect 5634 -1639 5664 -1636
rect 5634 -1642 5670 -1639
rect 5600 -1650 5616 -1648
rect 5374 -1662 5389 -1658
rect 5292 -1664 5389 -1662
rect 5417 -1664 5585 -1652
rect 5601 -1662 5616 -1658
rect 5634 -1661 5673 -1642
rect 5692 -1648 5699 -1647
rect 5698 -1655 5699 -1648
rect 5682 -1658 5683 -1655
rect 5698 -1658 5711 -1655
rect 5634 -1662 5664 -1661
rect 5673 -1662 5679 -1661
rect 5682 -1662 5711 -1658
rect 5601 -1663 5711 -1662
rect 5601 -1664 5717 -1663
rect 5276 -1672 5327 -1664
rect 5276 -1684 5301 -1672
rect 5308 -1684 5327 -1672
rect 5358 -1672 5408 -1664
rect 5358 -1680 5374 -1672
rect 5381 -1674 5408 -1672
rect 5417 -1674 5638 -1664
rect 5381 -1684 5638 -1674
rect 5667 -1672 5717 -1664
rect 5667 -1681 5683 -1672
rect 5276 -1692 5327 -1684
rect 5374 -1692 5638 -1684
rect 5664 -1684 5683 -1681
rect 5690 -1684 5717 -1672
rect 5664 -1692 5717 -1684
rect 5292 -1700 5293 -1692
rect 5308 -1700 5321 -1692
rect 5292 -1708 5308 -1700
rect 5289 -1715 5308 -1712
rect 5289 -1724 5311 -1715
rect 5262 -1734 5311 -1724
rect 5262 -1740 5292 -1734
rect 5311 -1739 5316 -1734
rect 5234 -1756 5308 -1740
rect 5326 -1748 5356 -1692
rect 5391 -1702 5599 -1692
rect 5634 -1696 5679 -1692
rect 5682 -1693 5683 -1692
rect 5698 -1693 5711 -1692
rect 5417 -1732 5606 -1702
rect 5432 -1735 5606 -1732
rect 5425 -1738 5606 -1735
rect 5234 -1758 5247 -1756
rect 5262 -1758 5296 -1756
rect 5234 -1774 5308 -1758
rect 5335 -1762 5348 -1748
rect 5363 -1762 5379 -1746
rect 5425 -1751 5436 -1738
rect 5218 -1796 5219 -1780
rect 5234 -1796 5247 -1774
rect 5262 -1796 5292 -1774
rect 5335 -1778 5397 -1762
rect 5425 -1769 5436 -1753
rect 5441 -1758 5451 -1738
rect 5461 -1758 5475 -1738
rect 5478 -1751 5487 -1738
rect 5503 -1751 5512 -1738
rect 5441 -1769 5475 -1758
rect 5478 -1769 5487 -1753
rect 5503 -1769 5512 -1753
rect 5519 -1758 5529 -1738
rect 5539 -1758 5553 -1738
rect 5554 -1751 5565 -1738
rect 5519 -1769 5553 -1758
rect 5554 -1769 5565 -1753
rect 5611 -1762 5627 -1746
rect 5634 -1748 5664 -1696
rect 5698 -1700 5699 -1693
rect 5683 -1708 5699 -1700
rect 5670 -1740 5683 -1721
rect 5698 -1740 5728 -1724
rect 5670 -1756 5744 -1740
rect 5670 -1758 5683 -1756
rect 5698 -1758 5732 -1756
rect 5335 -1780 5348 -1778
rect 5363 -1780 5397 -1778
rect 5335 -1796 5397 -1780
rect 5441 -1785 5457 -1778
rect 5519 -1785 5549 -1774
rect 5597 -1778 5643 -1762
rect 5670 -1774 5744 -1758
rect 5597 -1780 5631 -1778
rect 5596 -1796 5643 -1780
rect 5670 -1796 5683 -1774
rect 5698 -1796 5728 -1774
rect 5755 -1796 5756 -1780
rect 5771 -1796 5784 -1636
rect 5814 -1740 5827 -1636
rect 5872 -1658 5873 -1648
rect 5888 -1658 5901 -1648
rect 5872 -1662 5901 -1658
rect 5906 -1662 5936 -1636
rect 5954 -1650 5970 -1648
rect 6042 -1650 6093 -1636
rect 6043 -1652 6107 -1650
rect 6150 -1652 6165 -1636
rect 6214 -1639 6244 -1636
rect 6214 -1642 6250 -1639
rect 6180 -1650 6196 -1648
rect 5954 -1662 5969 -1658
rect 5872 -1664 5969 -1662
rect 5997 -1664 6165 -1652
rect 6181 -1662 6196 -1658
rect 6214 -1661 6253 -1642
rect 6272 -1648 6279 -1647
rect 6278 -1655 6279 -1648
rect 6262 -1658 6263 -1655
rect 6278 -1658 6291 -1655
rect 6214 -1662 6244 -1661
rect 6253 -1662 6259 -1661
rect 6262 -1662 6291 -1658
rect 6181 -1663 6291 -1662
rect 6181 -1664 6297 -1663
rect 5856 -1672 5907 -1664
rect 5856 -1684 5881 -1672
rect 5888 -1684 5907 -1672
rect 5938 -1672 5988 -1664
rect 5938 -1680 5954 -1672
rect 5961 -1674 5988 -1672
rect 5997 -1674 6218 -1664
rect 5961 -1684 6218 -1674
rect 6247 -1672 6297 -1664
rect 6247 -1681 6263 -1672
rect 5856 -1692 5907 -1684
rect 5954 -1692 6218 -1684
rect 6244 -1684 6263 -1681
rect 6270 -1684 6297 -1672
rect 6244 -1692 6297 -1684
rect 5872 -1700 5873 -1692
rect 5888 -1700 5901 -1692
rect 5872 -1708 5888 -1700
rect 5869 -1715 5888 -1712
rect 5869 -1724 5891 -1715
rect 5842 -1734 5891 -1724
rect 5842 -1740 5872 -1734
rect 5891 -1739 5896 -1734
rect 5814 -1756 5888 -1740
rect 5906 -1748 5936 -1692
rect 5971 -1702 6179 -1692
rect 6214 -1696 6259 -1692
rect 6262 -1693 6263 -1692
rect 6278 -1693 6291 -1692
rect 5997 -1732 6186 -1702
rect 6012 -1735 6186 -1732
rect 6005 -1738 6186 -1735
rect 5814 -1758 5827 -1756
rect 5842 -1758 5876 -1756
rect 5814 -1774 5888 -1758
rect 5915 -1762 5928 -1748
rect 5943 -1762 5959 -1746
rect 6005 -1751 6016 -1738
rect 5798 -1796 5799 -1780
rect 5814 -1796 5827 -1774
rect 5842 -1796 5872 -1774
rect 5915 -1778 5977 -1762
rect 6005 -1769 6016 -1753
rect 6021 -1758 6031 -1738
rect 6041 -1758 6055 -1738
rect 6058 -1751 6067 -1738
rect 6083 -1751 6092 -1738
rect 6021 -1769 6055 -1758
rect 6058 -1769 6067 -1753
rect 6083 -1769 6092 -1753
rect 6099 -1758 6109 -1738
rect 6119 -1758 6133 -1738
rect 6134 -1751 6145 -1738
rect 6099 -1769 6133 -1758
rect 6134 -1769 6145 -1753
rect 6191 -1762 6207 -1746
rect 6214 -1748 6244 -1696
rect 6278 -1700 6279 -1693
rect 6263 -1708 6279 -1700
rect 6250 -1740 6263 -1721
rect 6278 -1740 6308 -1724
rect 6250 -1756 6324 -1740
rect 6250 -1758 6263 -1756
rect 6278 -1758 6312 -1756
rect 5915 -1780 5928 -1778
rect 5943 -1780 5977 -1778
rect 5915 -1796 5977 -1780
rect 6021 -1785 6037 -1778
rect 6099 -1785 6129 -1774
rect 6177 -1778 6223 -1762
rect 6250 -1774 6324 -1758
rect 6177 -1780 6211 -1778
rect 6176 -1796 6223 -1780
rect 6250 -1796 6263 -1774
rect 6278 -1796 6308 -1774
rect 6335 -1796 6336 -1780
rect 6351 -1796 6364 -1636
rect 6394 -1740 6407 -1636
rect 6452 -1658 6453 -1648
rect 6468 -1658 6481 -1648
rect 6452 -1662 6481 -1658
rect 6486 -1662 6516 -1636
rect 6534 -1650 6550 -1648
rect 6622 -1650 6673 -1636
rect 6623 -1652 6687 -1650
rect 6730 -1652 6745 -1636
rect 6794 -1639 6824 -1636
rect 6794 -1642 6830 -1639
rect 6760 -1650 6776 -1648
rect 6534 -1662 6549 -1658
rect 6452 -1664 6549 -1662
rect 6577 -1664 6745 -1652
rect 6761 -1662 6776 -1658
rect 6794 -1661 6833 -1642
rect 6852 -1648 6859 -1647
rect 6858 -1655 6859 -1648
rect 6842 -1658 6843 -1655
rect 6858 -1658 6871 -1655
rect 6794 -1662 6824 -1661
rect 6833 -1662 6839 -1661
rect 6842 -1662 6871 -1658
rect 6761 -1663 6871 -1662
rect 6761 -1664 6877 -1663
rect 6436 -1672 6487 -1664
rect 6436 -1684 6461 -1672
rect 6468 -1684 6487 -1672
rect 6518 -1672 6568 -1664
rect 6518 -1680 6534 -1672
rect 6541 -1674 6568 -1672
rect 6577 -1674 6798 -1664
rect 6541 -1684 6798 -1674
rect 6827 -1672 6877 -1664
rect 6827 -1681 6843 -1672
rect 6436 -1692 6487 -1684
rect 6534 -1692 6798 -1684
rect 6824 -1684 6843 -1681
rect 6850 -1684 6877 -1672
rect 6824 -1692 6877 -1684
rect 6452 -1700 6453 -1692
rect 6468 -1700 6481 -1692
rect 6452 -1708 6468 -1700
rect 6449 -1715 6468 -1712
rect 6449 -1724 6471 -1715
rect 6422 -1734 6471 -1724
rect 6422 -1740 6452 -1734
rect 6471 -1739 6476 -1734
rect 6394 -1756 6468 -1740
rect 6486 -1748 6516 -1692
rect 6551 -1702 6759 -1692
rect 6794 -1696 6839 -1692
rect 6842 -1693 6843 -1692
rect 6858 -1693 6871 -1692
rect 6577 -1732 6766 -1702
rect 6592 -1735 6766 -1732
rect 6585 -1738 6766 -1735
rect 6394 -1758 6407 -1756
rect 6422 -1758 6456 -1756
rect 6394 -1774 6468 -1758
rect 6495 -1762 6508 -1748
rect 6523 -1762 6539 -1746
rect 6585 -1751 6596 -1738
rect 6378 -1796 6379 -1780
rect 6394 -1796 6407 -1774
rect 6422 -1796 6452 -1774
rect 6495 -1778 6557 -1762
rect 6585 -1769 6596 -1753
rect 6601 -1758 6611 -1738
rect 6621 -1758 6635 -1738
rect 6638 -1751 6647 -1738
rect 6663 -1751 6672 -1738
rect 6601 -1769 6635 -1758
rect 6638 -1769 6647 -1753
rect 6663 -1769 6672 -1753
rect 6679 -1758 6689 -1738
rect 6699 -1758 6713 -1738
rect 6714 -1751 6725 -1738
rect 6679 -1769 6713 -1758
rect 6714 -1769 6725 -1753
rect 6771 -1762 6787 -1746
rect 6794 -1748 6824 -1696
rect 6858 -1700 6859 -1693
rect 6843 -1708 6859 -1700
rect 6830 -1740 6843 -1721
rect 6858 -1740 6888 -1724
rect 6830 -1756 6904 -1740
rect 6830 -1758 6843 -1756
rect 6858 -1758 6892 -1756
rect 6495 -1780 6508 -1778
rect 6523 -1780 6557 -1778
rect 6495 -1796 6557 -1780
rect 6601 -1785 6617 -1778
rect 6679 -1785 6709 -1774
rect 6757 -1778 6803 -1762
rect 6830 -1774 6904 -1758
rect 6757 -1780 6791 -1778
rect 6756 -1796 6803 -1780
rect 6830 -1796 6843 -1774
rect 6858 -1796 6888 -1774
rect 6915 -1796 6916 -1780
rect 6931 -1796 6944 -1636
rect -8 -1804 33 -1796
rect -8 -1830 7 -1804
rect 14 -1830 33 -1804
rect 97 -1808 159 -1796
rect 171 -1808 246 -1796
rect 304 -1808 379 -1796
rect 391 -1808 422 -1796
rect 428 -1808 463 -1796
rect 97 -1810 259 -1808
rect -8 -1838 33 -1830
rect 115 -1834 128 -1810
rect 143 -1812 158 -1810
rect -2 -1848 -1 -1838
rect 14 -1848 27 -1838
rect 42 -1848 72 -1834
rect 115 -1848 158 -1834
rect 182 -1837 189 -1830
rect 192 -1834 259 -1810
rect 291 -1810 463 -1808
rect 261 -1832 289 -1828
rect 291 -1832 371 -1810
rect 392 -1812 407 -1810
rect 261 -1834 371 -1832
rect 192 -1838 371 -1834
rect 165 -1848 195 -1838
rect 197 -1848 350 -1838
rect 358 -1848 388 -1838
rect 392 -1848 422 -1834
rect 450 -1848 463 -1810
rect 535 -1804 570 -1796
rect 535 -1830 536 -1804
rect 543 -1830 570 -1804
rect 478 -1848 508 -1834
rect 535 -1838 570 -1830
rect 572 -1804 613 -1796
rect 572 -1830 587 -1804
rect 594 -1830 613 -1804
rect 677 -1808 739 -1796
rect 751 -1808 826 -1796
rect 884 -1808 959 -1796
rect 971 -1808 1002 -1796
rect 1008 -1808 1043 -1796
rect 677 -1810 839 -1808
rect 572 -1838 613 -1830
rect 695 -1834 708 -1810
rect 723 -1812 738 -1810
rect 535 -1848 536 -1838
rect 551 -1848 564 -1838
rect 578 -1848 579 -1838
rect 594 -1848 607 -1838
rect 622 -1848 652 -1834
rect 695 -1848 738 -1834
rect 762 -1837 769 -1830
rect 772 -1834 839 -1810
rect 871 -1810 1043 -1808
rect 841 -1832 869 -1828
rect 871 -1832 951 -1810
rect 972 -1812 987 -1810
rect 841 -1834 951 -1832
rect 772 -1838 951 -1834
rect 745 -1848 775 -1838
rect 777 -1848 930 -1838
rect 938 -1848 968 -1838
rect 972 -1848 1002 -1834
rect 1030 -1848 1043 -1810
rect 1115 -1804 1150 -1796
rect 1115 -1830 1116 -1804
rect 1123 -1830 1150 -1804
rect 1058 -1848 1088 -1834
rect 1115 -1838 1150 -1830
rect 1152 -1804 1193 -1796
rect 1152 -1830 1167 -1804
rect 1174 -1830 1193 -1804
rect 1257 -1808 1319 -1796
rect 1331 -1808 1406 -1796
rect 1464 -1808 1539 -1796
rect 3435 -1804 3470 -1796
rect 1257 -1810 1419 -1808
rect 1152 -1838 1193 -1830
rect 1275 -1834 1288 -1810
rect 1303 -1812 1318 -1810
rect 1115 -1848 1116 -1838
rect 1131 -1848 1144 -1838
rect 1158 -1848 1159 -1838
rect 1174 -1848 1187 -1838
rect 1202 -1848 1232 -1834
rect 1275 -1848 1318 -1834
rect 1342 -1837 1349 -1830
rect 1352 -1834 1419 -1810
rect 1451 -1810 1551 -1808
rect 1421 -1832 1449 -1828
rect 1451 -1832 1531 -1810
rect 1421 -1834 1531 -1832
rect 3435 -1830 3436 -1804
rect 3443 -1830 3470 -1804
rect 1352 -1838 1531 -1834
rect 1325 -1848 1355 -1838
rect 1357 -1848 1510 -1838
rect 1518 -1848 1548 -1838
rect 3379 -1848 3408 -1834
rect 3435 -1838 3470 -1830
rect 3472 -1804 3513 -1796
rect 3472 -1830 3487 -1804
rect 3494 -1830 3513 -1804
rect 3577 -1808 3639 -1796
rect 3651 -1808 3726 -1796
rect 3784 -1808 3859 -1796
rect 3871 -1808 3902 -1796
rect 3908 -1808 3943 -1796
rect 3577 -1810 3739 -1808
rect 3472 -1838 3513 -1830
rect 3595 -1834 3608 -1810
rect 3623 -1812 3638 -1810
rect 3435 -1848 3436 -1838
rect 3451 -1848 3464 -1838
rect 3478 -1848 3479 -1838
rect 3494 -1848 3507 -1838
rect 3522 -1848 3552 -1834
rect 3595 -1848 3638 -1834
rect 3662 -1837 3669 -1830
rect 3672 -1834 3739 -1810
rect 3771 -1810 3943 -1808
rect 3741 -1832 3769 -1828
rect 3771 -1832 3851 -1810
rect 3872 -1812 3887 -1810
rect 3741 -1834 3851 -1832
rect 3672 -1838 3851 -1834
rect 3645 -1848 3675 -1838
rect 3677 -1848 3830 -1838
rect 3838 -1848 3868 -1838
rect 3872 -1848 3902 -1834
rect 3930 -1848 3943 -1810
rect 4015 -1804 4050 -1796
rect 4015 -1830 4016 -1804
rect 4023 -1830 4050 -1804
rect 3958 -1848 3988 -1834
rect 4015 -1838 4050 -1830
rect 4052 -1804 4093 -1796
rect 4052 -1830 4067 -1804
rect 4074 -1830 4093 -1804
rect 4157 -1808 4219 -1796
rect 4231 -1808 4306 -1796
rect 4364 -1808 4439 -1796
rect 4451 -1808 4482 -1796
rect 4488 -1808 4523 -1796
rect 4157 -1810 4319 -1808
rect 4052 -1838 4093 -1830
rect 4175 -1834 4188 -1810
rect 4203 -1812 4218 -1810
rect 4015 -1848 4016 -1838
rect 4031 -1848 4044 -1838
rect 4058 -1848 4059 -1838
rect 4074 -1848 4087 -1838
rect 4102 -1848 4132 -1834
rect 4175 -1848 4218 -1834
rect 4242 -1837 4249 -1830
rect 4252 -1834 4319 -1810
rect 4351 -1810 4523 -1808
rect 4321 -1832 4349 -1828
rect 4351 -1832 4431 -1810
rect 4452 -1812 4467 -1810
rect 4321 -1834 4431 -1832
rect 4252 -1838 4431 -1834
rect 4225 -1848 4255 -1838
rect 4257 -1848 4410 -1838
rect 4418 -1848 4448 -1838
rect 4452 -1848 4482 -1834
rect 4510 -1848 4523 -1810
rect 4595 -1804 4630 -1796
rect 4595 -1830 4596 -1804
rect 4603 -1830 4630 -1804
rect 4538 -1848 4568 -1834
rect 4595 -1838 4630 -1830
rect 4632 -1804 4673 -1796
rect 4632 -1830 4647 -1804
rect 4654 -1830 4673 -1804
rect 4737 -1808 4799 -1796
rect 4811 -1808 4886 -1796
rect 4944 -1808 5019 -1796
rect 5031 -1808 5062 -1796
rect 5068 -1808 5103 -1796
rect 4737 -1810 4899 -1808
rect 4632 -1838 4673 -1830
rect 4755 -1834 4768 -1810
rect 4783 -1812 4798 -1810
rect 4832 -1828 4899 -1810
rect 4931 -1810 5103 -1808
rect 4931 -1828 5011 -1810
rect 5032 -1812 5047 -1810
rect 4595 -1848 4596 -1838
rect 4611 -1848 4624 -1838
rect 4638 -1848 4639 -1838
rect 4654 -1848 4667 -1838
rect 4682 -1848 4712 -1834
rect 4755 -1848 4798 -1834
rect 4822 -1837 4829 -1830
rect 4832 -1838 5011 -1828
rect 4805 -1848 4835 -1838
rect 4837 -1848 4990 -1838
rect 4998 -1848 5028 -1838
rect 5032 -1848 5062 -1834
rect 5090 -1848 5103 -1810
rect 5175 -1804 5210 -1796
rect 5175 -1830 5176 -1804
rect 5183 -1830 5210 -1804
rect 5118 -1848 5148 -1834
rect 5175 -1838 5210 -1830
rect 5212 -1804 5253 -1796
rect 5212 -1830 5227 -1804
rect 5234 -1830 5253 -1804
rect 5317 -1808 5379 -1796
rect 5391 -1808 5466 -1796
rect 5524 -1808 5599 -1796
rect 5611 -1808 5642 -1796
rect 5648 -1808 5683 -1796
rect 5317 -1810 5479 -1808
rect 5212 -1838 5253 -1830
rect 5335 -1834 5348 -1810
rect 5363 -1812 5378 -1810
rect 5412 -1828 5479 -1810
rect 5511 -1810 5683 -1808
rect 5511 -1828 5591 -1810
rect 5612 -1812 5627 -1810
rect 5175 -1848 5176 -1838
rect 5191 -1848 5204 -1838
rect 5218 -1848 5219 -1838
rect 5234 -1848 5247 -1838
rect 5262 -1848 5292 -1834
rect 5335 -1848 5378 -1834
rect 5402 -1837 5409 -1830
rect 5412 -1838 5591 -1828
rect 5385 -1848 5415 -1838
rect 5417 -1848 5570 -1838
rect 5578 -1848 5608 -1838
rect 5612 -1848 5642 -1834
rect 5670 -1848 5683 -1810
rect 5755 -1804 5790 -1796
rect 5755 -1830 5756 -1804
rect 5763 -1830 5790 -1804
rect 5698 -1848 5728 -1834
rect 5755 -1838 5790 -1830
rect 5792 -1804 5833 -1796
rect 5792 -1830 5807 -1804
rect 5814 -1830 5833 -1804
rect 5897 -1808 5959 -1796
rect 5971 -1808 6046 -1796
rect 6104 -1808 6179 -1796
rect 6191 -1808 6222 -1796
rect 6228 -1808 6263 -1796
rect 5897 -1810 6059 -1808
rect 5792 -1838 5833 -1830
rect 5915 -1834 5928 -1810
rect 5943 -1812 5958 -1810
rect 5992 -1828 6059 -1810
rect 6091 -1810 6263 -1808
rect 6091 -1828 6171 -1810
rect 6192 -1812 6207 -1810
rect 5755 -1848 5756 -1838
rect 5771 -1848 5784 -1838
rect 5798 -1848 5799 -1838
rect 5814 -1848 5827 -1838
rect 5842 -1848 5872 -1834
rect 5915 -1848 5958 -1834
rect 5982 -1837 5989 -1830
rect 5992 -1838 6171 -1828
rect 5965 -1848 5995 -1838
rect 5997 -1848 6150 -1838
rect 6158 -1848 6188 -1838
rect 6192 -1848 6222 -1834
rect 6250 -1848 6263 -1810
rect 6335 -1804 6370 -1796
rect 6335 -1830 6336 -1804
rect 6343 -1830 6370 -1804
rect 6278 -1848 6308 -1834
rect 6335 -1838 6370 -1830
rect 6372 -1804 6413 -1796
rect 6372 -1830 6387 -1804
rect 6394 -1830 6413 -1804
rect 6477 -1808 6539 -1796
rect 6551 -1808 6626 -1796
rect 6684 -1808 6759 -1796
rect 6771 -1808 6802 -1796
rect 6808 -1808 6843 -1796
rect 6477 -1810 6639 -1808
rect 6372 -1838 6413 -1830
rect 6495 -1834 6508 -1810
rect 6523 -1812 6538 -1810
rect 6572 -1828 6639 -1810
rect 6671 -1810 6843 -1808
rect 6671 -1828 6751 -1810
rect 6772 -1812 6787 -1810
rect 6335 -1848 6336 -1838
rect 6351 -1848 6364 -1838
rect 6378 -1848 6379 -1838
rect 6394 -1848 6407 -1838
rect 6422 -1848 6452 -1834
rect 6495 -1848 6538 -1834
rect 6562 -1837 6569 -1830
rect 6572 -1838 6751 -1828
rect 6545 -1848 6575 -1838
rect 6577 -1848 6730 -1838
rect 6738 -1848 6768 -1838
rect 6772 -1848 6802 -1834
rect 6830 -1848 6843 -1810
rect 6915 -1804 6950 -1796
rect 6915 -1830 6916 -1804
rect 6923 -1830 6950 -1804
rect 6858 -1848 6888 -1834
rect 6915 -1838 6950 -1830
rect 6915 -1848 6916 -1838
rect 6931 -1848 6944 -1838
rect -2 -1854 1551 -1848
rect -1 -1862 1551 -1854
rect 3379 -1862 6944 -1848
rect 14 -1892 27 -1862
rect 42 -1880 72 -1862
rect 115 -1876 129 -1862
rect 165 -1876 385 -1862
rect 116 -1878 129 -1876
rect 82 -1890 97 -1878
rect 79 -1892 101 -1890
rect 106 -1892 136 -1878
rect 197 -1880 350 -1876
rect 179 -1892 371 -1880
rect 414 -1892 444 -1878
rect 450 -1892 463 -1862
rect 478 -1880 508 -1862
rect 551 -1892 564 -1862
rect 594 -1892 607 -1862
rect 622 -1880 652 -1862
rect 695 -1876 709 -1862
rect 745 -1876 965 -1862
rect 696 -1878 709 -1876
rect 662 -1890 677 -1878
rect 659 -1892 681 -1890
rect 686 -1892 716 -1878
rect 777 -1880 930 -1876
rect 759 -1892 951 -1880
rect 994 -1892 1024 -1878
rect 1030 -1892 1043 -1862
rect 1058 -1880 1088 -1862
rect 1131 -1892 1144 -1862
rect 1174 -1892 1187 -1862
rect 1202 -1880 1232 -1862
rect 1275 -1876 1289 -1862
rect 1325 -1876 1545 -1862
rect 1276 -1878 1289 -1876
rect 1242 -1890 1257 -1878
rect 1239 -1892 1261 -1890
rect 1266 -1892 1296 -1878
rect 1357 -1880 1510 -1876
rect 3379 -1880 3408 -1862
rect 1339 -1892 1531 -1880
rect 3451 -1892 3464 -1862
rect 3494 -1892 3507 -1862
rect 3522 -1880 3552 -1862
rect 3595 -1876 3609 -1862
rect 3645 -1876 3865 -1862
rect 3596 -1878 3609 -1876
rect 3562 -1890 3577 -1878
rect 3559 -1892 3581 -1890
rect 3586 -1892 3616 -1878
rect 3677 -1880 3830 -1876
rect 3659 -1892 3851 -1880
rect 3894 -1892 3924 -1878
rect 3930 -1892 3943 -1862
rect 3958 -1880 3988 -1862
rect 4031 -1892 4044 -1862
rect 4074 -1892 4087 -1862
rect 4102 -1880 4132 -1862
rect 4175 -1876 4189 -1862
rect 4225 -1876 4445 -1862
rect 4176 -1878 4189 -1876
rect 4142 -1890 4157 -1878
rect 4139 -1892 4161 -1890
rect 4166 -1892 4196 -1878
rect 4257 -1880 4410 -1876
rect 4239 -1892 4431 -1880
rect 4474 -1892 4504 -1878
rect 4510 -1892 4523 -1862
rect 4538 -1880 4568 -1862
rect 4611 -1892 4624 -1862
rect 4654 -1892 4667 -1862
rect 4682 -1880 4712 -1862
rect 4755 -1876 4769 -1862
rect 4805 -1876 5025 -1862
rect 4756 -1878 4769 -1876
rect 4722 -1890 4737 -1878
rect 4719 -1892 4741 -1890
rect 4746 -1892 4776 -1878
rect 4837 -1880 4990 -1876
rect 4819 -1892 5011 -1880
rect 5054 -1892 5084 -1878
rect 5090 -1892 5103 -1862
rect 5118 -1880 5148 -1862
rect 5191 -1892 5204 -1862
rect 5234 -1892 5247 -1862
rect 5262 -1880 5292 -1862
rect 5335 -1876 5349 -1862
rect 5385 -1876 5605 -1862
rect 5336 -1878 5349 -1876
rect 5302 -1890 5317 -1878
rect 5299 -1892 5321 -1890
rect 5326 -1892 5356 -1878
rect 5417 -1880 5570 -1876
rect 5399 -1892 5591 -1880
rect 5634 -1892 5664 -1878
rect 5670 -1892 5683 -1862
rect 5698 -1880 5728 -1862
rect 5771 -1892 5784 -1862
rect 5814 -1892 5827 -1862
rect 5842 -1880 5872 -1862
rect 5915 -1876 5929 -1862
rect 5965 -1876 6185 -1862
rect 5916 -1878 5929 -1876
rect 5882 -1890 5897 -1878
rect 5879 -1892 5901 -1890
rect 5906 -1892 5936 -1878
rect 5997 -1880 6150 -1876
rect 5979 -1892 6171 -1880
rect 6214 -1892 6244 -1878
rect 6250 -1892 6263 -1862
rect 6278 -1880 6308 -1862
rect 6351 -1892 6364 -1862
rect 6394 -1892 6407 -1862
rect 6422 -1880 6452 -1862
rect 6495 -1876 6509 -1862
rect 6545 -1876 6765 -1862
rect 6496 -1878 6509 -1876
rect 6462 -1890 6477 -1878
rect 6459 -1892 6481 -1890
rect 6486 -1892 6516 -1878
rect 6577 -1880 6730 -1876
rect 6559 -1892 6751 -1880
rect 6794 -1892 6824 -1878
rect 6830 -1892 6843 -1862
rect 6858 -1880 6888 -1862
rect 6931 -1892 6944 -1862
rect -1 -1906 1551 -1892
rect 3379 -1906 6944 -1892
rect 14 -2010 27 -1906
rect 72 -1928 73 -1918
rect 88 -1928 101 -1918
rect 72 -1932 101 -1928
rect 106 -1932 136 -1906
rect 154 -1920 170 -1918
rect 242 -1920 295 -1906
rect 243 -1922 307 -1920
rect 154 -1932 169 -1928
rect 72 -1934 169 -1932
rect 56 -1942 107 -1934
rect 56 -1954 81 -1942
rect 88 -1954 107 -1942
rect 138 -1942 188 -1934
rect 138 -1950 154 -1942
rect 161 -1944 188 -1942
rect 197 -1942 212 -1938
rect 259 -1942 291 -1922
rect 350 -1934 365 -1906
rect 414 -1909 444 -1906
rect 414 -1912 450 -1909
rect 380 -1920 396 -1918
rect 381 -1932 396 -1928
rect 414 -1931 453 -1912
rect 472 -1918 479 -1917
rect 478 -1925 479 -1918
rect 462 -1928 463 -1925
rect 478 -1928 491 -1925
rect 414 -1932 444 -1931
rect 453 -1932 459 -1931
rect 462 -1932 491 -1928
rect 381 -1933 491 -1932
rect 381 -1934 497 -1933
rect 350 -1942 418 -1934
rect 197 -1944 266 -1942
rect 284 -1944 418 -1942
rect 161 -1948 233 -1944
rect 161 -1950 286 -1948
rect 161 -1954 233 -1950
rect 56 -1962 107 -1954
rect 154 -1958 233 -1954
rect 314 -1958 418 -1944
rect 447 -1942 497 -1934
rect 447 -1951 463 -1942
rect 154 -1962 418 -1958
rect 444 -1954 463 -1951
rect 470 -1954 497 -1942
rect 444 -1962 497 -1954
rect 72 -1970 73 -1962
rect 88 -1970 101 -1962
rect 72 -1978 88 -1970
rect 69 -1985 88 -1982
rect 69 -1994 91 -1985
rect 42 -2004 91 -1994
rect 42 -2010 72 -2004
rect 91 -2009 96 -2004
rect 14 -2026 88 -2010
rect 106 -2018 136 -1962
rect 171 -1972 379 -1962
rect 414 -1966 459 -1962
rect 462 -1963 463 -1962
rect 478 -1963 491 -1962
rect 338 -1976 386 -1972
rect 221 -1998 251 -1989
rect 314 -1996 329 -1989
rect 350 -1998 386 -1976
rect 197 -2002 386 -1998
rect 212 -2005 386 -2002
rect 205 -2008 386 -2005
rect 14 -2028 27 -2026
rect 42 -2028 76 -2026
rect 14 -2044 88 -2028
rect 115 -2032 128 -2018
rect 143 -2032 159 -2016
rect 205 -2021 216 -2008
rect -2 -2066 -1 -2050
rect 14 -2066 27 -2044
rect 42 -2066 72 -2044
rect 115 -2048 177 -2032
rect 205 -2039 216 -2023
rect 221 -2028 231 -2008
rect 241 -2028 255 -2008
rect 258 -2021 267 -2008
rect 283 -2021 292 -2008
rect 221 -2039 255 -2028
rect 258 -2039 267 -2023
rect 283 -2039 292 -2023
rect 299 -2028 309 -2008
rect 319 -2028 333 -2008
rect 334 -2021 345 -2008
rect 299 -2039 333 -2028
rect 334 -2039 345 -2023
rect 391 -2032 407 -2016
rect 414 -2018 444 -1966
rect 478 -1970 479 -1963
rect 463 -1978 479 -1970
rect 450 -2010 463 -1991
rect 478 -2010 508 -1994
rect 450 -2026 524 -2010
rect 450 -2028 463 -2026
rect 478 -2028 512 -2026
rect 115 -2050 128 -2048
rect 143 -2050 177 -2048
rect 115 -2066 177 -2050
rect 221 -2055 237 -2048
rect 299 -2055 329 -2044
rect 377 -2048 423 -2032
rect 450 -2044 524 -2028
rect 377 -2050 411 -2048
rect 376 -2066 423 -2050
rect 450 -2066 463 -2044
rect 478 -2066 508 -2044
rect 535 -2066 536 -2050
rect 551 -2066 564 -1906
rect 594 -2010 607 -1906
rect 652 -1928 653 -1918
rect 668 -1928 681 -1918
rect 652 -1932 681 -1928
rect 686 -1932 716 -1906
rect 734 -1920 750 -1918
rect 822 -1920 875 -1906
rect 823 -1922 887 -1920
rect 734 -1932 749 -1928
rect 652 -1934 749 -1932
rect 636 -1942 687 -1934
rect 636 -1954 661 -1942
rect 668 -1954 687 -1942
rect 718 -1942 768 -1934
rect 718 -1950 734 -1942
rect 741 -1944 768 -1942
rect 777 -1942 792 -1938
rect 839 -1942 871 -1922
rect 930 -1934 945 -1906
rect 994 -1909 1024 -1906
rect 994 -1912 1030 -1909
rect 960 -1920 976 -1918
rect 961 -1932 976 -1928
rect 994 -1931 1033 -1912
rect 1052 -1918 1059 -1917
rect 1058 -1925 1059 -1918
rect 1042 -1928 1043 -1925
rect 1058 -1928 1071 -1925
rect 994 -1932 1024 -1931
rect 1033 -1932 1039 -1931
rect 1042 -1932 1071 -1928
rect 961 -1933 1071 -1932
rect 961 -1934 1077 -1933
rect 930 -1942 998 -1934
rect 777 -1944 846 -1942
rect 864 -1944 998 -1942
rect 741 -1948 813 -1944
rect 741 -1950 866 -1948
rect 741 -1954 813 -1950
rect 636 -1962 687 -1954
rect 734 -1958 813 -1954
rect 894 -1958 998 -1944
rect 1027 -1942 1077 -1934
rect 1027 -1951 1043 -1942
rect 734 -1962 998 -1958
rect 1024 -1954 1043 -1951
rect 1050 -1954 1077 -1942
rect 1024 -1962 1077 -1954
rect 652 -1970 653 -1962
rect 668 -1970 681 -1962
rect 652 -1978 668 -1970
rect 649 -1985 668 -1982
rect 649 -1994 671 -1985
rect 622 -2004 671 -1994
rect 622 -2010 652 -2004
rect 671 -2009 676 -2004
rect 594 -2026 668 -2010
rect 686 -2018 716 -1962
rect 751 -1972 959 -1962
rect 994 -1966 1039 -1962
rect 1042 -1963 1043 -1962
rect 1058 -1963 1071 -1962
rect 918 -1976 966 -1972
rect 801 -1998 831 -1989
rect 894 -1996 909 -1989
rect 930 -1998 966 -1976
rect 777 -2002 966 -1998
rect 792 -2005 966 -2002
rect 785 -2008 966 -2005
rect 594 -2028 607 -2026
rect 622 -2028 656 -2026
rect 594 -2044 668 -2028
rect 695 -2032 708 -2018
rect 723 -2032 739 -2016
rect 785 -2021 796 -2008
rect 578 -2066 579 -2050
rect 594 -2066 607 -2044
rect 622 -2066 652 -2044
rect 695 -2048 757 -2032
rect 785 -2039 796 -2023
rect 801 -2028 811 -2008
rect 821 -2028 835 -2008
rect 838 -2021 847 -2008
rect 863 -2021 872 -2008
rect 801 -2039 835 -2028
rect 838 -2039 847 -2023
rect 863 -2039 872 -2023
rect 879 -2028 889 -2008
rect 899 -2028 913 -2008
rect 914 -2021 925 -2008
rect 879 -2039 913 -2028
rect 914 -2039 925 -2023
rect 971 -2032 987 -2016
rect 994 -2018 1024 -1966
rect 1058 -1970 1059 -1963
rect 1043 -1978 1059 -1970
rect 1030 -2010 1043 -1991
rect 1058 -2010 1088 -1994
rect 1030 -2026 1104 -2010
rect 1030 -2028 1043 -2026
rect 1058 -2028 1092 -2026
rect 695 -2050 708 -2048
rect 723 -2050 757 -2048
rect 695 -2066 757 -2050
rect 801 -2055 817 -2048
rect 879 -2055 909 -2044
rect 957 -2048 1003 -2032
rect 1030 -2044 1104 -2028
rect 957 -2050 991 -2048
rect 956 -2066 1003 -2050
rect 1030 -2066 1043 -2044
rect 1058 -2066 1088 -2044
rect 1115 -2066 1116 -2050
rect 1131 -2066 1144 -1906
rect 1174 -2010 1187 -1906
rect 1232 -1928 1233 -1918
rect 1248 -1928 1261 -1918
rect 1232 -1932 1261 -1928
rect 1266 -1932 1296 -1906
rect 1314 -1920 1330 -1918
rect 1402 -1920 1455 -1906
rect 1403 -1922 1467 -1920
rect 1314 -1932 1329 -1928
rect 1232 -1934 1329 -1932
rect 1216 -1942 1267 -1934
rect 1216 -1954 1241 -1942
rect 1248 -1954 1267 -1942
rect 1298 -1942 1348 -1934
rect 1298 -1950 1314 -1942
rect 1321 -1944 1348 -1942
rect 1357 -1942 1372 -1938
rect 1419 -1942 1451 -1922
rect 1510 -1934 1525 -1906
rect 1540 -1920 1551 -1918
rect 1541 -1934 1551 -1928
rect 1510 -1942 1551 -1934
rect 1357 -1944 1426 -1942
rect 1444 -1944 1551 -1942
rect 1321 -1948 1393 -1944
rect 1321 -1950 1446 -1948
rect 1321 -1954 1393 -1950
rect 1216 -1962 1267 -1954
rect 1314 -1958 1393 -1954
rect 1474 -1958 1551 -1944
rect 1314 -1962 1551 -1958
rect 3379 -1933 3391 -1925
rect 3379 -1962 3397 -1933
rect 1232 -1970 1233 -1962
rect 1248 -1970 1261 -1962
rect 1232 -1978 1248 -1970
rect 1229 -1985 1248 -1982
rect 1229 -1994 1251 -1985
rect 1202 -2004 1251 -1994
rect 1202 -2010 1232 -2004
rect 1251 -2009 1256 -2004
rect 1174 -2026 1248 -2010
rect 1266 -2018 1296 -1962
rect 1331 -1972 1539 -1962
rect 3379 -1963 3391 -1962
rect 1498 -1976 1546 -1972
rect 1381 -1998 1411 -1989
rect 1474 -1996 1489 -1989
rect 1510 -1998 1546 -1976
rect 1357 -2002 1546 -1998
rect 1372 -2005 1546 -2002
rect 1365 -2008 1546 -2005
rect 1174 -2028 1187 -2026
rect 1202 -2028 1236 -2026
rect 1174 -2044 1248 -2028
rect 1275 -2032 1288 -2018
rect 1303 -2032 1319 -2016
rect 1365 -2021 1376 -2008
rect 1158 -2066 1159 -2050
rect 1174 -2066 1187 -2044
rect 1202 -2066 1232 -2044
rect 1275 -2048 1337 -2032
rect 1365 -2039 1376 -2023
rect 1381 -2028 1391 -2008
rect 1401 -2028 1415 -2008
rect 1418 -2021 1427 -2008
rect 1443 -2021 1452 -2008
rect 1381 -2039 1415 -2028
rect 1418 -2039 1427 -2023
rect 1443 -2039 1452 -2023
rect 1459 -2028 1469 -2008
rect 1479 -2028 1493 -2008
rect 1494 -2021 1505 -2008
rect 3379 -2010 3408 -1994
rect 1459 -2039 1493 -2028
rect 1494 -2039 1505 -2023
rect 3379 -2026 3424 -2010
rect 3379 -2028 3412 -2026
rect 1275 -2050 1288 -2048
rect 1303 -2050 1337 -2048
rect 1275 -2066 1337 -2050
rect 1381 -2055 1397 -2048
rect 1459 -2055 1489 -2044
rect 1537 -2050 1551 -2032
rect 1536 -2066 1551 -2050
rect 3379 -2044 3424 -2028
rect 3379 -2066 3408 -2044
rect 3435 -2066 3436 -2050
rect 3451 -2066 3464 -1906
rect 3494 -2010 3507 -1906
rect 3552 -1928 3553 -1918
rect 3568 -1928 3581 -1918
rect 3552 -1932 3581 -1928
rect 3586 -1932 3616 -1906
rect 3634 -1920 3650 -1918
rect 3722 -1920 3775 -1906
rect 3723 -1922 3787 -1920
rect 3634 -1932 3649 -1928
rect 3552 -1934 3649 -1932
rect 3536 -1942 3587 -1934
rect 3536 -1954 3561 -1942
rect 3568 -1954 3587 -1942
rect 3618 -1942 3668 -1934
rect 3618 -1950 3634 -1942
rect 3641 -1944 3668 -1942
rect 3677 -1942 3692 -1938
rect 3739 -1942 3771 -1922
rect 3830 -1934 3845 -1906
rect 3894 -1909 3924 -1906
rect 3894 -1912 3930 -1909
rect 3860 -1920 3876 -1918
rect 3861 -1932 3876 -1928
rect 3894 -1931 3933 -1912
rect 3952 -1918 3959 -1917
rect 3958 -1925 3959 -1918
rect 3942 -1928 3943 -1925
rect 3958 -1928 3971 -1925
rect 3894 -1932 3924 -1931
rect 3933 -1932 3939 -1931
rect 3942 -1932 3971 -1928
rect 3861 -1933 3971 -1932
rect 3861 -1934 3977 -1933
rect 3830 -1942 3898 -1934
rect 3677 -1944 3746 -1942
rect 3764 -1944 3898 -1942
rect 3641 -1948 3713 -1944
rect 3641 -1950 3766 -1948
rect 3641 -1954 3713 -1950
rect 3536 -1962 3587 -1954
rect 3634 -1958 3713 -1954
rect 3794 -1958 3898 -1944
rect 3927 -1942 3977 -1934
rect 3927 -1951 3943 -1942
rect 3634 -1962 3898 -1958
rect 3924 -1954 3943 -1951
rect 3950 -1954 3977 -1942
rect 3924 -1962 3977 -1954
rect 3552 -1970 3553 -1962
rect 3568 -1970 3581 -1962
rect 3552 -1978 3568 -1970
rect 3549 -1985 3568 -1982
rect 3549 -1994 3571 -1985
rect 3522 -2004 3571 -1994
rect 3522 -2010 3552 -2004
rect 3571 -2009 3576 -2004
rect 3494 -2026 3568 -2010
rect 3586 -2018 3616 -1962
rect 3651 -1972 3859 -1962
rect 3894 -1966 3939 -1962
rect 3942 -1963 3943 -1962
rect 3958 -1963 3971 -1962
rect 3818 -1976 3866 -1972
rect 3701 -1998 3731 -1989
rect 3794 -1996 3809 -1989
rect 3830 -1998 3866 -1976
rect 3677 -2002 3866 -1998
rect 3692 -2005 3866 -2002
rect 3685 -2008 3866 -2005
rect 3494 -2028 3507 -2026
rect 3522 -2028 3556 -2026
rect 3494 -2044 3568 -2028
rect 3595 -2032 3608 -2018
rect 3623 -2032 3639 -2016
rect 3685 -2021 3696 -2008
rect 3478 -2066 3479 -2050
rect 3494 -2066 3507 -2044
rect 3522 -2066 3552 -2044
rect 3595 -2048 3657 -2032
rect 3685 -2039 3696 -2023
rect 3701 -2028 3711 -2008
rect 3721 -2028 3735 -2008
rect 3738 -2021 3747 -2008
rect 3763 -2021 3772 -2008
rect 3701 -2039 3735 -2028
rect 3738 -2039 3747 -2023
rect 3763 -2039 3772 -2023
rect 3779 -2028 3789 -2008
rect 3799 -2028 3813 -2008
rect 3814 -2021 3825 -2008
rect 3779 -2039 3813 -2028
rect 3814 -2039 3825 -2023
rect 3871 -2032 3887 -2016
rect 3894 -2018 3924 -1966
rect 3958 -1970 3959 -1963
rect 3943 -1978 3959 -1970
rect 3930 -2010 3943 -1991
rect 3958 -2010 3988 -1994
rect 3930 -2026 4004 -2010
rect 3930 -2028 3943 -2026
rect 3958 -2028 3992 -2026
rect 3595 -2050 3608 -2048
rect 3623 -2050 3657 -2048
rect 3595 -2066 3657 -2050
rect 3701 -2055 3717 -2048
rect 3779 -2055 3809 -2044
rect 3857 -2048 3903 -2032
rect 3930 -2044 4004 -2028
rect 3857 -2050 3891 -2048
rect 3856 -2066 3903 -2050
rect 3930 -2066 3943 -2044
rect 3958 -2066 3988 -2044
rect 4015 -2066 4016 -2050
rect 4031 -2066 4044 -1906
rect 4074 -2010 4087 -1906
rect 4132 -1928 4133 -1918
rect 4148 -1928 4161 -1918
rect 4132 -1932 4161 -1928
rect 4166 -1932 4196 -1906
rect 4214 -1920 4230 -1918
rect 4302 -1920 4355 -1906
rect 4303 -1922 4367 -1920
rect 4214 -1932 4229 -1928
rect 4132 -1934 4229 -1932
rect 4116 -1942 4167 -1934
rect 4116 -1954 4141 -1942
rect 4148 -1954 4167 -1942
rect 4198 -1942 4248 -1934
rect 4198 -1950 4214 -1942
rect 4221 -1944 4248 -1942
rect 4257 -1942 4272 -1938
rect 4319 -1942 4351 -1922
rect 4410 -1934 4425 -1906
rect 4474 -1909 4504 -1906
rect 4474 -1912 4510 -1909
rect 4440 -1920 4456 -1918
rect 4441 -1932 4456 -1928
rect 4474 -1931 4513 -1912
rect 4532 -1918 4539 -1917
rect 4538 -1925 4539 -1918
rect 4522 -1928 4523 -1925
rect 4538 -1928 4551 -1925
rect 4474 -1932 4504 -1931
rect 4513 -1932 4519 -1931
rect 4522 -1932 4551 -1928
rect 4441 -1933 4551 -1932
rect 4441 -1934 4557 -1933
rect 4410 -1942 4478 -1934
rect 4257 -1944 4326 -1942
rect 4344 -1944 4478 -1942
rect 4221 -1948 4293 -1944
rect 4221 -1950 4346 -1948
rect 4221 -1954 4293 -1950
rect 4116 -1962 4167 -1954
rect 4214 -1958 4293 -1954
rect 4374 -1958 4478 -1944
rect 4507 -1942 4557 -1934
rect 4507 -1951 4523 -1942
rect 4214 -1962 4478 -1958
rect 4504 -1954 4523 -1951
rect 4530 -1954 4557 -1942
rect 4504 -1962 4557 -1954
rect 4132 -1970 4133 -1962
rect 4148 -1970 4161 -1962
rect 4132 -1978 4148 -1970
rect 4129 -1985 4148 -1982
rect 4129 -1994 4151 -1985
rect 4102 -2004 4151 -1994
rect 4102 -2010 4132 -2004
rect 4151 -2009 4156 -2004
rect 4074 -2026 4148 -2010
rect 4166 -2018 4196 -1962
rect 4231 -1972 4439 -1962
rect 4474 -1966 4519 -1962
rect 4522 -1963 4523 -1962
rect 4538 -1963 4551 -1962
rect 4398 -1976 4446 -1972
rect 4281 -1998 4311 -1989
rect 4374 -1996 4389 -1989
rect 4410 -1998 4446 -1976
rect 4257 -2002 4446 -1998
rect 4272 -2005 4446 -2002
rect 4265 -2008 4446 -2005
rect 4074 -2028 4087 -2026
rect 4102 -2028 4136 -2026
rect 4074 -2044 4148 -2028
rect 4175 -2032 4188 -2018
rect 4203 -2032 4219 -2016
rect 4265 -2021 4276 -2008
rect 4058 -2066 4059 -2050
rect 4074 -2066 4087 -2044
rect 4102 -2066 4132 -2044
rect 4175 -2048 4237 -2032
rect 4265 -2039 4276 -2023
rect 4281 -2028 4291 -2008
rect 4301 -2028 4315 -2008
rect 4318 -2021 4327 -2008
rect 4343 -2021 4352 -2008
rect 4281 -2039 4315 -2028
rect 4318 -2039 4327 -2023
rect 4343 -2039 4352 -2023
rect 4359 -2028 4369 -2008
rect 4379 -2028 4393 -2008
rect 4394 -2021 4405 -2008
rect 4359 -2039 4393 -2028
rect 4394 -2039 4405 -2023
rect 4451 -2032 4467 -2016
rect 4474 -2018 4504 -1966
rect 4538 -1970 4539 -1963
rect 4523 -1978 4539 -1970
rect 4510 -2010 4523 -1991
rect 4538 -2010 4568 -1994
rect 4510 -2026 4584 -2010
rect 4510 -2028 4523 -2026
rect 4538 -2028 4572 -2026
rect 4175 -2050 4188 -2048
rect 4203 -2050 4237 -2048
rect 4175 -2066 4237 -2050
rect 4281 -2055 4297 -2048
rect 4359 -2055 4389 -2044
rect 4437 -2048 4483 -2032
rect 4510 -2044 4584 -2028
rect 4437 -2050 4471 -2048
rect 4436 -2066 4483 -2050
rect 4510 -2066 4523 -2044
rect 4538 -2066 4568 -2044
rect 4595 -2066 4596 -2050
rect 4611 -2066 4624 -1906
rect 4654 -2010 4667 -1906
rect 4712 -1928 4713 -1918
rect 4728 -1928 4741 -1918
rect 4712 -1932 4741 -1928
rect 4746 -1932 4776 -1906
rect 4794 -1920 4810 -1918
rect 4882 -1920 4933 -1906
rect 4883 -1922 4947 -1920
rect 4794 -1932 4809 -1928
rect 4712 -1934 4809 -1932
rect 4696 -1942 4747 -1934
rect 4696 -1954 4721 -1942
rect 4728 -1954 4747 -1942
rect 4778 -1942 4828 -1934
rect 4778 -1950 4794 -1942
rect 4801 -1944 4828 -1942
rect 4837 -1942 4852 -1938
rect 4899 -1942 4931 -1922
rect 4990 -1934 5005 -1906
rect 5054 -1909 5084 -1906
rect 5054 -1912 5090 -1909
rect 5020 -1920 5036 -1918
rect 5021 -1932 5036 -1928
rect 5054 -1931 5093 -1912
rect 5112 -1918 5119 -1917
rect 5118 -1925 5119 -1918
rect 5102 -1928 5103 -1925
rect 5118 -1928 5131 -1925
rect 5054 -1932 5084 -1931
rect 5093 -1932 5099 -1931
rect 5102 -1932 5131 -1928
rect 5021 -1933 5131 -1932
rect 5021 -1934 5137 -1933
rect 4990 -1942 5058 -1934
rect 4837 -1944 4906 -1942
rect 4924 -1944 5058 -1942
rect 4801 -1948 4873 -1944
rect 4801 -1950 4926 -1948
rect 4801 -1954 4873 -1950
rect 4696 -1962 4747 -1954
rect 4794 -1958 4873 -1954
rect 4954 -1958 5058 -1944
rect 5087 -1942 5137 -1934
rect 5087 -1951 5103 -1942
rect 4794 -1962 5058 -1958
rect 5084 -1954 5103 -1951
rect 5110 -1954 5137 -1942
rect 5084 -1962 5137 -1954
rect 4712 -1970 4713 -1962
rect 4728 -1970 4741 -1962
rect 4712 -1978 4728 -1970
rect 4709 -1985 4728 -1982
rect 4709 -1994 4731 -1985
rect 4682 -2004 4731 -1994
rect 4682 -2010 4712 -2004
rect 4731 -2009 4736 -2004
rect 4654 -2026 4728 -2010
rect 4746 -2018 4776 -1962
rect 4811 -1972 5019 -1962
rect 5054 -1966 5099 -1962
rect 5102 -1963 5103 -1962
rect 5118 -1963 5131 -1962
rect 4978 -1976 5026 -1972
rect 4861 -1998 4891 -1989
rect 4954 -1996 4969 -1989
rect 4990 -1998 5026 -1976
rect 4837 -2002 5026 -1998
rect 4852 -2005 5026 -2002
rect 4845 -2008 5026 -2005
rect 4654 -2028 4667 -2026
rect 4682 -2028 4716 -2026
rect 4654 -2044 4728 -2028
rect 4755 -2032 4768 -2018
rect 4783 -2032 4799 -2016
rect 4845 -2021 4856 -2008
rect 4638 -2066 4639 -2050
rect 4654 -2066 4667 -2044
rect 4682 -2066 4712 -2044
rect 4755 -2048 4817 -2032
rect 4845 -2039 4856 -2023
rect 4861 -2028 4871 -2008
rect 4881 -2028 4895 -2008
rect 4898 -2021 4907 -2008
rect 4923 -2021 4932 -2008
rect 4861 -2039 4895 -2028
rect 4898 -2039 4907 -2023
rect 4923 -2039 4932 -2023
rect 4939 -2028 4949 -2008
rect 4959 -2028 4973 -2008
rect 4974 -2021 4985 -2008
rect 4939 -2039 4973 -2028
rect 4974 -2039 4985 -2023
rect 5031 -2032 5047 -2016
rect 5054 -2018 5084 -1966
rect 5118 -1970 5119 -1963
rect 5103 -1978 5119 -1970
rect 5090 -2010 5103 -1991
rect 5118 -2010 5148 -1994
rect 5090 -2026 5164 -2010
rect 5090 -2028 5103 -2026
rect 5118 -2028 5152 -2026
rect 4755 -2050 4768 -2048
rect 4783 -2050 4817 -2048
rect 4755 -2066 4817 -2050
rect 4861 -2055 4877 -2048
rect 4939 -2055 4969 -2044
rect 5017 -2048 5063 -2032
rect 5090 -2044 5164 -2028
rect 5017 -2050 5051 -2048
rect 5016 -2066 5063 -2050
rect 5090 -2066 5103 -2044
rect 5118 -2066 5148 -2044
rect 5175 -2066 5176 -2050
rect 5191 -2066 5204 -1906
rect 5234 -2010 5247 -1906
rect 5292 -1928 5293 -1918
rect 5308 -1928 5321 -1918
rect 5292 -1932 5321 -1928
rect 5326 -1932 5356 -1906
rect 5374 -1920 5390 -1918
rect 5462 -1920 5513 -1906
rect 5463 -1922 5527 -1920
rect 5374 -1932 5389 -1928
rect 5292 -1934 5389 -1932
rect 5276 -1942 5327 -1934
rect 5276 -1954 5301 -1942
rect 5308 -1954 5327 -1942
rect 5358 -1942 5408 -1934
rect 5358 -1950 5374 -1942
rect 5381 -1944 5408 -1942
rect 5417 -1942 5432 -1938
rect 5479 -1942 5511 -1922
rect 5570 -1934 5585 -1906
rect 5634 -1909 5664 -1906
rect 5634 -1912 5670 -1909
rect 5600 -1920 5616 -1918
rect 5601 -1932 5616 -1928
rect 5634 -1931 5673 -1912
rect 5692 -1918 5699 -1917
rect 5698 -1925 5699 -1918
rect 5682 -1928 5683 -1925
rect 5698 -1928 5711 -1925
rect 5634 -1932 5664 -1931
rect 5673 -1932 5679 -1931
rect 5682 -1932 5711 -1928
rect 5601 -1933 5711 -1932
rect 5601 -1934 5717 -1933
rect 5570 -1942 5638 -1934
rect 5417 -1944 5486 -1942
rect 5504 -1944 5638 -1942
rect 5381 -1948 5453 -1944
rect 5381 -1950 5506 -1948
rect 5381 -1954 5453 -1950
rect 5276 -1962 5327 -1954
rect 5374 -1958 5453 -1954
rect 5534 -1958 5638 -1944
rect 5667 -1942 5717 -1934
rect 5667 -1951 5683 -1942
rect 5374 -1962 5638 -1958
rect 5664 -1954 5683 -1951
rect 5690 -1954 5717 -1942
rect 5664 -1962 5717 -1954
rect 5292 -1970 5293 -1962
rect 5308 -1970 5321 -1962
rect 5292 -1978 5308 -1970
rect 5289 -1985 5308 -1982
rect 5289 -1994 5311 -1985
rect 5262 -2004 5311 -1994
rect 5262 -2010 5292 -2004
rect 5311 -2009 5316 -2004
rect 5234 -2026 5308 -2010
rect 5326 -2018 5356 -1962
rect 5391 -1972 5599 -1962
rect 5634 -1966 5679 -1962
rect 5682 -1963 5683 -1962
rect 5698 -1963 5711 -1962
rect 5558 -1976 5606 -1972
rect 5441 -1998 5471 -1989
rect 5534 -1996 5549 -1989
rect 5570 -1998 5606 -1976
rect 5417 -2002 5606 -1998
rect 5432 -2005 5606 -2002
rect 5425 -2008 5606 -2005
rect 5234 -2028 5247 -2026
rect 5262 -2028 5296 -2026
rect 5234 -2044 5308 -2028
rect 5335 -2032 5348 -2018
rect 5363 -2032 5379 -2016
rect 5425 -2021 5436 -2008
rect 5218 -2066 5219 -2050
rect 5234 -2066 5247 -2044
rect 5262 -2066 5292 -2044
rect 5335 -2048 5397 -2032
rect 5425 -2039 5436 -2023
rect 5441 -2028 5451 -2008
rect 5461 -2028 5475 -2008
rect 5478 -2021 5487 -2008
rect 5503 -2021 5512 -2008
rect 5441 -2039 5475 -2028
rect 5478 -2039 5487 -2023
rect 5503 -2039 5512 -2023
rect 5519 -2028 5529 -2008
rect 5539 -2028 5553 -2008
rect 5554 -2021 5565 -2008
rect 5519 -2039 5553 -2028
rect 5554 -2039 5565 -2023
rect 5611 -2032 5627 -2016
rect 5634 -2018 5664 -1966
rect 5698 -1970 5699 -1963
rect 5683 -1978 5699 -1970
rect 5670 -2010 5683 -1991
rect 5698 -2010 5728 -1994
rect 5670 -2026 5744 -2010
rect 5670 -2028 5683 -2026
rect 5698 -2028 5732 -2026
rect 5335 -2050 5348 -2048
rect 5363 -2050 5397 -2048
rect 5335 -2066 5397 -2050
rect 5441 -2055 5457 -2048
rect 5519 -2055 5549 -2044
rect 5597 -2048 5643 -2032
rect 5670 -2044 5744 -2028
rect 5597 -2050 5631 -2048
rect 5596 -2066 5643 -2050
rect 5670 -2066 5683 -2044
rect 5698 -2066 5728 -2044
rect 5755 -2066 5756 -2050
rect 5771 -2066 5784 -1906
rect 5814 -2010 5827 -1906
rect 5872 -1928 5873 -1918
rect 5888 -1928 5901 -1918
rect 5872 -1932 5901 -1928
rect 5906 -1932 5936 -1906
rect 5954 -1920 5970 -1918
rect 6042 -1920 6093 -1906
rect 6043 -1922 6107 -1920
rect 5954 -1932 5969 -1928
rect 5872 -1934 5969 -1932
rect 5856 -1942 5907 -1934
rect 5856 -1954 5881 -1942
rect 5888 -1954 5907 -1942
rect 5938 -1942 5988 -1934
rect 5938 -1950 5954 -1942
rect 5961 -1944 5988 -1942
rect 5997 -1942 6012 -1938
rect 6059 -1942 6091 -1922
rect 6150 -1934 6165 -1906
rect 6214 -1909 6244 -1906
rect 6214 -1912 6250 -1909
rect 6180 -1920 6196 -1918
rect 6181 -1932 6196 -1928
rect 6214 -1931 6253 -1912
rect 6272 -1918 6279 -1917
rect 6278 -1925 6279 -1918
rect 6262 -1928 6263 -1925
rect 6278 -1928 6291 -1925
rect 6214 -1932 6244 -1931
rect 6253 -1932 6259 -1931
rect 6262 -1932 6291 -1928
rect 6181 -1933 6291 -1932
rect 6181 -1934 6297 -1933
rect 6150 -1942 6218 -1934
rect 5997 -1944 6066 -1942
rect 6084 -1944 6218 -1942
rect 5961 -1948 6033 -1944
rect 5961 -1950 6086 -1948
rect 5961 -1954 6033 -1950
rect 5856 -1962 5907 -1954
rect 5954 -1958 6033 -1954
rect 6114 -1958 6218 -1944
rect 6247 -1942 6297 -1934
rect 6247 -1951 6263 -1942
rect 5954 -1962 6218 -1958
rect 6244 -1954 6263 -1951
rect 6270 -1954 6297 -1942
rect 6244 -1962 6297 -1954
rect 5872 -1970 5873 -1962
rect 5888 -1970 5901 -1962
rect 5872 -1978 5888 -1970
rect 5869 -1985 5888 -1982
rect 5869 -1994 5891 -1985
rect 5842 -2004 5891 -1994
rect 5842 -2010 5872 -2004
rect 5891 -2009 5896 -2004
rect 5814 -2026 5888 -2010
rect 5906 -2018 5936 -1962
rect 5971 -1972 6179 -1962
rect 6214 -1966 6259 -1962
rect 6262 -1963 6263 -1962
rect 6278 -1963 6291 -1962
rect 6138 -1976 6186 -1972
rect 6021 -1998 6051 -1989
rect 6114 -1996 6129 -1989
rect 6150 -1998 6186 -1976
rect 5997 -2002 6186 -1998
rect 6012 -2005 6186 -2002
rect 6005 -2008 6186 -2005
rect 5814 -2028 5827 -2026
rect 5842 -2028 5876 -2026
rect 5814 -2044 5888 -2028
rect 5915 -2032 5928 -2018
rect 5943 -2032 5959 -2016
rect 6005 -2021 6016 -2008
rect 5798 -2066 5799 -2050
rect 5814 -2066 5827 -2044
rect 5842 -2066 5872 -2044
rect 5915 -2048 5977 -2032
rect 6005 -2039 6016 -2023
rect 6021 -2028 6031 -2008
rect 6041 -2028 6055 -2008
rect 6058 -2021 6067 -2008
rect 6083 -2021 6092 -2008
rect 6021 -2039 6055 -2028
rect 6058 -2039 6067 -2023
rect 6083 -2039 6092 -2023
rect 6099 -2028 6109 -2008
rect 6119 -2028 6133 -2008
rect 6134 -2021 6145 -2008
rect 6099 -2039 6133 -2028
rect 6134 -2039 6145 -2023
rect 6191 -2032 6207 -2016
rect 6214 -2018 6244 -1966
rect 6278 -1970 6279 -1963
rect 6263 -1978 6279 -1970
rect 6250 -2010 6263 -1991
rect 6278 -2010 6308 -1994
rect 6250 -2026 6324 -2010
rect 6250 -2028 6263 -2026
rect 6278 -2028 6312 -2026
rect 5915 -2050 5928 -2048
rect 5943 -2050 5977 -2048
rect 5915 -2066 5977 -2050
rect 6021 -2055 6037 -2048
rect 6099 -2055 6129 -2044
rect 6177 -2048 6223 -2032
rect 6250 -2044 6324 -2028
rect 6177 -2050 6211 -2048
rect 6176 -2066 6223 -2050
rect 6250 -2066 6263 -2044
rect 6278 -2066 6308 -2044
rect 6335 -2066 6336 -2050
rect 6351 -2066 6364 -1906
rect 6394 -2010 6407 -1906
rect 6452 -1928 6453 -1918
rect 6468 -1928 6481 -1918
rect 6452 -1932 6481 -1928
rect 6486 -1932 6516 -1906
rect 6534 -1920 6550 -1918
rect 6622 -1920 6673 -1906
rect 6623 -1922 6687 -1920
rect 6534 -1932 6549 -1928
rect 6452 -1934 6549 -1932
rect 6436 -1942 6487 -1934
rect 6436 -1954 6461 -1942
rect 6468 -1954 6487 -1942
rect 6518 -1942 6568 -1934
rect 6518 -1950 6534 -1942
rect 6541 -1944 6568 -1942
rect 6577 -1942 6592 -1938
rect 6639 -1942 6671 -1922
rect 6730 -1934 6745 -1906
rect 6794 -1909 6824 -1906
rect 6794 -1912 6830 -1909
rect 6760 -1920 6776 -1918
rect 6761 -1932 6776 -1928
rect 6794 -1931 6833 -1912
rect 6852 -1918 6859 -1917
rect 6858 -1925 6859 -1918
rect 6842 -1928 6843 -1925
rect 6858 -1928 6871 -1925
rect 6794 -1932 6824 -1931
rect 6833 -1932 6839 -1931
rect 6842 -1932 6871 -1928
rect 6761 -1933 6871 -1932
rect 6761 -1934 6877 -1933
rect 6730 -1942 6798 -1934
rect 6577 -1944 6646 -1942
rect 6664 -1944 6798 -1942
rect 6541 -1948 6613 -1944
rect 6541 -1950 6666 -1948
rect 6541 -1954 6613 -1950
rect 6436 -1962 6487 -1954
rect 6534 -1958 6613 -1954
rect 6694 -1958 6798 -1944
rect 6827 -1942 6877 -1934
rect 6827 -1951 6843 -1942
rect 6534 -1962 6798 -1958
rect 6824 -1954 6843 -1951
rect 6850 -1954 6877 -1942
rect 6824 -1962 6877 -1954
rect 6452 -1970 6453 -1962
rect 6468 -1970 6481 -1962
rect 6452 -1978 6468 -1970
rect 6449 -1985 6468 -1982
rect 6449 -1994 6471 -1985
rect 6422 -2004 6471 -1994
rect 6422 -2010 6452 -2004
rect 6471 -2009 6476 -2004
rect 6394 -2026 6468 -2010
rect 6486 -2018 6516 -1962
rect 6551 -1972 6759 -1962
rect 6794 -1966 6839 -1962
rect 6842 -1963 6843 -1962
rect 6858 -1963 6871 -1962
rect 6718 -1976 6766 -1972
rect 6601 -1998 6631 -1989
rect 6694 -1996 6709 -1989
rect 6730 -1998 6766 -1976
rect 6577 -2002 6766 -1998
rect 6592 -2005 6766 -2002
rect 6585 -2008 6766 -2005
rect 6394 -2028 6407 -2026
rect 6422 -2028 6456 -2026
rect 6394 -2044 6468 -2028
rect 6495 -2032 6508 -2018
rect 6523 -2032 6539 -2016
rect 6585 -2021 6596 -2008
rect 6378 -2066 6379 -2050
rect 6394 -2066 6407 -2044
rect 6422 -2066 6452 -2044
rect 6495 -2048 6557 -2032
rect 6585 -2039 6596 -2023
rect 6601 -2028 6611 -2008
rect 6621 -2028 6635 -2008
rect 6638 -2021 6647 -2008
rect 6663 -2021 6672 -2008
rect 6601 -2039 6635 -2028
rect 6638 -2039 6647 -2023
rect 6663 -2039 6672 -2023
rect 6679 -2028 6689 -2008
rect 6699 -2028 6713 -2008
rect 6714 -2021 6725 -2008
rect 6679 -2039 6713 -2028
rect 6714 -2039 6725 -2023
rect 6771 -2032 6787 -2016
rect 6794 -2018 6824 -1966
rect 6858 -1970 6859 -1963
rect 6843 -1978 6859 -1970
rect 6830 -2010 6843 -1991
rect 6858 -2010 6888 -1994
rect 6830 -2026 6904 -2010
rect 6830 -2028 6843 -2026
rect 6858 -2028 6892 -2026
rect 6495 -2050 6508 -2048
rect 6523 -2050 6557 -2048
rect 6495 -2066 6557 -2050
rect 6601 -2055 6617 -2048
rect 6679 -2055 6709 -2044
rect 6757 -2048 6803 -2032
rect 6830 -2044 6904 -2028
rect 6757 -2050 6791 -2048
rect 6756 -2066 6803 -2050
rect 6830 -2066 6843 -2044
rect 6858 -2066 6888 -2044
rect 6915 -2066 6916 -2050
rect 6931 -2066 6944 -1906
rect -8 -2074 33 -2066
rect -8 -2100 7 -2074
rect 14 -2100 33 -2074
rect 97 -2078 159 -2066
rect 171 -2078 246 -2066
rect 304 -2078 379 -2066
rect 391 -2078 422 -2066
rect 428 -2078 463 -2066
rect 97 -2080 259 -2078
rect -8 -2108 33 -2100
rect 115 -2108 128 -2080
rect 143 -2082 158 -2080
rect 182 -2107 189 -2100
rect 192 -2108 259 -2080
rect 291 -2080 463 -2078
rect 261 -2102 289 -2098
rect 291 -2102 371 -2080
rect 392 -2082 407 -2080
rect 261 -2104 371 -2102
rect 261 -2108 289 -2104
rect 291 -2108 371 -2104
rect -2 -2118 -1 -2108
rect 14 -2118 27 -2108
rect 42 -2118 72 -2108
rect 115 -2118 158 -2108
rect 165 -2118 173 -2108
rect 192 -2116 195 -2108
rect 259 -2116 291 -2108
rect 192 -2118 358 -2116
rect 377 -2118 388 -2108
rect 392 -2118 422 -2108
rect 450 -2118 463 -2080
rect 535 -2074 570 -2066
rect 535 -2100 536 -2074
rect 543 -2100 570 -2074
rect 535 -2108 570 -2100
rect 572 -2074 613 -2066
rect 572 -2100 587 -2074
rect 594 -2100 613 -2074
rect 677 -2078 739 -2066
rect 751 -2078 826 -2066
rect 884 -2078 959 -2066
rect 971 -2078 1002 -2066
rect 1008 -2078 1043 -2066
rect 677 -2080 839 -2078
rect 572 -2108 613 -2100
rect 695 -2108 708 -2080
rect 723 -2082 738 -2080
rect 762 -2107 769 -2100
rect 772 -2108 839 -2080
rect 871 -2080 1043 -2078
rect 841 -2102 869 -2098
rect 871 -2102 951 -2080
rect 972 -2082 987 -2080
rect 841 -2104 951 -2102
rect 841 -2108 869 -2104
rect 871 -2108 951 -2104
rect 478 -2118 508 -2108
rect 535 -2118 536 -2108
rect 551 -2118 564 -2108
rect 578 -2118 579 -2108
rect 594 -2118 607 -2108
rect 622 -2118 652 -2108
rect 695 -2118 738 -2108
rect 745 -2118 753 -2108
rect 772 -2116 775 -2108
rect 839 -2116 871 -2108
rect 772 -2118 938 -2116
rect 957 -2118 968 -2108
rect 972 -2118 1002 -2108
rect 1030 -2118 1043 -2080
rect 1115 -2074 1150 -2066
rect 1115 -2100 1116 -2074
rect 1123 -2100 1150 -2074
rect 1115 -2108 1150 -2100
rect 1152 -2074 1193 -2066
rect 1152 -2100 1167 -2074
rect 1174 -2100 1193 -2074
rect 1257 -2078 1319 -2066
rect 1331 -2078 1406 -2066
rect 1464 -2078 1539 -2066
rect 3435 -2074 3470 -2066
rect 1257 -2080 1419 -2078
rect 1152 -2108 1193 -2100
rect 1275 -2108 1288 -2080
rect 1303 -2082 1318 -2080
rect 1342 -2107 1349 -2100
rect 1352 -2108 1419 -2080
rect 1451 -2080 1551 -2078
rect 1421 -2102 1449 -2098
rect 1451 -2102 1531 -2080
rect 1421 -2104 1531 -2102
rect 1421 -2108 1449 -2104
rect 1451 -2108 1531 -2104
rect 3435 -2100 3436 -2074
rect 3443 -2100 3470 -2074
rect 3435 -2108 3470 -2100
rect 3472 -2074 3513 -2066
rect 3472 -2100 3487 -2074
rect 3494 -2100 3513 -2074
rect 3577 -2078 3639 -2066
rect 3651 -2078 3726 -2066
rect 3784 -2078 3859 -2066
rect 3871 -2078 3902 -2066
rect 3908 -2078 3943 -2066
rect 3577 -2080 3739 -2078
rect 3472 -2108 3513 -2100
rect 3595 -2108 3608 -2080
rect 3623 -2082 3638 -2080
rect 3662 -2107 3669 -2100
rect 3672 -2108 3739 -2080
rect 3771 -2080 3943 -2078
rect 3741 -2102 3769 -2098
rect 3771 -2102 3851 -2080
rect 3872 -2082 3887 -2080
rect 3741 -2104 3851 -2102
rect 3741 -2108 3769 -2104
rect 3771 -2108 3851 -2104
rect 1058 -2118 1088 -2108
rect 1115 -2118 1116 -2108
rect 1131 -2118 1144 -2108
rect 1158 -2118 1159 -2108
rect 1174 -2118 1187 -2108
rect 1202 -2118 1232 -2108
rect 1275 -2118 1318 -2108
rect 1325 -2118 1333 -2108
rect 1352 -2116 1355 -2108
rect 1419 -2116 1451 -2108
rect 1352 -2118 1518 -2116
rect 1537 -2118 1548 -2108
rect 3379 -2118 3408 -2108
rect 3435 -2118 3436 -2108
rect 3451 -2118 3464 -2108
rect 3478 -2118 3479 -2108
rect 3494 -2118 3507 -2108
rect 3522 -2118 3552 -2108
rect 3595 -2118 3638 -2108
rect 3645 -2118 3653 -2108
rect 3672 -2116 3675 -2108
rect 3739 -2116 3771 -2108
rect 3672 -2118 3838 -2116
rect 3857 -2118 3868 -2108
rect 3872 -2118 3902 -2108
rect 3930 -2118 3943 -2080
rect 4015 -2074 4050 -2066
rect 4015 -2100 4016 -2074
rect 4023 -2100 4050 -2074
rect 4015 -2108 4050 -2100
rect 4052 -2074 4093 -2066
rect 4052 -2100 4067 -2074
rect 4074 -2100 4093 -2074
rect 4157 -2078 4219 -2066
rect 4231 -2078 4306 -2066
rect 4364 -2078 4439 -2066
rect 4451 -2078 4482 -2066
rect 4488 -2078 4523 -2066
rect 4157 -2080 4319 -2078
rect 4052 -2108 4093 -2100
rect 4175 -2108 4188 -2080
rect 4203 -2082 4218 -2080
rect 4242 -2107 4249 -2100
rect 4252 -2108 4319 -2080
rect 4351 -2080 4523 -2078
rect 4321 -2102 4349 -2098
rect 4351 -2102 4431 -2080
rect 4452 -2082 4467 -2080
rect 4321 -2104 4431 -2102
rect 4321 -2108 4349 -2104
rect 4351 -2108 4431 -2104
rect 3958 -2118 3988 -2108
rect 4015 -2118 4016 -2108
rect 4031 -2118 4044 -2108
rect 4058 -2118 4059 -2108
rect 4074 -2118 4087 -2108
rect 4102 -2118 4132 -2108
rect 4175 -2118 4218 -2108
rect 4225 -2118 4233 -2108
rect 4252 -2116 4255 -2108
rect 4319 -2116 4351 -2108
rect 4252 -2118 4418 -2116
rect 4437 -2118 4448 -2108
rect 4452 -2118 4482 -2108
rect 4510 -2118 4523 -2080
rect 4595 -2074 4630 -2066
rect 4595 -2100 4596 -2074
rect 4603 -2100 4630 -2074
rect 4595 -2108 4630 -2100
rect 4632 -2074 4673 -2066
rect 4632 -2100 4647 -2074
rect 4654 -2100 4673 -2074
rect 4737 -2078 4799 -2066
rect 4811 -2078 4886 -2066
rect 4944 -2078 5019 -2066
rect 5031 -2078 5062 -2066
rect 5068 -2078 5103 -2066
rect 4737 -2080 4899 -2078
rect 4632 -2108 4673 -2100
rect 4755 -2108 4768 -2080
rect 4783 -2082 4798 -2080
rect 4832 -2098 4899 -2080
rect 4931 -2080 5103 -2078
rect 4931 -2098 5011 -2080
rect 5032 -2082 5047 -2080
rect 4822 -2107 4829 -2100
rect 4832 -2108 5011 -2098
rect 4538 -2118 4568 -2108
rect 4595 -2118 4596 -2108
rect 4611 -2118 4624 -2108
rect 4638 -2118 4639 -2108
rect 4654 -2118 4667 -2108
rect 4682 -2118 4712 -2108
rect 4755 -2118 4798 -2108
rect 4805 -2118 4813 -2108
rect 4832 -2116 4835 -2108
rect 4899 -2116 4931 -2108
rect 4832 -2118 4998 -2116
rect 5017 -2118 5028 -2108
rect 5032 -2118 5062 -2108
rect 5090 -2118 5103 -2080
rect 5175 -2074 5210 -2066
rect 5175 -2100 5176 -2074
rect 5183 -2100 5210 -2074
rect 5175 -2108 5210 -2100
rect 5212 -2074 5253 -2066
rect 5212 -2100 5227 -2074
rect 5234 -2100 5253 -2074
rect 5317 -2078 5379 -2066
rect 5391 -2078 5466 -2066
rect 5524 -2078 5599 -2066
rect 5611 -2078 5642 -2066
rect 5648 -2078 5683 -2066
rect 5317 -2080 5479 -2078
rect 5212 -2108 5253 -2100
rect 5335 -2108 5348 -2080
rect 5363 -2082 5378 -2080
rect 5412 -2098 5479 -2080
rect 5511 -2080 5683 -2078
rect 5511 -2098 5591 -2080
rect 5612 -2082 5627 -2080
rect 5402 -2107 5409 -2100
rect 5412 -2108 5591 -2098
rect 5118 -2118 5148 -2108
rect 5175 -2118 5176 -2108
rect 5191 -2118 5204 -2108
rect 5218 -2118 5219 -2108
rect 5234 -2118 5247 -2108
rect 5262 -2118 5292 -2108
rect 5335 -2118 5378 -2108
rect 5385 -2118 5393 -2108
rect 5412 -2116 5415 -2108
rect 5479 -2116 5511 -2108
rect 5412 -2118 5578 -2116
rect 5597 -2118 5608 -2108
rect 5612 -2118 5642 -2108
rect 5670 -2118 5683 -2080
rect 5755 -2074 5790 -2066
rect 5755 -2100 5756 -2074
rect 5763 -2100 5790 -2074
rect 5755 -2108 5790 -2100
rect 5792 -2074 5833 -2066
rect 5792 -2100 5807 -2074
rect 5814 -2100 5833 -2074
rect 5897 -2078 5959 -2066
rect 5971 -2078 6046 -2066
rect 6104 -2078 6179 -2066
rect 6191 -2078 6222 -2066
rect 6228 -2078 6263 -2066
rect 5897 -2080 6059 -2078
rect 5792 -2108 5833 -2100
rect 5915 -2108 5928 -2080
rect 5943 -2082 5958 -2080
rect 5992 -2098 6059 -2080
rect 6091 -2080 6263 -2078
rect 6091 -2098 6171 -2080
rect 6192 -2082 6207 -2080
rect 5982 -2107 5989 -2100
rect 5992 -2108 6171 -2098
rect 5698 -2118 5728 -2108
rect 5755 -2118 5756 -2108
rect 5771 -2118 5784 -2108
rect 5798 -2118 5799 -2108
rect 5814 -2118 5827 -2108
rect 5842 -2118 5872 -2108
rect 5915 -2118 5958 -2108
rect 5965 -2118 5973 -2108
rect 5992 -2116 5995 -2108
rect 6059 -2116 6091 -2108
rect 5992 -2118 6158 -2116
rect 6177 -2118 6188 -2108
rect 6192 -2118 6222 -2108
rect 6250 -2118 6263 -2080
rect 6335 -2074 6370 -2066
rect 6335 -2100 6336 -2074
rect 6343 -2100 6370 -2074
rect 6335 -2108 6370 -2100
rect 6372 -2074 6413 -2066
rect 6372 -2100 6387 -2074
rect 6394 -2100 6413 -2074
rect 6477 -2078 6539 -2066
rect 6551 -2078 6626 -2066
rect 6684 -2078 6759 -2066
rect 6771 -2078 6802 -2066
rect 6808 -2078 6843 -2066
rect 6477 -2080 6639 -2078
rect 6372 -2108 6413 -2100
rect 6495 -2108 6508 -2080
rect 6523 -2082 6538 -2080
rect 6572 -2098 6639 -2080
rect 6671 -2080 6843 -2078
rect 6671 -2098 6751 -2080
rect 6772 -2082 6787 -2080
rect 6562 -2107 6569 -2100
rect 6572 -2108 6751 -2098
rect 6278 -2118 6308 -2108
rect 6335 -2118 6336 -2108
rect 6351 -2118 6364 -2108
rect 6378 -2118 6379 -2108
rect 6394 -2118 6407 -2108
rect 6422 -2118 6452 -2108
rect 6495 -2118 6538 -2108
rect 6545 -2118 6553 -2108
rect 6572 -2116 6575 -2108
rect 6639 -2116 6671 -2108
rect 6572 -2118 6738 -2116
rect 6757 -2118 6768 -2108
rect 6772 -2118 6802 -2108
rect 6830 -2118 6843 -2080
rect 6915 -2074 6950 -2066
rect 6915 -2100 6916 -2074
rect 6923 -2100 6950 -2074
rect 6915 -2108 6950 -2100
rect 6858 -2118 6888 -2108
rect 6915 -2118 6916 -2108
rect 6931 -2118 6944 -2108
rect -2 -2124 1551 -2118
rect -1 -2132 1551 -2124
rect 3379 -2132 6944 -2118
rect 14 -2146 27 -2132
rect 42 -2150 72 -2132
rect 115 -2146 128 -2132
rect 165 -2145 173 -2132
rect 206 -2145 344 -2132
rect 377 -2145 385 -2132
rect 242 -2146 293 -2145
rect 450 -2146 463 -2132
rect 243 -2148 307 -2146
rect 478 -2150 508 -2132
rect 551 -2146 564 -2132
rect 594 -2146 607 -2132
rect 622 -2150 652 -2132
rect 695 -2146 708 -2132
rect 745 -2145 753 -2132
rect 786 -2145 924 -2132
rect 957 -2145 965 -2132
rect 822 -2146 873 -2145
rect 1030 -2146 1043 -2132
rect 823 -2148 887 -2146
rect 1058 -2150 1088 -2132
rect 1131 -2146 1144 -2132
rect 1174 -2146 1187 -2132
rect 1202 -2150 1232 -2132
rect 1275 -2146 1288 -2132
rect 1325 -2145 1333 -2132
rect 1366 -2145 1504 -2132
rect 1537 -2145 1545 -2132
rect 1402 -2146 1453 -2145
rect 1403 -2148 1467 -2146
rect 3379 -2150 3408 -2132
rect 3451 -2146 3464 -2132
rect 3494 -2146 3507 -2132
rect 3522 -2150 3552 -2132
rect 3595 -2146 3608 -2132
rect 3645 -2145 3653 -2132
rect 3686 -2145 3824 -2132
rect 3857 -2145 3865 -2132
rect 3722 -2146 3773 -2145
rect 3930 -2146 3943 -2132
rect 3723 -2148 3787 -2146
rect 3958 -2150 3988 -2132
rect 4031 -2146 4044 -2132
rect 4074 -2146 4087 -2132
rect 4102 -2150 4132 -2132
rect 4175 -2146 4188 -2132
rect 4225 -2145 4233 -2132
rect 4266 -2145 4404 -2132
rect 4437 -2145 4445 -2132
rect 4302 -2146 4353 -2145
rect 4510 -2146 4523 -2132
rect 4303 -2148 4367 -2146
rect 4538 -2150 4568 -2132
rect 4611 -2146 4624 -2132
rect 4654 -2146 4667 -2132
rect 4682 -2150 4712 -2132
rect 4755 -2146 4768 -2132
rect 4805 -2145 4813 -2132
rect 4846 -2145 4984 -2132
rect 5017 -2145 5025 -2132
rect 4882 -2146 4933 -2145
rect 5090 -2146 5103 -2132
rect 4899 -2148 4931 -2146
rect 5118 -2150 5148 -2132
rect 5191 -2146 5204 -2132
rect 5234 -2146 5247 -2132
rect 5262 -2150 5292 -2132
rect 5335 -2146 5348 -2132
rect 5385 -2145 5393 -2132
rect 5426 -2145 5564 -2132
rect 5597 -2145 5605 -2132
rect 5462 -2146 5513 -2145
rect 5670 -2146 5683 -2132
rect 5479 -2148 5511 -2146
rect 5698 -2150 5728 -2132
rect 5771 -2146 5784 -2132
rect 5814 -2146 5827 -2132
rect 5842 -2150 5872 -2132
rect 5915 -2146 5928 -2132
rect 5965 -2145 5973 -2132
rect 6006 -2145 6144 -2132
rect 6177 -2145 6185 -2132
rect 6042 -2146 6093 -2145
rect 6250 -2146 6263 -2132
rect 6059 -2148 6091 -2146
rect 6278 -2150 6308 -2132
rect 6351 -2146 6364 -2132
rect 6394 -2146 6407 -2132
rect 6422 -2150 6452 -2132
rect 6495 -2146 6508 -2132
rect 6545 -2145 6553 -2132
rect 6586 -2145 6724 -2132
rect 6757 -2145 6765 -2132
rect 6622 -2146 6673 -2145
rect 6830 -2146 6843 -2132
rect 6639 -2148 6671 -2146
rect 6858 -2150 6888 -2132
rect 6931 -2146 6944 -2132
<< nwell >>
rect 197 2048 350 2144
rect 777 2048 930 2144
rect 1357 2048 1510 2144
rect 1937 2048 2090 2144
rect 2517 2048 2670 2144
rect 3097 2048 3250 2144
rect 3677 2048 3830 2144
rect 4257 2048 4410 2144
rect 197 1778 350 1874
rect 777 1778 930 1874
rect 1357 1778 1510 1874
rect 1937 1778 2090 1874
rect 2517 1778 2670 1874
rect 3097 1778 3250 1874
rect 3677 1778 3830 1874
rect 4257 1778 4410 1874
rect 197 1508 350 1604
rect 777 1508 930 1604
rect 1357 1508 1510 1604
rect 1937 1508 2090 1604
rect 2517 1508 2670 1604
rect 3097 1508 3250 1604
rect 3677 1508 3830 1604
rect 4257 1508 4410 1604
rect 197 1238 350 1334
rect 777 1238 930 1334
rect 1357 1238 1510 1334
rect 1937 1238 2090 1334
rect 2517 1238 2670 1334
rect 3097 1238 3250 1334
rect 3677 1238 3830 1334
rect 4257 1238 4410 1334
rect 197 968 350 1064
rect 777 968 930 1064
rect 1357 968 1510 1064
rect 1937 968 2090 1064
rect 2517 968 2670 1064
rect 3097 968 3250 1064
rect 3677 968 3830 1064
rect 4257 968 4410 1064
rect 197 698 350 794
rect 777 698 930 794
rect 1357 698 1510 794
rect 1937 698 2090 794
rect 2517 698 2670 794
rect 3097 698 3250 794
rect 3677 698 3830 794
rect 4257 698 4410 794
rect 197 428 350 524
rect 777 428 930 524
rect 1357 428 1510 524
rect 1937 428 2090 524
rect 2517 428 2670 524
rect 3097 428 3250 524
rect 3677 428 3830 524
rect 4257 428 4410 524
rect 197 158 350 254
rect 777 158 930 254
rect 1357 158 1510 254
rect 1937 158 2090 254
rect 2517 158 2670 254
rect 3097 158 3250 254
rect 3677 158 3830 254
rect 4257 158 4410 254
rect 197 -112 350 -16
rect 777 -112 930 -16
rect 1357 -112 1510 -16
rect 1937 -112 2090 -16
rect 2517 -112 2670 -16
rect 3097 -112 3250 -16
rect 3677 -112 3830 -16
rect 4257 -112 4410 -16
rect 197 -382 350 -286
rect 777 -382 930 -286
rect 1357 -382 1510 -286
rect 1937 -382 2090 -286
rect 2517 -382 2670 -286
rect 3097 -382 3250 -286
rect 3677 -382 3830 -286
rect 4257 -382 4410 -286
rect 197 -652 350 -556
rect 777 -652 930 -556
rect 1357 -652 1510 -556
rect 1937 -652 2090 -556
rect 2517 -652 2670 -556
rect 3097 -652 3250 -556
rect 3677 -652 3830 -556
rect 4257 -652 4410 -556
rect 197 -922 350 -826
rect 777 -922 930 -826
rect 1357 -922 1510 -826
rect 1937 -922 2090 -826
rect 2517 -922 2670 -826
rect 3097 -922 3250 -826
rect 3677 -922 3830 -826
rect 4257 -922 4410 -826
rect 197 -1192 350 -1096
rect 777 -1192 930 -1096
rect 1357 -1192 1510 -1096
rect 1937 -1192 2090 -1096
rect 2517 -1192 2670 -1096
rect 3097 -1192 3250 -1096
rect 3677 -1192 3830 -1096
rect 4257 -1192 4410 -1096
rect 197 -1462 350 -1366
rect 777 -1462 930 -1366
rect 1357 -1462 1510 -1366
rect 1937 -1462 2090 -1366
rect 2517 -1462 2670 -1366
rect 3097 -1462 3250 -1366
rect 3677 -1462 3830 -1366
rect 4257 -1462 4410 -1366
rect 197 -1732 350 -1636
rect 777 -1732 930 -1636
rect 1357 -1732 1510 -1636
rect 1937 -1732 2090 -1636
rect 2517 -1732 2670 -1636
rect 3097 -1732 3250 -1636
rect 3677 -1732 3830 -1636
rect 4257 -1732 4410 -1636
rect 197 -2002 350 -1906
rect 777 -2002 930 -1906
rect 1357 -2002 1510 -1906
rect 1937 -2002 2090 -1906
rect 2517 -2002 2670 -1906
rect 3097 -2002 3250 -1906
rect 3677 -2002 3830 -1906
rect 4257 -2002 4410 -1906
rect 4837 2048 4990 2144
rect 5417 2048 5570 2144
rect 4837 1778 4990 1874
rect 5417 1778 5570 1874
rect 4837 1508 4990 1604
rect 5417 1508 5570 1604
rect 4837 1238 4990 1334
rect 5417 1238 5570 1334
rect 4837 968 4990 1064
rect 5417 968 5570 1064
rect 4837 698 4990 794
rect 5417 698 5570 794
rect 4837 428 4990 524
rect 5417 428 5570 524
rect 4837 158 4990 254
rect 5417 158 5570 254
rect 4837 -112 4990 -16
rect 5417 -112 5570 -16
rect 4837 -382 4990 -286
rect 5417 -382 5570 -286
rect 4837 -652 4990 -556
rect 5417 -652 5570 -556
rect 4837 -922 4990 -826
rect 5417 -922 5570 -826
rect 4837 -1192 4990 -1096
rect 5417 -1192 5570 -1096
rect 4837 -1462 4990 -1366
rect 5417 -1462 5570 -1366
rect 4837 -1732 4990 -1636
rect 5417 -1732 5570 -1636
rect 4837 -2002 4990 -1906
rect 5417 -2002 5570 -1906
rect 5997 2048 6150 2144
rect 6577 2048 6730 2144
rect 5997 1778 6150 1874
rect 6577 1778 6730 1874
rect 5997 1508 6150 1604
rect 6577 1508 6730 1604
rect 5997 1238 6150 1334
rect 6577 1238 6730 1334
rect 5997 968 6150 1064
rect 6577 968 6730 1064
rect 5997 698 6150 794
rect 6577 698 6730 794
rect 5997 428 6150 524
rect 6577 428 6730 524
rect 5997 158 6150 254
rect 6577 158 6730 254
rect 5997 -112 6150 -16
rect 6577 -112 6730 -16
rect 5997 -382 6150 -286
rect 6577 -382 6730 -286
rect 5997 -652 6150 -556
rect 6577 -652 6730 -556
rect 5997 -922 6150 -826
rect 6577 -922 6730 -826
rect 5997 -1192 6150 -1096
rect 6577 -1192 6730 -1096
rect 5997 -1462 6150 -1366
rect 6577 -1462 6730 -1366
rect 5997 -1732 6150 -1636
rect 6577 -1732 6730 -1636
rect 5997 -2002 6150 -1906
rect 6577 -2002 6730 -1906
<< pwell >>
rect -1 2002 169 2174
rect 381 2002 749 2174
rect 961 2002 1329 2174
rect 1541 2002 1909 2174
rect 2121 2002 2489 2174
rect 2701 2002 3069 2174
rect 3281 2002 3649 2174
rect 3861 2002 4229 2174
rect 4441 2002 4611 2174
rect -1 1904 4611 2002
rect -1 1732 169 1904
rect 381 1732 749 1904
rect 961 1732 1329 1904
rect 1541 1732 1909 1904
rect 2121 1732 2489 1904
rect 2701 1732 3069 1904
rect 3281 1732 3649 1904
rect 3861 1732 4229 1904
rect 4441 1732 4611 1904
rect -1 1634 4611 1732
rect -1 1462 169 1634
rect 381 1462 749 1634
rect 961 1462 1329 1634
rect 1541 1462 1909 1634
rect 2121 1462 2489 1634
rect 2701 1462 3069 1634
rect 3281 1462 3649 1634
rect 3861 1462 4229 1634
rect 4441 1462 4611 1634
rect -1 1364 4611 1462
rect -1 1192 169 1364
rect 381 1192 749 1364
rect 961 1192 1329 1364
rect 1541 1192 1909 1364
rect 2121 1192 2489 1364
rect 2701 1192 3069 1364
rect 3281 1192 3649 1364
rect 3861 1192 4229 1364
rect 4441 1192 4611 1364
rect -1 1094 4611 1192
rect -1 922 169 1094
rect 381 922 749 1094
rect 961 922 1329 1094
rect 1541 922 1909 1094
rect 2121 922 2489 1094
rect 2701 922 3069 1094
rect 3281 922 3649 1094
rect 3861 922 4229 1094
rect 4441 922 4611 1094
rect -1 824 4611 922
rect -1 652 169 824
rect 381 652 749 824
rect 961 652 1329 824
rect 1541 652 1909 824
rect 2121 652 2489 824
rect 2701 652 3069 824
rect 3281 652 3649 824
rect 3861 652 4229 824
rect 4441 652 4611 824
rect -1 554 4611 652
rect -1 382 169 554
rect 381 382 749 554
rect 961 382 1329 554
rect 1541 382 1909 554
rect 2121 382 2489 554
rect 2701 382 3069 554
rect 3281 382 3649 554
rect 3861 382 4229 554
rect 4441 382 4611 554
rect -1 284 4611 382
rect -1 112 169 284
rect 381 112 749 284
rect 961 112 1329 284
rect 1541 112 1909 284
rect 2121 112 2489 284
rect 2701 112 3069 284
rect 3281 112 3649 284
rect 3861 112 4229 284
rect 4441 112 4611 284
rect -1 14 4611 112
rect -1 -158 169 14
rect 381 -158 749 14
rect 961 -158 1329 14
rect 1541 -158 1909 14
rect 2121 -158 2489 14
rect 2701 -158 3069 14
rect 3281 -158 3649 14
rect 3861 -158 4229 14
rect 4441 -158 4611 14
rect -1 -256 4611 -158
rect -1 -428 169 -256
rect 381 -428 749 -256
rect 961 -428 1329 -256
rect 1541 -428 1909 -256
rect 2121 -428 2489 -256
rect 2701 -428 3069 -256
rect 3281 -428 3649 -256
rect 3861 -428 4229 -256
rect 4441 -428 4611 -256
rect -1 -526 4611 -428
rect -1 -698 169 -526
rect 381 -698 749 -526
rect 961 -698 1329 -526
rect 1541 -698 1909 -526
rect 2121 -698 2489 -526
rect 2701 -698 3069 -526
rect 3281 -698 3649 -526
rect 3861 -698 4229 -526
rect 4441 -698 4611 -526
rect -1 -796 4611 -698
rect -1 -968 169 -796
rect 381 -968 749 -796
rect 961 -968 1329 -796
rect 1541 -968 1909 -796
rect 2121 -968 2489 -796
rect 2701 -968 3069 -796
rect 3281 -968 3649 -796
rect 3861 -968 4229 -796
rect 4441 -968 4611 -796
rect -1 -1066 4611 -968
rect -1 -1238 169 -1066
rect 381 -1238 749 -1066
rect 961 -1238 1329 -1066
rect 1541 -1238 1909 -1066
rect 2121 -1238 2489 -1066
rect 2701 -1238 3069 -1066
rect 3281 -1238 3649 -1066
rect 3861 -1238 4229 -1066
rect 4441 -1238 4611 -1066
rect -1 -1336 4611 -1238
rect -1 -1508 169 -1336
rect 381 -1508 749 -1336
rect 961 -1508 1329 -1336
rect 1541 -1508 1909 -1336
rect 2121 -1508 2489 -1336
rect 2701 -1508 3069 -1336
rect 3281 -1508 3649 -1336
rect 3861 -1508 4229 -1336
rect 4441 -1508 4611 -1336
rect -1 -1606 4611 -1508
rect -1 -1778 169 -1606
rect 381 -1778 749 -1606
rect 961 -1778 1329 -1606
rect 1541 -1778 1909 -1606
rect 2121 -1778 2489 -1606
rect 2701 -1778 3069 -1606
rect 3281 -1778 3649 -1606
rect 3861 -1778 4229 -1606
rect 4441 -1778 4611 -1606
rect -1 -1876 4611 -1778
rect -1 -2048 169 -1876
rect 381 -2048 749 -1876
rect 961 -2048 1329 -1876
rect 1541 -2048 1909 -1876
rect 2121 -2048 2489 -1876
rect 2701 -2048 3069 -1876
rect 3281 -2048 3649 -1876
rect 3861 -2048 4229 -1876
rect 4441 -2048 4611 -1876
rect -1 -2146 4611 -2048
rect 4639 2002 4809 2174
rect 5021 2002 5389 2174
rect 5601 2002 5771 2174
rect 4639 1904 5771 2002
rect 4639 1732 4809 1904
rect 5021 1732 5389 1904
rect 5601 1732 5771 1904
rect 4639 1634 5771 1732
rect 4639 1462 4809 1634
rect 5021 1462 5389 1634
rect 5601 1462 5771 1634
rect 4639 1364 5771 1462
rect 4639 1192 4809 1364
rect 5021 1192 5389 1364
rect 5601 1192 5771 1364
rect 4639 1094 5771 1192
rect 4639 922 4809 1094
rect 5021 922 5389 1094
rect 5601 922 5771 1094
rect 4639 824 5771 922
rect 4639 652 4809 824
rect 5021 652 5389 824
rect 5601 652 5771 824
rect 4639 554 5771 652
rect 4639 382 4809 554
rect 5021 382 5389 554
rect 5601 382 5771 554
rect 4639 284 5771 382
rect 4639 112 4809 284
rect 5021 112 5389 284
rect 5601 112 5771 284
rect 4639 14 5771 112
rect 4639 -158 4809 14
rect 5021 -158 5389 14
rect 5601 -158 5771 14
rect 4639 -256 5771 -158
rect 4639 -428 4809 -256
rect 5021 -428 5389 -256
rect 5601 -428 5771 -256
rect 4639 -526 5771 -428
rect 4639 -698 4809 -526
rect 5021 -698 5389 -526
rect 5601 -698 5771 -526
rect 4639 -796 5771 -698
rect 4639 -968 4809 -796
rect 5021 -968 5389 -796
rect 5601 -968 5771 -796
rect 4639 -1066 5771 -968
rect 4639 -1238 4809 -1066
rect 5021 -1238 5389 -1066
rect 5601 -1238 5771 -1066
rect 4639 -1336 5771 -1238
rect 4639 -1508 4809 -1336
rect 5021 -1508 5389 -1336
rect 5601 -1508 5771 -1336
rect 4639 -1606 5771 -1508
rect 4639 -1778 4809 -1606
rect 5021 -1778 5389 -1606
rect 5601 -1778 5771 -1606
rect 4639 -1876 5771 -1778
rect 4639 -2048 4809 -1876
rect 5021 -2048 5389 -1876
rect 5601 -2048 5771 -1876
rect 4639 -2146 5771 -2048
rect 5799 2002 5969 2174
rect 6181 2002 6549 2174
rect 6761 2002 6931 2174
rect 5799 1904 6931 2002
rect 5799 1732 5969 1904
rect 6181 1732 6549 1904
rect 6761 1732 6931 1904
rect 5799 1634 6931 1732
rect 5799 1462 5969 1634
rect 6181 1462 6549 1634
rect 6761 1462 6931 1634
rect 5799 1364 6931 1462
rect 5799 1192 5969 1364
rect 6181 1192 6549 1364
rect 6761 1192 6931 1364
rect 5799 1094 6931 1192
rect 5799 922 5969 1094
rect 6181 922 6549 1094
rect 6761 922 6931 1094
rect 5799 824 6931 922
rect 5799 652 5969 824
rect 6181 652 6549 824
rect 6761 652 6931 824
rect 5799 554 6931 652
rect 5799 382 5969 554
rect 6181 382 6549 554
rect 6761 382 6931 554
rect 5799 284 6931 382
rect 5799 112 5969 284
rect 6181 112 6549 284
rect 6761 112 6931 284
rect 5799 14 6931 112
rect 5799 -158 5969 14
rect 6181 -158 6549 14
rect 6761 -158 6931 14
rect 5799 -256 6931 -158
rect 5799 -428 5969 -256
rect 6181 -428 6549 -256
rect 6761 -428 6931 -256
rect 5799 -526 6931 -428
rect 5799 -698 5969 -526
rect 6181 -698 6549 -526
rect 6761 -698 6931 -526
rect 5799 -796 6931 -698
rect 5799 -968 5969 -796
rect 6181 -968 6549 -796
rect 6761 -968 6931 -796
rect 5799 -1066 6931 -968
rect 5799 -1238 5969 -1066
rect 6181 -1238 6549 -1066
rect 6761 -1238 6931 -1066
rect 5799 -1336 6931 -1238
rect 5799 -1508 5969 -1336
rect 6181 -1508 6549 -1336
rect 6761 -1508 6931 -1336
rect 5799 -1606 6931 -1508
rect 5799 -1778 5969 -1606
rect 6181 -1778 6549 -1606
rect 6761 -1778 6931 -1606
rect 5799 -1876 6931 -1778
rect 5799 -2048 5969 -1876
rect 6181 -2048 6549 -1876
rect 6761 -2048 6931 -1876
rect 5799 -2146 6931 -2048
<< nmos >>
rect 106 2088 136 2116
rect 414 2088 444 2116
rect 686 2088 716 2116
rect 994 2088 1024 2116
rect 1266 2088 1296 2116
rect 1574 2088 1604 2116
rect 1846 2088 1876 2116
rect 2154 2088 2184 2116
rect 2426 2088 2456 2116
rect 2734 2088 2764 2116
rect 3006 2088 3036 2116
rect 3314 2088 3344 2116
rect 3586 2088 3616 2116
rect 3894 2088 3924 2116
rect 4166 2088 4196 2116
rect 4474 2088 4504 2116
rect 4746 2088 4776 2116
rect 5054 2088 5084 2116
rect 5326 2088 5356 2116
rect 5634 2088 5664 2116
rect 5906 2088 5936 2116
rect 6214 2088 6244 2116
rect 6486 2088 6516 2116
rect 6794 2088 6824 2116
rect 42 1942 72 1984
rect 478 1942 508 1984
rect 622 1942 652 1984
rect 1058 1942 1088 1984
rect 1202 1942 1232 1984
rect 1638 1942 1668 1984
rect 1782 1942 1812 1984
rect 2218 1942 2248 1984
rect 2362 1942 2392 1984
rect 2798 1942 2828 1984
rect 2942 1942 2972 1984
rect 3378 1942 3408 1984
rect 3522 1942 3552 1984
rect 3958 1942 3988 1984
rect 4102 1942 4132 1984
rect 4538 1942 4568 1984
rect 4682 1942 4712 1984
rect 5118 1942 5148 1984
rect 5262 1942 5292 1984
rect 5698 1942 5728 1984
rect 5842 1942 5872 1984
rect 6278 1942 6308 1984
rect 6422 1942 6452 1984
rect 6858 1942 6888 1984
rect 106 1818 136 1846
rect 414 1818 444 1846
rect 686 1818 716 1846
rect 994 1818 1024 1846
rect 1266 1818 1296 1846
rect 1574 1818 1604 1846
rect 1846 1818 1876 1846
rect 2154 1818 2184 1846
rect 2426 1818 2456 1846
rect 2734 1818 2764 1846
rect 3006 1818 3036 1846
rect 3314 1818 3344 1846
rect 3586 1818 3616 1846
rect 3894 1818 3924 1846
rect 4166 1818 4196 1846
rect 4474 1818 4504 1846
rect 4746 1818 4776 1846
rect 5054 1818 5084 1846
rect 5326 1818 5356 1846
rect 5634 1818 5664 1846
rect 5906 1818 5936 1846
rect 6214 1818 6244 1846
rect 6486 1818 6516 1846
rect 6794 1818 6824 1846
rect 42 1672 72 1714
rect 478 1672 508 1714
rect 622 1672 652 1714
rect 1058 1672 1088 1714
rect 1202 1672 1232 1714
rect 1638 1672 1668 1714
rect 1782 1672 1812 1714
rect 2218 1672 2248 1714
rect 2362 1672 2392 1714
rect 2798 1672 2828 1714
rect 2942 1672 2972 1714
rect 3378 1672 3408 1714
rect 3522 1672 3552 1714
rect 3958 1672 3988 1714
rect 4102 1672 4132 1714
rect 4538 1672 4568 1714
rect 4682 1672 4712 1714
rect 5118 1672 5148 1714
rect 5262 1672 5292 1714
rect 5698 1672 5728 1714
rect 5842 1672 5872 1714
rect 6278 1672 6308 1714
rect 6422 1672 6452 1714
rect 6858 1672 6888 1714
rect 106 1548 136 1576
rect 414 1548 444 1576
rect 686 1548 716 1576
rect 994 1548 1024 1576
rect 1266 1548 1296 1576
rect 1574 1548 1604 1576
rect 1846 1548 1876 1576
rect 2154 1548 2184 1576
rect 2426 1548 2456 1576
rect 2734 1548 2764 1576
rect 3006 1548 3036 1576
rect 3314 1548 3344 1576
rect 3586 1548 3616 1576
rect 3894 1548 3924 1576
rect 4166 1548 4196 1576
rect 4474 1548 4504 1576
rect 4746 1548 4776 1576
rect 5054 1548 5084 1576
rect 5326 1548 5356 1576
rect 5634 1548 5664 1576
rect 5906 1548 5936 1576
rect 6214 1548 6244 1576
rect 6486 1548 6516 1576
rect 6794 1548 6824 1576
rect 42 1402 72 1444
rect 478 1402 508 1444
rect 622 1402 652 1444
rect 1058 1402 1088 1444
rect 1202 1402 1232 1444
rect 1638 1402 1668 1444
rect 1782 1402 1812 1444
rect 2218 1402 2248 1444
rect 2362 1402 2392 1444
rect 2798 1402 2828 1444
rect 2942 1402 2972 1444
rect 3378 1402 3408 1444
rect 3522 1402 3552 1444
rect 3958 1402 3988 1444
rect 4102 1402 4132 1444
rect 4538 1402 4568 1444
rect 4682 1402 4712 1444
rect 5118 1402 5148 1444
rect 5262 1402 5292 1444
rect 5698 1402 5728 1444
rect 5842 1402 5872 1444
rect 6278 1402 6308 1444
rect 6422 1402 6452 1444
rect 6858 1402 6888 1444
rect 106 1278 136 1306
rect 414 1278 444 1306
rect 686 1278 716 1306
rect 994 1278 1024 1306
rect 1266 1278 1296 1306
rect 1574 1278 1604 1306
rect 1846 1278 1876 1306
rect 2154 1278 2184 1306
rect 2426 1278 2456 1306
rect 2734 1278 2764 1306
rect 3006 1278 3036 1306
rect 3314 1278 3344 1306
rect 3586 1278 3616 1306
rect 3894 1278 3924 1306
rect 4166 1278 4196 1306
rect 4474 1278 4504 1306
rect 4746 1278 4776 1306
rect 5054 1278 5084 1306
rect 5326 1278 5356 1306
rect 5634 1278 5664 1306
rect 5906 1278 5936 1306
rect 6214 1278 6244 1306
rect 6486 1278 6516 1306
rect 6794 1278 6824 1306
rect 42 1132 72 1174
rect 478 1132 508 1174
rect 622 1132 652 1174
rect 1058 1132 1088 1174
rect 1202 1132 1232 1174
rect 1638 1132 1668 1174
rect 1782 1132 1812 1174
rect 2218 1132 2248 1174
rect 2362 1132 2392 1174
rect 2798 1132 2828 1174
rect 2942 1132 2972 1174
rect 3378 1132 3408 1174
rect 3522 1132 3552 1174
rect 3958 1132 3988 1174
rect 4102 1132 4132 1174
rect 4538 1132 4568 1174
rect 4682 1132 4712 1174
rect 5118 1132 5148 1174
rect 5262 1132 5292 1174
rect 5698 1132 5728 1174
rect 5842 1132 5872 1174
rect 6278 1132 6308 1174
rect 6422 1132 6452 1174
rect 6858 1132 6888 1174
rect 106 1008 136 1036
rect 414 1008 444 1036
rect 686 1008 716 1036
rect 994 1008 1024 1036
rect 1266 1008 1296 1036
rect 1574 1008 1604 1036
rect 1846 1008 1876 1036
rect 2154 1008 2184 1036
rect 2426 1008 2456 1036
rect 2734 1008 2764 1036
rect 3006 1008 3036 1036
rect 3314 1008 3344 1036
rect 3586 1008 3616 1036
rect 3894 1008 3924 1036
rect 4166 1008 4196 1036
rect 4474 1008 4504 1036
rect 4746 1008 4776 1036
rect 5054 1008 5084 1036
rect 5326 1008 5356 1036
rect 5634 1008 5664 1036
rect 5906 1008 5936 1036
rect 6214 1008 6244 1036
rect 6486 1008 6516 1036
rect 6794 1008 6824 1036
rect 42 862 72 904
rect 478 862 508 904
rect 622 862 652 904
rect 1058 862 1088 904
rect 1202 862 1232 904
rect 1638 862 1668 904
rect 1782 862 1812 904
rect 2218 862 2248 904
rect 2362 862 2392 904
rect 2798 862 2828 904
rect 2942 862 2972 904
rect 3378 862 3408 904
rect 3522 862 3552 904
rect 3958 862 3988 904
rect 4102 862 4132 904
rect 4538 862 4568 904
rect 4682 862 4712 904
rect 5118 862 5148 904
rect 5262 862 5292 904
rect 5698 862 5728 904
rect 5842 862 5872 904
rect 6278 862 6308 904
rect 6422 862 6452 904
rect 6858 862 6888 904
rect 106 738 136 766
rect 414 738 444 766
rect 686 738 716 766
rect 994 738 1024 766
rect 1266 738 1296 766
rect 1574 738 1604 766
rect 1846 738 1876 766
rect 2154 738 2184 766
rect 2426 738 2456 766
rect 2734 738 2764 766
rect 3006 738 3036 766
rect 3314 738 3344 766
rect 3586 738 3616 766
rect 3894 738 3924 766
rect 4166 738 4196 766
rect 4474 738 4504 766
rect 4746 738 4776 766
rect 5054 738 5084 766
rect 5326 738 5356 766
rect 5634 738 5664 766
rect 5906 738 5936 766
rect 6214 738 6244 766
rect 6486 738 6516 766
rect 6794 738 6824 766
rect 42 592 72 634
rect 478 592 508 634
rect 622 592 652 634
rect 1058 592 1088 634
rect 1202 592 1232 634
rect 1638 592 1668 634
rect 1782 592 1812 634
rect 2218 592 2248 634
rect 2362 592 2392 634
rect 2798 592 2828 634
rect 2942 592 2972 634
rect 3378 592 3408 634
rect 3522 592 3552 634
rect 3958 592 3988 634
rect 4102 592 4132 634
rect 4538 592 4568 634
rect 4682 592 4712 634
rect 5118 592 5148 634
rect 5262 592 5292 634
rect 5698 592 5728 634
rect 5842 592 5872 634
rect 6278 592 6308 634
rect 6422 592 6452 634
rect 6858 592 6888 634
rect 106 468 136 496
rect 414 468 444 496
rect 686 468 716 496
rect 994 468 1024 496
rect 1266 468 1296 496
rect 1574 468 1604 496
rect 1846 468 1876 496
rect 2154 468 2184 496
rect 2426 468 2456 496
rect 2734 468 2764 496
rect 3006 468 3036 496
rect 3314 468 3344 496
rect 3586 468 3616 496
rect 3894 468 3924 496
rect 4166 468 4196 496
rect 4474 468 4504 496
rect 4746 468 4776 496
rect 5054 468 5084 496
rect 5326 468 5356 496
rect 5634 468 5664 496
rect 5906 468 5936 496
rect 6214 468 6244 496
rect 6486 468 6516 496
rect 6794 468 6824 496
rect 42 322 72 364
rect 478 322 508 364
rect 622 322 652 364
rect 1058 322 1088 364
rect 1202 322 1232 364
rect 1638 322 1668 364
rect 1782 322 1812 364
rect 2218 322 2248 364
rect 2362 322 2392 364
rect 2798 322 2828 364
rect 2942 322 2972 364
rect 3378 322 3408 364
rect 3522 322 3552 364
rect 3958 322 3988 364
rect 4102 322 4132 364
rect 4538 322 4568 364
rect 4682 322 4712 364
rect 5118 322 5148 364
rect 5262 322 5292 364
rect 5698 322 5728 364
rect 5842 322 5872 364
rect 6278 322 6308 364
rect 6422 322 6452 364
rect 6858 322 6888 364
rect 106 198 136 226
rect 414 198 444 226
rect 686 198 716 226
rect 994 198 1024 226
rect 1266 198 1296 226
rect 1574 198 1604 226
rect 1846 198 1876 226
rect 2154 198 2184 226
rect 2426 198 2456 226
rect 2734 198 2764 226
rect 3006 198 3036 226
rect 3314 198 3344 226
rect 3586 198 3616 226
rect 3894 198 3924 226
rect 4166 198 4196 226
rect 4474 198 4504 226
rect 4746 198 4776 226
rect 5054 198 5084 226
rect 5326 198 5356 226
rect 5634 198 5664 226
rect 5906 198 5936 226
rect 6214 198 6244 226
rect 6486 198 6516 226
rect 6794 198 6824 226
rect 42 52 72 94
rect 478 52 508 94
rect 622 52 652 94
rect 1058 52 1088 94
rect 1202 52 1232 94
rect 1638 52 1668 94
rect 1782 52 1812 94
rect 2218 52 2248 94
rect 2362 52 2392 94
rect 2798 52 2828 94
rect 2942 52 2972 94
rect 3378 52 3408 94
rect 3522 52 3552 94
rect 3958 52 3988 94
rect 4102 52 4132 94
rect 4538 52 4568 94
rect 4682 52 4712 94
rect 5118 52 5148 94
rect 5262 52 5292 94
rect 5698 52 5728 94
rect 5842 52 5872 94
rect 6278 52 6308 94
rect 6422 52 6452 94
rect 6858 52 6888 94
rect 106 -72 136 -44
rect 414 -72 444 -44
rect 686 -72 716 -44
rect 994 -72 1024 -44
rect 1266 -72 1296 -44
rect 1574 -72 1604 -44
rect 1846 -72 1876 -44
rect 2154 -72 2184 -44
rect 2426 -72 2456 -44
rect 2734 -72 2764 -44
rect 3006 -72 3036 -44
rect 3314 -72 3344 -44
rect 3586 -72 3616 -44
rect 3894 -72 3924 -44
rect 4166 -72 4196 -44
rect 4474 -72 4504 -44
rect 4746 -72 4776 -44
rect 5054 -72 5084 -44
rect 5326 -72 5356 -44
rect 5634 -72 5664 -44
rect 5906 -72 5936 -44
rect 6214 -72 6244 -44
rect 6486 -72 6516 -44
rect 6794 -72 6824 -44
rect 42 -218 72 -176
rect 478 -218 508 -176
rect 622 -218 652 -176
rect 1058 -218 1088 -176
rect 1202 -218 1232 -176
rect 1638 -218 1668 -176
rect 1782 -218 1812 -176
rect 2218 -218 2248 -176
rect 2362 -218 2392 -176
rect 2798 -218 2828 -176
rect 2942 -218 2972 -176
rect 3378 -218 3408 -176
rect 3522 -218 3552 -176
rect 3958 -218 3988 -176
rect 4102 -218 4132 -176
rect 4538 -218 4568 -176
rect 4682 -218 4712 -176
rect 5118 -218 5148 -176
rect 5262 -218 5292 -176
rect 5698 -218 5728 -176
rect 5842 -218 5872 -176
rect 6278 -218 6308 -176
rect 6422 -218 6452 -176
rect 6858 -218 6888 -176
rect 106 -342 136 -314
rect 414 -342 444 -314
rect 686 -342 716 -314
rect 994 -342 1024 -314
rect 1266 -342 1296 -314
rect 1574 -342 1604 -314
rect 1846 -342 1876 -314
rect 2154 -342 2184 -314
rect 2426 -342 2456 -314
rect 2734 -342 2764 -314
rect 3006 -342 3036 -314
rect 3314 -342 3344 -314
rect 3586 -342 3616 -314
rect 3894 -342 3924 -314
rect 4166 -342 4196 -314
rect 4474 -342 4504 -314
rect 4746 -342 4776 -314
rect 5054 -342 5084 -314
rect 5326 -342 5356 -314
rect 5634 -342 5664 -314
rect 5906 -342 5936 -314
rect 6214 -342 6244 -314
rect 6486 -342 6516 -314
rect 6794 -342 6824 -314
rect 42 -488 72 -446
rect 478 -488 508 -446
rect 622 -488 652 -446
rect 1058 -488 1088 -446
rect 1202 -488 1232 -446
rect 1638 -488 1668 -446
rect 1782 -488 1812 -446
rect 2218 -488 2248 -446
rect 2362 -488 2392 -446
rect 2798 -488 2828 -446
rect 2942 -488 2972 -446
rect 3378 -488 3408 -446
rect 3522 -488 3552 -446
rect 3958 -488 3988 -446
rect 4102 -488 4132 -446
rect 4538 -488 4568 -446
rect 4682 -488 4712 -446
rect 5118 -488 5148 -446
rect 5262 -488 5292 -446
rect 5698 -488 5728 -446
rect 5842 -488 5872 -446
rect 6278 -488 6308 -446
rect 6422 -488 6452 -446
rect 6858 -488 6888 -446
rect 106 -612 136 -584
rect 414 -612 444 -584
rect 686 -612 716 -584
rect 994 -612 1024 -584
rect 1266 -612 1296 -584
rect 1574 -612 1604 -584
rect 1846 -612 1876 -584
rect 2154 -612 2184 -584
rect 2426 -612 2456 -584
rect 2734 -612 2764 -584
rect 3006 -612 3036 -584
rect 3314 -612 3344 -584
rect 3586 -612 3616 -584
rect 3894 -612 3924 -584
rect 4166 -612 4196 -584
rect 4474 -612 4504 -584
rect 4746 -612 4776 -584
rect 5054 -612 5084 -584
rect 5326 -612 5356 -584
rect 5634 -612 5664 -584
rect 5906 -612 5936 -584
rect 6214 -612 6244 -584
rect 6486 -612 6516 -584
rect 6794 -612 6824 -584
rect 42 -758 72 -716
rect 478 -758 508 -716
rect 622 -758 652 -716
rect 1058 -758 1088 -716
rect 1202 -758 1232 -716
rect 1638 -758 1668 -716
rect 1782 -758 1812 -716
rect 2218 -758 2248 -716
rect 2362 -758 2392 -716
rect 2798 -758 2828 -716
rect 2942 -758 2972 -716
rect 3378 -758 3408 -716
rect 3522 -758 3552 -716
rect 3958 -758 3988 -716
rect 4102 -758 4132 -716
rect 4538 -758 4568 -716
rect 4682 -758 4712 -716
rect 5118 -758 5148 -716
rect 5262 -758 5292 -716
rect 5698 -758 5728 -716
rect 5842 -758 5872 -716
rect 6278 -758 6308 -716
rect 6422 -758 6452 -716
rect 6858 -758 6888 -716
rect 106 -882 136 -854
rect 414 -882 444 -854
rect 686 -882 716 -854
rect 994 -882 1024 -854
rect 1266 -882 1296 -854
rect 1574 -882 1604 -854
rect 1846 -882 1876 -854
rect 2154 -882 2184 -854
rect 2426 -882 2456 -854
rect 2734 -882 2764 -854
rect 3006 -882 3036 -854
rect 3314 -882 3344 -854
rect 3586 -882 3616 -854
rect 3894 -882 3924 -854
rect 4166 -882 4196 -854
rect 4474 -882 4504 -854
rect 4746 -882 4776 -854
rect 5054 -882 5084 -854
rect 5326 -882 5356 -854
rect 5634 -882 5664 -854
rect 5906 -882 5936 -854
rect 6214 -882 6244 -854
rect 6486 -882 6516 -854
rect 6794 -882 6824 -854
rect 42 -1028 72 -986
rect 478 -1028 508 -986
rect 622 -1028 652 -986
rect 1058 -1028 1088 -986
rect 1202 -1028 1232 -986
rect 1638 -1028 1668 -986
rect 1782 -1028 1812 -986
rect 2218 -1028 2248 -986
rect 2362 -1028 2392 -986
rect 2798 -1028 2828 -986
rect 2942 -1028 2972 -986
rect 3378 -1028 3408 -986
rect 3522 -1028 3552 -986
rect 3958 -1028 3988 -986
rect 4102 -1028 4132 -986
rect 4538 -1028 4568 -986
rect 4682 -1028 4712 -986
rect 5118 -1028 5148 -986
rect 5262 -1028 5292 -986
rect 5698 -1028 5728 -986
rect 5842 -1028 5872 -986
rect 6278 -1028 6308 -986
rect 6422 -1028 6452 -986
rect 6858 -1028 6888 -986
rect 106 -1152 136 -1124
rect 414 -1152 444 -1124
rect 686 -1152 716 -1124
rect 994 -1152 1024 -1124
rect 1266 -1152 1296 -1124
rect 1574 -1152 1604 -1124
rect 1846 -1152 1876 -1124
rect 2154 -1152 2184 -1124
rect 2426 -1152 2456 -1124
rect 2734 -1152 2764 -1124
rect 3006 -1152 3036 -1124
rect 3314 -1152 3344 -1124
rect 3586 -1152 3616 -1124
rect 3894 -1152 3924 -1124
rect 4166 -1152 4196 -1124
rect 4474 -1152 4504 -1124
rect 4746 -1152 4776 -1124
rect 5054 -1152 5084 -1124
rect 5326 -1152 5356 -1124
rect 5634 -1152 5664 -1124
rect 5906 -1152 5936 -1124
rect 6214 -1152 6244 -1124
rect 6486 -1152 6516 -1124
rect 6794 -1152 6824 -1124
rect 42 -1298 72 -1256
rect 478 -1298 508 -1256
rect 622 -1298 652 -1256
rect 1058 -1298 1088 -1256
rect 1202 -1298 1232 -1256
rect 1638 -1298 1668 -1256
rect 1782 -1298 1812 -1256
rect 2218 -1298 2248 -1256
rect 2362 -1298 2392 -1256
rect 2798 -1298 2828 -1256
rect 2942 -1298 2972 -1256
rect 3378 -1298 3408 -1256
rect 3522 -1298 3552 -1256
rect 3958 -1298 3988 -1256
rect 4102 -1298 4132 -1256
rect 4538 -1298 4568 -1256
rect 4682 -1298 4712 -1256
rect 5118 -1298 5148 -1256
rect 5262 -1298 5292 -1256
rect 5698 -1298 5728 -1256
rect 5842 -1298 5872 -1256
rect 6278 -1298 6308 -1256
rect 6422 -1298 6452 -1256
rect 6858 -1298 6888 -1256
rect 106 -1422 136 -1394
rect 414 -1422 444 -1394
rect 686 -1422 716 -1394
rect 994 -1422 1024 -1394
rect 1266 -1422 1296 -1394
rect 1574 -1422 1604 -1394
rect 1846 -1422 1876 -1394
rect 2154 -1422 2184 -1394
rect 2426 -1422 2456 -1394
rect 2734 -1422 2764 -1394
rect 3006 -1422 3036 -1394
rect 3314 -1422 3344 -1394
rect 3586 -1422 3616 -1394
rect 3894 -1422 3924 -1394
rect 4166 -1422 4196 -1394
rect 4474 -1422 4504 -1394
rect 4746 -1422 4776 -1394
rect 5054 -1422 5084 -1394
rect 5326 -1422 5356 -1394
rect 5634 -1422 5664 -1394
rect 5906 -1422 5936 -1394
rect 6214 -1422 6244 -1394
rect 6486 -1422 6516 -1394
rect 6794 -1422 6824 -1394
rect 42 -1568 72 -1526
rect 478 -1568 508 -1526
rect 622 -1568 652 -1526
rect 1058 -1568 1088 -1526
rect 1202 -1568 1232 -1526
rect 1638 -1568 1668 -1526
rect 1782 -1568 1812 -1526
rect 2218 -1568 2248 -1526
rect 2362 -1568 2392 -1526
rect 2798 -1568 2828 -1526
rect 2942 -1568 2972 -1526
rect 3378 -1568 3408 -1526
rect 3522 -1568 3552 -1526
rect 3958 -1568 3988 -1526
rect 4102 -1568 4132 -1526
rect 4538 -1568 4568 -1526
rect 4682 -1568 4712 -1526
rect 5118 -1568 5148 -1526
rect 5262 -1568 5292 -1526
rect 5698 -1568 5728 -1526
rect 5842 -1568 5872 -1526
rect 6278 -1568 6308 -1526
rect 6422 -1568 6452 -1526
rect 6858 -1568 6888 -1526
rect 106 -1692 136 -1664
rect 414 -1692 444 -1664
rect 686 -1692 716 -1664
rect 994 -1692 1024 -1664
rect 1266 -1692 1296 -1664
rect 1574 -1692 1604 -1664
rect 1846 -1692 1876 -1664
rect 2154 -1692 2184 -1664
rect 2426 -1692 2456 -1664
rect 2734 -1692 2764 -1664
rect 3006 -1692 3036 -1664
rect 3314 -1692 3344 -1664
rect 3586 -1692 3616 -1664
rect 3894 -1692 3924 -1664
rect 4166 -1692 4196 -1664
rect 4474 -1692 4504 -1664
rect 4746 -1692 4776 -1664
rect 5054 -1692 5084 -1664
rect 5326 -1692 5356 -1664
rect 5634 -1692 5664 -1664
rect 5906 -1692 5936 -1664
rect 6214 -1692 6244 -1664
rect 6486 -1692 6516 -1664
rect 6794 -1692 6824 -1664
rect 42 -1838 72 -1796
rect 478 -1838 508 -1796
rect 622 -1838 652 -1796
rect 1058 -1838 1088 -1796
rect 1202 -1838 1232 -1796
rect 1638 -1838 1668 -1796
rect 1782 -1838 1812 -1796
rect 2218 -1838 2248 -1796
rect 2362 -1838 2392 -1796
rect 2798 -1838 2828 -1796
rect 2942 -1838 2972 -1796
rect 3378 -1838 3408 -1796
rect 3522 -1838 3552 -1796
rect 3958 -1838 3988 -1796
rect 4102 -1838 4132 -1796
rect 4538 -1838 4568 -1796
rect 4682 -1838 4712 -1796
rect 5118 -1838 5148 -1796
rect 5262 -1838 5292 -1796
rect 5698 -1838 5728 -1796
rect 5842 -1838 5872 -1796
rect 6278 -1838 6308 -1796
rect 6422 -1838 6452 -1796
rect 6858 -1838 6888 -1796
rect 106 -1962 136 -1934
rect 414 -1962 444 -1934
rect 686 -1962 716 -1934
rect 994 -1962 1024 -1934
rect 1266 -1962 1296 -1934
rect 1574 -1962 1604 -1934
rect 1846 -1962 1876 -1934
rect 2154 -1962 2184 -1934
rect 2426 -1962 2456 -1934
rect 2734 -1962 2764 -1934
rect 3006 -1962 3036 -1934
rect 3314 -1962 3344 -1934
rect 3586 -1962 3616 -1934
rect 3894 -1962 3924 -1934
rect 4166 -1962 4196 -1934
rect 4474 -1962 4504 -1934
rect 4746 -1962 4776 -1934
rect 5054 -1962 5084 -1934
rect 5326 -1962 5356 -1934
rect 5634 -1962 5664 -1934
rect 5906 -1962 5936 -1934
rect 6214 -1962 6244 -1934
rect 6486 -1962 6516 -1934
rect 6794 -1962 6824 -1934
rect 42 -2108 72 -2066
rect 478 -2108 508 -2066
rect 622 -2108 652 -2066
rect 1058 -2108 1088 -2066
rect 1202 -2108 1232 -2066
rect 1638 -2108 1668 -2066
rect 1782 -2108 1812 -2066
rect 2218 -2108 2248 -2066
rect 2362 -2108 2392 -2066
rect 2798 -2108 2828 -2066
rect 2942 -2108 2972 -2066
rect 3378 -2108 3408 -2066
rect 3522 -2108 3552 -2066
rect 3958 -2108 3988 -2066
rect 4102 -2108 4132 -2066
rect 4538 -2108 4568 -2066
rect 4682 -2108 4712 -2066
rect 5118 -2108 5148 -2066
rect 5262 -2108 5292 -2066
rect 5698 -2108 5728 -2066
rect 5842 -2108 5872 -2066
rect 6278 -2108 6308 -2066
rect 6422 -2108 6452 -2066
rect 6858 -2108 6888 -2066
<< npd >>
rect 221 1942 251 1984
rect 299 1942 329 1984
rect 801 1942 831 1984
rect 879 1942 909 1984
rect 1381 1942 1411 1984
rect 1459 1942 1489 1984
rect 1961 1942 1991 1984
rect 2039 1942 2069 1984
rect 2541 1942 2571 1984
rect 2619 1942 2649 1984
rect 3121 1942 3151 1984
rect 3199 1942 3229 1984
rect 3701 1942 3731 1984
rect 3779 1942 3809 1984
rect 4281 1942 4311 1984
rect 4359 1942 4389 1984
rect 4861 1942 4891 1984
rect 4939 1942 4969 1984
rect 5441 1942 5471 1984
rect 5519 1942 5549 1984
rect 6021 1942 6051 1984
rect 6099 1942 6129 1984
rect 6601 1942 6631 1984
rect 6679 1942 6709 1984
rect 221 1672 251 1714
rect 299 1672 329 1714
rect 801 1672 831 1714
rect 879 1672 909 1714
rect 1381 1672 1411 1714
rect 1459 1672 1489 1714
rect 1961 1672 1991 1714
rect 2039 1672 2069 1714
rect 2541 1672 2571 1714
rect 2619 1672 2649 1714
rect 3121 1672 3151 1714
rect 3199 1672 3229 1714
rect 3701 1672 3731 1714
rect 3779 1672 3809 1714
rect 4281 1672 4311 1714
rect 4359 1672 4389 1714
rect 4861 1672 4891 1714
rect 4939 1672 4969 1714
rect 5441 1672 5471 1714
rect 5519 1672 5549 1714
rect 6021 1672 6051 1714
rect 6099 1672 6129 1714
rect 6601 1672 6631 1714
rect 6679 1672 6709 1714
rect 221 1402 251 1444
rect 299 1402 329 1444
rect 801 1402 831 1444
rect 879 1402 909 1444
rect 1381 1402 1411 1444
rect 1459 1402 1489 1444
rect 1961 1402 1991 1444
rect 2039 1402 2069 1444
rect 2541 1402 2571 1444
rect 2619 1402 2649 1444
rect 3121 1402 3151 1444
rect 3199 1402 3229 1444
rect 3701 1402 3731 1444
rect 3779 1402 3809 1444
rect 4281 1402 4311 1444
rect 4359 1402 4389 1444
rect 4861 1402 4891 1444
rect 4939 1402 4969 1444
rect 5441 1402 5471 1444
rect 5519 1402 5549 1444
rect 6021 1402 6051 1444
rect 6099 1402 6129 1444
rect 6601 1402 6631 1444
rect 6679 1402 6709 1444
rect 221 1132 251 1174
rect 299 1132 329 1174
rect 801 1132 831 1174
rect 879 1132 909 1174
rect 1381 1132 1411 1174
rect 1459 1132 1489 1174
rect 1961 1132 1991 1174
rect 2039 1132 2069 1174
rect 2541 1132 2571 1174
rect 2619 1132 2649 1174
rect 3121 1132 3151 1174
rect 3199 1132 3229 1174
rect 3701 1132 3731 1174
rect 3779 1132 3809 1174
rect 4281 1132 4311 1174
rect 4359 1132 4389 1174
rect 4861 1132 4891 1174
rect 4939 1132 4969 1174
rect 5441 1132 5471 1174
rect 5519 1132 5549 1174
rect 6021 1132 6051 1174
rect 6099 1132 6129 1174
rect 6601 1132 6631 1174
rect 6679 1132 6709 1174
rect 221 862 251 904
rect 299 862 329 904
rect 801 862 831 904
rect 879 862 909 904
rect 1381 862 1411 904
rect 1459 862 1489 904
rect 1961 862 1991 904
rect 2039 862 2069 904
rect 2541 862 2571 904
rect 2619 862 2649 904
rect 3121 862 3151 904
rect 3199 862 3229 904
rect 3701 862 3731 904
rect 3779 862 3809 904
rect 4281 862 4311 904
rect 4359 862 4389 904
rect 4861 862 4891 904
rect 4939 862 4969 904
rect 5441 862 5471 904
rect 5519 862 5549 904
rect 6021 862 6051 904
rect 6099 862 6129 904
rect 6601 862 6631 904
rect 6679 862 6709 904
rect 221 592 251 634
rect 299 592 329 634
rect 801 592 831 634
rect 879 592 909 634
rect 1381 592 1411 634
rect 1459 592 1489 634
rect 1961 592 1991 634
rect 2039 592 2069 634
rect 2541 592 2571 634
rect 2619 592 2649 634
rect 3121 592 3151 634
rect 3199 592 3229 634
rect 3701 592 3731 634
rect 3779 592 3809 634
rect 4281 592 4311 634
rect 4359 592 4389 634
rect 4861 592 4891 634
rect 4939 592 4969 634
rect 5441 592 5471 634
rect 5519 592 5549 634
rect 6021 592 6051 634
rect 6099 592 6129 634
rect 6601 592 6631 634
rect 6679 592 6709 634
rect 221 322 251 364
rect 299 322 329 364
rect 801 322 831 364
rect 879 322 909 364
rect 1381 322 1411 364
rect 1459 322 1489 364
rect 1961 322 1991 364
rect 2039 322 2069 364
rect 2541 322 2571 364
rect 2619 322 2649 364
rect 3121 322 3151 364
rect 3199 322 3229 364
rect 3701 322 3731 364
rect 3779 322 3809 364
rect 4281 322 4311 364
rect 4359 322 4389 364
rect 4861 322 4891 364
rect 4939 322 4969 364
rect 5441 322 5471 364
rect 5519 322 5549 364
rect 6021 322 6051 364
rect 6099 322 6129 364
rect 6601 322 6631 364
rect 6679 322 6709 364
rect 221 52 251 94
rect 299 52 329 94
rect 801 52 831 94
rect 879 52 909 94
rect 1381 52 1411 94
rect 1459 52 1489 94
rect 1961 52 1991 94
rect 2039 52 2069 94
rect 2541 52 2571 94
rect 2619 52 2649 94
rect 3121 52 3151 94
rect 3199 52 3229 94
rect 3701 52 3731 94
rect 3779 52 3809 94
rect 4281 52 4311 94
rect 4359 52 4389 94
rect 4861 52 4891 94
rect 4939 52 4969 94
rect 5441 52 5471 94
rect 5519 52 5549 94
rect 6021 52 6051 94
rect 6099 52 6129 94
rect 6601 52 6631 94
rect 6679 52 6709 94
rect 221 -218 251 -176
rect 299 -218 329 -176
rect 801 -218 831 -176
rect 879 -218 909 -176
rect 1381 -218 1411 -176
rect 1459 -218 1489 -176
rect 1961 -218 1991 -176
rect 2039 -218 2069 -176
rect 2541 -218 2571 -176
rect 2619 -218 2649 -176
rect 3121 -218 3151 -176
rect 3199 -218 3229 -176
rect 3701 -218 3731 -176
rect 3779 -218 3809 -176
rect 4281 -218 4311 -176
rect 4359 -218 4389 -176
rect 4861 -218 4891 -176
rect 4939 -218 4969 -176
rect 5441 -218 5471 -176
rect 5519 -218 5549 -176
rect 6021 -218 6051 -176
rect 6099 -218 6129 -176
rect 6601 -218 6631 -176
rect 6679 -218 6709 -176
rect 221 -488 251 -446
rect 299 -488 329 -446
rect 801 -488 831 -446
rect 879 -488 909 -446
rect 1381 -488 1411 -446
rect 1459 -488 1489 -446
rect 1961 -488 1991 -446
rect 2039 -488 2069 -446
rect 2541 -488 2571 -446
rect 2619 -488 2649 -446
rect 3121 -488 3151 -446
rect 3199 -488 3229 -446
rect 3701 -488 3731 -446
rect 3779 -488 3809 -446
rect 4281 -488 4311 -446
rect 4359 -488 4389 -446
rect 4861 -488 4891 -446
rect 4939 -488 4969 -446
rect 5441 -488 5471 -446
rect 5519 -488 5549 -446
rect 6021 -488 6051 -446
rect 6099 -488 6129 -446
rect 6601 -488 6631 -446
rect 6679 -488 6709 -446
rect 221 -758 251 -716
rect 299 -758 329 -716
rect 801 -758 831 -716
rect 879 -758 909 -716
rect 1381 -758 1411 -716
rect 1459 -758 1489 -716
rect 1961 -758 1991 -716
rect 2039 -758 2069 -716
rect 2541 -758 2571 -716
rect 2619 -758 2649 -716
rect 3121 -758 3151 -716
rect 3199 -758 3229 -716
rect 3701 -758 3731 -716
rect 3779 -758 3809 -716
rect 4281 -758 4311 -716
rect 4359 -758 4389 -716
rect 4861 -758 4891 -716
rect 4939 -758 4969 -716
rect 5441 -758 5471 -716
rect 5519 -758 5549 -716
rect 6021 -758 6051 -716
rect 6099 -758 6129 -716
rect 6601 -758 6631 -716
rect 6679 -758 6709 -716
rect 221 -1028 251 -986
rect 299 -1028 329 -986
rect 801 -1028 831 -986
rect 879 -1028 909 -986
rect 1381 -1028 1411 -986
rect 1459 -1028 1489 -986
rect 1961 -1028 1991 -986
rect 2039 -1028 2069 -986
rect 2541 -1028 2571 -986
rect 2619 -1028 2649 -986
rect 3121 -1028 3151 -986
rect 3199 -1028 3229 -986
rect 3701 -1028 3731 -986
rect 3779 -1028 3809 -986
rect 4281 -1028 4311 -986
rect 4359 -1028 4389 -986
rect 4861 -1028 4891 -986
rect 4939 -1028 4969 -986
rect 5441 -1028 5471 -986
rect 5519 -1028 5549 -986
rect 6021 -1028 6051 -986
rect 6099 -1028 6129 -986
rect 6601 -1028 6631 -986
rect 6679 -1028 6709 -986
rect 221 -1298 251 -1256
rect 299 -1298 329 -1256
rect 801 -1298 831 -1256
rect 879 -1298 909 -1256
rect 1381 -1298 1411 -1256
rect 1459 -1298 1489 -1256
rect 1961 -1298 1991 -1256
rect 2039 -1298 2069 -1256
rect 2541 -1298 2571 -1256
rect 2619 -1298 2649 -1256
rect 3121 -1298 3151 -1256
rect 3199 -1298 3229 -1256
rect 3701 -1298 3731 -1256
rect 3779 -1298 3809 -1256
rect 4281 -1298 4311 -1256
rect 4359 -1298 4389 -1256
rect 4861 -1298 4891 -1256
rect 4939 -1298 4969 -1256
rect 5441 -1298 5471 -1256
rect 5519 -1298 5549 -1256
rect 6021 -1298 6051 -1256
rect 6099 -1298 6129 -1256
rect 6601 -1298 6631 -1256
rect 6679 -1298 6709 -1256
rect 221 -1568 251 -1526
rect 299 -1568 329 -1526
rect 801 -1568 831 -1526
rect 879 -1568 909 -1526
rect 1381 -1568 1411 -1526
rect 1459 -1568 1489 -1526
rect 1961 -1568 1991 -1526
rect 2039 -1568 2069 -1526
rect 2541 -1568 2571 -1526
rect 2619 -1568 2649 -1526
rect 3121 -1568 3151 -1526
rect 3199 -1568 3229 -1526
rect 3701 -1568 3731 -1526
rect 3779 -1568 3809 -1526
rect 4281 -1568 4311 -1526
rect 4359 -1568 4389 -1526
rect 4861 -1568 4891 -1526
rect 4939 -1568 4969 -1526
rect 5441 -1568 5471 -1526
rect 5519 -1568 5549 -1526
rect 6021 -1568 6051 -1526
rect 6099 -1568 6129 -1526
rect 6601 -1568 6631 -1526
rect 6679 -1568 6709 -1526
rect 221 -1838 251 -1796
rect 299 -1838 329 -1796
rect 801 -1838 831 -1796
rect 879 -1838 909 -1796
rect 1381 -1838 1411 -1796
rect 1459 -1838 1489 -1796
rect 1961 -1838 1991 -1796
rect 2039 -1838 2069 -1796
rect 2541 -1838 2571 -1796
rect 2619 -1838 2649 -1796
rect 3121 -1838 3151 -1796
rect 3199 -1838 3229 -1796
rect 3701 -1838 3731 -1796
rect 3779 -1838 3809 -1796
rect 4281 -1838 4311 -1796
rect 4359 -1838 4389 -1796
rect 4861 -1838 4891 -1796
rect 4939 -1838 4969 -1796
rect 5441 -1838 5471 -1796
rect 5519 -1838 5549 -1796
rect 6021 -1838 6051 -1796
rect 6099 -1838 6129 -1796
rect 6601 -1838 6631 -1796
rect 6679 -1838 6709 -1796
rect 221 -2108 251 -2066
rect 299 -2108 329 -2066
rect 801 -2108 831 -2066
rect 879 -2108 909 -2066
rect 1381 -2108 1411 -2066
rect 1459 -2108 1489 -2066
rect 1961 -2108 1991 -2066
rect 2039 -2108 2069 -2066
rect 2541 -2108 2571 -2066
rect 2619 -2108 2649 -2066
rect 3121 -2108 3151 -2066
rect 3199 -2108 3229 -2066
rect 3701 -2108 3731 -2066
rect 3779 -2108 3809 -2066
rect 4281 -2108 4311 -2066
rect 4359 -2108 4389 -2066
rect 4861 -2108 4891 -2066
rect 4939 -2108 4969 -2066
rect 5441 -2108 5471 -2066
rect 5519 -2108 5549 -2066
rect 6021 -2108 6051 -2066
rect 6099 -2108 6129 -2066
rect 6601 -2108 6631 -2066
rect 6679 -2108 6709 -2066
<< npass >>
rect 128 1942 158 1970
rect 392 1942 422 1970
rect 708 1942 738 1970
rect 972 1942 1002 1970
rect 1288 1942 1318 1970
rect 1552 1942 1582 1970
rect 1868 1942 1898 1970
rect 2132 1942 2162 1970
rect 2448 1942 2478 1970
rect 2712 1942 2742 1970
rect 3028 1942 3058 1970
rect 3292 1942 3322 1970
rect 3608 1942 3638 1970
rect 3872 1942 3902 1970
rect 4188 1942 4218 1970
rect 4452 1942 4482 1970
rect 4768 1942 4798 1970
rect 5032 1942 5062 1970
rect 5348 1942 5378 1970
rect 5612 1942 5642 1970
rect 5928 1942 5958 1970
rect 6192 1942 6222 1970
rect 6508 1942 6538 1970
rect 6772 1942 6802 1970
rect 128 1672 158 1700
rect 392 1672 422 1700
rect 708 1672 738 1700
rect 972 1672 1002 1700
rect 1288 1672 1318 1700
rect 1552 1672 1582 1700
rect 1868 1672 1898 1700
rect 2132 1672 2162 1700
rect 2448 1672 2478 1700
rect 2712 1672 2742 1700
rect 3028 1672 3058 1700
rect 3292 1672 3322 1700
rect 3608 1672 3638 1700
rect 3872 1672 3902 1700
rect 4188 1672 4218 1700
rect 4452 1672 4482 1700
rect 4768 1672 4798 1700
rect 5032 1672 5062 1700
rect 5348 1672 5378 1700
rect 5612 1672 5642 1700
rect 5928 1672 5958 1700
rect 6192 1672 6222 1700
rect 6508 1672 6538 1700
rect 6772 1672 6802 1700
rect 128 1402 158 1430
rect 392 1402 422 1430
rect 708 1402 738 1430
rect 972 1402 1002 1430
rect 1288 1402 1318 1430
rect 1552 1402 1582 1430
rect 1868 1402 1898 1430
rect 2132 1402 2162 1430
rect 2448 1402 2478 1430
rect 2712 1402 2742 1430
rect 3028 1402 3058 1430
rect 3292 1402 3322 1430
rect 3608 1402 3638 1430
rect 3872 1402 3902 1430
rect 4188 1402 4218 1430
rect 4452 1402 4482 1430
rect 4768 1402 4798 1430
rect 5032 1402 5062 1430
rect 5348 1402 5378 1430
rect 5612 1402 5642 1430
rect 5928 1402 5958 1430
rect 6192 1402 6222 1430
rect 6508 1402 6538 1430
rect 6772 1402 6802 1430
rect 128 1132 158 1160
rect 392 1132 422 1160
rect 708 1132 738 1160
rect 972 1132 1002 1160
rect 1288 1132 1318 1160
rect 1552 1132 1582 1160
rect 1868 1132 1898 1160
rect 2132 1132 2162 1160
rect 2448 1132 2478 1160
rect 2712 1132 2742 1160
rect 3028 1132 3058 1160
rect 3292 1132 3322 1160
rect 3608 1132 3638 1160
rect 3872 1132 3902 1160
rect 4188 1132 4218 1160
rect 4452 1132 4482 1160
rect 4768 1132 4798 1160
rect 5032 1132 5062 1160
rect 5348 1132 5378 1160
rect 5612 1132 5642 1160
rect 5928 1132 5958 1160
rect 6192 1132 6222 1160
rect 6508 1132 6538 1160
rect 6772 1132 6802 1160
rect 128 862 158 890
rect 392 862 422 890
rect 708 862 738 890
rect 972 862 1002 890
rect 1288 862 1318 890
rect 1552 862 1582 890
rect 1868 862 1898 890
rect 2132 862 2162 890
rect 2448 862 2478 890
rect 2712 862 2742 890
rect 3028 862 3058 890
rect 3292 862 3322 890
rect 3608 862 3638 890
rect 3872 862 3902 890
rect 4188 862 4218 890
rect 4452 862 4482 890
rect 4768 862 4798 890
rect 5032 862 5062 890
rect 5348 862 5378 890
rect 5612 862 5642 890
rect 5928 862 5958 890
rect 6192 862 6222 890
rect 6508 862 6538 890
rect 6772 862 6802 890
rect 128 592 158 620
rect 392 592 422 620
rect 708 592 738 620
rect 972 592 1002 620
rect 1288 592 1318 620
rect 1552 592 1582 620
rect 1868 592 1898 620
rect 2132 592 2162 620
rect 2448 592 2478 620
rect 2712 592 2742 620
rect 3028 592 3058 620
rect 3292 592 3322 620
rect 3608 592 3638 620
rect 3872 592 3902 620
rect 4188 592 4218 620
rect 4452 592 4482 620
rect 4768 592 4798 620
rect 5032 592 5062 620
rect 5348 592 5378 620
rect 5612 592 5642 620
rect 5928 592 5958 620
rect 6192 592 6222 620
rect 6508 592 6538 620
rect 6772 592 6802 620
rect 128 322 158 350
rect 392 322 422 350
rect 708 322 738 350
rect 972 322 1002 350
rect 1288 322 1318 350
rect 1552 322 1582 350
rect 1868 322 1898 350
rect 2132 322 2162 350
rect 2448 322 2478 350
rect 2712 322 2742 350
rect 3028 322 3058 350
rect 3292 322 3322 350
rect 3608 322 3638 350
rect 3872 322 3902 350
rect 4188 322 4218 350
rect 4452 322 4482 350
rect 4768 322 4798 350
rect 5032 322 5062 350
rect 5348 322 5378 350
rect 5612 322 5642 350
rect 5928 322 5958 350
rect 6192 322 6222 350
rect 6508 322 6538 350
rect 6772 322 6802 350
rect 128 52 158 80
rect 392 52 422 80
rect 708 52 738 80
rect 972 52 1002 80
rect 1288 52 1318 80
rect 1552 52 1582 80
rect 1868 52 1898 80
rect 2132 52 2162 80
rect 2448 52 2478 80
rect 2712 52 2742 80
rect 3028 52 3058 80
rect 3292 52 3322 80
rect 3608 52 3638 80
rect 3872 52 3902 80
rect 4188 52 4218 80
rect 4452 52 4482 80
rect 4768 52 4798 80
rect 5032 52 5062 80
rect 5348 52 5378 80
rect 5612 52 5642 80
rect 5928 52 5958 80
rect 6192 52 6222 80
rect 6508 52 6538 80
rect 6772 52 6802 80
rect 128 -218 158 -190
rect 392 -218 422 -190
rect 708 -218 738 -190
rect 972 -218 1002 -190
rect 1288 -218 1318 -190
rect 1552 -218 1582 -190
rect 1868 -218 1898 -190
rect 2132 -218 2162 -190
rect 2448 -218 2478 -190
rect 2712 -218 2742 -190
rect 3028 -218 3058 -190
rect 3292 -218 3322 -190
rect 3608 -218 3638 -190
rect 3872 -218 3902 -190
rect 4188 -218 4218 -190
rect 4452 -218 4482 -190
rect 4768 -218 4798 -190
rect 5032 -218 5062 -190
rect 5348 -218 5378 -190
rect 5612 -218 5642 -190
rect 5928 -218 5958 -190
rect 6192 -218 6222 -190
rect 6508 -218 6538 -190
rect 6772 -218 6802 -190
rect 128 -488 158 -460
rect 392 -488 422 -460
rect 708 -488 738 -460
rect 972 -488 1002 -460
rect 1288 -488 1318 -460
rect 1552 -488 1582 -460
rect 1868 -488 1898 -460
rect 2132 -488 2162 -460
rect 2448 -488 2478 -460
rect 2712 -488 2742 -460
rect 3028 -488 3058 -460
rect 3292 -488 3322 -460
rect 3608 -488 3638 -460
rect 3872 -488 3902 -460
rect 4188 -488 4218 -460
rect 4452 -488 4482 -460
rect 4768 -488 4798 -460
rect 5032 -488 5062 -460
rect 5348 -488 5378 -460
rect 5612 -488 5642 -460
rect 5928 -488 5958 -460
rect 6192 -488 6222 -460
rect 6508 -488 6538 -460
rect 6772 -488 6802 -460
rect 128 -758 158 -730
rect 392 -758 422 -730
rect 708 -758 738 -730
rect 972 -758 1002 -730
rect 1288 -758 1318 -730
rect 1552 -758 1582 -730
rect 1868 -758 1898 -730
rect 2132 -758 2162 -730
rect 2448 -758 2478 -730
rect 2712 -758 2742 -730
rect 3028 -758 3058 -730
rect 3292 -758 3322 -730
rect 3608 -758 3638 -730
rect 3872 -758 3902 -730
rect 4188 -758 4218 -730
rect 4452 -758 4482 -730
rect 4768 -758 4798 -730
rect 5032 -758 5062 -730
rect 5348 -758 5378 -730
rect 5612 -758 5642 -730
rect 5928 -758 5958 -730
rect 6192 -758 6222 -730
rect 6508 -758 6538 -730
rect 6772 -758 6802 -730
rect 128 -1028 158 -1000
rect 392 -1028 422 -1000
rect 708 -1028 738 -1000
rect 972 -1028 1002 -1000
rect 1288 -1028 1318 -1000
rect 1552 -1028 1582 -1000
rect 1868 -1028 1898 -1000
rect 2132 -1028 2162 -1000
rect 2448 -1028 2478 -1000
rect 2712 -1028 2742 -1000
rect 3028 -1028 3058 -1000
rect 3292 -1028 3322 -1000
rect 3608 -1028 3638 -1000
rect 3872 -1028 3902 -1000
rect 4188 -1028 4218 -1000
rect 4452 -1028 4482 -1000
rect 4768 -1028 4798 -1000
rect 5032 -1028 5062 -1000
rect 5348 -1028 5378 -1000
rect 5612 -1028 5642 -1000
rect 5928 -1028 5958 -1000
rect 6192 -1028 6222 -1000
rect 6508 -1028 6538 -1000
rect 6772 -1028 6802 -1000
rect 128 -1298 158 -1270
rect 392 -1298 422 -1270
rect 708 -1298 738 -1270
rect 972 -1298 1002 -1270
rect 1288 -1298 1318 -1270
rect 1552 -1298 1582 -1270
rect 1868 -1298 1898 -1270
rect 2132 -1298 2162 -1270
rect 2448 -1298 2478 -1270
rect 2712 -1298 2742 -1270
rect 3028 -1298 3058 -1270
rect 3292 -1298 3322 -1270
rect 3608 -1298 3638 -1270
rect 3872 -1298 3902 -1270
rect 4188 -1298 4218 -1270
rect 4452 -1298 4482 -1270
rect 4768 -1298 4798 -1270
rect 5032 -1298 5062 -1270
rect 5348 -1298 5378 -1270
rect 5612 -1298 5642 -1270
rect 5928 -1298 5958 -1270
rect 6192 -1298 6222 -1270
rect 6508 -1298 6538 -1270
rect 6772 -1298 6802 -1270
rect 128 -1568 158 -1540
rect 392 -1568 422 -1540
rect 708 -1568 738 -1540
rect 972 -1568 1002 -1540
rect 1288 -1568 1318 -1540
rect 1552 -1568 1582 -1540
rect 1868 -1568 1898 -1540
rect 2132 -1568 2162 -1540
rect 2448 -1568 2478 -1540
rect 2712 -1568 2742 -1540
rect 3028 -1568 3058 -1540
rect 3292 -1568 3322 -1540
rect 3608 -1568 3638 -1540
rect 3872 -1568 3902 -1540
rect 4188 -1568 4218 -1540
rect 4452 -1568 4482 -1540
rect 4768 -1568 4798 -1540
rect 5032 -1568 5062 -1540
rect 5348 -1568 5378 -1540
rect 5612 -1568 5642 -1540
rect 5928 -1568 5958 -1540
rect 6192 -1568 6222 -1540
rect 6508 -1568 6538 -1540
rect 6772 -1568 6802 -1540
rect 128 -1838 158 -1810
rect 392 -1838 422 -1810
rect 708 -1838 738 -1810
rect 972 -1838 1002 -1810
rect 1288 -1838 1318 -1810
rect 1552 -1838 1582 -1810
rect 1868 -1838 1898 -1810
rect 2132 -1838 2162 -1810
rect 2448 -1838 2478 -1810
rect 2712 -1838 2742 -1810
rect 3028 -1838 3058 -1810
rect 3292 -1838 3322 -1810
rect 3608 -1838 3638 -1810
rect 3872 -1838 3902 -1810
rect 4188 -1838 4218 -1810
rect 4452 -1838 4482 -1810
rect 4768 -1838 4798 -1810
rect 5032 -1838 5062 -1810
rect 5348 -1838 5378 -1810
rect 5612 -1838 5642 -1810
rect 5928 -1838 5958 -1810
rect 6192 -1838 6222 -1810
rect 6508 -1838 6538 -1810
rect 6772 -1838 6802 -1810
rect 128 -2108 158 -2080
rect 392 -2108 422 -2080
rect 708 -2108 738 -2080
rect 972 -2108 1002 -2080
rect 1288 -2108 1318 -2080
rect 1552 -2108 1582 -2080
rect 1868 -2108 1898 -2080
rect 2132 -2108 2162 -2080
rect 2448 -2108 2478 -2080
rect 2712 -2108 2742 -2080
rect 3028 -2108 3058 -2080
rect 3292 -2108 3322 -2080
rect 3608 -2108 3638 -2080
rect 3872 -2108 3902 -2080
rect 4188 -2108 4218 -2080
rect 4452 -2108 4482 -2080
rect 4768 -2108 4798 -2080
rect 5032 -2108 5062 -2080
rect 5348 -2108 5378 -2080
rect 5612 -2108 5642 -2080
rect 5928 -2108 5958 -2080
rect 6192 -2108 6222 -2080
rect 6508 -2108 6538 -2080
rect 6772 -2108 6802 -2080
<< ppu >>
rect 221 2078 251 2106
rect 299 2078 329 2106
rect 801 2078 831 2106
rect 879 2078 909 2106
rect 1381 2078 1411 2106
rect 1459 2078 1489 2106
rect 1961 2078 1991 2106
rect 2039 2078 2069 2106
rect 2541 2078 2571 2106
rect 2619 2078 2649 2106
rect 3121 2078 3151 2106
rect 3199 2078 3229 2106
rect 3701 2078 3731 2106
rect 3779 2078 3809 2106
rect 4281 2078 4311 2106
rect 4359 2078 4389 2106
rect 4861 2078 4891 2106
rect 4939 2078 4969 2106
rect 5441 2078 5471 2106
rect 5519 2078 5549 2106
rect 6021 2078 6051 2106
rect 6099 2078 6129 2106
rect 6601 2078 6631 2106
rect 6679 2078 6709 2106
rect 221 1808 251 1836
rect 299 1808 329 1836
rect 801 1808 831 1836
rect 879 1808 909 1836
rect 1381 1808 1411 1836
rect 1459 1808 1489 1836
rect 1961 1808 1991 1836
rect 2039 1808 2069 1836
rect 2541 1808 2571 1836
rect 2619 1808 2649 1836
rect 3121 1808 3151 1836
rect 3199 1808 3229 1836
rect 3701 1808 3731 1836
rect 3779 1808 3809 1836
rect 4281 1808 4311 1836
rect 4359 1808 4389 1836
rect 4861 1808 4891 1836
rect 4939 1808 4969 1836
rect 5441 1808 5471 1836
rect 5519 1808 5549 1836
rect 6021 1808 6051 1836
rect 6099 1808 6129 1836
rect 6601 1808 6631 1836
rect 6679 1808 6709 1836
rect 221 1538 251 1566
rect 299 1538 329 1566
rect 801 1538 831 1566
rect 879 1538 909 1566
rect 1381 1538 1411 1566
rect 1459 1538 1489 1566
rect 1961 1538 1991 1566
rect 2039 1538 2069 1566
rect 2541 1538 2571 1566
rect 2619 1538 2649 1566
rect 3121 1538 3151 1566
rect 3199 1538 3229 1566
rect 3701 1538 3731 1566
rect 3779 1538 3809 1566
rect 4281 1538 4311 1566
rect 4359 1538 4389 1566
rect 4861 1538 4891 1566
rect 4939 1538 4969 1566
rect 5441 1538 5471 1566
rect 5519 1538 5549 1566
rect 6021 1538 6051 1566
rect 6099 1538 6129 1566
rect 6601 1538 6631 1566
rect 6679 1538 6709 1566
rect 221 1268 251 1296
rect 299 1268 329 1296
rect 801 1268 831 1296
rect 879 1268 909 1296
rect 1381 1268 1411 1296
rect 1459 1268 1489 1296
rect 1961 1268 1991 1296
rect 2039 1268 2069 1296
rect 2541 1268 2571 1296
rect 2619 1268 2649 1296
rect 3121 1268 3151 1296
rect 3199 1268 3229 1296
rect 3701 1268 3731 1296
rect 3779 1268 3809 1296
rect 4281 1268 4311 1296
rect 4359 1268 4389 1296
rect 4861 1268 4891 1296
rect 4939 1268 4969 1296
rect 5441 1268 5471 1296
rect 5519 1268 5549 1296
rect 6021 1268 6051 1296
rect 6099 1268 6129 1296
rect 6601 1268 6631 1296
rect 6679 1268 6709 1296
rect 221 998 251 1026
rect 299 998 329 1026
rect 801 998 831 1026
rect 879 998 909 1026
rect 1381 998 1411 1026
rect 1459 998 1489 1026
rect 1961 998 1991 1026
rect 2039 998 2069 1026
rect 2541 998 2571 1026
rect 2619 998 2649 1026
rect 3121 998 3151 1026
rect 3199 998 3229 1026
rect 3701 998 3731 1026
rect 3779 998 3809 1026
rect 4281 998 4311 1026
rect 4359 998 4389 1026
rect 4861 998 4891 1026
rect 4939 998 4969 1026
rect 5441 998 5471 1026
rect 5519 998 5549 1026
rect 6021 998 6051 1026
rect 6099 998 6129 1026
rect 6601 998 6631 1026
rect 6679 998 6709 1026
rect 221 728 251 756
rect 299 728 329 756
rect 801 728 831 756
rect 879 728 909 756
rect 1381 728 1411 756
rect 1459 728 1489 756
rect 1961 728 1991 756
rect 2039 728 2069 756
rect 2541 728 2571 756
rect 2619 728 2649 756
rect 3121 728 3151 756
rect 3199 728 3229 756
rect 3701 728 3731 756
rect 3779 728 3809 756
rect 4281 728 4311 756
rect 4359 728 4389 756
rect 4861 728 4891 756
rect 4939 728 4969 756
rect 5441 728 5471 756
rect 5519 728 5549 756
rect 6021 728 6051 756
rect 6099 728 6129 756
rect 6601 728 6631 756
rect 6679 728 6709 756
rect 221 458 251 486
rect 299 458 329 486
rect 801 458 831 486
rect 879 458 909 486
rect 1381 458 1411 486
rect 1459 458 1489 486
rect 1961 458 1991 486
rect 2039 458 2069 486
rect 2541 458 2571 486
rect 2619 458 2649 486
rect 3121 458 3151 486
rect 3199 458 3229 486
rect 3701 458 3731 486
rect 3779 458 3809 486
rect 4281 458 4311 486
rect 4359 458 4389 486
rect 4861 458 4891 486
rect 4939 458 4969 486
rect 5441 458 5471 486
rect 5519 458 5549 486
rect 6021 458 6051 486
rect 6099 458 6129 486
rect 6601 458 6631 486
rect 6679 458 6709 486
rect 221 188 251 216
rect 299 188 329 216
rect 801 188 831 216
rect 879 188 909 216
rect 1381 188 1411 216
rect 1459 188 1489 216
rect 1961 188 1991 216
rect 2039 188 2069 216
rect 2541 188 2571 216
rect 2619 188 2649 216
rect 3121 188 3151 216
rect 3199 188 3229 216
rect 3701 188 3731 216
rect 3779 188 3809 216
rect 4281 188 4311 216
rect 4359 188 4389 216
rect 4861 188 4891 216
rect 4939 188 4969 216
rect 5441 188 5471 216
rect 5519 188 5549 216
rect 6021 188 6051 216
rect 6099 188 6129 216
rect 6601 188 6631 216
rect 6679 188 6709 216
rect 221 -82 251 -54
rect 299 -82 329 -54
rect 801 -82 831 -54
rect 879 -82 909 -54
rect 1381 -82 1411 -54
rect 1459 -82 1489 -54
rect 1961 -82 1991 -54
rect 2039 -82 2069 -54
rect 2541 -82 2571 -54
rect 2619 -82 2649 -54
rect 3121 -82 3151 -54
rect 3199 -82 3229 -54
rect 3701 -82 3731 -54
rect 3779 -82 3809 -54
rect 4281 -82 4311 -54
rect 4359 -82 4389 -54
rect 4861 -82 4891 -54
rect 4939 -82 4969 -54
rect 5441 -82 5471 -54
rect 5519 -82 5549 -54
rect 6021 -82 6051 -54
rect 6099 -82 6129 -54
rect 6601 -82 6631 -54
rect 6679 -82 6709 -54
rect 221 -352 251 -324
rect 299 -352 329 -324
rect 801 -352 831 -324
rect 879 -352 909 -324
rect 1381 -352 1411 -324
rect 1459 -352 1489 -324
rect 1961 -352 1991 -324
rect 2039 -352 2069 -324
rect 2541 -352 2571 -324
rect 2619 -352 2649 -324
rect 3121 -352 3151 -324
rect 3199 -352 3229 -324
rect 3701 -352 3731 -324
rect 3779 -352 3809 -324
rect 4281 -352 4311 -324
rect 4359 -352 4389 -324
rect 4861 -352 4891 -324
rect 4939 -352 4969 -324
rect 5441 -352 5471 -324
rect 5519 -352 5549 -324
rect 6021 -352 6051 -324
rect 6099 -352 6129 -324
rect 6601 -352 6631 -324
rect 6679 -352 6709 -324
rect 221 -622 251 -594
rect 299 -622 329 -594
rect 801 -622 831 -594
rect 879 -622 909 -594
rect 1381 -622 1411 -594
rect 1459 -622 1489 -594
rect 1961 -622 1991 -594
rect 2039 -622 2069 -594
rect 2541 -622 2571 -594
rect 2619 -622 2649 -594
rect 3121 -622 3151 -594
rect 3199 -622 3229 -594
rect 3701 -622 3731 -594
rect 3779 -622 3809 -594
rect 4281 -622 4311 -594
rect 4359 -622 4389 -594
rect 4861 -622 4891 -594
rect 4939 -622 4969 -594
rect 5441 -622 5471 -594
rect 5519 -622 5549 -594
rect 6021 -622 6051 -594
rect 6099 -622 6129 -594
rect 6601 -622 6631 -594
rect 6679 -622 6709 -594
rect 221 -892 251 -864
rect 299 -892 329 -864
rect 801 -892 831 -864
rect 879 -892 909 -864
rect 1381 -892 1411 -864
rect 1459 -892 1489 -864
rect 1961 -892 1991 -864
rect 2039 -892 2069 -864
rect 2541 -892 2571 -864
rect 2619 -892 2649 -864
rect 3121 -892 3151 -864
rect 3199 -892 3229 -864
rect 3701 -892 3731 -864
rect 3779 -892 3809 -864
rect 4281 -892 4311 -864
rect 4359 -892 4389 -864
rect 4861 -892 4891 -864
rect 4939 -892 4969 -864
rect 5441 -892 5471 -864
rect 5519 -892 5549 -864
rect 6021 -892 6051 -864
rect 6099 -892 6129 -864
rect 6601 -892 6631 -864
rect 6679 -892 6709 -864
rect 221 -1162 251 -1134
rect 299 -1162 329 -1134
rect 801 -1162 831 -1134
rect 879 -1162 909 -1134
rect 1381 -1162 1411 -1134
rect 1459 -1162 1489 -1134
rect 1961 -1162 1991 -1134
rect 2039 -1162 2069 -1134
rect 2541 -1162 2571 -1134
rect 2619 -1162 2649 -1134
rect 3121 -1162 3151 -1134
rect 3199 -1162 3229 -1134
rect 3701 -1162 3731 -1134
rect 3779 -1162 3809 -1134
rect 4281 -1162 4311 -1134
rect 4359 -1162 4389 -1134
rect 4861 -1162 4891 -1134
rect 4939 -1162 4969 -1134
rect 5441 -1162 5471 -1134
rect 5519 -1162 5549 -1134
rect 6021 -1162 6051 -1134
rect 6099 -1162 6129 -1134
rect 6601 -1162 6631 -1134
rect 6679 -1162 6709 -1134
rect 221 -1432 251 -1404
rect 299 -1432 329 -1404
rect 801 -1432 831 -1404
rect 879 -1432 909 -1404
rect 1381 -1432 1411 -1404
rect 1459 -1432 1489 -1404
rect 1961 -1432 1991 -1404
rect 2039 -1432 2069 -1404
rect 2541 -1432 2571 -1404
rect 2619 -1432 2649 -1404
rect 3121 -1432 3151 -1404
rect 3199 -1432 3229 -1404
rect 3701 -1432 3731 -1404
rect 3779 -1432 3809 -1404
rect 4281 -1432 4311 -1404
rect 4359 -1432 4389 -1404
rect 4861 -1432 4891 -1404
rect 4939 -1432 4969 -1404
rect 5441 -1432 5471 -1404
rect 5519 -1432 5549 -1404
rect 6021 -1432 6051 -1404
rect 6099 -1432 6129 -1404
rect 6601 -1432 6631 -1404
rect 6679 -1432 6709 -1404
rect 221 -1702 251 -1674
rect 299 -1702 329 -1674
rect 801 -1702 831 -1674
rect 879 -1702 909 -1674
rect 1381 -1702 1411 -1674
rect 1459 -1702 1489 -1674
rect 1961 -1702 1991 -1674
rect 2039 -1702 2069 -1674
rect 2541 -1702 2571 -1674
rect 2619 -1702 2649 -1674
rect 3121 -1702 3151 -1674
rect 3199 -1702 3229 -1674
rect 3701 -1702 3731 -1674
rect 3779 -1702 3809 -1674
rect 4281 -1702 4311 -1674
rect 4359 -1702 4389 -1674
rect 4861 -1702 4891 -1674
rect 4939 -1702 4969 -1674
rect 5441 -1702 5471 -1674
rect 5519 -1702 5549 -1674
rect 6021 -1702 6051 -1674
rect 6099 -1702 6129 -1674
rect 6601 -1702 6631 -1674
rect 6679 -1702 6709 -1674
rect 221 -1972 251 -1944
rect 299 -1972 329 -1944
rect 801 -1972 831 -1944
rect 879 -1972 909 -1944
rect 1381 -1972 1411 -1944
rect 1459 -1972 1489 -1944
rect 1961 -1972 1991 -1944
rect 2039 -1972 2069 -1944
rect 2541 -1972 2571 -1944
rect 2619 -1972 2649 -1944
rect 3121 -1972 3151 -1944
rect 3199 -1972 3229 -1944
rect 3701 -1972 3731 -1944
rect 3779 -1972 3809 -1944
rect 4281 -1972 4311 -1944
rect 4359 -1972 4389 -1944
rect 4861 -1972 4891 -1944
rect 4939 -1972 4969 -1944
rect 5441 -1972 5471 -1944
rect 5519 -1972 5549 -1944
rect 6021 -1972 6051 -1944
rect 6099 -1972 6129 -1944
rect 6601 -1972 6631 -1944
rect 6679 -1972 6709 -1944
<< ndiff >>
rect 88 2088 106 2116
rect 136 2088 154 2116
rect 396 2088 414 2116
rect 444 2088 463 2116
rect 668 2088 686 2116
rect 716 2088 734 2116
rect 976 2088 994 2116
rect 1024 2088 1043 2116
rect 1248 2088 1266 2116
rect 1296 2088 1314 2116
rect 1556 2088 1574 2116
rect 1604 2088 1623 2116
rect 1828 2088 1846 2116
rect 1876 2088 1894 2116
rect 2136 2088 2154 2116
rect 2184 2088 2203 2116
rect 2408 2088 2426 2116
rect 2456 2088 2474 2116
rect 2716 2088 2734 2116
rect 2764 2088 2783 2116
rect 2988 2088 3006 2116
rect 3036 2088 3054 2116
rect 3296 2088 3314 2116
rect 3344 2088 3363 2116
rect 3568 2088 3586 2116
rect 3616 2088 3634 2116
rect 3876 2088 3894 2116
rect 3924 2088 3943 2116
rect 4148 2088 4166 2116
rect 4196 2088 4214 2116
rect 4456 2088 4474 2116
rect 4504 2088 4523 2116
rect 4728 2088 4746 2116
rect 4776 2088 4794 2116
rect 5036 2088 5054 2116
rect 5084 2088 5103 2116
rect 5308 2088 5326 2116
rect 5356 2088 5374 2116
rect 5616 2088 5634 2116
rect 5664 2088 5683 2116
rect 5888 2088 5906 2116
rect 5936 2088 5954 2116
rect 6196 2088 6214 2116
rect 6244 2088 6263 2116
rect 6468 2088 6486 2116
rect 6516 2088 6534 2116
rect 6776 2088 6794 2116
rect 6824 2088 6843 2116
rect 14 1942 42 1984
rect 72 1970 97 1984
rect 196 1974 221 1984
rect 72 1942 128 1970
rect 158 1942 192 1970
tri 206 1967 213 1974 ne
rect 213 1942 221 1974
rect 251 1942 299 1984
rect 329 1974 354 1984
rect 329 1942 337 1974
rect 453 1970 478 1984
rect 358 1942 392 1970
rect 422 1942 478 1970
rect 508 1942 536 1984
rect 594 1942 622 1984
rect 652 1970 677 1984
rect 776 1974 801 1984
rect 652 1942 708 1970
rect 738 1942 772 1970
tri 786 1967 793 1974 ne
rect 793 1942 801 1974
rect 831 1942 879 1984
rect 909 1974 934 1984
rect 909 1942 917 1974
rect 1033 1970 1058 1984
rect 938 1942 972 1970
rect 1002 1942 1058 1970
rect 1088 1942 1116 1984
rect 1174 1942 1202 1984
rect 1232 1970 1257 1984
rect 1356 1974 1381 1984
rect 1232 1942 1288 1970
rect 1318 1942 1352 1970
tri 1366 1967 1373 1974 ne
rect 1373 1942 1381 1974
rect 1411 1942 1459 1984
rect 1489 1974 1514 1984
rect 1489 1942 1497 1974
rect 1613 1970 1638 1984
rect 1518 1942 1552 1970
rect 1582 1942 1638 1970
rect 1668 1942 1696 1984
rect 1754 1942 1782 1984
rect 1812 1970 1837 1984
rect 1936 1974 1961 1984
rect 1812 1942 1868 1970
rect 1898 1942 1932 1970
tri 1946 1967 1953 1974 ne
rect 1953 1942 1961 1974
rect 1991 1942 2039 1984
rect 2069 1974 2094 1984
rect 2069 1942 2077 1974
rect 2193 1970 2218 1984
rect 2098 1942 2132 1970
rect 2162 1942 2218 1970
rect 2248 1942 2276 1984
rect 2334 1942 2362 1984
rect 2392 1970 2417 1984
rect 2516 1974 2541 1984
rect 2392 1942 2448 1970
rect 2478 1942 2512 1970
tri 2526 1967 2533 1974 ne
rect 2533 1942 2541 1974
rect 2571 1942 2619 1984
rect 2649 1974 2674 1984
rect 2649 1942 2657 1974
rect 2773 1970 2798 1984
rect 2678 1942 2712 1970
rect 2742 1942 2798 1970
rect 2828 1942 2856 1984
rect 2914 1942 2942 1984
rect 2972 1970 2997 1984
rect 3096 1974 3121 1984
rect 2972 1942 3028 1970
rect 3058 1942 3092 1970
tri 3106 1967 3113 1974 ne
rect 3113 1942 3121 1974
rect 3151 1942 3199 1984
rect 3229 1974 3254 1984
rect 3229 1942 3237 1974
rect 3353 1970 3378 1984
rect 3258 1942 3292 1970
rect 3322 1942 3378 1970
rect 3408 1942 3436 1984
rect 3494 1942 3522 1984
rect 3552 1970 3577 1984
rect 3676 1974 3701 1984
rect 3552 1942 3608 1970
rect 3638 1942 3672 1970
tri 3686 1967 3693 1974 ne
rect 3693 1942 3701 1974
rect 3731 1942 3779 1984
rect 3809 1974 3834 1984
rect 3809 1942 3817 1974
rect 3933 1970 3958 1984
rect 3838 1942 3872 1970
rect 3902 1942 3958 1970
rect 3988 1942 4016 1984
rect 4074 1942 4102 1984
rect 4132 1970 4157 1984
rect 4256 1974 4281 1984
rect 4132 1942 4188 1970
rect 4218 1942 4252 1970
tri 4266 1967 4273 1974 ne
rect 4273 1942 4281 1974
rect 4311 1942 4359 1984
rect 4389 1974 4414 1984
rect 4389 1942 4397 1974
rect 4513 1970 4538 1984
rect 4418 1942 4452 1970
rect 4482 1942 4538 1970
rect 4568 1942 4596 1984
rect 4654 1942 4682 1984
rect 4712 1970 4737 1984
rect 4836 1974 4861 1984
rect 4712 1942 4768 1970
rect 4798 1942 4832 1970
tri 4846 1967 4853 1974 ne
rect 4853 1942 4861 1974
rect 4891 1942 4939 1984
rect 4969 1974 4994 1984
rect 4969 1942 4977 1974
rect 5093 1970 5118 1984
rect 4998 1942 5032 1970
rect 5062 1942 5118 1970
rect 5148 1942 5176 1984
rect 5234 1942 5262 1984
rect 5292 1970 5317 1984
rect 5416 1974 5441 1984
rect 5292 1942 5348 1970
rect 5378 1942 5412 1970
tri 5426 1967 5433 1974 ne
rect 5433 1942 5441 1974
rect 5471 1942 5519 1984
rect 5549 1974 5574 1984
rect 5549 1942 5557 1974
rect 5673 1970 5698 1984
rect 5578 1942 5612 1970
rect 5642 1942 5698 1970
rect 5728 1942 5756 1984
rect 5814 1942 5842 1984
rect 5872 1970 5897 1984
rect 5996 1974 6021 1984
rect 5872 1942 5928 1970
rect 5958 1942 5992 1970
tri 6006 1967 6013 1974 ne
rect 6013 1942 6021 1974
rect 6051 1942 6099 1984
rect 6129 1974 6154 1984
rect 6129 1942 6137 1974
rect 6253 1970 6278 1984
rect 6158 1942 6192 1970
rect 6222 1942 6278 1970
rect 6308 1942 6336 1984
rect 6394 1942 6422 1984
rect 6452 1970 6477 1984
rect 6576 1974 6601 1984
rect 6452 1942 6508 1970
rect 6538 1942 6572 1970
tri 6586 1967 6593 1974 ne
rect 6593 1942 6601 1974
rect 6631 1942 6679 1984
rect 6709 1974 6734 1984
rect 6709 1942 6717 1974
rect 6833 1970 6858 1984
rect 6738 1942 6772 1970
rect 6802 1942 6858 1970
rect 6888 1942 6916 1984
rect 165 1918 192 1942
rect 259 1920 291 1942
rect 259 1918 261 1920
rect 289 1918 291 1920
rect 358 1918 385 1942
rect 165 1904 259 1918
rect 291 1904 385 1918
rect 745 1918 772 1942
rect 839 1920 871 1942
rect 839 1918 841 1920
rect 869 1918 871 1920
rect 938 1918 965 1942
rect 745 1904 839 1918
rect 871 1904 965 1918
rect 1325 1918 1352 1942
rect 1419 1920 1451 1942
rect 1419 1918 1421 1920
rect 1449 1918 1451 1920
rect 1518 1918 1545 1942
rect 1325 1904 1419 1918
rect 1451 1904 1545 1918
rect 1905 1918 1932 1942
rect 1999 1920 2031 1942
rect 1999 1918 2001 1920
rect 2029 1918 2031 1920
rect 2098 1918 2125 1942
rect 1905 1904 1999 1918
rect 2031 1904 2125 1918
rect 2485 1918 2512 1942
rect 2579 1920 2611 1942
rect 2579 1918 2581 1920
rect 2609 1918 2611 1920
rect 2678 1918 2705 1942
rect 2485 1904 2579 1918
rect 2611 1904 2705 1918
rect 3065 1918 3092 1942
rect 3159 1920 3191 1942
rect 3159 1918 3161 1920
rect 3189 1918 3191 1920
rect 3258 1918 3285 1942
rect 3065 1904 3159 1918
rect 3191 1904 3285 1918
rect 3645 1918 3672 1942
rect 3739 1920 3771 1942
rect 3739 1918 3741 1920
rect 3769 1918 3771 1920
rect 3838 1918 3865 1942
rect 3645 1904 3739 1918
rect 3771 1904 3865 1918
rect 4225 1918 4252 1942
rect 4319 1920 4351 1942
rect 4319 1918 4321 1920
rect 4349 1918 4351 1920
rect 4418 1918 4445 1942
rect 4225 1904 4319 1918
rect 4351 1904 4445 1918
rect 4805 1918 4832 1942
rect 4899 1920 4931 1942
rect 4899 1918 4901 1920
rect 4929 1918 4931 1920
rect 4998 1918 5025 1942
rect 4805 1904 4899 1918
rect 4931 1904 5025 1918
rect 5385 1918 5412 1942
rect 5479 1920 5511 1942
rect 5479 1918 5481 1920
rect 5509 1918 5511 1920
rect 5578 1918 5605 1942
rect 5385 1904 5479 1918
rect 5511 1904 5605 1918
rect 5965 1918 5992 1942
rect 6059 1920 6091 1942
rect 6059 1918 6061 1920
rect 6089 1918 6091 1920
rect 6158 1918 6185 1942
rect 5965 1904 6059 1918
rect 6091 1904 6185 1918
rect 6545 1918 6572 1942
rect 6639 1920 6671 1942
rect 6639 1918 6641 1920
rect 6669 1918 6671 1920
rect 6738 1918 6765 1942
rect 6545 1904 6639 1918
rect 6671 1904 6765 1918
rect 88 1818 106 1846
rect 136 1818 154 1846
rect 396 1818 414 1846
rect 444 1818 463 1846
rect 668 1818 686 1846
rect 716 1818 734 1846
rect 976 1818 994 1846
rect 1024 1818 1043 1846
rect 1248 1818 1266 1846
rect 1296 1818 1314 1846
rect 1556 1818 1574 1846
rect 1604 1818 1623 1846
rect 1828 1818 1846 1846
rect 1876 1818 1894 1846
rect 2136 1818 2154 1846
rect 2184 1818 2203 1846
rect 2408 1818 2426 1846
rect 2456 1818 2474 1846
rect 2716 1818 2734 1846
rect 2764 1818 2783 1846
rect 2988 1818 3006 1846
rect 3036 1818 3054 1846
rect 3296 1818 3314 1846
rect 3344 1818 3363 1846
rect 3568 1818 3586 1846
rect 3616 1818 3634 1846
rect 3876 1818 3894 1846
rect 3924 1818 3943 1846
rect 4148 1818 4166 1846
rect 4196 1818 4214 1846
rect 4456 1818 4474 1846
rect 4504 1818 4523 1846
rect 4728 1818 4746 1846
rect 4776 1818 4794 1846
rect 5036 1818 5054 1846
rect 5084 1818 5103 1846
rect 5308 1818 5326 1846
rect 5356 1818 5374 1846
rect 5616 1818 5634 1846
rect 5664 1818 5683 1846
rect 5888 1818 5906 1846
rect 5936 1818 5954 1846
rect 6196 1818 6214 1846
rect 6244 1818 6263 1846
rect 6468 1818 6486 1846
rect 6516 1818 6534 1846
rect 6776 1818 6794 1846
rect 6824 1818 6843 1846
rect 14 1672 42 1714
rect 72 1700 97 1714
rect 196 1704 221 1714
rect 72 1672 128 1700
rect 158 1672 192 1700
tri 206 1697 213 1704 ne
rect 213 1672 221 1704
rect 251 1672 299 1714
rect 329 1704 354 1714
rect 329 1672 337 1704
rect 453 1700 478 1714
rect 358 1672 392 1700
rect 422 1672 478 1700
rect 508 1672 536 1714
rect 594 1672 622 1714
rect 652 1700 677 1714
rect 776 1704 801 1714
rect 652 1672 708 1700
rect 738 1672 772 1700
tri 786 1697 793 1704 ne
rect 793 1672 801 1704
rect 831 1672 879 1714
rect 909 1704 934 1714
rect 909 1672 917 1704
rect 1033 1700 1058 1714
rect 938 1672 972 1700
rect 1002 1672 1058 1700
rect 1088 1672 1116 1714
rect 1174 1672 1202 1714
rect 1232 1700 1257 1714
rect 1356 1704 1381 1714
rect 1232 1672 1288 1700
rect 1318 1672 1352 1700
tri 1366 1697 1373 1704 ne
rect 1373 1672 1381 1704
rect 1411 1672 1459 1714
rect 1489 1704 1514 1714
rect 1489 1672 1497 1704
rect 1613 1700 1638 1714
rect 1518 1672 1552 1700
rect 1582 1672 1638 1700
rect 1668 1672 1696 1714
rect 1754 1672 1782 1714
rect 1812 1700 1837 1714
rect 1936 1704 1961 1714
rect 1812 1672 1868 1700
rect 1898 1672 1932 1700
tri 1946 1697 1953 1704 ne
rect 1953 1672 1961 1704
rect 1991 1672 2039 1714
rect 2069 1704 2094 1714
rect 2069 1672 2077 1704
rect 2193 1700 2218 1714
rect 2098 1672 2132 1700
rect 2162 1672 2218 1700
rect 2248 1672 2276 1714
rect 2334 1672 2362 1714
rect 2392 1700 2417 1714
rect 2516 1704 2541 1714
rect 2392 1672 2448 1700
rect 2478 1672 2512 1700
tri 2526 1697 2533 1704 ne
rect 2533 1672 2541 1704
rect 2571 1672 2619 1714
rect 2649 1704 2674 1714
rect 2649 1672 2657 1704
rect 2773 1700 2798 1714
rect 2678 1672 2712 1700
rect 2742 1672 2798 1700
rect 2828 1672 2856 1714
rect 2914 1672 2942 1714
rect 2972 1700 2997 1714
rect 3096 1704 3121 1714
rect 2972 1672 3028 1700
rect 3058 1672 3092 1700
tri 3106 1697 3113 1704 ne
rect 3113 1672 3121 1704
rect 3151 1672 3199 1714
rect 3229 1704 3254 1714
rect 3229 1672 3237 1704
rect 3353 1700 3378 1714
rect 3258 1672 3292 1700
rect 3322 1672 3378 1700
rect 3408 1672 3436 1714
rect 3494 1672 3522 1714
rect 3552 1700 3577 1714
rect 3676 1704 3701 1714
rect 3552 1672 3608 1700
rect 3638 1672 3672 1700
tri 3686 1697 3693 1704 ne
rect 3693 1672 3701 1704
rect 3731 1672 3779 1714
rect 3809 1704 3834 1714
rect 3809 1672 3817 1704
rect 3933 1700 3958 1714
rect 3838 1672 3872 1700
rect 3902 1672 3958 1700
rect 3988 1672 4016 1714
rect 4074 1672 4102 1714
rect 4132 1700 4157 1714
rect 4256 1704 4281 1714
rect 4132 1672 4188 1700
rect 4218 1672 4252 1700
tri 4266 1697 4273 1704 ne
rect 4273 1672 4281 1704
rect 4311 1672 4359 1714
rect 4389 1704 4414 1714
rect 4389 1672 4397 1704
rect 4513 1700 4538 1714
rect 4418 1672 4452 1700
rect 4482 1672 4538 1700
rect 4568 1672 4596 1714
rect 4654 1672 4682 1714
rect 4712 1700 4737 1714
rect 4836 1704 4861 1714
rect 4712 1672 4768 1700
rect 4798 1672 4832 1700
tri 4846 1697 4853 1704 ne
rect 4853 1672 4861 1704
rect 4891 1672 4939 1714
rect 4969 1704 4994 1714
rect 4969 1672 4977 1704
rect 5093 1700 5118 1714
rect 4998 1672 5032 1700
rect 5062 1672 5118 1700
rect 5148 1672 5176 1714
rect 5234 1672 5262 1714
rect 5292 1700 5317 1714
rect 5416 1704 5441 1714
rect 5292 1672 5348 1700
rect 5378 1672 5412 1700
tri 5426 1697 5433 1704 ne
rect 5433 1672 5441 1704
rect 5471 1672 5519 1714
rect 5549 1704 5574 1714
rect 5549 1672 5557 1704
rect 5673 1700 5698 1714
rect 5578 1672 5612 1700
rect 5642 1672 5698 1700
rect 5728 1672 5756 1714
rect 5814 1672 5842 1714
rect 5872 1700 5897 1714
rect 5996 1704 6021 1714
rect 5872 1672 5928 1700
rect 5958 1672 5992 1700
tri 6006 1697 6013 1704 ne
rect 6013 1672 6021 1704
rect 6051 1672 6099 1714
rect 6129 1704 6154 1714
rect 6129 1672 6137 1704
rect 6253 1700 6278 1714
rect 6158 1672 6192 1700
rect 6222 1672 6278 1700
rect 6308 1672 6336 1714
rect 6394 1672 6422 1714
rect 6452 1700 6477 1714
rect 6576 1704 6601 1714
rect 6452 1672 6508 1700
rect 6538 1672 6572 1700
tri 6586 1697 6593 1704 ne
rect 6593 1672 6601 1704
rect 6631 1672 6679 1714
rect 6709 1704 6734 1714
rect 6709 1672 6717 1704
rect 6833 1700 6858 1714
rect 6738 1672 6772 1700
rect 6802 1672 6858 1700
rect 6888 1672 6916 1714
rect 165 1648 192 1672
rect 259 1650 291 1672
rect 259 1648 261 1650
rect 289 1648 291 1650
rect 358 1648 385 1672
rect 165 1634 259 1648
rect 291 1634 385 1648
rect 745 1648 772 1672
rect 839 1650 871 1672
rect 839 1648 841 1650
rect 869 1648 871 1650
rect 938 1648 965 1672
rect 745 1634 839 1648
rect 871 1634 965 1648
rect 1325 1648 1352 1672
rect 1419 1650 1451 1672
rect 1419 1648 1421 1650
rect 1449 1648 1451 1650
rect 1518 1648 1545 1672
rect 1325 1634 1419 1648
rect 1451 1634 1545 1648
rect 1905 1648 1932 1672
rect 1999 1650 2031 1672
rect 1999 1648 2001 1650
rect 2029 1648 2031 1650
rect 2098 1648 2125 1672
rect 1905 1634 1999 1648
rect 2031 1634 2125 1648
rect 2485 1648 2512 1672
rect 2579 1650 2611 1672
rect 2579 1648 2581 1650
rect 2609 1648 2611 1650
rect 2678 1648 2705 1672
rect 2485 1634 2579 1648
rect 2611 1634 2705 1648
rect 3065 1648 3092 1672
rect 3159 1650 3191 1672
rect 3159 1648 3161 1650
rect 3189 1648 3191 1650
rect 3258 1648 3285 1672
rect 3065 1634 3159 1648
rect 3191 1634 3285 1648
rect 3645 1648 3672 1672
rect 3739 1650 3771 1672
rect 3739 1648 3741 1650
rect 3769 1648 3771 1650
rect 3838 1648 3865 1672
rect 3645 1634 3739 1648
rect 3771 1634 3865 1648
rect 4225 1648 4252 1672
rect 4319 1650 4351 1672
rect 4319 1648 4321 1650
rect 4349 1648 4351 1650
rect 4418 1648 4445 1672
rect 4225 1634 4319 1648
rect 4351 1634 4445 1648
rect 4805 1648 4832 1672
rect 4899 1650 4931 1672
rect 4899 1648 4901 1650
rect 4929 1648 4931 1650
rect 4998 1648 5025 1672
rect 4805 1634 4899 1648
rect 4931 1634 5025 1648
rect 5385 1648 5412 1672
rect 5479 1650 5511 1672
rect 5479 1648 5481 1650
rect 5509 1648 5511 1650
rect 5578 1648 5605 1672
rect 5385 1634 5479 1648
rect 5511 1634 5605 1648
rect 5965 1648 5992 1672
rect 6059 1650 6091 1672
rect 6059 1648 6061 1650
rect 6089 1648 6091 1650
rect 6158 1648 6185 1672
rect 5965 1634 6059 1648
rect 6091 1634 6185 1648
rect 6545 1648 6572 1672
rect 6639 1650 6671 1672
rect 6639 1648 6641 1650
rect 6669 1648 6671 1650
rect 6738 1648 6765 1672
rect 6545 1634 6639 1648
rect 6671 1634 6765 1648
rect 88 1548 106 1576
rect 136 1548 154 1576
rect 396 1548 414 1576
rect 444 1548 463 1576
rect 668 1548 686 1576
rect 716 1548 734 1576
rect 976 1548 994 1576
rect 1024 1548 1043 1576
rect 1248 1548 1266 1576
rect 1296 1548 1314 1576
rect 1556 1548 1574 1576
rect 1604 1548 1623 1576
rect 1828 1548 1846 1576
rect 1876 1548 1894 1576
rect 2136 1548 2154 1576
rect 2184 1548 2203 1576
rect 2408 1548 2426 1576
rect 2456 1548 2474 1576
rect 2716 1548 2734 1576
rect 2764 1548 2783 1576
rect 2988 1548 3006 1576
rect 3036 1548 3054 1576
rect 3296 1548 3314 1576
rect 3344 1548 3363 1576
rect 3568 1548 3586 1576
rect 3616 1548 3634 1576
rect 3876 1548 3894 1576
rect 3924 1548 3943 1576
rect 4148 1548 4166 1576
rect 4196 1548 4214 1576
rect 4456 1548 4474 1576
rect 4504 1548 4523 1576
rect 4728 1548 4746 1576
rect 4776 1548 4794 1576
rect 5036 1548 5054 1576
rect 5084 1548 5103 1576
rect 5308 1548 5326 1576
rect 5356 1548 5374 1576
rect 5616 1548 5634 1576
rect 5664 1548 5683 1576
rect 5888 1548 5906 1576
rect 5936 1548 5954 1576
rect 6196 1548 6214 1576
rect 6244 1548 6263 1576
rect 6468 1548 6486 1576
rect 6516 1548 6534 1576
rect 6776 1548 6794 1576
rect 6824 1548 6843 1576
rect 14 1402 42 1444
rect 72 1430 97 1444
rect 196 1434 221 1444
rect 72 1402 128 1430
rect 158 1402 192 1430
tri 206 1427 213 1434 ne
rect 213 1402 221 1434
rect 251 1402 299 1444
rect 329 1434 354 1444
rect 329 1402 337 1434
rect 453 1430 478 1444
rect 358 1402 392 1430
rect 422 1402 478 1430
rect 508 1402 536 1444
rect 594 1402 622 1444
rect 652 1430 677 1444
rect 776 1434 801 1444
rect 652 1402 708 1430
rect 738 1402 772 1430
tri 786 1427 793 1434 ne
rect 793 1402 801 1434
rect 831 1402 879 1444
rect 909 1434 934 1444
rect 909 1402 917 1434
rect 1033 1430 1058 1444
rect 938 1402 972 1430
rect 1002 1402 1058 1430
rect 1088 1402 1116 1444
rect 1174 1402 1202 1444
rect 1232 1430 1257 1444
rect 1356 1434 1381 1444
rect 1232 1402 1288 1430
rect 1318 1402 1352 1430
tri 1366 1427 1373 1434 ne
rect 1373 1402 1381 1434
rect 1411 1402 1459 1444
rect 1489 1434 1514 1444
rect 1489 1402 1497 1434
rect 1613 1430 1638 1444
rect 1518 1402 1552 1430
rect 1582 1402 1638 1430
rect 1668 1402 1696 1444
rect 1754 1402 1782 1444
rect 1812 1430 1837 1444
rect 1936 1434 1961 1444
rect 1812 1402 1868 1430
rect 1898 1402 1932 1430
tri 1946 1427 1953 1434 ne
rect 1953 1402 1961 1434
rect 1991 1402 2039 1444
rect 2069 1434 2094 1444
rect 2069 1402 2077 1434
rect 2193 1430 2218 1444
rect 2098 1402 2132 1430
rect 2162 1402 2218 1430
rect 2248 1402 2276 1444
rect 2334 1402 2362 1444
rect 2392 1430 2417 1444
rect 2516 1434 2541 1444
rect 2392 1402 2448 1430
rect 2478 1402 2512 1430
tri 2526 1427 2533 1434 ne
rect 2533 1402 2541 1434
rect 2571 1402 2619 1444
rect 2649 1434 2674 1444
rect 2649 1402 2657 1434
rect 2773 1430 2798 1444
rect 2678 1402 2712 1430
rect 2742 1402 2798 1430
rect 2828 1402 2856 1444
rect 2914 1402 2942 1444
rect 2972 1430 2997 1444
rect 3096 1434 3121 1444
rect 2972 1402 3028 1430
rect 3058 1402 3092 1430
tri 3106 1427 3113 1434 ne
rect 3113 1402 3121 1434
rect 3151 1402 3199 1444
rect 3229 1434 3254 1444
rect 3229 1402 3237 1434
rect 3353 1430 3378 1444
rect 3258 1402 3292 1430
rect 3322 1402 3378 1430
rect 3408 1402 3436 1444
rect 3494 1402 3522 1444
rect 3552 1430 3577 1444
rect 3676 1434 3701 1444
rect 3552 1402 3608 1430
rect 3638 1402 3672 1430
tri 3686 1427 3693 1434 ne
rect 3693 1402 3701 1434
rect 3731 1402 3779 1444
rect 3809 1434 3834 1444
rect 3809 1402 3817 1434
rect 3933 1430 3958 1444
rect 3838 1402 3872 1430
rect 3902 1402 3958 1430
rect 3988 1402 4016 1444
rect 4074 1402 4102 1444
rect 4132 1430 4157 1444
rect 4256 1434 4281 1444
rect 4132 1402 4188 1430
rect 4218 1402 4252 1430
tri 4266 1427 4273 1434 ne
rect 4273 1402 4281 1434
rect 4311 1402 4359 1444
rect 4389 1434 4414 1444
rect 4389 1402 4397 1434
rect 4513 1430 4538 1444
rect 4418 1402 4452 1430
rect 4482 1402 4538 1430
rect 4568 1402 4596 1444
rect 4654 1402 4682 1444
rect 4712 1430 4737 1444
rect 4836 1434 4861 1444
rect 4712 1402 4768 1430
rect 4798 1402 4832 1430
tri 4846 1427 4853 1434 ne
rect 4853 1402 4861 1434
rect 4891 1402 4939 1444
rect 4969 1434 4994 1444
rect 4969 1402 4977 1434
rect 5093 1430 5118 1444
rect 4998 1402 5032 1430
rect 5062 1402 5118 1430
rect 5148 1402 5176 1444
rect 5234 1402 5262 1444
rect 5292 1430 5317 1444
rect 5416 1434 5441 1444
rect 5292 1402 5348 1430
rect 5378 1402 5412 1430
tri 5426 1427 5433 1434 ne
rect 5433 1402 5441 1434
rect 5471 1402 5519 1444
rect 5549 1434 5574 1444
rect 5549 1402 5557 1434
rect 5673 1430 5698 1444
rect 5578 1402 5612 1430
rect 5642 1402 5698 1430
rect 5728 1402 5756 1444
rect 5814 1402 5842 1444
rect 5872 1430 5897 1444
rect 5996 1434 6021 1444
rect 5872 1402 5928 1430
rect 5958 1402 5992 1430
tri 6006 1427 6013 1434 ne
rect 6013 1402 6021 1434
rect 6051 1402 6099 1444
rect 6129 1434 6154 1444
rect 6129 1402 6137 1434
rect 6253 1430 6278 1444
rect 6158 1402 6192 1430
rect 6222 1402 6278 1430
rect 6308 1402 6336 1444
rect 6394 1402 6422 1444
rect 6452 1430 6477 1444
rect 6576 1434 6601 1444
rect 6452 1402 6508 1430
rect 6538 1402 6572 1430
tri 6586 1427 6593 1434 ne
rect 6593 1402 6601 1434
rect 6631 1402 6679 1444
rect 6709 1434 6734 1444
rect 6709 1402 6717 1434
rect 6833 1430 6858 1444
rect 6738 1402 6772 1430
rect 6802 1402 6858 1430
rect 6888 1402 6916 1444
rect 165 1378 192 1402
rect 259 1380 291 1402
rect 259 1378 261 1380
rect 289 1378 291 1380
rect 358 1378 385 1402
rect 165 1364 259 1378
rect 291 1364 385 1378
rect 745 1378 772 1402
rect 839 1380 871 1402
rect 839 1378 841 1380
rect 869 1378 871 1380
rect 938 1378 965 1402
rect 745 1364 839 1378
rect 871 1364 965 1378
rect 1325 1378 1352 1402
rect 1419 1380 1451 1402
rect 1419 1378 1421 1380
rect 1449 1378 1451 1380
rect 1518 1378 1545 1402
rect 1325 1364 1419 1378
rect 1451 1364 1545 1378
rect 1905 1378 1932 1402
rect 1999 1380 2031 1402
rect 1999 1378 2001 1380
rect 2029 1378 2031 1380
rect 2098 1378 2125 1402
rect 1905 1364 1999 1378
rect 2031 1364 2125 1378
rect 2485 1378 2512 1402
rect 2579 1380 2611 1402
rect 2579 1378 2581 1380
rect 2609 1378 2611 1380
rect 2678 1378 2705 1402
rect 2485 1364 2579 1378
rect 2611 1364 2705 1378
rect 3065 1378 3092 1402
rect 3159 1380 3191 1402
rect 3159 1378 3161 1380
rect 3189 1378 3191 1380
rect 3258 1378 3285 1402
rect 3065 1364 3159 1378
rect 3191 1364 3285 1378
rect 3645 1378 3672 1402
rect 3739 1380 3771 1402
rect 3739 1378 3741 1380
rect 3769 1378 3771 1380
rect 3838 1378 3865 1402
rect 3645 1364 3739 1378
rect 3771 1364 3865 1378
rect 4225 1378 4252 1402
rect 4319 1380 4351 1402
rect 4319 1378 4321 1380
rect 4349 1378 4351 1380
rect 4418 1378 4445 1402
rect 4225 1364 4319 1378
rect 4351 1364 4445 1378
rect 4805 1378 4832 1402
rect 4899 1380 4931 1402
rect 4899 1378 4901 1380
rect 4929 1378 4931 1380
rect 4998 1378 5025 1402
rect 4805 1364 4899 1378
rect 4931 1364 5025 1378
rect 5385 1378 5412 1402
rect 5479 1380 5511 1402
rect 5479 1378 5481 1380
rect 5509 1378 5511 1380
rect 5578 1378 5605 1402
rect 5385 1364 5479 1378
rect 5511 1364 5605 1378
rect 5965 1378 5992 1402
rect 6059 1380 6091 1402
rect 6059 1378 6061 1380
rect 6089 1378 6091 1380
rect 6158 1378 6185 1402
rect 5965 1364 6059 1378
rect 6091 1364 6185 1378
rect 6545 1378 6572 1402
rect 6639 1380 6671 1402
rect 6639 1378 6641 1380
rect 6669 1378 6671 1380
rect 6738 1378 6765 1402
rect 6545 1364 6639 1378
rect 6671 1364 6765 1378
rect 88 1278 106 1306
rect 136 1278 154 1306
rect 396 1278 414 1306
rect 444 1278 463 1306
rect 668 1278 686 1306
rect 716 1278 734 1306
rect 976 1278 994 1306
rect 1024 1278 1043 1306
rect 1248 1278 1266 1306
rect 1296 1278 1314 1306
rect 1556 1278 1574 1306
rect 1604 1278 1623 1306
rect 1828 1278 1846 1306
rect 1876 1278 1894 1306
rect 2136 1278 2154 1306
rect 2184 1278 2203 1306
rect 2408 1278 2426 1306
rect 2456 1278 2474 1306
rect 2716 1278 2734 1306
rect 2764 1278 2783 1306
rect 2988 1278 3006 1306
rect 3036 1278 3054 1306
rect 3296 1278 3314 1306
rect 3344 1278 3363 1306
rect 3568 1278 3586 1306
rect 3616 1278 3634 1306
rect 3876 1278 3894 1306
rect 3924 1278 3943 1306
rect 4148 1278 4166 1306
rect 4196 1278 4214 1306
rect 4456 1278 4474 1306
rect 4504 1278 4523 1306
rect 4728 1278 4746 1306
rect 4776 1278 4794 1306
rect 5036 1278 5054 1306
rect 5084 1278 5103 1306
rect 5308 1278 5326 1306
rect 5356 1278 5374 1306
rect 5616 1278 5634 1306
rect 5664 1278 5683 1306
rect 5888 1278 5906 1306
rect 5936 1278 5954 1306
rect 6196 1278 6214 1306
rect 6244 1278 6263 1306
rect 6468 1278 6486 1306
rect 6516 1278 6534 1306
rect 6776 1278 6794 1306
rect 6824 1278 6843 1306
rect 14 1132 42 1174
rect 72 1160 97 1174
rect 196 1164 221 1174
rect 72 1132 128 1160
rect 158 1132 192 1160
tri 206 1157 213 1164 ne
rect 213 1132 221 1164
rect 251 1132 299 1174
rect 329 1164 354 1174
rect 329 1132 337 1164
rect 453 1160 478 1174
rect 358 1132 392 1160
rect 422 1132 478 1160
rect 508 1132 536 1174
rect 594 1132 622 1174
rect 652 1160 677 1174
rect 776 1164 801 1174
rect 652 1132 708 1160
rect 738 1132 772 1160
tri 786 1157 793 1164 ne
rect 793 1132 801 1164
rect 831 1132 879 1174
rect 909 1164 934 1174
rect 909 1132 917 1164
rect 1033 1160 1058 1174
rect 938 1132 972 1160
rect 1002 1132 1058 1160
rect 1088 1132 1116 1174
rect 1174 1132 1202 1174
rect 1232 1160 1257 1174
rect 1356 1164 1381 1174
rect 1232 1132 1288 1160
rect 1318 1132 1352 1160
tri 1366 1157 1373 1164 ne
rect 1373 1132 1381 1164
rect 1411 1132 1459 1174
rect 1489 1164 1514 1174
rect 1489 1132 1497 1164
rect 1613 1160 1638 1174
rect 1518 1132 1552 1160
rect 1582 1132 1638 1160
rect 1668 1132 1696 1174
rect 1754 1132 1782 1174
rect 1812 1160 1837 1174
rect 1936 1164 1961 1174
rect 1812 1132 1868 1160
rect 1898 1132 1932 1160
tri 1946 1157 1953 1164 ne
rect 1953 1132 1961 1164
rect 1991 1132 2039 1174
rect 2069 1164 2094 1174
rect 2069 1132 2077 1164
rect 2193 1160 2218 1174
rect 2098 1132 2132 1160
rect 2162 1132 2218 1160
rect 2248 1132 2276 1174
rect 2334 1132 2362 1174
rect 2392 1160 2417 1174
rect 2516 1164 2541 1174
rect 2392 1132 2448 1160
rect 2478 1132 2512 1160
tri 2526 1157 2533 1164 ne
rect 2533 1132 2541 1164
rect 2571 1132 2619 1174
rect 2649 1164 2674 1174
rect 2649 1132 2657 1164
rect 2773 1160 2798 1174
rect 2678 1132 2712 1160
rect 2742 1132 2798 1160
rect 2828 1132 2856 1174
rect 2914 1132 2942 1174
rect 2972 1160 2997 1174
rect 3096 1164 3121 1174
rect 2972 1132 3028 1160
rect 3058 1132 3092 1160
tri 3106 1157 3113 1164 ne
rect 3113 1132 3121 1164
rect 3151 1132 3199 1174
rect 3229 1164 3254 1174
rect 3229 1132 3237 1164
rect 3353 1160 3378 1174
rect 3258 1132 3292 1160
rect 3322 1132 3378 1160
rect 3408 1132 3436 1174
rect 3494 1132 3522 1174
rect 3552 1160 3577 1174
rect 3676 1164 3701 1174
rect 3552 1132 3608 1160
rect 3638 1132 3672 1160
tri 3686 1157 3693 1164 ne
rect 3693 1132 3701 1164
rect 3731 1132 3779 1174
rect 3809 1164 3834 1174
rect 3809 1132 3817 1164
rect 3933 1160 3958 1174
rect 3838 1132 3872 1160
rect 3902 1132 3958 1160
rect 3988 1132 4016 1174
rect 4074 1132 4102 1174
rect 4132 1160 4157 1174
rect 4256 1164 4281 1174
rect 4132 1132 4188 1160
rect 4218 1132 4252 1160
tri 4266 1157 4273 1164 ne
rect 4273 1132 4281 1164
rect 4311 1132 4359 1174
rect 4389 1164 4414 1174
rect 4389 1132 4397 1164
rect 4513 1160 4538 1174
rect 4418 1132 4452 1160
rect 4482 1132 4538 1160
rect 4568 1132 4596 1174
rect 4654 1132 4682 1174
rect 4712 1160 4737 1174
rect 4836 1164 4861 1174
rect 4712 1132 4768 1160
rect 4798 1132 4832 1160
tri 4846 1157 4853 1164 ne
rect 4853 1132 4861 1164
rect 4891 1132 4939 1174
rect 4969 1164 4994 1174
rect 4969 1132 4977 1164
rect 5093 1160 5118 1174
rect 4998 1132 5032 1160
rect 5062 1132 5118 1160
rect 5148 1132 5176 1174
rect 5234 1132 5262 1174
rect 5292 1160 5317 1174
rect 5416 1164 5441 1174
rect 5292 1132 5348 1160
rect 5378 1132 5412 1160
tri 5426 1157 5433 1164 ne
rect 5433 1132 5441 1164
rect 5471 1132 5519 1174
rect 5549 1164 5574 1174
rect 5549 1132 5557 1164
rect 5673 1160 5698 1174
rect 5578 1132 5612 1160
rect 5642 1132 5698 1160
rect 5728 1132 5756 1174
rect 5814 1132 5842 1174
rect 5872 1160 5897 1174
rect 5996 1164 6021 1174
rect 5872 1132 5928 1160
rect 5958 1132 5992 1160
tri 6006 1157 6013 1164 ne
rect 6013 1132 6021 1164
rect 6051 1132 6099 1174
rect 6129 1164 6154 1174
rect 6129 1132 6137 1164
rect 6253 1160 6278 1174
rect 6158 1132 6192 1160
rect 6222 1132 6278 1160
rect 6308 1132 6336 1174
rect 6394 1132 6422 1174
rect 6452 1160 6477 1174
rect 6576 1164 6601 1174
rect 6452 1132 6508 1160
rect 6538 1132 6572 1160
tri 6586 1157 6593 1164 ne
rect 6593 1132 6601 1164
rect 6631 1132 6679 1174
rect 6709 1164 6734 1174
rect 6709 1132 6717 1164
rect 6833 1160 6858 1174
rect 6738 1132 6772 1160
rect 6802 1132 6858 1160
rect 6888 1132 6916 1174
rect 165 1108 192 1132
rect 259 1110 291 1132
rect 259 1108 261 1110
rect 289 1108 291 1110
rect 358 1108 385 1132
rect 165 1094 259 1108
rect 291 1094 385 1108
rect 745 1108 772 1132
rect 839 1110 871 1132
rect 839 1108 841 1110
rect 869 1108 871 1110
rect 938 1108 965 1132
rect 745 1094 839 1108
rect 871 1094 965 1108
rect 1325 1108 1352 1132
rect 1419 1110 1451 1132
rect 1419 1108 1421 1110
rect 1449 1108 1451 1110
rect 1518 1108 1545 1132
rect 1325 1094 1419 1108
rect 1451 1094 1545 1108
rect 1905 1108 1932 1132
rect 1999 1110 2031 1132
rect 1999 1108 2001 1110
rect 2029 1108 2031 1110
rect 2098 1108 2125 1132
rect 1905 1094 1999 1108
rect 2031 1094 2125 1108
rect 2485 1108 2512 1132
rect 2579 1110 2611 1132
rect 2579 1108 2581 1110
rect 2609 1108 2611 1110
rect 2678 1108 2705 1132
rect 2485 1094 2579 1108
rect 2611 1094 2705 1108
rect 3065 1108 3092 1132
rect 3159 1110 3191 1132
rect 3159 1108 3161 1110
rect 3189 1108 3191 1110
rect 3258 1108 3285 1132
rect 3065 1094 3159 1108
rect 3191 1094 3285 1108
rect 3645 1108 3672 1132
rect 3739 1110 3771 1132
rect 3739 1108 3741 1110
rect 3769 1108 3771 1110
rect 3838 1108 3865 1132
rect 3645 1094 3739 1108
rect 3771 1094 3865 1108
rect 4225 1108 4252 1132
rect 4319 1110 4351 1132
rect 4319 1108 4321 1110
rect 4349 1108 4351 1110
rect 4418 1108 4445 1132
rect 4225 1094 4319 1108
rect 4351 1094 4445 1108
rect 4805 1108 4832 1132
rect 4899 1110 4931 1132
rect 4899 1108 4901 1110
rect 4929 1108 4931 1110
rect 4998 1108 5025 1132
rect 4805 1094 4899 1108
rect 4931 1094 5025 1108
rect 5385 1108 5412 1132
rect 5479 1110 5511 1132
rect 5479 1108 5481 1110
rect 5509 1108 5511 1110
rect 5578 1108 5605 1132
rect 5385 1094 5479 1108
rect 5511 1094 5605 1108
rect 5965 1108 5992 1132
rect 6059 1110 6091 1132
rect 6059 1108 6061 1110
rect 6089 1108 6091 1110
rect 6158 1108 6185 1132
rect 5965 1094 6059 1108
rect 6091 1094 6185 1108
rect 6545 1108 6572 1132
rect 6639 1110 6671 1132
rect 6639 1108 6641 1110
rect 6669 1108 6671 1110
rect 6738 1108 6765 1132
rect 6545 1094 6639 1108
rect 6671 1094 6765 1108
rect 88 1008 106 1036
rect 136 1008 154 1036
rect 396 1008 414 1036
rect 444 1008 463 1036
rect 668 1008 686 1036
rect 716 1008 734 1036
rect 976 1008 994 1036
rect 1024 1008 1043 1036
rect 1248 1008 1266 1036
rect 1296 1008 1314 1036
rect 1556 1008 1574 1036
rect 1604 1008 1623 1036
rect 1828 1008 1846 1036
rect 1876 1008 1894 1036
rect 2136 1008 2154 1036
rect 2184 1008 2203 1036
rect 2408 1008 2426 1036
rect 2456 1008 2474 1036
rect 2716 1008 2734 1036
rect 2764 1008 2783 1036
rect 2988 1008 3006 1036
rect 3036 1008 3054 1036
rect 3296 1008 3314 1036
rect 3344 1008 3363 1036
rect 3568 1008 3586 1036
rect 3616 1008 3634 1036
rect 3876 1008 3894 1036
rect 3924 1008 3943 1036
rect 4148 1008 4166 1036
rect 4196 1008 4214 1036
rect 4456 1008 4474 1036
rect 4504 1008 4523 1036
rect 4728 1008 4746 1036
rect 4776 1008 4794 1036
rect 5036 1008 5054 1036
rect 5084 1008 5103 1036
rect 5308 1008 5326 1036
rect 5356 1008 5374 1036
rect 5616 1008 5634 1036
rect 5664 1008 5683 1036
rect 5888 1008 5906 1036
rect 5936 1008 5954 1036
rect 6196 1008 6214 1036
rect 6244 1008 6263 1036
rect 6468 1008 6486 1036
rect 6516 1008 6534 1036
rect 6776 1008 6794 1036
rect 6824 1008 6843 1036
rect 14 862 42 904
rect 72 890 97 904
rect 196 894 221 904
rect 72 862 128 890
rect 158 862 192 890
tri 206 887 213 894 ne
rect 213 862 221 894
rect 251 862 299 904
rect 329 894 354 904
rect 329 862 337 894
rect 453 890 478 904
rect 358 862 392 890
rect 422 862 478 890
rect 508 862 536 904
rect 594 862 622 904
rect 652 890 677 904
rect 776 894 801 904
rect 652 862 708 890
rect 738 862 772 890
tri 786 887 793 894 ne
rect 793 862 801 894
rect 831 862 879 904
rect 909 894 934 904
rect 909 862 917 894
rect 1033 890 1058 904
rect 938 862 972 890
rect 1002 862 1058 890
rect 1088 862 1116 904
rect 1174 862 1202 904
rect 1232 890 1257 904
rect 1356 894 1381 904
rect 1232 862 1288 890
rect 1318 862 1352 890
tri 1366 887 1373 894 ne
rect 1373 862 1381 894
rect 1411 862 1459 904
rect 1489 894 1514 904
rect 1489 862 1497 894
rect 1613 890 1638 904
rect 1518 862 1552 890
rect 1582 862 1638 890
rect 1668 862 1696 904
rect 1754 862 1782 904
rect 1812 890 1837 904
rect 1936 894 1961 904
rect 1812 862 1868 890
rect 1898 862 1932 890
tri 1946 887 1953 894 ne
rect 1953 862 1961 894
rect 1991 862 2039 904
rect 2069 894 2094 904
rect 2069 862 2077 894
rect 2193 890 2218 904
rect 2098 862 2132 890
rect 2162 862 2218 890
rect 2248 862 2276 904
rect 2334 862 2362 904
rect 2392 890 2417 904
rect 2516 894 2541 904
rect 2392 862 2448 890
rect 2478 862 2512 890
tri 2526 887 2533 894 ne
rect 2533 862 2541 894
rect 2571 862 2619 904
rect 2649 894 2674 904
rect 2649 862 2657 894
rect 2773 890 2798 904
rect 2678 862 2712 890
rect 2742 862 2798 890
rect 2828 862 2856 904
rect 2914 862 2942 904
rect 2972 890 2997 904
rect 3096 894 3121 904
rect 2972 862 3028 890
rect 3058 862 3092 890
tri 3106 887 3113 894 ne
rect 3113 862 3121 894
rect 3151 862 3199 904
rect 3229 894 3254 904
rect 3229 862 3237 894
rect 3353 890 3378 904
rect 3258 862 3292 890
rect 3322 862 3378 890
rect 3408 862 3436 904
rect 3494 862 3522 904
rect 3552 890 3577 904
rect 3676 894 3701 904
rect 3552 862 3608 890
rect 3638 862 3672 890
tri 3686 887 3693 894 ne
rect 3693 862 3701 894
rect 3731 862 3779 904
rect 3809 894 3834 904
rect 3809 862 3817 894
rect 3933 890 3958 904
rect 3838 862 3872 890
rect 3902 862 3958 890
rect 3988 862 4016 904
rect 4074 862 4102 904
rect 4132 890 4157 904
rect 4256 894 4281 904
rect 4132 862 4188 890
rect 4218 862 4252 890
tri 4266 887 4273 894 ne
rect 4273 862 4281 894
rect 4311 862 4359 904
rect 4389 894 4414 904
rect 4389 862 4397 894
rect 4513 890 4538 904
rect 4418 862 4452 890
rect 4482 862 4538 890
rect 4568 862 4596 904
rect 4654 862 4682 904
rect 4712 890 4737 904
rect 4836 894 4861 904
rect 4712 862 4768 890
rect 4798 862 4832 890
tri 4846 887 4853 894 ne
rect 4853 862 4861 894
rect 4891 862 4939 904
rect 4969 894 4994 904
rect 4969 862 4977 894
rect 5093 890 5118 904
rect 4998 862 5032 890
rect 5062 862 5118 890
rect 5148 862 5176 904
rect 5234 862 5262 904
rect 5292 890 5317 904
rect 5416 894 5441 904
rect 5292 862 5348 890
rect 5378 862 5412 890
tri 5426 887 5433 894 ne
rect 5433 862 5441 894
rect 5471 862 5519 904
rect 5549 894 5574 904
rect 5549 862 5557 894
rect 5673 890 5698 904
rect 5578 862 5612 890
rect 5642 862 5698 890
rect 5728 862 5756 904
rect 5814 862 5842 904
rect 5872 890 5897 904
rect 5996 894 6021 904
rect 5872 862 5928 890
rect 5958 862 5992 890
tri 6006 887 6013 894 ne
rect 6013 862 6021 894
rect 6051 862 6099 904
rect 6129 894 6154 904
rect 6129 862 6137 894
rect 6253 890 6278 904
rect 6158 862 6192 890
rect 6222 862 6278 890
rect 6308 862 6336 904
rect 6394 862 6422 904
rect 6452 890 6477 904
rect 6576 894 6601 904
rect 6452 862 6508 890
rect 6538 862 6572 890
tri 6586 887 6593 894 ne
rect 6593 862 6601 894
rect 6631 862 6679 904
rect 6709 894 6734 904
rect 6709 862 6717 894
rect 6833 890 6858 904
rect 6738 862 6772 890
rect 6802 862 6858 890
rect 6888 862 6916 904
rect 165 838 192 862
rect 259 840 291 862
rect 259 838 261 840
rect 289 838 291 840
rect 358 838 385 862
rect 165 824 259 838
rect 291 824 385 838
rect 745 838 772 862
rect 839 840 871 862
rect 839 838 841 840
rect 869 838 871 840
rect 938 838 965 862
rect 745 824 839 838
rect 871 824 965 838
rect 1325 838 1352 862
rect 1419 840 1451 862
rect 1419 838 1421 840
rect 1449 838 1451 840
rect 1518 838 1545 862
rect 1325 824 1419 838
rect 1451 824 1545 838
rect 1905 838 1932 862
rect 1999 840 2031 862
rect 1999 838 2001 840
rect 2029 838 2031 840
rect 2098 838 2125 862
rect 1905 824 1999 838
rect 2031 824 2125 838
rect 2485 838 2512 862
rect 2579 840 2611 862
rect 2579 838 2581 840
rect 2609 838 2611 840
rect 2678 838 2705 862
rect 2485 824 2579 838
rect 2611 824 2705 838
rect 3065 838 3092 862
rect 3159 840 3191 862
rect 3159 838 3161 840
rect 3189 838 3191 840
rect 3258 838 3285 862
rect 3065 824 3159 838
rect 3191 824 3285 838
rect 3645 838 3672 862
rect 3739 840 3771 862
rect 3739 838 3741 840
rect 3769 838 3771 840
rect 3838 838 3865 862
rect 3645 824 3739 838
rect 3771 824 3865 838
rect 4225 838 4252 862
rect 4319 840 4351 862
rect 4319 838 4321 840
rect 4349 838 4351 840
rect 4418 838 4445 862
rect 4225 824 4319 838
rect 4351 824 4445 838
rect 4805 838 4832 862
rect 4899 840 4931 862
rect 4899 838 4901 840
rect 4929 838 4931 840
rect 4998 838 5025 862
rect 4805 824 4899 838
rect 4931 824 5025 838
rect 5385 838 5412 862
rect 5479 840 5511 862
rect 5479 838 5481 840
rect 5509 838 5511 840
rect 5578 838 5605 862
rect 5385 824 5479 838
rect 5511 824 5605 838
rect 5965 838 5992 862
rect 6059 840 6091 862
rect 6059 838 6061 840
rect 6089 838 6091 840
rect 6158 838 6185 862
rect 5965 824 6059 838
rect 6091 824 6185 838
rect 6545 838 6572 862
rect 6639 840 6671 862
rect 6639 838 6641 840
rect 6669 838 6671 840
rect 6738 838 6765 862
rect 6545 824 6639 838
rect 6671 824 6765 838
rect 88 738 106 766
rect 136 738 154 766
rect 396 738 414 766
rect 444 738 463 766
rect 668 738 686 766
rect 716 738 734 766
rect 976 738 994 766
rect 1024 738 1043 766
rect 1248 738 1266 766
rect 1296 738 1314 766
rect 1556 738 1574 766
rect 1604 738 1623 766
rect 1828 738 1846 766
rect 1876 738 1894 766
rect 2136 738 2154 766
rect 2184 738 2203 766
rect 2408 738 2426 766
rect 2456 738 2474 766
rect 2716 738 2734 766
rect 2764 738 2783 766
rect 2988 738 3006 766
rect 3036 738 3054 766
rect 3296 738 3314 766
rect 3344 738 3363 766
rect 3568 738 3586 766
rect 3616 738 3634 766
rect 3876 738 3894 766
rect 3924 738 3943 766
rect 4148 738 4166 766
rect 4196 738 4214 766
rect 4456 738 4474 766
rect 4504 738 4523 766
rect 4728 738 4746 766
rect 4776 738 4794 766
rect 5036 738 5054 766
rect 5084 738 5103 766
rect 5308 738 5326 766
rect 5356 738 5374 766
rect 5616 738 5634 766
rect 5664 738 5683 766
rect 5888 738 5906 766
rect 5936 738 5954 766
rect 6196 738 6214 766
rect 6244 738 6263 766
rect 6468 738 6486 766
rect 6516 738 6534 766
rect 6776 738 6794 766
rect 6824 738 6843 766
rect 14 592 42 634
rect 72 620 97 634
rect 196 624 221 634
rect 72 592 128 620
rect 158 592 192 620
tri 206 617 213 624 ne
rect 213 592 221 624
rect 251 592 299 634
rect 329 624 354 634
rect 329 592 337 624
rect 453 620 478 634
rect 358 592 392 620
rect 422 592 478 620
rect 508 592 536 634
rect 594 592 622 634
rect 652 620 677 634
rect 776 624 801 634
rect 652 592 708 620
rect 738 592 772 620
tri 786 617 793 624 ne
rect 793 592 801 624
rect 831 592 879 634
rect 909 624 934 634
rect 909 592 917 624
rect 1033 620 1058 634
rect 938 592 972 620
rect 1002 592 1058 620
rect 1088 592 1116 634
rect 1174 592 1202 634
rect 1232 620 1257 634
rect 1356 624 1381 634
rect 1232 592 1288 620
rect 1318 592 1352 620
tri 1366 617 1373 624 ne
rect 1373 592 1381 624
rect 1411 592 1459 634
rect 1489 624 1514 634
rect 1489 592 1497 624
rect 1613 620 1638 634
rect 1518 592 1552 620
rect 1582 592 1638 620
rect 1668 592 1696 634
rect 1754 592 1782 634
rect 1812 620 1837 634
rect 1936 624 1961 634
rect 1812 592 1868 620
rect 1898 592 1932 620
tri 1946 617 1953 624 ne
rect 1953 592 1961 624
rect 1991 592 2039 634
rect 2069 624 2094 634
rect 2069 592 2077 624
rect 2193 620 2218 634
rect 2098 592 2132 620
rect 2162 592 2218 620
rect 2248 592 2276 634
rect 2334 592 2362 634
rect 2392 620 2417 634
rect 2516 624 2541 634
rect 2392 592 2448 620
rect 2478 592 2512 620
tri 2526 617 2533 624 ne
rect 2533 592 2541 624
rect 2571 592 2619 634
rect 2649 624 2674 634
rect 2649 592 2657 624
rect 2773 620 2798 634
rect 2678 592 2712 620
rect 2742 592 2798 620
rect 2828 592 2856 634
rect 2914 592 2942 634
rect 2972 620 2997 634
rect 3096 624 3121 634
rect 2972 592 3028 620
rect 3058 592 3092 620
tri 3106 617 3113 624 ne
rect 3113 592 3121 624
rect 3151 592 3199 634
rect 3229 624 3254 634
rect 3229 592 3237 624
rect 3353 620 3378 634
rect 3258 592 3292 620
rect 3322 592 3378 620
rect 3408 592 3436 634
rect 3494 592 3522 634
rect 3552 620 3577 634
rect 3676 624 3701 634
rect 3552 592 3608 620
rect 3638 592 3672 620
tri 3686 617 3693 624 ne
rect 3693 592 3701 624
rect 3731 592 3779 634
rect 3809 624 3834 634
rect 3809 592 3817 624
rect 3933 620 3958 634
rect 3838 592 3872 620
rect 3902 592 3958 620
rect 3988 592 4016 634
rect 4074 592 4102 634
rect 4132 620 4157 634
rect 4256 624 4281 634
rect 4132 592 4188 620
rect 4218 592 4252 620
tri 4266 617 4273 624 ne
rect 4273 592 4281 624
rect 4311 592 4359 634
rect 4389 624 4414 634
rect 4389 592 4397 624
rect 4513 620 4538 634
rect 4418 592 4452 620
rect 4482 592 4538 620
rect 4568 592 4596 634
rect 4654 592 4682 634
rect 4712 620 4737 634
rect 4836 624 4861 634
rect 4712 592 4768 620
rect 4798 592 4832 620
tri 4846 617 4853 624 ne
rect 4853 592 4861 624
rect 4891 592 4939 634
rect 4969 624 4994 634
rect 4969 592 4977 624
rect 5093 620 5118 634
rect 4998 592 5032 620
rect 5062 592 5118 620
rect 5148 592 5176 634
rect 5234 592 5262 634
rect 5292 620 5317 634
rect 5416 624 5441 634
rect 5292 592 5348 620
rect 5378 592 5412 620
tri 5426 617 5433 624 ne
rect 5433 592 5441 624
rect 5471 592 5519 634
rect 5549 624 5574 634
rect 5549 592 5557 624
rect 5673 620 5698 634
rect 5578 592 5612 620
rect 5642 592 5698 620
rect 5728 592 5756 634
rect 5814 592 5842 634
rect 5872 620 5897 634
rect 5996 624 6021 634
rect 5872 592 5928 620
rect 5958 592 5992 620
tri 6006 617 6013 624 ne
rect 6013 592 6021 624
rect 6051 592 6099 634
rect 6129 624 6154 634
rect 6129 592 6137 624
rect 6253 620 6278 634
rect 6158 592 6192 620
rect 6222 592 6278 620
rect 6308 592 6336 634
rect 6394 592 6422 634
rect 6452 620 6477 634
rect 6576 624 6601 634
rect 6452 592 6508 620
rect 6538 592 6572 620
tri 6586 617 6593 624 ne
rect 6593 592 6601 624
rect 6631 592 6679 634
rect 6709 624 6734 634
rect 6709 592 6717 624
rect 6833 620 6858 634
rect 6738 592 6772 620
rect 6802 592 6858 620
rect 6888 592 6916 634
rect 165 568 192 592
rect 259 570 291 592
rect 259 568 261 570
rect 289 568 291 570
rect 358 568 385 592
rect 165 554 259 568
rect 291 554 385 568
rect 745 568 772 592
rect 839 570 871 592
rect 839 568 841 570
rect 869 568 871 570
rect 938 568 965 592
rect 745 554 839 568
rect 871 554 965 568
rect 1325 568 1352 592
rect 1419 570 1451 592
rect 1419 568 1421 570
rect 1449 568 1451 570
rect 1518 568 1545 592
rect 1325 554 1419 568
rect 1451 554 1545 568
rect 1905 568 1932 592
rect 1999 570 2031 592
rect 1999 568 2001 570
rect 2029 568 2031 570
rect 2098 568 2125 592
rect 1905 554 1999 568
rect 2031 554 2125 568
rect 2485 568 2512 592
rect 2579 570 2611 592
rect 2579 568 2581 570
rect 2609 568 2611 570
rect 2678 568 2705 592
rect 2485 554 2579 568
rect 2611 554 2705 568
rect 3065 568 3092 592
rect 3159 570 3191 592
rect 3159 568 3161 570
rect 3189 568 3191 570
rect 3258 568 3285 592
rect 3065 554 3159 568
rect 3191 554 3285 568
rect 3645 568 3672 592
rect 3739 570 3771 592
rect 3739 568 3741 570
rect 3769 568 3771 570
rect 3838 568 3865 592
rect 3645 554 3739 568
rect 3771 554 3865 568
rect 4225 568 4252 592
rect 4319 570 4351 592
rect 4319 568 4321 570
rect 4349 568 4351 570
rect 4418 568 4445 592
rect 4225 554 4319 568
rect 4351 554 4445 568
rect 4805 568 4832 592
rect 4899 570 4931 592
rect 4899 568 4901 570
rect 4929 568 4931 570
rect 4998 568 5025 592
rect 4805 554 4899 568
rect 4931 554 5025 568
rect 5385 568 5412 592
rect 5479 570 5511 592
rect 5479 568 5481 570
rect 5509 568 5511 570
rect 5578 568 5605 592
rect 5385 554 5479 568
rect 5511 554 5605 568
rect 5965 568 5992 592
rect 6059 570 6091 592
rect 6059 568 6061 570
rect 6089 568 6091 570
rect 6158 568 6185 592
rect 5965 554 6059 568
rect 6091 554 6185 568
rect 6545 568 6572 592
rect 6639 570 6671 592
rect 6639 568 6641 570
rect 6669 568 6671 570
rect 6738 568 6765 592
rect 6545 554 6639 568
rect 6671 554 6765 568
rect 88 468 106 496
rect 136 468 154 496
rect 396 468 414 496
rect 444 468 463 496
rect 668 468 686 496
rect 716 468 734 496
rect 976 468 994 496
rect 1024 468 1043 496
rect 1248 468 1266 496
rect 1296 468 1314 496
rect 1556 468 1574 496
rect 1604 468 1623 496
rect 1828 468 1846 496
rect 1876 468 1894 496
rect 2136 468 2154 496
rect 2184 468 2203 496
rect 2408 468 2426 496
rect 2456 468 2474 496
rect 2716 468 2734 496
rect 2764 468 2783 496
rect 2988 468 3006 496
rect 3036 468 3054 496
rect 3296 468 3314 496
rect 3344 468 3363 496
rect 3568 468 3586 496
rect 3616 468 3634 496
rect 3876 468 3894 496
rect 3924 468 3943 496
rect 4148 468 4166 496
rect 4196 468 4214 496
rect 4456 468 4474 496
rect 4504 468 4523 496
rect 4728 468 4746 496
rect 4776 468 4794 496
rect 5036 468 5054 496
rect 5084 468 5103 496
rect 5308 468 5326 496
rect 5356 468 5374 496
rect 5616 468 5634 496
rect 5664 468 5683 496
rect 5888 468 5906 496
rect 5936 468 5954 496
rect 6196 468 6214 496
rect 6244 468 6263 496
rect 6468 468 6486 496
rect 6516 468 6534 496
rect 6776 468 6794 496
rect 6824 468 6843 496
rect 14 322 42 364
rect 72 350 97 364
rect 196 354 221 364
rect 72 322 128 350
rect 158 322 192 350
tri 206 347 213 354 ne
rect 213 322 221 354
rect 251 322 299 364
rect 329 354 354 364
rect 329 322 337 354
rect 453 350 478 364
rect 358 322 392 350
rect 422 322 478 350
rect 508 322 536 364
rect 594 322 622 364
rect 652 350 677 364
rect 776 354 801 364
rect 652 322 708 350
rect 738 322 772 350
tri 786 347 793 354 ne
rect 793 322 801 354
rect 831 322 879 364
rect 909 354 934 364
rect 909 322 917 354
rect 1033 350 1058 364
rect 938 322 972 350
rect 1002 322 1058 350
rect 1088 322 1116 364
rect 1174 322 1202 364
rect 1232 350 1257 364
rect 1356 354 1381 364
rect 1232 322 1288 350
rect 1318 322 1352 350
tri 1366 347 1373 354 ne
rect 1373 322 1381 354
rect 1411 322 1459 364
rect 1489 354 1514 364
rect 1489 322 1497 354
rect 1613 350 1638 364
rect 1518 322 1552 350
rect 1582 322 1638 350
rect 1668 322 1696 364
rect 1754 322 1782 364
rect 1812 350 1837 364
rect 1936 354 1961 364
rect 1812 322 1868 350
rect 1898 322 1932 350
tri 1946 347 1953 354 ne
rect 1953 322 1961 354
rect 1991 322 2039 364
rect 2069 354 2094 364
rect 2069 322 2077 354
rect 2193 350 2218 364
rect 2098 322 2132 350
rect 2162 322 2218 350
rect 2248 322 2276 364
rect 2334 322 2362 364
rect 2392 350 2417 364
rect 2516 354 2541 364
rect 2392 322 2448 350
rect 2478 322 2512 350
tri 2526 347 2533 354 ne
rect 2533 322 2541 354
rect 2571 322 2619 364
rect 2649 354 2674 364
rect 2649 322 2657 354
rect 2773 350 2798 364
rect 2678 322 2712 350
rect 2742 322 2798 350
rect 2828 322 2856 364
rect 2914 322 2942 364
rect 2972 350 2997 364
rect 3096 354 3121 364
rect 2972 322 3028 350
rect 3058 322 3092 350
tri 3106 347 3113 354 ne
rect 3113 322 3121 354
rect 3151 322 3199 364
rect 3229 354 3254 364
rect 3229 322 3237 354
rect 3353 350 3378 364
rect 3258 322 3292 350
rect 3322 322 3378 350
rect 3408 322 3436 364
rect 3494 322 3522 364
rect 3552 350 3577 364
rect 3676 354 3701 364
rect 3552 322 3608 350
rect 3638 322 3672 350
tri 3686 347 3693 354 ne
rect 3693 322 3701 354
rect 3731 322 3779 364
rect 3809 354 3834 364
rect 3809 322 3817 354
rect 3933 350 3958 364
rect 3838 322 3872 350
rect 3902 322 3958 350
rect 3988 322 4016 364
rect 4074 322 4102 364
rect 4132 350 4157 364
rect 4256 354 4281 364
rect 4132 322 4188 350
rect 4218 322 4252 350
tri 4266 347 4273 354 ne
rect 4273 322 4281 354
rect 4311 322 4359 364
rect 4389 354 4414 364
rect 4389 322 4397 354
rect 4513 350 4538 364
rect 4418 322 4452 350
rect 4482 322 4538 350
rect 4568 322 4596 364
rect 4654 322 4682 364
rect 4712 350 4737 364
rect 4836 354 4861 364
rect 4712 322 4768 350
rect 4798 322 4832 350
tri 4846 347 4853 354 ne
rect 4853 322 4861 354
rect 4891 322 4939 364
rect 4969 354 4994 364
rect 4969 322 4977 354
rect 5093 350 5118 364
rect 4998 322 5032 350
rect 5062 322 5118 350
rect 5148 322 5176 364
rect 5234 322 5262 364
rect 5292 350 5317 364
rect 5416 354 5441 364
rect 5292 322 5348 350
rect 5378 322 5412 350
tri 5426 347 5433 354 ne
rect 5433 322 5441 354
rect 5471 322 5519 364
rect 5549 354 5574 364
rect 5549 322 5557 354
rect 5673 350 5698 364
rect 5578 322 5612 350
rect 5642 322 5698 350
rect 5728 322 5756 364
rect 5814 322 5842 364
rect 5872 350 5897 364
rect 5996 354 6021 364
rect 5872 322 5928 350
rect 5958 322 5992 350
tri 6006 347 6013 354 ne
rect 6013 322 6021 354
rect 6051 322 6099 364
rect 6129 354 6154 364
rect 6129 322 6137 354
rect 6253 350 6278 364
rect 6158 322 6192 350
rect 6222 322 6278 350
rect 6308 322 6336 364
rect 6394 322 6422 364
rect 6452 350 6477 364
rect 6576 354 6601 364
rect 6452 322 6508 350
rect 6538 322 6572 350
tri 6586 347 6593 354 ne
rect 6593 322 6601 354
rect 6631 322 6679 364
rect 6709 354 6734 364
rect 6709 322 6717 354
rect 6833 350 6858 364
rect 6738 322 6772 350
rect 6802 322 6858 350
rect 6888 322 6916 364
rect 165 298 192 322
rect 259 300 291 322
rect 259 298 261 300
rect 289 298 291 300
rect 358 298 385 322
rect 165 284 259 298
rect 291 284 385 298
rect 745 298 772 322
rect 839 300 871 322
rect 839 298 841 300
rect 869 298 871 300
rect 938 298 965 322
rect 745 284 839 298
rect 871 284 965 298
rect 1325 298 1352 322
rect 1419 300 1451 322
rect 1419 298 1421 300
rect 1449 298 1451 300
rect 1518 298 1545 322
rect 1325 284 1419 298
rect 1451 284 1545 298
rect 1905 298 1932 322
rect 1999 300 2031 322
rect 1999 298 2001 300
rect 2029 298 2031 300
rect 2098 298 2125 322
rect 1905 284 1999 298
rect 2031 284 2125 298
rect 2485 298 2512 322
rect 2579 300 2611 322
rect 2579 298 2581 300
rect 2609 298 2611 300
rect 2678 298 2705 322
rect 2485 284 2579 298
rect 2611 284 2705 298
rect 3065 298 3092 322
rect 3159 300 3191 322
rect 3159 298 3161 300
rect 3189 298 3191 300
rect 3258 298 3285 322
rect 3065 284 3159 298
rect 3191 284 3285 298
rect 3645 298 3672 322
rect 3739 300 3771 322
rect 3739 298 3741 300
rect 3769 298 3771 300
rect 3838 298 3865 322
rect 3645 284 3739 298
rect 3771 284 3865 298
rect 4225 298 4252 322
rect 4319 300 4351 322
rect 4319 298 4321 300
rect 4349 298 4351 300
rect 4418 298 4445 322
rect 4225 284 4319 298
rect 4351 284 4445 298
rect 4805 298 4832 322
rect 4899 300 4931 322
rect 4899 298 4901 300
rect 4929 298 4931 300
rect 4998 298 5025 322
rect 4805 284 4899 298
rect 4931 284 5025 298
rect 5385 298 5412 322
rect 5479 300 5511 322
rect 5479 298 5481 300
rect 5509 298 5511 300
rect 5578 298 5605 322
rect 5385 284 5479 298
rect 5511 284 5605 298
rect 5965 298 5992 322
rect 6059 300 6091 322
rect 6059 298 6061 300
rect 6089 298 6091 300
rect 6158 298 6185 322
rect 5965 284 6059 298
rect 6091 284 6185 298
rect 6545 298 6572 322
rect 6639 300 6671 322
rect 6639 298 6641 300
rect 6669 298 6671 300
rect 6738 298 6765 322
rect 6545 284 6639 298
rect 6671 284 6765 298
rect 88 198 106 226
rect 136 198 154 226
rect 396 198 414 226
rect 444 198 463 226
rect 668 198 686 226
rect 716 198 734 226
rect 976 198 994 226
rect 1024 198 1043 226
rect 1248 198 1266 226
rect 1296 198 1314 226
rect 1556 198 1574 226
rect 1604 198 1623 226
rect 1828 198 1846 226
rect 1876 198 1894 226
rect 2136 198 2154 226
rect 2184 198 2203 226
rect 2408 198 2426 226
rect 2456 198 2474 226
rect 2716 198 2734 226
rect 2764 198 2783 226
rect 2988 198 3006 226
rect 3036 198 3054 226
rect 3296 198 3314 226
rect 3344 198 3363 226
rect 3568 198 3586 226
rect 3616 198 3634 226
rect 3876 198 3894 226
rect 3924 198 3943 226
rect 4148 198 4166 226
rect 4196 198 4214 226
rect 4456 198 4474 226
rect 4504 198 4523 226
rect 4728 198 4746 226
rect 4776 198 4794 226
rect 5036 198 5054 226
rect 5084 198 5103 226
rect 5308 198 5326 226
rect 5356 198 5374 226
rect 5616 198 5634 226
rect 5664 198 5683 226
rect 5888 198 5906 226
rect 5936 198 5954 226
rect 6196 198 6214 226
rect 6244 198 6263 226
rect 6468 198 6486 226
rect 6516 198 6534 226
rect 6776 198 6794 226
rect 6824 198 6843 226
rect 14 52 42 94
rect 72 80 97 94
rect 196 84 221 94
rect 72 52 128 80
rect 158 52 192 80
tri 206 77 213 84 ne
rect 213 52 221 84
rect 251 52 299 94
rect 329 84 354 94
rect 329 52 337 84
rect 453 80 478 94
rect 358 52 392 80
rect 422 52 478 80
rect 508 52 536 94
rect 594 52 622 94
rect 652 80 677 94
rect 776 84 801 94
rect 652 52 708 80
rect 738 52 772 80
tri 786 77 793 84 ne
rect 793 52 801 84
rect 831 52 879 94
rect 909 84 934 94
rect 909 52 917 84
rect 1033 80 1058 94
rect 938 52 972 80
rect 1002 52 1058 80
rect 1088 52 1116 94
rect 1174 52 1202 94
rect 1232 80 1257 94
rect 1356 84 1381 94
rect 1232 52 1288 80
rect 1318 52 1352 80
tri 1366 77 1373 84 ne
rect 1373 52 1381 84
rect 1411 52 1459 94
rect 1489 84 1514 94
rect 1489 52 1497 84
rect 1613 80 1638 94
rect 1518 52 1552 80
rect 1582 52 1638 80
rect 1668 52 1696 94
rect 1754 52 1782 94
rect 1812 80 1837 94
rect 1936 84 1961 94
rect 1812 52 1868 80
rect 1898 52 1932 80
tri 1946 77 1953 84 ne
rect 1953 52 1961 84
rect 1991 52 2039 94
rect 2069 84 2094 94
rect 2069 52 2077 84
rect 2193 80 2218 94
rect 2098 52 2132 80
rect 2162 52 2218 80
rect 2248 52 2276 94
rect 2334 52 2362 94
rect 2392 80 2417 94
rect 2516 84 2541 94
rect 2392 52 2448 80
rect 2478 52 2512 80
tri 2526 77 2533 84 ne
rect 2533 52 2541 84
rect 2571 52 2619 94
rect 2649 84 2674 94
rect 2649 52 2657 84
rect 2773 80 2798 94
rect 2678 52 2712 80
rect 2742 52 2798 80
rect 2828 52 2856 94
rect 2914 52 2942 94
rect 2972 80 2997 94
rect 3096 84 3121 94
rect 2972 52 3028 80
rect 3058 52 3092 80
tri 3106 77 3113 84 ne
rect 3113 52 3121 84
rect 3151 52 3199 94
rect 3229 84 3254 94
rect 3229 52 3237 84
rect 3353 80 3378 94
rect 3258 52 3292 80
rect 3322 52 3378 80
rect 3408 52 3436 94
rect 3494 52 3522 94
rect 3552 80 3577 94
rect 3676 84 3701 94
rect 3552 52 3608 80
rect 3638 52 3672 80
tri 3686 77 3693 84 ne
rect 3693 52 3701 84
rect 3731 52 3779 94
rect 3809 84 3834 94
rect 3809 52 3817 84
rect 3933 80 3958 94
rect 3838 52 3872 80
rect 3902 52 3958 80
rect 3988 52 4016 94
rect 4074 52 4102 94
rect 4132 80 4157 94
rect 4256 84 4281 94
rect 4132 52 4188 80
rect 4218 52 4252 80
tri 4266 77 4273 84 ne
rect 4273 52 4281 84
rect 4311 52 4359 94
rect 4389 84 4414 94
rect 4389 52 4397 84
rect 4513 80 4538 94
rect 4418 52 4452 80
rect 4482 52 4538 80
rect 4568 52 4596 94
rect 4654 52 4682 94
rect 4712 80 4737 94
rect 4836 84 4861 94
rect 4712 52 4768 80
rect 4798 52 4832 80
tri 4846 77 4853 84 ne
rect 4853 52 4861 84
rect 4891 52 4939 94
rect 4969 84 4994 94
rect 4969 52 4977 84
rect 5093 80 5118 94
rect 4998 52 5032 80
rect 5062 52 5118 80
rect 5148 52 5176 94
rect 5234 52 5262 94
rect 5292 80 5317 94
rect 5416 84 5441 94
rect 5292 52 5348 80
rect 5378 52 5412 80
tri 5426 77 5433 84 ne
rect 5433 52 5441 84
rect 5471 52 5519 94
rect 5549 84 5574 94
rect 5549 52 5557 84
rect 5673 80 5698 94
rect 5578 52 5612 80
rect 5642 52 5698 80
rect 5728 52 5756 94
rect 5814 52 5842 94
rect 5872 80 5897 94
rect 5996 84 6021 94
rect 5872 52 5928 80
rect 5958 52 5992 80
tri 6006 77 6013 84 ne
rect 6013 52 6021 84
rect 6051 52 6099 94
rect 6129 84 6154 94
rect 6129 52 6137 84
rect 6253 80 6278 94
rect 6158 52 6192 80
rect 6222 52 6278 80
rect 6308 52 6336 94
rect 6394 52 6422 94
rect 6452 80 6477 94
rect 6576 84 6601 94
rect 6452 52 6508 80
rect 6538 52 6572 80
tri 6586 77 6593 84 ne
rect 6593 52 6601 84
rect 6631 52 6679 94
rect 6709 84 6734 94
rect 6709 52 6717 84
rect 6833 80 6858 94
rect 6738 52 6772 80
rect 6802 52 6858 80
rect 6888 52 6916 94
rect 165 28 192 52
rect 259 30 291 52
rect 259 28 261 30
rect 289 28 291 30
rect 358 28 385 52
rect 165 14 259 28
rect 291 14 385 28
rect 745 28 772 52
rect 839 30 871 52
rect 839 28 841 30
rect 869 28 871 30
rect 938 28 965 52
rect 745 14 839 28
rect 871 14 965 28
rect 1325 28 1352 52
rect 1419 30 1451 52
rect 1419 28 1421 30
rect 1449 28 1451 30
rect 1518 28 1545 52
rect 1325 14 1419 28
rect 1451 14 1545 28
rect 1905 28 1932 52
rect 1999 30 2031 52
rect 1999 28 2001 30
rect 2029 28 2031 30
rect 2098 28 2125 52
rect 1905 14 1999 28
rect 2031 14 2125 28
rect 2485 28 2512 52
rect 2579 30 2611 52
rect 2579 28 2581 30
rect 2609 28 2611 30
rect 2678 28 2705 52
rect 2485 14 2579 28
rect 2611 14 2705 28
rect 3065 28 3092 52
rect 3159 30 3191 52
rect 3159 28 3161 30
rect 3189 28 3191 30
rect 3258 28 3285 52
rect 3065 14 3159 28
rect 3191 14 3285 28
rect 3645 28 3672 52
rect 3739 30 3771 52
rect 3739 28 3741 30
rect 3769 28 3771 30
rect 3838 28 3865 52
rect 3645 14 3739 28
rect 3771 14 3865 28
rect 4225 28 4252 52
rect 4319 30 4351 52
rect 4319 28 4321 30
rect 4349 28 4351 30
rect 4418 28 4445 52
rect 4225 14 4319 28
rect 4351 14 4445 28
rect 4805 28 4832 52
rect 4899 30 4931 52
rect 4899 28 4901 30
rect 4929 28 4931 30
rect 4998 28 5025 52
rect 4805 14 4899 28
rect 4931 14 5025 28
rect 5385 28 5412 52
rect 5479 30 5511 52
rect 5479 28 5481 30
rect 5509 28 5511 30
rect 5578 28 5605 52
rect 5385 14 5479 28
rect 5511 14 5605 28
rect 5965 28 5992 52
rect 6059 30 6091 52
rect 6059 28 6061 30
rect 6089 28 6091 30
rect 6158 28 6185 52
rect 5965 14 6059 28
rect 6091 14 6185 28
rect 6545 28 6572 52
rect 6639 30 6671 52
rect 6639 28 6641 30
rect 6669 28 6671 30
rect 6738 28 6765 52
rect 6545 14 6639 28
rect 6671 14 6765 28
rect 88 -72 106 -44
rect 136 -72 154 -44
rect 396 -72 414 -44
rect 444 -72 463 -44
rect 668 -72 686 -44
rect 716 -72 734 -44
rect 976 -72 994 -44
rect 1024 -72 1043 -44
rect 1248 -72 1266 -44
rect 1296 -72 1314 -44
rect 1556 -72 1574 -44
rect 1604 -72 1623 -44
rect 1828 -72 1846 -44
rect 1876 -72 1894 -44
rect 2136 -72 2154 -44
rect 2184 -72 2203 -44
rect 2408 -72 2426 -44
rect 2456 -72 2474 -44
rect 2716 -72 2734 -44
rect 2764 -72 2783 -44
rect 2988 -72 3006 -44
rect 3036 -72 3054 -44
rect 3296 -72 3314 -44
rect 3344 -72 3363 -44
rect 3568 -72 3586 -44
rect 3616 -72 3634 -44
rect 3876 -72 3894 -44
rect 3924 -72 3943 -44
rect 4148 -72 4166 -44
rect 4196 -72 4214 -44
rect 4456 -72 4474 -44
rect 4504 -72 4523 -44
rect 4728 -72 4746 -44
rect 4776 -72 4794 -44
rect 5036 -72 5054 -44
rect 5084 -72 5103 -44
rect 5308 -72 5326 -44
rect 5356 -72 5374 -44
rect 5616 -72 5634 -44
rect 5664 -72 5683 -44
rect 5888 -72 5906 -44
rect 5936 -72 5954 -44
rect 6196 -72 6214 -44
rect 6244 -72 6263 -44
rect 6468 -72 6486 -44
rect 6516 -72 6534 -44
rect 6776 -72 6794 -44
rect 6824 -72 6843 -44
rect 14 -218 42 -176
rect 72 -190 97 -176
rect 196 -186 221 -176
rect 72 -218 128 -190
rect 158 -218 192 -190
tri 206 -193 213 -186 ne
rect 213 -218 221 -186
rect 251 -218 299 -176
rect 329 -186 354 -176
rect 329 -218 337 -186
rect 453 -190 478 -176
rect 358 -218 392 -190
rect 422 -218 478 -190
rect 508 -218 536 -176
rect 594 -218 622 -176
rect 652 -190 677 -176
rect 776 -186 801 -176
rect 652 -218 708 -190
rect 738 -218 772 -190
tri 786 -193 793 -186 ne
rect 793 -218 801 -186
rect 831 -218 879 -176
rect 909 -186 934 -176
rect 909 -218 917 -186
rect 1033 -190 1058 -176
rect 938 -218 972 -190
rect 1002 -218 1058 -190
rect 1088 -218 1116 -176
rect 1174 -218 1202 -176
rect 1232 -190 1257 -176
rect 1356 -186 1381 -176
rect 1232 -218 1288 -190
rect 1318 -218 1352 -190
tri 1366 -193 1373 -186 ne
rect 1373 -218 1381 -186
rect 1411 -218 1459 -176
rect 1489 -186 1514 -176
rect 1489 -218 1497 -186
rect 1613 -190 1638 -176
rect 1518 -218 1552 -190
rect 1582 -218 1638 -190
rect 1668 -218 1696 -176
rect 1754 -218 1782 -176
rect 1812 -190 1837 -176
rect 1936 -186 1961 -176
rect 1812 -218 1868 -190
rect 1898 -218 1932 -190
tri 1946 -193 1953 -186 ne
rect 1953 -218 1961 -186
rect 1991 -218 2039 -176
rect 2069 -186 2094 -176
rect 2069 -218 2077 -186
rect 2193 -190 2218 -176
rect 2098 -218 2132 -190
rect 2162 -218 2218 -190
rect 2248 -218 2276 -176
rect 2334 -218 2362 -176
rect 2392 -190 2417 -176
rect 2516 -186 2541 -176
rect 2392 -218 2448 -190
rect 2478 -218 2512 -190
tri 2526 -193 2533 -186 ne
rect 2533 -218 2541 -186
rect 2571 -218 2619 -176
rect 2649 -186 2674 -176
rect 2649 -218 2657 -186
rect 2773 -190 2798 -176
rect 2678 -218 2712 -190
rect 2742 -218 2798 -190
rect 2828 -218 2856 -176
rect 2914 -218 2942 -176
rect 2972 -190 2997 -176
rect 3096 -186 3121 -176
rect 2972 -218 3028 -190
rect 3058 -218 3092 -190
tri 3106 -193 3113 -186 ne
rect 3113 -218 3121 -186
rect 3151 -218 3199 -176
rect 3229 -186 3254 -176
rect 3229 -218 3237 -186
rect 3353 -190 3378 -176
rect 3258 -218 3292 -190
rect 3322 -218 3378 -190
rect 3408 -218 3436 -176
rect 3494 -218 3522 -176
rect 3552 -190 3577 -176
rect 3676 -186 3701 -176
rect 3552 -218 3608 -190
rect 3638 -218 3672 -190
tri 3686 -193 3693 -186 ne
rect 3693 -218 3701 -186
rect 3731 -218 3779 -176
rect 3809 -186 3834 -176
rect 3809 -218 3817 -186
rect 3933 -190 3958 -176
rect 3838 -218 3872 -190
rect 3902 -218 3958 -190
rect 3988 -218 4016 -176
rect 4074 -218 4102 -176
rect 4132 -190 4157 -176
rect 4256 -186 4281 -176
rect 4132 -218 4188 -190
rect 4218 -218 4252 -190
tri 4266 -193 4273 -186 ne
rect 4273 -218 4281 -186
rect 4311 -218 4359 -176
rect 4389 -186 4414 -176
rect 4389 -218 4397 -186
rect 4513 -190 4538 -176
rect 4418 -218 4452 -190
rect 4482 -218 4538 -190
rect 4568 -218 4596 -176
rect 4654 -218 4682 -176
rect 4712 -190 4737 -176
rect 4836 -186 4861 -176
rect 4712 -218 4768 -190
rect 4798 -218 4832 -190
tri 4846 -193 4853 -186 ne
rect 4853 -218 4861 -186
rect 4891 -218 4939 -176
rect 4969 -186 4994 -176
rect 4969 -218 4977 -186
rect 5093 -190 5118 -176
rect 4998 -218 5032 -190
rect 5062 -218 5118 -190
rect 5148 -218 5176 -176
rect 5234 -218 5262 -176
rect 5292 -190 5317 -176
rect 5416 -186 5441 -176
rect 5292 -218 5348 -190
rect 5378 -218 5412 -190
tri 5426 -193 5433 -186 ne
rect 5433 -218 5441 -186
rect 5471 -218 5519 -176
rect 5549 -186 5574 -176
rect 5549 -218 5557 -186
rect 5673 -190 5698 -176
rect 5578 -218 5612 -190
rect 5642 -218 5698 -190
rect 5728 -218 5756 -176
rect 5814 -218 5842 -176
rect 5872 -190 5897 -176
rect 5996 -186 6021 -176
rect 5872 -218 5928 -190
rect 5958 -218 5992 -190
tri 6006 -193 6013 -186 ne
rect 6013 -218 6021 -186
rect 6051 -218 6099 -176
rect 6129 -186 6154 -176
rect 6129 -218 6137 -186
rect 6253 -190 6278 -176
rect 6158 -218 6192 -190
rect 6222 -218 6278 -190
rect 6308 -218 6336 -176
rect 6394 -218 6422 -176
rect 6452 -190 6477 -176
rect 6576 -186 6601 -176
rect 6452 -218 6508 -190
rect 6538 -218 6572 -190
tri 6586 -193 6593 -186 ne
rect 6593 -218 6601 -186
rect 6631 -218 6679 -176
rect 6709 -186 6734 -176
rect 6709 -218 6717 -186
rect 6833 -190 6858 -176
rect 6738 -218 6772 -190
rect 6802 -218 6858 -190
rect 6888 -218 6916 -176
rect 165 -242 192 -218
rect 259 -240 291 -218
rect 259 -242 261 -240
rect 289 -242 291 -240
rect 358 -242 385 -218
rect 165 -256 259 -242
rect 291 -256 385 -242
rect 745 -242 772 -218
rect 839 -240 871 -218
rect 839 -242 841 -240
rect 869 -242 871 -240
rect 938 -242 965 -218
rect 745 -256 839 -242
rect 871 -256 965 -242
rect 1325 -242 1352 -218
rect 1419 -240 1451 -218
rect 1419 -242 1421 -240
rect 1449 -242 1451 -240
rect 1518 -242 1545 -218
rect 1325 -256 1419 -242
rect 1451 -256 1545 -242
rect 1905 -242 1932 -218
rect 1999 -240 2031 -218
rect 1999 -242 2001 -240
rect 2029 -242 2031 -240
rect 2098 -242 2125 -218
rect 1905 -256 1999 -242
rect 2031 -256 2125 -242
rect 2485 -242 2512 -218
rect 2579 -240 2611 -218
rect 2579 -242 2581 -240
rect 2609 -242 2611 -240
rect 2678 -242 2705 -218
rect 2485 -256 2579 -242
rect 2611 -256 2705 -242
rect 3065 -242 3092 -218
rect 3159 -240 3191 -218
rect 3159 -242 3161 -240
rect 3189 -242 3191 -240
rect 3258 -242 3285 -218
rect 3065 -256 3159 -242
rect 3191 -256 3285 -242
rect 3645 -242 3672 -218
rect 3739 -240 3771 -218
rect 3739 -242 3741 -240
rect 3769 -242 3771 -240
rect 3838 -242 3865 -218
rect 3645 -256 3739 -242
rect 3771 -256 3865 -242
rect 4225 -242 4252 -218
rect 4319 -240 4351 -218
rect 4319 -242 4321 -240
rect 4349 -242 4351 -240
rect 4418 -242 4445 -218
rect 4225 -256 4319 -242
rect 4351 -256 4445 -242
rect 4805 -242 4832 -218
rect 4899 -240 4931 -218
rect 4899 -242 4901 -240
rect 4929 -242 4931 -240
rect 4998 -242 5025 -218
rect 4805 -256 4899 -242
rect 4931 -256 5025 -242
rect 5385 -242 5412 -218
rect 5479 -240 5511 -218
rect 5479 -242 5481 -240
rect 5509 -242 5511 -240
rect 5578 -242 5605 -218
rect 5385 -256 5479 -242
rect 5511 -256 5605 -242
rect 5965 -242 5992 -218
rect 6059 -240 6091 -218
rect 6059 -242 6061 -240
rect 6089 -242 6091 -240
rect 6158 -242 6185 -218
rect 5965 -256 6059 -242
rect 6091 -256 6185 -242
rect 6545 -242 6572 -218
rect 6639 -240 6671 -218
rect 6639 -242 6641 -240
rect 6669 -242 6671 -240
rect 6738 -242 6765 -218
rect 6545 -256 6639 -242
rect 6671 -256 6765 -242
rect 88 -342 106 -314
rect 136 -342 154 -314
rect 396 -342 414 -314
rect 444 -342 463 -314
rect 668 -342 686 -314
rect 716 -342 734 -314
rect 976 -342 994 -314
rect 1024 -342 1043 -314
rect 1248 -342 1266 -314
rect 1296 -342 1314 -314
rect 1556 -342 1574 -314
rect 1604 -342 1623 -314
rect 1828 -342 1846 -314
rect 1876 -342 1894 -314
rect 2136 -342 2154 -314
rect 2184 -342 2203 -314
rect 2408 -342 2426 -314
rect 2456 -342 2474 -314
rect 2716 -342 2734 -314
rect 2764 -342 2783 -314
rect 2988 -342 3006 -314
rect 3036 -342 3054 -314
rect 3296 -342 3314 -314
rect 3344 -342 3363 -314
rect 3568 -342 3586 -314
rect 3616 -342 3634 -314
rect 3876 -342 3894 -314
rect 3924 -342 3943 -314
rect 4148 -342 4166 -314
rect 4196 -342 4214 -314
rect 4456 -342 4474 -314
rect 4504 -342 4523 -314
rect 4728 -342 4746 -314
rect 4776 -342 4794 -314
rect 5036 -342 5054 -314
rect 5084 -342 5103 -314
rect 5308 -342 5326 -314
rect 5356 -342 5374 -314
rect 5616 -342 5634 -314
rect 5664 -342 5683 -314
rect 5888 -342 5906 -314
rect 5936 -342 5954 -314
rect 6196 -342 6214 -314
rect 6244 -342 6263 -314
rect 6468 -342 6486 -314
rect 6516 -342 6534 -314
rect 6776 -342 6794 -314
rect 6824 -342 6843 -314
rect 14 -488 42 -446
rect 72 -460 97 -446
rect 196 -456 221 -446
rect 72 -488 128 -460
rect 158 -488 192 -460
tri 206 -463 213 -456 ne
rect 213 -488 221 -456
rect 251 -488 299 -446
rect 329 -456 354 -446
rect 329 -488 337 -456
rect 453 -460 478 -446
rect 358 -488 392 -460
rect 422 -488 478 -460
rect 508 -488 536 -446
rect 594 -488 622 -446
rect 652 -460 677 -446
rect 776 -456 801 -446
rect 652 -488 708 -460
rect 738 -488 772 -460
tri 786 -463 793 -456 ne
rect 793 -488 801 -456
rect 831 -488 879 -446
rect 909 -456 934 -446
rect 909 -488 917 -456
rect 1033 -460 1058 -446
rect 938 -488 972 -460
rect 1002 -488 1058 -460
rect 1088 -488 1116 -446
rect 1174 -488 1202 -446
rect 1232 -460 1257 -446
rect 1356 -456 1381 -446
rect 1232 -488 1288 -460
rect 1318 -488 1352 -460
tri 1366 -463 1373 -456 ne
rect 1373 -488 1381 -456
rect 1411 -488 1459 -446
rect 1489 -456 1514 -446
rect 1489 -488 1497 -456
rect 1613 -460 1638 -446
rect 1518 -488 1552 -460
rect 1582 -488 1638 -460
rect 1668 -488 1696 -446
rect 1754 -488 1782 -446
rect 1812 -460 1837 -446
rect 1936 -456 1961 -446
rect 1812 -488 1868 -460
rect 1898 -488 1932 -460
tri 1946 -463 1953 -456 ne
rect 1953 -488 1961 -456
rect 1991 -488 2039 -446
rect 2069 -456 2094 -446
rect 2069 -488 2077 -456
rect 2193 -460 2218 -446
rect 2098 -488 2132 -460
rect 2162 -488 2218 -460
rect 2248 -488 2276 -446
rect 2334 -488 2362 -446
rect 2392 -460 2417 -446
rect 2516 -456 2541 -446
rect 2392 -488 2448 -460
rect 2478 -488 2512 -460
tri 2526 -463 2533 -456 ne
rect 2533 -488 2541 -456
rect 2571 -488 2619 -446
rect 2649 -456 2674 -446
rect 2649 -488 2657 -456
rect 2773 -460 2798 -446
rect 2678 -488 2712 -460
rect 2742 -488 2798 -460
rect 2828 -488 2856 -446
rect 2914 -488 2942 -446
rect 2972 -460 2997 -446
rect 3096 -456 3121 -446
rect 2972 -488 3028 -460
rect 3058 -488 3092 -460
tri 3106 -463 3113 -456 ne
rect 3113 -488 3121 -456
rect 3151 -488 3199 -446
rect 3229 -456 3254 -446
rect 3229 -488 3237 -456
rect 3353 -460 3378 -446
rect 3258 -488 3292 -460
rect 3322 -488 3378 -460
rect 3408 -488 3436 -446
rect 3494 -488 3522 -446
rect 3552 -460 3577 -446
rect 3676 -456 3701 -446
rect 3552 -488 3608 -460
rect 3638 -488 3672 -460
tri 3686 -463 3693 -456 ne
rect 3693 -488 3701 -456
rect 3731 -488 3779 -446
rect 3809 -456 3834 -446
rect 3809 -488 3817 -456
rect 3933 -460 3958 -446
rect 3838 -488 3872 -460
rect 3902 -488 3958 -460
rect 3988 -488 4016 -446
rect 4074 -488 4102 -446
rect 4132 -460 4157 -446
rect 4256 -456 4281 -446
rect 4132 -488 4188 -460
rect 4218 -488 4252 -460
tri 4266 -463 4273 -456 ne
rect 4273 -488 4281 -456
rect 4311 -488 4359 -446
rect 4389 -456 4414 -446
rect 4389 -488 4397 -456
rect 4513 -460 4538 -446
rect 4418 -488 4452 -460
rect 4482 -488 4538 -460
rect 4568 -488 4596 -446
rect 4654 -488 4682 -446
rect 4712 -460 4737 -446
rect 4836 -456 4861 -446
rect 4712 -488 4768 -460
rect 4798 -488 4832 -460
tri 4846 -463 4853 -456 ne
rect 4853 -488 4861 -456
rect 4891 -488 4939 -446
rect 4969 -456 4994 -446
rect 4969 -488 4977 -456
rect 5093 -460 5118 -446
rect 4998 -488 5032 -460
rect 5062 -488 5118 -460
rect 5148 -488 5176 -446
rect 5234 -488 5262 -446
rect 5292 -460 5317 -446
rect 5416 -456 5441 -446
rect 5292 -488 5348 -460
rect 5378 -488 5412 -460
tri 5426 -463 5433 -456 ne
rect 5433 -488 5441 -456
rect 5471 -488 5519 -446
rect 5549 -456 5574 -446
rect 5549 -488 5557 -456
rect 5673 -460 5698 -446
rect 5578 -488 5612 -460
rect 5642 -488 5698 -460
rect 5728 -488 5756 -446
rect 5814 -488 5842 -446
rect 5872 -460 5897 -446
rect 5996 -456 6021 -446
rect 5872 -488 5928 -460
rect 5958 -488 5992 -460
tri 6006 -463 6013 -456 ne
rect 6013 -488 6021 -456
rect 6051 -488 6099 -446
rect 6129 -456 6154 -446
rect 6129 -488 6137 -456
rect 6253 -460 6278 -446
rect 6158 -488 6192 -460
rect 6222 -488 6278 -460
rect 6308 -488 6336 -446
rect 6394 -488 6422 -446
rect 6452 -460 6477 -446
rect 6576 -456 6601 -446
rect 6452 -488 6508 -460
rect 6538 -488 6572 -460
tri 6586 -463 6593 -456 ne
rect 6593 -488 6601 -456
rect 6631 -488 6679 -446
rect 6709 -456 6734 -446
rect 6709 -488 6717 -456
rect 6833 -460 6858 -446
rect 6738 -488 6772 -460
rect 6802 -488 6858 -460
rect 6888 -488 6916 -446
rect 165 -512 192 -488
rect 259 -510 291 -488
rect 259 -512 261 -510
rect 289 -512 291 -510
rect 358 -512 385 -488
rect 165 -526 259 -512
rect 291 -526 385 -512
rect 745 -512 772 -488
rect 839 -510 871 -488
rect 839 -512 841 -510
rect 869 -512 871 -510
rect 938 -512 965 -488
rect 745 -526 839 -512
rect 871 -526 965 -512
rect 1325 -512 1352 -488
rect 1419 -510 1451 -488
rect 1419 -512 1421 -510
rect 1449 -512 1451 -510
rect 1518 -512 1545 -488
rect 1325 -526 1419 -512
rect 1451 -526 1545 -512
rect 1905 -512 1932 -488
rect 1999 -510 2031 -488
rect 1999 -512 2001 -510
rect 2029 -512 2031 -510
rect 2098 -512 2125 -488
rect 1905 -526 1999 -512
rect 2031 -526 2125 -512
rect 2485 -512 2512 -488
rect 2579 -510 2611 -488
rect 2579 -512 2581 -510
rect 2609 -512 2611 -510
rect 2678 -512 2705 -488
rect 2485 -526 2579 -512
rect 2611 -526 2705 -512
rect 3065 -512 3092 -488
rect 3159 -510 3191 -488
rect 3159 -512 3161 -510
rect 3189 -512 3191 -510
rect 3258 -512 3285 -488
rect 3065 -526 3159 -512
rect 3191 -526 3285 -512
rect 3645 -512 3672 -488
rect 3739 -510 3771 -488
rect 3739 -512 3741 -510
rect 3769 -512 3771 -510
rect 3838 -512 3865 -488
rect 3645 -526 3739 -512
rect 3771 -526 3865 -512
rect 4225 -512 4252 -488
rect 4319 -510 4351 -488
rect 4319 -512 4321 -510
rect 4349 -512 4351 -510
rect 4418 -512 4445 -488
rect 4225 -526 4319 -512
rect 4351 -526 4445 -512
rect 4805 -512 4832 -488
rect 4899 -510 4931 -488
rect 4899 -512 4901 -510
rect 4929 -512 4931 -510
rect 4998 -512 5025 -488
rect 4805 -526 4899 -512
rect 4931 -526 5025 -512
rect 5385 -512 5412 -488
rect 5479 -510 5511 -488
rect 5479 -512 5481 -510
rect 5509 -512 5511 -510
rect 5578 -512 5605 -488
rect 5385 -526 5479 -512
rect 5511 -526 5605 -512
rect 5965 -512 5992 -488
rect 6059 -510 6091 -488
rect 6059 -512 6061 -510
rect 6089 -512 6091 -510
rect 6158 -512 6185 -488
rect 5965 -526 6059 -512
rect 6091 -526 6185 -512
rect 6545 -512 6572 -488
rect 6639 -510 6671 -488
rect 6639 -512 6641 -510
rect 6669 -512 6671 -510
rect 6738 -512 6765 -488
rect 6545 -526 6639 -512
rect 6671 -526 6765 -512
rect 88 -612 106 -584
rect 136 -612 154 -584
rect 396 -612 414 -584
rect 444 -612 463 -584
rect 668 -612 686 -584
rect 716 -612 734 -584
rect 976 -612 994 -584
rect 1024 -612 1043 -584
rect 1248 -612 1266 -584
rect 1296 -612 1314 -584
rect 1556 -612 1574 -584
rect 1604 -612 1623 -584
rect 1828 -612 1846 -584
rect 1876 -612 1894 -584
rect 2136 -612 2154 -584
rect 2184 -612 2203 -584
rect 2408 -612 2426 -584
rect 2456 -612 2474 -584
rect 2716 -612 2734 -584
rect 2764 -612 2783 -584
rect 2988 -612 3006 -584
rect 3036 -612 3054 -584
rect 3296 -612 3314 -584
rect 3344 -612 3363 -584
rect 3568 -612 3586 -584
rect 3616 -612 3634 -584
rect 3876 -612 3894 -584
rect 3924 -612 3943 -584
rect 4148 -612 4166 -584
rect 4196 -612 4214 -584
rect 4456 -612 4474 -584
rect 4504 -612 4523 -584
rect 4728 -612 4746 -584
rect 4776 -612 4794 -584
rect 5036 -612 5054 -584
rect 5084 -612 5103 -584
rect 5308 -612 5326 -584
rect 5356 -612 5374 -584
rect 5616 -612 5634 -584
rect 5664 -612 5683 -584
rect 5888 -612 5906 -584
rect 5936 -612 5954 -584
rect 6196 -612 6214 -584
rect 6244 -612 6263 -584
rect 6468 -612 6486 -584
rect 6516 -612 6534 -584
rect 6776 -612 6794 -584
rect 6824 -612 6843 -584
rect 14 -758 42 -716
rect 72 -730 97 -716
rect 196 -726 221 -716
rect 72 -758 128 -730
rect 158 -758 192 -730
tri 206 -733 213 -726 ne
rect 213 -758 221 -726
rect 251 -758 299 -716
rect 329 -726 354 -716
rect 329 -758 337 -726
rect 453 -730 478 -716
rect 358 -758 392 -730
rect 422 -758 478 -730
rect 508 -758 536 -716
rect 594 -758 622 -716
rect 652 -730 677 -716
rect 776 -726 801 -716
rect 652 -758 708 -730
rect 738 -758 772 -730
tri 786 -733 793 -726 ne
rect 793 -758 801 -726
rect 831 -758 879 -716
rect 909 -726 934 -716
rect 909 -758 917 -726
rect 1033 -730 1058 -716
rect 938 -758 972 -730
rect 1002 -758 1058 -730
rect 1088 -758 1116 -716
rect 1174 -758 1202 -716
rect 1232 -730 1257 -716
rect 1356 -726 1381 -716
rect 1232 -758 1288 -730
rect 1318 -758 1352 -730
tri 1366 -733 1373 -726 ne
rect 1373 -758 1381 -726
rect 1411 -758 1459 -716
rect 1489 -726 1514 -716
rect 1489 -758 1497 -726
rect 1613 -730 1638 -716
rect 1518 -758 1552 -730
rect 1582 -758 1638 -730
rect 1668 -758 1696 -716
rect 1754 -758 1782 -716
rect 1812 -730 1837 -716
rect 1936 -726 1961 -716
rect 1812 -758 1868 -730
rect 1898 -758 1932 -730
tri 1946 -733 1953 -726 ne
rect 1953 -758 1961 -726
rect 1991 -758 2039 -716
rect 2069 -726 2094 -716
rect 2069 -758 2077 -726
rect 2193 -730 2218 -716
rect 2098 -758 2132 -730
rect 2162 -758 2218 -730
rect 2248 -758 2276 -716
rect 2334 -758 2362 -716
rect 2392 -730 2417 -716
rect 2516 -726 2541 -716
rect 2392 -758 2448 -730
rect 2478 -758 2512 -730
tri 2526 -733 2533 -726 ne
rect 2533 -758 2541 -726
rect 2571 -758 2619 -716
rect 2649 -726 2674 -716
rect 2649 -758 2657 -726
rect 2773 -730 2798 -716
rect 2678 -758 2712 -730
rect 2742 -758 2798 -730
rect 2828 -758 2856 -716
rect 2914 -758 2942 -716
rect 2972 -730 2997 -716
rect 3096 -726 3121 -716
rect 2972 -758 3028 -730
rect 3058 -758 3092 -730
tri 3106 -733 3113 -726 ne
rect 3113 -758 3121 -726
rect 3151 -758 3199 -716
rect 3229 -726 3254 -716
rect 3229 -758 3237 -726
rect 3353 -730 3378 -716
rect 3258 -758 3292 -730
rect 3322 -758 3378 -730
rect 3408 -758 3436 -716
rect 3494 -758 3522 -716
rect 3552 -730 3577 -716
rect 3676 -726 3701 -716
rect 3552 -758 3608 -730
rect 3638 -758 3672 -730
tri 3686 -733 3693 -726 ne
rect 3693 -758 3701 -726
rect 3731 -758 3779 -716
rect 3809 -726 3834 -716
rect 3809 -758 3817 -726
rect 3933 -730 3958 -716
rect 3838 -758 3872 -730
rect 3902 -758 3958 -730
rect 3988 -758 4016 -716
rect 4074 -758 4102 -716
rect 4132 -730 4157 -716
rect 4256 -726 4281 -716
rect 4132 -758 4188 -730
rect 4218 -758 4252 -730
tri 4266 -733 4273 -726 ne
rect 4273 -758 4281 -726
rect 4311 -758 4359 -716
rect 4389 -726 4414 -716
rect 4389 -758 4397 -726
rect 4513 -730 4538 -716
rect 4418 -758 4452 -730
rect 4482 -758 4538 -730
rect 4568 -758 4596 -716
rect 4654 -758 4682 -716
rect 4712 -730 4737 -716
rect 4836 -726 4861 -716
rect 4712 -758 4768 -730
rect 4798 -758 4832 -730
tri 4846 -733 4853 -726 ne
rect 4853 -758 4861 -726
rect 4891 -758 4939 -716
rect 4969 -726 4994 -716
rect 4969 -758 4977 -726
rect 5093 -730 5118 -716
rect 4998 -758 5032 -730
rect 5062 -758 5118 -730
rect 5148 -758 5176 -716
rect 5234 -758 5262 -716
rect 5292 -730 5317 -716
rect 5416 -726 5441 -716
rect 5292 -758 5348 -730
rect 5378 -758 5412 -730
tri 5426 -733 5433 -726 ne
rect 5433 -758 5441 -726
rect 5471 -758 5519 -716
rect 5549 -726 5574 -716
rect 5549 -758 5557 -726
rect 5673 -730 5698 -716
rect 5578 -758 5612 -730
rect 5642 -758 5698 -730
rect 5728 -758 5756 -716
rect 5814 -758 5842 -716
rect 5872 -730 5897 -716
rect 5996 -726 6021 -716
rect 5872 -758 5928 -730
rect 5958 -758 5992 -730
tri 6006 -733 6013 -726 ne
rect 6013 -758 6021 -726
rect 6051 -758 6099 -716
rect 6129 -726 6154 -716
rect 6129 -758 6137 -726
rect 6253 -730 6278 -716
rect 6158 -758 6192 -730
rect 6222 -758 6278 -730
rect 6308 -758 6336 -716
rect 6394 -758 6422 -716
rect 6452 -730 6477 -716
rect 6576 -726 6601 -716
rect 6452 -758 6508 -730
rect 6538 -758 6572 -730
tri 6586 -733 6593 -726 ne
rect 6593 -758 6601 -726
rect 6631 -758 6679 -716
rect 6709 -726 6734 -716
rect 6709 -758 6717 -726
rect 6833 -730 6858 -716
rect 6738 -758 6772 -730
rect 6802 -758 6858 -730
rect 6888 -758 6916 -716
rect 165 -782 192 -758
rect 259 -780 291 -758
rect 259 -782 261 -780
rect 289 -782 291 -780
rect 358 -782 385 -758
rect 165 -796 259 -782
rect 291 -796 385 -782
rect 745 -782 772 -758
rect 839 -780 871 -758
rect 839 -782 841 -780
rect 869 -782 871 -780
rect 938 -782 965 -758
rect 745 -796 839 -782
rect 871 -796 965 -782
rect 1325 -782 1352 -758
rect 1419 -780 1451 -758
rect 1419 -782 1421 -780
rect 1449 -782 1451 -780
rect 1518 -782 1545 -758
rect 1325 -796 1419 -782
rect 1451 -796 1545 -782
rect 1905 -782 1932 -758
rect 1999 -780 2031 -758
rect 1999 -782 2001 -780
rect 2029 -782 2031 -780
rect 2098 -782 2125 -758
rect 1905 -796 1999 -782
rect 2031 -796 2125 -782
rect 2485 -782 2512 -758
rect 2579 -780 2611 -758
rect 2579 -782 2581 -780
rect 2609 -782 2611 -780
rect 2678 -782 2705 -758
rect 2485 -796 2579 -782
rect 2611 -796 2705 -782
rect 3065 -782 3092 -758
rect 3159 -780 3191 -758
rect 3159 -782 3161 -780
rect 3189 -782 3191 -780
rect 3258 -782 3285 -758
rect 3065 -796 3159 -782
rect 3191 -796 3285 -782
rect 3645 -782 3672 -758
rect 3739 -780 3771 -758
rect 3739 -782 3741 -780
rect 3769 -782 3771 -780
rect 3838 -782 3865 -758
rect 3645 -796 3739 -782
rect 3771 -796 3865 -782
rect 4225 -782 4252 -758
rect 4319 -780 4351 -758
rect 4319 -782 4321 -780
rect 4349 -782 4351 -780
rect 4418 -782 4445 -758
rect 4225 -796 4319 -782
rect 4351 -796 4445 -782
rect 4805 -782 4832 -758
rect 4899 -780 4931 -758
rect 4899 -782 4901 -780
rect 4929 -782 4931 -780
rect 4998 -782 5025 -758
rect 4805 -796 4899 -782
rect 4931 -796 5025 -782
rect 5385 -782 5412 -758
rect 5479 -780 5511 -758
rect 5479 -782 5481 -780
rect 5509 -782 5511 -780
rect 5578 -782 5605 -758
rect 5385 -796 5479 -782
rect 5511 -796 5605 -782
rect 5965 -782 5992 -758
rect 6059 -780 6091 -758
rect 6059 -782 6061 -780
rect 6089 -782 6091 -780
rect 6158 -782 6185 -758
rect 5965 -796 6059 -782
rect 6091 -796 6185 -782
rect 6545 -782 6572 -758
rect 6639 -780 6671 -758
rect 6639 -782 6641 -780
rect 6669 -782 6671 -780
rect 6738 -782 6765 -758
rect 6545 -796 6639 -782
rect 6671 -796 6765 -782
rect 88 -882 106 -854
rect 136 -882 154 -854
rect 396 -882 414 -854
rect 444 -882 463 -854
rect 668 -882 686 -854
rect 716 -882 734 -854
rect 976 -882 994 -854
rect 1024 -882 1043 -854
rect 1248 -882 1266 -854
rect 1296 -882 1314 -854
rect 1556 -882 1574 -854
rect 1604 -882 1623 -854
rect 1828 -882 1846 -854
rect 1876 -882 1894 -854
rect 2136 -882 2154 -854
rect 2184 -882 2203 -854
rect 2408 -882 2426 -854
rect 2456 -882 2474 -854
rect 2716 -882 2734 -854
rect 2764 -882 2783 -854
rect 2988 -882 3006 -854
rect 3036 -882 3054 -854
rect 3296 -882 3314 -854
rect 3344 -882 3363 -854
rect 3568 -882 3586 -854
rect 3616 -882 3634 -854
rect 3876 -882 3894 -854
rect 3924 -882 3943 -854
rect 4148 -882 4166 -854
rect 4196 -882 4214 -854
rect 4456 -882 4474 -854
rect 4504 -882 4523 -854
rect 4728 -882 4746 -854
rect 4776 -882 4794 -854
rect 5036 -882 5054 -854
rect 5084 -882 5103 -854
rect 5308 -882 5326 -854
rect 5356 -882 5374 -854
rect 5616 -882 5634 -854
rect 5664 -882 5683 -854
rect 5888 -882 5906 -854
rect 5936 -882 5954 -854
rect 6196 -882 6214 -854
rect 6244 -882 6263 -854
rect 6468 -882 6486 -854
rect 6516 -882 6534 -854
rect 6776 -882 6794 -854
rect 6824 -882 6843 -854
rect 14 -1028 42 -986
rect 72 -1000 97 -986
rect 196 -996 221 -986
rect 72 -1028 128 -1000
rect 158 -1028 192 -1000
tri 206 -1003 213 -996 ne
rect 213 -1028 221 -996
rect 251 -1028 299 -986
rect 329 -996 354 -986
rect 329 -1028 337 -996
rect 453 -1000 478 -986
rect 358 -1028 392 -1000
rect 422 -1028 478 -1000
rect 508 -1028 536 -986
rect 594 -1028 622 -986
rect 652 -1000 677 -986
rect 776 -996 801 -986
rect 652 -1028 708 -1000
rect 738 -1028 772 -1000
tri 786 -1003 793 -996 ne
rect 793 -1028 801 -996
rect 831 -1028 879 -986
rect 909 -996 934 -986
rect 909 -1028 917 -996
rect 1033 -1000 1058 -986
rect 938 -1028 972 -1000
rect 1002 -1028 1058 -1000
rect 1088 -1028 1116 -986
rect 1174 -1028 1202 -986
rect 1232 -1000 1257 -986
rect 1356 -996 1381 -986
rect 1232 -1028 1288 -1000
rect 1318 -1028 1352 -1000
tri 1366 -1003 1373 -996 ne
rect 1373 -1028 1381 -996
rect 1411 -1028 1459 -986
rect 1489 -996 1514 -986
rect 1489 -1028 1497 -996
rect 1613 -1000 1638 -986
rect 1518 -1028 1552 -1000
rect 1582 -1028 1638 -1000
rect 1668 -1028 1696 -986
rect 1754 -1028 1782 -986
rect 1812 -1000 1837 -986
rect 1936 -996 1961 -986
rect 1812 -1028 1868 -1000
rect 1898 -1028 1932 -1000
tri 1946 -1003 1953 -996 ne
rect 1953 -1028 1961 -996
rect 1991 -1028 2039 -986
rect 2069 -996 2094 -986
rect 2069 -1028 2077 -996
rect 2193 -1000 2218 -986
rect 2098 -1028 2132 -1000
rect 2162 -1028 2218 -1000
rect 2248 -1028 2276 -986
rect 2334 -1028 2362 -986
rect 2392 -1000 2417 -986
rect 2516 -996 2541 -986
rect 2392 -1028 2448 -1000
rect 2478 -1028 2512 -1000
tri 2526 -1003 2533 -996 ne
rect 2533 -1028 2541 -996
rect 2571 -1028 2619 -986
rect 2649 -996 2674 -986
rect 2649 -1028 2657 -996
rect 2773 -1000 2798 -986
rect 2678 -1028 2712 -1000
rect 2742 -1028 2798 -1000
rect 2828 -1028 2856 -986
rect 2914 -1028 2942 -986
rect 2972 -1000 2997 -986
rect 3096 -996 3121 -986
rect 2972 -1028 3028 -1000
rect 3058 -1028 3092 -1000
tri 3106 -1003 3113 -996 ne
rect 3113 -1028 3121 -996
rect 3151 -1028 3199 -986
rect 3229 -996 3254 -986
rect 3229 -1028 3237 -996
rect 3353 -1000 3378 -986
rect 3258 -1028 3292 -1000
rect 3322 -1028 3378 -1000
rect 3408 -1028 3436 -986
rect 3494 -1028 3522 -986
rect 3552 -1000 3577 -986
rect 3676 -996 3701 -986
rect 3552 -1028 3608 -1000
rect 3638 -1028 3672 -1000
tri 3686 -1003 3693 -996 ne
rect 3693 -1028 3701 -996
rect 3731 -1028 3779 -986
rect 3809 -996 3834 -986
rect 3809 -1028 3817 -996
rect 3933 -1000 3958 -986
rect 3838 -1028 3872 -1000
rect 3902 -1028 3958 -1000
rect 3988 -1028 4016 -986
rect 4074 -1028 4102 -986
rect 4132 -1000 4157 -986
rect 4256 -996 4281 -986
rect 4132 -1028 4188 -1000
rect 4218 -1028 4252 -1000
tri 4266 -1003 4273 -996 ne
rect 4273 -1028 4281 -996
rect 4311 -1028 4359 -986
rect 4389 -996 4414 -986
rect 4389 -1028 4397 -996
rect 4513 -1000 4538 -986
rect 4418 -1028 4452 -1000
rect 4482 -1028 4538 -1000
rect 4568 -1028 4596 -986
rect 4654 -1028 4682 -986
rect 4712 -1000 4737 -986
rect 4836 -996 4861 -986
rect 4712 -1028 4768 -1000
rect 4798 -1028 4832 -1000
tri 4846 -1003 4853 -996 ne
rect 4853 -1028 4861 -996
rect 4891 -1028 4939 -986
rect 4969 -996 4994 -986
rect 4969 -1028 4977 -996
rect 5093 -1000 5118 -986
rect 4998 -1028 5032 -1000
rect 5062 -1028 5118 -1000
rect 5148 -1028 5176 -986
rect 5234 -1028 5262 -986
rect 5292 -1000 5317 -986
rect 5416 -996 5441 -986
rect 5292 -1028 5348 -1000
rect 5378 -1028 5412 -1000
tri 5426 -1003 5433 -996 ne
rect 5433 -1028 5441 -996
rect 5471 -1028 5519 -986
rect 5549 -996 5574 -986
rect 5549 -1028 5557 -996
rect 5673 -1000 5698 -986
rect 5578 -1028 5612 -1000
rect 5642 -1028 5698 -1000
rect 5728 -1028 5756 -986
rect 5814 -1028 5842 -986
rect 5872 -1000 5897 -986
rect 5996 -996 6021 -986
rect 5872 -1028 5928 -1000
rect 5958 -1028 5992 -1000
tri 6006 -1003 6013 -996 ne
rect 6013 -1028 6021 -996
rect 6051 -1028 6099 -986
rect 6129 -996 6154 -986
rect 6129 -1028 6137 -996
rect 6253 -1000 6278 -986
rect 6158 -1028 6192 -1000
rect 6222 -1028 6278 -1000
rect 6308 -1028 6336 -986
rect 6394 -1028 6422 -986
rect 6452 -1000 6477 -986
rect 6576 -996 6601 -986
rect 6452 -1028 6508 -1000
rect 6538 -1028 6572 -1000
tri 6586 -1003 6593 -996 ne
rect 6593 -1028 6601 -996
rect 6631 -1028 6679 -986
rect 6709 -996 6734 -986
rect 6709 -1028 6717 -996
rect 6833 -1000 6858 -986
rect 6738 -1028 6772 -1000
rect 6802 -1028 6858 -1000
rect 6888 -1028 6916 -986
rect 165 -1052 192 -1028
rect 259 -1050 291 -1028
rect 259 -1052 261 -1050
rect 289 -1052 291 -1050
rect 358 -1052 385 -1028
rect 165 -1066 259 -1052
rect 291 -1066 385 -1052
rect 745 -1052 772 -1028
rect 839 -1050 871 -1028
rect 839 -1052 841 -1050
rect 869 -1052 871 -1050
rect 938 -1052 965 -1028
rect 745 -1066 839 -1052
rect 871 -1066 965 -1052
rect 1325 -1052 1352 -1028
rect 1419 -1050 1451 -1028
rect 1419 -1052 1421 -1050
rect 1449 -1052 1451 -1050
rect 1518 -1052 1545 -1028
rect 1325 -1066 1419 -1052
rect 1451 -1066 1545 -1052
rect 1905 -1052 1932 -1028
rect 1999 -1050 2031 -1028
rect 1999 -1052 2001 -1050
rect 2029 -1052 2031 -1050
rect 2098 -1052 2125 -1028
rect 1905 -1066 1999 -1052
rect 2031 -1066 2125 -1052
rect 2485 -1052 2512 -1028
rect 2579 -1050 2611 -1028
rect 2579 -1052 2581 -1050
rect 2609 -1052 2611 -1050
rect 2678 -1052 2705 -1028
rect 2485 -1066 2579 -1052
rect 2611 -1066 2705 -1052
rect 3065 -1052 3092 -1028
rect 3159 -1050 3191 -1028
rect 3159 -1052 3161 -1050
rect 3189 -1052 3191 -1050
rect 3258 -1052 3285 -1028
rect 3065 -1066 3159 -1052
rect 3191 -1066 3285 -1052
rect 3645 -1052 3672 -1028
rect 3739 -1050 3771 -1028
rect 3739 -1052 3741 -1050
rect 3769 -1052 3771 -1050
rect 3838 -1052 3865 -1028
rect 3645 -1066 3739 -1052
rect 3771 -1066 3865 -1052
rect 4225 -1052 4252 -1028
rect 4319 -1050 4351 -1028
rect 4319 -1052 4321 -1050
rect 4349 -1052 4351 -1050
rect 4418 -1052 4445 -1028
rect 4225 -1066 4319 -1052
rect 4351 -1066 4445 -1052
rect 4805 -1052 4832 -1028
rect 4899 -1050 4931 -1028
rect 4899 -1052 4901 -1050
rect 4929 -1052 4931 -1050
rect 4998 -1052 5025 -1028
rect 4805 -1066 4899 -1052
rect 4931 -1066 5025 -1052
rect 5385 -1052 5412 -1028
rect 5479 -1050 5511 -1028
rect 5479 -1052 5481 -1050
rect 5509 -1052 5511 -1050
rect 5578 -1052 5605 -1028
rect 5385 -1066 5479 -1052
rect 5511 -1066 5605 -1052
rect 5965 -1052 5992 -1028
rect 6059 -1050 6091 -1028
rect 6059 -1052 6061 -1050
rect 6089 -1052 6091 -1050
rect 6158 -1052 6185 -1028
rect 5965 -1066 6059 -1052
rect 6091 -1066 6185 -1052
rect 6545 -1052 6572 -1028
rect 6639 -1050 6671 -1028
rect 6639 -1052 6641 -1050
rect 6669 -1052 6671 -1050
rect 6738 -1052 6765 -1028
rect 6545 -1066 6639 -1052
rect 6671 -1066 6765 -1052
rect 88 -1152 106 -1124
rect 136 -1152 154 -1124
rect 396 -1152 414 -1124
rect 444 -1152 463 -1124
rect 668 -1152 686 -1124
rect 716 -1152 734 -1124
rect 976 -1152 994 -1124
rect 1024 -1152 1043 -1124
rect 1248 -1152 1266 -1124
rect 1296 -1152 1314 -1124
rect 1556 -1152 1574 -1124
rect 1604 -1152 1623 -1124
rect 1828 -1152 1846 -1124
rect 1876 -1152 1894 -1124
rect 2136 -1152 2154 -1124
rect 2184 -1152 2203 -1124
rect 2408 -1152 2426 -1124
rect 2456 -1152 2474 -1124
rect 2716 -1152 2734 -1124
rect 2764 -1152 2783 -1124
rect 2988 -1152 3006 -1124
rect 3036 -1152 3054 -1124
rect 3296 -1152 3314 -1124
rect 3344 -1152 3363 -1124
rect 3568 -1152 3586 -1124
rect 3616 -1152 3634 -1124
rect 3876 -1152 3894 -1124
rect 3924 -1152 3943 -1124
rect 4148 -1152 4166 -1124
rect 4196 -1152 4214 -1124
rect 4456 -1152 4474 -1124
rect 4504 -1152 4523 -1124
rect 4728 -1152 4746 -1124
rect 4776 -1152 4794 -1124
rect 5036 -1152 5054 -1124
rect 5084 -1152 5103 -1124
rect 5308 -1152 5326 -1124
rect 5356 -1152 5374 -1124
rect 5616 -1152 5634 -1124
rect 5664 -1152 5683 -1124
rect 5888 -1152 5906 -1124
rect 5936 -1152 5954 -1124
rect 6196 -1152 6214 -1124
rect 6244 -1152 6263 -1124
rect 6468 -1152 6486 -1124
rect 6516 -1152 6534 -1124
rect 6776 -1152 6794 -1124
rect 6824 -1152 6843 -1124
rect 14 -1298 42 -1256
rect 72 -1270 97 -1256
rect 196 -1266 221 -1256
rect 72 -1298 128 -1270
rect 158 -1298 192 -1270
tri 206 -1273 213 -1266 ne
rect 213 -1298 221 -1266
rect 251 -1298 299 -1256
rect 329 -1266 354 -1256
rect 329 -1298 337 -1266
rect 453 -1270 478 -1256
rect 358 -1298 392 -1270
rect 422 -1298 478 -1270
rect 508 -1298 536 -1256
rect 594 -1298 622 -1256
rect 652 -1270 677 -1256
rect 776 -1266 801 -1256
rect 652 -1298 708 -1270
rect 738 -1298 772 -1270
tri 786 -1273 793 -1266 ne
rect 793 -1298 801 -1266
rect 831 -1298 879 -1256
rect 909 -1266 934 -1256
rect 909 -1298 917 -1266
rect 1033 -1270 1058 -1256
rect 938 -1298 972 -1270
rect 1002 -1298 1058 -1270
rect 1088 -1298 1116 -1256
rect 1174 -1298 1202 -1256
rect 1232 -1270 1257 -1256
rect 1356 -1266 1381 -1256
rect 1232 -1298 1288 -1270
rect 1318 -1298 1352 -1270
tri 1366 -1273 1373 -1266 ne
rect 1373 -1298 1381 -1266
rect 1411 -1298 1459 -1256
rect 1489 -1266 1514 -1256
rect 1489 -1298 1497 -1266
rect 1613 -1270 1638 -1256
rect 1518 -1298 1552 -1270
rect 1582 -1298 1638 -1270
rect 1668 -1298 1696 -1256
rect 1754 -1298 1782 -1256
rect 1812 -1270 1837 -1256
rect 1936 -1266 1961 -1256
rect 1812 -1298 1868 -1270
rect 1898 -1298 1932 -1270
tri 1946 -1273 1953 -1266 ne
rect 1953 -1298 1961 -1266
rect 1991 -1298 2039 -1256
rect 2069 -1266 2094 -1256
rect 2069 -1298 2077 -1266
rect 2193 -1270 2218 -1256
rect 2098 -1298 2132 -1270
rect 2162 -1298 2218 -1270
rect 2248 -1298 2276 -1256
rect 2334 -1298 2362 -1256
rect 2392 -1270 2417 -1256
rect 2516 -1266 2541 -1256
rect 2392 -1298 2448 -1270
rect 2478 -1298 2512 -1270
tri 2526 -1273 2533 -1266 ne
rect 2533 -1298 2541 -1266
rect 2571 -1298 2619 -1256
rect 2649 -1266 2674 -1256
rect 2649 -1298 2657 -1266
rect 2773 -1270 2798 -1256
rect 2678 -1298 2712 -1270
rect 2742 -1298 2798 -1270
rect 2828 -1298 2856 -1256
rect 2914 -1298 2942 -1256
rect 2972 -1270 2997 -1256
rect 3096 -1266 3121 -1256
rect 2972 -1298 3028 -1270
rect 3058 -1298 3092 -1270
tri 3106 -1273 3113 -1266 ne
rect 3113 -1298 3121 -1266
rect 3151 -1298 3199 -1256
rect 3229 -1266 3254 -1256
rect 3229 -1298 3237 -1266
rect 3353 -1270 3378 -1256
rect 3258 -1298 3292 -1270
rect 3322 -1298 3378 -1270
rect 3408 -1298 3436 -1256
rect 3494 -1298 3522 -1256
rect 3552 -1270 3577 -1256
rect 3676 -1266 3701 -1256
rect 3552 -1298 3608 -1270
rect 3638 -1298 3672 -1270
tri 3686 -1273 3693 -1266 ne
rect 3693 -1298 3701 -1266
rect 3731 -1298 3779 -1256
rect 3809 -1266 3834 -1256
rect 3809 -1298 3817 -1266
rect 3933 -1270 3958 -1256
rect 3838 -1298 3872 -1270
rect 3902 -1298 3958 -1270
rect 3988 -1298 4016 -1256
rect 4074 -1298 4102 -1256
rect 4132 -1270 4157 -1256
rect 4256 -1266 4281 -1256
rect 4132 -1298 4188 -1270
rect 4218 -1298 4252 -1270
tri 4266 -1273 4273 -1266 ne
rect 4273 -1298 4281 -1266
rect 4311 -1298 4359 -1256
rect 4389 -1266 4414 -1256
rect 4389 -1298 4397 -1266
rect 4513 -1270 4538 -1256
rect 4418 -1298 4452 -1270
rect 4482 -1298 4538 -1270
rect 4568 -1298 4596 -1256
rect 4654 -1298 4682 -1256
rect 4712 -1270 4737 -1256
rect 4836 -1266 4861 -1256
rect 4712 -1298 4768 -1270
rect 4798 -1298 4832 -1270
tri 4846 -1273 4853 -1266 ne
rect 4853 -1298 4861 -1266
rect 4891 -1298 4939 -1256
rect 4969 -1266 4994 -1256
rect 4969 -1298 4977 -1266
rect 5093 -1270 5118 -1256
rect 4998 -1298 5032 -1270
rect 5062 -1298 5118 -1270
rect 5148 -1298 5176 -1256
rect 5234 -1298 5262 -1256
rect 5292 -1270 5317 -1256
rect 5416 -1266 5441 -1256
rect 5292 -1298 5348 -1270
rect 5378 -1298 5412 -1270
tri 5426 -1273 5433 -1266 ne
rect 5433 -1298 5441 -1266
rect 5471 -1298 5519 -1256
rect 5549 -1266 5574 -1256
rect 5549 -1298 5557 -1266
rect 5673 -1270 5698 -1256
rect 5578 -1298 5612 -1270
rect 5642 -1298 5698 -1270
rect 5728 -1298 5756 -1256
rect 5814 -1298 5842 -1256
rect 5872 -1270 5897 -1256
rect 5996 -1266 6021 -1256
rect 5872 -1298 5928 -1270
rect 5958 -1298 5992 -1270
tri 6006 -1273 6013 -1266 ne
rect 6013 -1298 6021 -1266
rect 6051 -1298 6099 -1256
rect 6129 -1266 6154 -1256
rect 6129 -1298 6137 -1266
rect 6253 -1270 6278 -1256
rect 6158 -1298 6192 -1270
rect 6222 -1298 6278 -1270
rect 6308 -1298 6336 -1256
rect 6394 -1298 6422 -1256
rect 6452 -1270 6477 -1256
rect 6576 -1266 6601 -1256
rect 6452 -1298 6508 -1270
rect 6538 -1298 6572 -1270
tri 6586 -1273 6593 -1266 ne
rect 6593 -1298 6601 -1266
rect 6631 -1298 6679 -1256
rect 6709 -1266 6734 -1256
rect 6709 -1298 6717 -1266
rect 6833 -1270 6858 -1256
rect 6738 -1298 6772 -1270
rect 6802 -1298 6858 -1270
rect 6888 -1298 6916 -1256
rect 165 -1322 192 -1298
rect 259 -1320 291 -1298
rect 259 -1322 261 -1320
rect 289 -1322 291 -1320
rect 358 -1322 385 -1298
rect 165 -1336 259 -1322
rect 291 -1336 385 -1322
rect 745 -1322 772 -1298
rect 839 -1320 871 -1298
rect 839 -1322 841 -1320
rect 869 -1322 871 -1320
rect 938 -1322 965 -1298
rect 745 -1336 839 -1322
rect 871 -1336 965 -1322
rect 1325 -1322 1352 -1298
rect 1419 -1320 1451 -1298
rect 1419 -1322 1421 -1320
rect 1449 -1322 1451 -1320
rect 1518 -1322 1545 -1298
rect 1325 -1336 1419 -1322
rect 1451 -1336 1545 -1322
rect 1905 -1322 1932 -1298
rect 1999 -1320 2031 -1298
rect 1999 -1322 2001 -1320
rect 2029 -1322 2031 -1320
rect 2098 -1322 2125 -1298
rect 1905 -1336 1999 -1322
rect 2031 -1336 2125 -1322
rect 2485 -1322 2512 -1298
rect 2579 -1320 2611 -1298
rect 2579 -1322 2581 -1320
rect 2609 -1322 2611 -1320
rect 2678 -1322 2705 -1298
rect 2485 -1336 2579 -1322
rect 2611 -1336 2705 -1322
rect 3065 -1322 3092 -1298
rect 3159 -1320 3191 -1298
rect 3159 -1322 3161 -1320
rect 3189 -1322 3191 -1320
rect 3258 -1322 3285 -1298
rect 3065 -1336 3159 -1322
rect 3191 -1336 3285 -1322
rect 3645 -1322 3672 -1298
rect 3739 -1320 3771 -1298
rect 3739 -1322 3741 -1320
rect 3769 -1322 3771 -1320
rect 3838 -1322 3865 -1298
rect 3645 -1336 3739 -1322
rect 3771 -1336 3865 -1322
rect 4225 -1322 4252 -1298
rect 4319 -1320 4351 -1298
rect 4319 -1322 4321 -1320
rect 4349 -1322 4351 -1320
rect 4418 -1322 4445 -1298
rect 4225 -1336 4319 -1322
rect 4351 -1336 4445 -1322
rect 4805 -1322 4832 -1298
rect 4899 -1320 4931 -1298
rect 4899 -1322 4901 -1320
rect 4929 -1322 4931 -1320
rect 4998 -1322 5025 -1298
rect 4805 -1336 4899 -1322
rect 4931 -1336 5025 -1322
rect 5385 -1322 5412 -1298
rect 5479 -1320 5511 -1298
rect 5479 -1322 5481 -1320
rect 5509 -1322 5511 -1320
rect 5578 -1322 5605 -1298
rect 5385 -1336 5479 -1322
rect 5511 -1336 5605 -1322
rect 5965 -1322 5992 -1298
rect 6059 -1320 6091 -1298
rect 6059 -1322 6061 -1320
rect 6089 -1322 6091 -1320
rect 6158 -1322 6185 -1298
rect 5965 -1336 6059 -1322
rect 6091 -1336 6185 -1322
rect 6545 -1322 6572 -1298
rect 6639 -1320 6671 -1298
rect 6639 -1322 6641 -1320
rect 6669 -1322 6671 -1320
rect 6738 -1322 6765 -1298
rect 6545 -1336 6639 -1322
rect 6671 -1336 6765 -1322
rect 88 -1422 106 -1394
rect 136 -1422 154 -1394
rect 396 -1422 414 -1394
rect 444 -1422 463 -1394
rect 668 -1422 686 -1394
rect 716 -1422 734 -1394
rect 976 -1422 994 -1394
rect 1024 -1422 1043 -1394
rect 1248 -1422 1266 -1394
rect 1296 -1422 1314 -1394
rect 1556 -1422 1574 -1394
rect 1604 -1422 1623 -1394
rect 1828 -1422 1846 -1394
rect 1876 -1422 1894 -1394
rect 2136 -1422 2154 -1394
rect 2184 -1422 2203 -1394
rect 2408 -1422 2426 -1394
rect 2456 -1422 2474 -1394
rect 2716 -1422 2734 -1394
rect 2764 -1422 2783 -1394
rect 2988 -1422 3006 -1394
rect 3036 -1422 3054 -1394
rect 3296 -1422 3314 -1394
rect 3344 -1422 3363 -1394
rect 3568 -1422 3586 -1394
rect 3616 -1422 3634 -1394
rect 3876 -1422 3894 -1394
rect 3924 -1422 3943 -1394
rect 4148 -1422 4166 -1394
rect 4196 -1422 4214 -1394
rect 4456 -1422 4474 -1394
rect 4504 -1422 4523 -1394
rect 4728 -1422 4746 -1394
rect 4776 -1422 4794 -1394
rect 5036 -1422 5054 -1394
rect 5084 -1422 5103 -1394
rect 5308 -1422 5326 -1394
rect 5356 -1422 5374 -1394
rect 5616 -1422 5634 -1394
rect 5664 -1422 5683 -1394
rect 5888 -1422 5906 -1394
rect 5936 -1422 5954 -1394
rect 6196 -1422 6214 -1394
rect 6244 -1422 6263 -1394
rect 6468 -1422 6486 -1394
rect 6516 -1422 6534 -1394
rect 6776 -1422 6794 -1394
rect 6824 -1422 6843 -1394
rect 14 -1568 42 -1526
rect 72 -1540 97 -1526
rect 196 -1536 221 -1526
rect 72 -1568 128 -1540
rect 158 -1568 192 -1540
tri 206 -1543 213 -1536 ne
rect 213 -1568 221 -1536
rect 251 -1568 299 -1526
rect 329 -1536 354 -1526
rect 329 -1568 337 -1536
rect 453 -1540 478 -1526
rect 358 -1568 392 -1540
rect 422 -1568 478 -1540
rect 508 -1568 536 -1526
rect 594 -1568 622 -1526
rect 652 -1540 677 -1526
rect 776 -1536 801 -1526
rect 652 -1568 708 -1540
rect 738 -1568 772 -1540
tri 786 -1543 793 -1536 ne
rect 793 -1568 801 -1536
rect 831 -1568 879 -1526
rect 909 -1536 934 -1526
rect 909 -1568 917 -1536
rect 1033 -1540 1058 -1526
rect 938 -1568 972 -1540
rect 1002 -1568 1058 -1540
rect 1088 -1568 1116 -1526
rect 1174 -1568 1202 -1526
rect 1232 -1540 1257 -1526
rect 1356 -1536 1381 -1526
rect 1232 -1568 1288 -1540
rect 1318 -1568 1352 -1540
tri 1366 -1543 1373 -1536 ne
rect 1373 -1568 1381 -1536
rect 1411 -1568 1459 -1526
rect 1489 -1536 1514 -1526
rect 1489 -1568 1497 -1536
rect 1613 -1540 1638 -1526
rect 1518 -1568 1552 -1540
rect 1582 -1568 1638 -1540
rect 1668 -1568 1696 -1526
rect 1754 -1568 1782 -1526
rect 1812 -1540 1837 -1526
rect 1936 -1536 1961 -1526
rect 1812 -1568 1868 -1540
rect 1898 -1568 1932 -1540
tri 1946 -1543 1953 -1536 ne
rect 1953 -1568 1961 -1536
rect 1991 -1568 2039 -1526
rect 2069 -1536 2094 -1526
rect 2069 -1568 2077 -1536
rect 2193 -1540 2218 -1526
rect 2098 -1568 2132 -1540
rect 2162 -1568 2218 -1540
rect 2248 -1568 2276 -1526
rect 2334 -1568 2362 -1526
rect 2392 -1540 2417 -1526
rect 2516 -1536 2541 -1526
rect 2392 -1568 2448 -1540
rect 2478 -1568 2512 -1540
tri 2526 -1543 2533 -1536 ne
rect 2533 -1568 2541 -1536
rect 2571 -1568 2619 -1526
rect 2649 -1536 2674 -1526
rect 2649 -1568 2657 -1536
rect 2773 -1540 2798 -1526
rect 2678 -1568 2712 -1540
rect 2742 -1568 2798 -1540
rect 2828 -1568 2856 -1526
rect 2914 -1568 2942 -1526
rect 2972 -1540 2997 -1526
rect 3096 -1536 3121 -1526
rect 2972 -1568 3028 -1540
rect 3058 -1568 3092 -1540
tri 3106 -1543 3113 -1536 ne
rect 3113 -1568 3121 -1536
rect 3151 -1568 3199 -1526
rect 3229 -1536 3254 -1526
rect 3229 -1568 3237 -1536
rect 3353 -1540 3378 -1526
rect 3258 -1568 3292 -1540
rect 3322 -1568 3378 -1540
rect 3408 -1568 3436 -1526
rect 3494 -1568 3522 -1526
rect 3552 -1540 3577 -1526
rect 3676 -1536 3701 -1526
rect 3552 -1568 3608 -1540
rect 3638 -1568 3672 -1540
tri 3686 -1543 3693 -1536 ne
rect 3693 -1568 3701 -1536
rect 3731 -1568 3779 -1526
rect 3809 -1536 3834 -1526
rect 3809 -1568 3817 -1536
rect 3933 -1540 3958 -1526
rect 3838 -1568 3872 -1540
rect 3902 -1568 3958 -1540
rect 3988 -1568 4016 -1526
rect 4074 -1568 4102 -1526
rect 4132 -1540 4157 -1526
rect 4256 -1536 4281 -1526
rect 4132 -1568 4188 -1540
rect 4218 -1568 4252 -1540
tri 4266 -1543 4273 -1536 ne
rect 4273 -1568 4281 -1536
rect 4311 -1568 4359 -1526
rect 4389 -1536 4414 -1526
rect 4389 -1568 4397 -1536
rect 4513 -1540 4538 -1526
rect 4418 -1568 4452 -1540
rect 4482 -1568 4538 -1540
rect 4568 -1568 4596 -1526
rect 4654 -1568 4682 -1526
rect 4712 -1540 4737 -1526
rect 4836 -1536 4861 -1526
rect 4712 -1568 4768 -1540
rect 4798 -1568 4832 -1540
tri 4846 -1543 4853 -1536 ne
rect 4853 -1568 4861 -1536
rect 4891 -1568 4939 -1526
rect 4969 -1536 4994 -1526
rect 4969 -1568 4977 -1536
rect 5093 -1540 5118 -1526
rect 4998 -1568 5032 -1540
rect 5062 -1568 5118 -1540
rect 5148 -1568 5176 -1526
rect 5234 -1568 5262 -1526
rect 5292 -1540 5317 -1526
rect 5416 -1536 5441 -1526
rect 5292 -1568 5348 -1540
rect 5378 -1568 5412 -1540
tri 5426 -1543 5433 -1536 ne
rect 5433 -1568 5441 -1536
rect 5471 -1568 5519 -1526
rect 5549 -1536 5574 -1526
rect 5549 -1568 5557 -1536
rect 5673 -1540 5698 -1526
rect 5578 -1568 5612 -1540
rect 5642 -1568 5698 -1540
rect 5728 -1568 5756 -1526
rect 5814 -1568 5842 -1526
rect 5872 -1540 5897 -1526
rect 5996 -1536 6021 -1526
rect 5872 -1568 5928 -1540
rect 5958 -1568 5992 -1540
tri 6006 -1543 6013 -1536 ne
rect 6013 -1568 6021 -1536
rect 6051 -1568 6099 -1526
rect 6129 -1536 6154 -1526
rect 6129 -1568 6137 -1536
rect 6253 -1540 6278 -1526
rect 6158 -1568 6192 -1540
rect 6222 -1568 6278 -1540
rect 6308 -1568 6336 -1526
rect 6394 -1568 6422 -1526
rect 6452 -1540 6477 -1526
rect 6576 -1536 6601 -1526
rect 6452 -1568 6508 -1540
rect 6538 -1568 6572 -1540
tri 6586 -1543 6593 -1536 ne
rect 6593 -1568 6601 -1536
rect 6631 -1568 6679 -1526
rect 6709 -1536 6734 -1526
rect 6709 -1568 6717 -1536
rect 6833 -1540 6858 -1526
rect 6738 -1568 6772 -1540
rect 6802 -1568 6858 -1540
rect 6888 -1568 6916 -1526
rect 165 -1592 192 -1568
rect 259 -1590 291 -1568
rect 259 -1592 261 -1590
rect 289 -1592 291 -1590
rect 358 -1592 385 -1568
rect 165 -1606 259 -1592
rect 291 -1606 385 -1592
rect 745 -1592 772 -1568
rect 839 -1590 871 -1568
rect 839 -1592 841 -1590
rect 869 -1592 871 -1590
rect 938 -1592 965 -1568
rect 745 -1606 839 -1592
rect 871 -1606 965 -1592
rect 1325 -1592 1352 -1568
rect 1419 -1590 1451 -1568
rect 1419 -1592 1421 -1590
rect 1449 -1592 1451 -1590
rect 1518 -1592 1545 -1568
rect 1325 -1606 1419 -1592
rect 1451 -1606 1545 -1592
rect 1905 -1592 1932 -1568
rect 1999 -1590 2031 -1568
rect 1999 -1592 2001 -1590
rect 2029 -1592 2031 -1590
rect 2098 -1592 2125 -1568
rect 1905 -1606 1999 -1592
rect 2031 -1606 2125 -1592
rect 2485 -1592 2512 -1568
rect 2579 -1590 2611 -1568
rect 2579 -1592 2581 -1590
rect 2609 -1592 2611 -1590
rect 2678 -1592 2705 -1568
rect 2485 -1606 2579 -1592
rect 2611 -1606 2705 -1592
rect 3065 -1592 3092 -1568
rect 3159 -1590 3191 -1568
rect 3159 -1592 3161 -1590
rect 3189 -1592 3191 -1590
rect 3258 -1592 3285 -1568
rect 3065 -1606 3159 -1592
rect 3191 -1606 3285 -1592
rect 3645 -1592 3672 -1568
rect 3739 -1590 3771 -1568
rect 3739 -1592 3741 -1590
rect 3769 -1592 3771 -1590
rect 3838 -1592 3865 -1568
rect 3645 -1606 3739 -1592
rect 3771 -1606 3865 -1592
rect 4225 -1592 4252 -1568
rect 4319 -1590 4351 -1568
rect 4319 -1592 4321 -1590
rect 4349 -1592 4351 -1590
rect 4418 -1592 4445 -1568
rect 4225 -1606 4319 -1592
rect 4351 -1606 4445 -1592
rect 4805 -1592 4832 -1568
rect 4899 -1590 4931 -1568
rect 4899 -1592 4901 -1590
rect 4929 -1592 4931 -1590
rect 4998 -1592 5025 -1568
rect 4805 -1606 4899 -1592
rect 4931 -1606 5025 -1592
rect 5385 -1592 5412 -1568
rect 5479 -1590 5511 -1568
rect 5479 -1592 5481 -1590
rect 5509 -1592 5511 -1590
rect 5578 -1592 5605 -1568
rect 5385 -1606 5479 -1592
rect 5511 -1606 5605 -1592
rect 5965 -1592 5992 -1568
rect 6059 -1590 6091 -1568
rect 6059 -1592 6061 -1590
rect 6089 -1592 6091 -1590
rect 6158 -1592 6185 -1568
rect 5965 -1606 6059 -1592
rect 6091 -1606 6185 -1592
rect 6545 -1592 6572 -1568
rect 6639 -1590 6671 -1568
rect 6639 -1592 6641 -1590
rect 6669 -1592 6671 -1590
rect 6738 -1592 6765 -1568
rect 6545 -1606 6639 -1592
rect 6671 -1606 6765 -1592
rect 88 -1692 106 -1664
rect 136 -1692 154 -1664
rect 396 -1692 414 -1664
rect 444 -1692 463 -1664
rect 668 -1692 686 -1664
rect 716 -1692 734 -1664
rect 976 -1692 994 -1664
rect 1024 -1692 1043 -1664
rect 1248 -1692 1266 -1664
rect 1296 -1692 1314 -1664
rect 1556 -1692 1574 -1664
rect 1604 -1692 1623 -1664
rect 1828 -1692 1846 -1664
rect 1876 -1692 1894 -1664
rect 2136 -1692 2154 -1664
rect 2184 -1692 2203 -1664
rect 2408 -1692 2426 -1664
rect 2456 -1692 2474 -1664
rect 2716 -1692 2734 -1664
rect 2764 -1692 2783 -1664
rect 2988 -1692 3006 -1664
rect 3036 -1692 3054 -1664
rect 3296 -1692 3314 -1664
rect 3344 -1692 3363 -1664
rect 3568 -1692 3586 -1664
rect 3616 -1692 3634 -1664
rect 3876 -1692 3894 -1664
rect 3924 -1692 3943 -1664
rect 4148 -1692 4166 -1664
rect 4196 -1692 4214 -1664
rect 4456 -1692 4474 -1664
rect 4504 -1692 4523 -1664
rect 4728 -1692 4746 -1664
rect 4776 -1692 4794 -1664
rect 5036 -1692 5054 -1664
rect 5084 -1692 5103 -1664
rect 5308 -1692 5326 -1664
rect 5356 -1692 5374 -1664
rect 5616 -1692 5634 -1664
rect 5664 -1692 5683 -1664
rect 5888 -1692 5906 -1664
rect 5936 -1692 5954 -1664
rect 6196 -1692 6214 -1664
rect 6244 -1692 6263 -1664
rect 6468 -1692 6486 -1664
rect 6516 -1692 6534 -1664
rect 6776 -1692 6794 -1664
rect 6824 -1692 6843 -1664
rect 14 -1838 42 -1796
rect 72 -1810 97 -1796
rect 196 -1806 221 -1796
rect 72 -1838 128 -1810
rect 158 -1838 192 -1810
tri 206 -1813 213 -1806 ne
rect 213 -1838 221 -1806
rect 251 -1838 299 -1796
rect 329 -1806 354 -1796
rect 329 -1838 337 -1806
rect 453 -1810 478 -1796
rect 358 -1838 392 -1810
rect 422 -1838 478 -1810
rect 508 -1838 536 -1796
rect 594 -1838 622 -1796
rect 652 -1810 677 -1796
rect 776 -1806 801 -1796
rect 652 -1838 708 -1810
rect 738 -1838 772 -1810
tri 786 -1813 793 -1806 ne
rect 793 -1838 801 -1806
rect 831 -1838 879 -1796
rect 909 -1806 934 -1796
rect 909 -1838 917 -1806
rect 1033 -1810 1058 -1796
rect 938 -1838 972 -1810
rect 1002 -1838 1058 -1810
rect 1088 -1838 1116 -1796
rect 1174 -1838 1202 -1796
rect 1232 -1810 1257 -1796
rect 1356 -1806 1381 -1796
rect 1232 -1838 1288 -1810
rect 1318 -1838 1352 -1810
tri 1366 -1813 1373 -1806 ne
rect 1373 -1838 1381 -1806
rect 1411 -1838 1459 -1796
rect 1489 -1806 1514 -1796
rect 1489 -1838 1497 -1806
rect 1613 -1810 1638 -1796
rect 1518 -1838 1552 -1810
rect 1582 -1838 1638 -1810
rect 1668 -1838 1696 -1796
rect 1754 -1838 1782 -1796
rect 1812 -1810 1837 -1796
rect 1936 -1806 1961 -1796
rect 1812 -1838 1868 -1810
rect 1898 -1838 1932 -1810
tri 1946 -1813 1953 -1806 ne
rect 1953 -1838 1961 -1806
rect 1991 -1838 2039 -1796
rect 2069 -1806 2094 -1796
rect 2069 -1838 2077 -1806
rect 2193 -1810 2218 -1796
rect 2098 -1838 2132 -1810
rect 2162 -1838 2218 -1810
rect 2248 -1838 2276 -1796
rect 2334 -1838 2362 -1796
rect 2392 -1810 2417 -1796
rect 2516 -1806 2541 -1796
rect 2392 -1838 2448 -1810
rect 2478 -1838 2512 -1810
tri 2526 -1813 2533 -1806 ne
rect 2533 -1838 2541 -1806
rect 2571 -1838 2619 -1796
rect 2649 -1806 2674 -1796
rect 2649 -1838 2657 -1806
rect 2773 -1810 2798 -1796
rect 2678 -1838 2712 -1810
rect 2742 -1838 2798 -1810
rect 2828 -1838 2856 -1796
rect 2914 -1838 2942 -1796
rect 2972 -1810 2997 -1796
rect 3096 -1806 3121 -1796
rect 2972 -1838 3028 -1810
rect 3058 -1838 3092 -1810
tri 3106 -1813 3113 -1806 ne
rect 3113 -1838 3121 -1806
rect 3151 -1838 3199 -1796
rect 3229 -1806 3254 -1796
rect 3229 -1838 3237 -1806
rect 3353 -1810 3378 -1796
rect 3258 -1838 3292 -1810
rect 3322 -1838 3378 -1810
rect 3408 -1838 3436 -1796
rect 3494 -1838 3522 -1796
rect 3552 -1810 3577 -1796
rect 3676 -1806 3701 -1796
rect 3552 -1838 3608 -1810
rect 3638 -1838 3672 -1810
tri 3686 -1813 3693 -1806 ne
rect 3693 -1838 3701 -1806
rect 3731 -1838 3779 -1796
rect 3809 -1806 3834 -1796
rect 3809 -1838 3817 -1806
rect 3933 -1810 3958 -1796
rect 3838 -1838 3872 -1810
rect 3902 -1838 3958 -1810
rect 3988 -1838 4016 -1796
rect 4074 -1838 4102 -1796
rect 4132 -1810 4157 -1796
rect 4256 -1806 4281 -1796
rect 4132 -1838 4188 -1810
rect 4218 -1838 4252 -1810
tri 4266 -1813 4273 -1806 ne
rect 4273 -1838 4281 -1806
rect 4311 -1838 4359 -1796
rect 4389 -1806 4414 -1796
rect 4389 -1838 4397 -1806
rect 4513 -1810 4538 -1796
rect 4418 -1838 4452 -1810
rect 4482 -1838 4538 -1810
rect 4568 -1838 4596 -1796
rect 4654 -1838 4682 -1796
rect 4712 -1810 4737 -1796
rect 4836 -1806 4861 -1796
rect 4712 -1838 4768 -1810
rect 4798 -1838 4832 -1810
tri 4846 -1813 4853 -1806 ne
rect 4853 -1838 4861 -1806
rect 4891 -1838 4939 -1796
rect 4969 -1806 4994 -1796
rect 4969 -1838 4977 -1806
rect 5093 -1810 5118 -1796
rect 4998 -1838 5032 -1810
rect 5062 -1838 5118 -1810
rect 5148 -1838 5176 -1796
rect 5234 -1838 5262 -1796
rect 5292 -1810 5317 -1796
rect 5416 -1806 5441 -1796
rect 5292 -1838 5348 -1810
rect 5378 -1838 5412 -1810
tri 5426 -1813 5433 -1806 ne
rect 5433 -1838 5441 -1806
rect 5471 -1838 5519 -1796
rect 5549 -1806 5574 -1796
rect 5549 -1838 5557 -1806
rect 5673 -1810 5698 -1796
rect 5578 -1838 5612 -1810
rect 5642 -1838 5698 -1810
rect 5728 -1838 5756 -1796
rect 5814 -1838 5842 -1796
rect 5872 -1810 5897 -1796
rect 5996 -1806 6021 -1796
rect 5872 -1838 5928 -1810
rect 5958 -1838 5992 -1810
tri 6006 -1813 6013 -1806 ne
rect 6013 -1838 6021 -1806
rect 6051 -1838 6099 -1796
rect 6129 -1806 6154 -1796
rect 6129 -1838 6137 -1806
rect 6253 -1810 6278 -1796
rect 6158 -1838 6192 -1810
rect 6222 -1838 6278 -1810
rect 6308 -1838 6336 -1796
rect 6394 -1838 6422 -1796
rect 6452 -1810 6477 -1796
rect 6576 -1806 6601 -1796
rect 6452 -1838 6508 -1810
rect 6538 -1838 6572 -1810
tri 6586 -1813 6593 -1806 ne
rect 6593 -1838 6601 -1806
rect 6631 -1838 6679 -1796
rect 6709 -1806 6734 -1796
rect 6709 -1838 6717 -1806
rect 6833 -1810 6858 -1796
rect 6738 -1838 6772 -1810
rect 6802 -1838 6858 -1810
rect 6888 -1838 6916 -1796
rect 165 -1862 192 -1838
rect 259 -1860 291 -1838
rect 259 -1862 261 -1860
rect 289 -1862 291 -1860
rect 358 -1862 385 -1838
rect 165 -1876 259 -1862
rect 291 -1876 385 -1862
rect 745 -1862 772 -1838
rect 839 -1860 871 -1838
rect 839 -1862 841 -1860
rect 869 -1862 871 -1860
rect 938 -1862 965 -1838
rect 745 -1876 839 -1862
rect 871 -1876 965 -1862
rect 1325 -1862 1352 -1838
rect 1419 -1860 1451 -1838
rect 1419 -1862 1421 -1860
rect 1449 -1862 1451 -1860
rect 1518 -1862 1545 -1838
rect 1325 -1876 1419 -1862
rect 1451 -1876 1545 -1862
rect 1905 -1862 1932 -1838
rect 1999 -1860 2031 -1838
rect 1999 -1862 2001 -1860
rect 2029 -1862 2031 -1860
rect 2098 -1862 2125 -1838
rect 1905 -1876 1999 -1862
rect 2031 -1876 2125 -1862
rect 2485 -1862 2512 -1838
rect 2579 -1860 2611 -1838
rect 2579 -1862 2581 -1860
rect 2609 -1862 2611 -1860
rect 2678 -1862 2705 -1838
rect 2485 -1876 2579 -1862
rect 2611 -1876 2705 -1862
rect 3065 -1862 3092 -1838
rect 3159 -1860 3191 -1838
rect 3159 -1862 3161 -1860
rect 3189 -1862 3191 -1860
rect 3258 -1862 3285 -1838
rect 3065 -1876 3159 -1862
rect 3191 -1876 3285 -1862
rect 3645 -1862 3672 -1838
rect 3739 -1860 3771 -1838
rect 3739 -1862 3741 -1860
rect 3769 -1862 3771 -1860
rect 3838 -1862 3865 -1838
rect 3645 -1876 3739 -1862
rect 3771 -1876 3865 -1862
rect 4225 -1862 4252 -1838
rect 4319 -1860 4351 -1838
rect 4319 -1862 4321 -1860
rect 4349 -1862 4351 -1860
rect 4418 -1862 4445 -1838
rect 4225 -1876 4319 -1862
rect 4351 -1876 4445 -1862
rect 4805 -1862 4832 -1838
rect 4899 -1860 4931 -1838
rect 4899 -1862 4901 -1860
rect 4929 -1862 4931 -1860
rect 4998 -1862 5025 -1838
rect 4805 -1876 4899 -1862
rect 4931 -1876 5025 -1862
rect 5385 -1862 5412 -1838
rect 5479 -1860 5511 -1838
rect 5479 -1862 5481 -1860
rect 5509 -1862 5511 -1860
rect 5578 -1862 5605 -1838
rect 5385 -1876 5479 -1862
rect 5511 -1876 5605 -1862
rect 5965 -1862 5992 -1838
rect 6059 -1860 6091 -1838
rect 6059 -1862 6061 -1860
rect 6089 -1862 6091 -1860
rect 6158 -1862 6185 -1838
rect 5965 -1876 6059 -1862
rect 6091 -1876 6185 -1862
rect 6545 -1862 6572 -1838
rect 6639 -1860 6671 -1838
rect 6639 -1862 6641 -1860
rect 6669 -1862 6671 -1860
rect 6738 -1862 6765 -1838
rect 6545 -1876 6639 -1862
rect 6671 -1876 6765 -1862
rect 88 -1962 106 -1934
rect 136 -1962 154 -1934
rect 396 -1962 414 -1934
rect 444 -1962 463 -1934
rect 668 -1962 686 -1934
rect 716 -1962 734 -1934
rect 976 -1962 994 -1934
rect 1024 -1962 1043 -1934
rect 1248 -1962 1266 -1934
rect 1296 -1962 1314 -1934
rect 1556 -1962 1574 -1934
rect 1604 -1962 1623 -1934
rect 1828 -1962 1846 -1934
rect 1876 -1962 1894 -1934
rect 2136 -1962 2154 -1934
rect 2184 -1962 2203 -1934
rect 2408 -1962 2426 -1934
rect 2456 -1962 2474 -1934
rect 2716 -1962 2734 -1934
rect 2764 -1962 2783 -1934
rect 2988 -1962 3006 -1934
rect 3036 -1962 3054 -1934
rect 3296 -1962 3314 -1934
rect 3344 -1962 3363 -1934
rect 3568 -1962 3586 -1934
rect 3616 -1962 3634 -1934
rect 3876 -1962 3894 -1934
rect 3924 -1962 3943 -1934
rect 4148 -1962 4166 -1934
rect 4196 -1962 4214 -1934
rect 4456 -1962 4474 -1934
rect 4504 -1962 4523 -1934
rect 4728 -1962 4746 -1934
rect 4776 -1962 4794 -1934
rect 5036 -1962 5054 -1934
rect 5084 -1962 5103 -1934
rect 5308 -1962 5326 -1934
rect 5356 -1962 5374 -1934
rect 5616 -1962 5634 -1934
rect 5664 -1962 5683 -1934
rect 5888 -1962 5906 -1934
rect 5936 -1962 5954 -1934
rect 6196 -1962 6214 -1934
rect 6244 -1962 6263 -1934
rect 6468 -1962 6486 -1934
rect 6516 -1962 6534 -1934
rect 6776 -1962 6794 -1934
rect 6824 -1962 6843 -1934
rect 14 -2108 42 -2066
rect 72 -2080 97 -2066
rect 196 -2076 221 -2066
rect 72 -2108 128 -2080
rect 158 -2108 192 -2080
tri 206 -2083 213 -2076 ne
rect 213 -2108 221 -2076
rect 251 -2108 299 -2066
rect 329 -2076 354 -2066
rect 329 -2108 337 -2076
rect 453 -2080 478 -2066
rect 358 -2108 392 -2080
rect 422 -2108 478 -2080
rect 508 -2108 536 -2066
rect 594 -2108 622 -2066
rect 652 -2080 677 -2066
rect 776 -2076 801 -2066
rect 652 -2108 708 -2080
rect 738 -2108 772 -2080
tri 786 -2083 793 -2076 ne
rect 793 -2108 801 -2076
rect 831 -2108 879 -2066
rect 909 -2076 934 -2066
rect 909 -2108 917 -2076
rect 1033 -2080 1058 -2066
rect 938 -2108 972 -2080
rect 1002 -2108 1058 -2080
rect 1088 -2108 1116 -2066
rect 1174 -2108 1202 -2066
rect 1232 -2080 1257 -2066
rect 1356 -2076 1381 -2066
rect 1232 -2108 1288 -2080
rect 1318 -2108 1352 -2080
tri 1366 -2083 1373 -2076 ne
rect 1373 -2108 1381 -2076
rect 1411 -2108 1459 -2066
rect 1489 -2076 1514 -2066
rect 1489 -2108 1497 -2076
rect 1613 -2080 1638 -2066
rect 1518 -2108 1552 -2080
rect 1582 -2108 1638 -2080
rect 1668 -2108 1696 -2066
rect 1754 -2108 1782 -2066
rect 1812 -2080 1837 -2066
rect 1936 -2076 1961 -2066
rect 1812 -2108 1868 -2080
rect 1898 -2108 1932 -2080
tri 1946 -2083 1953 -2076 ne
rect 1953 -2108 1961 -2076
rect 1991 -2108 2039 -2066
rect 2069 -2076 2094 -2066
rect 2069 -2108 2077 -2076
rect 2193 -2080 2218 -2066
rect 2098 -2108 2132 -2080
rect 2162 -2108 2218 -2080
rect 2248 -2108 2276 -2066
rect 2334 -2108 2362 -2066
rect 2392 -2080 2417 -2066
rect 2516 -2076 2541 -2066
rect 2392 -2108 2448 -2080
rect 2478 -2108 2512 -2080
tri 2526 -2083 2533 -2076 ne
rect 2533 -2108 2541 -2076
rect 2571 -2108 2619 -2066
rect 2649 -2076 2674 -2066
rect 2649 -2108 2657 -2076
rect 2773 -2080 2798 -2066
rect 2678 -2108 2712 -2080
rect 2742 -2108 2798 -2080
rect 2828 -2108 2856 -2066
rect 2914 -2108 2942 -2066
rect 2972 -2080 2997 -2066
rect 3096 -2076 3121 -2066
rect 2972 -2108 3028 -2080
rect 3058 -2108 3092 -2080
tri 3106 -2083 3113 -2076 ne
rect 3113 -2108 3121 -2076
rect 3151 -2108 3199 -2066
rect 3229 -2076 3254 -2066
rect 3229 -2108 3237 -2076
rect 3353 -2080 3378 -2066
rect 3258 -2108 3292 -2080
rect 3322 -2108 3378 -2080
rect 3408 -2108 3436 -2066
rect 3494 -2108 3522 -2066
rect 3552 -2080 3577 -2066
rect 3676 -2076 3701 -2066
rect 3552 -2108 3608 -2080
rect 3638 -2108 3672 -2080
tri 3686 -2083 3693 -2076 ne
rect 3693 -2108 3701 -2076
rect 3731 -2108 3779 -2066
rect 3809 -2076 3834 -2066
rect 3809 -2108 3817 -2076
rect 3933 -2080 3958 -2066
rect 3838 -2108 3872 -2080
rect 3902 -2108 3958 -2080
rect 3988 -2108 4016 -2066
rect 4074 -2108 4102 -2066
rect 4132 -2080 4157 -2066
rect 4256 -2076 4281 -2066
rect 4132 -2108 4188 -2080
rect 4218 -2108 4252 -2080
tri 4266 -2083 4273 -2076 ne
rect 4273 -2108 4281 -2076
rect 4311 -2108 4359 -2066
rect 4389 -2076 4414 -2066
rect 4389 -2108 4397 -2076
rect 4513 -2080 4538 -2066
rect 4418 -2108 4452 -2080
rect 4482 -2108 4538 -2080
rect 4568 -2108 4596 -2066
rect 4654 -2108 4682 -2066
rect 4712 -2080 4737 -2066
rect 4836 -2076 4861 -2066
rect 4712 -2108 4768 -2080
rect 4798 -2108 4832 -2080
tri 4846 -2083 4853 -2076 ne
rect 4853 -2108 4861 -2076
rect 4891 -2108 4939 -2066
rect 4969 -2076 4994 -2066
rect 4969 -2108 4977 -2076
rect 5093 -2080 5118 -2066
rect 4998 -2108 5032 -2080
rect 5062 -2108 5118 -2080
rect 5148 -2108 5176 -2066
rect 5234 -2108 5262 -2066
rect 5292 -2080 5317 -2066
rect 5416 -2076 5441 -2066
rect 5292 -2108 5348 -2080
rect 5378 -2108 5412 -2080
tri 5426 -2083 5433 -2076 ne
rect 5433 -2108 5441 -2076
rect 5471 -2108 5519 -2066
rect 5549 -2076 5574 -2066
rect 5549 -2108 5557 -2076
rect 5673 -2080 5698 -2066
rect 5578 -2108 5612 -2080
rect 5642 -2108 5698 -2080
rect 5728 -2108 5756 -2066
rect 5814 -2108 5842 -2066
rect 5872 -2080 5897 -2066
rect 5996 -2076 6021 -2066
rect 5872 -2108 5928 -2080
rect 5958 -2108 5992 -2080
tri 6006 -2083 6013 -2076 ne
rect 6013 -2108 6021 -2076
rect 6051 -2108 6099 -2066
rect 6129 -2076 6154 -2066
rect 6129 -2108 6137 -2076
rect 6253 -2080 6278 -2066
rect 6158 -2108 6192 -2080
rect 6222 -2108 6278 -2080
rect 6308 -2108 6336 -2066
rect 6394 -2108 6422 -2066
rect 6452 -2080 6477 -2066
rect 6576 -2076 6601 -2066
rect 6452 -2108 6508 -2080
rect 6538 -2108 6572 -2080
tri 6586 -2083 6593 -2076 ne
rect 6593 -2108 6601 -2076
rect 6631 -2108 6679 -2066
rect 6709 -2076 6734 -2066
rect 6709 -2108 6717 -2076
rect 6833 -2080 6858 -2066
rect 6738 -2108 6772 -2080
rect 6802 -2108 6858 -2080
rect 6888 -2108 6916 -2066
rect 165 -2132 192 -2108
rect 259 -2130 291 -2108
rect 259 -2132 261 -2130
rect 289 -2132 291 -2130
rect 358 -2132 385 -2108
rect 165 -2146 259 -2132
rect 291 -2146 385 -2132
rect 745 -2132 772 -2108
rect 839 -2130 871 -2108
rect 839 -2132 841 -2130
rect 869 -2132 871 -2130
rect 938 -2132 965 -2108
rect 745 -2146 839 -2132
rect 871 -2146 965 -2132
rect 1325 -2132 1352 -2108
rect 1419 -2130 1451 -2108
rect 1419 -2132 1421 -2130
rect 1449 -2132 1451 -2130
rect 1518 -2132 1545 -2108
rect 1325 -2146 1419 -2132
rect 1451 -2146 1545 -2132
rect 1905 -2132 1932 -2108
rect 1999 -2130 2031 -2108
rect 1999 -2132 2001 -2130
rect 2029 -2132 2031 -2130
rect 2098 -2132 2125 -2108
rect 1905 -2146 1999 -2132
rect 2031 -2146 2125 -2132
rect 2485 -2132 2512 -2108
rect 2579 -2130 2611 -2108
rect 2579 -2132 2581 -2130
rect 2609 -2132 2611 -2130
rect 2678 -2132 2705 -2108
rect 2485 -2146 2579 -2132
rect 2611 -2146 2705 -2132
rect 3065 -2132 3092 -2108
rect 3159 -2130 3191 -2108
rect 3159 -2132 3161 -2130
rect 3189 -2132 3191 -2130
rect 3258 -2132 3285 -2108
rect 3065 -2146 3159 -2132
rect 3191 -2146 3285 -2132
rect 3645 -2132 3672 -2108
rect 3739 -2130 3771 -2108
rect 3739 -2132 3741 -2130
rect 3769 -2132 3771 -2130
rect 3838 -2132 3865 -2108
rect 3645 -2146 3739 -2132
rect 3771 -2146 3865 -2132
rect 4225 -2132 4252 -2108
rect 4319 -2130 4351 -2108
rect 4319 -2132 4321 -2130
rect 4349 -2132 4351 -2130
rect 4418 -2132 4445 -2108
rect 4225 -2146 4319 -2132
rect 4351 -2146 4445 -2132
rect 4805 -2132 4832 -2108
rect 4899 -2130 4931 -2108
rect 4899 -2132 4901 -2130
rect 4929 -2132 4931 -2130
rect 4998 -2132 5025 -2108
rect 4805 -2146 4899 -2132
rect 4931 -2146 5025 -2132
rect 5385 -2132 5412 -2108
rect 5479 -2130 5511 -2108
rect 5479 -2132 5481 -2130
rect 5509 -2132 5511 -2130
rect 5578 -2132 5605 -2108
rect 5385 -2146 5479 -2132
rect 5511 -2146 5605 -2132
rect 5965 -2132 5992 -2108
rect 6059 -2130 6091 -2108
rect 6059 -2132 6061 -2130
rect 6089 -2132 6091 -2130
rect 6158 -2132 6185 -2108
rect 5965 -2146 6059 -2132
rect 6091 -2146 6185 -2132
rect 6545 -2132 6572 -2108
rect 6639 -2130 6671 -2108
rect 6639 -2132 6641 -2130
rect 6669 -2132 6671 -2130
rect 6738 -2132 6765 -2108
rect 6545 -2146 6639 -2132
rect 6671 -2146 6765 -2132
<< pdiff >>
rect 259 2128 261 2130
rect 289 2128 291 2130
rect 259 2106 291 2128
rect 212 2078 221 2106
rect 251 2078 299 2106
rect 329 2078 338 2106
tri 338 2078 350 2090 sw
rect 839 2128 841 2130
rect 869 2128 871 2130
rect 839 2106 871 2128
rect 792 2078 801 2106
rect 831 2078 879 2106
rect 909 2078 918 2106
tri 918 2078 930 2090 sw
rect 1419 2128 1421 2130
rect 1449 2128 1451 2130
rect 1419 2106 1451 2128
rect 1372 2078 1381 2106
rect 1411 2078 1459 2106
rect 1489 2078 1498 2106
tri 1498 2078 1510 2090 sw
rect 1999 2128 2001 2130
rect 2029 2128 2031 2130
rect 1999 2106 2031 2128
rect 1952 2078 1961 2106
rect 1991 2078 2039 2106
rect 2069 2078 2078 2106
tri 2078 2078 2090 2090 sw
rect 2579 2128 2581 2130
rect 2609 2128 2611 2130
rect 2579 2106 2611 2128
rect 2532 2078 2541 2106
rect 2571 2078 2619 2106
rect 2649 2078 2658 2106
tri 2658 2078 2670 2090 sw
rect 3159 2128 3161 2130
rect 3189 2128 3191 2130
rect 3159 2106 3191 2128
rect 3112 2078 3121 2106
rect 3151 2078 3199 2106
rect 3229 2078 3238 2106
tri 3238 2078 3250 2090 sw
rect 3739 2128 3741 2130
rect 3769 2128 3771 2130
rect 3739 2106 3771 2128
rect 3692 2078 3701 2106
rect 3731 2078 3779 2106
rect 3809 2078 3818 2106
tri 3818 2078 3830 2090 sw
rect 4319 2128 4321 2130
rect 4349 2128 4351 2130
rect 4319 2106 4351 2128
rect 4272 2078 4281 2106
rect 4311 2078 4359 2106
rect 4389 2078 4398 2106
tri 4398 2078 4410 2090 sw
rect 4899 2128 4901 2130
rect 4929 2128 4931 2130
rect 4899 2106 4931 2128
rect 4852 2078 4861 2106
rect 4891 2078 4939 2106
rect 4969 2078 4978 2106
tri 4978 2078 4990 2090 sw
rect 5479 2128 5481 2130
rect 5509 2128 5511 2130
rect 5479 2106 5511 2128
rect 5432 2078 5441 2106
rect 5471 2078 5519 2106
rect 5549 2078 5558 2106
tri 5558 2078 5570 2090 sw
rect 6059 2128 6061 2130
rect 6089 2128 6091 2130
rect 6059 2106 6091 2128
rect 6012 2078 6021 2106
rect 6051 2078 6099 2106
rect 6129 2078 6138 2106
tri 6138 2078 6150 2090 sw
rect 6639 2128 6641 2130
rect 6669 2128 6671 2130
rect 6639 2106 6671 2128
rect 6592 2078 6601 2106
rect 6631 2078 6679 2106
rect 6709 2078 6718 2106
tri 6718 2078 6730 2090 sw
rect 259 1858 261 1860
rect 289 1858 291 1860
rect 259 1836 291 1858
rect 212 1808 221 1836
rect 251 1808 299 1836
rect 329 1808 338 1836
tri 338 1808 350 1820 sw
rect 839 1858 841 1860
rect 869 1858 871 1860
rect 839 1836 871 1858
rect 792 1808 801 1836
rect 831 1808 879 1836
rect 909 1808 918 1836
tri 918 1808 930 1820 sw
rect 1419 1858 1421 1860
rect 1449 1858 1451 1860
rect 1419 1836 1451 1858
rect 1372 1808 1381 1836
rect 1411 1808 1459 1836
rect 1489 1808 1498 1836
tri 1498 1808 1510 1820 sw
rect 1999 1858 2001 1860
rect 2029 1858 2031 1860
rect 1999 1836 2031 1858
rect 1952 1808 1961 1836
rect 1991 1808 2039 1836
rect 2069 1808 2078 1836
tri 2078 1808 2090 1820 sw
rect 2579 1858 2581 1860
rect 2609 1858 2611 1860
rect 2579 1836 2611 1858
rect 2532 1808 2541 1836
rect 2571 1808 2619 1836
rect 2649 1808 2658 1836
tri 2658 1808 2670 1820 sw
rect 3159 1858 3161 1860
rect 3189 1858 3191 1860
rect 3159 1836 3191 1858
rect 3112 1808 3121 1836
rect 3151 1808 3199 1836
rect 3229 1808 3238 1836
tri 3238 1808 3250 1820 sw
rect 3739 1858 3741 1860
rect 3769 1858 3771 1860
rect 3739 1836 3771 1858
rect 3692 1808 3701 1836
rect 3731 1808 3779 1836
rect 3809 1808 3818 1836
tri 3818 1808 3830 1820 sw
rect 4319 1858 4321 1860
rect 4349 1858 4351 1860
rect 4319 1836 4351 1858
rect 4272 1808 4281 1836
rect 4311 1808 4359 1836
rect 4389 1808 4398 1836
tri 4398 1808 4410 1820 sw
rect 4899 1858 4901 1860
rect 4929 1858 4931 1860
rect 4899 1836 4931 1858
rect 4852 1808 4861 1836
rect 4891 1808 4939 1836
rect 4969 1808 4978 1836
tri 4978 1808 4990 1820 sw
rect 5479 1858 5481 1860
rect 5509 1858 5511 1860
rect 5479 1836 5511 1858
rect 5432 1808 5441 1836
rect 5471 1808 5519 1836
rect 5549 1808 5558 1836
tri 5558 1808 5570 1820 sw
rect 6059 1858 6061 1860
rect 6089 1858 6091 1860
rect 6059 1836 6091 1858
rect 6012 1808 6021 1836
rect 6051 1808 6099 1836
rect 6129 1808 6138 1836
tri 6138 1808 6150 1820 sw
rect 6639 1858 6641 1860
rect 6669 1858 6671 1860
rect 6639 1836 6671 1858
rect 6592 1808 6601 1836
rect 6631 1808 6679 1836
rect 6709 1808 6718 1836
tri 6718 1808 6730 1820 sw
rect 259 1588 261 1590
rect 289 1588 291 1590
rect 259 1566 291 1588
rect 212 1538 221 1566
rect 251 1538 299 1566
rect 329 1538 338 1566
tri 338 1538 350 1550 sw
rect 839 1588 841 1590
rect 869 1588 871 1590
rect 839 1566 871 1588
rect 792 1538 801 1566
rect 831 1538 879 1566
rect 909 1538 918 1566
tri 918 1538 930 1550 sw
rect 1419 1588 1421 1590
rect 1449 1588 1451 1590
rect 1419 1566 1451 1588
rect 1372 1538 1381 1566
rect 1411 1538 1459 1566
rect 1489 1538 1498 1566
tri 1498 1538 1510 1550 sw
rect 1999 1588 2001 1590
rect 2029 1588 2031 1590
rect 1999 1566 2031 1588
rect 1952 1538 1961 1566
rect 1991 1538 2039 1566
rect 2069 1538 2078 1566
tri 2078 1538 2090 1550 sw
rect 2579 1588 2581 1590
rect 2609 1588 2611 1590
rect 2579 1566 2611 1588
rect 2532 1538 2541 1566
rect 2571 1538 2619 1566
rect 2649 1538 2658 1566
tri 2658 1538 2670 1550 sw
rect 3159 1588 3161 1590
rect 3189 1588 3191 1590
rect 3159 1566 3191 1588
rect 3112 1538 3121 1566
rect 3151 1538 3199 1566
rect 3229 1538 3238 1566
tri 3238 1538 3250 1550 sw
rect 3739 1588 3741 1590
rect 3769 1588 3771 1590
rect 3739 1566 3771 1588
rect 3692 1538 3701 1566
rect 3731 1538 3779 1566
rect 3809 1538 3818 1566
tri 3818 1538 3830 1550 sw
rect 4319 1588 4321 1590
rect 4349 1588 4351 1590
rect 4319 1566 4351 1588
rect 4272 1538 4281 1566
rect 4311 1538 4359 1566
rect 4389 1538 4398 1566
tri 4398 1538 4410 1550 sw
rect 4899 1588 4901 1590
rect 4929 1588 4931 1590
rect 4899 1566 4931 1588
rect 4852 1538 4861 1566
rect 4891 1538 4939 1566
rect 4969 1538 4978 1566
tri 4978 1538 4990 1550 sw
rect 5479 1588 5481 1590
rect 5509 1588 5511 1590
rect 5479 1566 5511 1588
rect 5432 1538 5441 1566
rect 5471 1538 5519 1566
rect 5549 1538 5558 1566
tri 5558 1538 5570 1550 sw
rect 6059 1588 6061 1590
rect 6089 1588 6091 1590
rect 6059 1566 6091 1588
rect 6012 1538 6021 1566
rect 6051 1538 6099 1566
rect 6129 1538 6138 1566
tri 6138 1538 6150 1550 sw
rect 6639 1588 6641 1590
rect 6669 1588 6671 1590
rect 6639 1566 6671 1588
rect 6592 1538 6601 1566
rect 6631 1538 6679 1566
rect 6709 1538 6718 1566
tri 6718 1538 6730 1550 sw
rect 259 1318 261 1320
rect 289 1318 291 1320
rect 259 1296 291 1318
rect 212 1268 221 1296
rect 251 1268 299 1296
rect 329 1268 338 1296
tri 338 1268 350 1280 sw
rect 839 1318 841 1320
rect 869 1318 871 1320
rect 839 1296 871 1318
rect 792 1268 801 1296
rect 831 1268 879 1296
rect 909 1268 918 1296
tri 918 1268 930 1280 sw
rect 1419 1318 1421 1320
rect 1449 1318 1451 1320
rect 1419 1296 1451 1318
rect 1372 1268 1381 1296
rect 1411 1268 1459 1296
rect 1489 1268 1498 1296
tri 1498 1268 1510 1280 sw
rect 1999 1318 2001 1320
rect 2029 1318 2031 1320
rect 1999 1296 2031 1318
rect 1952 1268 1961 1296
rect 1991 1268 2039 1296
rect 2069 1268 2078 1296
tri 2078 1268 2090 1280 sw
rect 2579 1318 2581 1320
rect 2609 1318 2611 1320
rect 2579 1296 2611 1318
rect 2532 1268 2541 1296
rect 2571 1268 2619 1296
rect 2649 1268 2658 1296
tri 2658 1268 2670 1280 sw
rect 3159 1318 3161 1320
rect 3189 1318 3191 1320
rect 3159 1296 3191 1318
rect 3112 1268 3121 1296
rect 3151 1268 3199 1296
rect 3229 1268 3238 1296
tri 3238 1268 3250 1280 sw
rect 3739 1318 3741 1320
rect 3769 1318 3771 1320
rect 3739 1296 3771 1318
rect 3692 1268 3701 1296
rect 3731 1268 3779 1296
rect 3809 1268 3818 1296
tri 3818 1268 3830 1280 sw
rect 4319 1318 4321 1320
rect 4349 1318 4351 1320
rect 4319 1296 4351 1318
rect 4272 1268 4281 1296
rect 4311 1268 4359 1296
rect 4389 1268 4398 1296
tri 4398 1268 4410 1280 sw
rect 4899 1318 4901 1320
rect 4929 1318 4931 1320
rect 4899 1296 4931 1318
rect 4852 1268 4861 1296
rect 4891 1268 4939 1296
rect 4969 1268 4978 1296
tri 4978 1268 4990 1280 sw
rect 5479 1318 5481 1320
rect 5509 1318 5511 1320
rect 5479 1296 5511 1318
rect 5432 1268 5441 1296
rect 5471 1268 5519 1296
rect 5549 1268 5558 1296
tri 5558 1268 5570 1280 sw
rect 6059 1318 6061 1320
rect 6089 1318 6091 1320
rect 6059 1296 6091 1318
rect 6012 1268 6021 1296
rect 6051 1268 6099 1296
rect 6129 1268 6138 1296
tri 6138 1268 6150 1280 sw
rect 6639 1318 6641 1320
rect 6669 1318 6671 1320
rect 6639 1296 6671 1318
rect 6592 1268 6601 1296
rect 6631 1268 6679 1296
rect 6709 1268 6718 1296
tri 6718 1268 6730 1280 sw
rect 259 1048 261 1050
rect 289 1048 291 1050
rect 259 1026 291 1048
rect 212 998 221 1026
rect 251 998 299 1026
rect 329 998 338 1026
tri 338 998 350 1010 sw
rect 839 1048 841 1050
rect 869 1048 871 1050
rect 839 1026 871 1048
rect 792 998 801 1026
rect 831 998 879 1026
rect 909 998 918 1026
tri 918 998 930 1010 sw
rect 1419 1048 1421 1050
rect 1449 1048 1451 1050
rect 1419 1026 1451 1048
rect 1372 998 1381 1026
rect 1411 998 1459 1026
rect 1489 998 1498 1026
tri 1498 998 1510 1010 sw
rect 1999 1048 2001 1050
rect 2029 1048 2031 1050
rect 1999 1026 2031 1048
rect 1952 998 1961 1026
rect 1991 998 2039 1026
rect 2069 998 2078 1026
tri 2078 998 2090 1010 sw
rect 2579 1048 2581 1050
rect 2609 1048 2611 1050
rect 2579 1026 2611 1048
rect 2532 998 2541 1026
rect 2571 998 2619 1026
rect 2649 998 2658 1026
tri 2658 998 2670 1010 sw
rect 3159 1048 3161 1050
rect 3189 1048 3191 1050
rect 3159 1026 3191 1048
rect 3112 998 3121 1026
rect 3151 998 3199 1026
rect 3229 998 3238 1026
tri 3238 998 3250 1010 sw
rect 3739 1048 3741 1050
rect 3769 1048 3771 1050
rect 3739 1026 3771 1048
rect 3692 998 3701 1026
rect 3731 998 3779 1026
rect 3809 998 3818 1026
tri 3818 998 3830 1010 sw
rect 4319 1048 4321 1050
rect 4349 1048 4351 1050
rect 4319 1026 4351 1048
rect 4272 998 4281 1026
rect 4311 998 4359 1026
rect 4389 998 4398 1026
tri 4398 998 4410 1010 sw
rect 4899 1048 4901 1050
rect 4929 1048 4931 1050
rect 4899 1026 4931 1048
rect 4852 998 4861 1026
rect 4891 998 4939 1026
rect 4969 998 4978 1026
tri 4978 998 4990 1010 sw
rect 5479 1048 5481 1050
rect 5509 1048 5511 1050
rect 5479 1026 5511 1048
rect 5432 998 5441 1026
rect 5471 998 5519 1026
rect 5549 998 5558 1026
tri 5558 998 5570 1010 sw
rect 6059 1048 6061 1050
rect 6089 1048 6091 1050
rect 6059 1026 6091 1048
rect 6012 998 6021 1026
rect 6051 998 6099 1026
rect 6129 998 6138 1026
tri 6138 998 6150 1010 sw
rect 6639 1048 6641 1050
rect 6669 1048 6671 1050
rect 6639 1026 6671 1048
rect 6592 998 6601 1026
rect 6631 998 6679 1026
rect 6709 998 6718 1026
tri 6718 998 6730 1010 sw
rect 259 778 261 780
rect 289 778 291 780
rect 259 756 291 778
rect 212 728 221 756
rect 251 728 299 756
rect 329 728 338 756
tri 338 728 350 740 sw
rect 839 778 841 780
rect 869 778 871 780
rect 839 756 871 778
rect 792 728 801 756
rect 831 728 879 756
rect 909 728 918 756
tri 918 728 930 740 sw
rect 1419 778 1421 780
rect 1449 778 1451 780
rect 1419 756 1451 778
rect 1372 728 1381 756
rect 1411 728 1459 756
rect 1489 728 1498 756
tri 1498 728 1510 740 sw
rect 1999 778 2001 780
rect 2029 778 2031 780
rect 1999 756 2031 778
rect 1952 728 1961 756
rect 1991 728 2039 756
rect 2069 728 2078 756
tri 2078 728 2090 740 sw
rect 2579 778 2581 780
rect 2609 778 2611 780
rect 2579 756 2611 778
rect 2532 728 2541 756
rect 2571 728 2619 756
rect 2649 728 2658 756
tri 2658 728 2670 740 sw
rect 3159 778 3161 780
rect 3189 778 3191 780
rect 3159 756 3191 778
rect 3112 728 3121 756
rect 3151 728 3199 756
rect 3229 728 3238 756
tri 3238 728 3250 740 sw
rect 3739 778 3741 780
rect 3769 778 3771 780
rect 3739 756 3771 778
rect 3692 728 3701 756
rect 3731 728 3779 756
rect 3809 728 3818 756
tri 3818 728 3830 740 sw
rect 4319 778 4321 780
rect 4349 778 4351 780
rect 4319 756 4351 778
rect 4272 728 4281 756
rect 4311 728 4359 756
rect 4389 728 4398 756
tri 4398 728 4410 740 sw
rect 4899 778 4901 780
rect 4929 778 4931 780
rect 4899 756 4931 778
rect 4852 728 4861 756
rect 4891 728 4939 756
rect 4969 728 4978 756
tri 4978 728 4990 740 sw
rect 5479 778 5481 780
rect 5509 778 5511 780
rect 5479 756 5511 778
rect 5432 728 5441 756
rect 5471 728 5519 756
rect 5549 728 5558 756
tri 5558 728 5570 740 sw
rect 6059 778 6061 780
rect 6089 778 6091 780
rect 6059 756 6091 778
rect 6012 728 6021 756
rect 6051 728 6099 756
rect 6129 728 6138 756
tri 6138 728 6150 740 sw
rect 6639 778 6641 780
rect 6669 778 6671 780
rect 6639 756 6671 778
rect 6592 728 6601 756
rect 6631 728 6679 756
rect 6709 728 6718 756
tri 6718 728 6730 740 sw
rect 259 508 261 510
rect 289 508 291 510
rect 259 486 291 508
rect 212 458 221 486
rect 251 458 299 486
rect 329 458 338 486
tri 338 458 350 470 sw
rect 839 508 841 510
rect 869 508 871 510
rect 839 486 871 508
rect 792 458 801 486
rect 831 458 879 486
rect 909 458 918 486
tri 918 458 930 470 sw
rect 1419 508 1421 510
rect 1449 508 1451 510
rect 1419 486 1451 508
rect 1372 458 1381 486
rect 1411 458 1459 486
rect 1489 458 1498 486
tri 1498 458 1510 470 sw
rect 1999 508 2001 510
rect 2029 508 2031 510
rect 1999 486 2031 508
rect 1952 458 1961 486
rect 1991 458 2039 486
rect 2069 458 2078 486
tri 2078 458 2090 470 sw
rect 2579 508 2581 510
rect 2609 508 2611 510
rect 2579 486 2611 508
rect 2532 458 2541 486
rect 2571 458 2619 486
rect 2649 458 2658 486
tri 2658 458 2670 470 sw
rect 3159 508 3161 510
rect 3189 508 3191 510
rect 3159 486 3191 508
rect 3112 458 3121 486
rect 3151 458 3199 486
rect 3229 458 3238 486
tri 3238 458 3250 470 sw
rect 3739 508 3741 510
rect 3769 508 3771 510
rect 3739 486 3771 508
rect 3692 458 3701 486
rect 3731 458 3779 486
rect 3809 458 3818 486
tri 3818 458 3830 470 sw
rect 4319 508 4321 510
rect 4349 508 4351 510
rect 4319 486 4351 508
rect 4272 458 4281 486
rect 4311 458 4359 486
rect 4389 458 4398 486
tri 4398 458 4410 470 sw
rect 4899 508 4901 510
rect 4929 508 4931 510
rect 4899 486 4931 508
rect 4852 458 4861 486
rect 4891 458 4939 486
rect 4969 458 4978 486
tri 4978 458 4990 470 sw
rect 5479 508 5481 510
rect 5509 508 5511 510
rect 5479 486 5511 508
rect 5432 458 5441 486
rect 5471 458 5519 486
rect 5549 458 5558 486
tri 5558 458 5570 470 sw
rect 6059 508 6061 510
rect 6089 508 6091 510
rect 6059 486 6091 508
rect 6012 458 6021 486
rect 6051 458 6099 486
rect 6129 458 6138 486
tri 6138 458 6150 470 sw
rect 6639 508 6641 510
rect 6669 508 6671 510
rect 6639 486 6671 508
rect 6592 458 6601 486
rect 6631 458 6679 486
rect 6709 458 6718 486
tri 6718 458 6730 470 sw
rect 259 238 261 240
rect 289 238 291 240
rect 259 216 291 238
rect 212 188 221 216
rect 251 188 299 216
rect 329 188 338 216
tri 338 188 350 200 sw
rect 839 238 841 240
rect 869 238 871 240
rect 839 216 871 238
rect 792 188 801 216
rect 831 188 879 216
rect 909 188 918 216
tri 918 188 930 200 sw
rect 1419 238 1421 240
rect 1449 238 1451 240
rect 1419 216 1451 238
rect 1372 188 1381 216
rect 1411 188 1459 216
rect 1489 188 1498 216
tri 1498 188 1510 200 sw
rect 1999 238 2001 240
rect 2029 238 2031 240
rect 1999 216 2031 238
rect 1952 188 1961 216
rect 1991 188 2039 216
rect 2069 188 2078 216
tri 2078 188 2090 200 sw
rect 2579 238 2581 240
rect 2609 238 2611 240
rect 2579 216 2611 238
rect 2532 188 2541 216
rect 2571 188 2619 216
rect 2649 188 2658 216
tri 2658 188 2670 200 sw
rect 3159 238 3161 240
rect 3189 238 3191 240
rect 3159 216 3191 238
rect 3112 188 3121 216
rect 3151 188 3199 216
rect 3229 188 3238 216
tri 3238 188 3250 200 sw
rect 3739 238 3741 240
rect 3769 238 3771 240
rect 3739 216 3771 238
rect 3692 188 3701 216
rect 3731 188 3779 216
rect 3809 188 3818 216
tri 3818 188 3830 200 sw
rect 4319 238 4321 240
rect 4349 238 4351 240
rect 4319 216 4351 238
rect 4272 188 4281 216
rect 4311 188 4359 216
rect 4389 188 4398 216
tri 4398 188 4410 200 sw
rect 4899 238 4901 240
rect 4929 238 4931 240
rect 4899 216 4931 238
rect 4852 188 4861 216
rect 4891 188 4939 216
rect 4969 188 4978 216
tri 4978 188 4990 200 sw
rect 5479 238 5481 240
rect 5509 238 5511 240
rect 5479 216 5511 238
rect 5432 188 5441 216
rect 5471 188 5519 216
rect 5549 188 5558 216
tri 5558 188 5570 200 sw
rect 6059 238 6061 240
rect 6089 238 6091 240
rect 6059 216 6091 238
rect 6012 188 6021 216
rect 6051 188 6099 216
rect 6129 188 6138 216
tri 6138 188 6150 200 sw
rect 6639 238 6641 240
rect 6669 238 6671 240
rect 6639 216 6671 238
rect 6592 188 6601 216
rect 6631 188 6679 216
rect 6709 188 6718 216
tri 6718 188 6730 200 sw
rect 259 -32 261 -30
rect 289 -32 291 -30
rect 259 -54 291 -32
rect 212 -82 221 -54
rect 251 -82 299 -54
rect 329 -82 338 -54
tri 338 -82 350 -70 sw
rect 839 -32 841 -30
rect 869 -32 871 -30
rect 839 -54 871 -32
rect 792 -82 801 -54
rect 831 -82 879 -54
rect 909 -82 918 -54
tri 918 -82 930 -70 sw
rect 1419 -32 1421 -30
rect 1449 -32 1451 -30
rect 1419 -54 1451 -32
rect 1372 -82 1381 -54
rect 1411 -82 1459 -54
rect 1489 -82 1498 -54
tri 1498 -82 1510 -70 sw
rect 1999 -32 2001 -30
rect 2029 -32 2031 -30
rect 1999 -54 2031 -32
rect 1952 -82 1961 -54
rect 1991 -82 2039 -54
rect 2069 -82 2078 -54
tri 2078 -82 2090 -70 sw
rect 2579 -32 2581 -30
rect 2609 -32 2611 -30
rect 2579 -54 2611 -32
rect 2532 -82 2541 -54
rect 2571 -82 2619 -54
rect 2649 -82 2658 -54
tri 2658 -82 2670 -70 sw
rect 3159 -32 3161 -30
rect 3189 -32 3191 -30
rect 3159 -54 3191 -32
rect 3112 -82 3121 -54
rect 3151 -82 3199 -54
rect 3229 -82 3238 -54
tri 3238 -82 3250 -70 sw
rect 3739 -32 3741 -30
rect 3769 -32 3771 -30
rect 3739 -54 3771 -32
rect 3692 -82 3701 -54
rect 3731 -82 3779 -54
rect 3809 -82 3818 -54
tri 3818 -82 3830 -70 sw
rect 4319 -32 4321 -30
rect 4349 -32 4351 -30
rect 4319 -54 4351 -32
rect 4272 -82 4281 -54
rect 4311 -82 4359 -54
rect 4389 -82 4398 -54
tri 4398 -82 4410 -70 sw
rect 4899 -32 4901 -30
rect 4929 -32 4931 -30
rect 4899 -54 4931 -32
rect 4852 -82 4861 -54
rect 4891 -82 4939 -54
rect 4969 -82 4978 -54
tri 4978 -82 4990 -70 sw
rect 5479 -32 5481 -30
rect 5509 -32 5511 -30
rect 5479 -54 5511 -32
rect 5432 -82 5441 -54
rect 5471 -82 5519 -54
rect 5549 -82 5558 -54
tri 5558 -82 5570 -70 sw
rect 6059 -32 6061 -30
rect 6089 -32 6091 -30
rect 6059 -54 6091 -32
rect 6012 -82 6021 -54
rect 6051 -82 6099 -54
rect 6129 -82 6138 -54
tri 6138 -82 6150 -70 sw
rect 6639 -32 6641 -30
rect 6669 -32 6671 -30
rect 6639 -54 6671 -32
rect 6592 -82 6601 -54
rect 6631 -82 6679 -54
rect 6709 -82 6718 -54
tri 6718 -82 6730 -70 sw
rect 259 -302 261 -300
rect 289 -302 291 -300
rect 259 -324 291 -302
rect 212 -352 221 -324
rect 251 -352 299 -324
rect 329 -352 338 -324
tri 338 -352 350 -340 sw
rect 839 -302 841 -300
rect 869 -302 871 -300
rect 839 -324 871 -302
rect 792 -352 801 -324
rect 831 -352 879 -324
rect 909 -352 918 -324
tri 918 -352 930 -340 sw
rect 1419 -302 1421 -300
rect 1449 -302 1451 -300
rect 1419 -324 1451 -302
rect 1372 -352 1381 -324
rect 1411 -352 1459 -324
rect 1489 -352 1498 -324
tri 1498 -352 1510 -340 sw
rect 1999 -302 2001 -300
rect 2029 -302 2031 -300
rect 1999 -324 2031 -302
rect 1952 -352 1961 -324
rect 1991 -352 2039 -324
rect 2069 -352 2078 -324
tri 2078 -352 2090 -340 sw
rect 2579 -302 2581 -300
rect 2609 -302 2611 -300
rect 2579 -324 2611 -302
rect 2532 -352 2541 -324
rect 2571 -352 2619 -324
rect 2649 -352 2658 -324
tri 2658 -352 2670 -340 sw
rect 3159 -302 3161 -300
rect 3189 -302 3191 -300
rect 3159 -324 3191 -302
rect 3112 -352 3121 -324
rect 3151 -352 3199 -324
rect 3229 -352 3238 -324
tri 3238 -352 3250 -340 sw
rect 3739 -302 3741 -300
rect 3769 -302 3771 -300
rect 3739 -324 3771 -302
rect 3692 -352 3701 -324
rect 3731 -352 3779 -324
rect 3809 -352 3818 -324
tri 3818 -352 3830 -340 sw
rect 4319 -302 4321 -300
rect 4349 -302 4351 -300
rect 4319 -324 4351 -302
rect 4272 -352 4281 -324
rect 4311 -352 4359 -324
rect 4389 -352 4398 -324
tri 4398 -352 4410 -340 sw
rect 4899 -302 4901 -300
rect 4929 -302 4931 -300
rect 4899 -324 4931 -302
rect 4852 -352 4861 -324
rect 4891 -352 4939 -324
rect 4969 -352 4978 -324
tri 4978 -352 4990 -340 sw
rect 5479 -302 5481 -300
rect 5509 -302 5511 -300
rect 5479 -324 5511 -302
rect 5432 -352 5441 -324
rect 5471 -352 5519 -324
rect 5549 -352 5558 -324
tri 5558 -352 5570 -340 sw
rect 6059 -302 6061 -300
rect 6089 -302 6091 -300
rect 6059 -324 6091 -302
rect 6012 -352 6021 -324
rect 6051 -352 6099 -324
rect 6129 -352 6138 -324
tri 6138 -352 6150 -340 sw
rect 6639 -302 6641 -300
rect 6669 -302 6671 -300
rect 6639 -324 6671 -302
rect 6592 -352 6601 -324
rect 6631 -352 6679 -324
rect 6709 -352 6718 -324
tri 6718 -352 6730 -340 sw
rect 259 -572 261 -570
rect 289 -572 291 -570
rect 259 -594 291 -572
rect 212 -622 221 -594
rect 251 -622 299 -594
rect 329 -622 338 -594
tri 338 -622 350 -610 sw
rect 839 -572 841 -570
rect 869 -572 871 -570
rect 839 -594 871 -572
rect 792 -622 801 -594
rect 831 -622 879 -594
rect 909 -622 918 -594
tri 918 -622 930 -610 sw
rect 1419 -572 1421 -570
rect 1449 -572 1451 -570
rect 1419 -594 1451 -572
rect 1372 -622 1381 -594
rect 1411 -622 1459 -594
rect 1489 -622 1498 -594
tri 1498 -622 1510 -610 sw
rect 1999 -572 2001 -570
rect 2029 -572 2031 -570
rect 1999 -594 2031 -572
rect 1952 -622 1961 -594
rect 1991 -622 2039 -594
rect 2069 -622 2078 -594
tri 2078 -622 2090 -610 sw
rect 2579 -572 2581 -570
rect 2609 -572 2611 -570
rect 2579 -594 2611 -572
rect 2532 -622 2541 -594
rect 2571 -622 2619 -594
rect 2649 -622 2658 -594
tri 2658 -622 2670 -610 sw
rect 3159 -572 3161 -570
rect 3189 -572 3191 -570
rect 3159 -594 3191 -572
rect 3112 -622 3121 -594
rect 3151 -622 3199 -594
rect 3229 -622 3238 -594
tri 3238 -622 3250 -610 sw
rect 3739 -572 3741 -570
rect 3769 -572 3771 -570
rect 3739 -594 3771 -572
rect 3692 -622 3701 -594
rect 3731 -622 3779 -594
rect 3809 -622 3818 -594
tri 3818 -622 3830 -610 sw
rect 4319 -572 4321 -570
rect 4349 -572 4351 -570
rect 4319 -594 4351 -572
rect 4272 -622 4281 -594
rect 4311 -622 4359 -594
rect 4389 -622 4398 -594
tri 4398 -622 4410 -610 sw
rect 4899 -572 4901 -570
rect 4929 -572 4931 -570
rect 4899 -594 4931 -572
rect 4852 -622 4861 -594
rect 4891 -622 4939 -594
rect 4969 -622 4978 -594
tri 4978 -622 4990 -610 sw
rect 5479 -572 5481 -570
rect 5509 -572 5511 -570
rect 5479 -594 5511 -572
rect 5432 -622 5441 -594
rect 5471 -622 5519 -594
rect 5549 -622 5558 -594
tri 5558 -622 5570 -610 sw
rect 6059 -572 6061 -570
rect 6089 -572 6091 -570
rect 6059 -594 6091 -572
rect 6012 -622 6021 -594
rect 6051 -622 6099 -594
rect 6129 -622 6138 -594
tri 6138 -622 6150 -610 sw
rect 6639 -572 6641 -570
rect 6669 -572 6671 -570
rect 6639 -594 6671 -572
rect 6592 -622 6601 -594
rect 6631 -622 6679 -594
rect 6709 -622 6718 -594
tri 6718 -622 6730 -610 sw
rect 259 -842 261 -840
rect 289 -842 291 -840
rect 259 -864 291 -842
rect 212 -892 221 -864
rect 251 -892 299 -864
rect 329 -892 338 -864
tri 338 -892 350 -880 sw
rect 839 -842 841 -840
rect 869 -842 871 -840
rect 839 -864 871 -842
rect 792 -892 801 -864
rect 831 -892 879 -864
rect 909 -892 918 -864
tri 918 -892 930 -880 sw
rect 1419 -842 1421 -840
rect 1449 -842 1451 -840
rect 1419 -864 1451 -842
rect 1372 -892 1381 -864
rect 1411 -892 1459 -864
rect 1489 -892 1498 -864
tri 1498 -892 1510 -880 sw
rect 1999 -842 2001 -840
rect 2029 -842 2031 -840
rect 1999 -864 2031 -842
rect 1952 -892 1961 -864
rect 1991 -892 2039 -864
rect 2069 -892 2078 -864
tri 2078 -892 2090 -880 sw
rect 2579 -842 2581 -840
rect 2609 -842 2611 -840
rect 2579 -864 2611 -842
rect 2532 -892 2541 -864
rect 2571 -892 2619 -864
rect 2649 -892 2658 -864
tri 2658 -892 2670 -880 sw
rect 3159 -842 3161 -840
rect 3189 -842 3191 -840
rect 3159 -864 3191 -842
rect 3112 -892 3121 -864
rect 3151 -892 3199 -864
rect 3229 -892 3238 -864
tri 3238 -892 3250 -880 sw
rect 3739 -842 3741 -840
rect 3769 -842 3771 -840
rect 3739 -864 3771 -842
rect 3692 -892 3701 -864
rect 3731 -892 3779 -864
rect 3809 -892 3818 -864
tri 3818 -892 3830 -880 sw
rect 4319 -842 4321 -840
rect 4349 -842 4351 -840
rect 4319 -864 4351 -842
rect 4272 -892 4281 -864
rect 4311 -892 4359 -864
rect 4389 -892 4398 -864
tri 4398 -892 4410 -880 sw
rect 4899 -842 4901 -840
rect 4929 -842 4931 -840
rect 4899 -864 4931 -842
rect 4852 -892 4861 -864
rect 4891 -892 4939 -864
rect 4969 -892 4978 -864
tri 4978 -892 4990 -880 sw
rect 5479 -842 5481 -840
rect 5509 -842 5511 -840
rect 5479 -864 5511 -842
rect 5432 -892 5441 -864
rect 5471 -892 5519 -864
rect 5549 -892 5558 -864
tri 5558 -892 5570 -880 sw
rect 6059 -842 6061 -840
rect 6089 -842 6091 -840
rect 6059 -864 6091 -842
rect 6012 -892 6021 -864
rect 6051 -892 6099 -864
rect 6129 -892 6138 -864
tri 6138 -892 6150 -880 sw
rect 6639 -842 6641 -840
rect 6669 -842 6671 -840
rect 6639 -864 6671 -842
rect 6592 -892 6601 -864
rect 6631 -892 6679 -864
rect 6709 -892 6718 -864
tri 6718 -892 6730 -880 sw
rect 259 -1112 261 -1110
rect 289 -1112 291 -1110
rect 259 -1134 291 -1112
rect 212 -1162 221 -1134
rect 251 -1162 299 -1134
rect 329 -1162 338 -1134
tri 338 -1162 350 -1150 sw
rect 839 -1112 841 -1110
rect 869 -1112 871 -1110
rect 839 -1134 871 -1112
rect 792 -1162 801 -1134
rect 831 -1162 879 -1134
rect 909 -1162 918 -1134
tri 918 -1162 930 -1150 sw
rect 1419 -1112 1421 -1110
rect 1449 -1112 1451 -1110
rect 1419 -1134 1451 -1112
rect 1372 -1162 1381 -1134
rect 1411 -1162 1459 -1134
rect 1489 -1162 1498 -1134
tri 1498 -1162 1510 -1150 sw
rect 1999 -1112 2001 -1110
rect 2029 -1112 2031 -1110
rect 1999 -1134 2031 -1112
rect 1952 -1162 1961 -1134
rect 1991 -1162 2039 -1134
rect 2069 -1162 2078 -1134
tri 2078 -1162 2090 -1150 sw
rect 2579 -1112 2581 -1110
rect 2609 -1112 2611 -1110
rect 2579 -1134 2611 -1112
rect 2532 -1162 2541 -1134
rect 2571 -1162 2619 -1134
rect 2649 -1162 2658 -1134
tri 2658 -1162 2670 -1150 sw
rect 3159 -1112 3161 -1110
rect 3189 -1112 3191 -1110
rect 3159 -1134 3191 -1112
rect 3112 -1162 3121 -1134
rect 3151 -1162 3199 -1134
rect 3229 -1162 3238 -1134
tri 3238 -1162 3250 -1150 sw
rect 3739 -1112 3741 -1110
rect 3769 -1112 3771 -1110
rect 3739 -1134 3771 -1112
rect 3692 -1162 3701 -1134
rect 3731 -1162 3779 -1134
rect 3809 -1162 3818 -1134
tri 3818 -1162 3830 -1150 sw
rect 4319 -1112 4321 -1110
rect 4349 -1112 4351 -1110
rect 4319 -1134 4351 -1112
rect 4272 -1162 4281 -1134
rect 4311 -1162 4359 -1134
rect 4389 -1162 4398 -1134
tri 4398 -1162 4410 -1150 sw
rect 4899 -1112 4901 -1110
rect 4929 -1112 4931 -1110
rect 4899 -1134 4931 -1112
rect 4852 -1162 4861 -1134
rect 4891 -1162 4939 -1134
rect 4969 -1162 4978 -1134
tri 4978 -1162 4990 -1150 sw
rect 5479 -1112 5481 -1110
rect 5509 -1112 5511 -1110
rect 5479 -1134 5511 -1112
rect 5432 -1162 5441 -1134
rect 5471 -1162 5519 -1134
rect 5549 -1162 5558 -1134
tri 5558 -1162 5570 -1150 sw
rect 6059 -1112 6061 -1110
rect 6089 -1112 6091 -1110
rect 6059 -1134 6091 -1112
rect 6012 -1162 6021 -1134
rect 6051 -1162 6099 -1134
rect 6129 -1162 6138 -1134
tri 6138 -1162 6150 -1150 sw
rect 6639 -1112 6641 -1110
rect 6669 -1112 6671 -1110
rect 6639 -1134 6671 -1112
rect 6592 -1162 6601 -1134
rect 6631 -1162 6679 -1134
rect 6709 -1162 6718 -1134
tri 6718 -1162 6730 -1150 sw
rect 259 -1382 261 -1380
rect 289 -1382 291 -1380
rect 259 -1404 291 -1382
rect 212 -1432 221 -1404
rect 251 -1432 299 -1404
rect 329 -1432 338 -1404
tri 338 -1432 350 -1420 sw
rect 839 -1382 841 -1380
rect 869 -1382 871 -1380
rect 839 -1404 871 -1382
rect 792 -1432 801 -1404
rect 831 -1432 879 -1404
rect 909 -1432 918 -1404
tri 918 -1432 930 -1420 sw
rect 1419 -1382 1421 -1380
rect 1449 -1382 1451 -1380
rect 1419 -1404 1451 -1382
rect 1372 -1432 1381 -1404
rect 1411 -1432 1459 -1404
rect 1489 -1432 1498 -1404
tri 1498 -1432 1510 -1420 sw
rect 1999 -1382 2001 -1380
rect 2029 -1382 2031 -1380
rect 1999 -1404 2031 -1382
rect 1952 -1432 1961 -1404
rect 1991 -1432 2039 -1404
rect 2069 -1432 2078 -1404
tri 2078 -1432 2090 -1420 sw
rect 2579 -1382 2581 -1380
rect 2609 -1382 2611 -1380
rect 2579 -1404 2611 -1382
rect 2532 -1432 2541 -1404
rect 2571 -1432 2619 -1404
rect 2649 -1432 2658 -1404
tri 2658 -1432 2670 -1420 sw
rect 3159 -1382 3161 -1380
rect 3189 -1382 3191 -1380
rect 3159 -1404 3191 -1382
rect 3112 -1432 3121 -1404
rect 3151 -1432 3199 -1404
rect 3229 -1432 3238 -1404
tri 3238 -1432 3250 -1420 sw
rect 3739 -1382 3741 -1380
rect 3769 -1382 3771 -1380
rect 3739 -1404 3771 -1382
rect 3692 -1432 3701 -1404
rect 3731 -1432 3779 -1404
rect 3809 -1432 3818 -1404
tri 3818 -1432 3830 -1420 sw
rect 4319 -1382 4321 -1380
rect 4349 -1382 4351 -1380
rect 4319 -1404 4351 -1382
rect 4272 -1432 4281 -1404
rect 4311 -1432 4359 -1404
rect 4389 -1432 4398 -1404
tri 4398 -1432 4410 -1420 sw
rect 4899 -1382 4901 -1380
rect 4929 -1382 4931 -1380
rect 4899 -1404 4931 -1382
rect 4852 -1432 4861 -1404
rect 4891 -1432 4939 -1404
rect 4969 -1432 4978 -1404
tri 4978 -1432 4990 -1420 sw
rect 5479 -1382 5481 -1380
rect 5509 -1382 5511 -1380
rect 5479 -1404 5511 -1382
rect 5432 -1432 5441 -1404
rect 5471 -1432 5519 -1404
rect 5549 -1432 5558 -1404
tri 5558 -1432 5570 -1420 sw
rect 6059 -1382 6061 -1380
rect 6089 -1382 6091 -1380
rect 6059 -1404 6091 -1382
rect 6012 -1432 6021 -1404
rect 6051 -1432 6099 -1404
rect 6129 -1432 6138 -1404
tri 6138 -1432 6150 -1420 sw
rect 6639 -1382 6641 -1380
rect 6669 -1382 6671 -1380
rect 6639 -1404 6671 -1382
rect 6592 -1432 6601 -1404
rect 6631 -1432 6679 -1404
rect 6709 -1432 6718 -1404
tri 6718 -1432 6730 -1420 sw
rect 259 -1652 261 -1650
rect 289 -1652 291 -1650
rect 259 -1674 291 -1652
rect 212 -1702 221 -1674
rect 251 -1702 299 -1674
rect 329 -1702 338 -1674
tri 338 -1702 350 -1690 sw
rect 839 -1652 841 -1650
rect 869 -1652 871 -1650
rect 839 -1674 871 -1652
rect 792 -1702 801 -1674
rect 831 -1702 879 -1674
rect 909 -1702 918 -1674
tri 918 -1702 930 -1690 sw
rect 1419 -1652 1421 -1650
rect 1449 -1652 1451 -1650
rect 1419 -1674 1451 -1652
rect 1372 -1702 1381 -1674
rect 1411 -1702 1459 -1674
rect 1489 -1702 1498 -1674
tri 1498 -1702 1510 -1690 sw
rect 1999 -1652 2001 -1650
rect 2029 -1652 2031 -1650
rect 1999 -1674 2031 -1652
rect 1952 -1702 1961 -1674
rect 1991 -1702 2039 -1674
rect 2069 -1702 2078 -1674
tri 2078 -1702 2090 -1690 sw
rect 2579 -1652 2581 -1650
rect 2609 -1652 2611 -1650
rect 2579 -1674 2611 -1652
rect 2532 -1702 2541 -1674
rect 2571 -1702 2619 -1674
rect 2649 -1702 2658 -1674
tri 2658 -1702 2670 -1690 sw
rect 3159 -1652 3161 -1650
rect 3189 -1652 3191 -1650
rect 3159 -1674 3191 -1652
rect 3112 -1702 3121 -1674
rect 3151 -1702 3199 -1674
rect 3229 -1702 3238 -1674
tri 3238 -1702 3250 -1690 sw
rect 3739 -1652 3741 -1650
rect 3769 -1652 3771 -1650
rect 3739 -1674 3771 -1652
rect 3692 -1702 3701 -1674
rect 3731 -1702 3779 -1674
rect 3809 -1702 3818 -1674
tri 3818 -1702 3830 -1690 sw
rect 4319 -1652 4321 -1650
rect 4349 -1652 4351 -1650
rect 4319 -1674 4351 -1652
rect 4272 -1702 4281 -1674
rect 4311 -1702 4359 -1674
rect 4389 -1702 4398 -1674
tri 4398 -1702 4410 -1690 sw
rect 4899 -1652 4901 -1650
rect 4929 -1652 4931 -1650
rect 4899 -1674 4931 -1652
rect 4852 -1702 4861 -1674
rect 4891 -1702 4939 -1674
rect 4969 -1702 4978 -1674
tri 4978 -1702 4990 -1690 sw
rect 5479 -1652 5481 -1650
rect 5509 -1652 5511 -1650
rect 5479 -1674 5511 -1652
rect 5432 -1702 5441 -1674
rect 5471 -1702 5519 -1674
rect 5549 -1702 5558 -1674
tri 5558 -1702 5570 -1690 sw
rect 6059 -1652 6061 -1650
rect 6089 -1652 6091 -1650
rect 6059 -1674 6091 -1652
rect 6012 -1702 6021 -1674
rect 6051 -1702 6099 -1674
rect 6129 -1702 6138 -1674
tri 6138 -1702 6150 -1690 sw
rect 6639 -1652 6641 -1650
rect 6669 -1652 6671 -1650
rect 6639 -1674 6671 -1652
rect 6592 -1702 6601 -1674
rect 6631 -1702 6679 -1674
rect 6709 -1702 6718 -1674
tri 6718 -1702 6730 -1690 sw
rect 259 -1922 261 -1920
rect 289 -1922 291 -1920
rect 259 -1944 291 -1922
rect 212 -1972 221 -1944
rect 251 -1972 299 -1944
rect 329 -1972 338 -1944
tri 338 -1972 350 -1960 sw
rect 839 -1922 841 -1920
rect 869 -1922 871 -1920
rect 839 -1944 871 -1922
rect 792 -1972 801 -1944
rect 831 -1972 879 -1944
rect 909 -1972 918 -1944
tri 918 -1972 930 -1960 sw
rect 1419 -1922 1421 -1920
rect 1449 -1922 1451 -1920
rect 1419 -1944 1451 -1922
rect 1372 -1972 1381 -1944
rect 1411 -1972 1459 -1944
rect 1489 -1972 1498 -1944
tri 1498 -1972 1510 -1960 sw
rect 1999 -1922 2001 -1920
rect 2029 -1922 2031 -1920
rect 1999 -1944 2031 -1922
rect 1952 -1972 1961 -1944
rect 1991 -1972 2039 -1944
rect 2069 -1972 2078 -1944
tri 2078 -1972 2090 -1960 sw
rect 2579 -1922 2581 -1920
rect 2609 -1922 2611 -1920
rect 2579 -1944 2611 -1922
rect 2532 -1972 2541 -1944
rect 2571 -1972 2619 -1944
rect 2649 -1972 2658 -1944
tri 2658 -1972 2670 -1960 sw
rect 3159 -1922 3161 -1920
rect 3189 -1922 3191 -1920
rect 3159 -1944 3191 -1922
rect 3112 -1972 3121 -1944
rect 3151 -1972 3199 -1944
rect 3229 -1972 3238 -1944
tri 3238 -1972 3250 -1960 sw
rect 3739 -1922 3741 -1920
rect 3769 -1922 3771 -1920
rect 3739 -1944 3771 -1922
rect 3692 -1972 3701 -1944
rect 3731 -1972 3779 -1944
rect 3809 -1972 3818 -1944
tri 3818 -1972 3830 -1960 sw
rect 4319 -1922 4321 -1920
rect 4349 -1922 4351 -1920
rect 4319 -1944 4351 -1922
rect 4272 -1972 4281 -1944
rect 4311 -1972 4359 -1944
rect 4389 -1972 4398 -1944
tri 4398 -1972 4410 -1960 sw
rect 4899 -1922 4901 -1920
rect 4929 -1922 4931 -1920
rect 4899 -1944 4931 -1922
rect 4852 -1972 4861 -1944
rect 4891 -1972 4939 -1944
rect 4969 -1972 4978 -1944
tri 4978 -1972 4990 -1960 sw
rect 5479 -1922 5481 -1920
rect 5509 -1922 5511 -1920
rect 5479 -1944 5511 -1922
rect 5432 -1972 5441 -1944
rect 5471 -1972 5519 -1944
rect 5549 -1972 5558 -1944
tri 5558 -1972 5570 -1960 sw
rect 6059 -1922 6061 -1920
rect 6089 -1922 6091 -1920
rect 6059 -1944 6091 -1922
rect 6012 -1972 6021 -1944
rect 6051 -1972 6099 -1944
rect 6129 -1972 6138 -1944
tri 6138 -1972 6150 -1960 sw
rect 6639 -1922 6641 -1920
rect 6669 -1922 6671 -1920
rect 6639 -1944 6671 -1922
rect 6592 -1972 6601 -1944
rect 6631 -1972 6679 -1944
rect 6709 -1972 6718 -1944
tri 6718 -1972 6730 -1960 sw
<< ndiffc >>
rect 73 2088 88 2116
rect 154 2088 169 2116
rect 381 2088 396 2116
rect 463 2088 478 2117
rect 653 2088 668 2116
rect 734 2088 749 2116
rect 961 2088 976 2116
rect 1043 2088 1058 2117
rect 1233 2088 1248 2116
rect 1314 2088 1329 2116
rect 1541 2088 1556 2116
rect 1623 2088 1638 2117
rect 1813 2088 1828 2116
rect 1894 2088 1909 2116
rect 2121 2088 2136 2116
rect 2203 2088 2218 2117
rect 2393 2088 2408 2116
rect 2474 2088 2489 2116
rect 2701 2088 2716 2116
rect 2783 2088 2798 2117
rect 2973 2088 2988 2116
rect 3054 2088 3069 2116
rect 3281 2088 3296 2116
rect 3363 2088 3378 2117
rect 3553 2088 3568 2116
rect 3634 2088 3649 2116
rect 3861 2088 3876 2116
rect 3943 2088 3958 2117
rect 4133 2088 4148 2116
rect 4214 2088 4229 2116
rect 4441 2088 4456 2116
rect 4523 2088 4538 2117
rect 4713 2088 4728 2116
rect 4794 2088 4809 2116
rect 5021 2088 5036 2116
rect 5103 2088 5118 2117
rect 5293 2088 5308 2116
rect 5374 2088 5389 2116
rect 5601 2088 5616 2116
rect 5683 2088 5698 2117
rect 5873 2088 5888 2116
rect 5954 2088 5969 2116
rect 6181 2088 6196 2116
rect 6263 2088 6278 2117
rect 6453 2088 6468 2116
rect 6534 2088 6549 2116
rect 6761 2088 6776 2116
rect 6843 2088 6858 2117
rect -1 1942 14 1984
rect 196 1967 206 1974
tri 206 1967 213 1974 sw
rect 196 1942 213 1967
rect 337 1942 354 1974
rect 536 1942 551 1984
rect 579 1942 594 1984
rect 776 1967 786 1974
tri 786 1967 793 1974 sw
rect 776 1942 793 1967
rect 917 1942 934 1974
rect 1116 1942 1131 1984
rect 1159 1942 1174 1984
rect 1356 1967 1366 1974
tri 1366 1967 1373 1974 sw
rect 1356 1942 1373 1967
rect 1497 1942 1514 1974
rect 1696 1942 1711 1984
rect 1739 1942 1754 1984
rect 1936 1967 1946 1974
tri 1946 1967 1953 1974 sw
rect 1936 1942 1953 1967
rect 2077 1942 2094 1974
rect 2276 1942 2291 1984
rect 2319 1942 2334 1984
rect 2516 1967 2526 1974
tri 2526 1967 2533 1974 sw
rect 2516 1942 2533 1967
rect 2657 1942 2674 1974
rect 2856 1942 2871 1984
rect 2899 1942 2914 1984
rect 3096 1967 3106 1974
tri 3106 1967 3113 1974 sw
rect 3096 1942 3113 1967
rect 3237 1942 3254 1974
rect 3436 1942 3451 1984
rect 3479 1942 3494 1984
rect 3676 1967 3686 1974
tri 3686 1967 3693 1974 sw
rect 3676 1942 3693 1967
rect 3817 1942 3834 1974
rect 4016 1942 4031 1984
rect 4059 1942 4074 1984
rect 4256 1967 4266 1974
tri 4266 1967 4273 1974 sw
rect 4256 1942 4273 1967
rect 4397 1942 4414 1974
rect 4596 1942 4611 1984
rect 4639 1942 4654 1984
rect 4836 1967 4846 1974
tri 4846 1967 4853 1974 sw
rect 4836 1942 4853 1967
rect 4977 1942 4994 1974
rect 5176 1942 5191 1984
rect 5219 1942 5234 1984
rect 5416 1967 5426 1974
tri 5426 1967 5433 1974 sw
rect 5416 1942 5433 1967
rect 5557 1942 5574 1974
rect 5756 1942 5771 1984
rect 5799 1942 5814 1984
rect 5996 1967 6006 1974
tri 6006 1967 6013 1974 sw
rect 5996 1942 6013 1967
rect 6137 1942 6154 1974
rect 6336 1942 6351 1984
rect 6379 1942 6394 1984
rect 6576 1967 6586 1974
tri 6586 1967 6593 1974 sw
rect 6576 1942 6593 1967
rect 6717 1942 6734 1974
rect 6916 1942 6931 1984
rect 259 1904 291 1918
rect 839 1904 871 1918
rect 1419 1904 1451 1918
rect 1999 1904 2031 1918
rect 2579 1904 2611 1918
rect 3159 1904 3191 1918
rect 3739 1904 3771 1918
rect 4319 1904 4351 1918
rect 4899 1904 4931 1918
rect 5479 1904 5511 1918
rect 6059 1904 6091 1918
rect 6639 1904 6671 1918
rect 73 1818 88 1846
rect 154 1818 169 1846
rect 381 1818 396 1846
rect 463 1818 478 1847
rect 653 1818 668 1846
rect 734 1818 749 1846
rect 961 1818 976 1846
rect 1043 1818 1058 1847
rect 1233 1818 1248 1846
rect 1314 1818 1329 1846
rect 1541 1818 1556 1846
rect 1623 1818 1638 1847
rect 1813 1818 1828 1846
rect 1894 1818 1909 1846
rect 2121 1818 2136 1846
rect 2203 1818 2218 1847
rect 2393 1818 2408 1846
rect 2474 1818 2489 1846
rect 2701 1818 2716 1846
rect 2783 1818 2798 1847
rect 2973 1818 2988 1846
rect 3054 1818 3069 1846
rect 3281 1818 3296 1846
rect 3363 1818 3378 1847
rect 3553 1818 3568 1846
rect 3634 1818 3649 1846
rect 3861 1818 3876 1846
rect 3943 1818 3958 1847
rect 4133 1818 4148 1846
rect 4214 1818 4229 1846
rect 4441 1818 4456 1846
rect 4523 1818 4538 1847
rect 4713 1818 4728 1846
rect 4794 1818 4809 1846
rect 5021 1818 5036 1846
rect 5103 1818 5118 1847
rect 5293 1818 5308 1846
rect 5374 1818 5389 1846
rect 5601 1818 5616 1846
rect 5683 1818 5698 1847
rect 5873 1818 5888 1846
rect 5954 1818 5969 1846
rect 6181 1818 6196 1846
rect 6263 1818 6278 1847
rect 6453 1818 6468 1846
rect 6534 1818 6549 1846
rect 6761 1818 6776 1846
rect 6843 1818 6858 1847
rect -1 1672 14 1714
rect 196 1697 206 1704
tri 206 1697 213 1704 sw
rect 196 1672 213 1697
rect 337 1672 354 1704
rect 536 1672 551 1714
rect 579 1672 594 1714
rect 776 1697 786 1704
tri 786 1697 793 1704 sw
rect 776 1672 793 1697
rect 917 1672 934 1704
rect 1116 1672 1131 1714
rect 1159 1672 1174 1714
rect 1356 1697 1366 1704
tri 1366 1697 1373 1704 sw
rect 1356 1672 1373 1697
rect 1497 1672 1514 1704
rect 1696 1672 1711 1714
rect 1739 1672 1754 1714
rect 1936 1697 1946 1704
tri 1946 1697 1953 1704 sw
rect 1936 1672 1953 1697
rect 2077 1672 2094 1704
rect 2276 1672 2291 1714
rect 2319 1672 2334 1714
rect 2516 1697 2526 1704
tri 2526 1697 2533 1704 sw
rect 2516 1672 2533 1697
rect 2657 1672 2674 1704
rect 2856 1672 2871 1714
rect 2899 1672 2914 1714
rect 3096 1697 3106 1704
tri 3106 1697 3113 1704 sw
rect 3096 1672 3113 1697
rect 3237 1672 3254 1704
rect 3436 1672 3451 1714
rect 3479 1672 3494 1714
rect 3676 1697 3686 1704
tri 3686 1697 3693 1704 sw
rect 3676 1672 3693 1697
rect 3817 1672 3834 1704
rect 4016 1672 4031 1714
rect 4059 1672 4074 1714
rect 4256 1697 4266 1704
tri 4266 1697 4273 1704 sw
rect 4256 1672 4273 1697
rect 4397 1672 4414 1704
rect 4596 1672 4611 1714
rect 4639 1672 4654 1714
rect 4836 1697 4846 1704
tri 4846 1697 4853 1704 sw
rect 4836 1672 4853 1697
rect 4977 1672 4994 1704
rect 5176 1672 5191 1714
rect 5219 1672 5234 1714
rect 5416 1697 5426 1704
tri 5426 1697 5433 1704 sw
rect 5416 1672 5433 1697
rect 5557 1672 5574 1704
rect 5756 1672 5771 1714
rect 5799 1672 5814 1714
rect 5996 1697 6006 1704
tri 6006 1697 6013 1704 sw
rect 5996 1672 6013 1697
rect 6137 1672 6154 1704
rect 6336 1672 6351 1714
rect 6379 1672 6394 1714
rect 6576 1697 6586 1704
tri 6586 1697 6593 1704 sw
rect 6576 1672 6593 1697
rect 6717 1672 6734 1704
rect 6916 1672 6931 1714
rect 259 1634 291 1648
rect 839 1634 871 1648
rect 1419 1634 1451 1648
rect 1999 1634 2031 1648
rect 2579 1634 2611 1648
rect 3159 1634 3191 1648
rect 3739 1634 3771 1648
rect 4319 1634 4351 1648
rect 4899 1634 4931 1648
rect 5479 1634 5511 1648
rect 6059 1634 6091 1648
rect 6639 1634 6671 1648
rect 73 1548 88 1576
rect 154 1548 169 1576
rect 381 1548 396 1576
rect 463 1548 478 1577
rect 653 1548 668 1576
rect 734 1548 749 1576
rect 961 1548 976 1576
rect 1043 1548 1058 1577
rect 1233 1548 1248 1576
rect 1314 1548 1329 1576
rect 1541 1548 1556 1576
rect 1623 1548 1638 1577
rect 1813 1548 1828 1576
rect 1894 1548 1909 1576
rect 2121 1548 2136 1576
rect 2203 1548 2218 1577
rect 2393 1548 2408 1576
rect 2474 1548 2489 1576
rect 2701 1548 2716 1576
rect 2783 1548 2798 1577
rect 2973 1548 2988 1576
rect 3054 1548 3069 1576
rect 3281 1548 3296 1576
rect 3363 1548 3378 1577
rect 3553 1548 3568 1576
rect 3634 1548 3649 1576
rect 3861 1548 3876 1576
rect 3943 1548 3958 1577
rect 4133 1548 4148 1576
rect 4214 1548 4229 1576
rect 4441 1548 4456 1576
rect 4523 1548 4538 1577
rect 4713 1548 4728 1576
rect 4794 1548 4809 1576
rect 5021 1548 5036 1576
rect 5103 1548 5118 1577
rect 5293 1548 5308 1576
rect 5374 1548 5389 1576
rect 5601 1548 5616 1576
rect 5683 1548 5698 1577
rect 5873 1548 5888 1576
rect 5954 1548 5969 1576
rect 6181 1548 6196 1576
rect 6263 1548 6278 1577
rect 6453 1548 6468 1576
rect 6534 1548 6549 1576
rect 6761 1548 6776 1576
rect 6843 1548 6858 1577
rect -1 1402 14 1444
rect 196 1427 206 1434
tri 206 1427 213 1434 sw
rect 196 1402 213 1427
rect 337 1402 354 1434
rect 536 1402 551 1444
rect 579 1402 594 1444
rect 776 1427 786 1434
tri 786 1427 793 1434 sw
rect 776 1402 793 1427
rect 917 1402 934 1434
rect 1116 1402 1131 1444
rect 1159 1402 1174 1444
rect 1356 1427 1366 1434
tri 1366 1427 1373 1434 sw
rect 1356 1402 1373 1427
rect 1497 1402 1514 1434
rect 1696 1402 1711 1444
rect 1739 1402 1754 1444
rect 1936 1427 1946 1434
tri 1946 1427 1953 1434 sw
rect 1936 1402 1953 1427
rect 2077 1402 2094 1434
rect 2276 1402 2291 1444
rect 2319 1402 2334 1444
rect 2516 1427 2526 1434
tri 2526 1427 2533 1434 sw
rect 2516 1402 2533 1427
rect 2657 1402 2674 1434
rect 2856 1402 2871 1444
rect 2899 1402 2914 1444
rect 3096 1427 3106 1434
tri 3106 1427 3113 1434 sw
rect 3096 1402 3113 1427
rect 3237 1402 3254 1434
rect 3436 1402 3451 1444
rect 3479 1402 3494 1444
rect 3676 1427 3686 1434
tri 3686 1427 3693 1434 sw
rect 3676 1402 3693 1427
rect 3817 1402 3834 1434
rect 4016 1402 4031 1444
rect 4059 1402 4074 1444
rect 4256 1427 4266 1434
tri 4266 1427 4273 1434 sw
rect 4256 1402 4273 1427
rect 4397 1402 4414 1434
rect 4596 1402 4611 1444
rect 4639 1402 4654 1444
rect 4836 1427 4846 1434
tri 4846 1427 4853 1434 sw
rect 4836 1402 4853 1427
rect 4977 1402 4994 1434
rect 5176 1402 5191 1444
rect 5219 1402 5234 1444
rect 5416 1427 5426 1434
tri 5426 1427 5433 1434 sw
rect 5416 1402 5433 1427
rect 5557 1402 5574 1434
rect 5756 1402 5771 1444
rect 5799 1402 5814 1444
rect 5996 1427 6006 1434
tri 6006 1427 6013 1434 sw
rect 5996 1402 6013 1427
rect 6137 1402 6154 1434
rect 6336 1402 6351 1444
rect 6379 1402 6394 1444
rect 6576 1427 6586 1434
tri 6586 1427 6593 1434 sw
rect 6576 1402 6593 1427
rect 6717 1402 6734 1434
rect 6916 1402 6931 1444
rect 259 1364 291 1378
rect 839 1364 871 1378
rect 1419 1364 1451 1378
rect 1999 1364 2031 1378
rect 2579 1364 2611 1378
rect 3159 1364 3191 1378
rect 3739 1364 3771 1378
rect 4319 1364 4351 1378
rect 4899 1364 4931 1378
rect 5479 1364 5511 1378
rect 6059 1364 6091 1378
rect 6639 1364 6671 1378
rect 73 1278 88 1306
rect 154 1278 169 1306
rect 381 1278 396 1306
rect 463 1278 478 1307
rect 653 1278 668 1306
rect 734 1278 749 1306
rect 961 1278 976 1306
rect 1043 1278 1058 1307
rect 1233 1278 1248 1306
rect 1314 1278 1329 1306
rect 1541 1278 1556 1306
rect 1623 1278 1638 1307
rect 1813 1278 1828 1306
rect 1894 1278 1909 1306
rect 2121 1278 2136 1306
rect 2203 1278 2218 1307
rect 2393 1278 2408 1306
rect 2474 1278 2489 1306
rect 2701 1278 2716 1306
rect 2783 1278 2798 1307
rect 2973 1278 2988 1306
rect 3054 1278 3069 1306
rect 3281 1278 3296 1306
rect 3363 1278 3378 1307
rect 3553 1278 3568 1306
rect 3634 1278 3649 1306
rect 3861 1278 3876 1306
rect 3943 1278 3958 1307
rect 4133 1278 4148 1306
rect 4214 1278 4229 1306
rect 4441 1278 4456 1306
rect 4523 1278 4538 1307
rect 4713 1278 4728 1306
rect 4794 1278 4809 1306
rect 5021 1278 5036 1306
rect 5103 1278 5118 1307
rect 5293 1278 5308 1306
rect 5374 1278 5389 1306
rect 5601 1278 5616 1306
rect 5683 1278 5698 1307
rect 5873 1278 5888 1306
rect 5954 1278 5969 1306
rect 6181 1278 6196 1306
rect 6263 1278 6278 1307
rect 6453 1278 6468 1306
rect 6534 1278 6549 1306
rect 6761 1278 6776 1306
rect 6843 1278 6858 1307
rect -1 1132 14 1174
rect 196 1157 206 1164
tri 206 1157 213 1164 sw
rect 196 1132 213 1157
rect 337 1132 354 1164
rect 536 1132 551 1174
rect 579 1132 594 1174
rect 776 1157 786 1164
tri 786 1157 793 1164 sw
rect 776 1132 793 1157
rect 917 1132 934 1164
rect 1116 1132 1131 1174
rect 1159 1132 1174 1174
rect 1356 1157 1366 1164
tri 1366 1157 1373 1164 sw
rect 1356 1132 1373 1157
rect 1497 1132 1514 1164
rect 1696 1132 1711 1174
rect 1739 1132 1754 1174
rect 1936 1157 1946 1164
tri 1946 1157 1953 1164 sw
rect 1936 1132 1953 1157
rect 2077 1132 2094 1164
rect 2276 1132 2291 1174
rect 2319 1132 2334 1174
rect 2516 1157 2526 1164
tri 2526 1157 2533 1164 sw
rect 2516 1132 2533 1157
rect 2657 1132 2674 1164
rect 2856 1132 2871 1174
rect 2899 1132 2914 1174
rect 3096 1157 3106 1164
tri 3106 1157 3113 1164 sw
rect 3096 1132 3113 1157
rect 3237 1132 3254 1164
rect 3436 1132 3451 1174
rect 3479 1132 3494 1174
rect 3676 1157 3686 1164
tri 3686 1157 3693 1164 sw
rect 3676 1132 3693 1157
rect 3817 1132 3834 1164
rect 4016 1132 4031 1174
rect 4059 1132 4074 1174
rect 4256 1157 4266 1164
tri 4266 1157 4273 1164 sw
rect 4256 1132 4273 1157
rect 4397 1132 4414 1164
rect 4596 1132 4611 1174
rect 4639 1132 4654 1174
rect 4836 1157 4846 1164
tri 4846 1157 4853 1164 sw
rect 4836 1132 4853 1157
rect 4977 1132 4994 1164
rect 5176 1132 5191 1174
rect 5219 1132 5234 1174
rect 5416 1157 5426 1164
tri 5426 1157 5433 1164 sw
rect 5416 1132 5433 1157
rect 5557 1132 5574 1164
rect 5756 1132 5771 1174
rect 5799 1132 5814 1174
rect 5996 1157 6006 1164
tri 6006 1157 6013 1164 sw
rect 5996 1132 6013 1157
rect 6137 1132 6154 1164
rect 6336 1132 6351 1174
rect 6379 1132 6394 1174
rect 6576 1157 6586 1164
tri 6586 1157 6593 1164 sw
rect 6576 1132 6593 1157
rect 6717 1132 6734 1164
rect 6916 1132 6931 1174
rect 259 1094 291 1108
rect 839 1094 871 1108
rect 1419 1094 1451 1108
rect 1999 1094 2031 1108
rect 2579 1094 2611 1108
rect 3159 1094 3191 1108
rect 3739 1094 3771 1108
rect 4319 1094 4351 1108
rect 4899 1094 4931 1108
rect 5479 1094 5511 1108
rect 6059 1094 6091 1108
rect 6639 1094 6671 1108
rect 73 1008 88 1036
rect 154 1008 169 1036
rect 381 1008 396 1036
rect 463 1008 478 1037
rect 653 1008 668 1036
rect 734 1008 749 1036
rect 961 1008 976 1036
rect 1043 1008 1058 1037
rect 1233 1008 1248 1036
rect 1314 1008 1329 1036
rect 1541 1008 1556 1036
rect 1623 1008 1638 1037
rect 1813 1008 1828 1036
rect 1894 1008 1909 1036
rect 2121 1008 2136 1036
rect 2203 1008 2218 1037
rect 2393 1008 2408 1036
rect 2474 1008 2489 1036
rect 2701 1008 2716 1036
rect 2783 1008 2798 1037
rect 2973 1008 2988 1036
rect 3054 1008 3069 1036
rect 3281 1008 3296 1036
rect 3363 1008 3378 1037
rect 3553 1008 3568 1036
rect 3634 1008 3649 1036
rect 3861 1008 3876 1036
rect 3943 1008 3958 1037
rect 4133 1008 4148 1036
rect 4214 1008 4229 1036
rect 4441 1008 4456 1036
rect 4523 1008 4538 1037
rect 4713 1008 4728 1036
rect 4794 1008 4809 1036
rect 5021 1008 5036 1036
rect 5103 1008 5118 1037
rect 5293 1008 5308 1036
rect 5374 1008 5389 1036
rect 5601 1008 5616 1036
rect 5683 1008 5698 1037
rect 5873 1008 5888 1036
rect 5954 1008 5969 1036
rect 6181 1008 6196 1036
rect 6263 1008 6278 1037
rect 6453 1008 6468 1036
rect 6534 1008 6549 1036
rect 6761 1008 6776 1036
rect 6843 1008 6858 1037
rect -1 862 14 904
rect 196 887 206 894
tri 206 887 213 894 sw
rect 196 862 213 887
rect 337 862 354 894
rect 536 862 551 904
rect 579 862 594 904
rect 776 887 786 894
tri 786 887 793 894 sw
rect 776 862 793 887
rect 917 862 934 894
rect 1116 862 1131 904
rect 1159 862 1174 904
rect 1356 887 1366 894
tri 1366 887 1373 894 sw
rect 1356 862 1373 887
rect 1497 862 1514 894
rect 1696 862 1711 904
rect 1739 862 1754 904
rect 1936 887 1946 894
tri 1946 887 1953 894 sw
rect 1936 862 1953 887
rect 2077 862 2094 894
rect 2276 862 2291 904
rect 2319 862 2334 904
rect 2516 887 2526 894
tri 2526 887 2533 894 sw
rect 2516 862 2533 887
rect 2657 862 2674 894
rect 2856 862 2871 904
rect 2899 862 2914 904
rect 3096 887 3106 894
tri 3106 887 3113 894 sw
rect 3096 862 3113 887
rect 3237 862 3254 894
rect 3436 862 3451 904
rect 3479 862 3494 904
rect 3676 887 3686 894
tri 3686 887 3693 894 sw
rect 3676 862 3693 887
rect 3817 862 3834 894
rect 4016 862 4031 904
rect 4059 862 4074 904
rect 4256 887 4266 894
tri 4266 887 4273 894 sw
rect 4256 862 4273 887
rect 4397 862 4414 894
rect 4596 862 4611 904
rect 4639 862 4654 904
rect 4836 887 4846 894
tri 4846 887 4853 894 sw
rect 4836 862 4853 887
rect 4977 862 4994 894
rect 5176 862 5191 904
rect 5219 862 5234 904
rect 5416 887 5426 894
tri 5426 887 5433 894 sw
rect 5416 862 5433 887
rect 5557 862 5574 894
rect 5756 862 5771 904
rect 5799 862 5814 904
rect 5996 887 6006 894
tri 6006 887 6013 894 sw
rect 5996 862 6013 887
rect 6137 862 6154 894
rect 6336 862 6351 904
rect 6379 862 6394 904
rect 6576 887 6586 894
tri 6586 887 6593 894 sw
rect 6576 862 6593 887
rect 6717 862 6734 894
rect 6916 862 6931 904
rect 259 824 291 838
rect 839 824 871 838
rect 1419 824 1451 838
rect 1999 824 2031 838
rect 2579 824 2611 838
rect 3159 824 3191 838
rect 3739 824 3771 838
rect 4319 824 4351 838
rect 4899 824 4931 838
rect 5479 824 5511 838
rect 6059 824 6091 838
rect 6639 824 6671 838
rect 73 738 88 766
rect 154 738 169 766
rect 381 738 396 766
rect 463 738 478 767
rect 653 738 668 766
rect 734 738 749 766
rect 961 738 976 766
rect 1043 738 1058 767
rect 1233 738 1248 766
rect 1314 738 1329 766
rect 1541 738 1556 766
rect 1623 738 1638 767
rect 1813 738 1828 766
rect 1894 738 1909 766
rect 2121 738 2136 766
rect 2203 738 2218 767
rect 2393 738 2408 766
rect 2474 738 2489 766
rect 2701 738 2716 766
rect 2783 738 2798 767
rect 2973 738 2988 766
rect 3054 738 3069 766
rect 3281 738 3296 766
rect 3363 738 3378 767
rect 3553 738 3568 766
rect 3634 738 3649 766
rect 3861 738 3876 766
rect 3943 738 3958 767
rect 4133 738 4148 766
rect 4214 738 4229 766
rect 4441 738 4456 766
rect 4523 738 4538 767
rect 4713 738 4728 766
rect 4794 738 4809 766
rect 5021 738 5036 766
rect 5103 738 5118 767
rect 5293 738 5308 766
rect 5374 738 5389 766
rect 5601 738 5616 766
rect 5683 738 5698 767
rect 5873 738 5888 766
rect 5954 738 5969 766
rect 6181 738 6196 766
rect 6263 738 6278 767
rect 6453 738 6468 766
rect 6534 738 6549 766
rect 6761 738 6776 766
rect 6843 738 6858 767
rect -1 592 14 634
rect 196 617 206 624
tri 206 617 213 624 sw
rect 196 592 213 617
rect 337 592 354 624
rect 536 592 551 634
rect 579 592 594 634
rect 776 617 786 624
tri 786 617 793 624 sw
rect 776 592 793 617
rect 917 592 934 624
rect 1116 592 1131 634
rect 1159 592 1174 634
rect 1356 617 1366 624
tri 1366 617 1373 624 sw
rect 1356 592 1373 617
rect 1497 592 1514 624
rect 1696 592 1711 634
rect 1739 592 1754 634
rect 1936 617 1946 624
tri 1946 617 1953 624 sw
rect 1936 592 1953 617
rect 2077 592 2094 624
rect 2276 592 2291 634
rect 2319 592 2334 634
rect 2516 617 2526 624
tri 2526 617 2533 624 sw
rect 2516 592 2533 617
rect 2657 592 2674 624
rect 2856 592 2871 634
rect 2899 592 2914 634
rect 3096 617 3106 624
tri 3106 617 3113 624 sw
rect 3096 592 3113 617
rect 3237 592 3254 624
rect 3436 592 3451 634
rect 3479 592 3494 634
rect 3676 617 3686 624
tri 3686 617 3693 624 sw
rect 3676 592 3693 617
rect 3817 592 3834 624
rect 4016 592 4031 634
rect 4059 592 4074 634
rect 4256 617 4266 624
tri 4266 617 4273 624 sw
rect 4256 592 4273 617
rect 4397 592 4414 624
rect 4596 592 4611 634
rect 4639 592 4654 634
rect 4836 617 4846 624
tri 4846 617 4853 624 sw
rect 4836 592 4853 617
rect 4977 592 4994 624
rect 5176 592 5191 634
rect 5219 592 5234 634
rect 5416 617 5426 624
tri 5426 617 5433 624 sw
rect 5416 592 5433 617
rect 5557 592 5574 624
rect 5756 592 5771 634
rect 5799 592 5814 634
rect 5996 617 6006 624
tri 6006 617 6013 624 sw
rect 5996 592 6013 617
rect 6137 592 6154 624
rect 6336 592 6351 634
rect 6379 592 6394 634
rect 6576 617 6586 624
tri 6586 617 6593 624 sw
rect 6576 592 6593 617
rect 6717 592 6734 624
rect 6916 592 6931 634
rect 259 554 291 568
rect 839 554 871 568
rect 1419 554 1451 568
rect 1999 554 2031 568
rect 2579 554 2611 568
rect 3159 554 3191 568
rect 3739 554 3771 568
rect 4319 554 4351 568
rect 4899 554 4931 568
rect 5479 554 5511 568
rect 6059 554 6091 568
rect 6639 554 6671 568
rect 73 468 88 496
rect 154 468 169 496
rect 381 468 396 496
rect 463 468 478 497
rect 653 468 668 496
rect 734 468 749 496
rect 961 468 976 496
rect 1043 468 1058 497
rect 1233 468 1248 496
rect 1314 468 1329 496
rect 1541 468 1556 496
rect 1623 468 1638 497
rect 1813 468 1828 496
rect 1894 468 1909 496
rect 2121 468 2136 496
rect 2203 468 2218 497
rect 2393 468 2408 496
rect 2474 468 2489 496
rect 2701 468 2716 496
rect 2783 468 2798 497
rect 2973 468 2988 496
rect 3054 468 3069 496
rect 3281 468 3296 496
rect 3363 468 3378 497
rect 3553 468 3568 496
rect 3634 468 3649 496
rect 3861 468 3876 496
rect 3943 468 3958 497
rect 4133 468 4148 496
rect 4214 468 4229 496
rect 4441 468 4456 496
rect 4523 468 4538 497
rect 4713 468 4728 496
rect 4794 468 4809 496
rect 5021 468 5036 496
rect 5103 468 5118 497
rect 5293 468 5308 496
rect 5374 468 5389 496
rect 5601 468 5616 496
rect 5683 468 5698 497
rect 5873 468 5888 496
rect 5954 468 5969 496
rect 6181 468 6196 496
rect 6263 468 6278 497
rect 6453 468 6468 496
rect 6534 468 6549 496
rect 6761 468 6776 496
rect 6843 468 6858 497
rect -1 322 14 364
rect 196 347 206 354
tri 206 347 213 354 sw
rect 196 322 213 347
rect 337 322 354 354
rect 536 322 551 364
rect 579 322 594 364
rect 776 347 786 354
tri 786 347 793 354 sw
rect 776 322 793 347
rect 917 322 934 354
rect 1116 322 1131 364
rect 1159 322 1174 364
rect 1356 347 1366 354
tri 1366 347 1373 354 sw
rect 1356 322 1373 347
rect 1497 322 1514 354
rect 1696 322 1711 364
rect 1739 322 1754 364
rect 1936 347 1946 354
tri 1946 347 1953 354 sw
rect 1936 322 1953 347
rect 2077 322 2094 354
rect 2276 322 2291 364
rect 2319 322 2334 364
rect 2516 347 2526 354
tri 2526 347 2533 354 sw
rect 2516 322 2533 347
rect 2657 322 2674 354
rect 2856 322 2871 364
rect 2899 322 2914 364
rect 3096 347 3106 354
tri 3106 347 3113 354 sw
rect 3096 322 3113 347
rect 3237 322 3254 354
rect 3436 322 3451 364
rect 3479 322 3494 364
rect 3676 347 3686 354
tri 3686 347 3693 354 sw
rect 3676 322 3693 347
rect 3817 322 3834 354
rect 4016 322 4031 364
rect 4059 322 4074 364
rect 4256 347 4266 354
tri 4266 347 4273 354 sw
rect 4256 322 4273 347
rect 4397 322 4414 354
rect 4596 322 4611 364
rect 4639 322 4654 364
rect 4836 347 4846 354
tri 4846 347 4853 354 sw
rect 4836 322 4853 347
rect 4977 322 4994 354
rect 5176 322 5191 364
rect 5219 322 5234 364
rect 5416 347 5426 354
tri 5426 347 5433 354 sw
rect 5416 322 5433 347
rect 5557 322 5574 354
rect 5756 322 5771 364
rect 5799 322 5814 364
rect 5996 347 6006 354
tri 6006 347 6013 354 sw
rect 5996 322 6013 347
rect 6137 322 6154 354
rect 6336 322 6351 364
rect 6379 322 6394 364
rect 6576 347 6586 354
tri 6586 347 6593 354 sw
rect 6576 322 6593 347
rect 6717 322 6734 354
rect 6916 322 6931 364
rect 259 284 291 298
rect 839 284 871 298
rect 1419 284 1451 298
rect 1999 284 2031 298
rect 2579 284 2611 298
rect 3159 284 3191 298
rect 3739 284 3771 298
rect 4319 284 4351 298
rect 4899 284 4931 298
rect 5479 284 5511 298
rect 6059 284 6091 298
rect 6639 284 6671 298
rect 73 198 88 226
rect 154 198 169 226
rect 381 198 396 226
rect 463 198 478 227
rect 653 198 668 226
rect 734 198 749 226
rect 961 198 976 226
rect 1043 198 1058 227
rect 1233 198 1248 226
rect 1314 198 1329 226
rect 1541 198 1556 226
rect 1623 198 1638 227
rect 1813 198 1828 226
rect 1894 198 1909 226
rect 2121 198 2136 226
rect 2203 198 2218 227
rect 2393 198 2408 226
rect 2474 198 2489 226
rect 2701 198 2716 226
rect 2783 198 2798 227
rect 2973 198 2988 226
rect 3054 198 3069 226
rect 3281 198 3296 226
rect 3363 198 3378 227
rect 3553 198 3568 226
rect 3634 198 3649 226
rect 3861 198 3876 226
rect 3943 198 3958 227
rect 4133 198 4148 226
rect 4214 198 4229 226
rect 4441 198 4456 226
rect 4523 198 4538 227
rect 4713 198 4728 226
rect 4794 198 4809 226
rect 5021 198 5036 226
rect 5103 198 5118 227
rect 5293 198 5308 226
rect 5374 198 5389 226
rect 5601 198 5616 226
rect 5683 198 5698 227
rect 5873 198 5888 226
rect 5954 198 5969 226
rect 6181 198 6196 226
rect 6263 198 6278 227
rect 6453 198 6468 226
rect 6534 198 6549 226
rect 6761 198 6776 226
rect 6843 198 6858 227
rect -1 52 14 94
rect 196 77 206 84
tri 206 77 213 84 sw
rect 196 52 213 77
rect 337 52 354 84
rect 536 52 551 94
rect 579 52 594 94
rect 776 77 786 84
tri 786 77 793 84 sw
rect 776 52 793 77
rect 917 52 934 84
rect 1116 52 1131 94
rect 1159 52 1174 94
rect 1356 77 1366 84
tri 1366 77 1373 84 sw
rect 1356 52 1373 77
rect 1497 52 1514 84
rect 1696 52 1711 94
rect 1739 52 1754 94
rect 1936 77 1946 84
tri 1946 77 1953 84 sw
rect 1936 52 1953 77
rect 2077 52 2094 84
rect 2276 52 2291 94
rect 2319 52 2334 94
rect 2516 77 2526 84
tri 2526 77 2533 84 sw
rect 2516 52 2533 77
rect 2657 52 2674 84
rect 2856 52 2871 94
rect 2899 52 2914 94
rect 3096 77 3106 84
tri 3106 77 3113 84 sw
rect 3096 52 3113 77
rect 3237 52 3254 84
rect 3436 52 3451 94
rect 3479 52 3494 94
rect 3676 77 3686 84
tri 3686 77 3693 84 sw
rect 3676 52 3693 77
rect 3817 52 3834 84
rect 4016 52 4031 94
rect 4059 52 4074 94
rect 4256 77 4266 84
tri 4266 77 4273 84 sw
rect 4256 52 4273 77
rect 4397 52 4414 84
rect 4596 52 4611 94
rect 4639 52 4654 94
rect 4836 77 4846 84
tri 4846 77 4853 84 sw
rect 4836 52 4853 77
rect 4977 52 4994 84
rect 5176 52 5191 94
rect 5219 52 5234 94
rect 5416 77 5426 84
tri 5426 77 5433 84 sw
rect 5416 52 5433 77
rect 5557 52 5574 84
rect 5756 52 5771 94
rect 5799 52 5814 94
rect 5996 77 6006 84
tri 6006 77 6013 84 sw
rect 5996 52 6013 77
rect 6137 52 6154 84
rect 6336 52 6351 94
rect 6379 52 6394 94
rect 6576 77 6586 84
tri 6586 77 6593 84 sw
rect 6576 52 6593 77
rect 6717 52 6734 84
rect 6916 52 6931 94
rect 259 14 291 28
rect 839 14 871 28
rect 1419 14 1451 28
rect 1999 14 2031 28
rect 2579 14 2611 28
rect 3159 14 3191 28
rect 3739 14 3771 28
rect 4319 14 4351 28
rect 4899 14 4931 28
rect 5479 14 5511 28
rect 6059 14 6091 28
rect 6639 14 6671 28
rect 73 -72 88 -44
rect 154 -72 169 -44
rect 381 -72 396 -44
rect 463 -72 478 -43
rect 653 -72 668 -44
rect 734 -72 749 -44
rect 961 -72 976 -44
rect 1043 -72 1058 -43
rect 1233 -72 1248 -44
rect 1314 -72 1329 -44
rect 1541 -72 1556 -44
rect 1623 -72 1638 -43
rect 1813 -72 1828 -44
rect 1894 -72 1909 -44
rect 2121 -72 2136 -44
rect 2203 -72 2218 -43
rect 2393 -72 2408 -44
rect 2474 -72 2489 -44
rect 2701 -72 2716 -44
rect 2783 -72 2798 -43
rect 2973 -72 2988 -44
rect 3054 -72 3069 -44
rect 3281 -72 3296 -44
rect 3363 -72 3378 -43
rect 3553 -72 3568 -44
rect 3634 -72 3649 -44
rect 3861 -72 3876 -44
rect 3943 -72 3958 -43
rect 4133 -72 4148 -44
rect 4214 -72 4229 -44
rect 4441 -72 4456 -44
rect 4523 -72 4538 -43
rect 4713 -72 4728 -44
rect 4794 -72 4809 -44
rect 5021 -72 5036 -44
rect 5103 -72 5118 -43
rect 5293 -72 5308 -44
rect 5374 -72 5389 -44
rect 5601 -72 5616 -44
rect 5683 -72 5698 -43
rect 5873 -72 5888 -44
rect 5954 -72 5969 -44
rect 6181 -72 6196 -44
rect 6263 -72 6278 -43
rect 6453 -72 6468 -44
rect 6534 -72 6549 -44
rect 6761 -72 6776 -44
rect 6843 -72 6858 -43
rect -1 -218 14 -176
rect 196 -193 206 -186
tri 206 -193 213 -186 sw
rect 196 -218 213 -193
rect 337 -218 354 -186
rect 536 -218 551 -176
rect 579 -218 594 -176
rect 776 -193 786 -186
tri 786 -193 793 -186 sw
rect 776 -218 793 -193
rect 917 -218 934 -186
rect 1116 -218 1131 -176
rect 1159 -218 1174 -176
rect 1356 -193 1366 -186
tri 1366 -193 1373 -186 sw
rect 1356 -218 1373 -193
rect 1497 -218 1514 -186
rect 1696 -218 1711 -176
rect 1739 -218 1754 -176
rect 1936 -193 1946 -186
tri 1946 -193 1953 -186 sw
rect 1936 -218 1953 -193
rect 2077 -218 2094 -186
rect 2276 -218 2291 -176
rect 2319 -218 2334 -176
rect 2516 -193 2526 -186
tri 2526 -193 2533 -186 sw
rect 2516 -218 2533 -193
rect 2657 -218 2674 -186
rect 2856 -218 2871 -176
rect 2899 -218 2914 -176
rect 3096 -193 3106 -186
tri 3106 -193 3113 -186 sw
rect 3096 -218 3113 -193
rect 3237 -218 3254 -186
rect 3436 -218 3451 -176
rect 3479 -218 3494 -176
rect 3676 -193 3686 -186
tri 3686 -193 3693 -186 sw
rect 3676 -218 3693 -193
rect 3817 -218 3834 -186
rect 4016 -218 4031 -176
rect 4059 -218 4074 -176
rect 4256 -193 4266 -186
tri 4266 -193 4273 -186 sw
rect 4256 -218 4273 -193
rect 4397 -218 4414 -186
rect 4596 -218 4611 -176
rect 4639 -218 4654 -176
rect 4836 -193 4846 -186
tri 4846 -193 4853 -186 sw
rect 4836 -218 4853 -193
rect 4977 -218 4994 -186
rect 5176 -218 5191 -176
rect 5219 -218 5234 -176
rect 5416 -193 5426 -186
tri 5426 -193 5433 -186 sw
rect 5416 -218 5433 -193
rect 5557 -218 5574 -186
rect 5756 -218 5771 -176
rect 5799 -218 5814 -176
rect 5996 -193 6006 -186
tri 6006 -193 6013 -186 sw
rect 5996 -218 6013 -193
rect 6137 -218 6154 -186
rect 6336 -218 6351 -176
rect 6379 -218 6394 -176
rect 6576 -193 6586 -186
tri 6586 -193 6593 -186 sw
rect 6576 -218 6593 -193
rect 6717 -218 6734 -186
rect 6916 -218 6931 -176
rect 259 -256 291 -242
rect 839 -256 871 -242
rect 1419 -256 1451 -242
rect 1999 -256 2031 -242
rect 2579 -256 2611 -242
rect 3159 -256 3191 -242
rect 3739 -256 3771 -242
rect 4319 -256 4351 -242
rect 4899 -256 4931 -242
rect 5479 -256 5511 -242
rect 6059 -256 6091 -242
rect 6639 -256 6671 -242
rect 73 -342 88 -314
rect 154 -342 169 -314
rect 381 -342 396 -314
rect 463 -342 478 -313
rect 653 -342 668 -314
rect 734 -342 749 -314
rect 961 -342 976 -314
rect 1043 -342 1058 -313
rect 1233 -342 1248 -314
rect 1314 -342 1329 -314
rect 1541 -342 1556 -314
rect 1623 -342 1638 -313
rect 1813 -342 1828 -314
rect 1894 -342 1909 -314
rect 2121 -342 2136 -314
rect 2203 -342 2218 -313
rect 2393 -342 2408 -314
rect 2474 -342 2489 -314
rect 2701 -342 2716 -314
rect 2783 -342 2798 -313
rect 2973 -342 2988 -314
rect 3054 -342 3069 -314
rect 3281 -342 3296 -314
rect 3363 -342 3378 -313
rect 3553 -342 3568 -314
rect 3634 -342 3649 -314
rect 3861 -342 3876 -314
rect 3943 -342 3958 -313
rect 4133 -342 4148 -314
rect 4214 -342 4229 -314
rect 4441 -342 4456 -314
rect 4523 -342 4538 -313
rect 4713 -342 4728 -314
rect 4794 -342 4809 -314
rect 5021 -342 5036 -314
rect 5103 -342 5118 -313
rect 5293 -342 5308 -314
rect 5374 -342 5389 -314
rect 5601 -342 5616 -314
rect 5683 -342 5698 -313
rect 5873 -342 5888 -314
rect 5954 -342 5969 -314
rect 6181 -342 6196 -314
rect 6263 -342 6278 -313
rect 6453 -342 6468 -314
rect 6534 -342 6549 -314
rect 6761 -342 6776 -314
rect 6843 -342 6858 -313
rect -1 -488 14 -446
rect 196 -463 206 -456
tri 206 -463 213 -456 sw
rect 196 -488 213 -463
rect 337 -488 354 -456
rect 536 -488 551 -446
rect 579 -488 594 -446
rect 776 -463 786 -456
tri 786 -463 793 -456 sw
rect 776 -488 793 -463
rect 917 -488 934 -456
rect 1116 -488 1131 -446
rect 1159 -488 1174 -446
rect 1356 -463 1366 -456
tri 1366 -463 1373 -456 sw
rect 1356 -488 1373 -463
rect 1497 -488 1514 -456
rect 1696 -488 1711 -446
rect 1739 -488 1754 -446
rect 1936 -463 1946 -456
tri 1946 -463 1953 -456 sw
rect 1936 -488 1953 -463
rect 2077 -488 2094 -456
rect 2276 -488 2291 -446
rect 2319 -488 2334 -446
rect 2516 -463 2526 -456
tri 2526 -463 2533 -456 sw
rect 2516 -488 2533 -463
rect 2657 -488 2674 -456
rect 2856 -488 2871 -446
rect 2899 -488 2914 -446
rect 3096 -463 3106 -456
tri 3106 -463 3113 -456 sw
rect 3096 -488 3113 -463
rect 3237 -488 3254 -456
rect 3436 -488 3451 -446
rect 3479 -488 3494 -446
rect 3676 -463 3686 -456
tri 3686 -463 3693 -456 sw
rect 3676 -488 3693 -463
rect 3817 -488 3834 -456
rect 4016 -488 4031 -446
rect 4059 -488 4074 -446
rect 4256 -463 4266 -456
tri 4266 -463 4273 -456 sw
rect 4256 -488 4273 -463
rect 4397 -488 4414 -456
rect 4596 -488 4611 -446
rect 4639 -488 4654 -446
rect 4836 -463 4846 -456
tri 4846 -463 4853 -456 sw
rect 4836 -488 4853 -463
rect 4977 -488 4994 -456
rect 5176 -488 5191 -446
rect 5219 -488 5234 -446
rect 5416 -463 5426 -456
tri 5426 -463 5433 -456 sw
rect 5416 -488 5433 -463
rect 5557 -488 5574 -456
rect 5756 -488 5771 -446
rect 5799 -488 5814 -446
rect 5996 -463 6006 -456
tri 6006 -463 6013 -456 sw
rect 5996 -488 6013 -463
rect 6137 -488 6154 -456
rect 6336 -488 6351 -446
rect 6379 -488 6394 -446
rect 6576 -463 6586 -456
tri 6586 -463 6593 -456 sw
rect 6576 -488 6593 -463
rect 6717 -488 6734 -456
rect 6916 -488 6931 -446
rect 259 -526 291 -512
rect 839 -526 871 -512
rect 1419 -526 1451 -512
rect 1999 -526 2031 -512
rect 2579 -526 2611 -512
rect 3159 -526 3191 -512
rect 3739 -526 3771 -512
rect 4319 -526 4351 -512
rect 4899 -526 4931 -512
rect 5479 -526 5511 -512
rect 6059 -526 6091 -512
rect 6639 -526 6671 -512
rect 73 -612 88 -584
rect 154 -612 169 -584
rect 381 -612 396 -584
rect 463 -612 478 -583
rect 653 -612 668 -584
rect 734 -612 749 -584
rect 961 -612 976 -584
rect 1043 -612 1058 -583
rect 1233 -612 1248 -584
rect 1314 -612 1329 -584
rect 1541 -612 1556 -584
rect 1623 -612 1638 -583
rect 1813 -612 1828 -584
rect 1894 -612 1909 -584
rect 2121 -612 2136 -584
rect 2203 -612 2218 -583
rect 2393 -612 2408 -584
rect 2474 -612 2489 -584
rect 2701 -612 2716 -584
rect 2783 -612 2798 -583
rect 2973 -612 2988 -584
rect 3054 -612 3069 -584
rect 3281 -612 3296 -584
rect 3363 -612 3378 -583
rect 3553 -612 3568 -584
rect 3634 -612 3649 -584
rect 3861 -612 3876 -584
rect 3943 -612 3958 -583
rect 4133 -612 4148 -584
rect 4214 -612 4229 -584
rect 4441 -612 4456 -584
rect 4523 -612 4538 -583
rect 4713 -612 4728 -584
rect 4794 -612 4809 -584
rect 5021 -612 5036 -584
rect 5103 -612 5118 -583
rect 5293 -612 5308 -584
rect 5374 -612 5389 -584
rect 5601 -612 5616 -584
rect 5683 -612 5698 -583
rect 5873 -612 5888 -584
rect 5954 -612 5969 -584
rect 6181 -612 6196 -584
rect 6263 -612 6278 -583
rect 6453 -612 6468 -584
rect 6534 -612 6549 -584
rect 6761 -612 6776 -584
rect 6843 -612 6858 -583
rect -1 -758 14 -716
rect 196 -733 206 -726
tri 206 -733 213 -726 sw
rect 196 -758 213 -733
rect 337 -758 354 -726
rect 536 -758 551 -716
rect 579 -758 594 -716
rect 776 -733 786 -726
tri 786 -733 793 -726 sw
rect 776 -758 793 -733
rect 917 -758 934 -726
rect 1116 -758 1131 -716
rect 1159 -758 1174 -716
rect 1356 -733 1366 -726
tri 1366 -733 1373 -726 sw
rect 1356 -758 1373 -733
rect 1497 -758 1514 -726
rect 1696 -758 1711 -716
rect 1739 -758 1754 -716
rect 1936 -733 1946 -726
tri 1946 -733 1953 -726 sw
rect 1936 -758 1953 -733
rect 2077 -758 2094 -726
rect 2276 -758 2291 -716
rect 2319 -758 2334 -716
rect 2516 -733 2526 -726
tri 2526 -733 2533 -726 sw
rect 2516 -758 2533 -733
rect 2657 -758 2674 -726
rect 2856 -758 2871 -716
rect 2899 -758 2914 -716
rect 3096 -733 3106 -726
tri 3106 -733 3113 -726 sw
rect 3096 -758 3113 -733
rect 3237 -758 3254 -726
rect 3436 -758 3451 -716
rect 3479 -758 3494 -716
rect 3676 -733 3686 -726
tri 3686 -733 3693 -726 sw
rect 3676 -758 3693 -733
rect 3817 -758 3834 -726
rect 4016 -758 4031 -716
rect 4059 -758 4074 -716
rect 4256 -733 4266 -726
tri 4266 -733 4273 -726 sw
rect 4256 -758 4273 -733
rect 4397 -758 4414 -726
rect 4596 -758 4611 -716
rect 4639 -758 4654 -716
rect 4836 -733 4846 -726
tri 4846 -733 4853 -726 sw
rect 4836 -758 4853 -733
rect 4977 -758 4994 -726
rect 5176 -758 5191 -716
rect 5219 -758 5234 -716
rect 5416 -733 5426 -726
tri 5426 -733 5433 -726 sw
rect 5416 -758 5433 -733
rect 5557 -758 5574 -726
rect 5756 -758 5771 -716
rect 5799 -758 5814 -716
rect 5996 -733 6006 -726
tri 6006 -733 6013 -726 sw
rect 5996 -758 6013 -733
rect 6137 -758 6154 -726
rect 6336 -758 6351 -716
rect 6379 -758 6394 -716
rect 6576 -733 6586 -726
tri 6586 -733 6593 -726 sw
rect 6576 -758 6593 -733
rect 6717 -758 6734 -726
rect 6916 -758 6931 -716
rect 259 -796 291 -782
rect 839 -796 871 -782
rect 1419 -796 1451 -782
rect 1999 -796 2031 -782
rect 2579 -796 2611 -782
rect 3159 -796 3191 -782
rect 3739 -796 3771 -782
rect 4319 -796 4351 -782
rect 4899 -796 4931 -782
rect 5479 -796 5511 -782
rect 6059 -796 6091 -782
rect 6639 -796 6671 -782
rect 73 -882 88 -854
rect 154 -882 169 -854
rect 381 -882 396 -854
rect 463 -882 478 -853
rect 653 -882 668 -854
rect 734 -882 749 -854
rect 961 -882 976 -854
rect 1043 -882 1058 -853
rect 1233 -882 1248 -854
rect 1314 -882 1329 -854
rect 1541 -882 1556 -854
rect 1623 -882 1638 -853
rect 1813 -882 1828 -854
rect 1894 -882 1909 -854
rect 2121 -882 2136 -854
rect 2203 -882 2218 -853
rect 2393 -882 2408 -854
rect 2474 -882 2489 -854
rect 2701 -882 2716 -854
rect 2783 -882 2798 -853
rect 2973 -882 2988 -854
rect 3054 -882 3069 -854
rect 3281 -882 3296 -854
rect 3363 -882 3378 -853
rect 3553 -882 3568 -854
rect 3634 -882 3649 -854
rect 3861 -882 3876 -854
rect 3943 -882 3958 -853
rect 4133 -882 4148 -854
rect 4214 -882 4229 -854
rect 4441 -882 4456 -854
rect 4523 -882 4538 -853
rect 4713 -882 4728 -854
rect 4794 -882 4809 -854
rect 5021 -882 5036 -854
rect 5103 -882 5118 -853
rect 5293 -882 5308 -854
rect 5374 -882 5389 -854
rect 5601 -882 5616 -854
rect 5683 -882 5698 -853
rect 5873 -882 5888 -854
rect 5954 -882 5969 -854
rect 6181 -882 6196 -854
rect 6263 -882 6278 -853
rect 6453 -882 6468 -854
rect 6534 -882 6549 -854
rect 6761 -882 6776 -854
rect 6843 -882 6858 -853
rect -1 -1028 14 -986
rect 196 -1003 206 -996
tri 206 -1003 213 -996 sw
rect 196 -1028 213 -1003
rect 337 -1028 354 -996
rect 536 -1028 551 -986
rect 579 -1028 594 -986
rect 776 -1003 786 -996
tri 786 -1003 793 -996 sw
rect 776 -1028 793 -1003
rect 917 -1028 934 -996
rect 1116 -1028 1131 -986
rect 1159 -1028 1174 -986
rect 1356 -1003 1366 -996
tri 1366 -1003 1373 -996 sw
rect 1356 -1028 1373 -1003
rect 1497 -1028 1514 -996
rect 1696 -1028 1711 -986
rect 1739 -1028 1754 -986
rect 1936 -1003 1946 -996
tri 1946 -1003 1953 -996 sw
rect 1936 -1028 1953 -1003
rect 2077 -1028 2094 -996
rect 2276 -1028 2291 -986
rect 2319 -1028 2334 -986
rect 2516 -1003 2526 -996
tri 2526 -1003 2533 -996 sw
rect 2516 -1028 2533 -1003
rect 2657 -1028 2674 -996
rect 2856 -1028 2871 -986
rect 2899 -1028 2914 -986
rect 3096 -1003 3106 -996
tri 3106 -1003 3113 -996 sw
rect 3096 -1028 3113 -1003
rect 3237 -1028 3254 -996
rect 3436 -1028 3451 -986
rect 3479 -1028 3494 -986
rect 3676 -1003 3686 -996
tri 3686 -1003 3693 -996 sw
rect 3676 -1028 3693 -1003
rect 3817 -1028 3834 -996
rect 4016 -1028 4031 -986
rect 4059 -1028 4074 -986
rect 4256 -1003 4266 -996
tri 4266 -1003 4273 -996 sw
rect 4256 -1028 4273 -1003
rect 4397 -1028 4414 -996
rect 4596 -1028 4611 -986
rect 4639 -1028 4654 -986
rect 4836 -1003 4846 -996
tri 4846 -1003 4853 -996 sw
rect 4836 -1028 4853 -1003
rect 4977 -1028 4994 -996
rect 5176 -1028 5191 -986
rect 5219 -1028 5234 -986
rect 5416 -1003 5426 -996
tri 5426 -1003 5433 -996 sw
rect 5416 -1028 5433 -1003
rect 5557 -1028 5574 -996
rect 5756 -1028 5771 -986
rect 5799 -1028 5814 -986
rect 5996 -1003 6006 -996
tri 6006 -1003 6013 -996 sw
rect 5996 -1028 6013 -1003
rect 6137 -1028 6154 -996
rect 6336 -1028 6351 -986
rect 6379 -1028 6394 -986
rect 6576 -1003 6586 -996
tri 6586 -1003 6593 -996 sw
rect 6576 -1028 6593 -1003
rect 6717 -1028 6734 -996
rect 6916 -1028 6931 -986
rect 259 -1066 291 -1052
rect 839 -1066 871 -1052
rect 1419 -1066 1451 -1052
rect 1999 -1066 2031 -1052
rect 2579 -1066 2611 -1052
rect 3159 -1066 3191 -1052
rect 3739 -1066 3771 -1052
rect 4319 -1066 4351 -1052
rect 4899 -1066 4931 -1052
rect 5479 -1066 5511 -1052
rect 6059 -1066 6091 -1052
rect 6639 -1066 6671 -1052
rect 73 -1152 88 -1124
rect 154 -1152 169 -1124
rect 381 -1152 396 -1124
rect 463 -1152 478 -1123
rect 653 -1152 668 -1124
rect 734 -1152 749 -1124
rect 961 -1152 976 -1124
rect 1043 -1152 1058 -1123
rect 1233 -1152 1248 -1124
rect 1314 -1152 1329 -1124
rect 1541 -1152 1556 -1124
rect 1623 -1152 1638 -1123
rect 1813 -1152 1828 -1124
rect 1894 -1152 1909 -1124
rect 2121 -1152 2136 -1124
rect 2203 -1152 2218 -1123
rect 2393 -1152 2408 -1124
rect 2474 -1152 2489 -1124
rect 2701 -1152 2716 -1124
rect 2783 -1152 2798 -1123
rect 2973 -1152 2988 -1124
rect 3054 -1152 3069 -1124
rect 3281 -1152 3296 -1124
rect 3363 -1152 3378 -1123
rect 3553 -1152 3568 -1124
rect 3634 -1152 3649 -1124
rect 3861 -1152 3876 -1124
rect 3943 -1152 3958 -1123
rect 4133 -1152 4148 -1124
rect 4214 -1152 4229 -1124
rect 4441 -1152 4456 -1124
rect 4523 -1152 4538 -1123
rect 4713 -1152 4728 -1124
rect 4794 -1152 4809 -1124
rect 5021 -1152 5036 -1124
rect 5103 -1152 5118 -1123
rect 5293 -1152 5308 -1124
rect 5374 -1152 5389 -1124
rect 5601 -1152 5616 -1124
rect 5683 -1152 5698 -1123
rect 5873 -1152 5888 -1124
rect 5954 -1152 5969 -1124
rect 6181 -1152 6196 -1124
rect 6263 -1152 6278 -1123
rect 6453 -1152 6468 -1124
rect 6534 -1152 6549 -1124
rect 6761 -1152 6776 -1124
rect 6843 -1152 6858 -1123
rect -1 -1298 14 -1256
rect 196 -1273 206 -1266
tri 206 -1273 213 -1266 sw
rect 196 -1298 213 -1273
rect 337 -1298 354 -1266
rect 536 -1298 551 -1256
rect 579 -1298 594 -1256
rect 776 -1273 786 -1266
tri 786 -1273 793 -1266 sw
rect 776 -1298 793 -1273
rect 917 -1298 934 -1266
rect 1116 -1298 1131 -1256
rect 1159 -1298 1174 -1256
rect 1356 -1273 1366 -1266
tri 1366 -1273 1373 -1266 sw
rect 1356 -1298 1373 -1273
rect 1497 -1298 1514 -1266
rect 1696 -1298 1711 -1256
rect 1739 -1298 1754 -1256
rect 1936 -1273 1946 -1266
tri 1946 -1273 1953 -1266 sw
rect 1936 -1298 1953 -1273
rect 2077 -1298 2094 -1266
rect 2276 -1298 2291 -1256
rect 2319 -1298 2334 -1256
rect 2516 -1273 2526 -1266
tri 2526 -1273 2533 -1266 sw
rect 2516 -1298 2533 -1273
rect 2657 -1298 2674 -1266
rect 2856 -1298 2871 -1256
rect 2899 -1298 2914 -1256
rect 3096 -1273 3106 -1266
tri 3106 -1273 3113 -1266 sw
rect 3096 -1298 3113 -1273
rect 3237 -1298 3254 -1266
rect 3436 -1298 3451 -1256
rect 3479 -1298 3494 -1256
rect 3676 -1273 3686 -1266
tri 3686 -1273 3693 -1266 sw
rect 3676 -1298 3693 -1273
rect 3817 -1298 3834 -1266
rect 4016 -1298 4031 -1256
rect 4059 -1298 4074 -1256
rect 4256 -1273 4266 -1266
tri 4266 -1273 4273 -1266 sw
rect 4256 -1298 4273 -1273
rect 4397 -1298 4414 -1266
rect 4596 -1298 4611 -1256
rect 4639 -1298 4654 -1256
rect 4836 -1273 4846 -1266
tri 4846 -1273 4853 -1266 sw
rect 4836 -1298 4853 -1273
rect 4977 -1298 4994 -1266
rect 5176 -1298 5191 -1256
rect 5219 -1298 5234 -1256
rect 5416 -1273 5426 -1266
tri 5426 -1273 5433 -1266 sw
rect 5416 -1298 5433 -1273
rect 5557 -1298 5574 -1266
rect 5756 -1298 5771 -1256
rect 5799 -1298 5814 -1256
rect 5996 -1273 6006 -1266
tri 6006 -1273 6013 -1266 sw
rect 5996 -1298 6013 -1273
rect 6137 -1298 6154 -1266
rect 6336 -1298 6351 -1256
rect 6379 -1298 6394 -1256
rect 6576 -1273 6586 -1266
tri 6586 -1273 6593 -1266 sw
rect 6576 -1298 6593 -1273
rect 6717 -1298 6734 -1266
rect 6916 -1298 6931 -1256
rect 259 -1336 291 -1322
rect 839 -1336 871 -1322
rect 1419 -1336 1451 -1322
rect 1999 -1336 2031 -1322
rect 2579 -1336 2611 -1322
rect 3159 -1336 3191 -1322
rect 3739 -1336 3771 -1322
rect 4319 -1336 4351 -1322
rect 4899 -1336 4931 -1322
rect 5479 -1336 5511 -1322
rect 6059 -1336 6091 -1322
rect 6639 -1336 6671 -1322
rect 73 -1422 88 -1394
rect 154 -1422 169 -1394
rect 381 -1422 396 -1394
rect 463 -1422 478 -1393
rect 653 -1422 668 -1394
rect 734 -1422 749 -1394
rect 961 -1422 976 -1394
rect 1043 -1422 1058 -1393
rect 1233 -1422 1248 -1394
rect 1314 -1422 1329 -1394
rect 1541 -1422 1556 -1394
rect 1623 -1422 1638 -1393
rect 1813 -1422 1828 -1394
rect 1894 -1422 1909 -1394
rect 2121 -1422 2136 -1394
rect 2203 -1422 2218 -1393
rect 2393 -1422 2408 -1394
rect 2474 -1422 2489 -1394
rect 2701 -1422 2716 -1394
rect 2783 -1422 2798 -1393
rect 2973 -1422 2988 -1394
rect 3054 -1422 3069 -1394
rect 3281 -1422 3296 -1394
rect 3363 -1422 3378 -1393
rect 3553 -1422 3568 -1394
rect 3634 -1422 3649 -1394
rect 3861 -1422 3876 -1394
rect 3943 -1422 3958 -1393
rect 4133 -1422 4148 -1394
rect 4214 -1422 4229 -1394
rect 4441 -1422 4456 -1394
rect 4523 -1422 4538 -1393
rect 4713 -1422 4728 -1394
rect 4794 -1422 4809 -1394
rect 5021 -1422 5036 -1394
rect 5103 -1422 5118 -1393
rect 5293 -1422 5308 -1394
rect 5374 -1422 5389 -1394
rect 5601 -1422 5616 -1394
rect 5683 -1422 5698 -1393
rect 5873 -1422 5888 -1394
rect 5954 -1422 5969 -1394
rect 6181 -1422 6196 -1394
rect 6263 -1422 6278 -1393
rect 6453 -1422 6468 -1394
rect 6534 -1422 6549 -1394
rect 6761 -1422 6776 -1394
rect 6843 -1422 6858 -1393
rect -1 -1568 14 -1526
rect 196 -1543 206 -1536
tri 206 -1543 213 -1536 sw
rect 196 -1568 213 -1543
rect 337 -1568 354 -1536
rect 536 -1568 551 -1526
rect 579 -1568 594 -1526
rect 776 -1543 786 -1536
tri 786 -1543 793 -1536 sw
rect 776 -1568 793 -1543
rect 917 -1568 934 -1536
rect 1116 -1568 1131 -1526
rect 1159 -1568 1174 -1526
rect 1356 -1543 1366 -1536
tri 1366 -1543 1373 -1536 sw
rect 1356 -1568 1373 -1543
rect 1497 -1568 1514 -1536
rect 1696 -1568 1711 -1526
rect 1739 -1568 1754 -1526
rect 1936 -1543 1946 -1536
tri 1946 -1543 1953 -1536 sw
rect 1936 -1568 1953 -1543
rect 2077 -1568 2094 -1536
rect 2276 -1568 2291 -1526
rect 2319 -1568 2334 -1526
rect 2516 -1543 2526 -1536
tri 2526 -1543 2533 -1536 sw
rect 2516 -1568 2533 -1543
rect 2657 -1568 2674 -1536
rect 2856 -1568 2871 -1526
rect 2899 -1568 2914 -1526
rect 3096 -1543 3106 -1536
tri 3106 -1543 3113 -1536 sw
rect 3096 -1568 3113 -1543
rect 3237 -1568 3254 -1536
rect 3436 -1568 3451 -1526
rect 3479 -1568 3494 -1526
rect 3676 -1543 3686 -1536
tri 3686 -1543 3693 -1536 sw
rect 3676 -1568 3693 -1543
rect 3817 -1568 3834 -1536
rect 4016 -1568 4031 -1526
rect 4059 -1568 4074 -1526
rect 4256 -1543 4266 -1536
tri 4266 -1543 4273 -1536 sw
rect 4256 -1568 4273 -1543
rect 4397 -1568 4414 -1536
rect 4596 -1568 4611 -1526
rect 4639 -1568 4654 -1526
rect 4836 -1543 4846 -1536
tri 4846 -1543 4853 -1536 sw
rect 4836 -1568 4853 -1543
rect 4977 -1568 4994 -1536
rect 5176 -1568 5191 -1526
rect 5219 -1568 5234 -1526
rect 5416 -1543 5426 -1536
tri 5426 -1543 5433 -1536 sw
rect 5416 -1568 5433 -1543
rect 5557 -1568 5574 -1536
rect 5756 -1568 5771 -1526
rect 5799 -1568 5814 -1526
rect 5996 -1543 6006 -1536
tri 6006 -1543 6013 -1536 sw
rect 5996 -1568 6013 -1543
rect 6137 -1568 6154 -1536
rect 6336 -1568 6351 -1526
rect 6379 -1568 6394 -1526
rect 6576 -1543 6586 -1536
tri 6586 -1543 6593 -1536 sw
rect 6576 -1568 6593 -1543
rect 6717 -1568 6734 -1536
rect 6916 -1568 6931 -1526
rect 259 -1606 291 -1592
rect 839 -1606 871 -1592
rect 1419 -1606 1451 -1592
rect 1999 -1606 2031 -1592
rect 2579 -1606 2611 -1592
rect 3159 -1606 3191 -1592
rect 3739 -1606 3771 -1592
rect 4319 -1606 4351 -1592
rect 4899 -1606 4931 -1592
rect 5479 -1606 5511 -1592
rect 6059 -1606 6091 -1592
rect 6639 -1606 6671 -1592
rect 73 -1692 88 -1664
rect 154 -1692 169 -1664
rect 381 -1692 396 -1664
rect 463 -1692 478 -1663
rect 653 -1692 668 -1664
rect 734 -1692 749 -1664
rect 961 -1692 976 -1664
rect 1043 -1692 1058 -1663
rect 1233 -1692 1248 -1664
rect 1314 -1692 1329 -1664
rect 1541 -1692 1556 -1664
rect 1623 -1692 1638 -1663
rect 1813 -1692 1828 -1664
rect 1894 -1692 1909 -1664
rect 2121 -1692 2136 -1664
rect 2203 -1692 2218 -1663
rect 2393 -1692 2408 -1664
rect 2474 -1692 2489 -1664
rect 2701 -1692 2716 -1664
rect 2783 -1692 2798 -1663
rect 2973 -1692 2988 -1664
rect 3054 -1692 3069 -1664
rect 3281 -1692 3296 -1664
rect 3363 -1692 3378 -1663
rect 3553 -1692 3568 -1664
rect 3634 -1692 3649 -1664
rect 3861 -1692 3876 -1664
rect 3943 -1692 3958 -1663
rect 4133 -1692 4148 -1664
rect 4214 -1692 4229 -1664
rect 4441 -1692 4456 -1664
rect 4523 -1692 4538 -1663
rect 4713 -1692 4728 -1664
rect 4794 -1692 4809 -1664
rect 5021 -1692 5036 -1664
rect 5103 -1692 5118 -1663
rect 5293 -1692 5308 -1664
rect 5374 -1692 5389 -1664
rect 5601 -1692 5616 -1664
rect 5683 -1692 5698 -1663
rect 5873 -1692 5888 -1664
rect 5954 -1692 5969 -1664
rect 6181 -1692 6196 -1664
rect 6263 -1692 6278 -1663
rect 6453 -1692 6468 -1664
rect 6534 -1692 6549 -1664
rect 6761 -1692 6776 -1664
rect 6843 -1692 6858 -1663
rect -1 -1838 14 -1796
rect 196 -1813 206 -1806
tri 206 -1813 213 -1806 sw
rect 196 -1838 213 -1813
rect 337 -1838 354 -1806
rect 536 -1838 551 -1796
rect 579 -1838 594 -1796
rect 776 -1813 786 -1806
tri 786 -1813 793 -1806 sw
rect 776 -1838 793 -1813
rect 917 -1838 934 -1806
rect 1116 -1838 1131 -1796
rect 1159 -1838 1174 -1796
rect 1356 -1813 1366 -1806
tri 1366 -1813 1373 -1806 sw
rect 1356 -1838 1373 -1813
rect 1497 -1838 1514 -1806
rect 1696 -1838 1711 -1796
rect 1739 -1838 1754 -1796
rect 1936 -1813 1946 -1806
tri 1946 -1813 1953 -1806 sw
rect 1936 -1838 1953 -1813
rect 2077 -1838 2094 -1806
rect 2276 -1838 2291 -1796
rect 2319 -1838 2334 -1796
rect 2516 -1813 2526 -1806
tri 2526 -1813 2533 -1806 sw
rect 2516 -1838 2533 -1813
rect 2657 -1838 2674 -1806
rect 2856 -1838 2871 -1796
rect 2899 -1838 2914 -1796
rect 3096 -1813 3106 -1806
tri 3106 -1813 3113 -1806 sw
rect 3096 -1838 3113 -1813
rect 3237 -1838 3254 -1806
rect 3436 -1838 3451 -1796
rect 3479 -1838 3494 -1796
rect 3676 -1813 3686 -1806
tri 3686 -1813 3693 -1806 sw
rect 3676 -1838 3693 -1813
rect 3817 -1838 3834 -1806
rect 4016 -1838 4031 -1796
rect 4059 -1838 4074 -1796
rect 4256 -1813 4266 -1806
tri 4266 -1813 4273 -1806 sw
rect 4256 -1838 4273 -1813
rect 4397 -1838 4414 -1806
rect 4596 -1838 4611 -1796
rect 4639 -1838 4654 -1796
rect 4836 -1813 4846 -1806
tri 4846 -1813 4853 -1806 sw
rect 4836 -1838 4853 -1813
rect 4977 -1838 4994 -1806
rect 5176 -1838 5191 -1796
rect 5219 -1838 5234 -1796
rect 5416 -1813 5426 -1806
tri 5426 -1813 5433 -1806 sw
rect 5416 -1838 5433 -1813
rect 5557 -1838 5574 -1806
rect 5756 -1838 5771 -1796
rect 5799 -1838 5814 -1796
rect 5996 -1813 6006 -1806
tri 6006 -1813 6013 -1806 sw
rect 5996 -1838 6013 -1813
rect 6137 -1838 6154 -1806
rect 6336 -1838 6351 -1796
rect 6379 -1838 6394 -1796
rect 6576 -1813 6586 -1806
tri 6586 -1813 6593 -1806 sw
rect 6576 -1838 6593 -1813
rect 6717 -1838 6734 -1806
rect 6916 -1838 6931 -1796
rect 259 -1876 291 -1862
rect 839 -1876 871 -1862
rect 1419 -1876 1451 -1862
rect 1999 -1876 2031 -1862
rect 2579 -1876 2611 -1862
rect 3159 -1876 3191 -1862
rect 3739 -1876 3771 -1862
rect 4319 -1876 4351 -1862
rect 4899 -1876 4931 -1862
rect 5479 -1876 5511 -1862
rect 6059 -1876 6091 -1862
rect 6639 -1876 6671 -1862
rect 73 -1962 88 -1934
rect 154 -1962 169 -1934
rect 381 -1962 396 -1934
rect 463 -1962 478 -1933
rect 653 -1962 668 -1934
rect 734 -1962 749 -1934
rect 961 -1962 976 -1934
rect 1043 -1962 1058 -1933
rect 1233 -1962 1248 -1934
rect 1314 -1962 1329 -1934
rect 1541 -1962 1556 -1934
rect 1623 -1962 1638 -1933
rect 1813 -1962 1828 -1934
rect 1894 -1962 1909 -1934
rect 2121 -1962 2136 -1934
rect 2203 -1962 2218 -1933
rect 2393 -1962 2408 -1934
rect 2474 -1962 2489 -1934
rect 2701 -1962 2716 -1934
rect 2783 -1962 2798 -1933
rect 2973 -1962 2988 -1934
rect 3054 -1962 3069 -1934
rect 3281 -1962 3296 -1934
rect 3363 -1962 3378 -1933
rect 3553 -1962 3568 -1934
rect 3634 -1962 3649 -1934
rect 3861 -1962 3876 -1934
rect 3943 -1962 3958 -1933
rect 4133 -1962 4148 -1934
rect 4214 -1962 4229 -1934
rect 4441 -1962 4456 -1934
rect 4523 -1962 4538 -1933
rect 4713 -1962 4728 -1934
rect 4794 -1962 4809 -1934
rect 5021 -1962 5036 -1934
rect 5103 -1962 5118 -1933
rect 5293 -1962 5308 -1934
rect 5374 -1962 5389 -1934
rect 5601 -1962 5616 -1934
rect 5683 -1962 5698 -1933
rect 5873 -1962 5888 -1934
rect 5954 -1962 5969 -1934
rect 6181 -1962 6196 -1934
rect 6263 -1962 6278 -1933
rect 6453 -1962 6468 -1934
rect 6534 -1962 6549 -1934
rect 6761 -1962 6776 -1934
rect 6843 -1962 6858 -1933
rect -1 -2108 14 -2066
rect 196 -2083 206 -2076
tri 206 -2083 213 -2076 sw
rect 196 -2108 213 -2083
rect 337 -2108 354 -2076
rect 536 -2108 551 -2066
rect 579 -2108 594 -2066
rect 776 -2083 786 -2076
tri 786 -2083 793 -2076 sw
rect 776 -2108 793 -2083
rect 917 -2108 934 -2076
rect 1116 -2108 1131 -2066
rect 1159 -2108 1174 -2066
rect 1356 -2083 1366 -2076
tri 1366 -2083 1373 -2076 sw
rect 1356 -2108 1373 -2083
rect 1497 -2108 1514 -2076
rect 1696 -2108 1711 -2066
rect 1739 -2108 1754 -2066
rect 1936 -2083 1946 -2076
tri 1946 -2083 1953 -2076 sw
rect 1936 -2108 1953 -2083
rect 2077 -2108 2094 -2076
rect 2276 -2108 2291 -2066
rect 2319 -2108 2334 -2066
rect 2516 -2083 2526 -2076
tri 2526 -2083 2533 -2076 sw
rect 2516 -2108 2533 -2083
rect 2657 -2108 2674 -2076
rect 2856 -2108 2871 -2066
rect 2899 -2108 2914 -2066
rect 3096 -2083 3106 -2076
tri 3106 -2083 3113 -2076 sw
rect 3096 -2108 3113 -2083
rect 3237 -2108 3254 -2076
rect 3436 -2108 3451 -2066
rect 3479 -2108 3494 -2066
rect 3676 -2083 3686 -2076
tri 3686 -2083 3693 -2076 sw
rect 3676 -2108 3693 -2083
rect 3817 -2108 3834 -2076
rect 4016 -2108 4031 -2066
rect 4059 -2108 4074 -2066
rect 4256 -2083 4266 -2076
tri 4266 -2083 4273 -2076 sw
rect 4256 -2108 4273 -2083
rect 4397 -2108 4414 -2076
rect 4596 -2108 4611 -2066
rect 4639 -2108 4654 -2066
rect 4836 -2083 4846 -2076
tri 4846 -2083 4853 -2076 sw
rect 4836 -2108 4853 -2083
rect 4977 -2108 4994 -2076
rect 5176 -2108 5191 -2066
rect 5219 -2108 5234 -2066
rect 5416 -2083 5426 -2076
tri 5426 -2083 5433 -2076 sw
rect 5416 -2108 5433 -2083
rect 5557 -2108 5574 -2076
rect 5756 -2108 5771 -2066
rect 5799 -2108 5814 -2066
rect 5996 -2083 6006 -2076
tri 6006 -2083 6013 -2076 sw
rect 5996 -2108 6013 -2083
rect 6137 -2108 6154 -2076
rect 6336 -2108 6351 -2066
rect 6379 -2108 6394 -2066
rect 6576 -2083 6586 -2076
tri 6586 -2083 6593 -2076 sw
rect 6576 -2108 6593 -2083
rect 6717 -2108 6734 -2076
rect 6916 -2108 6931 -2066
rect 259 -2146 291 -2132
rect 839 -2146 871 -2132
rect 1419 -2146 1451 -2132
rect 1999 -2146 2031 -2132
rect 2579 -2146 2611 -2132
rect 3159 -2146 3191 -2132
rect 3739 -2146 3771 -2132
rect 4319 -2146 4351 -2132
rect 4899 -2146 4931 -2132
rect 5479 -2146 5511 -2132
rect 6059 -2146 6091 -2132
rect 6639 -2146 6671 -2132
<< pdiffc >>
rect 259 2130 291 2144
rect 197 2078 212 2106
rect 338 2090 350 2106
tri 338 2078 350 2090 ne
rect 839 2130 871 2144
rect 777 2078 792 2106
rect 918 2090 930 2106
tri 918 2078 930 2090 ne
rect 1419 2130 1451 2144
rect 1357 2078 1372 2106
rect 1498 2090 1510 2106
tri 1498 2078 1510 2090 ne
rect 1999 2130 2031 2144
rect 1937 2078 1952 2106
rect 2078 2090 2090 2106
tri 2078 2078 2090 2090 ne
rect 2579 2130 2611 2144
rect 2517 2078 2532 2106
rect 2658 2090 2670 2106
tri 2658 2078 2670 2090 ne
rect 3159 2130 3191 2144
rect 3097 2078 3112 2106
rect 3238 2090 3250 2106
tri 3238 2078 3250 2090 ne
rect 3739 2130 3771 2144
rect 3677 2078 3692 2106
rect 3818 2090 3830 2106
tri 3818 2078 3830 2090 ne
rect 4319 2130 4351 2144
rect 4257 2078 4272 2106
rect 4398 2090 4410 2106
tri 4398 2078 4410 2090 ne
rect 4899 2130 4931 2144
rect 4837 2078 4852 2106
rect 4978 2090 4990 2106
tri 4978 2078 4990 2090 ne
rect 5479 2130 5511 2144
rect 5417 2078 5432 2106
rect 5558 2090 5570 2106
tri 5558 2078 5570 2090 ne
rect 6059 2130 6091 2144
rect 5997 2078 6012 2106
rect 6138 2090 6150 2106
tri 6138 2078 6150 2090 ne
rect 6639 2130 6671 2144
rect 6577 2078 6592 2106
rect 6718 2090 6730 2106
tri 6718 2078 6730 2090 ne
rect 259 1860 291 1874
rect 197 1808 212 1836
rect 338 1820 350 1836
tri 338 1808 350 1820 ne
rect 839 1860 871 1874
rect 777 1808 792 1836
rect 918 1820 930 1836
tri 918 1808 930 1820 ne
rect 1419 1860 1451 1874
rect 1357 1808 1372 1836
rect 1498 1820 1510 1836
tri 1498 1808 1510 1820 ne
rect 1999 1860 2031 1874
rect 1937 1808 1952 1836
rect 2078 1820 2090 1836
tri 2078 1808 2090 1820 ne
rect 2579 1860 2611 1874
rect 2517 1808 2532 1836
rect 2658 1820 2670 1836
tri 2658 1808 2670 1820 ne
rect 3159 1860 3191 1874
rect 3097 1808 3112 1836
rect 3238 1820 3250 1836
tri 3238 1808 3250 1820 ne
rect 3739 1860 3771 1874
rect 3677 1808 3692 1836
rect 3818 1820 3830 1836
tri 3818 1808 3830 1820 ne
rect 4319 1860 4351 1874
rect 4257 1808 4272 1836
rect 4398 1820 4410 1836
tri 4398 1808 4410 1820 ne
rect 4899 1860 4931 1874
rect 4837 1808 4852 1836
rect 4978 1820 4990 1836
tri 4978 1808 4990 1820 ne
rect 5479 1860 5511 1874
rect 5417 1808 5432 1836
rect 5558 1820 5570 1836
tri 5558 1808 5570 1820 ne
rect 6059 1860 6091 1874
rect 5997 1808 6012 1836
rect 6138 1820 6150 1836
tri 6138 1808 6150 1820 ne
rect 6639 1860 6671 1874
rect 6577 1808 6592 1836
rect 6718 1820 6730 1836
tri 6718 1808 6730 1820 ne
rect 259 1590 291 1604
rect 197 1538 212 1566
rect 338 1550 350 1566
tri 338 1538 350 1550 ne
rect 839 1590 871 1604
rect 777 1538 792 1566
rect 918 1550 930 1566
tri 918 1538 930 1550 ne
rect 1419 1590 1451 1604
rect 1357 1538 1372 1566
rect 1498 1550 1510 1566
tri 1498 1538 1510 1550 ne
rect 1999 1590 2031 1604
rect 1937 1538 1952 1566
rect 2078 1550 2090 1566
tri 2078 1538 2090 1550 ne
rect 2579 1590 2611 1604
rect 2517 1538 2532 1566
rect 2658 1550 2670 1566
tri 2658 1538 2670 1550 ne
rect 3159 1590 3191 1604
rect 3097 1538 3112 1566
rect 3238 1550 3250 1566
tri 3238 1538 3250 1550 ne
rect 3739 1590 3771 1604
rect 3677 1538 3692 1566
rect 3818 1550 3830 1566
tri 3818 1538 3830 1550 ne
rect 4319 1590 4351 1604
rect 4257 1538 4272 1566
rect 4398 1550 4410 1566
tri 4398 1538 4410 1550 ne
rect 4899 1590 4931 1604
rect 4837 1538 4852 1566
rect 4978 1550 4990 1566
tri 4978 1538 4990 1550 ne
rect 5479 1590 5511 1604
rect 5417 1538 5432 1566
rect 5558 1550 5570 1566
tri 5558 1538 5570 1550 ne
rect 6059 1590 6091 1604
rect 5997 1538 6012 1566
rect 6138 1550 6150 1566
tri 6138 1538 6150 1550 ne
rect 6639 1590 6671 1604
rect 6577 1538 6592 1566
rect 6718 1550 6730 1566
tri 6718 1538 6730 1550 ne
rect 259 1320 291 1334
rect 197 1268 212 1296
rect 338 1280 350 1296
tri 338 1268 350 1280 ne
rect 839 1320 871 1334
rect 777 1268 792 1296
rect 918 1280 930 1296
tri 918 1268 930 1280 ne
rect 1419 1320 1451 1334
rect 1357 1268 1372 1296
rect 1498 1280 1510 1296
tri 1498 1268 1510 1280 ne
rect 1999 1320 2031 1334
rect 1937 1268 1952 1296
rect 2078 1280 2090 1296
tri 2078 1268 2090 1280 ne
rect 2579 1320 2611 1334
rect 2517 1268 2532 1296
rect 2658 1280 2670 1296
tri 2658 1268 2670 1280 ne
rect 3159 1320 3191 1334
rect 3097 1268 3112 1296
rect 3238 1280 3250 1296
tri 3238 1268 3250 1280 ne
rect 3739 1320 3771 1334
rect 3677 1268 3692 1296
rect 3818 1280 3830 1296
tri 3818 1268 3830 1280 ne
rect 4319 1320 4351 1334
rect 4257 1268 4272 1296
rect 4398 1280 4410 1296
tri 4398 1268 4410 1280 ne
rect 4899 1320 4931 1334
rect 4837 1268 4852 1296
rect 4978 1280 4990 1296
tri 4978 1268 4990 1280 ne
rect 5479 1320 5511 1334
rect 5417 1268 5432 1296
rect 5558 1280 5570 1296
tri 5558 1268 5570 1280 ne
rect 6059 1320 6091 1334
rect 5997 1268 6012 1296
rect 6138 1280 6150 1296
tri 6138 1268 6150 1280 ne
rect 6639 1320 6671 1334
rect 6577 1268 6592 1296
rect 6718 1280 6730 1296
tri 6718 1268 6730 1280 ne
rect 259 1050 291 1064
rect 197 998 212 1026
rect 338 1010 350 1026
tri 338 998 350 1010 ne
rect 839 1050 871 1064
rect 777 998 792 1026
rect 918 1010 930 1026
tri 918 998 930 1010 ne
rect 1419 1050 1451 1064
rect 1357 998 1372 1026
rect 1498 1010 1510 1026
tri 1498 998 1510 1010 ne
rect 1999 1050 2031 1064
rect 1937 998 1952 1026
rect 2078 1010 2090 1026
tri 2078 998 2090 1010 ne
rect 2579 1050 2611 1064
rect 2517 998 2532 1026
rect 2658 1010 2670 1026
tri 2658 998 2670 1010 ne
rect 3159 1050 3191 1064
rect 3097 998 3112 1026
rect 3238 1010 3250 1026
tri 3238 998 3250 1010 ne
rect 3739 1050 3771 1064
rect 3677 998 3692 1026
rect 3818 1010 3830 1026
tri 3818 998 3830 1010 ne
rect 4319 1050 4351 1064
rect 4257 998 4272 1026
rect 4398 1010 4410 1026
tri 4398 998 4410 1010 ne
rect 4899 1050 4931 1064
rect 4837 998 4852 1026
rect 4978 1010 4990 1026
tri 4978 998 4990 1010 ne
rect 5479 1050 5511 1064
rect 5417 998 5432 1026
rect 5558 1010 5570 1026
tri 5558 998 5570 1010 ne
rect 6059 1050 6091 1064
rect 5997 998 6012 1026
rect 6138 1010 6150 1026
tri 6138 998 6150 1010 ne
rect 6639 1050 6671 1064
rect 6577 998 6592 1026
rect 6718 1010 6730 1026
tri 6718 998 6730 1010 ne
rect 259 780 291 794
rect 197 728 212 756
rect 338 740 350 756
tri 338 728 350 740 ne
rect 839 780 871 794
rect 777 728 792 756
rect 918 740 930 756
tri 918 728 930 740 ne
rect 1419 780 1451 794
rect 1357 728 1372 756
rect 1498 740 1510 756
tri 1498 728 1510 740 ne
rect 1999 780 2031 794
rect 1937 728 1952 756
rect 2078 740 2090 756
tri 2078 728 2090 740 ne
rect 2579 780 2611 794
rect 2517 728 2532 756
rect 2658 740 2670 756
tri 2658 728 2670 740 ne
rect 3159 780 3191 794
rect 3097 728 3112 756
rect 3238 740 3250 756
tri 3238 728 3250 740 ne
rect 3739 780 3771 794
rect 3677 728 3692 756
rect 3818 740 3830 756
tri 3818 728 3830 740 ne
rect 4319 780 4351 794
rect 4257 728 4272 756
rect 4398 740 4410 756
tri 4398 728 4410 740 ne
rect 4899 780 4931 794
rect 4837 728 4852 756
rect 4978 740 4990 756
tri 4978 728 4990 740 ne
rect 5479 780 5511 794
rect 5417 728 5432 756
rect 5558 740 5570 756
tri 5558 728 5570 740 ne
rect 6059 780 6091 794
rect 5997 728 6012 756
rect 6138 740 6150 756
tri 6138 728 6150 740 ne
rect 6639 780 6671 794
rect 6577 728 6592 756
rect 6718 740 6730 756
tri 6718 728 6730 740 ne
rect 259 510 291 524
rect 197 458 212 486
rect 338 470 350 486
tri 338 458 350 470 ne
rect 839 510 871 524
rect 777 458 792 486
rect 918 470 930 486
tri 918 458 930 470 ne
rect 1419 510 1451 524
rect 1357 458 1372 486
rect 1498 470 1510 486
tri 1498 458 1510 470 ne
rect 1999 510 2031 524
rect 1937 458 1952 486
rect 2078 470 2090 486
tri 2078 458 2090 470 ne
rect 2579 510 2611 524
rect 2517 458 2532 486
rect 2658 470 2670 486
tri 2658 458 2670 470 ne
rect 3159 510 3191 524
rect 3097 458 3112 486
rect 3238 470 3250 486
tri 3238 458 3250 470 ne
rect 3739 510 3771 524
rect 3677 458 3692 486
rect 3818 470 3830 486
tri 3818 458 3830 470 ne
rect 4319 510 4351 524
rect 4257 458 4272 486
rect 4398 470 4410 486
tri 4398 458 4410 470 ne
rect 4899 510 4931 524
rect 4837 458 4852 486
rect 4978 470 4990 486
tri 4978 458 4990 470 ne
rect 5479 510 5511 524
rect 5417 458 5432 486
rect 5558 470 5570 486
tri 5558 458 5570 470 ne
rect 6059 510 6091 524
rect 5997 458 6012 486
rect 6138 470 6150 486
tri 6138 458 6150 470 ne
rect 6639 510 6671 524
rect 6577 458 6592 486
rect 6718 470 6730 486
tri 6718 458 6730 470 ne
rect 259 240 291 254
rect 197 188 212 216
rect 338 200 350 216
tri 338 188 350 200 ne
rect 839 240 871 254
rect 777 188 792 216
rect 918 200 930 216
tri 918 188 930 200 ne
rect 1419 240 1451 254
rect 1357 188 1372 216
rect 1498 200 1510 216
tri 1498 188 1510 200 ne
rect 1999 240 2031 254
rect 1937 188 1952 216
rect 2078 200 2090 216
tri 2078 188 2090 200 ne
rect 2579 240 2611 254
rect 2517 188 2532 216
rect 2658 200 2670 216
tri 2658 188 2670 200 ne
rect 3159 240 3191 254
rect 3097 188 3112 216
rect 3238 200 3250 216
tri 3238 188 3250 200 ne
rect 3739 240 3771 254
rect 3677 188 3692 216
rect 3818 200 3830 216
tri 3818 188 3830 200 ne
rect 4319 240 4351 254
rect 4257 188 4272 216
rect 4398 200 4410 216
tri 4398 188 4410 200 ne
rect 4899 240 4931 254
rect 4837 188 4852 216
rect 4978 200 4990 216
tri 4978 188 4990 200 ne
rect 5479 240 5511 254
rect 5417 188 5432 216
rect 5558 200 5570 216
tri 5558 188 5570 200 ne
rect 6059 240 6091 254
rect 5997 188 6012 216
rect 6138 200 6150 216
tri 6138 188 6150 200 ne
rect 6639 240 6671 254
rect 6577 188 6592 216
rect 6718 200 6730 216
tri 6718 188 6730 200 ne
rect 259 -30 291 -16
rect 197 -82 212 -54
rect 338 -70 350 -54
tri 338 -82 350 -70 ne
rect 839 -30 871 -16
rect 777 -82 792 -54
rect 918 -70 930 -54
tri 918 -82 930 -70 ne
rect 1419 -30 1451 -16
rect 1357 -82 1372 -54
rect 1498 -70 1510 -54
tri 1498 -82 1510 -70 ne
rect 1999 -30 2031 -16
rect 1937 -82 1952 -54
rect 2078 -70 2090 -54
tri 2078 -82 2090 -70 ne
rect 2579 -30 2611 -16
rect 2517 -82 2532 -54
rect 2658 -70 2670 -54
tri 2658 -82 2670 -70 ne
rect 3159 -30 3191 -16
rect 3097 -82 3112 -54
rect 3238 -70 3250 -54
tri 3238 -82 3250 -70 ne
rect 3739 -30 3771 -16
rect 3677 -82 3692 -54
rect 3818 -70 3830 -54
tri 3818 -82 3830 -70 ne
rect 4319 -30 4351 -16
rect 4257 -82 4272 -54
rect 4398 -70 4410 -54
tri 4398 -82 4410 -70 ne
rect 4899 -30 4931 -16
rect 4837 -82 4852 -54
rect 4978 -70 4990 -54
tri 4978 -82 4990 -70 ne
rect 5479 -30 5511 -16
rect 5417 -82 5432 -54
rect 5558 -70 5570 -54
tri 5558 -82 5570 -70 ne
rect 6059 -30 6091 -16
rect 5997 -82 6012 -54
rect 6138 -70 6150 -54
tri 6138 -82 6150 -70 ne
rect 6639 -30 6671 -16
rect 6577 -82 6592 -54
rect 6718 -70 6730 -54
tri 6718 -82 6730 -70 ne
rect 259 -300 291 -286
rect 197 -352 212 -324
rect 338 -340 350 -324
tri 338 -352 350 -340 ne
rect 839 -300 871 -286
rect 777 -352 792 -324
rect 918 -340 930 -324
tri 918 -352 930 -340 ne
rect 1419 -300 1451 -286
rect 1357 -352 1372 -324
rect 1498 -340 1510 -324
tri 1498 -352 1510 -340 ne
rect 1999 -300 2031 -286
rect 1937 -352 1952 -324
rect 2078 -340 2090 -324
tri 2078 -352 2090 -340 ne
rect 2579 -300 2611 -286
rect 2517 -352 2532 -324
rect 2658 -340 2670 -324
tri 2658 -352 2670 -340 ne
rect 3159 -300 3191 -286
rect 3097 -352 3112 -324
rect 3238 -340 3250 -324
tri 3238 -352 3250 -340 ne
rect 3739 -300 3771 -286
rect 3677 -352 3692 -324
rect 3818 -340 3830 -324
tri 3818 -352 3830 -340 ne
rect 4319 -300 4351 -286
rect 4257 -352 4272 -324
rect 4398 -340 4410 -324
tri 4398 -352 4410 -340 ne
rect 4899 -300 4931 -286
rect 4837 -352 4852 -324
rect 4978 -340 4990 -324
tri 4978 -352 4990 -340 ne
rect 5479 -300 5511 -286
rect 5417 -352 5432 -324
rect 5558 -340 5570 -324
tri 5558 -352 5570 -340 ne
rect 6059 -300 6091 -286
rect 5997 -352 6012 -324
rect 6138 -340 6150 -324
tri 6138 -352 6150 -340 ne
rect 6639 -300 6671 -286
rect 6577 -352 6592 -324
rect 6718 -340 6730 -324
tri 6718 -352 6730 -340 ne
rect 259 -570 291 -556
rect 197 -622 212 -594
rect 338 -610 350 -594
tri 338 -622 350 -610 ne
rect 839 -570 871 -556
rect 777 -622 792 -594
rect 918 -610 930 -594
tri 918 -622 930 -610 ne
rect 1419 -570 1451 -556
rect 1357 -622 1372 -594
rect 1498 -610 1510 -594
tri 1498 -622 1510 -610 ne
rect 1999 -570 2031 -556
rect 1937 -622 1952 -594
rect 2078 -610 2090 -594
tri 2078 -622 2090 -610 ne
rect 2579 -570 2611 -556
rect 2517 -622 2532 -594
rect 2658 -610 2670 -594
tri 2658 -622 2670 -610 ne
rect 3159 -570 3191 -556
rect 3097 -622 3112 -594
rect 3238 -610 3250 -594
tri 3238 -622 3250 -610 ne
rect 3739 -570 3771 -556
rect 3677 -622 3692 -594
rect 3818 -610 3830 -594
tri 3818 -622 3830 -610 ne
rect 4319 -570 4351 -556
rect 4257 -622 4272 -594
rect 4398 -610 4410 -594
tri 4398 -622 4410 -610 ne
rect 4899 -570 4931 -556
rect 4837 -622 4852 -594
rect 4978 -610 4990 -594
tri 4978 -622 4990 -610 ne
rect 5479 -570 5511 -556
rect 5417 -622 5432 -594
rect 5558 -610 5570 -594
tri 5558 -622 5570 -610 ne
rect 6059 -570 6091 -556
rect 5997 -622 6012 -594
rect 6138 -610 6150 -594
tri 6138 -622 6150 -610 ne
rect 6639 -570 6671 -556
rect 6577 -622 6592 -594
rect 6718 -610 6730 -594
tri 6718 -622 6730 -610 ne
rect 259 -840 291 -826
rect 197 -892 212 -864
rect 338 -880 350 -864
tri 338 -892 350 -880 ne
rect 839 -840 871 -826
rect 777 -892 792 -864
rect 918 -880 930 -864
tri 918 -892 930 -880 ne
rect 1419 -840 1451 -826
rect 1357 -892 1372 -864
rect 1498 -880 1510 -864
tri 1498 -892 1510 -880 ne
rect 1999 -840 2031 -826
rect 1937 -892 1952 -864
rect 2078 -880 2090 -864
tri 2078 -892 2090 -880 ne
rect 2579 -840 2611 -826
rect 2517 -892 2532 -864
rect 2658 -880 2670 -864
tri 2658 -892 2670 -880 ne
rect 3159 -840 3191 -826
rect 3097 -892 3112 -864
rect 3238 -880 3250 -864
tri 3238 -892 3250 -880 ne
rect 3739 -840 3771 -826
rect 3677 -892 3692 -864
rect 3818 -880 3830 -864
tri 3818 -892 3830 -880 ne
rect 4319 -840 4351 -826
rect 4257 -892 4272 -864
rect 4398 -880 4410 -864
tri 4398 -892 4410 -880 ne
rect 4899 -840 4931 -826
rect 4837 -892 4852 -864
rect 4978 -880 4990 -864
tri 4978 -892 4990 -880 ne
rect 5479 -840 5511 -826
rect 5417 -892 5432 -864
rect 5558 -880 5570 -864
tri 5558 -892 5570 -880 ne
rect 6059 -840 6091 -826
rect 5997 -892 6012 -864
rect 6138 -880 6150 -864
tri 6138 -892 6150 -880 ne
rect 6639 -840 6671 -826
rect 6577 -892 6592 -864
rect 6718 -880 6730 -864
tri 6718 -892 6730 -880 ne
rect 259 -1110 291 -1096
rect 197 -1162 212 -1134
rect 338 -1150 350 -1134
tri 338 -1162 350 -1150 ne
rect 839 -1110 871 -1096
rect 777 -1162 792 -1134
rect 918 -1150 930 -1134
tri 918 -1162 930 -1150 ne
rect 1419 -1110 1451 -1096
rect 1357 -1162 1372 -1134
rect 1498 -1150 1510 -1134
tri 1498 -1162 1510 -1150 ne
rect 1999 -1110 2031 -1096
rect 1937 -1162 1952 -1134
rect 2078 -1150 2090 -1134
tri 2078 -1162 2090 -1150 ne
rect 2579 -1110 2611 -1096
rect 2517 -1162 2532 -1134
rect 2658 -1150 2670 -1134
tri 2658 -1162 2670 -1150 ne
rect 3159 -1110 3191 -1096
rect 3097 -1162 3112 -1134
rect 3238 -1150 3250 -1134
tri 3238 -1162 3250 -1150 ne
rect 3739 -1110 3771 -1096
rect 3677 -1162 3692 -1134
rect 3818 -1150 3830 -1134
tri 3818 -1162 3830 -1150 ne
rect 4319 -1110 4351 -1096
rect 4257 -1162 4272 -1134
rect 4398 -1150 4410 -1134
tri 4398 -1162 4410 -1150 ne
rect 4899 -1110 4931 -1096
rect 4837 -1162 4852 -1134
rect 4978 -1150 4990 -1134
tri 4978 -1162 4990 -1150 ne
rect 5479 -1110 5511 -1096
rect 5417 -1162 5432 -1134
rect 5558 -1150 5570 -1134
tri 5558 -1162 5570 -1150 ne
rect 6059 -1110 6091 -1096
rect 5997 -1162 6012 -1134
rect 6138 -1150 6150 -1134
tri 6138 -1162 6150 -1150 ne
rect 6639 -1110 6671 -1096
rect 6577 -1162 6592 -1134
rect 6718 -1150 6730 -1134
tri 6718 -1162 6730 -1150 ne
rect 259 -1380 291 -1366
rect 197 -1432 212 -1404
rect 338 -1420 350 -1404
tri 338 -1432 350 -1420 ne
rect 839 -1380 871 -1366
rect 777 -1432 792 -1404
rect 918 -1420 930 -1404
tri 918 -1432 930 -1420 ne
rect 1419 -1380 1451 -1366
rect 1357 -1432 1372 -1404
rect 1498 -1420 1510 -1404
tri 1498 -1432 1510 -1420 ne
rect 1999 -1380 2031 -1366
rect 1937 -1432 1952 -1404
rect 2078 -1420 2090 -1404
tri 2078 -1432 2090 -1420 ne
rect 2579 -1380 2611 -1366
rect 2517 -1432 2532 -1404
rect 2658 -1420 2670 -1404
tri 2658 -1432 2670 -1420 ne
rect 3159 -1380 3191 -1366
rect 3097 -1432 3112 -1404
rect 3238 -1420 3250 -1404
tri 3238 -1432 3250 -1420 ne
rect 3739 -1380 3771 -1366
rect 3677 -1432 3692 -1404
rect 3818 -1420 3830 -1404
tri 3818 -1432 3830 -1420 ne
rect 4319 -1380 4351 -1366
rect 4257 -1432 4272 -1404
rect 4398 -1420 4410 -1404
tri 4398 -1432 4410 -1420 ne
rect 4899 -1380 4931 -1366
rect 4837 -1432 4852 -1404
rect 4978 -1420 4990 -1404
tri 4978 -1432 4990 -1420 ne
rect 5479 -1380 5511 -1366
rect 5417 -1432 5432 -1404
rect 5558 -1420 5570 -1404
tri 5558 -1432 5570 -1420 ne
rect 6059 -1380 6091 -1366
rect 5997 -1432 6012 -1404
rect 6138 -1420 6150 -1404
tri 6138 -1432 6150 -1420 ne
rect 6639 -1380 6671 -1366
rect 6577 -1432 6592 -1404
rect 6718 -1420 6730 -1404
tri 6718 -1432 6730 -1420 ne
rect 259 -1650 291 -1636
rect 197 -1702 212 -1674
rect 338 -1690 350 -1674
tri 338 -1702 350 -1690 ne
rect 839 -1650 871 -1636
rect 777 -1702 792 -1674
rect 918 -1690 930 -1674
tri 918 -1702 930 -1690 ne
rect 1419 -1650 1451 -1636
rect 1357 -1702 1372 -1674
rect 1498 -1690 1510 -1674
tri 1498 -1702 1510 -1690 ne
rect 1999 -1650 2031 -1636
rect 1937 -1702 1952 -1674
rect 2078 -1690 2090 -1674
tri 2078 -1702 2090 -1690 ne
rect 2579 -1650 2611 -1636
rect 2517 -1702 2532 -1674
rect 2658 -1690 2670 -1674
tri 2658 -1702 2670 -1690 ne
rect 3159 -1650 3191 -1636
rect 3097 -1702 3112 -1674
rect 3238 -1690 3250 -1674
tri 3238 -1702 3250 -1690 ne
rect 3739 -1650 3771 -1636
rect 3677 -1702 3692 -1674
rect 3818 -1690 3830 -1674
tri 3818 -1702 3830 -1690 ne
rect 4319 -1650 4351 -1636
rect 4257 -1702 4272 -1674
rect 4398 -1690 4410 -1674
tri 4398 -1702 4410 -1690 ne
rect 4899 -1650 4931 -1636
rect 4837 -1702 4852 -1674
rect 4978 -1690 4990 -1674
tri 4978 -1702 4990 -1690 ne
rect 5479 -1650 5511 -1636
rect 5417 -1702 5432 -1674
rect 5558 -1690 5570 -1674
tri 5558 -1702 5570 -1690 ne
rect 6059 -1650 6091 -1636
rect 5997 -1702 6012 -1674
rect 6138 -1690 6150 -1674
tri 6138 -1702 6150 -1690 ne
rect 6639 -1650 6671 -1636
rect 6577 -1702 6592 -1674
rect 6718 -1690 6730 -1674
tri 6718 -1702 6730 -1690 ne
rect 259 -1920 291 -1906
rect 197 -1972 212 -1944
rect 338 -1960 350 -1944
tri 338 -1972 350 -1960 ne
rect 839 -1920 871 -1906
rect 777 -1972 792 -1944
rect 918 -1960 930 -1944
tri 918 -1972 930 -1960 ne
rect 1419 -1920 1451 -1906
rect 1357 -1972 1372 -1944
rect 1498 -1960 1510 -1944
tri 1498 -1972 1510 -1960 ne
rect 1999 -1920 2031 -1906
rect 1937 -1972 1952 -1944
rect 2078 -1960 2090 -1944
tri 2078 -1972 2090 -1960 ne
rect 2579 -1920 2611 -1906
rect 2517 -1972 2532 -1944
rect 2658 -1960 2670 -1944
tri 2658 -1972 2670 -1960 ne
rect 3159 -1920 3191 -1906
rect 3097 -1972 3112 -1944
rect 3238 -1960 3250 -1944
tri 3238 -1972 3250 -1960 ne
rect 3739 -1920 3771 -1906
rect 3677 -1972 3692 -1944
rect 3818 -1960 3830 -1944
tri 3818 -1972 3830 -1960 ne
rect 4319 -1920 4351 -1906
rect 4257 -1972 4272 -1944
rect 4398 -1960 4410 -1944
tri 4398 -1972 4410 -1960 ne
rect 4899 -1920 4931 -1906
rect 4837 -1972 4852 -1944
rect 4978 -1960 4990 -1944
tri 4978 -1972 4990 -1960 ne
rect 5479 -1920 5511 -1906
rect 5417 -1972 5432 -1944
rect 5558 -1960 5570 -1944
tri 5558 -1972 5570 -1960 ne
rect 6059 -1920 6091 -1906
rect 5997 -1972 6012 -1944
rect 6138 -1960 6150 -1944
tri 6138 -1972 6150 -1960 ne
rect 6639 -1920 6671 -1906
rect 6577 -1972 6592 -1944
rect 6718 -1960 6730 -1944
tri 6718 -1972 6730 -1960 ne
<< psubdiffcont >>
rect 261 1918 289 1920
rect 841 1918 869 1920
rect 1421 1918 1449 1920
rect 2001 1918 2029 1920
rect 2581 1918 2609 1920
rect 3161 1918 3189 1920
rect 3741 1918 3769 1920
rect 4321 1918 4349 1920
rect 4901 1918 4929 1920
rect 5481 1918 5509 1920
rect 6061 1918 6089 1920
rect 6641 1918 6669 1920
rect 261 1648 289 1650
rect 841 1648 869 1650
rect 1421 1648 1449 1650
rect 2001 1648 2029 1650
rect 2581 1648 2609 1650
rect 3161 1648 3189 1650
rect 3741 1648 3769 1650
rect 4321 1648 4349 1650
rect 4901 1648 4929 1650
rect 5481 1648 5509 1650
rect 6061 1648 6089 1650
rect 6641 1648 6669 1650
rect 261 1378 289 1380
rect 841 1378 869 1380
rect 1421 1378 1449 1380
rect 2001 1378 2029 1380
rect 2581 1378 2609 1380
rect 3161 1378 3189 1380
rect 3741 1378 3769 1380
rect 4321 1378 4349 1380
rect 4901 1378 4929 1380
rect 5481 1378 5509 1380
rect 6061 1378 6089 1380
rect 6641 1378 6669 1380
rect 261 1108 289 1110
rect 841 1108 869 1110
rect 1421 1108 1449 1110
rect 2001 1108 2029 1110
rect 2581 1108 2609 1110
rect 3161 1108 3189 1110
rect 3741 1108 3769 1110
rect 4321 1108 4349 1110
rect 4901 1108 4929 1110
rect 5481 1108 5509 1110
rect 6061 1108 6089 1110
rect 6641 1108 6669 1110
rect 261 838 289 840
rect 841 838 869 840
rect 1421 838 1449 840
rect 2001 838 2029 840
rect 2581 838 2609 840
rect 3161 838 3189 840
rect 3741 838 3769 840
rect 4321 838 4349 840
rect 4901 838 4929 840
rect 5481 838 5509 840
rect 6061 838 6089 840
rect 6641 838 6669 840
rect 261 568 289 570
rect 841 568 869 570
rect 1421 568 1449 570
rect 2001 568 2029 570
rect 2581 568 2609 570
rect 3161 568 3189 570
rect 3741 568 3769 570
rect 4321 568 4349 570
rect 4901 568 4929 570
rect 5481 568 5509 570
rect 6061 568 6089 570
rect 6641 568 6669 570
rect 261 298 289 300
rect 841 298 869 300
rect 1421 298 1449 300
rect 2001 298 2029 300
rect 2581 298 2609 300
rect 3161 298 3189 300
rect 3741 298 3769 300
rect 4321 298 4349 300
rect 4901 298 4929 300
rect 5481 298 5509 300
rect 6061 298 6089 300
rect 6641 298 6669 300
rect 261 28 289 30
rect 841 28 869 30
rect 1421 28 1449 30
rect 2001 28 2029 30
rect 2581 28 2609 30
rect 3161 28 3189 30
rect 3741 28 3769 30
rect 4321 28 4349 30
rect 4901 28 4929 30
rect 5481 28 5509 30
rect 6061 28 6089 30
rect 6641 28 6669 30
rect 261 -242 289 -240
rect 841 -242 869 -240
rect 1421 -242 1449 -240
rect 2001 -242 2029 -240
rect 2581 -242 2609 -240
rect 3161 -242 3189 -240
rect 3741 -242 3769 -240
rect 4321 -242 4349 -240
rect 4901 -242 4929 -240
rect 5481 -242 5509 -240
rect 6061 -242 6089 -240
rect 6641 -242 6669 -240
rect 261 -512 289 -510
rect 841 -512 869 -510
rect 1421 -512 1449 -510
rect 2001 -512 2029 -510
rect 2581 -512 2609 -510
rect 3161 -512 3189 -510
rect 3741 -512 3769 -510
rect 4321 -512 4349 -510
rect 4901 -512 4929 -510
rect 5481 -512 5509 -510
rect 6061 -512 6089 -510
rect 6641 -512 6669 -510
rect 261 -782 289 -780
rect 841 -782 869 -780
rect 1421 -782 1449 -780
rect 2001 -782 2029 -780
rect 2581 -782 2609 -780
rect 3161 -782 3189 -780
rect 3741 -782 3769 -780
rect 4321 -782 4349 -780
rect 4901 -782 4929 -780
rect 5481 -782 5509 -780
rect 6061 -782 6089 -780
rect 6641 -782 6669 -780
rect 261 -1052 289 -1050
rect 841 -1052 869 -1050
rect 1421 -1052 1449 -1050
rect 2001 -1052 2029 -1050
rect 2581 -1052 2609 -1050
rect 3161 -1052 3189 -1050
rect 3741 -1052 3769 -1050
rect 4321 -1052 4349 -1050
rect 4901 -1052 4929 -1050
rect 5481 -1052 5509 -1050
rect 6061 -1052 6089 -1050
rect 6641 -1052 6669 -1050
rect 261 -1322 289 -1320
rect 841 -1322 869 -1320
rect 1421 -1322 1449 -1320
rect 2001 -1322 2029 -1320
rect 2581 -1322 2609 -1320
rect 3161 -1322 3189 -1320
rect 3741 -1322 3769 -1320
rect 4321 -1322 4349 -1320
rect 4901 -1322 4929 -1320
rect 5481 -1322 5509 -1320
rect 6061 -1322 6089 -1320
rect 6641 -1322 6669 -1320
rect 261 -1592 289 -1590
rect 841 -1592 869 -1590
rect 1421 -1592 1449 -1590
rect 2001 -1592 2029 -1590
rect 2581 -1592 2609 -1590
rect 3161 -1592 3189 -1590
rect 3741 -1592 3769 -1590
rect 4321 -1592 4349 -1590
rect 4901 -1592 4929 -1590
rect 5481 -1592 5509 -1590
rect 6061 -1592 6089 -1590
rect 6641 -1592 6669 -1590
rect 261 -1862 289 -1860
rect 841 -1862 869 -1860
rect 1421 -1862 1449 -1860
rect 2001 -1862 2029 -1860
rect 2581 -1862 2609 -1860
rect 3161 -1862 3189 -1860
rect 3741 -1862 3769 -1860
rect 4321 -1862 4349 -1860
rect 4901 -1862 4929 -1860
rect 5481 -1862 5509 -1860
rect 6061 -1862 6089 -1860
rect 6641 -1862 6669 -1860
rect 261 -2132 289 -2130
rect 841 -2132 869 -2130
rect 1421 -2132 1449 -2130
rect 2001 -2132 2029 -2130
rect 2581 -2132 2609 -2130
rect 3161 -2132 3189 -2130
rect 3741 -2132 3769 -2130
rect 4321 -2132 4349 -2130
rect 4901 -2132 4929 -2130
rect 5481 -2132 5509 -2130
rect 6061 -2132 6089 -2130
rect 6641 -2132 6669 -2130
<< nsubdiffcont >>
rect 261 2128 289 2130
rect 841 2128 869 2130
rect 1421 2128 1449 2130
rect 2001 2128 2029 2130
rect 2581 2128 2609 2130
rect 3161 2128 3189 2130
rect 3741 2128 3769 2130
rect 4321 2128 4349 2130
rect 4901 2128 4929 2130
rect 5481 2128 5509 2130
rect 6061 2128 6089 2130
rect 6641 2128 6669 2130
rect 261 1858 289 1860
rect 841 1858 869 1860
rect 1421 1858 1449 1860
rect 2001 1858 2029 1860
rect 2581 1858 2609 1860
rect 3161 1858 3189 1860
rect 3741 1858 3769 1860
rect 4321 1858 4349 1860
rect 4901 1858 4929 1860
rect 5481 1858 5509 1860
rect 6061 1858 6089 1860
rect 6641 1858 6669 1860
rect 261 1588 289 1590
rect 841 1588 869 1590
rect 1421 1588 1449 1590
rect 2001 1588 2029 1590
rect 2581 1588 2609 1590
rect 3161 1588 3189 1590
rect 3741 1588 3769 1590
rect 4321 1588 4349 1590
rect 4901 1588 4929 1590
rect 5481 1588 5509 1590
rect 6061 1588 6089 1590
rect 6641 1588 6669 1590
rect 261 1318 289 1320
rect 841 1318 869 1320
rect 1421 1318 1449 1320
rect 2001 1318 2029 1320
rect 2581 1318 2609 1320
rect 3161 1318 3189 1320
rect 3741 1318 3769 1320
rect 4321 1318 4349 1320
rect 4901 1318 4929 1320
rect 5481 1318 5509 1320
rect 6061 1318 6089 1320
rect 6641 1318 6669 1320
rect 261 1048 289 1050
rect 841 1048 869 1050
rect 1421 1048 1449 1050
rect 2001 1048 2029 1050
rect 2581 1048 2609 1050
rect 3161 1048 3189 1050
rect 3741 1048 3769 1050
rect 4321 1048 4349 1050
rect 4901 1048 4929 1050
rect 5481 1048 5509 1050
rect 6061 1048 6089 1050
rect 6641 1048 6669 1050
rect 261 778 289 780
rect 841 778 869 780
rect 1421 778 1449 780
rect 2001 778 2029 780
rect 2581 778 2609 780
rect 3161 778 3189 780
rect 3741 778 3769 780
rect 4321 778 4349 780
rect 4901 778 4929 780
rect 5481 778 5509 780
rect 6061 778 6089 780
rect 6641 778 6669 780
rect 261 508 289 510
rect 841 508 869 510
rect 1421 508 1449 510
rect 2001 508 2029 510
rect 2581 508 2609 510
rect 3161 508 3189 510
rect 3741 508 3769 510
rect 4321 508 4349 510
rect 4901 508 4929 510
rect 5481 508 5509 510
rect 6061 508 6089 510
rect 6641 508 6669 510
rect 261 238 289 240
rect 841 238 869 240
rect 1421 238 1449 240
rect 2001 238 2029 240
rect 2581 238 2609 240
rect 3161 238 3189 240
rect 3741 238 3769 240
rect 4321 238 4349 240
rect 4901 238 4929 240
rect 5481 238 5509 240
rect 6061 238 6089 240
rect 6641 238 6669 240
rect 261 -32 289 -30
rect 841 -32 869 -30
rect 1421 -32 1449 -30
rect 2001 -32 2029 -30
rect 2581 -32 2609 -30
rect 3161 -32 3189 -30
rect 3741 -32 3769 -30
rect 4321 -32 4349 -30
rect 4901 -32 4929 -30
rect 5481 -32 5509 -30
rect 6061 -32 6089 -30
rect 6641 -32 6669 -30
rect 261 -302 289 -300
rect 841 -302 869 -300
rect 1421 -302 1449 -300
rect 2001 -302 2029 -300
rect 2581 -302 2609 -300
rect 3161 -302 3189 -300
rect 3741 -302 3769 -300
rect 4321 -302 4349 -300
rect 4901 -302 4929 -300
rect 5481 -302 5509 -300
rect 6061 -302 6089 -300
rect 6641 -302 6669 -300
rect 261 -572 289 -570
rect 841 -572 869 -570
rect 1421 -572 1449 -570
rect 2001 -572 2029 -570
rect 2581 -572 2609 -570
rect 3161 -572 3189 -570
rect 3741 -572 3769 -570
rect 4321 -572 4349 -570
rect 4901 -572 4929 -570
rect 5481 -572 5509 -570
rect 6061 -572 6089 -570
rect 6641 -572 6669 -570
rect 261 -842 289 -840
rect 841 -842 869 -840
rect 1421 -842 1449 -840
rect 2001 -842 2029 -840
rect 2581 -842 2609 -840
rect 3161 -842 3189 -840
rect 3741 -842 3769 -840
rect 4321 -842 4349 -840
rect 4901 -842 4929 -840
rect 5481 -842 5509 -840
rect 6061 -842 6089 -840
rect 6641 -842 6669 -840
rect 261 -1112 289 -1110
rect 841 -1112 869 -1110
rect 1421 -1112 1449 -1110
rect 2001 -1112 2029 -1110
rect 2581 -1112 2609 -1110
rect 3161 -1112 3189 -1110
rect 3741 -1112 3769 -1110
rect 4321 -1112 4349 -1110
rect 4901 -1112 4929 -1110
rect 5481 -1112 5509 -1110
rect 6061 -1112 6089 -1110
rect 6641 -1112 6669 -1110
rect 261 -1382 289 -1380
rect 841 -1382 869 -1380
rect 1421 -1382 1449 -1380
rect 2001 -1382 2029 -1380
rect 2581 -1382 2609 -1380
rect 3161 -1382 3189 -1380
rect 3741 -1382 3769 -1380
rect 4321 -1382 4349 -1380
rect 4901 -1382 4929 -1380
rect 5481 -1382 5509 -1380
rect 6061 -1382 6089 -1380
rect 6641 -1382 6669 -1380
rect 261 -1652 289 -1650
rect 841 -1652 869 -1650
rect 1421 -1652 1449 -1650
rect 2001 -1652 2029 -1650
rect 2581 -1652 2609 -1650
rect 3161 -1652 3189 -1650
rect 3741 -1652 3769 -1650
rect 4321 -1652 4349 -1650
rect 4901 -1652 4929 -1650
rect 5481 -1652 5509 -1650
rect 6061 -1652 6089 -1650
rect 6641 -1652 6669 -1650
rect 261 -1922 289 -1920
rect 841 -1922 869 -1920
rect 1421 -1922 1449 -1920
rect 2001 -1922 2029 -1920
rect 2581 -1922 2609 -1920
rect 3161 -1922 3189 -1920
rect 3741 -1922 3769 -1920
rect 4321 -1922 4349 -1920
rect 4901 -1922 4929 -1920
rect 5481 -1922 5509 -1920
rect 6061 -1922 6089 -1920
rect 6641 -1922 6669 -1920
<< poly >>
rect -1 2144 6931 2174
rect 106 2116 136 2144
rect 221 2106 251 2128
rect 299 2106 329 2128
rect 414 2116 444 2144
rect 106 2066 136 2088
rect 686 2116 716 2144
rect 801 2106 831 2128
rect 879 2106 909 2128
rect 994 2116 1024 2144
rect 221 2045 251 2078
rect 42 1984 72 2006
rect 128 1984 143 2018
rect 221 1984 251 2011
rect 299 2045 329 2078
rect 414 2066 444 2088
rect 686 2066 716 2088
rect 1266 2116 1296 2144
rect 1381 2106 1411 2128
rect 1459 2106 1489 2128
rect 1574 2116 1604 2144
rect 801 2045 831 2078
rect 299 1984 329 2011
rect 407 1984 422 2018
rect 478 1984 508 2006
rect 622 1984 652 2006
rect 708 1984 723 2018
rect 801 1984 831 2011
rect 879 2045 909 2078
rect 994 2066 1024 2088
rect 1266 2066 1296 2088
rect 1846 2116 1876 2144
rect 1961 2106 1991 2128
rect 2039 2106 2069 2128
rect 2154 2116 2184 2144
rect 1381 2045 1411 2078
rect 879 1984 909 2011
rect 987 1984 1002 2018
rect 1058 1984 1088 2006
rect 1202 1984 1232 2006
rect 1288 1984 1303 2018
rect 1381 1984 1411 2011
rect 1459 2045 1489 2078
rect 1574 2066 1604 2088
rect 1846 2066 1876 2088
rect 2426 2116 2456 2144
rect 2541 2106 2571 2128
rect 2619 2106 2649 2128
rect 2734 2116 2764 2144
rect 1961 2045 1991 2078
rect 1459 1984 1489 2011
rect 1567 1984 1582 2018
rect 1638 1984 1668 2006
rect 1782 1984 1812 2006
rect 1868 1984 1883 2018
rect 1961 1984 1991 2011
rect 2039 2045 2069 2078
rect 2154 2066 2184 2088
rect 2426 2066 2456 2088
rect 3006 2116 3036 2144
rect 3121 2106 3151 2128
rect 3199 2106 3229 2128
rect 3314 2116 3344 2144
rect 2541 2045 2571 2078
rect 2039 1984 2069 2011
rect 2147 1984 2162 2018
rect 2218 1984 2248 2006
rect 2362 1984 2392 2006
rect 2448 1984 2463 2018
rect 2541 1984 2571 2011
rect 2619 2045 2649 2078
rect 2734 2066 2764 2088
rect 3006 2066 3036 2088
rect 3586 2116 3616 2144
rect 3701 2106 3731 2128
rect 3779 2106 3809 2128
rect 3894 2116 3924 2144
rect 3121 2045 3151 2078
rect 2619 1984 2649 2011
rect 2727 1984 2742 2018
rect 2798 1984 2828 2006
rect 2942 1984 2972 2006
rect 3028 1984 3043 2018
rect 3121 1984 3151 2011
rect 3199 2045 3229 2078
rect 3314 2066 3344 2088
rect 3586 2066 3616 2088
rect 4166 2116 4196 2144
rect 4281 2106 4311 2128
rect 4359 2106 4389 2128
rect 4474 2116 4504 2144
rect 3701 2045 3731 2078
rect 3199 1984 3229 2011
rect 3307 1984 3322 2018
rect 3378 1984 3408 2006
rect 3522 1984 3552 2006
rect 3608 1984 3623 2018
rect 3701 1984 3731 2011
rect 3779 2045 3809 2078
rect 3894 2066 3924 2088
rect 4166 2066 4196 2088
rect 4746 2116 4776 2144
rect 4861 2106 4891 2128
rect 4939 2106 4969 2128
rect 5054 2116 5084 2144
rect 4281 2045 4311 2078
rect 3779 1984 3809 2011
rect 3887 1984 3902 2018
rect 3958 1984 3988 2006
rect 4102 1984 4132 2006
rect 4188 1984 4203 2018
rect 4281 1984 4311 2011
rect 4359 2045 4389 2078
rect 4474 2066 4504 2088
rect 4746 2066 4776 2088
rect 5326 2116 5356 2144
rect 5441 2106 5471 2128
rect 5519 2106 5549 2128
rect 5634 2116 5664 2144
rect 4861 2045 4891 2078
rect 4359 1984 4389 2011
rect 4467 1984 4482 2018
rect 4538 1984 4568 2006
rect 4682 1984 4712 2006
rect 4768 1984 4783 2018
rect 4861 1984 4891 2011
rect 4939 2045 4969 2078
rect 5054 2066 5084 2088
rect 5326 2066 5356 2088
rect 5906 2116 5936 2144
rect 6021 2106 6051 2128
rect 6099 2106 6129 2128
rect 6214 2116 6244 2144
rect 5441 2045 5471 2078
rect 4939 1984 4969 2011
rect 5047 1984 5062 2018
rect 5118 1984 5148 2006
rect 5262 1984 5292 2006
rect 5348 1984 5363 2018
rect 5441 1984 5471 2011
rect 5519 2045 5549 2078
rect 5634 2066 5664 2088
rect 5906 2066 5936 2088
rect 6486 2116 6516 2144
rect 6601 2106 6631 2128
rect 6679 2106 6709 2128
rect 6794 2116 6824 2144
rect 6021 2045 6051 2078
rect 5519 1984 5549 2011
rect 5627 1984 5642 2018
rect 5698 1984 5728 2006
rect 5842 1984 5872 2006
rect 5928 1984 5943 2018
rect 6021 1984 6051 2011
rect 6099 2045 6129 2078
rect 6214 2066 6244 2088
rect 6486 2066 6516 2088
rect 6601 2045 6631 2078
rect 6099 1984 6129 2011
rect 6207 1984 6222 2018
rect 6278 1984 6308 2006
rect 6422 1984 6452 2006
rect 6508 1984 6523 2018
rect 6601 1984 6631 2011
rect 6679 2045 6709 2078
rect 6794 2066 6824 2088
rect 6679 1984 6709 2011
rect 6787 1984 6802 2018
rect 6858 1984 6888 2006
rect 128 1970 158 1984
rect 392 1970 422 1984
rect 708 1970 738 1984
rect 972 1970 1002 1984
rect 1288 1970 1318 1984
rect 1552 1970 1582 1984
rect 1868 1970 1898 1984
rect 2132 1970 2162 1984
rect 2448 1970 2478 1984
rect 2712 1970 2742 1984
rect 3028 1970 3058 1984
rect 3292 1970 3322 1984
rect 3608 1970 3638 1984
rect 3872 1970 3902 1984
rect 4188 1970 4218 1984
rect 4452 1970 4482 1984
rect 4768 1970 4798 1984
rect 5032 1970 5062 1984
rect 5348 1970 5378 1984
rect 5612 1970 5642 1984
rect 5928 1970 5958 1984
rect 6192 1970 6222 1984
rect 6508 1970 6538 1984
rect 6772 1970 6802 1984
rect 42 1920 72 1942
rect 128 1920 158 1942
rect 221 1920 251 1942
rect 299 1920 329 1942
rect 392 1920 422 1942
rect 478 1920 508 1942
rect 622 1920 652 1942
rect 708 1920 738 1942
rect 801 1920 831 1942
rect 879 1920 909 1942
rect 972 1920 1002 1942
rect 1058 1920 1088 1942
rect 1202 1920 1232 1942
rect 1288 1920 1318 1942
rect 1381 1920 1411 1942
rect 1459 1920 1489 1942
rect 1552 1920 1582 1942
rect 1638 1920 1668 1942
rect 1782 1920 1812 1942
rect 1868 1920 1898 1942
rect 1961 1920 1991 1942
rect 2039 1920 2069 1942
rect 2132 1920 2162 1942
rect 2218 1920 2248 1942
rect 2362 1920 2392 1942
rect 2448 1920 2478 1942
rect 2541 1920 2571 1942
rect 2619 1920 2649 1942
rect 2712 1920 2742 1942
rect 2798 1920 2828 1942
rect 2942 1920 2972 1942
rect 3028 1920 3058 1942
rect 3121 1920 3151 1942
rect 3199 1920 3229 1942
rect 3292 1920 3322 1942
rect 3378 1920 3408 1942
rect 3522 1920 3552 1942
rect 3608 1920 3638 1942
rect 3701 1920 3731 1942
rect 3779 1920 3809 1942
rect 3872 1920 3902 1942
rect 3958 1920 3988 1942
rect 4102 1920 4132 1942
rect 4188 1920 4218 1942
rect 4281 1920 4311 1942
rect 4359 1920 4389 1942
rect 4452 1920 4482 1942
rect 4538 1920 4568 1942
rect 4682 1920 4712 1942
rect 4768 1920 4798 1942
rect 4861 1920 4891 1942
rect 4939 1920 4969 1942
rect 5032 1920 5062 1942
rect 5118 1920 5148 1942
rect 5262 1920 5292 1942
rect 5348 1920 5378 1942
rect 5441 1920 5471 1942
rect 5519 1920 5549 1942
rect 5612 1920 5642 1942
rect 5698 1920 5728 1942
rect 5842 1920 5872 1942
rect 5928 1920 5958 1942
rect 6021 1920 6051 1942
rect 6099 1920 6129 1942
rect 6192 1920 6222 1942
rect 6278 1920 6308 1942
rect 6422 1920 6452 1942
rect 6508 1920 6538 1942
rect 6601 1920 6631 1942
rect 6679 1920 6709 1942
rect 6772 1920 6802 1942
rect 6858 1920 6888 1942
rect -1 1874 6931 1904
rect 106 1846 136 1874
rect 221 1836 251 1858
rect 299 1836 329 1858
rect 414 1846 444 1874
rect 106 1796 136 1818
rect 686 1846 716 1874
rect 801 1836 831 1858
rect 879 1836 909 1858
rect 994 1846 1024 1874
rect 221 1775 251 1808
rect 42 1714 72 1736
rect 128 1714 143 1748
rect 221 1714 251 1741
rect 299 1775 329 1808
rect 414 1796 444 1818
rect 686 1796 716 1818
rect 1266 1846 1296 1874
rect 1381 1836 1411 1858
rect 1459 1836 1489 1858
rect 1574 1846 1604 1874
rect 801 1775 831 1808
rect 299 1714 329 1741
rect 407 1714 422 1748
rect 478 1714 508 1736
rect 622 1714 652 1736
rect 708 1714 723 1748
rect 801 1714 831 1741
rect 879 1775 909 1808
rect 994 1796 1024 1818
rect 1266 1796 1296 1818
rect 1846 1846 1876 1874
rect 1961 1836 1991 1858
rect 2039 1836 2069 1858
rect 2154 1846 2184 1874
rect 1381 1775 1411 1808
rect 879 1714 909 1741
rect 987 1714 1002 1748
rect 1058 1714 1088 1736
rect 1202 1714 1232 1736
rect 1288 1714 1303 1748
rect 1381 1714 1411 1741
rect 1459 1775 1489 1808
rect 1574 1796 1604 1818
rect 1846 1796 1876 1818
rect 2426 1846 2456 1874
rect 2541 1836 2571 1858
rect 2619 1836 2649 1858
rect 2734 1846 2764 1874
rect 1961 1775 1991 1808
rect 1459 1714 1489 1741
rect 1567 1714 1582 1748
rect 1638 1714 1668 1736
rect 1782 1714 1812 1736
rect 1868 1714 1883 1748
rect 1961 1714 1991 1741
rect 2039 1775 2069 1808
rect 2154 1796 2184 1818
rect 2426 1796 2456 1818
rect 3006 1846 3036 1874
rect 3121 1836 3151 1858
rect 3199 1836 3229 1858
rect 3314 1846 3344 1874
rect 2541 1775 2571 1808
rect 2039 1714 2069 1741
rect 2147 1714 2162 1748
rect 2218 1714 2248 1736
rect 2362 1714 2392 1736
rect 2448 1714 2463 1748
rect 2541 1714 2571 1741
rect 2619 1775 2649 1808
rect 2734 1796 2764 1818
rect 3006 1796 3036 1818
rect 3586 1846 3616 1874
rect 3701 1836 3731 1858
rect 3779 1836 3809 1858
rect 3894 1846 3924 1874
rect 3121 1775 3151 1808
rect 2619 1714 2649 1741
rect 2727 1714 2742 1748
rect 2798 1714 2828 1736
rect 2942 1714 2972 1736
rect 3028 1714 3043 1748
rect 3121 1714 3151 1741
rect 3199 1775 3229 1808
rect 3314 1796 3344 1818
rect 3586 1796 3616 1818
rect 4166 1846 4196 1874
rect 4281 1836 4311 1858
rect 4359 1836 4389 1858
rect 4474 1846 4504 1874
rect 3701 1775 3731 1808
rect 3199 1714 3229 1741
rect 3307 1714 3322 1748
rect 3378 1714 3408 1736
rect 3522 1714 3552 1736
rect 3608 1714 3623 1748
rect 3701 1714 3731 1741
rect 3779 1775 3809 1808
rect 3894 1796 3924 1818
rect 4166 1796 4196 1818
rect 4746 1846 4776 1874
rect 4861 1836 4891 1858
rect 4939 1836 4969 1858
rect 5054 1846 5084 1874
rect 4281 1775 4311 1808
rect 3779 1714 3809 1741
rect 3887 1714 3902 1748
rect 3958 1714 3988 1736
rect 4102 1714 4132 1736
rect 4188 1714 4203 1748
rect 4281 1714 4311 1741
rect 4359 1775 4389 1808
rect 4474 1796 4504 1818
rect 4746 1796 4776 1818
rect 5326 1846 5356 1874
rect 5441 1836 5471 1858
rect 5519 1836 5549 1858
rect 5634 1846 5664 1874
rect 4861 1775 4891 1808
rect 4359 1714 4389 1741
rect 4467 1714 4482 1748
rect 4538 1714 4568 1736
rect 4682 1714 4712 1736
rect 4768 1714 4783 1748
rect 4861 1714 4891 1741
rect 4939 1775 4969 1808
rect 5054 1796 5084 1818
rect 5326 1796 5356 1818
rect 5906 1846 5936 1874
rect 6021 1836 6051 1858
rect 6099 1836 6129 1858
rect 6214 1846 6244 1874
rect 5441 1775 5471 1808
rect 4939 1714 4969 1741
rect 5047 1714 5062 1748
rect 5118 1714 5148 1736
rect 5262 1714 5292 1736
rect 5348 1714 5363 1748
rect 5441 1714 5471 1741
rect 5519 1775 5549 1808
rect 5634 1796 5664 1818
rect 5906 1796 5936 1818
rect 6486 1846 6516 1874
rect 6601 1836 6631 1858
rect 6679 1836 6709 1858
rect 6794 1846 6824 1874
rect 6021 1775 6051 1808
rect 5519 1714 5549 1741
rect 5627 1714 5642 1748
rect 5698 1714 5728 1736
rect 5842 1714 5872 1736
rect 5928 1714 5943 1748
rect 6021 1714 6051 1741
rect 6099 1775 6129 1808
rect 6214 1796 6244 1818
rect 6486 1796 6516 1818
rect 6601 1775 6631 1808
rect 6099 1714 6129 1741
rect 6207 1714 6222 1748
rect 6278 1714 6308 1736
rect 6422 1714 6452 1736
rect 6508 1714 6523 1748
rect 6601 1714 6631 1741
rect 6679 1775 6709 1808
rect 6794 1796 6824 1818
rect 6679 1714 6709 1741
rect 6787 1714 6802 1748
rect 6858 1714 6888 1736
rect 128 1700 158 1714
rect 392 1700 422 1714
rect 708 1700 738 1714
rect 972 1700 1002 1714
rect 1288 1700 1318 1714
rect 1552 1700 1582 1714
rect 1868 1700 1898 1714
rect 2132 1700 2162 1714
rect 2448 1700 2478 1714
rect 2712 1700 2742 1714
rect 3028 1700 3058 1714
rect 3292 1700 3322 1714
rect 3608 1700 3638 1714
rect 3872 1700 3902 1714
rect 4188 1700 4218 1714
rect 4452 1700 4482 1714
rect 4768 1700 4798 1714
rect 5032 1700 5062 1714
rect 5348 1700 5378 1714
rect 5612 1700 5642 1714
rect 5928 1700 5958 1714
rect 6192 1700 6222 1714
rect 6508 1700 6538 1714
rect 6772 1700 6802 1714
rect 42 1650 72 1672
rect 128 1650 158 1672
rect 221 1650 251 1672
rect 299 1650 329 1672
rect 392 1650 422 1672
rect 478 1650 508 1672
rect 622 1650 652 1672
rect 708 1650 738 1672
rect 801 1650 831 1672
rect 879 1650 909 1672
rect 972 1650 1002 1672
rect 1058 1650 1088 1672
rect 1202 1650 1232 1672
rect 1288 1650 1318 1672
rect 1381 1650 1411 1672
rect 1459 1650 1489 1672
rect 1552 1650 1582 1672
rect 1638 1650 1668 1672
rect 1782 1650 1812 1672
rect 1868 1650 1898 1672
rect 1961 1650 1991 1672
rect 2039 1650 2069 1672
rect 2132 1650 2162 1672
rect 2218 1650 2248 1672
rect 2362 1650 2392 1672
rect 2448 1650 2478 1672
rect 2541 1650 2571 1672
rect 2619 1650 2649 1672
rect 2712 1650 2742 1672
rect 2798 1650 2828 1672
rect 2942 1650 2972 1672
rect 3028 1650 3058 1672
rect 3121 1650 3151 1672
rect 3199 1650 3229 1672
rect 3292 1650 3322 1672
rect 3378 1650 3408 1672
rect 3522 1650 3552 1672
rect 3608 1650 3638 1672
rect 3701 1650 3731 1672
rect 3779 1650 3809 1672
rect 3872 1650 3902 1672
rect 3958 1650 3988 1672
rect 4102 1650 4132 1672
rect 4188 1650 4218 1672
rect 4281 1650 4311 1672
rect 4359 1650 4389 1672
rect 4452 1650 4482 1672
rect 4538 1650 4568 1672
rect 4682 1650 4712 1672
rect 4768 1650 4798 1672
rect 4861 1650 4891 1672
rect 4939 1650 4969 1672
rect 5032 1650 5062 1672
rect 5118 1650 5148 1672
rect 5262 1650 5292 1672
rect 5348 1650 5378 1672
rect 5441 1650 5471 1672
rect 5519 1650 5549 1672
rect 5612 1650 5642 1672
rect 5698 1650 5728 1672
rect 5842 1650 5872 1672
rect 5928 1650 5958 1672
rect 6021 1650 6051 1672
rect 6099 1650 6129 1672
rect 6192 1650 6222 1672
rect 6278 1650 6308 1672
rect 6422 1650 6452 1672
rect 6508 1650 6538 1672
rect 6601 1650 6631 1672
rect 6679 1650 6709 1672
rect 6772 1650 6802 1672
rect 6858 1650 6888 1672
rect -1 1604 6931 1634
rect 106 1576 136 1604
rect 221 1566 251 1588
rect 299 1566 329 1588
rect 414 1576 444 1604
rect 106 1526 136 1548
rect 686 1576 716 1604
rect 801 1566 831 1588
rect 879 1566 909 1588
rect 994 1576 1024 1604
rect 221 1505 251 1538
rect 42 1444 72 1466
rect 128 1444 143 1478
rect 221 1444 251 1471
rect 299 1505 329 1538
rect 414 1526 444 1548
rect 686 1526 716 1548
rect 1266 1576 1296 1604
rect 1381 1566 1411 1588
rect 1459 1566 1489 1588
rect 1574 1576 1604 1604
rect 801 1505 831 1538
rect 299 1444 329 1471
rect 407 1444 422 1478
rect 478 1444 508 1466
rect 622 1444 652 1466
rect 708 1444 723 1478
rect 801 1444 831 1471
rect 879 1505 909 1538
rect 994 1526 1024 1548
rect 1266 1526 1296 1548
rect 1846 1576 1876 1604
rect 1961 1566 1991 1588
rect 2039 1566 2069 1588
rect 2154 1576 2184 1604
rect 1381 1505 1411 1538
rect 879 1444 909 1471
rect 987 1444 1002 1478
rect 1058 1444 1088 1466
rect 1202 1444 1232 1466
rect 1288 1444 1303 1478
rect 1381 1444 1411 1471
rect 1459 1505 1489 1538
rect 1574 1526 1604 1548
rect 1846 1526 1876 1548
rect 2426 1576 2456 1604
rect 2541 1566 2571 1588
rect 2619 1566 2649 1588
rect 2734 1576 2764 1604
rect 1961 1505 1991 1538
rect 1459 1444 1489 1471
rect 1567 1444 1582 1478
rect 1638 1444 1668 1466
rect 1782 1444 1812 1466
rect 1868 1444 1883 1478
rect 1961 1444 1991 1471
rect 2039 1505 2069 1538
rect 2154 1526 2184 1548
rect 2426 1526 2456 1548
rect 3006 1576 3036 1604
rect 3121 1566 3151 1588
rect 3199 1566 3229 1588
rect 3314 1576 3344 1604
rect 2541 1505 2571 1538
rect 2039 1444 2069 1471
rect 2147 1444 2162 1478
rect 2218 1444 2248 1466
rect 2362 1444 2392 1466
rect 2448 1444 2463 1478
rect 2541 1444 2571 1471
rect 2619 1505 2649 1538
rect 2734 1526 2764 1548
rect 3006 1526 3036 1548
rect 3586 1576 3616 1604
rect 3701 1566 3731 1588
rect 3779 1566 3809 1588
rect 3894 1576 3924 1604
rect 3121 1505 3151 1538
rect 2619 1444 2649 1471
rect 2727 1444 2742 1478
rect 2798 1444 2828 1466
rect 2942 1444 2972 1466
rect 3028 1444 3043 1478
rect 3121 1444 3151 1471
rect 3199 1505 3229 1538
rect 3314 1526 3344 1548
rect 3586 1526 3616 1548
rect 4166 1576 4196 1604
rect 4281 1566 4311 1588
rect 4359 1566 4389 1588
rect 4474 1576 4504 1604
rect 3701 1505 3731 1538
rect 3199 1444 3229 1471
rect 3307 1444 3322 1478
rect 3378 1444 3408 1466
rect 3522 1444 3552 1466
rect 3608 1444 3623 1478
rect 3701 1444 3731 1471
rect 3779 1505 3809 1538
rect 3894 1526 3924 1548
rect 4166 1526 4196 1548
rect 4746 1576 4776 1604
rect 4861 1566 4891 1588
rect 4939 1566 4969 1588
rect 5054 1576 5084 1604
rect 4281 1505 4311 1538
rect 3779 1444 3809 1471
rect 3887 1444 3902 1478
rect 3958 1444 3988 1466
rect 4102 1444 4132 1466
rect 4188 1444 4203 1478
rect 4281 1444 4311 1471
rect 4359 1505 4389 1538
rect 4474 1526 4504 1548
rect 4746 1526 4776 1548
rect 5326 1576 5356 1604
rect 5441 1566 5471 1588
rect 5519 1566 5549 1588
rect 5634 1576 5664 1604
rect 4861 1505 4891 1538
rect 4359 1444 4389 1471
rect 4467 1444 4482 1478
rect 4538 1444 4568 1466
rect 4682 1444 4712 1466
rect 4768 1444 4783 1478
rect 4861 1444 4891 1471
rect 4939 1505 4969 1538
rect 5054 1526 5084 1548
rect 5326 1526 5356 1548
rect 5906 1576 5936 1604
rect 6021 1566 6051 1588
rect 6099 1566 6129 1588
rect 6214 1576 6244 1604
rect 5441 1505 5471 1538
rect 4939 1444 4969 1471
rect 5047 1444 5062 1478
rect 5118 1444 5148 1466
rect 5262 1444 5292 1466
rect 5348 1444 5363 1478
rect 5441 1444 5471 1471
rect 5519 1505 5549 1538
rect 5634 1526 5664 1548
rect 5906 1526 5936 1548
rect 6486 1576 6516 1604
rect 6601 1566 6631 1588
rect 6679 1566 6709 1588
rect 6794 1576 6824 1604
rect 6021 1505 6051 1538
rect 5519 1444 5549 1471
rect 5627 1444 5642 1478
rect 5698 1444 5728 1466
rect 5842 1444 5872 1466
rect 5928 1444 5943 1478
rect 6021 1444 6051 1471
rect 6099 1505 6129 1538
rect 6214 1526 6244 1548
rect 6486 1526 6516 1548
rect 6601 1505 6631 1538
rect 6099 1444 6129 1471
rect 6207 1444 6222 1478
rect 6278 1444 6308 1466
rect 6422 1444 6452 1466
rect 6508 1444 6523 1478
rect 6601 1444 6631 1471
rect 6679 1505 6709 1538
rect 6794 1526 6824 1548
rect 6679 1444 6709 1471
rect 6787 1444 6802 1478
rect 6858 1444 6888 1466
rect 128 1430 158 1444
rect 392 1430 422 1444
rect 708 1430 738 1444
rect 972 1430 1002 1444
rect 1288 1430 1318 1444
rect 1552 1430 1582 1444
rect 1868 1430 1898 1444
rect 2132 1430 2162 1444
rect 2448 1430 2478 1444
rect 2712 1430 2742 1444
rect 3028 1430 3058 1444
rect 3292 1430 3322 1444
rect 3608 1430 3638 1444
rect 3872 1430 3902 1444
rect 4188 1430 4218 1444
rect 4452 1430 4482 1444
rect 4768 1430 4798 1444
rect 5032 1430 5062 1444
rect 5348 1430 5378 1444
rect 5612 1430 5642 1444
rect 5928 1430 5958 1444
rect 6192 1430 6222 1444
rect 6508 1430 6538 1444
rect 6772 1430 6802 1444
rect 42 1380 72 1402
rect 128 1380 158 1402
rect 221 1380 251 1402
rect 299 1380 329 1402
rect 392 1380 422 1402
rect 478 1380 508 1402
rect 622 1380 652 1402
rect 708 1380 738 1402
rect 801 1380 831 1402
rect 879 1380 909 1402
rect 972 1380 1002 1402
rect 1058 1380 1088 1402
rect 1202 1380 1232 1402
rect 1288 1380 1318 1402
rect 1381 1380 1411 1402
rect 1459 1380 1489 1402
rect 1552 1380 1582 1402
rect 1638 1380 1668 1402
rect 1782 1380 1812 1402
rect 1868 1380 1898 1402
rect 1961 1380 1991 1402
rect 2039 1380 2069 1402
rect 2132 1380 2162 1402
rect 2218 1380 2248 1402
rect 2362 1380 2392 1402
rect 2448 1380 2478 1402
rect 2541 1380 2571 1402
rect 2619 1380 2649 1402
rect 2712 1380 2742 1402
rect 2798 1380 2828 1402
rect 2942 1380 2972 1402
rect 3028 1380 3058 1402
rect 3121 1380 3151 1402
rect 3199 1380 3229 1402
rect 3292 1380 3322 1402
rect 3378 1380 3408 1402
rect 3522 1380 3552 1402
rect 3608 1380 3638 1402
rect 3701 1380 3731 1402
rect 3779 1380 3809 1402
rect 3872 1380 3902 1402
rect 3958 1380 3988 1402
rect 4102 1380 4132 1402
rect 4188 1380 4218 1402
rect 4281 1380 4311 1402
rect 4359 1380 4389 1402
rect 4452 1380 4482 1402
rect 4538 1380 4568 1402
rect 4682 1380 4712 1402
rect 4768 1380 4798 1402
rect 4861 1380 4891 1402
rect 4939 1380 4969 1402
rect 5032 1380 5062 1402
rect 5118 1380 5148 1402
rect 5262 1380 5292 1402
rect 5348 1380 5378 1402
rect 5441 1380 5471 1402
rect 5519 1380 5549 1402
rect 5612 1380 5642 1402
rect 5698 1380 5728 1402
rect 5842 1380 5872 1402
rect 5928 1380 5958 1402
rect 6021 1380 6051 1402
rect 6099 1380 6129 1402
rect 6192 1380 6222 1402
rect 6278 1380 6308 1402
rect 6422 1380 6452 1402
rect 6508 1380 6538 1402
rect 6601 1380 6631 1402
rect 6679 1380 6709 1402
rect 6772 1380 6802 1402
rect 6858 1380 6888 1402
rect -1 1334 6931 1364
rect 106 1306 136 1334
rect 221 1296 251 1318
rect 299 1296 329 1318
rect 414 1306 444 1334
rect 106 1256 136 1278
rect 686 1306 716 1334
rect 801 1296 831 1318
rect 879 1296 909 1318
rect 994 1306 1024 1334
rect 221 1235 251 1268
rect 42 1174 72 1196
rect 128 1174 143 1208
rect 221 1174 251 1201
rect 299 1235 329 1268
rect 414 1256 444 1278
rect 686 1256 716 1278
rect 1266 1306 1296 1334
rect 1381 1296 1411 1318
rect 1459 1296 1489 1318
rect 1574 1306 1604 1334
rect 801 1235 831 1268
rect 299 1174 329 1201
rect 407 1174 422 1208
rect 478 1174 508 1196
rect 622 1174 652 1196
rect 708 1174 723 1208
rect 801 1174 831 1201
rect 879 1235 909 1268
rect 994 1256 1024 1278
rect 1266 1256 1296 1278
rect 1846 1306 1876 1334
rect 1961 1296 1991 1318
rect 2039 1296 2069 1318
rect 2154 1306 2184 1334
rect 1381 1235 1411 1268
rect 879 1174 909 1201
rect 987 1174 1002 1208
rect 1058 1174 1088 1196
rect 1202 1174 1232 1196
rect 1288 1174 1303 1208
rect 1381 1174 1411 1201
rect 1459 1235 1489 1268
rect 1574 1256 1604 1278
rect 1846 1256 1876 1278
rect 2426 1306 2456 1334
rect 2541 1296 2571 1318
rect 2619 1296 2649 1318
rect 2734 1306 2764 1334
rect 1961 1235 1991 1268
rect 1459 1174 1489 1201
rect 1567 1174 1582 1208
rect 1638 1174 1668 1196
rect 1782 1174 1812 1196
rect 1868 1174 1883 1208
rect 1961 1174 1991 1201
rect 2039 1235 2069 1268
rect 2154 1256 2184 1278
rect 2426 1256 2456 1278
rect 3006 1306 3036 1334
rect 3121 1296 3151 1318
rect 3199 1296 3229 1318
rect 3314 1306 3344 1334
rect 2541 1235 2571 1268
rect 2039 1174 2069 1201
rect 2147 1174 2162 1208
rect 2218 1174 2248 1196
rect 2362 1174 2392 1196
rect 2448 1174 2463 1208
rect 2541 1174 2571 1201
rect 2619 1235 2649 1268
rect 2734 1256 2764 1278
rect 3006 1256 3036 1278
rect 3586 1306 3616 1334
rect 3701 1296 3731 1318
rect 3779 1296 3809 1318
rect 3894 1306 3924 1334
rect 3121 1235 3151 1268
rect 2619 1174 2649 1201
rect 2727 1174 2742 1208
rect 2798 1174 2828 1196
rect 2942 1174 2972 1196
rect 3028 1174 3043 1208
rect 3121 1174 3151 1201
rect 3199 1235 3229 1268
rect 3314 1256 3344 1278
rect 3586 1256 3616 1278
rect 4166 1306 4196 1334
rect 4281 1296 4311 1318
rect 4359 1296 4389 1318
rect 4474 1306 4504 1334
rect 3701 1235 3731 1268
rect 3199 1174 3229 1201
rect 3307 1174 3322 1208
rect 3378 1174 3408 1196
rect 3522 1174 3552 1196
rect 3608 1174 3623 1208
rect 3701 1174 3731 1201
rect 3779 1235 3809 1268
rect 3894 1256 3924 1278
rect 4166 1256 4196 1278
rect 4746 1306 4776 1334
rect 4861 1296 4891 1318
rect 4939 1296 4969 1318
rect 5054 1306 5084 1334
rect 4281 1235 4311 1268
rect 3779 1174 3809 1201
rect 3887 1174 3902 1208
rect 3958 1174 3988 1196
rect 4102 1174 4132 1196
rect 4188 1174 4203 1208
rect 4281 1174 4311 1201
rect 4359 1235 4389 1268
rect 4474 1256 4504 1278
rect 4746 1256 4776 1278
rect 5326 1306 5356 1334
rect 5441 1296 5471 1318
rect 5519 1296 5549 1318
rect 5634 1306 5664 1334
rect 4861 1235 4891 1268
rect 4359 1174 4389 1201
rect 4467 1174 4482 1208
rect 4538 1174 4568 1196
rect 4682 1174 4712 1196
rect 4768 1174 4783 1208
rect 4861 1174 4891 1201
rect 4939 1235 4969 1268
rect 5054 1256 5084 1278
rect 5326 1256 5356 1278
rect 5906 1306 5936 1334
rect 6021 1296 6051 1318
rect 6099 1296 6129 1318
rect 6214 1306 6244 1334
rect 5441 1235 5471 1268
rect 4939 1174 4969 1201
rect 5047 1174 5062 1208
rect 5118 1174 5148 1196
rect 5262 1174 5292 1196
rect 5348 1174 5363 1208
rect 5441 1174 5471 1201
rect 5519 1235 5549 1268
rect 5634 1256 5664 1278
rect 5906 1256 5936 1278
rect 6486 1306 6516 1334
rect 6601 1296 6631 1318
rect 6679 1296 6709 1318
rect 6794 1306 6824 1334
rect 6021 1235 6051 1268
rect 5519 1174 5549 1201
rect 5627 1174 5642 1208
rect 5698 1174 5728 1196
rect 5842 1174 5872 1196
rect 5928 1174 5943 1208
rect 6021 1174 6051 1201
rect 6099 1235 6129 1268
rect 6214 1256 6244 1278
rect 6486 1256 6516 1278
rect 6601 1235 6631 1268
rect 6099 1174 6129 1201
rect 6207 1174 6222 1208
rect 6278 1174 6308 1196
rect 6422 1174 6452 1196
rect 6508 1174 6523 1208
rect 6601 1174 6631 1201
rect 6679 1235 6709 1268
rect 6794 1256 6824 1278
rect 6679 1174 6709 1201
rect 6787 1174 6802 1208
rect 6858 1174 6888 1196
rect 128 1160 158 1174
rect 392 1160 422 1174
rect 708 1160 738 1174
rect 972 1160 1002 1174
rect 1288 1160 1318 1174
rect 1552 1160 1582 1174
rect 1868 1160 1898 1174
rect 2132 1160 2162 1174
rect 2448 1160 2478 1174
rect 2712 1160 2742 1174
rect 3028 1160 3058 1174
rect 3292 1160 3322 1174
rect 3608 1160 3638 1174
rect 3872 1160 3902 1174
rect 4188 1160 4218 1174
rect 4452 1160 4482 1174
rect 4768 1160 4798 1174
rect 5032 1160 5062 1174
rect 5348 1160 5378 1174
rect 5612 1160 5642 1174
rect 5928 1160 5958 1174
rect 6192 1160 6222 1174
rect 6508 1160 6538 1174
rect 6772 1160 6802 1174
rect 42 1110 72 1132
rect 128 1110 158 1132
rect 221 1110 251 1132
rect 299 1110 329 1132
rect 392 1110 422 1132
rect 478 1110 508 1132
rect 622 1110 652 1132
rect 708 1110 738 1132
rect 801 1110 831 1132
rect 879 1110 909 1132
rect 972 1110 1002 1132
rect 1058 1110 1088 1132
rect 1202 1110 1232 1132
rect 1288 1110 1318 1132
rect 1381 1110 1411 1132
rect 1459 1110 1489 1132
rect 1552 1110 1582 1132
rect 1638 1110 1668 1132
rect 1782 1110 1812 1132
rect 1868 1110 1898 1132
rect 1961 1110 1991 1132
rect 2039 1110 2069 1132
rect 2132 1110 2162 1132
rect 2218 1110 2248 1132
rect 2362 1110 2392 1132
rect 2448 1110 2478 1132
rect 2541 1110 2571 1132
rect 2619 1110 2649 1132
rect 2712 1110 2742 1132
rect 2798 1110 2828 1132
rect 2942 1110 2972 1132
rect 3028 1110 3058 1132
rect 3121 1110 3151 1132
rect 3199 1110 3229 1132
rect 3292 1110 3322 1132
rect 3378 1110 3408 1132
rect 3522 1110 3552 1132
rect 3608 1110 3638 1132
rect 3701 1110 3731 1132
rect 3779 1110 3809 1132
rect 3872 1110 3902 1132
rect 3958 1110 3988 1132
rect 4102 1110 4132 1132
rect 4188 1110 4218 1132
rect 4281 1110 4311 1132
rect 4359 1110 4389 1132
rect 4452 1110 4482 1132
rect 4538 1110 4568 1132
rect 4682 1110 4712 1132
rect 4768 1110 4798 1132
rect 4861 1110 4891 1132
rect 4939 1110 4969 1132
rect 5032 1110 5062 1132
rect 5118 1110 5148 1132
rect 5262 1110 5292 1132
rect 5348 1110 5378 1132
rect 5441 1110 5471 1132
rect 5519 1110 5549 1132
rect 5612 1110 5642 1132
rect 5698 1110 5728 1132
rect 5842 1110 5872 1132
rect 5928 1110 5958 1132
rect 6021 1110 6051 1132
rect 6099 1110 6129 1132
rect 6192 1110 6222 1132
rect 6278 1110 6308 1132
rect 6422 1110 6452 1132
rect 6508 1110 6538 1132
rect 6601 1110 6631 1132
rect 6679 1110 6709 1132
rect 6772 1110 6802 1132
rect 6858 1110 6888 1132
rect -1 1064 6931 1094
rect 106 1036 136 1064
rect 221 1026 251 1048
rect 299 1026 329 1048
rect 414 1036 444 1064
rect 106 986 136 1008
rect 686 1036 716 1064
rect 801 1026 831 1048
rect 879 1026 909 1048
rect 994 1036 1024 1064
rect 221 965 251 998
rect 42 904 72 926
rect 128 904 143 938
rect 221 904 251 931
rect 299 965 329 998
rect 414 986 444 1008
rect 686 986 716 1008
rect 1266 1036 1296 1064
rect 1381 1026 1411 1048
rect 1459 1026 1489 1048
rect 1574 1036 1604 1064
rect 801 965 831 998
rect 299 904 329 931
rect 407 904 422 938
rect 478 904 508 926
rect 622 904 652 926
rect 708 904 723 938
rect 801 904 831 931
rect 879 965 909 998
rect 994 986 1024 1008
rect 1266 986 1296 1008
rect 1846 1036 1876 1064
rect 1961 1026 1991 1048
rect 2039 1026 2069 1048
rect 2154 1036 2184 1064
rect 1381 965 1411 998
rect 879 904 909 931
rect 987 904 1002 938
rect 1058 904 1088 926
rect 1202 904 1232 926
rect 1288 904 1303 938
rect 1381 904 1411 931
rect 1459 965 1489 998
rect 1574 986 1604 1008
rect 1846 986 1876 1008
rect 2426 1036 2456 1064
rect 2541 1026 2571 1048
rect 2619 1026 2649 1048
rect 2734 1036 2764 1064
rect 1961 965 1991 998
rect 1459 904 1489 931
rect 1567 904 1582 938
rect 1638 904 1668 926
rect 1782 904 1812 926
rect 1868 904 1883 938
rect 1961 904 1991 931
rect 2039 965 2069 998
rect 2154 986 2184 1008
rect 2426 986 2456 1008
rect 3006 1036 3036 1064
rect 3121 1026 3151 1048
rect 3199 1026 3229 1048
rect 3314 1036 3344 1064
rect 2541 965 2571 998
rect 2039 904 2069 931
rect 2147 904 2162 938
rect 2218 904 2248 926
rect 2362 904 2392 926
rect 2448 904 2463 938
rect 2541 904 2571 931
rect 2619 965 2649 998
rect 2734 986 2764 1008
rect 3006 986 3036 1008
rect 3586 1036 3616 1064
rect 3701 1026 3731 1048
rect 3779 1026 3809 1048
rect 3894 1036 3924 1064
rect 3121 965 3151 998
rect 2619 904 2649 931
rect 2727 904 2742 938
rect 2798 904 2828 926
rect 2942 904 2972 926
rect 3028 904 3043 938
rect 3121 904 3151 931
rect 3199 965 3229 998
rect 3314 986 3344 1008
rect 3586 986 3616 1008
rect 4166 1036 4196 1064
rect 4281 1026 4311 1048
rect 4359 1026 4389 1048
rect 4474 1036 4504 1064
rect 3701 965 3731 998
rect 3199 904 3229 931
rect 3307 904 3322 938
rect 3378 904 3408 926
rect 3522 904 3552 926
rect 3608 904 3623 938
rect 3701 904 3731 931
rect 3779 965 3809 998
rect 3894 986 3924 1008
rect 4166 986 4196 1008
rect 4746 1036 4776 1064
rect 4861 1026 4891 1048
rect 4939 1026 4969 1048
rect 5054 1036 5084 1064
rect 4281 965 4311 998
rect 3779 904 3809 931
rect 3887 904 3902 938
rect 3958 904 3988 926
rect 4102 904 4132 926
rect 4188 904 4203 938
rect 4281 904 4311 931
rect 4359 965 4389 998
rect 4474 986 4504 1008
rect 4746 986 4776 1008
rect 5326 1036 5356 1064
rect 5441 1026 5471 1048
rect 5519 1026 5549 1048
rect 5634 1036 5664 1064
rect 4861 965 4891 998
rect 4359 904 4389 931
rect 4467 904 4482 938
rect 4538 904 4568 926
rect 4682 904 4712 926
rect 4768 904 4783 938
rect 4861 904 4891 931
rect 4939 965 4969 998
rect 5054 986 5084 1008
rect 5326 986 5356 1008
rect 5906 1036 5936 1064
rect 6021 1026 6051 1048
rect 6099 1026 6129 1048
rect 6214 1036 6244 1064
rect 5441 965 5471 998
rect 4939 904 4969 931
rect 5047 904 5062 938
rect 5118 904 5148 926
rect 5262 904 5292 926
rect 5348 904 5363 938
rect 5441 904 5471 931
rect 5519 965 5549 998
rect 5634 986 5664 1008
rect 5906 986 5936 1008
rect 6486 1036 6516 1064
rect 6601 1026 6631 1048
rect 6679 1026 6709 1048
rect 6794 1036 6824 1064
rect 6021 965 6051 998
rect 5519 904 5549 931
rect 5627 904 5642 938
rect 5698 904 5728 926
rect 5842 904 5872 926
rect 5928 904 5943 938
rect 6021 904 6051 931
rect 6099 965 6129 998
rect 6214 986 6244 1008
rect 6486 986 6516 1008
rect 6601 965 6631 998
rect 6099 904 6129 931
rect 6207 904 6222 938
rect 6278 904 6308 926
rect 6422 904 6452 926
rect 6508 904 6523 938
rect 6601 904 6631 931
rect 6679 965 6709 998
rect 6794 986 6824 1008
rect 6679 904 6709 931
rect 6787 904 6802 938
rect 6858 904 6888 926
rect 128 890 158 904
rect 392 890 422 904
rect 708 890 738 904
rect 972 890 1002 904
rect 1288 890 1318 904
rect 1552 890 1582 904
rect 1868 890 1898 904
rect 2132 890 2162 904
rect 2448 890 2478 904
rect 2712 890 2742 904
rect 3028 890 3058 904
rect 3292 890 3322 904
rect 3608 890 3638 904
rect 3872 890 3902 904
rect 4188 890 4218 904
rect 4452 890 4482 904
rect 4768 890 4798 904
rect 5032 890 5062 904
rect 5348 890 5378 904
rect 5612 890 5642 904
rect 5928 890 5958 904
rect 6192 890 6222 904
rect 6508 890 6538 904
rect 6772 890 6802 904
rect 42 840 72 862
rect 128 840 158 862
rect 221 840 251 862
rect 299 840 329 862
rect 392 840 422 862
rect 478 840 508 862
rect 622 840 652 862
rect 708 840 738 862
rect 801 840 831 862
rect 879 840 909 862
rect 972 840 1002 862
rect 1058 840 1088 862
rect 1202 840 1232 862
rect 1288 840 1318 862
rect 1381 840 1411 862
rect 1459 840 1489 862
rect 1552 840 1582 862
rect 1638 840 1668 862
rect 1782 840 1812 862
rect 1868 840 1898 862
rect 1961 840 1991 862
rect 2039 840 2069 862
rect 2132 840 2162 862
rect 2218 840 2248 862
rect 2362 840 2392 862
rect 2448 840 2478 862
rect 2541 840 2571 862
rect 2619 840 2649 862
rect 2712 840 2742 862
rect 2798 840 2828 862
rect 2942 840 2972 862
rect 3028 840 3058 862
rect 3121 840 3151 862
rect 3199 840 3229 862
rect 3292 840 3322 862
rect 3378 840 3408 862
rect 3522 840 3552 862
rect 3608 840 3638 862
rect 3701 840 3731 862
rect 3779 840 3809 862
rect 3872 840 3902 862
rect 3958 840 3988 862
rect 4102 840 4132 862
rect 4188 840 4218 862
rect 4281 840 4311 862
rect 4359 840 4389 862
rect 4452 840 4482 862
rect 4538 840 4568 862
rect 4682 840 4712 862
rect 4768 840 4798 862
rect 4861 840 4891 862
rect 4939 840 4969 862
rect 5032 840 5062 862
rect 5118 840 5148 862
rect 5262 840 5292 862
rect 5348 840 5378 862
rect 5441 840 5471 862
rect 5519 840 5549 862
rect 5612 840 5642 862
rect 5698 840 5728 862
rect 5842 840 5872 862
rect 5928 840 5958 862
rect 6021 840 6051 862
rect 6099 840 6129 862
rect 6192 840 6222 862
rect 6278 840 6308 862
rect 6422 840 6452 862
rect 6508 840 6538 862
rect 6601 840 6631 862
rect 6679 840 6709 862
rect 6772 840 6802 862
rect 6858 840 6888 862
rect -1 794 6931 824
rect 106 766 136 794
rect 221 756 251 778
rect 299 756 329 778
rect 414 766 444 794
rect 106 716 136 738
rect 686 766 716 794
rect 801 756 831 778
rect 879 756 909 778
rect 994 766 1024 794
rect 221 695 251 728
rect 42 634 72 656
rect 128 634 143 668
rect 221 634 251 661
rect 299 695 329 728
rect 414 716 444 738
rect 686 716 716 738
rect 1266 766 1296 794
rect 1381 756 1411 778
rect 1459 756 1489 778
rect 1574 766 1604 794
rect 801 695 831 728
rect 299 634 329 661
rect 407 634 422 668
rect 478 634 508 656
rect 622 634 652 656
rect 708 634 723 668
rect 801 634 831 661
rect 879 695 909 728
rect 994 716 1024 738
rect 1266 716 1296 738
rect 1846 766 1876 794
rect 1961 756 1991 778
rect 2039 756 2069 778
rect 2154 766 2184 794
rect 1381 695 1411 728
rect 879 634 909 661
rect 987 634 1002 668
rect 1058 634 1088 656
rect 1202 634 1232 656
rect 1288 634 1303 668
rect 1381 634 1411 661
rect 1459 695 1489 728
rect 1574 716 1604 738
rect 1846 716 1876 738
rect 2426 766 2456 794
rect 2541 756 2571 778
rect 2619 756 2649 778
rect 2734 766 2764 794
rect 1961 695 1991 728
rect 1459 634 1489 661
rect 1567 634 1582 668
rect 1638 634 1668 656
rect 1782 634 1812 656
rect 1868 634 1883 668
rect 1961 634 1991 661
rect 2039 695 2069 728
rect 2154 716 2184 738
rect 2426 716 2456 738
rect 3006 766 3036 794
rect 3121 756 3151 778
rect 3199 756 3229 778
rect 3314 766 3344 794
rect 2541 695 2571 728
rect 2039 634 2069 661
rect 2147 634 2162 668
rect 2218 634 2248 656
rect 2362 634 2392 656
rect 2448 634 2463 668
rect 2541 634 2571 661
rect 2619 695 2649 728
rect 2734 716 2764 738
rect 3006 716 3036 738
rect 3586 766 3616 794
rect 3701 756 3731 778
rect 3779 756 3809 778
rect 3894 766 3924 794
rect 3121 695 3151 728
rect 2619 634 2649 661
rect 2727 634 2742 668
rect 2798 634 2828 656
rect 2942 634 2972 656
rect 3028 634 3043 668
rect 3121 634 3151 661
rect 3199 695 3229 728
rect 3314 716 3344 738
rect 3586 716 3616 738
rect 4166 766 4196 794
rect 4281 756 4311 778
rect 4359 756 4389 778
rect 4474 766 4504 794
rect 3701 695 3731 728
rect 3199 634 3229 661
rect 3307 634 3322 668
rect 3378 634 3408 656
rect 3522 634 3552 656
rect 3608 634 3623 668
rect 3701 634 3731 661
rect 3779 695 3809 728
rect 3894 716 3924 738
rect 4166 716 4196 738
rect 4746 766 4776 794
rect 4861 756 4891 778
rect 4939 756 4969 778
rect 5054 766 5084 794
rect 4281 695 4311 728
rect 3779 634 3809 661
rect 3887 634 3902 668
rect 3958 634 3988 656
rect 4102 634 4132 656
rect 4188 634 4203 668
rect 4281 634 4311 661
rect 4359 695 4389 728
rect 4474 716 4504 738
rect 4746 716 4776 738
rect 5326 766 5356 794
rect 5441 756 5471 778
rect 5519 756 5549 778
rect 5634 766 5664 794
rect 4861 695 4891 728
rect 4359 634 4389 661
rect 4467 634 4482 668
rect 4538 634 4568 656
rect 4682 634 4712 656
rect 4768 634 4783 668
rect 4861 634 4891 661
rect 4939 695 4969 728
rect 5054 716 5084 738
rect 5326 716 5356 738
rect 5906 766 5936 794
rect 6021 756 6051 778
rect 6099 756 6129 778
rect 6214 766 6244 794
rect 5441 695 5471 728
rect 4939 634 4969 661
rect 5047 634 5062 668
rect 5118 634 5148 656
rect 5262 634 5292 656
rect 5348 634 5363 668
rect 5441 634 5471 661
rect 5519 695 5549 728
rect 5634 716 5664 738
rect 5906 716 5936 738
rect 6486 766 6516 794
rect 6601 756 6631 778
rect 6679 756 6709 778
rect 6794 766 6824 794
rect 6021 695 6051 728
rect 5519 634 5549 661
rect 5627 634 5642 668
rect 5698 634 5728 656
rect 5842 634 5872 656
rect 5928 634 5943 668
rect 6021 634 6051 661
rect 6099 695 6129 728
rect 6214 716 6244 738
rect 6486 716 6516 738
rect 6601 695 6631 728
rect 6099 634 6129 661
rect 6207 634 6222 668
rect 6278 634 6308 656
rect 6422 634 6452 656
rect 6508 634 6523 668
rect 6601 634 6631 661
rect 6679 695 6709 728
rect 6794 716 6824 738
rect 6679 634 6709 661
rect 6787 634 6802 668
rect 6858 634 6888 656
rect 128 620 158 634
rect 392 620 422 634
rect 708 620 738 634
rect 972 620 1002 634
rect 1288 620 1318 634
rect 1552 620 1582 634
rect 1868 620 1898 634
rect 2132 620 2162 634
rect 2448 620 2478 634
rect 2712 620 2742 634
rect 3028 620 3058 634
rect 3292 620 3322 634
rect 3608 620 3638 634
rect 3872 620 3902 634
rect 4188 620 4218 634
rect 4452 620 4482 634
rect 4768 620 4798 634
rect 5032 620 5062 634
rect 5348 620 5378 634
rect 5612 620 5642 634
rect 5928 620 5958 634
rect 6192 620 6222 634
rect 6508 620 6538 634
rect 6772 620 6802 634
rect 42 570 72 592
rect 128 570 158 592
rect 221 570 251 592
rect 299 570 329 592
rect 392 570 422 592
rect 478 570 508 592
rect 622 570 652 592
rect 708 570 738 592
rect 801 570 831 592
rect 879 570 909 592
rect 972 570 1002 592
rect 1058 570 1088 592
rect 1202 570 1232 592
rect 1288 570 1318 592
rect 1381 570 1411 592
rect 1459 570 1489 592
rect 1552 570 1582 592
rect 1638 570 1668 592
rect 1782 570 1812 592
rect 1868 570 1898 592
rect 1961 570 1991 592
rect 2039 570 2069 592
rect 2132 570 2162 592
rect 2218 570 2248 592
rect 2362 570 2392 592
rect 2448 570 2478 592
rect 2541 570 2571 592
rect 2619 570 2649 592
rect 2712 570 2742 592
rect 2798 570 2828 592
rect 2942 570 2972 592
rect 3028 570 3058 592
rect 3121 570 3151 592
rect 3199 570 3229 592
rect 3292 570 3322 592
rect 3378 570 3408 592
rect 3522 570 3552 592
rect 3608 570 3638 592
rect 3701 570 3731 592
rect 3779 570 3809 592
rect 3872 570 3902 592
rect 3958 570 3988 592
rect 4102 570 4132 592
rect 4188 570 4218 592
rect 4281 570 4311 592
rect 4359 570 4389 592
rect 4452 570 4482 592
rect 4538 570 4568 592
rect 4682 570 4712 592
rect 4768 570 4798 592
rect 4861 570 4891 592
rect 4939 570 4969 592
rect 5032 570 5062 592
rect 5118 570 5148 592
rect 5262 570 5292 592
rect 5348 570 5378 592
rect 5441 570 5471 592
rect 5519 570 5549 592
rect 5612 570 5642 592
rect 5698 570 5728 592
rect 5842 570 5872 592
rect 5928 570 5958 592
rect 6021 570 6051 592
rect 6099 570 6129 592
rect 6192 570 6222 592
rect 6278 570 6308 592
rect 6422 570 6452 592
rect 6508 570 6538 592
rect 6601 570 6631 592
rect 6679 570 6709 592
rect 6772 570 6802 592
rect 6858 570 6888 592
rect -1 524 6931 554
rect 106 496 136 524
rect 221 486 251 508
rect 299 486 329 508
rect 414 496 444 524
rect 106 446 136 468
rect 686 496 716 524
rect 801 486 831 508
rect 879 486 909 508
rect 994 496 1024 524
rect 221 425 251 458
rect 42 364 72 386
rect 128 364 143 398
rect 221 364 251 391
rect 299 425 329 458
rect 414 446 444 468
rect 686 446 716 468
rect 1266 496 1296 524
rect 1381 486 1411 508
rect 1459 486 1489 508
rect 1574 496 1604 524
rect 801 425 831 458
rect 299 364 329 391
rect 407 364 422 398
rect 478 364 508 386
rect 622 364 652 386
rect 708 364 723 398
rect 801 364 831 391
rect 879 425 909 458
rect 994 446 1024 468
rect 1266 446 1296 468
rect 1846 496 1876 524
rect 1961 486 1991 508
rect 2039 486 2069 508
rect 2154 496 2184 524
rect 1381 425 1411 458
rect 879 364 909 391
rect 987 364 1002 398
rect 1058 364 1088 386
rect 1202 364 1232 386
rect 1288 364 1303 398
rect 1381 364 1411 391
rect 1459 425 1489 458
rect 1574 446 1604 468
rect 1846 446 1876 468
rect 2426 496 2456 524
rect 2541 486 2571 508
rect 2619 486 2649 508
rect 2734 496 2764 524
rect 1961 425 1991 458
rect 1459 364 1489 391
rect 1567 364 1582 398
rect 1638 364 1668 386
rect 1782 364 1812 386
rect 1868 364 1883 398
rect 1961 364 1991 391
rect 2039 425 2069 458
rect 2154 446 2184 468
rect 2426 446 2456 468
rect 3006 496 3036 524
rect 3121 486 3151 508
rect 3199 486 3229 508
rect 3314 496 3344 524
rect 2541 425 2571 458
rect 2039 364 2069 391
rect 2147 364 2162 398
rect 2218 364 2248 386
rect 2362 364 2392 386
rect 2448 364 2463 398
rect 2541 364 2571 391
rect 2619 425 2649 458
rect 2734 446 2764 468
rect 3006 446 3036 468
rect 3586 496 3616 524
rect 3701 486 3731 508
rect 3779 486 3809 508
rect 3894 496 3924 524
rect 3121 425 3151 458
rect 2619 364 2649 391
rect 2727 364 2742 398
rect 2798 364 2828 386
rect 2942 364 2972 386
rect 3028 364 3043 398
rect 3121 364 3151 391
rect 3199 425 3229 458
rect 3314 446 3344 468
rect 3586 446 3616 468
rect 4166 496 4196 524
rect 4281 486 4311 508
rect 4359 486 4389 508
rect 4474 496 4504 524
rect 3701 425 3731 458
rect 3199 364 3229 391
rect 3307 364 3322 398
rect 3378 364 3408 386
rect 3522 364 3552 386
rect 3608 364 3623 398
rect 3701 364 3731 391
rect 3779 425 3809 458
rect 3894 446 3924 468
rect 4166 446 4196 468
rect 4746 496 4776 524
rect 4861 486 4891 508
rect 4939 486 4969 508
rect 5054 496 5084 524
rect 4281 425 4311 458
rect 3779 364 3809 391
rect 3887 364 3902 398
rect 3958 364 3988 386
rect 4102 364 4132 386
rect 4188 364 4203 398
rect 4281 364 4311 391
rect 4359 425 4389 458
rect 4474 446 4504 468
rect 4746 446 4776 468
rect 5326 496 5356 524
rect 5441 486 5471 508
rect 5519 486 5549 508
rect 5634 496 5664 524
rect 4861 425 4891 458
rect 4359 364 4389 391
rect 4467 364 4482 398
rect 4538 364 4568 386
rect 4682 364 4712 386
rect 4768 364 4783 398
rect 4861 364 4891 391
rect 4939 425 4969 458
rect 5054 446 5084 468
rect 5326 446 5356 468
rect 5906 496 5936 524
rect 6021 486 6051 508
rect 6099 486 6129 508
rect 6214 496 6244 524
rect 5441 425 5471 458
rect 4939 364 4969 391
rect 5047 364 5062 398
rect 5118 364 5148 386
rect 5262 364 5292 386
rect 5348 364 5363 398
rect 5441 364 5471 391
rect 5519 425 5549 458
rect 5634 446 5664 468
rect 5906 446 5936 468
rect 6486 496 6516 524
rect 6601 486 6631 508
rect 6679 486 6709 508
rect 6794 496 6824 524
rect 6021 425 6051 458
rect 5519 364 5549 391
rect 5627 364 5642 398
rect 5698 364 5728 386
rect 5842 364 5872 386
rect 5928 364 5943 398
rect 6021 364 6051 391
rect 6099 425 6129 458
rect 6214 446 6244 468
rect 6486 446 6516 468
rect 6601 425 6631 458
rect 6099 364 6129 391
rect 6207 364 6222 398
rect 6278 364 6308 386
rect 6422 364 6452 386
rect 6508 364 6523 398
rect 6601 364 6631 391
rect 6679 425 6709 458
rect 6794 446 6824 468
rect 6679 364 6709 391
rect 6787 364 6802 398
rect 6858 364 6888 386
rect 128 350 158 364
rect 392 350 422 364
rect 708 350 738 364
rect 972 350 1002 364
rect 1288 350 1318 364
rect 1552 350 1582 364
rect 1868 350 1898 364
rect 2132 350 2162 364
rect 2448 350 2478 364
rect 2712 350 2742 364
rect 3028 350 3058 364
rect 3292 350 3322 364
rect 3608 350 3638 364
rect 3872 350 3902 364
rect 4188 350 4218 364
rect 4452 350 4482 364
rect 4768 350 4798 364
rect 5032 350 5062 364
rect 5348 350 5378 364
rect 5612 350 5642 364
rect 5928 350 5958 364
rect 6192 350 6222 364
rect 6508 350 6538 364
rect 6772 350 6802 364
rect 42 300 72 322
rect 128 300 158 322
rect 221 300 251 322
rect 299 300 329 322
rect 392 300 422 322
rect 478 300 508 322
rect 622 300 652 322
rect 708 300 738 322
rect 801 300 831 322
rect 879 300 909 322
rect 972 300 1002 322
rect 1058 300 1088 322
rect 1202 300 1232 322
rect 1288 300 1318 322
rect 1381 300 1411 322
rect 1459 300 1489 322
rect 1552 300 1582 322
rect 1638 300 1668 322
rect 1782 300 1812 322
rect 1868 300 1898 322
rect 1961 300 1991 322
rect 2039 300 2069 322
rect 2132 300 2162 322
rect 2218 300 2248 322
rect 2362 300 2392 322
rect 2448 300 2478 322
rect 2541 300 2571 322
rect 2619 300 2649 322
rect 2712 300 2742 322
rect 2798 300 2828 322
rect 2942 300 2972 322
rect 3028 300 3058 322
rect 3121 300 3151 322
rect 3199 300 3229 322
rect 3292 300 3322 322
rect 3378 300 3408 322
rect 3522 300 3552 322
rect 3608 300 3638 322
rect 3701 300 3731 322
rect 3779 300 3809 322
rect 3872 300 3902 322
rect 3958 300 3988 322
rect 4102 300 4132 322
rect 4188 300 4218 322
rect 4281 300 4311 322
rect 4359 300 4389 322
rect 4452 300 4482 322
rect 4538 300 4568 322
rect 4682 300 4712 322
rect 4768 300 4798 322
rect 4861 300 4891 322
rect 4939 300 4969 322
rect 5032 300 5062 322
rect 5118 300 5148 322
rect 5262 300 5292 322
rect 5348 300 5378 322
rect 5441 300 5471 322
rect 5519 300 5549 322
rect 5612 300 5642 322
rect 5698 300 5728 322
rect 5842 300 5872 322
rect 5928 300 5958 322
rect 6021 300 6051 322
rect 6099 300 6129 322
rect 6192 300 6222 322
rect 6278 300 6308 322
rect 6422 300 6452 322
rect 6508 300 6538 322
rect 6601 300 6631 322
rect 6679 300 6709 322
rect 6772 300 6802 322
rect 6858 300 6888 322
rect -1 254 6931 284
rect 106 226 136 254
rect 221 216 251 238
rect 299 216 329 238
rect 414 226 444 254
rect 106 176 136 198
rect 686 226 716 254
rect 801 216 831 238
rect 879 216 909 238
rect 994 226 1024 254
rect 221 155 251 188
rect 42 94 72 116
rect 128 94 143 128
rect 221 94 251 121
rect 299 155 329 188
rect 414 176 444 198
rect 686 176 716 198
rect 1266 226 1296 254
rect 1381 216 1411 238
rect 1459 216 1489 238
rect 1574 226 1604 254
rect 801 155 831 188
rect 299 94 329 121
rect 407 94 422 128
rect 478 94 508 116
rect 622 94 652 116
rect 708 94 723 128
rect 801 94 831 121
rect 879 155 909 188
rect 994 176 1024 198
rect 1266 176 1296 198
rect 1846 226 1876 254
rect 1961 216 1991 238
rect 2039 216 2069 238
rect 2154 226 2184 254
rect 1381 155 1411 188
rect 879 94 909 121
rect 987 94 1002 128
rect 1058 94 1088 116
rect 1202 94 1232 116
rect 1288 94 1303 128
rect 1381 94 1411 121
rect 1459 155 1489 188
rect 1574 176 1604 198
rect 1846 176 1876 198
rect 2426 226 2456 254
rect 2541 216 2571 238
rect 2619 216 2649 238
rect 2734 226 2764 254
rect 1961 155 1991 188
rect 1459 94 1489 121
rect 1567 94 1582 128
rect 1638 94 1668 116
rect 1782 94 1812 116
rect 1868 94 1883 128
rect 1961 94 1991 121
rect 2039 155 2069 188
rect 2154 176 2184 198
rect 2426 176 2456 198
rect 3006 226 3036 254
rect 3121 216 3151 238
rect 3199 216 3229 238
rect 3314 226 3344 254
rect 2541 155 2571 188
rect 2039 94 2069 121
rect 2147 94 2162 128
rect 2218 94 2248 116
rect 2362 94 2392 116
rect 2448 94 2463 128
rect 2541 94 2571 121
rect 2619 155 2649 188
rect 2734 176 2764 198
rect 3006 176 3036 198
rect 3586 226 3616 254
rect 3701 216 3731 238
rect 3779 216 3809 238
rect 3894 226 3924 254
rect 3121 155 3151 188
rect 2619 94 2649 121
rect 2727 94 2742 128
rect 2798 94 2828 116
rect 2942 94 2972 116
rect 3028 94 3043 128
rect 3121 94 3151 121
rect 3199 155 3229 188
rect 3314 176 3344 198
rect 3586 176 3616 198
rect 4166 226 4196 254
rect 4281 216 4311 238
rect 4359 216 4389 238
rect 4474 226 4504 254
rect 3701 155 3731 188
rect 3199 94 3229 121
rect 3307 94 3322 128
rect 3378 94 3408 116
rect 3522 94 3552 116
rect 3608 94 3623 128
rect 3701 94 3731 121
rect 3779 155 3809 188
rect 3894 176 3924 198
rect 4166 176 4196 198
rect 4746 226 4776 254
rect 4861 216 4891 238
rect 4939 216 4969 238
rect 5054 226 5084 254
rect 4281 155 4311 188
rect 3779 94 3809 121
rect 3887 94 3902 128
rect 3958 94 3988 116
rect 4102 94 4132 116
rect 4188 94 4203 128
rect 4281 94 4311 121
rect 4359 155 4389 188
rect 4474 176 4504 198
rect 4746 176 4776 198
rect 5326 226 5356 254
rect 5441 216 5471 238
rect 5519 216 5549 238
rect 5634 226 5664 254
rect 4861 155 4891 188
rect 4359 94 4389 121
rect 4467 94 4482 128
rect 4538 94 4568 116
rect 4682 94 4712 116
rect 4768 94 4783 128
rect 4861 94 4891 121
rect 4939 155 4969 188
rect 5054 176 5084 198
rect 5326 176 5356 198
rect 5906 226 5936 254
rect 6021 216 6051 238
rect 6099 216 6129 238
rect 6214 226 6244 254
rect 5441 155 5471 188
rect 4939 94 4969 121
rect 5047 94 5062 128
rect 5118 94 5148 116
rect 5262 94 5292 116
rect 5348 94 5363 128
rect 5441 94 5471 121
rect 5519 155 5549 188
rect 5634 176 5664 198
rect 5906 176 5936 198
rect 6486 226 6516 254
rect 6601 216 6631 238
rect 6679 216 6709 238
rect 6794 226 6824 254
rect 6021 155 6051 188
rect 5519 94 5549 121
rect 5627 94 5642 128
rect 5698 94 5728 116
rect 5842 94 5872 116
rect 5928 94 5943 128
rect 6021 94 6051 121
rect 6099 155 6129 188
rect 6214 176 6244 198
rect 6486 176 6516 198
rect 6601 155 6631 188
rect 6099 94 6129 121
rect 6207 94 6222 128
rect 6278 94 6308 116
rect 6422 94 6452 116
rect 6508 94 6523 128
rect 6601 94 6631 121
rect 6679 155 6709 188
rect 6794 176 6824 198
rect 6679 94 6709 121
rect 6787 94 6802 128
rect 6858 94 6888 116
rect 128 80 158 94
rect 392 80 422 94
rect 708 80 738 94
rect 972 80 1002 94
rect 1288 80 1318 94
rect 1552 80 1582 94
rect 1868 80 1898 94
rect 2132 80 2162 94
rect 2448 80 2478 94
rect 2712 80 2742 94
rect 3028 80 3058 94
rect 3292 80 3322 94
rect 3608 80 3638 94
rect 3872 80 3902 94
rect 4188 80 4218 94
rect 4452 80 4482 94
rect 4768 80 4798 94
rect 5032 80 5062 94
rect 5348 80 5378 94
rect 5612 80 5642 94
rect 5928 80 5958 94
rect 6192 80 6222 94
rect 6508 80 6538 94
rect 6772 80 6802 94
rect 42 30 72 52
rect 128 30 158 52
rect 221 30 251 52
rect 299 30 329 52
rect 392 30 422 52
rect 478 30 508 52
rect 622 30 652 52
rect 708 30 738 52
rect 801 30 831 52
rect 879 30 909 52
rect 972 30 1002 52
rect 1058 30 1088 52
rect 1202 30 1232 52
rect 1288 30 1318 52
rect 1381 30 1411 52
rect 1459 30 1489 52
rect 1552 30 1582 52
rect 1638 30 1668 52
rect 1782 30 1812 52
rect 1868 30 1898 52
rect 1961 30 1991 52
rect 2039 30 2069 52
rect 2132 30 2162 52
rect 2218 30 2248 52
rect 2362 30 2392 52
rect 2448 30 2478 52
rect 2541 30 2571 52
rect 2619 30 2649 52
rect 2712 30 2742 52
rect 2798 30 2828 52
rect 2942 30 2972 52
rect 3028 30 3058 52
rect 3121 30 3151 52
rect 3199 30 3229 52
rect 3292 30 3322 52
rect 3378 30 3408 52
rect 3522 30 3552 52
rect 3608 30 3638 52
rect 3701 30 3731 52
rect 3779 30 3809 52
rect 3872 30 3902 52
rect 3958 30 3988 52
rect 4102 30 4132 52
rect 4188 30 4218 52
rect 4281 30 4311 52
rect 4359 30 4389 52
rect 4452 30 4482 52
rect 4538 30 4568 52
rect 4682 30 4712 52
rect 4768 30 4798 52
rect 4861 30 4891 52
rect 4939 30 4969 52
rect 5032 30 5062 52
rect 5118 30 5148 52
rect 5262 30 5292 52
rect 5348 30 5378 52
rect 5441 30 5471 52
rect 5519 30 5549 52
rect 5612 30 5642 52
rect 5698 30 5728 52
rect 5842 30 5872 52
rect 5928 30 5958 52
rect 6021 30 6051 52
rect 6099 30 6129 52
rect 6192 30 6222 52
rect 6278 30 6308 52
rect 6422 30 6452 52
rect 6508 30 6538 52
rect 6601 30 6631 52
rect 6679 30 6709 52
rect 6772 30 6802 52
rect 6858 30 6888 52
rect -1 -16 6931 14
rect 106 -44 136 -16
rect 221 -54 251 -32
rect 299 -54 329 -32
rect 414 -44 444 -16
rect 106 -94 136 -72
rect 686 -44 716 -16
rect 801 -54 831 -32
rect 879 -54 909 -32
rect 994 -44 1024 -16
rect 221 -115 251 -82
rect 42 -176 72 -154
rect 128 -176 143 -142
rect 221 -176 251 -149
rect 299 -115 329 -82
rect 414 -94 444 -72
rect 686 -94 716 -72
rect 1266 -44 1296 -16
rect 1381 -54 1411 -32
rect 1459 -54 1489 -32
rect 1574 -44 1604 -16
rect 801 -115 831 -82
rect 299 -176 329 -149
rect 407 -176 422 -142
rect 478 -176 508 -154
rect 622 -176 652 -154
rect 708 -176 723 -142
rect 801 -176 831 -149
rect 879 -115 909 -82
rect 994 -94 1024 -72
rect 1266 -94 1296 -72
rect 1846 -44 1876 -16
rect 1961 -54 1991 -32
rect 2039 -54 2069 -32
rect 2154 -44 2184 -16
rect 1381 -115 1411 -82
rect 879 -176 909 -149
rect 987 -176 1002 -142
rect 1058 -176 1088 -154
rect 1202 -176 1232 -154
rect 1288 -176 1303 -142
rect 1381 -176 1411 -149
rect 1459 -115 1489 -82
rect 1574 -94 1604 -72
rect 1846 -94 1876 -72
rect 2426 -44 2456 -16
rect 2541 -54 2571 -32
rect 2619 -54 2649 -32
rect 2734 -44 2764 -16
rect 1961 -115 1991 -82
rect 1459 -176 1489 -149
rect 1567 -176 1582 -142
rect 1638 -176 1668 -154
rect 1782 -176 1812 -154
rect 1868 -176 1883 -142
rect 1961 -176 1991 -149
rect 2039 -115 2069 -82
rect 2154 -94 2184 -72
rect 2426 -94 2456 -72
rect 3006 -44 3036 -16
rect 3121 -54 3151 -32
rect 3199 -54 3229 -32
rect 3314 -44 3344 -16
rect 2541 -115 2571 -82
rect 2039 -176 2069 -149
rect 2147 -176 2162 -142
rect 2218 -176 2248 -154
rect 2362 -176 2392 -154
rect 2448 -176 2463 -142
rect 2541 -176 2571 -149
rect 2619 -115 2649 -82
rect 2734 -94 2764 -72
rect 3006 -94 3036 -72
rect 3586 -44 3616 -16
rect 3701 -54 3731 -32
rect 3779 -54 3809 -32
rect 3894 -44 3924 -16
rect 3121 -115 3151 -82
rect 2619 -176 2649 -149
rect 2727 -176 2742 -142
rect 2798 -176 2828 -154
rect 2942 -176 2972 -154
rect 3028 -176 3043 -142
rect 3121 -176 3151 -149
rect 3199 -115 3229 -82
rect 3314 -94 3344 -72
rect 3586 -94 3616 -72
rect 4166 -44 4196 -16
rect 4281 -54 4311 -32
rect 4359 -54 4389 -32
rect 4474 -44 4504 -16
rect 3701 -115 3731 -82
rect 3199 -176 3229 -149
rect 3307 -176 3322 -142
rect 3378 -176 3408 -154
rect 3522 -176 3552 -154
rect 3608 -176 3623 -142
rect 3701 -176 3731 -149
rect 3779 -115 3809 -82
rect 3894 -94 3924 -72
rect 4166 -94 4196 -72
rect 4746 -44 4776 -16
rect 4861 -54 4891 -32
rect 4939 -54 4969 -32
rect 5054 -44 5084 -16
rect 4281 -115 4311 -82
rect 3779 -176 3809 -149
rect 3887 -176 3902 -142
rect 3958 -176 3988 -154
rect 4102 -176 4132 -154
rect 4188 -176 4203 -142
rect 4281 -176 4311 -149
rect 4359 -115 4389 -82
rect 4474 -94 4504 -72
rect 4746 -94 4776 -72
rect 5326 -44 5356 -16
rect 5441 -54 5471 -32
rect 5519 -54 5549 -32
rect 5634 -44 5664 -16
rect 4861 -115 4891 -82
rect 4359 -176 4389 -149
rect 4467 -176 4482 -142
rect 4538 -176 4568 -154
rect 4682 -176 4712 -154
rect 4768 -176 4783 -142
rect 4861 -176 4891 -149
rect 4939 -115 4969 -82
rect 5054 -94 5084 -72
rect 5326 -94 5356 -72
rect 5906 -44 5936 -16
rect 6021 -54 6051 -32
rect 6099 -54 6129 -32
rect 6214 -44 6244 -16
rect 5441 -115 5471 -82
rect 4939 -176 4969 -149
rect 5047 -176 5062 -142
rect 5118 -176 5148 -154
rect 5262 -176 5292 -154
rect 5348 -176 5363 -142
rect 5441 -176 5471 -149
rect 5519 -115 5549 -82
rect 5634 -94 5664 -72
rect 5906 -94 5936 -72
rect 6486 -44 6516 -16
rect 6601 -54 6631 -32
rect 6679 -54 6709 -32
rect 6794 -44 6824 -16
rect 6021 -115 6051 -82
rect 5519 -176 5549 -149
rect 5627 -176 5642 -142
rect 5698 -176 5728 -154
rect 5842 -176 5872 -154
rect 5928 -176 5943 -142
rect 6021 -176 6051 -149
rect 6099 -115 6129 -82
rect 6214 -94 6244 -72
rect 6486 -94 6516 -72
rect 6601 -115 6631 -82
rect 6099 -176 6129 -149
rect 6207 -176 6222 -142
rect 6278 -176 6308 -154
rect 6422 -176 6452 -154
rect 6508 -176 6523 -142
rect 6601 -176 6631 -149
rect 6679 -115 6709 -82
rect 6794 -94 6824 -72
rect 6679 -176 6709 -149
rect 6787 -176 6802 -142
rect 6858 -176 6888 -154
rect 128 -190 158 -176
rect 392 -190 422 -176
rect 708 -190 738 -176
rect 972 -190 1002 -176
rect 1288 -190 1318 -176
rect 1552 -190 1582 -176
rect 1868 -190 1898 -176
rect 2132 -190 2162 -176
rect 2448 -190 2478 -176
rect 2712 -190 2742 -176
rect 3028 -190 3058 -176
rect 3292 -190 3322 -176
rect 3608 -190 3638 -176
rect 3872 -190 3902 -176
rect 4188 -190 4218 -176
rect 4452 -190 4482 -176
rect 4768 -190 4798 -176
rect 5032 -190 5062 -176
rect 5348 -190 5378 -176
rect 5612 -190 5642 -176
rect 5928 -190 5958 -176
rect 6192 -190 6222 -176
rect 6508 -190 6538 -176
rect 6772 -190 6802 -176
rect 42 -240 72 -218
rect 128 -240 158 -218
rect 221 -240 251 -218
rect 299 -240 329 -218
rect 392 -240 422 -218
rect 478 -240 508 -218
rect 622 -240 652 -218
rect 708 -240 738 -218
rect 801 -240 831 -218
rect 879 -240 909 -218
rect 972 -240 1002 -218
rect 1058 -240 1088 -218
rect 1202 -240 1232 -218
rect 1288 -240 1318 -218
rect 1381 -240 1411 -218
rect 1459 -240 1489 -218
rect 1552 -240 1582 -218
rect 1638 -240 1668 -218
rect 1782 -240 1812 -218
rect 1868 -240 1898 -218
rect 1961 -240 1991 -218
rect 2039 -240 2069 -218
rect 2132 -240 2162 -218
rect 2218 -240 2248 -218
rect 2362 -240 2392 -218
rect 2448 -240 2478 -218
rect 2541 -240 2571 -218
rect 2619 -240 2649 -218
rect 2712 -240 2742 -218
rect 2798 -240 2828 -218
rect 2942 -240 2972 -218
rect 3028 -240 3058 -218
rect 3121 -240 3151 -218
rect 3199 -240 3229 -218
rect 3292 -240 3322 -218
rect 3378 -240 3408 -218
rect 3522 -240 3552 -218
rect 3608 -240 3638 -218
rect 3701 -240 3731 -218
rect 3779 -240 3809 -218
rect 3872 -240 3902 -218
rect 3958 -240 3988 -218
rect 4102 -240 4132 -218
rect 4188 -240 4218 -218
rect 4281 -240 4311 -218
rect 4359 -240 4389 -218
rect 4452 -240 4482 -218
rect 4538 -240 4568 -218
rect 4682 -240 4712 -218
rect 4768 -240 4798 -218
rect 4861 -240 4891 -218
rect 4939 -240 4969 -218
rect 5032 -240 5062 -218
rect 5118 -240 5148 -218
rect 5262 -240 5292 -218
rect 5348 -240 5378 -218
rect 5441 -240 5471 -218
rect 5519 -240 5549 -218
rect 5612 -240 5642 -218
rect 5698 -240 5728 -218
rect 5842 -240 5872 -218
rect 5928 -240 5958 -218
rect 6021 -240 6051 -218
rect 6099 -240 6129 -218
rect 6192 -240 6222 -218
rect 6278 -240 6308 -218
rect 6422 -240 6452 -218
rect 6508 -240 6538 -218
rect 6601 -240 6631 -218
rect 6679 -240 6709 -218
rect 6772 -240 6802 -218
rect 6858 -240 6888 -218
rect -1 -286 6931 -256
rect 106 -314 136 -286
rect 221 -324 251 -302
rect 299 -324 329 -302
rect 414 -314 444 -286
rect 106 -364 136 -342
rect 686 -314 716 -286
rect 801 -324 831 -302
rect 879 -324 909 -302
rect 994 -314 1024 -286
rect 221 -385 251 -352
rect 42 -446 72 -424
rect 128 -446 143 -412
rect 221 -446 251 -419
rect 299 -385 329 -352
rect 414 -364 444 -342
rect 686 -364 716 -342
rect 1266 -314 1296 -286
rect 1381 -324 1411 -302
rect 1459 -324 1489 -302
rect 1574 -314 1604 -286
rect 801 -385 831 -352
rect 299 -446 329 -419
rect 407 -446 422 -412
rect 478 -446 508 -424
rect 622 -446 652 -424
rect 708 -446 723 -412
rect 801 -446 831 -419
rect 879 -385 909 -352
rect 994 -364 1024 -342
rect 1266 -364 1296 -342
rect 1846 -314 1876 -286
rect 1961 -324 1991 -302
rect 2039 -324 2069 -302
rect 2154 -314 2184 -286
rect 1381 -385 1411 -352
rect 879 -446 909 -419
rect 987 -446 1002 -412
rect 1058 -446 1088 -424
rect 1202 -446 1232 -424
rect 1288 -446 1303 -412
rect 1381 -446 1411 -419
rect 1459 -385 1489 -352
rect 1574 -364 1604 -342
rect 1846 -364 1876 -342
rect 2426 -314 2456 -286
rect 2541 -324 2571 -302
rect 2619 -324 2649 -302
rect 2734 -314 2764 -286
rect 1961 -385 1991 -352
rect 1459 -446 1489 -419
rect 1567 -446 1582 -412
rect 1638 -446 1668 -424
rect 1782 -446 1812 -424
rect 1868 -446 1883 -412
rect 1961 -446 1991 -419
rect 2039 -385 2069 -352
rect 2154 -364 2184 -342
rect 2426 -364 2456 -342
rect 3006 -314 3036 -286
rect 3121 -324 3151 -302
rect 3199 -324 3229 -302
rect 3314 -314 3344 -286
rect 2541 -385 2571 -352
rect 2039 -446 2069 -419
rect 2147 -446 2162 -412
rect 2218 -446 2248 -424
rect 2362 -446 2392 -424
rect 2448 -446 2463 -412
rect 2541 -446 2571 -419
rect 2619 -385 2649 -352
rect 2734 -364 2764 -342
rect 3006 -364 3036 -342
rect 3586 -314 3616 -286
rect 3701 -324 3731 -302
rect 3779 -324 3809 -302
rect 3894 -314 3924 -286
rect 3121 -385 3151 -352
rect 2619 -446 2649 -419
rect 2727 -446 2742 -412
rect 2798 -446 2828 -424
rect 2942 -446 2972 -424
rect 3028 -446 3043 -412
rect 3121 -446 3151 -419
rect 3199 -385 3229 -352
rect 3314 -364 3344 -342
rect 3586 -364 3616 -342
rect 4166 -314 4196 -286
rect 4281 -324 4311 -302
rect 4359 -324 4389 -302
rect 4474 -314 4504 -286
rect 3701 -385 3731 -352
rect 3199 -446 3229 -419
rect 3307 -446 3322 -412
rect 3378 -446 3408 -424
rect 3522 -446 3552 -424
rect 3608 -446 3623 -412
rect 3701 -446 3731 -419
rect 3779 -385 3809 -352
rect 3894 -364 3924 -342
rect 4166 -364 4196 -342
rect 4746 -314 4776 -286
rect 4861 -324 4891 -302
rect 4939 -324 4969 -302
rect 5054 -314 5084 -286
rect 4281 -385 4311 -352
rect 3779 -446 3809 -419
rect 3887 -446 3902 -412
rect 3958 -446 3988 -424
rect 4102 -446 4132 -424
rect 4188 -446 4203 -412
rect 4281 -446 4311 -419
rect 4359 -385 4389 -352
rect 4474 -364 4504 -342
rect 4746 -364 4776 -342
rect 5326 -314 5356 -286
rect 5441 -324 5471 -302
rect 5519 -324 5549 -302
rect 5634 -314 5664 -286
rect 4861 -385 4891 -352
rect 4359 -446 4389 -419
rect 4467 -446 4482 -412
rect 4538 -446 4568 -424
rect 4682 -446 4712 -424
rect 4768 -446 4783 -412
rect 4861 -446 4891 -419
rect 4939 -385 4969 -352
rect 5054 -364 5084 -342
rect 5326 -364 5356 -342
rect 5906 -314 5936 -286
rect 6021 -324 6051 -302
rect 6099 -324 6129 -302
rect 6214 -314 6244 -286
rect 5441 -385 5471 -352
rect 4939 -446 4969 -419
rect 5047 -446 5062 -412
rect 5118 -446 5148 -424
rect 5262 -446 5292 -424
rect 5348 -446 5363 -412
rect 5441 -446 5471 -419
rect 5519 -385 5549 -352
rect 5634 -364 5664 -342
rect 5906 -364 5936 -342
rect 6486 -314 6516 -286
rect 6601 -324 6631 -302
rect 6679 -324 6709 -302
rect 6794 -314 6824 -286
rect 6021 -385 6051 -352
rect 5519 -446 5549 -419
rect 5627 -446 5642 -412
rect 5698 -446 5728 -424
rect 5842 -446 5872 -424
rect 5928 -446 5943 -412
rect 6021 -446 6051 -419
rect 6099 -385 6129 -352
rect 6214 -364 6244 -342
rect 6486 -364 6516 -342
rect 6601 -385 6631 -352
rect 6099 -446 6129 -419
rect 6207 -446 6222 -412
rect 6278 -446 6308 -424
rect 6422 -446 6452 -424
rect 6508 -446 6523 -412
rect 6601 -446 6631 -419
rect 6679 -385 6709 -352
rect 6794 -364 6824 -342
rect 6679 -446 6709 -419
rect 6787 -446 6802 -412
rect 6858 -446 6888 -424
rect 128 -460 158 -446
rect 392 -460 422 -446
rect 708 -460 738 -446
rect 972 -460 1002 -446
rect 1288 -460 1318 -446
rect 1552 -460 1582 -446
rect 1868 -460 1898 -446
rect 2132 -460 2162 -446
rect 2448 -460 2478 -446
rect 2712 -460 2742 -446
rect 3028 -460 3058 -446
rect 3292 -460 3322 -446
rect 3608 -460 3638 -446
rect 3872 -460 3902 -446
rect 4188 -460 4218 -446
rect 4452 -460 4482 -446
rect 4768 -460 4798 -446
rect 5032 -460 5062 -446
rect 5348 -460 5378 -446
rect 5612 -460 5642 -446
rect 5928 -460 5958 -446
rect 6192 -460 6222 -446
rect 6508 -460 6538 -446
rect 6772 -460 6802 -446
rect 42 -510 72 -488
rect 128 -510 158 -488
rect 221 -510 251 -488
rect 299 -510 329 -488
rect 392 -510 422 -488
rect 478 -510 508 -488
rect 622 -510 652 -488
rect 708 -510 738 -488
rect 801 -510 831 -488
rect 879 -510 909 -488
rect 972 -510 1002 -488
rect 1058 -510 1088 -488
rect 1202 -510 1232 -488
rect 1288 -510 1318 -488
rect 1381 -510 1411 -488
rect 1459 -510 1489 -488
rect 1552 -510 1582 -488
rect 1638 -510 1668 -488
rect 1782 -510 1812 -488
rect 1868 -510 1898 -488
rect 1961 -510 1991 -488
rect 2039 -510 2069 -488
rect 2132 -510 2162 -488
rect 2218 -510 2248 -488
rect 2362 -510 2392 -488
rect 2448 -510 2478 -488
rect 2541 -510 2571 -488
rect 2619 -510 2649 -488
rect 2712 -510 2742 -488
rect 2798 -510 2828 -488
rect 2942 -510 2972 -488
rect 3028 -510 3058 -488
rect 3121 -510 3151 -488
rect 3199 -510 3229 -488
rect 3292 -510 3322 -488
rect 3378 -510 3408 -488
rect 3522 -510 3552 -488
rect 3608 -510 3638 -488
rect 3701 -510 3731 -488
rect 3779 -510 3809 -488
rect 3872 -510 3902 -488
rect 3958 -510 3988 -488
rect 4102 -510 4132 -488
rect 4188 -510 4218 -488
rect 4281 -510 4311 -488
rect 4359 -510 4389 -488
rect 4452 -510 4482 -488
rect 4538 -510 4568 -488
rect 4682 -510 4712 -488
rect 4768 -510 4798 -488
rect 4861 -510 4891 -488
rect 4939 -510 4969 -488
rect 5032 -510 5062 -488
rect 5118 -510 5148 -488
rect 5262 -510 5292 -488
rect 5348 -510 5378 -488
rect 5441 -510 5471 -488
rect 5519 -510 5549 -488
rect 5612 -510 5642 -488
rect 5698 -510 5728 -488
rect 5842 -510 5872 -488
rect 5928 -510 5958 -488
rect 6021 -510 6051 -488
rect 6099 -510 6129 -488
rect 6192 -510 6222 -488
rect 6278 -510 6308 -488
rect 6422 -510 6452 -488
rect 6508 -510 6538 -488
rect 6601 -510 6631 -488
rect 6679 -510 6709 -488
rect 6772 -510 6802 -488
rect 6858 -510 6888 -488
rect -1 -556 6931 -526
rect 106 -584 136 -556
rect 221 -594 251 -572
rect 299 -594 329 -572
rect 414 -584 444 -556
rect 106 -634 136 -612
rect 686 -584 716 -556
rect 801 -594 831 -572
rect 879 -594 909 -572
rect 994 -584 1024 -556
rect 221 -655 251 -622
rect 42 -716 72 -694
rect 128 -716 143 -682
rect 221 -716 251 -689
rect 299 -655 329 -622
rect 414 -634 444 -612
rect 686 -634 716 -612
rect 1266 -584 1296 -556
rect 1381 -594 1411 -572
rect 1459 -594 1489 -572
rect 1574 -584 1604 -556
rect 801 -655 831 -622
rect 299 -716 329 -689
rect 407 -716 422 -682
rect 478 -716 508 -694
rect 622 -716 652 -694
rect 708 -716 723 -682
rect 801 -716 831 -689
rect 879 -655 909 -622
rect 994 -634 1024 -612
rect 1266 -634 1296 -612
rect 1846 -584 1876 -556
rect 1961 -594 1991 -572
rect 2039 -594 2069 -572
rect 2154 -584 2184 -556
rect 1381 -655 1411 -622
rect 879 -716 909 -689
rect 987 -716 1002 -682
rect 1058 -716 1088 -694
rect 1202 -716 1232 -694
rect 1288 -716 1303 -682
rect 1381 -716 1411 -689
rect 1459 -655 1489 -622
rect 1574 -634 1604 -612
rect 1846 -634 1876 -612
rect 2426 -584 2456 -556
rect 2541 -594 2571 -572
rect 2619 -594 2649 -572
rect 2734 -584 2764 -556
rect 1961 -655 1991 -622
rect 1459 -716 1489 -689
rect 1567 -716 1582 -682
rect 1638 -716 1668 -694
rect 1782 -716 1812 -694
rect 1868 -716 1883 -682
rect 1961 -716 1991 -689
rect 2039 -655 2069 -622
rect 2154 -634 2184 -612
rect 2426 -634 2456 -612
rect 3006 -584 3036 -556
rect 3121 -594 3151 -572
rect 3199 -594 3229 -572
rect 3314 -584 3344 -556
rect 2541 -655 2571 -622
rect 2039 -716 2069 -689
rect 2147 -716 2162 -682
rect 2218 -716 2248 -694
rect 2362 -716 2392 -694
rect 2448 -716 2463 -682
rect 2541 -716 2571 -689
rect 2619 -655 2649 -622
rect 2734 -634 2764 -612
rect 3006 -634 3036 -612
rect 3586 -584 3616 -556
rect 3701 -594 3731 -572
rect 3779 -594 3809 -572
rect 3894 -584 3924 -556
rect 3121 -655 3151 -622
rect 2619 -716 2649 -689
rect 2727 -716 2742 -682
rect 2798 -716 2828 -694
rect 2942 -716 2972 -694
rect 3028 -716 3043 -682
rect 3121 -716 3151 -689
rect 3199 -655 3229 -622
rect 3314 -634 3344 -612
rect 3586 -634 3616 -612
rect 4166 -584 4196 -556
rect 4281 -594 4311 -572
rect 4359 -594 4389 -572
rect 4474 -584 4504 -556
rect 3701 -655 3731 -622
rect 3199 -716 3229 -689
rect 3307 -716 3322 -682
rect 3378 -716 3408 -694
rect 3522 -716 3552 -694
rect 3608 -716 3623 -682
rect 3701 -716 3731 -689
rect 3779 -655 3809 -622
rect 3894 -634 3924 -612
rect 4166 -634 4196 -612
rect 4746 -584 4776 -556
rect 4861 -594 4891 -572
rect 4939 -594 4969 -572
rect 5054 -584 5084 -556
rect 4281 -655 4311 -622
rect 3779 -716 3809 -689
rect 3887 -716 3902 -682
rect 3958 -716 3988 -694
rect 4102 -716 4132 -694
rect 4188 -716 4203 -682
rect 4281 -716 4311 -689
rect 4359 -655 4389 -622
rect 4474 -634 4504 -612
rect 4746 -634 4776 -612
rect 5326 -584 5356 -556
rect 5441 -594 5471 -572
rect 5519 -594 5549 -572
rect 5634 -584 5664 -556
rect 4861 -655 4891 -622
rect 4359 -716 4389 -689
rect 4467 -716 4482 -682
rect 4538 -716 4568 -694
rect 4682 -716 4712 -694
rect 4768 -716 4783 -682
rect 4861 -716 4891 -689
rect 4939 -655 4969 -622
rect 5054 -634 5084 -612
rect 5326 -634 5356 -612
rect 5906 -584 5936 -556
rect 6021 -594 6051 -572
rect 6099 -594 6129 -572
rect 6214 -584 6244 -556
rect 5441 -655 5471 -622
rect 4939 -716 4969 -689
rect 5047 -716 5062 -682
rect 5118 -716 5148 -694
rect 5262 -716 5292 -694
rect 5348 -716 5363 -682
rect 5441 -716 5471 -689
rect 5519 -655 5549 -622
rect 5634 -634 5664 -612
rect 5906 -634 5936 -612
rect 6486 -584 6516 -556
rect 6601 -594 6631 -572
rect 6679 -594 6709 -572
rect 6794 -584 6824 -556
rect 6021 -655 6051 -622
rect 5519 -716 5549 -689
rect 5627 -716 5642 -682
rect 5698 -716 5728 -694
rect 5842 -716 5872 -694
rect 5928 -716 5943 -682
rect 6021 -716 6051 -689
rect 6099 -655 6129 -622
rect 6214 -634 6244 -612
rect 6486 -634 6516 -612
rect 6601 -655 6631 -622
rect 6099 -716 6129 -689
rect 6207 -716 6222 -682
rect 6278 -716 6308 -694
rect 6422 -716 6452 -694
rect 6508 -716 6523 -682
rect 6601 -716 6631 -689
rect 6679 -655 6709 -622
rect 6794 -634 6824 -612
rect 6679 -716 6709 -689
rect 6787 -716 6802 -682
rect 6858 -716 6888 -694
rect 128 -730 158 -716
rect 392 -730 422 -716
rect 708 -730 738 -716
rect 972 -730 1002 -716
rect 1288 -730 1318 -716
rect 1552 -730 1582 -716
rect 1868 -730 1898 -716
rect 2132 -730 2162 -716
rect 2448 -730 2478 -716
rect 2712 -730 2742 -716
rect 3028 -730 3058 -716
rect 3292 -730 3322 -716
rect 3608 -730 3638 -716
rect 3872 -730 3902 -716
rect 4188 -730 4218 -716
rect 4452 -730 4482 -716
rect 4768 -730 4798 -716
rect 5032 -730 5062 -716
rect 5348 -730 5378 -716
rect 5612 -730 5642 -716
rect 5928 -730 5958 -716
rect 6192 -730 6222 -716
rect 6508 -730 6538 -716
rect 6772 -730 6802 -716
rect 42 -780 72 -758
rect 128 -780 158 -758
rect 221 -780 251 -758
rect 299 -780 329 -758
rect 392 -780 422 -758
rect 478 -780 508 -758
rect 622 -780 652 -758
rect 708 -780 738 -758
rect 801 -780 831 -758
rect 879 -780 909 -758
rect 972 -780 1002 -758
rect 1058 -780 1088 -758
rect 1202 -780 1232 -758
rect 1288 -780 1318 -758
rect 1381 -780 1411 -758
rect 1459 -780 1489 -758
rect 1552 -780 1582 -758
rect 1638 -780 1668 -758
rect 1782 -780 1812 -758
rect 1868 -780 1898 -758
rect 1961 -780 1991 -758
rect 2039 -780 2069 -758
rect 2132 -780 2162 -758
rect 2218 -780 2248 -758
rect 2362 -780 2392 -758
rect 2448 -780 2478 -758
rect 2541 -780 2571 -758
rect 2619 -780 2649 -758
rect 2712 -780 2742 -758
rect 2798 -780 2828 -758
rect 2942 -780 2972 -758
rect 3028 -780 3058 -758
rect 3121 -780 3151 -758
rect 3199 -780 3229 -758
rect 3292 -780 3322 -758
rect 3378 -780 3408 -758
rect 3522 -780 3552 -758
rect 3608 -780 3638 -758
rect 3701 -780 3731 -758
rect 3779 -780 3809 -758
rect 3872 -780 3902 -758
rect 3958 -780 3988 -758
rect 4102 -780 4132 -758
rect 4188 -780 4218 -758
rect 4281 -780 4311 -758
rect 4359 -780 4389 -758
rect 4452 -780 4482 -758
rect 4538 -780 4568 -758
rect 4682 -780 4712 -758
rect 4768 -780 4798 -758
rect 4861 -780 4891 -758
rect 4939 -780 4969 -758
rect 5032 -780 5062 -758
rect 5118 -780 5148 -758
rect 5262 -780 5292 -758
rect 5348 -780 5378 -758
rect 5441 -780 5471 -758
rect 5519 -780 5549 -758
rect 5612 -780 5642 -758
rect 5698 -780 5728 -758
rect 5842 -780 5872 -758
rect 5928 -780 5958 -758
rect 6021 -780 6051 -758
rect 6099 -780 6129 -758
rect 6192 -780 6222 -758
rect 6278 -780 6308 -758
rect 6422 -780 6452 -758
rect 6508 -780 6538 -758
rect 6601 -780 6631 -758
rect 6679 -780 6709 -758
rect 6772 -780 6802 -758
rect 6858 -780 6888 -758
rect -1 -826 6931 -796
rect 106 -854 136 -826
rect 221 -864 251 -842
rect 299 -864 329 -842
rect 414 -854 444 -826
rect 106 -904 136 -882
rect 686 -854 716 -826
rect 801 -864 831 -842
rect 879 -864 909 -842
rect 994 -854 1024 -826
rect 221 -925 251 -892
rect 42 -986 72 -964
rect 128 -986 143 -952
rect 221 -986 251 -959
rect 299 -925 329 -892
rect 414 -904 444 -882
rect 686 -904 716 -882
rect 1266 -854 1296 -826
rect 1381 -864 1411 -842
rect 1459 -864 1489 -842
rect 1574 -854 1604 -826
rect 801 -925 831 -892
rect 299 -986 329 -959
rect 407 -986 422 -952
rect 478 -986 508 -964
rect 622 -986 652 -964
rect 708 -986 723 -952
rect 801 -986 831 -959
rect 879 -925 909 -892
rect 994 -904 1024 -882
rect 1266 -904 1296 -882
rect 1846 -854 1876 -826
rect 1961 -864 1991 -842
rect 2039 -864 2069 -842
rect 2154 -854 2184 -826
rect 1381 -925 1411 -892
rect 879 -986 909 -959
rect 987 -986 1002 -952
rect 1058 -986 1088 -964
rect 1202 -986 1232 -964
rect 1288 -986 1303 -952
rect 1381 -986 1411 -959
rect 1459 -925 1489 -892
rect 1574 -904 1604 -882
rect 1846 -904 1876 -882
rect 2426 -854 2456 -826
rect 2541 -864 2571 -842
rect 2619 -864 2649 -842
rect 2734 -854 2764 -826
rect 1961 -925 1991 -892
rect 1459 -986 1489 -959
rect 1567 -986 1582 -952
rect 1638 -986 1668 -964
rect 1782 -986 1812 -964
rect 1868 -986 1883 -952
rect 1961 -986 1991 -959
rect 2039 -925 2069 -892
rect 2154 -904 2184 -882
rect 2426 -904 2456 -882
rect 3006 -854 3036 -826
rect 3121 -864 3151 -842
rect 3199 -864 3229 -842
rect 3314 -854 3344 -826
rect 2541 -925 2571 -892
rect 2039 -986 2069 -959
rect 2147 -986 2162 -952
rect 2218 -986 2248 -964
rect 2362 -986 2392 -964
rect 2448 -986 2463 -952
rect 2541 -986 2571 -959
rect 2619 -925 2649 -892
rect 2734 -904 2764 -882
rect 3006 -904 3036 -882
rect 3586 -854 3616 -826
rect 3701 -864 3731 -842
rect 3779 -864 3809 -842
rect 3894 -854 3924 -826
rect 3121 -925 3151 -892
rect 2619 -986 2649 -959
rect 2727 -986 2742 -952
rect 2798 -986 2828 -964
rect 2942 -986 2972 -964
rect 3028 -986 3043 -952
rect 3121 -986 3151 -959
rect 3199 -925 3229 -892
rect 3314 -904 3344 -882
rect 3586 -904 3616 -882
rect 4166 -854 4196 -826
rect 4281 -864 4311 -842
rect 4359 -864 4389 -842
rect 4474 -854 4504 -826
rect 3701 -925 3731 -892
rect 3199 -986 3229 -959
rect 3307 -986 3322 -952
rect 3378 -986 3408 -964
rect 3522 -986 3552 -964
rect 3608 -986 3623 -952
rect 3701 -986 3731 -959
rect 3779 -925 3809 -892
rect 3894 -904 3924 -882
rect 4166 -904 4196 -882
rect 4746 -854 4776 -826
rect 4861 -864 4891 -842
rect 4939 -864 4969 -842
rect 5054 -854 5084 -826
rect 4281 -925 4311 -892
rect 3779 -986 3809 -959
rect 3887 -986 3902 -952
rect 3958 -986 3988 -964
rect 4102 -986 4132 -964
rect 4188 -986 4203 -952
rect 4281 -986 4311 -959
rect 4359 -925 4389 -892
rect 4474 -904 4504 -882
rect 4746 -904 4776 -882
rect 5326 -854 5356 -826
rect 5441 -864 5471 -842
rect 5519 -864 5549 -842
rect 5634 -854 5664 -826
rect 4861 -925 4891 -892
rect 4359 -986 4389 -959
rect 4467 -986 4482 -952
rect 4538 -986 4568 -964
rect 4682 -986 4712 -964
rect 4768 -986 4783 -952
rect 4861 -986 4891 -959
rect 4939 -925 4969 -892
rect 5054 -904 5084 -882
rect 5326 -904 5356 -882
rect 5906 -854 5936 -826
rect 6021 -864 6051 -842
rect 6099 -864 6129 -842
rect 6214 -854 6244 -826
rect 5441 -925 5471 -892
rect 4939 -986 4969 -959
rect 5047 -986 5062 -952
rect 5118 -986 5148 -964
rect 5262 -986 5292 -964
rect 5348 -986 5363 -952
rect 5441 -986 5471 -959
rect 5519 -925 5549 -892
rect 5634 -904 5664 -882
rect 5906 -904 5936 -882
rect 6486 -854 6516 -826
rect 6601 -864 6631 -842
rect 6679 -864 6709 -842
rect 6794 -854 6824 -826
rect 6021 -925 6051 -892
rect 5519 -986 5549 -959
rect 5627 -986 5642 -952
rect 5698 -986 5728 -964
rect 5842 -986 5872 -964
rect 5928 -986 5943 -952
rect 6021 -986 6051 -959
rect 6099 -925 6129 -892
rect 6214 -904 6244 -882
rect 6486 -904 6516 -882
rect 6601 -925 6631 -892
rect 6099 -986 6129 -959
rect 6207 -986 6222 -952
rect 6278 -986 6308 -964
rect 6422 -986 6452 -964
rect 6508 -986 6523 -952
rect 6601 -986 6631 -959
rect 6679 -925 6709 -892
rect 6794 -904 6824 -882
rect 6679 -986 6709 -959
rect 6787 -986 6802 -952
rect 6858 -986 6888 -964
rect 128 -1000 158 -986
rect 392 -1000 422 -986
rect 708 -1000 738 -986
rect 972 -1000 1002 -986
rect 1288 -1000 1318 -986
rect 1552 -1000 1582 -986
rect 1868 -1000 1898 -986
rect 2132 -1000 2162 -986
rect 2448 -1000 2478 -986
rect 2712 -1000 2742 -986
rect 3028 -1000 3058 -986
rect 3292 -1000 3322 -986
rect 3608 -1000 3638 -986
rect 3872 -1000 3902 -986
rect 4188 -1000 4218 -986
rect 4452 -1000 4482 -986
rect 4768 -1000 4798 -986
rect 5032 -1000 5062 -986
rect 5348 -1000 5378 -986
rect 5612 -1000 5642 -986
rect 5928 -1000 5958 -986
rect 6192 -1000 6222 -986
rect 6508 -1000 6538 -986
rect 6772 -1000 6802 -986
rect 42 -1050 72 -1028
rect 128 -1050 158 -1028
rect 221 -1050 251 -1028
rect 299 -1050 329 -1028
rect 392 -1050 422 -1028
rect 478 -1050 508 -1028
rect 622 -1050 652 -1028
rect 708 -1050 738 -1028
rect 801 -1050 831 -1028
rect 879 -1050 909 -1028
rect 972 -1050 1002 -1028
rect 1058 -1050 1088 -1028
rect 1202 -1050 1232 -1028
rect 1288 -1050 1318 -1028
rect 1381 -1050 1411 -1028
rect 1459 -1050 1489 -1028
rect 1552 -1050 1582 -1028
rect 1638 -1050 1668 -1028
rect 1782 -1050 1812 -1028
rect 1868 -1050 1898 -1028
rect 1961 -1050 1991 -1028
rect 2039 -1050 2069 -1028
rect 2132 -1050 2162 -1028
rect 2218 -1050 2248 -1028
rect 2362 -1050 2392 -1028
rect 2448 -1050 2478 -1028
rect 2541 -1050 2571 -1028
rect 2619 -1050 2649 -1028
rect 2712 -1050 2742 -1028
rect 2798 -1050 2828 -1028
rect 2942 -1050 2972 -1028
rect 3028 -1050 3058 -1028
rect 3121 -1050 3151 -1028
rect 3199 -1050 3229 -1028
rect 3292 -1050 3322 -1028
rect 3378 -1050 3408 -1028
rect 3522 -1050 3552 -1028
rect 3608 -1050 3638 -1028
rect 3701 -1050 3731 -1028
rect 3779 -1050 3809 -1028
rect 3872 -1050 3902 -1028
rect 3958 -1050 3988 -1028
rect 4102 -1050 4132 -1028
rect 4188 -1050 4218 -1028
rect 4281 -1050 4311 -1028
rect 4359 -1050 4389 -1028
rect 4452 -1050 4482 -1028
rect 4538 -1050 4568 -1028
rect 4682 -1050 4712 -1028
rect 4768 -1050 4798 -1028
rect 4861 -1050 4891 -1028
rect 4939 -1050 4969 -1028
rect 5032 -1050 5062 -1028
rect 5118 -1050 5148 -1028
rect 5262 -1050 5292 -1028
rect 5348 -1050 5378 -1028
rect 5441 -1050 5471 -1028
rect 5519 -1050 5549 -1028
rect 5612 -1050 5642 -1028
rect 5698 -1050 5728 -1028
rect 5842 -1050 5872 -1028
rect 5928 -1050 5958 -1028
rect 6021 -1050 6051 -1028
rect 6099 -1050 6129 -1028
rect 6192 -1050 6222 -1028
rect 6278 -1050 6308 -1028
rect 6422 -1050 6452 -1028
rect 6508 -1050 6538 -1028
rect 6601 -1050 6631 -1028
rect 6679 -1050 6709 -1028
rect 6772 -1050 6802 -1028
rect 6858 -1050 6888 -1028
rect -1 -1096 6931 -1066
rect 106 -1124 136 -1096
rect 221 -1134 251 -1112
rect 299 -1134 329 -1112
rect 414 -1124 444 -1096
rect 106 -1174 136 -1152
rect 686 -1124 716 -1096
rect 801 -1134 831 -1112
rect 879 -1134 909 -1112
rect 994 -1124 1024 -1096
rect 221 -1195 251 -1162
rect 42 -1256 72 -1234
rect 128 -1256 143 -1222
rect 221 -1256 251 -1229
rect 299 -1195 329 -1162
rect 414 -1174 444 -1152
rect 686 -1174 716 -1152
rect 1266 -1124 1296 -1096
rect 1381 -1134 1411 -1112
rect 1459 -1134 1489 -1112
rect 1574 -1124 1604 -1096
rect 801 -1195 831 -1162
rect 299 -1256 329 -1229
rect 407 -1256 422 -1222
rect 478 -1256 508 -1234
rect 622 -1256 652 -1234
rect 708 -1256 723 -1222
rect 801 -1256 831 -1229
rect 879 -1195 909 -1162
rect 994 -1174 1024 -1152
rect 1266 -1174 1296 -1152
rect 1846 -1124 1876 -1096
rect 1961 -1134 1991 -1112
rect 2039 -1134 2069 -1112
rect 2154 -1124 2184 -1096
rect 1381 -1195 1411 -1162
rect 879 -1256 909 -1229
rect 987 -1256 1002 -1222
rect 1058 -1256 1088 -1234
rect 1202 -1256 1232 -1234
rect 1288 -1256 1303 -1222
rect 1381 -1256 1411 -1229
rect 1459 -1195 1489 -1162
rect 1574 -1174 1604 -1152
rect 1846 -1174 1876 -1152
rect 2426 -1124 2456 -1096
rect 2541 -1134 2571 -1112
rect 2619 -1134 2649 -1112
rect 2734 -1124 2764 -1096
rect 1961 -1195 1991 -1162
rect 1459 -1256 1489 -1229
rect 1567 -1256 1582 -1222
rect 1638 -1256 1668 -1234
rect 1782 -1256 1812 -1234
rect 1868 -1256 1883 -1222
rect 1961 -1256 1991 -1229
rect 2039 -1195 2069 -1162
rect 2154 -1174 2184 -1152
rect 2426 -1174 2456 -1152
rect 3006 -1124 3036 -1096
rect 3121 -1134 3151 -1112
rect 3199 -1134 3229 -1112
rect 3314 -1124 3344 -1096
rect 2541 -1195 2571 -1162
rect 2039 -1256 2069 -1229
rect 2147 -1256 2162 -1222
rect 2218 -1256 2248 -1234
rect 2362 -1256 2392 -1234
rect 2448 -1256 2463 -1222
rect 2541 -1256 2571 -1229
rect 2619 -1195 2649 -1162
rect 2734 -1174 2764 -1152
rect 3006 -1174 3036 -1152
rect 3586 -1124 3616 -1096
rect 3701 -1134 3731 -1112
rect 3779 -1134 3809 -1112
rect 3894 -1124 3924 -1096
rect 3121 -1195 3151 -1162
rect 2619 -1256 2649 -1229
rect 2727 -1256 2742 -1222
rect 2798 -1256 2828 -1234
rect 2942 -1256 2972 -1234
rect 3028 -1256 3043 -1222
rect 3121 -1256 3151 -1229
rect 3199 -1195 3229 -1162
rect 3314 -1174 3344 -1152
rect 3586 -1174 3616 -1152
rect 4166 -1124 4196 -1096
rect 4281 -1134 4311 -1112
rect 4359 -1134 4389 -1112
rect 4474 -1124 4504 -1096
rect 3701 -1195 3731 -1162
rect 3199 -1256 3229 -1229
rect 3307 -1256 3322 -1222
rect 3378 -1256 3408 -1234
rect 3522 -1256 3552 -1234
rect 3608 -1256 3623 -1222
rect 3701 -1256 3731 -1229
rect 3779 -1195 3809 -1162
rect 3894 -1174 3924 -1152
rect 4166 -1174 4196 -1152
rect 4746 -1124 4776 -1096
rect 4861 -1134 4891 -1112
rect 4939 -1134 4969 -1112
rect 5054 -1124 5084 -1096
rect 4281 -1195 4311 -1162
rect 3779 -1256 3809 -1229
rect 3887 -1256 3902 -1222
rect 3958 -1256 3988 -1234
rect 4102 -1256 4132 -1234
rect 4188 -1256 4203 -1222
rect 4281 -1256 4311 -1229
rect 4359 -1195 4389 -1162
rect 4474 -1174 4504 -1152
rect 4746 -1174 4776 -1152
rect 5326 -1124 5356 -1096
rect 5441 -1134 5471 -1112
rect 5519 -1134 5549 -1112
rect 5634 -1124 5664 -1096
rect 4861 -1195 4891 -1162
rect 4359 -1256 4389 -1229
rect 4467 -1256 4482 -1222
rect 4538 -1256 4568 -1234
rect 4682 -1256 4712 -1234
rect 4768 -1256 4783 -1222
rect 4861 -1256 4891 -1229
rect 4939 -1195 4969 -1162
rect 5054 -1174 5084 -1152
rect 5326 -1174 5356 -1152
rect 5906 -1124 5936 -1096
rect 6021 -1134 6051 -1112
rect 6099 -1134 6129 -1112
rect 6214 -1124 6244 -1096
rect 5441 -1195 5471 -1162
rect 4939 -1256 4969 -1229
rect 5047 -1256 5062 -1222
rect 5118 -1256 5148 -1234
rect 5262 -1256 5292 -1234
rect 5348 -1256 5363 -1222
rect 5441 -1256 5471 -1229
rect 5519 -1195 5549 -1162
rect 5634 -1174 5664 -1152
rect 5906 -1174 5936 -1152
rect 6486 -1124 6516 -1096
rect 6601 -1134 6631 -1112
rect 6679 -1134 6709 -1112
rect 6794 -1124 6824 -1096
rect 6021 -1195 6051 -1162
rect 5519 -1256 5549 -1229
rect 5627 -1256 5642 -1222
rect 5698 -1256 5728 -1234
rect 5842 -1256 5872 -1234
rect 5928 -1256 5943 -1222
rect 6021 -1256 6051 -1229
rect 6099 -1195 6129 -1162
rect 6214 -1174 6244 -1152
rect 6486 -1174 6516 -1152
rect 6601 -1195 6631 -1162
rect 6099 -1256 6129 -1229
rect 6207 -1256 6222 -1222
rect 6278 -1256 6308 -1234
rect 6422 -1256 6452 -1234
rect 6508 -1256 6523 -1222
rect 6601 -1256 6631 -1229
rect 6679 -1195 6709 -1162
rect 6794 -1174 6824 -1152
rect 6679 -1256 6709 -1229
rect 6787 -1256 6802 -1222
rect 6858 -1256 6888 -1234
rect 128 -1270 158 -1256
rect 392 -1270 422 -1256
rect 708 -1270 738 -1256
rect 972 -1270 1002 -1256
rect 1288 -1270 1318 -1256
rect 1552 -1270 1582 -1256
rect 1868 -1270 1898 -1256
rect 2132 -1270 2162 -1256
rect 2448 -1270 2478 -1256
rect 2712 -1270 2742 -1256
rect 3028 -1270 3058 -1256
rect 3292 -1270 3322 -1256
rect 3608 -1270 3638 -1256
rect 3872 -1270 3902 -1256
rect 4188 -1270 4218 -1256
rect 4452 -1270 4482 -1256
rect 4768 -1270 4798 -1256
rect 5032 -1270 5062 -1256
rect 5348 -1270 5378 -1256
rect 5612 -1270 5642 -1256
rect 5928 -1270 5958 -1256
rect 6192 -1270 6222 -1256
rect 6508 -1270 6538 -1256
rect 6772 -1270 6802 -1256
rect 42 -1320 72 -1298
rect 128 -1320 158 -1298
rect 221 -1320 251 -1298
rect 299 -1320 329 -1298
rect 392 -1320 422 -1298
rect 478 -1320 508 -1298
rect 622 -1320 652 -1298
rect 708 -1320 738 -1298
rect 801 -1320 831 -1298
rect 879 -1320 909 -1298
rect 972 -1320 1002 -1298
rect 1058 -1320 1088 -1298
rect 1202 -1320 1232 -1298
rect 1288 -1320 1318 -1298
rect 1381 -1320 1411 -1298
rect 1459 -1320 1489 -1298
rect 1552 -1320 1582 -1298
rect 1638 -1320 1668 -1298
rect 1782 -1320 1812 -1298
rect 1868 -1320 1898 -1298
rect 1961 -1320 1991 -1298
rect 2039 -1320 2069 -1298
rect 2132 -1320 2162 -1298
rect 2218 -1320 2248 -1298
rect 2362 -1320 2392 -1298
rect 2448 -1320 2478 -1298
rect 2541 -1320 2571 -1298
rect 2619 -1320 2649 -1298
rect 2712 -1320 2742 -1298
rect 2798 -1320 2828 -1298
rect 2942 -1320 2972 -1298
rect 3028 -1320 3058 -1298
rect 3121 -1320 3151 -1298
rect 3199 -1320 3229 -1298
rect 3292 -1320 3322 -1298
rect 3378 -1320 3408 -1298
rect 3522 -1320 3552 -1298
rect 3608 -1320 3638 -1298
rect 3701 -1320 3731 -1298
rect 3779 -1320 3809 -1298
rect 3872 -1320 3902 -1298
rect 3958 -1320 3988 -1298
rect 4102 -1320 4132 -1298
rect 4188 -1320 4218 -1298
rect 4281 -1320 4311 -1298
rect 4359 -1320 4389 -1298
rect 4452 -1320 4482 -1298
rect 4538 -1320 4568 -1298
rect 4682 -1320 4712 -1298
rect 4768 -1320 4798 -1298
rect 4861 -1320 4891 -1298
rect 4939 -1320 4969 -1298
rect 5032 -1320 5062 -1298
rect 5118 -1320 5148 -1298
rect 5262 -1320 5292 -1298
rect 5348 -1320 5378 -1298
rect 5441 -1320 5471 -1298
rect 5519 -1320 5549 -1298
rect 5612 -1320 5642 -1298
rect 5698 -1320 5728 -1298
rect 5842 -1320 5872 -1298
rect 5928 -1320 5958 -1298
rect 6021 -1320 6051 -1298
rect 6099 -1320 6129 -1298
rect 6192 -1320 6222 -1298
rect 6278 -1320 6308 -1298
rect 6422 -1320 6452 -1298
rect 6508 -1320 6538 -1298
rect 6601 -1320 6631 -1298
rect 6679 -1320 6709 -1298
rect 6772 -1320 6802 -1298
rect 6858 -1320 6888 -1298
rect -1 -1366 6931 -1336
rect 106 -1394 136 -1366
rect 221 -1404 251 -1382
rect 299 -1404 329 -1382
rect 414 -1394 444 -1366
rect 106 -1444 136 -1422
rect 686 -1394 716 -1366
rect 801 -1404 831 -1382
rect 879 -1404 909 -1382
rect 994 -1394 1024 -1366
rect 221 -1465 251 -1432
rect 42 -1526 72 -1504
rect 128 -1526 143 -1492
rect 221 -1526 251 -1499
rect 299 -1465 329 -1432
rect 414 -1444 444 -1422
rect 686 -1444 716 -1422
rect 1266 -1394 1296 -1366
rect 1381 -1404 1411 -1382
rect 1459 -1404 1489 -1382
rect 1574 -1394 1604 -1366
rect 801 -1465 831 -1432
rect 299 -1526 329 -1499
rect 407 -1526 422 -1492
rect 478 -1526 508 -1504
rect 622 -1526 652 -1504
rect 708 -1526 723 -1492
rect 801 -1526 831 -1499
rect 879 -1465 909 -1432
rect 994 -1444 1024 -1422
rect 1266 -1444 1296 -1422
rect 1846 -1394 1876 -1366
rect 1961 -1404 1991 -1382
rect 2039 -1404 2069 -1382
rect 2154 -1394 2184 -1366
rect 1381 -1465 1411 -1432
rect 879 -1526 909 -1499
rect 987 -1526 1002 -1492
rect 1058 -1526 1088 -1504
rect 1202 -1526 1232 -1504
rect 1288 -1526 1303 -1492
rect 1381 -1526 1411 -1499
rect 1459 -1465 1489 -1432
rect 1574 -1444 1604 -1422
rect 1846 -1444 1876 -1422
rect 2426 -1394 2456 -1366
rect 2541 -1404 2571 -1382
rect 2619 -1404 2649 -1382
rect 2734 -1394 2764 -1366
rect 1961 -1465 1991 -1432
rect 1459 -1526 1489 -1499
rect 1567 -1526 1582 -1492
rect 1638 -1526 1668 -1504
rect 1782 -1526 1812 -1504
rect 1868 -1526 1883 -1492
rect 1961 -1526 1991 -1499
rect 2039 -1465 2069 -1432
rect 2154 -1444 2184 -1422
rect 2426 -1444 2456 -1422
rect 3006 -1394 3036 -1366
rect 3121 -1404 3151 -1382
rect 3199 -1404 3229 -1382
rect 3314 -1394 3344 -1366
rect 2541 -1465 2571 -1432
rect 2039 -1526 2069 -1499
rect 2147 -1526 2162 -1492
rect 2218 -1526 2248 -1504
rect 2362 -1526 2392 -1504
rect 2448 -1526 2463 -1492
rect 2541 -1526 2571 -1499
rect 2619 -1465 2649 -1432
rect 2734 -1444 2764 -1422
rect 3006 -1444 3036 -1422
rect 3586 -1394 3616 -1366
rect 3701 -1404 3731 -1382
rect 3779 -1404 3809 -1382
rect 3894 -1394 3924 -1366
rect 3121 -1465 3151 -1432
rect 2619 -1526 2649 -1499
rect 2727 -1526 2742 -1492
rect 2798 -1526 2828 -1504
rect 2942 -1526 2972 -1504
rect 3028 -1526 3043 -1492
rect 3121 -1526 3151 -1499
rect 3199 -1465 3229 -1432
rect 3314 -1444 3344 -1422
rect 3586 -1444 3616 -1422
rect 4166 -1394 4196 -1366
rect 4281 -1404 4311 -1382
rect 4359 -1404 4389 -1382
rect 4474 -1394 4504 -1366
rect 3701 -1465 3731 -1432
rect 3199 -1526 3229 -1499
rect 3307 -1526 3322 -1492
rect 3378 -1526 3408 -1504
rect 3522 -1526 3552 -1504
rect 3608 -1526 3623 -1492
rect 3701 -1526 3731 -1499
rect 3779 -1465 3809 -1432
rect 3894 -1444 3924 -1422
rect 4166 -1444 4196 -1422
rect 4746 -1394 4776 -1366
rect 4861 -1404 4891 -1382
rect 4939 -1404 4969 -1382
rect 5054 -1394 5084 -1366
rect 4281 -1465 4311 -1432
rect 3779 -1526 3809 -1499
rect 3887 -1526 3902 -1492
rect 3958 -1526 3988 -1504
rect 4102 -1526 4132 -1504
rect 4188 -1526 4203 -1492
rect 4281 -1526 4311 -1499
rect 4359 -1465 4389 -1432
rect 4474 -1444 4504 -1422
rect 4746 -1444 4776 -1422
rect 5326 -1394 5356 -1366
rect 5441 -1404 5471 -1382
rect 5519 -1404 5549 -1382
rect 5634 -1394 5664 -1366
rect 4861 -1465 4891 -1432
rect 4359 -1526 4389 -1499
rect 4467 -1526 4482 -1492
rect 4538 -1526 4568 -1504
rect 4682 -1526 4712 -1504
rect 4768 -1526 4783 -1492
rect 4861 -1526 4891 -1499
rect 4939 -1465 4969 -1432
rect 5054 -1444 5084 -1422
rect 5326 -1444 5356 -1422
rect 5906 -1394 5936 -1366
rect 6021 -1404 6051 -1382
rect 6099 -1404 6129 -1382
rect 6214 -1394 6244 -1366
rect 5441 -1465 5471 -1432
rect 4939 -1526 4969 -1499
rect 5047 -1526 5062 -1492
rect 5118 -1526 5148 -1504
rect 5262 -1526 5292 -1504
rect 5348 -1526 5363 -1492
rect 5441 -1526 5471 -1499
rect 5519 -1465 5549 -1432
rect 5634 -1444 5664 -1422
rect 5906 -1444 5936 -1422
rect 6486 -1394 6516 -1366
rect 6601 -1404 6631 -1382
rect 6679 -1404 6709 -1382
rect 6794 -1394 6824 -1366
rect 6021 -1465 6051 -1432
rect 5519 -1526 5549 -1499
rect 5627 -1526 5642 -1492
rect 5698 -1526 5728 -1504
rect 5842 -1526 5872 -1504
rect 5928 -1526 5943 -1492
rect 6021 -1526 6051 -1499
rect 6099 -1465 6129 -1432
rect 6214 -1444 6244 -1422
rect 6486 -1444 6516 -1422
rect 6601 -1465 6631 -1432
rect 6099 -1526 6129 -1499
rect 6207 -1526 6222 -1492
rect 6278 -1526 6308 -1504
rect 6422 -1526 6452 -1504
rect 6508 -1526 6523 -1492
rect 6601 -1526 6631 -1499
rect 6679 -1465 6709 -1432
rect 6794 -1444 6824 -1422
rect 6679 -1526 6709 -1499
rect 6787 -1526 6802 -1492
rect 6858 -1526 6888 -1504
rect 128 -1540 158 -1526
rect 392 -1540 422 -1526
rect 708 -1540 738 -1526
rect 972 -1540 1002 -1526
rect 1288 -1540 1318 -1526
rect 1552 -1540 1582 -1526
rect 1868 -1540 1898 -1526
rect 2132 -1540 2162 -1526
rect 2448 -1540 2478 -1526
rect 2712 -1540 2742 -1526
rect 3028 -1540 3058 -1526
rect 3292 -1540 3322 -1526
rect 3608 -1540 3638 -1526
rect 3872 -1540 3902 -1526
rect 4188 -1540 4218 -1526
rect 4452 -1540 4482 -1526
rect 4768 -1540 4798 -1526
rect 5032 -1540 5062 -1526
rect 5348 -1540 5378 -1526
rect 5612 -1540 5642 -1526
rect 5928 -1540 5958 -1526
rect 6192 -1540 6222 -1526
rect 6508 -1540 6538 -1526
rect 6772 -1540 6802 -1526
rect 42 -1590 72 -1568
rect 128 -1590 158 -1568
rect 221 -1590 251 -1568
rect 299 -1590 329 -1568
rect 392 -1590 422 -1568
rect 478 -1590 508 -1568
rect 622 -1590 652 -1568
rect 708 -1590 738 -1568
rect 801 -1590 831 -1568
rect 879 -1590 909 -1568
rect 972 -1590 1002 -1568
rect 1058 -1590 1088 -1568
rect 1202 -1590 1232 -1568
rect 1288 -1590 1318 -1568
rect 1381 -1590 1411 -1568
rect 1459 -1590 1489 -1568
rect 1552 -1590 1582 -1568
rect 1638 -1590 1668 -1568
rect 1782 -1590 1812 -1568
rect 1868 -1590 1898 -1568
rect 1961 -1590 1991 -1568
rect 2039 -1590 2069 -1568
rect 2132 -1590 2162 -1568
rect 2218 -1590 2248 -1568
rect 2362 -1590 2392 -1568
rect 2448 -1590 2478 -1568
rect 2541 -1590 2571 -1568
rect 2619 -1590 2649 -1568
rect 2712 -1590 2742 -1568
rect 2798 -1590 2828 -1568
rect 2942 -1590 2972 -1568
rect 3028 -1590 3058 -1568
rect 3121 -1590 3151 -1568
rect 3199 -1590 3229 -1568
rect 3292 -1590 3322 -1568
rect 3378 -1590 3408 -1568
rect 3522 -1590 3552 -1568
rect 3608 -1590 3638 -1568
rect 3701 -1590 3731 -1568
rect 3779 -1590 3809 -1568
rect 3872 -1590 3902 -1568
rect 3958 -1590 3988 -1568
rect 4102 -1590 4132 -1568
rect 4188 -1590 4218 -1568
rect 4281 -1590 4311 -1568
rect 4359 -1590 4389 -1568
rect 4452 -1590 4482 -1568
rect 4538 -1590 4568 -1568
rect 4682 -1590 4712 -1568
rect 4768 -1590 4798 -1568
rect 4861 -1590 4891 -1568
rect 4939 -1590 4969 -1568
rect 5032 -1590 5062 -1568
rect 5118 -1590 5148 -1568
rect 5262 -1590 5292 -1568
rect 5348 -1590 5378 -1568
rect 5441 -1590 5471 -1568
rect 5519 -1590 5549 -1568
rect 5612 -1590 5642 -1568
rect 5698 -1590 5728 -1568
rect 5842 -1590 5872 -1568
rect 5928 -1590 5958 -1568
rect 6021 -1590 6051 -1568
rect 6099 -1590 6129 -1568
rect 6192 -1590 6222 -1568
rect 6278 -1590 6308 -1568
rect 6422 -1590 6452 -1568
rect 6508 -1590 6538 -1568
rect 6601 -1590 6631 -1568
rect 6679 -1590 6709 -1568
rect 6772 -1590 6802 -1568
rect 6858 -1590 6888 -1568
rect -1 -1636 6931 -1606
rect 106 -1664 136 -1636
rect 221 -1674 251 -1652
rect 299 -1674 329 -1652
rect 414 -1664 444 -1636
rect 106 -1714 136 -1692
rect 686 -1664 716 -1636
rect 801 -1674 831 -1652
rect 879 -1674 909 -1652
rect 994 -1664 1024 -1636
rect 221 -1735 251 -1702
rect 42 -1796 72 -1774
rect 128 -1796 143 -1762
rect 221 -1796 251 -1769
rect 299 -1735 329 -1702
rect 414 -1714 444 -1692
rect 686 -1714 716 -1692
rect 1266 -1664 1296 -1636
rect 1381 -1674 1411 -1652
rect 1459 -1674 1489 -1652
rect 1574 -1664 1604 -1636
rect 801 -1735 831 -1702
rect 299 -1796 329 -1769
rect 407 -1796 422 -1762
rect 478 -1796 508 -1774
rect 622 -1796 652 -1774
rect 708 -1796 723 -1762
rect 801 -1796 831 -1769
rect 879 -1735 909 -1702
rect 994 -1714 1024 -1692
rect 1266 -1714 1296 -1692
rect 1846 -1664 1876 -1636
rect 1961 -1674 1991 -1652
rect 2039 -1674 2069 -1652
rect 2154 -1664 2184 -1636
rect 1381 -1735 1411 -1702
rect 879 -1796 909 -1769
rect 987 -1796 1002 -1762
rect 1058 -1796 1088 -1774
rect 1202 -1796 1232 -1774
rect 1288 -1796 1303 -1762
rect 1381 -1796 1411 -1769
rect 1459 -1735 1489 -1702
rect 1574 -1714 1604 -1692
rect 1846 -1714 1876 -1692
rect 2426 -1664 2456 -1636
rect 2541 -1674 2571 -1652
rect 2619 -1674 2649 -1652
rect 2734 -1664 2764 -1636
rect 1961 -1735 1991 -1702
rect 1459 -1796 1489 -1769
rect 1567 -1796 1582 -1762
rect 1638 -1796 1668 -1774
rect 1782 -1796 1812 -1774
rect 1868 -1796 1883 -1762
rect 1961 -1796 1991 -1769
rect 2039 -1735 2069 -1702
rect 2154 -1714 2184 -1692
rect 2426 -1714 2456 -1692
rect 3006 -1664 3036 -1636
rect 3121 -1674 3151 -1652
rect 3199 -1674 3229 -1652
rect 3314 -1664 3344 -1636
rect 2541 -1735 2571 -1702
rect 2039 -1796 2069 -1769
rect 2147 -1796 2162 -1762
rect 2218 -1796 2248 -1774
rect 2362 -1796 2392 -1774
rect 2448 -1796 2463 -1762
rect 2541 -1796 2571 -1769
rect 2619 -1735 2649 -1702
rect 2734 -1714 2764 -1692
rect 3006 -1714 3036 -1692
rect 3586 -1664 3616 -1636
rect 3701 -1674 3731 -1652
rect 3779 -1674 3809 -1652
rect 3894 -1664 3924 -1636
rect 3121 -1735 3151 -1702
rect 2619 -1796 2649 -1769
rect 2727 -1796 2742 -1762
rect 2798 -1796 2828 -1774
rect 2942 -1796 2972 -1774
rect 3028 -1796 3043 -1762
rect 3121 -1796 3151 -1769
rect 3199 -1735 3229 -1702
rect 3314 -1714 3344 -1692
rect 3586 -1714 3616 -1692
rect 4166 -1664 4196 -1636
rect 4281 -1674 4311 -1652
rect 4359 -1674 4389 -1652
rect 4474 -1664 4504 -1636
rect 3701 -1735 3731 -1702
rect 3199 -1796 3229 -1769
rect 3307 -1796 3322 -1762
rect 3378 -1796 3408 -1774
rect 3522 -1796 3552 -1774
rect 3608 -1796 3623 -1762
rect 3701 -1796 3731 -1769
rect 3779 -1735 3809 -1702
rect 3894 -1714 3924 -1692
rect 4166 -1714 4196 -1692
rect 4746 -1664 4776 -1636
rect 4861 -1674 4891 -1652
rect 4939 -1674 4969 -1652
rect 5054 -1664 5084 -1636
rect 4281 -1735 4311 -1702
rect 3779 -1796 3809 -1769
rect 3887 -1796 3902 -1762
rect 3958 -1796 3988 -1774
rect 4102 -1796 4132 -1774
rect 4188 -1796 4203 -1762
rect 4281 -1796 4311 -1769
rect 4359 -1735 4389 -1702
rect 4474 -1714 4504 -1692
rect 4746 -1714 4776 -1692
rect 5326 -1664 5356 -1636
rect 5441 -1674 5471 -1652
rect 5519 -1674 5549 -1652
rect 5634 -1664 5664 -1636
rect 4861 -1735 4891 -1702
rect 4359 -1796 4389 -1769
rect 4467 -1796 4482 -1762
rect 4538 -1796 4568 -1774
rect 4682 -1796 4712 -1774
rect 4768 -1796 4783 -1762
rect 4861 -1796 4891 -1769
rect 4939 -1735 4969 -1702
rect 5054 -1714 5084 -1692
rect 5326 -1714 5356 -1692
rect 5906 -1664 5936 -1636
rect 6021 -1674 6051 -1652
rect 6099 -1674 6129 -1652
rect 6214 -1664 6244 -1636
rect 5441 -1735 5471 -1702
rect 4939 -1796 4969 -1769
rect 5047 -1796 5062 -1762
rect 5118 -1796 5148 -1774
rect 5262 -1796 5292 -1774
rect 5348 -1796 5363 -1762
rect 5441 -1796 5471 -1769
rect 5519 -1735 5549 -1702
rect 5634 -1714 5664 -1692
rect 5906 -1714 5936 -1692
rect 6486 -1664 6516 -1636
rect 6601 -1674 6631 -1652
rect 6679 -1674 6709 -1652
rect 6794 -1664 6824 -1636
rect 6021 -1735 6051 -1702
rect 5519 -1796 5549 -1769
rect 5627 -1796 5642 -1762
rect 5698 -1796 5728 -1774
rect 5842 -1796 5872 -1774
rect 5928 -1796 5943 -1762
rect 6021 -1796 6051 -1769
rect 6099 -1735 6129 -1702
rect 6214 -1714 6244 -1692
rect 6486 -1714 6516 -1692
rect 6601 -1735 6631 -1702
rect 6099 -1796 6129 -1769
rect 6207 -1796 6222 -1762
rect 6278 -1796 6308 -1774
rect 6422 -1796 6452 -1774
rect 6508 -1796 6523 -1762
rect 6601 -1796 6631 -1769
rect 6679 -1735 6709 -1702
rect 6794 -1714 6824 -1692
rect 6679 -1796 6709 -1769
rect 6787 -1796 6802 -1762
rect 6858 -1796 6888 -1774
rect 128 -1810 158 -1796
rect 392 -1810 422 -1796
rect 708 -1810 738 -1796
rect 972 -1810 1002 -1796
rect 1288 -1810 1318 -1796
rect 1552 -1810 1582 -1796
rect 1868 -1810 1898 -1796
rect 2132 -1810 2162 -1796
rect 2448 -1810 2478 -1796
rect 2712 -1810 2742 -1796
rect 3028 -1810 3058 -1796
rect 3292 -1810 3322 -1796
rect 3608 -1810 3638 -1796
rect 3872 -1810 3902 -1796
rect 4188 -1810 4218 -1796
rect 4452 -1810 4482 -1796
rect 4768 -1810 4798 -1796
rect 5032 -1810 5062 -1796
rect 5348 -1810 5378 -1796
rect 5612 -1810 5642 -1796
rect 5928 -1810 5958 -1796
rect 6192 -1810 6222 -1796
rect 6508 -1810 6538 -1796
rect 6772 -1810 6802 -1796
rect 42 -1860 72 -1838
rect 128 -1860 158 -1838
rect 221 -1860 251 -1838
rect 299 -1860 329 -1838
rect 392 -1860 422 -1838
rect 478 -1860 508 -1838
rect 622 -1860 652 -1838
rect 708 -1860 738 -1838
rect 801 -1860 831 -1838
rect 879 -1860 909 -1838
rect 972 -1860 1002 -1838
rect 1058 -1860 1088 -1838
rect 1202 -1860 1232 -1838
rect 1288 -1860 1318 -1838
rect 1381 -1860 1411 -1838
rect 1459 -1860 1489 -1838
rect 1552 -1860 1582 -1838
rect 1638 -1860 1668 -1838
rect 1782 -1860 1812 -1838
rect 1868 -1860 1898 -1838
rect 1961 -1860 1991 -1838
rect 2039 -1860 2069 -1838
rect 2132 -1860 2162 -1838
rect 2218 -1860 2248 -1838
rect 2362 -1860 2392 -1838
rect 2448 -1860 2478 -1838
rect 2541 -1860 2571 -1838
rect 2619 -1860 2649 -1838
rect 2712 -1860 2742 -1838
rect 2798 -1860 2828 -1838
rect 2942 -1860 2972 -1838
rect 3028 -1860 3058 -1838
rect 3121 -1860 3151 -1838
rect 3199 -1860 3229 -1838
rect 3292 -1860 3322 -1838
rect 3378 -1860 3408 -1838
rect 3522 -1860 3552 -1838
rect 3608 -1860 3638 -1838
rect 3701 -1860 3731 -1838
rect 3779 -1860 3809 -1838
rect 3872 -1860 3902 -1838
rect 3958 -1860 3988 -1838
rect 4102 -1860 4132 -1838
rect 4188 -1860 4218 -1838
rect 4281 -1860 4311 -1838
rect 4359 -1860 4389 -1838
rect 4452 -1860 4482 -1838
rect 4538 -1860 4568 -1838
rect 4682 -1860 4712 -1838
rect 4768 -1860 4798 -1838
rect 4861 -1860 4891 -1838
rect 4939 -1860 4969 -1838
rect 5032 -1860 5062 -1838
rect 5118 -1860 5148 -1838
rect 5262 -1860 5292 -1838
rect 5348 -1860 5378 -1838
rect 5441 -1860 5471 -1838
rect 5519 -1860 5549 -1838
rect 5612 -1860 5642 -1838
rect 5698 -1860 5728 -1838
rect 5842 -1860 5872 -1838
rect 5928 -1860 5958 -1838
rect 6021 -1860 6051 -1838
rect 6099 -1860 6129 -1838
rect 6192 -1860 6222 -1838
rect 6278 -1860 6308 -1838
rect 6422 -1860 6452 -1838
rect 6508 -1860 6538 -1838
rect 6601 -1860 6631 -1838
rect 6679 -1860 6709 -1838
rect 6772 -1860 6802 -1838
rect 6858 -1860 6888 -1838
rect -1 -1906 6931 -1876
rect 106 -1934 136 -1906
rect 221 -1944 251 -1922
rect 299 -1944 329 -1922
rect 414 -1934 444 -1906
rect 106 -1984 136 -1962
rect 686 -1934 716 -1906
rect 801 -1944 831 -1922
rect 879 -1944 909 -1922
rect 994 -1934 1024 -1906
rect 221 -2005 251 -1972
rect 42 -2066 72 -2044
rect 128 -2066 143 -2032
rect 221 -2066 251 -2039
rect 299 -2005 329 -1972
rect 414 -1984 444 -1962
rect 686 -1984 716 -1962
rect 1266 -1934 1296 -1906
rect 1381 -1944 1411 -1922
rect 1459 -1944 1489 -1922
rect 1574 -1934 1604 -1906
rect 801 -2005 831 -1972
rect 299 -2066 329 -2039
rect 407 -2066 422 -2032
rect 478 -2066 508 -2044
rect 622 -2066 652 -2044
rect 708 -2066 723 -2032
rect 801 -2066 831 -2039
rect 879 -2005 909 -1972
rect 994 -1984 1024 -1962
rect 1266 -1984 1296 -1962
rect 1846 -1934 1876 -1906
rect 1961 -1944 1991 -1922
rect 2039 -1944 2069 -1922
rect 2154 -1934 2184 -1906
rect 1381 -2005 1411 -1972
rect 879 -2066 909 -2039
rect 987 -2066 1002 -2032
rect 1058 -2066 1088 -2044
rect 1202 -2066 1232 -2044
rect 1288 -2066 1303 -2032
rect 1381 -2066 1411 -2039
rect 1459 -2005 1489 -1972
rect 1574 -1984 1604 -1962
rect 1846 -1984 1876 -1962
rect 2426 -1934 2456 -1906
rect 2541 -1944 2571 -1922
rect 2619 -1944 2649 -1922
rect 2734 -1934 2764 -1906
rect 1961 -2005 1991 -1972
rect 1459 -2066 1489 -2039
rect 1567 -2066 1582 -2032
rect 1638 -2066 1668 -2044
rect 1782 -2066 1812 -2044
rect 1868 -2066 1883 -2032
rect 1961 -2066 1991 -2039
rect 2039 -2005 2069 -1972
rect 2154 -1984 2184 -1962
rect 2426 -1984 2456 -1962
rect 3006 -1934 3036 -1906
rect 3121 -1944 3151 -1922
rect 3199 -1944 3229 -1922
rect 3314 -1934 3344 -1906
rect 2541 -2005 2571 -1972
rect 2039 -2066 2069 -2039
rect 2147 -2066 2162 -2032
rect 2218 -2066 2248 -2044
rect 2362 -2066 2392 -2044
rect 2448 -2066 2463 -2032
rect 2541 -2066 2571 -2039
rect 2619 -2005 2649 -1972
rect 2734 -1984 2764 -1962
rect 3006 -1984 3036 -1962
rect 3586 -1934 3616 -1906
rect 3701 -1944 3731 -1922
rect 3779 -1944 3809 -1922
rect 3894 -1934 3924 -1906
rect 3121 -2005 3151 -1972
rect 2619 -2066 2649 -2039
rect 2727 -2066 2742 -2032
rect 2798 -2066 2828 -2044
rect 2942 -2066 2972 -2044
rect 3028 -2066 3043 -2032
rect 3121 -2066 3151 -2039
rect 3199 -2005 3229 -1972
rect 3314 -1984 3344 -1962
rect 3586 -1984 3616 -1962
rect 4166 -1934 4196 -1906
rect 4281 -1944 4311 -1922
rect 4359 -1944 4389 -1922
rect 4474 -1934 4504 -1906
rect 3701 -2005 3731 -1972
rect 3199 -2066 3229 -2039
rect 3307 -2066 3322 -2032
rect 3378 -2066 3408 -2044
rect 3522 -2066 3552 -2044
rect 3608 -2066 3623 -2032
rect 3701 -2066 3731 -2039
rect 3779 -2005 3809 -1972
rect 3894 -1984 3924 -1962
rect 4166 -1984 4196 -1962
rect 4746 -1934 4776 -1906
rect 4861 -1944 4891 -1922
rect 4939 -1944 4969 -1922
rect 5054 -1934 5084 -1906
rect 4281 -2005 4311 -1972
rect 3779 -2066 3809 -2039
rect 3887 -2066 3902 -2032
rect 3958 -2066 3988 -2044
rect 4102 -2066 4132 -2044
rect 4188 -2066 4203 -2032
rect 4281 -2066 4311 -2039
rect 4359 -2005 4389 -1972
rect 4474 -1984 4504 -1962
rect 4746 -1984 4776 -1962
rect 5326 -1934 5356 -1906
rect 5441 -1944 5471 -1922
rect 5519 -1944 5549 -1922
rect 5634 -1934 5664 -1906
rect 4861 -2005 4891 -1972
rect 4359 -2066 4389 -2039
rect 4467 -2066 4482 -2032
rect 4538 -2066 4568 -2044
rect 4682 -2066 4712 -2044
rect 4768 -2066 4783 -2032
rect 4861 -2066 4891 -2039
rect 4939 -2005 4969 -1972
rect 5054 -1984 5084 -1962
rect 5326 -1984 5356 -1962
rect 5906 -1934 5936 -1906
rect 6021 -1944 6051 -1922
rect 6099 -1944 6129 -1922
rect 6214 -1934 6244 -1906
rect 5441 -2005 5471 -1972
rect 4939 -2066 4969 -2039
rect 5047 -2066 5062 -2032
rect 5118 -2066 5148 -2044
rect 5262 -2066 5292 -2044
rect 5348 -2066 5363 -2032
rect 5441 -2066 5471 -2039
rect 5519 -2005 5549 -1972
rect 5634 -1984 5664 -1962
rect 5906 -1984 5936 -1962
rect 6486 -1934 6516 -1906
rect 6601 -1944 6631 -1922
rect 6679 -1944 6709 -1922
rect 6794 -1934 6824 -1906
rect 6021 -2005 6051 -1972
rect 5519 -2066 5549 -2039
rect 5627 -2066 5642 -2032
rect 5698 -2066 5728 -2044
rect 5842 -2066 5872 -2044
rect 5928 -2066 5943 -2032
rect 6021 -2066 6051 -2039
rect 6099 -2005 6129 -1972
rect 6214 -1984 6244 -1962
rect 6486 -1984 6516 -1962
rect 6601 -2005 6631 -1972
rect 6099 -2066 6129 -2039
rect 6207 -2066 6222 -2032
rect 6278 -2066 6308 -2044
rect 6422 -2066 6452 -2044
rect 6508 -2066 6523 -2032
rect 6601 -2066 6631 -2039
rect 6679 -2005 6709 -1972
rect 6794 -1984 6824 -1962
rect 6679 -2066 6709 -2039
rect 6787 -2066 6802 -2032
rect 6858 -2066 6888 -2044
rect 128 -2080 158 -2066
rect 392 -2080 422 -2066
rect 708 -2080 738 -2066
rect 972 -2080 1002 -2066
rect 1288 -2080 1318 -2066
rect 1552 -2080 1582 -2066
rect 1868 -2080 1898 -2066
rect 2132 -2080 2162 -2066
rect 2448 -2080 2478 -2066
rect 2712 -2080 2742 -2066
rect 3028 -2080 3058 -2066
rect 3292 -2080 3322 -2066
rect 3608 -2080 3638 -2066
rect 3872 -2080 3902 -2066
rect 4188 -2080 4218 -2066
rect 4452 -2080 4482 -2066
rect 4768 -2080 4798 -2066
rect 5032 -2080 5062 -2066
rect 5348 -2080 5378 -2066
rect 5612 -2080 5642 -2066
rect 5928 -2080 5958 -2066
rect 6192 -2080 6222 -2066
rect 6508 -2080 6538 -2066
rect 6772 -2080 6802 -2066
rect 42 -2130 72 -2108
rect 128 -2130 158 -2108
rect 221 -2130 251 -2108
rect 299 -2130 329 -2108
rect 392 -2130 422 -2108
rect 478 -2130 508 -2108
rect 622 -2130 652 -2108
rect 708 -2130 738 -2108
rect 801 -2130 831 -2108
rect 879 -2130 909 -2108
rect 972 -2130 1002 -2108
rect 1058 -2130 1088 -2108
rect 1202 -2130 1232 -2108
rect 1288 -2130 1318 -2108
rect 1381 -2130 1411 -2108
rect 1459 -2130 1489 -2108
rect 1552 -2130 1582 -2108
rect 1638 -2130 1668 -2108
rect 1782 -2130 1812 -2108
rect 1868 -2130 1898 -2108
rect 1961 -2130 1991 -2108
rect 2039 -2130 2069 -2108
rect 2132 -2130 2162 -2108
rect 2218 -2130 2248 -2108
rect 2362 -2130 2392 -2108
rect 2448 -2130 2478 -2108
rect 2541 -2130 2571 -2108
rect 2619 -2130 2649 -2108
rect 2712 -2130 2742 -2108
rect 2798 -2130 2828 -2108
rect 2942 -2130 2972 -2108
rect 3028 -2130 3058 -2108
rect 3121 -2130 3151 -2108
rect 3199 -2130 3229 -2108
rect 3292 -2130 3322 -2108
rect 3378 -2130 3408 -2108
rect 3522 -2130 3552 -2108
rect 3608 -2130 3638 -2108
rect 3701 -2130 3731 -2108
rect 3779 -2130 3809 -2108
rect 3872 -2130 3902 -2108
rect 3958 -2130 3988 -2108
rect 4102 -2130 4132 -2108
rect 4188 -2130 4218 -2108
rect 4281 -2130 4311 -2108
rect 4359 -2130 4389 -2108
rect 4452 -2130 4482 -2108
rect 4538 -2130 4568 -2108
rect 4682 -2130 4712 -2108
rect 4768 -2130 4798 -2108
rect 4861 -2130 4891 -2108
rect 4939 -2130 4969 -2108
rect 5032 -2130 5062 -2108
rect 5118 -2130 5148 -2108
rect 5262 -2130 5292 -2108
rect 5348 -2130 5378 -2108
rect 5441 -2130 5471 -2108
rect 5519 -2130 5549 -2108
rect 5612 -2130 5642 -2108
rect 5698 -2130 5728 -2108
rect 5842 -2130 5872 -2108
rect 5928 -2130 5958 -2108
rect 6021 -2130 6051 -2108
rect 6099 -2130 6129 -2108
rect 6192 -2130 6222 -2108
rect 6278 -2130 6308 -2108
rect 6422 -2130 6452 -2108
rect 6508 -2130 6538 -2108
rect 6601 -2130 6631 -2108
rect 6679 -2130 6709 -2108
rect 6772 -2130 6802 -2108
rect 6858 -2130 6888 -2108
<< polycont >>
rect 42 2006 72 2040
rect 143 1984 173 2018
rect 221 2011 251 2045
rect 299 2011 329 2045
rect 377 1984 407 2018
rect 478 2006 508 2040
rect 622 2006 652 2040
rect 723 1984 753 2018
rect 801 2011 831 2045
rect 879 2011 909 2045
rect 957 1984 987 2018
rect 1058 2006 1088 2040
rect 1202 2006 1232 2040
rect 1303 1984 1333 2018
rect 1381 2011 1411 2045
rect 1459 2011 1489 2045
rect 1537 1984 1567 2018
rect 1638 2006 1668 2040
rect 1782 2006 1812 2040
rect 1883 1984 1913 2018
rect 1961 2011 1991 2045
rect 2039 2011 2069 2045
rect 2117 1984 2147 2018
rect 2218 2006 2248 2040
rect 2362 2006 2392 2040
rect 2463 1984 2493 2018
rect 2541 2011 2571 2045
rect 2619 2011 2649 2045
rect 2697 1984 2727 2018
rect 2798 2006 2828 2040
rect 2942 2006 2972 2040
rect 3043 1984 3073 2018
rect 3121 2011 3151 2045
rect 3199 2011 3229 2045
rect 3277 1984 3307 2018
rect 3378 2006 3408 2040
rect 3522 2006 3552 2040
rect 3623 1984 3653 2018
rect 3701 2011 3731 2045
rect 3779 2011 3809 2045
rect 3857 1984 3887 2018
rect 3958 2006 3988 2040
rect 4102 2006 4132 2040
rect 4203 1984 4233 2018
rect 4281 2011 4311 2045
rect 4359 2011 4389 2045
rect 4437 1984 4467 2018
rect 4538 2006 4568 2040
rect 4682 2006 4712 2040
rect 4783 1984 4813 2018
rect 4861 2011 4891 2045
rect 4939 2011 4969 2045
rect 5017 1984 5047 2018
rect 5118 2006 5148 2040
rect 5262 2006 5292 2040
rect 5363 1984 5393 2018
rect 5441 2011 5471 2045
rect 5519 2011 5549 2045
rect 5597 1984 5627 2018
rect 5698 2006 5728 2040
rect 5842 2006 5872 2040
rect 5943 1984 5973 2018
rect 6021 2011 6051 2045
rect 6099 2011 6129 2045
rect 6177 1984 6207 2018
rect 6278 2006 6308 2040
rect 6422 2006 6452 2040
rect 6523 1984 6553 2018
rect 6601 2011 6631 2045
rect 6679 2011 6709 2045
rect 6757 1984 6787 2018
rect 6858 2006 6888 2040
rect 42 1736 72 1770
rect 143 1714 173 1748
rect 221 1741 251 1775
rect 299 1741 329 1775
rect 377 1714 407 1748
rect 478 1736 508 1770
rect 622 1736 652 1770
rect 723 1714 753 1748
rect 801 1741 831 1775
rect 879 1741 909 1775
rect 957 1714 987 1748
rect 1058 1736 1088 1770
rect 1202 1736 1232 1770
rect 1303 1714 1333 1748
rect 1381 1741 1411 1775
rect 1459 1741 1489 1775
rect 1537 1714 1567 1748
rect 1638 1736 1668 1770
rect 1782 1736 1812 1770
rect 1883 1714 1913 1748
rect 1961 1741 1991 1775
rect 2039 1741 2069 1775
rect 2117 1714 2147 1748
rect 2218 1736 2248 1770
rect 2362 1736 2392 1770
rect 2463 1714 2493 1748
rect 2541 1741 2571 1775
rect 2619 1741 2649 1775
rect 2697 1714 2727 1748
rect 2798 1736 2828 1770
rect 2942 1736 2972 1770
rect 3043 1714 3073 1748
rect 3121 1741 3151 1775
rect 3199 1741 3229 1775
rect 3277 1714 3307 1748
rect 3378 1736 3408 1770
rect 3522 1736 3552 1770
rect 3623 1714 3653 1748
rect 3701 1741 3731 1775
rect 3779 1741 3809 1775
rect 3857 1714 3887 1748
rect 3958 1736 3988 1770
rect 4102 1736 4132 1770
rect 4203 1714 4233 1748
rect 4281 1741 4311 1775
rect 4359 1741 4389 1775
rect 4437 1714 4467 1748
rect 4538 1736 4568 1770
rect 4682 1736 4712 1770
rect 4783 1714 4813 1748
rect 4861 1741 4891 1775
rect 4939 1741 4969 1775
rect 5017 1714 5047 1748
rect 5118 1736 5148 1770
rect 5262 1736 5292 1770
rect 5363 1714 5393 1748
rect 5441 1741 5471 1775
rect 5519 1741 5549 1775
rect 5597 1714 5627 1748
rect 5698 1736 5728 1770
rect 5842 1736 5872 1770
rect 5943 1714 5973 1748
rect 6021 1741 6051 1775
rect 6099 1741 6129 1775
rect 6177 1714 6207 1748
rect 6278 1736 6308 1770
rect 6422 1736 6452 1770
rect 6523 1714 6553 1748
rect 6601 1741 6631 1775
rect 6679 1741 6709 1775
rect 6757 1714 6787 1748
rect 6858 1736 6888 1770
rect 42 1466 72 1500
rect 143 1444 173 1478
rect 221 1471 251 1505
rect 299 1471 329 1505
rect 377 1444 407 1478
rect 478 1466 508 1500
rect 622 1466 652 1500
rect 723 1444 753 1478
rect 801 1471 831 1505
rect 879 1471 909 1505
rect 957 1444 987 1478
rect 1058 1466 1088 1500
rect 1202 1466 1232 1500
rect 1303 1444 1333 1478
rect 1381 1471 1411 1505
rect 1459 1471 1489 1505
rect 1537 1444 1567 1478
rect 1638 1466 1668 1500
rect 1782 1466 1812 1500
rect 1883 1444 1913 1478
rect 1961 1471 1991 1505
rect 2039 1471 2069 1505
rect 2117 1444 2147 1478
rect 2218 1466 2248 1500
rect 2362 1466 2392 1500
rect 2463 1444 2493 1478
rect 2541 1471 2571 1505
rect 2619 1471 2649 1505
rect 2697 1444 2727 1478
rect 2798 1466 2828 1500
rect 2942 1466 2972 1500
rect 3043 1444 3073 1478
rect 3121 1471 3151 1505
rect 3199 1471 3229 1505
rect 3277 1444 3307 1478
rect 3378 1466 3408 1500
rect 3522 1466 3552 1500
rect 3623 1444 3653 1478
rect 3701 1471 3731 1505
rect 3779 1471 3809 1505
rect 3857 1444 3887 1478
rect 3958 1466 3988 1500
rect 4102 1466 4132 1500
rect 4203 1444 4233 1478
rect 4281 1471 4311 1505
rect 4359 1471 4389 1505
rect 4437 1444 4467 1478
rect 4538 1466 4568 1500
rect 4682 1466 4712 1500
rect 4783 1444 4813 1478
rect 4861 1471 4891 1505
rect 4939 1471 4969 1505
rect 5017 1444 5047 1478
rect 5118 1466 5148 1500
rect 5262 1466 5292 1500
rect 5363 1444 5393 1478
rect 5441 1471 5471 1505
rect 5519 1471 5549 1505
rect 5597 1444 5627 1478
rect 5698 1466 5728 1500
rect 5842 1466 5872 1500
rect 5943 1444 5973 1478
rect 6021 1471 6051 1505
rect 6099 1471 6129 1505
rect 6177 1444 6207 1478
rect 6278 1466 6308 1500
rect 6422 1466 6452 1500
rect 6523 1444 6553 1478
rect 6601 1471 6631 1505
rect 6679 1471 6709 1505
rect 6757 1444 6787 1478
rect 6858 1466 6888 1500
rect 42 1196 72 1230
rect 143 1174 173 1208
rect 221 1201 251 1235
rect 299 1201 329 1235
rect 377 1174 407 1208
rect 478 1196 508 1230
rect 622 1196 652 1230
rect 723 1174 753 1208
rect 801 1201 831 1235
rect 879 1201 909 1235
rect 957 1174 987 1208
rect 1058 1196 1088 1230
rect 1202 1196 1232 1230
rect 1303 1174 1333 1208
rect 1381 1201 1411 1235
rect 1459 1201 1489 1235
rect 1537 1174 1567 1208
rect 1638 1196 1668 1230
rect 1782 1196 1812 1230
rect 1883 1174 1913 1208
rect 1961 1201 1991 1235
rect 2039 1201 2069 1235
rect 2117 1174 2147 1208
rect 2218 1196 2248 1230
rect 2362 1196 2392 1230
rect 2463 1174 2493 1208
rect 2541 1201 2571 1235
rect 2619 1201 2649 1235
rect 2697 1174 2727 1208
rect 2798 1196 2828 1230
rect 2942 1196 2972 1230
rect 3043 1174 3073 1208
rect 3121 1201 3151 1235
rect 3199 1201 3229 1235
rect 3277 1174 3307 1208
rect 3378 1196 3408 1230
rect 3522 1196 3552 1230
rect 3623 1174 3653 1208
rect 3701 1201 3731 1235
rect 3779 1201 3809 1235
rect 3857 1174 3887 1208
rect 3958 1196 3988 1230
rect 4102 1196 4132 1230
rect 4203 1174 4233 1208
rect 4281 1201 4311 1235
rect 4359 1201 4389 1235
rect 4437 1174 4467 1208
rect 4538 1196 4568 1230
rect 4682 1196 4712 1230
rect 4783 1174 4813 1208
rect 4861 1201 4891 1235
rect 4939 1201 4969 1235
rect 5017 1174 5047 1208
rect 5118 1196 5148 1230
rect 5262 1196 5292 1230
rect 5363 1174 5393 1208
rect 5441 1201 5471 1235
rect 5519 1201 5549 1235
rect 5597 1174 5627 1208
rect 5698 1196 5728 1230
rect 5842 1196 5872 1230
rect 5943 1174 5973 1208
rect 6021 1201 6051 1235
rect 6099 1201 6129 1235
rect 6177 1174 6207 1208
rect 6278 1196 6308 1230
rect 6422 1196 6452 1230
rect 6523 1174 6553 1208
rect 6601 1201 6631 1235
rect 6679 1201 6709 1235
rect 6757 1174 6787 1208
rect 6858 1196 6888 1230
rect 42 926 72 960
rect 143 904 173 938
rect 221 931 251 965
rect 299 931 329 965
rect 377 904 407 938
rect 478 926 508 960
rect 622 926 652 960
rect 723 904 753 938
rect 801 931 831 965
rect 879 931 909 965
rect 957 904 987 938
rect 1058 926 1088 960
rect 1202 926 1232 960
rect 1303 904 1333 938
rect 1381 931 1411 965
rect 1459 931 1489 965
rect 1537 904 1567 938
rect 1638 926 1668 960
rect 1782 926 1812 960
rect 1883 904 1913 938
rect 1961 931 1991 965
rect 2039 931 2069 965
rect 2117 904 2147 938
rect 2218 926 2248 960
rect 2362 926 2392 960
rect 2463 904 2493 938
rect 2541 931 2571 965
rect 2619 931 2649 965
rect 2697 904 2727 938
rect 2798 926 2828 960
rect 2942 926 2972 960
rect 3043 904 3073 938
rect 3121 931 3151 965
rect 3199 931 3229 965
rect 3277 904 3307 938
rect 3378 926 3408 960
rect 3522 926 3552 960
rect 3623 904 3653 938
rect 3701 931 3731 965
rect 3779 931 3809 965
rect 3857 904 3887 938
rect 3958 926 3988 960
rect 4102 926 4132 960
rect 4203 904 4233 938
rect 4281 931 4311 965
rect 4359 931 4389 965
rect 4437 904 4467 938
rect 4538 926 4568 960
rect 4682 926 4712 960
rect 4783 904 4813 938
rect 4861 931 4891 965
rect 4939 931 4969 965
rect 5017 904 5047 938
rect 5118 926 5148 960
rect 5262 926 5292 960
rect 5363 904 5393 938
rect 5441 931 5471 965
rect 5519 931 5549 965
rect 5597 904 5627 938
rect 5698 926 5728 960
rect 5842 926 5872 960
rect 5943 904 5973 938
rect 6021 931 6051 965
rect 6099 931 6129 965
rect 6177 904 6207 938
rect 6278 926 6308 960
rect 6422 926 6452 960
rect 6523 904 6553 938
rect 6601 931 6631 965
rect 6679 931 6709 965
rect 6757 904 6787 938
rect 6858 926 6888 960
rect 42 656 72 690
rect 143 634 173 668
rect 221 661 251 695
rect 299 661 329 695
rect 377 634 407 668
rect 478 656 508 690
rect 622 656 652 690
rect 723 634 753 668
rect 801 661 831 695
rect 879 661 909 695
rect 957 634 987 668
rect 1058 656 1088 690
rect 1202 656 1232 690
rect 1303 634 1333 668
rect 1381 661 1411 695
rect 1459 661 1489 695
rect 1537 634 1567 668
rect 1638 656 1668 690
rect 1782 656 1812 690
rect 1883 634 1913 668
rect 1961 661 1991 695
rect 2039 661 2069 695
rect 2117 634 2147 668
rect 2218 656 2248 690
rect 2362 656 2392 690
rect 2463 634 2493 668
rect 2541 661 2571 695
rect 2619 661 2649 695
rect 2697 634 2727 668
rect 2798 656 2828 690
rect 2942 656 2972 690
rect 3043 634 3073 668
rect 3121 661 3151 695
rect 3199 661 3229 695
rect 3277 634 3307 668
rect 3378 656 3408 690
rect 3522 656 3552 690
rect 3623 634 3653 668
rect 3701 661 3731 695
rect 3779 661 3809 695
rect 3857 634 3887 668
rect 3958 656 3988 690
rect 4102 656 4132 690
rect 4203 634 4233 668
rect 4281 661 4311 695
rect 4359 661 4389 695
rect 4437 634 4467 668
rect 4538 656 4568 690
rect 4682 656 4712 690
rect 4783 634 4813 668
rect 4861 661 4891 695
rect 4939 661 4969 695
rect 5017 634 5047 668
rect 5118 656 5148 690
rect 5262 656 5292 690
rect 5363 634 5393 668
rect 5441 661 5471 695
rect 5519 661 5549 695
rect 5597 634 5627 668
rect 5698 656 5728 690
rect 5842 656 5872 690
rect 5943 634 5973 668
rect 6021 661 6051 695
rect 6099 661 6129 695
rect 6177 634 6207 668
rect 6278 656 6308 690
rect 6422 656 6452 690
rect 6523 634 6553 668
rect 6601 661 6631 695
rect 6679 661 6709 695
rect 6757 634 6787 668
rect 6858 656 6888 690
rect 42 386 72 420
rect 143 364 173 398
rect 221 391 251 425
rect 299 391 329 425
rect 377 364 407 398
rect 478 386 508 420
rect 622 386 652 420
rect 723 364 753 398
rect 801 391 831 425
rect 879 391 909 425
rect 957 364 987 398
rect 1058 386 1088 420
rect 1202 386 1232 420
rect 1303 364 1333 398
rect 1381 391 1411 425
rect 1459 391 1489 425
rect 1537 364 1567 398
rect 1638 386 1668 420
rect 1782 386 1812 420
rect 1883 364 1913 398
rect 1961 391 1991 425
rect 2039 391 2069 425
rect 2117 364 2147 398
rect 2218 386 2248 420
rect 2362 386 2392 420
rect 2463 364 2493 398
rect 2541 391 2571 425
rect 2619 391 2649 425
rect 2697 364 2727 398
rect 2798 386 2828 420
rect 2942 386 2972 420
rect 3043 364 3073 398
rect 3121 391 3151 425
rect 3199 391 3229 425
rect 3277 364 3307 398
rect 3378 386 3408 420
rect 3522 386 3552 420
rect 3623 364 3653 398
rect 3701 391 3731 425
rect 3779 391 3809 425
rect 3857 364 3887 398
rect 3958 386 3988 420
rect 4102 386 4132 420
rect 4203 364 4233 398
rect 4281 391 4311 425
rect 4359 391 4389 425
rect 4437 364 4467 398
rect 4538 386 4568 420
rect 4682 386 4712 420
rect 4783 364 4813 398
rect 4861 391 4891 425
rect 4939 391 4969 425
rect 5017 364 5047 398
rect 5118 386 5148 420
rect 5262 386 5292 420
rect 5363 364 5393 398
rect 5441 391 5471 425
rect 5519 391 5549 425
rect 5597 364 5627 398
rect 5698 386 5728 420
rect 5842 386 5872 420
rect 5943 364 5973 398
rect 6021 391 6051 425
rect 6099 391 6129 425
rect 6177 364 6207 398
rect 6278 386 6308 420
rect 6422 386 6452 420
rect 6523 364 6553 398
rect 6601 391 6631 425
rect 6679 391 6709 425
rect 6757 364 6787 398
rect 6858 386 6888 420
rect 42 116 72 150
rect 143 94 173 128
rect 221 121 251 155
rect 299 121 329 155
rect 377 94 407 128
rect 478 116 508 150
rect 622 116 652 150
rect 723 94 753 128
rect 801 121 831 155
rect 879 121 909 155
rect 957 94 987 128
rect 1058 116 1088 150
rect 1202 116 1232 150
rect 1303 94 1333 128
rect 1381 121 1411 155
rect 1459 121 1489 155
rect 1537 94 1567 128
rect 1638 116 1668 150
rect 1782 116 1812 150
rect 1883 94 1913 128
rect 1961 121 1991 155
rect 2039 121 2069 155
rect 2117 94 2147 128
rect 2218 116 2248 150
rect 2362 116 2392 150
rect 2463 94 2493 128
rect 2541 121 2571 155
rect 2619 121 2649 155
rect 2697 94 2727 128
rect 2798 116 2828 150
rect 2942 116 2972 150
rect 3043 94 3073 128
rect 3121 121 3151 155
rect 3199 121 3229 155
rect 3277 94 3307 128
rect 3378 116 3408 150
rect 3522 116 3552 150
rect 3623 94 3653 128
rect 3701 121 3731 155
rect 3779 121 3809 155
rect 3857 94 3887 128
rect 3958 116 3988 150
rect 4102 116 4132 150
rect 4203 94 4233 128
rect 4281 121 4311 155
rect 4359 121 4389 155
rect 4437 94 4467 128
rect 4538 116 4568 150
rect 4682 116 4712 150
rect 4783 94 4813 128
rect 4861 121 4891 155
rect 4939 121 4969 155
rect 5017 94 5047 128
rect 5118 116 5148 150
rect 5262 116 5292 150
rect 5363 94 5393 128
rect 5441 121 5471 155
rect 5519 121 5549 155
rect 5597 94 5627 128
rect 5698 116 5728 150
rect 5842 116 5872 150
rect 5943 94 5973 128
rect 6021 121 6051 155
rect 6099 121 6129 155
rect 6177 94 6207 128
rect 6278 116 6308 150
rect 6422 116 6452 150
rect 6523 94 6553 128
rect 6601 121 6631 155
rect 6679 121 6709 155
rect 6757 94 6787 128
rect 6858 116 6888 150
rect 42 -154 72 -120
rect 143 -176 173 -142
rect 221 -149 251 -115
rect 299 -149 329 -115
rect 377 -176 407 -142
rect 478 -154 508 -120
rect 622 -154 652 -120
rect 723 -176 753 -142
rect 801 -149 831 -115
rect 879 -149 909 -115
rect 957 -176 987 -142
rect 1058 -154 1088 -120
rect 1202 -154 1232 -120
rect 1303 -176 1333 -142
rect 1381 -149 1411 -115
rect 1459 -149 1489 -115
rect 1537 -176 1567 -142
rect 1638 -154 1668 -120
rect 1782 -154 1812 -120
rect 1883 -176 1913 -142
rect 1961 -149 1991 -115
rect 2039 -149 2069 -115
rect 2117 -176 2147 -142
rect 2218 -154 2248 -120
rect 2362 -154 2392 -120
rect 2463 -176 2493 -142
rect 2541 -149 2571 -115
rect 2619 -149 2649 -115
rect 2697 -176 2727 -142
rect 2798 -154 2828 -120
rect 2942 -154 2972 -120
rect 3043 -176 3073 -142
rect 3121 -149 3151 -115
rect 3199 -149 3229 -115
rect 3277 -176 3307 -142
rect 3378 -154 3408 -120
rect 3522 -154 3552 -120
rect 3623 -176 3653 -142
rect 3701 -149 3731 -115
rect 3779 -149 3809 -115
rect 3857 -176 3887 -142
rect 3958 -154 3988 -120
rect 4102 -154 4132 -120
rect 4203 -176 4233 -142
rect 4281 -149 4311 -115
rect 4359 -149 4389 -115
rect 4437 -176 4467 -142
rect 4538 -154 4568 -120
rect 4682 -154 4712 -120
rect 4783 -176 4813 -142
rect 4861 -149 4891 -115
rect 4939 -149 4969 -115
rect 5017 -176 5047 -142
rect 5118 -154 5148 -120
rect 5262 -154 5292 -120
rect 5363 -176 5393 -142
rect 5441 -149 5471 -115
rect 5519 -149 5549 -115
rect 5597 -176 5627 -142
rect 5698 -154 5728 -120
rect 5842 -154 5872 -120
rect 5943 -176 5973 -142
rect 6021 -149 6051 -115
rect 6099 -149 6129 -115
rect 6177 -176 6207 -142
rect 6278 -154 6308 -120
rect 6422 -154 6452 -120
rect 6523 -176 6553 -142
rect 6601 -149 6631 -115
rect 6679 -149 6709 -115
rect 6757 -176 6787 -142
rect 6858 -154 6888 -120
rect 42 -424 72 -390
rect 143 -446 173 -412
rect 221 -419 251 -385
rect 299 -419 329 -385
rect 377 -446 407 -412
rect 478 -424 508 -390
rect 622 -424 652 -390
rect 723 -446 753 -412
rect 801 -419 831 -385
rect 879 -419 909 -385
rect 957 -446 987 -412
rect 1058 -424 1088 -390
rect 1202 -424 1232 -390
rect 1303 -446 1333 -412
rect 1381 -419 1411 -385
rect 1459 -419 1489 -385
rect 1537 -446 1567 -412
rect 1638 -424 1668 -390
rect 1782 -424 1812 -390
rect 1883 -446 1913 -412
rect 1961 -419 1991 -385
rect 2039 -419 2069 -385
rect 2117 -446 2147 -412
rect 2218 -424 2248 -390
rect 2362 -424 2392 -390
rect 2463 -446 2493 -412
rect 2541 -419 2571 -385
rect 2619 -419 2649 -385
rect 2697 -446 2727 -412
rect 2798 -424 2828 -390
rect 2942 -424 2972 -390
rect 3043 -446 3073 -412
rect 3121 -419 3151 -385
rect 3199 -419 3229 -385
rect 3277 -446 3307 -412
rect 3378 -424 3408 -390
rect 3522 -424 3552 -390
rect 3623 -446 3653 -412
rect 3701 -419 3731 -385
rect 3779 -419 3809 -385
rect 3857 -446 3887 -412
rect 3958 -424 3988 -390
rect 4102 -424 4132 -390
rect 4203 -446 4233 -412
rect 4281 -419 4311 -385
rect 4359 -419 4389 -385
rect 4437 -446 4467 -412
rect 4538 -424 4568 -390
rect 4682 -424 4712 -390
rect 4783 -446 4813 -412
rect 4861 -419 4891 -385
rect 4939 -419 4969 -385
rect 5017 -446 5047 -412
rect 5118 -424 5148 -390
rect 5262 -424 5292 -390
rect 5363 -446 5393 -412
rect 5441 -419 5471 -385
rect 5519 -419 5549 -385
rect 5597 -446 5627 -412
rect 5698 -424 5728 -390
rect 5842 -424 5872 -390
rect 5943 -446 5973 -412
rect 6021 -419 6051 -385
rect 6099 -419 6129 -385
rect 6177 -446 6207 -412
rect 6278 -424 6308 -390
rect 6422 -424 6452 -390
rect 6523 -446 6553 -412
rect 6601 -419 6631 -385
rect 6679 -419 6709 -385
rect 6757 -446 6787 -412
rect 6858 -424 6888 -390
rect 42 -694 72 -660
rect 143 -716 173 -682
rect 221 -689 251 -655
rect 299 -689 329 -655
rect 377 -716 407 -682
rect 478 -694 508 -660
rect 622 -694 652 -660
rect 723 -716 753 -682
rect 801 -689 831 -655
rect 879 -689 909 -655
rect 957 -716 987 -682
rect 1058 -694 1088 -660
rect 1202 -694 1232 -660
rect 1303 -716 1333 -682
rect 1381 -689 1411 -655
rect 1459 -689 1489 -655
rect 1537 -716 1567 -682
rect 1638 -694 1668 -660
rect 1782 -694 1812 -660
rect 1883 -716 1913 -682
rect 1961 -689 1991 -655
rect 2039 -689 2069 -655
rect 2117 -716 2147 -682
rect 2218 -694 2248 -660
rect 2362 -694 2392 -660
rect 2463 -716 2493 -682
rect 2541 -689 2571 -655
rect 2619 -689 2649 -655
rect 2697 -716 2727 -682
rect 2798 -694 2828 -660
rect 2942 -694 2972 -660
rect 3043 -716 3073 -682
rect 3121 -689 3151 -655
rect 3199 -689 3229 -655
rect 3277 -716 3307 -682
rect 3378 -694 3408 -660
rect 3522 -694 3552 -660
rect 3623 -716 3653 -682
rect 3701 -689 3731 -655
rect 3779 -689 3809 -655
rect 3857 -716 3887 -682
rect 3958 -694 3988 -660
rect 4102 -694 4132 -660
rect 4203 -716 4233 -682
rect 4281 -689 4311 -655
rect 4359 -689 4389 -655
rect 4437 -716 4467 -682
rect 4538 -694 4568 -660
rect 4682 -694 4712 -660
rect 4783 -716 4813 -682
rect 4861 -689 4891 -655
rect 4939 -689 4969 -655
rect 5017 -716 5047 -682
rect 5118 -694 5148 -660
rect 5262 -694 5292 -660
rect 5363 -716 5393 -682
rect 5441 -689 5471 -655
rect 5519 -689 5549 -655
rect 5597 -716 5627 -682
rect 5698 -694 5728 -660
rect 5842 -694 5872 -660
rect 5943 -716 5973 -682
rect 6021 -689 6051 -655
rect 6099 -689 6129 -655
rect 6177 -716 6207 -682
rect 6278 -694 6308 -660
rect 6422 -694 6452 -660
rect 6523 -716 6553 -682
rect 6601 -689 6631 -655
rect 6679 -689 6709 -655
rect 6757 -716 6787 -682
rect 6858 -694 6888 -660
rect 42 -964 72 -930
rect 143 -986 173 -952
rect 221 -959 251 -925
rect 299 -959 329 -925
rect 377 -986 407 -952
rect 478 -964 508 -930
rect 622 -964 652 -930
rect 723 -986 753 -952
rect 801 -959 831 -925
rect 879 -959 909 -925
rect 957 -986 987 -952
rect 1058 -964 1088 -930
rect 1202 -964 1232 -930
rect 1303 -986 1333 -952
rect 1381 -959 1411 -925
rect 1459 -959 1489 -925
rect 1537 -986 1567 -952
rect 1638 -964 1668 -930
rect 1782 -964 1812 -930
rect 1883 -986 1913 -952
rect 1961 -959 1991 -925
rect 2039 -959 2069 -925
rect 2117 -986 2147 -952
rect 2218 -964 2248 -930
rect 2362 -964 2392 -930
rect 2463 -986 2493 -952
rect 2541 -959 2571 -925
rect 2619 -959 2649 -925
rect 2697 -986 2727 -952
rect 2798 -964 2828 -930
rect 2942 -964 2972 -930
rect 3043 -986 3073 -952
rect 3121 -959 3151 -925
rect 3199 -959 3229 -925
rect 3277 -986 3307 -952
rect 3378 -964 3408 -930
rect 3522 -964 3552 -930
rect 3623 -986 3653 -952
rect 3701 -959 3731 -925
rect 3779 -959 3809 -925
rect 3857 -986 3887 -952
rect 3958 -964 3988 -930
rect 4102 -964 4132 -930
rect 4203 -986 4233 -952
rect 4281 -959 4311 -925
rect 4359 -959 4389 -925
rect 4437 -986 4467 -952
rect 4538 -964 4568 -930
rect 4682 -964 4712 -930
rect 4783 -986 4813 -952
rect 4861 -959 4891 -925
rect 4939 -959 4969 -925
rect 5017 -986 5047 -952
rect 5118 -964 5148 -930
rect 5262 -964 5292 -930
rect 5363 -986 5393 -952
rect 5441 -959 5471 -925
rect 5519 -959 5549 -925
rect 5597 -986 5627 -952
rect 5698 -964 5728 -930
rect 5842 -964 5872 -930
rect 5943 -986 5973 -952
rect 6021 -959 6051 -925
rect 6099 -959 6129 -925
rect 6177 -986 6207 -952
rect 6278 -964 6308 -930
rect 6422 -964 6452 -930
rect 6523 -986 6553 -952
rect 6601 -959 6631 -925
rect 6679 -959 6709 -925
rect 6757 -986 6787 -952
rect 6858 -964 6888 -930
rect 42 -1234 72 -1200
rect 143 -1256 173 -1222
rect 221 -1229 251 -1195
rect 299 -1229 329 -1195
rect 377 -1256 407 -1222
rect 478 -1234 508 -1200
rect 622 -1234 652 -1200
rect 723 -1256 753 -1222
rect 801 -1229 831 -1195
rect 879 -1229 909 -1195
rect 957 -1256 987 -1222
rect 1058 -1234 1088 -1200
rect 1202 -1234 1232 -1200
rect 1303 -1256 1333 -1222
rect 1381 -1229 1411 -1195
rect 1459 -1229 1489 -1195
rect 1537 -1256 1567 -1222
rect 1638 -1234 1668 -1200
rect 1782 -1234 1812 -1200
rect 1883 -1256 1913 -1222
rect 1961 -1229 1991 -1195
rect 2039 -1229 2069 -1195
rect 2117 -1256 2147 -1222
rect 2218 -1234 2248 -1200
rect 2362 -1234 2392 -1200
rect 2463 -1256 2493 -1222
rect 2541 -1229 2571 -1195
rect 2619 -1229 2649 -1195
rect 2697 -1256 2727 -1222
rect 2798 -1234 2828 -1200
rect 2942 -1234 2972 -1200
rect 3043 -1256 3073 -1222
rect 3121 -1229 3151 -1195
rect 3199 -1229 3229 -1195
rect 3277 -1256 3307 -1222
rect 3378 -1234 3408 -1200
rect 3522 -1234 3552 -1200
rect 3623 -1256 3653 -1222
rect 3701 -1229 3731 -1195
rect 3779 -1229 3809 -1195
rect 3857 -1256 3887 -1222
rect 3958 -1234 3988 -1200
rect 4102 -1234 4132 -1200
rect 4203 -1256 4233 -1222
rect 4281 -1229 4311 -1195
rect 4359 -1229 4389 -1195
rect 4437 -1256 4467 -1222
rect 4538 -1234 4568 -1200
rect 4682 -1234 4712 -1200
rect 4783 -1256 4813 -1222
rect 4861 -1229 4891 -1195
rect 4939 -1229 4969 -1195
rect 5017 -1256 5047 -1222
rect 5118 -1234 5148 -1200
rect 5262 -1234 5292 -1200
rect 5363 -1256 5393 -1222
rect 5441 -1229 5471 -1195
rect 5519 -1229 5549 -1195
rect 5597 -1256 5627 -1222
rect 5698 -1234 5728 -1200
rect 5842 -1234 5872 -1200
rect 5943 -1256 5973 -1222
rect 6021 -1229 6051 -1195
rect 6099 -1229 6129 -1195
rect 6177 -1256 6207 -1222
rect 6278 -1234 6308 -1200
rect 6422 -1234 6452 -1200
rect 6523 -1256 6553 -1222
rect 6601 -1229 6631 -1195
rect 6679 -1229 6709 -1195
rect 6757 -1256 6787 -1222
rect 6858 -1234 6888 -1200
rect 42 -1504 72 -1470
rect 143 -1526 173 -1492
rect 221 -1499 251 -1465
rect 299 -1499 329 -1465
rect 377 -1526 407 -1492
rect 478 -1504 508 -1470
rect 622 -1504 652 -1470
rect 723 -1526 753 -1492
rect 801 -1499 831 -1465
rect 879 -1499 909 -1465
rect 957 -1526 987 -1492
rect 1058 -1504 1088 -1470
rect 1202 -1504 1232 -1470
rect 1303 -1526 1333 -1492
rect 1381 -1499 1411 -1465
rect 1459 -1499 1489 -1465
rect 1537 -1526 1567 -1492
rect 1638 -1504 1668 -1470
rect 1782 -1504 1812 -1470
rect 1883 -1526 1913 -1492
rect 1961 -1499 1991 -1465
rect 2039 -1499 2069 -1465
rect 2117 -1526 2147 -1492
rect 2218 -1504 2248 -1470
rect 2362 -1504 2392 -1470
rect 2463 -1526 2493 -1492
rect 2541 -1499 2571 -1465
rect 2619 -1499 2649 -1465
rect 2697 -1526 2727 -1492
rect 2798 -1504 2828 -1470
rect 2942 -1504 2972 -1470
rect 3043 -1526 3073 -1492
rect 3121 -1499 3151 -1465
rect 3199 -1499 3229 -1465
rect 3277 -1526 3307 -1492
rect 3378 -1504 3408 -1470
rect 3522 -1504 3552 -1470
rect 3623 -1526 3653 -1492
rect 3701 -1499 3731 -1465
rect 3779 -1499 3809 -1465
rect 3857 -1526 3887 -1492
rect 3958 -1504 3988 -1470
rect 4102 -1504 4132 -1470
rect 4203 -1526 4233 -1492
rect 4281 -1499 4311 -1465
rect 4359 -1499 4389 -1465
rect 4437 -1526 4467 -1492
rect 4538 -1504 4568 -1470
rect 4682 -1504 4712 -1470
rect 4783 -1526 4813 -1492
rect 4861 -1499 4891 -1465
rect 4939 -1499 4969 -1465
rect 5017 -1526 5047 -1492
rect 5118 -1504 5148 -1470
rect 5262 -1504 5292 -1470
rect 5363 -1526 5393 -1492
rect 5441 -1499 5471 -1465
rect 5519 -1499 5549 -1465
rect 5597 -1526 5627 -1492
rect 5698 -1504 5728 -1470
rect 5842 -1504 5872 -1470
rect 5943 -1526 5973 -1492
rect 6021 -1499 6051 -1465
rect 6099 -1499 6129 -1465
rect 6177 -1526 6207 -1492
rect 6278 -1504 6308 -1470
rect 6422 -1504 6452 -1470
rect 6523 -1526 6553 -1492
rect 6601 -1499 6631 -1465
rect 6679 -1499 6709 -1465
rect 6757 -1526 6787 -1492
rect 6858 -1504 6888 -1470
rect 42 -1774 72 -1740
rect 143 -1796 173 -1762
rect 221 -1769 251 -1735
rect 299 -1769 329 -1735
rect 377 -1796 407 -1762
rect 478 -1774 508 -1740
rect 622 -1774 652 -1740
rect 723 -1796 753 -1762
rect 801 -1769 831 -1735
rect 879 -1769 909 -1735
rect 957 -1796 987 -1762
rect 1058 -1774 1088 -1740
rect 1202 -1774 1232 -1740
rect 1303 -1796 1333 -1762
rect 1381 -1769 1411 -1735
rect 1459 -1769 1489 -1735
rect 1537 -1796 1567 -1762
rect 1638 -1774 1668 -1740
rect 1782 -1774 1812 -1740
rect 1883 -1796 1913 -1762
rect 1961 -1769 1991 -1735
rect 2039 -1769 2069 -1735
rect 2117 -1796 2147 -1762
rect 2218 -1774 2248 -1740
rect 2362 -1774 2392 -1740
rect 2463 -1796 2493 -1762
rect 2541 -1769 2571 -1735
rect 2619 -1769 2649 -1735
rect 2697 -1796 2727 -1762
rect 2798 -1774 2828 -1740
rect 2942 -1774 2972 -1740
rect 3043 -1796 3073 -1762
rect 3121 -1769 3151 -1735
rect 3199 -1769 3229 -1735
rect 3277 -1796 3307 -1762
rect 3378 -1774 3408 -1740
rect 3522 -1774 3552 -1740
rect 3623 -1796 3653 -1762
rect 3701 -1769 3731 -1735
rect 3779 -1769 3809 -1735
rect 3857 -1796 3887 -1762
rect 3958 -1774 3988 -1740
rect 4102 -1774 4132 -1740
rect 4203 -1796 4233 -1762
rect 4281 -1769 4311 -1735
rect 4359 -1769 4389 -1735
rect 4437 -1796 4467 -1762
rect 4538 -1774 4568 -1740
rect 4682 -1774 4712 -1740
rect 4783 -1796 4813 -1762
rect 4861 -1769 4891 -1735
rect 4939 -1769 4969 -1735
rect 5017 -1796 5047 -1762
rect 5118 -1774 5148 -1740
rect 5262 -1774 5292 -1740
rect 5363 -1796 5393 -1762
rect 5441 -1769 5471 -1735
rect 5519 -1769 5549 -1735
rect 5597 -1796 5627 -1762
rect 5698 -1774 5728 -1740
rect 5842 -1774 5872 -1740
rect 5943 -1796 5973 -1762
rect 6021 -1769 6051 -1735
rect 6099 -1769 6129 -1735
rect 6177 -1796 6207 -1762
rect 6278 -1774 6308 -1740
rect 6422 -1774 6452 -1740
rect 6523 -1796 6553 -1762
rect 6601 -1769 6631 -1735
rect 6679 -1769 6709 -1735
rect 6757 -1796 6787 -1762
rect 6858 -1774 6888 -1740
rect 42 -2044 72 -2010
rect 143 -2066 173 -2032
rect 221 -2039 251 -2005
rect 299 -2039 329 -2005
rect 377 -2066 407 -2032
rect 478 -2044 508 -2010
rect 622 -2044 652 -2010
rect 723 -2066 753 -2032
rect 801 -2039 831 -2005
rect 879 -2039 909 -2005
rect 957 -2066 987 -2032
rect 1058 -2044 1088 -2010
rect 1202 -2044 1232 -2010
rect 1303 -2066 1333 -2032
rect 1381 -2039 1411 -2005
rect 1459 -2039 1489 -2005
rect 1537 -2066 1567 -2032
rect 1638 -2044 1668 -2010
rect 1782 -2044 1812 -2010
rect 1883 -2066 1913 -2032
rect 1961 -2039 1991 -2005
rect 2039 -2039 2069 -2005
rect 2117 -2066 2147 -2032
rect 2218 -2044 2248 -2010
rect 2362 -2044 2392 -2010
rect 2463 -2066 2493 -2032
rect 2541 -2039 2571 -2005
rect 2619 -2039 2649 -2005
rect 2697 -2066 2727 -2032
rect 2798 -2044 2828 -2010
rect 2942 -2044 2972 -2010
rect 3043 -2066 3073 -2032
rect 3121 -2039 3151 -2005
rect 3199 -2039 3229 -2005
rect 3277 -2066 3307 -2032
rect 3378 -2044 3408 -2010
rect 3522 -2044 3552 -2010
rect 3623 -2066 3653 -2032
rect 3701 -2039 3731 -2005
rect 3779 -2039 3809 -2005
rect 3857 -2066 3887 -2032
rect 3958 -2044 3988 -2010
rect 4102 -2044 4132 -2010
rect 4203 -2066 4233 -2032
rect 4281 -2039 4311 -2005
rect 4359 -2039 4389 -2005
rect 4437 -2066 4467 -2032
rect 4538 -2044 4568 -2010
rect 4682 -2044 4712 -2010
rect 4783 -2066 4813 -2032
rect 4861 -2039 4891 -2005
rect 4939 -2039 4969 -2005
rect 5017 -2066 5047 -2032
rect 5118 -2044 5148 -2010
rect 5262 -2044 5292 -2010
rect 5363 -2066 5393 -2032
rect 5441 -2039 5471 -2005
rect 5519 -2039 5549 -2005
rect 5597 -2066 5627 -2032
rect 5698 -2044 5728 -2010
rect 5842 -2044 5872 -2010
rect 5943 -2066 5973 -2032
rect 6021 -2039 6051 -2005
rect 6099 -2039 6129 -2005
rect 6177 -2066 6207 -2032
rect 6278 -2044 6308 -2010
rect 6422 -2044 6452 -2010
rect 6523 -2066 6553 -2032
rect 6601 -2039 6631 -2005
rect 6679 -2039 6709 -2005
rect 6757 -2066 6787 -2032
rect 6858 -2044 6888 -2010
<< corelocali >>
rect -1 1984 14 2174
tri 79 2138 101 2160 se
rect 101 2153 116 2174
tri 101 2138 116 2153 nw
rect 435 2153 450 2174
tri 73 2132 79 2138 se
rect 79 2132 88 2138
rect 73 2116 88 2132
tri 88 2125 101 2138 nw
rect 242 2130 259 2144
rect 291 2130 308 2144
tri 435 2138 450 2153 ne
tri 450 2138 472 2160 sw
rect 73 2080 88 2088
rect 154 2116 214 2130
rect 169 2106 214 2116
rect 169 2088 197 2106
tri 73 2065 88 2080 ne
tri 88 2065 110 2087 sw
rect 154 2078 197 2088
rect 212 2102 214 2106
rect 336 2116 396 2130
tri 450 2125 463 2138 ne
rect 463 2132 472 2138
tri 472 2132 478 2138 sw
rect 336 2106 381 2116
rect 212 2078 286 2102
rect 154 2074 286 2078
tri 286 2074 314 2102 sw
rect 336 2092 338 2106
tri 336 2090 338 2092 ne
rect 350 2088 381 2106
rect 350 2078 396 2088
rect 463 2117 478 2132
tri 88 2053 100 2065 ne
rect 100 2060 110 2065
tri 110 2060 115 2065 sw
rect -1 1714 14 1942
rect 100 1904 115 2060
rect 154 2018 182 2074
tri 274 2056 292 2074 ne
rect 292 2054 314 2074
tri 314 2054 334 2074 sw
tri 350 2060 368 2078 ne
rect 173 1984 182 2018
rect 216 2045 258 2046
rect 216 2011 221 2045
rect 251 2011 258 2045
rect 216 2002 258 2011
rect 292 2045 334 2054
rect 292 2011 299 2045
rect 329 2011 334 2045
rect 292 2006 334 2011
rect 368 2018 396 2078
tri 441 2065 463 2087 se
rect 463 2080 478 2088
tri 463 2065 478 2080 nw
tri 435 2059 441 2065 se
rect 441 2059 450 2065
rect 154 1974 182 1984
tri 182 1974 206 1998 sw
rect 154 1942 196 1974
tri 213 1966 214 1967 sw
rect 213 1942 214 1966
tri 216 1965 253 2002 ne
rect 253 1974 258 2002
tri 258 1974 284 2000 sw
rect 368 1984 377 2018
rect 368 1974 396 1984
rect 253 1965 337 1974
tri 253 1946 272 1965 ne
rect 272 1946 337 1965
rect 154 1920 214 1942
rect 336 1942 337 1946
rect 354 1942 396 1974
rect 336 1920 396 1942
rect 242 1904 259 1918
rect 291 1904 308 1918
tri 79 1868 101 1890 se
rect 101 1883 116 1904
tri 101 1868 116 1883 nw
rect 435 1883 450 2059
tri 450 2052 463 2065 nw
rect 536 1984 551 2174
tri 73 1862 79 1868 se
rect 79 1862 88 1868
rect 73 1846 88 1862
tri 88 1855 101 1868 nw
rect 242 1860 259 1874
rect 291 1860 308 1874
tri 435 1868 450 1883 ne
tri 450 1868 472 1890 sw
rect 73 1810 88 1818
rect 154 1846 214 1860
rect 169 1836 214 1846
rect 169 1818 197 1836
tri 73 1795 88 1810 ne
tri 88 1795 110 1817 sw
rect 154 1808 197 1818
rect 212 1832 214 1836
rect 336 1846 396 1860
tri 450 1855 463 1868 ne
rect 463 1862 472 1868
tri 472 1862 478 1868 sw
rect 336 1836 381 1846
rect 212 1808 286 1832
rect 154 1804 286 1808
tri 286 1804 314 1832 sw
rect 336 1822 338 1836
tri 336 1820 338 1822 ne
rect 350 1818 381 1836
rect 350 1808 396 1818
rect 463 1847 478 1862
tri 88 1783 100 1795 ne
rect 100 1790 110 1795
tri 110 1790 115 1795 sw
rect -1 1444 14 1672
rect 100 1634 115 1790
rect 154 1748 182 1804
tri 274 1786 292 1804 ne
rect 292 1784 314 1804
tri 314 1784 334 1804 sw
tri 350 1790 368 1808 ne
rect 173 1714 182 1748
rect 216 1775 258 1776
rect 216 1741 221 1775
rect 251 1741 258 1775
rect 216 1732 258 1741
rect 292 1775 334 1784
rect 292 1741 299 1775
rect 329 1741 334 1775
rect 292 1736 334 1741
rect 368 1748 396 1808
tri 441 1795 463 1817 se
rect 463 1810 478 1818
tri 463 1795 478 1810 nw
tri 435 1789 441 1795 se
rect 441 1789 450 1795
rect 154 1704 182 1714
tri 182 1704 206 1728 sw
rect 154 1672 196 1704
tri 213 1696 214 1697 sw
rect 213 1672 214 1696
tri 216 1695 253 1732 ne
rect 253 1704 258 1732
tri 258 1704 284 1730 sw
rect 368 1714 377 1748
rect 368 1704 396 1714
rect 253 1695 337 1704
tri 253 1676 272 1695 ne
rect 272 1676 337 1695
rect 154 1650 214 1672
rect 336 1672 337 1676
rect 354 1672 396 1704
rect 336 1650 396 1672
rect 242 1634 259 1648
rect 291 1634 308 1648
tri 79 1598 101 1620 se
rect 101 1613 116 1634
tri 101 1598 116 1613 nw
rect 435 1613 450 1789
tri 450 1782 463 1795 nw
rect 536 1714 551 1942
tri 73 1592 79 1598 se
rect 79 1592 88 1598
rect 73 1576 88 1592
tri 88 1585 101 1598 nw
rect 242 1590 259 1604
rect 291 1590 308 1604
tri 435 1598 450 1613 ne
tri 450 1598 472 1620 sw
rect 73 1540 88 1548
rect 154 1576 214 1590
rect 169 1566 214 1576
rect 169 1548 197 1566
tri 73 1525 88 1540 ne
tri 88 1525 110 1547 sw
rect 154 1538 197 1548
rect 212 1562 214 1566
rect 336 1576 396 1590
tri 450 1585 463 1598 ne
rect 463 1592 472 1598
tri 472 1592 478 1598 sw
rect 336 1566 381 1576
rect 212 1538 286 1562
rect 154 1534 286 1538
tri 286 1534 314 1562 sw
rect 336 1552 338 1566
tri 336 1550 338 1552 ne
rect 350 1548 381 1566
rect 350 1538 396 1548
rect 463 1577 478 1592
tri 88 1513 100 1525 ne
rect 100 1520 110 1525
tri 110 1520 115 1525 sw
rect -1 1174 14 1402
rect 100 1364 115 1520
rect 154 1478 182 1534
tri 274 1516 292 1534 ne
rect 292 1514 314 1534
tri 314 1514 334 1534 sw
tri 350 1520 368 1538 ne
rect 173 1444 182 1478
rect 216 1505 258 1506
rect 216 1471 221 1505
rect 251 1471 258 1505
rect 216 1462 258 1471
rect 292 1505 334 1514
rect 292 1471 299 1505
rect 329 1471 334 1505
rect 292 1466 334 1471
rect 368 1478 396 1538
tri 441 1525 463 1547 se
rect 463 1540 478 1548
tri 463 1525 478 1540 nw
tri 435 1519 441 1525 se
rect 441 1519 450 1525
rect 154 1434 182 1444
tri 182 1434 206 1458 sw
rect 154 1402 196 1434
tri 213 1426 214 1427 sw
rect 213 1402 214 1426
tri 216 1425 253 1462 ne
rect 253 1434 258 1462
tri 258 1434 284 1460 sw
rect 368 1444 377 1478
rect 368 1434 396 1444
rect 253 1425 337 1434
tri 253 1406 272 1425 ne
rect 272 1406 337 1425
rect 154 1380 214 1402
rect 336 1402 337 1406
rect 354 1402 396 1434
rect 336 1380 396 1402
rect 242 1364 259 1378
rect 291 1364 308 1378
tri 79 1328 101 1350 se
rect 101 1343 116 1364
tri 101 1328 116 1343 nw
rect 435 1343 450 1519
tri 450 1512 463 1525 nw
rect 536 1444 551 1672
tri 73 1322 79 1328 se
rect 79 1322 88 1328
rect 73 1306 88 1322
tri 88 1315 101 1328 nw
rect 242 1320 259 1334
rect 291 1320 308 1334
tri 435 1328 450 1343 ne
tri 450 1328 472 1350 sw
rect 73 1270 88 1278
rect 154 1306 214 1320
rect 169 1296 214 1306
rect 169 1278 197 1296
tri 73 1255 88 1270 ne
tri 88 1255 110 1277 sw
rect 154 1268 197 1278
rect 212 1292 214 1296
rect 336 1306 396 1320
tri 450 1315 463 1328 ne
rect 463 1322 472 1328
tri 472 1322 478 1328 sw
rect 336 1296 381 1306
rect 212 1268 286 1292
rect 154 1264 286 1268
tri 286 1264 314 1292 sw
rect 336 1282 338 1296
tri 336 1280 338 1282 ne
rect 350 1278 381 1296
rect 350 1268 396 1278
rect 463 1307 478 1322
tri 88 1243 100 1255 ne
rect 100 1250 110 1255
tri 110 1250 115 1255 sw
rect -1 904 14 1132
rect 100 1094 115 1250
rect 154 1208 182 1264
tri 274 1246 292 1264 ne
rect 292 1244 314 1264
tri 314 1244 334 1264 sw
tri 350 1250 368 1268 ne
rect 173 1174 182 1208
rect 216 1235 258 1236
rect 216 1201 221 1235
rect 251 1201 258 1235
rect 216 1192 258 1201
rect 292 1235 334 1244
rect 292 1201 299 1235
rect 329 1201 334 1235
rect 292 1196 334 1201
rect 368 1208 396 1268
tri 441 1255 463 1277 se
rect 463 1270 478 1278
tri 463 1255 478 1270 nw
tri 435 1249 441 1255 se
rect 441 1249 450 1255
rect 154 1164 182 1174
tri 182 1164 206 1188 sw
rect 154 1132 196 1164
tri 213 1156 214 1157 sw
rect 213 1132 214 1156
tri 216 1155 253 1192 ne
rect 253 1164 258 1192
tri 258 1164 284 1190 sw
rect 368 1174 377 1208
rect 368 1164 396 1174
rect 253 1155 337 1164
tri 253 1136 272 1155 ne
rect 272 1136 337 1155
rect 154 1110 214 1132
rect 336 1132 337 1136
rect 354 1132 396 1164
rect 336 1110 396 1132
rect 242 1094 259 1108
rect 291 1094 308 1108
tri 79 1058 101 1080 se
rect 101 1073 116 1094
tri 101 1058 116 1073 nw
rect 435 1073 450 1249
tri 450 1242 463 1255 nw
rect 536 1174 551 1402
tri 73 1052 79 1058 se
rect 79 1052 88 1058
rect 73 1036 88 1052
tri 88 1045 101 1058 nw
rect 242 1050 259 1064
rect 291 1050 308 1064
tri 435 1058 450 1073 ne
tri 450 1058 472 1080 sw
rect 73 1000 88 1008
rect 154 1036 214 1050
rect 169 1026 214 1036
rect 169 1008 197 1026
tri 73 985 88 1000 ne
tri 88 985 110 1007 sw
rect 154 998 197 1008
rect 212 1022 214 1026
rect 336 1036 396 1050
tri 450 1045 463 1058 ne
rect 463 1052 472 1058
tri 472 1052 478 1058 sw
rect 336 1026 381 1036
rect 212 998 286 1022
rect 154 994 286 998
tri 286 994 314 1022 sw
rect 336 1012 338 1026
tri 336 1010 338 1012 ne
rect 350 1008 381 1026
rect 350 998 396 1008
rect 463 1037 478 1052
tri 88 973 100 985 ne
rect 100 980 110 985
tri 110 980 115 985 sw
rect -1 634 14 862
rect 100 824 115 980
rect 154 938 182 994
tri 274 976 292 994 ne
rect 292 974 314 994
tri 314 974 334 994 sw
tri 350 980 368 998 ne
rect 173 904 182 938
rect 216 965 258 966
rect 216 931 221 965
rect 251 931 258 965
rect 216 922 258 931
rect 292 965 334 974
rect 292 931 299 965
rect 329 931 334 965
rect 292 926 334 931
rect 368 938 396 998
tri 441 985 463 1007 se
rect 463 1000 478 1008
tri 463 985 478 1000 nw
tri 435 979 441 985 se
rect 441 979 450 985
rect 154 894 182 904
tri 182 894 206 918 sw
rect 154 862 196 894
tri 213 886 214 887 sw
rect 213 862 214 886
tri 216 885 253 922 ne
rect 253 894 258 922
tri 258 894 284 920 sw
rect 368 904 377 938
rect 368 894 396 904
rect 253 885 337 894
tri 253 866 272 885 ne
rect 272 866 337 885
rect 154 840 214 862
rect 336 862 337 866
rect 354 862 396 894
rect 336 840 396 862
rect 242 824 259 838
rect 291 824 308 838
tri 79 788 101 810 se
rect 101 803 116 824
tri 101 788 116 803 nw
rect 435 803 450 979
tri 450 972 463 985 nw
rect 536 904 551 1132
tri 73 782 79 788 se
rect 79 782 88 788
rect 73 766 88 782
tri 88 775 101 788 nw
rect 242 780 259 794
rect 291 780 308 794
tri 435 788 450 803 ne
tri 450 788 472 810 sw
rect 73 730 88 738
rect 154 766 214 780
rect 169 756 214 766
rect 169 738 197 756
tri 73 715 88 730 ne
tri 88 715 110 737 sw
rect 154 728 197 738
rect 212 752 214 756
rect 336 766 396 780
tri 450 775 463 788 ne
rect 463 782 472 788
tri 472 782 478 788 sw
rect 336 756 381 766
rect 212 728 286 752
rect 154 724 286 728
tri 286 724 314 752 sw
rect 336 742 338 756
tri 336 740 338 742 ne
rect 350 738 381 756
rect 350 728 396 738
rect 463 767 478 782
tri 88 703 100 715 ne
rect 100 710 110 715
tri 110 710 115 715 sw
rect -1 364 14 592
rect 100 554 115 710
rect 154 668 182 724
tri 274 706 292 724 ne
rect 292 704 314 724
tri 314 704 334 724 sw
tri 350 710 368 728 ne
rect 173 634 182 668
rect 216 695 258 696
rect 216 661 221 695
rect 251 661 258 695
rect 216 652 258 661
rect 292 695 334 704
rect 292 661 299 695
rect 329 661 334 695
rect 292 656 334 661
rect 368 668 396 728
tri 441 715 463 737 se
rect 463 730 478 738
tri 463 715 478 730 nw
tri 435 709 441 715 se
rect 441 709 450 715
rect 154 624 182 634
tri 182 624 206 648 sw
rect 154 592 196 624
tri 213 616 214 617 sw
rect 213 592 214 616
tri 216 615 253 652 ne
rect 253 624 258 652
tri 258 624 284 650 sw
rect 368 634 377 668
rect 368 624 396 634
rect 253 615 337 624
tri 253 596 272 615 ne
rect 272 596 337 615
rect 154 570 214 592
rect 336 592 337 596
rect 354 592 396 624
rect 336 570 396 592
rect 242 554 259 568
rect 291 554 308 568
tri 79 518 101 540 se
rect 101 533 116 554
tri 101 518 116 533 nw
rect 435 533 450 709
tri 450 702 463 715 nw
rect 536 634 551 862
tri 73 512 79 518 se
rect 79 512 88 518
rect 73 496 88 512
tri 88 505 101 518 nw
rect 242 510 259 524
rect 291 510 308 524
tri 435 518 450 533 ne
tri 450 518 472 540 sw
rect 73 460 88 468
rect 154 496 214 510
rect 169 486 214 496
rect 169 468 197 486
tri 73 445 88 460 ne
tri 88 445 110 467 sw
rect 154 458 197 468
rect 212 482 214 486
rect 336 496 396 510
tri 450 505 463 518 ne
rect 463 512 472 518
tri 472 512 478 518 sw
rect 336 486 381 496
rect 212 458 286 482
rect 154 454 286 458
tri 286 454 314 482 sw
rect 336 472 338 486
tri 336 470 338 472 ne
rect 350 468 381 486
rect 350 458 396 468
rect 463 497 478 512
tri 88 433 100 445 ne
rect 100 440 110 445
tri 110 440 115 445 sw
rect -1 94 14 322
rect 100 284 115 440
rect 154 398 182 454
tri 274 436 292 454 ne
rect 292 434 314 454
tri 314 434 334 454 sw
tri 350 440 368 458 ne
rect 173 364 182 398
rect 216 425 258 426
rect 216 391 221 425
rect 251 391 258 425
rect 216 382 258 391
rect 292 425 334 434
rect 292 391 299 425
rect 329 391 334 425
rect 292 386 334 391
rect 368 398 396 458
tri 441 445 463 467 se
rect 463 460 478 468
tri 463 445 478 460 nw
tri 435 439 441 445 se
rect 441 439 450 445
rect 154 354 182 364
tri 182 354 206 378 sw
rect 154 322 196 354
tri 213 346 214 347 sw
rect 213 322 214 346
tri 216 345 253 382 ne
rect 253 354 258 382
tri 258 354 284 380 sw
rect 368 364 377 398
rect 368 354 396 364
rect 253 345 337 354
tri 253 326 272 345 ne
rect 272 326 337 345
rect 154 300 214 322
rect 336 322 337 326
rect 354 322 396 354
rect 336 300 396 322
rect 242 284 259 298
rect 291 284 308 298
tri 79 248 101 270 se
rect 101 263 116 284
tri 101 248 116 263 nw
rect 435 263 450 439
tri 450 432 463 445 nw
rect 536 364 551 592
tri 73 242 79 248 se
rect 79 242 88 248
rect 73 226 88 242
tri 88 235 101 248 nw
rect 242 240 259 254
rect 291 240 308 254
tri 435 248 450 263 ne
tri 450 248 472 270 sw
rect 73 190 88 198
rect 154 226 214 240
rect 169 216 214 226
rect 169 198 197 216
tri 73 175 88 190 ne
tri 88 175 110 197 sw
rect 154 188 197 198
rect 212 212 214 216
rect 336 226 396 240
tri 450 235 463 248 ne
rect 463 242 472 248
tri 472 242 478 248 sw
rect 336 216 381 226
rect 212 188 286 212
rect 154 184 286 188
tri 286 184 314 212 sw
rect 336 202 338 216
tri 336 200 338 202 ne
rect 350 198 381 216
rect 350 188 396 198
rect 463 227 478 242
tri 88 163 100 175 ne
rect 100 170 110 175
tri 110 170 115 175 sw
rect -1 -176 14 52
rect 100 14 115 170
rect 154 128 182 184
tri 274 166 292 184 ne
rect 292 164 314 184
tri 314 164 334 184 sw
tri 350 170 368 188 ne
rect 173 94 182 128
rect 216 155 258 156
rect 216 121 221 155
rect 251 121 258 155
rect 216 112 258 121
rect 292 155 334 164
rect 292 121 299 155
rect 329 121 334 155
rect 292 116 334 121
rect 368 128 396 188
tri 441 175 463 197 se
rect 463 190 478 198
tri 463 175 478 190 nw
tri 435 169 441 175 se
rect 441 169 450 175
rect 154 84 182 94
tri 182 84 206 108 sw
rect 154 52 196 84
tri 213 76 214 77 sw
rect 213 52 214 76
tri 216 75 253 112 ne
rect 253 84 258 112
tri 258 84 284 110 sw
rect 368 94 377 128
rect 368 84 396 94
rect 253 75 337 84
tri 253 56 272 75 ne
rect 272 56 337 75
rect 154 30 214 52
rect 336 52 337 56
rect 354 52 396 84
rect 336 30 396 52
rect 242 14 259 28
rect 291 14 308 28
tri 79 -22 101 0 se
rect 101 -7 116 14
tri 101 -22 116 -7 nw
rect 435 -7 450 169
tri 450 162 463 175 nw
rect 536 94 551 322
tri 73 -28 79 -22 se
rect 79 -28 88 -22
rect 73 -44 88 -28
tri 88 -35 101 -22 nw
rect 242 -30 259 -16
rect 291 -30 308 -16
tri 435 -22 450 -7 ne
tri 450 -22 472 0 sw
rect 73 -80 88 -72
rect 154 -44 214 -30
rect 169 -54 214 -44
rect 169 -72 197 -54
tri 73 -95 88 -80 ne
tri 88 -95 110 -73 sw
rect 154 -82 197 -72
rect 212 -58 214 -54
rect 336 -44 396 -30
tri 450 -35 463 -22 ne
rect 463 -28 472 -22
tri 472 -28 478 -22 sw
rect 336 -54 381 -44
rect 212 -82 286 -58
rect 154 -86 286 -82
tri 286 -86 314 -58 sw
rect 336 -68 338 -54
tri 336 -70 338 -68 ne
rect 350 -72 381 -54
rect 350 -82 396 -72
rect 463 -43 478 -28
tri 88 -107 100 -95 ne
rect 100 -100 110 -95
tri 110 -100 115 -95 sw
rect -1 -446 14 -218
rect 100 -256 115 -100
rect 154 -142 182 -86
tri 274 -104 292 -86 ne
rect 292 -106 314 -86
tri 314 -106 334 -86 sw
tri 350 -100 368 -82 ne
rect 173 -176 182 -142
rect 216 -115 258 -114
rect 216 -149 221 -115
rect 251 -149 258 -115
rect 216 -158 258 -149
rect 292 -115 334 -106
rect 292 -149 299 -115
rect 329 -149 334 -115
rect 292 -154 334 -149
rect 368 -142 396 -82
tri 441 -95 463 -73 se
rect 463 -80 478 -72
tri 463 -95 478 -80 nw
tri 435 -101 441 -95 se
rect 441 -101 450 -95
rect 154 -186 182 -176
tri 182 -186 206 -162 sw
rect 154 -218 196 -186
tri 213 -194 214 -193 sw
rect 213 -218 214 -194
tri 216 -195 253 -158 ne
rect 253 -186 258 -158
tri 258 -186 284 -160 sw
rect 368 -176 377 -142
rect 368 -186 396 -176
rect 253 -195 337 -186
tri 253 -214 272 -195 ne
rect 272 -214 337 -195
rect 154 -240 214 -218
rect 336 -218 337 -214
rect 354 -218 396 -186
rect 336 -240 396 -218
rect 242 -256 259 -242
rect 291 -256 308 -242
tri 79 -292 101 -270 se
rect 101 -277 116 -256
tri 101 -292 116 -277 nw
rect 435 -277 450 -101
tri 450 -108 463 -95 nw
rect 536 -176 551 52
tri 73 -298 79 -292 se
rect 79 -298 88 -292
rect 73 -314 88 -298
tri 88 -305 101 -292 nw
rect 242 -300 259 -286
rect 291 -300 308 -286
tri 435 -292 450 -277 ne
tri 450 -292 472 -270 sw
rect 73 -350 88 -342
rect 154 -314 214 -300
rect 169 -324 214 -314
rect 169 -342 197 -324
tri 73 -365 88 -350 ne
tri 88 -365 110 -343 sw
rect 154 -352 197 -342
rect 212 -328 214 -324
rect 336 -314 396 -300
tri 450 -305 463 -292 ne
rect 463 -298 472 -292
tri 472 -298 478 -292 sw
rect 336 -324 381 -314
rect 212 -352 286 -328
rect 154 -356 286 -352
tri 286 -356 314 -328 sw
rect 336 -338 338 -324
tri 336 -340 338 -338 ne
rect 350 -342 381 -324
rect 350 -352 396 -342
rect 463 -313 478 -298
tri 88 -377 100 -365 ne
rect 100 -370 110 -365
tri 110 -370 115 -365 sw
rect -1 -716 14 -488
rect 100 -526 115 -370
rect 154 -412 182 -356
tri 274 -374 292 -356 ne
rect 292 -376 314 -356
tri 314 -376 334 -356 sw
tri 350 -370 368 -352 ne
rect 173 -446 182 -412
rect 216 -385 258 -384
rect 216 -419 221 -385
rect 251 -419 258 -385
rect 216 -428 258 -419
rect 292 -385 334 -376
rect 292 -419 299 -385
rect 329 -419 334 -385
rect 292 -424 334 -419
rect 368 -412 396 -352
tri 441 -365 463 -343 se
rect 463 -350 478 -342
tri 463 -365 478 -350 nw
tri 435 -371 441 -365 se
rect 441 -371 450 -365
rect 154 -456 182 -446
tri 182 -456 206 -432 sw
rect 154 -488 196 -456
tri 213 -464 214 -463 sw
rect 213 -488 214 -464
tri 216 -465 253 -428 ne
rect 253 -456 258 -428
tri 258 -456 284 -430 sw
rect 368 -446 377 -412
rect 368 -456 396 -446
rect 253 -465 337 -456
tri 253 -484 272 -465 ne
rect 272 -484 337 -465
rect 154 -510 214 -488
rect 336 -488 337 -484
rect 354 -488 396 -456
rect 336 -510 396 -488
rect 242 -526 259 -512
rect 291 -526 308 -512
tri 79 -562 101 -540 se
rect 101 -547 116 -526
tri 101 -562 116 -547 nw
rect 435 -547 450 -371
tri 450 -378 463 -365 nw
rect 536 -446 551 -218
tri 73 -568 79 -562 se
rect 79 -568 88 -562
rect 73 -584 88 -568
tri 88 -575 101 -562 nw
rect 242 -570 259 -556
rect 291 -570 308 -556
tri 435 -562 450 -547 ne
tri 450 -562 472 -540 sw
rect 73 -620 88 -612
rect 154 -584 214 -570
rect 169 -594 214 -584
rect 169 -612 197 -594
tri 73 -635 88 -620 ne
tri 88 -635 110 -613 sw
rect 154 -622 197 -612
rect 212 -598 214 -594
rect 336 -584 396 -570
tri 450 -575 463 -562 ne
rect 463 -568 472 -562
tri 472 -568 478 -562 sw
rect 336 -594 381 -584
rect 212 -622 286 -598
rect 154 -626 286 -622
tri 286 -626 314 -598 sw
rect 336 -608 338 -594
tri 336 -610 338 -608 ne
rect 350 -612 381 -594
rect 350 -622 396 -612
rect 463 -583 478 -568
tri 88 -647 100 -635 ne
rect 100 -640 110 -635
tri 110 -640 115 -635 sw
rect -1 -986 14 -758
rect 100 -796 115 -640
rect 154 -682 182 -626
tri 274 -644 292 -626 ne
rect 292 -646 314 -626
tri 314 -646 334 -626 sw
tri 350 -640 368 -622 ne
rect 173 -716 182 -682
rect 216 -655 258 -654
rect 216 -689 221 -655
rect 251 -689 258 -655
rect 216 -698 258 -689
rect 292 -655 334 -646
rect 292 -689 299 -655
rect 329 -689 334 -655
rect 292 -694 334 -689
rect 368 -682 396 -622
tri 441 -635 463 -613 se
rect 463 -620 478 -612
tri 463 -635 478 -620 nw
tri 435 -641 441 -635 se
rect 441 -641 450 -635
rect 154 -726 182 -716
tri 182 -726 206 -702 sw
rect 154 -758 196 -726
tri 213 -734 214 -733 sw
rect 213 -758 214 -734
tri 216 -735 253 -698 ne
rect 253 -726 258 -698
tri 258 -726 284 -700 sw
rect 368 -716 377 -682
rect 368 -726 396 -716
rect 253 -735 337 -726
tri 253 -754 272 -735 ne
rect 272 -754 337 -735
rect 154 -780 214 -758
rect 336 -758 337 -754
rect 354 -758 396 -726
rect 336 -780 396 -758
rect 242 -796 259 -782
rect 291 -796 308 -782
tri 79 -832 101 -810 se
rect 101 -817 116 -796
tri 101 -832 116 -817 nw
rect 435 -817 450 -641
tri 450 -648 463 -635 nw
rect 536 -716 551 -488
tri 73 -838 79 -832 se
rect 79 -838 88 -832
rect 73 -854 88 -838
tri 88 -845 101 -832 nw
rect 242 -840 259 -826
rect 291 -840 308 -826
tri 435 -832 450 -817 ne
tri 450 -832 472 -810 sw
rect 73 -890 88 -882
rect 154 -854 214 -840
rect 169 -864 214 -854
rect 169 -882 197 -864
tri 73 -905 88 -890 ne
tri 88 -905 110 -883 sw
rect 154 -892 197 -882
rect 212 -868 214 -864
rect 336 -854 396 -840
tri 450 -845 463 -832 ne
rect 463 -838 472 -832
tri 472 -838 478 -832 sw
rect 336 -864 381 -854
rect 212 -892 286 -868
rect 154 -896 286 -892
tri 286 -896 314 -868 sw
rect 336 -878 338 -864
tri 336 -880 338 -878 ne
rect 350 -882 381 -864
rect 350 -892 396 -882
rect 463 -853 478 -838
tri 88 -917 100 -905 ne
rect 100 -910 110 -905
tri 110 -910 115 -905 sw
rect -1 -1256 14 -1028
rect 100 -1066 115 -910
rect 154 -952 182 -896
tri 274 -914 292 -896 ne
rect 292 -916 314 -896
tri 314 -916 334 -896 sw
tri 350 -910 368 -892 ne
rect 173 -986 182 -952
rect 216 -925 258 -924
rect 216 -959 221 -925
rect 251 -959 258 -925
rect 216 -968 258 -959
rect 292 -925 334 -916
rect 292 -959 299 -925
rect 329 -959 334 -925
rect 292 -964 334 -959
rect 368 -952 396 -892
tri 441 -905 463 -883 se
rect 463 -890 478 -882
tri 463 -905 478 -890 nw
tri 435 -911 441 -905 se
rect 441 -911 450 -905
rect 154 -996 182 -986
tri 182 -996 206 -972 sw
rect 154 -1028 196 -996
tri 213 -1004 214 -1003 sw
rect 213 -1028 214 -1004
tri 216 -1005 253 -968 ne
rect 253 -996 258 -968
tri 258 -996 284 -970 sw
rect 368 -986 377 -952
rect 368 -996 396 -986
rect 253 -1005 337 -996
tri 253 -1024 272 -1005 ne
rect 272 -1024 337 -1005
rect 154 -1050 214 -1028
rect 336 -1028 337 -1024
rect 354 -1028 396 -996
rect 336 -1050 396 -1028
rect 242 -1066 259 -1052
rect 291 -1066 308 -1052
tri 79 -1102 101 -1080 se
rect 101 -1087 116 -1066
tri 101 -1102 116 -1087 nw
rect 435 -1087 450 -911
tri 450 -918 463 -905 nw
rect 536 -986 551 -758
tri 73 -1108 79 -1102 se
rect 79 -1108 88 -1102
rect 73 -1124 88 -1108
tri 88 -1115 101 -1102 nw
rect 242 -1110 259 -1096
rect 291 -1110 308 -1096
tri 435 -1102 450 -1087 ne
tri 450 -1102 472 -1080 sw
rect 73 -1160 88 -1152
rect 154 -1124 214 -1110
rect 169 -1134 214 -1124
rect 169 -1152 197 -1134
tri 73 -1175 88 -1160 ne
tri 88 -1175 110 -1153 sw
rect 154 -1162 197 -1152
rect 212 -1138 214 -1134
rect 336 -1124 396 -1110
tri 450 -1115 463 -1102 ne
rect 463 -1108 472 -1102
tri 472 -1108 478 -1102 sw
rect 336 -1134 381 -1124
rect 212 -1162 286 -1138
rect 154 -1166 286 -1162
tri 286 -1166 314 -1138 sw
rect 336 -1148 338 -1134
tri 336 -1150 338 -1148 ne
rect 350 -1152 381 -1134
rect 350 -1162 396 -1152
rect 463 -1123 478 -1108
tri 88 -1187 100 -1175 ne
rect 100 -1180 110 -1175
tri 110 -1180 115 -1175 sw
rect -1 -1526 14 -1298
rect 100 -1336 115 -1180
rect 154 -1222 182 -1166
tri 274 -1184 292 -1166 ne
rect 292 -1186 314 -1166
tri 314 -1186 334 -1166 sw
tri 350 -1180 368 -1162 ne
rect 173 -1256 182 -1222
rect 216 -1195 258 -1194
rect 216 -1229 221 -1195
rect 251 -1229 258 -1195
rect 216 -1238 258 -1229
rect 292 -1195 334 -1186
rect 292 -1229 299 -1195
rect 329 -1229 334 -1195
rect 292 -1234 334 -1229
rect 368 -1222 396 -1162
tri 441 -1175 463 -1153 se
rect 463 -1160 478 -1152
tri 463 -1175 478 -1160 nw
tri 435 -1181 441 -1175 se
rect 441 -1181 450 -1175
rect 154 -1266 182 -1256
tri 182 -1266 206 -1242 sw
rect 154 -1298 196 -1266
tri 213 -1274 214 -1273 sw
rect 213 -1298 214 -1274
tri 216 -1275 253 -1238 ne
rect 253 -1266 258 -1238
tri 258 -1266 284 -1240 sw
rect 368 -1256 377 -1222
rect 368 -1266 396 -1256
rect 253 -1275 337 -1266
tri 253 -1294 272 -1275 ne
rect 272 -1294 337 -1275
rect 154 -1320 214 -1298
rect 336 -1298 337 -1294
rect 354 -1298 396 -1266
rect 336 -1320 396 -1298
rect 242 -1336 259 -1322
rect 291 -1336 308 -1322
tri 79 -1372 101 -1350 se
rect 101 -1357 116 -1336
tri 101 -1372 116 -1357 nw
rect 435 -1357 450 -1181
tri 450 -1188 463 -1175 nw
rect 536 -1256 551 -1028
tri 73 -1378 79 -1372 se
rect 79 -1378 88 -1372
rect 73 -1394 88 -1378
tri 88 -1385 101 -1372 nw
rect 242 -1380 259 -1366
rect 291 -1380 308 -1366
tri 435 -1372 450 -1357 ne
tri 450 -1372 472 -1350 sw
rect 73 -1430 88 -1422
rect 154 -1394 214 -1380
rect 169 -1404 214 -1394
rect 169 -1422 197 -1404
tri 73 -1445 88 -1430 ne
tri 88 -1445 110 -1423 sw
rect 154 -1432 197 -1422
rect 212 -1408 214 -1404
rect 336 -1394 396 -1380
tri 450 -1385 463 -1372 ne
rect 463 -1378 472 -1372
tri 472 -1378 478 -1372 sw
rect 336 -1404 381 -1394
rect 212 -1432 286 -1408
rect 154 -1436 286 -1432
tri 286 -1436 314 -1408 sw
rect 336 -1418 338 -1404
tri 336 -1420 338 -1418 ne
rect 350 -1422 381 -1404
rect 350 -1432 396 -1422
rect 463 -1393 478 -1378
tri 88 -1457 100 -1445 ne
rect 100 -1450 110 -1445
tri 110 -1450 115 -1445 sw
rect -1 -1796 14 -1568
rect 100 -1606 115 -1450
rect 154 -1492 182 -1436
tri 274 -1454 292 -1436 ne
rect 292 -1456 314 -1436
tri 314 -1456 334 -1436 sw
tri 350 -1450 368 -1432 ne
rect 173 -1526 182 -1492
rect 216 -1465 258 -1464
rect 216 -1499 221 -1465
rect 251 -1499 258 -1465
rect 216 -1508 258 -1499
rect 292 -1465 334 -1456
rect 292 -1499 299 -1465
rect 329 -1499 334 -1465
rect 292 -1504 334 -1499
rect 368 -1492 396 -1432
tri 441 -1445 463 -1423 se
rect 463 -1430 478 -1422
tri 463 -1445 478 -1430 nw
tri 435 -1451 441 -1445 se
rect 441 -1451 450 -1445
rect 154 -1536 182 -1526
tri 182 -1536 206 -1512 sw
rect 154 -1568 196 -1536
tri 213 -1544 214 -1543 sw
rect 213 -1568 214 -1544
tri 216 -1545 253 -1508 ne
rect 253 -1536 258 -1508
tri 258 -1536 284 -1510 sw
rect 368 -1526 377 -1492
rect 368 -1536 396 -1526
rect 253 -1545 337 -1536
tri 253 -1564 272 -1545 ne
rect 272 -1564 337 -1545
rect 154 -1590 214 -1568
rect 336 -1568 337 -1564
rect 354 -1568 396 -1536
rect 336 -1590 396 -1568
rect 242 -1606 259 -1592
rect 291 -1606 308 -1592
tri 79 -1642 101 -1620 se
rect 101 -1627 116 -1606
tri 101 -1642 116 -1627 nw
rect 435 -1627 450 -1451
tri 450 -1458 463 -1445 nw
rect 536 -1526 551 -1298
tri 73 -1648 79 -1642 se
rect 79 -1648 88 -1642
rect 73 -1664 88 -1648
tri 88 -1655 101 -1642 nw
rect 242 -1650 259 -1636
rect 291 -1650 308 -1636
tri 435 -1642 450 -1627 ne
tri 450 -1642 472 -1620 sw
rect 73 -1700 88 -1692
rect 154 -1664 214 -1650
rect 169 -1674 214 -1664
rect 169 -1692 197 -1674
tri 73 -1715 88 -1700 ne
tri 88 -1715 110 -1693 sw
rect 154 -1702 197 -1692
rect 212 -1678 214 -1674
rect 336 -1664 396 -1650
tri 450 -1655 463 -1642 ne
rect 463 -1648 472 -1642
tri 472 -1648 478 -1642 sw
rect 336 -1674 381 -1664
rect 212 -1702 286 -1678
rect 154 -1706 286 -1702
tri 286 -1706 314 -1678 sw
rect 336 -1688 338 -1674
tri 336 -1690 338 -1688 ne
rect 350 -1692 381 -1674
rect 350 -1702 396 -1692
rect 463 -1663 478 -1648
tri 88 -1727 100 -1715 ne
rect 100 -1720 110 -1715
tri 110 -1720 115 -1715 sw
rect -1 -2066 14 -1838
rect 100 -1876 115 -1720
rect 154 -1762 182 -1706
tri 274 -1724 292 -1706 ne
rect 292 -1726 314 -1706
tri 314 -1726 334 -1706 sw
tri 350 -1720 368 -1702 ne
rect 173 -1796 182 -1762
rect 216 -1735 258 -1734
rect 216 -1769 221 -1735
rect 251 -1769 258 -1735
rect 216 -1778 258 -1769
rect 292 -1735 334 -1726
rect 292 -1769 299 -1735
rect 329 -1769 334 -1735
rect 292 -1774 334 -1769
rect 368 -1762 396 -1702
tri 441 -1715 463 -1693 se
rect 463 -1700 478 -1692
tri 463 -1715 478 -1700 nw
tri 435 -1721 441 -1715 se
rect 441 -1721 450 -1715
rect 154 -1806 182 -1796
tri 182 -1806 206 -1782 sw
rect 154 -1838 196 -1806
tri 213 -1814 214 -1813 sw
rect 213 -1838 214 -1814
tri 216 -1815 253 -1778 ne
rect 253 -1806 258 -1778
tri 258 -1806 284 -1780 sw
rect 368 -1796 377 -1762
rect 368 -1806 396 -1796
rect 253 -1815 337 -1806
tri 253 -1834 272 -1815 ne
rect 272 -1834 337 -1815
rect 154 -1860 214 -1838
rect 336 -1838 337 -1834
rect 354 -1838 396 -1806
rect 336 -1860 396 -1838
rect 242 -1876 259 -1862
rect 291 -1876 308 -1862
tri 79 -1912 101 -1890 se
rect 101 -1897 116 -1876
tri 101 -1912 116 -1897 nw
rect 435 -1897 450 -1721
tri 450 -1728 463 -1715 nw
rect 536 -1796 551 -1568
tri 73 -1918 79 -1912 se
rect 79 -1918 88 -1912
rect 73 -1934 88 -1918
tri 88 -1925 101 -1912 nw
rect 242 -1920 259 -1906
rect 291 -1920 308 -1906
tri 435 -1912 450 -1897 ne
tri 450 -1912 472 -1890 sw
rect 73 -1970 88 -1962
rect 154 -1934 214 -1920
rect 169 -1944 214 -1934
rect 169 -1962 197 -1944
tri 73 -1985 88 -1970 ne
tri 88 -1985 110 -1963 sw
rect 154 -1972 197 -1962
rect 212 -1948 214 -1944
rect 336 -1934 396 -1920
tri 450 -1925 463 -1912 ne
rect 463 -1918 472 -1912
tri 472 -1918 478 -1912 sw
rect 336 -1944 381 -1934
rect 212 -1972 286 -1948
rect 154 -1976 286 -1972
tri 286 -1976 314 -1948 sw
rect 336 -1958 338 -1944
tri 336 -1960 338 -1958 ne
rect 350 -1962 381 -1944
rect 350 -1972 396 -1962
rect 463 -1933 478 -1918
tri 88 -1997 100 -1985 ne
rect 100 -1990 110 -1985
tri 110 -1990 115 -1985 sw
rect -1 -2146 14 -2108
rect 100 -2146 115 -1990
rect 154 -2032 182 -1976
tri 274 -1994 292 -1976 ne
rect 292 -1996 314 -1976
tri 314 -1996 334 -1976 sw
tri 350 -1990 368 -1972 ne
rect 173 -2066 182 -2032
rect 216 -2005 258 -2004
rect 216 -2039 221 -2005
rect 251 -2039 258 -2005
rect 216 -2048 258 -2039
rect 292 -2005 334 -1996
rect 292 -2039 299 -2005
rect 329 -2039 334 -2005
rect 292 -2044 334 -2039
rect 368 -2032 396 -1972
tri 441 -1985 463 -1963 se
rect 463 -1970 478 -1962
tri 463 -1985 478 -1970 nw
tri 435 -1991 441 -1985 se
rect 441 -1991 450 -1985
rect 154 -2076 182 -2066
tri 182 -2076 206 -2052 sw
rect 154 -2108 196 -2076
tri 213 -2084 214 -2083 sw
rect 213 -2108 214 -2084
tri 216 -2085 253 -2048 ne
rect 253 -2076 258 -2048
tri 258 -2076 284 -2050 sw
rect 368 -2066 377 -2032
rect 368 -2076 396 -2066
rect 253 -2085 337 -2076
tri 253 -2104 272 -2085 ne
rect 272 -2104 337 -2085
rect 154 -2130 214 -2108
rect 336 -2108 337 -2104
rect 354 -2108 396 -2076
rect 336 -2130 396 -2108
rect 242 -2146 259 -2132
rect 291 -2146 308 -2132
rect 435 -2146 450 -1991
tri 450 -1998 463 -1985 nw
rect 536 -2066 551 -1838
rect 536 -2146 551 -2108
rect 579 1984 594 2174
tri 659 2138 681 2160 se
rect 681 2153 696 2174
tri 681 2138 696 2153 nw
rect 1015 2153 1030 2174
tri 653 2132 659 2138 se
rect 659 2132 668 2138
rect 653 2116 668 2132
tri 668 2125 681 2138 nw
rect 822 2130 839 2144
rect 871 2130 888 2144
tri 1015 2138 1030 2153 ne
tri 1030 2138 1052 2160 sw
rect 653 2080 668 2088
rect 734 2116 794 2130
rect 749 2106 794 2116
rect 749 2088 777 2106
tri 653 2065 668 2080 ne
tri 668 2065 690 2087 sw
rect 734 2078 777 2088
rect 792 2102 794 2106
rect 916 2116 976 2130
tri 1030 2125 1043 2138 ne
rect 1043 2132 1052 2138
tri 1052 2132 1058 2138 sw
rect 916 2106 961 2116
rect 792 2078 866 2102
rect 734 2074 866 2078
tri 866 2074 894 2102 sw
rect 916 2092 918 2106
tri 916 2090 918 2092 ne
rect 930 2088 961 2106
rect 930 2078 976 2088
rect 1043 2117 1058 2132
tri 668 2053 680 2065 ne
rect 680 2060 690 2065
tri 690 2060 695 2065 sw
rect 579 1714 594 1942
rect 680 1904 695 2060
rect 734 2018 762 2074
tri 854 2056 872 2074 ne
rect 872 2054 894 2074
tri 894 2054 914 2074 sw
tri 930 2060 948 2078 ne
rect 753 1984 762 2018
rect 796 2045 838 2046
rect 796 2011 801 2045
rect 831 2011 838 2045
rect 796 2002 838 2011
rect 872 2045 914 2054
rect 872 2011 879 2045
rect 909 2011 914 2045
rect 872 2006 914 2011
rect 948 2018 976 2078
tri 1021 2065 1043 2087 se
rect 1043 2080 1058 2088
tri 1043 2065 1058 2080 nw
tri 1015 2059 1021 2065 se
rect 1021 2059 1030 2065
rect 734 1974 762 1984
tri 762 1974 786 1998 sw
rect 734 1942 776 1974
tri 793 1966 794 1967 sw
rect 793 1942 794 1966
tri 796 1965 833 2002 ne
rect 833 1974 838 2002
tri 838 1974 864 2000 sw
rect 948 1984 957 2018
rect 948 1974 976 1984
rect 833 1965 917 1974
tri 833 1946 852 1965 ne
rect 852 1946 917 1965
rect 734 1920 794 1942
rect 916 1942 917 1946
rect 934 1942 976 1974
rect 916 1920 976 1942
rect 822 1904 839 1918
rect 871 1904 888 1918
tri 659 1868 681 1890 se
rect 681 1883 696 1904
tri 681 1868 696 1883 nw
rect 1015 1883 1030 2059
tri 1030 2052 1043 2065 nw
rect 1116 1984 1131 2174
tri 653 1862 659 1868 se
rect 659 1862 668 1868
rect 653 1846 668 1862
tri 668 1855 681 1868 nw
rect 822 1860 839 1874
rect 871 1860 888 1874
tri 1015 1868 1030 1883 ne
tri 1030 1868 1052 1890 sw
rect 653 1810 668 1818
rect 734 1846 794 1860
rect 749 1836 794 1846
rect 749 1818 777 1836
tri 653 1795 668 1810 ne
tri 668 1795 690 1817 sw
rect 734 1808 777 1818
rect 792 1832 794 1836
rect 916 1846 976 1860
tri 1030 1855 1043 1868 ne
rect 1043 1862 1052 1868
tri 1052 1862 1058 1868 sw
rect 916 1836 961 1846
rect 792 1808 866 1832
rect 734 1804 866 1808
tri 866 1804 894 1832 sw
rect 916 1822 918 1836
tri 916 1820 918 1822 ne
rect 930 1818 961 1836
rect 930 1808 976 1818
rect 1043 1847 1058 1862
tri 668 1783 680 1795 ne
rect 680 1790 690 1795
tri 690 1790 695 1795 sw
rect 579 1444 594 1672
rect 680 1634 695 1790
rect 734 1748 762 1804
tri 854 1786 872 1804 ne
rect 872 1784 894 1804
tri 894 1784 914 1804 sw
tri 930 1790 948 1808 ne
rect 753 1714 762 1748
rect 796 1775 838 1776
rect 796 1741 801 1775
rect 831 1741 838 1775
rect 796 1732 838 1741
rect 872 1775 914 1784
rect 872 1741 879 1775
rect 909 1741 914 1775
rect 872 1736 914 1741
rect 948 1748 976 1808
tri 1021 1795 1043 1817 se
rect 1043 1810 1058 1818
tri 1043 1795 1058 1810 nw
tri 1015 1789 1021 1795 se
rect 1021 1789 1030 1795
rect 734 1704 762 1714
tri 762 1704 786 1728 sw
rect 734 1672 776 1704
tri 793 1696 794 1697 sw
rect 793 1672 794 1696
tri 796 1695 833 1732 ne
rect 833 1704 838 1732
tri 838 1704 864 1730 sw
rect 948 1714 957 1748
rect 948 1704 976 1714
rect 833 1695 917 1704
tri 833 1676 852 1695 ne
rect 852 1676 917 1695
rect 734 1650 794 1672
rect 916 1672 917 1676
rect 934 1672 976 1704
rect 916 1650 976 1672
rect 822 1634 839 1648
rect 871 1634 888 1648
tri 659 1598 681 1620 se
rect 681 1613 696 1634
tri 681 1598 696 1613 nw
rect 1015 1613 1030 1789
tri 1030 1782 1043 1795 nw
rect 1116 1714 1131 1942
tri 653 1592 659 1598 se
rect 659 1592 668 1598
rect 653 1576 668 1592
tri 668 1585 681 1598 nw
rect 822 1590 839 1604
rect 871 1590 888 1604
tri 1015 1598 1030 1613 ne
tri 1030 1598 1052 1620 sw
rect 653 1540 668 1548
rect 734 1576 794 1590
rect 749 1566 794 1576
rect 749 1548 777 1566
tri 653 1525 668 1540 ne
tri 668 1525 690 1547 sw
rect 734 1538 777 1548
rect 792 1562 794 1566
rect 916 1576 976 1590
tri 1030 1585 1043 1598 ne
rect 1043 1592 1052 1598
tri 1052 1592 1058 1598 sw
rect 916 1566 961 1576
rect 792 1538 866 1562
rect 734 1534 866 1538
tri 866 1534 894 1562 sw
rect 916 1552 918 1566
tri 916 1550 918 1552 ne
rect 930 1548 961 1566
rect 930 1538 976 1548
rect 1043 1577 1058 1592
tri 668 1513 680 1525 ne
rect 680 1520 690 1525
tri 690 1520 695 1525 sw
rect 579 1174 594 1402
rect 680 1364 695 1520
rect 734 1478 762 1534
tri 854 1516 872 1534 ne
rect 872 1514 894 1534
tri 894 1514 914 1534 sw
tri 930 1520 948 1538 ne
rect 753 1444 762 1478
rect 796 1505 838 1506
rect 796 1471 801 1505
rect 831 1471 838 1505
rect 796 1462 838 1471
rect 872 1505 914 1514
rect 872 1471 879 1505
rect 909 1471 914 1505
rect 872 1466 914 1471
rect 948 1478 976 1538
tri 1021 1525 1043 1547 se
rect 1043 1540 1058 1548
tri 1043 1525 1058 1540 nw
tri 1015 1519 1021 1525 se
rect 1021 1519 1030 1525
rect 734 1434 762 1444
tri 762 1434 786 1458 sw
rect 734 1402 776 1434
tri 793 1426 794 1427 sw
rect 793 1402 794 1426
tri 796 1425 833 1462 ne
rect 833 1434 838 1462
tri 838 1434 864 1460 sw
rect 948 1444 957 1478
rect 948 1434 976 1444
rect 833 1425 917 1434
tri 833 1406 852 1425 ne
rect 852 1406 917 1425
rect 734 1380 794 1402
rect 916 1402 917 1406
rect 934 1402 976 1434
rect 916 1380 976 1402
rect 822 1364 839 1378
rect 871 1364 888 1378
tri 659 1328 681 1350 se
rect 681 1343 696 1364
tri 681 1328 696 1343 nw
rect 1015 1343 1030 1519
tri 1030 1512 1043 1525 nw
rect 1116 1444 1131 1672
tri 653 1322 659 1328 se
rect 659 1322 668 1328
rect 653 1306 668 1322
tri 668 1315 681 1328 nw
rect 822 1320 839 1334
rect 871 1320 888 1334
tri 1015 1328 1030 1343 ne
tri 1030 1328 1052 1350 sw
rect 653 1270 668 1278
rect 734 1306 794 1320
rect 749 1296 794 1306
rect 749 1278 777 1296
tri 653 1255 668 1270 ne
tri 668 1255 690 1277 sw
rect 734 1268 777 1278
rect 792 1292 794 1296
rect 916 1306 976 1320
tri 1030 1315 1043 1328 ne
rect 1043 1322 1052 1328
tri 1052 1322 1058 1328 sw
rect 916 1296 961 1306
rect 792 1268 866 1292
rect 734 1264 866 1268
tri 866 1264 894 1292 sw
rect 916 1282 918 1296
tri 916 1280 918 1282 ne
rect 930 1278 961 1296
rect 930 1268 976 1278
rect 1043 1307 1058 1322
tri 668 1243 680 1255 ne
rect 680 1250 690 1255
tri 690 1250 695 1255 sw
rect 579 904 594 1132
rect 680 1094 695 1250
rect 734 1208 762 1264
tri 854 1246 872 1264 ne
rect 872 1244 894 1264
tri 894 1244 914 1264 sw
tri 930 1250 948 1268 ne
rect 753 1174 762 1208
rect 796 1235 838 1236
rect 796 1201 801 1235
rect 831 1201 838 1235
rect 796 1192 838 1201
rect 872 1235 914 1244
rect 872 1201 879 1235
rect 909 1201 914 1235
rect 872 1196 914 1201
rect 948 1208 976 1268
tri 1021 1255 1043 1277 se
rect 1043 1270 1058 1278
tri 1043 1255 1058 1270 nw
tri 1015 1249 1021 1255 se
rect 1021 1249 1030 1255
rect 734 1164 762 1174
tri 762 1164 786 1188 sw
rect 734 1132 776 1164
tri 793 1156 794 1157 sw
rect 793 1132 794 1156
tri 796 1155 833 1192 ne
rect 833 1164 838 1192
tri 838 1164 864 1190 sw
rect 948 1174 957 1208
rect 948 1164 976 1174
rect 833 1155 917 1164
tri 833 1136 852 1155 ne
rect 852 1136 917 1155
rect 734 1110 794 1132
rect 916 1132 917 1136
rect 934 1132 976 1164
rect 916 1110 976 1132
rect 822 1094 839 1108
rect 871 1094 888 1108
tri 659 1058 681 1080 se
rect 681 1073 696 1094
tri 681 1058 696 1073 nw
rect 1015 1073 1030 1249
tri 1030 1242 1043 1255 nw
rect 1116 1174 1131 1402
tri 653 1052 659 1058 se
rect 659 1052 668 1058
rect 653 1036 668 1052
tri 668 1045 681 1058 nw
rect 822 1050 839 1064
rect 871 1050 888 1064
tri 1015 1058 1030 1073 ne
tri 1030 1058 1052 1080 sw
rect 653 1000 668 1008
rect 734 1036 794 1050
rect 749 1026 794 1036
rect 749 1008 777 1026
tri 653 985 668 1000 ne
tri 668 985 690 1007 sw
rect 734 998 777 1008
rect 792 1022 794 1026
rect 916 1036 976 1050
tri 1030 1045 1043 1058 ne
rect 1043 1052 1052 1058
tri 1052 1052 1058 1058 sw
rect 916 1026 961 1036
rect 792 998 866 1022
rect 734 994 866 998
tri 866 994 894 1022 sw
rect 916 1012 918 1026
tri 916 1010 918 1012 ne
rect 930 1008 961 1026
rect 930 998 976 1008
rect 1043 1037 1058 1052
tri 668 973 680 985 ne
rect 680 980 690 985
tri 690 980 695 985 sw
rect 579 634 594 862
rect 680 824 695 980
rect 734 938 762 994
tri 854 976 872 994 ne
rect 872 974 894 994
tri 894 974 914 994 sw
tri 930 980 948 998 ne
rect 753 904 762 938
rect 796 965 838 966
rect 796 931 801 965
rect 831 931 838 965
rect 796 922 838 931
rect 872 965 914 974
rect 872 931 879 965
rect 909 931 914 965
rect 872 926 914 931
rect 948 938 976 998
tri 1021 985 1043 1007 se
rect 1043 1000 1058 1008
tri 1043 985 1058 1000 nw
tri 1015 979 1021 985 se
rect 1021 979 1030 985
rect 734 894 762 904
tri 762 894 786 918 sw
rect 734 862 776 894
tri 793 886 794 887 sw
rect 793 862 794 886
tri 796 885 833 922 ne
rect 833 894 838 922
tri 838 894 864 920 sw
rect 948 904 957 938
rect 948 894 976 904
rect 833 885 917 894
tri 833 866 852 885 ne
rect 852 866 917 885
rect 734 840 794 862
rect 916 862 917 866
rect 934 862 976 894
rect 916 840 976 862
rect 822 824 839 838
rect 871 824 888 838
tri 659 788 681 810 se
rect 681 803 696 824
tri 681 788 696 803 nw
rect 1015 803 1030 979
tri 1030 972 1043 985 nw
rect 1116 904 1131 1132
tri 653 782 659 788 se
rect 659 782 668 788
rect 653 766 668 782
tri 668 775 681 788 nw
rect 822 780 839 794
rect 871 780 888 794
tri 1015 788 1030 803 ne
tri 1030 788 1052 810 sw
rect 653 730 668 738
rect 734 766 794 780
rect 749 756 794 766
rect 749 738 777 756
tri 653 715 668 730 ne
tri 668 715 690 737 sw
rect 734 728 777 738
rect 792 752 794 756
rect 916 766 976 780
tri 1030 775 1043 788 ne
rect 1043 782 1052 788
tri 1052 782 1058 788 sw
rect 916 756 961 766
rect 792 728 866 752
rect 734 724 866 728
tri 866 724 894 752 sw
rect 916 742 918 756
tri 916 740 918 742 ne
rect 930 738 961 756
rect 930 728 976 738
rect 1043 767 1058 782
tri 668 703 680 715 ne
rect 680 710 690 715
tri 690 710 695 715 sw
rect 579 364 594 592
rect 680 554 695 710
rect 734 668 762 724
tri 854 706 872 724 ne
rect 872 704 894 724
tri 894 704 914 724 sw
tri 930 710 948 728 ne
rect 753 634 762 668
rect 796 695 838 696
rect 796 661 801 695
rect 831 661 838 695
rect 796 652 838 661
rect 872 695 914 704
rect 872 661 879 695
rect 909 661 914 695
rect 872 656 914 661
rect 948 668 976 728
tri 1021 715 1043 737 se
rect 1043 730 1058 738
tri 1043 715 1058 730 nw
tri 1015 709 1021 715 se
rect 1021 709 1030 715
rect 734 624 762 634
tri 762 624 786 648 sw
rect 734 592 776 624
tri 793 616 794 617 sw
rect 793 592 794 616
tri 796 615 833 652 ne
rect 833 624 838 652
tri 838 624 864 650 sw
rect 948 634 957 668
rect 948 624 976 634
rect 833 615 917 624
tri 833 596 852 615 ne
rect 852 596 917 615
rect 734 570 794 592
rect 916 592 917 596
rect 934 592 976 624
rect 916 570 976 592
rect 822 554 839 568
rect 871 554 888 568
tri 659 518 681 540 se
rect 681 533 696 554
tri 681 518 696 533 nw
rect 1015 533 1030 709
tri 1030 702 1043 715 nw
rect 1116 634 1131 862
tri 653 512 659 518 se
rect 659 512 668 518
rect 653 496 668 512
tri 668 505 681 518 nw
rect 822 510 839 524
rect 871 510 888 524
tri 1015 518 1030 533 ne
tri 1030 518 1052 540 sw
rect 653 460 668 468
rect 734 496 794 510
rect 749 486 794 496
rect 749 468 777 486
tri 653 445 668 460 ne
tri 668 445 690 467 sw
rect 734 458 777 468
rect 792 482 794 486
rect 916 496 976 510
tri 1030 505 1043 518 ne
rect 1043 512 1052 518
tri 1052 512 1058 518 sw
rect 916 486 961 496
rect 792 458 866 482
rect 734 454 866 458
tri 866 454 894 482 sw
rect 916 472 918 486
tri 916 470 918 472 ne
rect 930 468 961 486
rect 930 458 976 468
rect 1043 497 1058 512
tri 668 433 680 445 ne
rect 680 440 690 445
tri 690 440 695 445 sw
rect 579 94 594 322
rect 680 284 695 440
rect 734 398 762 454
tri 854 436 872 454 ne
rect 872 434 894 454
tri 894 434 914 454 sw
tri 930 440 948 458 ne
rect 753 364 762 398
rect 796 425 838 426
rect 796 391 801 425
rect 831 391 838 425
rect 796 382 838 391
rect 872 425 914 434
rect 872 391 879 425
rect 909 391 914 425
rect 872 386 914 391
rect 948 398 976 458
tri 1021 445 1043 467 se
rect 1043 460 1058 468
tri 1043 445 1058 460 nw
tri 1015 439 1021 445 se
rect 1021 439 1030 445
rect 734 354 762 364
tri 762 354 786 378 sw
rect 734 322 776 354
tri 793 346 794 347 sw
rect 793 322 794 346
tri 796 345 833 382 ne
rect 833 354 838 382
tri 838 354 864 380 sw
rect 948 364 957 398
rect 948 354 976 364
rect 833 345 917 354
tri 833 326 852 345 ne
rect 852 326 917 345
rect 734 300 794 322
rect 916 322 917 326
rect 934 322 976 354
rect 916 300 976 322
rect 822 284 839 298
rect 871 284 888 298
tri 659 248 681 270 se
rect 681 263 696 284
tri 681 248 696 263 nw
rect 1015 263 1030 439
tri 1030 432 1043 445 nw
rect 1116 364 1131 592
tri 653 242 659 248 se
rect 659 242 668 248
rect 653 226 668 242
tri 668 235 681 248 nw
rect 822 240 839 254
rect 871 240 888 254
tri 1015 248 1030 263 ne
tri 1030 248 1052 270 sw
rect 653 190 668 198
rect 734 226 794 240
rect 749 216 794 226
rect 749 198 777 216
tri 653 175 668 190 ne
tri 668 175 690 197 sw
rect 734 188 777 198
rect 792 212 794 216
rect 916 226 976 240
tri 1030 235 1043 248 ne
rect 1043 242 1052 248
tri 1052 242 1058 248 sw
rect 916 216 961 226
rect 792 188 866 212
rect 734 184 866 188
tri 866 184 894 212 sw
rect 916 202 918 216
tri 916 200 918 202 ne
rect 930 198 961 216
rect 930 188 976 198
rect 1043 227 1058 242
tri 668 163 680 175 ne
rect 680 170 690 175
tri 690 170 695 175 sw
rect 579 -176 594 52
rect 680 14 695 170
rect 734 128 762 184
tri 854 166 872 184 ne
rect 872 164 894 184
tri 894 164 914 184 sw
tri 930 170 948 188 ne
rect 753 94 762 128
rect 796 155 838 156
rect 796 121 801 155
rect 831 121 838 155
rect 796 112 838 121
rect 872 155 914 164
rect 872 121 879 155
rect 909 121 914 155
rect 872 116 914 121
rect 948 128 976 188
tri 1021 175 1043 197 se
rect 1043 190 1058 198
tri 1043 175 1058 190 nw
tri 1015 169 1021 175 se
rect 1021 169 1030 175
rect 734 84 762 94
tri 762 84 786 108 sw
rect 734 52 776 84
tri 793 76 794 77 sw
rect 793 52 794 76
tri 796 75 833 112 ne
rect 833 84 838 112
tri 838 84 864 110 sw
rect 948 94 957 128
rect 948 84 976 94
rect 833 75 917 84
tri 833 56 852 75 ne
rect 852 56 917 75
rect 734 30 794 52
rect 916 52 917 56
rect 934 52 976 84
rect 916 30 976 52
rect 822 14 839 28
rect 871 14 888 28
tri 659 -22 681 0 se
rect 681 -7 696 14
tri 681 -22 696 -7 nw
rect 1015 -7 1030 169
tri 1030 162 1043 175 nw
rect 1116 94 1131 322
tri 653 -28 659 -22 se
rect 659 -28 668 -22
rect 653 -44 668 -28
tri 668 -35 681 -22 nw
rect 822 -30 839 -16
rect 871 -30 888 -16
tri 1015 -22 1030 -7 ne
tri 1030 -22 1052 0 sw
rect 653 -80 668 -72
rect 734 -44 794 -30
rect 749 -54 794 -44
rect 749 -72 777 -54
tri 653 -95 668 -80 ne
tri 668 -95 690 -73 sw
rect 734 -82 777 -72
rect 792 -58 794 -54
rect 916 -44 976 -30
tri 1030 -35 1043 -22 ne
rect 1043 -28 1052 -22
tri 1052 -28 1058 -22 sw
rect 916 -54 961 -44
rect 792 -82 866 -58
rect 734 -86 866 -82
tri 866 -86 894 -58 sw
rect 916 -68 918 -54
tri 916 -70 918 -68 ne
rect 930 -72 961 -54
rect 930 -82 976 -72
rect 1043 -43 1058 -28
tri 668 -107 680 -95 ne
rect 680 -100 690 -95
tri 690 -100 695 -95 sw
rect 579 -446 594 -218
rect 680 -256 695 -100
rect 734 -142 762 -86
tri 854 -104 872 -86 ne
rect 872 -106 894 -86
tri 894 -106 914 -86 sw
tri 930 -100 948 -82 ne
rect 753 -176 762 -142
rect 796 -115 838 -114
rect 796 -149 801 -115
rect 831 -149 838 -115
rect 796 -158 838 -149
rect 872 -115 914 -106
rect 872 -149 879 -115
rect 909 -149 914 -115
rect 872 -154 914 -149
rect 948 -142 976 -82
tri 1021 -95 1043 -73 se
rect 1043 -80 1058 -72
tri 1043 -95 1058 -80 nw
tri 1015 -101 1021 -95 se
rect 1021 -101 1030 -95
rect 734 -186 762 -176
tri 762 -186 786 -162 sw
rect 734 -218 776 -186
tri 793 -194 794 -193 sw
rect 793 -218 794 -194
tri 796 -195 833 -158 ne
rect 833 -186 838 -158
tri 838 -186 864 -160 sw
rect 948 -176 957 -142
rect 948 -186 976 -176
rect 833 -195 917 -186
tri 833 -214 852 -195 ne
rect 852 -214 917 -195
rect 734 -240 794 -218
rect 916 -218 917 -214
rect 934 -218 976 -186
rect 916 -240 976 -218
rect 822 -256 839 -242
rect 871 -256 888 -242
tri 659 -292 681 -270 se
rect 681 -277 696 -256
tri 681 -292 696 -277 nw
rect 1015 -277 1030 -101
tri 1030 -108 1043 -95 nw
rect 1116 -176 1131 52
tri 653 -298 659 -292 se
rect 659 -298 668 -292
rect 653 -314 668 -298
tri 668 -305 681 -292 nw
rect 822 -300 839 -286
rect 871 -300 888 -286
tri 1015 -292 1030 -277 ne
tri 1030 -292 1052 -270 sw
rect 653 -350 668 -342
rect 734 -314 794 -300
rect 749 -324 794 -314
rect 749 -342 777 -324
tri 653 -365 668 -350 ne
tri 668 -365 690 -343 sw
rect 734 -352 777 -342
rect 792 -328 794 -324
rect 916 -314 976 -300
tri 1030 -305 1043 -292 ne
rect 1043 -298 1052 -292
tri 1052 -298 1058 -292 sw
rect 916 -324 961 -314
rect 792 -352 866 -328
rect 734 -356 866 -352
tri 866 -356 894 -328 sw
rect 916 -338 918 -324
tri 916 -340 918 -338 ne
rect 930 -342 961 -324
rect 930 -352 976 -342
rect 1043 -313 1058 -298
tri 668 -377 680 -365 ne
rect 680 -370 690 -365
tri 690 -370 695 -365 sw
rect 579 -716 594 -488
rect 680 -526 695 -370
rect 734 -412 762 -356
tri 854 -374 872 -356 ne
rect 872 -376 894 -356
tri 894 -376 914 -356 sw
tri 930 -370 948 -352 ne
rect 753 -446 762 -412
rect 796 -385 838 -384
rect 796 -419 801 -385
rect 831 -419 838 -385
rect 796 -428 838 -419
rect 872 -385 914 -376
rect 872 -419 879 -385
rect 909 -419 914 -385
rect 872 -424 914 -419
rect 948 -412 976 -352
tri 1021 -365 1043 -343 se
rect 1043 -350 1058 -342
tri 1043 -365 1058 -350 nw
tri 1015 -371 1021 -365 se
rect 1021 -371 1030 -365
rect 734 -456 762 -446
tri 762 -456 786 -432 sw
rect 734 -488 776 -456
tri 793 -464 794 -463 sw
rect 793 -488 794 -464
tri 796 -465 833 -428 ne
rect 833 -456 838 -428
tri 838 -456 864 -430 sw
rect 948 -446 957 -412
rect 948 -456 976 -446
rect 833 -465 917 -456
tri 833 -484 852 -465 ne
rect 852 -484 917 -465
rect 734 -510 794 -488
rect 916 -488 917 -484
rect 934 -488 976 -456
rect 916 -510 976 -488
rect 822 -526 839 -512
rect 871 -526 888 -512
tri 659 -562 681 -540 se
rect 681 -547 696 -526
tri 681 -562 696 -547 nw
rect 1015 -547 1030 -371
tri 1030 -378 1043 -365 nw
rect 1116 -446 1131 -218
tri 653 -568 659 -562 se
rect 659 -568 668 -562
rect 653 -584 668 -568
tri 668 -575 681 -562 nw
rect 822 -570 839 -556
rect 871 -570 888 -556
tri 1015 -562 1030 -547 ne
tri 1030 -562 1052 -540 sw
rect 653 -620 668 -612
rect 734 -584 794 -570
rect 749 -594 794 -584
rect 749 -612 777 -594
tri 653 -635 668 -620 ne
tri 668 -635 690 -613 sw
rect 734 -622 777 -612
rect 792 -598 794 -594
rect 916 -584 976 -570
tri 1030 -575 1043 -562 ne
rect 1043 -568 1052 -562
tri 1052 -568 1058 -562 sw
rect 916 -594 961 -584
rect 792 -622 866 -598
rect 734 -626 866 -622
tri 866 -626 894 -598 sw
rect 916 -608 918 -594
tri 916 -610 918 -608 ne
rect 930 -612 961 -594
rect 930 -622 976 -612
rect 1043 -583 1058 -568
tri 668 -647 680 -635 ne
rect 680 -640 690 -635
tri 690 -640 695 -635 sw
rect 579 -986 594 -758
rect 680 -796 695 -640
rect 734 -682 762 -626
tri 854 -644 872 -626 ne
rect 872 -646 894 -626
tri 894 -646 914 -626 sw
tri 930 -640 948 -622 ne
rect 753 -716 762 -682
rect 796 -655 838 -654
rect 796 -689 801 -655
rect 831 -689 838 -655
rect 796 -698 838 -689
rect 872 -655 914 -646
rect 872 -689 879 -655
rect 909 -689 914 -655
rect 872 -694 914 -689
rect 948 -682 976 -622
tri 1021 -635 1043 -613 se
rect 1043 -620 1058 -612
tri 1043 -635 1058 -620 nw
tri 1015 -641 1021 -635 se
rect 1021 -641 1030 -635
rect 734 -726 762 -716
tri 762 -726 786 -702 sw
rect 734 -758 776 -726
tri 793 -734 794 -733 sw
rect 793 -758 794 -734
tri 796 -735 833 -698 ne
rect 833 -726 838 -698
tri 838 -726 864 -700 sw
rect 948 -716 957 -682
rect 948 -726 976 -716
rect 833 -735 917 -726
tri 833 -754 852 -735 ne
rect 852 -754 917 -735
rect 734 -780 794 -758
rect 916 -758 917 -754
rect 934 -758 976 -726
rect 916 -780 976 -758
rect 822 -796 839 -782
rect 871 -796 888 -782
tri 659 -832 681 -810 se
rect 681 -817 696 -796
tri 681 -832 696 -817 nw
rect 1015 -817 1030 -641
tri 1030 -648 1043 -635 nw
rect 1116 -716 1131 -488
tri 653 -838 659 -832 se
rect 659 -838 668 -832
rect 653 -854 668 -838
tri 668 -845 681 -832 nw
rect 822 -840 839 -826
rect 871 -840 888 -826
tri 1015 -832 1030 -817 ne
tri 1030 -832 1052 -810 sw
rect 653 -890 668 -882
rect 734 -854 794 -840
rect 749 -864 794 -854
rect 749 -882 777 -864
tri 653 -905 668 -890 ne
tri 668 -905 690 -883 sw
rect 734 -892 777 -882
rect 792 -868 794 -864
rect 916 -854 976 -840
tri 1030 -845 1043 -832 ne
rect 1043 -838 1052 -832
tri 1052 -838 1058 -832 sw
rect 916 -864 961 -854
rect 792 -892 866 -868
rect 734 -896 866 -892
tri 866 -896 894 -868 sw
rect 916 -878 918 -864
tri 916 -880 918 -878 ne
rect 930 -882 961 -864
rect 930 -892 976 -882
rect 1043 -853 1058 -838
tri 668 -917 680 -905 ne
rect 680 -910 690 -905
tri 690 -910 695 -905 sw
rect 579 -1256 594 -1028
rect 680 -1066 695 -910
rect 734 -952 762 -896
tri 854 -914 872 -896 ne
rect 872 -916 894 -896
tri 894 -916 914 -896 sw
tri 930 -910 948 -892 ne
rect 753 -986 762 -952
rect 796 -925 838 -924
rect 796 -959 801 -925
rect 831 -959 838 -925
rect 796 -968 838 -959
rect 872 -925 914 -916
rect 872 -959 879 -925
rect 909 -959 914 -925
rect 872 -964 914 -959
rect 948 -952 976 -892
tri 1021 -905 1043 -883 se
rect 1043 -890 1058 -882
tri 1043 -905 1058 -890 nw
tri 1015 -911 1021 -905 se
rect 1021 -911 1030 -905
rect 734 -996 762 -986
tri 762 -996 786 -972 sw
rect 734 -1028 776 -996
tri 793 -1004 794 -1003 sw
rect 793 -1028 794 -1004
tri 796 -1005 833 -968 ne
rect 833 -996 838 -968
tri 838 -996 864 -970 sw
rect 948 -986 957 -952
rect 948 -996 976 -986
rect 833 -1005 917 -996
tri 833 -1024 852 -1005 ne
rect 852 -1024 917 -1005
rect 734 -1050 794 -1028
rect 916 -1028 917 -1024
rect 934 -1028 976 -996
rect 916 -1050 976 -1028
rect 822 -1066 839 -1052
rect 871 -1066 888 -1052
tri 659 -1102 681 -1080 se
rect 681 -1087 696 -1066
tri 681 -1102 696 -1087 nw
rect 1015 -1087 1030 -911
tri 1030 -918 1043 -905 nw
rect 1116 -986 1131 -758
tri 653 -1108 659 -1102 se
rect 659 -1108 668 -1102
rect 653 -1124 668 -1108
tri 668 -1115 681 -1102 nw
rect 822 -1110 839 -1096
rect 871 -1110 888 -1096
tri 1015 -1102 1030 -1087 ne
tri 1030 -1102 1052 -1080 sw
rect 653 -1160 668 -1152
rect 734 -1124 794 -1110
rect 749 -1134 794 -1124
rect 749 -1152 777 -1134
tri 653 -1175 668 -1160 ne
tri 668 -1175 690 -1153 sw
rect 734 -1162 777 -1152
rect 792 -1138 794 -1134
rect 916 -1124 976 -1110
tri 1030 -1115 1043 -1102 ne
rect 1043 -1108 1052 -1102
tri 1052 -1108 1058 -1102 sw
rect 916 -1134 961 -1124
rect 792 -1162 866 -1138
rect 734 -1166 866 -1162
tri 866 -1166 894 -1138 sw
rect 916 -1148 918 -1134
tri 916 -1150 918 -1148 ne
rect 930 -1152 961 -1134
rect 930 -1162 976 -1152
rect 1043 -1123 1058 -1108
tri 668 -1187 680 -1175 ne
rect 680 -1180 690 -1175
tri 690 -1180 695 -1175 sw
rect 579 -1526 594 -1298
rect 680 -1336 695 -1180
rect 734 -1222 762 -1166
tri 854 -1184 872 -1166 ne
rect 872 -1186 894 -1166
tri 894 -1186 914 -1166 sw
tri 930 -1180 948 -1162 ne
rect 753 -1256 762 -1222
rect 796 -1195 838 -1194
rect 796 -1229 801 -1195
rect 831 -1229 838 -1195
rect 796 -1238 838 -1229
rect 872 -1195 914 -1186
rect 872 -1229 879 -1195
rect 909 -1229 914 -1195
rect 872 -1234 914 -1229
rect 948 -1222 976 -1162
tri 1021 -1175 1043 -1153 se
rect 1043 -1160 1058 -1152
tri 1043 -1175 1058 -1160 nw
tri 1015 -1181 1021 -1175 se
rect 1021 -1181 1030 -1175
rect 734 -1266 762 -1256
tri 762 -1266 786 -1242 sw
rect 734 -1298 776 -1266
tri 793 -1274 794 -1273 sw
rect 793 -1298 794 -1274
tri 796 -1275 833 -1238 ne
rect 833 -1266 838 -1238
tri 838 -1266 864 -1240 sw
rect 948 -1256 957 -1222
rect 948 -1266 976 -1256
rect 833 -1275 917 -1266
tri 833 -1294 852 -1275 ne
rect 852 -1294 917 -1275
rect 734 -1320 794 -1298
rect 916 -1298 917 -1294
rect 934 -1298 976 -1266
rect 916 -1320 976 -1298
rect 822 -1336 839 -1322
rect 871 -1336 888 -1322
tri 659 -1372 681 -1350 se
rect 681 -1357 696 -1336
tri 681 -1372 696 -1357 nw
rect 1015 -1357 1030 -1181
tri 1030 -1188 1043 -1175 nw
rect 1116 -1256 1131 -1028
tri 653 -1378 659 -1372 se
rect 659 -1378 668 -1372
rect 653 -1394 668 -1378
tri 668 -1385 681 -1372 nw
rect 822 -1380 839 -1366
rect 871 -1380 888 -1366
tri 1015 -1372 1030 -1357 ne
tri 1030 -1372 1052 -1350 sw
rect 653 -1430 668 -1422
rect 734 -1394 794 -1380
rect 749 -1404 794 -1394
rect 749 -1422 777 -1404
tri 653 -1445 668 -1430 ne
tri 668 -1445 690 -1423 sw
rect 734 -1432 777 -1422
rect 792 -1408 794 -1404
rect 916 -1394 976 -1380
tri 1030 -1385 1043 -1372 ne
rect 1043 -1378 1052 -1372
tri 1052 -1378 1058 -1372 sw
rect 916 -1404 961 -1394
rect 792 -1432 866 -1408
rect 734 -1436 866 -1432
tri 866 -1436 894 -1408 sw
rect 916 -1418 918 -1404
tri 916 -1420 918 -1418 ne
rect 930 -1422 961 -1404
rect 930 -1432 976 -1422
rect 1043 -1393 1058 -1378
tri 668 -1457 680 -1445 ne
rect 680 -1450 690 -1445
tri 690 -1450 695 -1445 sw
rect 579 -1796 594 -1568
rect 680 -1606 695 -1450
rect 734 -1492 762 -1436
tri 854 -1454 872 -1436 ne
rect 872 -1456 894 -1436
tri 894 -1456 914 -1436 sw
tri 930 -1450 948 -1432 ne
rect 753 -1526 762 -1492
rect 796 -1465 838 -1464
rect 796 -1499 801 -1465
rect 831 -1499 838 -1465
rect 796 -1508 838 -1499
rect 872 -1465 914 -1456
rect 872 -1499 879 -1465
rect 909 -1499 914 -1465
rect 872 -1504 914 -1499
rect 948 -1492 976 -1432
tri 1021 -1445 1043 -1423 se
rect 1043 -1430 1058 -1422
tri 1043 -1445 1058 -1430 nw
tri 1015 -1451 1021 -1445 se
rect 1021 -1451 1030 -1445
rect 734 -1536 762 -1526
tri 762 -1536 786 -1512 sw
rect 734 -1568 776 -1536
tri 793 -1544 794 -1543 sw
rect 793 -1568 794 -1544
tri 796 -1545 833 -1508 ne
rect 833 -1536 838 -1508
tri 838 -1536 864 -1510 sw
rect 948 -1526 957 -1492
rect 948 -1536 976 -1526
rect 833 -1545 917 -1536
tri 833 -1564 852 -1545 ne
rect 852 -1564 917 -1545
rect 734 -1590 794 -1568
rect 916 -1568 917 -1564
rect 934 -1568 976 -1536
rect 916 -1590 976 -1568
rect 822 -1606 839 -1592
rect 871 -1606 888 -1592
tri 659 -1642 681 -1620 se
rect 681 -1627 696 -1606
tri 681 -1642 696 -1627 nw
rect 1015 -1627 1030 -1451
tri 1030 -1458 1043 -1445 nw
rect 1116 -1526 1131 -1298
tri 653 -1648 659 -1642 se
rect 659 -1648 668 -1642
rect 653 -1664 668 -1648
tri 668 -1655 681 -1642 nw
rect 822 -1650 839 -1636
rect 871 -1650 888 -1636
tri 1015 -1642 1030 -1627 ne
tri 1030 -1642 1052 -1620 sw
rect 653 -1700 668 -1692
rect 734 -1664 794 -1650
rect 749 -1674 794 -1664
rect 749 -1692 777 -1674
tri 653 -1715 668 -1700 ne
tri 668 -1715 690 -1693 sw
rect 734 -1702 777 -1692
rect 792 -1678 794 -1674
rect 916 -1664 976 -1650
tri 1030 -1655 1043 -1642 ne
rect 1043 -1648 1052 -1642
tri 1052 -1648 1058 -1642 sw
rect 916 -1674 961 -1664
rect 792 -1702 866 -1678
rect 734 -1706 866 -1702
tri 866 -1706 894 -1678 sw
rect 916 -1688 918 -1674
tri 916 -1690 918 -1688 ne
rect 930 -1692 961 -1674
rect 930 -1702 976 -1692
rect 1043 -1663 1058 -1648
tri 668 -1727 680 -1715 ne
rect 680 -1720 690 -1715
tri 690 -1720 695 -1715 sw
rect 579 -2066 594 -1838
rect 680 -1876 695 -1720
rect 734 -1762 762 -1706
tri 854 -1724 872 -1706 ne
rect 872 -1726 894 -1706
tri 894 -1726 914 -1706 sw
tri 930 -1720 948 -1702 ne
rect 753 -1796 762 -1762
rect 796 -1735 838 -1734
rect 796 -1769 801 -1735
rect 831 -1769 838 -1735
rect 796 -1778 838 -1769
rect 872 -1735 914 -1726
rect 872 -1769 879 -1735
rect 909 -1769 914 -1735
rect 872 -1774 914 -1769
rect 948 -1762 976 -1702
tri 1021 -1715 1043 -1693 se
rect 1043 -1700 1058 -1692
tri 1043 -1715 1058 -1700 nw
tri 1015 -1721 1021 -1715 se
rect 1021 -1721 1030 -1715
rect 734 -1806 762 -1796
tri 762 -1806 786 -1782 sw
rect 734 -1838 776 -1806
tri 793 -1814 794 -1813 sw
rect 793 -1838 794 -1814
tri 796 -1815 833 -1778 ne
rect 833 -1806 838 -1778
tri 838 -1806 864 -1780 sw
rect 948 -1796 957 -1762
rect 948 -1806 976 -1796
rect 833 -1815 917 -1806
tri 833 -1834 852 -1815 ne
rect 852 -1834 917 -1815
rect 734 -1860 794 -1838
rect 916 -1838 917 -1834
rect 934 -1838 976 -1806
rect 916 -1860 976 -1838
rect 822 -1876 839 -1862
rect 871 -1876 888 -1862
tri 659 -1912 681 -1890 se
rect 681 -1897 696 -1876
tri 681 -1912 696 -1897 nw
rect 1015 -1897 1030 -1721
tri 1030 -1728 1043 -1715 nw
rect 1116 -1796 1131 -1568
tri 653 -1918 659 -1912 se
rect 659 -1918 668 -1912
rect 653 -1934 668 -1918
tri 668 -1925 681 -1912 nw
rect 822 -1920 839 -1906
rect 871 -1920 888 -1906
tri 1015 -1912 1030 -1897 ne
tri 1030 -1912 1052 -1890 sw
rect 653 -1970 668 -1962
rect 734 -1934 794 -1920
rect 749 -1944 794 -1934
rect 749 -1962 777 -1944
tri 653 -1985 668 -1970 ne
tri 668 -1985 690 -1963 sw
rect 734 -1972 777 -1962
rect 792 -1948 794 -1944
rect 916 -1934 976 -1920
tri 1030 -1925 1043 -1912 ne
rect 1043 -1918 1052 -1912
tri 1052 -1918 1058 -1912 sw
rect 916 -1944 961 -1934
rect 792 -1972 866 -1948
rect 734 -1976 866 -1972
tri 866 -1976 894 -1948 sw
rect 916 -1958 918 -1944
tri 916 -1960 918 -1958 ne
rect 930 -1962 961 -1944
rect 930 -1972 976 -1962
rect 1043 -1933 1058 -1918
tri 668 -1997 680 -1985 ne
rect 680 -1990 690 -1985
tri 690 -1990 695 -1985 sw
rect 579 -2146 594 -2108
rect 680 -2146 695 -1990
rect 734 -2032 762 -1976
tri 854 -1994 872 -1976 ne
rect 872 -1996 894 -1976
tri 894 -1996 914 -1976 sw
tri 930 -1990 948 -1972 ne
rect 753 -2066 762 -2032
rect 796 -2005 838 -2004
rect 796 -2039 801 -2005
rect 831 -2039 838 -2005
rect 796 -2048 838 -2039
rect 872 -2005 914 -1996
rect 872 -2039 879 -2005
rect 909 -2039 914 -2005
rect 872 -2044 914 -2039
rect 948 -2032 976 -1972
tri 1021 -1985 1043 -1963 se
rect 1043 -1970 1058 -1962
tri 1043 -1985 1058 -1970 nw
tri 1015 -1991 1021 -1985 se
rect 1021 -1991 1030 -1985
rect 734 -2076 762 -2066
tri 762 -2076 786 -2052 sw
rect 734 -2108 776 -2076
tri 793 -2084 794 -2083 sw
rect 793 -2108 794 -2084
tri 796 -2085 833 -2048 ne
rect 833 -2076 838 -2048
tri 838 -2076 864 -2050 sw
rect 948 -2066 957 -2032
rect 948 -2076 976 -2066
rect 833 -2085 917 -2076
tri 833 -2104 852 -2085 ne
rect 852 -2104 917 -2085
rect 734 -2130 794 -2108
rect 916 -2108 917 -2104
rect 934 -2108 976 -2076
rect 916 -2130 976 -2108
rect 822 -2146 839 -2132
rect 871 -2146 888 -2132
rect 1015 -2146 1030 -1991
tri 1030 -1998 1043 -1985 nw
rect 1116 -2066 1131 -1838
rect 1116 -2146 1131 -2108
rect 1159 1984 1174 2174
tri 1239 2138 1261 2160 se
rect 1261 2153 1276 2174
tri 1261 2138 1276 2153 nw
rect 1595 2153 1610 2174
tri 1233 2132 1239 2138 se
rect 1239 2132 1248 2138
rect 1233 2116 1248 2132
tri 1248 2125 1261 2138 nw
rect 1402 2130 1419 2144
rect 1451 2130 1468 2144
tri 1595 2138 1610 2153 ne
tri 1610 2138 1632 2160 sw
rect 1233 2080 1248 2088
rect 1314 2116 1374 2130
rect 1329 2106 1374 2116
rect 1329 2088 1357 2106
tri 1233 2065 1248 2080 ne
tri 1248 2065 1270 2087 sw
rect 1314 2078 1357 2088
rect 1372 2102 1374 2106
rect 1496 2116 1556 2130
tri 1610 2125 1623 2138 ne
rect 1623 2132 1632 2138
tri 1632 2132 1638 2138 sw
rect 1496 2106 1541 2116
rect 1372 2078 1446 2102
rect 1314 2074 1446 2078
tri 1446 2074 1474 2102 sw
rect 1496 2092 1498 2106
tri 1496 2090 1498 2092 ne
rect 1510 2088 1541 2106
rect 1510 2078 1556 2088
rect 1623 2117 1638 2132
tri 1248 2053 1260 2065 ne
rect 1260 2060 1270 2065
tri 1270 2060 1275 2065 sw
rect 1159 1714 1174 1942
rect 1260 1904 1275 2060
rect 1314 2018 1342 2074
tri 1434 2056 1452 2074 ne
rect 1452 2054 1474 2074
tri 1474 2054 1494 2074 sw
tri 1510 2060 1528 2078 ne
rect 1333 1984 1342 2018
rect 1376 2045 1418 2046
rect 1376 2011 1381 2045
rect 1411 2011 1418 2045
rect 1376 2002 1418 2011
rect 1452 2045 1494 2054
rect 1452 2011 1459 2045
rect 1489 2011 1494 2045
rect 1452 2006 1494 2011
rect 1528 2018 1556 2078
tri 1601 2065 1623 2087 se
rect 1623 2080 1638 2088
tri 1623 2065 1638 2080 nw
tri 1595 2059 1601 2065 se
rect 1601 2059 1610 2065
rect 1314 1974 1342 1984
tri 1342 1974 1366 1998 sw
rect 1314 1942 1356 1974
tri 1373 1966 1374 1967 sw
rect 1373 1942 1374 1966
tri 1376 1965 1413 2002 ne
rect 1413 1974 1418 2002
tri 1418 1974 1444 2000 sw
rect 1528 1984 1537 2018
rect 1528 1974 1556 1984
rect 1413 1965 1497 1974
tri 1413 1946 1432 1965 ne
rect 1432 1946 1497 1965
rect 1314 1920 1374 1942
rect 1496 1942 1497 1946
rect 1514 1942 1556 1974
rect 1496 1920 1556 1942
rect 1402 1904 1419 1918
rect 1451 1904 1468 1918
tri 1239 1868 1261 1890 se
rect 1261 1883 1276 1904
tri 1261 1868 1276 1883 nw
rect 1595 1883 1610 2059
tri 1610 2052 1623 2065 nw
rect 1696 1984 1711 2174
tri 1233 1862 1239 1868 se
rect 1239 1862 1248 1868
rect 1233 1846 1248 1862
tri 1248 1855 1261 1868 nw
rect 1402 1860 1419 1874
rect 1451 1860 1468 1874
tri 1595 1868 1610 1883 ne
tri 1610 1868 1632 1890 sw
rect 1233 1810 1248 1818
rect 1314 1846 1374 1860
rect 1329 1836 1374 1846
rect 1329 1818 1357 1836
tri 1233 1795 1248 1810 ne
tri 1248 1795 1270 1817 sw
rect 1314 1808 1357 1818
rect 1372 1832 1374 1836
rect 1496 1846 1556 1860
tri 1610 1855 1623 1868 ne
rect 1623 1862 1632 1868
tri 1632 1862 1638 1868 sw
rect 1496 1836 1541 1846
rect 1372 1808 1446 1832
rect 1314 1804 1446 1808
tri 1446 1804 1474 1832 sw
rect 1496 1822 1498 1836
tri 1496 1820 1498 1822 ne
rect 1510 1818 1541 1836
rect 1510 1808 1556 1818
rect 1623 1847 1638 1862
tri 1248 1783 1260 1795 ne
rect 1260 1790 1270 1795
tri 1270 1790 1275 1795 sw
rect 1159 1444 1174 1672
rect 1260 1634 1275 1790
rect 1314 1748 1342 1804
tri 1434 1786 1452 1804 ne
rect 1452 1784 1474 1804
tri 1474 1784 1494 1804 sw
tri 1510 1790 1528 1808 ne
rect 1333 1714 1342 1748
rect 1376 1775 1418 1776
rect 1376 1741 1381 1775
rect 1411 1741 1418 1775
rect 1376 1732 1418 1741
rect 1452 1775 1494 1784
rect 1452 1741 1459 1775
rect 1489 1741 1494 1775
rect 1452 1736 1494 1741
rect 1528 1748 1556 1808
tri 1601 1795 1623 1817 se
rect 1623 1810 1638 1818
tri 1623 1795 1638 1810 nw
tri 1595 1789 1601 1795 se
rect 1601 1789 1610 1795
rect 1314 1704 1342 1714
tri 1342 1704 1366 1728 sw
rect 1314 1672 1356 1704
tri 1373 1696 1374 1697 sw
rect 1373 1672 1374 1696
tri 1376 1695 1413 1732 ne
rect 1413 1704 1418 1732
tri 1418 1704 1444 1730 sw
rect 1528 1714 1537 1748
rect 1528 1704 1556 1714
rect 1413 1695 1497 1704
tri 1413 1676 1432 1695 ne
rect 1432 1676 1497 1695
rect 1314 1650 1374 1672
rect 1496 1672 1497 1676
rect 1514 1672 1556 1704
rect 1496 1650 1556 1672
rect 1402 1634 1419 1648
rect 1451 1634 1468 1648
tri 1239 1598 1261 1620 se
rect 1261 1613 1276 1634
tri 1261 1598 1276 1613 nw
rect 1595 1613 1610 1789
tri 1610 1782 1623 1795 nw
rect 1696 1714 1711 1942
tri 1233 1592 1239 1598 se
rect 1239 1592 1248 1598
rect 1233 1576 1248 1592
tri 1248 1585 1261 1598 nw
rect 1402 1590 1419 1604
rect 1451 1590 1468 1604
tri 1595 1598 1610 1613 ne
tri 1610 1598 1632 1620 sw
rect 1233 1540 1248 1548
rect 1314 1576 1374 1590
rect 1329 1566 1374 1576
rect 1329 1548 1357 1566
tri 1233 1525 1248 1540 ne
tri 1248 1525 1270 1547 sw
rect 1314 1538 1357 1548
rect 1372 1562 1374 1566
rect 1496 1576 1556 1590
tri 1610 1585 1623 1598 ne
rect 1623 1592 1632 1598
tri 1632 1592 1638 1598 sw
rect 1496 1566 1541 1576
rect 1372 1538 1446 1562
rect 1314 1534 1446 1538
tri 1446 1534 1474 1562 sw
rect 1496 1552 1498 1566
tri 1496 1550 1498 1552 ne
rect 1510 1548 1541 1566
rect 1510 1538 1556 1548
rect 1623 1577 1638 1592
tri 1248 1513 1260 1525 ne
rect 1260 1520 1270 1525
tri 1270 1520 1275 1525 sw
rect 1159 1174 1174 1402
rect 1260 1364 1275 1520
rect 1314 1478 1342 1534
tri 1434 1516 1452 1534 ne
rect 1452 1514 1474 1534
tri 1474 1514 1494 1534 sw
tri 1510 1520 1528 1538 ne
rect 1333 1444 1342 1478
rect 1376 1505 1418 1506
rect 1376 1471 1381 1505
rect 1411 1471 1418 1505
rect 1376 1462 1418 1471
rect 1452 1505 1494 1514
rect 1452 1471 1459 1505
rect 1489 1471 1494 1505
rect 1452 1466 1494 1471
rect 1528 1478 1556 1538
tri 1601 1525 1623 1547 se
rect 1623 1540 1638 1548
tri 1623 1525 1638 1540 nw
tri 1595 1519 1601 1525 se
rect 1601 1519 1610 1525
rect 1314 1434 1342 1444
tri 1342 1434 1366 1458 sw
rect 1314 1402 1356 1434
tri 1373 1426 1374 1427 sw
rect 1373 1402 1374 1426
tri 1376 1425 1413 1462 ne
rect 1413 1434 1418 1462
tri 1418 1434 1444 1460 sw
rect 1528 1444 1537 1478
rect 1528 1434 1556 1444
rect 1413 1425 1497 1434
tri 1413 1406 1432 1425 ne
rect 1432 1406 1497 1425
rect 1314 1380 1374 1402
rect 1496 1402 1497 1406
rect 1514 1402 1556 1434
rect 1496 1380 1556 1402
rect 1402 1364 1419 1378
rect 1451 1364 1468 1378
tri 1239 1328 1261 1350 se
rect 1261 1343 1276 1364
tri 1261 1328 1276 1343 nw
rect 1595 1343 1610 1519
tri 1610 1512 1623 1525 nw
rect 1696 1444 1711 1672
tri 1233 1322 1239 1328 se
rect 1239 1322 1248 1328
rect 1233 1306 1248 1322
tri 1248 1315 1261 1328 nw
rect 1402 1320 1419 1334
rect 1451 1320 1468 1334
tri 1595 1328 1610 1343 ne
tri 1610 1328 1632 1350 sw
rect 1233 1270 1248 1278
rect 1314 1306 1374 1320
rect 1329 1296 1374 1306
rect 1329 1278 1357 1296
tri 1233 1255 1248 1270 ne
tri 1248 1255 1270 1277 sw
rect 1314 1268 1357 1278
rect 1372 1292 1374 1296
rect 1496 1306 1556 1320
tri 1610 1315 1623 1328 ne
rect 1623 1322 1632 1328
tri 1632 1322 1638 1328 sw
rect 1496 1296 1541 1306
rect 1372 1268 1446 1292
rect 1314 1264 1446 1268
tri 1446 1264 1474 1292 sw
rect 1496 1282 1498 1296
tri 1496 1280 1498 1282 ne
rect 1510 1278 1541 1296
rect 1510 1268 1556 1278
rect 1623 1307 1638 1322
tri 1248 1243 1260 1255 ne
rect 1260 1250 1270 1255
tri 1270 1250 1275 1255 sw
rect 1159 904 1174 1132
rect 1260 1094 1275 1250
rect 1314 1208 1342 1264
tri 1434 1246 1452 1264 ne
rect 1452 1244 1474 1264
tri 1474 1244 1494 1264 sw
tri 1510 1250 1528 1268 ne
rect 1333 1174 1342 1208
rect 1376 1235 1418 1236
rect 1376 1201 1381 1235
rect 1411 1201 1418 1235
rect 1376 1192 1418 1201
rect 1452 1235 1494 1244
rect 1452 1201 1459 1235
rect 1489 1201 1494 1235
rect 1452 1196 1494 1201
rect 1528 1208 1556 1268
tri 1601 1255 1623 1277 se
rect 1623 1270 1638 1278
tri 1623 1255 1638 1270 nw
tri 1595 1249 1601 1255 se
rect 1601 1249 1610 1255
rect 1314 1164 1342 1174
tri 1342 1164 1366 1188 sw
rect 1314 1132 1356 1164
tri 1373 1156 1374 1157 sw
rect 1373 1132 1374 1156
tri 1376 1155 1413 1192 ne
rect 1413 1164 1418 1192
tri 1418 1164 1444 1190 sw
rect 1528 1174 1537 1208
rect 1528 1164 1556 1174
rect 1413 1155 1497 1164
tri 1413 1136 1432 1155 ne
rect 1432 1136 1497 1155
rect 1314 1110 1374 1132
rect 1496 1132 1497 1136
rect 1514 1132 1556 1164
rect 1496 1110 1556 1132
rect 1402 1094 1419 1108
rect 1451 1094 1468 1108
tri 1239 1058 1261 1080 se
rect 1261 1073 1276 1094
tri 1261 1058 1276 1073 nw
rect 1595 1073 1610 1249
tri 1610 1242 1623 1255 nw
rect 1696 1174 1711 1402
tri 1233 1052 1239 1058 se
rect 1239 1052 1248 1058
rect 1233 1036 1248 1052
tri 1248 1045 1261 1058 nw
rect 1402 1050 1419 1064
rect 1451 1050 1468 1064
tri 1595 1058 1610 1073 ne
tri 1610 1058 1632 1080 sw
rect 1233 1000 1248 1008
rect 1314 1036 1374 1050
rect 1329 1026 1374 1036
rect 1329 1008 1357 1026
tri 1233 985 1248 1000 ne
tri 1248 985 1270 1007 sw
rect 1314 998 1357 1008
rect 1372 1022 1374 1026
rect 1496 1036 1556 1050
tri 1610 1045 1623 1058 ne
rect 1623 1052 1632 1058
tri 1632 1052 1638 1058 sw
rect 1496 1026 1541 1036
rect 1372 998 1446 1022
rect 1314 994 1446 998
tri 1446 994 1474 1022 sw
rect 1496 1012 1498 1026
tri 1496 1010 1498 1012 ne
rect 1510 1008 1541 1026
rect 1510 998 1556 1008
rect 1623 1037 1638 1052
tri 1248 973 1260 985 ne
rect 1260 980 1270 985
tri 1270 980 1275 985 sw
rect 1159 634 1174 862
rect 1260 824 1275 980
rect 1314 938 1342 994
tri 1434 976 1452 994 ne
rect 1452 974 1474 994
tri 1474 974 1494 994 sw
tri 1510 980 1528 998 ne
rect 1333 904 1342 938
rect 1376 965 1418 966
rect 1376 931 1381 965
rect 1411 931 1418 965
rect 1376 922 1418 931
rect 1452 965 1494 974
rect 1452 931 1459 965
rect 1489 931 1494 965
rect 1452 926 1494 931
rect 1528 938 1556 998
tri 1601 985 1623 1007 se
rect 1623 1000 1638 1008
tri 1623 985 1638 1000 nw
tri 1595 979 1601 985 se
rect 1601 979 1610 985
rect 1314 894 1342 904
tri 1342 894 1366 918 sw
rect 1314 862 1356 894
tri 1373 886 1374 887 sw
rect 1373 862 1374 886
tri 1376 885 1413 922 ne
rect 1413 894 1418 922
tri 1418 894 1444 920 sw
rect 1528 904 1537 938
rect 1528 894 1556 904
rect 1413 885 1497 894
tri 1413 866 1432 885 ne
rect 1432 866 1497 885
rect 1314 840 1374 862
rect 1496 862 1497 866
rect 1514 862 1556 894
rect 1496 840 1556 862
rect 1402 824 1419 838
rect 1451 824 1468 838
tri 1239 788 1261 810 se
rect 1261 803 1276 824
tri 1261 788 1276 803 nw
rect 1595 803 1610 979
tri 1610 972 1623 985 nw
rect 1696 904 1711 1132
tri 1233 782 1239 788 se
rect 1239 782 1248 788
rect 1233 766 1248 782
tri 1248 775 1261 788 nw
rect 1402 780 1419 794
rect 1451 780 1468 794
tri 1595 788 1610 803 ne
tri 1610 788 1632 810 sw
rect 1233 730 1248 738
rect 1314 766 1374 780
rect 1329 756 1374 766
rect 1329 738 1357 756
tri 1233 715 1248 730 ne
tri 1248 715 1270 737 sw
rect 1314 728 1357 738
rect 1372 752 1374 756
rect 1496 766 1556 780
tri 1610 775 1623 788 ne
rect 1623 782 1632 788
tri 1632 782 1638 788 sw
rect 1496 756 1541 766
rect 1372 728 1446 752
rect 1314 724 1446 728
tri 1446 724 1474 752 sw
rect 1496 742 1498 756
tri 1496 740 1498 742 ne
rect 1510 738 1541 756
rect 1510 728 1556 738
rect 1623 767 1638 782
tri 1248 703 1260 715 ne
rect 1260 710 1270 715
tri 1270 710 1275 715 sw
rect 1159 364 1174 592
rect 1260 554 1275 710
rect 1314 668 1342 724
tri 1434 706 1452 724 ne
rect 1452 704 1474 724
tri 1474 704 1494 724 sw
tri 1510 710 1528 728 ne
rect 1333 634 1342 668
rect 1376 695 1418 696
rect 1376 661 1381 695
rect 1411 661 1418 695
rect 1376 652 1418 661
rect 1452 695 1494 704
rect 1452 661 1459 695
rect 1489 661 1494 695
rect 1452 656 1494 661
rect 1528 668 1556 728
tri 1601 715 1623 737 se
rect 1623 730 1638 738
tri 1623 715 1638 730 nw
tri 1595 709 1601 715 se
rect 1601 709 1610 715
rect 1314 624 1342 634
tri 1342 624 1366 648 sw
rect 1314 592 1356 624
tri 1373 616 1374 617 sw
rect 1373 592 1374 616
tri 1376 615 1413 652 ne
rect 1413 624 1418 652
tri 1418 624 1444 650 sw
rect 1528 634 1537 668
rect 1528 624 1556 634
rect 1413 615 1497 624
tri 1413 596 1432 615 ne
rect 1432 596 1497 615
rect 1314 570 1374 592
rect 1496 592 1497 596
rect 1514 592 1556 624
rect 1496 570 1556 592
rect 1402 554 1419 568
rect 1451 554 1468 568
tri 1239 518 1261 540 se
rect 1261 533 1276 554
tri 1261 518 1276 533 nw
rect 1595 533 1610 709
tri 1610 702 1623 715 nw
rect 1696 634 1711 862
tri 1233 512 1239 518 se
rect 1239 512 1248 518
rect 1233 496 1248 512
tri 1248 505 1261 518 nw
rect 1402 510 1419 524
rect 1451 510 1468 524
tri 1595 518 1610 533 ne
tri 1610 518 1632 540 sw
rect 1233 460 1248 468
rect 1314 496 1374 510
rect 1329 486 1374 496
rect 1329 468 1357 486
tri 1233 445 1248 460 ne
tri 1248 445 1270 467 sw
rect 1314 458 1357 468
rect 1372 482 1374 486
rect 1496 496 1556 510
tri 1610 505 1623 518 ne
rect 1623 512 1632 518
tri 1632 512 1638 518 sw
rect 1496 486 1541 496
rect 1372 458 1446 482
rect 1314 454 1446 458
tri 1446 454 1474 482 sw
rect 1496 472 1498 486
tri 1496 470 1498 472 ne
rect 1510 468 1541 486
rect 1510 458 1556 468
rect 1623 497 1638 512
tri 1248 433 1260 445 ne
rect 1260 440 1270 445
tri 1270 440 1275 445 sw
rect 1159 94 1174 322
rect 1260 284 1275 440
rect 1314 398 1342 454
tri 1434 436 1452 454 ne
rect 1452 434 1474 454
tri 1474 434 1494 454 sw
tri 1510 440 1528 458 ne
rect 1333 364 1342 398
rect 1376 425 1418 426
rect 1376 391 1381 425
rect 1411 391 1418 425
rect 1376 382 1418 391
rect 1452 425 1494 434
rect 1452 391 1459 425
rect 1489 391 1494 425
rect 1452 386 1494 391
rect 1528 398 1556 458
tri 1601 445 1623 467 se
rect 1623 460 1638 468
tri 1623 445 1638 460 nw
tri 1595 439 1601 445 se
rect 1601 439 1610 445
rect 1314 354 1342 364
tri 1342 354 1366 378 sw
rect 1314 322 1356 354
tri 1373 346 1374 347 sw
rect 1373 322 1374 346
tri 1376 345 1413 382 ne
rect 1413 354 1418 382
tri 1418 354 1444 380 sw
rect 1528 364 1537 398
rect 1528 354 1556 364
rect 1413 345 1497 354
tri 1413 326 1432 345 ne
rect 1432 326 1497 345
rect 1314 300 1374 322
rect 1496 322 1497 326
rect 1514 322 1556 354
rect 1496 300 1556 322
rect 1402 284 1419 298
rect 1451 284 1468 298
tri 1239 248 1261 270 se
rect 1261 263 1276 284
tri 1261 248 1276 263 nw
rect 1595 263 1610 439
tri 1610 432 1623 445 nw
rect 1696 364 1711 592
tri 1233 242 1239 248 se
rect 1239 242 1248 248
rect 1233 226 1248 242
tri 1248 235 1261 248 nw
rect 1402 240 1419 254
rect 1451 240 1468 254
tri 1595 248 1610 263 ne
tri 1610 248 1632 270 sw
rect 1233 190 1248 198
rect 1314 226 1374 240
rect 1329 216 1374 226
rect 1329 198 1357 216
tri 1233 175 1248 190 ne
tri 1248 175 1270 197 sw
rect 1314 188 1357 198
rect 1372 212 1374 216
rect 1496 226 1556 240
tri 1610 235 1623 248 ne
rect 1623 242 1632 248
tri 1632 242 1638 248 sw
rect 1496 216 1541 226
rect 1372 188 1446 212
rect 1314 184 1446 188
tri 1446 184 1474 212 sw
rect 1496 202 1498 216
tri 1496 200 1498 202 ne
rect 1510 198 1541 216
rect 1510 188 1556 198
rect 1623 227 1638 242
tri 1248 163 1260 175 ne
rect 1260 170 1270 175
tri 1270 170 1275 175 sw
rect 1159 -176 1174 52
rect 1260 14 1275 170
rect 1314 128 1342 184
tri 1434 166 1452 184 ne
rect 1452 164 1474 184
tri 1474 164 1494 184 sw
tri 1510 170 1528 188 ne
rect 1333 94 1342 128
rect 1376 155 1418 156
rect 1376 121 1381 155
rect 1411 121 1418 155
rect 1376 112 1418 121
rect 1452 155 1494 164
rect 1452 121 1459 155
rect 1489 121 1494 155
rect 1452 116 1494 121
rect 1528 128 1556 188
tri 1601 175 1623 197 se
rect 1623 190 1638 198
tri 1623 175 1638 190 nw
tri 1595 169 1601 175 se
rect 1601 169 1610 175
rect 1314 84 1342 94
tri 1342 84 1366 108 sw
rect 1314 52 1356 84
tri 1373 76 1374 77 sw
rect 1373 52 1374 76
tri 1376 75 1413 112 ne
rect 1413 84 1418 112
tri 1418 84 1444 110 sw
rect 1528 94 1537 128
rect 1528 84 1556 94
rect 1413 75 1497 84
tri 1413 56 1432 75 ne
rect 1432 56 1497 75
rect 1314 30 1374 52
rect 1496 52 1497 56
rect 1514 52 1556 84
rect 1496 30 1556 52
rect 1402 14 1419 28
rect 1451 14 1468 28
tri 1239 -22 1261 0 se
rect 1261 -7 1276 14
tri 1261 -22 1276 -7 nw
rect 1595 -7 1610 169
tri 1610 162 1623 175 nw
rect 1696 94 1711 322
tri 1233 -28 1239 -22 se
rect 1239 -28 1248 -22
rect 1233 -44 1248 -28
tri 1248 -35 1261 -22 nw
rect 1402 -30 1419 -16
rect 1451 -30 1468 -16
tri 1595 -22 1610 -7 ne
tri 1610 -22 1632 0 sw
rect 1233 -80 1248 -72
rect 1314 -44 1374 -30
rect 1329 -54 1374 -44
rect 1329 -72 1357 -54
tri 1233 -95 1248 -80 ne
tri 1248 -95 1270 -73 sw
rect 1314 -82 1357 -72
rect 1372 -58 1374 -54
rect 1496 -44 1556 -30
tri 1610 -35 1623 -22 ne
rect 1623 -28 1632 -22
tri 1632 -28 1638 -22 sw
rect 1496 -54 1541 -44
rect 1372 -82 1446 -58
rect 1314 -86 1446 -82
tri 1446 -86 1474 -58 sw
rect 1496 -68 1498 -54
tri 1496 -70 1498 -68 ne
rect 1510 -72 1541 -54
rect 1510 -82 1556 -72
rect 1623 -43 1638 -28
tri 1248 -107 1260 -95 ne
rect 1260 -100 1270 -95
tri 1270 -100 1275 -95 sw
rect 1159 -446 1174 -218
rect 1260 -256 1275 -100
rect 1314 -142 1342 -86
tri 1434 -104 1452 -86 ne
rect 1452 -106 1474 -86
tri 1474 -106 1494 -86 sw
tri 1510 -100 1528 -82 ne
rect 1333 -176 1342 -142
rect 1376 -115 1418 -114
rect 1376 -149 1381 -115
rect 1411 -149 1418 -115
rect 1376 -158 1418 -149
rect 1452 -115 1494 -106
rect 1452 -149 1459 -115
rect 1489 -149 1494 -115
rect 1452 -154 1494 -149
rect 1528 -142 1556 -82
tri 1601 -95 1623 -73 se
rect 1623 -80 1638 -72
tri 1623 -95 1638 -80 nw
tri 1595 -101 1601 -95 se
rect 1601 -101 1610 -95
rect 1314 -186 1342 -176
tri 1342 -186 1366 -162 sw
rect 1314 -218 1356 -186
tri 1373 -194 1374 -193 sw
rect 1373 -218 1374 -194
tri 1376 -195 1413 -158 ne
rect 1413 -186 1418 -158
tri 1418 -186 1444 -160 sw
rect 1528 -176 1537 -142
rect 1528 -186 1556 -176
rect 1413 -195 1497 -186
tri 1413 -214 1432 -195 ne
rect 1432 -214 1497 -195
rect 1314 -240 1374 -218
rect 1496 -218 1497 -214
rect 1514 -218 1556 -186
rect 1496 -240 1556 -218
rect 1402 -256 1419 -242
rect 1451 -256 1468 -242
tri 1239 -292 1261 -270 se
rect 1261 -277 1276 -256
tri 1261 -292 1276 -277 nw
rect 1595 -277 1610 -101
tri 1610 -108 1623 -95 nw
rect 1696 -176 1711 52
tri 1233 -298 1239 -292 se
rect 1239 -298 1248 -292
rect 1233 -314 1248 -298
tri 1248 -305 1261 -292 nw
rect 1402 -300 1419 -286
rect 1451 -300 1468 -286
tri 1595 -292 1610 -277 ne
tri 1610 -292 1632 -270 sw
rect 1233 -350 1248 -342
rect 1314 -314 1374 -300
rect 1329 -324 1374 -314
rect 1329 -342 1357 -324
tri 1233 -365 1248 -350 ne
tri 1248 -365 1270 -343 sw
rect 1314 -352 1357 -342
rect 1372 -328 1374 -324
rect 1496 -314 1556 -300
tri 1610 -305 1623 -292 ne
rect 1623 -298 1632 -292
tri 1632 -298 1638 -292 sw
rect 1496 -324 1541 -314
rect 1372 -352 1446 -328
rect 1314 -356 1446 -352
tri 1446 -356 1474 -328 sw
rect 1496 -338 1498 -324
tri 1496 -340 1498 -338 ne
rect 1510 -342 1541 -324
rect 1510 -352 1556 -342
rect 1623 -313 1638 -298
tri 1248 -377 1260 -365 ne
rect 1260 -370 1270 -365
tri 1270 -370 1275 -365 sw
rect 1159 -716 1174 -488
rect 1260 -526 1275 -370
rect 1314 -412 1342 -356
tri 1434 -374 1452 -356 ne
rect 1452 -376 1474 -356
tri 1474 -376 1494 -356 sw
tri 1510 -370 1528 -352 ne
rect 1333 -446 1342 -412
rect 1376 -385 1418 -384
rect 1376 -419 1381 -385
rect 1411 -419 1418 -385
rect 1376 -428 1418 -419
rect 1452 -385 1494 -376
rect 1452 -419 1459 -385
rect 1489 -419 1494 -385
rect 1452 -424 1494 -419
rect 1528 -412 1556 -352
tri 1601 -365 1623 -343 se
rect 1623 -350 1638 -342
tri 1623 -365 1638 -350 nw
tri 1595 -371 1601 -365 se
rect 1601 -371 1610 -365
rect 1314 -456 1342 -446
tri 1342 -456 1366 -432 sw
rect 1314 -488 1356 -456
tri 1373 -464 1374 -463 sw
rect 1373 -488 1374 -464
tri 1376 -465 1413 -428 ne
rect 1413 -456 1418 -428
tri 1418 -456 1444 -430 sw
rect 1528 -446 1537 -412
rect 1528 -456 1556 -446
rect 1413 -465 1497 -456
tri 1413 -484 1432 -465 ne
rect 1432 -484 1497 -465
rect 1314 -510 1374 -488
rect 1496 -488 1497 -484
rect 1514 -488 1556 -456
rect 1496 -510 1556 -488
rect 1402 -526 1419 -512
rect 1451 -526 1468 -512
tri 1239 -562 1261 -540 se
rect 1261 -547 1276 -526
tri 1261 -562 1276 -547 nw
rect 1595 -547 1610 -371
tri 1610 -378 1623 -365 nw
rect 1696 -446 1711 -218
tri 1233 -568 1239 -562 se
rect 1239 -568 1248 -562
rect 1233 -584 1248 -568
tri 1248 -575 1261 -562 nw
rect 1402 -570 1419 -556
rect 1451 -570 1468 -556
tri 1595 -562 1610 -547 ne
tri 1610 -562 1632 -540 sw
rect 1233 -620 1248 -612
rect 1314 -584 1374 -570
rect 1329 -594 1374 -584
rect 1329 -612 1357 -594
tri 1233 -635 1248 -620 ne
tri 1248 -635 1270 -613 sw
rect 1314 -622 1357 -612
rect 1372 -598 1374 -594
rect 1496 -584 1556 -570
tri 1610 -575 1623 -562 ne
rect 1623 -568 1632 -562
tri 1632 -568 1638 -562 sw
rect 1496 -594 1541 -584
rect 1372 -622 1446 -598
rect 1314 -626 1446 -622
tri 1446 -626 1474 -598 sw
rect 1496 -608 1498 -594
tri 1496 -610 1498 -608 ne
rect 1510 -612 1541 -594
rect 1510 -622 1556 -612
rect 1623 -583 1638 -568
tri 1248 -647 1260 -635 ne
rect 1260 -640 1270 -635
tri 1270 -640 1275 -635 sw
rect 1159 -986 1174 -758
rect 1260 -796 1275 -640
rect 1314 -682 1342 -626
tri 1434 -644 1452 -626 ne
rect 1452 -646 1474 -626
tri 1474 -646 1494 -626 sw
tri 1510 -640 1528 -622 ne
rect 1333 -716 1342 -682
rect 1376 -655 1418 -654
rect 1376 -689 1381 -655
rect 1411 -689 1418 -655
rect 1376 -698 1418 -689
rect 1452 -655 1494 -646
rect 1452 -689 1459 -655
rect 1489 -689 1494 -655
rect 1452 -694 1494 -689
rect 1528 -682 1556 -622
tri 1601 -635 1623 -613 se
rect 1623 -620 1638 -612
tri 1623 -635 1638 -620 nw
tri 1595 -641 1601 -635 se
rect 1601 -641 1610 -635
rect 1314 -726 1342 -716
tri 1342 -726 1366 -702 sw
rect 1314 -758 1356 -726
tri 1373 -734 1374 -733 sw
rect 1373 -758 1374 -734
tri 1376 -735 1413 -698 ne
rect 1413 -726 1418 -698
tri 1418 -726 1444 -700 sw
rect 1528 -716 1537 -682
rect 1528 -726 1556 -716
rect 1413 -735 1497 -726
tri 1413 -754 1432 -735 ne
rect 1432 -754 1497 -735
rect 1314 -780 1374 -758
rect 1496 -758 1497 -754
rect 1514 -758 1556 -726
rect 1496 -780 1556 -758
rect 1402 -796 1419 -782
rect 1451 -796 1468 -782
tri 1239 -832 1261 -810 se
rect 1261 -817 1276 -796
tri 1261 -832 1276 -817 nw
rect 1595 -817 1610 -641
tri 1610 -648 1623 -635 nw
rect 1696 -716 1711 -488
tri 1233 -838 1239 -832 se
rect 1239 -838 1248 -832
rect 1233 -854 1248 -838
tri 1248 -845 1261 -832 nw
rect 1402 -840 1419 -826
rect 1451 -840 1468 -826
tri 1595 -832 1610 -817 ne
tri 1610 -832 1632 -810 sw
rect 1233 -890 1248 -882
rect 1314 -854 1374 -840
rect 1329 -864 1374 -854
rect 1329 -882 1357 -864
tri 1233 -905 1248 -890 ne
tri 1248 -905 1270 -883 sw
rect 1314 -892 1357 -882
rect 1372 -868 1374 -864
rect 1496 -854 1556 -840
tri 1610 -845 1623 -832 ne
rect 1623 -838 1632 -832
tri 1632 -838 1638 -832 sw
rect 1496 -864 1541 -854
rect 1372 -892 1446 -868
rect 1314 -896 1446 -892
tri 1446 -896 1474 -868 sw
rect 1496 -878 1498 -864
tri 1496 -880 1498 -878 ne
rect 1510 -882 1541 -864
rect 1510 -892 1556 -882
rect 1623 -853 1638 -838
tri 1248 -917 1260 -905 ne
rect 1260 -910 1270 -905
tri 1270 -910 1275 -905 sw
rect 1159 -1256 1174 -1028
rect 1260 -1066 1275 -910
rect 1314 -952 1342 -896
tri 1434 -914 1452 -896 ne
rect 1452 -916 1474 -896
tri 1474 -916 1494 -896 sw
tri 1510 -910 1528 -892 ne
rect 1333 -986 1342 -952
rect 1376 -925 1418 -924
rect 1376 -959 1381 -925
rect 1411 -959 1418 -925
rect 1376 -968 1418 -959
rect 1452 -925 1494 -916
rect 1452 -959 1459 -925
rect 1489 -959 1494 -925
rect 1452 -964 1494 -959
rect 1528 -952 1556 -892
tri 1601 -905 1623 -883 se
rect 1623 -890 1638 -882
tri 1623 -905 1638 -890 nw
tri 1595 -911 1601 -905 se
rect 1601 -911 1610 -905
rect 1314 -996 1342 -986
tri 1342 -996 1366 -972 sw
rect 1314 -1028 1356 -996
tri 1373 -1004 1374 -1003 sw
rect 1373 -1028 1374 -1004
tri 1376 -1005 1413 -968 ne
rect 1413 -996 1418 -968
tri 1418 -996 1444 -970 sw
rect 1528 -986 1537 -952
rect 1528 -996 1556 -986
rect 1413 -1005 1497 -996
tri 1413 -1024 1432 -1005 ne
rect 1432 -1024 1497 -1005
rect 1314 -1050 1374 -1028
rect 1496 -1028 1497 -1024
rect 1514 -1028 1556 -996
rect 1496 -1050 1556 -1028
rect 1402 -1066 1419 -1052
rect 1451 -1066 1468 -1052
tri 1239 -1102 1261 -1080 se
rect 1261 -1087 1276 -1066
tri 1261 -1102 1276 -1087 nw
rect 1595 -1087 1610 -911
tri 1610 -918 1623 -905 nw
rect 1696 -986 1711 -758
tri 1233 -1108 1239 -1102 se
rect 1239 -1108 1248 -1102
rect 1233 -1124 1248 -1108
tri 1248 -1115 1261 -1102 nw
rect 1402 -1110 1419 -1096
rect 1451 -1110 1468 -1096
tri 1595 -1102 1610 -1087 ne
tri 1610 -1102 1632 -1080 sw
rect 1233 -1160 1248 -1152
rect 1314 -1124 1374 -1110
rect 1329 -1134 1374 -1124
rect 1329 -1152 1357 -1134
tri 1233 -1175 1248 -1160 ne
tri 1248 -1175 1270 -1153 sw
rect 1314 -1162 1357 -1152
rect 1372 -1138 1374 -1134
rect 1496 -1124 1556 -1110
tri 1610 -1115 1623 -1102 ne
rect 1623 -1108 1632 -1102
tri 1632 -1108 1638 -1102 sw
rect 1496 -1134 1541 -1124
rect 1372 -1162 1446 -1138
rect 1314 -1166 1446 -1162
tri 1446 -1166 1474 -1138 sw
rect 1496 -1148 1498 -1134
tri 1496 -1150 1498 -1148 ne
rect 1510 -1152 1541 -1134
rect 1510 -1162 1556 -1152
rect 1623 -1123 1638 -1108
tri 1248 -1187 1260 -1175 ne
rect 1260 -1180 1270 -1175
tri 1270 -1180 1275 -1175 sw
rect 1159 -1526 1174 -1298
rect 1260 -1336 1275 -1180
rect 1314 -1222 1342 -1166
tri 1434 -1184 1452 -1166 ne
rect 1452 -1186 1474 -1166
tri 1474 -1186 1494 -1166 sw
tri 1510 -1180 1528 -1162 ne
rect 1333 -1256 1342 -1222
rect 1376 -1195 1418 -1194
rect 1376 -1229 1381 -1195
rect 1411 -1229 1418 -1195
rect 1376 -1238 1418 -1229
rect 1452 -1195 1494 -1186
rect 1452 -1229 1459 -1195
rect 1489 -1229 1494 -1195
rect 1452 -1234 1494 -1229
rect 1528 -1222 1556 -1162
tri 1601 -1175 1623 -1153 se
rect 1623 -1160 1638 -1152
tri 1623 -1175 1638 -1160 nw
tri 1595 -1181 1601 -1175 se
rect 1601 -1181 1610 -1175
rect 1314 -1266 1342 -1256
tri 1342 -1266 1366 -1242 sw
rect 1314 -1298 1356 -1266
tri 1373 -1274 1374 -1273 sw
rect 1373 -1298 1374 -1274
tri 1376 -1275 1413 -1238 ne
rect 1413 -1266 1418 -1238
tri 1418 -1266 1444 -1240 sw
rect 1528 -1256 1537 -1222
rect 1528 -1266 1556 -1256
rect 1413 -1275 1497 -1266
tri 1413 -1294 1432 -1275 ne
rect 1432 -1294 1497 -1275
rect 1314 -1320 1374 -1298
rect 1496 -1298 1497 -1294
rect 1514 -1298 1556 -1266
rect 1496 -1320 1556 -1298
rect 1402 -1336 1419 -1322
rect 1451 -1336 1468 -1322
tri 1239 -1372 1261 -1350 se
rect 1261 -1357 1276 -1336
tri 1261 -1372 1276 -1357 nw
rect 1595 -1357 1610 -1181
tri 1610 -1188 1623 -1175 nw
rect 1696 -1256 1711 -1028
tri 1233 -1378 1239 -1372 se
rect 1239 -1378 1248 -1372
rect 1233 -1394 1248 -1378
tri 1248 -1385 1261 -1372 nw
rect 1402 -1380 1419 -1366
rect 1451 -1380 1468 -1366
tri 1595 -1372 1610 -1357 ne
tri 1610 -1372 1632 -1350 sw
rect 1233 -1430 1248 -1422
rect 1314 -1394 1374 -1380
rect 1329 -1404 1374 -1394
rect 1329 -1422 1357 -1404
tri 1233 -1445 1248 -1430 ne
tri 1248 -1445 1270 -1423 sw
rect 1314 -1432 1357 -1422
rect 1372 -1408 1374 -1404
rect 1496 -1394 1556 -1380
tri 1610 -1385 1623 -1372 ne
rect 1623 -1378 1632 -1372
tri 1632 -1378 1638 -1372 sw
rect 1496 -1404 1541 -1394
rect 1372 -1432 1446 -1408
rect 1314 -1436 1446 -1432
tri 1446 -1436 1474 -1408 sw
rect 1496 -1418 1498 -1404
tri 1496 -1420 1498 -1418 ne
rect 1510 -1422 1541 -1404
rect 1510 -1432 1556 -1422
rect 1623 -1393 1638 -1378
tri 1248 -1457 1260 -1445 ne
rect 1260 -1450 1270 -1445
tri 1270 -1450 1275 -1445 sw
rect 1159 -1796 1174 -1568
rect 1260 -1606 1275 -1450
rect 1314 -1492 1342 -1436
tri 1434 -1454 1452 -1436 ne
rect 1452 -1456 1474 -1436
tri 1474 -1456 1494 -1436 sw
tri 1510 -1450 1528 -1432 ne
rect 1333 -1526 1342 -1492
rect 1376 -1465 1418 -1464
rect 1376 -1499 1381 -1465
rect 1411 -1499 1418 -1465
rect 1376 -1508 1418 -1499
rect 1452 -1465 1494 -1456
rect 1452 -1499 1459 -1465
rect 1489 -1499 1494 -1465
rect 1452 -1504 1494 -1499
rect 1528 -1492 1556 -1432
tri 1601 -1445 1623 -1423 se
rect 1623 -1430 1638 -1422
tri 1623 -1445 1638 -1430 nw
tri 1595 -1451 1601 -1445 se
rect 1601 -1451 1610 -1445
rect 1314 -1536 1342 -1526
tri 1342 -1536 1366 -1512 sw
rect 1314 -1568 1356 -1536
tri 1373 -1544 1374 -1543 sw
rect 1373 -1568 1374 -1544
tri 1376 -1545 1413 -1508 ne
rect 1413 -1536 1418 -1508
tri 1418 -1536 1444 -1510 sw
rect 1528 -1526 1537 -1492
rect 1528 -1536 1556 -1526
rect 1413 -1545 1497 -1536
tri 1413 -1564 1432 -1545 ne
rect 1432 -1564 1497 -1545
rect 1314 -1590 1374 -1568
rect 1496 -1568 1497 -1564
rect 1514 -1568 1556 -1536
rect 1496 -1590 1556 -1568
rect 1402 -1606 1419 -1592
rect 1451 -1606 1468 -1592
tri 1239 -1642 1261 -1620 se
rect 1261 -1627 1276 -1606
tri 1261 -1642 1276 -1627 nw
rect 1595 -1627 1610 -1451
tri 1610 -1458 1623 -1445 nw
rect 1696 -1526 1711 -1298
tri 1233 -1648 1239 -1642 se
rect 1239 -1648 1248 -1642
rect 1233 -1664 1248 -1648
tri 1248 -1655 1261 -1642 nw
rect 1402 -1650 1419 -1636
rect 1451 -1650 1468 -1636
tri 1595 -1642 1610 -1627 ne
tri 1610 -1642 1632 -1620 sw
rect 1233 -1700 1248 -1692
rect 1314 -1664 1374 -1650
rect 1329 -1674 1374 -1664
rect 1329 -1692 1357 -1674
tri 1233 -1715 1248 -1700 ne
tri 1248 -1715 1270 -1693 sw
rect 1314 -1702 1357 -1692
rect 1372 -1678 1374 -1674
rect 1496 -1664 1556 -1650
tri 1610 -1655 1623 -1642 ne
rect 1623 -1648 1632 -1642
tri 1632 -1648 1638 -1642 sw
rect 1496 -1674 1541 -1664
rect 1372 -1702 1446 -1678
rect 1314 -1706 1446 -1702
tri 1446 -1706 1474 -1678 sw
rect 1496 -1688 1498 -1674
tri 1496 -1690 1498 -1688 ne
rect 1510 -1692 1541 -1674
rect 1510 -1702 1556 -1692
rect 1623 -1663 1638 -1648
tri 1248 -1727 1260 -1715 ne
rect 1260 -1720 1270 -1715
tri 1270 -1720 1275 -1715 sw
rect 1159 -2066 1174 -1838
rect 1260 -1876 1275 -1720
rect 1314 -1762 1342 -1706
tri 1434 -1724 1452 -1706 ne
rect 1452 -1726 1474 -1706
tri 1474 -1726 1494 -1706 sw
tri 1510 -1720 1528 -1702 ne
rect 1333 -1796 1342 -1762
rect 1376 -1735 1418 -1734
rect 1376 -1769 1381 -1735
rect 1411 -1769 1418 -1735
rect 1376 -1778 1418 -1769
rect 1452 -1735 1494 -1726
rect 1452 -1769 1459 -1735
rect 1489 -1769 1494 -1735
rect 1452 -1774 1494 -1769
rect 1528 -1762 1556 -1702
tri 1601 -1715 1623 -1693 se
rect 1623 -1700 1638 -1692
tri 1623 -1715 1638 -1700 nw
tri 1595 -1721 1601 -1715 se
rect 1601 -1721 1610 -1715
rect 1314 -1806 1342 -1796
tri 1342 -1806 1366 -1782 sw
rect 1314 -1838 1356 -1806
tri 1373 -1814 1374 -1813 sw
rect 1373 -1838 1374 -1814
tri 1376 -1815 1413 -1778 ne
rect 1413 -1806 1418 -1778
tri 1418 -1806 1444 -1780 sw
rect 1528 -1796 1537 -1762
rect 1528 -1806 1556 -1796
rect 1413 -1815 1497 -1806
tri 1413 -1834 1432 -1815 ne
rect 1432 -1834 1497 -1815
rect 1314 -1860 1374 -1838
rect 1496 -1838 1497 -1834
rect 1514 -1838 1556 -1806
rect 1496 -1860 1556 -1838
rect 1402 -1876 1419 -1862
rect 1451 -1876 1468 -1862
tri 1239 -1912 1261 -1890 se
rect 1261 -1897 1276 -1876
tri 1261 -1912 1276 -1897 nw
rect 1595 -1897 1610 -1721
tri 1610 -1728 1623 -1715 nw
rect 1696 -1796 1711 -1568
tri 1233 -1918 1239 -1912 se
rect 1239 -1918 1248 -1912
rect 1233 -1934 1248 -1918
tri 1248 -1925 1261 -1912 nw
rect 1402 -1920 1419 -1906
rect 1451 -1920 1468 -1906
tri 1595 -1912 1610 -1897 ne
tri 1610 -1912 1632 -1890 sw
rect 1233 -1970 1248 -1962
rect 1314 -1934 1374 -1920
rect 1329 -1944 1374 -1934
rect 1329 -1962 1357 -1944
tri 1233 -1985 1248 -1970 ne
tri 1248 -1985 1270 -1963 sw
rect 1314 -1972 1357 -1962
rect 1372 -1948 1374 -1944
rect 1496 -1934 1556 -1920
tri 1610 -1925 1623 -1912 ne
rect 1623 -1918 1632 -1912
tri 1632 -1918 1638 -1912 sw
rect 1496 -1944 1541 -1934
rect 1372 -1972 1446 -1948
rect 1314 -1976 1446 -1972
tri 1446 -1976 1474 -1948 sw
rect 1496 -1958 1498 -1944
tri 1496 -1960 1498 -1958 ne
rect 1510 -1962 1541 -1944
rect 1510 -1972 1556 -1962
rect 1623 -1933 1638 -1918
tri 1248 -1997 1260 -1985 ne
rect 1260 -1990 1270 -1985
tri 1270 -1990 1275 -1985 sw
rect 1159 -2146 1174 -2108
rect 1260 -2146 1275 -1990
rect 1314 -2032 1342 -1976
tri 1434 -1994 1452 -1976 ne
rect 1452 -1996 1474 -1976
tri 1474 -1996 1494 -1976 sw
tri 1510 -1990 1528 -1972 ne
rect 1333 -2066 1342 -2032
rect 1376 -2005 1418 -2004
rect 1376 -2039 1381 -2005
rect 1411 -2039 1418 -2005
rect 1376 -2048 1418 -2039
rect 1452 -2005 1494 -1996
rect 1452 -2039 1459 -2005
rect 1489 -2039 1494 -2005
rect 1452 -2044 1494 -2039
rect 1528 -2032 1556 -1972
tri 1601 -1985 1623 -1963 se
rect 1623 -1970 1638 -1962
tri 1623 -1985 1638 -1970 nw
tri 1595 -1991 1601 -1985 se
rect 1601 -1991 1610 -1985
rect 1314 -2076 1342 -2066
tri 1342 -2076 1366 -2052 sw
rect 1314 -2108 1356 -2076
tri 1373 -2084 1374 -2083 sw
rect 1373 -2108 1374 -2084
tri 1376 -2085 1413 -2048 ne
rect 1413 -2076 1418 -2048
tri 1418 -2076 1444 -2050 sw
rect 1528 -2066 1537 -2032
rect 1528 -2076 1556 -2066
rect 1413 -2085 1497 -2076
tri 1413 -2104 1432 -2085 ne
rect 1432 -2104 1497 -2085
rect 1314 -2130 1374 -2108
rect 1496 -2108 1497 -2104
rect 1514 -2108 1556 -2076
rect 1496 -2130 1556 -2108
rect 1402 -2146 1419 -2132
rect 1451 -2146 1468 -2132
rect 1595 -2146 1610 -1991
tri 1610 -1998 1623 -1985 nw
rect 1696 -2066 1711 -1838
rect 1696 -2146 1711 -2108
rect 1739 1984 1754 2174
tri 1819 2138 1841 2160 se
rect 1841 2153 1856 2174
tri 1841 2138 1856 2153 nw
rect 2175 2153 2190 2174
tri 1813 2132 1819 2138 se
rect 1819 2132 1828 2138
rect 1813 2116 1828 2132
tri 1828 2125 1841 2138 nw
rect 1982 2130 1999 2144
rect 2031 2130 2048 2144
tri 2175 2138 2190 2153 ne
tri 2190 2138 2212 2160 sw
rect 1813 2080 1828 2088
rect 1894 2116 1954 2130
rect 1909 2106 1954 2116
rect 1909 2088 1937 2106
tri 1813 2065 1828 2080 ne
tri 1828 2065 1850 2087 sw
rect 1894 2078 1937 2088
rect 1952 2102 1954 2106
rect 2076 2116 2136 2130
tri 2190 2125 2203 2138 ne
rect 2203 2132 2212 2138
tri 2212 2132 2218 2138 sw
rect 2076 2106 2121 2116
rect 1952 2078 2026 2102
rect 1894 2074 2026 2078
tri 2026 2074 2054 2102 sw
rect 2076 2092 2078 2106
tri 2076 2090 2078 2092 ne
rect 2090 2088 2121 2106
rect 2090 2078 2136 2088
rect 2203 2117 2218 2132
tri 1828 2053 1840 2065 ne
rect 1840 2060 1850 2065
tri 1850 2060 1855 2065 sw
rect 1739 1714 1754 1942
rect 1840 1904 1855 2060
rect 1894 2018 1922 2074
tri 2014 2056 2032 2074 ne
rect 2032 2054 2054 2074
tri 2054 2054 2074 2074 sw
tri 2090 2060 2108 2078 ne
rect 1913 1984 1922 2018
rect 1956 2045 1998 2046
rect 1956 2011 1961 2045
rect 1991 2011 1998 2045
rect 1956 2002 1998 2011
rect 2032 2045 2074 2054
rect 2032 2011 2039 2045
rect 2069 2011 2074 2045
rect 2032 2006 2074 2011
rect 2108 2018 2136 2078
tri 2181 2065 2203 2087 se
rect 2203 2080 2218 2088
tri 2203 2065 2218 2080 nw
tri 2175 2059 2181 2065 se
rect 2181 2059 2190 2065
rect 1894 1974 1922 1984
tri 1922 1974 1946 1998 sw
rect 1894 1942 1936 1974
tri 1953 1966 1954 1967 sw
rect 1953 1942 1954 1966
tri 1956 1965 1993 2002 ne
rect 1993 1974 1998 2002
tri 1998 1974 2024 2000 sw
rect 2108 1984 2117 2018
rect 2108 1974 2136 1984
rect 1993 1965 2077 1974
tri 1993 1946 2012 1965 ne
rect 2012 1946 2077 1965
rect 1894 1920 1954 1942
rect 2076 1942 2077 1946
rect 2094 1942 2136 1974
rect 2076 1920 2136 1942
rect 1982 1904 1999 1918
rect 2031 1904 2048 1918
tri 1819 1868 1841 1890 se
rect 1841 1883 1856 1904
tri 1841 1868 1856 1883 nw
rect 2175 1883 2190 2059
tri 2190 2052 2203 2065 nw
rect 2276 1984 2291 2174
tri 1813 1862 1819 1868 se
rect 1819 1862 1828 1868
rect 1813 1846 1828 1862
tri 1828 1855 1841 1868 nw
rect 1982 1860 1999 1874
rect 2031 1860 2048 1874
tri 2175 1868 2190 1883 ne
tri 2190 1868 2212 1890 sw
rect 1813 1810 1828 1818
rect 1894 1846 1954 1860
rect 1909 1836 1954 1846
rect 1909 1818 1937 1836
tri 1813 1795 1828 1810 ne
tri 1828 1795 1850 1817 sw
rect 1894 1808 1937 1818
rect 1952 1832 1954 1836
rect 2076 1846 2136 1860
tri 2190 1855 2203 1868 ne
rect 2203 1862 2212 1868
tri 2212 1862 2218 1868 sw
rect 2076 1836 2121 1846
rect 1952 1808 2026 1832
rect 1894 1804 2026 1808
tri 2026 1804 2054 1832 sw
rect 2076 1822 2078 1836
tri 2076 1820 2078 1822 ne
rect 2090 1818 2121 1836
rect 2090 1808 2136 1818
rect 2203 1847 2218 1862
tri 1828 1783 1840 1795 ne
rect 1840 1790 1850 1795
tri 1850 1790 1855 1795 sw
rect 1739 1444 1754 1672
rect 1840 1634 1855 1790
rect 1894 1748 1922 1804
tri 2014 1786 2032 1804 ne
rect 2032 1784 2054 1804
tri 2054 1784 2074 1804 sw
tri 2090 1790 2108 1808 ne
rect 1913 1714 1922 1748
rect 1956 1775 1998 1776
rect 1956 1741 1961 1775
rect 1991 1741 1998 1775
rect 1956 1732 1998 1741
rect 2032 1775 2074 1784
rect 2032 1741 2039 1775
rect 2069 1741 2074 1775
rect 2032 1736 2074 1741
rect 2108 1748 2136 1808
tri 2181 1795 2203 1817 se
rect 2203 1810 2218 1818
tri 2203 1795 2218 1810 nw
tri 2175 1789 2181 1795 se
rect 2181 1789 2190 1795
rect 1894 1704 1922 1714
tri 1922 1704 1946 1728 sw
rect 1894 1672 1936 1704
tri 1953 1696 1954 1697 sw
rect 1953 1672 1954 1696
tri 1956 1695 1993 1732 ne
rect 1993 1704 1998 1732
tri 1998 1704 2024 1730 sw
rect 2108 1714 2117 1748
rect 2108 1704 2136 1714
rect 1993 1695 2077 1704
tri 1993 1676 2012 1695 ne
rect 2012 1676 2077 1695
rect 1894 1650 1954 1672
rect 2076 1672 2077 1676
rect 2094 1672 2136 1704
rect 2076 1650 2136 1672
rect 1982 1634 1999 1648
rect 2031 1634 2048 1648
tri 1819 1598 1841 1620 se
rect 1841 1613 1856 1634
tri 1841 1598 1856 1613 nw
rect 2175 1613 2190 1789
tri 2190 1782 2203 1795 nw
rect 2276 1714 2291 1942
tri 1813 1592 1819 1598 se
rect 1819 1592 1828 1598
rect 1813 1576 1828 1592
tri 1828 1585 1841 1598 nw
rect 1982 1590 1999 1604
rect 2031 1590 2048 1604
tri 2175 1598 2190 1613 ne
tri 2190 1598 2212 1620 sw
rect 1813 1540 1828 1548
rect 1894 1576 1954 1590
rect 1909 1566 1954 1576
rect 1909 1548 1937 1566
tri 1813 1525 1828 1540 ne
tri 1828 1525 1850 1547 sw
rect 1894 1538 1937 1548
rect 1952 1562 1954 1566
rect 2076 1576 2136 1590
tri 2190 1585 2203 1598 ne
rect 2203 1592 2212 1598
tri 2212 1592 2218 1598 sw
rect 2076 1566 2121 1576
rect 1952 1538 2026 1562
rect 1894 1534 2026 1538
tri 2026 1534 2054 1562 sw
rect 2076 1552 2078 1566
tri 2076 1550 2078 1552 ne
rect 2090 1548 2121 1566
rect 2090 1538 2136 1548
rect 2203 1577 2218 1592
tri 1828 1513 1840 1525 ne
rect 1840 1520 1850 1525
tri 1850 1520 1855 1525 sw
rect 1739 1174 1754 1402
rect 1840 1364 1855 1520
rect 1894 1478 1922 1534
tri 2014 1516 2032 1534 ne
rect 2032 1514 2054 1534
tri 2054 1514 2074 1534 sw
tri 2090 1520 2108 1538 ne
rect 1913 1444 1922 1478
rect 1956 1505 1998 1506
rect 1956 1471 1961 1505
rect 1991 1471 1998 1505
rect 1956 1462 1998 1471
rect 2032 1505 2074 1514
rect 2032 1471 2039 1505
rect 2069 1471 2074 1505
rect 2032 1466 2074 1471
rect 2108 1478 2136 1538
tri 2181 1525 2203 1547 se
rect 2203 1540 2218 1548
tri 2203 1525 2218 1540 nw
tri 2175 1519 2181 1525 se
rect 2181 1519 2190 1525
rect 1894 1434 1922 1444
tri 1922 1434 1946 1458 sw
rect 1894 1402 1936 1434
tri 1953 1426 1954 1427 sw
rect 1953 1402 1954 1426
tri 1956 1425 1993 1462 ne
rect 1993 1434 1998 1462
tri 1998 1434 2024 1460 sw
rect 2108 1444 2117 1478
rect 2108 1434 2136 1444
rect 1993 1425 2077 1434
tri 1993 1406 2012 1425 ne
rect 2012 1406 2077 1425
rect 1894 1380 1954 1402
rect 2076 1402 2077 1406
rect 2094 1402 2136 1434
rect 2076 1380 2136 1402
rect 1982 1364 1999 1378
rect 2031 1364 2048 1378
tri 1819 1328 1841 1350 se
rect 1841 1343 1856 1364
tri 1841 1328 1856 1343 nw
rect 2175 1343 2190 1519
tri 2190 1512 2203 1525 nw
rect 2276 1444 2291 1672
tri 1813 1322 1819 1328 se
rect 1819 1322 1828 1328
rect 1813 1306 1828 1322
tri 1828 1315 1841 1328 nw
rect 1982 1320 1999 1334
rect 2031 1320 2048 1334
tri 2175 1328 2190 1343 ne
tri 2190 1328 2212 1350 sw
rect 1813 1270 1828 1278
rect 1894 1306 1954 1320
rect 1909 1296 1954 1306
rect 1909 1278 1937 1296
tri 1813 1255 1828 1270 ne
tri 1828 1255 1850 1277 sw
rect 1894 1268 1937 1278
rect 1952 1292 1954 1296
rect 2076 1306 2136 1320
tri 2190 1315 2203 1328 ne
rect 2203 1322 2212 1328
tri 2212 1322 2218 1328 sw
rect 2076 1296 2121 1306
rect 1952 1268 2026 1292
rect 1894 1264 2026 1268
tri 2026 1264 2054 1292 sw
rect 2076 1282 2078 1296
tri 2076 1280 2078 1282 ne
rect 2090 1278 2121 1296
rect 2090 1268 2136 1278
rect 2203 1307 2218 1322
tri 1828 1243 1840 1255 ne
rect 1840 1250 1850 1255
tri 1850 1250 1855 1255 sw
rect 1739 904 1754 1132
rect 1840 1094 1855 1250
rect 1894 1208 1922 1264
tri 2014 1246 2032 1264 ne
rect 2032 1244 2054 1264
tri 2054 1244 2074 1264 sw
tri 2090 1250 2108 1268 ne
rect 1913 1174 1922 1208
rect 1956 1235 1998 1236
rect 1956 1201 1961 1235
rect 1991 1201 1998 1235
rect 1956 1192 1998 1201
rect 2032 1235 2074 1244
rect 2032 1201 2039 1235
rect 2069 1201 2074 1235
rect 2032 1196 2074 1201
rect 2108 1208 2136 1268
tri 2181 1255 2203 1277 se
rect 2203 1270 2218 1278
tri 2203 1255 2218 1270 nw
tri 2175 1249 2181 1255 se
rect 2181 1249 2190 1255
rect 1894 1164 1922 1174
tri 1922 1164 1946 1188 sw
rect 1894 1132 1936 1164
tri 1953 1156 1954 1157 sw
rect 1953 1132 1954 1156
tri 1956 1155 1993 1192 ne
rect 1993 1164 1998 1192
tri 1998 1164 2024 1190 sw
rect 2108 1174 2117 1208
rect 2108 1164 2136 1174
rect 1993 1155 2077 1164
tri 1993 1136 2012 1155 ne
rect 2012 1136 2077 1155
rect 1894 1110 1954 1132
rect 2076 1132 2077 1136
rect 2094 1132 2136 1164
rect 2076 1110 2136 1132
rect 1982 1094 1999 1108
rect 2031 1094 2048 1108
tri 1819 1058 1841 1080 se
rect 1841 1073 1856 1094
tri 1841 1058 1856 1073 nw
rect 2175 1073 2190 1249
tri 2190 1242 2203 1255 nw
rect 2276 1174 2291 1402
tri 1813 1052 1819 1058 se
rect 1819 1052 1828 1058
rect 1813 1036 1828 1052
tri 1828 1045 1841 1058 nw
rect 1982 1050 1999 1064
rect 2031 1050 2048 1064
tri 2175 1058 2190 1073 ne
tri 2190 1058 2212 1080 sw
rect 1813 1000 1828 1008
rect 1894 1036 1954 1050
rect 1909 1026 1954 1036
rect 1909 1008 1937 1026
tri 1813 985 1828 1000 ne
tri 1828 985 1850 1007 sw
rect 1894 998 1937 1008
rect 1952 1022 1954 1026
rect 2076 1036 2136 1050
tri 2190 1045 2203 1058 ne
rect 2203 1052 2212 1058
tri 2212 1052 2218 1058 sw
rect 2076 1026 2121 1036
rect 1952 998 2026 1022
rect 1894 994 2026 998
tri 2026 994 2054 1022 sw
rect 2076 1012 2078 1026
tri 2076 1010 2078 1012 ne
rect 2090 1008 2121 1026
rect 2090 998 2136 1008
rect 2203 1037 2218 1052
tri 1828 973 1840 985 ne
rect 1840 980 1850 985
tri 1850 980 1855 985 sw
rect 1739 634 1754 862
rect 1840 824 1855 980
rect 1894 938 1922 994
tri 2014 976 2032 994 ne
rect 2032 974 2054 994
tri 2054 974 2074 994 sw
tri 2090 980 2108 998 ne
rect 1913 904 1922 938
rect 1956 965 1998 966
rect 1956 931 1961 965
rect 1991 931 1998 965
rect 1956 922 1998 931
rect 2032 965 2074 974
rect 2032 931 2039 965
rect 2069 931 2074 965
rect 2032 926 2074 931
rect 2108 938 2136 998
tri 2181 985 2203 1007 se
rect 2203 1000 2218 1008
tri 2203 985 2218 1000 nw
tri 2175 979 2181 985 se
rect 2181 979 2190 985
rect 1894 894 1922 904
tri 1922 894 1946 918 sw
rect 1894 862 1936 894
tri 1953 886 1954 887 sw
rect 1953 862 1954 886
tri 1956 885 1993 922 ne
rect 1993 894 1998 922
tri 1998 894 2024 920 sw
rect 2108 904 2117 938
rect 2108 894 2136 904
rect 1993 885 2077 894
tri 1993 866 2012 885 ne
rect 2012 866 2077 885
rect 1894 840 1954 862
rect 2076 862 2077 866
rect 2094 862 2136 894
rect 2076 840 2136 862
rect 1982 824 1999 838
rect 2031 824 2048 838
tri 1819 788 1841 810 se
rect 1841 803 1856 824
tri 1841 788 1856 803 nw
rect 2175 803 2190 979
tri 2190 972 2203 985 nw
rect 2276 904 2291 1132
tri 1813 782 1819 788 se
rect 1819 782 1828 788
rect 1813 766 1828 782
tri 1828 775 1841 788 nw
rect 1982 780 1999 794
rect 2031 780 2048 794
tri 2175 788 2190 803 ne
tri 2190 788 2212 810 sw
rect 1813 730 1828 738
rect 1894 766 1954 780
rect 1909 756 1954 766
rect 1909 738 1937 756
tri 1813 715 1828 730 ne
tri 1828 715 1850 737 sw
rect 1894 728 1937 738
rect 1952 752 1954 756
rect 2076 766 2136 780
tri 2190 775 2203 788 ne
rect 2203 782 2212 788
tri 2212 782 2218 788 sw
rect 2076 756 2121 766
rect 1952 728 2026 752
rect 1894 724 2026 728
tri 2026 724 2054 752 sw
rect 2076 742 2078 756
tri 2076 740 2078 742 ne
rect 2090 738 2121 756
rect 2090 728 2136 738
rect 2203 767 2218 782
tri 1828 703 1840 715 ne
rect 1840 710 1850 715
tri 1850 710 1855 715 sw
rect 1739 364 1754 592
rect 1840 554 1855 710
rect 1894 668 1922 724
tri 2014 706 2032 724 ne
rect 2032 704 2054 724
tri 2054 704 2074 724 sw
tri 2090 710 2108 728 ne
rect 1913 634 1922 668
rect 1956 695 1998 696
rect 1956 661 1961 695
rect 1991 661 1998 695
rect 1956 652 1998 661
rect 2032 695 2074 704
rect 2032 661 2039 695
rect 2069 661 2074 695
rect 2032 656 2074 661
rect 2108 668 2136 728
tri 2181 715 2203 737 se
rect 2203 730 2218 738
tri 2203 715 2218 730 nw
tri 2175 709 2181 715 se
rect 2181 709 2190 715
rect 1894 624 1922 634
tri 1922 624 1946 648 sw
rect 1894 592 1936 624
tri 1953 616 1954 617 sw
rect 1953 592 1954 616
tri 1956 615 1993 652 ne
rect 1993 624 1998 652
tri 1998 624 2024 650 sw
rect 2108 634 2117 668
rect 2108 624 2136 634
rect 1993 615 2077 624
tri 1993 596 2012 615 ne
rect 2012 596 2077 615
rect 1894 570 1954 592
rect 2076 592 2077 596
rect 2094 592 2136 624
rect 2076 570 2136 592
rect 1982 554 1999 568
rect 2031 554 2048 568
tri 1819 518 1841 540 se
rect 1841 533 1856 554
tri 1841 518 1856 533 nw
rect 2175 533 2190 709
tri 2190 702 2203 715 nw
rect 2276 634 2291 862
tri 1813 512 1819 518 se
rect 1819 512 1828 518
rect 1813 496 1828 512
tri 1828 505 1841 518 nw
rect 1982 510 1999 524
rect 2031 510 2048 524
tri 2175 518 2190 533 ne
tri 2190 518 2212 540 sw
rect 1813 460 1828 468
rect 1894 496 1954 510
rect 1909 486 1954 496
rect 1909 468 1937 486
tri 1813 445 1828 460 ne
tri 1828 445 1850 467 sw
rect 1894 458 1937 468
rect 1952 482 1954 486
rect 2076 496 2136 510
tri 2190 505 2203 518 ne
rect 2203 512 2212 518
tri 2212 512 2218 518 sw
rect 2076 486 2121 496
rect 1952 458 2026 482
rect 1894 454 2026 458
tri 2026 454 2054 482 sw
rect 2076 472 2078 486
tri 2076 470 2078 472 ne
rect 2090 468 2121 486
rect 2090 458 2136 468
rect 2203 497 2218 512
tri 1828 433 1840 445 ne
rect 1840 440 1850 445
tri 1850 440 1855 445 sw
rect 1739 94 1754 322
rect 1840 284 1855 440
rect 1894 398 1922 454
tri 2014 436 2032 454 ne
rect 2032 434 2054 454
tri 2054 434 2074 454 sw
tri 2090 440 2108 458 ne
rect 1913 364 1922 398
rect 1956 425 1998 426
rect 1956 391 1961 425
rect 1991 391 1998 425
rect 1956 382 1998 391
rect 2032 425 2074 434
rect 2032 391 2039 425
rect 2069 391 2074 425
rect 2032 386 2074 391
rect 2108 398 2136 458
tri 2181 445 2203 467 se
rect 2203 460 2218 468
tri 2203 445 2218 460 nw
tri 2175 439 2181 445 se
rect 2181 439 2190 445
rect 1894 354 1922 364
tri 1922 354 1946 378 sw
rect 1894 322 1936 354
tri 1953 346 1954 347 sw
rect 1953 322 1954 346
tri 1956 345 1993 382 ne
rect 1993 354 1998 382
tri 1998 354 2024 380 sw
rect 2108 364 2117 398
rect 2108 354 2136 364
rect 1993 345 2077 354
tri 1993 326 2012 345 ne
rect 2012 326 2077 345
rect 1894 300 1954 322
rect 2076 322 2077 326
rect 2094 322 2136 354
rect 2076 300 2136 322
rect 1982 284 1999 298
rect 2031 284 2048 298
tri 1819 248 1841 270 se
rect 1841 263 1856 284
tri 1841 248 1856 263 nw
rect 2175 263 2190 439
tri 2190 432 2203 445 nw
rect 2276 364 2291 592
tri 1813 242 1819 248 se
rect 1819 242 1828 248
rect 1813 226 1828 242
tri 1828 235 1841 248 nw
rect 1982 240 1999 254
rect 2031 240 2048 254
tri 2175 248 2190 263 ne
tri 2190 248 2212 270 sw
rect 1813 190 1828 198
rect 1894 226 1954 240
rect 1909 216 1954 226
rect 1909 198 1937 216
tri 1813 175 1828 190 ne
tri 1828 175 1850 197 sw
rect 1894 188 1937 198
rect 1952 212 1954 216
rect 2076 226 2136 240
tri 2190 235 2203 248 ne
rect 2203 242 2212 248
tri 2212 242 2218 248 sw
rect 2076 216 2121 226
rect 1952 188 2026 212
rect 1894 184 2026 188
tri 2026 184 2054 212 sw
rect 2076 202 2078 216
tri 2076 200 2078 202 ne
rect 2090 198 2121 216
rect 2090 188 2136 198
rect 2203 227 2218 242
tri 1828 163 1840 175 ne
rect 1840 170 1850 175
tri 1850 170 1855 175 sw
rect 1739 -176 1754 52
rect 1840 14 1855 170
rect 1894 128 1922 184
tri 2014 166 2032 184 ne
rect 2032 164 2054 184
tri 2054 164 2074 184 sw
tri 2090 170 2108 188 ne
rect 1913 94 1922 128
rect 1956 155 1998 156
rect 1956 121 1961 155
rect 1991 121 1998 155
rect 1956 112 1998 121
rect 2032 155 2074 164
rect 2032 121 2039 155
rect 2069 121 2074 155
rect 2032 116 2074 121
rect 2108 128 2136 188
tri 2181 175 2203 197 se
rect 2203 190 2218 198
tri 2203 175 2218 190 nw
tri 2175 169 2181 175 se
rect 2181 169 2190 175
rect 1894 84 1922 94
tri 1922 84 1946 108 sw
rect 1894 52 1936 84
tri 1953 76 1954 77 sw
rect 1953 52 1954 76
tri 1956 75 1993 112 ne
rect 1993 84 1998 112
tri 1998 84 2024 110 sw
rect 2108 94 2117 128
rect 2108 84 2136 94
rect 1993 75 2077 84
tri 1993 56 2012 75 ne
rect 2012 56 2077 75
rect 1894 30 1954 52
rect 2076 52 2077 56
rect 2094 52 2136 84
rect 2076 30 2136 52
rect 1982 14 1999 28
rect 2031 14 2048 28
tri 1819 -22 1841 0 se
rect 1841 -7 1856 14
tri 1841 -22 1856 -7 nw
rect 2175 -7 2190 169
tri 2190 162 2203 175 nw
rect 2276 94 2291 322
tri 1813 -28 1819 -22 se
rect 1819 -28 1828 -22
rect 1813 -44 1828 -28
tri 1828 -35 1841 -22 nw
rect 1982 -30 1999 -16
rect 2031 -30 2048 -16
tri 2175 -22 2190 -7 ne
tri 2190 -22 2212 0 sw
rect 1813 -80 1828 -72
rect 1894 -44 1954 -30
rect 1909 -54 1954 -44
rect 1909 -72 1937 -54
tri 1813 -95 1828 -80 ne
tri 1828 -95 1850 -73 sw
rect 1894 -82 1937 -72
rect 1952 -58 1954 -54
rect 2076 -44 2136 -30
tri 2190 -35 2203 -22 ne
rect 2203 -28 2212 -22
tri 2212 -28 2218 -22 sw
rect 2076 -54 2121 -44
rect 1952 -82 2026 -58
rect 1894 -86 2026 -82
tri 2026 -86 2054 -58 sw
rect 2076 -68 2078 -54
tri 2076 -70 2078 -68 ne
rect 2090 -72 2121 -54
rect 2090 -82 2136 -72
rect 2203 -43 2218 -28
tri 1828 -107 1840 -95 ne
rect 1840 -100 1850 -95
tri 1850 -100 1855 -95 sw
rect 1739 -446 1754 -218
rect 1840 -256 1855 -100
rect 1894 -142 1922 -86
tri 2014 -104 2032 -86 ne
rect 2032 -106 2054 -86
tri 2054 -106 2074 -86 sw
tri 2090 -100 2108 -82 ne
rect 1913 -176 1922 -142
rect 1956 -115 1998 -114
rect 1956 -149 1961 -115
rect 1991 -149 1998 -115
rect 1956 -158 1998 -149
rect 2032 -115 2074 -106
rect 2032 -149 2039 -115
rect 2069 -149 2074 -115
rect 2032 -154 2074 -149
rect 2108 -142 2136 -82
tri 2181 -95 2203 -73 se
rect 2203 -80 2218 -72
tri 2203 -95 2218 -80 nw
tri 2175 -101 2181 -95 se
rect 2181 -101 2190 -95
rect 1894 -186 1922 -176
tri 1922 -186 1946 -162 sw
rect 1894 -218 1936 -186
tri 1953 -194 1954 -193 sw
rect 1953 -218 1954 -194
tri 1956 -195 1993 -158 ne
rect 1993 -186 1998 -158
tri 1998 -186 2024 -160 sw
rect 2108 -176 2117 -142
rect 2108 -186 2136 -176
rect 1993 -195 2077 -186
tri 1993 -214 2012 -195 ne
rect 2012 -214 2077 -195
rect 1894 -240 1954 -218
rect 2076 -218 2077 -214
rect 2094 -218 2136 -186
rect 2076 -240 2136 -218
rect 1982 -256 1999 -242
rect 2031 -256 2048 -242
tri 1819 -292 1841 -270 se
rect 1841 -277 1856 -256
tri 1841 -292 1856 -277 nw
rect 2175 -277 2190 -101
tri 2190 -108 2203 -95 nw
rect 2276 -176 2291 52
tri 1813 -298 1819 -292 se
rect 1819 -298 1828 -292
rect 1813 -314 1828 -298
tri 1828 -305 1841 -292 nw
rect 1982 -300 1999 -286
rect 2031 -300 2048 -286
tri 2175 -292 2190 -277 ne
tri 2190 -292 2212 -270 sw
rect 1813 -350 1828 -342
rect 1894 -314 1954 -300
rect 1909 -324 1954 -314
rect 1909 -342 1937 -324
tri 1813 -365 1828 -350 ne
tri 1828 -365 1850 -343 sw
rect 1894 -352 1937 -342
rect 1952 -328 1954 -324
rect 2076 -314 2136 -300
tri 2190 -305 2203 -292 ne
rect 2203 -298 2212 -292
tri 2212 -298 2218 -292 sw
rect 2076 -324 2121 -314
rect 1952 -352 2026 -328
rect 1894 -356 2026 -352
tri 2026 -356 2054 -328 sw
rect 2076 -338 2078 -324
tri 2076 -340 2078 -338 ne
rect 2090 -342 2121 -324
rect 2090 -352 2136 -342
rect 2203 -313 2218 -298
tri 1828 -377 1840 -365 ne
rect 1840 -370 1850 -365
tri 1850 -370 1855 -365 sw
rect 1739 -716 1754 -488
rect 1840 -526 1855 -370
rect 1894 -412 1922 -356
tri 2014 -374 2032 -356 ne
rect 2032 -376 2054 -356
tri 2054 -376 2074 -356 sw
tri 2090 -370 2108 -352 ne
rect 1913 -446 1922 -412
rect 1956 -385 1998 -384
rect 1956 -419 1961 -385
rect 1991 -419 1998 -385
rect 1956 -428 1998 -419
rect 2032 -385 2074 -376
rect 2032 -419 2039 -385
rect 2069 -419 2074 -385
rect 2032 -424 2074 -419
rect 2108 -412 2136 -352
tri 2181 -365 2203 -343 se
rect 2203 -350 2218 -342
tri 2203 -365 2218 -350 nw
tri 2175 -371 2181 -365 se
rect 2181 -371 2190 -365
rect 1894 -456 1922 -446
tri 1922 -456 1946 -432 sw
rect 1894 -488 1936 -456
tri 1953 -464 1954 -463 sw
rect 1953 -488 1954 -464
tri 1956 -465 1993 -428 ne
rect 1993 -456 1998 -428
tri 1998 -456 2024 -430 sw
rect 2108 -446 2117 -412
rect 2108 -456 2136 -446
rect 1993 -465 2077 -456
tri 1993 -484 2012 -465 ne
rect 2012 -484 2077 -465
rect 1894 -510 1954 -488
rect 2076 -488 2077 -484
rect 2094 -488 2136 -456
rect 2076 -510 2136 -488
rect 1982 -526 1999 -512
rect 2031 -526 2048 -512
tri 1819 -562 1841 -540 se
rect 1841 -547 1856 -526
tri 1841 -562 1856 -547 nw
rect 2175 -547 2190 -371
tri 2190 -378 2203 -365 nw
rect 2276 -446 2291 -218
tri 1813 -568 1819 -562 se
rect 1819 -568 1828 -562
rect 1813 -584 1828 -568
tri 1828 -575 1841 -562 nw
rect 1982 -570 1999 -556
rect 2031 -570 2048 -556
tri 2175 -562 2190 -547 ne
tri 2190 -562 2212 -540 sw
rect 1813 -620 1828 -612
rect 1894 -584 1954 -570
rect 1909 -594 1954 -584
rect 1909 -612 1937 -594
tri 1813 -635 1828 -620 ne
tri 1828 -635 1850 -613 sw
rect 1894 -622 1937 -612
rect 1952 -598 1954 -594
rect 2076 -584 2136 -570
tri 2190 -575 2203 -562 ne
rect 2203 -568 2212 -562
tri 2212 -568 2218 -562 sw
rect 2076 -594 2121 -584
rect 1952 -622 2026 -598
rect 1894 -626 2026 -622
tri 2026 -626 2054 -598 sw
rect 2076 -608 2078 -594
tri 2076 -610 2078 -608 ne
rect 2090 -612 2121 -594
rect 2090 -622 2136 -612
rect 2203 -583 2218 -568
tri 1828 -647 1840 -635 ne
rect 1840 -640 1850 -635
tri 1850 -640 1855 -635 sw
rect 1739 -986 1754 -758
rect 1840 -796 1855 -640
rect 1894 -682 1922 -626
tri 2014 -644 2032 -626 ne
rect 2032 -646 2054 -626
tri 2054 -646 2074 -626 sw
tri 2090 -640 2108 -622 ne
rect 1913 -716 1922 -682
rect 1956 -655 1998 -654
rect 1956 -689 1961 -655
rect 1991 -689 1998 -655
rect 1956 -698 1998 -689
rect 2032 -655 2074 -646
rect 2032 -689 2039 -655
rect 2069 -689 2074 -655
rect 2032 -694 2074 -689
rect 2108 -682 2136 -622
tri 2181 -635 2203 -613 se
rect 2203 -620 2218 -612
tri 2203 -635 2218 -620 nw
tri 2175 -641 2181 -635 se
rect 2181 -641 2190 -635
rect 1894 -726 1922 -716
tri 1922 -726 1946 -702 sw
rect 1894 -758 1936 -726
tri 1953 -734 1954 -733 sw
rect 1953 -758 1954 -734
tri 1956 -735 1993 -698 ne
rect 1993 -726 1998 -698
tri 1998 -726 2024 -700 sw
rect 2108 -716 2117 -682
rect 2108 -726 2136 -716
rect 1993 -735 2077 -726
tri 1993 -754 2012 -735 ne
rect 2012 -754 2077 -735
rect 1894 -780 1954 -758
rect 2076 -758 2077 -754
rect 2094 -758 2136 -726
rect 2076 -780 2136 -758
rect 1982 -796 1999 -782
rect 2031 -796 2048 -782
tri 1819 -832 1841 -810 se
rect 1841 -817 1856 -796
tri 1841 -832 1856 -817 nw
rect 2175 -817 2190 -641
tri 2190 -648 2203 -635 nw
rect 2276 -716 2291 -488
tri 1813 -838 1819 -832 se
rect 1819 -838 1828 -832
rect 1813 -854 1828 -838
tri 1828 -845 1841 -832 nw
rect 1982 -840 1999 -826
rect 2031 -840 2048 -826
tri 2175 -832 2190 -817 ne
tri 2190 -832 2212 -810 sw
rect 1813 -890 1828 -882
rect 1894 -854 1954 -840
rect 1909 -864 1954 -854
rect 1909 -882 1937 -864
tri 1813 -905 1828 -890 ne
tri 1828 -905 1850 -883 sw
rect 1894 -892 1937 -882
rect 1952 -868 1954 -864
rect 2076 -854 2136 -840
tri 2190 -845 2203 -832 ne
rect 2203 -838 2212 -832
tri 2212 -838 2218 -832 sw
rect 2076 -864 2121 -854
rect 1952 -892 2026 -868
rect 1894 -896 2026 -892
tri 2026 -896 2054 -868 sw
rect 2076 -878 2078 -864
tri 2076 -880 2078 -878 ne
rect 2090 -882 2121 -864
rect 2090 -892 2136 -882
rect 2203 -853 2218 -838
tri 1828 -917 1840 -905 ne
rect 1840 -910 1850 -905
tri 1850 -910 1855 -905 sw
rect 1739 -1256 1754 -1028
rect 1840 -1066 1855 -910
rect 1894 -952 1922 -896
tri 2014 -914 2032 -896 ne
rect 2032 -916 2054 -896
tri 2054 -916 2074 -896 sw
tri 2090 -910 2108 -892 ne
rect 1913 -986 1922 -952
rect 1956 -925 1998 -924
rect 1956 -959 1961 -925
rect 1991 -959 1998 -925
rect 1956 -968 1998 -959
rect 2032 -925 2074 -916
rect 2032 -959 2039 -925
rect 2069 -959 2074 -925
rect 2032 -964 2074 -959
rect 2108 -952 2136 -892
tri 2181 -905 2203 -883 se
rect 2203 -890 2218 -882
tri 2203 -905 2218 -890 nw
tri 2175 -911 2181 -905 se
rect 2181 -911 2190 -905
rect 1894 -996 1922 -986
tri 1922 -996 1946 -972 sw
rect 1894 -1028 1936 -996
tri 1953 -1004 1954 -1003 sw
rect 1953 -1028 1954 -1004
tri 1956 -1005 1993 -968 ne
rect 1993 -996 1998 -968
tri 1998 -996 2024 -970 sw
rect 2108 -986 2117 -952
rect 2108 -996 2136 -986
rect 1993 -1005 2077 -996
tri 1993 -1024 2012 -1005 ne
rect 2012 -1024 2077 -1005
rect 1894 -1050 1954 -1028
rect 2076 -1028 2077 -1024
rect 2094 -1028 2136 -996
rect 2076 -1050 2136 -1028
rect 1982 -1066 1999 -1052
rect 2031 -1066 2048 -1052
tri 1819 -1102 1841 -1080 se
rect 1841 -1087 1856 -1066
tri 1841 -1102 1856 -1087 nw
rect 2175 -1087 2190 -911
tri 2190 -918 2203 -905 nw
rect 2276 -986 2291 -758
tri 1813 -1108 1819 -1102 se
rect 1819 -1108 1828 -1102
rect 1813 -1124 1828 -1108
tri 1828 -1115 1841 -1102 nw
rect 1982 -1110 1999 -1096
rect 2031 -1110 2048 -1096
tri 2175 -1102 2190 -1087 ne
tri 2190 -1102 2212 -1080 sw
rect 1813 -1160 1828 -1152
rect 1894 -1124 1954 -1110
rect 1909 -1134 1954 -1124
rect 1909 -1152 1937 -1134
tri 1813 -1175 1828 -1160 ne
tri 1828 -1175 1850 -1153 sw
rect 1894 -1162 1937 -1152
rect 1952 -1138 1954 -1134
rect 2076 -1124 2136 -1110
tri 2190 -1115 2203 -1102 ne
rect 2203 -1108 2212 -1102
tri 2212 -1108 2218 -1102 sw
rect 2076 -1134 2121 -1124
rect 1952 -1162 2026 -1138
rect 1894 -1166 2026 -1162
tri 2026 -1166 2054 -1138 sw
rect 2076 -1148 2078 -1134
tri 2076 -1150 2078 -1148 ne
rect 2090 -1152 2121 -1134
rect 2090 -1162 2136 -1152
rect 2203 -1123 2218 -1108
tri 1828 -1187 1840 -1175 ne
rect 1840 -1180 1850 -1175
tri 1850 -1180 1855 -1175 sw
rect 1739 -1526 1754 -1298
rect 1840 -1336 1855 -1180
rect 1894 -1222 1922 -1166
tri 2014 -1184 2032 -1166 ne
rect 2032 -1186 2054 -1166
tri 2054 -1186 2074 -1166 sw
tri 2090 -1180 2108 -1162 ne
rect 1913 -1256 1922 -1222
rect 1956 -1195 1998 -1194
rect 1956 -1229 1961 -1195
rect 1991 -1229 1998 -1195
rect 1956 -1238 1998 -1229
rect 2032 -1195 2074 -1186
rect 2032 -1229 2039 -1195
rect 2069 -1229 2074 -1195
rect 2032 -1234 2074 -1229
rect 2108 -1222 2136 -1162
tri 2181 -1175 2203 -1153 se
rect 2203 -1160 2218 -1152
tri 2203 -1175 2218 -1160 nw
tri 2175 -1181 2181 -1175 se
rect 2181 -1181 2190 -1175
rect 1894 -1266 1922 -1256
tri 1922 -1266 1946 -1242 sw
rect 1894 -1298 1936 -1266
tri 1953 -1274 1954 -1273 sw
rect 1953 -1298 1954 -1274
tri 1956 -1275 1993 -1238 ne
rect 1993 -1266 1998 -1238
tri 1998 -1266 2024 -1240 sw
rect 2108 -1256 2117 -1222
rect 2108 -1266 2136 -1256
rect 1993 -1275 2077 -1266
tri 1993 -1294 2012 -1275 ne
rect 2012 -1294 2077 -1275
rect 1894 -1320 1954 -1298
rect 2076 -1298 2077 -1294
rect 2094 -1298 2136 -1266
rect 2076 -1320 2136 -1298
rect 1982 -1336 1999 -1322
rect 2031 -1336 2048 -1322
tri 1819 -1372 1841 -1350 se
rect 1841 -1357 1856 -1336
tri 1841 -1372 1856 -1357 nw
rect 2175 -1357 2190 -1181
tri 2190 -1188 2203 -1175 nw
rect 2276 -1256 2291 -1028
tri 1813 -1378 1819 -1372 se
rect 1819 -1378 1828 -1372
rect 1813 -1394 1828 -1378
tri 1828 -1385 1841 -1372 nw
rect 1982 -1380 1999 -1366
rect 2031 -1380 2048 -1366
tri 2175 -1372 2190 -1357 ne
tri 2190 -1372 2212 -1350 sw
rect 1813 -1430 1828 -1422
rect 1894 -1394 1954 -1380
rect 1909 -1404 1954 -1394
rect 1909 -1422 1937 -1404
tri 1813 -1445 1828 -1430 ne
tri 1828 -1445 1850 -1423 sw
rect 1894 -1432 1937 -1422
rect 1952 -1408 1954 -1404
rect 2076 -1394 2136 -1380
tri 2190 -1385 2203 -1372 ne
rect 2203 -1378 2212 -1372
tri 2212 -1378 2218 -1372 sw
rect 2076 -1404 2121 -1394
rect 1952 -1432 2026 -1408
rect 1894 -1436 2026 -1432
tri 2026 -1436 2054 -1408 sw
rect 2076 -1418 2078 -1404
tri 2076 -1420 2078 -1418 ne
rect 2090 -1422 2121 -1404
rect 2090 -1432 2136 -1422
rect 2203 -1393 2218 -1378
tri 1828 -1457 1840 -1445 ne
rect 1840 -1450 1850 -1445
tri 1850 -1450 1855 -1445 sw
rect 1739 -1796 1754 -1568
rect 1840 -1606 1855 -1450
rect 1894 -1492 1922 -1436
tri 2014 -1454 2032 -1436 ne
rect 2032 -1456 2054 -1436
tri 2054 -1456 2074 -1436 sw
tri 2090 -1450 2108 -1432 ne
rect 1913 -1526 1922 -1492
rect 1956 -1465 1998 -1464
rect 1956 -1499 1961 -1465
rect 1991 -1499 1998 -1465
rect 1956 -1508 1998 -1499
rect 2032 -1465 2074 -1456
rect 2032 -1499 2039 -1465
rect 2069 -1499 2074 -1465
rect 2032 -1504 2074 -1499
rect 2108 -1492 2136 -1432
tri 2181 -1445 2203 -1423 se
rect 2203 -1430 2218 -1422
tri 2203 -1445 2218 -1430 nw
tri 2175 -1451 2181 -1445 se
rect 2181 -1451 2190 -1445
rect 1894 -1536 1922 -1526
tri 1922 -1536 1946 -1512 sw
rect 1894 -1568 1936 -1536
tri 1953 -1544 1954 -1543 sw
rect 1953 -1568 1954 -1544
tri 1956 -1545 1993 -1508 ne
rect 1993 -1536 1998 -1508
tri 1998 -1536 2024 -1510 sw
rect 2108 -1526 2117 -1492
rect 2108 -1536 2136 -1526
rect 1993 -1545 2077 -1536
tri 1993 -1564 2012 -1545 ne
rect 2012 -1564 2077 -1545
rect 1894 -1590 1954 -1568
rect 2076 -1568 2077 -1564
rect 2094 -1568 2136 -1536
rect 2076 -1590 2136 -1568
rect 1982 -1606 1999 -1592
rect 2031 -1606 2048 -1592
tri 1819 -1642 1841 -1620 se
rect 1841 -1627 1856 -1606
tri 1841 -1642 1856 -1627 nw
rect 2175 -1627 2190 -1451
tri 2190 -1458 2203 -1445 nw
rect 2276 -1526 2291 -1298
tri 1813 -1648 1819 -1642 se
rect 1819 -1648 1828 -1642
rect 1813 -1664 1828 -1648
tri 1828 -1655 1841 -1642 nw
rect 1982 -1650 1999 -1636
rect 2031 -1650 2048 -1636
tri 2175 -1642 2190 -1627 ne
tri 2190 -1642 2212 -1620 sw
rect 1813 -1700 1828 -1692
rect 1894 -1664 1954 -1650
rect 1909 -1674 1954 -1664
rect 1909 -1692 1937 -1674
tri 1813 -1715 1828 -1700 ne
tri 1828 -1715 1850 -1693 sw
rect 1894 -1702 1937 -1692
rect 1952 -1678 1954 -1674
rect 2076 -1664 2136 -1650
tri 2190 -1655 2203 -1642 ne
rect 2203 -1648 2212 -1642
tri 2212 -1648 2218 -1642 sw
rect 2076 -1674 2121 -1664
rect 1952 -1702 2026 -1678
rect 1894 -1706 2026 -1702
tri 2026 -1706 2054 -1678 sw
rect 2076 -1688 2078 -1674
tri 2076 -1690 2078 -1688 ne
rect 2090 -1692 2121 -1674
rect 2090 -1702 2136 -1692
rect 2203 -1663 2218 -1648
tri 1828 -1727 1840 -1715 ne
rect 1840 -1720 1850 -1715
tri 1850 -1720 1855 -1715 sw
rect 1739 -2066 1754 -1838
rect 1840 -1876 1855 -1720
rect 1894 -1762 1922 -1706
tri 2014 -1724 2032 -1706 ne
rect 2032 -1726 2054 -1706
tri 2054 -1726 2074 -1706 sw
tri 2090 -1720 2108 -1702 ne
rect 1913 -1796 1922 -1762
rect 1956 -1735 1998 -1734
rect 1956 -1769 1961 -1735
rect 1991 -1769 1998 -1735
rect 1956 -1778 1998 -1769
rect 2032 -1735 2074 -1726
rect 2032 -1769 2039 -1735
rect 2069 -1769 2074 -1735
rect 2032 -1774 2074 -1769
rect 2108 -1762 2136 -1702
tri 2181 -1715 2203 -1693 se
rect 2203 -1700 2218 -1692
tri 2203 -1715 2218 -1700 nw
tri 2175 -1721 2181 -1715 se
rect 2181 -1721 2190 -1715
rect 1894 -1806 1922 -1796
tri 1922 -1806 1946 -1782 sw
rect 1894 -1838 1936 -1806
tri 1953 -1814 1954 -1813 sw
rect 1953 -1838 1954 -1814
tri 1956 -1815 1993 -1778 ne
rect 1993 -1806 1998 -1778
tri 1998 -1806 2024 -1780 sw
rect 2108 -1796 2117 -1762
rect 2108 -1806 2136 -1796
rect 1993 -1815 2077 -1806
tri 1993 -1834 2012 -1815 ne
rect 2012 -1834 2077 -1815
rect 1894 -1860 1954 -1838
rect 2076 -1838 2077 -1834
rect 2094 -1838 2136 -1806
rect 2076 -1860 2136 -1838
rect 1982 -1876 1999 -1862
rect 2031 -1876 2048 -1862
tri 1819 -1912 1841 -1890 se
rect 1841 -1897 1856 -1876
tri 1841 -1912 1856 -1897 nw
rect 2175 -1897 2190 -1721
tri 2190 -1728 2203 -1715 nw
rect 2276 -1796 2291 -1568
tri 1813 -1918 1819 -1912 se
rect 1819 -1918 1828 -1912
rect 1813 -1934 1828 -1918
tri 1828 -1925 1841 -1912 nw
rect 1982 -1920 1999 -1906
rect 2031 -1920 2048 -1906
tri 2175 -1912 2190 -1897 ne
tri 2190 -1912 2212 -1890 sw
rect 1813 -1970 1828 -1962
rect 1894 -1934 1954 -1920
rect 1909 -1944 1954 -1934
rect 1909 -1962 1937 -1944
tri 1813 -1985 1828 -1970 ne
tri 1828 -1985 1850 -1963 sw
rect 1894 -1972 1937 -1962
rect 1952 -1948 1954 -1944
rect 2076 -1934 2136 -1920
tri 2190 -1925 2203 -1912 ne
rect 2203 -1918 2212 -1912
tri 2212 -1918 2218 -1912 sw
rect 2076 -1944 2121 -1934
rect 1952 -1972 2026 -1948
rect 1894 -1976 2026 -1972
tri 2026 -1976 2054 -1948 sw
rect 2076 -1958 2078 -1944
tri 2076 -1960 2078 -1958 ne
rect 2090 -1962 2121 -1944
rect 2090 -1972 2136 -1962
rect 2203 -1933 2218 -1918
tri 1828 -1997 1840 -1985 ne
rect 1840 -1990 1850 -1985
tri 1850 -1990 1855 -1985 sw
rect 1739 -2146 1754 -2108
rect 1840 -2146 1855 -1990
rect 1894 -2032 1922 -1976
tri 2014 -1994 2032 -1976 ne
rect 2032 -1996 2054 -1976
tri 2054 -1996 2074 -1976 sw
tri 2090 -1990 2108 -1972 ne
rect 1913 -2066 1922 -2032
rect 1956 -2005 1998 -2004
rect 1956 -2039 1961 -2005
rect 1991 -2039 1998 -2005
rect 1956 -2048 1998 -2039
rect 2032 -2005 2074 -1996
rect 2032 -2039 2039 -2005
rect 2069 -2039 2074 -2005
rect 2032 -2044 2074 -2039
rect 2108 -2032 2136 -1972
tri 2181 -1985 2203 -1963 se
rect 2203 -1970 2218 -1962
tri 2203 -1985 2218 -1970 nw
tri 2175 -1991 2181 -1985 se
rect 2181 -1991 2190 -1985
rect 1894 -2076 1922 -2066
tri 1922 -2076 1946 -2052 sw
rect 1894 -2108 1936 -2076
tri 1953 -2084 1954 -2083 sw
rect 1953 -2108 1954 -2084
tri 1956 -2085 1993 -2048 ne
rect 1993 -2076 1998 -2048
tri 1998 -2076 2024 -2050 sw
rect 2108 -2066 2117 -2032
rect 2108 -2076 2136 -2066
rect 1993 -2085 2077 -2076
tri 1993 -2104 2012 -2085 ne
rect 2012 -2104 2077 -2085
rect 1894 -2130 1954 -2108
rect 2076 -2108 2077 -2104
rect 2094 -2108 2136 -2076
rect 2076 -2130 2136 -2108
rect 1982 -2146 1999 -2132
rect 2031 -2146 2048 -2132
rect 2175 -2146 2190 -1991
tri 2190 -1998 2203 -1985 nw
rect 2276 -2066 2291 -1838
rect 2276 -2146 2291 -2108
rect 2319 1984 2334 2174
tri 2399 2138 2421 2160 se
rect 2421 2153 2436 2174
tri 2421 2138 2436 2153 nw
rect 2755 2153 2770 2174
tri 2393 2132 2399 2138 se
rect 2399 2132 2408 2138
rect 2393 2116 2408 2132
tri 2408 2125 2421 2138 nw
rect 2562 2130 2579 2144
rect 2611 2130 2628 2144
tri 2755 2138 2770 2153 ne
tri 2770 2138 2792 2160 sw
rect 2393 2080 2408 2088
rect 2474 2116 2534 2130
rect 2489 2106 2534 2116
rect 2489 2088 2517 2106
tri 2393 2065 2408 2080 ne
tri 2408 2065 2430 2087 sw
rect 2474 2078 2517 2088
rect 2532 2102 2534 2106
rect 2656 2116 2716 2130
tri 2770 2125 2783 2138 ne
rect 2783 2132 2792 2138
tri 2792 2132 2798 2138 sw
rect 2656 2106 2701 2116
rect 2532 2078 2606 2102
rect 2474 2074 2606 2078
tri 2606 2074 2634 2102 sw
rect 2656 2092 2658 2106
tri 2656 2090 2658 2092 ne
rect 2670 2088 2701 2106
rect 2670 2078 2716 2088
rect 2783 2117 2798 2132
tri 2408 2053 2420 2065 ne
rect 2420 2060 2430 2065
tri 2430 2060 2435 2065 sw
rect 2319 1714 2334 1942
rect 2420 1904 2435 2060
rect 2474 2018 2502 2074
tri 2594 2056 2612 2074 ne
rect 2612 2054 2634 2074
tri 2634 2054 2654 2074 sw
tri 2670 2060 2688 2078 ne
rect 2493 1984 2502 2018
rect 2536 2045 2578 2046
rect 2536 2011 2541 2045
rect 2571 2011 2578 2045
rect 2536 2002 2578 2011
rect 2612 2045 2654 2054
rect 2612 2011 2619 2045
rect 2649 2011 2654 2045
rect 2612 2006 2654 2011
rect 2688 2018 2716 2078
tri 2761 2065 2783 2087 se
rect 2783 2080 2798 2088
tri 2783 2065 2798 2080 nw
tri 2755 2059 2761 2065 se
rect 2761 2059 2770 2065
rect 2474 1974 2502 1984
tri 2502 1974 2526 1998 sw
rect 2474 1942 2516 1974
tri 2533 1966 2534 1967 sw
rect 2533 1942 2534 1966
tri 2536 1965 2573 2002 ne
rect 2573 1974 2578 2002
tri 2578 1974 2604 2000 sw
rect 2688 1984 2697 2018
rect 2688 1974 2716 1984
rect 2573 1965 2657 1974
tri 2573 1946 2592 1965 ne
rect 2592 1946 2657 1965
rect 2474 1920 2534 1942
rect 2656 1942 2657 1946
rect 2674 1942 2716 1974
rect 2656 1920 2716 1942
rect 2562 1904 2579 1918
rect 2611 1904 2628 1918
tri 2399 1868 2421 1890 se
rect 2421 1883 2436 1904
tri 2421 1868 2436 1883 nw
rect 2755 1883 2770 2059
tri 2770 2052 2783 2065 nw
rect 2856 1984 2871 2174
tri 2393 1862 2399 1868 se
rect 2399 1862 2408 1868
rect 2393 1846 2408 1862
tri 2408 1855 2421 1868 nw
rect 2562 1860 2579 1874
rect 2611 1860 2628 1874
tri 2755 1868 2770 1883 ne
tri 2770 1868 2792 1890 sw
rect 2393 1810 2408 1818
rect 2474 1846 2534 1860
rect 2489 1836 2534 1846
rect 2489 1818 2517 1836
tri 2393 1795 2408 1810 ne
tri 2408 1795 2430 1817 sw
rect 2474 1808 2517 1818
rect 2532 1832 2534 1836
rect 2656 1846 2716 1860
tri 2770 1855 2783 1868 ne
rect 2783 1862 2792 1868
tri 2792 1862 2798 1868 sw
rect 2656 1836 2701 1846
rect 2532 1808 2606 1832
rect 2474 1804 2606 1808
tri 2606 1804 2634 1832 sw
rect 2656 1822 2658 1836
tri 2656 1820 2658 1822 ne
rect 2670 1818 2701 1836
rect 2670 1808 2716 1818
rect 2783 1847 2798 1862
tri 2408 1783 2420 1795 ne
rect 2420 1790 2430 1795
tri 2430 1790 2435 1795 sw
rect 2319 1444 2334 1672
rect 2420 1634 2435 1790
rect 2474 1748 2502 1804
tri 2594 1786 2612 1804 ne
rect 2612 1784 2634 1804
tri 2634 1784 2654 1804 sw
tri 2670 1790 2688 1808 ne
rect 2493 1714 2502 1748
rect 2536 1775 2578 1776
rect 2536 1741 2541 1775
rect 2571 1741 2578 1775
rect 2536 1732 2578 1741
rect 2612 1775 2654 1784
rect 2612 1741 2619 1775
rect 2649 1741 2654 1775
rect 2612 1736 2654 1741
rect 2688 1748 2716 1808
tri 2761 1795 2783 1817 se
rect 2783 1810 2798 1818
tri 2783 1795 2798 1810 nw
tri 2755 1789 2761 1795 se
rect 2761 1789 2770 1795
rect 2474 1704 2502 1714
tri 2502 1704 2526 1728 sw
rect 2474 1672 2516 1704
tri 2533 1696 2534 1697 sw
rect 2533 1672 2534 1696
tri 2536 1695 2573 1732 ne
rect 2573 1704 2578 1732
tri 2578 1704 2604 1730 sw
rect 2688 1714 2697 1748
rect 2688 1704 2716 1714
rect 2573 1695 2657 1704
tri 2573 1676 2592 1695 ne
rect 2592 1676 2657 1695
rect 2474 1650 2534 1672
rect 2656 1672 2657 1676
rect 2674 1672 2716 1704
rect 2656 1650 2716 1672
rect 2562 1634 2579 1648
rect 2611 1634 2628 1648
tri 2399 1598 2421 1620 se
rect 2421 1613 2436 1634
tri 2421 1598 2436 1613 nw
rect 2755 1613 2770 1789
tri 2770 1782 2783 1795 nw
rect 2856 1714 2871 1942
tri 2393 1592 2399 1598 se
rect 2399 1592 2408 1598
rect 2393 1576 2408 1592
tri 2408 1585 2421 1598 nw
rect 2562 1590 2579 1604
rect 2611 1590 2628 1604
tri 2755 1598 2770 1613 ne
tri 2770 1598 2792 1620 sw
rect 2393 1540 2408 1548
rect 2474 1576 2534 1590
rect 2489 1566 2534 1576
rect 2489 1548 2517 1566
tri 2393 1525 2408 1540 ne
tri 2408 1525 2430 1547 sw
rect 2474 1538 2517 1548
rect 2532 1562 2534 1566
rect 2656 1576 2716 1590
tri 2770 1585 2783 1598 ne
rect 2783 1592 2792 1598
tri 2792 1592 2798 1598 sw
rect 2656 1566 2701 1576
rect 2532 1538 2606 1562
rect 2474 1534 2606 1538
tri 2606 1534 2634 1562 sw
rect 2656 1552 2658 1566
tri 2656 1550 2658 1552 ne
rect 2670 1548 2701 1566
rect 2670 1538 2716 1548
rect 2783 1577 2798 1592
tri 2408 1513 2420 1525 ne
rect 2420 1520 2430 1525
tri 2430 1520 2435 1525 sw
rect 2319 1174 2334 1402
rect 2420 1364 2435 1520
rect 2474 1478 2502 1534
tri 2594 1516 2612 1534 ne
rect 2612 1514 2634 1534
tri 2634 1514 2654 1534 sw
tri 2670 1520 2688 1538 ne
rect 2493 1444 2502 1478
rect 2536 1505 2578 1506
rect 2536 1471 2541 1505
rect 2571 1471 2578 1505
rect 2536 1462 2578 1471
rect 2612 1505 2654 1514
rect 2612 1471 2619 1505
rect 2649 1471 2654 1505
rect 2612 1466 2654 1471
rect 2688 1478 2716 1538
tri 2761 1525 2783 1547 se
rect 2783 1540 2798 1548
tri 2783 1525 2798 1540 nw
tri 2755 1519 2761 1525 se
rect 2761 1519 2770 1525
rect 2474 1434 2502 1444
tri 2502 1434 2526 1458 sw
rect 2474 1402 2516 1434
tri 2533 1426 2534 1427 sw
rect 2533 1402 2534 1426
tri 2536 1425 2573 1462 ne
rect 2573 1434 2578 1462
tri 2578 1434 2604 1460 sw
rect 2688 1444 2697 1478
rect 2688 1434 2716 1444
rect 2573 1425 2657 1434
tri 2573 1406 2592 1425 ne
rect 2592 1406 2657 1425
rect 2474 1380 2534 1402
rect 2656 1402 2657 1406
rect 2674 1402 2716 1434
rect 2656 1380 2716 1402
rect 2562 1364 2579 1378
rect 2611 1364 2628 1378
tri 2399 1328 2421 1350 se
rect 2421 1343 2436 1364
tri 2421 1328 2436 1343 nw
rect 2755 1343 2770 1519
tri 2770 1512 2783 1525 nw
rect 2856 1444 2871 1672
tri 2393 1322 2399 1328 se
rect 2399 1322 2408 1328
rect 2393 1306 2408 1322
tri 2408 1315 2421 1328 nw
rect 2562 1320 2579 1334
rect 2611 1320 2628 1334
tri 2755 1328 2770 1343 ne
tri 2770 1328 2792 1350 sw
rect 2393 1270 2408 1278
rect 2474 1306 2534 1320
rect 2489 1296 2534 1306
rect 2489 1278 2517 1296
tri 2393 1255 2408 1270 ne
tri 2408 1255 2430 1277 sw
rect 2474 1268 2517 1278
rect 2532 1292 2534 1296
rect 2656 1306 2716 1320
tri 2770 1315 2783 1328 ne
rect 2783 1322 2792 1328
tri 2792 1322 2798 1328 sw
rect 2656 1296 2701 1306
rect 2532 1268 2606 1292
rect 2474 1264 2606 1268
tri 2606 1264 2634 1292 sw
rect 2656 1282 2658 1296
tri 2656 1280 2658 1282 ne
rect 2670 1278 2701 1296
rect 2670 1268 2716 1278
rect 2783 1307 2798 1322
tri 2408 1243 2420 1255 ne
rect 2420 1250 2430 1255
tri 2430 1250 2435 1255 sw
rect 2319 904 2334 1132
rect 2420 1094 2435 1250
rect 2474 1208 2502 1264
tri 2594 1246 2612 1264 ne
rect 2612 1244 2634 1264
tri 2634 1244 2654 1264 sw
tri 2670 1250 2688 1268 ne
rect 2493 1174 2502 1208
rect 2536 1235 2578 1236
rect 2536 1201 2541 1235
rect 2571 1201 2578 1235
rect 2536 1192 2578 1201
rect 2612 1235 2654 1244
rect 2612 1201 2619 1235
rect 2649 1201 2654 1235
rect 2612 1196 2654 1201
rect 2688 1208 2716 1268
tri 2761 1255 2783 1277 se
rect 2783 1270 2798 1278
tri 2783 1255 2798 1270 nw
tri 2755 1249 2761 1255 se
rect 2761 1249 2770 1255
rect 2474 1164 2502 1174
tri 2502 1164 2526 1188 sw
rect 2474 1132 2516 1164
tri 2533 1156 2534 1157 sw
rect 2533 1132 2534 1156
tri 2536 1155 2573 1192 ne
rect 2573 1164 2578 1192
tri 2578 1164 2604 1190 sw
rect 2688 1174 2697 1208
rect 2688 1164 2716 1174
rect 2573 1155 2657 1164
tri 2573 1136 2592 1155 ne
rect 2592 1136 2657 1155
rect 2474 1110 2534 1132
rect 2656 1132 2657 1136
rect 2674 1132 2716 1164
rect 2656 1110 2716 1132
rect 2562 1094 2579 1108
rect 2611 1094 2628 1108
tri 2399 1058 2421 1080 se
rect 2421 1073 2436 1094
tri 2421 1058 2436 1073 nw
rect 2755 1073 2770 1249
tri 2770 1242 2783 1255 nw
rect 2856 1174 2871 1402
tri 2393 1052 2399 1058 se
rect 2399 1052 2408 1058
rect 2393 1036 2408 1052
tri 2408 1045 2421 1058 nw
rect 2562 1050 2579 1064
rect 2611 1050 2628 1064
tri 2755 1058 2770 1073 ne
tri 2770 1058 2792 1080 sw
rect 2393 1000 2408 1008
rect 2474 1036 2534 1050
rect 2489 1026 2534 1036
rect 2489 1008 2517 1026
tri 2393 985 2408 1000 ne
tri 2408 985 2430 1007 sw
rect 2474 998 2517 1008
rect 2532 1022 2534 1026
rect 2656 1036 2716 1050
tri 2770 1045 2783 1058 ne
rect 2783 1052 2792 1058
tri 2792 1052 2798 1058 sw
rect 2656 1026 2701 1036
rect 2532 998 2606 1022
rect 2474 994 2606 998
tri 2606 994 2634 1022 sw
rect 2656 1012 2658 1026
tri 2656 1010 2658 1012 ne
rect 2670 1008 2701 1026
rect 2670 998 2716 1008
rect 2783 1037 2798 1052
tri 2408 973 2420 985 ne
rect 2420 980 2430 985
tri 2430 980 2435 985 sw
rect 2319 634 2334 862
rect 2420 824 2435 980
rect 2474 938 2502 994
tri 2594 976 2612 994 ne
rect 2612 974 2634 994
tri 2634 974 2654 994 sw
tri 2670 980 2688 998 ne
rect 2493 904 2502 938
rect 2536 965 2578 966
rect 2536 931 2541 965
rect 2571 931 2578 965
rect 2536 922 2578 931
rect 2612 965 2654 974
rect 2612 931 2619 965
rect 2649 931 2654 965
rect 2612 926 2654 931
rect 2688 938 2716 998
tri 2761 985 2783 1007 se
rect 2783 1000 2798 1008
tri 2783 985 2798 1000 nw
tri 2755 979 2761 985 se
rect 2761 979 2770 985
rect 2474 894 2502 904
tri 2502 894 2526 918 sw
rect 2474 862 2516 894
tri 2533 886 2534 887 sw
rect 2533 862 2534 886
tri 2536 885 2573 922 ne
rect 2573 894 2578 922
tri 2578 894 2604 920 sw
rect 2688 904 2697 938
rect 2688 894 2716 904
rect 2573 885 2657 894
tri 2573 866 2592 885 ne
rect 2592 866 2657 885
rect 2474 840 2534 862
rect 2656 862 2657 866
rect 2674 862 2716 894
rect 2656 840 2716 862
rect 2562 824 2579 838
rect 2611 824 2628 838
tri 2399 788 2421 810 se
rect 2421 803 2436 824
tri 2421 788 2436 803 nw
rect 2755 803 2770 979
tri 2770 972 2783 985 nw
rect 2856 904 2871 1132
tri 2393 782 2399 788 se
rect 2399 782 2408 788
rect 2393 766 2408 782
tri 2408 775 2421 788 nw
rect 2562 780 2579 794
rect 2611 780 2628 794
tri 2755 788 2770 803 ne
tri 2770 788 2792 810 sw
rect 2393 730 2408 738
rect 2474 766 2534 780
rect 2489 756 2534 766
rect 2489 738 2517 756
tri 2393 715 2408 730 ne
tri 2408 715 2430 737 sw
rect 2474 728 2517 738
rect 2532 752 2534 756
rect 2656 766 2716 780
tri 2770 775 2783 788 ne
rect 2783 782 2792 788
tri 2792 782 2798 788 sw
rect 2656 756 2701 766
rect 2532 728 2606 752
rect 2474 724 2606 728
tri 2606 724 2634 752 sw
rect 2656 742 2658 756
tri 2656 740 2658 742 ne
rect 2670 738 2701 756
rect 2670 728 2716 738
rect 2783 767 2798 782
tri 2408 703 2420 715 ne
rect 2420 710 2430 715
tri 2430 710 2435 715 sw
rect 2319 364 2334 592
rect 2420 554 2435 710
rect 2474 668 2502 724
tri 2594 706 2612 724 ne
rect 2612 704 2634 724
tri 2634 704 2654 724 sw
tri 2670 710 2688 728 ne
rect 2493 634 2502 668
rect 2536 695 2578 696
rect 2536 661 2541 695
rect 2571 661 2578 695
rect 2536 652 2578 661
rect 2612 695 2654 704
rect 2612 661 2619 695
rect 2649 661 2654 695
rect 2612 656 2654 661
rect 2688 668 2716 728
tri 2761 715 2783 737 se
rect 2783 730 2798 738
tri 2783 715 2798 730 nw
tri 2755 709 2761 715 se
rect 2761 709 2770 715
rect 2474 624 2502 634
tri 2502 624 2526 648 sw
rect 2474 592 2516 624
tri 2533 616 2534 617 sw
rect 2533 592 2534 616
tri 2536 615 2573 652 ne
rect 2573 624 2578 652
tri 2578 624 2604 650 sw
rect 2688 634 2697 668
rect 2688 624 2716 634
rect 2573 615 2657 624
tri 2573 596 2592 615 ne
rect 2592 596 2657 615
rect 2474 570 2534 592
rect 2656 592 2657 596
rect 2674 592 2716 624
rect 2656 570 2716 592
rect 2562 554 2579 568
rect 2611 554 2628 568
tri 2399 518 2421 540 se
rect 2421 533 2436 554
tri 2421 518 2436 533 nw
rect 2755 533 2770 709
tri 2770 702 2783 715 nw
rect 2856 634 2871 862
tri 2393 512 2399 518 se
rect 2399 512 2408 518
rect 2393 496 2408 512
tri 2408 505 2421 518 nw
rect 2562 510 2579 524
rect 2611 510 2628 524
tri 2755 518 2770 533 ne
tri 2770 518 2792 540 sw
rect 2393 460 2408 468
rect 2474 496 2534 510
rect 2489 486 2534 496
rect 2489 468 2517 486
tri 2393 445 2408 460 ne
tri 2408 445 2430 467 sw
rect 2474 458 2517 468
rect 2532 482 2534 486
rect 2656 496 2716 510
tri 2770 505 2783 518 ne
rect 2783 512 2792 518
tri 2792 512 2798 518 sw
rect 2656 486 2701 496
rect 2532 458 2606 482
rect 2474 454 2606 458
tri 2606 454 2634 482 sw
rect 2656 472 2658 486
tri 2656 470 2658 472 ne
rect 2670 468 2701 486
rect 2670 458 2716 468
rect 2783 497 2798 512
tri 2408 433 2420 445 ne
rect 2420 440 2430 445
tri 2430 440 2435 445 sw
rect 2319 94 2334 322
rect 2420 284 2435 440
rect 2474 398 2502 454
tri 2594 436 2612 454 ne
rect 2612 434 2634 454
tri 2634 434 2654 454 sw
tri 2670 440 2688 458 ne
rect 2493 364 2502 398
rect 2536 425 2578 426
rect 2536 391 2541 425
rect 2571 391 2578 425
rect 2536 382 2578 391
rect 2612 425 2654 434
rect 2612 391 2619 425
rect 2649 391 2654 425
rect 2612 386 2654 391
rect 2688 398 2716 458
tri 2761 445 2783 467 se
rect 2783 460 2798 468
tri 2783 445 2798 460 nw
tri 2755 439 2761 445 se
rect 2761 439 2770 445
rect 2474 354 2502 364
tri 2502 354 2526 378 sw
rect 2474 322 2516 354
tri 2533 346 2534 347 sw
rect 2533 322 2534 346
tri 2536 345 2573 382 ne
rect 2573 354 2578 382
tri 2578 354 2604 380 sw
rect 2688 364 2697 398
rect 2688 354 2716 364
rect 2573 345 2657 354
tri 2573 326 2592 345 ne
rect 2592 326 2657 345
rect 2474 300 2534 322
rect 2656 322 2657 326
rect 2674 322 2716 354
rect 2656 300 2716 322
rect 2562 284 2579 298
rect 2611 284 2628 298
tri 2399 248 2421 270 se
rect 2421 263 2436 284
tri 2421 248 2436 263 nw
rect 2755 263 2770 439
tri 2770 432 2783 445 nw
rect 2856 364 2871 592
tri 2393 242 2399 248 se
rect 2399 242 2408 248
rect 2393 226 2408 242
tri 2408 235 2421 248 nw
rect 2562 240 2579 254
rect 2611 240 2628 254
tri 2755 248 2770 263 ne
tri 2770 248 2792 270 sw
rect 2393 190 2408 198
rect 2474 226 2534 240
rect 2489 216 2534 226
rect 2489 198 2517 216
tri 2393 175 2408 190 ne
tri 2408 175 2430 197 sw
rect 2474 188 2517 198
rect 2532 212 2534 216
rect 2656 226 2716 240
tri 2770 235 2783 248 ne
rect 2783 242 2792 248
tri 2792 242 2798 248 sw
rect 2656 216 2701 226
rect 2532 188 2606 212
rect 2474 184 2606 188
tri 2606 184 2634 212 sw
rect 2656 202 2658 216
tri 2656 200 2658 202 ne
rect 2670 198 2701 216
rect 2670 188 2716 198
rect 2783 227 2798 242
tri 2408 163 2420 175 ne
rect 2420 170 2430 175
tri 2430 170 2435 175 sw
rect 2319 -176 2334 52
rect 2420 14 2435 170
rect 2474 128 2502 184
tri 2594 166 2612 184 ne
rect 2612 164 2634 184
tri 2634 164 2654 184 sw
tri 2670 170 2688 188 ne
rect 2493 94 2502 128
rect 2536 155 2578 156
rect 2536 121 2541 155
rect 2571 121 2578 155
rect 2536 112 2578 121
rect 2612 155 2654 164
rect 2612 121 2619 155
rect 2649 121 2654 155
rect 2612 116 2654 121
rect 2688 128 2716 188
tri 2761 175 2783 197 se
rect 2783 190 2798 198
tri 2783 175 2798 190 nw
tri 2755 169 2761 175 se
rect 2761 169 2770 175
rect 2474 84 2502 94
tri 2502 84 2526 108 sw
rect 2474 52 2516 84
tri 2533 76 2534 77 sw
rect 2533 52 2534 76
tri 2536 75 2573 112 ne
rect 2573 84 2578 112
tri 2578 84 2604 110 sw
rect 2688 94 2697 128
rect 2688 84 2716 94
rect 2573 75 2657 84
tri 2573 56 2592 75 ne
rect 2592 56 2657 75
rect 2474 30 2534 52
rect 2656 52 2657 56
rect 2674 52 2716 84
rect 2656 30 2716 52
rect 2562 14 2579 28
rect 2611 14 2628 28
tri 2399 -22 2421 0 se
rect 2421 -7 2436 14
tri 2421 -22 2436 -7 nw
rect 2755 -7 2770 169
tri 2770 162 2783 175 nw
rect 2856 94 2871 322
tri 2393 -28 2399 -22 se
rect 2399 -28 2408 -22
rect 2393 -44 2408 -28
tri 2408 -35 2421 -22 nw
rect 2562 -30 2579 -16
rect 2611 -30 2628 -16
tri 2755 -22 2770 -7 ne
tri 2770 -22 2792 0 sw
rect 2393 -80 2408 -72
rect 2474 -44 2534 -30
rect 2489 -54 2534 -44
rect 2489 -72 2517 -54
tri 2393 -95 2408 -80 ne
tri 2408 -95 2430 -73 sw
rect 2474 -82 2517 -72
rect 2532 -58 2534 -54
rect 2656 -44 2716 -30
tri 2770 -35 2783 -22 ne
rect 2783 -28 2792 -22
tri 2792 -28 2798 -22 sw
rect 2656 -54 2701 -44
rect 2532 -82 2606 -58
rect 2474 -86 2606 -82
tri 2606 -86 2634 -58 sw
rect 2656 -68 2658 -54
tri 2656 -70 2658 -68 ne
rect 2670 -72 2701 -54
rect 2670 -82 2716 -72
rect 2783 -43 2798 -28
tri 2408 -107 2420 -95 ne
rect 2420 -100 2430 -95
tri 2430 -100 2435 -95 sw
rect 2319 -446 2334 -218
rect 2420 -256 2435 -100
rect 2474 -142 2502 -86
tri 2594 -104 2612 -86 ne
rect 2612 -106 2634 -86
tri 2634 -106 2654 -86 sw
tri 2670 -100 2688 -82 ne
rect 2493 -176 2502 -142
rect 2536 -115 2578 -114
rect 2536 -149 2541 -115
rect 2571 -149 2578 -115
rect 2536 -158 2578 -149
rect 2612 -115 2654 -106
rect 2612 -149 2619 -115
rect 2649 -149 2654 -115
rect 2612 -154 2654 -149
rect 2688 -142 2716 -82
tri 2761 -95 2783 -73 se
rect 2783 -80 2798 -72
tri 2783 -95 2798 -80 nw
tri 2755 -101 2761 -95 se
rect 2761 -101 2770 -95
rect 2474 -186 2502 -176
tri 2502 -186 2526 -162 sw
rect 2474 -218 2516 -186
tri 2533 -194 2534 -193 sw
rect 2533 -218 2534 -194
tri 2536 -195 2573 -158 ne
rect 2573 -186 2578 -158
tri 2578 -186 2604 -160 sw
rect 2688 -176 2697 -142
rect 2688 -186 2716 -176
rect 2573 -195 2657 -186
tri 2573 -214 2592 -195 ne
rect 2592 -214 2657 -195
rect 2474 -240 2534 -218
rect 2656 -218 2657 -214
rect 2674 -218 2716 -186
rect 2656 -240 2716 -218
rect 2562 -256 2579 -242
rect 2611 -256 2628 -242
tri 2399 -292 2421 -270 se
rect 2421 -277 2436 -256
tri 2421 -292 2436 -277 nw
rect 2755 -277 2770 -101
tri 2770 -108 2783 -95 nw
rect 2856 -176 2871 52
tri 2393 -298 2399 -292 se
rect 2399 -298 2408 -292
rect 2393 -314 2408 -298
tri 2408 -305 2421 -292 nw
rect 2562 -300 2579 -286
rect 2611 -300 2628 -286
tri 2755 -292 2770 -277 ne
tri 2770 -292 2792 -270 sw
rect 2393 -350 2408 -342
rect 2474 -314 2534 -300
rect 2489 -324 2534 -314
rect 2489 -342 2517 -324
tri 2393 -365 2408 -350 ne
tri 2408 -365 2430 -343 sw
rect 2474 -352 2517 -342
rect 2532 -328 2534 -324
rect 2656 -314 2716 -300
tri 2770 -305 2783 -292 ne
rect 2783 -298 2792 -292
tri 2792 -298 2798 -292 sw
rect 2656 -324 2701 -314
rect 2532 -352 2606 -328
rect 2474 -356 2606 -352
tri 2606 -356 2634 -328 sw
rect 2656 -338 2658 -324
tri 2656 -340 2658 -338 ne
rect 2670 -342 2701 -324
rect 2670 -352 2716 -342
rect 2783 -313 2798 -298
tri 2408 -377 2420 -365 ne
rect 2420 -370 2430 -365
tri 2430 -370 2435 -365 sw
rect 2319 -716 2334 -488
rect 2420 -526 2435 -370
rect 2474 -412 2502 -356
tri 2594 -374 2612 -356 ne
rect 2612 -376 2634 -356
tri 2634 -376 2654 -356 sw
tri 2670 -370 2688 -352 ne
rect 2493 -446 2502 -412
rect 2536 -385 2578 -384
rect 2536 -419 2541 -385
rect 2571 -419 2578 -385
rect 2536 -428 2578 -419
rect 2612 -385 2654 -376
rect 2612 -419 2619 -385
rect 2649 -419 2654 -385
rect 2612 -424 2654 -419
rect 2688 -412 2716 -352
tri 2761 -365 2783 -343 se
rect 2783 -350 2798 -342
tri 2783 -365 2798 -350 nw
tri 2755 -371 2761 -365 se
rect 2761 -371 2770 -365
rect 2474 -456 2502 -446
tri 2502 -456 2526 -432 sw
rect 2474 -488 2516 -456
tri 2533 -464 2534 -463 sw
rect 2533 -488 2534 -464
tri 2536 -465 2573 -428 ne
rect 2573 -456 2578 -428
tri 2578 -456 2604 -430 sw
rect 2688 -446 2697 -412
rect 2688 -456 2716 -446
rect 2573 -465 2657 -456
tri 2573 -484 2592 -465 ne
rect 2592 -484 2657 -465
rect 2474 -510 2534 -488
rect 2656 -488 2657 -484
rect 2674 -488 2716 -456
rect 2656 -510 2716 -488
rect 2562 -526 2579 -512
rect 2611 -526 2628 -512
tri 2399 -562 2421 -540 se
rect 2421 -547 2436 -526
tri 2421 -562 2436 -547 nw
rect 2755 -547 2770 -371
tri 2770 -378 2783 -365 nw
rect 2856 -446 2871 -218
tri 2393 -568 2399 -562 se
rect 2399 -568 2408 -562
rect 2393 -584 2408 -568
tri 2408 -575 2421 -562 nw
rect 2562 -570 2579 -556
rect 2611 -570 2628 -556
tri 2755 -562 2770 -547 ne
tri 2770 -562 2792 -540 sw
rect 2393 -620 2408 -612
rect 2474 -584 2534 -570
rect 2489 -594 2534 -584
rect 2489 -612 2517 -594
tri 2393 -635 2408 -620 ne
tri 2408 -635 2430 -613 sw
rect 2474 -622 2517 -612
rect 2532 -598 2534 -594
rect 2656 -584 2716 -570
tri 2770 -575 2783 -562 ne
rect 2783 -568 2792 -562
tri 2792 -568 2798 -562 sw
rect 2656 -594 2701 -584
rect 2532 -622 2606 -598
rect 2474 -626 2606 -622
tri 2606 -626 2634 -598 sw
rect 2656 -608 2658 -594
tri 2656 -610 2658 -608 ne
rect 2670 -612 2701 -594
rect 2670 -622 2716 -612
rect 2783 -583 2798 -568
tri 2408 -647 2420 -635 ne
rect 2420 -640 2430 -635
tri 2430 -640 2435 -635 sw
rect 2319 -986 2334 -758
rect 2420 -796 2435 -640
rect 2474 -682 2502 -626
tri 2594 -644 2612 -626 ne
rect 2612 -646 2634 -626
tri 2634 -646 2654 -626 sw
tri 2670 -640 2688 -622 ne
rect 2493 -716 2502 -682
rect 2536 -655 2578 -654
rect 2536 -689 2541 -655
rect 2571 -689 2578 -655
rect 2536 -698 2578 -689
rect 2612 -655 2654 -646
rect 2612 -689 2619 -655
rect 2649 -689 2654 -655
rect 2612 -694 2654 -689
rect 2688 -682 2716 -622
tri 2761 -635 2783 -613 se
rect 2783 -620 2798 -612
tri 2783 -635 2798 -620 nw
tri 2755 -641 2761 -635 se
rect 2761 -641 2770 -635
rect 2474 -726 2502 -716
tri 2502 -726 2526 -702 sw
rect 2474 -758 2516 -726
tri 2533 -734 2534 -733 sw
rect 2533 -758 2534 -734
tri 2536 -735 2573 -698 ne
rect 2573 -726 2578 -698
tri 2578 -726 2604 -700 sw
rect 2688 -716 2697 -682
rect 2688 -726 2716 -716
rect 2573 -735 2657 -726
tri 2573 -754 2592 -735 ne
rect 2592 -754 2657 -735
rect 2474 -780 2534 -758
rect 2656 -758 2657 -754
rect 2674 -758 2716 -726
rect 2656 -780 2716 -758
rect 2562 -796 2579 -782
rect 2611 -796 2628 -782
tri 2399 -832 2421 -810 se
rect 2421 -817 2436 -796
tri 2421 -832 2436 -817 nw
rect 2755 -817 2770 -641
tri 2770 -648 2783 -635 nw
rect 2856 -716 2871 -488
tri 2393 -838 2399 -832 se
rect 2399 -838 2408 -832
rect 2393 -854 2408 -838
tri 2408 -845 2421 -832 nw
rect 2562 -840 2579 -826
rect 2611 -840 2628 -826
tri 2755 -832 2770 -817 ne
tri 2770 -832 2792 -810 sw
rect 2393 -890 2408 -882
rect 2474 -854 2534 -840
rect 2489 -864 2534 -854
rect 2489 -882 2517 -864
tri 2393 -905 2408 -890 ne
tri 2408 -905 2430 -883 sw
rect 2474 -892 2517 -882
rect 2532 -868 2534 -864
rect 2656 -854 2716 -840
tri 2770 -845 2783 -832 ne
rect 2783 -838 2792 -832
tri 2792 -838 2798 -832 sw
rect 2656 -864 2701 -854
rect 2532 -892 2606 -868
rect 2474 -896 2606 -892
tri 2606 -896 2634 -868 sw
rect 2656 -878 2658 -864
tri 2656 -880 2658 -878 ne
rect 2670 -882 2701 -864
rect 2670 -892 2716 -882
rect 2783 -853 2798 -838
tri 2408 -917 2420 -905 ne
rect 2420 -910 2430 -905
tri 2430 -910 2435 -905 sw
rect 2319 -1256 2334 -1028
rect 2420 -1066 2435 -910
rect 2474 -952 2502 -896
tri 2594 -914 2612 -896 ne
rect 2612 -916 2634 -896
tri 2634 -916 2654 -896 sw
tri 2670 -910 2688 -892 ne
rect 2493 -986 2502 -952
rect 2536 -925 2578 -924
rect 2536 -959 2541 -925
rect 2571 -959 2578 -925
rect 2536 -968 2578 -959
rect 2612 -925 2654 -916
rect 2612 -959 2619 -925
rect 2649 -959 2654 -925
rect 2612 -964 2654 -959
rect 2688 -952 2716 -892
tri 2761 -905 2783 -883 se
rect 2783 -890 2798 -882
tri 2783 -905 2798 -890 nw
tri 2755 -911 2761 -905 se
rect 2761 -911 2770 -905
rect 2474 -996 2502 -986
tri 2502 -996 2526 -972 sw
rect 2474 -1028 2516 -996
tri 2533 -1004 2534 -1003 sw
rect 2533 -1028 2534 -1004
tri 2536 -1005 2573 -968 ne
rect 2573 -996 2578 -968
tri 2578 -996 2604 -970 sw
rect 2688 -986 2697 -952
rect 2688 -996 2716 -986
rect 2573 -1005 2657 -996
tri 2573 -1024 2592 -1005 ne
rect 2592 -1024 2657 -1005
rect 2474 -1050 2534 -1028
rect 2656 -1028 2657 -1024
rect 2674 -1028 2716 -996
rect 2656 -1050 2716 -1028
rect 2562 -1066 2579 -1052
rect 2611 -1066 2628 -1052
tri 2399 -1102 2421 -1080 se
rect 2421 -1087 2436 -1066
tri 2421 -1102 2436 -1087 nw
rect 2755 -1087 2770 -911
tri 2770 -918 2783 -905 nw
rect 2856 -986 2871 -758
tri 2393 -1108 2399 -1102 se
rect 2399 -1108 2408 -1102
rect 2393 -1124 2408 -1108
tri 2408 -1115 2421 -1102 nw
rect 2562 -1110 2579 -1096
rect 2611 -1110 2628 -1096
tri 2755 -1102 2770 -1087 ne
tri 2770 -1102 2792 -1080 sw
rect 2393 -1160 2408 -1152
rect 2474 -1124 2534 -1110
rect 2489 -1134 2534 -1124
rect 2489 -1152 2517 -1134
tri 2393 -1175 2408 -1160 ne
tri 2408 -1175 2430 -1153 sw
rect 2474 -1162 2517 -1152
rect 2532 -1138 2534 -1134
rect 2656 -1124 2716 -1110
tri 2770 -1115 2783 -1102 ne
rect 2783 -1108 2792 -1102
tri 2792 -1108 2798 -1102 sw
rect 2656 -1134 2701 -1124
rect 2532 -1162 2606 -1138
rect 2474 -1166 2606 -1162
tri 2606 -1166 2634 -1138 sw
rect 2656 -1148 2658 -1134
tri 2656 -1150 2658 -1148 ne
rect 2670 -1152 2701 -1134
rect 2670 -1162 2716 -1152
rect 2783 -1123 2798 -1108
tri 2408 -1187 2420 -1175 ne
rect 2420 -1180 2430 -1175
tri 2430 -1180 2435 -1175 sw
rect 2319 -1526 2334 -1298
rect 2420 -1336 2435 -1180
rect 2474 -1222 2502 -1166
tri 2594 -1184 2612 -1166 ne
rect 2612 -1186 2634 -1166
tri 2634 -1186 2654 -1166 sw
tri 2670 -1180 2688 -1162 ne
rect 2493 -1256 2502 -1222
rect 2536 -1195 2578 -1194
rect 2536 -1229 2541 -1195
rect 2571 -1229 2578 -1195
rect 2536 -1238 2578 -1229
rect 2612 -1195 2654 -1186
rect 2612 -1229 2619 -1195
rect 2649 -1229 2654 -1195
rect 2612 -1234 2654 -1229
rect 2688 -1222 2716 -1162
tri 2761 -1175 2783 -1153 se
rect 2783 -1160 2798 -1152
tri 2783 -1175 2798 -1160 nw
tri 2755 -1181 2761 -1175 se
rect 2761 -1181 2770 -1175
rect 2474 -1266 2502 -1256
tri 2502 -1266 2526 -1242 sw
rect 2474 -1298 2516 -1266
tri 2533 -1274 2534 -1273 sw
rect 2533 -1298 2534 -1274
tri 2536 -1275 2573 -1238 ne
rect 2573 -1266 2578 -1238
tri 2578 -1266 2604 -1240 sw
rect 2688 -1256 2697 -1222
rect 2688 -1266 2716 -1256
rect 2573 -1275 2657 -1266
tri 2573 -1294 2592 -1275 ne
rect 2592 -1294 2657 -1275
rect 2474 -1320 2534 -1298
rect 2656 -1298 2657 -1294
rect 2674 -1298 2716 -1266
rect 2656 -1320 2716 -1298
rect 2562 -1336 2579 -1322
rect 2611 -1336 2628 -1322
tri 2399 -1372 2421 -1350 se
rect 2421 -1357 2436 -1336
tri 2421 -1372 2436 -1357 nw
rect 2755 -1357 2770 -1181
tri 2770 -1188 2783 -1175 nw
rect 2856 -1256 2871 -1028
tri 2393 -1378 2399 -1372 se
rect 2399 -1378 2408 -1372
rect 2393 -1394 2408 -1378
tri 2408 -1385 2421 -1372 nw
rect 2562 -1380 2579 -1366
rect 2611 -1380 2628 -1366
tri 2755 -1372 2770 -1357 ne
tri 2770 -1372 2792 -1350 sw
rect 2393 -1430 2408 -1422
rect 2474 -1394 2534 -1380
rect 2489 -1404 2534 -1394
rect 2489 -1422 2517 -1404
tri 2393 -1445 2408 -1430 ne
tri 2408 -1445 2430 -1423 sw
rect 2474 -1432 2517 -1422
rect 2532 -1408 2534 -1404
rect 2656 -1394 2716 -1380
tri 2770 -1385 2783 -1372 ne
rect 2783 -1378 2792 -1372
tri 2792 -1378 2798 -1372 sw
rect 2656 -1404 2701 -1394
rect 2532 -1432 2606 -1408
rect 2474 -1436 2606 -1432
tri 2606 -1436 2634 -1408 sw
rect 2656 -1418 2658 -1404
tri 2656 -1420 2658 -1418 ne
rect 2670 -1422 2701 -1404
rect 2670 -1432 2716 -1422
rect 2783 -1393 2798 -1378
tri 2408 -1457 2420 -1445 ne
rect 2420 -1450 2430 -1445
tri 2430 -1450 2435 -1445 sw
rect 2319 -1796 2334 -1568
rect 2420 -1606 2435 -1450
rect 2474 -1492 2502 -1436
tri 2594 -1454 2612 -1436 ne
rect 2612 -1456 2634 -1436
tri 2634 -1456 2654 -1436 sw
tri 2670 -1450 2688 -1432 ne
rect 2493 -1526 2502 -1492
rect 2536 -1465 2578 -1464
rect 2536 -1499 2541 -1465
rect 2571 -1499 2578 -1465
rect 2536 -1508 2578 -1499
rect 2612 -1465 2654 -1456
rect 2612 -1499 2619 -1465
rect 2649 -1499 2654 -1465
rect 2612 -1504 2654 -1499
rect 2688 -1492 2716 -1432
tri 2761 -1445 2783 -1423 se
rect 2783 -1430 2798 -1422
tri 2783 -1445 2798 -1430 nw
tri 2755 -1451 2761 -1445 se
rect 2761 -1451 2770 -1445
rect 2474 -1536 2502 -1526
tri 2502 -1536 2526 -1512 sw
rect 2474 -1568 2516 -1536
tri 2533 -1544 2534 -1543 sw
rect 2533 -1568 2534 -1544
tri 2536 -1545 2573 -1508 ne
rect 2573 -1536 2578 -1508
tri 2578 -1536 2604 -1510 sw
rect 2688 -1526 2697 -1492
rect 2688 -1536 2716 -1526
rect 2573 -1545 2657 -1536
tri 2573 -1564 2592 -1545 ne
rect 2592 -1564 2657 -1545
rect 2474 -1590 2534 -1568
rect 2656 -1568 2657 -1564
rect 2674 -1568 2716 -1536
rect 2656 -1590 2716 -1568
rect 2562 -1606 2579 -1592
rect 2611 -1606 2628 -1592
tri 2399 -1642 2421 -1620 se
rect 2421 -1627 2436 -1606
tri 2421 -1642 2436 -1627 nw
rect 2755 -1627 2770 -1451
tri 2770 -1458 2783 -1445 nw
rect 2856 -1526 2871 -1298
tri 2393 -1648 2399 -1642 se
rect 2399 -1648 2408 -1642
rect 2393 -1664 2408 -1648
tri 2408 -1655 2421 -1642 nw
rect 2562 -1650 2579 -1636
rect 2611 -1650 2628 -1636
tri 2755 -1642 2770 -1627 ne
tri 2770 -1642 2792 -1620 sw
rect 2393 -1700 2408 -1692
rect 2474 -1664 2534 -1650
rect 2489 -1674 2534 -1664
rect 2489 -1692 2517 -1674
tri 2393 -1715 2408 -1700 ne
tri 2408 -1715 2430 -1693 sw
rect 2474 -1702 2517 -1692
rect 2532 -1678 2534 -1674
rect 2656 -1664 2716 -1650
tri 2770 -1655 2783 -1642 ne
rect 2783 -1648 2792 -1642
tri 2792 -1648 2798 -1642 sw
rect 2656 -1674 2701 -1664
rect 2532 -1702 2606 -1678
rect 2474 -1706 2606 -1702
tri 2606 -1706 2634 -1678 sw
rect 2656 -1688 2658 -1674
tri 2656 -1690 2658 -1688 ne
rect 2670 -1692 2701 -1674
rect 2670 -1702 2716 -1692
rect 2783 -1663 2798 -1648
tri 2408 -1727 2420 -1715 ne
rect 2420 -1720 2430 -1715
tri 2430 -1720 2435 -1715 sw
rect 2319 -2066 2334 -1838
rect 2420 -1876 2435 -1720
rect 2474 -1762 2502 -1706
tri 2594 -1724 2612 -1706 ne
rect 2612 -1726 2634 -1706
tri 2634 -1726 2654 -1706 sw
tri 2670 -1720 2688 -1702 ne
rect 2493 -1796 2502 -1762
rect 2536 -1735 2578 -1734
rect 2536 -1769 2541 -1735
rect 2571 -1769 2578 -1735
rect 2536 -1778 2578 -1769
rect 2612 -1735 2654 -1726
rect 2612 -1769 2619 -1735
rect 2649 -1769 2654 -1735
rect 2612 -1774 2654 -1769
rect 2688 -1762 2716 -1702
tri 2761 -1715 2783 -1693 se
rect 2783 -1700 2798 -1692
tri 2783 -1715 2798 -1700 nw
tri 2755 -1721 2761 -1715 se
rect 2761 -1721 2770 -1715
rect 2474 -1806 2502 -1796
tri 2502 -1806 2526 -1782 sw
rect 2474 -1838 2516 -1806
tri 2533 -1814 2534 -1813 sw
rect 2533 -1838 2534 -1814
tri 2536 -1815 2573 -1778 ne
rect 2573 -1806 2578 -1778
tri 2578 -1806 2604 -1780 sw
rect 2688 -1796 2697 -1762
rect 2688 -1806 2716 -1796
rect 2573 -1815 2657 -1806
tri 2573 -1834 2592 -1815 ne
rect 2592 -1834 2657 -1815
rect 2474 -1860 2534 -1838
rect 2656 -1838 2657 -1834
rect 2674 -1838 2716 -1806
rect 2656 -1860 2716 -1838
rect 2562 -1876 2579 -1862
rect 2611 -1876 2628 -1862
tri 2399 -1912 2421 -1890 se
rect 2421 -1897 2436 -1876
tri 2421 -1912 2436 -1897 nw
rect 2755 -1897 2770 -1721
tri 2770 -1728 2783 -1715 nw
rect 2856 -1796 2871 -1568
tri 2393 -1918 2399 -1912 se
rect 2399 -1918 2408 -1912
rect 2393 -1934 2408 -1918
tri 2408 -1925 2421 -1912 nw
rect 2562 -1920 2579 -1906
rect 2611 -1920 2628 -1906
tri 2755 -1912 2770 -1897 ne
tri 2770 -1912 2792 -1890 sw
rect 2393 -1970 2408 -1962
rect 2474 -1934 2534 -1920
rect 2489 -1944 2534 -1934
rect 2489 -1962 2517 -1944
tri 2393 -1985 2408 -1970 ne
tri 2408 -1985 2430 -1963 sw
rect 2474 -1972 2517 -1962
rect 2532 -1948 2534 -1944
rect 2656 -1934 2716 -1920
tri 2770 -1925 2783 -1912 ne
rect 2783 -1918 2792 -1912
tri 2792 -1918 2798 -1912 sw
rect 2656 -1944 2701 -1934
rect 2532 -1972 2606 -1948
rect 2474 -1976 2606 -1972
tri 2606 -1976 2634 -1948 sw
rect 2656 -1958 2658 -1944
tri 2656 -1960 2658 -1958 ne
rect 2670 -1962 2701 -1944
rect 2670 -1972 2716 -1962
rect 2783 -1933 2798 -1918
tri 2408 -1997 2420 -1985 ne
rect 2420 -1990 2430 -1985
tri 2430 -1990 2435 -1985 sw
rect 2319 -2146 2334 -2108
rect 2420 -2146 2435 -1990
rect 2474 -2032 2502 -1976
tri 2594 -1994 2612 -1976 ne
rect 2612 -1996 2634 -1976
tri 2634 -1996 2654 -1976 sw
tri 2670 -1990 2688 -1972 ne
rect 2493 -2066 2502 -2032
rect 2536 -2005 2578 -2004
rect 2536 -2039 2541 -2005
rect 2571 -2039 2578 -2005
rect 2536 -2048 2578 -2039
rect 2612 -2005 2654 -1996
rect 2612 -2039 2619 -2005
rect 2649 -2039 2654 -2005
rect 2612 -2044 2654 -2039
rect 2688 -2032 2716 -1972
tri 2761 -1985 2783 -1963 se
rect 2783 -1970 2798 -1962
tri 2783 -1985 2798 -1970 nw
tri 2755 -1991 2761 -1985 se
rect 2761 -1991 2770 -1985
rect 2474 -2076 2502 -2066
tri 2502 -2076 2526 -2052 sw
rect 2474 -2108 2516 -2076
tri 2533 -2084 2534 -2083 sw
rect 2533 -2108 2534 -2084
tri 2536 -2085 2573 -2048 ne
rect 2573 -2076 2578 -2048
tri 2578 -2076 2604 -2050 sw
rect 2688 -2066 2697 -2032
rect 2688 -2076 2716 -2066
rect 2573 -2085 2657 -2076
tri 2573 -2104 2592 -2085 ne
rect 2592 -2104 2657 -2085
rect 2474 -2130 2534 -2108
rect 2656 -2108 2657 -2104
rect 2674 -2108 2716 -2076
rect 2656 -2130 2716 -2108
rect 2562 -2146 2579 -2132
rect 2611 -2146 2628 -2132
rect 2755 -2146 2770 -1991
tri 2770 -1998 2783 -1985 nw
rect 2856 -2066 2871 -1838
rect 2856 -2146 2871 -2108
rect 2899 1984 2914 2174
tri 2979 2138 3001 2160 se
rect 3001 2153 3016 2174
tri 3001 2138 3016 2153 nw
rect 3335 2153 3350 2174
tri 2973 2132 2979 2138 se
rect 2979 2132 2988 2138
rect 2973 2116 2988 2132
tri 2988 2125 3001 2138 nw
rect 3142 2130 3159 2144
rect 3191 2130 3208 2144
tri 3335 2138 3350 2153 ne
tri 3350 2138 3372 2160 sw
rect 2973 2080 2988 2088
rect 3054 2116 3114 2130
rect 3069 2106 3114 2116
rect 3069 2088 3097 2106
tri 2973 2065 2988 2080 ne
tri 2988 2065 3010 2087 sw
rect 3054 2078 3097 2088
rect 3112 2102 3114 2106
rect 3236 2116 3296 2130
tri 3350 2125 3363 2138 ne
rect 3363 2132 3372 2138
tri 3372 2132 3378 2138 sw
rect 3236 2106 3281 2116
rect 3112 2078 3186 2102
rect 3054 2074 3186 2078
tri 3186 2074 3214 2102 sw
rect 3236 2092 3238 2106
tri 3236 2090 3238 2092 ne
rect 3250 2088 3281 2106
rect 3250 2078 3296 2088
rect 3363 2117 3378 2132
tri 2988 2053 3000 2065 ne
rect 3000 2060 3010 2065
tri 3010 2060 3015 2065 sw
rect 2899 1714 2914 1942
rect 3000 1904 3015 2060
rect 3054 2018 3082 2074
tri 3174 2056 3192 2074 ne
rect 3192 2054 3214 2074
tri 3214 2054 3234 2074 sw
tri 3250 2060 3268 2078 ne
rect 3073 1984 3082 2018
rect 3116 2045 3158 2046
rect 3116 2011 3121 2045
rect 3151 2011 3158 2045
rect 3116 2002 3158 2011
rect 3192 2045 3234 2054
rect 3192 2011 3199 2045
rect 3229 2011 3234 2045
rect 3192 2006 3234 2011
rect 3268 2018 3296 2078
tri 3341 2065 3363 2087 se
rect 3363 2080 3378 2088
tri 3363 2065 3378 2080 nw
tri 3335 2059 3341 2065 se
rect 3341 2059 3350 2065
rect 3054 1974 3082 1984
tri 3082 1974 3106 1998 sw
rect 3054 1942 3096 1974
tri 3113 1966 3114 1967 sw
rect 3113 1942 3114 1966
tri 3116 1965 3153 2002 ne
rect 3153 1974 3158 2002
tri 3158 1974 3184 2000 sw
rect 3268 1984 3277 2018
rect 3268 1974 3296 1984
rect 3153 1965 3237 1974
tri 3153 1946 3172 1965 ne
rect 3172 1946 3237 1965
rect 3054 1920 3114 1942
rect 3236 1942 3237 1946
rect 3254 1942 3296 1974
rect 3236 1920 3296 1942
rect 3142 1904 3159 1918
rect 3191 1904 3208 1918
tri 2979 1868 3001 1890 se
rect 3001 1883 3016 1904
tri 3001 1868 3016 1883 nw
rect 3335 1883 3350 2059
tri 3350 2052 3363 2065 nw
rect 3436 1984 3451 2174
tri 2973 1862 2979 1868 se
rect 2979 1862 2988 1868
rect 2973 1846 2988 1862
tri 2988 1855 3001 1868 nw
rect 3142 1860 3159 1874
rect 3191 1860 3208 1874
tri 3335 1868 3350 1883 ne
tri 3350 1868 3372 1890 sw
rect 2973 1810 2988 1818
rect 3054 1846 3114 1860
rect 3069 1836 3114 1846
rect 3069 1818 3097 1836
tri 2973 1795 2988 1810 ne
tri 2988 1795 3010 1817 sw
rect 3054 1808 3097 1818
rect 3112 1832 3114 1836
rect 3236 1846 3296 1860
tri 3350 1855 3363 1868 ne
rect 3363 1862 3372 1868
tri 3372 1862 3378 1868 sw
rect 3236 1836 3281 1846
rect 3112 1808 3186 1832
rect 3054 1804 3186 1808
tri 3186 1804 3214 1832 sw
rect 3236 1822 3238 1836
tri 3236 1820 3238 1822 ne
rect 3250 1818 3281 1836
rect 3250 1808 3296 1818
rect 3363 1847 3378 1862
tri 2988 1783 3000 1795 ne
rect 3000 1790 3010 1795
tri 3010 1790 3015 1795 sw
rect 2899 1444 2914 1672
rect 3000 1634 3015 1790
rect 3054 1748 3082 1804
tri 3174 1786 3192 1804 ne
rect 3192 1784 3214 1804
tri 3214 1784 3234 1804 sw
tri 3250 1790 3268 1808 ne
rect 3073 1714 3082 1748
rect 3116 1775 3158 1776
rect 3116 1741 3121 1775
rect 3151 1741 3158 1775
rect 3116 1732 3158 1741
rect 3192 1775 3234 1784
rect 3192 1741 3199 1775
rect 3229 1741 3234 1775
rect 3192 1736 3234 1741
rect 3268 1748 3296 1808
tri 3341 1795 3363 1817 se
rect 3363 1810 3378 1818
tri 3363 1795 3378 1810 nw
tri 3335 1789 3341 1795 se
rect 3341 1789 3350 1795
rect 3054 1704 3082 1714
tri 3082 1704 3106 1728 sw
rect 3054 1672 3096 1704
tri 3113 1696 3114 1697 sw
rect 3113 1672 3114 1696
tri 3116 1695 3153 1732 ne
rect 3153 1704 3158 1732
tri 3158 1704 3184 1730 sw
rect 3268 1714 3277 1748
rect 3268 1704 3296 1714
rect 3153 1695 3237 1704
tri 3153 1676 3172 1695 ne
rect 3172 1676 3237 1695
rect 3054 1650 3114 1672
rect 3236 1672 3237 1676
rect 3254 1672 3296 1704
rect 3236 1650 3296 1672
rect 3142 1634 3159 1648
rect 3191 1634 3208 1648
tri 2979 1598 3001 1620 se
rect 3001 1613 3016 1634
tri 3001 1598 3016 1613 nw
rect 3335 1613 3350 1789
tri 3350 1782 3363 1795 nw
rect 3436 1714 3451 1942
tri 2973 1592 2979 1598 se
rect 2979 1592 2988 1598
rect 2973 1576 2988 1592
tri 2988 1585 3001 1598 nw
rect 3142 1590 3159 1604
rect 3191 1590 3208 1604
tri 3335 1598 3350 1613 ne
tri 3350 1598 3372 1620 sw
rect 2973 1540 2988 1548
rect 3054 1576 3114 1590
rect 3069 1566 3114 1576
rect 3069 1548 3097 1566
tri 2973 1525 2988 1540 ne
tri 2988 1525 3010 1547 sw
rect 3054 1538 3097 1548
rect 3112 1562 3114 1566
rect 3236 1576 3296 1590
tri 3350 1585 3363 1598 ne
rect 3363 1592 3372 1598
tri 3372 1592 3378 1598 sw
rect 3236 1566 3281 1576
rect 3112 1538 3186 1562
rect 3054 1534 3186 1538
tri 3186 1534 3214 1562 sw
rect 3236 1552 3238 1566
tri 3236 1550 3238 1552 ne
rect 3250 1548 3281 1566
rect 3250 1538 3296 1548
rect 3363 1577 3378 1592
tri 2988 1513 3000 1525 ne
rect 3000 1520 3010 1525
tri 3010 1520 3015 1525 sw
rect 2899 1174 2914 1402
rect 3000 1364 3015 1520
rect 3054 1478 3082 1534
tri 3174 1516 3192 1534 ne
rect 3192 1514 3214 1534
tri 3214 1514 3234 1534 sw
tri 3250 1520 3268 1538 ne
rect 3073 1444 3082 1478
rect 3116 1505 3158 1506
rect 3116 1471 3121 1505
rect 3151 1471 3158 1505
rect 3116 1462 3158 1471
rect 3192 1505 3234 1514
rect 3192 1471 3199 1505
rect 3229 1471 3234 1505
rect 3192 1466 3234 1471
rect 3268 1478 3296 1538
tri 3341 1525 3363 1547 se
rect 3363 1540 3378 1548
tri 3363 1525 3378 1540 nw
tri 3335 1519 3341 1525 se
rect 3341 1519 3350 1525
rect 3054 1434 3082 1444
tri 3082 1434 3106 1458 sw
rect 3054 1402 3096 1434
tri 3113 1426 3114 1427 sw
rect 3113 1402 3114 1426
tri 3116 1425 3153 1462 ne
rect 3153 1434 3158 1462
tri 3158 1434 3184 1460 sw
rect 3268 1444 3277 1478
rect 3268 1434 3296 1444
rect 3153 1425 3237 1434
tri 3153 1406 3172 1425 ne
rect 3172 1406 3237 1425
rect 3054 1380 3114 1402
rect 3236 1402 3237 1406
rect 3254 1402 3296 1434
rect 3236 1380 3296 1402
rect 3142 1364 3159 1378
rect 3191 1364 3208 1378
tri 2979 1328 3001 1350 se
rect 3001 1343 3016 1364
tri 3001 1328 3016 1343 nw
rect 3335 1343 3350 1519
tri 3350 1512 3363 1525 nw
rect 3436 1444 3451 1672
tri 2973 1322 2979 1328 se
rect 2979 1322 2988 1328
rect 2973 1306 2988 1322
tri 2988 1315 3001 1328 nw
rect 3142 1320 3159 1334
rect 3191 1320 3208 1334
tri 3335 1328 3350 1343 ne
tri 3350 1328 3372 1350 sw
rect 2973 1270 2988 1278
rect 3054 1306 3114 1320
rect 3069 1296 3114 1306
rect 3069 1278 3097 1296
tri 2973 1255 2988 1270 ne
tri 2988 1255 3010 1277 sw
rect 3054 1268 3097 1278
rect 3112 1292 3114 1296
rect 3236 1306 3296 1320
tri 3350 1315 3363 1328 ne
rect 3363 1322 3372 1328
tri 3372 1322 3378 1328 sw
rect 3236 1296 3281 1306
rect 3112 1268 3186 1292
rect 3054 1264 3186 1268
tri 3186 1264 3214 1292 sw
rect 3236 1282 3238 1296
tri 3236 1280 3238 1282 ne
rect 3250 1278 3281 1296
rect 3250 1268 3296 1278
rect 3363 1307 3378 1322
tri 2988 1243 3000 1255 ne
rect 3000 1250 3010 1255
tri 3010 1250 3015 1255 sw
rect 2899 904 2914 1132
rect 3000 1094 3015 1250
rect 3054 1208 3082 1264
tri 3174 1246 3192 1264 ne
rect 3192 1244 3214 1264
tri 3214 1244 3234 1264 sw
tri 3250 1250 3268 1268 ne
rect 3073 1174 3082 1208
rect 3116 1235 3158 1236
rect 3116 1201 3121 1235
rect 3151 1201 3158 1235
rect 3116 1192 3158 1201
rect 3192 1235 3234 1244
rect 3192 1201 3199 1235
rect 3229 1201 3234 1235
rect 3192 1196 3234 1201
rect 3268 1208 3296 1268
tri 3341 1255 3363 1277 se
rect 3363 1270 3378 1278
tri 3363 1255 3378 1270 nw
tri 3335 1249 3341 1255 se
rect 3341 1249 3350 1255
rect 3054 1164 3082 1174
tri 3082 1164 3106 1188 sw
rect 3054 1132 3096 1164
tri 3113 1156 3114 1157 sw
rect 3113 1132 3114 1156
tri 3116 1155 3153 1192 ne
rect 3153 1164 3158 1192
tri 3158 1164 3184 1190 sw
rect 3268 1174 3277 1208
rect 3268 1164 3296 1174
rect 3153 1155 3237 1164
tri 3153 1136 3172 1155 ne
rect 3172 1136 3237 1155
rect 3054 1110 3114 1132
rect 3236 1132 3237 1136
rect 3254 1132 3296 1164
rect 3236 1110 3296 1132
rect 3142 1094 3159 1108
rect 3191 1094 3208 1108
tri 2979 1058 3001 1080 se
rect 3001 1073 3016 1094
tri 3001 1058 3016 1073 nw
rect 3335 1073 3350 1249
tri 3350 1242 3363 1255 nw
rect 3436 1174 3451 1402
tri 2973 1052 2979 1058 se
rect 2979 1052 2988 1058
rect 2973 1036 2988 1052
tri 2988 1045 3001 1058 nw
rect 3142 1050 3159 1064
rect 3191 1050 3208 1064
tri 3335 1058 3350 1073 ne
tri 3350 1058 3372 1080 sw
rect 2973 1000 2988 1008
rect 3054 1036 3114 1050
rect 3069 1026 3114 1036
rect 3069 1008 3097 1026
tri 2973 985 2988 1000 ne
tri 2988 985 3010 1007 sw
rect 3054 998 3097 1008
rect 3112 1022 3114 1026
rect 3236 1036 3296 1050
tri 3350 1045 3363 1058 ne
rect 3363 1052 3372 1058
tri 3372 1052 3378 1058 sw
rect 3236 1026 3281 1036
rect 3112 998 3186 1022
rect 3054 994 3186 998
tri 3186 994 3214 1022 sw
rect 3236 1012 3238 1026
tri 3236 1010 3238 1012 ne
rect 3250 1008 3281 1026
rect 3250 998 3296 1008
rect 3363 1037 3378 1052
tri 2988 973 3000 985 ne
rect 3000 980 3010 985
tri 3010 980 3015 985 sw
rect 2899 634 2914 862
rect 3000 824 3015 980
rect 3054 938 3082 994
tri 3174 976 3192 994 ne
rect 3192 974 3214 994
tri 3214 974 3234 994 sw
tri 3250 980 3268 998 ne
rect 3073 904 3082 938
rect 3116 965 3158 966
rect 3116 931 3121 965
rect 3151 931 3158 965
rect 3116 922 3158 931
rect 3192 965 3234 974
rect 3192 931 3199 965
rect 3229 931 3234 965
rect 3192 926 3234 931
rect 3268 938 3296 998
tri 3341 985 3363 1007 se
rect 3363 1000 3378 1008
tri 3363 985 3378 1000 nw
tri 3335 979 3341 985 se
rect 3341 979 3350 985
rect 3054 894 3082 904
tri 3082 894 3106 918 sw
rect 3054 862 3096 894
tri 3113 886 3114 887 sw
rect 3113 862 3114 886
tri 3116 885 3153 922 ne
rect 3153 894 3158 922
tri 3158 894 3184 920 sw
rect 3268 904 3277 938
rect 3268 894 3296 904
rect 3153 885 3237 894
tri 3153 866 3172 885 ne
rect 3172 866 3237 885
rect 3054 840 3114 862
rect 3236 862 3237 866
rect 3254 862 3296 894
rect 3236 840 3296 862
rect 3142 824 3159 838
rect 3191 824 3208 838
tri 2979 788 3001 810 se
rect 3001 803 3016 824
tri 3001 788 3016 803 nw
rect 3335 803 3350 979
tri 3350 972 3363 985 nw
rect 3436 904 3451 1132
tri 2973 782 2979 788 se
rect 2979 782 2988 788
rect 2973 766 2988 782
tri 2988 775 3001 788 nw
rect 3142 780 3159 794
rect 3191 780 3208 794
tri 3335 788 3350 803 ne
tri 3350 788 3372 810 sw
rect 2973 730 2988 738
rect 3054 766 3114 780
rect 3069 756 3114 766
rect 3069 738 3097 756
tri 2973 715 2988 730 ne
tri 2988 715 3010 737 sw
rect 3054 728 3097 738
rect 3112 752 3114 756
rect 3236 766 3296 780
tri 3350 775 3363 788 ne
rect 3363 782 3372 788
tri 3372 782 3378 788 sw
rect 3236 756 3281 766
rect 3112 728 3186 752
rect 3054 724 3186 728
tri 3186 724 3214 752 sw
rect 3236 742 3238 756
tri 3236 740 3238 742 ne
rect 3250 738 3281 756
rect 3250 728 3296 738
rect 3363 767 3378 782
tri 2988 703 3000 715 ne
rect 3000 710 3010 715
tri 3010 710 3015 715 sw
rect 2899 364 2914 592
rect 3000 554 3015 710
rect 3054 668 3082 724
tri 3174 706 3192 724 ne
rect 3192 704 3214 724
tri 3214 704 3234 724 sw
tri 3250 710 3268 728 ne
rect 3073 634 3082 668
rect 3116 695 3158 696
rect 3116 661 3121 695
rect 3151 661 3158 695
rect 3116 652 3158 661
rect 3192 695 3234 704
rect 3192 661 3199 695
rect 3229 661 3234 695
rect 3192 656 3234 661
rect 3268 668 3296 728
tri 3341 715 3363 737 se
rect 3363 730 3378 738
tri 3363 715 3378 730 nw
tri 3335 709 3341 715 se
rect 3341 709 3350 715
rect 3054 624 3082 634
tri 3082 624 3106 648 sw
rect 3054 592 3096 624
tri 3113 616 3114 617 sw
rect 3113 592 3114 616
tri 3116 615 3153 652 ne
rect 3153 624 3158 652
tri 3158 624 3184 650 sw
rect 3268 634 3277 668
rect 3268 624 3296 634
rect 3153 615 3237 624
tri 3153 596 3172 615 ne
rect 3172 596 3237 615
rect 3054 570 3114 592
rect 3236 592 3237 596
rect 3254 592 3296 624
rect 3236 570 3296 592
rect 3142 554 3159 568
rect 3191 554 3208 568
tri 2979 518 3001 540 se
rect 3001 533 3016 554
tri 3001 518 3016 533 nw
rect 3335 533 3350 709
tri 3350 702 3363 715 nw
rect 3436 634 3451 862
tri 2973 512 2979 518 se
rect 2979 512 2988 518
rect 2973 496 2988 512
tri 2988 505 3001 518 nw
rect 3142 510 3159 524
rect 3191 510 3208 524
tri 3335 518 3350 533 ne
tri 3350 518 3372 540 sw
rect 2973 460 2988 468
rect 3054 496 3114 510
rect 3069 486 3114 496
rect 3069 468 3097 486
tri 2973 445 2988 460 ne
tri 2988 445 3010 467 sw
rect 3054 458 3097 468
rect 3112 482 3114 486
rect 3236 496 3296 510
tri 3350 505 3363 518 ne
rect 3363 512 3372 518
tri 3372 512 3378 518 sw
rect 3236 486 3281 496
rect 3112 458 3186 482
rect 3054 454 3186 458
tri 3186 454 3214 482 sw
rect 3236 472 3238 486
tri 3236 470 3238 472 ne
rect 3250 468 3281 486
rect 3250 458 3296 468
rect 3363 497 3378 512
tri 2988 433 3000 445 ne
rect 3000 440 3010 445
tri 3010 440 3015 445 sw
rect 2899 94 2914 322
rect 3000 284 3015 440
rect 3054 398 3082 454
tri 3174 436 3192 454 ne
rect 3192 434 3214 454
tri 3214 434 3234 454 sw
tri 3250 440 3268 458 ne
rect 3073 364 3082 398
rect 3116 425 3158 426
rect 3116 391 3121 425
rect 3151 391 3158 425
rect 3116 382 3158 391
rect 3192 425 3234 434
rect 3192 391 3199 425
rect 3229 391 3234 425
rect 3192 386 3234 391
rect 3268 398 3296 458
tri 3341 445 3363 467 se
rect 3363 460 3378 468
tri 3363 445 3378 460 nw
tri 3335 439 3341 445 se
rect 3341 439 3350 445
rect 3054 354 3082 364
tri 3082 354 3106 378 sw
rect 3054 322 3096 354
tri 3113 346 3114 347 sw
rect 3113 322 3114 346
tri 3116 345 3153 382 ne
rect 3153 354 3158 382
tri 3158 354 3184 380 sw
rect 3268 364 3277 398
rect 3268 354 3296 364
rect 3153 345 3237 354
tri 3153 326 3172 345 ne
rect 3172 326 3237 345
rect 3054 300 3114 322
rect 3236 322 3237 326
rect 3254 322 3296 354
rect 3236 300 3296 322
rect 3142 284 3159 298
rect 3191 284 3208 298
tri 2979 248 3001 270 se
rect 3001 263 3016 284
tri 3001 248 3016 263 nw
rect 3335 263 3350 439
tri 3350 432 3363 445 nw
rect 3436 364 3451 592
tri 2973 242 2979 248 se
rect 2979 242 2988 248
rect 2973 226 2988 242
tri 2988 235 3001 248 nw
rect 3142 240 3159 254
rect 3191 240 3208 254
tri 3335 248 3350 263 ne
tri 3350 248 3372 270 sw
rect 2973 190 2988 198
rect 3054 226 3114 240
rect 3069 216 3114 226
rect 3069 198 3097 216
tri 2973 175 2988 190 ne
tri 2988 175 3010 197 sw
rect 3054 188 3097 198
rect 3112 212 3114 216
rect 3236 226 3296 240
tri 3350 235 3363 248 ne
rect 3363 242 3372 248
tri 3372 242 3378 248 sw
rect 3236 216 3281 226
rect 3112 188 3186 212
rect 3054 184 3186 188
tri 3186 184 3214 212 sw
rect 3236 202 3238 216
tri 3236 200 3238 202 ne
rect 3250 198 3281 216
rect 3250 188 3296 198
rect 3363 227 3378 242
tri 2988 163 3000 175 ne
rect 3000 170 3010 175
tri 3010 170 3015 175 sw
rect 2899 -176 2914 52
rect 3000 14 3015 170
rect 3054 128 3082 184
tri 3174 166 3192 184 ne
rect 3192 164 3214 184
tri 3214 164 3234 184 sw
tri 3250 170 3268 188 ne
rect 3073 94 3082 128
rect 3116 155 3158 156
rect 3116 121 3121 155
rect 3151 121 3158 155
rect 3116 112 3158 121
rect 3192 155 3234 164
rect 3192 121 3199 155
rect 3229 121 3234 155
rect 3192 116 3234 121
rect 3268 128 3296 188
tri 3341 175 3363 197 se
rect 3363 190 3378 198
tri 3363 175 3378 190 nw
tri 3335 169 3341 175 se
rect 3341 169 3350 175
rect 3054 84 3082 94
tri 3082 84 3106 108 sw
rect 3054 52 3096 84
tri 3113 76 3114 77 sw
rect 3113 52 3114 76
tri 3116 75 3153 112 ne
rect 3153 84 3158 112
tri 3158 84 3184 110 sw
rect 3268 94 3277 128
rect 3268 84 3296 94
rect 3153 75 3237 84
tri 3153 56 3172 75 ne
rect 3172 56 3237 75
rect 3054 30 3114 52
rect 3236 52 3237 56
rect 3254 52 3296 84
rect 3236 30 3296 52
rect 3142 14 3159 28
rect 3191 14 3208 28
tri 2979 -22 3001 0 se
rect 3001 -7 3016 14
tri 3001 -22 3016 -7 nw
rect 3335 -7 3350 169
tri 3350 162 3363 175 nw
rect 3436 94 3451 322
tri 2973 -28 2979 -22 se
rect 2979 -28 2988 -22
rect 2973 -44 2988 -28
tri 2988 -35 3001 -22 nw
rect 3142 -30 3159 -16
rect 3191 -30 3208 -16
tri 3335 -22 3350 -7 ne
tri 3350 -22 3372 0 sw
rect 2973 -80 2988 -72
rect 3054 -44 3114 -30
rect 3069 -54 3114 -44
rect 3069 -72 3097 -54
tri 2973 -95 2988 -80 ne
tri 2988 -95 3010 -73 sw
rect 3054 -82 3097 -72
rect 3112 -58 3114 -54
rect 3236 -44 3296 -30
tri 3350 -35 3363 -22 ne
rect 3363 -28 3372 -22
tri 3372 -28 3378 -22 sw
rect 3236 -54 3281 -44
rect 3112 -82 3186 -58
rect 3054 -86 3186 -82
tri 3186 -86 3214 -58 sw
rect 3236 -68 3238 -54
tri 3236 -70 3238 -68 ne
rect 3250 -72 3281 -54
rect 3250 -82 3296 -72
rect 3363 -43 3378 -28
tri 2988 -107 3000 -95 ne
rect 3000 -100 3010 -95
tri 3010 -100 3015 -95 sw
rect 2899 -446 2914 -218
rect 3000 -256 3015 -100
rect 3054 -142 3082 -86
tri 3174 -104 3192 -86 ne
rect 3192 -106 3214 -86
tri 3214 -106 3234 -86 sw
tri 3250 -100 3268 -82 ne
rect 3073 -176 3082 -142
rect 3116 -115 3158 -114
rect 3116 -149 3121 -115
rect 3151 -149 3158 -115
rect 3116 -158 3158 -149
rect 3192 -115 3234 -106
rect 3192 -149 3199 -115
rect 3229 -149 3234 -115
rect 3192 -154 3234 -149
rect 3268 -142 3296 -82
tri 3341 -95 3363 -73 se
rect 3363 -80 3378 -72
tri 3363 -95 3378 -80 nw
tri 3335 -101 3341 -95 se
rect 3341 -101 3350 -95
rect 3054 -186 3082 -176
tri 3082 -186 3106 -162 sw
rect 3054 -218 3096 -186
tri 3113 -194 3114 -193 sw
rect 3113 -218 3114 -194
tri 3116 -195 3153 -158 ne
rect 3153 -186 3158 -158
tri 3158 -186 3184 -160 sw
rect 3268 -176 3277 -142
rect 3268 -186 3296 -176
rect 3153 -195 3237 -186
tri 3153 -214 3172 -195 ne
rect 3172 -214 3237 -195
rect 3054 -240 3114 -218
rect 3236 -218 3237 -214
rect 3254 -218 3296 -186
rect 3236 -240 3296 -218
rect 3142 -256 3159 -242
rect 3191 -256 3208 -242
tri 2979 -292 3001 -270 se
rect 3001 -277 3016 -256
tri 3001 -292 3016 -277 nw
rect 3335 -277 3350 -101
tri 3350 -108 3363 -95 nw
rect 3436 -176 3451 52
tri 2973 -298 2979 -292 se
rect 2979 -298 2988 -292
rect 2973 -314 2988 -298
tri 2988 -305 3001 -292 nw
rect 3142 -300 3159 -286
rect 3191 -300 3208 -286
tri 3335 -292 3350 -277 ne
tri 3350 -292 3372 -270 sw
rect 2973 -350 2988 -342
rect 3054 -314 3114 -300
rect 3069 -324 3114 -314
rect 3069 -342 3097 -324
tri 2973 -365 2988 -350 ne
tri 2988 -365 3010 -343 sw
rect 3054 -352 3097 -342
rect 3112 -328 3114 -324
rect 3236 -314 3296 -300
tri 3350 -305 3363 -292 ne
rect 3363 -298 3372 -292
tri 3372 -298 3378 -292 sw
rect 3236 -324 3281 -314
rect 3112 -352 3186 -328
rect 3054 -356 3186 -352
tri 3186 -356 3214 -328 sw
rect 3236 -338 3238 -324
tri 3236 -340 3238 -338 ne
rect 3250 -342 3281 -324
rect 3250 -352 3296 -342
rect 3363 -313 3378 -298
tri 2988 -377 3000 -365 ne
rect 3000 -370 3010 -365
tri 3010 -370 3015 -365 sw
rect 2899 -716 2914 -488
rect 3000 -526 3015 -370
rect 3054 -412 3082 -356
tri 3174 -374 3192 -356 ne
rect 3192 -376 3214 -356
tri 3214 -376 3234 -356 sw
tri 3250 -370 3268 -352 ne
rect 3073 -446 3082 -412
rect 3116 -385 3158 -384
rect 3116 -419 3121 -385
rect 3151 -419 3158 -385
rect 3116 -428 3158 -419
rect 3192 -385 3234 -376
rect 3192 -419 3199 -385
rect 3229 -419 3234 -385
rect 3192 -424 3234 -419
rect 3268 -412 3296 -352
tri 3341 -365 3363 -343 se
rect 3363 -350 3378 -342
tri 3363 -365 3378 -350 nw
tri 3335 -371 3341 -365 se
rect 3341 -371 3350 -365
rect 3054 -456 3082 -446
tri 3082 -456 3106 -432 sw
rect 3054 -488 3096 -456
tri 3113 -464 3114 -463 sw
rect 3113 -488 3114 -464
tri 3116 -465 3153 -428 ne
rect 3153 -456 3158 -428
tri 3158 -456 3184 -430 sw
rect 3268 -446 3277 -412
rect 3268 -456 3296 -446
rect 3153 -465 3237 -456
tri 3153 -484 3172 -465 ne
rect 3172 -484 3237 -465
rect 3054 -510 3114 -488
rect 3236 -488 3237 -484
rect 3254 -488 3296 -456
rect 3236 -510 3296 -488
rect 3142 -526 3159 -512
rect 3191 -526 3208 -512
tri 2979 -562 3001 -540 se
rect 3001 -547 3016 -526
tri 3001 -562 3016 -547 nw
rect 3335 -547 3350 -371
tri 3350 -378 3363 -365 nw
rect 3436 -446 3451 -218
tri 2973 -568 2979 -562 se
rect 2979 -568 2988 -562
rect 2973 -584 2988 -568
tri 2988 -575 3001 -562 nw
rect 3142 -570 3159 -556
rect 3191 -570 3208 -556
tri 3335 -562 3350 -547 ne
tri 3350 -562 3372 -540 sw
rect 2973 -620 2988 -612
rect 3054 -584 3114 -570
rect 3069 -594 3114 -584
rect 3069 -612 3097 -594
tri 2973 -635 2988 -620 ne
tri 2988 -635 3010 -613 sw
rect 3054 -622 3097 -612
rect 3112 -598 3114 -594
rect 3236 -584 3296 -570
tri 3350 -575 3363 -562 ne
rect 3363 -568 3372 -562
tri 3372 -568 3378 -562 sw
rect 3236 -594 3281 -584
rect 3112 -622 3186 -598
rect 3054 -626 3186 -622
tri 3186 -626 3214 -598 sw
rect 3236 -608 3238 -594
tri 3236 -610 3238 -608 ne
rect 3250 -612 3281 -594
rect 3250 -622 3296 -612
rect 3363 -583 3378 -568
tri 2988 -647 3000 -635 ne
rect 3000 -640 3010 -635
tri 3010 -640 3015 -635 sw
rect 2899 -986 2914 -758
rect 3000 -796 3015 -640
rect 3054 -682 3082 -626
tri 3174 -644 3192 -626 ne
rect 3192 -646 3214 -626
tri 3214 -646 3234 -626 sw
tri 3250 -640 3268 -622 ne
rect 3073 -716 3082 -682
rect 3116 -655 3158 -654
rect 3116 -689 3121 -655
rect 3151 -689 3158 -655
rect 3116 -698 3158 -689
rect 3192 -655 3234 -646
rect 3192 -689 3199 -655
rect 3229 -689 3234 -655
rect 3192 -694 3234 -689
rect 3268 -682 3296 -622
tri 3341 -635 3363 -613 se
rect 3363 -620 3378 -612
tri 3363 -635 3378 -620 nw
tri 3335 -641 3341 -635 se
rect 3341 -641 3350 -635
rect 3054 -726 3082 -716
tri 3082 -726 3106 -702 sw
rect 3054 -758 3096 -726
tri 3113 -734 3114 -733 sw
rect 3113 -758 3114 -734
tri 3116 -735 3153 -698 ne
rect 3153 -726 3158 -698
tri 3158 -726 3184 -700 sw
rect 3268 -716 3277 -682
rect 3268 -726 3296 -716
rect 3153 -735 3237 -726
tri 3153 -754 3172 -735 ne
rect 3172 -754 3237 -735
rect 3054 -780 3114 -758
rect 3236 -758 3237 -754
rect 3254 -758 3296 -726
rect 3236 -780 3296 -758
rect 3142 -796 3159 -782
rect 3191 -796 3208 -782
tri 2979 -832 3001 -810 se
rect 3001 -817 3016 -796
tri 3001 -832 3016 -817 nw
rect 3335 -817 3350 -641
tri 3350 -648 3363 -635 nw
rect 3436 -716 3451 -488
tri 2973 -838 2979 -832 se
rect 2979 -838 2988 -832
rect 2973 -854 2988 -838
tri 2988 -845 3001 -832 nw
rect 3142 -840 3159 -826
rect 3191 -840 3208 -826
tri 3335 -832 3350 -817 ne
tri 3350 -832 3372 -810 sw
rect 2973 -890 2988 -882
rect 3054 -854 3114 -840
rect 3069 -864 3114 -854
rect 3069 -882 3097 -864
tri 2973 -905 2988 -890 ne
tri 2988 -905 3010 -883 sw
rect 3054 -892 3097 -882
rect 3112 -868 3114 -864
rect 3236 -854 3296 -840
tri 3350 -845 3363 -832 ne
rect 3363 -838 3372 -832
tri 3372 -838 3378 -832 sw
rect 3236 -864 3281 -854
rect 3112 -892 3186 -868
rect 3054 -896 3186 -892
tri 3186 -896 3214 -868 sw
rect 3236 -878 3238 -864
tri 3236 -880 3238 -878 ne
rect 3250 -882 3281 -864
rect 3250 -892 3296 -882
rect 3363 -853 3378 -838
tri 2988 -917 3000 -905 ne
rect 3000 -910 3010 -905
tri 3010 -910 3015 -905 sw
rect 2899 -1256 2914 -1028
rect 3000 -1066 3015 -910
rect 3054 -952 3082 -896
tri 3174 -914 3192 -896 ne
rect 3192 -916 3214 -896
tri 3214 -916 3234 -896 sw
tri 3250 -910 3268 -892 ne
rect 3073 -986 3082 -952
rect 3116 -925 3158 -924
rect 3116 -959 3121 -925
rect 3151 -959 3158 -925
rect 3116 -968 3158 -959
rect 3192 -925 3234 -916
rect 3192 -959 3199 -925
rect 3229 -959 3234 -925
rect 3192 -964 3234 -959
rect 3268 -952 3296 -892
tri 3341 -905 3363 -883 se
rect 3363 -890 3378 -882
tri 3363 -905 3378 -890 nw
tri 3335 -911 3341 -905 se
rect 3341 -911 3350 -905
rect 3054 -996 3082 -986
tri 3082 -996 3106 -972 sw
rect 3054 -1028 3096 -996
tri 3113 -1004 3114 -1003 sw
rect 3113 -1028 3114 -1004
tri 3116 -1005 3153 -968 ne
rect 3153 -996 3158 -968
tri 3158 -996 3184 -970 sw
rect 3268 -986 3277 -952
rect 3268 -996 3296 -986
rect 3153 -1005 3237 -996
tri 3153 -1024 3172 -1005 ne
rect 3172 -1024 3237 -1005
rect 3054 -1050 3114 -1028
rect 3236 -1028 3237 -1024
rect 3254 -1028 3296 -996
rect 3236 -1050 3296 -1028
rect 3142 -1066 3159 -1052
rect 3191 -1066 3208 -1052
tri 2979 -1102 3001 -1080 se
rect 3001 -1087 3016 -1066
tri 3001 -1102 3016 -1087 nw
rect 3335 -1087 3350 -911
tri 3350 -918 3363 -905 nw
rect 3436 -986 3451 -758
tri 2973 -1108 2979 -1102 se
rect 2979 -1108 2988 -1102
rect 2973 -1124 2988 -1108
tri 2988 -1115 3001 -1102 nw
rect 3142 -1110 3159 -1096
rect 3191 -1110 3208 -1096
tri 3335 -1102 3350 -1087 ne
tri 3350 -1102 3372 -1080 sw
rect 2973 -1160 2988 -1152
rect 3054 -1124 3114 -1110
rect 3069 -1134 3114 -1124
rect 3069 -1152 3097 -1134
tri 2973 -1175 2988 -1160 ne
tri 2988 -1175 3010 -1153 sw
rect 3054 -1162 3097 -1152
rect 3112 -1138 3114 -1134
rect 3236 -1124 3296 -1110
tri 3350 -1115 3363 -1102 ne
rect 3363 -1108 3372 -1102
tri 3372 -1108 3378 -1102 sw
rect 3236 -1134 3281 -1124
rect 3112 -1162 3186 -1138
rect 3054 -1166 3186 -1162
tri 3186 -1166 3214 -1138 sw
rect 3236 -1148 3238 -1134
tri 3236 -1150 3238 -1148 ne
rect 3250 -1152 3281 -1134
rect 3250 -1162 3296 -1152
rect 3363 -1123 3378 -1108
tri 2988 -1187 3000 -1175 ne
rect 3000 -1180 3010 -1175
tri 3010 -1180 3015 -1175 sw
rect 2899 -1526 2914 -1298
rect 3000 -1336 3015 -1180
rect 3054 -1222 3082 -1166
tri 3174 -1184 3192 -1166 ne
rect 3192 -1186 3214 -1166
tri 3214 -1186 3234 -1166 sw
tri 3250 -1180 3268 -1162 ne
rect 3073 -1256 3082 -1222
rect 3116 -1195 3158 -1194
rect 3116 -1229 3121 -1195
rect 3151 -1229 3158 -1195
rect 3116 -1238 3158 -1229
rect 3192 -1195 3234 -1186
rect 3192 -1229 3199 -1195
rect 3229 -1229 3234 -1195
rect 3192 -1234 3234 -1229
rect 3268 -1222 3296 -1162
tri 3341 -1175 3363 -1153 se
rect 3363 -1160 3378 -1152
tri 3363 -1175 3378 -1160 nw
tri 3335 -1181 3341 -1175 se
rect 3341 -1181 3350 -1175
rect 3054 -1266 3082 -1256
tri 3082 -1266 3106 -1242 sw
rect 3054 -1298 3096 -1266
tri 3113 -1274 3114 -1273 sw
rect 3113 -1298 3114 -1274
tri 3116 -1275 3153 -1238 ne
rect 3153 -1266 3158 -1238
tri 3158 -1266 3184 -1240 sw
rect 3268 -1256 3277 -1222
rect 3268 -1266 3296 -1256
rect 3153 -1275 3237 -1266
tri 3153 -1294 3172 -1275 ne
rect 3172 -1294 3237 -1275
rect 3054 -1320 3114 -1298
rect 3236 -1298 3237 -1294
rect 3254 -1298 3296 -1266
rect 3236 -1320 3296 -1298
rect 3142 -1336 3159 -1322
rect 3191 -1336 3208 -1322
tri 2979 -1372 3001 -1350 se
rect 3001 -1357 3016 -1336
tri 3001 -1372 3016 -1357 nw
rect 3335 -1357 3350 -1181
tri 3350 -1188 3363 -1175 nw
rect 3436 -1256 3451 -1028
tri 2973 -1378 2979 -1372 se
rect 2979 -1378 2988 -1372
rect 2973 -1394 2988 -1378
tri 2988 -1385 3001 -1372 nw
rect 3142 -1380 3159 -1366
rect 3191 -1380 3208 -1366
tri 3335 -1372 3350 -1357 ne
tri 3350 -1372 3372 -1350 sw
rect 2973 -1430 2988 -1422
rect 3054 -1394 3114 -1380
rect 3069 -1404 3114 -1394
rect 3069 -1422 3097 -1404
tri 2973 -1445 2988 -1430 ne
tri 2988 -1445 3010 -1423 sw
rect 3054 -1432 3097 -1422
rect 3112 -1408 3114 -1404
rect 3236 -1394 3296 -1380
tri 3350 -1385 3363 -1372 ne
rect 3363 -1378 3372 -1372
tri 3372 -1378 3378 -1372 sw
rect 3236 -1404 3281 -1394
rect 3112 -1432 3186 -1408
rect 3054 -1436 3186 -1432
tri 3186 -1436 3214 -1408 sw
rect 3236 -1418 3238 -1404
tri 3236 -1420 3238 -1418 ne
rect 3250 -1422 3281 -1404
rect 3250 -1432 3296 -1422
rect 3363 -1393 3378 -1378
tri 2988 -1457 3000 -1445 ne
rect 3000 -1450 3010 -1445
tri 3010 -1450 3015 -1445 sw
rect 2899 -1796 2914 -1568
rect 3000 -1606 3015 -1450
rect 3054 -1492 3082 -1436
tri 3174 -1454 3192 -1436 ne
rect 3192 -1456 3214 -1436
tri 3214 -1456 3234 -1436 sw
tri 3250 -1450 3268 -1432 ne
rect 3073 -1526 3082 -1492
rect 3116 -1465 3158 -1464
rect 3116 -1499 3121 -1465
rect 3151 -1499 3158 -1465
rect 3116 -1508 3158 -1499
rect 3192 -1465 3234 -1456
rect 3192 -1499 3199 -1465
rect 3229 -1499 3234 -1465
rect 3192 -1504 3234 -1499
rect 3268 -1492 3296 -1432
tri 3341 -1445 3363 -1423 se
rect 3363 -1430 3378 -1422
tri 3363 -1445 3378 -1430 nw
tri 3335 -1451 3341 -1445 se
rect 3341 -1451 3350 -1445
rect 3054 -1536 3082 -1526
tri 3082 -1536 3106 -1512 sw
rect 3054 -1568 3096 -1536
tri 3113 -1544 3114 -1543 sw
rect 3113 -1568 3114 -1544
tri 3116 -1545 3153 -1508 ne
rect 3153 -1536 3158 -1508
tri 3158 -1536 3184 -1510 sw
rect 3268 -1526 3277 -1492
rect 3268 -1536 3296 -1526
rect 3153 -1545 3237 -1536
tri 3153 -1564 3172 -1545 ne
rect 3172 -1564 3237 -1545
rect 3054 -1590 3114 -1568
rect 3236 -1568 3237 -1564
rect 3254 -1568 3296 -1536
rect 3236 -1590 3296 -1568
rect 3142 -1606 3159 -1592
rect 3191 -1606 3208 -1592
tri 2979 -1642 3001 -1620 se
rect 3001 -1627 3016 -1606
tri 3001 -1642 3016 -1627 nw
rect 3335 -1627 3350 -1451
tri 3350 -1458 3363 -1445 nw
rect 3436 -1526 3451 -1298
tri 2973 -1648 2979 -1642 se
rect 2979 -1648 2988 -1642
rect 2973 -1664 2988 -1648
tri 2988 -1655 3001 -1642 nw
rect 3142 -1650 3159 -1636
rect 3191 -1650 3208 -1636
tri 3335 -1642 3350 -1627 ne
tri 3350 -1642 3372 -1620 sw
rect 2973 -1700 2988 -1692
rect 3054 -1664 3114 -1650
rect 3069 -1674 3114 -1664
rect 3069 -1692 3097 -1674
tri 2973 -1715 2988 -1700 ne
tri 2988 -1715 3010 -1693 sw
rect 3054 -1702 3097 -1692
rect 3112 -1678 3114 -1674
rect 3236 -1664 3296 -1650
tri 3350 -1655 3363 -1642 ne
rect 3363 -1648 3372 -1642
tri 3372 -1648 3378 -1642 sw
rect 3236 -1674 3281 -1664
rect 3112 -1702 3186 -1678
rect 3054 -1706 3186 -1702
tri 3186 -1706 3214 -1678 sw
rect 3236 -1688 3238 -1674
tri 3236 -1690 3238 -1688 ne
rect 3250 -1692 3281 -1674
rect 3250 -1702 3296 -1692
rect 3363 -1663 3378 -1648
tri 2988 -1727 3000 -1715 ne
rect 3000 -1720 3010 -1715
tri 3010 -1720 3015 -1715 sw
rect 2899 -2066 2914 -1838
rect 3000 -1876 3015 -1720
rect 3054 -1762 3082 -1706
tri 3174 -1724 3192 -1706 ne
rect 3192 -1726 3214 -1706
tri 3214 -1726 3234 -1706 sw
tri 3250 -1720 3268 -1702 ne
rect 3073 -1796 3082 -1762
rect 3116 -1735 3158 -1734
rect 3116 -1769 3121 -1735
rect 3151 -1769 3158 -1735
rect 3116 -1778 3158 -1769
rect 3192 -1735 3234 -1726
rect 3192 -1769 3199 -1735
rect 3229 -1769 3234 -1735
rect 3192 -1774 3234 -1769
rect 3268 -1762 3296 -1702
tri 3341 -1715 3363 -1693 se
rect 3363 -1700 3378 -1692
tri 3363 -1715 3378 -1700 nw
tri 3335 -1721 3341 -1715 se
rect 3341 -1721 3350 -1715
rect 3054 -1806 3082 -1796
tri 3082 -1806 3106 -1782 sw
rect 3054 -1838 3096 -1806
tri 3113 -1814 3114 -1813 sw
rect 3113 -1838 3114 -1814
tri 3116 -1815 3153 -1778 ne
rect 3153 -1806 3158 -1778
tri 3158 -1806 3184 -1780 sw
rect 3268 -1796 3277 -1762
rect 3268 -1806 3296 -1796
rect 3153 -1815 3237 -1806
tri 3153 -1834 3172 -1815 ne
rect 3172 -1834 3237 -1815
rect 3054 -1860 3114 -1838
rect 3236 -1838 3237 -1834
rect 3254 -1838 3296 -1806
rect 3236 -1860 3296 -1838
rect 3142 -1876 3159 -1862
rect 3191 -1876 3208 -1862
tri 2979 -1912 3001 -1890 se
rect 3001 -1897 3016 -1876
tri 3001 -1912 3016 -1897 nw
rect 3335 -1897 3350 -1721
tri 3350 -1728 3363 -1715 nw
rect 3436 -1796 3451 -1568
tri 2973 -1918 2979 -1912 se
rect 2979 -1918 2988 -1912
rect 2973 -1934 2988 -1918
tri 2988 -1925 3001 -1912 nw
rect 3142 -1920 3159 -1906
rect 3191 -1920 3208 -1906
tri 3335 -1912 3350 -1897 ne
tri 3350 -1912 3372 -1890 sw
rect 2973 -1970 2988 -1962
rect 3054 -1934 3114 -1920
rect 3069 -1944 3114 -1934
rect 3069 -1962 3097 -1944
tri 2973 -1985 2988 -1970 ne
tri 2988 -1985 3010 -1963 sw
rect 3054 -1972 3097 -1962
rect 3112 -1948 3114 -1944
rect 3236 -1934 3296 -1920
tri 3350 -1925 3363 -1912 ne
rect 3363 -1918 3372 -1912
tri 3372 -1918 3378 -1912 sw
rect 3236 -1944 3281 -1934
rect 3112 -1972 3186 -1948
rect 3054 -1976 3186 -1972
tri 3186 -1976 3214 -1948 sw
rect 3236 -1958 3238 -1944
tri 3236 -1960 3238 -1958 ne
rect 3250 -1962 3281 -1944
rect 3250 -1972 3296 -1962
rect 3363 -1933 3378 -1918
tri 2988 -1997 3000 -1985 ne
rect 3000 -1990 3010 -1985
tri 3010 -1990 3015 -1985 sw
rect 2899 -2146 2914 -2108
rect 3000 -2146 3015 -1990
rect 3054 -2032 3082 -1976
tri 3174 -1994 3192 -1976 ne
rect 3192 -1996 3214 -1976
tri 3214 -1996 3234 -1976 sw
tri 3250 -1990 3268 -1972 ne
rect 3073 -2066 3082 -2032
rect 3116 -2005 3158 -2004
rect 3116 -2039 3121 -2005
rect 3151 -2039 3158 -2005
rect 3116 -2048 3158 -2039
rect 3192 -2005 3234 -1996
rect 3192 -2039 3199 -2005
rect 3229 -2039 3234 -2005
rect 3192 -2044 3234 -2039
rect 3268 -2032 3296 -1972
tri 3341 -1985 3363 -1963 se
rect 3363 -1970 3378 -1962
tri 3363 -1985 3378 -1970 nw
tri 3335 -1991 3341 -1985 se
rect 3341 -1991 3350 -1985
rect 3054 -2076 3082 -2066
tri 3082 -2076 3106 -2052 sw
rect 3054 -2108 3096 -2076
tri 3113 -2084 3114 -2083 sw
rect 3113 -2108 3114 -2084
tri 3116 -2085 3153 -2048 ne
rect 3153 -2076 3158 -2048
tri 3158 -2076 3184 -2050 sw
rect 3268 -2066 3277 -2032
rect 3268 -2076 3296 -2066
rect 3153 -2085 3237 -2076
tri 3153 -2104 3172 -2085 ne
rect 3172 -2104 3237 -2085
rect 3054 -2130 3114 -2108
rect 3236 -2108 3237 -2104
rect 3254 -2108 3296 -2076
rect 3236 -2130 3296 -2108
rect 3142 -2146 3159 -2132
rect 3191 -2146 3208 -2132
rect 3335 -2146 3350 -1991
tri 3350 -1998 3363 -1985 nw
rect 3436 -2066 3451 -1838
rect 3436 -2146 3451 -2108
rect 3479 1984 3494 2174
tri 3559 2138 3581 2160 se
rect 3581 2153 3596 2174
tri 3581 2138 3596 2153 nw
rect 3915 2153 3930 2174
tri 3553 2132 3559 2138 se
rect 3559 2132 3568 2138
rect 3553 2116 3568 2132
tri 3568 2125 3581 2138 nw
rect 3722 2130 3739 2144
rect 3771 2130 3788 2144
tri 3915 2138 3930 2153 ne
tri 3930 2138 3952 2160 sw
rect 3553 2080 3568 2088
rect 3634 2116 3694 2130
rect 3649 2106 3694 2116
rect 3649 2088 3677 2106
tri 3553 2065 3568 2080 ne
tri 3568 2065 3590 2087 sw
rect 3634 2078 3677 2088
rect 3692 2102 3694 2106
rect 3816 2116 3876 2130
tri 3930 2125 3943 2138 ne
rect 3943 2132 3952 2138
tri 3952 2132 3958 2138 sw
rect 3816 2106 3861 2116
rect 3692 2078 3766 2102
rect 3634 2074 3766 2078
tri 3766 2074 3794 2102 sw
rect 3816 2092 3818 2106
tri 3816 2090 3818 2092 ne
rect 3830 2088 3861 2106
rect 3830 2078 3876 2088
rect 3943 2117 3958 2132
tri 3568 2053 3580 2065 ne
rect 3580 2060 3590 2065
tri 3590 2060 3595 2065 sw
rect 3479 1714 3494 1942
rect 3580 1904 3595 2060
rect 3634 2018 3662 2074
tri 3754 2056 3772 2074 ne
rect 3772 2054 3794 2074
tri 3794 2054 3814 2074 sw
tri 3830 2060 3848 2078 ne
rect 3653 1984 3662 2018
rect 3696 2045 3738 2046
rect 3696 2011 3701 2045
rect 3731 2011 3738 2045
rect 3696 2002 3738 2011
rect 3772 2045 3814 2054
rect 3772 2011 3779 2045
rect 3809 2011 3814 2045
rect 3772 2006 3814 2011
rect 3848 2018 3876 2078
tri 3921 2065 3943 2087 se
rect 3943 2080 3958 2088
tri 3943 2065 3958 2080 nw
tri 3915 2059 3921 2065 se
rect 3921 2059 3930 2065
rect 3634 1974 3662 1984
tri 3662 1974 3686 1998 sw
rect 3634 1942 3676 1974
tri 3693 1966 3694 1967 sw
rect 3693 1942 3694 1966
tri 3696 1965 3733 2002 ne
rect 3733 1974 3738 2002
tri 3738 1974 3764 2000 sw
rect 3848 1984 3857 2018
rect 3848 1974 3876 1984
rect 3733 1965 3817 1974
tri 3733 1946 3752 1965 ne
rect 3752 1946 3817 1965
rect 3634 1920 3694 1942
rect 3816 1942 3817 1946
rect 3834 1942 3876 1974
rect 3816 1920 3876 1942
rect 3722 1904 3739 1918
rect 3771 1904 3788 1918
tri 3559 1868 3581 1890 se
rect 3581 1883 3596 1904
tri 3581 1868 3596 1883 nw
rect 3915 1883 3930 2059
tri 3930 2052 3943 2065 nw
rect 4016 1984 4031 2174
tri 3553 1862 3559 1868 se
rect 3559 1862 3568 1868
rect 3553 1846 3568 1862
tri 3568 1855 3581 1868 nw
rect 3722 1860 3739 1874
rect 3771 1860 3788 1874
tri 3915 1868 3930 1883 ne
tri 3930 1868 3952 1890 sw
rect 3553 1810 3568 1818
rect 3634 1846 3694 1860
rect 3649 1836 3694 1846
rect 3649 1818 3677 1836
tri 3553 1795 3568 1810 ne
tri 3568 1795 3590 1817 sw
rect 3634 1808 3677 1818
rect 3692 1832 3694 1836
rect 3816 1846 3876 1860
tri 3930 1855 3943 1868 ne
rect 3943 1862 3952 1868
tri 3952 1862 3958 1868 sw
rect 3816 1836 3861 1846
rect 3692 1808 3766 1832
rect 3634 1804 3766 1808
tri 3766 1804 3794 1832 sw
rect 3816 1822 3818 1836
tri 3816 1820 3818 1822 ne
rect 3830 1818 3861 1836
rect 3830 1808 3876 1818
rect 3943 1847 3958 1862
tri 3568 1783 3580 1795 ne
rect 3580 1790 3590 1795
tri 3590 1790 3595 1795 sw
rect 3479 1444 3494 1672
rect 3580 1634 3595 1790
rect 3634 1748 3662 1804
tri 3754 1786 3772 1804 ne
rect 3772 1784 3794 1804
tri 3794 1784 3814 1804 sw
tri 3830 1790 3848 1808 ne
rect 3653 1714 3662 1748
rect 3696 1775 3738 1776
rect 3696 1741 3701 1775
rect 3731 1741 3738 1775
rect 3696 1732 3738 1741
rect 3772 1775 3814 1784
rect 3772 1741 3779 1775
rect 3809 1741 3814 1775
rect 3772 1736 3814 1741
rect 3848 1748 3876 1808
tri 3921 1795 3943 1817 se
rect 3943 1810 3958 1818
tri 3943 1795 3958 1810 nw
tri 3915 1789 3921 1795 se
rect 3921 1789 3930 1795
rect 3634 1704 3662 1714
tri 3662 1704 3686 1728 sw
rect 3634 1672 3676 1704
tri 3693 1696 3694 1697 sw
rect 3693 1672 3694 1696
tri 3696 1695 3733 1732 ne
rect 3733 1704 3738 1732
tri 3738 1704 3764 1730 sw
rect 3848 1714 3857 1748
rect 3848 1704 3876 1714
rect 3733 1695 3817 1704
tri 3733 1676 3752 1695 ne
rect 3752 1676 3817 1695
rect 3634 1650 3694 1672
rect 3816 1672 3817 1676
rect 3834 1672 3876 1704
rect 3816 1650 3876 1672
rect 3722 1634 3739 1648
rect 3771 1634 3788 1648
tri 3559 1598 3581 1620 se
rect 3581 1613 3596 1634
tri 3581 1598 3596 1613 nw
rect 3915 1613 3930 1789
tri 3930 1782 3943 1795 nw
rect 4016 1714 4031 1942
tri 3553 1592 3559 1598 se
rect 3559 1592 3568 1598
rect 3553 1576 3568 1592
tri 3568 1585 3581 1598 nw
rect 3722 1590 3739 1604
rect 3771 1590 3788 1604
tri 3915 1598 3930 1613 ne
tri 3930 1598 3952 1620 sw
rect 3553 1540 3568 1548
rect 3634 1576 3694 1590
rect 3649 1566 3694 1576
rect 3649 1548 3677 1566
tri 3553 1525 3568 1540 ne
tri 3568 1525 3590 1547 sw
rect 3634 1538 3677 1548
rect 3692 1562 3694 1566
rect 3816 1576 3876 1590
tri 3930 1585 3943 1598 ne
rect 3943 1592 3952 1598
tri 3952 1592 3958 1598 sw
rect 3816 1566 3861 1576
rect 3692 1538 3766 1562
rect 3634 1534 3766 1538
tri 3766 1534 3794 1562 sw
rect 3816 1552 3818 1566
tri 3816 1550 3818 1552 ne
rect 3830 1548 3861 1566
rect 3830 1538 3876 1548
rect 3943 1577 3958 1592
tri 3568 1513 3580 1525 ne
rect 3580 1520 3590 1525
tri 3590 1520 3595 1525 sw
rect 3479 1174 3494 1402
rect 3580 1364 3595 1520
rect 3634 1478 3662 1534
tri 3754 1516 3772 1534 ne
rect 3772 1514 3794 1534
tri 3794 1514 3814 1534 sw
tri 3830 1520 3848 1538 ne
rect 3653 1444 3662 1478
rect 3696 1505 3738 1506
rect 3696 1471 3701 1505
rect 3731 1471 3738 1505
rect 3696 1462 3738 1471
rect 3772 1505 3814 1514
rect 3772 1471 3779 1505
rect 3809 1471 3814 1505
rect 3772 1466 3814 1471
rect 3848 1478 3876 1538
tri 3921 1525 3943 1547 se
rect 3943 1540 3958 1548
tri 3943 1525 3958 1540 nw
tri 3915 1519 3921 1525 se
rect 3921 1519 3930 1525
rect 3634 1434 3662 1444
tri 3662 1434 3686 1458 sw
rect 3634 1402 3676 1434
tri 3693 1426 3694 1427 sw
rect 3693 1402 3694 1426
tri 3696 1425 3733 1462 ne
rect 3733 1434 3738 1462
tri 3738 1434 3764 1460 sw
rect 3848 1444 3857 1478
rect 3848 1434 3876 1444
rect 3733 1425 3817 1434
tri 3733 1406 3752 1425 ne
rect 3752 1406 3817 1425
rect 3634 1380 3694 1402
rect 3816 1402 3817 1406
rect 3834 1402 3876 1434
rect 3816 1380 3876 1402
rect 3722 1364 3739 1378
rect 3771 1364 3788 1378
tri 3559 1328 3581 1350 se
rect 3581 1343 3596 1364
tri 3581 1328 3596 1343 nw
rect 3915 1343 3930 1519
tri 3930 1512 3943 1525 nw
rect 4016 1444 4031 1672
tri 3553 1322 3559 1328 se
rect 3559 1322 3568 1328
rect 3553 1306 3568 1322
tri 3568 1315 3581 1328 nw
rect 3722 1320 3739 1334
rect 3771 1320 3788 1334
tri 3915 1328 3930 1343 ne
tri 3930 1328 3952 1350 sw
rect 3553 1270 3568 1278
rect 3634 1306 3694 1320
rect 3649 1296 3694 1306
rect 3649 1278 3677 1296
tri 3553 1255 3568 1270 ne
tri 3568 1255 3590 1277 sw
rect 3634 1268 3677 1278
rect 3692 1292 3694 1296
rect 3816 1306 3876 1320
tri 3930 1315 3943 1328 ne
rect 3943 1322 3952 1328
tri 3952 1322 3958 1328 sw
rect 3816 1296 3861 1306
rect 3692 1268 3766 1292
rect 3634 1264 3766 1268
tri 3766 1264 3794 1292 sw
rect 3816 1282 3818 1296
tri 3816 1280 3818 1282 ne
rect 3830 1278 3861 1296
rect 3830 1268 3876 1278
rect 3943 1307 3958 1322
tri 3568 1243 3580 1255 ne
rect 3580 1250 3590 1255
tri 3590 1250 3595 1255 sw
rect 3479 904 3494 1132
rect 3580 1094 3595 1250
rect 3634 1208 3662 1264
tri 3754 1246 3772 1264 ne
rect 3772 1244 3794 1264
tri 3794 1244 3814 1264 sw
tri 3830 1250 3848 1268 ne
rect 3653 1174 3662 1208
rect 3696 1235 3738 1236
rect 3696 1201 3701 1235
rect 3731 1201 3738 1235
rect 3696 1192 3738 1201
rect 3772 1235 3814 1244
rect 3772 1201 3779 1235
rect 3809 1201 3814 1235
rect 3772 1196 3814 1201
rect 3848 1208 3876 1268
tri 3921 1255 3943 1277 se
rect 3943 1270 3958 1278
tri 3943 1255 3958 1270 nw
tri 3915 1249 3921 1255 se
rect 3921 1249 3930 1255
rect 3634 1164 3662 1174
tri 3662 1164 3686 1188 sw
rect 3634 1132 3676 1164
tri 3693 1156 3694 1157 sw
rect 3693 1132 3694 1156
tri 3696 1155 3733 1192 ne
rect 3733 1164 3738 1192
tri 3738 1164 3764 1190 sw
rect 3848 1174 3857 1208
rect 3848 1164 3876 1174
rect 3733 1155 3817 1164
tri 3733 1136 3752 1155 ne
rect 3752 1136 3817 1155
rect 3634 1110 3694 1132
rect 3816 1132 3817 1136
rect 3834 1132 3876 1164
rect 3816 1110 3876 1132
rect 3722 1094 3739 1108
rect 3771 1094 3788 1108
tri 3559 1058 3581 1080 se
rect 3581 1073 3596 1094
tri 3581 1058 3596 1073 nw
rect 3915 1073 3930 1249
tri 3930 1242 3943 1255 nw
rect 4016 1174 4031 1402
tri 3553 1052 3559 1058 se
rect 3559 1052 3568 1058
rect 3553 1036 3568 1052
tri 3568 1045 3581 1058 nw
rect 3722 1050 3739 1064
rect 3771 1050 3788 1064
tri 3915 1058 3930 1073 ne
tri 3930 1058 3952 1080 sw
rect 3553 1000 3568 1008
rect 3634 1036 3694 1050
rect 3649 1026 3694 1036
rect 3649 1008 3677 1026
tri 3553 985 3568 1000 ne
tri 3568 985 3590 1007 sw
rect 3634 998 3677 1008
rect 3692 1022 3694 1026
rect 3816 1036 3876 1050
tri 3930 1045 3943 1058 ne
rect 3943 1052 3952 1058
tri 3952 1052 3958 1058 sw
rect 3816 1026 3861 1036
rect 3692 998 3766 1022
rect 3634 994 3766 998
tri 3766 994 3794 1022 sw
rect 3816 1012 3818 1026
tri 3816 1010 3818 1012 ne
rect 3830 1008 3861 1026
rect 3830 998 3876 1008
rect 3943 1037 3958 1052
tri 3568 973 3580 985 ne
rect 3580 980 3590 985
tri 3590 980 3595 985 sw
rect 3479 634 3494 862
rect 3580 824 3595 980
rect 3634 938 3662 994
tri 3754 976 3772 994 ne
rect 3772 974 3794 994
tri 3794 974 3814 994 sw
tri 3830 980 3848 998 ne
rect 3653 904 3662 938
rect 3696 965 3738 966
rect 3696 931 3701 965
rect 3731 931 3738 965
rect 3696 922 3738 931
rect 3772 965 3814 974
rect 3772 931 3779 965
rect 3809 931 3814 965
rect 3772 926 3814 931
rect 3848 938 3876 998
tri 3921 985 3943 1007 se
rect 3943 1000 3958 1008
tri 3943 985 3958 1000 nw
tri 3915 979 3921 985 se
rect 3921 979 3930 985
rect 3634 894 3662 904
tri 3662 894 3686 918 sw
rect 3634 862 3676 894
tri 3693 886 3694 887 sw
rect 3693 862 3694 886
tri 3696 885 3733 922 ne
rect 3733 894 3738 922
tri 3738 894 3764 920 sw
rect 3848 904 3857 938
rect 3848 894 3876 904
rect 3733 885 3817 894
tri 3733 866 3752 885 ne
rect 3752 866 3817 885
rect 3634 840 3694 862
rect 3816 862 3817 866
rect 3834 862 3876 894
rect 3816 840 3876 862
rect 3722 824 3739 838
rect 3771 824 3788 838
tri 3559 788 3581 810 se
rect 3581 803 3596 824
tri 3581 788 3596 803 nw
rect 3915 803 3930 979
tri 3930 972 3943 985 nw
rect 4016 904 4031 1132
tri 3553 782 3559 788 se
rect 3559 782 3568 788
rect 3553 766 3568 782
tri 3568 775 3581 788 nw
rect 3722 780 3739 794
rect 3771 780 3788 794
tri 3915 788 3930 803 ne
tri 3930 788 3952 810 sw
rect 3553 730 3568 738
rect 3634 766 3694 780
rect 3649 756 3694 766
rect 3649 738 3677 756
tri 3553 715 3568 730 ne
tri 3568 715 3590 737 sw
rect 3634 728 3677 738
rect 3692 752 3694 756
rect 3816 766 3876 780
tri 3930 775 3943 788 ne
rect 3943 782 3952 788
tri 3952 782 3958 788 sw
rect 3816 756 3861 766
rect 3692 728 3766 752
rect 3634 724 3766 728
tri 3766 724 3794 752 sw
rect 3816 742 3818 756
tri 3816 740 3818 742 ne
rect 3830 738 3861 756
rect 3830 728 3876 738
rect 3943 767 3958 782
tri 3568 703 3580 715 ne
rect 3580 710 3590 715
tri 3590 710 3595 715 sw
rect 3479 364 3494 592
rect 3580 554 3595 710
rect 3634 668 3662 724
tri 3754 706 3772 724 ne
rect 3772 704 3794 724
tri 3794 704 3814 724 sw
tri 3830 710 3848 728 ne
rect 3653 634 3662 668
rect 3696 695 3738 696
rect 3696 661 3701 695
rect 3731 661 3738 695
rect 3696 652 3738 661
rect 3772 695 3814 704
rect 3772 661 3779 695
rect 3809 661 3814 695
rect 3772 656 3814 661
rect 3848 668 3876 728
tri 3921 715 3943 737 se
rect 3943 730 3958 738
tri 3943 715 3958 730 nw
tri 3915 709 3921 715 se
rect 3921 709 3930 715
rect 3634 624 3662 634
tri 3662 624 3686 648 sw
rect 3634 592 3676 624
tri 3693 616 3694 617 sw
rect 3693 592 3694 616
tri 3696 615 3733 652 ne
rect 3733 624 3738 652
tri 3738 624 3764 650 sw
rect 3848 634 3857 668
rect 3848 624 3876 634
rect 3733 615 3817 624
tri 3733 596 3752 615 ne
rect 3752 596 3817 615
rect 3634 570 3694 592
rect 3816 592 3817 596
rect 3834 592 3876 624
rect 3816 570 3876 592
rect 3722 554 3739 568
rect 3771 554 3788 568
tri 3559 518 3581 540 se
rect 3581 533 3596 554
tri 3581 518 3596 533 nw
rect 3915 533 3930 709
tri 3930 702 3943 715 nw
rect 4016 634 4031 862
tri 3553 512 3559 518 se
rect 3559 512 3568 518
rect 3553 496 3568 512
tri 3568 505 3581 518 nw
rect 3722 510 3739 524
rect 3771 510 3788 524
tri 3915 518 3930 533 ne
tri 3930 518 3952 540 sw
rect 3553 460 3568 468
rect 3634 496 3694 510
rect 3649 486 3694 496
rect 3649 468 3677 486
tri 3553 445 3568 460 ne
tri 3568 445 3590 467 sw
rect 3634 458 3677 468
rect 3692 482 3694 486
rect 3816 496 3876 510
tri 3930 505 3943 518 ne
rect 3943 512 3952 518
tri 3952 512 3958 518 sw
rect 3816 486 3861 496
rect 3692 458 3766 482
rect 3634 454 3766 458
tri 3766 454 3794 482 sw
rect 3816 472 3818 486
tri 3816 470 3818 472 ne
rect 3830 468 3861 486
rect 3830 458 3876 468
rect 3943 497 3958 512
tri 3568 433 3580 445 ne
rect 3580 440 3590 445
tri 3590 440 3595 445 sw
rect 3479 94 3494 322
rect 3580 284 3595 440
rect 3634 398 3662 454
tri 3754 436 3772 454 ne
rect 3772 434 3794 454
tri 3794 434 3814 454 sw
tri 3830 440 3848 458 ne
rect 3653 364 3662 398
rect 3696 425 3738 426
rect 3696 391 3701 425
rect 3731 391 3738 425
rect 3696 382 3738 391
rect 3772 425 3814 434
rect 3772 391 3779 425
rect 3809 391 3814 425
rect 3772 386 3814 391
rect 3848 398 3876 458
tri 3921 445 3943 467 se
rect 3943 460 3958 468
tri 3943 445 3958 460 nw
tri 3915 439 3921 445 se
rect 3921 439 3930 445
rect 3634 354 3662 364
tri 3662 354 3686 378 sw
rect 3634 322 3676 354
tri 3693 346 3694 347 sw
rect 3693 322 3694 346
tri 3696 345 3733 382 ne
rect 3733 354 3738 382
tri 3738 354 3764 380 sw
rect 3848 364 3857 398
rect 3848 354 3876 364
rect 3733 345 3817 354
tri 3733 326 3752 345 ne
rect 3752 326 3817 345
rect 3634 300 3694 322
rect 3816 322 3817 326
rect 3834 322 3876 354
rect 3816 300 3876 322
rect 3722 284 3739 298
rect 3771 284 3788 298
tri 3559 248 3581 270 se
rect 3581 263 3596 284
tri 3581 248 3596 263 nw
rect 3915 263 3930 439
tri 3930 432 3943 445 nw
rect 4016 364 4031 592
tri 3553 242 3559 248 se
rect 3559 242 3568 248
rect 3553 226 3568 242
tri 3568 235 3581 248 nw
rect 3722 240 3739 254
rect 3771 240 3788 254
tri 3915 248 3930 263 ne
tri 3930 248 3952 270 sw
rect 3553 190 3568 198
rect 3634 226 3694 240
rect 3649 216 3694 226
rect 3649 198 3677 216
tri 3553 175 3568 190 ne
tri 3568 175 3590 197 sw
rect 3634 188 3677 198
rect 3692 212 3694 216
rect 3816 226 3876 240
tri 3930 235 3943 248 ne
rect 3943 242 3952 248
tri 3952 242 3958 248 sw
rect 3816 216 3861 226
rect 3692 188 3766 212
rect 3634 184 3766 188
tri 3766 184 3794 212 sw
rect 3816 202 3818 216
tri 3816 200 3818 202 ne
rect 3830 198 3861 216
rect 3830 188 3876 198
rect 3943 227 3958 242
tri 3568 163 3580 175 ne
rect 3580 170 3590 175
tri 3590 170 3595 175 sw
rect 3479 -176 3494 52
rect 3580 14 3595 170
rect 3634 128 3662 184
tri 3754 166 3772 184 ne
rect 3772 164 3794 184
tri 3794 164 3814 184 sw
tri 3830 170 3848 188 ne
rect 3653 94 3662 128
rect 3696 155 3738 156
rect 3696 121 3701 155
rect 3731 121 3738 155
rect 3696 112 3738 121
rect 3772 155 3814 164
rect 3772 121 3779 155
rect 3809 121 3814 155
rect 3772 116 3814 121
rect 3848 128 3876 188
tri 3921 175 3943 197 se
rect 3943 190 3958 198
tri 3943 175 3958 190 nw
tri 3915 169 3921 175 se
rect 3921 169 3930 175
rect 3634 84 3662 94
tri 3662 84 3686 108 sw
rect 3634 52 3676 84
tri 3693 76 3694 77 sw
rect 3693 52 3694 76
tri 3696 75 3733 112 ne
rect 3733 84 3738 112
tri 3738 84 3764 110 sw
rect 3848 94 3857 128
rect 3848 84 3876 94
rect 3733 75 3817 84
tri 3733 56 3752 75 ne
rect 3752 56 3817 75
rect 3634 30 3694 52
rect 3816 52 3817 56
rect 3834 52 3876 84
rect 3816 30 3876 52
rect 3722 14 3739 28
rect 3771 14 3788 28
tri 3559 -22 3581 0 se
rect 3581 -7 3596 14
tri 3581 -22 3596 -7 nw
rect 3915 -7 3930 169
tri 3930 162 3943 175 nw
rect 4016 94 4031 322
tri 3553 -28 3559 -22 se
rect 3559 -28 3568 -22
rect 3553 -44 3568 -28
tri 3568 -35 3581 -22 nw
rect 3722 -30 3739 -16
rect 3771 -30 3788 -16
tri 3915 -22 3930 -7 ne
tri 3930 -22 3952 0 sw
rect 3553 -80 3568 -72
rect 3634 -44 3694 -30
rect 3649 -54 3694 -44
rect 3649 -72 3677 -54
tri 3553 -95 3568 -80 ne
tri 3568 -95 3590 -73 sw
rect 3634 -82 3677 -72
rect 3692 -58 3694 -54
rect 3816 -44 3876 -30
tri 3930 -35 3943 -22 ne
rect 3943 -28 3952 -22
tri 3952 -28 3958 -22 sw
rect 3816 -54 3861 -44
rect 3692 -82 3766 -58
rect 3634 -86 3766 -82
tri 3766 -86 3794 -58 sw
rect 3816 -68 3818 -54
tri 3816 -70 3818 -68 ne
rect 3830 -72 3861 -54
rect 3830 -82 3876 -72
rect 3943 -43 3958 -28
tri 3568 -107 3580 -95 ne
rect 3580 -100 3590 -95
tri 3590 -100 3595 -95 sw
rect 3479 -446 3494 -218
rect 3580 -256 3595 -100
rect 3634 -142 3662 -86
tri 3754 -104 3772 -86 ne
rect 3772 -106 3794 -86
tri 3794 -106 3814 -86 sw
tri 3830 -100 3848 -82 ne
rect 3653 -176 3662 -142
rect 3696 -115 3738 -114
rect 3696 -149 3701 -115
rect 3731 -149 3738 -115
rect 3696 -158 3738 -149
rect 3772 -115 3814 -106
rect 3772 -149 3779 -115
rect 3809 -149 3814 -115
rect 3772 -154 3814 -149
rect 3848 -142 3876 -82
tri 3921 -95 3943 -73 se
rect 3943 -80 3958 -72
tri 3943 -95 3958 -80 nw
tri 3915 -101 3921 -95 se
rect 3921 -101 3930 -95
rect 3634 -186 3662 -176
tri 3662 -186 3686 -162 sw
rect 3634 -218 3676 -186
tri 3693 -194 3694 -193 sw
rect 3693 -218 3694 -194
tri 3696 -195 3733 -158 ne
rect 3733 -186 3738 -158
tri 3738 -186 3764 -160 sw
rect 3848 -176 3857 -142
rect 3848 -186 3876 -176
rect 3733 -195 3817 -186
tri 3733 -214 3752 -195 ne
rect 3752 -214 3817 -195
rect 3634 -240 3694 -218
rect 3816 -218 3817 -214
rect 3834 -218 3876 -186
rect 3816 -240 3876 -218
rect 3722 -256 3739 -242
rect 3771 -256 3788 -242
tri 3559 -292 3581 -270 se
rect 3581 -277 3596 -256
tri 3581 -292 3596 -277 nw
rect 3915 -277 3930 -101
tri 3930 -108 3943 -95 nw
rect 4016 -176 4031 52
tri 3553 -298 3559 -292 se
rect 3559 -298 3568 -292
rect 3553 -314 3568 -298
tri 3568 -305 3581 -292 nw
rect 3722 -300 3739 -286
rect 3771 -300 3788 -286
tri 3915 -292 3930 -277 ne
tri 3930 -292 3952 -270 sw
rect 3553 -350 3568 -342
rect 3634 -314 3694 -300
rect 3649 -324 3694 -314
rect 3649 -342 3677 -324
tri 3553 -365 3568 -350 ne
tri 3568 -365 3590 -343 sw
rect 3634 -352 3677 -342
rect 3692 -328 3694 -324
rect 3816 -314 3876 -300
tri 3930 -305 3943 -292 ne
rect 3943 -298 3952 -292
tri 3952 -298 3958 -292 sw
rect 3816 -324 3861 -314
rect 3692 -352 3766 -328
rect 3634 -356 3766 -352
tri 3766 -356 3794 -328 sw
rect 3816 -338 3818 -324
tri 3816 -340 3818 -338 ne
rect 3830 -342 3861 -324
rect 3830 -352 3876 -342
rect 3943 -313 3958 -298
tri 3568 -377 3580 -365 ne
rect 3580 -370 3590 -365
tri 3590 -370 3595 -365 sw
rect 3479 -716 3494 -488
rect 3580 -526 3595 -370
rect 3634 -412 3662 -356
tri 3754 -374 3772 -356 ne
rect 3772 -376 3794 -356
tri 3794 -376 3814 -356 sw
tri 3830 -370 3848 -352 ne
rect 3653 -446 3662 -412
rect 3696 -385 3738 -384
rect 3696 -419 3701 -385
rect 3731 -419 3738 -385
rect 3696 -428 3738 -419
rect 3772 -385 3814 -376
rect 3772 -419 3779 -385
rect 3809 -419 3814 -385
rect 3772 -424 3814 -419
rect 3848 -412 3876 -352
tri 3921 -365 3943 -343 se
rect 3943 -350 3958 -342
tri 3943 -365 3958 -350 nw
tri 3915 -371 3921 -365 se
rect 3921 -371 3930 -365
rect 3634 -456 3662 -446
tri 3662 -456 3686 -432 sw
rect 3634 -488 3676 -456
tri 3693 -464 3694 -463 sw
rect 3693 -488 3694 -464
tri 3696 -465 3733 -428 ne
rect 3733 -456 3738 -428
tri 3738 -456 3764 -430 sw
rect 3848 -446 3857 -412
rect 3848 -456 3876 -446
rect 3733 -465 3817 -456
tri 3733 -484 3752 -465 ne
rect 3752 -484 3817 -465
rect 3634 -510 3694 -488
rect 3816 -488 3817 -484
rect 3834 -488 3876 -456
rect 3816 -510 3876 -488
rect 3722 -526 3739 -512
rect 3771 -526 3788 -512
tri 3559 -562 3581 -540 se
rect 3581 -547 3596 -526
tri 3581 -562 3596 -547 nw
rect 3915 -547 3930 -371
tri 3930 -378 3943 -365 nw
rect 4016 -446 4031 -218
tri 3553 -568 3559 -562 se
rect 3559 -568 3568 -562
rect 3553 -584 3568 -568
tri 3568 -575 3581 -562 nw
rect 3722 -570 3739 -556
rect 3771 -570 3788 -556
tri 3915 -562 3930 -547 ne
tri 3930 -562 3952 -540 sw
rect 3553 -620 3568 -612
rect 3634 -584 3694 -570
rect 3649 -594 3694 -584
rect 3649 -612 3677 -594
tri 3553 -635 3568 -620 ne
tri 3568 -635 3590 -613 sw
rect 3634 -622 3677 -612
rect 3692 -598 3694 -594
rect 3816 -584 3876 -570
tri 3930 -575 3943 -562 ne
rect 3943 -568 3952 -562
tri 3952 -568 3958 -562 sw
rect 3816 -594 3861 -584
rect 3692 -622 3766 -598
rect 3634 -626 3766 -622
tri 3766 -626 3794 -598 sw
rect 3816 -608 3818 -594
tri 3816 -610 3818 -608 ne
rect 3830 -612 3861 -594
rect 3830 -622 3876 -612
rect 3943 -583 3958 -568
tri 3568 -647 3580 -635 ne
rect 3580 -640 3590 -635
tri 3590 -640 3595 -635 sw
rect 3479 -986 3494 -758
rect 3580 -796 3595 -640
rect 3634 -682 3662 -626
tri 3754 -644 3772 -626 ne
rect 3772 -646 3794 -626
tri 3794 -646 3814 -626 sw
tri 3830 -640 3848 -622 ne
rect 3653 -716 3662 -682
rect 3696 -655 3738 -654
rect 3696 -689 3701 -655
rect 3731 -689 3738 -655
rect 3696 -698 3738 -689
rect 3772 -655 3814 -646
rect 3772 -689 3779 -655
rect 3809 -689 3814 -655
rect 3772 -694 3814 -689
rect 3848 -682 3876 -622
tri 3921 -635 3943 -613 se
rect 3943 -620 3958 -612
tri 3943 -635 3958 -620 nw
tri 3915 -641 3921 -635 se
rect 3921 -641 3930 -635
rect 3634 -726 3662 -716
tri 3662 -726 3686 -702 sw
rect 3634 -758 3676 -726
tri 3693 -734 3694 -733 sw
rect 3693 -758 3694 -734
tri 3696 -735 3733 -698 ne
rect 3733 -726 3738 -698
tri 3738 -726 3764 -700 sw
rect 3848 -716 3857 -682
rect 3848 -726 3876 -716
rect 3733 -735 3817 -726
tri 3733 -754 3752 -735 ne
rect 3752 -754 3817 -735
rect 3634 -780 3694 -758
rect 3816 -758 3817 -754
rect 3834 -758 3876 -726
rect 3816 -780 3876 -758
rect 3722 -796 3739 -782
rect 3771 -796 3788 -782
tri 3559 -832 3581 -810 se
rect 3581 -817 3596 -796
tri 3581 -832 3596 -817 nw
rect 3915 -817 3930 -641
tri 3930 -648 3943 -635 nw
rect 4016 -716 4031 -488
tri 3553 -838 3559 -832 se
rect 3559 -838 3568 -832
rect 3553 -854 3568 -838
tri 3568 -845 3581 -832 nw
rect 3722 -840 3739 -826
rect 3771 -840 3788 -826
tri 3915 -832 3930 -817 ne
tri 3930 -832 3952 -810 sw
rect 3553 -890 3568 -882
rect 3634 -854 3694 -840
rect 3649 -864 3694 -854
rect 3649 -882 3677 -864
tri 3553 -905 3568 -890 ne
tri 3568 -905 3590 -883 sw
rect 3634 -892 3677 -882
rect 3692 -868 3694 -864
rect 3816 -854 3876 -840
tri 3930 -845 3943 -832 ne
rect 3943 -838 3952 -832
tri 3952 -838 3958 -832 sw
rect 3816 -864 3861 -854
rect 3692 -892 3766 -868
rect 3634 -896 3766 -892
tri 3766 -896 3794 -868 sw
rect 3816 -878 3818 -864
tri 3816 -880 3818 -878 ne
rect 3830 -882 3861 -864
rect 3830 -892 3876 -882
rect 3943 -853 3958 -838
tri 3568 -917 3580 -905 ne
rect 3580 -910 3590 -905
tri 3590 -910 3595 -905 sw
rect 3479 -1256 3494 -1028
rect 3580 -1066 3595 -910
rect 3634 -952 3662 -896
tri 3754 -914 3772 -896 ne
rect 3772 -916 3794 -896
tri 3794 -916 3814 -896 sw
tri 3830 -910 3848 -892 ne
rect 3653 -986 3662 -952
rect 3696 -925 3738 -924
rect 3696 -959 3701 -925
rect 3731 -959 3738 -925
rect 3696 -968 3738 -959
rect 3772 -925 3814 -916
rect 3772 -959 3779 -925
rect 3809 -959 3814 -925
rect 3772 -964 3814 -959
rect 3848 -952 3876 -892
tri 3921 -905 3943 -883 se
rect 3943 -890 3958 -882
tri 3943 -905 3958 -890 nw
tri 3915 -911 3921 -905 se
rect 3921 -911 3930 -905
rect 3634 -996 3662 -986
tri 3662 -996 3686 -972 sw
rect 3634 -1028 3676 -996
tri 3693 -1004 3694 -1003 sw
rect 3693 -1028 3694 -1004
tri 3696 -1005 3733 -968 ne
rect 3733 -996 3738 -968
tri 3738 -996 3764 -970 sw
rect 3848 -986 3857 -952
rect 3848 -996 3876 -986
rect 3733 -1005 3817 -996
tri 3733 -1024 3752 -1005 ne
rect 3752 -1024 3817 -1005
rect 3634 -1050 3694 -1028
rect 3816 -1028 3817 -1024
rect 3834 -1028 3876 -996
rect 3816 -1050 3876 -1028
rect 3722 -1066 3739 -1052
rect 3771 -1066 3788 -1052
tri 3559 -1102 3581 -1080 se
rect 3581 -1087 3596 -1066
tri 3581 -1102 3596 -1087 nw
rect 3915 -1087 3930 -911
tri 3930 -918 3943 -905 nw
rect 4016 -986 4031 -758
tri 3553 -1108 3559 -1102 se
rect 3559 -1108 3568 -1102
rect 3553 -1124 3568 -1108
tri 3568 -1115 3581 -1102 nw
rect 3722 -1110 3739 -1096
rect 3771 -1110 3788 -1096
tri 3915 -1102 3930 -1087 ne
tri 3930 -1102 3952 -1080 sw
rect 3553 -1160 3568 -1152
rect 3634 -1124 3694 -1110
rect 3649 -1134 3694 -1124
rect 3649 -1152 3677 -1134
tri 3553 -1175 3568 -1160 ne
tri 3568 -1175 3590 -1153 sw
rect 3634 -1162 3677 -1152
rect 3692 -1138 3694 -1134
rect 3816 -1124 3876 -1110
tri 3930 -1115 3943 -1102 ne
rect 3943 -1108 3952 -1102
tri 3952 -1108 3958 -1102 sw
rect 3816 -1134 3861 -1124
rect 3692 -1162 3766 -1138
rect 3634 -1166 3766 -1162
tri 3766 -1166 3794 -1138 sw
rect 3816 -1148 3818 -1134
tri 3816 -1150 3818 -1148 ne
rect 3830 -1152 3861 -1134
rect 3830 -1162 3876 -1152
rect 3943 -1123 3958 -1108
tri 3568 -1187 3580 -1175 ne
rect 3580 -1180 3590 -1175
tri 3590 -1180 3595 -1175 sw
rect 3479 -1526 3494 -1298
rect 3580 -1336 3595 -1180
rect 3634 -1222 3662 -1166
tri 3754 -1184 3772 -1166 ne
rect 3772 -1186 3794 -1166
tri 3794 -1186 3814 -1166 sw
tri 3830 -1180 3848 -1162 ne
rect 3653 -1256 3662 -1222
rect 3696 -1195 3738 -1194
rect 3696 -1229 3701 -1195
rect 3731 -1229 3738 -1195
rect 3696 -1238 3738 -1229
rect 3772 -1195 3814 -1186
rect 3772 -1229 3779 -1195
rect 3809 -1229 3814 -1195
rect 3772 -1234 3814 -1229
rect 3848 -1222 3876 -1162
tri 3921 -1175 3943 -1153 se
rect 3943 -1160 3958 -1152
tri 3943 -1175 3958 -1160 nw
tri 3915 -1181 3921 -1175 se
rect 3921 -1181 3930 -1175
rect 3634 -1266 3662 -1256
tri 3662 -1266 3686 -1242 sw
rect 3634 -1298 3676 -1266
tri 3693 -1274 3694 -1273 sw
rect 3693 -1298 3694 -1274
tri 3696 -1275 3733 -1238 ne
rect 3733 -1266 3738 -1238
tri 3738 -1266 3764 -1240 sw
rect 3848 -1256 3857 -1222
rect 3848 -1266 3876 -1256
rect 3733 -1275 3817 -1266
tri 3733 -1294 3752 -1275 ne
rect 3752 -1294 3817 -1275
rect 3634 -1320 3694 -1298
rect 3816 -1298 3817 -1294
rect 3834 -1298 3876 -1266
rect 3816 -1320 3876 -1298
rect 3722 -1336 3739 -1322
rect 3771 -1336 3788 -1322
tri 3559 -1372 3581 -1350 se
rect 3581 -1357 3596 -1336
tri 3581 -1372 3596 -1357 nw
rect 3915 -1357 3930 -1181
tri 3930 -1188 3943 -1175 nw
rect 4016 -1256 4031 -1028
tri 3553 -1378 3559 -1372 se
rect 3559 -1378 3568 -1372
rect 3553 -1394 3568 -1378
tri 3568 -1385 3581 -1372 nw
rect 3722 -1380 3739 -1366
rect 3771 -1380 3788 -1366
tri 3915 -1372 3930 -1357 ne
tri 3930 -1372 3952 -1350 sw
rect 3553 -1430 3568 -1422
rect 3634 -1394 3694 -1380
rect 3649 -1404 3694 -1394
rect 3649 -1422 3677 -1404
tri 3553 -1445 3568 -1430 ne
tri 3568 -1445 3590 -1423 sw
rect 3634 -1432 3677 -1422
rect 3692 -1408 3694 -1404
rect 3816 -1394 3876 -1380
tri 3930 -1385 3943 -1372 ne
rect 3943 -1378 3952 -1372
tri 3952 -1378 3958 -1372 sw
rect 3816 -1404 3861 -1394
rect 3692 -1432 3766 -1408
rect 3634 -1436 3766 -1432
tri 3766 -1436 3794 -1408 sw
rect 3816 -1418 3818 -1404
tri 3816 -1420 3818 -1418 ne
rect 3830 -1422 3861 -1404
rect 3830 -1432 3876 -1422
rect 3943 -1393 3958 -1378
tri 3568 -1457 3580 -1445 ne
rect 3580 -1450 3590 -1445
tri 3590 -1450 3595 -1445 sw
rect 3479 -1796 3494 -1568
rect 3580 -1606 3595 -1450
rect 3634 -1492 3662 -1436
tri 3754 -1454 3772 -1436 ne
rect 3772 -1456 3794 -1436
tri 3794 -1456 3814 -1436 sw
tri 3830 -1450 3848 -1432 ne
rect 3653 -1526 3662 -1492
rect 3696 -1465 3738 -1464
rect 3696 -1499 3701 -1465
rect 3731 -1499 3738 -1465
rect 3696 -1508 3738 -1499
rect 3772 -1465 3814 -1456
rect 3772 -1499 3779 -1465
rect 3809 -1499 3814 -1465
rect 3772 -1504 3814 -1499
rect 3848 -1492 3876 -1432
tri 3921 -1445 3943 -1423 se
rect 3943 -1430 3958 -1422
tri 3943 -1445 3958 -1430 nw
tri 3915 -1451 3921 -1445 se
rect 3921 -1451 3930 -1445
rect 3634 -1536 3662 -1526
tri 3662 -1536 3686 -1512 sw
rect 3634 -1568 3676 -1536
tri 3693 -1544 3694 -1543 sw
rect 3693 -1568 3694 -1544
tri 3696 -1545 3733 -1508 ne
rect 3733 -1536 3738 -1508
tri 3738 -1536 3764 -1510 sw
rect 3848 -1526 3857 -1492
rect 3848 -1536 3876 -1526
rect 3733 -1545 3817 -1536
tri 3733 -1564 3752 -1545 ne
rect 3752 -1564 3817 -1545
rect 3634 -1590 3694 -1568
rect 3816 -1568 3817 -1564
rect 3834 -1568 3876 -1536
rect 3816 -1590 3876 -1568
rect 3722 -1606 3739 -1592
rect 3771 -1606 3788 -1592
tri 3559 -1642 3581 -1620 se
rect 3581 -1627 3596 -1606
tri 3581 -1642 3596 -1627 nw
rect 3915 -1627 3930 -1451
tri 3930 -1458 3943 -1445 nw
rect 4016 -1526 4031 -1298
tri 3553 -1648 3559 -1642 se
rect 3559 -1648 3568 -1642
rect 3553 -1664 3568 -1648
tri 3568 -1655 3581 -1642 nw
rect 3722 -1650 3739 -1636
rect 3771 -1650 3788 -1636
tri 3915 -1642 3930 -1627 ne
tri 3930 -1642 3952 -1620 sw
rect 3553 -1700 3568 -1692
rect 3634 -1664 3694 -1650
rect 3649 -1674 3694 -1664
rect 3649 -1692 3677 -1674
tri 3553 -1715 3568 -1700 ne
tri 3568 -1715 3590 -1693 sw
rect 3634 -1702 3677 -1692
rect 3692 -1678 3694 -1674
rect 3816 -1664 3876 -1650
tri 3930 -1655 3943 -1642 ne
rect 3943 -1648 3952 -1642
tri 3952 -1648 3958 -1642 sw
rect 3816 -1674 3861 -1664
rect 3692 -1702 3766 -1678
rect 3634 -1706 3766 -1702
tri 3766 -1706 3794 -1678 sw
rect 3816 -1688 3818 -1674
tri 3816 -1690 3818 -1688 ne
rect 3830 -1692 3861 -1674
rect 3830 -1702 3876 -1692
rect 3943 -1663 3958 -1648
tri 3568 -1727 3580 -1715 ne
rect 3580 -1720 3590 -1715
tri 3590 -1720 3595 -1715 sw
rect 3479 -2066 3494 -1838
rect 3580 -1876 3595 -1720
rect 3634 -1762 3662 -1706
tri 3754 -1724 3772 -1706 ne
rect 3772 -1726 3794 -1706
tri 3794 -1726 3814 -1706 sw
tri 3830 -1720 3848 -1702 ne
rect 3653 -1796 3662 -1762
rect 3696 -1735 3738 -1734
rect 3696 -1769 3701 -1735
rect 3731 -1769 3738 -1735
rect 3696 -1778 3738 -1769
rect 3772 -1735 3814 -1726
rect 3772 -1769 3779 -1735
rect 3809 -1769 3814 -1735
rect 3772 -1774 3814 -1769
rect 3848 -1762 3876 -1702
tri 3921 -1715 3943 -1693 se
rect 3943 -1700 3958 -1692
tri 3943 -1715 3958 -1700 nw
tri 3915 -1721 3921 -1715 se
rect 3921 -1721 3930 -1715
rect 3634 -1806 3662 -1796
tri 3662 -1806 3686 -1782 sw
rect 3634 -1838 3676 -1806
tri 3693 -1814 3694 -1813 sw
rect 3693 -1838 3694 -1814
tri 3696 -1815 3733 -1778 ne
rect 3733 -1806 3738 -1778
tri 3738 -1806 3764 -1780 sw
rect 3848 -1796 3857 -1762
rect 3848 -1806 3876 -1796
rect 3733 -1815 3817 -1806
tri 3733 -1834 3752 -1815 ne
rect 3752 -1834 3817 -1815
rect 3634 -1860 3694 -1838
rect 3816 -1838 3817 -1834
rect 3834 -1838 3876 -1806
rect 3816 -1860 3876 -1838
rect 3722 -1876 3739 -1862
rect 3771 -1876 3788 -1862
tri 3559 -1912 3581 -1890 se
rect 3581 -1897 3596 -1876
tri 3581 -1912 3596 -1897 nw
rect 3915 -1897 3930 -1721
tri 3930 -1728 3943 -1715 nw
rect 4016 -1796 4031 -1568
tri 3553 -1918 3559 -1912 se
rect 3559 -1918 3568 -1912
rect 3553 -1934 3568 -1918
tri 3568 -1925 3581 -1912 nw
rect 3722 -1920 3739 -1906
rect 3771 -1920 3788 -1906
tri 3915 -1912 3930 -1897 ne
tri 3930 -1912 3952 -1890 sw
rect 3553 -1970 3568 -1962
rect 3634 -1934 3694 -1920
rect 3649 -1944 3694 -1934
rect 3649 -1962 3677 -1944
tri 3553 -1985 3568 -1970 ne
tri 3568 -1985 3590 -1963 sw
rect 3634 -1972 3677 -1962
rect 3692 -1948 3694 -1944
rect 3816 -1934 3876 -1920
tri 3930 -1925 3943 -1912 ne
rect 3943 -1918 3952 -1912
tri 3952 -1918 3958 -1912 sw
rect 3816 -1944 3861 -1934
rect 3692 -1972 3766 -1948
rect 3634 -1976 3766 -1972
tri 3766 -1976 3794 -1948 sw
rect 3816 -1958 3818 -1944
tri 3816 -1960 3818 -1958 ne
rect 3830 -1962 3861 -1944
rect 3830 -1972 3876 -1962
rect 3943 -1933 3958 -1918
tri 3568 -1997 3580 -1985 ne
rect 3580 -1990 3590 -1985
tri 3590 -1990 3595 -1985 sw
rect 3479 -2146 3494 -2108
rect 3580 -2146 3595 -1990
rect 3634 -2032 3662 -1976
tri 3754 -1994 3772 -1976 ne
rect 3772 -1996 3794 -1976
tri 3794 -1996 3814 -1976 sw
tri 3830 -1990 3848 -1972 ne
rect 3653 -2066 3662 -2032
rect 3696 -2005 3738 -2004
rect 3696 -2039 3701 -2005
rect 3731 -2039 3738 -2005
rect 3696 -2048 3738 -2039
rect 3772 -2005 3814 -1996
rect 3772 -2039 3779 -2005
rect 3809 -2039 3814 -2005
rect 3772 -2044 3814 -2039
rect 3848 -2032 3876 -1972
tri 3921 -1985 3943 -1963 se
rect 3943 -1970 3958 -1962
tri 3943 -1985 3958 -1970 nw
tri 3915 -1991 3921 -1985 se
rect 3921 -1991 3930 -1985
rect 3634 -2076 3662 -2066
tri 3662 -2076 3686 -2052 sw
rect 3634 -2108 3676 -2076
tri 3693 -2084 3694 -2083 sw
rect 3693 -2108 3694 -2084
tri 3696 -2085 3733 -2048 ne
rect 3733 -2076 3738 -2048
tri 3738 -2076 3764 -2050 sw
rect 3848 -2066 3857 -2032
rect 3848 -2076 3876 -2066
rect 3733 -2085 3817 -2076
tri 3733 -2104 3752 -2085 ne
rect 3752 -2104 3817 -2085
rect 3634 -2130 3694 -2108
rect 3816 -2108 3817 -2104
rect 3834 -2108 3876 -2076
rect 3816 -2130 3876 -2108
rect 3722 -2146 3739 -2132
rect 3771 -2146 3788 -2132
rect 3915 -2146 3930 -1991
tri 3930 -1998 3943 -1985 nw
rect 4016 -2066 4031 -1838
rect 4016 -2146 4031 -2108
rect 4059 1984 4074 2174
tri 4139 2138 4161 2160 se
rect 4161 2153 4176 2174
tri 4161 2138 4176 2153 nw
rect 4495 2153 4510 2174
tri 4133 2132 4139 2138 se
rect 4139 2132 4148 2138
rect 4133 2116 4148 2132
tri 4148 2125 4161 2138 nw
rect 4302 2130 4319 2144
rect 4351 2130 4368 2144
tri 4495 2138 4510 2153 ne
tri 4510 2138 4532 2160 sw
rect 4133 2080 4148 2088
rect 4214 2116 4274 2130
rect 4229 2106 4274 2116
rect 4229 2088 4257 2106
tri 4133 2065 4148 2080 ne
tri 4148 2065 4170 2087 sw
rect 4214 2078 4257 2088
rect 4272 2102 4274 2106
rect 4396 2116 4456 2130
tri 4510 2125 4523 2138 ne
rect 4523 2132 4532 2138
tri 4532 2132 4538 2138 sw
rect 4396 2106 4441 2116
rect 4272 2078 4346 2102
rect 4214 2074 4346 2078
tri 4346 2074 4374 2102 sw
rect 4396 2092 4398 2106
tri 4396 2090 4398 2092 ne
rect 4410 2088 4441 2106
rect 4410 2078 4456 2088
rect 4523 2117 4538 2132
tri 4148 2053 4160 2065 ne
rect 4160 2060 4170 2065
tri 4170 2060 4175 2065 sw
rect 4059 1714 4074 1942
rect 4160 1904 4175 2060
rect 4214 2018 4242 2074
tri 4334 2056 4352 2074 ne
rect 4352 2054 4374 2074
tri 4374 2054 4394 2074 sw
tri 4410 2060 4428 2078 ne
rect 4233 1984 4242 2018
rect 4276 2045 4318 2046
rect 4276 2011 4281 2045
rect 4311 2011 4318 2045
rect 4276 2002 4318 2011
rect 4352 2045 4394 2054
rect 4352 2011 4359 2045
rect 4389 2011 4394 2045
rect 4352 2006 4394 2011
rect 4428 2018 4456 2078
tri 4501 2065 4523 2087 se
rect 4523 2080 4538 2088
tri 4523 2065 4538 2080 nw
tri 4495 2059 4501 2065 se
rect 4501 2059 4510 2065
rect 4214 1974 4242 1984
tri 4242 1974 4266 1998 sw
rect 4214 1942 4256 1974
tri 4273 1966 4274 1967 sw
rect 4273 1942 4274 1966
tri 4276 1965 4313 2002 ne
rect 4313 1974 4318 2002
tri 4318 1974 4344 2000 sw
rect 4428 1984 4437 2018
rect 4428 1974 4456 1984
rect 4313 1965 4397 1974
tri 4313 1946 4332 1965 ne
rect 4332 1946 4397 1965
rect 4214 1920 4274 1942
rect 4396 1942 4397 1946
rect 4414 1942 4456 1974
rect 4396 1920 4456 1942
rect 4302 1904 4319 1918
rect 4351 1904 4368 1918
tri 4139 1868 4161 1890 se
rect 4161 1883 4176 1904
tri 4161 1868 4176 1883 nw
rect 4495 1883 4510 2059
tri 4510 2052 4523 2065 nw
rect 4596 1984 4611 2174
tri 4133 1862 4139 1868 se
rect 4139 1862 4148 1868
rect 4133 1846 4148 1862
tri 4148 1855 4161 1868 nw
rect 4302 1860 4319 1874
rect 4351 1860 4368 1874
tri 4495 1868 4510 1883 ne
tri 4510 1868 4532 1890 sw
rect 4133 1810 4148 1818
rect 4214 1846 4274 1860
rect 4229 1836 4274 1846
rect 4229 1818 4257 1836
tri 4133 1795 4148 1810 ne
tri 4148 1795 4170 1817 sw
rect 4214 1808 4257 1818
rect 4272 1832 4274 1836
rect 4396 1846 4456 1860
tri 4510 1855 4523 1868 ne
rect 4523 1862 4532 1868
tri 4532 1862 4538 1868 sw
rect 4396 1836 4441 1846
rect 4272 1808 4346 1832
rect 4214 1804 4346 1808
tri 4346 1804 4374 1832 sw
rect 4396 1822 4398 1836
tri 4396 1820 4398 1822 ne
rect 4410 1818 4441 1836
rect 4410 1808 4456 1818
rect 4523 1847 4538 1862
tri 4148 1783 4160 1795 ne
rect 4160 1790 4170 1795
tri 4170 1790 4175 1795 sw
rect 4059 1444 4074 1672
rect 4160 1634 4175 1790
rect 4214 1748 4242 1804
tri 4334 1786 4352 1804 ne
rect 4352 1784 4374 1804
tri 4374 1784 4394 1804 sw
tri 4410 1790 4428 1808 ne
rect 4233 1714 4242 1748
rect 4276 1775 4318 1776
rect 4276 1741 4281 1775
rect 4311 1741 4318 1775
rect 4276 1732 4318 1741
rect 4352 1775 4394 1784
rect 4352 1741 4359 1775
rect 4389 1741 4394 1775
rect 4352 1736 4394 1741
rect 4428 1748 4456 1808
tri 4501 1795 4523 1817 se
rect 4523 1810 4538 1818
tri 4523 1795 4538 1810 nw
tri 4495 1789 4501 1795 se
rect 4501 1789 4510 1795
rect 4214 1704 4242 1714
tri 4242 1704 4266 1728 sw
rect 4214 1672 4256 1704
tri 4273 1696 4274 1697 sw
rect 4273 1672 4274 1696
tri 4276 1695 4313 1732 ne
rect 4313 1704 4318 1732
tri 4318 1704 4344 1730 sw
rect 4428 1714 4437 1748
rect 4428 1704 4456 1714
rect 4313 1695 4397 1704
tri 4313 1676 4332 1695 ne
rect 4332 1676 4397 1695
rect 4214 1650 4274 1672
rect 4396 1672 4397 1676
rect 4414 1672 4456 1704
rect 4396 1650 4456 1672
rect 4302 1634 4319 1648
rect 4351 1634 4368 1648
tri 4139 1598 4161 1620 se
rect 4161 1613 4176 1634
tri 4161 1598 4176 1613 nw
rect 4495 1613 4510 1789
tri 4510 1782 4523 1795 nw
rect 4596 1714 4611 1942
tri 4133 1592 4139 1598 se
rect 4139 1592 4148 1598
rect 4133 1576 4148 1592
tri 4148 1585 4161 1598 nw
rect 4302 1590 4319 1604
rect 4351 1590 4368 1604
tri 4495 1598 4510 1613 ne
tri 4510 1598 4532 1620 sw
rect 4133 1540 4148 1548
rect 4214 1576 4274 1590
rect 4229 1566 4274 1576
rect 4229 1548 4257 1566
tri 4133 1525 4148 1540 ne
tri 4148 1525 4170 1547 sw
rect 4214 1538 4257 1548
rect 4272 1562 4274 1566
rect 4396 1576 4456 1590
tri 4510 1585 4523 1598 ne
rect 4523 1592 4532 1598
tri 4532 1592 4538 1598 sw
rect 4396 1566 4441 1576
rect 4272 1538 4346 1562
rect 4214 1534 4346 1538
tri 4346 1534 4374 1562 sw
rect 4396 1552 4398 1566
tri 4396 1550 4398 1552 ne
rect 4410 1548 4441 1566
rect 4410 1538 4456 1548
rect 4523 1577 4538 1592
tri 4148 1513 4160 1525 ne
rect 4160 1520 4170 1525
tri 4170 1520 4175 1525 sw
rect 4059 1174 4074 1402
rect 4160 1364 4175 1520
rect 4214 1478 4242 1534
tri 4334 1516 4352 1534 ne
rect 4352 1514 4374 1534
tri 4374 1514 4394 1534 sw
tri 4410 1520 4428 1538 ne
rect 4233 1444 4242 1478
rect 4276 1505 4318 1506
rect 4276 1471 4281 1505
rect 4311 1471 4318 1505
rect 4276 1462 4318 1471
rect 4352 1505 4394 1514
rect 4352 1471 4359 1505
rect 4389 1471 4394 1505
rect 4352 1466 4394 1471
rect 4428 1478 4456 1538
tri 4501 1525 4523 1547 se
rect 4523 1540 4538 1548
tri 4523 1525 4538 1540 nw
tri 4495 1519 4501 1525 se
rect 4501 1519 4510 1525
rect 4214 1434 4242 1444
tri 4242 1434 4266 1458 sw
rect 4214 1402 4256 1434
tri 4273 1426 4274 1427 sw
rect 4273 1402 4274 1426
tri 4276 1425 4313 1462 ne
rect 4313 1434 4318 1462
tri 4318 1434 4344 1460 sw
rect 4428 1444 4437 1478
rect 4428 1434 4456 1444
rect 4313 1425 4397 1434
tri 4313 1406 4332 1425 ne
rect 4332 1406 4397 1425
rect 4214 1380 4274 1402
rect 4396 1402 4397 1406
rect 4414 1402 4456 1434
rect 4396 1380 4456 1402
rect 4302 1364 4319 1378
rect 4351 1364 4368 1378
tri 4139 1328 4161 1350 se
rect 4161 1343 4176 1364
tri 4161 1328 4176 1343 nw
rect 4495 1343 4510 1519
tri 4510 1512 4523 1525 nw
rect 4596 1444 4611 1672
tri 4133 1322 4139 1328 se
rect 4139 1322 4148 1328
rect 4133 1306 4148 1322
tri 4148 1315 4161 1328 nw
rect 4302 1320 4319 1334
rect 4351 1320 4368 1334
tri 4495 1328 4510 1343 ne
tri 4510 1328 4532 1350 sw
rect 4133 1270 4148 1278
rect 4214 1306 4274 1320
rect 4229 1296 4274 1306
rect 4229 1278 4257 1296
tri 4133 1255 4148 1270 ne
tri 4148 1255 4170 1277 sw
rect 4214 1268 4257 1278
rect 4272 1292 4274 1296
rect 4396 1306 4456 1320
tri 4510 1315 4523 1328 ne
rect 4523 1322 4532 1328
tri 4532 1322 4538 1328 sw
rect 4396 1296 4441 1306
rect 4272 1268 4346 1292
rect 4214 1264 4346 1268
tri 4346 1264 4374 1292 sw
rect 4396 1282 4398 1296
tri 4396 1280 4398 1282 ne
rect 4410 1278 4441 1296
rect 4410 1268 4456 1278
rect 4523 1307 4538 1322
tri 4148 1243 4160 1255 ne
rect 4160 1250 4170 1255
tri 4170 1250 4175 1255 sw
rect 4059 904 4074 1132
rect 4160 1094 4175 1250
rect 4214 1208 4242 1264
tri 4334 1246 4352 1264 ne
rect 4352 1244 4374 1264
tri 4374 1244 4394 1264 sw
tri 4410 1250 4428 1268 ne
rect 4233 1174 4242 1208
rect 4276 1235 4318 1236
rect 4276 1201 4281 1235
rect 4311 1201 4318 1235
rect 4276 1192 4318 1201
rect 4352 1235 4394 1244
rect 4352 1201 4359 1235
rect 4389 1201 4394 1235
rect 4352 1196 4394 1201
rect 4428 1208 4456 1268
tri 4501 1255 4523 1277 se
rect 4523 1270 4538 1278
tri 4523 1255 4538 1270 nw
tri 4495 1249 4501 1255 se
rect 4501 1249 4510 1255
rect 4214 1164 4242 1174
tri 4242 1164 4266 1188 sw
rect 4214 1132 4256 1164
tri 4273 1156 4274 1157 sw
rect 4273 1132 4274 1156
tri 4276 1155 4313 1192 ne
rect 4313 1164 4318 1192
tri 4318 1164 4344 1190 sw
rect 4428 1174 4437 1208
rect 4428 1164 4456 1174
rect 4313 1155 4397 1164
tri 4313 1136 4332 1155 ne
rect 4332 1136 4397 1155
rect 4214 1110 4274 1132
rect 4396 1132 4397 1136
rect 4414 1132 4456 1164
rect 4396 1110 4456 1132
rect 4302 1094 4319 1108
rect 4351 1094 4368 1108
tri 4139 1058 4161 1080 se
rect 4161 1073 4176 1094
tri 4161 1058 4176 1073 nw
rect 4495 1073 4510 1249
tri 4510 1242 4523 1255 nw
rect 4596 1174 4611 1402
tri 4133 1052 4139 1058 se
rect 4139 1052 4148 1058
rect 4133 1036 4148 1052
tri 4148 1045 4161 1058 nw
rect 4302 1050 4319 1064
rect 4351 1050 4368 1064
tri 4495 1058 4510 1073 ne
tri 4510 1058 4532 1080 sw
rect 4133 1000 4148 1008
rect 4214 1036 4274 1050
rect 4229 1026 4274 1036
rect 4229 1008 4257 1026
tri 4133 985 4148 1000 ne
tri 4148 985 4170 1007 sw
rect 4214 998 4257 1008
rect 4272 1022 4274 1026
rect 4396 1036 4456 1050
tri 4510 1045 4523 1058 ne
rect 4523 1052 4532 1058
tri 4532 1052 4538 1058 sw
rect 4396 1026 4441 1036
rect 4272 998 4346 1022
rect 4214 994 4346 998
tri 4346 994 4374 1022 sw
rect 4396 1012 4398 1026
tri 4396 1010 4398 1012 ne
rect 4410 1008 4441 1026
rect 4410 998 4456 1008
rect 4523 1037 4538 1052
tri 4148 973 4160 985 ne
rect 4160 980 4170 985
tri 4170 980 4175 985 sw
rect 4059 634 4074 862
rect 4160 824 4175 980
rect 4214 938 4242 994
tri 4334 976 4352 994 ne
rect 4352 974 4374 994
tri 4374 974 4394 994 sw
tri 4410 980 4428 998 ne
rect 4233 904 4242 938
rect 4276 965 4318 966
rect 4276 931 4281 965
rect 4311 931 4318 965
rect 4276 922 4318 931
rect 4352 965 4394 974
rect 4352 931 4359 965
rect 4389 931 4394 965
rect 4352 926 4394 931
rect 4428 938 4456 998
tri 4501 985 4523 1007 se
rect 4523 1000 4538 1008
tri 4523 985 4538 1000 nw
tri 4495 979 4501 985 se
rect 4501 979 4510 985
rect 4214 894 4242 904
tri 4242 894 4266 918 sw
rect 4214 862 4256 894
tri 4273 886 4274 887 sw
rect 4273 862 4274 886
tri 4276 885 4313 922 ne
rect 4313 894 4318 922
tri 4318 894 4344 920 sw
rect 4428 904 4437 938
rect 4428 894 4456 904
rect 4313 885 4397 894
tri 4313 866 4332 885 ne
rect 4332 866 4397 885
rect 4214 840 4274 862
rect 4396 862 4397 866
rect 4414 862 4456 894
rect 4396 840 4456 862
rect 4302 824 4319 838
rect 4351 824 4368 838
tri 4139 788 4161 810 se
rect 4161 803 4176 824
tri 4161 788 4176 803 nw
rect 4495 803 4510 979
tri 4510 972 4523 985 nw
rect 4596 904 4611 1132
tri 4133 782 4139 788 se
rect 4139 782 4148 788
rect 4133 766 4148 782
tri 4148 775 4161 788 nw
rect 4302 780 4319 794
rect 4351 780 4368 794
tri 4495 788 4510 803 ne
tri 4510 788 4532 810 sw
rect 4133 730 4148 738
rect 4214 766 4274 780
rect 4229 756 4274 766
rect 4229 738 4257 756
tri 4133 715 4148 730 ne
tri 4148 715 4170 737 sw
rect 4214 728 4257 738
rect 4272 752 4274 756
rect 4396 766 4456 780
tri 4510 775 4523 788 ne
rect 4523 782 4532 788
tri 4532 782 4538 788 sw
rect 4396 756 4441 766
rect 4272 728 4346 752
rect 4214 724 4346 728
tri 4346 724 4374 752 sw
rect 4396 742 4398 756
tri 4396 740 4398 742 ne
rect 4410 738 4441 756
rect 4410 728 4456 738
rect 4523 767 4538 782
tri 4148 703 4160 715 ne
rect 4160 710 4170 715
tri 4170 710 4175 715 sw
rect 4059 364 4074 592
rect 4160 554 4175 710
rect 4214 668 4242 724
tri 4334 706 4352 724 ne
rect 4352 704 4374 724
tri 4374 704 4394 724 sw
tri 4410 710 4428 728 ne
rect 4233 634 4242 668
rect 4276 695 4318 696
rect 4276 661 4281 695
rect 4311 661 4318 695
rect 4276 652 4318 661
rect 4352 695 4394 704
rect 4352 661 4359 695
rect 4389 661 4394 695
rect 4352 656 4394 661
rect 4428 668 4456 728
tri 4501 715 4523 737 se
rect 4523 730 4538 738
tri 4523 715 4538 730 nw
tri 4495 709 4501 715 se
rect 4501 709 4510 715
rect 4214 624 4242 634
tri 4242 624 4266 648 sw
rect 4214 592 4256 624
tri 4273 616 4274 617 sw
rect 4273 592 4274 616
tri 4276 615 4313 652 ne
rect 4313 624 4318 652
tri 4318 624 4344 650 sw
rect 4428 634 4437 668
rect 4428 624 4456 634
rect 4313 615 4397 624
tri 4313 596 4332 615 ne
rect 4332 596 4397 615
rect 4214 570 4274 592
rect 4396 592 4397 596
rect 4414 592 4456 624
rect 4396 570 4456 592
rect 4302 554 4319 568
rect 4351 554 4368 568
tri 4139 518 4161 540 se
rect 4161 533 4176 554
tri 4161 518 4176 533 nw
rect 4495 533 4510 709
tri 4510 702 4523 715 nw
rect 4596 634 4611 862
tri 4133 512 4139 518 se
rect 4139 512 4148 518
rect 4133 496 4148 512
tri 4148 505 4161 518 nw
rect 4302 510 4319 524
rect 4351 510 4368 524
tri 4495 518 4510 533 ne
tri 4510 518 4532 540 sw
rect 4133 460 4148 468
rect 4214 496 4274 510
rect 4229 486 4274 496
rect 4229 468 4257 486
tri 4133 445 4148 460 ne
tri 4148 445 4170 467 sw
rect 4214 458 4257 468
rect 4272 482 4274 486
rect 4396 496 4456 510
tri 4510 505 4523 518 ne
rect 4523 512 4532 518
tri 4532 512 4538 518 sw
rect 4396 486 4441 496
rect 4272 458 4346 482
rect 4214 454 4346 458
tri 4346 454 4374 482 sw
rect 4396 472 4398 486
tri 4396 470 4398 472 ne
rect 4410 468 4441 486
rect 4410 458 4456 468
rect 4523 497 4538 512
tri 4148 433 4160 445 ne
rect 4160 440 4170 445
tri 4170 440 4175 445 sw
rect 4059 94 4074 322
rect 4160 284 4175 440
rect 4214 398 4242 454
tri 4334 436 4352 454 ne
rect 4352 434 4374 454
tri 4374 434 4394 454 sw
tri 4410 440 4428 458 ne
rect 4233 364 4242 398
rect 4276 425 4318 426
rect 4276 391 4281 425
rect 4311 391 4318 425
rect 4276 382 4318 391
rect 4352 425 4394 434
rect 4352 391 4359 425
rect 4389 391 4394 425
rect 4352 386 4394 391
rect 4428 398 4456 458
tri 4501 445 4523 467 se
rect 4523 460 4538 468
tri 4523 445 4538 460 nw
tri 4495 439 4501 445 se
rect 4501 439 4510 445
rect 4214 354 4242 364
tri 4242 354 4266 378 sw
rect 4214 322 4256 354
tri 4273 346 4274 347 sw
rect 4273 322 4274 346
tri 4276 345 4313 382 ne
rect 4313 354 4318 382
tri 4318 354 4344 380 sw
rect 4428 364 4437 398
rect 4428 354 4456 364
rect 4313 345 4397 354
tri 4313 326 4332 345 ne
rect 4332 326 4397 345
rect 4214 300 4274 322
rect 4396 322 4397 326
rect 4414 322 4456 354
rect 4396 300 4456 322
rect 4302 284 4319 298
rect 4351 284 4368 298
tri 4139 248 4161 270 se
rect 4161 263 4176 284
tri 4161 248 4176 263 nw
rect 4495 263 4510 439
tri 4510 432 4523 445 nw
rect 4596 364 4611 592
tri 4133 242 4139 248 se
rect 4139 242 4148 248
rect 4133 226 4148 242
tri 4148 235 4161 248 nw
rect 4302 240 4319 254
rect 4351 240 4368 254
tri 4495 248 4510 263 ne
tri 4510 248 4532 270 sw
rect 4133 190 4148 198
rect 4214 226 4274 240
rect 4229 216 4274 226
rect 4229 198 4257 216
tri 4133 175 4148 190 ne
tri 4148 175 4170 197 sw
rect 4214 188 4257 198
rect 4272 212 4274 216
rect 4396 226 4456 240
tri 4510 235 4523 248 ne
rect 4523 242 4532 248
tri 4532 242 4538 248 sw
rect 4396 216 4441 226
rect 4272 188 4346 212
rect 4214 184 4346 188
tri 4346 184 4374 212 sw
rect 4396 202 4398 216
tri 4396 200 4398 202 ne
rect 4410 198 4441 216
rect 4410 188 4456 198
rect 4523 227 4538 242
tri 4148 163 4160 175 ne
rect 4160 170 4170 175
tri 4170 170 4175 175 sw
rect 4059 -176 4074 52
rect 4160 14 4175 170
rect 4214 128 4242 184
tri 4334 166 4352 184 ne
rect 4352 164 4374 184
tri 4374 164 4394 184 sw
tri 4410 170 4428 188 ne
rect 4233 94 4242 128
rect 4276 155 4318 156
rect 4276 121 4281 155
rect 4311 121 4318 155
rect 4276 112 4318 121
rect 4352 155 4394 164
rect 4352 121 4359 155
rect 4389 121 4394 155
rect 4352 116 4394 121
rect 4428 128 4456 188
tri 4501 175 4523 197 se
rect 4523 190 4538 198
tri 4523 175 4538 190 nw
tri 4495 169 4501 175 se
rect 4501 169 4510 175
rect 4214 84 4242 94
tri 4242 84 4266 108 sw
rect 4214 52 4256 84
tri 4273 76 4274 77 sw
rect 4273 52 4274 76
tri 4276 75 4313 112 ne
rect 4313 84 4318 112
tri 4318 84 4344 110 sw
rect 4428 94 4437 128
rect 4428 84 4456 94
rect 4313 75 4397 84
tri 4313 56 4332 75 ne
rect 4332 56 4397 75
rect 4214 30 4274 52
rect 4396 52 4397 56
rect 4414 52 4456 84
rect 4396 30 4456 52
rect 4302 14 4319 28
rect 4351 14 4368 28
tri 4139 -22 4161 0 se
rect 4161 -7 4176 14
tri 4161 -22 4176 -7 nw
rect 4495 -7 4510 169
tri 4510 162 4523 175 nw
rect 4596 94 4611 322
tri 4133 -28 4139 -22 se
rect 4139 -28 4148 -22
rect 4133 -44 4148 -28
tri 4148 -35 4161 -22 nw
rect 4302 -30 4319 -16
rect 4351 -30 4368 -16
tri 4495 -22 4510 -7 ne
tri 4510 -22 4532 0 sw
rect 4133 -80 4148 -72
rect 4214 -44 4274 -30
rect 4229 -54 4274 -44
rect 4229 -72 4257 -54
tri 4133 -95 4148 -80 ne
tri 4148 -95 4170 -73 sw
rect 4214 -82 4257 -72
rect 4272 -58 4274 -54
rect 4396 -44 4456 -30
tri 4510 -35 4523 -22 ne
rect 4523 -28 4532 -22
tri 4532 -28 4538 -22 sw
rect 4396 -54 4441 -44
rect 4272 -82 4346 -58
rect 4214 -86 4346 -82
tri 4346 -86 4374 -58 sw
rect 4396 -68 4398 -54
tri 4396 -70 4398 -68 ne
rect 4410 -72 4441 -54
rect 4410 -82 4456 -72
rect 4523 -43 4538 -28
tri 4148 -107 4160 -95 ne
rect 4160 -100 4170 -95
tri 4170 -100 4175 -95 sw
rect 4059 -446 4074 -218
rect 4160 -256 4175 -100
rect 4214 -142 4242 -86
tri 4334 -104 4352 -86 ne
rect 4352 -106 4374 -86
tri 4374 -106 4394 -86 sw
tri 4410 -100 4428 -82 ne
rect 4233 -176 4242 -142
rect 4276 -115 4318 -114
rect 4276 -149 4281 -115
rect 4311 -149 4318 -115
rect 4276 -158 4318 -149
rect 4352 -115 4394 -106
rect 4352 -149 4359 -115
rect 4389 -149 4394 -115
rect 4352 -154 4394 -149
rect 4428 -142 4456 -82
tri 4501 -95 4523 -73 se
rect 4523 -80 4538 -72
tri 4523 -95 4538 -80 nw
tri 4495 -101 4501 -95 se
rect 4501 -101 4510 -95
rect 4214 -186 4242 -176
tri 4242 -186 4266 -162 sw
rect 4214 -218 4256 -186
tri 4273 -194 4274 -193 sw
rect 4273 -218 4274 -194
tri 4276 -195 4313 -158 ne
rect 4313 -186 4318 -158
tri 4318 -186 4344 -160 sw
rect 4428 -176 4437 -142
rect 4428 -186 4456 -176
rect 4313 -195 4397 -186
tri 4313 -214 4332 -195 ne
rect 4332 -214 4397 -195
rect 4214 -240 4274 -218
rect 4396 -218 4397 -214
rect 4414 -218 4456 -186
rect 4396 -240 4456 -218
rect 4302 -256 4319 -242
rect 4351 -256 4368 -242
tri 4139 -292 4161 -270 se
rect 4161 -277 4176 -256
tri 4161 -292 4176 -277 nw
rect 4495 -277 4510 -101
tri 4510 -108 4523 -95 nw
rect 4596 -176 4611 52
tri 4133 -298 4139 -292 se
rect 4139 -298 4148 -292
rect 4133 -314 4148 -298
tri 4148 -305 4161 -292 nw
rect 4302 -300 4319 -286
rect 4351 -300 4368 -286
tri 4495 -292 4510 -277 ne
tri 4510 -292 4532 -270 sw
rect 4133 -350 4148 -342
rect 4214 -314 4274 -300
rect 4229 -324 4274 -314
rect 4229 -342 4257 -324
tri 4133 -365 4148 -350 ne
tri 4148 -365 4170 -343 sw
rect 4214 -352 4257 -342
rect 4272 -328 4274 -324
rect 4396 -314 4456 -300
tri 4510 -305 4523 -292 ne
rect 4523 -298 4532 -292
tri 4532 -298 4538 -292 sw
rect 4396 -324 4441 -314
rect 4272 -352 4346 -328
rect 4214 -356 4346 -352
tri 4346 -356 4374 -328 sw
rect 4396 -338 4398 -324
tri 4396 -340 4398 -338 ne
rect 4410 -342 4441 -324
rect 4410 -352 4456 -342
rect 4523 -313 4538 -298
tri 4148 -377 4160 -365 ne
rect 4160 -370 4170 -365
tri 4170 -370 4175 -365 sw
rect 4059 -716 4074 -488
rect 4160 -526 4175 -370
rect 4214 -412 4242 -356
tri 4334 -374 4352 -356 ne
rect 4352 -376 4374 -356
tri 4374 -376 4394 -356 sw
tri 4410 -370 4428 -352 ne
rect 4233 -446 4242 -412
rect 4276 -385 4318 -384
rect 4276 -419 4281 -385
rect 4311 -419 4318 -385
rect 4276 -428 4318 -419
rect 4352 -385 4394 -376
rect 4352 -419 4359 -385
rect 4389 -419 4394 -385
rect 4352 -424 4394 -419
rect 4428 -412 4456 -352
tri 4501 -365 4523 -343 se
rect 4523 -350 4538 -342
tri 4523 -365 4538 -350 nw
tri 4495 -371 4501 -365 se
rect 4501 -371 4510 -365
rect 4214 -456 4242 -446
tri 4242 -456 4266 -432 sw
rect 4214 -488 4256 -456
tri 4273 -464 4274 -463 sw
rect 4273 -488 4274 -464
tri 4276 -465 4313 -428 ne
rect 4313 -456 4318 -428
tri 4318 -456 4344 -430 sw
rect 4428 -446 4437 -412
rect 4428 -456 4456 -446
rect 4313 -465 4397 -456
tri 4313 -484 4332 -465 ne
rect 4332 -484 4397 -465
rect 4214 -510 4274 -488
rect 4396 -488 4397 -484
rect 4414 -488 4456 -456
rect 4396 -510 4456 -488
rect 4302 -526 4319 -512
rect 4351 -526 4368 -512
tri 4139 -562 4161 -540 se
rect 4161 -547 4176 -526
tri 4161 -562 4176 -547 nw
rect 4495 -547 4510 -371
tri 4510 -378 4523 -365 nw
rect 4596 -446 4611 -218
tri 4133 -568 4139 -562 se
rect 4139 -568 4148 -562
rect 4133 -584 4148 -568
tri 4148 -575 4161 -562 nw
rect 4302 -570 4319 -556
rect 4351 -570 4368 -556
tri 4495 -562 4510 -547 ne
tri 4510 -562 4532 -540 sw
rect 4133 -620 4148 -612
rect 4214 -584 4274 -570
rect 4229 -594 4274 -584
rect 4229 -612 4257 -594
tri 4133 -635 4148 -620 ne
tri 4148 -635 4170 -613 sw
rect 4214 -622 4257 -612
rect 4272 -598 4274 -594
rect 4396 -584 4456 -570
tri 4510 -575 4523 -562 ne
rect 4523 -568 4532 -562
tri 4532 -568 4538 -562 sw
rect 4396 -594 4441 -584
rect 4272 -622 4346 -598
rect 4214 -626 4346 -622
tri 4346 -626 4374 -598 sw
rect 4396 -608 4398 -594
tri 4396 -610 4398 -608 ne
rect 4410 -612 4441 -594
rect 4410 -622 4456 -612
rect 4523 -583 4538 -568
tri 4148 -647 4160 -635 ne
rect 4160 -640 4170 -635
tri 4170 -640 4175 -635 sw
rect 4059 -986 4074 -758
rect 4160 -796 4175 -640
rect 4214 -682 4242 -626
tri 4334 -644 4352 -626 ne
rect 4352 -646 4374 -626
tri 4374 -646 4394 -626 sw
tri 4410 -640 4428 -622 ne
rect 4233 -716 4242 -682
rect 4276 -655 4318 -654
rect 4276 -689 4281 -655
rect 4311 -689 4318 -655
rect 4276 -698 4318 -689
rect 4352 -655 4394 -646
rect 4352 -689 4359 -655
rect 4389 -689 4394 -655
rect 4352 -694 4394 -689
rect 4428 -682 4456 -622
tri 4501 -635 4523 -613 se
rect 4523 -620 4538 -612
tri 4523 -635 4538 -620 nw
tri 4495 -641 4501 -635 se
rect 4501 -641 4510 -635
rect 4214 -726 4242 -716
tri 4242 -726 4266 -702 sw
rect 4214 -758 4256 -726
tri 4273 -734 4274 -733 sw
rect 4273 -758 4274 -734
tri 4276 -735 4313 -698 ne
rect 4313 -726 4318 -698
tri 4318 -726 4344 -700 sw
rect 4428 -716 4437 -682
rect 4428 -726 4456 -716
rect 4313 -735 4397 -726
tri 4313 -754 4332 -735 ne
rect 4332 -754 4397 -735
rect 4214 -780 4274 -758
rect 4396 -758 4397 -754
rect 4414 -758 4456 -726
rect 4396 -780 4456 -758
rect 4302 -796 4319 -782
rect 4351 -796 4368 -782
tri 4139 -832 4161 -810 se
rect 4161 -817 4176 -796
tri 4161 -832 4176 -817 nw
rect 4495 -817 4510 -641
tri 4510 -648 4523 -635 nw
rect 4596 -716 4611 -488
tri 4133 -838 4139 -832 se
rect 4139 -838 4148 -832
rect 4133 -854 4148 -838
tri 4148 -845 4161 -832 nw
rect 4302 -840 4319 -826
rect 4351 -840 4368 -826
tri 4495 -832 4510 -817 ne
tri 4510 -832 4532 -810 sw
rect 4133 -890 4148 -882
rect 4214 -854 4274 -840
rect 4229 -864 4274 -854
rect 4229 -882 4257 -864
tri 4133 -905 4148 -890 ne
tri 4148 -905 4170 -883 sw
rect 4214 -892 4257 -882
rect 4272 -868 4274 -864
rect 4396 -854 4456 -840
tri 4510 -845 4523 -832 ne
rect 4523 -838 4532 -832
tri 4532 -838 4538 -832 sw
rect 4396 -864 4441 -854
rect 4272 -892 4346 -868
rect 4214 -896 4346 -892
tri 4346 -896 4374 -868 sw
rect 4396 -878 4398 -864
tri 4396 -880 4398 -878 ne
rect 4410 -882 4441 -864
rect 4410 -892 4456 -882
rect 4523 -853 4538 -838
tri 4148 -917 4160 -905 ne
rect 4160 -910 4170 -905
tri 4170 -910 4175 -905 sw
rect 4059 -1256 4074 -1028
rect 4160 -1066 4175 -910
rect 4214 -952 4242 -896
tri 4334 -914 4352 -896 ne
rect 4352 -916 4374 -896
tri 4374 -916 4394 -896 sw
tri 4410 -910 4428 -892 ne
rect 4233 -986 4242 -952
rect 4276 -925 4318 -924
rect 4276 -959 4281 -925
rect 4311 -959 4318 -925
rect 4276 -968 4318 -959
rect 4352 -925 4394 -916
rect 4352 -959 4359 -925
rect 4389 -959 4394 -925
rect 4352 -964 4394 -959
rect 4428 -952 4456 -892
tri 4501 -905 4523 -883 se
rect 4523 -890 4538 -882
tri 4523 -905 4538 -890 nw
tri 4495 -911 4501 -905 se
rect 4501 -911 4510 -905
rect 4214 -996 4242 -986
tri 4242 -996 4266 -972 sw
rect 4214 -1028 4256 -996
tri 4273 -1004 4274 -1003 sw
rect 4273 -1028 4274 -1004
tri 4276 -1005 4313 -968 ne
rect 4313 -996 4318 -968
tri 4318 -996 4344 -970 sw
rect 4428 -986 4437 -952
rect 4428 -996 4456 -986
rect 4313 -1005 4397 -996
tri 4313 -1024 4332 -1005 ne
rect 4332 -1024 4397 -1005
rect 4214 -1050 4274 -1028
rect 4396 -1028 4397 -1024
rect 4414 -1028 4456 -996
rect 4396 -1050 4456 -1028
rect 4302 -1066 4319 -1052
rect 4351 -1066 4368 -1052
tri 4139 -1102 4161 -1080 se
rect 4161 -1087 4176 -1066
tri 4161 -1102 4176 -1087 nw
rect 4495 -1087 4510 -911
tri 4510 -918 4523 -905 nw
rect 4596 -986 4611 -758
tri 4133 -1108 4139 -1102 se
rect 4139 -1108 4148 -1102
rect 4133 -1124 4148 -1108
tri 4148 -1115 4161 -1102 nw
rect 4302 -1110 4319 -1096
rect 4351 -1110 4368 -1096
tri 4495 -1102 4510 -1087 ne
tri 4510 -1102 4532 -1080 sw
rect 4133 -1160 4148 -1152
rect 4214 -1124 4274 -1110
rect 4229 -1134 4274 -1124
rect 4229 -1152 4257 -1134
tri 4133 -1175 4148 -1160 ne
tri 4148 -1175 4170 -1153 sw
rect 4214 -1162 4257 -1152
rect 4272 -1138 4274 -1134
rect 4396 -1124 4456 -1110
tri 4510 -1115 4523 -1102 ne
rect 4523 -1108 4532 -1102
tri 4532 -1108 4538 -1102 sw
rect 4396 -1134 4441 -1124
rect 4272 -1162 4346 -1138
rect 4214 -1166 4346 -1162
tri 4346 -1166 4374 -1138 sw
rect 4396 -1148 4398 -1134
tri 4396 -1150 4398 -1148 ne
rect 4410 -1152 4441 -1134
rect 4410 -1162 4456 -1152
rect 4523 -1123 4538 -1108
tri 4148 -1187 4160 -1175 ne
rect 4160 -1180 4170 -1175
tri 4170 -1180 4175 -1175 sw
rect 4059 -1526 4074 -1298
rect 4160 -1336 4175 -1180
rect 4214 -1222 4242 -1166
tri 4334 -1184 4352 -1166 ne
rect 4352 -1186 4374 -1166
tri 4374 -1186 4394 -1166 sw
tri 4410 -1180 4428 -1162 ne
rect 4233 -1256 4242 -1222
rect 4276 -1195 4318 -1194
rect 4276 -1229 4281 -1195
rect 4311 -1229 4318 -1195
rect 4276 -1238 4318 -1229
rect 4352 -1195 4394 -1186
rect 4352 -1229 4359 -1195
rect 4389 -1229 4394 -1195
rect 4352 -1234 4394 -1229
rect 4428 -1222 4456 -1162
tri 4501 -1175 4523 -1153 se
rect 4523 -1160 4538 -1152
tri 4523 -1175 4538 -1160 nw
tri 4495 -1181 4501 -1175 se
rect 4501 -1181 4510 -1175
rect 4214 -1266 4242 -1256
tri 4242 -1266 4266 -1242 sw
rect 4214 -1298 4256 -1266
tri 4273 -1274 4274 -1273 sw
rect 4273 -1298 4274 -1274
tri 4276 -1275 4313 -1238 ne
rect 4313 -1266 4318 -1238
tri 4318 -1266 4344 -1240 sw
rect 4428 -1256 4437 -1222
rect 4428 -1266 4456 -1256
rect 4313 -1275 4397 -1266
tri 4313 -1294 4332 -1275 ne
rect 4332 -1294 4397 -1275
rect 4214 -1320 4274 -1298
rect 4396 -1298 4397 -1294
rect 4414 -1298 4456 -1266
rect 4396 -1320 4456 -1298
rect 4302 -1336 4319 -1322
rect 4351 -1336 4368 -1322
tri 4139 -1372 4161 -1350 se
rect 4161 -1357 4176 -1336
tri 4161 -1372 4176 -1357 nw
rect 4495 -1357 4510 -1181
tri 4510 -1188 4523 -1175 nw
rect 4596 -1256 4611 -1028
tri 4133 -1378 4139 -1372 se
rect 4139 -1378 4148 -1372
rect 4133 -1394 4148 -1378
tri 4148 -1385 4161 -1372 nw
rect 4302 -1380 4319 -1366
rect 4351 -1380 4368 -1366
tri 4495 -1372 4510 -1357 ne
tri 4510 -1372 4532 -1350 sw
rect 4133 -1430 4148 -1422
rect 4214 -1394 4274 -1380
rect 4229 -1404 4274 -1394
rect 4229 -1422 4257 -1404
tri 4133 -1445 4148 -1430 ne
tri 4148 -1445 4170 -1423 sw
rect 4214 -1432 4257 -1422
rect 4272 -1408 4274 -1404
rect 4396 -1394 4456 -1380
tri 4510 -1385 4523 -1372 ne
rect 4523 -1378 4532 -1372
tri 4532 -1378 4538 -1372 sw
rect 4396 -1404 4441 -1394
rect 4272 -1432 4346 -1408
rect 4214 -1436 4346 -1432
tri 4346 -1436 4374 -1408 sw
rect 4396 -1418 4398 -1404
tri 4396 -1420 4398 -1418 ne
rect 4410 -1422 4441 -1404
rect 4410 -1432 4456 -1422
rect 4523 -1393 4538 -1378
tri 4148 -1457 4160 -1445 ne
rect 4160 -1450 4170 -1445
tri 4170 -1450 4175 -1445 sw
rect 4059 -1796 4074 -1568
rect 4160 -1606 4175 -1450
rect 4214 -1492 4242 -1436
tri 4334 -1454 4352 -1436 ne
rect 4352 -1456 4374 -1436
tri 4374 -1456 4394 -1436 sw
tri 4410 -1450 4428 -1432 ne
rect 4233 -1526 4242 -1492
rect 4276 -1465 4318 -1464
rect 4276 -1499 4281 -1465
rect 4311 -1499 4318 -1465
rect 4276 -1508 4318 -1499
rect 4352 -1465 4394 -1456
rect 4352 -1499 4359 -1465
rect 4389 -1499 4394 -1465
rect 4352 -1504 4394 -1499
rect 4428 -1492 4456 -1432
tri 4501 -1445 4523 -1423 se
rect 4523 -1430 4538 -1422
tri 4523 -1445 4538 -1430 nw
tri 4495 -1451 4501 -1445 se
rect 4501 -1451 4510 -1445
rect 4214 -1536 4242 -1526
tri 4242 -1536 4266 -1512 sw
rect 4214 -1568 4256 -1536
tri 4273 -1544 4274 -1543 sw
rect 4273 -1568 4274 -1544
tri 4276 -1545 4313 -1508 ne
rect 4313 -1536 4318 -1508
tri 4318 -1536 4344 -1510 sw
rect 4428 -1526 4437 -1492
rect 4428 -1536 4456 -1526
rect 4313 -1545 4397 -1536
tri 4313 -1564 4332 -1545 ne
rect 4332 -1564 4397 -1545
rect 4214 -1590 4274 -1568
rect 4396 -1568 4397 -1564
rect 4414 -1568 4456 -1536
rect 4396 -1590 4456 -1568
rect 4302 -1606 4319 -1592
rect 4351 -1606 4368 -1592
tri 4139 -1642 4161 -1620 se
rect 4161 -1627 4176 -1606
tri 4161 -1642 4176 -1627 nw
rect 4495 -1627 4510 -1451
tri 4510 -1458 4523 -1445 nw
rect 4596 -1526 4611 -1298
tri 4133 -1648 4139 -1642 se
rect 4139 -1648 4148 -1642
rect 4133 -1664 4148 -1648
tri 4148 -1655 4161 -1642 nw
rect 4302 -1650 4319 -1636
rect 4351 -1650 4368 -1636
tri 4495 -1642 4510 -1627 ne
tri 4510 -1642 4532 -1620 sw
rect 4133 -1700 4148 -1692
rect 4214 -1664 4274 -1650
rect 4229 -1674 4274 -1664
rect 4229 -1692 4257 -1674
tri 4133 -1715 4148 -1700 ne
tri 4148 -1715 4170 -1693 sw
rect 4214 -1702 4257 -1692
rect 4272 -1678 4274 -1674
rect 4396 -1664 4456 -1650
tri 4510 -1655 4523 -1642 ne
rect 4523 -1648 4532 -1642
tri 4532 -1648 4538 -1642 sw
rect 4396 -1674 4441 -1664
rect 4272 -1702 4346 -1678
rect 4214 -1706 4346 -1702
tri 4346 -1706 4374 -1678 sw
rect 4396 -1688 4398 -1674
tri 4396 -1690 4398 -1688 ne
rect 4410 -1692 4441 -1674
rect 4410 -1702 4456 -1692
rect 4523 -1663 4538 -1648
tri 4148 -1727 4160 -1715 ne
rect 4160 -1720 4170 -1715
tri 4170 -1720 4175 -1715 sw
rect 4059 -2066 4074 -1838
rect 4160 -1876 4175 -1720
rect 4214 -1762 4242 -1706
tri 4334 -1724 4352 -1706 ne
rect 4352 -1726 4374 -1706
tri 4374 -1726 4394 -1706 sw
tri 4410 -1720 4428 -1702 ne
rect 4233 -1796 4242 -1762
rect 4276 -1735 4318 -1734
rect 4276 -1769 4281 -1735
rect 4311 -1769 4318 -1735
rect 4276 -1778 4318 -1769
rect 4352 -1735 4394 -1726
rect 4352 -1769 4359 -1735
rect 4389 -1769 4394 -1735
rect 4352 -1774 4394 -1769
rect 4428 -1762 4456 -1702
tri 4501 -1715 4523 -1693 se
rect 4523 -1700 4538 -1692
tri 4523 -1715 4538 -1700 nw
tri 4495 -1721 4501 -1715 se
rect 4501 -1721 4510 -1715
rect 4214 -1806 4242 -1796
tri 4242 -1806 4266 -1782 sw
rect 4214 -1838 4256 -1806
tri 4273 -1814 4274 -1813 sw
rect 4273 -1838 4274 -1814
tri 4276 -1815 4313 -1778 ne
rect 4313 -1806 4318 -1778
tri 4318 -1806 4344 -1780 sw
rect 4428 -1796 4437 -1762
rect 4428 -1806 4456 -1796
rect 4313 -1815 4397 -1806
tri 4313 -1834 4332 -1815 ne
rect 4332 -1834 4397 -1815
rect 4214 -1860 4274 -1838
rect 4396 -1838 4397 -1834
rect 4414 -1838 4456 -1806
rect 4396 -1860 4456 -1838
rect 4302 -1876 4319 -1862
rect 4351 -1876 4368 -1862
tri 4139 -1912 4161 -1890 se
rect 4161 -1897 4176 -1876
tri 4161 -1912 4176 -1897 nw
rect 4495 -1897 4510 -1721
tri 4510 -1728 4523 -1715 nw
rect 4596 -1796 4611 -1568
tri 4133 -1918 4139 -1912 se
rect 4139 -1918 4148 -1912
rect 4133 -1934 4148 -1918
tri 4148 -1925 4161 -1912 nw
rect 4302 -1920 4319 -1906
rect 4351 -1920 4368 -1906
tri 4495 -1912 4510 -1897 ne
tri 4510 -1912 4532 -1890 sw
rect 4133 -1970 4148 -1962
rect 4214 -1934 4274 -1920
rect 4229 -1944 4274 -1934
rect 4229 -1962 4257 -1944
tri 4133 -1985 4148 -1970 ne
tri 4148 -1985 4170 -1963 sw
rect 4214 -1972 4257 -1962
rect 4272 -1948 4274 -1944
rect 4396 -1934 4456 -1920
tri 4510 -1925 4523 -1912 ne
rect 4523 -1918 4532 -1912
tri 4532 -1918 4538 -1912 sw
rect 4396 -1944 4441 -1934
rect 4272 -1972 4346 -1948
rect 4214 -1976 4346 -1972
tri 4346 -1976 4374 -1948 sw
rect 4396 -1958 4398 -1944
tri 4396 -1960 4398 -1958 ne
rect 4410 -1962 4441 -1944
rect 4410 -1972 4456 -1962
rect 4523 -1933 4538 -1918
tri 4148 -1997 4160 -1985 ne
rect 4160 -1990 4170 -1985
tri 4170 -1990 4175 -1985 sw
rect 4059 -2146 4074 -2108
rect 4160 -2146 4175 -1990
rect 4214 -2032 4242 -1976
tri 4334 -1994 4352 -1976 ne
rect 4352 -1996 4374 -1976
tri 4374 -1996 4394 -1976 sw
tri 4410 -1990 4428 -1972 ne
rect 4233 -2066 4242 -2032
rect 4276 -2005 4318 -2004
rect 4276 -2039 4281 -2005
rect 4311 -2039 4318 -2005
rect 4276 -2048 4318 -2039
rect 4352 -2005 4394 -1996
rect 4352 -2039 4359 -2005
rect 4389 -2039 4394 -2005
rect 4352 -2044 4394 -2039
rect 4428 -2032 4456 -1972
tri 4501 -1985 4523 -1963 se
rect 4523 -1970 4538 -1962
tri 4523 -1985 4538 -1970 nw
tri 4495 -1991 4501 -1985 se
rect 4501 -1991 4510 -1985
rect 4214 -2076 4242 -2066
tri 4242 -2076 4266 -2052 sw
rect 4214 -2108 4256 -2076
tri 4273 -2084 4274 -2083 sw
rect 4273 -2108 4274 -2084
tri 4276 -2085 4313 -2048 ne
rect 4313 -2076 4318 -2048
tri 4318 -2076 4344 -2050 sw
rect 4428 -2066 4437 -2032
rect 4428 -2076 4456 -2066
rect 4313 -2085 4397 -2076
tri 4313 -2104 4332 -2085 ne
rect 4332 -2104 4397 -2085
rect 4214 -2130 4274 -2108
rect 4396 -2108 4397 -2104
rect 4414 -2108 4456 -2076
rect 4396 -2130 4456 -2108
rect 4302 -2146 4319 -2132
rect 4351 -2146 4368 -2132
rect 4495 -2146 4510 -1991
tri 4510 -1998 4523 -1985 nw
rect 4596 -2066 4611 -1838
rect 4596 -2146 4611 -2108
rect 4639 1984 4654 2174
tri 4719 2138 4741 2160 se
rect 4741 2153 4756 2174
tri 4741 2138 4756 2153 nw
rect 5075 2153 5090 2174
tri 4713 2132 4719 2138 se
rect 4719 2132 4728 2138
rect 4713 2116 4728 2132
tri 4728 2125 4741 2138 nw
rect 4882 2130 4899 2144
rect 4931 2130 4948 2144
tri 5075 2138 5090 2153 ne
tri 5090 2138 5112 2160 sw
rect 4713 2080 4728 2088
rect 4794 2116 4854 2130
rect 4809 2106 4854 2116
rect 4809 2088 4837 2106
tri 4713 2065 4728 2080 ne
tri 4728 2065 4750 2087 sw
rect 4794 2078 4837 2088
rect 4852 2102 4854 2106
rect 4976 2116 5036 2130
tri 5090 2125 5103 2138 ne
rect 5103 2132 5112 2138
tri 5112 2132 5118 2138 sw
rect 4976 2106 5021 2116
rect 4852 2078 4926 2102
rect 4794 2074 4926 2078
tri 4926 2074 4954 2102 sw
rect 4976 2092 4978 2106
tri 4976 2090 4978 2092 ne
rect 4990 2088 5021 2106
rect 4990 2078 5036 2088
rect 5103 2117 5118 2132
tri 4728 2053 4740 2065 ne
rect 4740 2060 4750 2065
tri 4750 2060 4755 2065 sw
rect 4639 1714 4654 1942
rect 4740 1904 4755 2060
rect 4794 2018 4822 2074
tri 4914 2056 4932 2074 ne
rect 4932 2054 4954 2074
tri 4954 2054 4974 2074 sw
tri 4990 2060 5008 2078 ne
rect 4813 1984 4822 2018
rect 4856 2045 4898 2046
rect 4856 2011 4861 2045
rect 4891 2011 4898 2045
rect 4856 2002 4898 2011
rect 4932 2045 4974 2054
rect 4932 2011 4939 2045
rect 4969 2011 4974 2045
rect 4932 2006 4974 2011
rect 5008 2018 5036 2078
tri 5081 2065 5103 2087 se
rect 5103 2080 5118 2088
tri 5103 2065 5118 2080 nw
tri 5075 2059 5081 2065 se
rect 5081 2059 5090 2065
rect 4794 1974 4822 1984
tri 4822 1974 4846 1998 sw
rect 4794 1942 4836 1974
tri 4853 1966 4854 1967 sw
rect 4853 1942 4854 1966
tri 4856 1965 4893 2002 ne
rect 4893 1974 4898 2002
tri 4898 1974 4924 2000 sw
rect 5008 1984 5017 2018
rect 5008 1974 5036 1984
rect 4893 1965 4977 1974
tri 4893 1946 4912 1965 ne
rect 4912 1946 4977 1965
rect 4794 1920 4854 1942
rect 4976 1942 4977 1946
rect 4994 1942 5036 1974
rect 4976 1920 5036 1942
rect 4882 1904 4899 1918
rect 4931 1904 4948 1918
tri 4719 1868 4741 1890 se
rect 4741 1883 4756 1904
tri 4741 1868 4756 1883 nw
rect 5075 1883 5090 2059
tri 5090 2052 5103 2065 nw
rect 5176 1984 5191 2174
tri 4713 1862 4719 1868 se
rect 4719 1862 4728 1868
rect 4713 1846 4728 1862
tri 4728 1855 4741 1868 nw
rect 4882 1860 4899 1874
rect 4931 1860 4948 1874
tri 5075 1868 5090 1883 ne
tri 5090 1868 5112 1890 sw
rect 4713 1810 4728 1818
rect 4794 1846 4854 1860
rect 4809 1836 4854 1846
rect 4809 1818 4837 1836
tri 4713 1795 4728 1810 ne
tri 4728 1795 4750 1817 sw
rect 4794 1808 4837 1818
rect 4852 1832 4854 1836
rect 4976 1846 5036 1860
tri 5090 1855 5103 1868 ne
rect 5103 1862 5112 1868
tri 5112 1862 5118 1868 sw
rect 4976 1836 5021 1846
rect 4852 1808 4926 1832
rect 4794 1804 4926 1808
tri 4926 1804 4954 1832 sw
rect 4976 1822 4978 1836
tri 4976 1820 4978 1822 ne
rect 4990 1818 5021 1836
rect 4990 1808 5036 1818
rect 5103 1847 5118 1862
tri 4728 1783 4740 1795 ne
rect 4740 1790 4750 1795
tri 4750 1790 4755 1795 sw
rect 4639 1444 4654 1672
rect 4740 1682 4755 1790
rect 4794 1748 4822 1804
tri 4914 1786 4932 1804 ne
rect 4932 1784 4954 1804
tri 4954 1784 4974 1804 sw
tri 4990 1790 5008 1808 ne
rect 4813 1714 4822 1748
rect 4856 1775 4898 1776
rect 4856 1741 4861 1775
rect 4891 1741 4898 1775
rect 4856 1732 4898 1741
rect 4932 1775 4974 1784
rect 4932 1741 4939 1775
rect 4969 1741 4974 1775
rect 4932 1736 4974 1741
rect 5008 1748 5036 1808
tri 5081 1795 5103 1817 se
rect 5103 1810 5118 1818
tri 5103 1795 5118 1810 nw
tri 5075 1789 5081 1795 se
rect 5081 1789 5090 1795
rect 4794 1704 4822 1714
tri 4822 1704 4846 1728 sw
rect 4740 1634 4756 1682
rect 4794 1672 4836 1704
tri 4853 1696 4854 1697 sw
rect 4853 1672 4854 1696
tri 4856 1695 4893 1732 ne
rect 4893 1704 4898 1732
tri 4898 1704 4924 1730 sw
rect 5008 1714 5017 1748
rect 5008 1704 5036 1714
rect 4893 1695 4977 1704
tri 4893 1676 4912 1695 ne
rect 4912 1676 4977 1695
rect 4794 1650 4854 1672
rect 4976 1672 4977 1676
rect 4994 1672 5036 1704
rect 4976 1650 5036 1672
rect 4882 1634 4899 1648
rect 4931 1634 4948 1648
tri 4719 1598 4741 1620 se
rect 4741 1613 4756 1634
tri 4741 1598 4756 1613 nw
rect 5075 1613 5090 1789
tri 5090 1782 5103 1795 nw
rect 5176 1714 5191 1942
tri 4713 1592 4719 1598 se
rect 4719 1592 4728 1598
rect 4713 1576 4728 1592
tri 4728 1585 4741 1598 nw
rect 4882 1590 4899 1604
rect 4931 1590 4948 1604
tri 5075 1598 5090 1613 ne
tri 5090 1598 5112 1620 sw
rect 4713 1540 4728 1548
rect 4794 1576 4854 1590
rect 4809 1566 4854 1576
rect 4809 1548 4837 1566
tri 4713 1525 4728 1540 ne
tri 4728 1525 4750 1547 sw
rect 4794 1538 4837 1548
rect 4852 1562 4854 1566
rect 4976 1576 5036 1590
tri 5090 1585 5103 1598 ne
rect 5103 1592 5112 1598
tri 5112 1592 5118 1598 sw
rect 4976 1566 5021 1576
rect 4852 1538 4926 1562
rect 4794 1534 4926 1538
tri 4926 1534 4954 1562 sw
rect 4976 1552 4978 1566
tri 4976 1550 4978 1552 ne
rect 4990 1548 5021 1566
rect 4990 1538 5036 1548
rect 5103 1577 5118 1592
tri 4728 1513 4740 1525 ne
rect 4740 1520 4750 1525
tri 4750 1520 4755 1525 sw
rect 4639 1174 4654 1402
rect 4740 1364 4755 1520
rect 4794 1478 4822 1534
tri 4914 1516 4932 1534 ne
rect 4932 1514 4954 1534
tri 4954 1514 4974 1534 sw
tri 4990 1520 5008 1538 ne
rect 4813 1444 4822 1478
rect 4856 1505 4898 1506
rect 4856 1471 4861 1505
rect 4891 1471 4898 1505
rect 4856 1462 4898 1471
rect 4932 1505 4974 1514
rect 4932 1471 4939 1505
rect 4969 1471 4974 1505
rect 4932 1466 4974 1471
rect 5008 1478 5036 1538
tri 5081 1525 5103 1547 se
rect 5103 1540 5118 1548
tri 5103 1525 5118 1540 nw
tri 5075 1519 5081 1525 se
rect 5081 1519 5090 1525
rect 4794 1434 4822 1444
tri 4822 1434 4846 1458 sw
rect 4794 1402 4836 1434
tri 4853 1426 4854 1427 sw
rect 4853 1402 4854 1426
tri 4856 1425 4893 1462 ne
rect 4893 1434 4898 1462
tri 4898 1434 4924 1460 sw
rect 5008 1444 5017 1478
rect 5008 1434 5036 1444
rect 4893 1425 4977 1434
tri 4893 1406 4912 1425 ne
rect 4912 1406 4977 1425
rect 4794 1380 4854 1402
rect 4976 1402 4977 1406
rect 4994 1402 5036 1434
rect 4976 1380 5036 1402
rect 4882 1364 4899 1378
rect 4931 1364 4948 1378
tri 4719 1328 4741 1350 se
rect 4741 1343 4756 1364
tri 4741 1328 4756 1343 nw
rect 5075 1343 5090 1519
tri 5090 1512 5103 1525 nw
rect 5176 1444 5191 1672
tri 4713 1322 4719 1328 se
rect 4719 1322 4728 1328
rect 4713 1306 4728 1322
tri 4728 1315 4741 1328 nw
rect 4882 1320 4899 1334
rect 4931 1320 4948 1334
tri 5075 1328 5090 1343 ne
tri 5090 1328 5112 1350 sw
rect 4713 1270 4728 1278
rect 4794 1306 4854 1320
rect 4809 1296 4854 1306
rect 4809 1278 4837 1296
tri 4713 1255 4728 1270 ne
tri 4728 1255 4750 1277 sw
rect 4794 1268 4837 1278
rect 4852 1292 4854 1296
rect 4976 1306 5036 1320
tri 5090 1315 5103 1328 ne
rect 5103 1322 5112 1328
tri 5112 1322 5118 1328 sw
rect 4976 1296 5021 1306
rect 4852 1268 4926 1292
rect 4794 1264 4926 1268
tri 4926 1264 4954 1292 sw
rect 4976 1282 4978 1296
tri 4976 1280 4978 1282 ne
rect 4990 1278 5021 1296
rect 4990 1268 5036 1278
rect 5103 1307 5118 1322
tri 4728 1243 4740 1255 ne
rect 4740 1250 4750 1255
tri 4750 1250 4755 1255 sw
rect 4639 904 4654 1132
rect 4740 1142 4755 1250
rect 4794 1208 4822 1264
tri 4914 1246 4932 1264 ne
rect 4932 1244 4954 1264
tri 4954 1244 4974 1264 sw
tri 4990 1250 5008 1268 ne
rect 4813 1174 4822 1208
rect 4856 1235 4898 1236
rect 4856 1201 4861 1235
rect 4891 1201 4898 1235
rect 4856 1192 4898 1201
rect 4932 1235 4974 1244
rect 4932 1201 4939 1235
rect 4969 1201 4974 1235
rect 4932 1196 4974 1201
rect 5008 1208 5036 1268
tri 5081 1255 5103 1277 se
rect 5103 1270 5118 1278
tri 5103 1255 5118 1270 nw
tri 5075 1249 5081 1255 se
rect 5081 1249 5090 1255
rect 4794 1164 4822 1174
tri 4822 1164 4846 1188 sw
rect 4740 1094 4756 1142
rect 4794 1132 4836 1164
tri 4853 1156 4854 1157 sw
rect 4853 1132 4854 1156
tri 4856 1155 4893 1192 ne
rect 4893 1164 4898 1192
tri 4898 1164 4924 1190 sw
rect 5008 1174 5017 1208
rect 5008 1164 5036 1174
rect 4893 1155 4977 1164
tri 4893 1136 4912 1155 ne
rect 4912 1136 4977 1155
rect 4794 1110 4854 1132
rect 4976 1132 4977 1136
rect 4994 1132 5036 1164
rect 4976 1110 5036 1132
rect 4882 1094 4899 1108
rect 4931 1094 4948 1108
tri 4719 1058 4741 1080 se
rect 4741 1073 4756 1094
tri 4741 1058 4756 1073 nw
rect 5075 1073 5090 1249
tri 5090 1242 5103 1255 nw
rect 5176 1174 5191 1402
tri 4713 1052 4719 1058 se
rect 4719 1052 4728 1058
rect 4713 1036 4728 1052
tri 4728 1045 4741 1058 nw
rect 4882 1050 4899 1064
rect 4931 1050 4948 1064
tri 5075 1058 5090 1073 ne
tri 5090 1058 5112 1080 sw
rect 4713 1000 4728 1008
rect 4794 1036 4854 1050
rect 4809 1026 4854 1036
rect 4809 1008 4837 1026
tri 4713 985 4728 1000 ne
tri 4728 985 4750 1007 sw
rect 4794 998 4837 1008
rect 4852 1022 4854 1026
rect 4976 1036 5036 1050
tri 5090 1045 5103 1058 ne
rect 5103 1052 5112 1058
tri 5112 1052 5118 1058 sw
rect 4976 1026 5021 1036
rect 4852 998 4926 1022
rect 4794 994 4926 998
tri 4926 994 4954 1022 sw
rect 4976 1012 4978 1026
tri 4976 1010 4978 1012 ne
rect 4990 1008 5021 1026
rect 4990 998 5036 1008
rect 5103 1037 5118 1052
tri 4728 973 4740 985 ne
rect 4740 980 4750 985
tri 4750 980 4755 985 sw
rect 4639 634 4654 862
rect 4740 824 4755 980
rect 4794 938 4822 994
tri 4914 976 4932 994 ne
rect 4932 974 4954 994
tri 4954 974 4974 994 sw
tri 4990 980 5008 998 ne
rect 4813 904 4822 938
rect 4856 965 4898 966
rect 4856 931 4861 965
rect 4891 931 4898 965
rect 4856 922 4898 931
rect 4932 965 4974 974
rect 4932 931 4939 965
rect 4969 931 4974 965
rect 4932 926 4974 931
rect 5008 938 5036 998
tri 5081 985 5103 1007 se
rect 5103 1000 5118 1008
tri 5103 985 5118 1000 nw
tri 5075 979 5081 985 se
rect 5081 979 5090 985
rect 4794 894 4822 904
tri 4822 894 4846 918 sw
rect 4794 862 4836 894
tri 4853 886 4854 887 sw
rect 4853 862 4854 886
tri 4856 885 4893 922 ne
rect 4893 894 4898 922
tri 4898 894 4924 920 sw
rect 5008 904 5017 938
rect 5008 894 5036 904
rect 4893 885 4977 894
tri 4893 866 4912 885 ne
rect 4912 866 4977 885
rect 4794 840 4854 862
rect 4976 862 4977 866
rect 4994 862 5036 894
rect 4976 840 5036 862
rect 4882 824 4899 838
rect 4931 824 4948 838
tri 4719 788 4741 810 se
rect 4741 803 4756 824
tri 4741 788 4756 803 nw
rect 5075 803 5090 979
tri 5090 972 5103 985 nw
rect 5176 904 5191 1132
tri 4713 782 4719 788 se
rect 4719 782 4728 788
rect 4713 766 4728 782
tri 4728 775 4741 788 nw
rect 4882 780 4899 794
rect 4931 780 4948 794
tri 5075 788 5090 803 ne
tri 5090 788 5112 810 sw
rect 4713 730 4728 738
rect 4794 766 4854 780
rect 4809 756 4854 766
rect 4809 738 4837 756
tri 4713 715 4728 730 ne
tri 4728 715 4750 737 sw
rect 4794 728 4837 738
rect 4852 752 4854 756
rect 4976 766 5036 780
tri 5090 775 5103 788 ne
rect 5103 782 5112 788
tri 5112 782 5118 788 sw
rect 4976 756 5021 766
rect 4852 728 4926 752
rect 4794 724 4926 728
tri 4926 724 4954 752 sw
rect 4976 742 4978 756
tri 4976 740 4978 742 ne
rect 4990 738 5021 756
rect 4990 728 5036 738
rect 5103 767 5118 782
tri 4728 703 4740 715 ne
rect 4740 710 4750 715
tri 4750 710 4755 715 sw
rect 4639 364 4654 592
rect 4740 602 4755 710
rect 4794 668 4822 724
tri 4914 706 4932 724 ne
rect 4932 704 4954 724
tri 4954 704 4974 724 sw
tri 4990 710 5008 728 ne
rect 4813 634 4822 668
rect 4856 695 4898 696
rect 4856 661 4861 695
rect 4891 661 4898 695
rect 4856 652 4898 661
rect 4932 695 4974 704
rect 4932 661 4939 695
rect 4969 661 4974 695
rect 4932 656 4974 661
rect 5008 668 5036 728
tri 5081 715 5103 737 se
rect 5103 730 5118 738
tri 5103 715 5118 730 nw
tri 5075 709 5081 715 se
rect 5081 709 5090 715
rect 4794 624 4822 634
tri 4822 624 4846 648 sw
rect 4740 554 4756 602
rect 4794 592 4836 624
tri 4853 616 4854 617 sw
rect 4853 592 4854 616
tri 4856 615 4893 652 ne
rect 4893 624 4898 652
tri 4898 624 4924 650 sw
rect 5008 634 5017 668
rect 5008 624 5036 634
rect 4893 615 4977 624
tri 4893 596 4912 615 ne
rect 4912 596 4977 615
rect 4794 570 4854 592
rect 4976 592 4977 596
rect 4994 592 5036 624
rect 4976 570 5036 592
rect 4882 554 4899 568
rect 4931 554 4948 568
tri 4719 518 4741 540 se
rect 4741 533 4756 554
tri 4741 518 4756 533 nw
rect 5075 533 5090 709
tri 5090 702 5103 715 nw
rect 5176 634 5191 862
tri 4713 512 4719 518 se
rect 4719 512 4728 518
rect 4713 496 4728 512
tri 4728 505 4741 518 nw
rect 4882 510 4899 524
rect 4931 510 4948 524
tri 5075 518 5090 533 ne
tri 5090 518 5112 540 sw
rect 4713 460 4728 468
rect 4794 496 4854 510
rect 4809 486 4854 496
rect 4809 468 4837 486
tri 4713 445 4728 460 ne
tri 4728 445 4750 467 sw
rect 4794 458 4837 468
rect 4852 482 4854 486
rect 4976 496 5036 510
tri 5090 505 5103 518 ne
rect 5103 512 5112 518
tri 5112 512 5118 518 sw
rect 4976 486 5021 496
rect 4852 458 4926 482
rect 4794 454 4926 458
tri 4926 454 4954 482 sw
rect 4976 472 4978 486
tri 4976 470 4978 472 ne
rect 4990 468 5021 486
rect 4990 458 5036 468
rect 5103 497 5118 512
tri 4728 433 4740 445 ne
rect 4740 440 4750 445
tri 4750 440 4755 445 sw
rect 4639 94 4654 322
rect 4740 284 4755 440
rect 4794 398 4822 454
tri 4914 436 4932 454 ne
rect 4932 434 4954 454
tri 4954 434 4974 454 sw
tri 4990 440 5008 458 ne
rect 4813 364 4822 398
rect 4856 425 4898 426
rect 4856 391 4861 425
rect 4891 391 4898 425
rect 4856 382 4898 391
rect 4932 425 4974 434
rect 4932 391 4939 425
rect 4969 391 4974 425
rect 4932 386 4974 391
rect 5008 398 5036 458
tri 5081 445 5103 467 se
rect 5103 460 5118 468
tri 5103 445 5118 460 nw
tri 5075 439 5081 445 se
rect 5081 439 5090 445
rect 4794 354 4822 364
tri 4822 354 4846 378 sw
rect 4794 322 4836 354
tri 4853 346 4854 347 sw
rect 4853 322 4854 346
tri 4856 345 4893 382 ne
rect 4893 354 4898 382
tri 4898 354 4924 380 sw
rect 5008 364 5017 398
rect 5008 354 5036 364
rect 4893 345 4977 354
tri 4893 326 4912 345 ne
rect 4912 326 4977 345
rect 4794 300 4854 322
rect 4976 322 4977 326
rect 4994 322 5036 354
rect 4976 300 5036 322
rect 4882 284 4899 298
rect 4931 284 4948 298
tri 4719 248 4741 270 se
rect 4741 263 4756 284
tri 4741 248 4756 263 nw
rect 5075 263 5090 439
tri 5090 432 5103 445 nw
rect 5176 364 5191 592
tri 4713 242 4719 248 se
rect 4719 242 4728 248
rect 4713 226 4728 242
tri 4728 235 4741 248 nw
rect 4882 240 4899 254
rect 4931 240 4948 254
tri 5075 248 5090 263 ne
tri 5090 248 5112 270 sw
rect 4713 190 4728 198
rect 4794 226 4854 240
rect 4809 216 4854 226
rect 4809 198 4837 216
tri 4713 175 4728 190 ne
tri 4728 175 4750 197 sw
rect 4794 188 4837 198
rect 4852 212 4854 216
rect 4976 226 5036 240
tri 5090 235 5103 248 ne
rect 5103 242 5112 248
tri 5112 242 5118 248 sw
rect 4976 216 5021 226
rect 4852 188 4926 212
rect 4794 184 4926 188
tri 4926 184 4954 212 sw
rect 4976 202 4978 216
tri 4976 200 4978 202 ne
rect 4990 198 5021 216
rect 4990 188 5036 198
rect 5103 227 5118 242
tri 4728 163 4740 175 ne
rect 4740 170 4750 175
tri 4750 170 4755 175 sw
rect 4639 -176 4654 52
rect 4740 62 4755 170
rect 4794 128 4822 184
tri 4914 166 4932 184 ne
rect 4932 164 4954 184
tri 4954 164 4974 184 sw
tri 4990 170 5008 188 ne
rect 4813 94 4822 128
rect 4856 155 4898 156
rect 4856 121 4861 155
rect 4891 121 4898 155
rect 4856 112 4898 121
rect 4932 155 4974 164
rect 4932 121 4939 155
rect 4969 121 4974 155
rect 4932 116 4974 121
rect 5008 128 5036 188
tri 5081 175 5103 197 se
rect 5103 190 5118 198
tri 5103 175 5118 190 nw
tri 5075 169 5081 175 se
rect 5081 169 5090 175
rect 4794 84 4822 94
tri 4822 84 4846 108 sw
rect 4740 14 4756 62
rect 4794 52 4836 84
tri 4853 76 4854 77 sw
rect 4853 52 4854 76
tri 4856 75 4893 112 ne
rect 4893 84 4898 112
tri 4898 84 4924 110 sw
rect 5008 94 5017 128
rect 5008 84 5036 94
rect 4893 75 4977 84
tri 4893 56 4912 75 ne
rect 4912 56 4977 75
rect 4794 30 4854 52
rect 4976 52 4977 56
rect 4994 52 5036 84
rect 4976 30 5036 52
rect 4882 14 4899 28
rect 4931 14 4948 28
tri 4719 -22 4741 0 se
rect 4741 -7 4756 14
tri 4741 -22 4756 -7 nw
rect 5075 -7 5090 169
tri 5090 162 5103 175 nw
rect 5176 94 5191 322
tri 4713 -28 4719 -22 se
rect 4719 -28 4728 -22
rect 4713 -44 4728 -28
tri 4728 -35 4741 -22 nw
rect 4882 -30 4899 -16
rect 4931 -30 4948 -16
tri 5075 -22 5090 -7 ne
tri 5090 -22 5112 0 sw
rect 4713 -80 4728 -72
rect 4794 -44 4854 -30
rect 4809 -54 4854 -44
rect 4809 -72 4837 -54
tri 4713 -95 4728 -80 ne
tri 4728 -95 4750 -73 sw
rect 4794 -82 4837 -72
rect 4852 -58 4854 -54
rect 4976 -44 5036 -30
tri 5090 -35 5103 -22 ne
rect 5103 -28 5112 -22
tri 5112 -28 5118 -22 sw
rect 4976 -54 5021 -44
rect 4852 -82 4926 -58
rect 4794 -86 4926 -82
tri 4926 -86 4954 -58 sw
rect 4976 -68 4978 -54
tri 4976 -70 4978 -68 ne
rect 4990 -72 5021 -54
rect 4990 -82 5036 -72
rect 5103 -43 5118 -28
tri 4728 -107 4740 -95 ne
rect 4740 -100 4750 -95
tri 4750 -100 4755 -95 sw
rect 4639 -446 4654 -218
rect 4740 -256 4755 -100
rect 4794 -142 4822 -86
tri 4914 -104 4932 -86 ne
rect 4932 -106 4954 -86
tri 4954 -106 4974 -86 sw
tri 4990 -100 5008 -82 ne
rect 4813 -176 4822 -142
rect 4856 -115 4898 -114
rect 4856 -149 4861 -115
rect 4891 -149 4898 -115
rect 4856 -158 4898 -149
rect 4932 -115 4974 -106
rect 4932 -149 4939 -115
rect 4969 -149 4974 -115
rect 4932 -154 4974 -149
rect 5008 -142 5036 -82
tri 5081 -95 5103 -73 se
rect 5103 -80 5118 -72
tri 5103 -95 5118 -80 nw
tri 5075 -101 5081 -95 se
rect 5081 -101 5090 -95
rect 4794 -186 4822 -176
tri 4822 -186 4846 -162 sw
rect 4794 -218 4836 -186
tri 4853 -194 4854 -193 sw
rect 4853 -218 4854 -194
tri 4856 -195 4893 -158 ne
rect 4893 -186 4898 -158
tri 4898 -186 4924 -160 sw
rect 5008 -176 5017 -142
rect 5008 -186 5036 -176
rect 4893 -195 4977 -186
tri 4893 -214 4912 -195 ne
rect 4912 -214 4977 -195
rect 4794 -240 4854 -218
rect 4976 -218 4977 -214
rect 4994 -218 5036 -186
rect 4976 -240 5036 -218
rect 4882 -256 4899 -242
rect 4931 -256 4948 -242
tri 4719 -292 4741 -270 se
rect 4741 -277 4756 -256
tri 4741 -292 4756 -277 nw
rect 5075 -277 5090 -101
tri 5090 -108 5103 -95 nw
rect 5176 -176 5191 52
tri 4713 -298 4719 -292 se
rect 4719 -298 4728 -292
rect 4713 -314 4728 -298
tri 4728 -305 4741 -292 nw
rect 4882 -300 4899 -286
rect 4931 -300 4948 -286
tri 5075 -292 5090 -277 ne
tri 5090 -292 5112 -270 sw
rect 4713 -350 4728 -342
rect 4794 -314 4854 -300
rect 4809 -324 4854 -314
rect 4809 -342 4837 -324
tri 4713 -365 4728 -350 ne
tri 4728 -365 4750 -343 sw
rect 4794 -352 4837 -342
rect 4852 -328 4854 -324
rect 4976 -314 5036 -300
tri 5090 -305 5103 -292 ne
rect 5103 -298 5112 -292
tri 5112 -298 5118 -292 sw
rect 4976 -324 5021 -314
rect 4852 -352 4926 -328
rect 4794 -356 4926 -352
tri 4926 -356 4954 -328 sw
rect 4976 -338 4978 -324
tri 4976 -340 4978 -338 ne
rect 4990 -342 5021 -324
rect 4990 -352 5036 -342
rect 5103 -313 5118 -298
tri 4728 -377 4740 -365 ne
rect 4740 -370 4750 -365
tri 4750 -370 4755 -365 sw
rect 4639 -716 4654 -488
rect 4740 -478 4755 -370
rect 4794 -412 4822 -356
tri 4914 -374 4932 -356 ne
rect 4932 -376 4954 -356
tri 4954 -376 4974 -356 sw
tri 4990 -370 5008 -352 ne
rect 4813 -446 4822 -412
rect 4856 -385 4898 -384
rect 4856 -419 4861 -385
rect 4891 -419 4898 -385
rect 4856 -428 4898 -419
rect 4932 -385 4974 -376
rect 4932 -419 4939 -385
rect 4969 -419 4974 -385
rect 4932 -424 4974 -419
rect 5008 -412 5036 -352
tri 5081 -365 5103 -343 se
rect 5103 -350 5118 -342
tri 5103 -365 5118 -350 nw
tri 5075 -371 5081 -365 se
rect 5081 -371 5090 -365
rect 4794 -456 4822 -446
tri 4822 -456 4846 -432 sw
rect 4740 -526 4756 -478
rect 4794 -488 4836 -456
tri 4853 -464 4854 -463 sw
rect 4853 -488 4854 -464
tri 4856 -465 4893 -428 ne
rect 4893 -456 4898 -428
tri 4898 -456 4924 -430 sw
rect 5008 -446 5017 -412
rect 5008 -456 5036 -446
rect 4893 -465 4977 -456
tri 4893 -484 4912 -465 ne
rect 4912 -484 4977 -465
rect 4794 -510 4854 -488
rect 4976 -488 4977 -484
rect 4994 -488 5036 -456
rect 4976 -510 5036 -488
rect 4882 -526 4899 -512
rect 4931 -526 4948 -512
tri 4719 -562 4741 -540 se
rect 4741 -547 4756 -526
tri 4741 -562 4756 -547 nw
rect 5075 -547 5090 -371
tri 5090 -378 5103 -365 nw
rect 5176 -446 5191 -218
tri 4713 -568 4719 -562 se
rect 4719 -568 4728 -562
rect 4713 -584 4728 -568
tri 4728 -575 4741 -562 nw
rect 4882 -570 4899 -556
rect 4931 -570 4948 -556
tri 5075 -562 5090 -547 ne
tri 5090 -562 5112 -540 sw
rect 4713 -620 4728 -612
rect 4794 -584 4854 -570
rect 4809 -594 4854 -584
rect 4809 -612 4837 -594
tri 4713 -635 4728 -620 ne
tri 4728 -635 4750 -613 sw
rect 4794 -622 4837 -612
rect 4852 -598 4854 -594
rect 4976 -584 5036 -570
tri 5090 -575 5103 -562 ne
rect 5103 -568 5112 -562
tri 5112 -568 5118 -562 sw
rect 4976 -594 5021 -584
rect 4852 -622 4926 -598
rect 4794 -626 4926 -622
tri 4926 -626 4954 -598 sw
rect 4976 -608 4978 -594
tri 4976 -610 4978 -608 ne
rect 4990 -612 5021 -594
rect 4990 -622 5036 -612
rect 5103 -583 5118 -568
tri 4728 -647 4740 -635 ne
rect 4740 -640 4750 -635
tri 4750 -640 4755 -635 sw
rect 4639 -986 4654 -758
rect 4740 -796 4755 -640
rect 4794 -682 4822 -626
tri 4914 -644 4932 -626 ne
rect 4932 -646 4954 -626
tri 4954 -646 4974 -626 sw
tri 4990 -640 5008 -622 ne
rect 4813 -716 4822 -682
rect 4856 -655 4898 -654
rect 4856 -689 4861 -655
rect 4891 -689 4898 -655
rect 4856 -698 4898 -689
rect 4932 -655 4974 -646
rect 4932 -689 4939 -655
rect 4969 -689 4974 -655
rect 4932 -694 4974 -689
rect 5008 -682 5036 -622
tri 5081 -635 5103 -613 se
rect 5103 -620 5118 -612
tri 5103 -635 5118 -620 nw
tri 5075 -641 5081 -635 se
rect 5081 -641 5090 -635
rect 4794 -726 4822 -716
tri 4822 -726 4846 -702 sw
rect 4794 -758 4836 -726
tri 4853 -734 4854 -733 sw
rect 4853 -758 4854 -734
tri 4856 -735 4893 -698 ne
rect 4893 -726 4898 -698
tri 4898 -726 4924 -700 sw
rect 5008 -716 5017 -682
rect 5008 -726 5036 -716
rect 4893 -735 4977 -726
tri 4893 -754 4912 -735 ne
rect 4912 -754 4977 -735
rect 4794 -780 4854 -758
rect 4976 -758 4977 -754
rect 4994 -758 5036 -726
rect 4976 -780 5036 -758
rect 4882 -796 4899 -782
rect 4931 -796 4948 -782
tri 4719 -832 4741 -810 se
rect 4741 -817 4756 -796
tri 4741 -832 4756 -817 nw
rect 5075 -817 5090 -641
tri 5090 -648 5103 -635 nw
rect 5176 -716 5191 -488
tri 4713 -838 4719 -832 se
rect 4719 -838 4728 -832
rect 4713 -854 4728 -838
tri 4728 -845 4741 -832 nw
rect 4882 -840 4899 -826
rect 4931 -840 4948 -826
tri 5075 -832 5090 -817 ne
tri 5090 -832 5112 -810 sw
rect 4713 -890 4728 -882
rect 4794 -854 4854 -840
rect 4809 -864 4854 -854
rect 4809 -882 4837 -864
tri 4713 -905 4728 -890 ne
tri 4728 -905 4750 -883 sw
rect 4794 -892 4837 -882
rect 4852 -868 4854 -864
rect 4976 -854 5036 -840
tri 5090 -845 5103 -832 ne
rect 5103 -838 5112 -832
tri 5112 -838 5118 -832 sw
rect 4976 -864 5021 -854
rect 4852 -892 4926 -868
rect 4794 -896 4926 -892
tri 4926 -896 4954 -868 sw
rect 4976 -878 4978 -864
tri 4976 -880 4978 -878 ne
rect 4990 -882 5021 -864
rect 4990 -892 5036 -882
rect 5103 -853 5118 -838
tri 4728 -917 4740 -905 ne
rect 4740 -910 4750 -905
tri 4750 -910 4755 -905 sw
rect 4639 -1256 4654 -1028
rect 4740 -1018 4755 -910
rect 4794 -952 4822 -896
tri 4914 -914 4932 -896 ne
rect 4932 -916 4954 -896
tri 4954 -916 4974 -896 sw
tri 4990 -910 5008 -892 ne
rect 4813 -986 4822 -952
rect 4856 -925 4898 -924
rect 4856 -959 4861 -925
rect 4891 -959 4898 -925
rect 4856 -968 4898 -959
rect 4932 -925 4974 -916
rect 4932 -959 4939 -925
rect 4969 -959 4974 -925
rect 4932 -964 4974 -959
rect 5008 -952 5036 -892
tri 5081 -905 5103 -883 se
rect 5103 -890 5118 -882
tri 5103 -905 5118 -890 nw
tri 5075 -911 5081 -905 se
rect 5081 -911 5090 -905
rect 4794 -996 4822 -986
tri 4822 -996 4846 -972 sw
rect 4740 -1066 4756 -1018
rect 4794 -1028 4836 -996
tri 4853 -1004 4854 -1003 sw
rect 4853 -1028 4854 -1004
tri 4856 -1005 4893 -968 ne
rect 4893 -996 4898 -968
tri 4898 -996 4924 -970 sw
rect 5008 -986 5017 -952
rect 5008 -996 5036 -986
rect 4893 -1005 4977 -996
tri 4893 -1024 4912 -1005 ne
rect 4912 -1024 4977 -1005
rect 4794 -1050 4854 -1028
rect 4976 -1028 4977 -1024
rect 4994 -1028 5036 -996
rect 4976 -1050 5036 -1028
rect 4882 -1066 4899 -1052
rect 4931 -1066 4948 -1052
tri 4719 -1102 4741 -1080 se
rect 4741 -1087 4756 -1066
tri 4741 -1102 4756 -1087 nw
rect 5075 -1087 5090 -911
tri 5090 -918 5103 -905 nw
rect 5176 -986 5191 -758
tri 4713 -1108 4719 -1102 se
rect 4719 -1108 4728 -1102
rect 4713 -1124 4728 -1108
tri 4728 -1115 4741 -1102 nw
rect 4882 -1110 4899 -1096
rect 4931 -1110 4948 -1096
tri 5075 -1102 5090 -1087 ne
tri 5090 -1102 5112 -1080 sw
rect 4713 -1160 4728 -1152
rect 4794 -1124 4854 -1110
rect 4809 -1134 4854 -1124
rect 4809 -1152 4837 -1134
tri 4713 -1175 4728 -1160 ne
tri 4728 -1175 4750 -1153 sw
rect 4794 -1162 4837 -1152
rect 4852 -1138 4854 -1134
rect 4976 -1124 5036 -1110
tri 5090 -1115 5103 -1102 ne
rect 5103 -1108 5112 -1102
tri 5112 -1108 5118 -1102 sw
rect 4976 -1134 5021 -1124
rect 4852 -1162 4926 -1138
rect 4794 -1166 4926 -1162
tri 4926 -1166 4954 -1138 sw
rect 4976 -1148 4978 -1134
tri 4976 -1150 4978 -1148 ne
rect 4990 -1152 5021 -1134
rect 4990 -1162 5036 -1152
rect 5103 -1123 5118 -1108
tri 4728 -1187 4740 -1175 ne
rect 4740 -1180 4750 -1175
tri 4750 -1180 4755 -1175 sw
rect 4639 -1526 4654 -1298
rect 4740 -1336 4755 -1180
rect 4794 -1222 4822 -1166
tri 4914 -1184 4932 -1166 ne
rect 4932 -1186 4954 -1166
tri 4954 -1186 4974 -1166 sw
tri 4990 -1180 5008 -1162 ne
rect 4813 -1256 4822 -1222
rect 4856 -1195 4898 -1194
rect 4856 -1229 4861 -1195
rect 4891 -1229 4898 -1195
rect 4856 -1238 4898 -1229
rect 4932 -1195 4974 -1186
rect 4932 -1229 4939 -1195
rect 4969 -1229 4974 -1195
rect 4932 -1234 4974 -1229
rect 5008 -1222 5036 -1162
tri 5081 -1175 5103 -1153 se
rect 5103 -1160 5118 -1152
tri 5103 -1175 5118 -1160 nw
tri 5075 -1181 5081 -1175 se
rect 5081 -1181 5090 -1175
rect 4794 -1266 4822 -1256
tri 4822 -1266 4846 -1242 sw
rect 4794 -1298 4836 -1266
tri 4853 -1274 4854 -1273 sw
rect 4853 -1298 4854 -1274
tri 4856 -1275 4893 -1238 ne
rect 4893 -1266 4898 -1238
tri 4898 -1266 4924 -1240 sw
rect 5008 -1256 5017 -1222
rect 5008 -1266 5036 -1256
rect 4893 -1275 4977 -1266
tri 4893 -1294 4912 -1275 ne
rect 4912 -1294 4977 -1275
rect 4794 -1320 4854 -1298
rect 4976 -1298 4977 -1294
rect 4994 -1298 5036 -1266
rect 4976 -1320 5036 -1298
rect 4882 -1336 4899 -1322
rect 4931 -1336 4948 -1322
tri 4719 -1372 4741 -1350 se
rect 4741 -1357 4756 -1336
tri 4741 -1372 4756 -1357 nw
rect 5075 -1357 5090 -1181
tri 5090 -1188 5103 -1175 nw
rect 5176 -1256 5191 -1028
tri 4713 -1378 4719 -1372 se
rect 4719 -1378 4728 -1372
rect 4713 -1394 4728 -1378
tri 4728 -1385 4741 -1372 nw
rect 4882 -1380 4899 -1366
rect 4931 -1380 4948 -1366
tri 5075 -1372 5090 -1357 ne
tri 5090 -1372 5112 -1350 sw
rect 4713 -1430 4728 -1422
rect 4794 -1394 4854 -1380
rect 4809 -1404 4854 -1394
rect 4809 -1422 4837 -1404
tri 4713 -1445 4728 -1430 ne
tri 4728 -1445 4750 -1423 sw
rect 4794 -1432 4837 -1422
rect 4852 -1408 4854 -1404
rect 4976 -1394 5036 -1380
tri 5090 -1385 5103 -1372 ne
rect 5103 -1378 5112 -1372
tri 5112 -1378 5118 -1372 sw
rect 4976 -1404 5021 -1394
rect 4852 -1432 4926 -1408
rect 4794 -1436 4926 -1432
tri 4926 -1436 4954 -1408 sw
rect 4976 -1418 4978 -1404
tri 4976 -1420 4978 -1418 ne
rect 4990 -1422 5021 -1404
rect 4990 -1432 5036 -1422
rect 5103 -1393 5118 -1378
tri 4728 -1457 4740 -1445 ne
rect 4740 -1450 4750 -1445
tri 4750 -1450 4755 -1445 sw
rect 4639 -1796 4654 -1568
rect 4740 -1558 4755 -1450
rect 4794 -1492 4822 -1436
tri 4914 -1454 4932 -1436 ne
rect 4932 -1456 4954 -1436
tri 4954 -1456 4974 -1436 sw
tri 4990 -1450 5008 -1432 ne
rect 4813 -1526 4822 -1492
rect 4856 -1465 4898 -1464
rect 4856 -1499 4861 -1465
rect 4891 -1499 4898 -1465
rect 4856 -1508 4898 -1499
rect 4932 -1465 4974 -1456
rect 4932 -1499 4939 -1465
rect 4969 -1499 4974 -1465
rect 4932 -1504 4974 -1499
rect 5008 -1492 5036 -1432
tri 5081 -1445 5103 -1423 se
rect 5103 -1430 5118 -1422
tri 5103 -1445 5118 -1430 nw
tri 5075 -1451 5081 -1445 se
rect 5081 -1451 5090 -1445
rect 4794 -1536 4822 -1526
tri 4822 -1536 4846 -1512 sw
rect 4740 -1606 4756 -1558
rect 4794 -1568 4836 -1536
tri 4853 -1544 4854 -1543 sw
rect 4853 -1568 4854 -1544
tri 4856 -1545 4893 -1508 ne
rect 4893 -1536 4898 -1508
tri 4898 -1536 4924 -1510 sw
rect 5008 -1526 5017 -1492
rect 5008 -1536 5036 -1526
rect 4893 -1545 4977 -1536
tri 4893 -1564 4912 -1545 ne
rect 4912 -1564 4977 -1545
rect 4794 -1590 4854 -1568
rect 4976 -1568 4977 -1564
rect 4994 -1568 5036 -1536
rect 4976 -1590 5036 -1568
rect 4882 -1606 4899 -1592
rect 4931 -1606 4948 -1592
tri 4719 -1642 4741 -1620 se
rect 4741 -1627 4756 -1606
tri 4741 -1642 4756 -1627 nw
rect 5075 -1627 5090 -1451
tri 5090 -1458 5103 -1445 nw
rect 5176 -1526 5191 -1298
tri 4713 -1648 4719 -1642 se
rect 4719 -1648 4728 -1642
rect 4713 -1664 4728 -1648
tri 4728 -1655 4741 -1642 nw
rect 4882 -1650 4899 -1636
rect 4931 -1650 4948 -1636
tri 5075 -1642 5090 -1627 ne
tri 5090 -1642 5112 -1620 sw
rect 4713 -1700 4728 -1692
rect 4794 -1664 4854 -1650
rect 4809 -1674 4854 -1664
rect 4809 -1692 4837 -1674
tri 4713 -1715 4728 -1700 ne
tri 4728 -1715 4750 -1693 sw
rect 4794 -1702 4837 -1692
rect 4852 -1678 4854 -1674
rect 4976 -1664 5036 -1650
tri 5090 -1655 5103 -1642 ne
rect 5103 -1648 5112 -1642
tri 5112 -1648 5118 -1642 sw
rect 4976 -1674 5021 -1664
rect 4852 -1702 4926 -1678
rect 4794 -1706 4926 -1702
tri 4926 -1706 4954 -1678 sw
rect 4976 -1688 4978 -1674
tri 4976 -1690 4978 -1688 ne
rect 4990 -1692 5021 -1674
rect 4990 -1702 5036 -1692
rect 5103 -1663 5118 -1648
tri 4728 -1727 4740 -1715 ne
rect 4740 -1720 4750 -1715
tri 4750 -1720 4755 -1715 sw
rect 4639 -2066 4654 -1838
rect 4740 -1876 4755 -1720
rect 4794 -1762 4822 -1706
tri 4914 -1724 4932 -1706 ne
rect 4932 -1726 4954 -1706
tri 4954 -1726 4974 -1706 sw
tri 4990 -1720 5008 -1702 ne
rect 4813 -1796 4822 -1762
rect 4856 -1735 4898 -1734
rect 4856 -1769 4861 -1735
rect 4891 -1769 4898 -1735
rect 4856 -1778 4898 -1769
rect 4932 -1735 4974 -1726
rect 4932 -1769 4939 -1735
rect 4969 -1769 4974 -1735
rect 4932 -1774 4974 -1769
rect 5008 -1762 5036 -1702
tri 5081 -1715 5103 -1693 se
rect 5103 -1700 5118 -1692
tri 5103 -1715 5118 -1700 nw
tri 5075 -1721 5081 -1715 se
rect 5081 -1721 5090 -1715
rect 4794 -1806 4822 -1796
tri 4822 -1806 4846 -1782 sw
rect 4794 -1838 4836 -1806
tri 4853 -1814 4854 -1813 sw
rect 4853 -1838 4854 -1814
tri 4856 -1815 4893 -1778 ne
rect 4893 -1806 4898 -1778
tri 4898 -1806 4924 -1780 sw
rect 5008 -1796 5017 -1762
rect 5008 -1806 5036 -1796
rect 4893 -1815 4977 -1806
tri 4893 -1834 4912 -1815 ne
rect 4912 -1834 4977 -1815
rect 4794 -1860 4854 -1838
rect 4976 -1838 4977 -1834
rect 4994 -1838 5036 -1806
rect 4976 -1860 5036 -1838
rect 4882 -1876 4899 -1862
rect 4931 -1876 4948 -1862
tri 4719 -1912 4741 -1890 se
rect 4741 -1897 4756 -1876
tri 4741 -1912 4756 -1897 nw
rect 5075 -1897 5090 -1721
tri 5090 -1728 5103 -1715 nw
rect 5176 -1796 5191 -1568
tri 4713 -1918 4719 -1912 se
rect 4719 -1918 4728 -1912
rect 4713 -1934 4728 -1918
tri 4728 -1925 4741 -1912 nw
rect 4882 -1920 4899 -1906
rect 4931 -1920 4948 -1906
tri 5075 -1912 5090 -1897 ne
tri 5090 -1912 5112 -1890 sw
rect 4713 -1970 4728 -1962
rect 4794 -1934 4854 -1920
rect 4809 -1944 4854 -1934
rect 4809 -1962 4837 -1944
tri 4713 -1985 4728 -1970 ne
tri 4728 -1985 4750 -1963 sw
rect 4794 -1972 4837 -1962
rect 4852 -1948 4854 -1944
rect 4976 -1934 5036 -1920
tri 5090 -1925 5103 -1912 ne
rect 5103 -1918 5112 -1912
tri 5112 -1918 5118 -1912 sw
rect 4976 -1944 5021 -1934
rect 4852 -1972 4926 -1948
rect 4794 -1976 4926 -1972
tri 4926 -1976 4954 -1948 sw
rect 4976 -1958 4978 -1944
tri 4976 -1960 4978 -1958 ne
rect 4990 -1962 5021 -1944
rect 4990 -1972 5036 -1962
rect 5103 -1933 5118 -1918
tri 4728 -1997 4740 -1985 ne
rect 4740 -1990 4750 -1985
tri 4750 -1990 4755 -1985 sw
rect 4639 -2146 4654 -2108
rect 4740 -2146 4755 -1990
rect 4794 -2032 4822 -1976
tri 4914 -1994 4932 -1976 ne
rect 4932 -1996 4954 -1976
tri 4954 -1996 4974 -1976 sw
tri 4990 -1990 5008 -1972 ne
rect 4813 -2066 4822 -2032
rect 4856 -2005 4898 -2004
rect 4856 -2039 4861 -2005
rect 4891 -2039 4898 -2005
rect 4856 -2048 4898 -2039
rect 4932 -2005 4974 -1996
rect 4932 -2039 4939 -2005
rect 4969 -2039 4974 -2005
rect 4932 -2044 4974 -2039
rect 5008 -2032 5036 -1972
tri 5081 -1985 5103 -1963 se
rect 5103 -1970 5118 -1962
tri 5103 -1985 5118 -1970 nw
tri 5075 -1991 5081 -1985 se
rect 5081 -1991 5090 -1985
rect 4794 -2076 4822 -2066
tri 4822 -2076 4846 -2052 sw
rect 4794 -2108 4836 -2076
tri 4853 -2084 4854 -2083 sw
rect 4853 -2108 4854 -2084
tri 4856 -2085 4893 -2048 ne
rect 4893 -2076 4898 -2048
tri 4898 -2076 4924 -2050 sw
rect 5008 -2066 5017 -2032
rect 5008 -2076 5036 -2066
rect 4893 -2085 4977 -2076
tri 4893 -2104 4912 -2085 ne
rect 4912 -2104 4977 -2085
rect 4794 -2130 4854 -2108
rect 4976 -2108 4977 -2104
rect 4994 -2108 5036 -2076
rect 4976 -2130 5036 -2108
rect 4882 -2146 4899 -2132
rect 4931 -2146 4948 -2132
rect 5075 -2146 5090 -1991
tri 5090 -1998 5103 -1985 nw
rect 5176 -2066 5191 -1838
rect 5176 -2146 5191 -2108
rect 5219 1984 5234 2174
tri 5299 2138 5321 2160 se
rect 5321 2153 5336 2174
tri 5321 2138 5336 2153 nw
rect 5655 2153 5670 2174
tri 5293 2132 5299 2138 se
rect 5299 2132 5308 2138
rect 5293 2116 5308 2132
tri 5308 2125 5321 2138 nw
rect 5462 2130 5479 2144
rect 5511 2130 5528 2144
tri 5655 2138 5670 2153 ne
tri 5670 2138 5692 2160 sw
rect 5293 2080 5308 2088
rect 5374 2116 5434 2130
rect 5389 2106 5434 2116
rect 5389 2088 5417 2106
tri 5293 2065 5308 2080 ne
tri 5308 2065 5330 2087 sw
rect 5374 2078 5417 2088
rect 5432 2102 5434 2106
rect 5556 2116 5616 2130
tri 5670 2125 5683 2138 ne
rect 5683 2132 5692 2138
tri 5692 2132 5698 2138 sw
rect 5556 2106 5601 2116
rect 5432 2078 5506 2102
rect 5374 2074 5506 2078
tri 5506 2074 5534 2102 sw
rect 5556 2092 5558 2106
tri 5556 2090 5558 2092 ne
rect 5570 2088 5601 2106
rect 5570 2078 5616 2088
rect 5683 2117 5698 2132
tri 5308 2053 5320 2065 ne
rect 5320 2060 5330 2065
tri 5330 2060 5335 2065 sw
rect 5219 1714 5234 1942
rect 5320 1904 5335 2060
rect 5374 2018 5402 2074
tri 5494 2056 5512 2074 ne
rect 5512 2054 5534 2074
tri 5534 2054 5554 2074 sw
tri 5570 2060 5588 2078 ne
rect 5393 1984 5402 2018
rect 5436 2045 5478 2046
rect 5436 2011 5441 2045
rect 5471 2011 5478 2045
rect 5436 2002 5478 2011
rect 5512 2045 5554 2054
rect 5512 2011 5519 2045
rect 5549 2011 5554 2045
rect 5512 2006 5554 2011
rect 5588 2018 5616 2078
tri 5661 2065 5683 2087 se
rect 5683 2080 5698 2088
tri 5683 2065 5698 2080 nw
tri 5655 2059 5661 2065 se
rect 5661 2059 5670 2065
rect 5374 1974 5402 1984
tri 5402 1974 5426 1998 sw
rect 5374 1942 5416 1974
tri 5433 1966 5434 1967 sw
rect 5433 1942 5434 1966
tri 5436 1965 5473 2002 ne
rect 5473 1974 5478 2002
tri 5478 1974 5504 2000 sw
rect 5588 1984 5597 2018
rect 5588 1974 5616 1984
rect 5473 1965 5557 1974
tri 5473 1946 5492 1965 ne
rect 5492 1946 5557 1965
rect 5374 1920 5434 1942
rect 5556 1942 5557 1946
rect 5574 1942 5616 1974
rect 5556 1920 5616 1942
rect 5462 1904 5479 1918
rect 5511 1904 5528 1918
tri 5299 1868 5321 1890 se
rect 5321 1883 5336 1904
tri 5321 1868 5336 1883 nw
rect 5655 1883 5670 2059
tri 5670 2052 5683 2065 nw
rect 5756 1984 5771 2174
tri 5293 1862 5299 1868 se
rect 5299 1862 5308 1868
rect 5293 1846 5308 1862
tri 5308 1855 5321 1868 nw
rect 5462 1860 5479 1874
rect 5511 1860 5528 1874
tri 5655 1868 5670 1883 ne
tri 5670 1868 5692 1890 sw
rect 5293 1810 5308 1818
rect 5374 1846 5434 1860
rect 5389 1836 5434 1846
rect 5389 1818 5417 1836
tri 5293 1795 5308 1810 ne
tri 5308 1795 5330 1817 sw
rect 5374 1808 5417 1818
rect 5432 1832 5434 1836
rect 5556 1846 5616 1860
tri 5670 1855 5683 1868 ne
rect 5683 1862 5692 1868
tri 5692 1862 5698 1868 sw
rect 5556 1836 5601 1846
rect 5432 1808 5506 1832
rect 5374 1804 5506 1808
tri 5506 1804 5534 1832 sw
rect 5556 1822 5558 1836
tri 5556 1820 5558 1822 ne
rect 5570 1818 5601 1836
rect 5570 1808 5616 1818
rect 5683 1847 5698 1862
tri 5308 1783 5320 1795 ne
rect 5320 1790 5330 1795
tri 5330 1790 5335 1795 sw
rect 5219 1444 5234 1672
rect 5320 1682 5335 1790
rect 5374 1748 5402 1804
tri 5494 1786 5512 1804 ne
rect 5512 1784 5534 1804
tri 5534 1784 5554 1804 sw
tri 5570 1790 5588 1808 ne
rect 5393 1714 5402 1748
rect 5436 1775 5478 1776
rect 5436 1741 5441 1775
rect 5471 1741 5478 1775
rect 5436 1732 5478 1741
rect 5512 1775 5554 1784
rect 5512 1741 5519 1775
rect 5549 1741 5554 1775
rect 5512 1736 5554 1741
rect 5588 1748 5616 1808
tri 5661 1795 5683 1817 se
rect 5683 1810 5698 1818
tri 5683 1795 5698 1810 nw
tri 5655 1789 5661 1795 se
rect 5661 1789 5670 1795
rect 5374 1704 5402 1714
tri 5402 1704 5426 1728 sw
rect 5320 1634 5336 1682
rect 5374 1672 5416 1704
tri 5433 1696 5434 1697 sw
rect 5433 1672 5434 1696
tri 5436 1695 5473 1732 ne
rect 5473 1704 5478 1732
tri 5478 1704 5504 1730 sw
rect 5588 1714 5597 1748
rect 5588 1704 5616 1714
rect 5473 1695 5557 1704
tri 5473 1676 5492 1695 ne
rect 5492 1676 5557 1695
rect 5374 1650 5434 1672
rect 5556 1672 5557 1676
rect 5574 1672 5616 1704
rect 5556 1650 5616 1672
rect 5462 1634 5479 1648
rect 5511 1634 5528 1648
tri 5299 1598 5321 1620 se
rect 5321 1613 5336 1634
tri 5321 1598 5336 1613 nw
rect 5655 1613 5670 1789
tri 5670 1782 5683 1795 nw
rect 5756 1714 5771 1942
tri 5293 1592 5299 1598 se
rect 5299 1592 5308 1598
rect 5293 1576 5308 1592
tri 5308 1585 5321 1598 nw
rect 5462 1590 5479 1604
rect 5511 1590 5528 1604
tri 5655 1598 5670 1613 ne
tri 5670 1598 5692 1620 sw
rect 5293 1540 5308 1548
rect 5374 1576 5434 1590
rect 5389 1566 5434 1576
rect 5389 1548 5417 1566
tri 5293 1525 5308 1540 ne
tri 5308 1525 5330 1547 sw
rect 5374 1538 5417 1548
rect 5432 1562 5434 1566
rect 5556 1576 5616 1590
tri 5670 1585 5683 1598 ne
rect 5683 1592 5692 1598
tri 5692 1592 5698 1598 sw
rect 5556 1566 5601 1576
rect 5432 1538 5506 1562
rect 5374 1534 5506 1538
tri 5506 1534 5534 1562 sw
rect 5556 1552 5558 1566
tri 5556 1550 5558 1552 ne
rect 5570 1548 5601 1566
rect 5570 1538 5616 1548
rect 5683 1577 5698 1592
tri 5308 1513 5320 1525 ne
rect 5320 1520 5330 1525
tri 5330 1520 5335 1525 sw
rect 5219 1174 5234 1402
rect 5320 1364 5335 1520
rect 5374 1478 5402 1534
tri 5494 1516 5512 1534 ne
rect 5512 1514 5534 1534
tri 5534 1514 5554 1534 sw
tri 5570 1520 5588 1538 ne
rect 5393 1444 5402 1478
rect 5436 1505 5478 1506
rect 5436 1471 5441 1505
rect 5471 1471 5478 1505
rect 5436 1462 5478 1471
rect 5512 1505 5554 1514
rect 5512 1471 5519 1505
rect 5549 1471 5554 1505
rect 5512 1466 5554 1471
rect 5588 1478 5616 1538
tri 5661 1525 5683 1547 se
rect 5683 1540 5698 1548
tri 5683 1525 5698 1540 nw
tri 5655 1519 5661 1525 se
rect 5661 1519 5670 1525
rect 5374 1434 5402 1444
tri 5402 1434 5426 1458 sw
rect 5374 1402 5416 1434
tri 5433 1426 5434 1427 sw
rect 5433 1402 5434 1426
tri 5436 1425 5473 1462 ne
rect 5473 1434 5478 1462
tri 5478 1434 5504 1460 sw
rect 5588 1444 5597 1478
rect 5588 1434 5616 1444
rect 5473 1425 5557 1434
tri 5473 1406 5492 1425 ne
rect 5492 1406 5557 1425
rect 5374 1380 5434 1402
rect 5556 1402 5557 1406
rect 5574 1402 5616 1434
rect 5556 1380 5616 1402
rect 5462 1364 5479 1378
rect 5511 1364 5528 1378
tri 5299 1328 5321 1350 se
rect 5321 1343 5336 1364
tri 5321 1328 5336 1343 nw
rect 5655 1343 5670 1519
tri 5670 1512 5683 1525 nw
rect 5756 1444 5771 1672
tri 5293 1322 5299 1328 se
rect 5299 1322 5308 1328
rect 5293 1306 5308 1322
tri 5308 1315 5321 1328 nw
rect 5462 1320 5479 1334
rect 5511 1320 5528 1334
tri 5655 1328 5670 1343 ne
tri 5670 1328 5692 1350 sw
rect 5293 1270 5308 1278
rect 5374 1306 5434 1320
rect 5389 1296 5434 1306
rect 5389 1278 5417 1296
tri 5293 1255 5308 1270 ne
tri 5308 1255 5330 1277 sw
rect 5374 1268 5417 1278
rect 5432 1292 5434 1296
rect 5556 1306 5616 1320
tri 5670 1315 5683 1328 ne
rect 5683 1322 5692 1328
tri 5692 1322 5698 1328 sw
rect 5556 1296 5601 1306
rect 5432 1268 5506 1292
rect 5374 1264 5506 1268
tri 5506 1264 5534 1292 sw
rect 5556 1282 5558 1296
tri 5556 1280 5558 1282 ne
rect 5570 1278 5601 1296
rect 5570 1268 5616 1278
rect 5683 1307 5698 1322
tri 5308 1243 5320 1255 ne
rect 5320 1250 5330 1255
tri 5330 1250 5335 1255 sw
rect 5219 904 5234 1132
rect 5320 1142 5335 1250
rect 5374 1208 5402 1264
tri 5494 1246 5512 1264 ne
rect 5512 1244 5534 1264
tri 5534 1244 5554 1264 sw
tri 5570 1250 5588 1268 ne
rect 5393 1174 5402 1208
rect 5436 1235 5478 1236
rect 5436 1201 5441 1235
rect 5471 1201 5478 1235
rect 5436 1192 5478 1201
rect 5512 1235 5554 1244
rect 5512 1201 5519 1235
rect 5549 1201 5554 1235
rect 5512 1196 5554 1201
rect 5588 1208 5616 1268
tri 5661 1255 5683 1277 se
rect 5683 1270 5698 1278
tri 5683 1255 5698 1270 nw
tri 5655 1249 5661 1255 se
rect 5661 1249 5670 1255
rect 5374 1164 5402 1174
tri 5402 1164 5426 1188 sw
rect 5320 1094 5336 1142
rect 5374 1132 5416 1164
tri 5433 1156 5434 1157 sw
rect 5433 1132 5434 1156
tri 5436 1155 5473 1192 ne
rect 5473 1164 5478 1192
tri 5478 1164 5504 1190 sw
rect 5588 1174 5597 1208
rect 5588 1164 5616 1174
rect 5473 1155 5557 1164
tri 5473 1136 5492 1155 ne
rect 5492 1136 5557 1155
rect 5374 1110 5434 1132
rect 5556 1132 5557 1136
rect 5574 1132 5616 1164
rect 5556 1110 5616 1132
rect 5462 1094 5479 1108
rect 5511 1094 5528 1108
tri 5299 1058 5321 1080 se
rect 5321 1073 5336 1094
tri 5321 1058 5336 1073 nw
rect 5655 1073 5670 1249
tri 5670 1242 5683 1255 nw
rect 5756 1174 5771 1402
tri 5293 1052 5299 1058 se
rect 5299 1052 5308 1058
rect 5293 1036 5308 1052
tri 5308 1045 5321 1058 nw
rect 5462 1050 5479 1064
rect 5511 1050 5528 1064
tri 5655 1058 5670 1073 ne
tri 5670 1058 5692 1080 sw
rect 5293 1000 5308 1008
rect 5374 1036 5434 1050
rect 5389 1026 5434 1036
rect 5389 1008 5417 1026
tri 5293 985 5308 1000 ne
tri 5308 985 5330 1007 sw
rect 5374 998 5417 1008
rect 5432 1022 5434 1026
rect 5556 1036 5616 1050
tri 5670 1045 5683 1058 ne
rect 5683 1052 5692 1058
tri 5692 1052 5698 1058 sw
rect 5556 1026 5601 1036
rect 5432 998 5506 1022
rect 5374 994 5506 998
tri 5506 994 5534 1022 sw
rect 5556 1012 5558 1026
tri 5556 1010 5558 1012 ne
rect 5570 1008 5601 1026
rect 5570 998 5616 1008
rect 5683 1037 5698 1052
tri 5308 973 5320 985 ne
rect 5320 980 5330 985
tri 5330 980 5335 985 sw
rect 5219 634 5234 862
rect 5320 824 5335 980
rect 5374 938 5402 994
tri 5494 976 5512 994 ne
rect 5512 974 5534 994
tri 5534 974 5554 994 sw
tri 5570 980 5588 998 ne
rect 5393 904 5402 938
rect 5436 965 5478 966
rect 5436 931 5441 965
rect 5471 931 5478 965
rect 5436 922 5478 931
rect 5512 965 5554 974
rect 5512 931 5519 965
rect 5549 931 5554 965
rect 5512 926 5554 931
rect 5588 938 5616 998
tri 5661 985 5683 1007 se
rect 5683 1000 5698 1008
tri 5683 985 5698 1000 nw
tri 5655 979 5661 985 se
rect 5661 979 5670 985
rect 5374 894 5402 904
tri 5402 894 5426 918 sw
rect 5374 862 5416 894
tri 5433 886 5434 887 sw
rect 5433 862 5434 886
tri 5436 885 5473 922 ne
rect 5473 894 5478 922
tri 5478 894 5504 920 sw
rect 5588 904 5597 938
rect 5588 894 5616 904
rect 5473 885 5557 894
tri 5473 866 5492 885 ne
rect 5492 866 5557 885
rect 5374 840 5434 862
rect 5556 862 5557 866
rect 5574 862 5616 894
rect 5556 840 5616 862
rect 5462 824 5479 838
rect 5511 824 5528 838
tri 5299 788 5321 810 se
rect 5321 803 5336 824
tri 5321 788 5336 803 nw
rect 5655 803 5670 979
tri 5670 972 5683 985 nw
rect 5756 904 5771 1132
tri 5293 782 5299 788 se
rect 5299 782 5308 788
rect 5293 766 5308 782
tri 5308 775 5321 788 nw
rect 5462 780 5479 794
rect 5511 780 5528 794
tri 5655 788 5670 803 ne
tri 5670 788 5692 810 sw
rect 5293 730 5308 738
rect 5374 766 5434 780
rect 5389 756 5434 766
rect 5389 738 5417 756
tri 5293 715 5308 730 ne
tri 5308 715 5330 737 sw
rect 5374 728 5417 738
rect 5432 752 5434 756
rect 5556 766 5616 780
tri 5670 775 5683 788 ne
rect 5683 782 5692 788
tri 5692 782 5698 788 sw
rect 5556 756 5601 766
rect 5432 728 5506 752
rect 5374 724 5506 728
tri 5506 724 5534 752 sw
rect 5556 742 5558 756
tri 5556 740 5558 742 ne
rect 5570 738 5601 756
rect 5570 728 5616 738
rect 5683 767 5698 782
tri 5308 703 5320 715 ne
rect 5320 710 5330 715
tri 5330 710 5335 715 sw
rect 5219 364 5234 592
rect 5320 602 5335 710
rect 5374 668 5402 724
tri 5494 706 5512 724 ne
rect 5512 704 5534 724
tri 5534 704 5554 724 sw
tri 5570 710 5588 728 ne
rect 5393 634 5402 668
rect 5436 695 5478 696
rect 5436 661 5441 695
rect 5471 661 5478 695
rect 5436 652 5478 661
rect 5512 695 5554 704
rect 5512 661 5519 695
rect 5549 661 5554 695
rect 5512 656 5554 661
rect 5588 668 5616 728
tri 5661 715 5683 737 se
rect 5683 730 5698 738
tri 5683 715 5698 730 nw
tri 5655 709 5661 715 se
rect 5661 709 5670 715
rect 5374 624 5402 634
tri 5402 624 5426 648 sw
rect 5320 554 5336 602
rect 5374 592 5416 624
tri 5433 616 5434 617 sw
rect 5433 592 5434 616
tri 5436 615 5473 652 ne
rect 5473 624 5478 652
tri 5478 624 5504 650 sw
rect 5588 634 5597 668
rect 5588 624 5616 634
rect 5473 615 5557 624
tri 5473 596 5492 615 ne
rect 5492 596 5557 615
rect 5374 570 5434 592
rect 5556 592 5557 596
rect 5574 592 5616 624
rect 5556 570 5616 592
rect 5462 554 5479 568
rect 5511 554 5528 568
tri 5299 518 5321 540 se
rect 5321 533 5336 554
tri 5321 518 5336 533 nw
rect 5655 533 5670 709
tri 5670 702 5683 715 nw
rect 5756 634 5771 862
tri 5293 512 5299 518 se
rect 5299 512 5308 518
rect 5293 496 5308 512
tri 5308 505 5321 518 nw
rect 5462 510 5479 524
rect 5511 510 5528 524
tri 5655 518 5670 533 ne
tri 5670 518 5692 540 sw
rect 5293 460 5308 468
rect 5374 496 5434 510
rect 5389 486 5434 496
rect 5389 468 5417 486
tri 5293 445 5308 460 ne
tri 5308 445 5330 467 sw
rect 5374 458 5417 468
rect 5432 482 5434 486
rect 5556 496 5616 510
tri 5670 505 5683 518 ne
rect 5683 512 5692 518
tri 5692 512 5698 518 sw
rect 5556 486 5601 496
rect 5432 458 5506 482
rect 5374 454 5506 458
tri 5506 454 5534 482 sw
rect 5556 472 5558 486
tri 5556 470 5558 472 ne
rect 5570 468 5601 486
rect 5570 458 5616 468
rect 5683 497 5698 512
tri 5308 433 5320 445 ne
rect 5320 440 5330 445
tri 5330 440 5335 445 sw
rect 5219 94 5234 322
rect 5320 284 5335 440
rect 5374 398 5402 454
tri 5494 436 5512 454 ne
rect 5512 434 5534 454
tri 5534 434 5554 454 sw
tri 5570 440 5588 458 ne
rect 5393 364 5402 398
rect 5436 425 5478 426
rect 5436 391 5441 425
rect 5471 391 5478 425
rect 5436 382 5478 391
rect 5512 425 5554 434
rect 5512 391 5519 425
rect 5549 391 5554 425
rect 5512 386 5554 391
rect 5588 398 5616 458
tri 5661 445 5683 467 se
rect 5683 460 5698 468
tri 5683 445 5698 460 nw
tri 5655 439 5661 445 se
rect 5661 439 5670 445
rect 5374 354 5402 364
tri 5402 354 5426 378 sw
rect 5374 322 5416 354
tri 5433 346 5434 347 sw
rect 5433 322 5434 346
tri 5436 345 5473 382 ne
rect 5473 354 5478 382
tri 5478 354 5504 380 sw
rect 5588 364 5597 398
rect 5588 354 5616 364
rect 5473 345 5557 354
tri 5473 326 5492 345 ne
rect 5492 326 5557 345
rect 5374 300 5434 322
rect 5556 322 5557 326
rect 5574 322 5616 354
rect 5556 300 5616 322
rect 5462 284 5479 298
rect 5511 284 5528 298
tri 5299 248 5321 270 se
rect 5321 263 5336 284
tri 5321 248 5336 263 nw
rect 5655 263 5670 439
tri 5670 432 5683 445 nw
rect 5756 364 5771 592
tri 5293 242 5299 248 se
rect 5299 242 5308 248
rect 5293 226 5308 242
tri 5308 235 5321 248 nw
rect 5462 240 5479 254
rect 5511 240 5528 254
tri 5655 248 5670 263 ne
tri 5670 248 5692 270 sw
rect 5293 190 5308 198
rect 5374 226 5434 240
rect 5389 216 5434 226
rect 5389 198 5417 216
tri 5293 175 5308 190 ne
tri 5308 175 5330 197 sw
rect 5374 188 5417 198
rect 5432 212 5434 216
rect 5556 226 5616 240
tri 5670 235 5683 248 ne
rect 5683 242 5692 248
tri 5692 242 5698 248 sw
rect 5556 216 5601 226
rect 5432 188 5506 212
rect 5374 184 5506 188
tri 5506 184 5534 212 sw
rect 5556 202 5558 216
tri 5556 200 5558 202 ne
rect 5570 198 5601 216
rect 5570 188 5616 198
rect 5683 227 5698 242
tri 5308 163 5320 175 ne
rect 5320 170 5330 175
tri 5330 170 5335 175 sw
rect 5219 -176 5234 52
rect 5320 62 5335 170
rect 5374 128 5402 184
tri 5494 166 5512 184 ne
rect 5512 164 5534 184
tri 5534 164 5554 184 sw
tri 5570 170 5588 188 ne
rect 5393 94 5402 128
rect 5436 155 5478 156
rect 5436 121 5441 155
rect 5471 121 5478 155
rect 5436 112 5478 121
rect 5512 155 5554 164
rect 5512 121 5519 155
rect 5549 121 5554 155
rect 5512 116 5554 121
rect 5588 128 5616 188
tri 5661 175 5683 197 se
rect 5683 190 5698 198
tri 5683 175 5698 190 nw
tri 5655 169 5661 175 se
rect 5661 169 5670 175
rect 5374 84 5402 94
tri 5402 84 5426 108 sw
rect 5320 14 5336 62
rect 5374 52 5416 84
tri 5433 76 5434 77 sw
rect 5433 52 5434 76
tri 5436 75 5473 112 ne
rect 5473 84 5478 112
tri 5478 84 5504 110 sw
rect 5588 94 5597 128
rect 5588 84 5616 94
rect 5473 75 5557 84
tri 5473 56 5492 75 ne
rect 5492 56 5557 75
rect 5374 30 5434 52
rect 5556 52 5557 56
rect 5574 52 5616 84
rect 5556 30 5616 52
rect 5462 14 5479 28
rect 5511 14 5528 28
tri 5299 -22 5321 0 se
rect 5321 -7 5336 14
tri 5321 -22 5336 -7 nw
rect 5655 -7 5670 169
tri 5670 162 5683 175 nw
rect 5756 94 5771 322
tri 5293 -28 5299 -22 se
rect 5299 -28 5308 -22
rect 5293 -44 5308 -28
tri 5308 -35 5321 -22 nw
rect 5462 -30 5479 -16
rect 5511 -30 5528 -16
tri 5655 -22 5670 -7 ne
tri 5670 -22 5692 0 sw
rect 5293 -80 5308 -72
rect 5374 -44 5434 -30
rect 5389 -54 5434 -44
rect 5389 -72 5417 -54
tri 5293 -95 5308 -80 ne
tri 5308 -95 5330 -73 sw
rect 5374 -82 5417 -72
rect 5432 -58 5434 -54
rect 5556 -44 5616 -30
tri 5670 -35 5683 -22 ne
rect 5683 -28 5692 -22
tri 5692 -28 5698 -22 sw
rect 5556 -54 5601 -44
rect 5432 -82 5506 -58
rect 5374 -86 5506 -82
tri 5506 -86 5534 -58 sw
rect 5556 -68 5558 -54
tri 5556 -70 5558 -68 ne
rect 5570 -72 5601 -54
rect 5570 -82 5616 -72
rect 5683 -43 5698 -28
tri 5308 -107 5320 -95 ne
rect 5320 -100 5330 -95
tri 5330 -100 5335 -95 sw
rect 5219 -446 5234 -218
rect 5320 -256 5335 -100
rect 5374 -142 5402 -86
tri 5494 -104 5512 -86 ne
rect 5512 -106 5534 -86
tri 5534 -106 5554 -86 sw
tri 5570 -100 5588 -82 ne
rect 5393 -176 5402 -142
rect 5436 -115 5478 -114
rect 5436 -149 5441 -115
rect 5471 -149 5478 -115
rect 5436 -158 5478 -149
rect 5512 -115 5554 -106
rect 5512 -149 5519 -115
rect 5549 -149 5554 -115
rect 5512 -154 5554 -149
rect 5588 -142 5616 -82
tri 5661 -95 5683 -73 se
rect 5683 -80 5698 -72
tri 5683 -95 5698 -80 nw
tri 5655 -101 5661 -95 se
rect 5661 -101 5670 -95
rect 5374 -186 5402 -176
tri 5402 -186 5426 -162 sw
rect 5374 -218 5416 -186
tri 5433 -194 5434 -193 sw
rect 5433 -218 5434 -194
tri 5436 -195 5473 -158 ne
rect 5473 -186 5478 -158
tri 5478 -186 5504 -160 sw
rect 5588 -176 5597 -142
rect 5588 -186 5616 -176
rect 5473 -195 5557 -186
tri 5473 -214 5492 -195 ne
rect 5492 -214 5557 -195
rect 5374 -240 5434 -218
rect 5556 -218 5557 -214
rect 5574 -218 5616 -186
rect 5556 -240 5616 -218
rect 5462 -256 5479 -242
rect 5511 -256 5528 -242
tri 5299 -292 5321 -270 se
rect 5321 -277 5336 -256
tri 5321 -292 5336 -277 nw
rect 5655 -277 5670 -101
tri 5670 -108 5683 -95 nw
rect 5756 -176 5771 52
tri 5293 -298 5299 -292 se
rect 5299 -298 5308 -292
rect 5293 -314 5308 -298
tri 5308 -305 5321 -292 nw
rect 5462 -300 5479 -286
rect 5511 -300 5528 -286
tri 5655 -292 5670 -277 ne
tri 5670 -292 5692 -270 sw
rect 5293 -350 5308 -342
rect 5374 -314 5434 -300
rect 5389 -324 5434 -314
rect 5389 -342 5417 -324
tri 5293 -365 5308 -350 ne
tri 5308 -365 5330 -343 sw
rect 5374 -352 5417 -342
rect 5432 -328 5434 -324
rect 5556 -314 5616 -300
tri 5670 -305 5683 -292 ne
rect 5683 -298 5692 -292
tri 5692 -298 5698 -292 sw
rect 5556 -324 5601 -314
rect 5432 -352 5506 -328
rect 5374 -356 5506 -352
tri 5506 -356 5534 -328 sw
rect 5556 -338 5558 -324
tri 5556 -340 5558 -338 ne
rect 5570 -342 5601 -324
rect 5570 -352 5616 -342
rect 5683 -313 5698 -298
tri 5308 -377 5320 -365 ne
rect 5320 -370 5330 -365
tri 5330 -370 5335 -365 sw
rect 5219 -716 5234 -488
rect 5320 -478 5335 -370
rect 5374 -412 5402 -356
tri 5494 -374 5512 -356 ne
rect 5512 -376 5534 -356
tri 5534 -376 5554 -356 sw
tri 5570 -370 5588 -352 ne
rect 5393 -446 5402 -412
rect 5436 -385 5478 -384
rect 5436 -419 5441 -385
rect 5471 -419 5478 -385
rect 5436 -428 5478 -419
rect 5512 -385 5554 -376
rect 5512 -419 5519 -385
rect 5549 -419 5554 -385
rect 5512 -424 5554 -419
rect 5588 -412 5616 -352
tri 5661 -365 5683 -343 se
rect 5683 -350 5698 -342
tri 5683 -365 5698 -350 nw
tri 5655 -371 5661 -365 se
rect 5661 -371 5670 -365
rect 5374 -456 5402 -446
tri 5402 -456 5426 -432 sw
rect 5320 -526 5336 -478
rect 5374 -488 5416 -456
tri 5433 -464 5434 -463 sw
rect 5433 -488 5434 -464
tri 5436 -465 5473 -428 ne
rect 5473 -456 5478 -428
tri 5478 -456 5504 -430 sw
rect 5588 -446 5597 -412
rect 5588 -456 5616 -446
rect 5473 -465 5557 -456
tri 5473 -484 5492 -465 ne
rect 5492 -484 5557 -465
rect 5374 -510 5434 -488
rect 5556 -488 5557 -484
rect 5574 -488 5616 -456
rect 5556 -510 5616 -488
rect 5462 -526 5479 -512
rect 5511 -526 5528 -512
tri 5299 -562 5321 -540 se
rect 5321 -547 5336 -526
tri 5321 -562 5336 -547 nw
rect 5655 -547 5670 -371
tri 5670 -378 5683 -365 nw
rect 5756 -446 5771 -218
tri 5293 -568 5299 -562 se
rect 5299 -568 5308 -562
rect 5293 -584 5308 -568
tri 5308 -575 5321 -562 nw
rect 5462 -570 5479 -556
rect 5511 -570 5528 -556
tri 5655 -562 5670 -547 ne
tri 5670 -562 5692 -540 sw
rect 5293 -620 5308 -612
rect 5374 -584 5434 -570
rect 5389 -594 5434 -584
rect 5389 -612 5417 -594
tri 5293 -635 5308 -620 ne
tri 5308 -635 5330 -613 sw
rect 5374 -622 5417 -612
rect 5432 -598 5434 -594
rect 5556 -584 5616 -570
tri 5670 -575 5683 -562 ne
rect 5683 -568 5692 -562
tri 5692 -568 5698 -562 sw
rect 5556 -594 5601 -584
rect 5432 -622 5506 -598
rect 5374 -626 5506 -622
tri 5506 -626 5534 -598 sw
rect 5556 -608 5558 -594
tri 5556 -610 5558 -608 ne
rect 5570 -612 5601 -594
rect 5570 -622 5616 -612
rect 5683 -583 5698 -568
tri 5308 -647 5320 -635 ne
rect 5320 -640 5330 -635
tri 5330 -640 5335 -635 sw
rect 5219 -986 5234 -758
rect 5320 -796 5335 -640
rect 5374 -682 5402 -626
tri 5494 -644 5512 -626 ne
rect 5512 -646 5534 -626
tri 5534 -646 5554 -626 sw
tri 5570 -640 5588 -622 ne
rect 5393 -716 5402 -682
rect 5436 -655 5478 -654
rect 5436 -689 5441 -655
rect 5471 -689 5478 -655
rect 5436 -698 5478 -689
rect 5512 -655 5554 -646
rect 5512 -689 5519 -655
rect 5549 -689 5554 -655
rect 5512 -694 5554 -689
rect 5588 -682 5616 -622
tri 5661 -635 5683 -613 se
rect 5683 -620 5698 -612
tri 5683 -635 5698 -620 nw
tri 5655 -641 5661 -635 se
rect 5661 -641 5670 -635
rect 5374 -726 5402 -716
tri 5402 -726 5426 -702 sw
rect 5374 -758 5416 -726
tri 5433 -734 5434 -733 sw
rect 5433 -758 5434 -734
tri 5436 -735 5473 -698 ne
rect 5473 -726 5478 -698
tri 5478 -726 5504 -700 sw
rect 5588 -716 5597 -682
rect 5588 -726 5616 -716
rect 5473 -735 5557 -726
tri 5473 -754 5492 -735 ne
rect 5492 -754 5557 -735
rect 5374 -780 5434 -758
rect 5556 -758 5557 -754
rect 5574 -758 5616 -726
rect 5556 -780 5616 -758
rect 5462 -796 5479 -782
rect 5511 -796 5528 -782
tri 5299 -832 5321 -810 se
rect 5321 -817 5336 -796
tri 5321 -832 5336 -817 nw
rect 5655 -817 5670 -641
tri 5670 -648 5683 -635 nw
rect 5756 -716 5771 -488
tri 5293 -838 5299 -832 se
rect 5299 -838 5308 -832
rect 5293 -854 5308 -838
tri 5308 -845 5321 -832 nw
rect 5462 -840 5479 -826
rect 5511 -840 5528 -826
tri 5655 -832 5670 -817 ne
tri 5670 -832 5692 -810 sw
rect 5293 -890 5308 -882
rect 5374 -854 5434 -840
rect 5389 -864 5434 -854
rect 5389 -882 5417 -864
tri 5293 -905 5308 -890 ne
tri 5308 -905 5330 -883 sw
rect 5374 -892 5417 -882
rect 5432 -868 5434 -864
rect 5556 -854 5616 -840
tri 5670 -845 5683 -832 ne
rect 5683 -838 5692 -832
tri 5692 -838 5698 -832 sw
rect 5556 -864 5601 -854
rect 5432 -892 5506 -868
rect 5374 -896 5506 -892
tri 5506 -896 5534 -868 sw
rect 5556 -878 5558 -864
tri 5556 -880 5558 -878 ne
rect 5570 -882 5601 -864
rect 5570 -892 5616 -882
rect 5683 -853 5698 -838
tri 5308 -917 5320 -905 ne
rect 5320 -910 5330 -905
tri 5330 -910 5335 -905 sw
rect 5219 -1256 5234 -1028
rect 5320 -1018 5335 -910
rect 5374 -952 5402 -896
tri 5494 -914 5512 -896 ne
rect 5512 -916 5534 -896
tri 5534 -916 5554 -896 sw
tri 5570 -910 5588 -892 ne
rect 5393 -986 5402 -952
rect 5436 -925 5478 -924
rect 5436 -959 5441 -925
rect 5471 -959 5478 -925
rect 5436 -968 5478 -959
rect 5512 -925 5554 -916
rect 5512 -959 5519 -925
rect 5549 -959 5554 -925
rect 5512 -964 5554 -959
rect 5588 -952 5616 -892
tri 5661 -905 5683 -883 se
rect 5683 -890 5698 -882
tri 5683 -905 5698 -890 nw
tri 5655 -911 5661 -905 se
rect 5661 -911 5670 -905
rect 5374 -996 5402 -986
tri 5402 -996 5426 -972 sw
rect 5320 -1066 5336 -1018
rect 5374 -1028 5416 -996
tri 5433 -1004 5434 -1003 sw
rect 5433 -1028 5434 -1004
tri 5436 -1005 5473 -968 ne
rect 5473 -996 5478 -968
tri 5478 -996 5504 -970 sw
rect 5588 -986 5597 -952
rect 5588 -996 5616 -986
rect 5473 -1005 5557 -996
tri 5473 -1024 5492 -1005 ne
rect 5492 -1024 5557 -1005
rect 5374 -1050 5434 -1028
rect 5556 -1028 5557 -1024
rect 5574 -1028 5616 -996
rect 5556 -1050 5616 -1028
rect 5462 -1066 5479 -1052
rect 5511 -1066 5528 -1052
tri 5299 -1102 5321 -1080 se
rect 5321 -1087 5336 -1066
tri 5321 -1102 5336 -1087 nw
rect 5655 -1087 5670 -911
tri 5670 -918 5683 -905 nw
rect 5756 -986 5771 -758
tri 5293 -1108 5299 -1102 se
rect 5299 -1108 5308 -1102
rect 5293 -1124 5308 -1108
tri 5308 -1115 5321 -1102 nw
rect 5462 -1110 5479 -1096
rect 5511 -1110 5528 -1096
tri 5655 -1102 5670 -1087 ne
tri 5670 -1102 5692 -1080 sw
rect 5293 -1160 5308 -1152
rect 5374 -1124 5434 -1110
rect 5389 -1134 5434 -1124
rect 5389 -1152 5417 -1134
tri 5293 -1175 5308 -1160 ne
tri 5308 -1175 5330 -1153 sw
rect 5374 -1162 5417 -1152
rect 5432 -1138 5434 -1134
rect 5556 -1124 5616 -1110
tri 5670 -1115 5683 -1102 ne
rect 5683 -1108 5692 -1102
tri 5692 -1108 5698 -1102 sw
rect 5556 -1134 5601 -1124
rect 5432 -1162 5506 -1138
rect 5374 -1166 5506 -1162
tri 5506 -1166 5534 -1138 sw
rect 5556 -1148 5558 -1134
tri 5556 -1150 5558 -1148 ne
rect 5570 -1152 5601 -1134
rect 5570 -1162 5616 -1152
rect 5683 -1123 5698 -1108
tri 5308 -1187 5320 -1175 ne
rect 5320 -1180 5330 -1175
tri 5330 -1180 5335 -1175 sw
rect 5219 -1526 5234 -1298
rect 5320 -1336 5335 -1180
rect 5374 -1222 5402 -1166
tri 5494 -1184 5512 -1166 ne
rect 5512 -1186 5534 -1166
tri 5534 -1186 5554 -1166 sw
tri 5570 -1180 5588 -1162 ne
rect 5393 -1256 5402 -1222
rect 5436 -1195 5478 -1194
rect 5436 -1229 5441 -1195
rect 5471 -1229 5478 -1195
rect 5436 -1238 5478 -1229
rect 5512 -1195 5554 -1186
rect 5512 -1229 5519 -1195
rect 5549 -1229 5554 -1195
rect 5512 -1234 5554 -1229
rect 5588 -1222 5616 -1162
tri 5661 -1175 5683 -1153 se
rect 5683 -1160 5698 -1152
tri 5683 -1175 5698 -1160 nw
tri 5655 -1181 5661 -1175 se
rect 5661 -1181 5670 -1175
rect 5374 -1266 5402 -1256
tri 5402 -1266 5426 -1242 sw
rect 5374 -1298 5416 -1266
tri 5433 -1274 5434 -1273 sw
rect 5433 -1298 5434 -1274
tri 5436 -1275 5473 -1238 ne
rect 5473 -1266 5478 -1238
tri 5478 -1266 5504 -1240 sw
rect 5588 -1256 5597 -1222
rect 5588 -1266 5616 -1256
rect 5473 -1275 5557 -1266
tri 5473 -1294 5492 -1275 ne
rect 5492 -1294 5557 -1275
rect 5374 -1320 5434 -1298
rect 5556 -1298 5557 -1294
rect 5574 -1298 5616 -1266
rect 5556 -1320 5616 -1298
rect 5462 -1336 5479 -1322
rect 5511 -1336 5528 -1322
tri 5299 -1372 5321 -1350 se
rect 5321 -1357 5336 -1336
tri 5321 -1372 5336 -1357 nw
rect 5655 -1357 5670 -1181
tri 5670 -1188 5683 -1175 nw
rect 5756 -1256 5771 -1028
tri 5293 -1378 5299 -1372 se
rect 5299 -1378 5308 -1372
rect 5293 -1394 5308 -1378
tri 5308 -1385 5321 -1372 nw
rect 5462 -1380 5479 -1366
rect 5511 -1380 5528 -1366
tri 5655 -1372 5670 -1357 ne
tri 5670 -1372 5692 -1350 sw
rect 5293 -1430 5308 -1422
rect 5374 -1394 5434 -1380
rect 5389 -1404 5434 -1394
rect 5389 -1422 5417 -1404
tri 5293 -1445 5308 -1430 ne
tri 5308 -1445 5330 -1423 sw
rect 5374 -1432 5417 -1422
rect 5432 -1408 5434 -1404
rect 5556 -1394 5616 -1380
tri 5670 -1385 5683 -1372 ne
rect 5683 -1378 5692 -1372
tri 5692 -1378 5698 -1372 sw
rect 5556 -1404 5601 -1394
rect 5432 -1432 5506 -1408
rect 5374 -1436 5506 -1432
tri 5506 -1436 5534 -1408 sw
rect 5556 -1418 5558 -1404
tri 5556 -1420 5558 -1418 ne
rect 5570 -1422 5601 -1404
rect 5570 -1432 5616 -1422
rect 5683 -1393 5698 -1378
tri 5308 -1457 5320 -1445 ne
rect 5320 -1450 5330 -1445
tri 5330 -1450 5335 -1445 sw
rect 5219 -1796 5234 -1568
rect 5320 -1558 5335 -1450
rect 5374 -1492 5402 -1436
tri 5494 -1454 5512 -1436 ne
rect 5512 -1456 5534 -1436
tri 5534 -1456 5554 -1436 sw
tri 5570 -1450 5588 -1432 ne
rect 5393 -1526 5402 -1492
rect 5436 -1465 5478 -1464
rect 5436 -1499 5441 -1465
rect 5471 -1499 5478 -1465
rect 5436 -1508 5478 -1499
rect 5512 -1465 5554 -1456
rect 5512 -1499 5519 -1465
rect 5549 -1499 5554 -1465
rect 5512 -1504 5554 -1499
rect 5588 -1492 5616 -1432
tri 5661 -1445 5683 -1423 se
rect 5683 -1430 5698 -1422
tri 5683 -1445 5698 -1430 nw
tri 5655 -1451 5661 -1445 se
rect 5661 -1451 5670 -1445
rect 5374 -1536 5402 -1526
tri 5402 -1536 5426 -1512 sw
rect 5320 -1606 5336 -1558
rect 5374 -1568 5416 -1536
tri 5433 -1544 5434 -1543 sw
rect 5433 -1568 5434 -1544
tri 5436 -1545 5473 -1508 ne
rect 5473 -1536 5478 -1508
tri 5478 -1536 5504 -1510 sw
rect 5588 -1526 5597 -1492
rect 5588 -1536 5616 -1526
rect 5473 -1545 5557 -1536
tri 5473 -1564 5492 -1545 ne
rect 5492 -1564 5557 -1545
rect 5374 -1590 5434 -1568
rect 5556 -1568 5557 -1564
rect 5574 -1568 5616 -1536
rect 5556 -1590 5616 -1568
rect 5462 -1606 5479 -1592
rect 5511 -1606 5528 -1592
tri 5299 -1642 5321 -1620 se
rect 5321 -1627 5336 -1606
tri 5321 -1642 5336 -1627 nw
rect 5655 -1627 5670 -1451
tri 5670 -1458 5683 -1445 nw
rect 5756 -1526 5771 -1298
tri 5293 -1648 5299 -1642 se
rect 5299 -1648 5308 -1642
rect 5293 -1664 5308 -1648
tri 5308 -1655 5321 -1642 nw
rect 5462 -1650 5479 -1636
rect 5511 -1650 5528 -1636
tri 5655 -1642 5670 -1627 ne
tri 5670 -1642 5692 -1620 sw
rect 5293 -1700 5308 -1692
rect 5374 -1664 5434 -1650
rect 5389 -1674 5434 -1664
rect 5389 -1692 5417 -1674
tri 5293 -1715 5308 -1700 ne
tri 5308 -1715 5330 -1693 sw
rect 5374 -1702 5417 -1692
rect 5432 -1678 5434 -1674
rect 5556 -1664 5616 -1650
tri 5670 -1655 5683 -1642 ne
rect 5683 -1648 5692 -1642
tri 5692 -1648 5698 -1642 sw
rect 5556 -1674 5601 -1664
rect 5432 -1702 5506 -1678
rect 5374 -1706 5506 -1702
tri 5506 -1706 5534 -1678 sw
rect 5556 -1688 5558 -1674
tri 5556 -1690 5558 -1688 ne
rect 5570 -1692 5601 -1674
rect 5570 -1702 5616 -1692
rect 5683 -1663 5698 -1648
tri 5308 -1727 5320 -1715 ne
rect 5320 -1720 5330 -1715
tri 5330 -1720 5335 -1715 sw
rect 5219 -2066 5234 -1838
rect 5320 -1876 5335 -1720
rect 5374 -1762 5402 -1706
tri 5494 -1724 5512 -1706 ne
rect 5512 -1726 5534 -1706
tri 5534 -1726 5554 -1706 sw
tri 5570 -1720 5588 -1702 ne
rect 5393 -1796 5402 -1762
rect 5436 -1735 5478 -1734
rect 5436 -1769 5441 -1735
rect 5471 -1769 5478 -1735
rect 5436 -1778 5478 -1769
rect 5512 -1735 5554 -1726
rect 5512 -1769 5519 -1735
rect 5549 -1769 5554 -1735
rect 5512 -1774 5554 -1769
rect 5588 -1762 5616 -1702
tri 5661 -1715 5683 -1693 se
rect 5683 -1700 5698 -1692
tri 5683 -1715 5698 -1700 nw
tri 5655 -1721 5661 -1715 se
rect 5661 -1721 5670 -1715
rect 5374 -1806 5402 -1796
tri 5402 -1806 5426 -1782 sw
rect 5374 -1838 5416 -1806
tri 5433 -1814 5434 -1813 sw
rect 5433 -1838 5434 -1814
tri 5436 -1815 5473 -1778 ne
rect 5473 -1806 5478 -1778
tri 5478 -1806 5504 -1780 sw
rect 5588 -1796 5597 -1762
rect 5588 -1806 5616 -1796
rect 5473 -1815 5557 -1806
tri 5473 -1834 5492 -1815 ne
rect 5492 -1834 5557 -1815
rect 5374 -1860 5434 -1838
rect 5556 -1838 5557 -1834
rect 5574 -1838 5616 -1806
rect 5556 -1860 5616 -1838
rect 5462 -1876 5479 -1862
rect 5511 -1876 5528 -1862
tri 5299 -1912 5321 -1890 se
rect 5321 -1897 5336 -1876
tri 5321 -1912 5336 -1897 nw
rect 5655 -1897 5670 -1721
tri 5670 -1728 5683 -1715 nw
rect 5756 -1796 5771 -1568
tri 5293 -1918 5299 -1912 se
rect 5299 -1918 5308 -1912
rect 5293 -1934 5308 -1918
tri 5308 -1925 5321 -1912 nw
rect 5462 -1920 5479 -1906
rect 5511 -1920 5528 -1906
tri 5655 -1912 5670 -1897 ne
tri 5670 -1912 5692 -1890 sw
rect 5293 -1970 5308 -1962
rect 5374 -1934 5434 -1920
rect 5389 -1944 5434 -1934
rect 5389 -1962 5417 -1944
tri 5293 -1985 5308 -1970 ne
tri 5308 -1985 5330 -1963 sw
rect 5374 -1972 5417 -1962
rect 5432 -1948 5434 -1944
rect 5556 -1934 5616 -1920
tri 5670 -1925 5683 -1912 ne
rect 5683 -1918 5692 -1912
tri 5692 -1918 5698 -1912 sw
rect 5556 -1944 5601 -1934
rect 5432 -1972 5506 -1948
rect 5374 -1976 5506 -1972
tri 5506 -1976 5534 -1948 sw
rect 5556 -1958 5558 -1944
tri 5556 -1960 5558 -1958 ne
rect 5570 -1962 5601 -1944
rect 5570 -1972 5616 -1962
rect 5683 -1933 5698 -1918
tri 5308 -1997 5320 -1985 ne
rect 5320 -1990 5330 -1985
tri 5330 -1990 5335 -1985 sw
rect 5219 -2146 5234 -2108
rect 5320 -2146 5335 -1990
rect 5374 -2032 5402 -1976
tri 5494 -1994 5512 -1976 ne
rect 5512 -1996 5534 -1976
tri 5534 -1996 5554 -1976 sw
tri 5570 -1990 5588 -1972 ne
rect 5393 -2066 5402 -2032
rect 5436 -2005 5478 -2004
rect 5436 -2039 5441 -2005
rect 5471 -2039 5478 -2005
rect 5436 -2048 5478 -2039
rect 5512 -2005 5554 -1996
rect 5512 -2039 5519 -2005
rect 5549 -2039 5554 -2005
rect 5512 -2044 5554 -2039
rect 5588 -2032 5616 -1972
tri 5661 -1985 5683 -1963 se
rect 5683 -1970 5698 -1962
tri 5683 -1985 5698 -1970 nw
tri 5655 -1991 5661 -1985 se
rect 5661 -1991 5670 -1985
rect 5374 -2076 5402 -2066
tri 5402 -2076 5426 -2052 sw
rect 5374 -2108 5416 -2076
tri 5433 -2084 5434 -2083 sw
rect 5433 -2108 5434 -2084
tri 5436 -2085 5473 -2048 ne
rect 5473 -2076 5478 -2048
tri 5478 -2076 5504 -2050 sw
rect 5588 -2066 5597 -2032
rect 5588 -2076 5616 -2066
rect 5473 -2085 5557 -2076
tri 5473 -2104 5492 -2085 ne
rect 5492 -2104 5557 -2085
rect 5374 -2130 5434 -2108
rect 5556 -2108 5557 -2104
rect 5574 -2108 5616 -2076
rect 5556 -2130 5616 -2108
rect 5462 -2146 5479 -2132
rect 5511 -2146 5528 -2132
rect 5655 -2146 5670 -1991
tri 5670 -1998 5683 -1985 nw
rect 5756 -2066 5771 -1838
rect 5756 -2146 5771 -2108
rect 5799 1984 5814 2174
tri 5879 2138 5901 2160 se
rect 5901 2153 5916 2174
tri 5901 2138 5916 2153 nw
rect 6235 2153 6250 2174
tri 5873 2132 5879 2138 se
rect 5879 2132 5888 2138
rect 5873 2116 5888 2132
tri 5888 2125 5901 2138 nw
rect 6042 2130 6059 2144
rect 6091 2130 6108 2144
tri 6235 2138 6250 2153 ne
tri 6250 2138 6272 2160 sw
rect 5873 2080 5888 2088
rect 5954 2116 6014 2130
rect 5969 2106 6014 2116
rect 5969 2088 5997 2106
tri 5873 2065 5888 2080 ne
tri 5888 2065 5910 2087 sw
rect 5954 2078 5997 2088
rect 6012 2102 6014 2106
rect 6136 2116 6196 2130
tri 6250 2125 6263 2138 ne
rect 6263 2132 6272 2138
tri 6272 2132 6278 2138 sw
rect 6136 2106 6181 2116
rect 6012 2078 6086 2102
rect 5954 2074 6086 2078
tri 6086 2074 6114 2102 sw
rect 6136 2092 6138 2106
tri 6136 2090 6138 2092 ne
rect 6150 2088 6181 2106
rect 6150 2078 6196 2088
rect 6263 2117 6278 2132
tri 5888 2053 5900 2065 ne
rect 5900 2060 5910 2065
tri 5910 2060 5915 2065 sw
rect 5799 1714 5814 1942
rect 5900 1904 5915 2060
rect 5954 2018 5982 2074
tri 6074 2056 6092 2074 ne
rect 6092 2054 6114 2074
tri 6114 2054 6134 2074 sw
tri 6150 2060 6168 2078 ne
rect 5973 1984 5982 2018
rect 6016 2045 6058 2046
rect 6016 2011 6021 2045
rect 6051 2011 6058 2045
rect 6016 2002 6058 2011
rect 6092 2045 6134 2054
rect 6092 2011 6099 2045
rect 6129 2011 6134 2045
rect 6092 2006 6134 2011
rect 6168 2018 6196 2078
tri 6241 2065 6263 2087 se
rect 6263 2080 6278 2088
tri 6263 2065 6278 2080 nw
tri 6235 2059 6241 2065 se
rect 6241 2059 6250 2065
rect 5954 1974 5982 1984
tri 5982 1974 6006 1998 sw
rect 5954 1942 5996 1974
tri 6013 1966 6014 1967 sw
rect 6013 1942 6014 1966
tri 6016 1965 6053 2002 ne
rect 6053 1974 6058 2002
tri 6058 1974 6084 2000 sw
rect 6168 1984 6177 2018
rect 6168 1974 6196 1984
rect 6053 1965 6137 1974
tri 6053 1946 6072 1965 ne
rect 6072 1946 6137 1965
rect 5954 1920 6014 1942
rect 6136 1942 6137 1946
rect 6154 1942 6196 1974
rect 6136 1920 6196 1942
rect 6042 1904 6059 1918
rect 6091 1904 6108 1918
tri 5879 1868 5901 1890 se
rect 5901 1883 5916 1904
tri 5901 1868 5916 1883 nw
rect 6235 1883 6250 2059
tri 6250 2052 6263 2065 nw
rect 6336 1984 6351 2174
tri 5873 1862 5879 1868 se
rect 5879 1862 5888 1868
rect 5873 1846 5888 1862
tri 5888 1855 5901 1868 nw
rect 6042 1860 6059 1874
rect 6091 1860 6108 1874
tri 6235 1868 6250 1883 ne
tri 6250 1868 6272 1890 sw
rect 5873 1810 5888 1818
rect 5954 1846 6014 1860
rect 5969 1836 6014 1846
rect 5969 1818 5997 1836
tri 5873 1795 5888 1810 ne
tri 5888 1795 5910 1817 sw
rect 5954 1808 5997 1818
rect 6012 1832 6014 1836
rect 6136 1846 6196 1860
tri 6250 1855 6263 1868 ne
rect 6263 1862 6272 1868
tri 6272 1862 6278 1868 sw
rect 6136 1836 6181 1846
rect 6012 1808 6086 1832
rect 5954 1804 6086 1808
tri 6086 1804 6114 1832 sw
rect 6136 1822 6138 1836
tri 6136 1820 6138 1822 ne
rect 6150 1818 6181 1836
rect 6150 1808 6196 1818
rect 6263 1847 6278 1862
tri 5888 1783 5900 1795 ne
rect 5900 1790 5910 1795
tri 5910 1790 5915 1795 sw
rect 5799 1444 5814 1672
rect 5900 1682 5915 1790
rect 5954 1748 5982 1804
tri 6074 1786 6092 1804 ne
rect 6092 1784 6114 1804
tri 6114 1784 6134 1804 sw
tri 6150 1790 6168 1808 ne
rect 5973 1714 5982 1748
rect 6016 1775 6058 1776
rect 6016 1741 6021 1775
rect 6051 1741 6058 1775
rect 6016 1732 6058 1741
rect 6092 1775 6134 1784
rect 6092 1741 6099 1775
rect 6129 1741 6134 1775
rect 6092 1736 6134 1741
rect 6168 1748 6196 1808
tri 6241 1795 6263 1817 se
rect 6263 1810 6278 1818
tri 6263 1795 6278 1810 nw
tri 6235 1789 6241 1795 se
rect 6241 1789 6250 1795
rect 5954 1704 5982 1714
tri 5982 1704 6006 1728 sw
rect 5900 1634 5916 1682
rect 5954 1672 5996 1704
tri 6013 1696 6014 1697 sw
rect 6013 1672 6014 1696
tri 6016 1695 6053 1732 ne
rect 6053 1704 6058 1732
tri 6058 1704 6084 1730 sw
rect 6168 1714 6177 1748
rect 6168 1704 6196 1714
rect 6053 1695 6137 1704
tri 6053 1676 6072 1695 ne
rect 6072 1676 6137 1695
rect 5954 1650 6014 1672
rect 6136 1672 6137 1676
rect 6154 1672 6196 1704
rect 6136 1650 6196 1672
rect 6042 1634 6059 1648
rect 6091 1634 6108 1648
tri 5879 1598 5901 1620 se
rect 5901 1613 5916 1634
tri 5901 1598 5916 1613 nw
rect 6235 1613 6250 1789
tri 6250 1782 6263 1795 nw
rect 6336 1714 6351 1942
tri 5873 1592 5879 1598 se
rect 5879 1592 5888 1598
rect 5873 1576 5888 1592
tri 5888 1585 5901 1598 nw
rect 6042 1590 6059 1604
rect 6091 1590 6108 1604
tri 6235 1598 6250 1613 ne
tri 6250 1598 6272 1620 sw
rect 5873 1540 5888 1548
rect 5954 1576 6014 1590
rect 5969 1566 6014 1576
rect 5969 1548 5997 1566
tri 5873 1525 5888 1540 ne
tri 5888 1525 5910 1547 sw
rect 5954 1538 5997 1548
rect 6012 1562 6014 1566
rect 6136 1576 6196 1590
tri 6250 1585 6263 1598 ne
rect 6263 1592 6272 1598
tri 6272 1592 6278 1598 sw
rect 6136 1566 6181 1576
rect 6012 1538 6086 1562
rect 5954 1534 6086 1538
tri 6086 1534 6114 1562 sw
rect 6136 1552 6138 1566
tri 6136 1550 6138 1552 ne
rect 6150 1548 6181 1566
rect 6150 1538 6196 1548
rect 6263 1577 6278 1592
tri 5888 1513 5900 1525 ne
rect 5900 1520 5910 1525
tri 5910 1520 5915 1525 sw
rect 5799 1174 5814 1402
rect 5900 1364 5915 1520
rect 5954 1478 5982 1534
tri 6074 1516 6092 1534 ne
rect 6092 1514 6114 1534
tri 6114 1514 6134 1534 sw
tri 6150 1520 6168 1538 ne
rect 5973 1444 5982 1478
rect 6016 1505 6058 1506
rect 6016 1471 6021 1505
rect 6051 1471 6058 1505
rect 6016 1462 6058 1471
rect 6092 1505 6134 1514
rect 6092 1471 6099 1505
rect 6129 1471 6134 1505
rect 6092 1466 6134 1471
rect 6168 1478 6196 1538
tri 6241 1525 6263 1547 se
rect 6263 1540 6278 1548
tri 6263 1525 6278 1540 nw
tri 6235 1519 6241 1525 se
rect 6241 1519 6250 1525
rect 5954 1434 5982 1444
tri 5982 1434 6006 1458 sw
rect 5954 1402 5996 1434
tri 6013 1426 6014 1427 sw
rect 6013 1402 6014 1426
tri 6016 1425 6053 1462 ne
rect 6053 1434 6058 1462
tri 6058 1434 6084 1460 sw
rect 6168 1444 6177 1478
rect 6168 1434 6196 1444
rect 6053 1425 6137 1434
tri 6053 1406 6072 1425 ne
rect 6072 1406 6137 1425
rect 5954 1380 6014 1402
rect 6136 1402 6137 1406
rect 6154 1402 6196 1434
rect 6136 1380 6196 1402
rect 6042 1364 6059 1378
rect 6091 1364 6108 1378
tri 5879 1328 5901 1350 se
rect 5901 1343 5916 1364
tri 5901 1328 5916 1343 nw
rect 6235 1343 6250 1519
tri 6250 1512 6263 1525 nw
rect 6336 1444 6351 1672
tri 5873 1322 5879 1328 se
rect 5879 1322 5888 1328
rect 5873 1306 5888 1322
tri 5888 1315 5901 1328 nw
rect 6042 1320 6059 1334
rect 6091 1320 6108 1334
tri 6235 1328 6250 1343 ne
tri 6250 1328 6272 1350 sw
rect 5873 1270 5888 1278
rect 5954 1306 6014 1320
rect 5969 1296 6014 1306
rect 5969 1278 5997 1296
tri 5873 1255 5888 1270 ne
tri 5888 1255 5910 1277 sw
rect 5954 1268 5997 1278
rect 6012 1292 6014 1296
rect 6136 1306 6196 1320
tri 6250 1315 6263 1328 ne
rect 6263 1322 6272 1328
tri 6272 1322 6278 1328 sw
rect 6136 1296 6181 1306
rect 6012 1268 6086 1292
rect 5954 1264 6086 1268
tri 6086 1264 6114 1292 sw
rect 6136 1282 6138 1296
tri 6136 1280 6138 1282 ne
rect 6150 1278 6181 1296
rect 6150 1268 6196 1278
rect 6263 1307 6278 1322
tri 5888 1243 5900 1255 ne
rect 5900 1250 5910 1255
tri 5910 1250 5915 1255 sw
rect 5799 904 5814 1132
rect 5900 1142 5915 1250
rect 5954 1208 5982 1264
tri 6074 1246 6092 1264 ne
rect 6092 1244 6114 1264
tri 6114 1244 6134 1264 sw
tri 6150 1250 6168 1268 ne
rect 5973 1174 5982 1208
rect 6016 1235 6058 1236
rect 6016 1201 6021 1235
rect 6051 1201 6058 1235
rect 6016 1192 6058 1201
rect 6092 1235 6134 1244
rect 6092 1201 6099 1235
rect 6129 1201 6134 1235
rect 6092 1196 6134 1201
rect 6168 1208 6196 1268
tri 6241 1255 6263 1277 se
rect 6263 1270 6278 1278
tri 6263 1255 6278 1270 nw
tri 6235 1249 6241 1255 se
rect 6241 1249 6250 1255
rect 5954 1164 5982 1174
tri 5982 1164 6006 1188 sw
rect 5900 1094 5916 1142
rect 5954 1132 5996 1164
tri 6013 1156 6014 1157 sw
rect 6013 1132 6014 1156
tri 6016 1155 6053 1192 ne
rect 6053 1164 6058 1192
tri 6058 1164 6084 1190 sw
rect 6168 1174 6177 1208
rect 6168 1164 6196 1174
rect 6053 1155 6137 1164
tri 6053 1136 6072 1155 ne
rect 6072 1136 6137 1155
rect 5954 1110 6014 1132
rect 6136 1132 6137 1136
rect 6154 1132 6196 1164
rect 6136 1110 6196 1132
rect 6042 1094 6059 1108
rect 6091 1094 6108 1108
tri 5879 1058 5901 1080 se
rect 5901 1073 5916 1094
tri 5901 1058 5916 1073 nw
rect 6235 1073 6250 1249
tri 6250 1242 6263 1255 nw
rect 6336 1174 6351 1402
tri 5873 1052 5879 1058 se
rect 5879 1052 5888 1058
rect 5873 1036 5888 1052
tri 5888 1045 5901 1058 nw
rect 6042 1050 6059 1064
rect 6091 1050 6108 1064
tri 6235 1058 6250 1073 ne
tri 6250 1058 6272 1080 sw
rect 5873 1000 5888 1008
rect 5954 1036 6014 1050
rect 5969 1026 6014 1036
rect 5969 1008 5997 1026
tri 5873 985 5888 1000 ne
tri 5888 985 5910 1007 sw
rect 5954 998 5997 1008
rect 6012 1022 6014 1026
rect 6136 1036 6196 1050
tri 6250 1045 6263 1058 ne
rect 6263 1052 6272 1058
tri 6272 1052 6278 1058 sw
rect 6136 1026 6181 1036
rect 6012 998 6086 1022
rect 5954 994 6086 998
tri 6086 994 6114 1022 sw
rect 6136 1012 6138 1026
tri 6136 1010 6138 1012 ne
rect 6150 1008 6181 1026
rect 6150 998 6196 1008
rect 6263 1037 6278 1052
tri 5888 973 5900 985 ne
rect 5900 980 5910 985
tri 5910 980 5915 985 sw
rect 5799 634 5814 862
rect 5900 824 5915 980
rect 5954 938 5982 994
tri 6074 976 6092 994 ne
rect 6092 974 6114 994
tri 6114 974 6134 994 sw
tri 6150 980 6168 998 ne
rect 5973 904 5982 938
rect 6016 965 6058 966
rect 6016 931 6021 965
rect 6051 931 6058 965
rect 6016 922 6058 931
rect 6092 965 6134 974
rect 6092 931 6099 965
rect 6129 931 6134 965
rect 6092 926 6134 931
rect 6168 938 6196 998
tri 6241 985 6263 1007 se
rect 6263 1000 6278 1008
tri 6263 985 6278 1000 nw
tri 6235 979 6241 985 se
rect 6241 979 6250 985
rect 5954 894 5982 904
tri 5982 894 6006 918 sw
rect 5954 862 5996 894
tri 6013 886 6014 887 sw
rect 6013 862 6014 886
tri 6016 885 6053 922 ne
rect 6053 894 6058 922
tri 6058 894 6084 920 sw
rect 6168 904 6177 938
rect 6168 894 6196 904
rect 6053 885 6137 894
tri 6053 866 6072 885 ne
rect 6072 866 6137 885
rect 5954 840 6014 862
rect 6136 862 6137 866
rect 6154 862 6196 894
rect 6136 840 6196 862
rect 6042 824 6059 838
rect 6091 824 6108 838
tri 5879 788 5901 810 se
rect 5901 803 5916 824
tri 5901 788 5916 803 nw
rect 6235 803 6250 979
tri 6250 972 6263 985 nw
rect 6336 904 6351 1132
tri 5873 782 5879 788 se
rect 5879 782 5888 788
rect 5873 766 5888 782
tri 5888 775 5901 788 nw
rect 6042 780 6059 794
rect 6091 780 6108 794
tri 6235 788 6250 803 ne
tri 6250 788 6272 810 sw
rect 5873 730 5888 738
rect 5954 766 6014 780
rect 5969 756 6014 766
rect 5969 738 5997 756
tri 5873 715 5888 730 ne
tri 5888 715 5910 737 sw
rect 5954 728 5997 738
rect 6012 752 6014 756
rect 6136 766 6196 780
tri 6250 775 6263 788 ne
rect 6263 782 6272 788
tri 6272 782 6278 788 sw
rect 6136 756 6181 766
rect 6012 728 6086 752
rect 5954 724 6086 728
tri 6086 724 6114 752 sw
rect 6136 742 6138 756
tri 6136 740 6138 742 ne
rect 6150 738 6181 756
rect 6150 728 6196 738
rect 6263 767 6278 782
tri 5888 703 5900 715 ne
rect 5900 710 5910 715
tri 5910 710 5915 715 sw
rect 5799 364 5814 592
rect 5900 602 5915 710
rect 5954 668 5982 724
tri 6074 706 6092 724 ne
rect 6092 704 6114 724
tri 6114 704 6134 724 sw
tri 6150 710 6168 728 ne
rect 5973 634 5982 668
rect 6016 695 6058 696
rect 6016 661 6021 695
rect 6051 661 6058 695
rect 6016 652 6058 661
rect 6092 695 6134 704
rect 6092 661 6099 695
rect 6129 661 6134 695
rect 6092 656 6134 661
rect 6168 668 6196 728
tri 6241 715 6263 737 se
rect 6263 730 6278 738
tri 6263 715 6278 730 nw
tri 6235 709 6241 715 se
rect 6241 709 6250 715
rect 5954 624 5982 634
tri 5982 624 6006 648 sw
rect 5900 554 5916 602
rect 5954 592 5996 624
tri 6013 616 6014 617 sw
rect 6013 592 6014 616
tri 6016 615 6053 652 ne
rect 6053 624 6058 652
tri 6058 624 6084 650 sw
rect 6168 634 6177 668
rect 6168 624 6196 634
rect 6053 615 6137 624
tri 6053 596 6072 615 ne
rect 6072 596 6137 615
rect 5954 570 6014 592
rect 6136 592 6137 596
rect 6154 592 6196 624
rect 6136 570 6196 592
rect 6042 554 6059 568
rect 6091 554 6108 568
tri 5879 518 5901 540 se
rect 5901 533 5916 554
tri 5901 518 5916 533 nw
rect 6235 533 6250 709
tri 6250 702 6263 715 nw
rect 6336 634 6351 862
tri 5873 512 5879 518 se
rect 5879 512 5888 518
rect 5873 496 5888 512
tri 5888 505 5901 518 nw
rect 6042 510 6059 524
rect 6091 510 6108 524
tri 6235 518 6250 533 ne
tri 6250 518 6272 540 sw
rect 5873 460 5888 468
rect 5954 496 6014 510
rect 5969 486 6014 496
rect 5969 468 5997 486
tri 5873 445 5888 460 ne
tri 5888 445 5910 467 sw
rect 5954 458 5997 468
rect 6012 482 6014 486
rect 6136 496 6196 510
tri 6250 505 6263 518 ne
rect 6263 512 6272 518
tri 6272 512 6278 518 sw
rect 6136 486 6181 496
rect 6012 458 6086 482
rect 5954 454 6086 458
tri 6086 454 6114 482 sw
rect 6136 472 6138 486
tri 6136 470 6138 472 ne
rect 6150 468 6181 486
rect 6150 458 6196 468
rect 6263 497 6278 512
tri 5888 433 5900 445 ne
rect 5900 440 5910 445
tri 5910 440 5915 445 sw
rect 5799 94 5814 322
rect 5900 284 5915 440
rect 5954 398 5982 454
tri 6074 436 6092 454 ne
rect 6092 434 6114 454
tri 6114 434 6134 454 sw
tri 6150 440 6168 458 ne
rect 5973 364 5982 398
rect 6016 425 6058 426
rect 6016 391 6021 425
rect 6051 391 6058 425
rect 6016 382 6058 391
rect 6092 425 6134 434
rect 6092 391 6099 425
rect 6129 391 6134 425
rect 6092 386 6134 391
rect 6168 398 6196 458
tri 6241 445 6263 467 se
rect 6263 460 6278 468
tri 6263 445 6278 460 nw
tri 6235 439 6241 445 se
rect 6241 439 6250 445
rect 5954 354 5982 364
tri 5982 354 6006 378 sw
rect 5954 322 5996 354
tri 6013 346 6014 347 sw
rect 6013 322 6014 346
tri 6016 345 6053 382 ne
rect 6053 354 6058 382
tri 6058 354 6084 380 sw
rect 6168 364 6177 398
rect 6168 354 6196 364
rect 6053 345 6137 354
tri 6053 326 6072 345 ne
rect 6072 326 6137 345
rect 5954 300 6014 322
rect 6136 322 6137 326
rect 6154 322 6196 354
rect 6136 300 6196 322
rect 6042 284 6059 298
rect 6091 284 6108 298
tri 5879 248 5901 270 se
rect 5901 263 5916 284
tri 5901 248 5916 263 nw
rect 6235 263 6250 439
tri 6250 432 6263 445 nw
rect 6336 364 6351 592
tri 5873 242 5879 248 se
rect 5879 242 5888 248
rect 5873 226 5888 242
tri 5888 235 5901 248 nw
rect 6042 240 6059 254
rect 6091 240 6108 254
tri 6235 248 6250 263 ne
tri 6250 248 6272 270 sw
rect 5873 190 5888 198
rect 5954 226 6014 240
rect 5969 216 6014 226
rect 5969 198 5997 216
tri 5873 175 5888 190 ne
tri 5888 175 5910 197 sw
rect 5954 188 5997 198
rect 6012 212 6014 216
rect 6136 226 6196 240
tri 6250 235 6263 248 ne
rect 6263 242 6272 248
tri 6272 242 6278 248 sw
rect 6136 216 6181 226
rect 6012 188 6086 212
rect 5954 184 6086 188
tri 6086 184 6114 212 sw
rect 6136 202 6138 216
tri 6136 200 6138 202 ne
rect 6150 198 6181 216
rect 6150 188 6196 198
rect 6263 227 6278 242
tri 5888 163 5900 175 ne
rect 5900 170 5910 175
tri 5910 170 5915 175 sw
rect 5799 -176 5814 52
rect 5900 62 5915 170
rect 5954 128 5982 184
tri 6074 166 6092 184 ne
rect 6092 164 6114 184
tri 6114 164 6134 184 sw
tri 6150 170 6168 188 ne
rect 5973 94 5982 128
rect 6016 155 6058 156
rect 6016 121 6021 155
rect 6051 121 6058 155
rect 6016 112 6058 121
rect 6092 155 6134 164
rect 6092 121 6099 155
rect 6129 121 6134 155
rect 6092 116 6134 121
rect 6168 128 6196 188
tri 6241 175 6263 197 se
rect 6263 190 6278 198
tri 6263 175 6278 190 nw
tri 6235 169 6241 175 se
rect 6241 169 6250 175
rect 5954 84 5982 94
tri 5982 84 6006 108 sw
rect 5900 14 5916 62
rect 5954 52 5996 84
tri 6013 76 6014 77 sw
rect 6013 52 6014 76
tri 6016 75 6053 112 ne
rect 6053 84 6058 112
tri 6058 84 6084 110 sw
rect 6168 94 6177 128
rect 6168 84 6196 94
rect 6053 75 6137 84
tri 6053 56 6072 75 ne
rect 6072 56 6137 75
rect 5954 30 6014 52
rect 6136 52 6137 56
rect 6154 52 6196 84
rect 6136 30 6196 52
rect 6042 14 6059 28
rect 6091 14 6108 28
tri 5879 -22 5901 0 se
rect 5901 -7 5916 14
tri 5901 -22 5916 -7 nw
rect 6235 -7 6250 169
tri 6250 162 6263 175 nw
rect 6336 94 6351 322
tri 5873 -28 5879 -22 se
rect 5879 -28 5888 -22
rect 5873 -44 5888 -28
tri 5888 -35 5901 -22 nw
rect 6042 -30 6059 -16
rect 6091 -30 6108 -16
tri 6235 -22 6250 -7 ne
tri 6250 -22 6272 0 sw
rect 5873 -80 5888 -72
rect 5954 -44 6014 -30
rect 5969 -54 6014 -44
rect 5969 -72 5997 -54
tri 5873 -95 5888 -80 ne
tri 5888 -95 5910 -73 sw
rect 5954 -82 5997 -72
rect 6012 -58 6014 -54
rect 6136 -44 6196 -30
tri 6250 -35 6263 -22 ne
rect 6263 -28 6272 -22
tri 6272 -28 6278 -22 sw
rect 6136 -54 6181 -44
rect 6012 -82 6086 -58
rect 5954 -86 6086 -82
tri 6086 -86 6114 -58 sw
rect 6136 -68 6138 -54
tri 6136 -70 6138 -68 ne
rect 6150 -72 6181 -54
rect 6150 -82 6196 -72
rect 6263 -43 6278 -28
tri 5888 -107 5900 -95 ne
rect 5900 -100 5910 -95
tri 5910 -100 5915 -95 sw
rect 5799 -446 5814 -218
rect 5900 -256 5915 -100
rect 5954 -142 5982 -86
tri 6074 -104 6092 -86 ne
rect 6092 -106 6114 -86
tri 6114 -106 6134 -86 sw
tri 6150 -100 6168 -82 ne
rect 5973 -176 5982 -142
rect 6016 -115 6058 -114
rect 6016 -149 6021 -115
rect 6051 -149 6058 -115
rect 6016 -158 6058 -149
rect 6092 -115 6134 -106
rect 6092 -149 6099 -115
rect 6129 -149 6134 -115
rect 6092 -154 6134 -149
rect 6168 -142 6196 -82
tri 6241 -95 6263 -73 se
rect 6263 -80 6278 -72
tri 6263 -95 6278 -80 nw
tri 6235 -101 6241 -95 se
rect 6241 -101 6250 -95
rect 5954 -186 5982 -176
tri 5982 -186 6006 -162 sw
rect 5954 -218 5996 -186
tri 6013 -194 6014 -193 sw
rect 6013 -218 6014 -194
tri 6016 -195 6053 -158 ne
rect 6053 -186 6058 -158
tri 6058 -186 6084 -160 sw
rect 6168 -176 6177 -142
rect 6168 -186 6196 -176
rect 6053 -195 6137 -186
tri 6053 -214 6072 -195 ne
rect 6072 -214 6137 -195
rect 5954 -240 6014 -218
rect 6136 -218 6137 -214
rect 6154 -218 6196 -186
rect 6136 -240 6196 -218
rect 6042 -256 6059 -242
rect 6091 -256 6108 -242
tri 5879 -292 5901 -270 se
rect 5901 -277 5916 -256
tri 5901 -292 5916 -277 nw
rect 6235 -277 6250 -101
tri 6250 -108 6263 -95 nw
rect 6336 -176 6351 52
tri 5873 -298 5879 -292 se
rect 5879 -298 5888 -292
rect 5873 -314 5888 -298
tri 5888 -305 5901 -292 nw
rect 6042 -300 6059 -286
rect 6091 -300 6108 -286
tri 6235 -292 6250 -277 ne
tri 6250 -292 6272 -270 sw
rect 5873 -350 5888 -342
rect 5954 -314 6014 -300
rect 5969 -324 6014 -314
rect 5969 -342 5997 -324
tri 5873 -365 5888 -350 ne
tri 5888 -365 5910 -343 sw
rect 5954 -352 5997 -342
rect 6012 -328 6014 -324
rect 6136 -314 6196 -300
tri 6250 -305 6263 -292 ne
rect 6263 -298 6272 -292
tri 6272 -298 6278 -292 sw
rect 6136 -324 6181 -314
rect 6012 -352 6086 -328
rect 5954 -356 6086 -352
tri 6086 -356 6114 -328 sw
rect 6136 -338 6138 -324
tri 6136 -340 6138 -338 ne
rect 6150 -342 6181 -324
rect 6150 -352 6196 -342
rect 6263 -313 6278 -298
tri 5888 -377 5900 -365 ne
rect 5900 -370 5910 -365
tri 5910 -370 5915 -365 sw
rect 5799 -716 5814 -488
rect 5900 -478 5915 -370
rect 5954 -412 5982 -356
tri 6074 -374 6092 -356 ne
rect 6092 -376 6114 -356
tri 6114 -376 6134 -356 sw
tri 6150 -370 6168 -352 ne
rect 5973 -446 5982 -412
rect 6016 -385 6058 -384
rect 6016 -419 6021 -385
rect 6051 -419 6058 -385
rect 6016 -428 6058 -419
rect 6092 -385 6134 -376
rect 6092 -419 6099 -385
rect 6129 -419 6134 -385
rect 6092 -424 6134 -419
rect 6168 -412 6196 -352
tri 6241 -365 6263 -343 se
rect 6263 -350 6278 -342
tri 6263 -365 6278 -350 nw
tri 6235 -371 6241 -365 se
rect 6241 -371 6250 -365
rect 5954 -456 5982 -446
tri 5982 -456 6006 -432 sw
rect 5900 -526 5916 -478
rect 5954 -488 5996 -456
tri 6013 -464 6014 -463 sw
rect 6013 -488 6014 -464
tri 6016 -465 6053 -428 ne
rect 6053 -456 6058 -428
tri 6058 -456 6084 -430 sw
rect 6168 -446 6177 -412
rect 6168 -456 6196 -446
rect 6053 -465 6137 -456
tri 6053 -484 6072 -465 ne
rect 6072 -484 6137 -465
rect 5954 -510 6014 -488
rect 6136 -488 6137 -484
rect 6154 -488 6196 -456
rect 6136 -510 6196 -488
rect 6042 -526 6059 -512
rect 6091 -526 6108 -512
tri 5879 -562 5901 -540 se
rect 5901 -547 5916 -526
tri 5901 -562 5916 -547 nw
rect 6235 -547 6250 -371
tri 6250 -378 6263 -365 nw
rect 6336 -446 6351 -218
tri 5873 -568 5879 -562 se
rect 5879 -568 5888 -562
rect 5873 -584 5888 -568
tri 5888 -575 5901 -562 nw
rect 6042 -570 6059 -556
rect 6091 -570 6108 -556
tri 6235 -562 6250 -547 ne
tri 6250 -562 6272 -540 sw
rect 5873 -620 5888 -612
rect 5954 -584 6014 -570
rect 5969 -594 6014 -584
rect 5969 -612 5997 -594
tri 5873 -635 5888 -620 ne
tri 5888 -635 5910 -613 sw
rect 5954 -622 5997 -612
rect 6012 -598 6014 -594
rect 6136 -584 6196 -570
tri 6250 -575 6263 -562 ne
rect 6263 -568 6272 -562
tri 6272 -568 6278 -562 sw
rect 6136 -594 6181 -584
rect 6012 -622 6086 -598
rect 5954 -626 6086 -622
tri 6086 -626 6114 -598 sw
rect 6136 -608 6138 -594
tri 6136 -610 6138 -608 ne
rect 6150 -612 6181 -594
rect 6150 -622 6196 -612
rect 6263 -583 6278 -568
tri 5888 -647 5900 -635 ne
rect 5900 -640 5910 -635
tri 5910 -640 5915 -635 sw
rect 5799 -986 5814 -758
rect 5900 -796 5915 -640
rect 5954 -682 5982 -626
tri 6074 -644 6092 -626 ne
rect 6092 -646 6114 -626
tri 6114 -646 6134 -626 sw
tri 6150 -640 6168 -622 ne
rect 5973 -716 5982 -682
rect 6016 -655 6058 -654
rect 6016 -689 6021 -655
rect 6051 -689 6058 -655
rect 6016 -698 6058 -689
rect 6092 -655 6134 -646
rect 6092 -689 6099 -655
rect 6129 -689 6134 -655
rect 6092 -694 6134 -689
rect 6168 -682 6196 -622
tri 6241 -635 6263 -613 se
rect 6263 -620 6278 -612
tri 6263 -635 6278 -620 nw
tri 6235 -641 6241 -635 se
rect 6241 -641 6250 -635
rect 5954 -726 5982 -716
tri 5982 -726 6006 -702 sw
rect 5954 -758 5996 -726
tri 6013 -734 6014 -733 sw
rect 6013 -758 6014 -734
tri 6016 -735 6053 -698 ne
rect 6053 -726 6058 -698
tri 6058 -726 6084 -700 sw
rect 6168 -716 6177 -682
rect 6168 -726 6196 -716
rect 6053 -735 6137 -726
tri 6053 -754 6072 -735 ne
rect 6072 -754 6137 -735
rect 5954 -780 6014 -758
rect 6136 -758 6137 -754
rect 6154 -758 6196 -726
rect 6136 -780 6196 -758
rect 6042 -796 6059 -782
rect 6091 -796 6108 -782
tri 5879 -832 5901 -810 se
rect 5901 -817 5916 -796
tri 5901 -832 5916 -817 nw
rect 6235 -817 6250 -641
tri 6250 -648 6263 -635 nw
rect 6336 -716 6351 -488
tri 5873 -838 5879 -832 se
rect 5879 -838 5888 -832
rect 5873 -854 5888 -838
tri 5888 -845 5901 -832 nw
rect 6042 -840 6059 -826
rect 6091 -840 6108 -826
tri 6235 -832 6250 -817 ne
tri 6250 -832 6272 -810 sw
rect 5873 -890 5888 -882
rect 5954 -854 6014 -840
rect 5969 -864 6014 -854
rect 5969 -882 5997 -864
tri 5873 -905 5888 -890 ne
tri 5888 -905 5910 -883 sw
rect 5954 -892 5997 -882
rect 6012 -868 6014 -864
rect 6136 -854 6196 -840
tri 6250 -845 6263 -832 ne
rect 6263 -838 6272 -832
tri 6272 -838 6278 -832 sw
rect 6136 -864 6181 -854
rect 6012 -892 6086 -868
rect 5954 -896 6086 -892
tri 6086 -896 6114 -868 sw
rect 6136 -878 6138 -864
tri 6136 -880 6138 -878 ne
rect 6150 -882 6181 -864
rect 6150 -892 6196 -882
rect 6263 -853 6278 -838
tri 5888 -917 5900 -905 ne
rect 5900 -910 5910 -905
tri 5910 -910 5915 -905 sw
rect 5799 -1256 5814 -1028
rect 5900 -1018 5915 -910
rect 5954 -952 5982 -896
tri 6074 -914 6092 -896 ne
rect 6092 -916 6114 -896
tri 6114 -916 6134 -896 sw
tri 6150 -910 6168 -892 ne
rect 5973 -986 5982 -952
rect 6016 -925 6058 -924
rect 6016 -959 6021 -925
rect 6051 -959 6058 -925
rect 6016 -968 6058 -959
rect 6092 -925 6134 -916
rect 6092 -959 6099 -925
rect 6129 -959 6134 -925
rect 6092 -964 6134 -959
rect 6168 -952 6196 -892
tri 6241 -905 6263 -883 se
rect 6263 -890 6278 -882
tri 6263 -905 6278 -890 nw
tri 6235 -911 6241 -905 se
rect 6241 -911 6250 -905
rect 5954 -996 5982 -986
tri 5982 -996 6006 -972 sw
rect 5900 -1066 5916 -1018
rect 5954 -1028 5996 -996
tri 6013 -1004 6014 -1003 sw
rect 6013 -1028 6014 -1004
tri 6016 -1005 6053 -968 ne
rect 6053 -996 6058 -968
tri 6058 -996 6084 -970 sw
rect 6168 -986 6177 -952
rect 6168 -996 6196 -986
rect 6053 -1005 6137 -996
tri 6053 -1024 6072 -1005 ne
rect 6072 -1024 6137 -1005
rect 5954 -1050 6014 -1028
rect 6136 -1028 6137 -1024
rect 6154 -1028 6196 -996
rect 6136 -1050 6196 -1028
rect 6042 -1066 6059 -1052
rect 6091 -1066 6108 -1052
tri 5879 -1102 5901 -1080 se
rect 5901 -1087 5916 -1066
tri 5901 -1102 5916 -1087 nw
rect 6235 -1087 6250 -911
tri 6250 -918 6263 -905 nw
rect 6336 -986 6351 -758
tri 5873 -1108 5879 -1102 se
rect 5879 -1108 5888 -1102
rect 5873 -1124 5888 -1108
tri 5888 -1115 5901 -1102 nw
rect 6042 -1110 6059 -1096
rect 6091 -1110 6108 -1096
tri 6235 -1102 6250 -1087 ne
tri 6250 -1102 6272 -1080 sw
rect 5873 -1160 5888 -1152
rect 5954 -1124 6014 -1110
rect 5969 -1134 6014 -1124
rect 5969 -1152 5997 -1134
tri 5873 -1175 5888 -1160 ne
tri 5888 -1175 5910 -1153 sw
rect 5954 -1162 5997 -1152
rect 6012 -1138 6014 -1134
rect 6136 -1124 6196 -1110
tri 6250 -1115 6263 -1102 ne
rect 6263 -1108 6272 -1102
tri 6272 -1108 6278 -1102 sw
rect 6136 -1134 6181 -1124
rect 6012 -1162 6086 -1138
rect 5954 -1166 6086 -1162
tri 6086 -1166 6114 -1138 sw
rect 6136 -1148 6138 -1134
tri 6136 -1150 6138 -1148 ne
rect 6150 -1152 6181 -1134
rect 6150 -1162 6196 -1152
rect 6263 -1123 6278 -1108
tri 5888 -1187 5900 -1175 ne
rect 5900 -1180 5910 -1175
tri 5910 -1180 5915 -1175 sw
rect 5799 -1526 5814 -1298
rect 5900 -1336 5915 -1180
rect 5954 -1222 5982 -1166
tri 6074 -1184 6092 -1166 ne
rect 6092 -1186 6114 -1166
tri 6114 -1186 6134 -1166 sw
tri 6150 -1180 6168 -1162 ne
rect 5973 -1256 5982 -1222
rect 6016 -1195 6058 -1194
rect 6016 -1229 6021 -1195
rect 6051 -1229 6058 -1195
rect 6016 -1238 6058 -1229
rect 6092 -1195 6134 -1186
rect 6092 -1229 6099 -1195
rect 6129 -1229 6134 -1195
rect 6092 -1234 6134 -1229
rect 6168 -1222 6196 -1162
tri 6241 -1175 6263 -1153 se
rect 6263 -1160 6278 -1152
tri 6263 -1175 6278 -1160 nw
tri 6235 -1181 6241 -1175 se
rect 6241 -1181 6250 -1175
rect 5954 -1266 5982 -1256
tri 5982 -1266 6006 -1242 sw
rect 5954 -1298 5996 -1266
tri 6013 -1274 6014 -1273 sw
rect 6013 -1298 6014 -1274
tri 6016 -1275 6053 -1238 ne
rect 6053 -1266 6058 -1238
tri 6058 -1266 6084 -1240 sw
rect 6168 -1256 6177 -1222
rect 6168 -1266 6196 -1256
rect 6053 -1275 6137 -1266
tri 6053 -1294 6072 -1275 ne
rect 6072 -1294 6137 -1275
rect 5954 -1320 6014 -1298
rect 6136 -1298 6137 -1294
rect 6154 -1298 6196 -1266
rect 6136 -1320 6196 -1298
rect 6042 -1336 6059 -1322
rect 6091 -1336 6108 -1322
tri 5879 -1372 5901 -1350 se
rect 5901 -1357 5916 -1336
tri 5901 -1372 5916 -1357 nw
rect 6235 -1357 6250 -1181
tri 6250 -1188 6263 -1175 nw
rect 6336 -1256 6351 -1028
tri 5873 -1378 5879 -1372 se
rect 5879 -1378 5888 -1372
rect 5873 -1394 5888 -1378
tri 5888 -1385 5901 -1372 nw
rect 6042 -1380 6059 -1366
rect 6091 -1380 6108 -1366
tri 6235 -1372 6250 -1357 ne
tri 6250 -1372 6272 -1350 sw
rect 5873 -1430 5888 -1422
rect 5954 -1394 6014 -1380
rect 5969 -1404 6014 -1394
rect 5969 -1422 5997 -1404
tri 5873 -1445 5888 -1430 ne
tri 5888 -1445 5910 -1423 sw
rect 5954 -1432 5997 -1422
rect 6012 -1408 6014 -1404
rect 6136 -1394 6196 -1380
tri 6250 -1385 6263 -1372 ne
rect 6263 -1378 6272 -1372
tri 6272 -1378 6278 -1372 sw
rect 6136 -1404 6181 -1394
rect 6012 -1432 6086 -1408
rect 5954 -1436 6086 -1432
tri 6086 -1436 6114 -1408 sw
rect 6136 -1418 6138 -1404
tri 6136 -1420 6138 -1418 ne
rect 6150 -1422 6181 -1404
rect 6150 -1432 6196 -1422
rect 6263 -1393 6278 -1378
tri 5888 -1457 5900 -1445 ne
rect 5900 -1450 5910 -1445
tri 5910 -1450 5915 -1445 sw
rect 5799 -1796 5814 -1568
rect 5900 -1558 5915 -1450
rect 5954 -1492 5982 -1436
tri 6074 -1454 6092 -1436 ne
rect 6092 -1456 6114 -1436
tri 6114 -1456 6134 -1436 sw
tri 6150 -1450 6168 -1432 ne
rect 5973 -1526 5982 -1492
rect 6016 -1465 6058 -1464
rect 6016 -1499 6021 -1465
rect 6051 -1499 6058 -1465
rect 6016 -1508 6058 -1499
rect 6092 -1465 6134 -1456
rect 6092 -1499 6099 -1465
rect 6129 -1499 6134 -1465
rect 6092 -1504 6134 -1499
rect 6168 -1492 6196 -1432
tri 6241 -1445 6263 -1423 se
rect 6263 -1430 6278 -1422
tri 6263 -1445 6278 -1430 nw
tri 6235 -1451 6241 -1445 se
rect 6241 -1451 6250 -1445
rect 5954 -1536 5982 -1526
tri 5982 -1536 6006 -1512 sw
rect 5900 -1606 5916 -1558
rect 5954 -1568 5996 -1536
tri 6013 -1544 6014 -1543 sw
rect 6013 -1568 6014 -1544
tri 6016 -1545 6053 -1508 ne
rect 6053 -1536 6058 -1508
tri 6058 -1536 6084 -1510 sw
rect 6168 -1526 6177 -1492
rect 6168 -1536 6196 -1526
rect 6053 -1545 6137 -1536
tri 6053 -1564 6072 -1545 ne
rect 6072 -1564 6137 -1545
rect 5954 -1590 6014 -1568
rect 6136 -1568 6137 -1564
rect 6154 -1568 6196 -1536
rect 6136 -1590 6196 -1568
rect 6042 -1606 6059 -1592
rect 6091 -1606 6108 -1592
tri 5879 -1642 5901 -1620 se
rect 5901 -1627 5916 -1606
tri 5901 -1642 5916 -1627 nw
rect 6235 -1627 6250 -1451
tri 6250 -1458 6263 -1445 nw
rect 6336 -1526 6351 -1298
tri 5873 -1648 5879 -1642 se
rect 5879 -1648 5888 -1642
rect 5873 -1664 5888 -1648
tri 5888 -1655 5901 -1642 nw
rect 6042 -1650 6059 -1636
rect 6091 -1650 6108 -1636
tri 6235 -1642 6250 -1627 ne
tri 6250 -1642 6272 -1620 sw
rect 5873 -1700 5888 -1692
rect 5954 -1664 6014 -1650
rect 5969 -1674 6014 -1664
rect 5969 -1692 5997 -1674
tri 5873 -1715 5888 -1700 ne
tri 5888 -1715 5910 -1693 sw
rect 5954 -1702 5997 -1692
rect 6012 -1678 6014 -1674
rect 6136 -1664 6196 -1650
tri 6250 -1655 6263 -1642 ne
rect 6263 -1648 6272 -1642
tri 6272 -1648 6278 -1642 sw
rect 6136 -1674 6181 -1664
rect 6012 -1702 6086 -1678
rect 5954 -1706 6086 -1702
tri 6086 -1706 6114 -1678 sw
rect 6136 -1688 6138 -1674
tri 6136 -1690 6138 -1688 ne
rect 6150 -1692 6181 -1674
rect 6150 -1702 6196 -1692
rect 6263 -1663 6278 -1648
tri 5888 -1727 5900 -1715 ne
rect 5900 -1720 5910 -1715
tri 5910 -1720 5915 -1715 sw
rect 5799 -2066 5814 -1838
rect 5900 -1876 5915 -1720
rect 5954 -1762 5982 -1706
tri 6074 -1724 6092 -1706 ne
rect 6092 -1726 6114 -1706
tri 6114 -1726 6134 -1706 sw
tri 6150 -1720 6168 -1702 ne
rect 5973 -1796 5982 -1762
rect 6016 -1735 6058 -1734
rect 6016 -1769 6021 -1735
rect 6051 -1769 6058 -1735
rect 6016 -1778 6058 -1769
rect 6092 -1735 6134 -1726
rect 6092 -1769 6099 -1735
rect 6129 -1769 6134 -1735
rect 6092 -1774 6134 -1769
rect 6168 -1762 6196 -1702
tri 6241 -1715 6263 -1693 se
rect 6263 -1700 6278 -1692
tri 6263 -1715 6278 -1700 nw
tri 6235 -1721 6241 -1715 se
rect 6241 -1721 6250 -1715
rect 5954 -1806 5982 -1796
tri 5982 -1806 6006 -1782 sw
rect 5954 -1838 5996 -1806
tri 6013 -1814 6014 -1813 sw
rect 6013 -1838 6014 -1814
tri 6016 -1815 6053 -1778 ne
rect 6053 -1806 6058 -1778
tri 6058 -1806 6084 -1780 sw
rect 6168 -1796 6177 -1762
rect 6168 -1806 6196 -1796
rect 6053 -1815 6137 -1806
tri 6053 -1834 6072 -1815 ne
rect 6072 -1834 6137 -1815
rect 5954 -1860 6014 -1838
rect 6136 -1838 6137 -1834
rect 6154 -1838 6196 -1806
rect 6136 -1860 6196 -1838
rect 6042 -1876 6059 -1862
rect 6091 -1876 6108 -1862
tri 5879 -1912 5901 -1890 se
rect 5901 -1897 5916 -1876
tri 5901 -1912 5916 -1897 nw
rect 6235 -1897 6250 -1721
tri 6250 -1728 6263 -1715 nw
rect 6336 -1796 6351 -1568
tri 5873 -1918 5879 -1912 se
rect 5879 -1918 5888 -1912
rect 5873 -1934 5888 -1918
tri 5888 -1925 5901 -1912 nw
rect 6042 -1920 6059 -1906
rect 6091 -1920 6108 -1906
tri 6235 -1912 6250 -1897 ne
tri 6250 -1912 6272 -1890 sw
rect 5873 -1970 5888 -1962
rect 5954 -1934 6014 -1920
rect 5969 -1944 6014 -1934
rect 5969 -1962 5997 -1944
tri 5873 -1985 5888 -1970 ne
tri 5888 -1985 5910 -1963 sw
rect 5954 -1972 5997 -1962
rect 6012 -1948 6014 -1944
rect 6136 -1934 6196 -1920
tri 6250 -1925 6263 -1912 ne
rect 6263 -1918 6272 -1912
tri 6272 -1918 6278 -1912 sw
rect 6136 -1944 6181 -1934
rect 6012 -1972 6086 -1948
rect 5954 -1976 6086 -1972
tri 6086 -1976 6114 -1948 sw
rect 6136 -1958 6138 -1944
tri 6136 -1960 6138 -1958 ne
rect 6150 -1962 6181 -1944
rect 6150 -1972 6196 -1962
rect 6263 -1933 6278 -1918
tri 5888 -1997 5900 -1985 ne
rect 5900 -1990 5910 -1985
tri 5910 -1990 5915 -1985 sw
rect 5799 -2146 5814 -2108
rect 5900 -2146 5915 -1990
rect 5954 -2032 5982 -1976
tri 6074 -1994 6092 -1976 ne
rect 6092 -1996 6114 -1976
tri 6114 -1996 6134 -1976 sw
tri 6150 -1990 6168 -1972 ne
rect 5973 -2066 5982 -2032
rect 6016 -2005 6058 -2004
rect 6016 -2039 6021 -2005
rect 6051 -2039 6058 -2005
rect 6016 -2048 6058 -2039
rect 6092 -2005 6134 -1996
rect 6092 -2039 6099 -2005
rect 6129 -2039 6134 -2005
rect 6092 -2044 6134 -2039
rect 6168 -2032 6196 -1972
tri 6241 -1985 6263 -1963 se
rect 6263 -1970 6278 -1962
tri 6263 -1985 6278 -1970 nw
tri 6235 -1991 6241 -1985 se
rect 6241 -1991 6250 -1985
rect 5954 -2076 5982 -2066
tri 5982 -2076 6006 -2052 sw
rect 5954 -2108 5996 -2076
tri 6013 -2084 6014 -2083 sw
rect 6013 -2108 6014 -2084
tri 6016 -2085 6053 -2048 ne
rect 6053 -2076 6058 -2048
tri 6058 -2076 6084 -2050 sw
rect 6168 -2066 6177 -2032
rect 6168 -2076 6196 -2066
rect 6053 -2085 6137 -2076
tri 6053 -2104 6072 -2085 ne
rect 6072 -2104 6137 -2085
rect 5954 -2130 6014 -2108
rect 6136 -2108 6137 -2104
rect 6154 -2108 6196 -2076
rect 6136 -2130 6196 -2108
rect 6042 -2146 6059 -2132
rect 6091 -2146 6108 -2132
rect 6235 -2146 6250 -1991
tri 6250 -1998 6263 -1985 nw
rect 6336 -2066 6351 -1838
rect 6336 -2146 6351 -2108
rect 6379 1984 6394 2174
tri 6459 2138 6481 2160 se
rect 6481 2153 6496 2174
tri 6481 2138 6496 2153 nw
rect 6815 2153 6830 2174
tri 6453 2132 6459 2138 se
rect 6459 2132 6468 2138
rect 6453 2116 6468 2132
tri 6468 2125 6481 2138 nw
rect 6622 2130 6639 2144
rect 6671 2130 6688 2144
tri 6815 2138 6830 2153 ne
tri 6830 2138 6852 2160 sw
rect 6453 2080 6468 2088
rect 6534 2116 6594 2130
rect 6549 2106 6594 2116
rect 6549 2088 6577 2106
tri 6453 2065 6468 2080 ne
tri 6468 2065 6490 2087 sw
rect 6534 2078 6577 2088
rect 6592 2102 6594 2106
rect 6716 2116 6776 2130
tri 6830 2125 6843 2138 ne
rect 6843 2132 6852 2138
tri 6852 2132 6858 2138 sw
rect 6716 2106 6761 2116
rect 6592 2078 6666 2102
rect 6534 2074 6666 2078
tri 6666 2074 6694 2102 sw
rect 6716 2092 6718 2106
tri 6716 2090 6718 2092 ne
rect 6730 2088 6761 2106
rect 6730 2078 6776 2088
rect 6843 2117 6858 2132
tri 6468 2053 6480 2065 ne
rect 6480 2060 6490 2065
tri 6490 2060 6495 2065 sw
rect 6379 1714 6394 1942
rect 6480 1904 6495 2060
rect 6534 2018 6562 2074
tri 6654 2056 6672 2074 ne
rect 6672 2054 6694 2074
tri 6694 2054 6714 2074 sw
tri 6730 2060 6748 2078 ne
rect 6553 1984 6562 2018
rect 6596 2045 6638 2046
rect 6596 2011 6601 2045
rect 6631 2011 6638 2045
rect 6596 2002 6638 2011
rect 6672 2045 6714 2054
rect 6672 2011 6679 2045
rect 6709 2011 6714 2045
rect 6672 2006 6714 2011
rect 6748 2018 6776 2078
tri 6821 2065 6843 2087 se
rect 6843 2080 6858 2088
tri 6843 2065 6858 2080 nw
tri 6815 2059 6821 2065 se
rect 6821 2059 6830 2065
rect 6534 1974 6562 1984
tri 6562 1974 6586 1998 sw
rect 6534 1942 6576 1974
tri 6593 1966 6594 1967 sw
rect 6593 1942 6594 1966
tri 6596 1965 6633 2002 ne
rect 6633 1974 6638 2002
tri 6638 1974 6664 2000 sw
rect 6748 1984 6757 2018
rect 6748 1974 6776 1984
rect 6633 1965 6717 1974
tri 6633 1946 6652 1965 ne
rect 6652 1946 6717 1965
rect 6534 1920 6594 1942
rect 6716 1942 6717 1946
rect 6734 1942 6776 1974
rect 6716 1920 6776 1942
rect 6622 1904 6639 1918
rect 6671 1904 6688 1918
tri 6459 1868 6481 1890 se
rect 6481 1883 6496 1904
tri 6481 1868 6496 1883 nw
rect 6815 1883 6830 2059
tri 6830 2052 6843 2065 nw
rect 6916 1984 6931 2174
tri 6453 1862 6459 1868 se
rect 6459 1862 6468 1868
rect 6453 1846 6468 1862
tri 6468 1855 6481 1868 nw
rect 6622 1860 6639 1874
rect 6671 1860 6688 1874
tri 6815 1868 6830 1883 ne
tri 6830 1868 6852 1890 sw
rect 6453 1810 6468 1818
rect 6534 1846 6594 1860
rect 6549 1836 6594 1846
rect 6549 1818 6577 1836
tri 6453 1795 6468 1810 ne
tri 6468 1795 6490 1817 sw
rect 6534 1808 6577 1818
rect 6592 1832 6594 1836
rect 6716 1846 6776 1860
tri 6830 1855 6843 1868 ne
rect 6843 1862 6852 1868
tri 6852 1862 6858 1868 sw
rect 6716 1836 6761 1846
rect 6592 1808 6666 1832
rect 6534 1804 6666 1808
tri 6666 1804 6694 1832 sw
rect 6716 1822 6718 1836
tri 6716 1820 6718 1822 ne
rect 6730 1818 6761 1836
rect 6730 1808 6776 1818
rect 6843 1847 6858 1862
tri 6468 1783 6480 1795 ne
rect 6480 1790 6490 1795
tri 6490 1790 6495 1795 sw
rect 6379 1444 6394 1672
rect 6480 1682 6495 1790
rect 6534 1748 6562 1804
tri 6654 1786 6672 1804 ne
rect 6672 1784 6694 1804
tri 6694 1784 6714 1804 sw
tri 6730 1790 6748 1808 ne
rect 6553 1714 6562 1748
rect 6596 1775 6638 1776
rect 6596 1741 6601 1775
rect 6631 1741 6638 1775
rect 6596 1732 6638 1741
rect 6672 1775 6714 1784
rect 6672 1741 6679 1775
rect 6709 1741 6714 1775
rect 6672 1736 6714 1741
rect 6748 1748 6776 1808
tri 6821 1795 6843 1817 se
rect 6843 1810 6858 1818
tri 6843 1795 6858 1810 nw
tri 6815 1789 6821 1795 se
rect 6821 1789 6830 1795
rect 6534 1704 6562 1714
tri 6562 1704 6586 1728 sw
rect 6480 1634 6496 1682
rect 6534 1672 6576 1704
tri 6593 1696 6594 1697 sw
rect 6593 1672 6594 1696
tri 6596 1695 6633 1732 ne
rect 6633 1704 6638 1732
tri 6638 1704 6664 1730 sw
rect 6748 1714 6757 1748
rect 6748 1704 6776 1714
rect 6633 1695 6717 1704
tri 6633 1676 6652 1695 ne
rect 6652 1676 6717 1695
rect 6534 1650 6594 1672
rect 6716 1672 6717 1676
rect 6734 1672 6776 1704
rect 6716 1650 6776 1672
rect 6622 1634 6639 1648
rect 6671 1634 6688 1648
tri 6459 1598 6481 1620 se
rect 6481 1613 6496 1634
tri 6481 1598 6496 1613 nw
rect 6815 1613 6830 1789
tri 6830 1782 6843 1795 nw
rect 6916 1714 6931 1942
tri 6453 1592 6459 1598 se
rect 6459 1592 6468 1598
rect 6453 1576 6468 1592
tri 6468 1585 6481 1598 nw
rect 6622 1590 6639 1604
rect 6671 1590 6688 1604
tri 6815 1598 6830 1613 ne
tri 6830 1598 6852 1620 sw
rect 6453 1540 6468 1548
rect 6534 1576 6594 1590
rect 6549 1566 6594 1576
rect 6549 1548 6577 1566
tri 6453 1525 6468 1540 ne
tri 6468 1525 6490 1547 sw
rect 6534 1538 6577 1548
rect 6592 1562 6594 1566
rect 6716 1576 6776 1590
tri 6830 1585 6843 1598 ne
rect 6843 1592 6852 1598
tri 6852 1592 6858 1598 sw
rect 6716 1566 6761 1576
rect 6592 1538 6666 1562
rect 6534 1534 6666 1538
tri 6666 1534 6694 1562 sw
rect 6716 1552 6718 1566
tri 6716 1550 6718 1552 ne
rect 6730 1548 6761 1566
rect 6730 1538 6776 1548
rect 6843 1577 6858 1592
tri 6468 1513 6480 1525 ne
rect 6480 1520 6490 1525
tri 6490 1520 6495 1525 sw
rect 6379 1174 6394 1402
rect 6480 1364 6495 1520
rect 6534 1478 6562 1534
tri 6654 1516 6672 1534 ne
rect 6672 1514 6694 1534
tri 6694 1514 6714 1534 sw
tri 6730 1520 6748 1538 ne
rect 6553 1444 6562 1478
rect 6596 1505 6638 1506
rect 6596 1471 6601 1505
rect 6631 1471 6638 1505
rect 6596 1462 6638 1471
rect 6672 1505 6714 1514
rect 6672 1471 6679 1505
rect 6709 1471 6714 1505
rect 6672 1466 6714 1471
rect 6748 1478 6776 1538
tri 6821 1525 6843 1547 se
rect 6843 1540 6858 1548
tri 6843 1525 6858 1540 nw
tri 6815 1519 6821 1525 se
rect 6821 1519 6830 1525
rect 6534 1434 6562 1444
tri 6562 1434 6586 1458 sw
rect 6534 1402 6576 1434
tri 6593 1426 6594 1427 sw
rect 6593 1402 6594 1426
tri 6596 1425 6633 1462 ne
rect 6633 1434 6638 1462
tri 6638 1434 6664 1460 sw
rect 6748 1444 6757 1478
rect 6748 1434 6776 1444
rect 6633 1425 6717 1434
tri 6633 1406 6652 1425 ne
rect 6652 1406 6717 1425
rect 6534 1380 6594 1402
rect 6716 1402 6717 1406
rect 6734 1402 6776 1434
rect 6716 1380 6776 1402
rect 6622 1364 6639 1378
rect 6671 1364 6688 1378
tri 6459 1328 6481 1350 se
rect 6481 1343 6496 1364
tri 6481 1328 6496 1343 nw
rect 6815 1343 6830 1519
tri 6830 1512 6843 1525 nw
rect 6916 1444 6931 1672
tri 6453 1322 6459 1328 se
rect 6459 1322 6468 1328
rect 6453 1306 6468 1322
tri 6468 1315 6481 1328 nw
rect 6622 1320 6639 1334
rect 6671 1320 6688 1334
tri 6815 1328 6830 1343 ne
tri 6830 1328 6852 1350 sw
rect 6453 1270 6468 1278
rect 6534 1306 6594 1320
rect 6549 1296 6594 1306
rect 6549 1278 6577 1296
tri 6453 1255 6468 1270 ne
tri 6468 1255 6490 1277 sw
rect 6534 1268 6577 1278
rect 6592 1292 6594 1296
rect 6716 1306 6776 1320
tri 6830 1315 6843 1328 ne
rect 6843 1322 6852 1328
tri 6852 1322 6858 1328 sw
rect 6716 1296 6761 1306
rect 6592 1268 6666 1292
rect 6534 1264 6666 1268
tri 6666 1264 6694 1292 sw
rect 6716 1282 6718 1296
tri 6716 1280 6718 1282 ne
rect 6730 1278 6761 1296
rect 6730 1268 6776 1278
rect 6843 1307 6858 1322
tri 6468 1243 6480 1255 ne
rect 6480 1250 6490 1255
tri 6490 1250 6495 1255 sw
rect 6379 904 6394 1132
rect 6480 1142 6495 1250
rect 6534 1208 6562 1264
tri 6654 1246 6672 1264 ne
rect 6672 1244 6694 1264
tri 6694 1244 6714 1264 sw
tri 6730 1250 6748 1268 ne
rect 6553 1174 6562 1208
rect 6596 1235 6638 1236
rect 6596 1201 6601 1235
rect 6631 1201 6638 1235
rect 6596 1192 6638 1201
rect 6672 1235 6714 1244
rect 6672 1201 6679 1235
rect 6709 1201 6714 1235
rect 6672 1196 6714 1201
rect 6748 1208 6776 1268
tri 6821 1255 6843 1277 se
rect 6843 1270 6858 1278
tri 6843 1255 6858 1270 nw
tri 6815 1249 6821 1255 se
rect 6821 1249 6830 1255
rect 6534 1164 6562 1174
tri 6562 1164 6586 1188 sw
rect 6480 1094 6496 1142
rect 6534 1132 6576 1164
tri 6593 1156 6594 1157 sw
rect 6593 1132 6594 1156
tri 6596 1155 6633 1192 ne
rect 6633 1164 6638 1192
tri 6638 1164 6664 1190 sw
rect 6748 1174 6757 1208
rect 6748 1164 6776 1174
rect 6633 1155 6717 1164
tri 6633 1136 6652 1155 ne
rect 6652 1136 6717 1155
rect 6534 1110 6594 1132
rect 6716 1132 6717 1136
rect 6734 1132 6776 1164
rect 6716 1110 6776 1132
rect 6622 1094 6639 1108
rect 6671 1094 6688 1108
tri 6459 1058 6481 1080 se
rect 6481 1073 6496 1094
tri 6481 1058 6496 1073 nw
rect 6815 1073 6830 1249
tri 6830 1242 6843 1255 nw
rect 6916 1174 6931 1402
tri 6453 1052 6459 1058 se
rect 6459 1052 6468 1058
rect 6453 1036 6468 1052
tri 6468 1045 6481 1058 nw
rect 6622 1050 6639 1064
rect 6671 1050 6688 1064
tri 6815 1058 6830 1073 ne
tri 6830 1058 6852 1080 sw
rect 6453 1000 6468 1008
rect 6534 1036 6594 1050
rect 6549 1026 6594 1036
rect 6549 1008 6577 1026
tri 6453 985 6468 1000 ne
tri 6468 985 6490 1007 sw
rect 6534 998 6577 1008
rect 6592 1022 6594 1026
rect 6716 1036 6776 1050
tri 6830 1045 6843 1058 ne
rect 6843 1052 6852 1058
tri 6852 1052 6858 1058 sw
rect 6716 1026 6761 1036
rect 6592 998 6666 1022
rect 6534 994 6666 998
tri 6666 994 6694 1022 sw
rect 6716 1012 6718 1026
tri 6716 1010 6718 1012 ne
rect 6730 1008 6761 1026
rect 6730 998 6776 1008
rect 6843 1037 6858 1052
tri 6468 973 6480 985 ne
rect 6480 980 6490 985
tri 6490 980 6495 985 sw
rect 6379 634 6394 862
rect 6480 824 6495 980
rect 6534 938 6562 994
tri 6654 976 6672 994 ne
rect 6672 974 6694 994
tri 6694 974 6714 994 sw
tri 6730 980 6748 998 ne
rect 6553 904 6562 938
rect 6596 965 6638 966
rect 6596 931 6601 965
rect 6631 931 6638 965
rect 6596 922 6638 931
rect 6672 965 6714 974
rect 6672 931 6679 965
rect 6709 931 6714 965
rect 6672 926 6714 931
rect 6748 938 6776 998
tri 6821 985 6843 1007 se
rect 6843 1000 6858 1008
tri 6843 985 6858 1000 nw
tri 6815 979 6821 985 se
rect 6821 979 6830 985
rect 6534 894 6562 904
tri 6562 894 6586 918 sw
rect 6534 862 6576 894
tri 6593 886 6594 887 sw
rect 6593 862 6594 886
tri 6596 885 6633 922 ne
rect 6633 894 6638 922
tri 6638 894 6664 920 sw
rect 6748 904 6757 938
rect 6748 894 6776 904
rect 6633 885 6717 894
tri 6633 866 6652 885 ne
rect 6652 866 6717 885
rect 6534 840 6594 862
rect 6716 862 6717 866
rect 6734 862 6776 894
rect 6716 840 6776 862
rect 6622 824 6639 838
rect 6671 824 6688 838
tri 6459 788 6481 810 se
rect 6481 803 6496 824
tri 6481 788 6496 803 nw
rect 6815 803 6830 979
tri 6830 972 6843 985 nw
rect 6916 904 6931 1132
tri 6453 782 6459 788 se
rect 6459 782 6468 788
rect 6453 766 6468 782
tri 6468 775 6481 788 nw
rect 6622 780 6639 794
rect 6671 780 6688 794
tri 6815 788 6830 803 ne
tri 6830 788 6852 810 sw
rect 6453 730 6468 738
rect 6534 766 6594 780
rect 6549 756 6594 766
rect 6549 738 6577 756
tri 6453 715 6468 730 ne
tri 6468 715 6490 737 sw
rect 6534 728 6577 738
rect 6592 752 6594 756
rect 6716 766 6776 780
tri 6830 775 6843 788 ne
rect 6843 782 6852 788
tri 6852 782 6858 788 sw
rect 6716 756 6761 766
rect 6592 728 6666 752
rect 6534 724 6666 728
tri 6666 724 6694 752 sw
rect 6716 742 6718 756
tri 6716 740 6718 742 ne
rect 6730 738 6761 756
rect 6730 728 6776 738
rect 6843 767 6858 782
tri 6468 703 6480 715 ne
rect 6480 710 6490 715
tri 6490 710 6495 715 sw
rect 6379 364 6394 592
rect 6480 602 6495 710
rect 6534 668 6562 724
tri 6654 706 6672 724 ne
rect 6672 704 6694 724
tri 6694 704 6714 724 sw
tri 6730 710 6748 728 ne
rect 6553 634 6562 668
rect 6596 695 6638 696
rect 6596 661 6601 695
rect 6631 661 6638 695
rect 6596 652 6638 661
rect 6672 695 6714 704
rect 6672 661 6679 695
rect 6709 661 6714 695
rect 6672 656 6714 661
rect 6748 668 6776 728
tri 6821 715 6843 737 se
rect 6843 730 6858 738
tri 6843 715 6858 730 nw
tri 6815 709 6821 715 se
rect 6821 709 6830 715
rect 6534 624 6562 634
tri 6562 624 6586 648 sw
rect 6480 554 6496 602
rect 6534 592 6576 624
tri 6593 616 6594 617 sw
rect 6593 592 6594 616
tri 6596 615 6633 652 ne
rect 6633 624 6638 652
tri 6638 624 6664 650 sw
rect 6748 634 6757 668
rect 6748 624 6776 634
rect 6633 615 6717 624
tri 6633 596 6652 615 ne
rect 6652 596 6717 615
rect 6534 570 6594 592
rect 6716 592 6717 596
rect 6734 592 6776 624
rect 6716 570 6776 592
rect 6622 554 6639 568
rect 6671 554 6688 568
tri 6459 518 6481 540 se
rect 6481 533 6496 554
tri 6481 518 6496 533 nw
rect 6815 533 6830 709
tri 6830 702 6843 715 nw
rect 6916 634 6931 862
tri 6453 512 6459 518 se
rect 6459 512 6468 518
rect 6453 496 6468 512
tri 6468 505 6481 518 nw
rect 6622 510 6639 524
rect 6671 510 6688 524
tri 6815 518 6830 533 ne
tri 6830 518 6852 540 sw
rect 6453 460 6468 468
rect 6534 496 6594 510
rect 6549 486 6594 496
rect 6549 468 6577 486
tri 6453 445 6468 460 ne
tri 6468 445 6490 467 sw
rect 6534 458 6577 468
rect 6592 482 6594 486
rect 6716 496 6776 510
tri 6830 505 6843 518 ne
rect 6843 512 6852 518
tri 6852 512 6858 518 sw
rect 6716 486 6761 496
rect 6592 458 6666 482
rect 6534 454 6666 458
tri 6666 454 6694 482 sw
rect 6716 472 6718 486
tri 6716 470 6718 472 ne
rect 6730 468 6761 486
rect 6730 458 6776 468
rect 6843 497 6858 512
tri 6468 433 6480 445 ne
rect 6480 440 6490 445
tri 6490 440 6495 445 sw
rect 6379 94 6394 322
rect 6480 284 6495 440
rect 6534 398 6562 454
tri 6654 436 6672 454 ne
rect 6672 434 6694 454
tri 6694 434 6714 454 sw
tri 6730 440 6748 458 ne
rect 6553 364 6562 398
rect 6596 425 6638 426
rect 6596 391 6601 425
rect 6631 391 6638 425
rect 6596 382 6638 391
rect 6672 425 6714 434
rect 6672 391 6679 425
rect 6709 391 6714 425
rect 6672 386 6714 391
rect 6748 398 6776 458
tri 6821 445 6843 467 se
rect 6843 460 6858 468
tri 6843 445 6858 460 nw
tri 6815 439 6821 445 se
rect 6821 439 6830 445
rect 6534 354 6562 364
tri 6562 354 6586 378 sw
rect 6534 322 6576 354
tri 6593 346 6594 347 sw
rect 6593 322 6594 346
tri 6596 345 6633 382 ne
rect 6633 354 6638 382
tri 6638 354 6664 380 sw
rect 6748 364 6757 398
rect 6748 354 6776 364
rect 6633 345 6717 354
tri 6633 326 6652 345 ne
rect 6652 326 6717 345
rect 6534 300 6594 322
rect 6716 322 6717 326
rect 6734 322 6776 354
rect 6716 300 6776 322
rect 6622 284 6639 298
rect 6671 284 6688 298
tri 6459 248 6481 270 se
rect 6481 263 6496 284
tri 6481 248 6496 263 nw
rect 6815 263 6830 439
tri 6830 432 6843 445 nw
rect 6916 364 6931 592
tri 6453 242 6459 248 se
rect 6459 242 6468 248
rect 6453 226 6468 242
tri 6468 235 6481 248 nw
rect 6622 240 6639 254
rect 6671 240 6688 254
tri 6815 248 6830 263 ne
tri 6830 248 6852 270 sw
rect 6453 190 6468 198
rect 6534 226 6594 240
rect 6549 216 6594 226
rect 6549 198 6577 216
tri 6453 175 6468 190 ne
tri 6468 175 6490 197 sw
rect 6534 188 6577 198
rect 6592 212 6594 216
rect 6716 226 6776 240
tri 6830 235 6843 248 ne
rect 6843 242 6852 248
tri 6852 242 6858 248 sw
rect 6716 216 6761 226
rect 6592 188 6666 212
rect 6534 184 6666 188
tri 6666 184 6694 212 sw
rect 6716 202 6718 216
tri 6716 200 6718 202 ne
rect 6730 198 6761 216
rect 6730 188 6776 198
rect 6843 227 6858 242
tri 6468 163 6480 175 ne
rect 6480 170 6490 175
tri 6490 170 6495 175 sw
rect 6379 -176 6394 52
rect 6480 62 6495 170
rect 6534 128 6562 184
tri 6654 166 6672 184 ne
rect 6672 164 6694 184
tri 6694 164 6714 184 sw
tri 6730 170 6748 188 ne
rect 6553 94 6562 128
rect 6596 155 6638 156
rect 6596 121 6601 155
rect 6631 121 6638 155
rect 6596 112 6638 121
rect 6672 155 6714 164
rect 6672 121 6679 155
rect 6709 121 6714 155
rect 6672 116 6714 121
rect 6748 128 6776 188
tri 6821 175 6843 197 se
rect 6843 190 6858 198
tri 6843 175 6858 190 nw
tri 6815 169 6821 175 se
rect 6821 169 6830 175
rect 6534 84 6562 94
tri 6562 84 6586 108 sw
rect 6480 14 6496 62
rect 6534 52 6576 84
tri 6593 76 6594 77 sw
rect 6593 52 6594 76
tri 6596 75 6633 112 ne
rect 6633 84 6638 112
tri 6638 84 6664 110 sw
rect 6748 94 6757 128
rect 6748 84 6776 94
rect 6633 75 6717 84
tri 6633 56 6652 75 ne
rect 6652 56 6717 75
rect 6534 30 6594 52
rect 6716 52 6717 56
rect 6734 52 6776 84
rect 6716 30 6776 52
rect 6622 14 6639 28
rect 6671 14 6688 28
tri 6459 -22 6481 0 se
rect 6481 -7 6496 14
tri 6481 -22 6496 -7 nw
rect 6815 -7 6830 169
tri 6830 162 6843 175 nw
rect 6916 94 6931 322
tri 6453 -28 6459 -22 se
rect 6459 -28 6468 -22
rect 6453 -44 6468 -28
tri 6468 -35 6481 -22 nw
rect 6622 -30 6639 -16
rect 6671 -30 6688 -16
tri 6815 -22 6830 -7 ne
tri 6830 -22 6852 0 sw
rect 6453 -80 6468 -72
rect 6534 -44 6594 -30
rect 6549 -54 6594 -44
rect 6549 -72 6577 -54
tri 6453 -95 6468 -80 ne
tri 6468 -95 6490 -73 sw
rect 6534 -82 6577 -72
rect 6592 -58 6594 -54
rect 6716 -44 6776 -30
tri 6830 -35 6843 -22 ne
rect 6843 -28 6852 -22
tri 6852 -28 6858 -22 sw
rect 6716 -54 6761 -44
rect 6592 -82 6666 -58
rect 6534 -86 6666 -82
tri 6666 -86 6694 -58 sw
rect 6716 -68 6718 -54
tri 6716 -70 6718 -68 ne
rect 6730 -72 6761 -54
rect 6730 -82 6776 -72
rect 6843 -43 6858 -28
tri 6468 -107 6480 -95 ne
rect 6480 -100 6490 -95
tri 6490 -100 6495 -95 sw
rect 6379 -446 6394 -218
rect 6480 -256 6495 -100
rect 6534 -142 6562 -86
tri 6654 -104 6672 -86 ne
rect 6672 -106 6694 -86
tri 6694 -106 6714 -86 sw
tri 6730 -100 6748 -82 ne
rect 6553 -176 6562 -142
rect 6596 -115 6638 -114
rect 6596 -149 6601 -115
rect 6631 -149 6638 -115
rect 6596 -158 6638 -149
rect 6672 -115 6714 -106
rect 6672 -149 6679 -115
rect 6709 -149 6714 -115
rect 6672 -154 6714 -149
rect 6748 -142 6776 -82
tri 6821 -95 6843 -73 se
rect 6843 -80 6858 -72
tri 6843 -95 6858 -80 nw
tri 6815 -101 6821 -95 se
rect 6821 -101 6830 -95
rect 6534 -186 6562 -176
tri 6562 -186 6586 -162 sw
rect 6534 -218 6576 -186
tri 6593 -194 6594 -193 sw
rect 6593 -218 6594 -194
tri 6596 -195 6633 -158 ne
rect 6633 -186 6638 -158
tri 6638 -186 6664 -160 sw
rect 6748 -176 6757 -142
rect 6748 -186 6776 -176
rect 6633 -195 6717 -186
tri 6633 -214 6652 -195 ne
rect 6652 -214 6717 -195
rect 6534 -240 6594 -218
rect 6716 -218 6717 -214
rect 6734 -218 6776 -186
rect 6716 -240 6776 -218
rect 6622 -256 6639 -242
rect 6671 -256 6688 -242
tri 6459 -292 6481 -270 se
rect 6481 -277 6496 -256
tri 6481 -292 6496 -277 nw
rect 6815 -277 6830 -101
tri 6830 -108 6843 -95 nw
rect 6916 -176 6931 52
tri 6453 -298 6459 -292 se
rect 6459 -298 6468 -292
rect 6453 -314 6468 -298
tri 6468 -305 6481 -292 nw
rect 6622 -300 6639 -286
rect 6671 -300 6688 -286
tri 6815 -292 6830 -277 ne
tri 6830 -292 6852 -270 sw
rect 6453 -350 6468 -342
rect 6534 -314 6594 -300
rect 6549 -324 6594 -314
rect 6549 -342 6577 -324
tri 6453 -365 6468 -350 ne
tri 6468 -365 6490 -343 sw
rect 6534 -352 6577 -342
rect 6592 -328 6594 -324
rect 6716 -314 6776 -300
tri 6830 -305 6843 -292 ne
rect 6843 -298 6852 -292
tri 6852 -298 6858 -292 sw
rect 6716 -324 6761 -314
rect 6592 -352 6666 -328
rect 6534 -356 6666 -352
tri 6666 -356 6694 -328 sw
rect 6716 -338 6718 -324
tri 6716 -340 6718 -338 ne
rect 6730 -342 6761 -324
rect 6730 -352 6776 -342
rect 6843 -313 6858 -298
tri 6468 -377 6480 -365 ne
rect 6480 -370 6490 -365
tri 6490 -370 6495 -365 sw
rect 6379 -716 6394 -488
rect 6480 -478 6495 -370
rect 6534 -412 6562 -356
tri 6654 -374 6672 -356 ne
rect 6672 -376 6694 -356
tri 6694 -376 6714 -356 sw
tri 6730 -370 6748 -352 ne
rect 6553 -446 6562 -412
rect 6596 -385 6638 -384
rect 6596 -419 6601 -385
rect 6631 -419 6638 -385
rect 6596 -428 6638 -419
rect 6672 -385 6714 -376
rect 6672 -419 6679 -385
rect 6709 -419 6714 -385
rect 6672 -424 6714 -419
rect 6748 -412 6776 -352
tri 6821 -365 6843 -343 se
rect 6843 -350 6858 -342
tri 6843 -365 6858 -350 nw
tri 6815 -371 6821 -365 se
rect 6821 -371 6830 -365
rect 6534 -456 6562 -446
tri 6562 -456 6586 -432 sw
rect 6480 -526 6496 -478
rect 6534 -488 6576 -456
tri 6593 -464 6594 -463 sw
rect 6593 -488 6594 -464
tri 6596 -465 6633 -428 ne
rect 6633 -456 6638 -428
tri 6638 -456 6664 -430 sw
rect 6748 -446 6757 -412
rect 6748 -456 6776 -446
rect 6633 -465 6717 -456
tri 6633 -484 6652 -465 ne
rect 6652 -484 6717 -465
rect 6534 -510 6594 -488
rect 6716 -488 6717 -484
rect 6734 -488 6776 -456
rect 6716 -510 6776 -488
rect 6622 -526 6639 -512
rect 6671 -526 6688 -512
tri 6459 -562 6481 -540 se
rect 6481 -547 6496 -526
tri 6481 -562 6496 -547 nw
rect 6815 -547 6830 -371
tri 6830 -378 6843 -365 nw
rect 6916 -446 6931 -218
tri 6453 -568 6459 -562 se
rect 6459 -568 6468 -562
rect 6453 -584 6468 -568
tri 6468 -575 6481 -562 nw
rect 6622 -570 6639 -556
rect 6671 -570 6688 -556
tri 6815 -562 6830 -547 ne
tri 6830 -562 6852 -540 sw
rect 6453 -620 6468 -612
rect 6534 -584 6594 -570
rect 6549 -594 6594 -584
rect 6549 -612 6577 -594
tri 6453 -635 6468 -620 ne
tri 6468 -635 6490 -613 sw
rect 6534 -622 6577 -612
rect 6592 -598 6594 -594
rect 6716 -584 6776 -570
tri 6830 -575 6843 -562 ne
rect 6843 -568 6852 -562
tri 6852 -568 6858 -562 sw
rect 6716 -594 6761 -584
rect 6592 -622 6666 -598
rect 6534 -626 6666 -622
tri 6666 -626 6694 -598 sw
rect 6716 -608 6718 -594
tri 6716 -610 6718 -608 ne
rect 6730 -612 6761 -594
rect 6730 -622 6776 -612
rect 6843 -583 6858 -568
tri 6468 -647 6480 -635 ne
rect 6480 -640 6490 -635
tri 6490 -640 6495 -635 sw
rect 6379 -986 6394 -758
rect 6480 -796 6495 -640
rect 6534 -682 6562 -626
tri 6654 -644 6672 -626 ne
rect 6672 -646 6694 -626
tri 6694 -646 6714 -626 sw
tri 6730 -640 6748 -622 ne
rect 6553 -716 6562 -682
rect 6596 -655 6638 -654
rect 6596 -689 6601 -655
rect 6631 -689 6638 -655
rect 6596 -698 6638 -689
rect 6672 -655 6714 -646
rect 6672 -689 6679 -655
rect 6709 -689 6714 -655
rect 6672 -694 6714 -689
rect 6748 -682 6776 -622
tri 6821 -635 6843 -613 se
rect 6843 -620 6858 -612
tri 6843 -635 6858 -620 nw
tri 6815 -641 6821 -635 se
rect 6821 -641 6830 -635
rect 6534 -726 6562 -716
tri 6562 -726 6586 -702 sw
rect 6534 -758 6576 -726
tri 6593 -734 6594 -733 sw
rect 6593 -758 6594 -734
tri 6596 -735 6633 -698 ne
rect 6633 -726 6638 -698
tri 6638 -726 6664 -700 sw
rect 6748 -716 6757 -682
rect 6748 -726 6776 -716
rect 6633 -735 6717 -726
tri 6633 -754 6652 -735 ne
rect 6652 -754 6717 -735
rect 6534 -780 6594 -758
rect 6716 -758 6717 -754
rect 6734 -758 6776 -726
rect 6716 -780 6776 -758
rect 6622 -796 6639 -782
rect 6671 -796 6688 -782
tri 6459 -832 6481 -810 se
rect 6481 -817 6496 -796
tri 6481 -832 6496 -817 nw
rect 6815 -817 6830 -641
tri 6830 -648 6843 -635 nw
rect 6916 -716 6931 -488
tri 6453 -838 6459 -832 se
rect 6459 -838 6468 -832
rect 6453 -854 6468 -838
tri 6468 -845 6481 -832 nw
rect 6622 -840 6639 -826
rect 6671 -840 6688 -826
tri 6815 -832 6830 -817 ne
tri 6830 -832 6852 -810 sw
rect 6453 -890 6468 -882
rect 6534 -854 6594 -840
rect 6549 -864 6594 -854
rect 6549 -882 6577 -864
tri 6453 -905 6468 -890 ne
tri 6468 -905 6490 -883 sw
rect 6534 -892 6577 -882
rect 6592 -868 6594 -864
rect 6716 -854 6776 -840
tri 6830 -845 6843 -832 ne
rect 6843 -838 6852 -832
tri 6852 -838 6858 -832 sw
rect 6716 -864 6761 -854
rect 6592 -892 6666 -868
rect 6534 -896 6666 -892
tri 6666 -896 6694 -868 sw
rect 6716 -878 6718 -864
tri 6716 -880 6718 -878 ne
rect 6730 -882 6761 -864
rect 6730 -892 6776 -882
rect 6843 -853 6858 -838
tri 6468 -917 6480 -905 ne
rect 6480 -910 6490 -905
tri 6490 -910 6495 -905 sw
rect 6379 -1256 6394 -1028
rect 6480 -1018 6495 -910
rect 6534 -952 6562 -896
tri 6654 -914 6672 -896 ne
rect 6672 -916 6694 -896
tri 6694 -916 6714 -896 sw
tri 6730 -910 6748 -892 ne
rect 6553 -986 6562 -952
rect 6596 -925 6638 -924
rect 6596 -959 6601 -925
rect 6631 -959 6638 -925
rect 6596 -968 6638 -959
rect 6672 -925 6714 -916
rect 6672 -959 6679 -925
rect 6709 -959 6714 -925
rect 6672 -964 6714 -959
rect 6748 -952 6776 -892
tri 6821 -905 6843 -883 se
rect 6843 -890 6858 -882
tri 6843 -905 6858 -890 nw
tri 6815 -911 6821 -905 se
rect 6821 -911 6830 -905
rect 6534 -996 6562 -986
tri 6562 -996 6586 -972 sw
rect 6480 -1066 6496 -1018
rect 6534 -1028 6576 -996
tri 6593 -1004 6594 -1003 sw
rect 6593 -1028 6594 -1004
tri 6596 -1005 6633 -968 ne
rect 6633 -996 6638 -968
tri 6638 -996 6664 -970 sw
rect 6748 -986 6757 -952
rect 6748 -996 6776 -986
rect 6633 -1005 6717 -996
tri 6633 -1024 6652 -1005 ne
rect 6652 -1024 6717 -1005
rect 6534 -1050 6594 -1028
rect 6716 -1028 6717 -1024
rect 6734 -1028 6776 -996
rect 6716 -1050 6776 -1028
rect 6622 -1066 6639 -1052
rect 6671 -1066 6688 -1052
tri 6459 -1102 6481 -1080 se
rect 6481 -1087 6496 -1066
tri 6481 -1102 6496 -1087 nw
rect 6815 -1087 6830 -911
tri 6830 -918 6843 -905 nw
rect 6916 -986 6931 -758
tri 6453 -1108 6459 -1102 se
rect 6459 -1108 6468 -1102
rect 6453 -1124 6468 -1108
tri 6468 -1115 6481 -1102 nw
rect 6622 -1110 6639 -1096
rect 6671 -1110 6688 -1096
tri 6815 -1102 6830 -1087 ne
tri 6830 -1102 6852 -1080 sw
rect 6453 -1160 6468 -1152
rect 6534 -1124 6594 -1110
rect 6549 -1134 6594 -1124
rect 6549 -1152 6577 -1134
tri 6453 -1175 6468 -1160 ne
tri 6468 -1175 6490 -1153 sw
rect 6534 -1162 6577 -1152
rect 6592 -1138 6594 -1134
rect 6716 -1124 6776 -1110
tri 6830 -1115 6843 -1102 ne
rect 6843 -1108 6852 -1102
tri 6852 -1108 6858 -1102 sw
rect 6716 -1134 6761 -1124
rect 6592 -1162 6666 -1138
rect 6534 -1166 6666 -1162
tri 6666 -1166 6694 -1138 sw
rect 6716 -1148 6718 -1134
tri 6716 -1150 6718 -1148 ne
rect 6730 -1152 6761 -1134
rect 6730 -1162 6776 -1152
rect 6843 -1123 6858 -1108
tri 6468 -1187 6480 -1175 ne
rect 6480 -1180 6490 -1175
tri 6490 -1180 6495 -1175 sw
rect 6379 -1526 6394 -1298
rect 6480 -1336 6495 -1180
rect 6534 -1222 6562 -1166
tri 6654 -1184 6672 -1166 ne
rect 6672 -1186 6694 -1166
tri 6694 -1186 6714 -1166 sw
tri 6730 -1180 6748 -1162 ne
rect 6553 -1256 6562 -1222
rect 6596 -1195 6638 -1194
rect 6596 -1229 6601 -1195
rect 6631 -1229 6638 -1195
rect 6596 -1238 6638 -1229
rect 6672 -1195 6714 -1186
rect 6672 -1229 6679 -1195
rect 6709 -1229 6714 -1195
rect 6672 -1234 6714 -1229
rect 6748 -1222 6776 -1162
tri 6821 -1175 6843 -1153 se
rect 6843 -1160 6858 -1152
tri 6843 -1175 6858 -1160 nw
tri 6815 -1181 6821 -1175 se
rect 6821 -1181 6830 -1175
rect 6534 -1266 6562 -1256
tri 6562 -1266 6586 -1242 sw
rect 6534 -1298 6576 -1266
tri 6593 -1274 6594 -1273 sw
rect 6593 -1298 6594 -1274
tri 6596 -1275 6633 -1238 ne
rect 6633 -1266 6638 -1238
tri 6638 -1266 6664 -1240 sw
rect 6748 -1256 6757 -1222
rect 6748 -1266 6776 -1256
rect 6633 -1275 6717 -1266
tri 6633 -1294 6652 -1275 ne
rect 6652 -1294 6717 -1275
rect 6534 -1320 6594 -1298
rect 6716 -1298 6717 -1294
rect 6734 -1298 6776 -1266
rect 6716 -1320 6776 -1298
rect 6622 -1336 6639 -1322
rect 6671 -1336 6688 -1322
tri 6459 -1372 6481 -1350 se
rect 6481 -1357 6496 -1336
tri 6481 -1372 6496 -1357 nw
rect 6815 -1357 6830 -1181
tri 6830 -1188 6843 -1175 nw
rect 6916 -1256 6931 -1028
tri 6453 -1378 6459 -1372 se
rect 6459 -1378 6468 -1372
rect 6453 -1394 6468 -1378
tri 6468 -1385 6481 -1372 nw
rect 6622 -1380 6639 -1366
rect 6671 -1380 6688 -1366
tri 6815 -1372 6830 -1357 ne
tri 6830 -1372 6852 -1350 sw
rect 6453 -1430 6468 -1422
rect 6534 -1394 6594 -1380
rect 6549 -1404 6594 -1394
rect 6549 -1422 6577 -1404
tri 6453 -1445 6468 -1430 ne
tri 6468 -1445 6490 -1423 sw
rect 6534 -1432 6577 -1422
rect 6592 -1408 6594 -1404
rect 6716 -1394 6776 -1380
tri 6830 -1385 6843 -1372 ne
rect 6843 -1378 6852 -1372
tri 6852 -1378 6858 -1372 sw
rect 6716 -1404 6761 -1394
rect 6592 -1432 6666 -1408
rect 6534 -1436 6666 -1432
tri 6666 -1436 6694 -1408 sw
rect 6716 -1418 6718 -1404
tri 6716 -1420 6718 -1418 ne
rect 6730 -1422 6761 -1404
rect 6730 -1432 6776 -1422
rect 6843 -1393 6858 -1378
tri 6468 -1457 6480 -1445 ne
rect 6480 -1450 6490 -1445
tri 6490 -1450 6495 -1445 sw
rect 6379 -1796 6394 -1568
rect 6480 -1558 6495 -1450
rect 6534 -1492 6562 -1436
tri 6654 -1454 6672 -1436 ne
rect 6672 -1456 6694 -1436
tri 6694 -1456 6714 -1436 sw
tri 6730 -1450 6748 -1432 ne
rect 6553 -1526 6562 -1492
rect 6596 -1465 6638 -1464
rect 6596 -1499 6601 -1465
rect 6631 -1499 6638 -1465
rect 6596 -1508 6638 -1499
rect 6672 -1465 6714 -1456
rect 6672 -1499 6679 -1465
rect 6709 -1499 6714 -1465
rect 6672 -1504 6714 -1499
rect 6748 -1492 6776 -1432
tri 6821 -1445 6843 -1423 se
rect 6843 -1430 6858 -1422
tri 6843 -1445 6858 -1430 nw
tri 6815 -1451 6821 -1445 se
rect 6821 -1451 6830 -1445
rect 6534 -1536 6562 -1526
tri 6562 -1536 6586 -1512 sw
rect 6480 -1606 6496 -1558
rect 6534 -1568 6576 -1536
tri 6593 -1544 6594 -1543 sw
rect 6593 -1568 6594 -1544
tri 6596 -1545 6633 -1508 ne
rect 6633 -1536 6638 -1508
tri 6638 -1536 6664 -1510 sw
rect 6748 -1526 6757 -1492
rect 6748 -1536 6776 -1526
rect 6633 -1545 6717 -1536
tri 6633 -1564 6652 -1545 ne
rect 6652 -1564 6717 -1545
rect 6534 -1590 6594 -1568
rect 6716 -1568 6717 -1564
rect 6734 -1568 6776 -1536
rect 6716 -1590 6776 -1568
rect 6622 -1606 6639 -1592
rect 6671 -1606 6688 -1592
tri 6459 -1642 6481 -1620 se
rect 6481 -1627 6496 -1606
tri 6481 -1642 6496 -1627 nw
rect 6815 -1627 6830 -1451
tri 6830 -1458 6843 -1445 nw
rect 6916 -1526 6931 -1298
tri 6453 -1648 6459 -1642 se
rect 6459 -1648 6468 -1642
rect 6453 -1664 6468 -1648
tri 6468 -1655 6481 -1642 nw
rect 6622 -1650 6639 -1636
rect 6671 -1650 6688 -1636
tri 6815 -1642 6830 -1627 ne
tri 6830 -1642 6852 -1620 sw
rect 6453 -1700 6468 -1692
rect 6534 -1664 6594 -1650
rect 6549 -1674 6594 -1664
rect 6549 -1692 6577 -1674
tri 6453 -1715 6468 -1700 ne
tri 6468 -1715 6490 -1693 sw
rect 6534 -1702 6577 -1692
rect 6592 -1678 6594 -1674
rect 6716 -1664 6776 -1650
tri 6830 -1655 6843 -1642 ne
rect 6843 -1648 6852 -1642
tri 6852 -1648 6858 -1642 sw
rect 6716 -1674 6761 -1664
rect 6592 -1702 6666 -1678
rect 6534 -1706 6666 -1702
tri 6666 -1706 6694 -1678 sw
rect 6716 -1688 6718 -1674
tri 6716 -1690 6718 -1688 ne
rect 6730 -1692 6761 -1674
rect 6730 -1702 6776 -1692
rect 6843 -1663 6858 -1648
tri 6468 -1727 6480 -1715 ne
rect 6480 -1720 6490 -1715
tri 6490 -1720 6495 -1715 sw
rect 6379 -2066 6394 -1838
rect 6480 -1876 6495 -1720
rect 6534 -1762 6562 -1706
tri 6654 -1724 6672 -1706 ne
rect 6672 -1726 6694 -1706
tri 6694 -1726 6714 -1706 sw
tri 6730 -1720 6748 -1702 ne
rect 6553 -1796 6562 -1762
rect 6596 -1735 6638 -1734
rect 6596 -1769 6601 -1735
rect 6631 -1769 6638 -1735
rect 6596 -1778 6638 -1769
rect 6672 -1735 6714 -1726
rect 6672 -1769 6679 -1735
rect 6709 -1769 6714 -1735
rect 6672 -1774 6714 -1769
rect 6748 -1762 6776 -1702
tri 6821 -1715 6843 -1693 se
rect 6843 -1700 6858 -1692
tri 6843 -1715 6858 -1700 nw
tri 6815 -1721 6821 -1715 se
rect 6821 -1721 6830 -1715
rect 6534 -1806 6562 -1796
tri 6562 -1806 6586 -1782 sw
rect 6534 -1838 6576 -1806
tri 6593 -1814 6594 -1813 sw
rect 6593 -1838 6594 -1814
tri 6596 -1815 6633 -1778 ne
rect 6633 -1806 6638 -1778
tri 6638 -1806 6664 -1780 sw
rect 6748 -1796 6757 -1762
rect 6748 -1806 6776 -1796
rect 6633 -1815 6717 -1806
tri 6633 -1834 6652 -1815 ne
rect 6652 -1834 6717 -1815
rect 6534 -1860 6594 -1838
rect 6716 -1838 6717 -1834
rect 6734 -1838 6776 -1806
rect 6716 -1860 6776 -1838
rect 6622 -1876 6639 -1862
rect 6671 -1876 6688 -1862
tri 6459 -1912 6481 -1890 se
rect 6481 -1897 6496 -1876
tri 6481 -1912 6496 -1897 nw
rect 6815 -1897 6830 -1721
tri 6830 -1728 6843 -1715 nw
rect 6916 -1796 6931 -1568
tri 6453 -1918 6459 -1912 se
rect 6459 -1918 6468 -1912
rect 6453 -1934 6468 -1918
tri 6468 -1925 6481 -1912 nw
rect 6622 -1920 6639 -1906
rect 6671 -1920 6688 -1906
tri 6815 -1912 6830 -1897 ne
tri 6830 -1912 6852 -1890 sw
rect 6453 -1970 6468 -1962
rect 6534 -1934 6594 -1920
rect 6549 -1944 6594 -1934
rect 6549 -1962 6577 -1944
tri 6453 -1985 6468 -1970 ne
tri 6468 -1985 6490 -1963 sw
rect 6534 -1972 6577 -1962
rect 6592 -1948 6594 -1944
rect 6716 -1934 6776 -1920
tri 6830 -1925 6843 -1912 ne
rect 6843 -1918 6852 -1912
tri 6852 -1918 6858 -1912 sw
rect 6716 -1944 6761 -1934
rect 6592 -1972 6666 -1948
rect 6534 -1976 6666 -1972
tri 6666 -1976 6694 -1948 sw
rect 6716 -1958 6718 -1944
tri 6716 -1960 6718 -1958 ne
rect 6730 -1962 6761 -1944
rect 6730 -1972 6776 -1962
rect 6843 -1933 6858 -1918
tri 6468 -1997 6480 -1985 ne
rect 6480 -1990 6490 -1985
tri 6490 -1990 6495 -1985 sw
rect 6379 -2146 6394 -2108
rect 6480 -2146 6495 -1990
rect 6534 -2032 6562 -1976
tri 6654 -1994 6672 -1976 ne
rect 6672 -1996 6694 -1976
tri 6694 -1996 6714 -1976 sw
tri 6730 -1990 6748 -1972 ne
rect 6553 -2066 6562 -2032
rect 6596 -2005 6638 -2004
rect 6596 -2039 6601 -2005
rect 6631 -2039 6638 -2005
rect 6596 -2048 6638 -2039
rect 6672 -2005 6714 -1996
rect 6672 -2039 6679 -2005
rect 6709 -2039 6714 -2005
rect 6672 -2044 6714 -2039
rect 6748 -2032 6776 -1972
tri 6821 -1985 6843 -1963 se
rect 6843 -1970 6858 -1962
tri 6843 -1985 6858 -1970 nw
tri 6815 -1991 6821 -1985 se
rect 6821 -1991 6830 -1985
rect 6534 -2076 6562 -2066
tri 6562 -2076 6586 -2052 sw
rect 6534 -2108 6576 -2076
tri 6593 -2084 6594 -2083 sw
rect 6593 -2108 6594 -2084
tri 6596 -2085 6633 -2048 ne
rect 6633 -2076 6638 -2048
tri 6638 -2076 6664 -2050 sw
rect 6748 -2066 6757 -2032
rect 6748 -2076 6776 -2066
rect 6633 -2085 6717 -2076
tri 6633 -2104 6652 -2085 ne
rect 6652 -2104 6717 -2085
rect 6534 -2130 6594 -2108
rect 6716 -2108 6717 -2104
rect 6734 -2108 6776 -2076
rect 6716 -2130 6776 -2108
rect 6622 -2146 6639 -2132
rect 6671 -2146 6688 -2132
rect 6815 -2146 6830 -1991
tri 6830 -1998 6843 -1985 nw
rect 6916 -2066 6931 -1838
rect 6916 -2146 6931 -2108
<< viali >>
rect 259 2130 291 2144
rect 42 2006 72 2040
rect 259 1904 291 1918
rect 478 2006 508 2040
rect 259 1860 291 1874
rect 42 1736 72 1770
rect 259 1634 291 1648
rect 478 1736 508 1770
rect 259 1590 291 1604
rect 42 1466 72 1500
rect 259 1364 291 1378
rect 478 1466 508 1500
rect 259 1320 291 1334
rect 42 1196 72 1230
rect 259 1094 291 1108
rect 478 1196 508 1230
rect 259 1050 291 1064
rect 42 926 72 960
rect 259 824 291 838
rect 478 926 508 960
rect 259 780 291 794
rect 42 656 72 690
rect 259 554 291 568
rect 478 656 508 690
rect 259 510 291 524
rect 42 386 72 420
rect 259 284 291 298
rect 478 386 508 420
rect 259 240 291 254
rect 42 116 72 150
rect 259 14 291 28
rect 478 116 508 150
rect 259 -30 291 -16
rect 42 -154 72 -120
rect 259 -256 291 -242
rect 478 -154 508 -120
rect 259 -300 291 -286
rect 42 -424 72 -390
rect 259 -526 291 -512
rect 478 -424 508 -390
rect 259 -570 291 -556
rect 42 -694 72 -660
rect 259 -796 291 -782
rect 478 -694 508 -660
rect 259 -840 291 -826
rect 42 -964 72 -930
rect 259 -1066 291 -1052
rect 478 -964 508 -930
rect 259 -1110 291 -1096
rect 42 -1234 72 -1200
rect 259 -1336 291 -1322
rect 478 -1234 508 -1200
rect 259 -1380 291 -1366
rect 42 -1504 72 -1470
rect 259 -1606 291 -1592
rect 478 -1504 508 -1470
rect 259 -1650 291 -1636
rect 42 -1774 72 -1740
rect 259 -1876 291 -1862
rect 478 -1774 508 -1740
rect 259 -1920 291 -1906
rect 42 -2044 72 -2010
rect 259 -2146 291 -2132
rect 478 -2044 508 -2010
rect 839 2130 871 2144
rect 622 2006 652 2040
rect 839 1904 871 1918
rect 1058 2006 1088 2040
rect 839 1860 871 1874
rect 622 1736 652 1770
rect 839 1634 871 1648
rect 1058 1736 1088 1770
rect 839 1590 871 1604
rect 622 1466 652 1500
rect 839 1364 871 1378
rect 1058 1466 1088 1500
rect 839 1320 871 1334
rect 622 1196 652 1230
rect 839 1094 871 1108
rect 1058 1196 1088 1230
rect 839 1050 871 1064
rect 622 926 652 960
rect 839 824 871 838
rect 1058 926 1088 960
rect 839 780 871 794
rect 622 656 652 690
rect 839 554 871 568
rect 1058 656 1088 690
rect 839 510 871 524
rect 622 386 652 420
rect 839 284 871 298
rect 1058 386 1088 420
rect 839 240 871 254
rect 622 116 652 150
rect 839 14 871 28
rect 1058 116 1088 150
rect 839 -30 871 -16
rect 622 -154 652 -120
rect 839 -256 871 -242
rect 1058 -154 1088 -120
rect 839 -300 871 -286
rect 622 -424 652 -390
rect 839 -526 871 -512
rect 1058 -424 1088 -390
rect 839 -570 871 -556
rect 622 -694 652 -660
rect 839 -796 871 -782
rect 1058 -694 1088 -660
rect 839 -840 871 -826
rect 622 -964 652 -930
rect 839 -1066 871 -1052
rect 1058 -964 1088 -930
rect 839 -1110 871 -1096
rect 622 -1234 652 -1200
rect 839 -1336 871 -1322
rect 1058 -1234 1088 -1200
rect 839 -1380 871 -1366
rect 622 -1504 652 -1470
rect 839 -1606 871 -1592
rect 1058 -1504 1088 -1470
rect 839 -1650 871 -1636
rect 622 -1774 652 -1740
rect 839 -1876 871 -1862
rect 1058 -1774 1088 -1740
rect 839 -1920 871 -1906
rect 622 -2044 652 -2010
rect 839 -2146 871 -2132
rect 1058 -2044 1088 -2010
rect 1419 2130 1451 2144
rect 1202 2006 1232 2040
rect 1419 1904 1451 1918
rect 1638 2006 1668 2040
rect 1419 1860 1451 1874
rect 1202 1736 1232 1770
rect 1419 1634 1451 1648
rect 1638 1736 1668 1770
rect 1419 1590 1451 1604
rect 1202 1466 1232 1500
rect 1419 1364 1451 1378
rect 1638 1466 1668 1500
rect 1419 1320 1451 1334
rect 1202 1196 1232 1230
rect 1419 1094 1451 1108
rect 1638 1196 1668 1230
rect 1419 1050 1451 1064
rect 1202 926 1232 960
rect 1419 824 1451 838
rect 1638 926 1668 960
rect 1419 780 1451 794
rect 1202 656 1232 690
rect 1419 554 1451 568
rect 1638 656 1668 690
rect 1419 510 1451 524
rect 1202 386 1232 420
rect 1419 284 1451 298
rect 1638 386 1668 420
rect 1419 240 1451 254
rect 1202 116 1232 150
rect 1419 14 1451 28
rect 1638 116 1668 150
rect 1419 -30 1451 -16
rect 1202 -154 1232 -120
rect 1419 -256 1451 -242
rect 1638 -154 1668 -120
rect 1419 -300 1451 -286
rect 1202 -424 1232 -390
rect 1419 -526 1451 -512
rect 1638 -424 1668 -390
rect 1419 -570 1451 -556
rect 1202 -694 1232 -660
rect 1419 -796 1451 -782
rect 1638 -694 1668 -660
rect 1419 -840 1451 -826
rect 1202 -964 1232 -930
rect 1419 -1066 1451 -1052
rect 1638 -964 1668 -930
rect 1419 -1110 1451 -1096
rect 1202 -1234 1232 -1200
rect 1419 -1336 1451 -1322
rect 1638 -1234 1668 -1200
rect 1419 -1380 1451 -1366
rect 1202 -1504 1232 -1470
rect 1419 -1606 1451 -1592
rect 1638 -1504 1668 -1470
rect 1419 -1650 1451 -1636
rect 1202 -1774 1232 -1740
rect 1419 -1876 1451 -1862
rect 1638 -1774 1668 -1740
rect 1419 -1920 1451 -1906
rect 1202 -2044 1232 -2010
rect 1419 -2146 1451 -2132
rect 1638 -2044 1668 -2010
rect 1999 2130 2031 2144
rect 1782 2006 1812 2040
rect 1999 1904 2031 1918
rect 2218 2006 2248 2040
rect 1999 1860 2031 1874
rect 1782 1736 1812 1770
rect 1999 1634 2031 1648
rect 2218 1736 2248 1770
rect 1999 1590 2031 1604
rect 1782 1466 1812 1500
rect 1999 1364 2031 1378
rect 2218 1466 2248 1500
rect 1999 1320 2031 1334
rect 1782 1196 1812 1230
rect 1999 1094 2031 1108
rect 2218 1196 2248 1230
rect 1999 1050 2031 1064
rect 1782 926 1812 960
rect 1999 824 2031 838
rect 2218 926 2248 960
rect 1999 780 2031 794
rect 1782 656 1812 690
rect 1999 554 2031 568
rect 2218 656 2248 690
rect 1999 510 2031 524
rect 1782 386 1812 420
rect 1999 284 2031 298
rect 2218 386 2248 420
rect 1999 240 2031 254
rect 1782 116 1812 150
rect 1999 14 2031 28
rect 2218 116 2248 150
rect 1999 -30 2031 -16
rect 1782 -154 1812 -120
rect 1999 -256 2031 -242
rect 2218 -154 2248 -120
rect 1999 -300 2031 -286
rect 1782 -424 1812 -390
rect 1999 -526 2031 -512
rect 2218 -424 2248 -390
rect 1999 -570 2031 -556
rect 1782 -694 1812 -660
rect 1999 -796 2031 -782
rect 2218 -694 2248 -660
rect 1999 -840 2031 -826
rect 1782 -964 1812 -930
rect 1999 -1066 2031 -1052
rect 2218 -964 2248 -930
rect 1999 -1110 2031 -1096
rect 1782 -1234 1812 -1200
rect 1999 -1336 2031 -1322
rect 2218 -1234 2248 -1200
rect 1999 -1380 2031 -1366
rect 1782 -1504 1812 -1470
rect 1999 -1606 2031 -1592
rect 2218 -1504 2248 -1470
rect 1999 -1650 2031 -1636
rect 1782 -1774 1812 -1740
rect 1999 -1876 2031 -1862
rect 2218 -1774 2248 -1740
rect 1999 -1920 2031 -1906
rect 1782 -2044 1812 -2010
rect 1999 -2146 2031 -2132
rect 2218 -2044 2248 -2010
rect 2579 2130 2611 2144
rect 2362 2006 2392 2040
rect 2579 1904 2611 1918
rect 2798 2006 2828 2040
rect 2579 1860 2611 1874
rect 2362 1736 2392 1770
rect 2579 1634 2611 1648
rect 2798 1736 2828 1770
rect 2579 1590 2611 1604
rect 2362 1466 2392 1500
rect 2579 1364 2611 1378
rect 2798 1466 2828 1500
rect 2579 1320 2611 1334
rect 2362 1196 2392 1230
rect 2579 1094 2611 1108
rect 2798 1196 2828 1230
rect 2579 1050 2611 1064
rect 2362 926 2392 960
rect 2579 824 2611 838
rect 2798 926 2828 960
rect 2579 780 2611 794
rect 2362 656 2392 690
rect 2579 554 2611 568
rect 2798 656 2828 690
rect 2579 510 2611 524
rect 2362 386 2392 420
rect 2579 284 2611 298
rect 2798 386 2828 420
rect 2579 240 2611 254
rect 2362 116 2392 150
rect 2579 14 2611 28
rect 2798 116 2828 150
rect 2579 -30 2611 -16
rect 2362 -154 2392 -120
rect 2579 -256 2611 -242
rect 2798 -154 2828 -120
rect 2579 -300 2611 -286
rect 2362 -424 2392 -390
rect 2579 -526 2611 -512
rect 2798 -424 2828 -390
rect 2579 -570 2611 -556
rect 2362 -694 2392 -660
rect 2579 -796 2611 -782
rect 2798 -694 2828 -660
rect 2579 -840 2611 -826
rect 2362 -964 2392 -930
rect 2579 -1066 2611 -1052
rect 2798 -964 2828 -930
rect 2579 -1110 2611 -1096
rect 2362 -1234 2392 -1200
rect 2579 -1336 2611 -1322
rect 2798 -1234 2828 -1200
rect 2579 -1380 2611 -1366
rect 2362 -1504 2392 -1470
rect 2579 -1606 2611 -1592
rect 2798 -1504 2828 -1470
rect 2579 -1650 2611 -1636
rect 2362 -1774 2392 -1740
rect 2579 -1876 2611 -1862
rect 2798 -1774 2828 -1740
rect 2579 -1920 2611 -1906
rect 2362 -2044 2392 -2010
rect 2579 -2146 2611 -2132
rect 2798 -2044 2828 -2010
rect 3159 2130 3191 2144
rect 2942 2006 2972 2040
rect 3159 1904 3191 1918
rect 3378 2006 3408 2040
rect 3159 1860 3191 1874
rect 2942 1736 2972 1770
rect 3159 1634 3191 1648
rect 3378 1736 3408 1770
rect 3159 1590 3191 1604
rect 2942 1466 2972 1500
rect 3159 1364 3191 1378
rect 3378 1466 3408 1500
rect 3159 1320 3191 1334
rect 2942 1196 2972 1230
rect 3159 1094 3191 1108
rect 3378 1196 3408 1230
rect 3159 1050 3191 1064
rect 2942 926 2972 960
rect 3159 824 3191 838
rect 3378 926 3408 960
rect 3159 780 3191 794
rect 2942 656 2972 690
rect 3159 554 3191 568
rect 3378 656 3408 690
rect 3159 510 3191 524
rect 2942 386 2972 420
rect 3159 284 3191 298
rect 3378 386 3408 420
rect 3159 240 3191 254
rect 2942 116 2972 150
rect 3159 14 3191 28
rect 3378 116 3408 150
rect 3159 -30 3191 -16
rect 2942 -154 2972 -120
rect 3159 -256 3191 -242
rect 3378 -154 3408 -120
rect 3159 -300 3191 -286
rect 2942 -424 2972 -390
rect 3159 -526 3191 -512
rect 3378 -424 3408 -390
rect 3159 -570 3191 -556
rect 2942 -694 2972 -660
rect 3159 -796 3191 -782
rect 3378 -694 3408 -660
rect 3159 -840 3191 -826
rect 2942 -964 2972 -930
rect 3159 -1066 3191 -1052
rect 3378 -964 3408 -930
rect 3159 -1110 3191 -1096
rect 2942 -1234 2972 -1200
rect 3159 -1336 3191 -1322
rect 3378 -1234 3408 -1200
rect 3159 -1380 3191 -1366
rect 2942 -1504 2972 -1470
rect 3159 -1606 3191 -1592
rect 3378 -1504 3408 -1470
rect 3159 -1650 3191 -1636
rect 2942 -1774 2972 -1740
rect 3159 -1876 3191 -1862
rect 3378 -1774 3408 -1740
rect 3159 -1920 3191 -1906
rect 2942 -2044 2972 -2010
rect 3159 -2146 3191 -2132
rect 3378 -2044 3408 -2010
rect 3739 2130 3771 2144
rect 3522 2006 3552 2040
rect 3739 1904 3771 1918
rect 3958 2006 3988 2040
rect 3739 1860 3771 1874
rect 3522 1736 3552 1770
rect 3739 1634 3771 1648
rect 3958 1736 3988 1770
rect 3739 1590 3771 1604
rect 3522 1466 3552 1500
rect 3739 1364 3771 1378
rect 3958 1466 3988 1500
rect 3739 1320 3771 1334
rect 3522 1196 3552 1230
rect 3739 1094 3771 1108
rect 3958 1196 3988 1230
rect 3739 1050 3771 1064
rect 3522 926 3552 960
rect 3739 824 3771 838
rect 3958 926 3988 960
rect 3739 780 3771 794
rect 3522 656 3552 690
rect 3739 554 3771 568
rect 3958 656 3988 690
rect 3739 510 3771 524
rect 3522 386 3552 420
rect 3739 284 3771 298
rect 3958 386 3988 420
rect 3739 240 3771 254
rect 3522 116 3552 150
rect 3739 14 3771 28
rect 3958 116 3988 150
rect 3739 -30 3771 -16
rect 3522 -154 3552 -120
rect 3739 -256 3771 -242
rect 3958 -154 3988 -120
rect 3739 -300 3771 -286
rect 3522 -424 3552 -390
rect 3739 -526 3771 -512
rect 3958 -424 3988 -390
rect 3739 -570 3771 -556
rect 3522 -694 3552 -660
rect 3739 -796 3771 -782
rect 3958 -694 3988 -660
rect 3739 -840 3771 -826
rect 3522 -964 3552 -930
rect 3739 -1066 3771 -1052
rect 3958 -964 3988 -930
rect 3739 -1110 3771 -1096
rect 3522 -1234 3552 -1200
rect 3739 -1336 3771 -1322
rect 3958 -1234 3988 -1200
rect 3739 -1380 3771 -1366
rect 3522 -1504 3552 -1470
rect 3739 -1606 3771 -1592
rect 3958 -1504 3988 -1470
rect 3739 -1650 3771 -1636
rect 3522 -1774 3552 -1740
rect 3739 -1876 3771 -1862
rect 3958 -1774 3988 -1740
rect 3739 -1920 3771 -1906
rect 3522 -2044 3552 -2010
rect 3739 -2146 3771 -2132
rect 3958 -2044 3988 -2010
rect 4319 2130 4351 2144
rect 4102 2006 4132 2040
rect 4319 1904 4351 1918
rect 4538 2006 4568 2040
rect 4319 1860 4351 1874
rect 4102 1736 4132 1770
rect 4319 1634 4351 1648
rect 4538 1736 4568 1770
rect 4319 1590 4351 1604
rect 4102 1466 4132 1500
rect 4319 1364 4351 1378
rect 4538 1466 4568 1500
rect 4319 1320 4351 1334
rect 4102 1196 4132 1230
rect 4319 1094 4351 1108
rect 4538 1196 4568 1230
rect 4319 1050 4351 1064
rect 4102 926 4132 960
rect 4319 824 4351 838
rect 4538 926 4568 960
rect 4319 780 4351 794
rect 4102 656 4132 690
rect 4319 554 4351 568
rect 4538 656 4568 690
rect 4319 510 4351 524
rect 4102 386 4132 420
rect 4319 284 4351 298
rect 4538 386 4568 420
rect 4319 240 4351 254
rect 4102 116 4132 150
rect 4319 14 4351 28
rect 4538 116 4568 150
rect 4319 -30 4351 -16
rect 4102 -154 4132 -120
rect 4319 -256 4351 -242
rect 4538 -154 4568 -120
rect 4319 -300 4351 -286
rect 4102 -424 4132 -390
rect 4319 -526 4351 -512
rect 4538 -424 4568 -390
rect 4319 -570 4351 -556
rect 4102 -694 4132 -660
rect 4319 -796 4351 -782
rect 4538 -694 4568 -660
rect 4319 -840 4351 -826
rect 4102 -964 4132 -930
rect 4319 -1066 4351 -1052
rect 4538 -964 4568 -930
rect 4319 -1110 4351 -1096
rect 4102 -1234 4132 -1200
rect 4319 -1336 4351 -1322
rect 4538 -1234 4568 -1200
rect 4319 -1380 4351 -1366
rect 4102 -1504 4132 -1470
rect 4319 -1606 4351 -1592
rect 4538 -1504 4568 -1470
rect 4319 -1650 4351 -1636
rect 4102 -1774 4132 -1740
rect 4319 -1876 4351 -1862
rect 4538 -1774 4568 -1740
rect 4319 -1920 4351 -1906
rect 4102 -2044 4132 -2010
rect 4319 -2146 4351 -2132
rect 4538 -2044 4568 -2010
rect 4899 2130 4931 2144
rect 4682 2006 4712 2040
rect 4899 1904 4931 1918
rect 5118 2006 5148 2040
rect 4899 1860 4931 1874
rect 4682 1736 4712 1770
rect 4899 1634 4931 1648
rect 5118 1736 5148 1770
rect 4899 1590 4931 1604
rect 4682 1466 4712 1500
rect 4899 1364 4931 1378
rect 5118 1466 5148 1500
rect 4899 1320 4931 1334
rect 4682 1196 4712 1230
rect 4899 1094 4931 1108
rect 5118 1196 5148 1230
rect 4899 1050 4931 1064
rect 4682 926 4712 960
rect 4899 824 4931 838
rect 5118 926 5148 960
rect 4899 780 4931 794
rect 4682 656 4712 690
rect 4899 554 4931 568
rect 5118 656 5148 690
rect 4899 510 4931 524
rect 4682 386 4712 420
rect 4899 284 4931 298
rect 5118 386 5148 420
rect 4899 240 4931 254
rect 4682 116 4712 150
rect 4899 14 4931 28
rect 5118 116 5148 150
rect 4899 -30 4931 -16
rect 4682 -154 4712 -120
rect 4899 -256 4931 -242
rect 5118 -154 5148 -120
rect 4899 -300 4931 -286
rect 4682 -424 4712 -390
rect 4899 -526 4931 -512
rect 5118 -424 5148 -390
rect 4899 -570 4931 -556
rect 4682 -694 4712 -660
rect 4899 -796 4931 -782
rect 5118 -694 5148 -660
rect 4899 -840 4931 -826
rect 4682 -964 4712 -930
rect 4899 -1066 4931 -1052
rect 5118 -964 5148 -930
rect 4899 -1110 4931 -1096
rect 4682 -1234 4712 -1200
rect 4899 -1336 4931 -1322
rect 5118 -1234 5148 -1200
rect 4899 -1380 4931 -1366
rect 4682 -1504 4712 -1470
rect 4899 -1606 4931 -1592
rect 5118 -1504 5148 -1470
rect 4899 -1650 4931 -1636
rect 4682 -1774 4712 -1740
rect 4899 -1876 4931 -1862
rect 5118 -1774 5148 -1740
rect 4899 -1920 4931 -1906
rect 4682 -2044 4712 -2010
rect 4899 -2146 4931 -2132
rect 5118 -2044 5148 -2010
rect 5479 2130 5511 2144
rect 5262 2006 5292 2040
rect 5479 1904 5511 1918
rect 5698 2006 5728 2040
rect 5479 1860 5511 1874
rect 5262 1736 5292 1770
rect 5479 1634 5511 1648
rect 5698 1736 5728 1770
rect 5479 1590 5511 1604
rect 5262 1466 5292 1500
rect 5479 1364 5511 1378
rect 5698 1466 5728 1500
rect 5479 1320 5511 1334
rect 5262 1196 5292 1230
rect 5479 1094 5511 1108
rect 5698 1196 5728 1230
rect 5479 1050 5511 1064
rect 5262 926 5292 960
rect 5479 824 5511 838
rect 5698 926 5728 960
rect 5479 780 5511 794
rect 5262 656 5292 690
rect 5479 554 5511 568
rect 5698 656 5728 690
rect 5479 510 5511 524
rect 5262 386 5292 420
rect 5479 284 5511 298
rect 5698 386 5728 420
rect 5479 240 5511 254
rect 5262 116 5292 150
rect 5479 14 5511 28
rect 5698 116 5728 150
rect 5479 -30 5511 -16
rect 5262 -154 5292 -120
rect 5479 -256 5511 -242
rect 5698 -154 5728 -120
rect 5479 -300 5511 -286
rect 5262 -424 5292 -390
rect 5479 -526 5511 -512
rect 5698 -424 5728 -390
rect 5479 -570 5511 -556
rect 5262 -694 5292 -660
rect 5479 -796 5511 -782
rect 5698 -694 5728 -660
rect 5479 -840 5511 -826
rect 5262 -964 5292 -930
rect 5479 -1066 5511 -1052
rect 5698 -964 5728 -930
rect 5479 -1110 5511 -1096
rect 5262 -1234 5292 -1200
rect 5479 -1336 5511 -1322
rect 5698 -1234 5728 -1200
rect 5479 -1380 5511 -1366
rect 5262 -1504 5292 -1470
rect 5479 -1606 5511 -1592
rect 5698 -1504 5728 -1470
rect 5479 -1650 5511 -1636
rect 5262 -1774 5292 -1740
rect 5479 -1876 5511 -1862
rect 5698 -1774 5728 -1740
rect 5479 -1920 5511 -1906
rect 5262 -2044 5292 -2010
rect 5479 -2146 5511 -2132
rect 5698 -2044 5728 -2010
rect 6059 2130 6091 2144
rect 5842 2006 5872 2040
rect 6059 1904 6091 1918
rect 6278 2006 6308 2040
rect 6059 1860 6091 1874
rect 5842 1736 5872 1770
rect 6059 1634 6091 1648
rect 6278 1736 6308 1770
rect 6059 1590 6091 1604
rect 5842 1466 5872 1500
rect 6059 1364 6091 1378
rect 6278 1466 6308 1500
rect 6059 1320 6091 1334
rect 5842 1196 5872 1230
rect 6059 1094 6091 1108
rect 6278 1196 6308 1230
rect 6059 1050 6091 1064
rect 5842 926 5872 960
rect 6059 824 6091 838
rect 6278 926 6308 960
rect 6059 780 6091 794
rect 5842 656 5872 690
rect 6059 554 6091 568
rect 6278 656 6308 690
rect 6059 510 6091 524
rect 5842 386 5872 420
rect 6059 284 6091 298
rect 6278 386 6308 420
rect 6059 240 6091 254
rect 5842 116 5872 150
rect 6059 14 6091 28
rect 6278 116 6308 150
rect 6059 -30 6091 -16
rect 5842 -154 5872 -120
rect 6059 -256 6091 -242
rect 6278 -154 6308 -120
rect 6059 -300 6091 -286
rect 5842 -424 5872 -390
rect 6059 -526 6091 -512
rect 6278 -424 6308 -390
rect 6059 -570 6091 -556
rect 5842 -694 5872 -660
rect 6059 -796 6091 -782
rect 6278 -694 6308 -660
rect 6059 -840 6091 -826
rect 5842 -964 5872 -930
rect 6059 -1066 6091 -1052
rect 6278 -964 6308 -930
rect 6059 -1110 6091 -1096
rect 5842 -1234 5872 -1200
rect 6059 -1336 6091 -1322
rect 6278 -1234 6308 -1200
rect 6059 -1380 6091 -1366
rect 5842 -1504 5872 -1470
rect 6059 -1606 6091 -1592
rect 6278 -1504 6308 -1470
rect 6059 -1650 6091 -1636
rect 5842 -1774 5872 -1740
rect 6059 -1876 6091 -1862
rect 6278 -1774 6308 -1740
rect 6059 -1920 6091 -1906
rect 5842 -2044 5872 -2010
rect 6059 -2146 6091 -2132
rect 6278 -2044 6308 -2010
rect 6639 2130 6671 2144
rect 6422 2006 6452 2040
rect 6639 1904 6671 1918
rect 6858 2006 6888 2040
rect 6639 1860 6671 1874
rect 6422 1736 6452 1770
rect 6639 1634 6671 1648
rect 6858 1736 6888 1770
rect 6639 1590 6671 1604
rect 6422 1466 6452 1500
rect 6639 1364 6671 1378
rect 6858 1466 6888 1500
rect 6639 1320 6671 1334
rect 6422 1196 6452 1230
rect 6639 1094 6671 1108
rect 6858 1196 6888 1230
rect 6639 1050 6671 1064
rect 6422 926 6452 960
rect 6639 824 6671 838
rect 6858 926 6888 960
rect 6639 780 6671 794
rect 6422 656 6452 690
rect 6639 554 6671 568
rect 6858 656 6888 690
rect 6639 510 6671 524
rect 6422 386 6452 420
rect 6639 284 6671 298
rect 6858 386 6888 420
rect 6639 240 6671 254
rect 6422 116 6452 150
rect 6639 14 6671 28
rect 6858 116 6888 150
rect 6639 -30 6671 -16
rect 6422 -154 6452 -120
rect 6639 -256 6671 -242
rect 6858 -154 6888 -120
rect 6639 -300 6671 -286
rect 6422 -424 6452 -390
rect 6639 -526 6671 -512
rect 6858 -424 6888 -390
rect 6639 -570 6671 -556
rect 6422 -694 6452 -660
rect 6639 -796 6671 -782
rect 6858 -694 6888 -660
rect 6639 -840 6671 -826
rect 6422 -964 6452 -930
rect 6639 -1066 6671 -1052
rect 6858 -964 6888 -930
rect 6639 -1110 6671 -1096
rect 6422 -1234 6452 -1200
rect 6639 -1336 6671 -1322
rect 6858 -1234 6888 -1200
rect 6639 -1380 6671 -1366
rect 6422 -1504 6452 -1470
rect 6639 -1606 6671 -1592
rect 6858 -1504 6888 -1470
rect 6639 -1650 6671 -1636
rect 6422 -1774 6452 -1740
rect 6639 -1876 6671 -1862
rect 6858 -1774 6888 -1740
rect 6639 -1920 6671 -1906
rect 6422 -2044 6452 -2010
rect 6639 -2146 6671 -2132
rect 6858 -2044 6888 -2010
<< metal1 >>
rect -1 2130 259 2144
rect 291 2130 839 2144
rect 871 2130 1419 2144
rect 1451 2130 1999 2144
rect 2031 2130 2579 2144
rect 2611 2130 3159 2144
rect 3191 2130 3739 2144
rect 3771 2130 4319 2144
rect 4351 2130 4899 2144
rect 4931 2130 5479 2144
rect 5511 2130 6059 2144
rect 6091 2130 6639 2144
rect 6671 2130 6931 2144
rect -1 2006 42 2040
rect 72 2006 478 2040
rect 508 2006 622 2040
rect 652 2006 1058 2040
rect 1088 2006 1202 2040
rect 1232 2006 1638 2040
rect 1668 2006 1782 2040
rect 1812 2006 2218 2040
rect 2248 2006 2362 2040
rect 2392 2006 2798 2040
rect 2828 2006 2942 2040
rect 2972 2006 3378 2040
rect 3408 2006 3522 2040
rect 3552 2006 3958 2040
rect 3988 2006 4102 2040
rect 4132 2006 4538 2040
rect 4568 2006 4682 2040
rect 4712 2006 5118 2040
rect 5148 2006 5262 2040
rect 5292 2006 5698 2040
rect 5728 2006 5842 2040
rect 5872 2006 6278 2040
rect 6308 2006 6422 2040
rect 6452 2006 6858 2040
rect 6888 2006 6931 2040
rect -1 1904 259 1918
rect 291 1904 839 1918
rect 871 1904 1419 1918
rect 1451 1904 1999 1918
rect 2031 1904 2579 1918
rect 2611 1904 3159 1918
rect 3191 1904 3739 1918
rect 3771 1904 4319 1918
rect 4351 1904 4899 1918
rect 4931 1904 5479 1918
rect 5511 1904 6059 1918
rect 6091 1904 6639 1918
rect 6671 1904 6931 1918
rect -1 1860 259 1874
rect 291 1860 839 1874
rect 871 1860 1419 1874
rect 1451 1860 1999 1874
rect 2031 1860 2579 1874
rect 2611 1860 3159 1874
rect 3191 1860 3739 1874
rect 3771 1860 4319 1874
rect 4351 1860 4899 1874
rect 4931 1860 5479 1874
rect 5511 1860 6059 1874
rect 6091 1860 6639 1874
rect 6671 1860 6931 1874
rect -1 1736 42 1770
rect 72 1736 478 1770
rect 508 1736 622 1770
rect 652 1736 1058 1770
rect 1088 1736 1202 1770
rect 1232 1736 1638 1770
rect 1668 1736 1782 1770
rect 1812 1736 2218 1770
rect 2248 1736 2362 1770
rect 2392 1736 2798 1770
rect 2828 1736 2942 1770
rect 2972 1736 3378 1770
rect 3408 1736 3522 1770
rect 3552 1736 3958 1770
rect 3988 1736 4102 1770
rect 4132 1736 4538 1770
rect 4568 1736 4682 1770
rect 4712 1736 5118 1770
rect 5148 1736 5262 1770
rect 5292 1736 5698 1770
rect 5728 1736 5842 1770
rect 5872 1736 6278 1770
rect 6308 1736 6422 1770
rect 6452 1736 6858 1770
rect 6888 1736 6931 1770
rect -1 1634 259 1648
rect 291 1634 839 1648
rect 871 1634 1419 1648
rect 1451 1634 1999 1648
rect 2031 1634 2579 1648
rect 2611 1634 3159 1648
rect 3191 1634 3739 1648
rect 3771 1634 4319 1648
rect 4351 1634 4899 1648
rect 4931 1634 5479 1648
rect 5511 1634 6059 1648
rect 6091 1634 6639 1648
rect 6671 1634 6931 1648
rect -1 1590 259 1604
rect 291 1590 839 1604
rect 871 1590 1419 1604
rect 1451 1590 1999 1604
rect 2031 1590 2579 1604
rect 2611 1590 3159 1604
rect 3191 1590 3739 1604
rect 3771 1590 4319 1604
rect 4351 1590 4899 1604
rect 4931 1590 5479 1604
rect 5511 1590 6059 1604
rect 6091 1590 6639 1604
rect 6671 1590 6931 1604
rect -1 1466 42 1500
rect 72 1466 478 1500
rect 508 1466 622 1500
rect 652 1466 1058 1500
rect 1088 1466 1202 1500
rect 1232 1466 1638 1500
rect 1668 1466 1782 1500
rect 1812 1466 2218 1500
rect 2248 1466 2362 1500
rect 2392 1466 2798 1500
rect 2828 1466 2942 1500
rect 2972 1466 3378 1500
rect 3408 1466 3522 1500
rect 3552 1466 3958 1500
rect 3988 1466 4102 1500
rect 4132 1466 4538 1500
rect 4591 1466 4682 1500
rect 4712 1466 5118 1500
rect 5148 1466 5262 1500
rect 5292 1466 5698 1500
rect 5728 1466 5842 1500
rect 5872 1466 6278 1500
rect 6308 1466 6422 1500
rect 6452 1466 6858 1500
rect 6888 1466 6931 1500
rect -1 1364 259 1378
rect 291 1364 839 1378
rect 871 1364 1419 1378
rect 1451 1364 1999 1378
rect 2031 1364 2579 1378
rect 2611 1364 3159 1378
rect 3191 1364 3739 1378
rect 3771 1364 4319 1378
rect 4351 1364 4899 1378
rect 4931 1364 5479 1378
rect 5511 1364 6059 1378
rect 6091 1364 6639 1378
rect 6671 1364 6931 1378
rect -1 1320 259 1334
rect 291 1320 839 1334
rect 871 1320 1419 1334
rect 1451 1320 1999 1334
rect 2031 1320 2579 1334
rect 2611 1320 3159 1334
rect 3191 1320 3739 1334
rect 3771 1320 4319 1334
rect 4351 1320 4899 1334
rect 4931 1320 5479 1334
rect 5511 1320 6059 1334
rect 6091 1320 6639 1334
rect 6671 1320 6931 1334
rect -1 1196 42 1230
rect 72 1196 478 1230
rect 508 1196 622 1230
rect 652 1196 1058 1230
rect 1088 1196 1202 1230
rect 1232 1196 1638 1230
rect 1668 1196 1782 1230
rect 1812 1196 2218 1230
rect 2248 1196 2362 1230
rect 2392 1196 2798 1230
rect 2828 1196 2942 1230
rect 2972 1196 3378 1230
rect 3408 1196 3522 1230
rect 3552 1196 3958 1230
rect 3988 1196 4102 1230
rect 4132 1196 4538 1230
rect 4591 1196 4682 1230
rect 4712 1196 5118 1230
rect 5148 1196 5262 1230
rect 5292 1196 5698 1230
rect 5728 1196 5842 1230
rect 5872 1196 6278 1230
rect 6308 1196 6422 1230
rect 6452 1196 6858 1230
rect 6888 1196 6931 1230
rect -1 1094 259 1108
rect 291 1094 839 1108
rect 871 1094 1419 1108
rect 1451 1094 1999 1108
rect 2031 1094 2579 1108
rect 2611 1094 3159 1108
rect 3191 1094 3739 1108
rect 3771 1094 4319 1108
rect 4351 1094 4899 1108
rect 4931 1094 5479 1108
rect 5511 1094 6059 1108
rect 6091 1094 6639 1108
rect 6671 1094 6931 1108
rect -1 1050 259 1064
rect 291 1050 839 1064
rect 871 1050 1419 1064
rect 1451 1050 1999 1064
rect 2031 1050 2579 1064
rect 2611 1050 3159 1064
rect 3191 1050 3739 1064
rect 3771 1050 4319 1064
rect 4351 1050 4899 1064
rect 4931 1050 5479 1064
rect 5511 1050 6059 1064
rect 6091 1050 6639 1064
rect 6671 1050 6931 1064
rect -1 926 42 960
rect 72 926 478 960
rect 508 926 622 960
rect 652 926 1058 960
rect 1088 926 1202 960
rect 1232 926 1638 960
rect 1668 926 1782 960
rect 1812 926 2218 960
rect 2248 926 2362 960
rect 2392 926 2798 960
rect 2828 926 2942 960
rect 2972 926 3378 960
rect 3408 926 3522 960
rect 3552 926 3958 960
rect 3988 926 4102 960
rect 4132 926 4538 960
rect 4591 926 4682 960
rect 4712 926 5118 960
rect 5148 926 5262 960
rect 5292 926 5698 960
rect 5728 926 5842 960
rect 5872 926 6278 960
rect 6308 926 6422 960
rect 6452 926 6858 960
rect 6888 926 6931 960
rect -1 824 259 838
rect 291 824 839 838
rect 871 824 1419 838
rect 1451 824 1999 838
rect 2031 824 2579 838
rect 2611 824 3159 838
rect 3191 824 3739 838
rect 3771 824 4319 838
rect 4351 824 4899 838
rect 4931 824 5479 838
rect 5511 824 6059 838
rect 6091 824 6639 838
rect 6671 824 6931 838
rect -1 780 259 794
rect 291 780 839 794
rect 871 780 1419 794
rect 1451 780 1999 794
rect 2031 780 2579 794
rect 2611 780 3159 794
rect 3191 780 3739 794
rect 3771 780 4319 794
rect 4351 780 4899 794
rect 4931 780 5479 794
rect 5511 780 6059 794
rect 6091 780 6639 794
rect 6671 780 6931 794
rect -1 656 42 690
rect 72 656 478 690
rect 508 656 622 690
rect 652 656 1058 690
rect 1088 656 1202 690
rect 1232 656 1638 690
rect 1668 656 1782 690
rect 1812 656 2218 690
rect 2248 656 2362 690
rect 2392 656 2798 690
rect 2828 656 2942 690
rect 2972 656 3378 690
rect 3408 656 3522 690
rect 3552 656 3958 690
rect 3988 656 4102 690
rect 4132 656 4538 690
rect 4591 656 4682 690
rect 4712 656 5118 690
rect 5148 656 5262 690
rect 5292 656 5698 690
rect 5728 656 5842 690
rect 5872 656 6278 690
rect 6308 656 6422 690
rect 6452 656 6858 690
rect 6888 656 6931 690
rect -1 554 259 568
rect 291 554 839 568
rect 871 554 1419 568
rect 1451 554 1999 568
rect 2031 554 2579 568
rect 2611 554 3159 568
rect 3191 554 3739 568
rect 3771 554 4319 568
rect 4351 554 4899 568
rect 4931 554 5479 568
rect 5511 554 6059 568
rect 6091 554 6639 568
rect 6671 554 6931 568
rect -1 510 259 524
rect 291 510 839 524
rect 871 510 1419 524
rect 1451 510 1999 524
rect 2031 510 2579 524
rect 2611 510 3159 524
rect 3191 510 3739 524
rect 3771 510 4319 524
rect 4351 510 4899 524
rect 4931 510 5479 524
rect 5511 510 6059 524
rect 6091 510 6639 524
rect 6671 510 6931 524
rect -1 386 42 420
rect 72 386 478 420
rect 508 386 622 420
rect 652 386 1058 420
rect 1088 386 1202 420
rect 1232 386 1638 420
rect 1668 386 1782 420
rect 1812 386 2218 420
rect 2248 386 2362 420
rect 2392 386 2798 420
rect 2828 386 2942 420
rect 2972 386 3378 420
rect 3408 386 3522 420
rect 3552 386 3958 420
rect 3988 386 4102 420
rect 4132 386 4538 420
rect 4591 386 4682 420
rect 4712 386 5118 420
rect 5148 386 5262 420
rect 5292 386 5698 420
rect 5728 386 5842 420
rect 5872 386 6278 420
rect 6308 386 6422 420
rect 6452 386 6858 420
rect 6888 386 6931 420
rect -1 284 259 298
rect 291 284 839 298
rect 871 284 1419 298
rect 1451 284 1999 298
rect 2031 284 2579 298
rect 2611 284 3159 298
rect 3191 284 3739 298
rect 3771 284 4319 298
rect 4351 284 4899 298
rect 4931 284 5479 298
rect 5511 284 6059 298
rect 6091 284 6639 298
rect 6671 284 6931 298
rect -1 240 259 254
rect 291 240 839 254
rect 871 240 1419 254
rect 1451 240 1999 254
rect 2031 240 2579 254
rect 2611 240 3159 254
rect 3191 240 3739 254
rect 3771 240 4319 254
rect 4351 240 4899 254
rect 4931 240 5479 254
rect 5511 240 6059 254
rect 6091 240 6639 254
rect 6671 240 6931 254
rect -1 116 42 150
rect 72 116 478 150
rect 508 116 622 150
rect 652 116 1058 150
rect 1088 116 1202 150
rect 1232 116 1638 150
rect 1668 116 1782 150
rect 1812 116 2218 150
rect 2248 116 2362 150
rect 2392 116 2798 150
rect 2828 116 2942 150
rect 2972 116 3378 150
rect 3408 116 3522 150
rect 3552 116 3958 150
rect 3988 116 4102 150
rect 4132 116 4538 150
rect 4591 116 4682 150
rect 4712 116 5118 150
rect 5148 116 5262 150
rect 5292 116 5698 150
rect 5728 116 5842 150
rect 5872 116 6278 150
rect 6308 116 6422 150
rect 6452 116 6858 150
rect 6888 116 6931 150
rect -1 14 259 28
rect 291 14 839 28
rect 871 14 1419 28
rect 1451 14 1999 28
rect 2031 14 2579 28
rect 2611 14 3159 28
rect 3191 14 3739 28
rect 3771 14 4319 28
rect 4351 14 4899 28
rect 4931 14 5479 28
rect 5511 14 6059 28
rect 6091 14 6639 28
rect 6671 14 6931 28
rect -1 -30 259 -16
rect 291 -30 839 -16
rect 871 -30 1419 -16
rect 1451 -30 1999 -16
rect 2031 -30 2579 -16
rect 2611 -30 3159 -16
rect 3191 -30 3739 -16
rect 3771 -30 4319 -16
rect 4351 -30 4899 -16
rect 4931 -30 5479 -16
rect 5511 -30 6059 -16
rect 6091 -30 6639 -16
rect 6671 -30 6931 -16
rect -1 -154 42 -120
rect 72 -154 478 -120
rect 508 -154 622 -120
rect 652 -154 1058 -120
rect 1088 -154 1202 -120
rect 1232 -154 1638 -120
rect 1668 -154 1782 -120
rect 1812 -154 2218 -120
rect 2248 -154 2362 -120
rect 2392 -154 2798 -120
rect 2828 -154 2942 -120
rect 2972 -154 3378 -120
rect 3408 -154 3522 -120
rect 3552 -154 3958 -120
rect 3988 -154 4102 -120
rect 4132 -154 4538 -120
rect 4591 -154 4682 -120
rect 4712 -154 5118 -120
rect 5148 -154 5262 -120
rect 5292 -154 5698 -120
rect 5728 -154 5842 -120
rect 5872 -154 6278 -120
rect 6308 -154 6422 -120
rect 6452 -154 6858 -120
rect 6888 -154 6931 -120
rect -1 -256 259 -242
rect 291 -256 839 -242
rect 871 -256 1419 -242
rect 1451 -256 1999 -242
rect 2031 -256 2579 -242
rect 2611 -256 3159 -242
rect 3191 -256 3739 -242
rect 3771 -256 4319 -242
rect 4351 -256 4899 -242
rect 4931 -256 5479 -242
rect 5511 -256 6059 -242
rect 6091 -256 6639 -242
rect 6671 -256 6931 -242
rect -1 -300 259 -286
rect 291 -300 839 -286
rect 871 -300 1419 -286
rect 1451 -300 1999 -286
rect 2031 -300 2579 -286
rect 2611 -300 3159 -286
rect 3191 -300 3739 -286
rect 3771 -300 4319 -286
rect 4351 -300 4899 -286
rect 4931 -300 5479 -286
rect 5511 -300 6059 -286
rect 6091 -300 6639 -286
rect 6671 -300 6931 -286
rect -1 -424 42 -390
rect 72 -424 478 -390
rect 508 -424 622 -390
rect 652 -424 1058 -390
rect 1088 -424 1202 -390
rect 1232 -424 1638 -390
rect 1668 -424 1782 -390
rect 1812 -424 2218 -390
rect 2248 -424 2362 -390
rect 2392 -424 2798 -390
rect 2828 -424 2942 -390
rect 2972 -424 3378 -390
rect 3408 -424 3522 -390
rect 3552 -424 3958 -390
rect 3988 -424 4102 -390
rect 4132 -424 4538 -390
rect 4591 -424 4682 -390
rect 4712 -424 5118 -390
rect 5148 -424 5262 -390
rect 5292 -424 5698 -390
rect 5728 -424 5842 -390
rect 5872 -424 6278 -390
rect 6308 -424 6422 -390
rect 6452 -424 6858 -390
rect 6888 -424 6931 -390
rect -1 -526 259 -512
rect 291 -526 839 -512
rect 871 -526 1419 -512
rect 1451 -526 1999 -512
rect 2031 -526 2579 -512
rect 2611 -526 3159 -512
rect 3191 -526 3739 -512
rect 3771 -526 4319 -512
rect 4351 -526 4899 -512
rect 4931 -526 5479 -512
rect 5511 -526 6059 -512
rect 6091 -526 6639 -512
rect 6671 -526 6931 -512
rect -1 -570 259 -556
rect 291 -570 839 -556
rect 871 -570 1419 -556
rect 1451 -570 1999 -556
rect 2031 -570 2579 -556
rect 2611 -570 3159 -556
rect 3191 -570 3739 -556
rect 3771 -570 4319 -556
rect 4351 -570 4899 -556
rect 4931 -570 5479 -556
rect 5511 -570 6059 -556
rect 6091 -570 6639 -556
rect 6671 -570 6931 -556
rect -1 -694 42 -660
rect 72 -694 478 -660
rect 508 -694 622 -660
rect 652 -694 1058 -660
rect 1088 -694 1202 -660
rect 1232 -694 1638 -660
rect 1668 -694 1782 -660
rect 1812 -694 2218 -660
rect 2248 -694 2362 -660
rect 2392 -694 2798 -660
rect 2828 -694 2942 -660
rect 2972 -694 3378 -660
rect 3408 -694 3522 -660
rect 3552 -694 3958 -660
rect 3988 -694 4102 -660
rect 4132 -694 4538 -660
rect 4591 -694 4682 -660
rect 4712 -694 5118 -660
rect 5148 -694 5262 -660
rect 5292 -694 5698 -660
rect 5728 -694 5842 -660
rect 5872 -694 6278 -660
rect 6308 -694 6422 -660
rect 6452 -694 6858 -660
rect 6888 -694 6931 -660
rect -1 -796 259 -782
rect 291 -796 839 -782
rect 871 -796 1419 -782
rect 1451 -796 1999 -782
rect 2031 -796 2579 -782
rect 2611 -796 3159 -782
rect 3191 -796 3739 -782
rect 3771 -796 4319 -782
rect 4351 -796 4899 -782
rect 4931 -796 5479 -782
rect 5511 -796 6059 -782
rect 6091 -796 6639 -782
rect 6671 -796 6931 -782
rect -1 -840 259 -826
rect 291 -840 839 -826
rect 871 -840 1419 -826
rect 1451 -840 1999 -826
rect 2031 -840 2579 -826
rect 2611 -840 3159 -826
rect 3191 -840 3739 -826
rect 3771 -840 4319 -826
rect 4351 -840 4899 -826
rect 4931 -840 5479 -826
rect 5511 -840 6059 -826
rect 6091 -840 6639 -826
rect 6671 -840 6931 -826
rect -1 -964 42 -930
rect 72 -964 478 -930
rect 508 -964 622 -930
rect 652 -964 1058 -930
rect 1088 -964 1202 -930
rect 1232 -964 1638 -930
rect 1668 -964 1782 -930
rect 1812 -964 2218 -930
rect 2248 -964 2362 -930
rect 2392 -964 2798 -930
rect 2828 -964 2942 -930
rect 2972 -964 3378 -930
rect 3408 -964 3522 -930
rect 3552 -964 3958 -930
rect 3988 -964 4102 -930
rect 4132 -964 4538 -930
rect 4591 -964 4682 -930
rect 4712 -964 5118 -930
rect 5148 -964 5262 -930
rect 5292 -964 5698 -930
rect 5728 -964 5842 -930
rect 5872 -964 6278 -930
rect 6308 -964 6422 -930
rect 6452 -964 6858 -930
rect 6888 -964 6931 -930
rect -1 -1066 259 -1052
rect 291 -1066 839 -1052
rect 871 -1066 1419 -1052
rect 1451 -1066 1999 -1052
rect 2031 -1066 2579 -1052
rect 2611 -1066 3159 -1052
rect 3191 -1066 3739 -1052
rect 3771 -1066 4319 -1052
rect 4351 -1066 4899 -1052
rect 4931 -1066 5479 -1052
rect 5511 -1066 6059 -1052
rect 6091 -1066 6639 -1052
rect 6671 -1066 6931 -1052
rect -1 -1110 259 -1096
rect 291 -1110 839 -1096
rect 871 -1110 1419 -1096
rect 1451 -1110 1999 -1096
rect 2031 -1110 2579 -1096
rect 2611 -1110 3159 -1096
rect 3191 -1110 3739 -1096
rect 3771 -1110 4319 -1096
rect 4351 -1110 4899 -1096
rect 4931 -1110 5479 -1096
rect 5511 -1110 6059 -1096
rect 6091 -1110 6639 -1096
rect 6671 -1110 6931 -1096
rect -1 -1234 42 -1200
rect 72 -1234 478 -1200
rect 508 -1234 622 -1200
rect 652 -1234 1058 -1200
rect 1088 -1234 1202 -1200
rect 1232 -1234 1638 -1200
rect 1668 -1234 1782 -1200
rect 1812 -1234 2218 -1200
rect 2248 -1234 2362 -1200
rect 2392 -1234 2798 -1200
rect 2828 -1234 2942 -1200
rect 2972 -1234 3378 -1200
rect 3408 -1234 3522 -1200
rect 3552 -1234 3958 -1200
rect 3988 -1234 4102 -1200
rect 4132 -1234 4538 -1200
rect 4591 -1234 4682 -1200
rect 4712 -1234 5118 -1200
rect 5148 -1234 5262 -1200
rect 5292 -1234 5698 -1200
rect 5728 -1234 5842 -1200
rect 5872 -1234 6278 -1200
rect 6308 -1234 6422 -1200
rect 6452 -1234 6858 -1200
rect 6888 -1234 6931 -1200
rect -1 -1336 259 -1322
rect 291 -1336 839 -1322
rect 871 -1336 1419 -1322
rect 1451 -1336 1999 -1322
rect 2031 -1336 2579 -1322
rect 2611 -1336 3159 -1322
rect 3191 -1336 3739 -1322
rect 3771 -1336 4319 -1322
rect 4351 -1336 4899 -1322
rect 4931 -1336 5479 -1322
rect 5511 -1336 6059 -1322
rect 6091 -1336 6639 -1322
rect 6671 -1336 6931 -1322
rect -1 -1380 259 -1366
rect 291 -1380 839 -1366
rect 871 -1380 1419 -1366
rect 1451 -1380 1999 -1366
rect 2031 -1380 2579 -1366
rect 2611 -1380 3159 -1366
rect 3191 -1380 3739 -1366
rect 3771 -1380 4319 -1366
rect 4351 -1380 4899 -1366
rect 4931 -1380 5479 -1366
rect 5511 -1380 6059 -1366
rect 6091 -1380 6639 -1366
rect 6671 -1380 6931 -1366
rect -1 -1504 42 -1470
rect 72 -1504 478 -1470
rect 508 -1504 622 -1470
rect 652 -1504 1058 -1470
rect 1088 -1504 1202 -1470
rect 1232 -1504 1638 -1470
rect 1668 -1504 1782 -1470
rect 1812 -1504 2218 -1470
rect 2248 -1504 2362 -1470
rect 2392 -1504 2798 -1470
rect 2828 -1504 2942 -1470
rect 2972 -1504 3378 -1470
rect 3408 -1504 3522 -1470
rect 3552 -1504 3958 -1470
rect 3988 -1504 4102 -1470
rect 4132 -1504 4538 -1470
rect 4591 -1504 4682 -1470
rect 4712 -1504 5118 -1470
rect 5148 -1504 5262 -1470
rect 5292 -1504 5698 -1470
rect 5728 -1504 5842 -1470
rect 5872 -1504 6278 -1470
rect 6308 -1504 6422 -1470
rect 6452 -1504 6858 -1470
rect 6888 -1504 6931 -1470
rect -1 -1606 259 -1592
rect 291 -1606 839 -1592
rect 871 -1606 1419 -1592
rect 1451 -1606 1999 -1592
rect 2031 -1606 2579 -1592
rect 2611 -1606 3159 -1592
rect 3191 -1606 3739 -1592
rect 3771 -1606 4319 -1592
rect 4351 -1606 4899 -1592
rect 4931 -1606 5479 -1592
rect 5511 -1606 6059 -1592
rect 6091 -1606 6639 -1592
rect 6671 -1606 6931 -1592
rect -1 -1650 259 -1636
rect 291 -1650 839 -1636
rect 871 -1650 1419 -1636
rect 1451 -1650 1999 -1636
rect 2031 -1650 2579 -1636
rect 2611 -1650 3159 -1636
rect 3191 -1650 3739 -1636
rect 3771 -1650 4319 -1636
rect 4351 -1650 4899 -1636
rect 4931 -1650 5479 -1636
rect 5511 -1650 6059 -1636
rect 6091 -1650 6639 -1636
rect 6671 -1650 6931 -1636
rect -1 -1774 42 -1740
rect 72 -1774 478 -1740
rect 508 -1774 622 -1740
rect 652 -1774 1058 -1740
rect 1088 -1774 1202 -1740
rect 1232 -1774 1638 -1740
rect 1668 -1774 1782 -1740
rect 1812 -1774 2218 -1740
rect 2248 -1774 2362 -1740
rect 2392 -1774 2798 -1740
rect 2828 -1774 2942 -1740
rect 2972 -1774 3378 -1740
rect 3408 -1774 3522 -1740
rect 3552 -1774 3958 -1740
rect 3988 -1774 4102 -1740
rect 4132 -1774 4538 -1740
rect 4591 -1774 4682 -1740
rect 4712 -1774 5118 -1740
rect 5148 -1774 5262 -1740
rect 5292 -1774 5698 -1740
rect 5728 -1774 5842 -1740
rect 5872 -1774 6278 -1740
rect 6308 -1774 6422 -1740
rect 6452 -1774 6858 -1740
rect 6888 -1774 6931 -1740
rect -1 -1876 259 -1862
rect 291 -1876 839 -1862
rect 871 -1876 1419 -1862
rect 1451 -1876 1999 -1862
rect 2031 -1876 2579 -1862
rect 2611 -1876 3159 -1862
rect 3191 -1876 3739 -1862
rect 3771 -1876 4319 -1862
rect 4351 -1876 4899 -1862
rect 4931 -1876 5479 -1862
rect 5511 -1876 6059 -1862
rect 6091 -1876 6639 -1862
rect 6671 -1876 6931 -1862
rect -1 -1920 259 -1906
rect 291 -1920 839 -1906
rect 871 -1920 1419 -1906
rect 1451 -1920 1999 -1906
rect 2031 -1920 2579 -1906
rect 2611 -1920 3159 -1906
rect 3191 -1920 3739 -1906
rect 3771 -1920 4319 -1906
rect 4351 -1920 4899 -1906
rect 4931 -1920 5479 -1906
rect 5511 -1920 6059 -1906
rect 6091 -1920 6639 -1906
rect 6671 -1920 6931 -1906
rect -1 -2044 42 -2010
rect 72 -2044 478 -2010
rect 508 -2044 622 -2010
rect 652 -2044 1058 -2010
rect 1088 -2044 1202 -2010
rect 1232 -2044 1638 -2010
rect 1668 -2044 1782 -2010
rect 1812 -2044 2218 -2010
rect 2248 -2044 2362 -2010
rect 2392 -2044 2798 -2010
rect 2828 -2044 2942 -2010
rect 2972 -2044 3378 -2010
rect 3408 -2044 3522 -2010
rect 3552 -2044 3958 -2010
rect 3988 -2044 4102 -2010
rect 4132 -2044 4538 -2010
rect 4591 -2044 4682 -2010
rect 4712 -2044 5118 -2010
rect 5148 -2044 5262 -2010
rect 5292 -2044 5698 -2010
rect 5728 -2044 5842 -2010
rect 5872 -2044 6278 -2010
rect 6308 -2044 6422 -2010
rect 6452 -2044 6858 -2010
rect 6888 -2044 6931 -2010
rect -1 -2146 259 -2132
rect 291 -2146 839 -2132
rect 871 -2146 1419 -2132
rect 1451 -2146 1999 -2132
rect 2031 -2146 2579 -2132
rect 2611 -2146 3159 -2132
rect 3191 -2146 3739 -2132
rect 3771 -2146 4319 -2132
rect 4351 -2146 4899 -2132
rect 4931 -2146 5479 -2132
rect 5511 -2146 6059 -2132
rect 6091 -2146 6639 -2132
rect 6671 -2146 6931 -2132
<< labels >>
rlabel poly -1 2144 6931 2174 1 WWL_0
port 1 n
rlabel metal1 73 2088 88 2116 1 WBLb_0
port 2 n
rlabel metal1 463 2088 478 2117 1 WBL_0
port 3 n
rlabel metal1 259 2130 291 2144 1 VDD
port 4 n
rlabel metal1 -1 1942 14 1984 1 RBL1_0
port 5 n
rlabel metal1 536 1942 551 1984 1 RBL0_0
port 6 n
rlabel metal1 42 2006 72 2040 1 RWL_0
port 7 n
rlabel metal1 259 1904 291 1918 1 GND
port 8 n
rlabel metal1 -1 2006 14 2040 1 RWL_0
port 7 n
rlabel poly -1 1874 6931 1904 1 WWL_1
port 9 n
rlabel poly -1 1874 14 1904 1 WWL_1
port 9 n
rlabel metal1 73 1818 88 1846 1 WBLb_1
port 10 n
rlabel metal1 463 1818 478 1847 1 WBL_1
port 11 n
rlabel metal1 -1 1672 14 1714 1 RBL1_1
port 12 n
rlabel metal1 536 1672 551 1714 1 RBL0_1
port 13 n
rlabel metal1 259 1860 291 1874 1 VDD
port 4 n
rlabel metal1 259 1634 291 1648 1 GND
port 8 n
rlabel metal1 42 1736 72 1770 1 RWL_1
port 14 n
rlabel metal1 -1 1736 14 1770 1 RWL_1
port 14 n
rlabel poly -1 1604 6931 1634 1 WWL_2
port 15 n
rlabel metal1 -1 1604 14 1634 1 WWL_2
port 15 n
rlabel metal1 73 1548 88 1576 1 WBLb_2
port 16 n
rlabel metal1 42 1466 72 1500 1 RWL_2
port 17 n
rlabel metal1 -1 1466 14 1500 1 RWL_2
port 17 n
rlabel metal1 -1 1402 14 1444 1 RBL1_2
port 18 n
rlabel metal1 259 1590 291 1604 1 VDD
port 4 n
rlabel metal1 259 1364 291 1378 1 GND
port 8 n
rlabel metal1 463 1548 478 1577 1 WBL_2
port 19 n
rlabel metal1 536 1402 551 1444 1 RBL0_2
port 20 n
rlabel poly -1 1334 6931 1364 1 WWL_3
port 21 n
rlabel metal1 -1 1334 14 1364 1 WWL_3
port 21 n
rlabel metal1 73 1278 88 1306 1 WBLb_3
port 22 n
rlabel metal1 259 1320 291 1334 1 VDD
port 4 n
rlabel metal1 42 1196 72 1230 1 RWL_3
port 23 n
rlabel metal1 -1 1196 14 1230 1 RWL_3
port 23 n
rlabel metal1 259 1094 291 1108 1 GND
port 8 n
rlabel metal1 463 1278 478 1307 1 WBL_3
port 25 n
rlabel metal1 536 1132 551 1174 1 RBL0_3
port 26 n
rlabel poly -1 1064 6931 1094 1 WWL_4
port 27 n
rlabel metal1 73 1008 88 1036 1 WBLb_4
port 28 n
rlabel metal1 42 926 72 960 1 RWL_4
port 29 n
rlabel metal1 -1 1064 14 1094 1 WWL_4
port 27 n
rlabel metal1 -1 1132 14 1174 1 RBL1_3
port 24 n
rlabel metal1 -1 926 14 960 1 RWL_4
port 29 n
rlabel metal1 -1 862 14 904 1 RBL1_4
port 30 n
rlabel metal1 259 1050 291 1064 1 VDD
port 4 n
rlabel metal1 259 824 291 838 1 GND
port 8 n
rlabel metal1 463 1008 478 1037 1 WBL_4
port 31 n
rlabel metal1 536 862 551 904 1 RBL0_4
port 32 n
rlabel poly -1 794 6931 824 1 WWL_5
port 33 n
rlabel metal1 -1 794 14 824 1 WWL_5
port 33 n
rlabel metal1 73 738 88 766 1 WBLb_5
port 34 n
rlabel metal1 42 656 72 690 1 RWL_5
port 35 n
rlabel metal1 -1 656 14 690 1 RWL_5
port 35 n
rlabel metal1 -1 592 14 634 1 RBL1_5
port 36 n
rlabel metal1 259 780 291 794 1 VDD
port 4 n
rlabel metal1 259 554 291 568 1 GND
port 8 n
rlabel metal1 463 738 478 767 1 WBL_5
port 37 n
rlabel metal1 536 592 551 634 1 RBL0_5
port 38 n
rlabel poly -1 524 6931 554 1 WWL_6
port 39 n
rlabel metal1 -1 524 14 554 1 WWL_6
port 39 n
rlabel metal1 73 468 88 496 1 WBLb_6
port 40 n
rlabel metal1 -1 322 14 364 1 RBL1_6
port 41 n
rlabel metal1 259 510 291 524 1 VDD
port 4 n
rlabel metal1 259 284 291 298 1 GND
port 8 n
rlabel metal1 463 468 478 497 1 WBL_6
port 42 n
rlabel metal1 536 322 551 364 1 RBL0_6
port 43 n
rlabel poly -1 254 6931 284 1 WWL_7
port 44 n
rlabel poly -1 254 14 284 1 WWL_7
port 44 n
rlabel metal1 73 198 88 226 1 WBLb_7
port 45 n
rlabel metal1 259 240 291 254 1 VDD
port 4 n
rlabel metal1 463 198 478 227 1 WBL_7
port 46 n
rlabel metal1 536 52 551 94 1 RBL0_7
port 47 n
rlabel metal1 259 14 291 28 1 GND
port 8 n
rlabel metal1 -1 52 14 94 1 RBL1_7
port 48 n
rlabel poly -1 -16 6931 14 1 WWL_8
port 49 n
rlabel poly -1 -16 14 14 1 WWL_8
port 49 n
rlabel metal1 73 -72 88 -44 1 WBLb_8
port 50 n
rlabel metal1 -1 -218 14 -176 1 RBL1_8
port 51 n
rlabel metal1 259 -30 291 -16 1 VDD
port 4 n
rlabel metal1 463 -72 478 -43 1 WBL_8
port 52 n
rlabel metal1 536 -218 551 -176 1 RBL0_8
port 53 n
rlabel metal1 259 -256 291 -242 1 GND
port 8 n
rlabel poly -1 -286 6931 -256 1 WWL_9
port 54 n
rlabel poly -1 -286 14 -256 1 WWL_9
port 54 n
rlabel metal1 73 -342 88 -314 1 WBLb_9
port 55 n
rlabel metal1 -1 -488 14 -446 1 RBL1_9
port 56 n
rlabel metal1 259 -526 291 -512 1 GND
port 8 n
rlabel metal1 259 -300 291 -286 1 VDD
port 4 n
rlabel metal1 463 -342 478 -313 1 WBL_9
port 57 n
rlabel metal1 536 -488 551 -446 1 RBL0_9
port 58 n
rlabel poly -1 -556 6931 -526 1 WWL_10
port 59 n
rlabel poly -1 -556 14 -526 1 WWL_10
port 59 n
rlabel metal1 73 -612 88 -584 1 WBLb_10
port 60 n
rlabel metal1 259 -570 291 -556 1 VDD
port 4 n
rlabel metal1 463 -612 478 -583 1 WBL_10
port 61 n
rlabel metal1 536 -758 551 -716 1 RBL0_10
port 62 n
rlabel metal1 259 -796 291 -782 1 GND
port 8 n
rlabel metal1 -1 -758 14 -716 1 RBL1_10
port 63 n
rlabel poly -1 -826 6931 -796 1 WWL_11
port 64 n
rlabel metal1 -1 -826 14 -796 1 WWL_11
port 64 n
rlabel metal1 73 -882 88 -854 1 WBLb_11
port 65 n
rlabel metal1 -1 -1028 14 -986 1 RBL1_11
port 66 n
rlabel metal1 259 -1066 291 -1052 1 GND
port 8 n
rlabel metal1 259 -840 291 -826 1 VDD
port 4 n
rlabel metal1 463 -882 478 -853 1 WBL_11
port 67 n
rlabel metal1 536 -1028 551 -986 1 RBL0_11
port 68 n
rlabel poly -1 -1096 6931 -1066 1 WWL_12
port 69 n
rlabel poly -1 -1096 14 -1066 1 WWL_12
port 69 n
rlabel metal1 73 -1152 88 -1124 1 WBLb_12
port 70 n
rlabel metal1 -1 -1298 14 -1256 1 RBL1_12
port 71 n
rlabel metal1 259 -1110 291 -1096 1 VDD
port 4 n
rlabel metal1 259 -1336 291 -1322 1 GND
port 8 n
rlabel metal1 463 -1152 478 -1123 1 WBL_12
port 72 n
rlabel metal1 536 -1298 551 -1256 1 RBL0_12
port 73 n
rlabel poly -1 -1366 6931 -1336 1 WWL_13
port 74 n
rlabel poly -1 -1366 14 -1336 1 WWL_13
port 74 n
rlabel metal1 73 -1422 88 -1394 1 WBLb_13
port 75 n
rlabel metal1 -1 -1568 14 -1526 1 RBL1_13
port 76 n
rlabel metal1 259 -1380 291 -1366 1 VDD
port 4 n
rlabel metal1 463 -1422 478 -1393 1 WBL_13
port 77 n
rlabel metal1 536 -1568 551 -1526 1 RBL0_13
port 78 n
rlabel metal1 259 -1606 291 -1592 1 GND
port 8 n
rlabel poly -1 -1636 6931 -1606 1 WWL_14
port 79 n
rlabel poly -1 -1636 14 -1606 1 WWL_14
port 79 n
rlabel metal1 73 -1692 88 -1664 1 WBLb_14
port 80 n
rlabel metal1 -1 -1838 14 -1796 1 RBL1_14
port 81 n
rlabel metal1 259 -1650 291 -1636 1 VDD
port 4 n
rlabel metal1 463 -1692 478 -1663 1 WBL_14
port 82 n
rlabel metal1 536 -1838 551 -1796 1 RBL0_14
port 83 n
rlabel metal1 259 -1876 291 -1862 1 GND
port 8 n
rlabel poly -1 -1906 6931 -1876 1 WWL_15
port 84 n
rlabel poly -1 -1906 14 -1876 1 WWL_15
port 84 n
rlabel metal1 -1 -2108 14 -2066 1 RBL1_15
port 86 n
rlabel metal1 73 -1962 88 -1934 1 WBLb_15
port 85 n
rlabel metal1 259 -2146 291 -2132 1 GND
port 8 n
rlabel metal1 259 -1920 291 -1906 1 VDD
port 4 n
rlabel metal1 463 -1962 478 -1933 1 WBL_15
port 87 n
rlabel metal1 536 -2108 551 -2066 1 RBL0_15
port 88 n
<< end >>
