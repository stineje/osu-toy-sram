** sch_path: /home/rjridle/osu-toy-sram/custom_layout/10T_toy_xschem.sch
.subckt 10T_toy_xschem WWL RWL0 RWL1 WBL WBLb RBL0 RBL1 VDD GND
*.PININFO WWL:I RWL0:I RWL1:I WBL:I WBLb:I RBL0:O RBL1:O
XM1 net1 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 
XM2 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1
XM3 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM4 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1
XM5 net2 WWL WBL GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 
XM6 WBLb WWL net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 
XM7 net3 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 
XM8 RBL0 RWL0 net3 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM9 net4 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 
XM10 RBL1 RWL1 net4 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1
.ends

.end
