magic
tech sky130A
magscale 1 2
timestamp 1667336911
<< error_s >>
rect 15 1064 28 1080
rect 117 1078 130 1080
rect 83 1064 98 1078
rect 107 1064 137 1078
rect 198 1076 351 1122
rect 180 1064 372 1076
rect 415 1064 445 1078
rect 451 1064 464 1080
rect 552 1064 565 1080
rect 595 1064 608 1080
rect 697 1078 710 1080
rect 663 1064 678 1078
rect 687 1064 717 1078
rect 778 1076 931 1122
rect 760 1064 952 1076
rect 995 1064 1025 1078
rect 1031 1064 1044 1080
rect 1132 1064 1145 1080
rect 1175 1064 1188 1080
rect 1277 1078 1290 1080
rect 1243 1064 1258 1078
rect 1267 1064 1297 1078
rect 1358 1076 1511 1122
rect 1340 1064 1532 1076
rect 1575 1064 1605 1078
rect 1611 1064 1624 1080
rect 1712 1064 1725 1080
rect 1755 1064 1768 1080
rect 1857 1078 1870 1080
rect 1823 1064 1838 1078
rect 1847 1064 1877 1078
rect 1938 1076 2091 1122
rect 1920 1064 2112 1076
rect 2155 1064 2185 1078
rect 2191 1064 2204 1080
rect 2292 1064 2305 1080
rect 2335 1064 2348 1080
rect 2437 1078 2450 1080
rect 2403 1064 2418 1078
rect 2427 1064 2457 1078
rect 2518 1076 2671 1122
rect 2500 1064 2692 1076
rect 2735 1064 2765 1078
rect 2771 1064 2784 1080
rect 2872 1064 2885 1080
rect 2915 1064 2928 1080
rect 3017 1078 3030 1080
rect 2983 1064 2998 1078
rect 3007 1064 3037 1078
rect 3098 1076 3251 1122
rect 3080 1064 3272 1076
rect 3315 1064 3345 1078
rect 3351 1064 3364 1080
rect 3452 1064 3465 1080
rect 3495 1064 3508 1080
rect 3597 1078 3610 1080
rect 3563 1064 3578 1078
rect 3587 1064 3617 1078
rect 3678 1076 3831 1122
rect 3660 1064 3852 1076
rect 3895 1064 3925 1078
rect 3931 1064 3944 1080
rect 4032 1064 4045 1080
rect 4075 1064 4088 1080
rect 4177 1078 4190 1080
rect 4143 1064 4158 1078
rect 4167 1064 4197 1078
rect 4258 1076 4411 1122
rect 4240 1064 4432 1076
rect 4475 1064 4505 1078
rect 4511 1064 4524 1080
rect 4612 1064 4625 1080
rect 0 1050 4625 1064
rect 15 946 28 1050
rect 73 1028 74 1038
rect 89 1028 102 1038
rect 73 1024 102 1028
rect 107 1024 137 1050
rect 155 1036 171 1038
rect 243 1036 296 1050
rect 244 1034 308 1036
rect 351 1034 366 1050
rect 415 1047 445 1050
rect 415 1044 451 1047
rect 381 1036 397 1038
rect 155 1024 170 1028
rect 73 1022 170 1024
rect 198 1022 366 1034
rect 382 1024 397 1028
rect 415 1025 454 1044
rect 473 1038 480 1039
rect 479 1031 480 1038
rect 463 1028 464 1031
rect 479 1028 492 1031
rect 415 1024 445 1025
rect 454 1024 460 1025
rect 463 1024 492 1028
rect 382 1023 492 1024
rect 382 1022 498 1023
rect 57 1014 108 1022
rect 57 1002 82 1014
rect 89 1002 108 1014
rect 139 1014 189 1022
rect 139 1006 155 1014
rect 162 1012 189 1014
rect 198 1012 419 1022
rect 162 1002 419 1012
rect 448 1014 498 1022
rect 448 1005 464 1014
rect 57 994 108 1002
rect 155 994 419 1002
rect 445 1002 464 1005
rect 471 1002 498 1014
rect 445 994 498 1002
rect 73 986 74 994
rect 89 986 102 994
rect 73 978 89 986
rect 70 971 89 974
rect 70 962 92 971
rect 43 952 92 962
rect 43 946 73 952
rect 92 947 97 952
rect 15 930 89 946
rect 107 938 137 994
rect 172 984 380 994
rect 415 990 460 994
rect 463 993 464 994
rect 479 993 492 994
rect 198 954 387 984
rect 213 951 387 954
rect 206 948 387 951
rect 15 928 28 930
rect 43 928 77 930
rect 15 912 89 928
rect 116 924 129 938
rect 144 924 160 940
rect 206 935 217 948
rect -1 890 0 906
rect 15 890 28 912
rect 43 890 73 912
rect 116 908 178 924
rect 206 917 217 933
rect 222 928 232 948
rect 242 928 256 948
rect 259 935 268 948
rect 284 935 293 948
rect 222 917 256 928
rect 259 917 268 933
rect 284 917 293 933
rect 300 928 310 948
rect 320 928 334 948
rect 335 935 346 948
rect 300 917 334 928
rect 335 917 346 933
rect 392 924 408 940
rect 415 938 445 990
rect 479 986 480 993
rect 464 978 480 986
rect 451 946 464 965
rect 479 946 509 962
rect 451 930 525 946
rect 451 928 464 930
rect 479 928 513 930
rect 116 906 129 908
rect 144 906 178 908
rect 116 890 178 906
rect 222 901 238 904
rect 300 901 330 912
rect 378 908 424 924
rect 451 912 525 928
rect 378 906 412 908
rect 377 890 424 906
rect 451 890 464 912
rect 479 890 509 912
rect 536 890 537 906
rect 552 890 565 1050
rect 595 946 608 1050
rect 653 1028 654 1038
rect 669 1028 682 1038
rect 653 1024 682 1028
rect 687 1024 717 1050
rect 735 1036 751 1038
rect 823 1036 876 1050
rect 824 1034 888 1036
rect 931 1034 946 1050
rect 995 1047 1025 1050
rect 995 1044 1031 1047
rect 961 1036 977 1038
rect 735 1024 750 1028
rect 653 1022 750 1024
rect 778 1022 946 1034
rect 962 1024 977 1028
rect 995 1025 1034 1044
rect 1053 1038 1060 1039
rect 1059 1031 1060 1038
rect 1043 1028 1044 1031
rect 1059 1028 1072 1031
rect 995 1024 1025 1025
rect 1034 1024 1040 1025
rect 1043 1024 1072 1028
rect 962 1023 1072 1024
rect 962 1022 1078 1023
rect 637 1014 688 1022
rect 637 1002 662 1014
rect 669 1002 688 1014
rect 719 1014 769 1022
rect 719 1006 735 1014
rect 742 1012 769 1014
rect 778 1012 999 1022
rect 742 1002 999 1012
rect 1028 1014 1078 1022
rect 1028 1005 1044 1014
rect 637 994 688 1002
rect 735 994 999 1002
rect 1025 1002 1044 1005
rect 1051 1002 1078 1014
rect 1025 994 1078 1002
rect 653 986 654 994
rect 669 986 682 994
rect 653 978 669 986
rect 650 971 669 974
rect 650 962 672 971
rect 623 952 672 962
rect 623 946 653 952
rect 672 947 677 952
rect 595 930 669 946
rect 687 938 717 994
rect 752 984 960 994
rect 995 990 1040 994
rect 1043 993 1044 994
rect 1059 993 1072 994
rect 778 954 967 984
rect 793 951 967 954
rect 786 948 967 951
rect 595 928 608 930
rect 623 928 657 930
rect 595 912 669 928
rect 696 924 709 938
rect 724 924 740 940
rect 786 935 797 948
rect 579 890 580 906
rect 595 890 608 912
rect 623 890 653 912
rect 696 908 758 924
rect 786 917 797 933
rect 802 928 812 948
rect 822 928 836 948
rect 839 935 848 948
rect 864 935 873 948
rect 802 917 836 928
rect 839 917 848 933
rect 864 917 873 933
rect 880 928 890 948
rect 900 928 914 948
rect 915 935 926 948
rect 880 917 914 928
rect 915 917 926 933
rect 972 924 988 940
rect 995 938 1025 990
rect 1059 986 1060 993
rect 1044 978 1060 986
rect 1031 946 1044 965
rect 1059 946 1089 962
rect 1031 930 1105 946
rect 1031 928 1044 930
rect 1059 928 1093 930
rect 696 906 709 908
rect 724 906 758 908
rect 696 890 758 906
rect 802 901 818 904
rect 880 901 910 912
rect 958 908 1004 924
rect 1031 912 1105 928
rect 958 906 992 908
rect 957 890 1004 906
rect 1031 890 1044 912
rect 1059 890 1089 912
rect 1116 890 1117 906
rect 1132 890 1145 1050
rect 1175 946 1188 1050
rect 1233 1028 1234 1038
rect 1249 1028 1262 1038
rect 1233 1024 1262 1028
rect 1267 1024 1297 1050
rect 1315 1036 1331 1038
rect 1403 1036 1456 1050
rect 1404 1034 1468 1036
rect 1511 1034 1526 1050
rect 1575 1047 1605 1050
rect 1575 1044 1611 1047
rect 1541 1036 1557 1038
rect 1315 1024 1330 1028
rect 1233 1022 1330 1024
rect 1358 1022 1526 1034
rect 1542 1024 1557 1028
rect 1575 1025 1614 1044
rect 1633 1038 1640 1039
rect 1639 1031 1640 1038
rect 1623 1028 1624 1031
rect 1639 1028 1652 1031
rect 1575 1024 1605 1025
rect 1614 1024 1620 1025
rect 1623 1024 1652 1028
rect 1542 1023 1652 1024
rect 1542 1022 1658 1023
rect 1217 1014 1268 1022
rect 1217 1002 1242 1014
rect 1249 1002 1268 1014
rect 1299 1014 1349 1022
rect 1299 1006 1315 1014
rect 1322 1012 1349 1014
rect 1358 1012 1579 1022
rect 1322 1002 1579 1012
rect 1608 1014 1658 1022
rect 1608 1005 1624 1014
rect 1217 994 1268 1002
rect 1315 994 1579 1002
rect 1605 1002 1624 1005
rect 1631 1002 1658 1014
rect 1605 994 1658 1002
rect 1233 986 1234 994
rect 1249 986 1262 994
rect 1233 978 1249 986
rect 1230 971 1249 974
rect 1230 962 1252 971
rect 1203 952 1252 962
rect 1203 946 1233 952
rect 1252 947 1257 952
rect 1175 930 1249 946
rect 1267 938 1297 994
rect 1332 984 1540 994
rect 1575 990 1620 994
rect 1623 993 1624 994
rect 1639 993 1652 994
rect 1358 954 1547 984
rect 1373 951 1547 954
rect 1366 948 1547 951
rect 1175 928 1188 930
rect 1203 928 1237 930
rect 1175 912 1249 928
rect 1276 924 1289 938
rect 1304 924 1320 940
rect 1366 935 1377 948
rect 1159 890 1160 906
rect 1175 890 1188 912
rect 1203 890 1233 912
rect 1276 908 1338 924
rect 1366 917 1377 933
rect 1382 928 1392 948
rect 1402 928 1416 948
rect 1419 935 1428 948
rect 1444 935 1453 948
rect 1382 917 1416 928
rect 1419 917 1428 933
rect 1444 917 1453 933
rect 1460 928 1470 948
rect 1480 928 1494 948
rect 1495 935 1506 948
rect 1460 917 1494 928
rect 1495 917 1506 933
rect 1552 924 1568 940
rect 1575 938 1605 990
rect 1639 986 1640 993
rect 1624 978 1640 986
rect 1611 946 1624 965
rect 1639 946 1669 962
rect 1611 930 1685 946
rect 1611 928 1624 930
rect 1639 928 1673 930
rect 1276 906 1289 908
rect 1304 906 1338 908
rect 1276 890 1338 906
rect 1382 901 1398 904
rect 1460 901 1490 912
rect 1538 908 1584 924
rect 1611 912 1685 928
rect 1538 906 1572 908
rect 1537 890 1584 906
rect 1611 890 1624 912
rect 1639 890 1669 912
rect 1696 890 1697 906
rect 1712 890 1725 1050
rect 1755 946 1768 1050
rect 1813 1028 1814 1038
rect 1829 1028 1842 1038
rect 1813 1024 1842 1028
rect 1847 1024 1877 1050
rect 1895 1036 1911 1038
rect 1983 1036 2036 1050
rect 1984 1034 2048 1036
rect 2091 1034 2106 1050
rect 2155 1047 2185 1050
rect 2155 1044 2191 1047
rect 2121 1036 2137 1038
rect 1895 1024 1910 1028
rect 1813 1022 1910 1024
rect 1938 1022 2106 1034
rect 2122 1024 2137 1028
rect 2155 1025 2194 1044
rect 2213 1038 2220 1039
rect 2219 1031 2220 1038
rect 2203 1028 2204 1031
rect 2219 1028 2232 1031
rect 2155 1024 2185 1025
rect 2194 1024 2200 1025
rect 2203 1024 2232 1028
rect 2122 1023 2232 1024
rect 2122 1022 2238 1023
rect 1797 1014 1848 1022
rect 1797 1002 1822 1014
rect 1829 1002 1848 1014
rect 1879 1014 1929 1022
rect 1879 1006 1895 1014
rect 1902 1012 1929 1014
rect 1938 1012 2159 1022
rect 1902 1002 2159 1012
rect 2188 1014 2238 1022
rect 2188 1005 2204 1014
rect 1797 994 1848 1002
rect 1895 994 2159 1002
rect 2185 1002 2204 1005
rect 2211 1002 2238 1014
rect 2185 994 2238 1002
rect 1813 986 1814 994
rect 1829 986 1842 994
rect 1813 978 1829 986
rect 1810 971 1829 974
rect 1810 962 1832 971
rect 1783 952 1832 962
rect 1783 946 1813 952
rect 1832 947 1837 952
rect 1755 930 1829 946
rect 1847 938 1877 994
rect 1912 984 2120 994
rect 2155 990 2200 994
rect 2203 993 2204 994
rect 2219 993 2232 994
rect 1938 954 2127 984
rect 1953 951 2127 954
rect 1946 948 2127 951
rect 1755 928 1768 930
rect 1783 928 1817 930
rect 1755 912 1829 928
rect 1856 924 1869 938
rect 1884 924 1900 940
rect 1946 935 1957 948
rect 1739 890 1740 906
rect 1755 890 1768 912
rect 1783 890 1813 912
rect 1856 908 1918 924
rect 1946 917 1957 933
rect 1962 928 1972 948
rect 1982 928 1996 948
rect 1999 935 2008 948
rect 2024 935 2033 948
rect 1962 917 1996 928
rect 1999 917 2008 933
rect 2024 917 2033 933
rect 2040 928 2050 948
rect 2060 928 2074 948
rect 2075 935 2086 948
rect 2040 917 2074 928
rect 2075 917 2086 933
rect 2132 924 2148 940
rect 2155 938 2185 990
rect 2219 986 2220 993
rect 2204 978 2220 986
rect 2191 946 2204 965
rect 2219 946 2249 962
rect 2191 930 2265 946
rect 2191 928 2204 930
rect 2219 928 2253 930
rect 1856 906 1869 908
rect 1884 906 1918 908
rect 1856 890 1918 906
rect 1962 901 1978 904
rect 2040 901 2070 912
rect 2118 908 2164 924
rect 2191 912 2265 928
rect 2118 906 2152 908
rect 2117 890 2164 906
rect 2191 890 2204 912
rect 2219 890 2249 912
rect 2276 890 2277 906
rect 2292 890 2305 1050
rect 2335 946 2348 1050
rect 2393 1028 2394 1038
rect 2409 1028 2422 1038
rect 2393 1024 2422 1028
rect 2427 1024 2457 1050
rect 2475 1036 2491 1038
rect 2563 1036 2616 1050
rect 2564 1034 2628 1036
rect 2671 1034 2686 1050
rect 2735 1047 2765 1050
rect 2735 1044 2771 1047
rect 2701 1036 2717 1038
rect 2475 1024 2490 1028
rect 2393 1022 2490 1024
rect 2518 1022 2686 1034
rect 2702 1024 2717 1028
rect 2735 1025 2774 1044
rect 2793 1038 2800 1039
rect 2799 1031 2800 1038
rect 2783 1028 2784 1031
rect 2799 1028 2812 1031
rect 2735 1024 2765 1025
rect 2774 1024 2780 1025
rect 2783 1024 2812 1028
rect 2702 1023 2812 1024
rect 2702 1022 2818 1023
rect 2377 1014 2428 1022
rect 2377 1002 2402 1014
rect 2409 1002 2428 1014
rect 2459 1014 2509 1022
rect 2459 1006 2475 1014
rect 2482 1012 2509 1014
rect 2518 1012 2739 1022
rect 2482 1002 2739 1012
rect 2768 1014 2818 1022
rect 2768 1005 2784 1014
rect 2377 994 2428 1002
rect 2475 994 2739 1002
rect 2765 1002 2784 1005
rect 2791 1002 2818 1014
rect 2765 994 2818 1002
rect 2393 986 2394 994
rect 2409 986 2422 994
rect 2393 978 2409 986
rect 2390 971 2409 974
rect 2390 962 2412 971
rect 2363 952 2412 962
rect 2363 946 2393 952
rect 2412 947 2417 952
rect 2335 930 2409 946
rect 2427 938 2457 994
rect 2492 984 2700 994
rect 2735 990 2780 994
rect 2783 993 2784 994
rect 2799 993 2812 994
rect 2518 954 2707 984
rect 2533 951 2707 954
rect 2526 948 2707 951
rect 2335 928 2348 930
rect 2363 928 2397 930
rect 2335 912 2409 928
rect 2436 924 2449 938
rect 2464 924 2480 940
rect 2526 935 2537 948
rect 2319 890 2320 906
rect 2335 890 2348 912
rect 2363 890 2393 912
rect 2436 908 2498 924
rect 2526 917 2537 933
rect 2542 928 2552 948
rect 2562 928 2576 948
rect 2579 935 2588 948
rect 2604 935 2613 948
rect 2542 917 2576 928
rect 2579 917 2588 933
rect 2604 917 2613 933
rect 2620 928 2630 948
rect 2640 928 2654 948
rect 2655 935 2666 948
rect 2620 917 2654 928
rect 2655 917 2666 933
rect 2712 924 2728 940
rect 2735 938 2765 990
rect 2799 986 2800 993
rect 2784 978 2800 986
rect 2771 946 2784 965
rect 2799 946 2829 962
rect 2771 930 2845 946
rect 2771 928 2784 930
rect 2799 928 2833 930
rect 2436 906 2449 908
rect 2464 906 2498 908
rect 2436 890 2498 906
rect 2542 901 2558 904
rect 2620 901 2650 912
rect 2698 908 2744 924
rect 2771 912 2845 928
rect 2698 906 2732 908
rect 2697 890 2744 906
rect 2771 890 2784 912
rect 2799 890 2829 912
rect 2856 890 2857 906
rect 2872 890 2885 1050
rect 2915 946 2928 1050
rect 2973 1028 2974 1038
rect 2989 1028 3002 1038
rect 2973 1024 3002 1028
rect 3007 1024 3037 1050
rect 3055 1036 3071 1038
rect 3143 1036 3196 1050
rect 3144 1034 3208 1036
rect 3251 1034 3266 1050
rect 3315 1047 3345 1050
rect 3315 1044 3351 1047
rect 3281 1036 3297 1038
rect 3055 1024 3070 1028
rect 2973 1022 3070 1024
rect 3098 1022 3266 1034
rect 3282 1024 3297 1028
rect 3315 1025 3354 1044
rect 3373 1038 3380 1039
rect 3379 1031 3380 1038
rect 3363 1028 3364 1031
rect 3379 1028 3392 1031
rect 3315 1024 3345 1025
rect 3354 1024 3360 1025
rect 3363 1024 3392 1028
rect 3282 1023 3392 1024
rect 3282 1022 3398 1023
rect 2957 1014 3008 1022
rect 2957 1002 2982 1014
rect 2989 1002 3008 1014
rect 3039 1014 3089 1022
rect 3039 1006 3055 1014
rect 3062 1012 3089 1014
rect 3098 1012 3319 1022
rect 3062 1002 3319 1012
rect 3348 1014 3398 1022
rect 3348 1005 3364 1014
rect 2957 994 3008 1002
rect 3055 994 3319 1002
rect 3345 1002 3364 1005
rect 3371 1002 3398 1014
rect 3345 994 3398 1002
rect 2973 986 2974 994
rect 2989 986 3002 994
rect 2973 978 2989 986
rect 2970 971 2989 974
rect 2970 962 2992 971
rect 2943 952 2992 962
rect 2943 946 2973 952
rect 2992 947 2997 952
rect 2915 930 2989 946
rect 3007 938 3037 994
rect 3072 984 3280 994
rect 3315 990 3360 994
rect 3363 993 3364 994
rect 3379 993 3392 994
rect 3098 954 3287 984
rect 3113 951 3287 954
rect 3106 948 3287 951
rect 2915 928 2928 930
rect 2943 928 2977 930
rect 2915 912 2989 928
rect 3016 924 3029 938
rect 3044 924 3060 940
rect 3106 935 3117 948
rect 2899 890 2900 906
rect 2915 890 2928 912
rect 2943 890 2973 912
rect 3016 908 3078 924
rect 3106 917 3117 933
rect 3122 928 3132 948
rect 3142 928 3156 948
rect 3159 935 3168 948
rect 3184 935 3193 948
rect 3122 917 3156 928
rect 3159 917 3168 933
rect 3184 917 3193 933
rect 3200 928 3210 948
rect 3220 928 3234 948
rect 3235 935 3246 948
rect 3200 917 3234 928
rect 3235 917 3246 933
rect 3292 924 3308 940
rect 3315 938 3345 990
rect 3379 986 3380 993
rect 3364 978 3380 986
rect 3351 946 3364 965
rect 3379 946 3409 962
rect 3351 930 3425 946
rect 3351 928 3364 930
rect 3379 928 3413 930
rect 3016 906 3029 908
rect 3044 906 3078 908
rect 3016 890 3078 906
rect 3122 901 3138 904
rect 3200 901 3230 912
rect 3278 908 3324 924
rect 3351 912 3425 928
rect 3278 906 3312 908
rect 3277 890 3324 906
rect 3351 890 3364 912
rect 3379 890 3409 912
rect 3436 890 3437 906
rect 3452 890 3465 1050
rect 3495 946 3508 1050
rect 3553 1028 3554 1038
rect 3569 1028 3582 1038
rect 3553 1024 3582 1028
rect 3587 1024 3617 1050
rect 3635 1036 3651 1038
rect 3723 1036 3776 1050
rect 3724 1034 3788 1036
rect 3831 1034 3846 1050
rect 3895 1047 3925 1050
rect 3895 1044 3931 1047
rect 3861 1036 3877 1038
rect 3635 1024 3650 1028
rect 3553 1022 3650 1024
rect 3678 1022 3846 1034
rect 3862 1024 3877 1028
rect 3895 1025 3934 1044
rect 3953 1038 3960 1039
rect 3959 1031 3960 1038
rect 3943 1028 3944 1031
rect 3959 1028 3972 1031
rect 3895 1024 3925 1025
rect 3934 1024 3940 1025
rect 3943 1024 3972 1028
rect 3862 1023 3972 1024
rect 3862 1022 3978 1023
rect 3537 1014 3588 1022
rect 3537 1002 3562 1014
rect 3569 1002 3588 1014
rect 3619 1014 3669 1022
rect 3619 1006 3635 1014
rect 3642 1012 3669 1014
rect 3678 1012 3899 1022
rect 3642 1002 3899 1012
rect 3928 1014 3978 1022
rect 3928 1005 3944 1014
rect 3537 994 3588 1002
rect 3635 994 3899 1002
rect 3925 1002 3944 1005
rect 3951 1002 3978 1014
rect 3925 994 3978 1002
rect 3553 986 3554 994
rect 3569 986 3582 994
rect 3553 978 3569 986
rect 3550 971 3569 974
rect 3550 962 3572 971
rect 3523 952 3572 962
rect 3523 946 3553 952
rect 3572 947 3577 952
rect 3495 930 3569 946
rect 3587 938 3617 994
rect 3652 984 3860 994
rect 3895 990 3940 994
rect 3943 993 3944 994
rect 3959 993 3972 994
rect 3678 954 3867 984
rect 3693 951 3867 954
rect 3686 948 3867 951
rect 3495 928 3508 930
rect 3523 928 3557 930
rect 3495 912 3569 928
rect 3596 924 3609 938
rect 3624 924 3640 940
rect 3686 935 3697 948
rect 3479 890 3480 906
rect 3495 890 3508 912
rect 3523 890 3553 912
rect 3596 908 3658 924
rect 3686 917 3697 933
rect 3702 928 3712 948
rect 3722 928 3736 948
rect 3739 935 3748 948
rect 3764 935 3773 948
rect 3702 917 3736 928
rect 3739 917 3748 933
rect 3764 917 3773 933
rect 3780 928 3790 948
rect 3800 928 3814 948
rect 3815 935 3826 948
rect 3780 917 3814 928
rect 3815 917 3826 933
rect 3872 924 3888 940
rect 3895 938 3925 990
rect 3959 986 3960 993
rect 3944 978 3960 986
rect 3931 946 3944 965
rect 3959 946 3989 962
rect 3931 930 4005 946
rect 3931 928 3944 930
rect 3959 928 3993 930
rect 3596 906 3609 908
rect 3624 906 3658 908
rect 3596 890 3658 906
rect 3702 901 3718 904
rect 3780 901 3810 912
rect 3858 908 3904 924
rect 3931 912 4005 928
rect 3858 906 3892 908
rect 3857 890 3904 906
rect 3931 890 3944 912
rect 3959 890 3989 912
rect 4016 890 4017 906
rect 4032 890 4045 1050
rect 4075 946 4088 1050
rect 4133 1028 4134 1038
rect 4149 1028 4162 1038
rect 4133 1024 4162 1028
rect 4167 1024 4197 1050
rect 4215 1036 4231 1038
rect 4303 1036 4356 1050
rect 4304 1034 4368 1036
rect 4411 1034 4426 1050
rect 4475 1047 4505 1050
rect 4475 1044 4511 1047
rect 4441 1036 4457 1038
rect 4215 1024 4230 1028
rect 4133 1022 4230 1024
rect 4258 1022 4426 1034
rect 4442 1024 4457 1028
rect 4475 1025 4514 1044
rect 4533 1038 4540 1039
rect 4539 1031 4540 1038
rect 4523 1028 4524 1031
rect 4539 1028 4552 1031
rect 4475 1024 4505 1025
rect 4514 1024 4520 1025
rect 4523 1024 4552 1028
rect 4442 1023 4552 1024
rect 4442 1022 4558 1023
rect 4117 1014 4168 1022
rect 4117 1002 4142 1014
rect 4149 1002 4168 1014
rect 4199 1014 4249 1022
rect 4199 1006 4215 1014
rect 4222 1012 4249 1014
rect 4258 1012 4479 1022
rect 4222 1002 4479 1012
rect 4508 1014 4558 1022
rect 4508 1005 4524 1014
rect 4117 994 4168 1002
rect 4215 994 4479 1002
rect 4505 1002 4524 1005
rect 4531 1002 4558 1014
rect 4505 994 4558 1002
rect 4133 986 4134 994
rect 4149 986 4162 994
rect 4133 978 4149 986
rect 4130 971 4149 974
rect 4130 962 4152 971
rect 4103 952 4152 962
rect 4103 946 4133 952
rect 4152 947 4157 952
rect 4075 930 4149 946
rect 4167 938 4197 994
rect 4232 984 4440 994
rect 4475 990 4520 994
rect 4523 993 4524 994
rect 4539 993 4552 994
rect 4258 954 4447 984
rect 4273 951 4447 954
rect 4266 948 4447 951
rect 4075 928 4088 930
rect 4103 928 4137 930
rect 4075 912 4149 928
rect 4176 924 4189 938
rect 4204 924 4220 940
rect 4266 935 4277 948
rect 4059 890 4060 906
rect 4075 890 4088 912
rect 4103 890 4133 912
rect 4176 908 4238 924
rect 4266 917 4277 933
rect 4282 928 4292 948
rect 4302 928 4316 948
rect 4319 935 4328 948
rect 4344 935 4353 948
rect 4282 917 4316 928
rect 4319 917 4328 933
rect 4344 917 4353 933
rect 4360 928 4370 948
rect 4380 928 4394 948
rect 4395 935 4406 948
rect 4360 917 4394 928
rect 4395 917 4406 933
rect 4452 924 4468 940
rect 4475 938 4505 990
rect 4539 986 4540 993
rect 4524 978 4540 986
rect 4511 946 4524 965
rect 4539 946 4569 962
rect 4511 930 4585 946
rect 4511 928 4524 930
rect 4539 928 4573 930
rect 4176 906 4189 908
rect 4204 906 4238 908
rect 4176 890 4238 906
rect 4282 901 4298 904
rect 4360 901 4390 912
rect 4438 908 4484 924
rect 4511 912 4585 928
rect 4438 906 4472 908
rect 4437 890 4484 906
rect 4511 890 4524 912
rect 4539 890 4569 912
rect 4596 890 4597 906
rect 4612 890 4625 1050
rect -7 882 34 890
rect -7 856 8 882
rect 15 856 34 882
rect 98 878 160 890
rect 172 878 247 890
rect 305 878 380 890
rect 392 878 423 890
rect 429 878 464 890
rect 98 876 260 878
rect -7 848 34 856
rect 116 852 129 876
rect 144 874 159 876
rect -1 838 0 848
rect 15 838 28 848
rect 43 838 73 852
rect 116 838 159 852
rect 183 849 190 856
rect 193 852 260 876
rect 292 876 464 878
rect 262 854 290 858
rect 292 854 372 876
rect 393 874 408 876
rect 262 852 372 854
rect 193 848 372 852
rect 166 838 196 848
rect 198 838 351 848
rect 359 838 389 848
rect 393 838 423 852
rect 451 838 464 876
rect 536 882 571 890
rect 536 856 537 882
rect 544 856 571 882
rect 479 838 509 852
rect 536 848 571 856
rect 573 882 614 890
rect 573 856 588 882
rect 595 856 614 882
rect 678 878 740 890
rect 752 878 827 890
rect 885 878 960 890
rect 972 878 1003 890
rect 1009 878 1044 890
rect 678 876 840 878
rect 573 848 614 856
rect 696 852 709 876
rect 724 874 739 876
rect 536 838 537 848
rect 552 838 565 848
rect 579 838 580 848
rect 595 838 608 848
rect 623 838 653 852
rect 696 838 739 852
rect 763 849 770 856
rect 773 852 840 876
rect 872 876 1044 878
rect 842 854 870 858
rect 872 854 952 876
rect 973 874 988 876
rect 842 852 952 854
rect 773 848 952 852
rect 746 838 776 848
rect 778 838 931 848
rect 939 838 969 848
rect 973 838 1003 852
rect 1031 838 1044 876
rect 1116 882 1151 890
rect 1116 856 1117 882
rect 1124 856 1151 882
rect 1059 838 1089 852
rect 1116 848 1151 856
rect 1153 882 1194 890
rect 1153 856 1168 882
rect 1175 856 1194 882
rect 1258 878 1320 890
rect 1332 878 1407 890
rect 1465 878 1540 890
rect 1552 878 1583 890
rect 1589 878 1624 890
rect 1258 876 1420 878
rect 1153 848 1194 856
rect 1276 852 1289 876
rect 1304 874 1319 876
rect 1116 838 1117 848
rect 1132 838 1145 848
rect 1159 838 1160 848
rect 1175 838 1188 848
rect 1203 838 1233 852
rect 1276 838 1319 852
rect 1343 849 1350 856
rect 1353 852 1420 876
rect 1452 876 1624 878
rect 1422 854 1450 858
rect 1452 854 1532 876
rect 1553 874 1568 876
rect 1422 852 1532 854
rect 1353 848 1532 852
rect 1326 838 1356 848
rect 1358 838 1511 848
rect 1519 838 1549 848
rect 1553 838 1583 852
rect 1611 838 1624 876
rect 1696 882 1731 890
rect 1696 856 1697 882
rect 1704 856 1731 882
rect 1639 838 1669 852
rect 1696 848 1731 856
rect 1733 882 1774 890
rect 1733 856 1748 882
rect 1755 856 1774 882
rect 1838 878 1900 890
rect 1912 878 1987 890
rect 2045 878 2120 890
rect 2132 878 2163 890
rect 2169 878 2204 890
rect 1838 876 2000 878
rect 1733 848 1774 856
rect 1856 852 1869 876
rect 1884 874 1899 876
rect 1696 838 1697 848
rect 1712 838 1725 848
rect 1739 838 1740 848
rect 1755 838 1768 848
rect 1783 838 1813 852
rect 1856 838 1899 852
rect 1923 849 1930 856
rect 1933 852 2000 876
rect 2032 876 2204 878
rect 2002 854 2030 858
rect 2032 854 2112 876
rect 2133 874 2148 876
rect 2002 852 2112 854
rect 1933 848 2112 852
rect 1906 838 1936 848
rect 1938 838 2091 848
rect 2099 838 2129 848
rect 2133 838 2163 852
rect 2191 838 2204 876
rect 2276 882 2311 890
rect 2276 856 2277 882
rect 2284 856 2311 882
rect 2219 838 2249 852
rect 2276 848 2311 856
rect 2313 882 2354 890
rect 2313 856 2328 882
rect 2335 856 2354 882
rect 2418 878 2480 890
rect 2492 878 2567 890
rect 2625 878 2700 890
rect 2712 878 2743 890
rect 2749 878 2784 890
rect 2418 876 2580 878
rect 2313 848 2354 856
rect 2436 852 2449 876
rect 2464 874 2479 876
rect 2276 838 2277 848
rect 2292 838 2305 848
rect 2319 838 2320 848
rect 2335 838 2348 848
rect 2363 838 2393 852
rect 2436 838 2479 852
rect 2503 849 2510 856
rect 2513 852 2580 876
rect 2612 876 2784 878
rect 2582 854 2610 858
rect 2612 854 2692 876
rect 2713 874 2728 876
rect 2582 852 2692 854
rect 2513 848 2692 852
rect 2486 838 2516 848
rect 2518 838 2671 848
rect 2679 838 2709 848
rect 2713 838 2743 852
rect 2771 838 2784 876
rect 2856 882 2891 890
rect 2856 856 2857 882
rect 2864 856 2891 882
rect 2799 838 2829 852
rect 2856 848 2891 856
rect 2893 882 2934 890
rect 2893 856 2908 882
rect 2915 856 2934 882
rect 2998 878 3060 890
rect 3072 878 3147 890
rect 3205 878 3280 890
rect 3292 878 3323 890
rect 3329 878 3364 890
rect 2998 876 3160 878
rect 2893 848 2934 856
rect 3016 852 3029 876
rect 3044 874 3059 876
rect 2856 838 2857 848
rect 2872 838 2885 848
rect 2899 838 2900 848
rect 2915 838 2928 848
rect 2943 838 2973 852
rect 3016 838 3059 852
rect 3083 849 3090 856
rect 3093 852 3160 876
rect 3192 876 3364 878
rect 3162 854 3190 858
rect 3192 854 3272 876
rect 3293 874 3308 876
rect 3162 852 3272 854
rect 3093 848 3272 852
rect 3066 838 3096 848
rect 3098 838 3251 848
rect 3259 838 3289 848
rect 3293 838 3323 852
rect 3351 838 3364 876
rect 3436 882 3471 890
rect 3436 856 3437 882
rect 3444 856 3471 882
rect 3379 838 3409 852
rect 3436 848 3471 856
rect 3473 882 3514 890
rect 3473 856 3488 882
rect 3495 856 3514 882
rect 3578 878 3640 890
rect 3652 878 3727 890
rect 3785 878 3860 890
rect 3872 878 3903 890
rect 3909 878 3944 890
rect 3578 876 3740 878
rect 3473 848 3514 856
rect 3596 852 3609 876
rect 3624 874 3639 876
rect 3436 838 3437 848
rect 3452 838 3465 848
rect 3479 838 3480 848
rect 3495 838 3508 848
rect 3523 838 3553 852
rect 3596 838 3639 852
rect 3663 849 3670 856
rect 3673 852 3740 876
rect 3772 876 3944 878
rect 3742 854 3770 858
rect 3772 854 3852 876
rect 3873 874 3888 876
rect 3742 852 3852 854
rect 3673 848 3852 852
rect 3646 838 3676 848
rect 3678 838 3831 848
rect 3839 838 3869 848
rect 3873 838 3903 852
rect 3931 838 3944 876
rect 4016 882 4051 890
rect 4016 856 4017 882
rect 4024 856 4051 882
rect 3959 838 3989 852
rect 4016 848 4051 856
rect 4053 882 4094 890
rect 4053 856 4068 882
rect 4075 856 4094 882
rect 4158 878 4220 890
rect 4232 878 4307 890
rect 4365 878 4440 890
rect 4452 878 4483 890
rect 4489 878 4524 890
rect 4158 876 4320 878
rect 4053 848 4094 856
rect 4176 852 4189 876
rect 4204 874 4219 876
rect 4016 838 4017 848
rect 4032 838 4045 848
rect 4059 838 4060 848
rect 4075 838 4088 848
rect 4103 838 4133 852
rect 4176 838 4219 852
rect 4243 849 4250 856
rect 4253 852 4320 876
rect 4352 876 4524 878
rect 4322 854 4350 858
rect 4352 854 4432 876
rect 4453 874 4468 876
rect 4322 852 4432 854
rect 4253 848 4432 852
rect 4226 838 4256 848
rect 4258 838 4411 848
rect 4419 838 4449 848
rect 4453 838 4483 852
rect 4511 838 4524 876
rect 4596 882 4631 890
rect 4596 856 4597 882
rect 4604 856 4631 882
rect 4539 838 4569 852
rect 4596 848 4631 856
rect 4596 838 4597 848
rect 4612 838 4625 848
rect -1 832 4625 838
rect 0 824 4625 832
rect 15 794 28 824
rect 43 806 73 824
rect 116 810 130 824
rect 166 810 386 824
rect 117 808 130 810
rect 83 796 98 808
rect 80 794 102 796
rect 107 794 137 808
rect 198 806 351 810
rect 180 794 372 806
rect 415 794 445 808
rect 451 794 464 824
rect 479 806 509 824
rect 552 794 565 824
rect 595 794 608 824
rect 623 806 653 824
rect 696 810 710 824
rect 746 810 966 824
rect 697 808 710 810
rect 663 796 678 808
rect 660 794 682 796
rect 687 794 717 808
rect 778 806 931 810
rect 760 794 952 806
rect 995 794 1025 808
rect 1031 794 1044 824
rect 1059 806 1089 824
rect 1132 794 1145 824
rect 1175 794 1188 824
rect 1203 806 1233 824
rect 1276 810 1290 824
rect 1326 810 1546 824
rect 1277 808 1290 810
rect 1243 796 1258 808
rect 1240 794 1262 796
rect 1267 794 1297 808
rect 1358 806 1511 810
rect 1340 794 1532 806
rect 1575 794 1605 808
rect 1611 794 1624 824
rect 1639 806 1669 824
rect 1712 794 1725 824
rect 1755 794 1768 824
rect 1783 806 1813 824
rect 1856 810 1870 824
rect 1906 810 2126 824
rect 1857 808 1870 810
rect 1823 796 1838 808
rect 1820 794 1842 796
rect 1847 794 1877 808
rect 1938 806 2091 810
rect 1920 794 2112 806
rect 2155 794 2185 808
rect 2191 794 2204 824
rect 2219 806 2249 824
rect 2292 794 2305 824
rect 2335 794 2348 824
rect 2363 806 2393 824
rect 2436 810 2450 824
rect 2486 810 2706 824
rect 2437 808 2450 810
rect 2403 796 2418 808
rect 2400 794 2422 796
rect 2427 794 2457 808
rect 2518 806 2671 810
rect 2500 794 2692 806
rect 2735 794 2765 808
rect 2771 794 2784 824
rect 2799 806 2829 824
rect 2872 794 2885 824
rect 2915 794 2928 824
rect 2943 806 2973 824
rect 3016 810 3030 824
rect 3066 810 3286 824
rect 3017 808 3030 810
rect 2983 796 2998 808
rect 2980 794 3002 796
rect 3007 794 3037 808
rect 3098 806 3251 810
rect 3080 794 3272 806
rect 3315 794 3345 808
rect 3351 794 3364 824
rect 3379 806 3409 824
rect 3452 794 3465 824
rect 3495 794 3508 824
rect 3523 806 3553 824
rect 3596 810 3610 824
rect 3646 810 3866 824
rect 3597 808 3610 810
rect 3563 796 3578 808
rect 3560 794 3582 796
rect 3587 794 3617 808
rect 3678 806 3831 810
rect 3660 794 3852 806
rect 3895 794 3925 808
rect 3931 794 3944 824
rect 3959 806 3989 824
rect 4032 794 4045 824
rect 4075 794 4088 824
rect 4103 806 4133 824
rect 4176 810 4190 824
rect 4226 810 4446 824
rect 4177 808 4190 810
rect 4143 796 4158 808
rect 4140 794 4162 796
rect 4167 794 4197 808
rect 4258 806 4411 810
rect 4240 794 4432 806
rect 4475 794 4505 808
rect 4511 794 4524 824
rect 4539 806 4569 824
rect 4612 794 4625 824
rect 0 780 4625 794
rect 15 676 28 780
rect 73 758 74 768
rect 89 758 102 768
rect 73 754 102 758
rect 107 754 137 780
rect 155 766 171 768
rect 243 766 296 780
rect 244 764 308 766
rect 351 764 366 780
rect 415 777 445 780
rect 415 774 451 777
rect 381 766 397 768
rect 155 754 170 758
rect 73 752 170 754
rect 198 752 366 764
rect 382 754 397 758
rect 415 755 454 774
rect 473 768 480 769
rect 479 761 480 768
rect 463 758 464 761
rect 479 758 492 761
rect 415 754 445 755
rect 454 754 460 755
rect 463 754 492 758
rect 382 753 492 754
rect 382 752 498 753
rect 57 744 108 752
rect 57 732 82 744
rect 89 732 108 744
rect 139 744 189 752
rect 139 736 155 744
rect 162 742 189 744
rect 198 742 419 752
rect 162 732 419 742
rect 448 744 498 752
rect 448 735 464 744
rect 57 724 108 732
rect 155 724 419 732
rect 445 732 464 735
rect 471 732 498 744
rect 445 724 498 732
rect 73 716 74 724
rect 89 716 102 724
rect 73 708 89 716
rect 70 701 89 704
rect 70 692 92 701
rect 43 682 92 692
rect 43 676 73 682
rect 92 677 97 682
rect 15 660 89 676
rect 107 668 137 724
rect 172 714 380 724
rect 415 720 460 724
rect 463 723 464 724
rect 479 723 492 724
rect 198 684 387 714
rect 213 681 387 684
rect 206 678 387 681
rect 15 658 28 660
rect 43 658 77 660
rect 15 642 89 658
rect 116 654 129 668
rect 144 654 160 670
rect 206 665 217 678
rect -1 620 0 636
rect 15 620 28 642
rect 43 620 73 642
rect 116 638 178 654
rect 206 647 217 663
rect 222 658 232 678
rect 242 658 256 678
rect 259 665 268 678
rect 284 665 293 678
rect 222 647 256 658
rect 259 647 268 663
rect 284 647 293 663
rect 300 658 310 678
rect 320 658 334 678
rect 335 665 346 678
rect 300 647 334 658
rect 335 647 346 663
rect 392 654 408 670
rect 415 668 445 720
rect 479 716 480 723
rect 464 708 480 716
rect 451 676 464 695
rect 479 676 509 692
rect 451 660 525 676
rect 451 658 464 660
rect 479 658 513 660
rect 116 636 129 638
rect 144 636 178 638
rect 116 620 178 636
rect 222 631 238 634
rect 300 631 330 642
rect 378 638 424 654
rect 451 642 525 658
rect 378 636 412 638
rect 377 620 424 636
rect 451 620 464 642
rect 479 620 509 642
rect 536 620 537 636
rect 552 620 565 780
rect 595 676 608 780
rect 653 758 654 768
rect 669 758 682 768
rect 653 754 682 758
rect 687 754 717 780
rect 735 766 751 768
rect 823 766 876 780
rect 824 764 888 766
rect 931 764 946 780
rect 995 777 1025 780
rect 995 774 1031 777
rect 961 766 977 768
rect 735 754 750 758
rect 653 752 750 754
rect 778 752 946 764
rect 962 754 977 758
rect 995 755 1034 774
rect 1053 768 1060 769
rect 1059 761 1060 768
rect 1043 758 1044 761
rect 1059 758 1072 761
rect 995 754 1025 755
rect 1034 754 1040 755
rect 1043 754 1072 758
rect 962 753 1072 754
rect 962 752 1078 753
rect 637 744 688 752
rect 637 732 662 744
rect 669 732 688 744
rect 719 744 769 752
rect 719 736 735 744
rect 742 742 769 744
rect 778 742 999 752
rect 742 732 999 742
rect 1028 744 1078 752
rect 1028 735 1044 744
rect 637 724 688 732
rect 735 724 999 732
rect 1025 732 1044 735
rect 1051 732 1078 744
rect 1025 724 1078 732
rect 653 716 654 724
rect 669 716 682 724
rect 653 708 669 716
rect 650 701 669 704
rect 650 692 672 701
rect 623 682 672 692
rect 623 676 653 682
rect 672 677 677 682
rect 595 660 669 676
rect 687 668 717 724
rect 752 714 960 724
rect 995 720 1040 724
rect 1043 723 1044 724
rect 1059 723 1072 724
rect 778 684 967 714
rect 793 681 967 684
rect 786 678 967 681
rect 595 658 608 660
rect 623 658 657 660
rect 595 642 669 658
rect 696 654 709 668
rect 724 654 740 670
rect 786 665 797 678
rect 579 620 580 636
rect 595 620 608 642
rect 623 620 653 642
rect 696 638 758 654
rect 786 647 797 663
rect 802 658 812 678
rect 822 658 836 678
rect 839 665 848 678
rect 864 665 873 678
rect 802 647 836 658
rect 839 647 848 663
rect 864 647 873 663
rect 880 658 890 678
rect 900 658 914 678
rect 915 665 926 678
rect 880 647 914 658
rect 915 647 926 663
rect 972 654 988 670
rect 995 668 1025 720
rect 1059 716 1060 723
rect 1044 708 1060 716
rect 1031 676 1044 695
rect 1059 676 1089 692
rect 1031 660 1105 676
rect 1031 658 1044 660
rect 1059 658 1093 660
rect 696 636 709 638
rect 724 636 758 638
rect 696 620 758 636
rect 802 631 818 634
rect 880 631 910 642
rect 958 638 1004 654
rect 1031 642 1105 658
rect 958 636 992 638
rect 957 620 1004 636
rect 1031 620 1044 642
rect 1059 620 1089 642
rect 1116 620 1117 636
rect 1132 620 1145 780
rect 1175 676 1188 780
rect 1233 758 1234 768
rect 1249 758 1262 768
rect 1233 754 1262 758
rect 1267 754 1297 780
rect 1315 766 1331 768
rect 1403 766 1456 780
rect 1404 764 1468 766
rect 1511 764 1526 780
rect 1575 777 1605 780
rect 1575 774 1611 777
rect 1541 766 1557 768
rect 1315 754 1330 758
rect 1233 752 1330 754
rect 1358 752 1526 764
rect 1542 754 1557 758
rect 1575 755 1614 774
rect 1633 768 1640 769
rect 1639 761 1640 768
rect 1623 758 1624 761
rect 1639 758 1652 761
rect 1575 754 1605 755
rect 1614 754 1620 755
rect 1623 754 1652 758
rect 1542 753 1652 754
rect 1542 752 1658 753
rect 1217 744 1268 752
rect 1217 732 1242 744
rect 1249 732 1268 744
rect 1299 744 1349 752
rect 1299 736 1315 744
rect 1322 742 1349 744
rect 1358 742 1579 752
rect 1322 732 1579 742
rect 1608 744 1658 752
rect 1608 735 1624 744
rect 1217 724 1268 732
rect 1315 724 1579 732
rect 1605 732 1624 735
rect 1631 732 1658 744
rect 1605 724 1658 732
rect 1233 716 1234 724
rect 1249 716 1262 724
rect 1233 708 1249 716
rect 1230 701 1249 704
rect 1230 692 1252 701
rect 1203 682 1252 692
rect 1203 676 1233 682
rect 1252 677 1257 682
rect 1175 660 1249 676
rect 1267 668 1297 724
rect 1332 714 1540 724
rect 1575 720 1620 724
rect 1623 723 1624 724
rect 1639 723 1652 724
rect 1358 684 1547 714
rect 1373 681 1547 684
rect 1366 678 1547 681
rect 1175 658 1188 660
rect 1203 658 1237 660
rect 1175 642 1249 658
rect 1276 654 1289 668
rect 1304 654 1320 670
rect 1366 665 1377 678
rect 1159 620 1160 636
rect 1175 620 1188 642
rect 1203 620 1233 642
rect 1276 638 1338 654
rect 1366 647 1377 663
rect 1382 658 1392 678
rect 1402 658 1416 678
rect 1419 665 1428 678
rect 1444 665 1453 678
rect 1382 647 1416 658
rect 1419 647 1428 663
rect 1444 647 1453 663
rect 1460 658 1470 678
rect 1480 658 1494 678
rect 1495 665 1506 678
rect 1460 647 1494 658
rect 1495 647 1506 663
rect 1552 654 1568 670
rect 1575 668 1605 720
rect 1639 716 1640 723
rect 1624 708 1640 716
rect 1611 676 1624 695
rect 1639 676 1669 692
rect 1611 660 1685 676
rect 1611 658 1624 660
rect 1639 658 1673 660
rect 1276 636 1289 638
rect 1304 636 1338 638
rect 1276 620 1338 636
rect 1382 631 1398 634
rect 1460 631 1490 642
rect 1538 638 1584 654
rect 1611 642 1685 658
rect 1538 636 1572 638
rect 1537 620 1584 636
rect 1611 620 1624 642
rect 1639 620 1669 642
rect 1696 620 1697 636
rect 1712 620 1725 780
rect 1755 676 1768 780
rect 1813 758 1814 768
rect 1829 758 1842 768
rect 1813 754 1842 758
rect 1847 754 1877 780
rect 1895 766 1911 768
rect 1983 766 2036 780
rect 1984 764 2048 766
rect 2091 764 2106 780
rect 2155 777 2185 780
rect 2155 774 2191 777
rect 2121 766 2137 768
rect 1895 754 1910 758
rect 1813 752 1910 754
rect 1938 752 2106 764
rect 2122 754 2137 758
rect 2155 755 2194 774
rect 2213 768 2220 769
rect 2219 761 2220 768
rect 2203 758 2204 761
rect 2219 758 2232 761
rect 2155 754 2185 755
rect 2194 754 2200 755
rect 2203 754 2232 758
rect 2122 753 2232 754
rect 2122 752 2238 753
rect 1797 744 1848 752
rect 1797 732 1822 744
rect 1829 732 1848 744
rect 1879 744 1929 752
rect 1879 736 1895 744
rect 1902 742 1929 744
rect 1938 742 2159 752
rect 1902 732 2159 742
rect 2188 744 2238 752
rect 2188 735 2204 744
rect 1797 724 1848 732
rect 1895 724 2159 732
rect 2185 732 2204 735
rect 2211 732 2238 744
rect 2185 724 2238 732
rect 1813 716 1814 724
rect 1829 716 1842 724
rect 1813 708 1829 716
rect 1810 701 1829 704
rect 1810 692 1832 701
rect 1783 682 1832 692
rect 1783 676 1813 682
rect 1832 677 1837 682
rect 1755 660 1829 676
rect 1847 668 1877 724
rect 1912 714 2120 724
rect 2155 720 2200 724
rect 2203 723 2204 724
rect 2219 723 2232 724
rect 1938 684 2127 714
rect 1953 681 2127 684
rect 1946 678 2127 681
rect 1755 658 1768 660
rect 1783 658 1817 660
rect 1755 642 1829 658
rect 1856 654 1869 668
rect 1884 654 1900 670
rect 1946 665 1957 678
rect 1739 620 1740 636
rect 1755 620 1768 642
rect 1783 620 1813 642
rect 1856 638 1918 654
rect 1946 647 1957 663
rect 1962 658 1972 678
rect 1982 658 1996 678
rect 1999 665 2008 678
rect 2024 665 2033 678
rect 1962 647 1996 658
rect 1999 647 2008 663
rect 2024 647 2033 663
rect 2040 658 2050 678
rect 2060 658 2074 678
rect 2075 665 2086 678
rect 2040 647 2074 658
rect 2075 647 2086 663
rect 2132 654 2148 670
rect 2155 668 2185 720
rect 2219 716 2220 723
rect 2204 708 2220 716
rect 2191 676 2204 695
rect 2219 676 2249 692
rect 2191 660 2265 676
rect 2191 658 2204 660
rect 2219 658 2253 660
rect 1856 636 1869 638
rect 1884 636 1918 638
rect 1856 620 1918 636
rect 1962 631 1978 634
rect 2040 631 2070 642
rect 2118 638 2164 654
rect 2191 642 2265 658
rect 2118 636 2152 638
rect 2117 620 2164 636
rect 2191 620 2204 642
rect 2219 620 2249 642
rect 2276 620 2277 636
rect 2292 620 2305 780
rect 2335 676 2348 780
rect 2393 758 2394 768
rect 2409 758 2422 768
rect 2393 754 2422 758
rect 2427 754 2457 780
rect 2475 766 2491 768
rect 2563 766 2616 780
rect 2564 764 2628 766
rect 2671 764 2686 780
rect 2735 777 2765 780
rect 2735 774 2771 777
rect 2701 766 2717 768
rect 2475 754 2490 758
rect 2393 752 2490 754
rect 2518 752 2686 764
rect 2702 754 2717 758
rect 2735 755 2774 774
rect 2793 768 2800 769
rect 2799 761 2800 768
rect 2783 758 2784 761
rect 2799 758 2812 761
rect 2735 754 2765 755
rect 2774 754 2780 755
rect 2783 754 2812 758
rect 2702 753 2812 754
rect 2702 752 2818 753
rect 2377 744 2428 752
rect 2377 732 2402 744
rect 2409 732 2428 744
rect 2459 744 2509 752
rect 2459 736 2475 744
rect 2482 742 2509 744
rect 2518 742 2739 752
rect 2482 732 2739 742
rect 2768 744 2818 752
rect 2768 735 2784 744
rect 2377 724 2428 732
rect 2475 724 2739 732
rect 2765 732 2784 735
rect 2791 732 2818 744
rect 2765 724 2818 732
rect 2393 716 2394 724
rect 2409 716 2422 724
rect 2393 708 2409 716
rect 2390 701 2409 704
rect 2390 692 2412 701
rect 2363 682 2412 692
rect 2363 676 2393 682
rect 2412 677 2417 682
rect 2335 660 2409 676
rect 2427 668 2457 724
rect 2492 714 2700 724
rect 2735 720 2780 724
rect 2783 723 2784 724
rect 2799 723 2812 724
rect 2518 684 2707 714
rect 2533 681 2707 684
rect 2526 678 2707 681
rect 2335 658 2348 660
rect 2363 658 2397 660
rect 2335 642 2409 658
rect 2436 654 2449 668
rect 2464 654 2480 670
rect 2526 665 2537 678
rect 2319 620 2320 636
rect 2335 620 2348 642
rect 2363 620 2393 642
rect 2436 638 2498 654
rect 2526 647 2537 663
rect 2542 658 2552 678
rect 2562 658 2576 678
rect 2579 665 2588 678
rect 2604 665 2613 678
rect 2542 647 2576 658
rect 2579 647 2588 663
rect 2604 647 2613 663
rect 2620 658 2630 678
rect 2640 658 2654 678
rect 2655 665 2666 678
rect 2620 647 2654 658
rect 2655 647 2666 663
rect 2712 654 2728 670
rect 2735 668 2765 720
rect 2799 716 2800 723
rect 2784 708 2800 716
rect 2771 676 2784 695
rect 2799 676 2829 692
rect 2771 660 2845 676
rect 2771 658 2784 660
rect 2799 658 2833 660
rect 2436 636 2449 638
rect 2464 636 2498 638
rect 2436 620 2498 636
rect 2542 631 2558 634
rect 2620 631 2650 642
rect 2698 638 2744 654
rect 2771 642 2845 658
rect 2698 636 2732 638
rect 2697 620 2744 636
rect 2771 620 2784 642
rect 2799 620 2829 642
rect 2856 620 2857 636
rect 2872 620 2885 780
rect 2915 676 2928 780
rect 2973 758 2974 768
rect 2989 758 3002 768
rect 2973 754 3002 758
rect 3007 754 3037 780
rect 3055 766 3071 768
rect 3143 766 3196 780
rect 3144 764 3208 766
rect 3251 764 3266 780
rect 3315 777 3345 780
rect 3315 774 3351 777
rect 3281 766 3297 768
rect 3055 754 3070 758
rect 2973 752 3070 754
rect 3098 752 3266 764
rect 3282 754 3297 758
rect 3315 755 3354 774
rect 3373 768 3380 769
rect 3379 761 3380 768
rect 3363 758 3364 761
rect 3379 758 3392 761
rect 3315 754 3345 755
rect 3354 754 3360 755
rect 3363 754 3392 758
rect 3282 753 3392 754
rect 3282 752 3398 753
rect 2957 744 3008 752
rect 2957 732 2982 744
rect 2989 732 3008 744
rect 3039 744 3089 752
rect 3039 736 3055 744
rect 3062 742 3089 744
rect 3098 742 3319 752
rect 3062 732 3319 742
rect 3348 744 3398 752
rect 3348 735 3364 744
rect 2957 724 3008 732
rect 3055 724 3319 732
rect 3345 732 3364 735
rect 3371 732 3398 744
rect 3345 724 3398 732
rect 2973 716 2974 724
rect 2989 716 3002 724
rect 2973 708 2989 716
rect 2970 701 2989 704
rect 2970 692 2992 701
rect 2943 682 2992 692
rect 2943 676 2973 682
rect 2992 677 2997 682
rect 2915 660 2989 676
rect 3007 668 3037 724
rect 3072 714 3280 724
rect 3315 720 3360 724
rect 3363 723 3364 724
rect 3379 723 3392 724
rect 3098 684 3287 714
rect 3113 681 3287 684
rect 3106 678 3287 681
rect 2915 658 2928 660
rect 2943 658 2977 660
rect 2915 642 2989 658
rect 3016 654 3029 668
rect 3044 654 3060 670
rect 3106 665 3117 678
rect 2899 620 2900 636
rect 2915 620 2928 642
rect 2943 620 2973 642
rect 3016 638 3078 654
rect 3106 647 3117 663
rect 3122 658 3132 678
rect 3142 658 3156 678
rect 3159 665 3168 678
rect 3184 665 3193 678
rect 3122 647 3156 658
rect 3159 647 3168 663
rect 3184 647 3193 663
rect 3200 658 3210 678
rect 3220 658 3234 678
rect 3235 665 3246 678
rect 3200 647 3234 658
rect 3235 647 3246 663
rect 3292 654 3308 670
rect 3315 668 3345 720
rect 3379 716 3380 723
rect 3364 708 3380 716
rect 3351 676 3364 695
rect 3379 676 3409 692
rect 3351 660 3425 676
rect 3351 658 3364 660
rect 3379 658 3413 660
rect 3016 636 3029 638
rect 3044 636 3078 638
rect 3016 620 3078 636
rect 3122 631 3138 634
rect 3200 631 3230 642
rect 3278 638 3324 654
rect 3351 642 3425 658
rect 3278 636 3312 638
rect 3277 620 3324 636
rect 3351 620 3364 642
rect 3379 620 3409 642
rect 3436 620 3437 636
rect 3452 620 3465 780
rect 3495 676 3508 780
rect 3553 758 3554 768
rect 3569 758 3582 768
rect 3553 754 3582 758
rect 3587 754 3617 780
rect 3635 766 3651 768
rect 3723 766 3776 780
rect 3724 764 3788 766
rect 3831 764 3846 780
rect 3895 777 3925 780
rect 3895 774 3931 777
rect 3861 766 3877 768
rect 3635 754 3650 758
rect 3553 752 3650 754
rect 3678 752 3846 764
rect 3862 754 3877 758
rect 3895 755 3934 774
rect 3953 768 3960 769
rect 3959 761 3960 768
rect 3943 758 3944 761
rect 3959 758 3972 761
rect 3895 754 3925 755
rect 3934 754 3940 755
rect 3943 754 3972 758
rect 3862 753 3972 754
rect 3862 752 3978 753
rect 3537 744 3588 752
rect 3537 732 3562 744
rect 3569 732 3588 744
rect 3619 744 3669 752
rect 3619 736 3635 744
rect 3642 742 3669 744
rect 3678 742 3899 752
rect 3642 732 3899 742
rect 3928 744 3978 752
rect 3928 735 3944 744
rect 3537 724 3588 732
rect 3635 724 3899 732
rect 3925 732 3944 735
rect 3951 732 3978 744
rect 3925 724 3978 732
rect 3553 716 3554 724
rect 3569 716 3582 724
rect 3553 708 3569 716
rect 3550 701 3569 704
rect 3550 692 3572 701
rect 3523 682 3572 692
rect 3523 676 3553 682
rect 3572 677 3577 682
rect 3495 660 3569 676
rect 3587 668 3617 724
rect 3652 714 3860 724
rect 3895 720 3940 724
rect 3943 723 3944 724
rect 3959 723 3972 724
rect 3678 684 3867 714
rect 3693 681 3867 684
rect 3686 678 3867 681
rect 3495 658 3508 660
rect 3523 658 3557 660
rect 3495 642 3569 658
rect 3596 654 3609 668
rect 3624 654 3640 670
rect 3686 665 3697 678
rect 3479 620 3480 636
rect 3495 620 3508 642
rect 3523 620 3553 642
rect 3596 638 3658 654
rect 3686 647 3697 663
rect 3702 658 3712 678
rect 3722 658 3736 678
rect 3739 665 3748 678
rect 3764 665 3773 678
rect 3702 647 3736 658
rect 3739 647 3748 663
rect 3764 647 3773 663
rect 3780 658 3790 678
rect 3800 658 3814 678
rect 3815 665 3826 678
rect 3780 647 3814 658
rect 3815 647 3826 663
rect 3872 654 3888 670
rect 3895 668 3925 720
rect 3959 716 3960 723
rect 3944 708 3960 716
rect 3931 676 3944 695
rect 3959 676 3989 692
rect 3931 660 4005 676
rect 3931 658 3944 660
rect 3959 658 3993 660
rect 3596 636 3609 638
rect 3624 636 3658 638
rect 3596 620 3658 636
rect 3702 631 3718 634
rect 3780 631 3810 642
rect 3858 638 3904 654
rect 3931 642 4005 658
rect 3858 636 3892 638
rect 3857 620 3904 636
rect 3931 620 3944 642
rect 3959 620 3989 642
rect 4016 620 4017 636
rect 4032 620 4045 780
rect 4075 676 4088 780
rect 4133 758 4134 768
rect 4149 758 4162 768
rect 4133 754 4162 758
rect 4167 754 4197 780
rect 4215 766 4231 768
rect 4303 766 4356 780
rect 4304 764 4368 766
rect 4411 764 4426 780
rect 4475 777 4505 780
rect 4475 774 4511 777
rect 4441 766 4457 768
rect 4215 754 4230 758
rect 4133 752 4230 754
rect 4258 752 4426 764
rect 4442 754 4457 758
rect 4475 755 4514 774
rect 4533 768 4540 769
rect 4539 761 4540 768
rect 4523 758 4524 761
rect 4539 758 4552 761
rect 4475 754 4505 755
rect 4514 754 4520 755
rect 4523 754 4552 758
rect 4442 753 4552 754
rect 4442 752 4558 753
rect 4117 744 4168 752
rect 4117 732 4142 744
rect 4149 732 4168 744
rect 4199 744 4249 752
rect 4199 736 4215 744
rect 4222 742 4249 744
rect 4258 742 4479 752
rect 4222 732 4479 742
rect 4508 744 4558 752
rect 4508 735 4524 744
rect 4117 724 4168 732
rect 4215 724 4479 732
rect 4505 732 4524 735
rect 4531 732 4558 744
rect 4505 724 4558 732
rect 4133 716 4134 724
rect 4149 716 4162 724
rect 4133 708 4149 716
rect 4130 701 4149 704
rect 4130 692 4152 701
rect 4103 682 4152 692
rect 4103 676 4133 682
rect 4152 677 4157 682
rect 4075 660 4149 676
rect 4167 668 4197 724
rect 4232 714 4440 724
rect 4475 720 4520 724
rect 4523 723 4524 724
rect 4539 723 4552 724
rect 4258 684 4447 714
rect 4273 681 4447 684
rect 4266 678 4447 681
rect 4075 658 4088 660
rect 4103 658 4137 660
rect 4075 642 4149 658
rect 4176 654 4189 668
rect 4204 654 4220 670
rect 4266 665 4277 678
rect 4059 620 4060 636
rect 4075 620 4088 642
rect 4103 620 4133 642
rect 4176 638 4238 654
rect 4266 647 4277 663
rect 4282 658 4292 678
rect 4302 658 4316 678
rect 4319 665 4328 678
rect 4344 665 4353 678
rect 4282 647 4316 658
rect 4319 647 4328 663
rect 4344 647 4353 663
rect 4360 658 4370 678
rect 4380 658 4394 678
rect 4395 665 4406 678
rect 4360 647 4394 658
rect 4395 647 4406 663
rect 4452 654 4468 670
rect 4475 668 4505 720
rect 4539 716 4540 723
rect 4524 708 4540 716
rect 4511 676 4524 695
rect 4539 676 4569 692
rect 4511 660 4585 676
rect 4511 658 4524 660
rect 4539 658 4573 660
rect 4176 636 4189 638
rect 4204 636 4238 638
rect 4176 620 4238 636
rect 4282 631 4298 634
rect 4360 631 4390 642
rect 4438 638 4484 654
rect 4511 642 4585 658
rect 4438 636 4472 638
rect 4437 620 4484 636
rect 4511 620 4524 642
rect 4539 620 4569 642
rect 4596 620 4597 636
rect 4612 620 4625 780
rect -7 612 34 620
rect -7 586 8 612
rect 15 586 34 612
rect 98 608 160 620
rect 172 608 247 620
rect 305 608 380 620
rect 392 608 423 620
rect 429 608 464 620
rect 98 606 260 608
rect -7 578 34 586
rect 116 582 129 606
rect 144 604 159 606
rect -1 568 0 578
rect 15 568 28 578
rect 43 568 73 582
rect 116 568 159 582
rect 183 579 190 586
rect 193 582 260 606
rect 292 606 464 608
rect 262 584 290 588
rect 292 584 372 606
rect 393 604 408 606
rect 262 582 372 584
rect 193 578 372 582
rect 166 568 196 578
rect 198 568 351 578
rect 359 568 389 578
rect 393 568 423 582
rect 451 568 464 606
rect 536 612 571 620
rect 536 586 537 612
rect 544 586 571 612
rect 479 568 509 582
rect 536 578 571 586
rect 573 612 614 620
rect 573 586 588 612
rect 595 586 614 612
rect 678 608 740 620
rect 752 608 827 620
rect 885 608 960 620
rect 972 608 1003 620
rect 1009 608 1044 620
rect 678 606 840 608
rect 573 578 614 586
rect 696 582 709 606
rect 724 604 739 606
rect 536 568 537 578
rect 552 568 565 578
rect 579 568 580 578
rect 595 568 608 578
rect 623 568 653 582
rect 696 568 739 582
rect 763 579 770 586
rect 773 582 840 606
rect 872 606 1044 608
rect 842 584 870 588
rect 872 584 952 606
rect 973 604 988 606
rect 842 582 952 584
rect 773 578 952 582
rect 746 568 776 578
rect 778 568 931 578
rect 939 568 969 578
rect 973 568 1003 582
rect 1031 568 1044 606
rect 1116 612 1151 620
rect 1116 586 1117 612
rect 1124 586 1151 612
rect 1059 568 1089 582
rect 1116 578 1151 586
rect 1153 612 1194 620
rect 1153 586 1168 612
rect 1175 586 1194 612
rect 1258 608 1320 620
rect 1332 608 1407 620
rect 1465 608 1540 620
rect 1552 608 1583 620
rect 1589 608 1624 620
rect 1258 606 1420 608
rect 1153 578 1194 586
rect 1276 582 1289 606
rect 1304 604 1319 606
rect 1116 568 1117 578
rect 1132 568 1145 578
rect 1159 568 1160 578
rect 1175 568 1188 578
rect 1203 568 1233 582
rect 1276 568 1319 582
rect 1343 579 1350 586
rect 1353 582 1420 606
rect 1452 606 1624 608
rect 1422 584 1450 588
rect 1452 584 1532 606
rect 1553 604 1568 606
rect 1422 582 1532 584
rect 1353 578 1532 582
rect 1326 568 1356 578
rect 1358 568 1511 578
rect 1519 568 1549 578
rect 1553 568 1583 582
rect 1611 568 1624 606
rect 1696 612 1731 620
rect 1696 586 1697 612
rect 1704 586 1731 612
rect 1639 568 1669 582
rect 1696 578 1731 586
rect 1733 612 1774 620
rect 1733 586 1748 612
rect 1755 586 1774 612
rect 1838 608 1900 620
rect 1912 608 1987 620
rect 2045 608 2120 620
rect 2132 608 2163 620
rect 2169 608 2204 620
rect 1838 606 2000 608
rect 1733 578 1774 586
rect 1856 582 1869 606
rect 1884 604 1899 606
rect 1696 568 1697 578
rect 1712 568 1725 578
rect 1739 568 1740 578
rect 1755 568 1768 578
rect 1783 568 1813 582
rect 1856 568 1899 582
rect 1923 579 1930 586
rect 1933 582 2000 606
rect 2032 606 2204 608
rect 2002 584 2030 588
rect 2032 584 2112 606
rect 2133 604 2148 606
rect 2002 582 2112 584
rect 1933 578 2112 582
rect 1906 568 1936 578
rect 1938 568 2091 578
rect 2099 568 2129 578
rect 2133 568 2163 582
rect 2191 568 2204 606
rect 2276 612 2311 620
rect 2276 586 2277 612
rect 2284 586 2311 612
rect 2219 568 2249 582
rect 2276 578 2311 586
rect 2313 612 2354 620
rect 2313 586 2328 612
rect 2335 586 2354 612
rect 2418 608 2480 620
rect 2492 608 2567 620
rect 2625 608 2700 620
rect 2712 608 2743 620
rect 2749 608 2784 620
rect 2418 606 2580 608
rect 2313 578 2354 586
rect 2436 582 2449 606
rect 2464 604 2479 606
rect 2276 568 2277 578
rect 2292 568 2305 578
rect 2319 568 2320 578
rect 2335 568 2348 578
rect 2363 568 2393 582
rect 2436 568 2479 582
rect 2503 579 2510 586
rect 2513 582 2580 606
rect 2612 606 2784 608
rect 2582 584 2610 588
rect 2612 584 2692 606
rect 2713 604 2728 606
rect 2582 582 2692 584
rect 2513 578 2692 582
rect 2486 568 2516 578
rect 2518 568 2671 578
rect 2679 568 2709 578
rect 2713 568 2743 582
rect 2771 568 2784 606
rect 2856 612 2891 620
rect 2856 586 2857 612
rect 2864 586 2891 612
rect 2799 568 2829 582
rect 2856 578 2891 586
rect 2893 612 2934 620
rect 2893 586 2908 612
rect 2915 586 2934 612
rect 2998 608 3060 620
rect 3072 608 3147 620
rect 3205 608 3280 620
rect 3292 608 3323 620
rect 3329 608 3364 620
rect 2998 606 3160 608
rect 2893 578 2934 586
rect 3016 582 3029 606
rect 3044 604 3059 606
rect 2856 568 2857 578
rect 2872 568 2885 578
rect 2899 568 2900 578
rect 2915 568 2928 578
rect 2943 568 2973 582
rect 3016 568 3059 582
rect 3083 579 3090 586
rect 3093 582 3160 606
rect 3192 606 3364 608
rect 3162 584 3190 588
rect 3192 584 3272 606
rect 3293 604 3308 606
rect 3162 582 3272 584
rect 3093 578 3272 582
rect 3066 568 3096 578
rect 3098 568 3251 578
rect 3259 568 3289 578
rect 3293 568 3323 582
rect 3351 568 3364 606
rect 3436 612 3471 620
rect 3436 586 3437 612
rect 3444 586 3471 612
rect 3379 568 3409 582
rect 3436 578 3471 586
rect 3473 612 3514 620
rect 3473 586 3488 612
rect 3495 586 3514 612
rect 3578 608 3640 620
rect 3652 608 3727 620
rect 3785 608 3860 620
rect 3872 608 3903 620
rect 3909 608 3944 620
rect 3578 606 3740 608
rect 3473 578 3514 586
rect 3596 582 3609 606
rect 3624 604 3639 606
rect 3436 568 3437 578
rect 3452 568 3465 578
rect 3479 568 3480 578
rect 3495 568 3508 578
rect 3523 568 3553 582
rect 3596 568 3639 582
rect 3663 579 3670 586
rect 3673 582 3740 606
rect 3772 606 3944 608
rect 3742 584 3770 588
rect 3772 584 3852 606
rect 3873 604 3888 606
rect 3742 582 3852 584
rect 3673 578 3852 582
rect 3646 568 3676 578
rect 3678 568 3831 578
rect 3839 568 3869 578
rect 3873 568 3903 582
rect 3931 568 3944 606
rect 4016 612 4051 620
rect 4016 586 4017 612
rect 4024 586 4051 612
rect 3959 568 3989 582
rect 4016 578 4051 586
rect 4053 612 4094 620
rect 4053 586 4068 612
rect 4075 586 4094 612
rect 4158 608 4220 620
rect 4232 608 4307 620
rect 4365 608 4440 620
rect 4452 608 4483 620
rect 4489 608 4524 620
rect 4158 606 4320 608
rect 4053 578 4094 586
rect 4176 582 4189 606
rect 4204 604 4219 606
rect 4016 568 4017 578
rect 4032 568 4045 578
rect 4059 568 4060 578
rect 4075 568 4088 578
rect 4103 568 4133 582
rect 4176 568 4219 582
rect 4243 579 4250 586
rect 4253 582 4320 606
rect 4352 606 4524 608
rect 4322 584 4350 588
rect 4352 584 4432 606
rect 4453 604 4468 606
rect 4322 582 4432 584
rect 4253 578 4432 582
rect 4226 568 4256 578
rect 4258 568 4411 578
rect 4419 568 4449 578
rect 4453 568 4483 582
rect 4511 568 4524 606
rect 4596 612 4631 620
rect 4596 586 4597 612
rect 4604 586 4631 612
rect 4539 568 4569 582
rect 4596 578 4631 586
rect 4596 568 4597 578
rect 4612 568 4625 578
rect -1 562 4625 568
rect 0 554 4625 562
rect 15 524 28 554
rect 43 536 73 554
rect 116 540 130 554
rect 166 540 386 554
rect 117 538 130 540
rect 83 526 98 538
rect 80 524 102 526
rect 107 524 137 538
rect 198 536 351 540
rect 180 524 372 536
rect 415 524 445 538
rect 451 524 464 554
rect 479 536 509 554
rect 552 524 565 554
rect 595 524 608 554
rect 623 536 653 554
rect 696 540 710 554
rect 746 540 966 554
rect 697 538 710 540
rect 663 526 678 538
rect 660 524 682 526
rect 687 524 717 538
rect 778 536 931 540
rect 760 524 952 536
rect 995 524 1025 538
rect 1031 524 1044 554
rect 1059 536 1089 554
rect 1132 524 1145 554
rect 1175 524 1188 554
rect 1203 536 1233 554
rect 1276 540 1290 554
rect 1326 540 1546 554
rect 1277 538 1290 540
rect 1243 526 1258 538
rect 1240 524 1262 526
rect 1267 524 1297 538
rect 1358 536 1511 540
rect 1340 524 1532 536
rect 1575 524 1605 538
rect 1611 524 1624 554
rect 1639 536 1669 554
rect 1712 524 1725 554
rect 1755 524 1768 554
rect 1783 536 1813 554
rect 1856 540 1870 554
rect 1906 540 2126 554
rect 1857 538 1870 540
rect 1823 526 1838 538
rect 1820 524 1842 526
rect 1847 524 1877 538
rect 1938 536 2091 540
rect 1920 524 2112 536
rect 2155 524 2185 538
rect 2191 524 2204 554
rect 2219 536 2249 554
rect 2292 524 2305 554
rect 2335 524 2348 554
rect 2363 536 2393 554
rect 2436 540 2450 554
rect 2486 540 2706 554
rect 2437 538 2450 540
rect 2403 526 2418 538
rect 2400 524 2422 526
rect 2427 524 2457 538
rect 2518 536 2671 540
rect 2500 524 2692 536
rect 2735 524 2765 538
rect 2771 524 2784 554
rect 2799 536 2829 554
rect 2872 524 2885 554
rect 2915 524 2928 554
rect 2943 536 2973 554
rect 3016 540 3030 554
rect 3066 540 3286 554
rect 3017 538 3030 540
rect 2983 526 2998 538
rect 2980 524 3002 526
rect 3007 524 3037 538
rect 3098 536 3251 540
rect 3080 524 3272 536
rect 3315 524 3345 538
rect 3351 524 3364 554
rect 3379 536 3409 554
rect 3452 524 3465 554
rect 3495 524 3508 554
rect 3523 536 3553 554
rect 3596 540 3610 554
rect 3646 540 3866 554
rect 3597 538 3610 540
rect 3563 526 3578 538
rect 3560 524 3582 526
rect 3587 524 3617 538
rect 3678 536 3831 540
rect 3660 524 3852 536
rect 3895 524 3925 538
rect 3931 524 3944 554
rect 3959 536 3989 554
rect 4032 524 4045 554
rect 4075 524 4088 554
rect 4103 536 4133 554
rect 4176 540 4190 554
rect 4226 540 4446 554
rect 4177 538 4190 540
rect 4143 526 4158 538
rect 4140 524 4162 526
rect 4167 524 4197 538
rect 4258 536 4411 540
rect 4240 524 4432 536
rect 4475 524 4505 538
rect 4511 524 4524 554
rect 4539 536 4569 554
rect 4612 524 4625 554
rect 0 510 4625 524
rect 15 406 28 510
rect 73 488 74 498
rect 89 488 102 498
rect 73 484 102 488
rect 107 484 137 510
rect 155 496 171 498
rect 243 496 296 510
rect 244 494 308 496
rect 351 494 366 510
rect 415 507 445 510
rect 415 504 451 507
rect 381 496 397 498
rect 155 484 170 488
rect 73 482 170 484
rect 198 482 366 494
rect 382 484 397 488
rect 415 485 454 504
rect 473 498 480 499
rect 479 491 480 498
rect 463 488 464 491
rect 479 488 492 491
rect 415 484 445 485
rect 454 484 460 485
rect 463 484 492 488
rect 382 483 492 484
rect 382 482 498 483
rect 57 474 108 482
rect 57 462 82 474
rect 89 462 108 474
rect 139 474 189 482
rect 139 466 155 474
rect 162 472 189 474
rect 198 472 419 482
rect 162 462 419 472
rect 448 474 498 482
rect 448 465 464 474
rect 57 454 108 462
rect 155 454 419 462
rect 445 462 464 465
rect 471 462 498 474
rect 445 454 498 462
rect 73 446 74 454
rect 89 446 102 454
rect 73 438 89 446
rect 70 431 89 434
rect 70 422 92 431
rect 43 412 92 422
rect 43 406 73 412
rect 92 407 97 412
rect 15 390 89 406
rect 107 398 137 454
rect 172 444 380 454
rect 415 450 460 454
rect 463 453 464 454
rect 479 453 492 454
rect 198 414 387 444
rect 213 411 387 414
rect 206 408 387 411
rect 15 388 28 390
rect 43 388 77 390
rect 15 372 89 388
rect 116 384 129 398
rect 144 384 160 400
rect 206 395 217 408
rect -1 350 0 366
rect 15 350 28 372
rect 43 350 73 372
rect 116 368 178 384
rect 206 377 217 393
rect 222 388 232 408
rect 242 388 256 408
rect 259 395 268 408
rect 284 395 293 408
rect 222 377 256 388
rect 259 377 268 393
rect 284 377 293 393
rect 300 388 310 408
rect 320 388 334 408
rect 335 395 346 408
rect 300 377 334 388
rect 335 377 346 393
rect 392 384 408 400
rect 415 398 445 450
rect 479 446 480 453
rect 464 438 480 446
rect 451 406 464 425
rect 479 406 509 422
rect 451 390 525 406
rect 451 388 464 390
rect 479 388 513 390
rect 116 366 129 368
rect 144 366 178 368
rect 116 350 178 366
rect 222 361 238 364
rect 300 361 330 372
rect 378 368 424 384
rect 451 372 525 388
rect 378 366 412 368
rect 377 350 424 366
rect 451 350 464 372
rect 479 350 509 372
rect 536 350 537 366
rect 552 350 565 510
rect 595 406 608 510
rect 653 488 654 498
rect 669 488 682 498
rect 653 484 682 488
rect 687 484 717 510
rect 735 496 751 498
rect 823 496 876 510
rect 824 494 888 496
rect 931 494 946 510
rect 995 507 1025 510
rect 995 504 1031 507
rect 961 496 977 498
rect 735 484 750 488
rect 653 482 750 484
rect 778 482 946 494
rect 962 484 977 488
rect 995 485 1034 504
rect 1053 498 1060 499
rect 1059 491 1060 498
rect 1043 488 1044 491
rect 1059 488 1072 491
rect 995 484 1025 485
rect 1034 484 1040 485
rect 1043 484 1072 488
rect 962 483 1072 484
rect 962 482 1078 483
rect 637 474 688 482
rect 637 462 662 474
rect 669 462 688 474
rect 719 474 769 482
rect 719 466 735 474
rect 742 472 769 474
rect 778 472 999 482
rect 742 462 999 472
rect 1028 474 1078 482
rect 1028 465 1044 474
rect 637 454 688 462
rect 735 454 999 462
rect 1025 462 1044 465
rect 1051 462 1078 474
rect 1025 454 1078 462
rect 653 446 654 454
rect 669 446 682 454
rect 653 438 669 446
rect 650 431 669 434
rect 650 422 672 431
rect 623 412 672 422
rect 623 406 653 412
rect 672 407 677 412
rect 595 390 669 406
rect 687 398 717 454
rect 752 444 960 454
rect 995 450 1040 454
rect 1043 453 1044 454
rect 1059 453 1072 454
rect 778 414 967 444
rect 793 411 967 414
rect 786 408 967 411
rect 595 388 608 390
rect 623 388 657 390
rect 595 372 669 388
rect 696 384 709 398
rect 724 384 740 400
rect 786 395 797 408
rect 579 350 580 366
rect 595 350 608 372
rect 623 350 653 372
rect 696 368 758 384
rect 786 377 797 393
rect 802 388 812 408
rect 822 388 836 408
rect 839 395 848 408
rect 864 395 873 408
rect 802 377 836 388
rect 839 377 848 393
rect 864 377 873 393
rect 880 388 890 408
rect 900 388 914 408
rect 915 395 926 408
rect 880 377 914 388
rect 915 377 926 393
rect 972 384 988 400
rect 995 398 1025 450
rect 1059 446 1060 453
rect 1044 438 1060 446
rect 1031 406 1044 425
rect 1059 406 1089 422
rect 1031 390 1105 406
rect 1031 388 1044 390
rect 1059 388 1093 390
rect 696 366 709 368
rect 724 366 758 368
rect 696 350 758 366
rect 802 361 818 364
rect 880 361 910 372
rect 958 368 1004 384
rect 1031 372 1105 388
rect 958 366 992 368
rect 957 350 1004 366
rect 1031 350 1044 372
rect 1059 350 1089 372
rect 1116 350 1117 366
rect 1132 350 1145 510
rect 1175 406 1188 510
rect 1233 488 1234 498
rect 1249 488 1262 498
rect 1233 484 1262 488
rect 1267 484 1297 510
rect 1315 496 1331 498
rect 1403 496 1456 510
rect 1404 494 1468 496
rect 1511 494 1526 510
rect 1575 507 1605 510
rect 1575 504 1611 507
rect 1541 496 1557 498
rect 1315 484 1330 488
rect 1233 482 1330 484
rect 1358 482 1526 494
rect 1542 484 1557 488
rect 1575 485 1614 504
rect 1633 498 1640 499
rect 1639 491 1640 498
rect 1623 488 1624 491
rect 1639 488 1652 491
rect 1575 484 1605 485
rect 1614 484 1620 485
rect 1623 484 1652 488
rect 1542 483 1652 484
rect 1542 482 1658 483
rect 1217 474 1268 482
rect 1217 462 1242 474
rect 1249 462 1268 474
rect 1299 474 1349 482
rect 1299 466 1315 474
rect 1322 472 1349 474
rect 1358 472 1579 482
rect 1322 462 1579 472
rect 1608 474 1658 482
rect 1608 465 1624 474
rect 1217 454 1268 462
rect 1315 454 1579 462
rect 1605 462 1624 465
rect 1631 462 1658 474
rect 1605 454 1658 462
rect 1233 446 1234 454
rect 1249 446 1262 454
rect 1233 438 1249 446
rect 1230 431 1249 434
rect 1230 422 1252 431
rect 1203 412 1252 422
rect 1203 406 1233 412
rect 1252 407 1257 412
rect 1175 390 1249 406
rect 1267 398 1297 454
rect 1332 444 1540 454
rect 1575 450 1620 454
rect 1623 453 1624 454
rect 1639 453 1652 454
rect 1358 414 1547 444
rect 1373 411 1547 414
rect 1366 408 1547 411
rect 1175 388 1188 390
rect 1203 388 1237 390
rect 1175 372 1249 388
rect 1276 384 1289 398
rect 1304 384 1320 400
rect 1366 395 1377 408
rect 1159 350 1160 366
rect 1175 350 1188 372
rect 1203 350 1233 372
rect 1276 368 1338 384
rect 1366 377 1377 393
rect 1382 388 1392 408
rect 1402 388 1416 408
rect 1419 395 1428 408
rect 1444 395 1453 408
rect 1382 377 1416 388
rect 1419 377 1428 393
rect 1444 377 1453 393
rect 1460 388 1470 408
rect 1480 388 1494 408
rect 1495 395 1506 408
rect 1460 377 1494 388
rect 1495 377 1506 393
rect 1552 384 1568 400
rect 1575 398 1605 450
rect 1639 446 1640 453
rect 1624 438 1640 446
rect 1611 406 1624 425
rect 1639 406 1669 422
rect 1611 390 1685 406
rect 1611 388 1624 390
rect 1639 388 1673 390
rect 1276 366 1289 368
rect 1304 366 1338 368
rect 1276 350 1338 366
rect 1382 361 1398 364
rect 1460 361 1490 372
rect 1538 368 1584 384
rect 1611 372 1685 388
rect 1538 366 1572 368
rect 1537 350 1584 366
rect 1611 350 1624 372
rect 1639 350 1669 372
rect 1696 350 1697 366
rect 1712 350 1725 510
rect 1755 406 1768 510
rect 1813 488 1814 498
rect 1829 488 1842 498
rect 1813 484 1842 488
rect 1847 484 1877 510
rect 1895 496 1911 498
rect 1983 496 2036 510
rect 1984 494 2048 496
rect 2091 494 2106 510
rect 2155 507 2185 510
rect 2155 504 2191 507
rect 2121 496 2137 498
rect 1895 484 1910 488
rect 1813 482 1910 484
rect 1938 482 2106 494
rect 2122 484 2137 488
rect 2155 485 2194 504
rect 2213 498 2220 499
rect 2219 491 2220 498
rect 2203 488 2204 491
rect 2219 488 2232 491
rect 2155 484 2185 485
rect 2194 484 2200 485
rect 2203 484 2232 488
rect 2122 483 2232 484
rect 2122 482 2238 483
rect 1797 474 1848 482
rect 1797 462 1822 474
rect 1829 462 1848 474
rect 1879 474 1929 482
rect 1879 466 1895 474
rect 1902 472 1929 474
rect 1938 472 2159 482
rect 1902 462 2159 472
rect 2188 474 2238 482
rect 2188 465 2204 474
rect 1797 454 1848 462
rect 1895 454 2159 462
rect 2185 462 2204 465
rect 2211 462 2238 474
rect 2185 454 2238 462
rect 1813 446 1814 454
rect 1829 446 1842 454
rect 1813 438 1829 446
rect 1810 431 1829 434
rect 1810 422 1832 431
rect 1783 412 1832 422
rect 1783 406 1813 412
rect 1832 407 1837 412
rect 1755 390 1829 406
rect 1847 398 1877 454
rect 1912 444 2120 454
rect 2155 450 2200 454
rect 2203 453 2204 454
rect 2219 453 2232 454
rect 1938 414 2127 444
rect 1953 411 2127 414
rect 1946 408 2127 411
rect 1755 388 1768 390
rect 1783 388 1817 390
rect 1755 372 1829 388
rect 1856 384 1869 398
rect 1884 384 1900 400
rect 1946 395 1957 408
rect 1739 350 1740 366
rect 1755 350 1768 372
rect 1783 350 1813 372
rect 1856 368 1918 384
rect 1946 377 1957 393
rect 1962 388 1972 408
rect 1982 388 1996 408
rect 1999 395 2008 408
rect 2024 395 2033 408
rect 1962 377 1996 388
rect 1999 377 2008 393
rect 2024 377 2033 393
rect 2040 388 2050 408
rect 2060 388 2074 408
rect 2075 395 2086 408
rect 2040 377 2074 388
rect 2075 377 2086 393
rect 2132 384 2148 400
rect 2155 398 2185 450
rect 2219 446 2220 453
rect 2204 438 2220 446
rect 2191 406 2204 425
rect 2219 406 2249 422
rect 2191 390 2265 406
rect 2191 388 2204 390
rect 2219 388 2253 390
rect 1856 366 1869 368
rect 1884 366 1918 368
rect 1856 350 1918 366
rect 1962 361 1978 364
rect 2040 361 2070 372
rect 2118 368 2164 384
rect 2191 372 2265 388
rect 2118 366 2152 368
rect 2117 350 2164 366
rect 2191 350 2204 372
rect 2219 350 2249 372
rect 2276 350 2277 366
rect 2292 350 2305 510
rect 2335 406 2348 510
rect 2393 488 2394 498
rect 2409 488 2422 498
rect 2393 484 2422 488
rect 2427 484 2457 510
rect 2475 496 2491 498
rect 2563 496 2616 510
rect 2564 494 2628 496
rect 2671 494 2686 510
rect 2735 507 2765 510
rect 2735 504 2771 507
rect 2701 496 2717 498
rect 2475 484 2490 488
rect 2393 482 2490 484
rect 2518 482 2686 494
rect 2702 484 2717 488
rect 2735 485 2774 504
rect 2793 498 2800 499
rect 2799 491 2800 498
rect 2783 488 2784 491
rect 2799 488 2812 491
rect 2735 484 2765 485
rect 2774 484 2780 485
rect 2783 484 2812 488
rect 2702 483 2812 484
rect 2702 482 2818 483
rect 2377 474 2428 482
rect 2377 462 2402 474
rect 2409 462 2428 474
rect 2459 474 2509 482
rect 2459 466 2475 474
rect 2482 472 2509 474
rect 2518 472 2739 482
rect 2482 462 2739 472
rect 2768 474 2818 482
rect 2768 465 2784 474
rect 2377 454 2428 462
rect 2475 454 2739 462
rect 2765 462 2784 465
rect 2791 462 2818 474
rect 2765 454 2818 462
rect 2393 446 2394 454
rect 2409 446 2422 454
rect 2393 438 2409 446
rect 2390 431 2409 434
rect 2390 422 2412 431
rect 2363 412 2412 422
rect 2363 406 2393 412
rect 2412 407 2417 412
rect 2335 390 2409 406
rect 2427 398 2457 454
rect 2492 444 2700 454
rect 2735 450 2780 454
rect 2783 453 2784 454
rect 2799 453 2812 454
rect 2518 414 2707 444
rect 2533 411 2707 414
rect 2526 408 2707 411
rect 2335 388 2348 390
rect 2363 388 2397 390
rect 2335 372 2409 388
rect 2436 384 2449 398
rect 2464 384 2480 400
rect 2526 395 2537 408
rect 2319 350 2320 366
rect 2335 350 2348 372
rect 2363 350 2393 372
rect 2436 368 2498 384
rect 2526 377 2537 393
rect 2542 388 2552 408
rect 2562 388 2576 408
rect 2579 395 2588 408
rect 2604 395 2613 408
rect 2542 377 2576 388
rect 2579 377 2588 393
rect 2604 377 2613 393
rect 2620 388 2630 408
rect 2640 388 2654 408
rect 2655 395 2666 408
rect 2620 377 2654 388
rect 2655 377 2666 393
rect 2712 384 2728 400
rect 2735 398 2765 450
rect 2799 446 2800 453
rect 2784 438 2800 446
rect 2771 406 2784 425
rect 2799 406 2829 422
rect 2771 390 2845 406
rect 2771 388 2784 390
rect 2799 388 2833 390
rect 2436 366 2449 368
rect 2464 366 2498 368
rect 2436 350 2498 366
rect 2542 361 2558 364
rect 2620 361 2650 372
rect 2698 368 2744 384
rect 2771 372 2845 388
rect 2698 366 2732 368
rect 2697 350 2744 366
rect 2771 350 2784 372
rect 2799 350 2829 372
rect 2856 350 2857 366
rect 2872 350 2885 510
rect 2915 406 2928 510
rect 2973 488 2974 498
rect 2989 488 3002 498
rect 2973 484 3002 488
rect 3007 484 3037 510
rect 3055 496 3071 498
rect 3143 496 3196 510
rect 3144 494 3208 496
rect 3251 494 3266 510
rect 3315 507 3345 510
rect 3315 504 3351 507
rect 3281 496 3297 498
rect 3055 484 3070 488
rect 2973 482 3070 484
rect 3098 482 3266 494
rect 3282 484 3297 488
rect 3315 485 3354 504
rect 3373 498 3380 499
rect 3379 491 3380 498
rect 3363 488 3364 491
rect 3379 488 3392 491
rect 3315 484 3345 485
rect 3354 484 3360 485
rect 3363 484 3392 488
rect 3282 483 3392 484
rect 3282 482 3398 483
rect 2957 474 3008 482
rect 2957 462 2982 474
rect 2989 462 3008 474
rect 3039 474 3089 482
rect 3039 466 3055 474
rect 3062 472 3089 474
rect 3098 472 3319 482
rect 3062 462 3319 472
rect 3348 474 3398 482
rect 3348 465 3364 474
rect 2957 454 3008 462
rect 3055 454 3319 462
rect 3345 462 3364 465
rect 3371 462 3398 474
rect 3345 454 3398 462
rect 2973 446 2974 454
rect 2989 446 3002 454
rect 2973 438 2989 446
rect 2970 431 2989 434
rect 2970 422 2992 431
rect 2943 412 2992 422
rect 2943 406 2973 412
rect 2992 407 2997 412
rect 2915 390 2989 406
rect 3007 398 3037 454
rect 3072 444 3280 454
rect 3315 450 3360 454
rect 3363 453 3364 454
rect 3379 453 3392 454
rect 3098 414 3287 444
rect 3113 411 3287 414
rect 3106 408 3287 411
rect 2915 388 2928 390
rect 2943 388 2977 390
rect 2915 372 2989 388
rect 3016 384 3029 398
rect 3044 384 3060 400
rect 3106 395 3117 408
rect 2899 350 2900 366
rect 2915 350 2928 372
rect 2943 350 2973 372
rect 3016 368 3078 384
rect 3106 377 3117 393
rect 3122 388 3132 408
rect 3142 388 3156 408
rect 3159 395 3168 408
rect 3184 395 3193 408
rect 3122 377 3156 388
rect 3159 377 3168 393
rect 3184 377 3193 393
rect 3200 388 3210 408
rect 3220 388 3234 408
rect 3235 395 3246 408
rect 3200 377 3234 388
rect 3235 377 3246 393
rect 3292 384 3308 400
rect 3315 398 3345 450
rect 3379 446 3380 453
rect 3364 438 3380 446
rect 3351 406 3364 425
rect 3379 406 3409 422
rect 3351 390 3425 406
rect 3351 388 3364 390
rect 3379 388 3413 390
rect 3016 366 3029 368
rect 3044 366 3078 368
rect 3016 350 3078 366
rect 3122 361 3138 364
rect 3200 361 3230 372
rect 3278 368 3324 384
rect 3351 372 3425 388
rect 3278 366 3312 368
rect 3277 350 3324 366
rect 3351 350 3364 372
rect 3379 350 3409 372
rect 3436 350 3437 366
rect 3452 350 3465 510
rect 3495 406 3508 510
rect 3553 488 3554 498
rect 3569 488 3582 498
rect 3553 484 3582 488
rect 3587 484 3617 510
rect 3635 496 3651 498
rect 3723 496 3776 510
rect 3724 494 3788 496
rect 3831 494 3846 510
rect 3895 507 3925 510
rect 3895 504 3931 507
rect 3861 496 3877 498
rect 3635 484 3650 488
rect 3553 482 3650 484
rect 3678 482 3846 494
rect 3862 484 3877 488
rect 3895 485 3934 504
rect 3953 498 3960 499
rect 3959 491 3960 498
rect 3943 488 3944 491
rect 3959 488 3972 491
rect 3895 484 3925 485
rect 3934 484 3940 485
rect 3943 484 3972 488
rect 3862 483 3972 484
rect 3862 482 3978 483
rect 3537 474 3588 482
rect 3537 462 3562 474
rect 3569 462 3588 474
rect 3619 474 3669 482
rect 3619 466 3635 474
rect 3642 472 3669 474
rect 3678 472 3899 482
rect 3642 462 3899 472
rect 3928 474 3978 482
rect 3928 465 3944 474
rect 3537 454 3588 462
rect 3635 454 3899 462
rect 3925 462 3944 465
rect 3951 462 3978 474
rect 3925 454 3978 462
rect 3553 446 3554 454
rect 3569 446 3582 454
rect 3553 438 3569 446
rect 3550 431 3569 434
rect 3550 422 3572 431
rect 3523 412 3572 422
rect 3523 406 3553 412
rect 3572 407 3577 412
rect 3495 390 3569 406
rect 3587 398 3617 454
rect 3652 444 3860 454
rect 3895 450 3940 454
rect 3943 453 3944 454
rect 3959 453 3972 454
rect 3678 414 3867 444
rect 3693 411 3867 414
rect 3686 408 3867 411
rect 3495 388 3508 390
rect 3523 388 3557 390
rect 3495 372 3569 388
rect 3596 384 3609 398
rect 3624 384 3640 400
rect 3686 395 3697 408
rect 3479 350 3480 366
rect 3495 350 3508 372
rect 3523 350 3553 372
rect 3596 368 3658 384
rect 3686 377 3697 393
rect 3702 388 3712 408
rect 3722 388 3736 408
rect 3739 395 3748 408
rect 3764 395 3773 408
rect 3702 377 3736 388
rect 3739 377 3748 393
rect 3764 377 3773 393
rect 3780 388 3790 408
rect 3800 388 3814 408
rect 3815 395 3826 408
rect 3780 377 3814 388
rect 3815 377 3826 393
rect 3872 384 3888 400
rect 3895 398 3925 450
rect 3959 446 3960 453
rect 3944 438 3960 446
rect 3931 406 3944 425
rect 3959 406 3989 422
rect 3931 390 4005 406
rect 3931 388 3944 390
rect 3959 388 3993 390
rect 3596 366 3609 368
rect 3624 366 3658 368
rect 3596 350 3658 366
rect 3702 361 3718 364
rect 3780 361 3810 372
rect 3858 368 3904 384
rect 3931 372 4005 388
rect 3858 366 3892 368
rect 3857 350 3904 366
rect 3931 350 3944 372
rect 3959 350 3989 372
rect 4016 350 4017 366
rect 4032 350 4045 510
rect 4075 406 4088 510
rect 4133 488 4134 498
rect 4149 488 4162 498
rect 4133 484 4162 488
rect 4167 484 4197 510
rect 4215 496 4231 498
rect 4303 496 4356 510
rect 4304 494 4368 496
rect 4411 494 4426 510
rect 4475 507 4505 510
rect 4475 504 4511 507
rect 4441 496 4457 498
rect 4215 484 4230 488
rect 4133 482 4230 484
rect 4258 482 4426 494
rect 4442 484 4457 488
rect 4475 485 4514 504
rect 4533 498 4540 499
rect 4539 491 4540 498
rect 4523 488 4524 491
rect 4539 488 4552 491
rect 4475 484 4505 485
rect 4514 484 4520 485
rect 4523 484 4552 488
rect 4442 483 4552 484
rect 4442 482 4558 483
rect 4117 474 4168 482
rect 4117 462 4142 474
rect 4149 462 4168 474
rect 4199 474 4249 482
rect 4199 466 4215 474
rect 4222 472 4249 474
rect 4258 472 4479 482
rect 4222 462 4479 472
rect 4508 474 4558 482
rect 4508 465 4524 474
rect 4117 454 4168 462
rect 4215 454 4479 462
rect 4505 462 4524 465
rect 4531 462 4558 474
rect 4505 454 4558 462
rect 4133 446 4134 454
rect 4149 446 4162 454
rect 4133 438 4149 446
rect 4130 431 4149 434
rect 4130 422 4152 431
rect 4103 412 4152 422
rect 4103 406 4133 412
rect 4152 407 4157 412
rect 4075 390 4149 406
rect 4167 398 4197 454
rect 4232 444 4440 454
rect 4475 450 4520 454
rect 4523 453 4524 454
rect 4539 453 4552 454
rect 4258 414 4447 444
rect 4273 411 4447 414
rect 4266 408 4447 411
rect 4075 388 4088 390
rect 4103 388 4137 390
rect 4075 372 4149 388
rect 4176 384 4189 398
rect 4204 384 4220 400
rect 4266 395 4277 408
rect 4059 350 4060 366
rect 4075 350 4088 372
rect 4103 350 4133 372
rect 4176 368 4238 384
rect 4266 377 4277 393
rect 4282 388 4292 408
rect 4302 388 4316 408
rect 4319 395 4328 408
rect 4344 395 4353 408
rect 4282 377 4316 388
rect 4319 377 4328 393
rect 4344 377 4353 393
rect 4360 388 4370 408
rect 4380 388 4394 408
rect 4395 395 4406 408
rect 4360 377 4394 388
rect 4395 377 4406 393
rect 4452 384 4468 400
rect 4475 398 4505 450
rect 4539 446 4540 453
rect 4524 438 4540 446
rect 4511 406 4524 425
rect 4539 406 4569 422
rect 4511 390 4585 406
rect 4511 388 4524 390
rect 4539 388 4573 390
rect 4176 366 4189 368
rect 4204 366 4238 368
rect 4176 350 4238 366
rect 4282 361 4298 364
rect 4360 361 4390 372
rect 4438 368 4484 384
rect 4511 372 4585 388
rect 4438 366 4472 368
rect 4437 350 4484 366
rect 4511 350 4524 372
rect 4539 350 4569 372
rect 4596 350 4597 366
rect 4612 350 4625 510
rect -7 342 34 350
rect -7 316 8 342
rect 15 316 34 342
rect 98 338 160 350
rect 172 338 247 350
rect 305 338 380 350
rect 392 338 423 350
rect 429 338 464 350
rect 98 336 260 338
rect -7 308 34 316
rect 116 312 129 336
rect 144 334 159 336
rect -1 298 0 308
rect 15 298 28 308
rect 43 298 73 312
rect 116 298 159 312
rect 183 309 190 316
rect 193 312 260 336
rect 292 336 464 338
rect 262 314 290 318
rect 292 314 372 336
rect 393 334 408 336
rect 262 312 372 314
rect 193 308 372 312
rect 166 298 196 308
rect 198 298 351 308
rect 359 298 389 308
rect 393 298 423 312
rect 451 298 464 336
rect 536 342 571 350
rect 536 316 537 342
rect 544 316 571 342
rect 479 298 509 312
rect 536 308 571 316
rect 573 342 614 350
rect 573 316 588 342
rect 595 316 614 342
rect 678 338 740 350
rect 752 338 827 350
rect 885 338 960 350
rect 972 338 1003 350
rect 1009 338 1044 350
rect 678 336 840 338
rect 573 308 614 316
rect 696 312 709 336
rect 724 334 739 336
rect 536 298 537 308
rect 552 298 565 308
rect 579 298 580 308
rect 595 298 608 308
rect 623 298 653 312
rect 696 298 739 312
rect 763 309 770 316
rect 773 312 840 336
rect 872 336 1044 338
rect 842 314 870 318
rect 872 314 952 336
rect 973 334 988 336
rect 842 312 952 314
rect 773 308 952 312
rect 746 298 776 308
rect 778 298 931 308
rect 939 298 969 308
rect 973 298 1003 312
rect 1031 298 1044 336
rect 1116 342 1151 350
rect 1116 316 1117 342
rect 1124 316 1151 342
rect 1059 298 1089 312
rect 1116 308 1151 316
rect 1153 342 1194 350
rect 1153 316 1168 342
rect 1175 316 1194 342
rect 1258 338 1320 350
rect 1332 338 1407 350
rect 1465 338 1540 350
rect 1552 338 1583 350
rect 1589 338 1624 350
rect 1258 336 1420 338
rect 1153 308 1194 316
rect 1276 312 1289 336
rect 1304 334 1319 336
rect 1116 298 1117 308
rect 1132 298 1145 308
rect 1159 298 1160 308
rect 1175 298 1188 308
rect 1203 298 1233 312
rect 1276 298 1319 312
rect 1343 309 1350 316
rect 1353 312 1420 336
rect 1452 336 1624 338
rect 1422 314 1450 318
rect 1452 314 1532 336
rect 1553 334 1568 336
rect 1422 312 1532 314
rect 1353 308 1532 312
rect 1326 298 1356 308
rect 1358 298 1511 308
rect 1519 298 1549 308
rect 1553 298 1583 312
rect 1611 298 1624 336
rect 1696 342 1731 350
rect 1696 316 1697 342
rect 1704 316 1731 342
rect 1639 298 1669 312
rect 1696 308 1731 316
rect 1733 342 1774 350
rect 1733 316 1748 342
rect 1755 316 1774 342
rect 1838 338 1900 350
rect 1912 338 1987 350
rect 2045 338 2120 350
rect 2132 338 2163 350
rect 2169 338 2204 350
rect 1838 336 2000 338
rect 1733 308 1774 316
rect 1856 312 1869 336
rect 1884 334 1899 336
rect 1696 298 1697 308
rect 1712 298 1725 308
rect 1739 298 1740 308
rect 1755 298 1768 308
rect 1783 298 1813 312
rect 1856 298 1899 312
rect 1923 309 1930 316
rect 1933 312 2000 336
rect 2032 336 2204 338
rect 2002 314 2030 318
rect 2032 314 2112 336
rect 2133 334 2148 336
rect 2002 312 2112 314
rect 1933 308 2112 312
rect 1906 298 1936 308
rect 1938 298 2091 308
rect 2099 298 2129 308
rect 2133 298 2163 312
rect 2191 298 2204 336
rect 2276 342 2311 350
rect 2276 316 2277 342
rect 2284 316 2311 342
rect 2219 298 2249 312
rect 2276 308 2311 316
rect 2313 342 2354 350
rect 2313 316 2328 342
rect 2335 316 2354 342
rect 2418 338 2480 350
rect 2492 338 2567 350
rect 2625 338 2700 350
rect 2712 338 2743 350
rect 2749 338 2784 350
rect 2418 336 2580 338
rect 2313 308 2354 316
rect 2436 312 2449 336
rect 2464 334 2479 336
rect 2276 298 2277 308
rect 2292 298 2305 308
rect 2319 298 2320 308
rect 2335 298 2348 308
rect 2363 298 2393 312
rect 2436 298 2479 312
rect 2503 309 2510 316
rect 2513 312 2580 336
rect 2612 336 2784 338
rect 2582 314 2610 318
rect 2612 314 2692 336
rect 2713 334 2728 336
rect 2582 312 2692 314
rect 2513 308 2692 312
rect 2486 298 2516 308
rect 2518 298 2671 308
rect 2679 298 2709 308
rect 2713 298 2743 312
rect 2771 298 2784 336
rect 2856 342 2891 350
rect 2856 316 2857 342
rect 2864 316 2891 342
rect 2799 298 2829 312
rect 2856 308 2891 316
rect 2893 342 2934 350
rect 2893 316 2908 342
rect 2915 316 2934 342
rect 2998 338 3060 350
rect 3072 338 3147 350
rect 3205 338 3280 350
rect 3292 338 3323 350
rect 3329 338 3364 350
rect 2998 336 3160 338
rect 2893 308 2934 316
rect 3016 312 3029 336
rect 3044 334 3059 336
rect 2856 298 2857 308
rect 2872 298 2885 308
rect 2899 298 2900 308
rect 2915 298 2928 308
rect 2943 298 2973 312
rect 3016 298 3059 312
rect 3083 309 3090 316
rect 3093 312 3160 336
rect 3192 336 3364 338
rect 3162 314 3190 318
rect 3192 314 3272 336
rect 3293 334 3308 336
rect 3162 312 3272 314
rect 3093 308 3272 312
rect 3066 298 3096 308
rect 3098 298 3251 308
rect 3259 298 3289 308
rect 3293 298 3323 312
rect 3351 298 3364 336
rect 3436 342 3471 350
rect 3436 316 3437 342
rect 3444 316 3471 342
rect 3379 298 3409 312
rect 3436 308 3471 316
rect 3473 342 3514 350
rect 3473 316 3488 342
rect 3495 316 3514 342
rect 3578 338 3640 350
rect 3652 338 3727 350
rect 3785 338 3860 350
rect 3872 338 3903 350
rect 3909 338 3944 350
rect 3578 336 3740 338
rect 3473 308 3514 316
rect 3596 312 3609 336
rect 3624 334 3639 336
rect 3436 298 3437 308
rect 3452 298 3465 308
rect 3479 298 3480 308
rect 3495 298 3508 308
rect 3523 298 3553 312
rect 3596 298 3639 312
rect 3663 309 3670 316
rect 3673 312 3740 336
rect 3772 336 3944 338
rect 3742 314 3770 318
rect 3772 314 3852 336
rect 3873 334 3888 336
rect 3742 312 3852 314
rect 3673 308 3852 312
rect 3646 298 3676 308
rect 3678 298 3831 308
rect 3839 298 3869 308
rect 3873 298 3903 312
rect 3931 298 3944 336
rect 4016 342 4051 350
rect 4016 316 4017 342
rect 4024 316 4051 342
rect 3959 298 3989 312
rect 4016 308 4051 316
rect 4053 342 4094 350
rect 4053 316 4068 342
rect 4075 316 4094 342
rect 4158 338 4220 350
rect 4232 338 4307 350
rect 4365 338 4440 350
rect 4452 338 4483 350
rect 4489 338 4524 350
rect 4158 336 4320 338
rect 4053 308 4094 316
rect 4176 312 4189 336
rect 4204 334 4219 336
rect 4016 298 4017 308
rect 4032 298 4045 308
rect 4059 298 4060 308
rect 4075 298 4088 308
rect 4103 298 4133 312
rect 4176 298 4219 312
rect 4243 309 4250 316
rect 4253 312 4320 336
rect 4352 336 4524 338
rect 4322 314 4350 318
rect 4352 314 4432 336
rect 4453 334 4468 336
rect 4322 312 4432 314
rect 4253 308 4432 312
rect 4226 298 4256 308
rect 4258 298 4411 308
rect 4419 298 4449 308
rect 4453 298 4483 312
rect 4511 298 4524 336
rect 4596 342 4631 350
rect 4596 316 4597 342
rect 4604 316 4631 342
rect 4539 298 4569 312
rect 4596 308 4631 316
rect 4596 298 4597 308
rect 4612 298 4625 308
rect -1 292 4625 298
rect 0 284 4625 292
rect 15 254 28 284
rect 43 266 73 284
rect 116 270 130 284
rect 166 270 386 284
rect 117 268 130 270
rect 83 256 98 268
rect 80 254 102 256
rect 107 254 137 268
rect 198 266 351 270
rect 180 254 372 266
rect 415 254 445 268
rect 451 254 464 284
rect 479 266 509 284
rect 552 254 565 284
rect 595 254 608 284
rect 623 266 653 284
rect 696 270 710 284
rect 746 270 966 284
rect 697 268 710 270
rect 663 256 678 268
rect 660 254 682 256
rect 687 254 717 268
rect 778 266 931 270
rect 760 254 952 266
rect 995 254 1025 268
rect 1031 254 1044 284
rect 1059 266 1089 284
rect 1132 254 1145 284
rect 1175 254 1188 284
rect 1203 266 1233 284
rect 1276 270 1290 284
rect 1326 270 1546 284
rect 1277 268 1290 270
rect 1243 256 1258 268
rect 1240 254 1262 256
rect 1267 254 1297 268
rect 1358 266 1511 270
rect 1340 254 1532 266
rect 1575 254 1605 268
rect 1611 254 1624 284
rect 1639 266 1669 284
rect 1712 254 1725 284
rect 1755 254 1768 284
rect 1783 266 1813 284
rect 1856 270 1870 284
rect 1906 270 2126 284
rect 1857 268 1870 270
rect 1823 256 1838 268
rect 1820 254 1842 256
rect 1847 254 1877 268
rect 1938 266 2091 270
rect 1920 254 2112 266
rect 2155 254 2185 268
rect 2191 254 2204 284
rect 2219 266 2249 284
rect 2292 254 2305 284
rect 2335 254 2348 284
rect 2363 266 2393 284
rect 2436 270 2450 284
rect 2486 270 2706 284
rect 2437 268 2450 270
rect 2403 256 2418 268
rect 2400 254 2422 256
rect 2427 254 2457 268
rect 2518 266 2671 270
rect 2500 254 2692 266
rect 2735 254 2765 268
rect 2771 254 2784 284
rect 2799 266 2829 284
rect 2872 254 2885 284
rect 2915 254 2928 284
rect 2943 266 2973 284
rect 3016 270 3030 284
rect 3066 270 3286 284
rect 3017 268 3030 270
rect 2983 256 2998 268
rect 2980 254 3002 256
rect 3007 254 3037 268
rect 3098 266 3251 270
rect 3080 254 3272 266
rect 3315 254 3345 268
rect 3351 254 3364 284
rect 3379 266 3409 284
rect 3452 254 3465 284
rect 3495 254 3508 284
rect 3523 266 3553 284
rect 3596 270 3610 284
rect 3646 270 3866 284
rect 3597 268 3610 270
rect 3563 256 3578 268
rect 3560 254 3582 256
rect 3587 254 3617 268
rect 3678 266 3831 270
rect 3660 254 3852 266
rect 3895 254 3925 268
rect 3931 254 3944 284
rect 3959 266 3989 284
rect 4032 254 4045 284
rect 4075 254 4088 284
rect 4103 266 4133 284
rect 4176 270 4190 284
rect 4226 270 4446 284
rect 4177 268 4190 270
rect 4143 256 4158 268
rect 4140 254 4162 256
rect 4167 254 4197 268
rect 4258 266 4411 270
rect 4240 254 4432 266
rect 4475 254 4505 268
rect 4511 254 4524 284
rect 4539 266 4569 284
rect 4612 254 4625 284
rect 0 240 4625 254
rect 15 136 28 240
rect 73 218 74 228
rect 89 218 102 228
rect 73 214 102 218
rect 107 214 137 240
rect 155 226 171 228
rect 243 226 296 240
rect 244 224 308 226
rect 351 224 366 240
rect 415 237 445 240
rect 415 234 451 237
rect 381 226 397 228
rect 155 214 170 218
rect 73 212 170 214
rect 198 212 366 224
rect 382 214 397 218
rect 415 215 454 234
rect 473 228 480 229
rect 479 221 480 228
rect 463 218 464 221
rect 479 218 492 221
rect 415 214 445 215
rect 454 214 460 215
rect 463 214 492 218
rect 382 213 492 214
rect 382 212 498 213
rect 57 204 108 212
rect 57 192 82 204
rect 89 192 108 204
rect 139 204 189 212
rect 139 196 155 204
rect 162 202 189 204
rect 198 202 419 212
rect 162 192 419 202
rect 448 204 498 212
rect 448 195 464 204
rect 57 184 108 192
rect 155 184 419 192
rect 445 192 464 195
rect 471 192 498 204
rect 445 184 498 192
rect 73 176 74 184
rect 89 176 102 184
rect 73 168 89 176
rect 70 161 89 164
rect 70 152 92 161
rect 43 142 92 152
rect 43 136 73 142
rect 92 137 97 142
rect 15 120 89 136
rect 107 128 137 184
rect 172 174 380 184
rect 415 180 460 184
rect 463 183 464 184
rect 479 183 492 184
rect 198 144 387 174
rect 213 141 387 144
rect 206 138 387 141
rect 15 118 28 120
rect 43 118 77 120
rect 15 102 89 118
rect 116 114 129 128
rect 144 114 160 130
rect 206 125 217 138
rect -1 80 0 96
rect 15 80 28 102
rect 43 80 73 102
rect 116 98 178 114
rect 206 107 217 123
rect 222 118 232 138
rect 242 118 256 138
rect 259 125 268 138
rect 284 125 293 138
rect 222 107 256 118
rect 259 107 268 123
rect 284 107 293 123
rect 300 118 310 138
rect 320 118 334 138
rect 335 125 346 138
rect 300 107 334 118
rect 335 107 346 123
rect 392 114 408 130
rect 415 128 445 180
rect 479 176 480 183
rect 464 168 480 176
rect 451 136 464 155
rect 479 136 509 152
rect 451 120 525 136
rect 451 118 464 120
rect 479 118 513 120
rect 116 96 129 98
rect 144 96 178 98
rect 116 80 178 96
rect 222 91 238 94
rect 300 91 330 102
rect 378 98 424 114
rect 451 102 525 118
rect 378 96 412 98
rect 377 80 424 96
rect 451 80 464 102
rect 479 80 509 102
rect 536 80 537 96
rect 552 80 565 240
rect 595 136 608 240
rect 653 218 654 228
rect 669 218 682 228
rect 653 214 682 218
rect 687 214 717 240
rect 735 226 751 228
rect 823 226 876 240
rect 824 224 888 226
rect 931 224 946 240
rect 995 237 1025 240
rect 995 234 1031 237
rect 961 226 977 228
rect 735 214 750 218
rect 653 212 750 214
rect 778 212 946 224
rect 962 214 977 218
rect 995 215 1034 234
rect 1053 228 1060 229
rect 1059 221 1060 228
rect 1043 218 1044 221
rect 1059 218 1072 221
rect 995 214 1025 215
rect 1034 214 1040 215
rect 1043 214 1072 218
rect 962 213 1072 214
rect 962 212 1078 213
rect 637 204 688 212
rect 637 192 662 204
rect 669 192 688 204
rect 719 204 769 212
rect 719 196 735 204
rect 742 202 769 204
rect 778 202 999 212
rect 742 192 999 202
rect 1028 204 1078 212
rect 1028 195 1044 204
rect 637 184 688 192
rect 735 184 999 192
rect 1025 192 1044 195
rect 1051 192 1078 204
rect 1025 184 1078 192
rect 653 176 654 184
rect 669 176 682 184
rect 653 168 669 176
rect 650 161 669 164
rect 650 152 672 161
rect 623 142 672 152
rect 623 136 653 142
rect 672 137 677 142
rect 595 120 669 136
rect 687 128 717 184
rect 752 174 960 184
rect 995 180 1040 184
rect 1043 183 1044 184
rect 1059 183 1072 184
rect 778 144 967 174
rect 793 141 967 144
rect 786 138 967 141
rect 595 118 608 120
rect 623 118 657 120
rect 595 102 669 118
rect 696 114 709 128
rect 724 114 740 130
rect 786 125 797 138
rect 579 80 580 96
rect 595 80 608 102
rect 623 80 653 102
rect 696 98 758 114
rect 786 107 797 123
rect 802 118 812 138
rect 822 118 836 138
rect 839 125 848 138
rect 864 125 873 138
rect 802 107 836 118
rect 839 107 848 123
rect 864 107 873 123
rect 880 118 890 138
rect 900 118 914 138
rect 915 125 926 138
rect 880 107 914 118
rect 915 107 926 123
rect 972 114 988 130
rect 995 128 1025 180
rect 1059 176 1060 183
rect 1044 168 1060 176
rect 1031 136 1044 155
rect 1059 136 1089 152
rect 1031 120 1105 136
rect 1031 118 1044 120
rect 1059 118 1093 120
rect 696 96 709 98
rect 724 96 758 98
rect 696 80 758 96
rect 802 91 818 94
rect 880 91 910 102
rect 958 98 1004 114
rect 1031 102 1105 118
rect 958 96 992 98
rect 957 80 1004 96
rect 1031 80 1044 102
rect 1059 80 1089 102
rect 1116 80 1117 96
rect 1132 80 1145 240
rect 1175 136 1188 240
rect 1233 218 1234 228
rect 1249 218 1262 228
rect 1233 214 1262 218
rect 1267 214 1297 240
rect 1315 226 1331 228
rect 1403 226 1456 240
rect 1404 224 1468 226
rect 1511 224 1526 240
rect 1575 237 1605 240
rect 1575 234 1611 237
rect 1541 226 1557 228
rect 1315 214 1330 218
rect 1233 212 1330 214
rect 1358 212 1526 224
rect 1542 214 1557 218
rect 1575 215 1614 234
rect 1633 228 1640 229
rect 1639 221 1640 228
rect 1623 218 1624 221
rect 1639 218 1652 221
rect 1575 214 1605 215
rect 1614 214 1620 215
rect 1623 214 1652 218
rect 1542 213 1652 214
rect 1542 212 1658 213
rect 1217 204 1268 212
rect 1217 192 1242 204
rect 1249 192 1268 204
rect 1299 204 1349 212
rect 1299 196 1315 204
rect 1322 202 1349 204
rect 1358 202 1579 212
rect 1322 192 1579 202
rect 1608 204 1658 212
rect 1608 195 1624 204
rect 1217 184 1268 192
rect 1315 184 1579 192
rect 1605 192 1624 195
rect 1631 192 1658 204
rect 1605 184 1658 192
rect 1233 176 1234 184
rect 1249 176 1262 184
rect 1233 168 1249 176
rect 1230 161 1249 164
rect 1230 152 1252 161
rect 1203 142 1252 152
rect 1203 136 1233 142
rect 1252 137 1257 142
rect 1175 120 1249 136
rect 1267 128 1297 184
rect 1332 174 1540 184
rect 1575 180 1620 184
rect 1623 183 1624 184
rect 1639 183 1652 184
rect 1358 144 1547 174
rect 1373 141 1547 144
rect 1366 138 1547 141
rect 1175 118 1188 120
rect 1203 118 1237 120
rect 1175 102 1249 118
rect 1276 114 1289 128
rect 1304 114 1320 130
rect 1366 125 1377 138
rect 1159 80 1160 96
rect 1175 80 1188 102
rect 1203 80 1233 102
rect 1276 98 1338 114
rect 1366 107 1377 123
rect 1382 118 1392 138
rect 1402 118 1416 138
rect 1419 125 1428 138
rect 1444 125 1453 138
rect 1382 107 1416 118
rect 1419 107 1428 123
rect 1444 107 1453 123
rect 1460 118 1470 138
rect 1480 118 1494 138
rect 1495 125 1506 138
rect 1460 107 1494 118
rect 1495 107 1506 123
rect 1552 114 1568 130
rect 1575 128 1605 180
rect 1639 176 1640 183
rect 1624 168 1640 176
rect 1611 136 1624 155
rect 1639 136 1669 152
rect 1611 120 1685 136
rect 1611 118 1624 120
rect 1639 118 1673 120
rect 1276 96 1289 98
rect 1304 96 1338 98
rect 1276 80 1338 96
rect 1382 91 1398 94
rect 1460 91 1490 102
rect 1538 98 1584 114
rect 1611 102 1685 118
rect 1538 96 1572 98
rect 1537 80 1584 96
rect 1611 80 1624 102
rect 1639 80 1669 102
rect 1696 80 1697 96
rect 1712 80 1725 240
rect 1755 136 1768 240
rect 1813 218 1814 228
rect 1829 218 1842 228
rect 1813 214 1842 218
rect 1847 214 1877 240
rect 1895 226 1911 228
rect 1983 226 2036 240
rect 1984 224 2048 226
rect 2091 224 2106 240
rect 2155 237 2185 240
rect 2155 234 2191 237
rect 2121 226 2137 228
rect 1895 214 1910 218
rect 1813 212 1910 214
rect 1938 212 2106 224
rect 2122 214 2137 218
rect 2155 215 2194 234
rect 2213 228 2220 229
rect 2219 221 2220 228
rect 2203 218 2204 221
rect 2219 218 2232 221
rect 2155 214 2185 215
rect 2194 214 2200 215
rect 2203 214 2232 218
rect 2122 213 2232 214
rect 2122 212 2238 213
rect 1797 204 1848 212
rect 1797 192 1822 204
rect 1829 192 1848 204
rect 1879 204 1929 212
rect 1879 196 1895 204
rect 1902 202 1929 204
rect 1938 202 2159 212
rect 1902 192 2159 202
rect 2188 204 2238 212
rect 2188 195 2204 204
rect 1797 184 1848 192
rect 1895 184 2159 192
rect 2185 192 2204 195
rect 2211 192 2238 204
rect 2185 184 2238 192
rect 1813 176 1814 184
rect 1829 176 1842 184
rect 1813 168 1829 176
rect 1810 161 1829 164
rect 1810 152 1832 161
rect 1783 142 1832 152
rect 1783 136 1813 142
rect 1832 137 1837 142
rect 1755 120 1829 136
rect 1847 128 1877 184
rect 1912 174 2120 184
rect 2155 180 2200 184
rect 2203 183 2204 184
rect 2219 183 2232 184
rect 1938 144 2127 174
rect 1953 141 2127 144
rect 1946 138 2127 141
rect 1755 118 1768 120
rect 1783 118 1817 120
rect 1755 102 1829 118
rect 1856 114 1869 128
rect 1884 114 1900 130
rect 1946 125 1957 138
rect 1739 80 1740 96
rect 1755 80 1768 102
rect 1783 80 1813 102
rect 1856 98 1918 114
rect 1946 107 1957 123
rect 1962 118 1972 138
rect 1982 118 1996 138
rect 1999 125 2008 138
rect 2024 125 2033 138
rect 1962 107 1996 118
rect 1999 107 2008 123
rect 2024 107 2033 123
rect 2040 118 2050 138
rect 2060 118 2074 138
rect 2075 125 2086 138
rect 2040 107 2074 118
rect 2075 107 2086 123
rect 2132 114 2148 130
rect 2155 128 2185 180
rect 2219 176 2220 183
rect 2204 168 2220 176
rect 2191 136 2204 155
rect 2219 136 2249 152
rect 2191 120 2265 136
rect 2191 118 2204 120
rect 2219 118 2253 120
rect 1856 96 1869 98
rect 1884 96 1918 98
rect 1856 80 1918 96
rect 1962 91 1978 94
rect 2040 91 2070 102
rect 2118 98 2164 114
rect 2191 102 2265 118
rect 2118 96 2152 98
rect 2117 80 2164 96
rect 2191 80 2204 102
rect 2219 80 2249 102
rect 2276 80 2277 96
rect 2292 80 2305 240
rect 2335 136 2348 240
rect 2393 218 2394 228
rect 2409 218 2422 228
rect 2393 214 2422 218
rect 2427 214 2457 240
rect 2475 226 2491 228
rect 2563 226 2616 240
rect 2564 224 2628 226
rect 2671 224 2686 240
rect 2735 237 2765 240
rect 2735 234 2771 237
rect 2701 226 2717 228
rect 2475 214 2490 218
rect 2393 212 2490 214
rect 2518 212 2686 224
rect 2702 214 2717 218
rect 2735 215 2774 234
rect 2793 228 2800 229
rect 2799 221 2800 228
rect 2783 218 2784 221
rect 2799 218 2812 221
rect 2735 214 2765 215
rect 2774 214 2780 215
rect 2783 214 2812 218
rect 2702 213 2812 214
rect 2702 212 2818 213
rect 2377 204 2428 212
rect 2377 192 2402 204
rect 2409 192 2428 204
rect 2459 204 2509 212
rect 2459 196 2475 204
rect 2482 202 2509 204
rect 2518 202 2739 212
rect 2482 192 2739 202
rect 2768 204 2818 212
rect 2768 195 2784 204
rect 2377 184 2428 192
rect 2475 184 2739 192
rect 2765 192 2784 195
rect 2791 192 2818 204
rect 2765 184 2818 192
rect 2393 176 2394 184
rect 2409 176 2422 184
rect 2393 168 2409 176
rect 2390 161 2409 164
rect 2390 152 2412 161
rect 2363 142 2412 152
rect 2363 136 2393 142
rect 2412 137 2417 142
rect 2335 120 2409 136
rect 2427 128 2457 184
rect 2492 174 2700 184
rect 2735 180 2780 184
rect 2783 183 2784 184
rect 2799 183 2812 184
rect 2518 144 2707 174
rect 2533 141 2707 144
rect 2526 138 2707 141
rect 2335 118 2348 120
rect 2363 118 2397 120
rect 2335 102 2409 118
rect 2436 114 2449 128
rect 2464 114 2480 130
rect 2526 125 2537 138
rect 2319 80 2320 96
rect 2335 80 2348 102
rect 2363 80 2393 102
rect 2436 98 2498 114
rect 2526 107 2537 123
rect 2542 118 2552 138
rect 2562 118 2576 138
rect 2579 125 2588 138
rect 2604 125 2613 138
rect 2542 107 2576 118
rect 2579 107 2588 123
rect 2604 107 2613 123
rect 2620 118 2630 138
rect 2640 118 2654 138
rect 2655 125 2666 138
rect 2620 107 2654 118
rect 2655 107 2666 123
rect 2712 114 2728 130
rect 2735 128 2765 180
rect 2799 176 2800 183
rect 2784 168 2800 176
rect 2771 136 2784 155
rect 2799 136 2829 152
rect 2771 120 2845 136
rect 2771 118 2784 120
rect 2799 118 2833 120
rect 2436 96 2449 98
rect 2464 96 2498 98
rect 2436 80 2498 96
rect 2542 91 2558 94
rect 2620 91 2650 102
rect 2698 98 2744 114
rect 2771 102 2845 118
rect 2698 96 2732 98
rect 2697 80 2744 96
rect 2771 80 2784 102
rect 2799 80 2829 102
rect 2856 80 2857 96
rect 2872 80 2885 240
rect 2915 136 2928 240
rect 2973 218 2974 228
rect 2989 218 3002 228
rect 2973 214 3002 218
rect 3007 214 3037 240
rect 3055 226 3071 228
rect 3143 226 3196 240
rect 3144 224 3208 226
rect 3251 224 3266 240
rect 3315 237 3345 240
rect 3315 234 3351 237
rect 3281 226 3297 228
rect 3055 214 3070 218
rect 2973 212 3070 214
rect 3098 212 3266 224
rect 3282 214 3297 218
rect 3315 215 3354 234
rect 3373 228 3380 229
rect 3379 221 3380 228
rect 3363 218 3364 221
rect 3379 218 3392 221
rect 3315 214 3345 215
rect 3354 214 3360 215
rect 3363 214 3392 218
rect 3282 213 3392 214
rect 3282 212 3398 213
rect 2957 204 3008 212
rect 2957 192 2982 204
rect 2989 192 3008 204
rect 3039 204 3089 212
rect 3039 196 3055 204
rect 3062 202 3089 204
rect 3098 202 3319 212
rect 3062 192 3319 202
rect 3348 204 3398 212
rect 3348 195 3364 204
rect 2957 184 3008 192
rect 3055 184 3319 192
rect 3345 192 3364 195
rect 3371 192 3398 204
rect 3345 184 3398 192
rect 2973 176 2974 184
rect 2989 176 3002 184
rect 2973 168 2989 176
rect 2970 161 2989 164
rect 2970 152 2992 161
rect 2943 142 2992 152
rect 2943 136 2973 142
rect 2992 137 2997 142
rect 2915 120 2989 136
rect 3007 128 3037 184
rect 3072 174 3280 184
rect 3315 180 3360 184
rect 3363 183 3364 184
rect 3379 183 3392 184
rect 3098 144 3287 174
rect 3113 141 3287 144
rect 3106 138 3287 141
rect 2915 118 2928 120
rect 2943 118 2977 120
rect 2915 102 2989 118
rect 3016 114 3029 128
rect 3044 114 3060 130
rect 3106 125 3117 138
rect 2899 80 2900 96
rect 2915 80 2928 102
rect 2943 80 2973 102
rect 3016 98 3078 114
rect 3106 107 3117 123
rect 3122 118 3132 138
rect 3142 118 3156 138
rect 3159 125 3168 138
rect 3184 125 3193 138
rect 3122 107 3156 118
rect 3159 107 3168 123
rect 3184 107 3193 123
rect 3200 118 3210 138
rect 3220 118 3234 138
rect 3235 125 3246 138
rect 3200 107 3234 118
rect 3235 107 3246 123
rect 3292 114 3308 130
rect 3315 128 3345 180
rect 3379 176 3380 183
rect 3364 168 3380 176
rect 3351 136 3364 155
rect 3379 136 3409 152
rect 3351 120 3425 136
rect 3351 118 3364 120
rect 3379 118 3413 120
rect 3016 96 3029 98
rect 3044 96 3078 98
rect 3016 80 3078 96
rect 3122 91 3138 94
rect 3200 91 3230 102
rect 3278 98 3324 114
rect 3351 102 3425 118
rect 3278 96 3312 98
rect 3277 80 3324 96
rect 3351 80 3364 102
rect 3379 80 3409 102
rect 3436 80 3437 96
rect 3452 80 3465 240
rect 3495 136 3508 240
rect 3553 218 3554 228
rect 3569 218 3582 228
rect 3553 214 3582 218
rect 3587 214 3617 240
rect 3635 226 3651 228
rect 3723 226 3776 240
rect 3724 224 3788 226
rect 3831 224 3846 240
rect 3895 237 3925 240
rect 3895 234 3931 237
rect 3861 226 3877 228
rect 3635 214 3650 218
rect 3553 212 3650 214
rect 3678 212 3846 224
rect 3862 214 3877 218
rect 3895 215 3934 234
rect 3953 228 3960 229
rect 3959 221 3960 228
rect 3943 218 3944 221
rect 3959 218 3972 221
rect 3895 214 3925 215
rect 3934 214 3940 215
rect 3943 214 3972 218
rect 3862 213 3972 214
rect 3862 212 3978 213
rect 3537 204 3588 212
rect 3537 192 3562 204
rect 3569 192 3588 204
rect 3619 204 3669 212
rect 3619 196 3635 204
rect 3642 202 3669 204
rect 3678 202 3899 212
rect 3642 192 3899 202
rect 3928 204 3978 212
rect 3928 195 3944 204
rect 3537 184 3588 192
rect 3635 184 3899 192
rect 3925 192 3944 195
rect 3951 192 3978 204
rect 3925 184 3978 192
rect 3553 176 3554 184
rect 3569 176 3582 184
rect 3553 168 3569 176
rect 3550 161 3569 164
rect 3550 152 3572 161
rect 3523 142 3572 152
rect 3523 136 3553 142
rect 3572 137 3577 142
rect 3495 120 3569 136
rect 3587 128 3617 184
rect 3652 174 3860 184
rect 3895 180 3940 184
rect 3943 183 3944 184
rect 3959 183 3972 184
rect 3678 144 3867 174
rect 3693 141 3867 144
rect 3686 138 3867 141
rect 3495 118 3508 120
rect 3523 118 3557 120
rect 3495 102 3569 118
rect 3596 114 3609 128
rect 3624 114 3640 130
rect 3686 125 3697 138
rect 3479 80 3480 96
rect 3495 80 3508 102
rect 3523 80 3553 102
rect 3596 98 3658 114
rect 3686 107 3697 123
rect 3702 118 3712 138
rect 3722 118 3736 138
rect 3739 125 3748 138
rect 3764 125 3773 138
rect 3702 107 3736 118
rect 3739 107 3748 123
rect 3764 107 3773 123
rect 3780 118 3790 138
rect 3800 118 3814 138
rect 3815 125 3826 138
rect 3780 107 3814 118
rect 3815 107 3826 123
rect 3872 114 3888 130
rect 3895 128 3925 180
rect 3959 176 3960 183
rect 3944 168 3960 176
rect 3931 136 3944 155
rect 3959 136 3989 152
rect 3931 120 4005 136
rect 3931 118 3944 120
rect 3959 118 3993 120
rect 3596 96 3609 98
rect 3624 96 3658 98
rect 3596 80 3658 96
rect 3702 91 3718 94
rect 3780 91 3810 102
rect 3858 98 3904 114
rect 3931 102 4005 118
rect 3858 96 3892 98
rect 3857 80 3904 96
rect 3931 80 3944 102
rect 3959 80 3989 102
rect 4016 80 4017 96
rect 4032 80 4045 240
rect 4075 136 4088 240
rect 4133 218 4134 228
rect 4149 218 4162 228
rect 4133 214 4162 218
rect 4167 214 4197 240
rect 4215 226 4231 228
rect 4303 226 4356 240
rect 4304 224 4368 226
rect 4411 224 4426 240
rect 4475 237 4505 240
rect 4475 234 4511 237
rect 4441 226 4457 228
rect 4215 214 4230 218
rect 4133 212 4230 214
rect 4258 212 4426 224
rect 4442 214 4457 218
rect 4475 215 4514 234
rect 4533 228 4540 229
rect 4539 221 4540 228
rect 4523 218 4524 221
rect 4539 218 4552 221
rect 4475 214 4505 215
rect 4514 214 4520 215
rect 4523 214 4552 218
rect 4442 213 4552 214
rect 4442 212 4558 213
rect 4117 204 4168 212
rect 4117 192 4142 204
rect 4149 192 4168 204
rect 4199 204 4249 212
rect 4199 196 4215 204
rect 4222 202 4249 204
rect 4258 202 4479 212
rect 4222 192 4479 202
rect 4508 204 4558 212
rect 4508 195 4524 204
rect 4117 184 4168 192
rect 4215 184 4479 192
rect 4505 192 4524 195
rect 4531 192 4558 204
rect 4505 184 4558 192
rect 4133 176 4134 184
rect 4149 176 4162 184
rect 4133 168 4149 176
rect 4130 161 4149 164
rect 4130 152 4152 161
rect 4103 142 4152 152
rect 4103 136 4133 142
rect 4152 137 4157 142
rect 4075 120 4149 136
rect 4167 128 4197 184
rect 4232 174 4440 184
rect 4475 180 4520 184
rect 4523 183 4524 184
rect 4539 183 4552 184
rect 4258 144 4447 174
rect 4273 141 4447 144
rect 4266 138 4447 141
rect 4075 118 4088 120
rect 4103 118 4137 120
rect 4075 102 4149 118
rect 4176 114 4189 128
rect 4204 114 4220 130
rect 4266 125 4277 138
rect 4059 80 4060 96
rect 4075 80 4088 102
rect 4103 80 4133 102
rect 4176 98 4238 114
rect 4266 107 4277 123
rect 4282 118 4292 138
rect 4302 118 4316 138
rect 4319 125 4328 138
rect 4344 125 4353 138
rect 4282 107 4316 118
rect 4319 107 4328 123
rect 4344 107 4353 123
rect 4360 118 4370 138
rect 4380 118 4394 138
rect 4395 125 4406 138
rect 4360 107 4394 118
rect 4395 107 4406 123
rect 4452 114 4468 130
rect 4475 128 4505 180
rect 4539 176 4540 183
rect 4524 168 4540 176
rect 4511 136 4524 155
rect 4539 136 4569 152
rect 4511 120 4585 136
rect 4511 118 4524 120
rect 4539 118 4573 120
rect 4176 96 4189 98
rect 4204 96 4238 98
rect 4176 80 4238 96
rect 4282 91 4298 94
rect 4360 91 4390 102
rect 4438 98 4484 114
rect 4511 102 4585 118
rect 4438 96 4472 98
rect 4437 80 4484 96
rect 4511 80 4524 102
rect 4539 80 4569 102
rect 4596 80 4597 96
rect 4612 80 4625 240
rect -7 72 34 80
rect -7 46 8 72
rect 15 46 34 72
rect 98 68 160 80
rect 172 68 247 80
rect 305 68 380 80
rect 392 68 423 80
rect 429 68 464 80
rect 98 66 260 68
rect -7 38 34 46
rect 116 42 129 66
rect 144 64 159 66
rect -1 28 0 38
rect 15 28 28 38
rect 43 28 73 42
rect 116 28 159 42
rect 183 39 190 46
rect 193 42 260 66
rect 292 66 464 68
rect 262 44 290 48
rect 292 44 372 66
rect 393 64 408 66
rect 262 42 372 44
rect 193 38 372 42
rect 166 28 196 38
rect 198 28 351 38
rect 359 28 389 38
rect 393 28 423 42
rect 451 28 464 66
rect 536 72 571 80
rect 536 46 537 72
rect 544 46 571 72
rect 479 28 509 42
rect 536 38 571 46
rect 573 72 614 80
rect 573 46 588 72
rect 595 46 614 72
rect 678 68 740 80
rect 752 68 827 80
rect 885 68 960 80
rect 972 68 1003 80
rect 1009 68 1044 80
rect 678 66 840 68
rect 573 38 614 46
rect 696 42 709 66
rect 724 64 739 66
rect 536 28 537 38
rect 552 28 565 38
rect 579 28 580 38
rect 595 28 608 38
rect 623 28 653 42
rect 696 28 739 42
rect 763 39 770 46
rect 773 42 840 66
rect 872 66 1044 68
rect 842 44 870 48
rect 872 44 952 66
rect 973 64 988 66
rect 842 42 952 44
rect 773 38 952 42
rect 746 28 776 38
rect 778 28 931 38
rect 939 28 969 38
rect 973 28 1003 42
rect 1031 28 1044 66
rect 1116 72 1151 80
rect 1116 46 1117 72
rect 1124 46 1151 72
rect 1059 28 1089 42
rect 1116 38 1151 46
rect 1153 72 1194 80
rect 1153 46 1168 72
rect 1175 46 1194 72
rect 1258 68 1320 80
rect 1332 68 1407 80
rect 1465 68 1540 80
rect 1552 68 1583 80
rect 1589 68 1624 80
rect 1258 66 1420 68
rect 1153 38 1194 46
rect 1276 42 1289 66
rect 1304 64 1319 66
rect 1116 28 1117 38
rect 1132 28 1145 38
rect 1159 28 1160 38
rect 1175 28 1188 38
rect 1203 28 1233 42
rect 1276 28 1319 42
rect 1343 39 1350 46
rect 1353 42 1420 66
rect 1452 66 1624 68
rect 1422 44 1450 48
rect 1452 44 1532 66
rect 1553 64 1568 66
rect 1422 42 1532 44
rect 1353 38 1532 42
rect 1326 28 1356 38
rect 1358 28 1511 38
rect 1519 28 1549 38
rect 1553 28 1583 42
rect 1611 28 1624 66
rect 1696 72 1731 80
rect 1696 46 1697 72
rect 1704 46 1731 72
rect 1639 28 1669 42
rect 1696 38 1731 46
rect 1733 72 1774 80
rect 1733 46 1748 72
rect 1755 46 1774 72
rect 1838 68 1900 80
rect 1912 68 1987 80
rect 2045 68 2120 80
rect 2132 68 2163 80
rect 2169 68 2204 80
rect 1838 66 2000 68
rect 1733 38 1774 46
rect 1856 42 1869 66
rect 1884 64 1899 66
rect 1696 28 1697 38
rect 1712 28 1725 38
rect 1739 28 1740 38
rect 1755 28 1768 38
rect 1783 28 1813 42
rect 1856 28 1899 42
rect 1923 39 1930 46
rect 1933 42 2000 66
rect 2032 66 2204 68
rect 2002 44 2030 48
rect 2032 44 2112 66
rect 2133 64 2148 66
rect 2002 42 2112 44
rect 1933 38 2112 42
rect 1906 28 1936 38
rect 1938 28 2091 38
rect 2099 28 2129 38
rect 2133 28 2163 42
rect 2191 28 2204 66
rect 2276 72 2311 80
rect 2276 46 2277 72
rect 2284 46 2311 72
rect 2219 28 2249 42
rect 2276 38 2311 46
rect 2313 72 2354 80
rect 2313 46 2328 72
rect 2335 46 2354 72
rect 2418 68 2480 80
rect 2492 68 2567 80
rect 2625 68 2700 80
rect 2712 68 2743 80
rect 2749 68 2784 80
rect 2418 66 2580 68
rect 2313 38 2354 46
rect 2436 42 2449 66
rect 2464 64 2479 66
rect 2276 28 2277 38
rect 2292 28 2305 38
rect 2319 28 2320 38
rect 2335 28 2348 38
rect 2363 28 2393 42
rect 2436 28 2479 42
rect 2503 39 2510 46
rect 2513 42 2580 66
rect 2612 66 2784 68
rect 2582 44 2610 48
rect 2612 44 2692 66
rect 2713 64 2728 66
rect 2582 42 2692 44
rect 2513 38 2692 42
rect 2486 28 2516 38
rect 2518 28 2671 38
rect 2679 28 2709 38
rect 2713 28 2743 42
rect 2771 28 2784 66
rect 2856 72 2891 80
rect 2856 46 2857 72
rect 2864 46 2891 72
rect 2799 28 2829 42
rect 2856 38 2891 46
rect 2893 72 2934 80
rect 2893 46 2908 72
rect 2915 46 2934 72
rect 2998 68 3060 80
rect 3072 68 3147 80
rect 3205 68 3280 80
rect 3292 68 3323 80
rect 3329 68 3364 80
rect 2998 66 3160 68
rect 2893 38 2934 46
rect 3016 42 3029 66
rect 3044 64 3059 66
rect 2856 28 2857 38
rect 2872 28 2885 38
rect 2899 28 2900 38
rect 2915 28 2928 38
rect 2943 28 2973 42
rect 3016 28 3059 42
rect 3083 39 3090 46
rect 3093 42 3160 66
rect 3192 66 3364 68
rect 3162 44 3190 48
rect 3192 44 3272 66
rect 3293 64 3308 66
rect 3162 42 3272 44
rect 3093 38 3272 42
rect 3066 28 3096 38
rect 3098 28 3251 38
rect 3259 28 3289 38
rect 3293 28 3323 42
rect 3351 28 3364 66
rect 3436 72 3471 80
rect 3436 46 3437 72
rect 3444 46 3471 72
rect 3379 28 3409 42
rect 3436 38 3471 46
rect 3473 72 3514 80
rect 3473 46 3488 72
rect 3495 46 3514 72
rect 3578 68 3640 80
rect 3652 68 3727 80
rect 3785 68 3860 80
rect 3872 68 3903 80
rect 3909 68 3944 80
rect 3578 66 3740 68
rect 3473 38 3514 46
rect 3596 42 3609 66
rect 3624 64 3639 66
rect 3436 28 3437 38
rect 3452 28 3465 38
rect 3479 28 3480 38
rect 3495 28 3508 38
rect 3523 28 3553 42
rect 3596 28 3639 42
rect 3663 39 3670 46
rect 3673 42 3740 66
rect 3772 66 3944 68
rect 3742 44 3770 48
rect 3772 44 3852 66
rect 3873 64 3888 66
rect 3742 42 3852 44
rect 3673 38 3852 42
rect 3646 28 3676 38
rect 3678 28 3831 38
rect 3839 28 3869 38
rect 3873 28 3903 42
rect 3931 28 3944 66
rect 4016 72 4051 80
rect 4016 46 4017 72
rect 4024 46 4051 72
rect 3959 28 3989 42
rect 4016 38 4051 46
rect 4053 72 4094 80
rect 4053 46 4068 72
rect 4075 46 4094 72
rect 4158 68 4220 80
rect 4232 68 4307 80
rect 4365 68 4440 80
rect 4452 68 4483 80
rect 4489 68 4524 80
rect 4158 66 4320 68
rect 4053 38 4094 46
rect 4176 42 4189 66
rect 4204 64 4219 66
rect 4016 28 4017 38
rect 4032 28 4045 38
rect 4059 28 4060 38
rect 4075 28 4088 38
rect 4103 28 4133 42
rect 4176 28 4219 42
rect 4243 39 4250 46
rect 4253 42 4320 66
rect 4352 66 4524 68
rect 4322 44 4350 48
rect 4352 44 4432 66
rect 4453 64 4468 66
rect 4322 42 4432 44
rect 4253 38 4432 42
rect 4226 28 4256 38
rect 4258 28 4411 38
rect 4419 28 4449 38
rect 4453 28 4483 42
rect 4511 28 4524 66
rect 4596 72 4631 80
rect 4596 46 4597 72
rect 4604 46 4631 72
rect 4539 28 4569 42
rect 4596 38 4631 46
rect 4596 28 4597 38
rect 4612 28 4625 38
rect -1 22 4625 28
rect 0 14 4625 22
rect 15 -16 28 14
rect 43 -4 73 14
rect 116 0 130 14
rect 166 0 386 14
rect 117 -2 130 0
rect 83 -14 98 -2
rect 80 -16 102 -14
rect 107 -16 137 -2
rect 198 -4 351 0
rect 180 -16 372 -4
rect 415 -16 445 -2
rect 451 -16 464 14
rect 479 -4 509 14
rect 552 -16 565 14
rect 595 -16 608 14
rect 623 -4 653 14
rect 696 0 710 14
rect 746 0 966 14
rect 697 -2 710 0
rect 663 -14 678 -2
rect 660 -16 682 -14
rect 687 -16 717 -2
rect 778 -4 931 0
rect 760 -16 952 -4
rect 995 -16 1025 -2
rect 1031 -16 1044 14
rect 1059 -4 1089 14
rect 1132 -16 1145 14
rect 1175 -16 1188 14
rect 1203 -4 1233 14
rect 1276 0 1290 14
rect 1326 0 1546 14
rect 1277 -2 1290 0
rect 1243 -14 1258 -2
rect 1240 -16 1262 -14
rect 1267 -16 1297 -2
rect 1358 -4 1511 0
rect 1340 -16 1532 -4
rect 1575 -16 1605 -2
rect 1611 -16 1624 14
rect 1639 -4 1669 14
rect 1712 -16 1725 14
rect 1755 -16 1768 14
rect 1783 -4 1813 14
rect 1856 0 1870 14
rect 1906 0 2126 14
rect 1857 -2 1870 0
rect 1823 -14 1838 -2
rect 1820 -16 1842 -14
rect 1847 -16 1877 -2
rect 1938 -4 2091 0
rect 1920 -16 2112 -4
rect 2155 -16 2185 -2
rect 2191 -16 2204 14
rect 2219 -4 2249 14
rect 2292 -16 2305 14
rect 2335 -16 2348 14
rect 2363 -4 2393 14
rect 2436 0 2450 14
rect 2486 0 2706 14
rect 2437 -2 2450 0
rect 2403 -14 2418 -2
rect 2400 -16 2422 -14
rect 2427 -16 2457 -2
rect 2518 -4 2671 0
rect 2500 -16 2692 -4
rect 2735 -16 2765 -2
rect 2771 -16 2784 14
rect 2799 -4 2829 14
rect 2872 -16 2885 14
rect 2915 -16 2928 14
rect 2943 -4 2973 14
rect 3016 0 3030 14
rect 3066 0 3286 14
rect 3017 -2 3030 0
rect 2983 -14 2998 -2
rect 2980 -16 3002 -14
rect 3007 -16 3037 -2
rect 3098 -4 3251 0
rect 3080 -16 3272 -4
rect 3315 -16 3345 -2
rect 3351 -16 3364 14
rect 3379 -4 3409 14
rect 3452 -16 3465 14
rect 3495 -16 3508 14
rect 3523 -4 3553 14
rect 3596 0 3610 14
rect 3646 0 3866 14
rect 3597 -2 3610 0
rect 3563 -14 3578 -2
rect 3560 -16 3582 -14
rect 3587 -16 3617 -2
rect 3678 -4 3831 0
rect 3660 -16 3852 -4
rect 3895 -16 3925 -2
rect 3931 -16 3944 14
rect 3959 -4 3989 14
rect 4032 -16 4045 14
rect 4075 -16 4088 14
rect 4103 -4 4133 14
rect 4176 0 4190 14
rect 4226 0 4446 14
rect 4177 -2 4190 0
rect 4143 -14 4158 -2
rect 4140 -16 4162 -14
rect 4167 -16 4197 -2
rect 4258 -4 4411 0
rect 4240 -16 4432 -4
rect 4475 -16 4505 -2
rect 4511 -16 4524 14
rect 4539 -4 4569 14
rect 4612 -16 4625 14
rect 0 -30 4625 -16
rect 15 -134 28 -30
rect 73 -52 74 -42
rect 89 -52 102 -42
rect 73 -56 102 -52
rect 107 -56 137 -30
rect 155 -44 171 -42
rect 243 -44 296 -30
rect 244 -46 308 -44
rect 351 -46 366 -30
rect 415 -33 445 -30
rect 415 -36 451 -33
rect 381 -44 397 -42
rect 155 -56 170 -52
rect 73 -58 170 -56
rect 198 -58 366 -46
rect 382 -56 397 -52
rect 415 -55 454 -36
rect 473 -42 480 -41
rect 479 -49 480 -42
rect 463 -52 464 -49
rect 479 -52 492 -49
rect 415 -56 445 -55
rect 454 -56 460 -55
rect 463 -56 492 -52
rect 382 -57 492 -56
rect 382 -58 498 -57
rect 57 -66 108 -58
rect 57 -78 82 -66
rect 89 -78 108 -66
rect 139 -66 189 -58
rect 139 -74 155 -66
rect 162 -68 189 -66
rect 198 -68 419 -58
rect 162 -78 419 -68
rect 448 -66 498 -58
rect 448 -75 464 -66
rect 57 -86 108 -78
rect 155 -86 419 -78
rect 445 -78 464 -75
rect 471 -78 498 -66
rect 445 -86 498 -78
rect 73 -94 74 -86
rect 89 -94 102 -86
rect 73 -102 89 -94
rect 70 -109 89 -106
rect 70 -118 92 -109
rect 43 -128 92 -118
rect 43 -134 73 -128
rect 92 -133 97 -128
rect 15 -150 89 -134
rect 107 -142 137 -86
rect 172 -96 380 -86
rect 415 -90 460 -86
rect 463 -87 464 -86
rect 479 -87 492 -86
rect 198 -126 387 -96
rect 213 -129 387 -126
rect 206 -132 387 -129
rect 15 -152 28 -150
rect 43 -152 77 -150
rect 15 -168 89 -152
rect 116 -156 129 -142
rect 144 -156 160 -140
rect 206 -145 217 -132
rect -1 -190 0 -174
rect 15 -190 28 -168
rect 43 -190 73 -168
rect 116 -172 178 -156
rect 206 -163 217 -147
rect 222 -152 232 -132
rect 242 -152 256 -132
rect 259 -145 268 -132
rect 284 -145 293 -132
rect 222 -163 256 -152
rect 259 -163 268 -147
rect 284 -163 293 -147
rect 300 -152 310 -132
rect 320 -152 334 -132
rect 335 -145 346 -132
rect 300 -163 334 -152
rect 335 -163 346 -147
rect 392 -156 408 -140
rect 415 -142 445 -90
rect 479 -94 480 -87
rect 464 -102 480 -94
rect 451 -134 464 -115
rect 479 -134 509 -118
rect 451 -150 525 -134
rect 451 -152 464 -150
rect 479 -152 513 -150
rect 116 -174 129 -172
rect 144 -174 178 -172
rect 116 -190 178 -174
rect 222 -179 238 -176
rect 300 -179 330 -168
rect 378 -172 424 -156
rect 451 -168 525 -152
rect 378 -174 412 -172
rect 377 -190 424 -174
rect 451 -190 464 -168
rect 479 -190 509 -168
rect 536 -190 537 -174
rect 552 -190 565 -30
rect 595 -134 608 -30
rect 653 -52 654 -42
rect 669 -52 682 -42
rect 653 -56 682 -52
rect 687 -56 717 -30
rect 735 -44 751 -42
rect 823 -44 876 -30
rect 824 -46 888 -44
rect 931 -46 946 -30
rect 995 -33 1025 -30
rect 995 -36 1031 -33
rect 961 -44 977 -42
rect 735 -56 750 -52
rect 653 -58 750 -56
rect 778 -58 946 -46
rect 962 -56 977 -52
rect 995 -55 1034 -36
rect 1053 -42 1060 -41
rect 1059 -49 1060 -42
rect 1043 -52 1044 -49
rect 1059 -52 1072 -49
rect 995 -56 1025 -55
rect 1034 -56 1040 -55
rect 1043 -56 1072 -52
rect 962 -57 1072 -56
rect 962 -58 1078 -57
rect 637 -66 688 -58
rect 637 -78 662 -66
rect 669 -78 688 -66
rect 719 -66 769 -58
rect 719 -74 735 -66
rect 742 -68 769 -66
rect 778 -68 999 -58
rect 742 -78 999 -68
rect 1028 -66 1078 -58
rect 1028 -75 1044 -66
rect 637 -86 688 -78
rect 735 -86 999 -78
rect 1025 -78 1044 -75
rect 1051 -78 1078 -66
rect 1025 -86 1078 -78
rect 653 -94 654 -86
rect 669 -94 682 -86
rect 653 -102 669 -94
rect 650 -109 669 -106
rect 650 -118 672 -109
rect 623 -128 672 -118
rect 623 -134 653 -128
rect 672 -133 677 -128
rect 595 -150 669 -134
rect 687 -142 717 -86
rect 752 -96 960 -86
rect 995 -90 1040 -86
rect 1043 -87 1044 -86
rect 1059 -87 1072 -86
rect 778 -126 967 -96
rect 793 -129 967 -126
rect 786 -132 967 -129
rect 595 -152 608 -150
rect 623 -152 657 -150
rect 595 -168 669 -152
rect 696 -156 709 -142
rect 724 -156 740 -140
rect 786 -145 797 -132
rect 579 -190 580 -174
rect 595 -190 608 -168
rect 623 -190 653 -168
rect 696 -172 758 -156
rect 786 -163 797 -147
rect 802 -152 812 -132
rect 822 -152 836 -132
rect 839 -145 848 -132
rect 864 -145 873 -132
rect 802 -163 836 -152
rect 839 -163 848 -147
rect 864 -163 873 -147
rect 880 -152 890 -132
rect 900 -152 914 -132
rect 915 -145 926 -132
rect 880 -163 914 -152
rect 915 -163 926 -147
rect 972 -156 988 -140
rect 995 -142 1025 -90
rect 1059 -94 1060 -87
rect 1044 -102 1060 -94
rect 1031 -134 1044 -115
rect 1059 -134 1089 -118
rect 1031 -150 1105 -134
rect 1031 -152 1044 -150
rect 1059 -152 1093 -150
rect 696 -174 709 -172
rect 724 -174 758 -172
rect 696 -190 758 -174
rect 802 -179 818 -176
rect 880 -179 910 -168
rect 958 -172 1004 -156
rect 1031 -168 1105 -152
rect 958 -174 992 -172
rect 957 -190 1004 -174
rect 1031 -190 1044 -168
rect 1059 -190 1089 -168
rect 1116 -190 1117 -174
rect 1132 -190 1145 -30
rect 1175 -134 1188 -30
rect 1233 -52 1234 -42
rect 1249 -52 1262 -42
rect 1233 -56 1262 -52
rect 1267 -56 1297 -30
rect 1315 -44 1331 -42
rect 1403 -44 1456 -30
rect 1404 -46 1468 -44
rect 1511 -46 1526 -30
rect 1575 -33 1605 -30
rect 1575 -36 1611 -33
rect 1541 -44 1557 -42
rect 1315 -56 1330 -52
rect 1233 -58 1330 -56
rect 1358 -58 1526 -46
rect 1542 -56 1557 -52
rect 1575 -55 1614 -36
rect 1633 -42 1640 -41
rect 1639 -49 1640 -42
rect 1623 -52 1624 -49
rect 1639 -52 1652 -49
rect 1575 -56 1605 -55
rect 1614 -56 1620 -55
rect 1623 -56 1652 -52
rect 1542 -57 1652 -56
rect 1542 -58 1658 -57
rect 1217 -66 1268 -58
rect 1217 -78 1242 -66
rect 1249 -78 1268 -66
rect 1299 -66 1349 -58
rect 1299 -74 1315 -66
rect 1322 -68 1349 -66
rect 1358 -68 1579 -58
rect 1322 -78 1579 -68
rect 1608 -66 1658 -58
rect 1608 -75 1624 -66
rect 1217 -86 1268 -78
rect 1315 -86 1579 -78
rect 1605 -78 1624 -75
rect 1631 -78 1658 -66
rect 1605 -86 1658 -78
rect 1233 -94 1234 -86
rect 1249 -94 1262 -86
rect 1233 -102 1249 -94
rect 1230 -109 1249 -106
rect 1230 -118 1252 -109
rect 1203 -128 1252 -118
rect 1203 -134 1233 -128
rect 1252 -133 1257 -128
rect 1175 -150 1249 -134
rect 1267 -142 1297 -86
rect 1332 -96 1540 -86
rect 1575 -90 1620 -86
rect 1623 -87 1624 -86
rect 1639 -87 1652 -86
rect 1358 -126 1547 -96
rect 1373 -129 1547 -126
rect 1366 -132 1547 -129
rect 1175 -152 1188 -150
rect 1203 -152 1237 -150
rect 1175 -168 1249 -152
rect 1276 -156 1289 -142
rect 1304 -156 1320 -140
rect 1366 -145 1377 -132
rect 1159 -190 1160 -174
rect 1175 -190 1188 -168
rect 1203 -190 1233 -168
rect 1276 -172 1338 -156
rect 1366 -163 1377 -147
rect 1382 -152 1392 -132
rect 1402 -152 1416 -132
rect 1419 -145 1428 -132
rect 1444 -145 1453 -132
rect 1382 -163 1416 -152
rect 1419 -163 1428 -147
rect 1444 -163 1453 -147
rect 1460 -152 1470 -132
rect 1480 -152 1494 -132
rect 1495 -145 1506 -132
rect 1460 -163 1494 -152
rect 1495 -163 1506 -147
rect 1552 -156 1568 -140
rect 1575 -142 1605 -90
rect 1639 -94 1640 -87
rect 1624 -102 1640 -94
rect 1611 -134 1624 -115
rect 1639 -134 1669 -118
rect 1611 -150 1685 -134
rect 1611 -152 1624 -150
rect 1639 -152 1673 -150
rect 1276 -174 1289 -172
rect 1304 -174 1338 -172
rect 1276 -190 1338 -174
rect 1382 -179 1398 -176
rect 1460 -179 1490 -168
rect 1538 -172 1584 -156
rect 1611 -168 1685 -152
rect 1538 -174 1572 -172
rect 1537 -190 1584 -174
rect 1611 -190 1624 -168
rect 1639 -190 1669 -168
rect 1696 -190 1697 -174
rect 1712 -190 1725 -30
rect 1755 -134 1768 -30
rect 1813 -52 1814 -42
rect 1829 -52 1842 -42
rect 1813 -56 1842 -52
rect 1847 -56 1877 -30
rect 1895 -44 1911 -42
rect 1983 -44 2036 -30
rect 1984 -46 2048 -44
rect 2091 -46 2106 -30
rect 2155 -33 2185 -30
rect 2155 -36 2191 -33
rect 2121 -44 2137 -42
rect 1895 -56 1910 -52
rect 1813 -58 1910 -56
rect 1938 -58 2106 -46
rect 2122 -56 2137 -52
rect 2155 -55 2194 -36
rect 2213 -42 2220 -41
rect 2219 -49 2220 -42
rect 2203 -52 2204 -49
rect 2219 -52 2232 -49
rect 2155 -56 2185 -55
rect 2194 -56 2200 -55
rect 2203 -56 2232 -52
rect 2122 -57 2232 -56
rect 2122 -58 2238 -57
rect 1797 -66 1848 -58
rect 1797 -78 1822 -66
rect 1829 -78 1848 -66
rect 1879 -66 1929 -58
rect 1879 -74 1895 -66
rect 1902 -68 1929 -66
rect 1938 -68 2159 -58
rect 1902 -78 2159 -68
rect 2188 -66 2238 -58
rect 2188 -75 2204 -66
rect 1797 -86 1848 -78
rect 1895 -86 2159 -78
rect 2185 -78 2204 -75
rect 2211 -78 2238 -66
rect 2185 -86 2238 -78
rect 1813 -94 1814 -86
rect 1829 -94 1842 -86
rect 1813 -102 1829 -94
rect 1810 -109 1829 -106
rect 1810 -118 1832 -109
rect 1783 -128 1832 -118
rect 1783 -134 1813 -128
rect 1832 -133 1837 -128
rect 1755 -150 1829 -134
rect 1847 -142 1877 -86
rect 1912 -96 2120 -86
rect 2155 -90 2200 -86
rect 2203 -87 2204 -86
rect 2219 -87 2232 -86
rect 1938 -126 2127 -96
rect 1953 -129 2127 -126
rect 1946 -132 2127 -129
rect 1755 -152 1768 -150
rect 1783 -152 1817 -150
rect 1755 -168 1829 -152
rect 1856 -156 1869 -142
rect 1884 -156 1900 -140
rect 1946 -145 1957 -132
rect 1739 -190 1740 -174
rect 1755 -190 1768 -168
rect 1783 -190 1813 -168
rect 1856 -172 1918 -156
rect 1946 -163 1957 -147
rect 1962 -152 1972 -132
rect 1982 -152 1996 -132
rect 1999 -145 2008 -132
rect 2024 -145 2033 -132
rect 1962 -163 1996 -152
rect 1999 -163 2008 -147
rect 2024 -163 2033 -147
rect 2040 -152 2050 -132
rect 2060 -152 2074 -132
rect 2075 -145 2086 -132
rect 2040 -163 2074 -152
rect 2075 -163 2086 -147
rect 2132 -156 2148 -140
rect 2155 -142 2185 -90
rect 2219 -94 2220 -87
rect 2204 -102 2220 -94
rect 2191 -134 2204 -115
rect 2219 -134 2249 -118
rect 2191 -150 2265 -134
rect 2191 -152 2204 -150
rect 2219 -152 2253 -150
rect 1856 -174 1869 -172
rect 1884 -174 1918 -172
rect 1856 -190 1918 -174
rect 1962 -179 1978 -176
rect 2040 -179 2070 -168
rect 2118 -172 2164 -156
rect 2191 -168 2265 -152
rect 2118 -174 2152 -172
rect 2117 -190 2164 -174
rect 2191 -190 2204 -168
rect 2219 -190 2249 -168
rect 2276 -190 2277 -174
rect 2292 -190 2305 -30
rect 2335 -134 2348 -30
rect 2393 -52 2394 -42
rect 2409 -52 2422 -42
rect 2393 -56 2422 -52
rect 2427 -56 2457 -30
rect 2475 -44 2491 -42
rect 2563 -44 2616 -30
rect 2564 -46 2628 -44
rect 2671 -46 2686 -30
rect 2735 -33 2765 -30
rect 2735 -36 2771 -33
rect 2701 -44 2717 -42
rect 2475 -56 2490 -52
rect 2393 -58 2490 -56
rect 2518 -58 2686 -46
rect 2702 -56 2717 -52
rect 2735 -55 2774 -36
rect 2793 -42 2800 -41
rect 2799 -49 2800 -42
rect 2783 -52 2784 -49
rect 2799 -52 2812 -49
rect 2735 -56 2765 -55
rect 2774 -56 2780 -55
rect 2783 -56 2812 -52
rect 2702 -57 2812 -56
rect 2702 -58 2818 -57
rect 2377 -66 2428 -58
rect 2377 -78 2402 -66
rect 2409 -78 2428 -66
rect 2459 -66 2509 -58
rect 2459 -74 2475 -66
rect 2482 -68 2509 -66
rect 2518 -68 2739 -58
rect 2482 -78 2739 -68
rect 2768 -66 2818 -58
rect 2768 -75 2784 -66
rect 2377 -86 2428 -78
rect 2475 -86 2739 -78
rect 2765 -78 2784 -75
rect 2791 -78 2818 -66
rect 2765 -86 2818 -78
rect 2393 -94 2394 -86
rect 2409 -94 2422 -86
rect 2393 -102 2409 -94
rect 2390 -109 2409 -106
rect 2390 -118 2412 -109
rect 2363 -128 2412 -118
rect 2363 -134 2393 -128
rect 2412 -133 2417 -128
rect 2335 -150 2409 -134
rect 2427 -142 2457 -86
rect 2492 -96 2700 -86
rect 2735 -90 2780 -86
rect 2783 -87 2784 -86
rect 2799 -87 2812 -86
rect 2518 -126 2707 -96
rect 2533 -129 2707 -126
rect 2526 -132 2707 -129
rect 2335 -152 2348 -150
rect 2363 -152 2397 -150
rect 2335 -168 2409 -152
rect 2436 -156 2449 -142
rect 2464 -156 2480 -140
rect 2526 -145 2537 -132
rect 2319 -190 2320 -174
rect 2335 -190 2348 -168
rect 2363 -190 2393 -168
rect 2436 -172 2498 -156
rect 2526 -163 2537 -147
rect 2542 -152 2552 -132
rect 2562 -152 2576 -132
rect 2579 -145 2588 -132
rect 2604 -145 2613 -132
rect 2542 -163 2576 -152
rect 2579 -163 2588 -147
rect 2604 -163 2613 -147
rect 2620 -152 2630 -132
rect 2640 -152 2654 -132
rect 2655 -145 2666 -132
rect 2620 -163 2654 -152
rect 2655 -163 2666 -147
rect 2712 -156 2728 -140
rect 2735 -142 2765 -90
rect 2799 -94 2800 -87
rect 2784 -102 2800 -94
rect 2771 -134 2784 -115
rect 2799 -134 2829 -118
rect 2771 -150 2845 -134
rect 2771 -152 2784 -150
rect 2799 -152 2833 -150
rect 2436 -174 2449 -172
rect 2464 -174 2498 -172
rect 2436 -190 2498 -174
rect 2542 -179 2558 -176
rect 2620 -179 2650 -168
rect 2698 -172 2744 -156
rect 2771 -168 2845 -152
rect 2698 -174 2732 -172
rect 2697 -190 2744 -174
rect 2771 -190 2784 -168
rect 2799 -190 2829 -168
rect 2856 -190 2857 -174
rect 2872 -190 2885 -30
rect 2915 -134 2928 -30
rect 2973 -52 2974 -42
rect 2989 -52 3002 -42
rect 2973 -56 3002 -52
rect 3007 -56 3037 -30
rect 3055 -44 3071 -42
rect 3143 -44 3196 -30
rect 3144 -46 3208 -44
rect 3251 -46 3266 -30
rect 3315 -33 3345 -30
rect 3315 -36 3351 -33
rect 3281 -44 3297 -42
rect 3055 -56 3070 -52
rect 2973 -58 3070 -56
rect 3098 -58 3266 -46
rect 3282 -56 3297 -52
rect 3315 -55 3354 -36
rect 3373 -42 3380 -41
rect 3379 -49 3380 -42
rect 3363 -52 3364 -49
rect 3379 -52 3392 -49
rect 3315 -56 3345 -55
rect 3354 -56 3360 -55
rect 3363 -56 3392 -52
rect 3282 -57 3392 -56
rect 3282 -58 3398 -57
rect 2957 -66 3008 -58
rect 2957 -78 2982 -66
rect 2989 -78 3008 -66
rect 3039 -66 3089 -58
rect 3039 -74 3055 -66
rect 3062 -68 3089 -66
rect 3098 -68 3319 -58
rect 3062 -78 3319 -68
rect 3348 -66 3398 -58
rect 3348 -75 3364 -66
rect 2957 -86 3008 -78
rect 3055 -86 3319 -78
rect 3345 -78 3364 -75
rect 3371 -78 3398 -66
rect 3345 -86 3398 -78
rect 2973 -94 2974 -86
rect 2989 -94 3002 -86
rect 2973 -102 2989 -94
rect 2970 -109 2989 -106
rect 2970 -118 2992 -109
rect 2943 -128 2992 -118
rect 2943 -134 2973 -128
rect 2992 -133 2997 -128
rect 2915 -150 2989 -134
rect 3007 -142 3037 -86
rect 3072 -96 3280 -86
rect 3315 -90 3360 -86
rect 3363 -87 3364 -86
rect 3379 -87 3392 -86
rect 3098 -126 3287 -96
rect 3113 -129 3287 -126
rect 3106 -132 3287 -129
rect 2915 -152 2928 -150
rect 2943 -152 2977 -150
rect 2915 -168 2989 -152
rect 3016 -156 3029 -142
rect 3044 -156 3060 -140
rect 3106 -145 3117 -132
rect 2899 -190 2900 -174
rect 2915 -190 2928 -168
rect 2943 -190 2973 -168
rect 3016 -172 3078 -156
rect 3106 -163 3117 -147
rect 3122 -152 3132 -132
rect 3142 -152 3156 -132
rect 3159 -145 3168 -132
rect 3184 -145 3193 -132
rect 3122 -163 3156 -152
rect 3159 -163 3168 -147
rect 3184 -163 3193 -147
rect 3200 -152 3210 -132
rect 3220 -152 3234 -132
rect 3235 -145 3246 -132
rect 3200 -163 3234 -152
rect 3235 -163 3246 -147
rect 3292 -156 3308 -140
rect 3315 -142 3345 -90
rect 3379 -94 3380 -87
rect 3364 -102 3380 -94
rect 3351 -134 3364 -115
rect 3379 -134 3409 -118
rect 3351 -150 3425 -134
rect 3351 -152 3364 -150
rect 3379 -152 3413 -150
rect 3016 -174 3029 -172
rect 3044 -174 3078 -172
rect 3016 -190 3078 -174
rect 3122 -179 3138 -176
rect 3200 -179 3230 -168
rect 3278 -172 3324 -156
rect 3351 -168 3425 -152
rect 3278 -174 3312 -172
rect 3277 -190 3324 -174
rect 3351 -190 3364 -168
rect 3379 -190 3409 -168
rect 3436 -190 3437 -174
rect 3452 -190 3465 -30
rect 3495 -134 3508 -30
rect 3553 -52 3554 -42
rect 3569 -52 3582 -42
rect 3553 -56 3582 -52
rect 3587 -56 3617 -30
rect 3635 -44 3651 -42
rect 3723 -44 3776 -30
rect 3724 -46 3788 -44
rect 3831 -46 3846 -30
rect 3895 -33 3925 -30
rect 3895 -36 3931 -33
rect 3861 -44 3877 -42
rect 3635 -56 3650 -52
rect 3553 -58 3650 -56
rect 3678 -58 3846 -46
rect 3862 -56 3877 -52
rect 3895 -55 3934 -36
rect 3953 -42 3960 -41
rect 3959 -49 3960 -42
rect 3943 -52 3944 -49
rect 3959 -52 3972 -49
rect 3895 -56 3925 -55
rect 3934 -56 3940 -55
rect 3943 -56 3972 -52
rect 3862 -57 3972 -56
rect 3862 -58 3978 -57
rect 3537 -66 3588 -58
rect 3537 -78 3562 -66
rect 3569 -78 3588 -66
rect 3619 -66 3669 -58
rect 3619 -74 3635 -66
rect 3642 -68 3669 -66
rect 3678 -68 3899 -58
rect 3642 -78 3899 -68
rect 3928 -66 3978 -58
rect 3928 -75 3944 -66
rect 3537 -86 3588 -78
rect 3635 -86 3899 -78
rect 3925 -78 3944 -75
rect 3951 -78 3978 -66
rect 3925 -86 3978 -78
rect 3553 -94 3554 -86
rect 3569 -94 3582 -86
rect 3553 -102 3569 -94
rect 3550 -109 3569 -106
rect 3550 -118 3572 -109
rect 3523 -128 3572 -118
rect 3523 -134 3553 -128
rect 3572 -133 3577 -128
rect 3495 -150 3569 -134
rect 3587 -142 3617 -86
rect 3652 -96 3860 -86
rect 3895 -90 3940 -86
rect 3943 -87 3944 -86
rect 3959 -87 3972 -86
rect 3678 -126 3867 -96
rect 3693 -129 3867 -126
rect 3686 -132 3867 -129
rect 3495 -152 3508 -150
rect 3523 -152 3557 -150
rect 3495 -168 3569 -152
rect 3596 -156 3609 -142
rect 3624 -156 3640 -140
rect 3686 -145 3697 -132
rect 3479 -190 3480 -174
rect 3495 -190 3508 -168
rect 3523 -190 3553 -168
rect 3596 -172 3658 -156
rect 3686 -163 3697 -147
rect 3702 -152 3712 -132
rect 3722 -152 3736 -132
rect 3739 -145 3748 -132
rect 3764 -145 3773 -132
rect 3702 -163 3736 -152
rect 3739 -163 3748 -147
rect 3764 -163 3773 -147
rect 3780 -152 3790 -132
rect 3800 -152 3814 -132
rect 3815 -145 3826 -132
rect 3780 -163 3814 -152
rect 3815 -163 3826 -147
rect 3872 -156 3888 -140
rect 3895 -142 3925 -90
rect 3959 -94 3960 -87
rect 3944 -102 3960 -94
rect 3931 -134 3944 -115
rect 3959 -134 3989 -118
rect 3931 -150 4005 -134
rect 3931 -152 3944 -150
rect 3959 -152 3993 -150
rect 3596 -174 3609 -172
rect 3624 -174 3658 -172
rect 3596 -190 3658 -174
rect 3702 -179 3718 -176
rect 3780 -179 3810 -168
rect 3858 -172 3904 -156
rect 3931 -168 4005 -152
rect 3858 -174 3892 -172
rect 3857 -190 3904 -174
rect 3931 -190 3944 -168
rect 3959 -190 3989 -168
rect 4016 -190 4017 -174
rect 4032 -190 4045 -30
rect 4075 -134 4088 -30
rect 4133 -52 4134 -42
rect 4149 -52 4162 -42
rect 4133 -56 4162 -52
rect 4167 -56 4197 -30
rect 4215 -44 4231 -42
rect 4303 -44 4356 -30
rect 4304 -46 4368 -44
rect 4411 -46 4426 -30
rect 4475 -33 4505 -30
rect 4475 -36 4511 -33
rect 4441 -44 4457 -42
rect 4215 -56 4230 -52
rect 4133 -58 4230 -56
rect 4258 -58 4426 -46
rect 4442 -56 4457 -52
rect 4475 -55 4514 -36
rect 4533 -42 4540 -41
rect 4539 -49 4540 -42
rect 4523 -52 4524 -49
rect 4539 -52 4552 -49
rect 4475 -56 4505 -55
rect 4514 -56 4520 -55
rect 4523 -56 4552 -52
rect 4442 -57 4552 -56
rect 4442 -58 4558 -57
rect 4117 -66 4168 -58
rect 4117 -78 4142 -66
rect 4149 -78 4168 -66
rect 4199 -66 4249 -58
rect 4199 -74 4215 -66
rect 4222 -68 4249 -66
rect 4258 -68 4479 -58
rect 4222 -78 4479 -68
rect 4508 -66 4558 -58
rect 4508 -75 4524 -66
rect 4117 -86 4168 -78
rect 4215 -86 4479 -78
rect 4505 -78 4524 -75
rect 4531 -78 4558 -66
rect 4505 -86 4558 -78
rect 4133 -94 4134 -86
rect 4149 -94 4162 -86
rect 4133 -102 4149 -94
rect 4130 -109 4149 -106
rect 4130 -118 4152 -109
rect 4103 -128 4152 -118
rect 4103 -134 4133 -128
rect 4152 -133 4157 -128
rect 4075 -150 4149 -134
rect 4167 -142 4197 -86
rect 4232 -96 4440 -86
rect 4475 -90 4520 -86
rect 4523 -87 4524 -86
rect 4539 -87 4552 -86
rect 4258 -126 4447 -96
rect 4273 -129 4447 -126
rect 4266 -132 4447 -129
rect 4075 -152 4088 -150
rect 4103 -152 4137 -150
rect 4075 -168 4149 -152
rect 4176 -156 4189 -142
rect 4204 -156 4220 -140
rect 4266 -145 4277 -132
rect 4059 -190 4060 -174
rect 4075 -190 4088 -168
rect 4103 -190 4133 -168
rect 4176 -172 4238 -156
rect 4266 -163 4277 -147
rect 4282 -152 4292 -132
rect 4302 -152 4316 -132
rect 4319 -145 4328 -132
rect 4344 -145 4353 -132
rect 4282 -163 4316 -152
rect 4319 -163 4328 -147
rect 4344 -163 4353 -147
rect 4360 -152 4370 -132
rect 4380 -152 4394 -132
rect 4395 -145 4406 -132
rect 4360 -163 4394 -152
rect 4395 -163 4406 -147
rect 4452 -156 4468 -140
rect 4475 -142 4505 -90
rect 4539 -94 4540 -87
rect 4524 -102 4540 -94
rect 4511 -134 4524 -115
rect 4539 -134 4569 -118
rect 4511 -150 4585 -134
rect 4511 -152 4524 -150
rect 4539 -152 4573 -150
rect 4176 -174 4189 -172
rect 4204 -174 4238 -172
rect 4176 -190 4238 -174
rect 4282 -179 4298 -176
rect 4360 -179 4390 -168
rect 4438 -172 4484 -156
rect 4511 -168 4585 -152
rect 4438 -174 4472 -172
rect 4437 -190 4484 -174
rect 4511 -190 4524 -168
rect 4539 -190 4569 -168
rect 4596 -190 4597 -174
rect 4612 -190 4625 -30
rect -7 -198 34 -190
rect -7 -224 8 -198
rect 15 -224 34 -198
rect 98 -202 160 -190
rect 172 -202 247 -190
rect 305 -202 380 -190
rect 392 -202 423 -190
rect 429 -202 464 -190
rect 98 -204 260 -202
rect -7 -232 34 -224
rect 116 -228 129 -204
rect 144 -206 159 -204
rect -1 -242 0 -232
rect 15 -242 28 -232
rect 43 -242 73 -228
rect 116 -242 159 -228
rect 183 -231 190 -224
rect 193 -228 260 -204
rect 292 -204 464 -202
rect 262 -226 290 -222
rect 292 -226 372 -204
rect 393 -206 408 -204
rect 262 -228 372 -226
rect 193 -232 372 -228
rect 166 -242 196 -232
rect 198 -242 351 -232
rect 359 -242 389 -232
rect 393 -242 423 -228
rect 451 -242 464 -204
rect 536 -198 571 -190
rect 536 -224 537 -198
rect 544 -224 571 -198
rect 479 -242 509 -228
rect 536 -232 571 -224
rect 573 -198 614 -190
rect 573 -224 588 -198
rect 595 -224 614 -198
rect 678 -202 740 -190
rect 752 -202 827 -190
rect 885 -202 960 -190
rect 972 -202 1003 -190
rect 1009 -202 1044 -190
rect 678 -204 840 -202
rect 573 -232 614 -224
rect 696 -228 709 -204
rect 724 -206 739 -204
rect 536 -242 537 -232
rect 552 -242 565 -232
rect 579 -242 580 -232
rect 595 -242 608 -232
rect 623 -242 653 -228
rect 696 -242 739 -228
rect 763 -231 770 -224
rect 773 -228 840 -204
rect 872 -204 1044 -202
rect 842 -226 870 -222
rect 872 -226 952 -204
rect 973 -206 988 -204
rect 842 -228 952 -226
rect 773 -232 952 -228
rect 746 -242 776 -232
rect 778 -242 931 -232
rect 939 -242 969 -232
rect 973 -242 1003 -228
rect 1031 -242 1044 -204
rect 1116 -198 1151 -190
rect 1116 -224 1117 -198
rect 1124 -224 1151 -198
rect 1059 -242 1089 -228
rect 1116 -232 1151 -224
rect 1153 -198 1194 -190
rect 1153 -224 1168 -198
rect 1175 -224 1194 -198
rect 1258 -202 1320 -190
rect 1332 -202 1407 -190
rect 1465 -202 1540 -190
rect 1552 -202 1583 -190
rect 1589 -202 1624 -190
rect 1258 -204 1420 -202
rect 1153 -232 1194 -224
rect 1276 -228 1289 -204
rect 1304 -206 1319 -204
rect 1116 -242 1117 -232
rect 1132 -242 1145 -232
rect 1159 -242 1160 -232
rect 1175 -242 1188 -232
rect 1203 -242 1233 -228
rect 1276 -242 1319 -228
rect 1343 -231 1350 -224
rect 1353 -228 1420 -204
rect 1452 -204 1624 -202
rect 1422 -226 1450 -222
rect 1452 -226 1532 -204
rect 1553 -206 1568 -204
rect 1422 -228 1532 -226
rect 1353 -232 1532 -228
rect 1326 -242 1356 -232
rect 1358 -242 1511 -232
rect 1519 -242 1549 -232
rect 1553 -242 1583 -228
rect 1611 -242 1624 -204
rect 1696 -198 1731 -190
rect 1696 -224 1697 -198
rect 1704 -224 1731 -198
rect 1639 -242 1669 -228
rect 1696 -232 1731 -224
rect 1733 -198 1774 -190
rect 1733 -224 1748 -198
rect 1755 -224 1774 -198
rect 1838 -202 1900 -190
rect 1912 -202 1987 -190
rect 2045 -202 2120 -190
rect 2132 -202 2163 -190
rect 2169 -202 2204 -190
rect 1838 -204 2000 -202
rect 1733 -232 1774 -224
rect 1856 -228 1869 -204
rect 1884 -206 1899 -204
rect 1696 -242 1697 -232
rect 1712 -242 1725 -232
rect 1739 -242 1740 -232
rect 1755 -242 1768 -232
rect 1783 -242 1813 -228
rect 1856 -242 1899 -228
rect 1923 -231 1930 -224
rect 1933 -228 2000 -204
rect 2032 -204 2204 -202
rect 2002 -226 2030 -222
rect 2032 -226 2112 -204
rect 2133 -206 2148 -204
rect 2002 -228 2112 -226
rect 1933 -232 2112 -228
rect 1906 -242 1936 -232
rect 1938 -242 2091 -232
rect 2099 -242 2129 -232
rect 2133 -242 2163 -228
rect 2191 -242 2204 -204
rect 2276 -198 2311 -190
rect 2276 -224 2277 -198
rect 2284 -224 2311 -198
rect 2219 -242 2249 -228
rect 2276 -232 2311 -224
rect 2313 -198 2354 -190
rect 2313 -224 2328 -198
rect 2335 -224 2354 -198
rect 2418 -202 2480 -190
rect 2492 -202 2567 -190
rect 2625 -202 2700 -190
rect 2712 -202 2743 -190
rect 2749 -202 2784 -190
rect 2418 -204 2580 -202
rect 2313 -232 2354 -224
rect 2436 -228 2449 -204
rect 2464 -206 2479 -204
rect 2276 -242 2277 -232
rect 2292 -242 2305 -232
rect 2319 -242 2320 -232
rect 2335 -242 2348 -232
rect 2363 -242 2393 -228
rect 2436 -242 2479 -228
rect 2503 -231 2510 -224
rect 2513 -228 2580 -204
rect 2612 -204 2784 -202
rect 2582 -226 2610 -222
rect 2612 -226 2692 -204
rect 2713 -206 2728 -204
rect 2582 -228 2692 -226
rect 2513 -232 2692 -228
rect 2486 -242 2516 -232
rect 2518 -242 2671 -232
rect 2679 -242 2709 -232
rect 2713 -242 2743 -228
rect 2771 -242 2784 -204
rect 2856 -198 2891 -190
rect 2856 -224 2857 -198
rect 2864 -224 2891 -198
rect 2799 -242 2829 -228
rect 2856 -232 2891 -224
rect 2893 -198 2934 -190
rect 2893 -224 2908 -198
rect 2915 -224 2934 -198
rect 2998 -202 3060 -190
rect 3072 -202 3147 -190
rect 3205 -202 3280 -190
rect 3292 -202 3323 -190
rect 3329 -202 3364 -190
rect 2998 -204 3160 -202
rect 2893 -232 2934 -224
rect 3016 -228 3029 -204
rect 3044 -206 3059 -204
rect 2856 -242 2857 -232
rect 2872 -242 2885 -232
rect 2899 -242 2900 -232
rect 2915 -242 2928 -232
rect 2943 -242 2973 -228
rect 3016 -242 3059 -228
rect 3083 -231 3090 -224
rect 3093 -228 3160 -204
rect 3192 -204 3364 -202
rect 3162 -226 3190 -222
rect 3192 -226 3272 -204
rect 3293 -206 3308 -204
rect 3162 -228 3272 -226
rect 3093 -232 3272 -228
rect 3066 -242 3096 -232
rect 3098 -242 3251 -232
rect 3259 -242 3289 -232
rect 3293 -242 3323 -228
rect 3351 -242 3364 -204
rect 3436 -198 3471 -190
rect 3436 -224 3437 -198
rect 3444 -224 3471 -198
rect 3379 -242 3409 -228
rect 3436 -232 3471 -224
rect 3473 -198 3514 -190
rect 3473 -224 3488 -198
rect 3495 -224 3514 -198
rect 3578 -202 3640 -190
rect 3652 -202 3727 -190
rect 3785 -202 3860 -190
rect 3872 -202 3903 -190
rect 3909 -202 3944 -190
rect 3578 -204 3740 -202
rect 3473 -232 3514 -224
rect 3596 -228 3609 -204
rect 3624 -206 3639 -204
rect 3436 -242 3437 -232
rect 3452 -242 3465 -232
rect 3479 -242 3480 -232
rect 3495 -242 3508 -232
rect 3523 -242 3553 -228
rect 3596 -242 3639 -228
rect 3663 -231 3670 -224
rect 3673 -228 3740 -204
rect 3772 -204 3944 -202
rect 3742 -226 3770 -222
rect 3772 -226 3852 -204
rect 3873 -206 3888 -204
rect 3742 -228 3852 -226
rect 3673 -232 3852 -228
rect 3646 -242 3676 -232
rect 3678 -242 3831 -232
rect 3839 -242 3869 -232
rect 3873 -242 3903 -228
rect 3931 -242 3944 -204
rect 4016 -198 4051 -190
rect 4016 -224 4017 -198
rect 4024 -224 4051 -198
rect 3959 -242 3989 -228
rect 4016 -232 4051 -224
rect 4053 -198 4094 -190
rect 4053 -224 4068 -198
rect 4075 -224 4094 -198
rect 4158 -202 4220 -190
rect 4232 -202 4307 -190
rect 4365 -202 4440 -190
rect 4452 -202 4483 -190
rect 4489 -202 4524 -190
rect 4158 -204 4320 -202
rect 4053 -232 4094 -224
rect 4176 -228 4189 -204
rect 4204 -206 4219 -204
rect 4016 -242 4017 -232
rect 4032 -242 4045 -232
rect 4059 -242 4060 -232
rect 4075 -242 4088 -232
rect 4103 -242 4133 -228
rect 4176 -242 4219 -228
rect 4243 -231 4250 -224
rect 4253 -228 4320 -204
rect 4352 -204 4524 -202
rect 4322 -226 4350 -222
rect 4352 -226 4432 -204
rect 4453 -206 4468 -204
rect 4322 -228 4432 -226
rect 4253 -232 4432 -228
rect 4226 -242 4256 -232
rect 4258 -242 4411 -232
rect 4419 -242 4449 -232
rect 4453 -242 4483 -228
rect 4511 -242 4524 -204
rect 4596 -198 4631 -190
rect 4596 -224 4597 -198
rect 4604 -224 4631 -198
rect 4539 -242 4569 -228
rect 4596 -232 4631 -224
rect 4596 -242 4597 -232
rect 4612 -242 4625 -232
rect -1 -248 4625 -242
rect 0 -256 4625 -248
rect 15 -286 28 -256
rect 43 -274 73 -256
rect 116 -270 130 -256
rect 166 -270 386 -256
rect 117 -272 130 -270
rect 83 -284 98 -272
rect 80 -286 102 -284
rect 107 -286 137 -272
rect 198 -274 351 -270
rect 180 -286 372 -274
rect 415 -286 445 -272
rect 451 -286 464 -256
rect 479 -274 509 -256
rect 552 -286 565 -256
rect 595 -286 608 -256
rect 623 -274 653 -256
rect 696 -270 710 -256
rect 746 -270 966 -256
rect 697 -272 710 -270
rect 663 -284 678 -272
rect 660 -286 682 -284
rect 687 -286 717 -272
rect 778 -274 931 -270
rect 760 -286 952 -274
rect 995 -286 1025 -272
rect 1031 -286 1044 -256
rect 1059 -274 1089 -256
rect 1132 -286 1145 -256
rect 1175 -286 1188 -256
rect 1203 -274 1233 -256
rect 1276 -270 1290 -256
rect 1326 -270 1546 -256
rect 1277 -272 1290 -270
rect 1243 -284 1258 -272
rect 1240 -286 1262 -284
rect 1267 -286 1297 -272
rect 1358 -274 1511 -270
rect 1340 -286 1532 -274
rect 1575 -286 1605 -272
rect 1611 -286 1624 -256
rect 1639 -274 1669 -256
rect 1712 -286 1725 -256
rect 1755 -286 1768 -256
rect 1783 -274 1813 -256
rect 1856 -270 1870 -256
rect 1906 -270 2126 -256
rect 1857 -272 1870 -270
rect 1823 -284 1838 -272
rect 1820 -286 1842 -284
rect 1847 -286 1877 -272
rect 1938 -274 2091 -270
rect 1920 -286 2112 -274
rect 2155 -286 2185 -272
rect 2191 -286 2204 -256
rect 2219 -274 2249 -256
rect 2292 -286 2305 -256
rect 2335 -286 2348 -256
rect 2363 -274 2393 -256
rect 2436 -270 2450 -256
rect 2486 -270 2706 -256
rect 2437 -272 2450 -270
rect 2403 -284 2418 -272
rect 2400 -286 2422 -284
rect 2427 -286 2457 -272
rect 2518 -274 2671 -270
rect 2500 -286 2692 -274
rect 2735 -286 2765 -272
rect 2771 -286 2784 -256
rect 2799 -274 2829 -256
rect 2872 -286 2885 -256
rect 2915 -286 2928 -256
rect 2943 -274 2973 -256
rect 3016 -270 3030 -256
rect 3066 -270 3286 -256
rect 3017 -272 3030 -270
rect 2983 -284 2998 -272
rect 2980 -286 3002 -284
rect 3007 -286 3037 -272
rect 3098 -274 3251 -270
rect 3080 -286 3272 -274
rect 3315 -286 3345 -272
rect 3351 -286 3364 -256
rect 3379 -274 3409 -256
rect 3452 -286 3465 -256
rect 3495 -286 3508 -256
rect 3523 -274 3553 -256
rect 3596 -270 3610 -256
rect 3646 -270 3866 -256
rect 3597 -272 3610 -270
rect 3563 -284 3578 -272
rect 3560 -286 3582 -284
rect 3587 -286 3617 -272
rect 3678 -274 3831 -270
rect 3660 -286 3852 -274
rect 3895 -286 3925 -272
rect 3931 -286 3944 -256
rect 3959 -274 3989 -256
rect 4032 -286 4045 -256
rect 4075 -286 4088 -256
rect 4103 -274 4133 -256
rect 4176 -270 4190 -256
rect 4226 -270 4446 -256
rect 4177 -272 4190 -270
rect 4143 -284 4158 -272
rect 4140 -286 4162 -284
rect 4167 -286 4197 -272
rect 4258 -274 4411 -270
rect 4240 -286 4432 -274
rect 4475 -286 4505 -272
rect 4511 -286 4524 -256
rect 4539 -274 4569 -256
rect 4612 -286 4625 -256
rect 0 -300 4625 -286
rect 15 -404 28 -300
rect 73 -322 74 -312
rect 89 -322 102 -312
rect 73 -326 102 -322
rect 107 -326 137 -300
rect 155 -314 171 -312
rect 243 -314 296 -300
rect 244 -316 308 -314
rect 351 -316 366 -300
rect 415 -303 445 -300
rect 415 -306 451 -303
rect 381 -314 397 -312
rect 155 -326 170 -322
rect 73 -328 170 -326
rect 198 -328 366 -316
rect 382 -326 397 -322
rect 415 -325 454 -306
rect 473 -312 480 -311
rect 479 -319 480 -312
rect 463 -322 464 -319
rect 479 -322 492 -319
rect 415 -326 445 -325
rect 454 -326 460 -325
rect 463 -326 492 -322
rect 382 -327 492 -326
rect 382 -328 498 -327
rect 57 -336 108 -328
rect 57 -348 82 -336
rect 89 -348 108 -336
rect 139 -336 189 -328
rect 139 -344 155 -336
rect 162 -338 189 -336
rect 198 -338 419 -328
rect 162 -348 419 -338
rect 448 -336 498 -328
rect 448 -345 464 -336
rect 57 -356 108 -348
rect 155 -356 419 -348
rect 445 -348 464 -345
rect 471 -348 498 -336
rect 445 -356 498 -348
rect 73 -364 74 -356
rect 89 -364 102 -356
rect 73 -372 89 -364
rect 70 -379 89 -376
rect 70 -388 92 -379
rect 43 -398 92 -388
rect 43 -404 73 -398
rect 92 -403 97 -398
rect 15 -420 89 -404
rect 107 -412 137 -356
rect 172 -366 380 -356
rect 415 -360 460 -356
rect 463 -357 464 -356
rect 479 -357 492 -356
rect 198 -396 387 -366
rect 213 -399 387 -396
rect 206 -402 387 -399
rect 15 -422 28 -420
rect 43 -422 77 -420
rect 15 -438 89 -422
rect 116 -426 129 -412
rect 144 -426 160 -410
rect 206 -415 217 -402
rect -1 -460 0 -444
rect 15 -460 28 -438
rect 43 -460 73 -438
rect 116 -442 178 -426
rect 206 -433 217 -417
rect 222 -422 232 -402
rect 242 -422 256 -402
rect 259 -415 268 -402
rect 284 -415 293 -402
rect 222 -433 256 -422
rect 259 -433 268 -417
rect 284 -433 293 -417
rect 300 -422 310 -402
rect 320 -422 334 -402
rect 335 -415 346 -402
rect 300 -433 334 -422
rect 335 -433 346 -417
rect 392 -426 408 -410
rect 415 -412 445 -360
rect 479 -364 480 -357
rect 464 -372 480 -364
rect 451 -404 464 -385
rect 479 -404 509 -388
rect 451 -420 525 -404
rect 451 -422 464 -420
rect 479 -422 513 -420
rect 116 -444 129 -442
rect 144 -444 178 -442
rect 116 -460 178 -444
rect 222 -449 238 -446
rect 300 -449 330 -438
rect 378 -442 424 -426
rect 451 -438 525 -422
rect 378 -444 412 -442
rect 377 -460 424 -444
rect 451 -460 464 -438
rect 479 -460 509 -438
rect 536 -460 537 -444
rect 552 -460 565 -300
rect 595 -404 608 -300
rect 653 -322 654 -312
rect 669 -322 682 -312
rect 653 -326 682 -322
rect 687 -326 717 -300
rect 735 -314 751 -312
rect 823 -314 876 -300
rect 824 -316 888 -314
rect 931 -316 946 -300
rect 995 -303 1025 -300
rect 995 -306 1031 -303
rect 961 -314 977 -312
rect 735 -326 750 -322
rect 653 -328 750 -326
rect 778 -328 946 -316
rect 962 -326 977 -322
rect 995 -325 1034 -306
rect 1053 -312 1060 -311
rect 1059 -319 1060 -312
rect 1043 -322 1044 -319
rect 1059 -322 1072 -319
rect 995 -326 1025 -325
rect 1034 -326 1040 -325
rect 1043 -326 1072 -322
rect 962 -327 1072 -326
rect 962 -328 1078 -327
rect 637 -336 688 -328
rect 637 -348 662 -336
rect 669 -348 688 -336
rect 719 -336 769 -328
rect 719 -344 735 -336
rect 742 -338 769 -336
rect 778 -338 999 -328
rect 742 -348 999 -338
rect 1028 -336 1078 -328
rect 1028 -345 1044 -336
rect 637 -356 688 -348
rect 735 -356 999 -348
rect 1025 -348 1044 -345
rect 1051 -348 1078 -336
rect 1025 -356 1078 -348
rect 653 -364 654 -356
rect 669 -364 682 -356
rect 653 -372 669 -364
rect 650 -379 669 -376
rect 650 -388 672 -379
rect 623 -398 672 -388
rect 623 -404 653 -398
rect 672 -403 677 -398
rect 595 -420 669 -404
rect 687 -412 717 -356
rect 752 -366 960 -356
rect 995 -360 1040 -356
rect 1043 -357 1044 -356
rect 1059 -357 1072 -356
rect 778 -396 967 -366
rect 793 -399 967 -396
rect 786 -402 967 -399
rect 595 -422 608 -420
rect 623 -422 657 -420
rect 595 -438 669 -422
rect 696 -426 709 -412
rect 724 -426 740 -410
rect 786 -415 797 -402
rect 579 -460 580 -444
rect 595 -460 608 -438
rect 623 -460 653 -438
rect 696 -442 758 -426
rect 786 -433 797 -417
rect 802 -422 812 -402
rect 822 -422 836 -402
rect 839 -415 848 -402
rect 864 -415 873 -402
rect 802 -433 836 -422
rect 839 -433 848 -417
rect 864 -433 873 -417
rect 880 -422 890 -402
rect 900 -422 914 -402
rect 915 -415 926 -402
rect 880 -433 914 -422
rect 915 -433 926 -417
rect 972 -426 988 -410
rect 995 -412 1025 -360
rect 1059 -364 1060 -357
rect 1044 -372 1060 -364
rect 1031 -404 1044 -385
rect 1059 -404 1089 -388
rect 1031 -420 1105 -404
rect 1031 -422 1044 -420
rect 1059 -422 1093 -420
rect 696 -444 709 -442
rect 724 -444 758 -442
rect 696 -460 758 -444
rect 802 -449 818 -446
rect 880 -449 910 -438
rect 958 -442 1004 -426
rect 1031 -438 1105 -422
rect 958 -444 992 -442
rect 957 -460 1004 -444
rect 1031 -460 1044 -438
rect 1059 -460 1089 -438
rect 1116 -460 1117 -444
rect 1132 -460 1145 -300
rect 1175 -404 1188 -300
rect 1233 -322 1234 -312
rect 1249 -322 1262 -312
rect 1233 -326 1262 -322
rect 1267 -326 1297 -300
rect 1315 -314 1331 -312
rect 1403 -314 1456 -300
rect 1404 -316 1468 -314
rect 1511 -316 1526 -300
rect 1575 -303 1605 -300
rect 1575 -306 1611 -303
rect 1541 -314 1557 -312
rect 1315 -326 1330 -322
rect 1233 -328 1330 -326
rect 1358 -328 1526 -316
rect 1542 -326 1557 -322
rect 1575 -325 1614 -306
rect 1633 -312 1640 -311
rect 1639 -319 1640 -312
rect 1623 -322 1624 -319
rect 1639 -322 1652 -319
rect 1575 -326 1605 -325
rect 1614 -326 1620 -325
rect 1623 -326 1652 -322
rect 1542 -327 1652 -326
rect 1542 -328 1658 -327
rect 1217 -336 1268 -328
rect 1217 -348 1242 -336
rect 1249 -348 1268 -336
rect 1299 -336 1349 -328
rect 1299 -344 1315 -336
rect 1322 -338 1349 -336
rect 1358 -338 1579 -328
rect 1322 -348 1579 -338
rect 1608 -336 1658 -328
rect 1608 -345 1624 -336
rect 1217 -356 1268 -348
rect 1315 -356 1579 -348
rect 1605 -348 1624 -345
rect 1631 -348 1658 -336
rect 1605 -356 1658 -348
rect 1233 -364 1234 -356
rect 1249 -364 1262 -356
rect 1233 -372 1249 -364
rect 1230 -379 1249 -376
rect 1230 -388 1252 -379
rect 1203 -398 1252 -388
rect 1203 -404 1233 -398
rect 1252 -403 1257 -398
rect 1175 -420 1249 -404
rect 1267 -412 1297 -356
rect 1332 -366 1540 -356
rect 1575 -360 1620 -356
rect 1623 -357 1624 -356
rect 1639 -357 1652 -356
rect 1358 -396 1547 -366
rect 1373 -399 1547 -396
rect 1366 -402 1547 -399
rect 1175 -422 1188 -420
rect 1203 -422 1237 -420
rect 1175 -438 1249 -422
rect 1276 -426 1289 -412
rect 1304 -426 1320 -410
rect 1366 -415 1377 -402
rect 1159 -460 1160 -444
rect 1175 -460 1188 -438
rect 1203 -460 1233 -438
rect 1276 -442 1338 -426
rect 1366 -433 1377 -417
rect 1382 -422 1392 -402
rect 1402 -422 1416 -402
rect 1419 -415 1428 -402
rect 1444 -415 1453 -402
rect 1382 -433 1416 -422
rect 1419 -433 1428 -417
rect 1444 -433 1453 -417
rect 1460 -422 1470 -402
rect 1480 -422 1494 -402
rect 1495 -415 1506 -402
rect 1460 -433 1494 -422
rect 1495 -433 1506 -417
rect 1552 -426 1568 -410
rect 1575 -412 1605 -360
rect 1639 -364 1640 -357
rect 1624 -372 1640 -364
rect 1611 -404 1624 -385
rect 1639 -404 1669 -388
rect 1611 -420 1685 -404
rect 1611 -422 1624 -420
rect 1639 -422 1673 -420
rect 1276 -444 1289 -442
rect 1304 -444 1338 -442
rect 1276 -460 1338 -444
rect 1382 -449 1398 -446
rect 1460 -449 1490 -438
rect 1538 -442 1584 -426
rect 1611 -438 1685 -422
rect 1538 -444 1572 -442
rect 1537 -460 1584 -444
rect 1611 -460 1624 -438
rect 1639 -460 1669 -438
rect 1696 -460 1697 -444
rect 1712 -460 1725 -300
rect 1755 -404 1768 -300
rect 1813 -322 1814 -312
rect 1829 -322 1842 -312
rect 1813 -326 1842 -322
rect 1847 -326 1877 -300
rect 1895 -314 1911 -312
rect 1983 -314 2036 -300
rect 1984 -316 2048 -314
rect 2091 -316 2106 -300
rect 2155 -303 2185 -300
rect 2155 -306 2191 -303
rect 2121 -314 2137 -312
rect 1895 -326 1910 -322
rect 1813 -328 1910 -326
rect 1938 -328 2106 -316
rect 2122 -326 2137 -322
rect 2155 -325 2194 -306
rect 2213 -312 2220 -311
rect 2219 -319 2220 -312
rect 2203 -322 2204 -319
rect 2219 -322 2232 -319
rect 2155 -326 2185 -325
rect 2194 -326 2200 -325
rect 2203 -326 2232 -322
rect 2122 -327 2232 -326
rect 2122 -328 2238 -327
rect 1797 -336 1848 -328
rect 1797 -348 1822 -336
rect 1829 -348 1848 -336
rect 1879 -336 1929 -328
rect 1879 -344 1895 -336
rect 1902 -338 1929 -336
rect 1938 -338 2159 -328
rect 1902 -348 2159 -338
rect 2188 -336 2238 -328
rect 2188 -345 2204 -336
rect 1797 -356 1848 -348
rect 1895 -356 2159 -348
rect 2185 -348 2204 -345
rect 2211 -348 2238 -336
rect 2185 -356 2238 -348
rect 1813 -364 1814 -356
rect 1829 -364 1842 -356
rect 1813 -372 1829 -364
rect 1810 -379 1829 -376
rect 1810 -388 1832 -379
rect 1783 -398 1832 -388
rect 1783 -404 1813 -398
rect 1832 -403 1837 -398
rect 1755 -420 1829 -404
rect 1847 -412 1877 -356
rect 1912 -366 2120 -356
rect 2155 -360 2200 -356
rect 2203 -357 2204 -356
rect 2219 -357 2232 -356
rect 1938 -396 2127 -366
rect 1953 -399 2127 -396
rect 1946 -402 2127 -399
rect 1755 -422 1768 -420
rect 1783 -422 1817 -420
rect 1755 -438 1829 -422
rect 1856 -426 1869 -412
rect 1884 -426 1900 -410
rect 1946 -415 1957 -402
rect 1739 -460 1740 -444
rect 1755 -460 1768 -438
rect 1783 -460 1813 -438
rect 1856 -442 1918 -426
rect 1946 -433 1957 -417
rect 1962 -422 1972 -402
rect 1982 -422 1996 -402
rect 1999 -415 2008 -402
rect 2024 -415 2033 -402
rect 1962 -433 1996 -422
rect 1999 -433 2008 -417
rect 2024 -433 2033 -417
rect 2040 -422 2050 -402
rect 2060 -422 2074 -402
rect 2075 -415 2086 -402
rect 2040 -433 2074 -422
rect 2075 -433 2086 -417
rect 2132 -426 2148 -410
rect 2155 -412 2185 -360
rect 2219 -364 2220 -357
rect 2204 -372 2220 -364
rect 2191 -404 2204 -385
rect 2219 -404 2249 -388
rect 2191 -420 2265 -404
rect 2191 -422 2204 -420
rect 2219 -422 2253 -420
rect 1856 -444 1869 -442
rect 1884 -444 1918 -442
rect 1856 -460 1918 -444
rect 1962 -449 1978 -446
rect 2040 -449 2070 -438
rect 2118 -442 2164 -426
rect 2191 -438 2265 -422
rect 2118 -444 2152 -442
rect 2117 -460 2164 -444
rect 2191 -460 2204 -438
rect 2219 -460 2249 -438
rect 2276 -460 2277 -444
rect 2292 -460 2305 -300
rect 2335 -404 2348 -300
rect 2393 -322 2394 -312
rect 2409 -322 2422 -312
rect 2393 -326 2422 -322
rect 2427 -326 2457 -300
rect 2475 -314 2491 -312
rect 2563 -314 2616 -300
rect 2564 -316 2628 -314
rect 2671 -316 2686 -300
rect 2735 -303 2765 -300
rect 2735 -306 2771 -303
rect 2701 -314 2717 -312
rect 2475 -326 2490 -322
rect 2393 -328 2490 -326
rect 2518 -328 2686 -316
rect 2702 -326 2717 -322
rect 2735 -325 2774 -306
rect 2793 -312 2800 -311
rect 2799 -319 2800 -312
rect 2783 -322 2784 -319
rect 2799 -322 2812 -319
rect 2735 -326 2765 -325
rect 2774 -326 2780 -325
rect 2783 -326 2812 -322
rect 2702 -327 2812 -326
rect 2702 -328 2818 -327
rect 2377 -336 2428 -328
rect 2377 -348 2402 -336
rect 2409 -348 2428 -336
rect 2459 -336 2509 -328
rect 2459 -344 2475 -336
rect 2482 -338 2509 -336
rect 2518 -338 2739 -328
rect 2482 -348 2739 -338
rect 2768 -336 2818 -328
rect 2768 -345 2784 -336
rect 2377 -356 2428 -348
rect 2475 -356 2739 -348
rect 2765 -348 2784 -345
rect 2791 -348 2818 -336
rect 2765 -356 2818 -348
rect 2393 -364 2394 -356
rect 2409 -364 2422 -356
rect 2393 -372 2409 -364
rect 2390 -379 2409 -376
rect 2390 -388 2412 -379
rect 2363 -398 2412 -388
rect 2363 -404 2393 -398
rect 2412 -403 2417 -398
rect 2335 -420 2409 -404
rect 2427 -412 2457 -356
rect 2492 -366 2700 -356
rect 2735 -360 2780 -356
rect 2783 -357 2784 -356
rect 2799 -357 2812 -356
rect 2518 -396 2707 -366
rect 2533 -399 2707 -396
rect 2526 -402 2707 -399
rect 2335 -422 2348 -420
rect 2363 -422 2397 -420
rect 2335 -438 2409 -422
rect 2436 -426 2449 -412
rect 2464 -426 2480 -410
rect 2526 -415 2537 -402
rect 2319 -460 2320 -444
rect 2335 -460 2348 -438
rect 2363 -460 2393 -438
rect 2436 -442 2498 -426
rect 2526 -433 2537 -417
rect 2542 -422 2552 -402
rect 2562 -422 2576 -402
rect 2579 -415 2588 -402
rect 2604 -415 2613 -402
rect 2542 -433 2576 -422
rect 2579 -433 2588 -417
rect 2604 -433 2613 -417
rect 2620 -422 2630 -402
rect 2640 -422 2654 -402
rect 2655 -415 2666 -402
rect 2620 -433 2654 -422
rect 2655 -433 2666 -417
rect 2712 -426 2728 -410
rect 2735 -412 2765 -360
rect 2799 -364 2800 -357
rect 2784 -372 2800 -364
rect 2771 -404 2784 -385
rect 2799 -404 2829 -388
rect 2771 -420 2845 -404
rect 2771 -422 2784 -420
rect 2799 -422 2833 -420
rect 2436 -444 2449 -442
rect 2464 -444 2498 -442
rect 2436 -460 2498 -444
rect 2542 -449 2558 -446
rect 2620 -449 2650 -438
rect 2698 -442 2744 -426
rect 2771 -438 2845 -422
rect 2698 -444 2732 -442
rect 2697 -460 2744 -444
rect 2771 -460 2784 -438
rect 2799 -460 2829 -438
rect 2856 -460 2857 -444
rect 2872 -460 2885 -300
rect 2915 -404 2928 -300
rect 2973 -322 2974 -312
rect 2989 -322 3002 -312
rect 2973 -326 3002 -322
rect 3007 -326 3037 -300
rect 3055 -314 3071 -312
rect 3143 -314 3196 -300
rect 3144 -316 3208 -314
rect 3251 -316 3266 -300
rect 3315 -303 3345 -300
rect 3315 -306 3351 -303
rect 3281 -314 3297 -312
rect 3055 -326 3070 -322
rect 2973 -328 3070 -326
rect 3098 -328 3266 -316
rect 3282 -326 3297 -322
rect 3315 -325 3354 -306
rect 3373 -312 3380 -311
rect 3379 -319 3380 -312
rect 3363 -322 3364 -319
rect 3379 -322 3392 -319
rect 3315 -326 3345 -325
rect 3354 -326 3360 -325
rect 3363 -326 3392 -322
rect 3282 -327 3392 -326
rect 3282 -328 3398 -327
rect 2957 -336 3008 -328
rect 2957 -348 2982 -336
rect 2989 -348 3008 -336
rect 3039 -336 3089 -328
rect 3039 -344 3055 -336
rect 3062 -338 3089 -336
rect 3098 -338 3319 -328
rect 3062 -348 3319 -338
rect 3348 -336 3398 -328
rect 3348 -345 3364 -336
rect 2957 -356 3008 -348
rect 3055 -356 3319 -348
rect 3345 -348 3364 -345
rect 3371 -348 3398 -336
rect 3345 -356 3398 -348
rect 2973 -364 2974 -356
rect 2989 -364 3002 -356
rect 2973 -372 2989 -364
rect 2970 -379 2989 -376
rect 2970 -388 2992 -379
rect 2943 -398 2992 -388
rect 2943 -404 2973 -398
rect 2992 -403 2997 -398
rect 2915 -420 2989 -404
rect 3007 -412 3037 -356
rect 3072 -366 3280 -356
rect 3315 -360 3360 -356
rect 3363 -357 3364 -356
rect 3379 -357 3392 -356
rect 3098 -396 3287 -366
rect 3113 -399 3287 -396
rect 3106 -402 3287 -399
rect 2915 -422 2928 -420
rect 2943 -422 2977 -420
rect 2915 -438 2989 -422
rect 3016 -426 3029 -412
rect 3044 -426 3060 -410
rect 3106 -415 3117 -402
rect 2899 -460 2900 -444
rect 2915 -460 2928 -438
rect 2943 -460 2973 -438
rect 3016 -442 3078 -426
rect 3106 -433 3117 -417
rect 3122 -422 3132 -402
rect 3142 -422 3156 -402
rect 3159 -415 3168 -402
rect 3184 -415 3193 -402
rect 3122 -433 3156 -422
rect 3159 -433 3168 -417
rect 3184 -433 3193 -417
rect 3200 -422 3210 -402
rect 3220 -422 3234 -402
rect 3235 -415 3246 -402
rect 3200 -433 3234 -422
rect 3235 -433 3246 -417
rect 3292 -426 3308 -410
rect 3315 -412 3345 -360
rect 3379 -364 3380 -357
rect 3364 -372 3380 -364
rect 3351 -404 3364 -385
rect 3379 -404 3409 -388
rect 3351 -420 3425 -404
rect 3351 -422 3364 -420
rect 3379 -422 3413 -420
rect 3016 -444 3029 -442
rect 3044 -444 3078 -442
rect 3016 -460 3078 -444
rect 3122 -449 3138 -446
rect 3200 -449 3230 -438
rect 3278 -442 3324 -426
rect 3351 -438 3425 -422
rect 3278 -444 3312 -442
rect 3277 -460 3324 -444
rect 3351 -460 3364 -438
rect 3379 -460 3409 -438
rect 3436 -460 3437 -444
rect 3452 -460 3465 -300
rect 3495 -404 3508 -300
rect 3553 -322 3554 -312
rect 3569 -322 3582 -312
rect 3553 -326 3582 -322
rect 3587 -326 3617 -300
rect 3635 -314 3651 -312
rect 3723 -314 3776 -300
rect 3724 -316 3788 -314
rect 3831 -316 3846 -300
rect 3895 -303 3925 -300
rect 3895 -306 3931 -303
rect 3861 -314 3877 -312
rect 3635 -326 3650 -322
rect 3553 -328 3650 -326
rect 3678 -328 3846 -316
rect 3862 -326 3877 -322
rect 3895 -325 3934 -306
rect 3953 -312 3960 -311
rect 3959 -319 3960 -312
rect 3943 -322 3944 -319
rect 3959 -322 3972 -319
rect 3895 -326 3925 -325
rect 3934 -326 3940 -325
rect 3943 -326 3972 -322
rect 3862 -327 3972 -326
rect 3862 -328 3978 -327
rect 3537 -336 3588 -328
rect 3537 -348 3562 -336
rect 3569 -348 3588 -336
rect 3619 -336 3669 -328
rect 3619 -344 3635 -336
rect 3642 -338 3669 -336
rect 3678 -338 3899 -328
rect 3642 -348 3899 -338
rect 3928 -336 3978 -328
rect 3928 -345 3944 -336
rect 3537 -356 3588 -348
rect 3635 -356 3899 -348
rect 3925 -348 3944 -345
rect 3951 -348 3978 -336
rect 3925 -356 3978 -348
rect 3553 -364 3554 -356
rect 3569 -364 3582 -356
rect 3553 -372 3569 -364
rect 3550 -379 3569 -376
rect 3550 -388 3572 -379
rect 3523 -398 3572 -388
rect 3523 -404 3553 -398
rect 3572 -403 3577 -398
rect 3495 -420 3569 -404
rect 3587 -412 3617 -356
rect 3652 -366 3860 -356
rect 3895 -360 3940 -356
rect 3943 -357 3944 -356
rect 3959 -357 3972 -356
rect 3678 -396 3867 -366
rect 3693 -399 3867 -396
rect 3686 -402 3867 -399
rect 3495 -422 3508 -420
rect 3523 -422 3557 -420
rect 3495 -438 3569 -422
rect 3596 -426 3609 -412
rect 3624 -426 3640 -410
rect 3686 -415 3697 -402
rect 3479 -460 3480 -444
rect 3495 -460 3508 -438
rect 3523 -460 3553 -438
rect 3596 -442 3658 -426
rect 3686 -433 3697 -417
rect 3702 -422 3712 -402
rect 3722 -422 3736 -402
rect 3739 -415 3748 -402
rect 3764 -415 3773 -402
rect 3702 -433 3736 -422
rect 3739 -433 3748 -417
rect 3764 -433 3773 -417
rect 3780 -422 3790 -402
rect 3800 -422 3814 -402
rect 3815 -415 3826 -402
rect 3780 -433 3814 -422
rect 3815 -433 3826 -417
rect 3872 -426 3888 -410
rect 3895 -412 3925 -360
rect 3959 -364 3960 -357
rect 3944 -372 3960 -364
rect 3931 -404 3944 -385
rect 3959 -404 3989 -388
rect 3931 -420 4005 -404
rect 3931 -422 3944 -420
rect 3959 -422 3993 -420
rect 3596 -444 3609 -442
rect 3624 -444 3658 -442
rect 3596 -460 3658 -444
rect 3702 -449 3718 -446
rect 3780 -449 3810 -438
rect 3858 -442 3904 -426
rect 3931 -438 4005 -422
rect 3858 -444 3892 -442
rect 3857 -460 3904 -444
rect 3931 -460 3944 -438
rect 3959 -460 3989 -438
rect 4016 -460 4017 -444
rect 4032 -460 4045 -300
rect 4075 -404 4088 -300
rect 4133 -322 4134 -312
rect 4149 -322 4162 -312
rect 4133 -326 4162 -322
rect 4167 -326 4197 -300
rect 4215 -314 4231 -312
rect 4303 -314 4356 -300
rect 4304 -316 4368 -314
rect 4411 -316 4426 -300
rect 4475 -303 4505 -300
rect 4475 -306 4511 -303
rect 4441 -314 4457 -312
rect 4215 -326 4230 -322
rect 4133 -328 4230 -326
rect 4258 -328 4426 -316
rect 4442 -326 4457 -322
rect 4475 -325 4514 -306
rect 4533 -312 4540 -311
rect 4539 -319 4540 -312
rect 4523 -322 4524 -319
rect 4539 -322 4552 -319
rect 4475 -326 4505 -325
rect 4514 -326 4520 -325
rect 4523 -326 4552 -322
rect 4442 -327 4552 -326
rect 4442 -328 4558 -327
rect 4117 -336 4168 -328
rect 4117 -348 4142 -336
rect 4149 -348 4168 -336
rect 4199 -336 4249 -328
rect 4199 -344 4215 -336
rect 4222 -338 4249 -336
rect 4258 -338 4479 -328
rect 4222 -348 4479 -338
rect 4508 -336 4558 -328
rect 4508 -345 4524 -336
rect 4117 -356 4168 -348
rect 4215 -356 4479 -348
rect 4505 -348 4524 -345
rect 4531 -348 4558 -336
rect 4505 -356 4558 -348
rect 4133 -364 4134 -356
rect 4149 -364 4162 -356
rect 4133 -372 4149 -364
rect 4130 -379 4149 -376
rect 4130 -388 4152 -379
rect 4103 -398 4152 -388
rect 4103 -404 4133 -398
rect 4152 -403 4157 -398
rect 4075 -420 4149 -404
rect 4167 -412 4197 -356
rect 4232 -366 4440 -356
rect 4475 -360 4520 -356
rect 4523 -357 4524 -356
rect 4539 -357 4552 -356
rect 4258 -396 4447 -366
rect 4273 -399 4447 -396
rect 4266 -402 4447 -399
rect 4075 -422 4088 -420
rect 4103 -422 4137 -420
rect 4075 -438 4149 -422
rect 4176 -426 4189 -412
rect 4204 -426 4220 -410
rect 4266 -415 4277 -402
rect 4059 -460 4060 -444
rect 4075 -460 4088 -438
rect 4103 -460 4133 -438
rect 4176 -442 4238 -426
rect 4266 -433 4277 -417
rect 4282 -422 4292 -402
rect 4302 -422 4316 -402
rect 4319 -415 4328 -402
rect 4344 -415 4353 -402
rect 4282 -433 4316 -422
rect 4319 -433 4328 -417
rect 4344 -433 4353 -417
rect 4360 -422 4370 -402
rect 4380 -422 4394 -402
rect 4395 -415 4406 -402
rect 4360 -433 4394 -422
rect 4395 -433 4406 -417
rect 4452 -426 4468 -410
rect 4475 -412 4505 -360
rect 4539 -364 4540 -357
rect 4524 -372 4540 -364
rect 4511 -404 4524 -385
rect 4539 -404 4569 -388
rect 4511 -420 4585 -404
rect 4511 -422 4524 -420
rect 4539 -422 4573 -420
rect 4176 -444 4189 -442
rect 4204 -444 4238 -442
rect 4176 -460 4238 -444
rect 4282 -449 4298 -446
rect 4360 -449 4390 -438
rect 4438 -442 4484 -426
rect 4511 -438 4585 -422
rect 4438 -444 4472 -442
rect 4437 -460 4484 -444
rect 4511 -460 4524 -438
rect 4539 -460 4569 -438
rect 4596 -460 4597 -444
rect 4612 -460 4625 -300
rect -7 -468 34 -460
rect -7 -494 8 -468
rect 15 -494 34 -468
rect 98 -472 160 -460
rect 172 -472 247 -460
rect 305 -472 380 -460
rect 392 -472 423 -460
rect 429 -472 464 -460
rect 98 -474 260 -472
rect -7 -502 34 -494
rect 116 -498 129 -474
rect 144 -476 159 -474
rect -1 -512 0 -502
rect 15 -512 28 -502
rect 43 -512 73 -498
rect 116 -512 159 -498
rect 183 -501 190 -494
rect 193 -498 260 -474
rect 292 -474 464 -472
rect 262 -496 290 -492
rect 292 -496 372 -474
rect 393 -476 408 -474
rect 262 -498 372 -496
rect 193 -502 372 -498
rect 166 -512 196 -502
rect 198 -512 351 -502
rect 359 -512 389 -502
rect 393 -512 423 -498
rect 451 -512 464 -474
rect 536 -468 571 -460
rect 536 -494 537 -468
rect 544 -494 571 -468
rect 479 -512 509 -498
rect 536 -502 571 -494
rect 573 -468 614 -460
rect 573 -494 588 -468
rect 595 -494 614 -468
rect 678 -472 740 -460
rect 752 -472 827 -460
rect 885 -472 960 -460
rect 972 -472 1003 -460
rect 1009 -472 1044 -460
rect 678 -474 840 -472
rect 573 -502 614 -494
rect 696 -498 709 -474
rect 724 -476 739 -474
rect 536 -512 537 -502
rect 552 -512 565 -502
rect 579 -512 580 -502
rect 595 -512 608 -502
rect 623 -512 653 -498
rect 696 -512 739 -498
rect 763 -501 770 -494
rect 773 -498 840 -474
rect 872 -474 1044 -472
rect 842 -496 870 -492
rect 872 -496 952 -474
rect 973 -476 988 -474
rect 842 -498 952 -496
rect 773 -502 952 -498
rect 746 -512 776 -502
rect 778 -512 931 -502
rect 939 -512 969 -502
rect 973 -512 1003 -498
rect 1031 -512 1044 -474
rect 1116 -468 1151 -460
rect 1116 -494 1117 -468
rect 1124 -494 1151 -468
rect 1059 -512 1089 -498
rect 1116 -502 1151 -494
rect 1153 -468 1194 -460
rect 1153 -494 1168 -468
rect 1175 -494 1194 -468
rect 1258 -472 1320 -460
rect 1332 -472 1407 -460
rect 1465 -472 1540 -460
rect 1552 -472 1583 -460
rect 1589 -472 1624 -460
rect 1258 -474 1420 -472
rect 1153 -502 1194 -494
rect 1276 -498 1289 -474
rect 1304 -476 1319 -474
rect 1116 -512 1117 -502
rect 1132 -512 1145 -502
rect 1159 -512 1160 -502
rect 1175 -512 1188 -502
rect 1203 -512 1233 -498
rect 1276 -512 1319 -498
rect 1343 -501 1350 -494
rect 1353 -498 1420 -474
rect 1452 -474 1624 -472
rect 1422 -496 1450 -492
rect 1452 -496 1532 -474
rect 1553 -476 1568 -474
rect 1422 -498 1532 -496
rect 1353 -502 1532 -498
rect 1326 -512 1356 -502
rect 1358 -512 1511 -502
rect 1519 -512 1549 -502
rect 1553 -512 1583 -498
rect 1611 -512 1624 -474
rect 1696 -468 1731 -460
rect 1696 -494 1697 -468
rect 1704 -494 1731 -468
rect 1639 -512 1669 -498
rect 1696 -502 1731 -494
rect 1733 -468 1774 -460
rect 1733 -494 1748 -468
rect 1755 -494 1774 -468
rect 1838 -472 1900 -460
rect 1912 -472 1987 -460
rect 2045 -472 2120 -460
rect 2132 -472 2163 -460
rect 2169 -472 2204 -460
rect 1838 -474 2000 -472
rect 1733 -502 1774 -494
rect 1856 -498 1869 -474
rect 1884 -476 1899 -474
rect 1696 -512 1697 -502
rect 1712 -512 1725 -502
rect 1739 -512 1740 -502
rect 1755 -512 1768 -502
rect 1783 -512 1813 -498
rect 1856 -512 1899 -498
rect 1923 -501 1930 -494
rect 1933 -498 2000 -474
rect 2032 -474 2204 -472
rect 2002 -496 2030 -492
rect 2032 -496 2112 -474
rect 2133 -476 2148 -474
rect 2002 -498 2112 -496
rect 1933 -502 2112 -498
rect 1906 -512 1936 -502
rect 1938 -512 2091 -502
rect 2099 -512 2129 -502
rect 2133 -512 2163 -498
rect 2191 -512 2204 -474
rect 2276 -468 2311 -460
rect 2276 -494 2277 -468
rect 2284 -494 2311 -468
rect 2219 -512 2249 -498
rect 2276 -502 2311 -494
rect 2313 -468 2354 -460
rect 2313 -494 2328 -468
rect 2335 -494 2354 -468
rect 2418 -472 2480 -460
rect 2492 -472 2567 -460
rect 2625 -472 2700 -460
rect 2712 -472 2743 -460
rect 2749 -472 2784 -460
rect 2418 -474 2580 -472
rect 2313 -502 2354 -494
rect 2436 -498 2449 -474
rect 2464 -476 2479 -474
rect 2276 -512 2277 -502
rect 2292 -512 2305 -502
rect 2319 -512 2320 -502
rect 2335 -512 2348 -502
rect 2363 -512 2393 -498
rect 2436 -512 2479 -498
rect 2503 -501 2510 -494
rect 2513 -498 2580 -474
rect 2612 -474 2784 -472
rect 2582 -496 2610 -492
rect 2612 -496 2692 -474
rect 2713 -476 2728 -474
rect 2582 -498 2692 -496
rect 2513 -502 2692 -498
rect 2486 -512 2516 -502
rect 2518 -512 2671 -502
rect 2679 -512 2709 -502
rect 2713 -512 2743 -498
rect 2771 -512 2784 -474
rect 2856 -468 2891 -460
rect 2856 -494 2857 -468
rect 2864 -494 2891 -468
rect 2799 -512 2829 -498
rect 2856 -502 2891 -494
rect 2893 -468 2934 -460
rect 2893 -494 2908 -468
rect 2915 -494 2934 -468
rect 2998 -472 3060 -460
rect 3072 -472 3147 -460
rect 3205 -472 3280 -460
rect 3292 -472 3323 -460
rect 3329 -472 3364 -460
rect 2998 -474 3160 -472
rect 2893 -502 2934 -494
rect 3016 -498 3029 -474
rect 3044 -476 3059 -474
rect 2856 -512 2857 -502
rect 2872 -512 2885 -502
rect 2899 -512 2900 -502
rect 2915 -512 2928 -502
rect 2943 -512 2973 -498
rect 3016 -512 3059 -498
rect 3083 -501 3090 -494
rect 3093 -498 3160 -474
rect 3192 -474 3364 -472
rect 3162 -496 3190 -492
rect 3192 -496 3272 -474
rect 3293 -476 3308 -474
rect 3162 -498 3272 -496
rect 3093 -502 3272 -498
rect 3066 -512 3096 -502
rect 3098 -512 3251 -502
rect 3259 -512 3289 -502
rect 3293 -512 3323 -498
rect 3351 -512 3364 -474
rect 3436 -468 3471 -460
rect 3436 -494 3437 -468
rect 3444 -494 3471 -468
rect 3379 -512 3409 -498
rect 3436 -502 3471 -494
rect 3473 -468 3514 -460
rect 3473 -494 3488 -468
rect 3495 -494 3514 -468
rect 3578 -472 3640 -460
rect 3652 -472 3727 -460
rect 3785 -472 3860 -460
rect 3872 -472 3903 -460
rect 3909 -472 3944 -460
rect 3578 -474 3740 -472
rect 3473 -502 3514 -494
rect 3596 -498 3609 -474
rect 3624 -476 3639 -474
rect 3436 -512 3437 -502
rect 3452 -512 3465 -502
rect 3479 -512 3480 -502
rect 3495 -512 3508 -502
rect 3523 -512 3553 -498
rect 3596 -512 3639 -498
rect 3663 -501 3670 -494
rect 3673 -498 3740 -474
rect 3772 -474 3944 -472
rect 3742 -496 3770 -492
rect 3772 -496 3852 -474
rect 3873 -476 3888 -474
rect 3742 -498 3852 -496
rect 3673 -502 3852 -498
rect 3646 -512 3676 -502
rect 3678 -512 3831 -502
rect 3839 -512 3869 -502
rect 3873 -512 3903 -498
rect 3931 -512 3944 -474
rect 4016 -468 4051 -460
rect 4016 -494 4017 -468
rect 4024 -494 4051 -468
rect 3959 -512 3989 -498
rect 4016 -502 4051 -494
rect 4053 -468 4094 -460
rect 4053 -494 4068 -468
rect 4075 -494 4094 -468
rect 4158 -472 4220 -460
rect 4232 -472 4307 -460
rect 4365 -472 4440 -460
rect 4452 -472 4483 -460
rect 4489 -472 4524 -460
rect 4158 -474 4320 -472
rect 4053 -502 4094 -494
rect 4176 -498 4189 -474
rect 4204 -476 4219 -474
rect 4016 -512 4017 -502
rect 4032 -512 4045 -502
rect 4059 -512 4060 -502
rect 4075 -512 4088 -502
rect 4103 -512 4133 -498
rect 4176 -512 4219 -498
rect 4243 -501 4250 -494
rect 4253 -498 4320 -474
rect 4352 -474 4524 -472
rect 4322 -496 4350 -492
rect 4352 -496 4432 -474
rect 4453 -476 4468 -474
rect 4322 -498 4432 -496
rect 4253 -502 4432 -498
rect 4226 -512 4256 -502
rect 4258 -512 4411 -502
rect 4419 -512 4449 -502
rect 4453 -512 4483 -498
rect 4511 -512 4524 -474
rect 4596 -468 4631 -460
rect 4596 -494 4597 -468
rect 4604 -494 4631 -468
rect 4539 -512 4569 -498
rect 4596 -502 4631 -494
rect 4596 -512 4597 -502
rect 4612 -512 4625 -502
rect -1 -518 4625 -512
rect 0 -526 4625 -518
rect 15 -556 28 -526
rect 43 -544 73 -526
rect 116 -540 130 -526
rect 166 -540 386 -526
rect 117 -542 130 -540
rect 83 -554 98 -542
rect 80 -556 102 -554
rect 107 -556 137 -542
rect 198 -544 351 -540
rect 180 -556 372 -544
rect 415 -556 445 -542
rect 451 -556 464 -526
rect 479 -544 509 -526
rect 552 -556 565 -526
rect 595 -556 608 -526
rect 623 -544 653 -526
rect 696 -540 710 -526
rect 746 -540 966 -526
rect 697 -542 710 -540
rect 663 -554 678 -542
rect 660 -556 682 -554
rect 687 -556 717 -542
rect 778 -544 931 -540
rect 760 -556 952 -544
rect 995 -556 1025 -542
rect 1031 -556 1044 -526
rect 1059 -544 1089 -526
rect 1132 -556 1145 -526
rect 1175 -556 1188 -526
rect 1203 -544 1233 -526
rect 1276 -540 1290 -526
rect 1326 -540 1546 -526
rect 1277 -542 1290 -540
rect 1243 -554 1258 -542
rect 1240 -556 1262 -554
rect 1267 -556 1297 -542
rect 1358 -544 1511 -540
rect 1340 -556 1532 -544
rect 1575 -556 1605 -542
rect 1611 -556 1624 -526
rect 1639 -544 1669 -526
rect 1712 -556 1725 -526
rect 1755 -556 1768 -526
rect 1783 -544 1813 -526
rect 1856 -540 1870 -526
rect 1906 -540 2126 -526
rect 1857 -542 1870 -540
rect 1823 -554 1838 -542
rect 1820 -556 1842 -554
rect 1847 -556 1877 -542
rect 1938 -544 2091 -540
rect 1920 -556 2112 -544
rect 2155 -556 2185 -542
rect 2191 -556 2204 -526
rect 2219 -544 2249 -526
rect 2292 -556 2305 -526
rect 2335 -556 2348 -526
rect 2363 -544 2393 -526
rect 2436 -540 2450 -526
rect 2486 -540 2706 -526
rect 2437 -542 2450 -540
rect 2403 -554 2418 -542
rect 2400 -556 2422 -554
rect 2427 -556 2457 -542
rect 2518 -544 2671 -540
rect 2500 -556 2692 -544
rect 2735 -556 2765 -542
rect 2771 -556 2784 -526
rect 2799 -544 2829 -526
rect 2872 -556 2885 -526
rect 2915 -556 2928 -526
rect 2943 -544 2973 -526
rect 3016 -540 3030 -526
rect 3066 -540 3286 -526
rect 3017 -542 3030 -540
rect 2983 -554 2998 -542
rect 2980 -556 3002 -554
rect 3007 -556 3037 -542
rect 3098 -544 3251 -540
rect 3080 -556 3272 -544
rect 3315 -556 3345 -542
rect 3351 -556 3364 -526
rect 3379 -544 3409 -526
rect 3452 -556 3465 -526
rect 3495 -556 3508 -526
rect 3523 -544 3553 -526
rect 3596 -540 3610 -526
rect 3646 -540 3866 -526
rect 3597 -542 3610 -540
rect 3563 -554 3578 -542
rect 3560 -556 3582 -554
rect 3587 -556 3617 -542
rect 3678 -544 3831 -540
rect 3660 -556 3852 -544
rect 3895 -556 3925 -542
rect 3931 -556 3944 -526
rect 3959 -544 3989 -526
rect 4032 -556 4045 -526
rect 4075 -556 4088 -526
rect 4103 -544 4133 -526
rect 4176 -540 4190 -526
rect 4226 -540 4446 -526
rect 4177 -542 4190 -540
rect 4143 -554 4158 -542
rect 4140 -556 4162 -554
rect 4167 -556 4197 -542
rect 4258 -544 4411 -540
rect 4240 -556 4432 -544
rect 4475 -556 4505 -542
rect 4511 -556 4524 -526
rect 4539 -544 4569 -526
rect 4612 -556 4625 -526
rect 0 -570 4625 -556
rect 15 -674 28 -570
rect 73 -592 74 -582
rect 89 -592 102 -582
rect 73 -596 102 -592
rect 107 -596 137 -570
rect 155 -584 171 -582
rect 243 -584 296 -570
rect 244 -586 308 -584
rect 351 -586 366 -570
rect 415 -573 445 -570
rect 415 -576 451 -573
rect 381 -584 397 -582
rect 155 -596 170 -592
rect 73 -598 170 -596
rect 198 -598 366 -586
rect 382 -596 397 -592
rect 415 -595 454 -576
rect 473 -582 480 -581
rect 479 -589 480 -582
rect 463 -592 464 -589
rect 479 -592 492 -589
rect 415 -596 445 -595
rect 454 -596 460 -595
rect 463 -596 492 -592
rect 382 -597 492 -596
rect 382 -598 498 -597
rect 57 -606 108 -598
rect 57 -618 82 -606
rect 89 -618 108 -606
rect 139 -606 189 -598
rect 139 -614 155 -606
rect 162 -608 189 -606
rect 198 -608 419 -598
rect 162 -618 419 -608
rect 448 -606 498 -598
rect 448 -615 464 -606
rect 57 -626 108 -618
rect 155 -626 419 -618
rect 445 -618 464 -615
rect 471 -618 498 -606
rect 445 -626 498 -618
rect 73 -634 74 -626
rect 89 -634 102 -626
rect 73 -642 89 -634
rect 70 -649 89 -646
rect 70 -658 92 -649
rect 43 -668 92 -658
rect 43 -674 73 -668
rect 92 -673 97 -668
rect 15 -690 89 -674
rect 107 -682 137 -626
rect 172 -636 380 -626
rect 415 -630 460 -626
rect 463 -627 464 -626
rect 479 -627 492 -626
rect 198 -666 387 -636
rect 213 -669 387 -666
rect 206 -672 387 -669
rect 15 -692 28 -690
rect 43 -692 77 -690
rect 15 -708 89 -692
rect 116 -696 129 -682
rect 144 -696 160 -680
rect 206 -685 217 -672
rect -1 -730 0 -714
rect 15 -730 28 -708
rect 43 -730 73 -708
rect 116 -712 178 -696
rect 206 -703 217 -687
rect 222 -692 232 -672
rect 242 -692 256 -672
rect 259 -685 268 -672
rect 284 -685 293 -672
rect 222 -703 256 -692
rect 259 -703 268 -687
rect 284 -703 293 -687
rect 300 -692 310 -672
rect 320 -692 334 -672
rect 335 -685 346 -672
rect 300 -703 334 -692
rect 335 -703 346 -687
rect 392 -696 408 -680
rect 415 -682 445 -630
rect 479 -634 480 -627
rect 464 -642 480 -634
rect 451 -674 464 -655
rect 479 -674 509 -658
rect 451 -690 525 -674
rect 451 -692 464 -690
rect 479 -692 513 -690
rect 116 -714 129 -712
rect 144 -714 178 -712
rect 116 -730 178 -714
rect 222 -719 238 -716
rect 300 -719 330 -708
rect 378 -712 424 -696
rect 451 -708 525 -692
rect 378 -714 412 -712
rect 377 -730 424 -714
rect 451 -730 464 -708
rect 479 -730 509 -708
rect 536 -730 537 -714
rect 552 -730 565 -570
rect 595 -674 608 -570
rect 653 -592 654 -582
rect 669 -592 682 -582
rect 653 -596 682 -592
rect 687 -596 717 -570
rect 735 -584 751 -582
rect 823 -584 876 -570
rect 824 -586 888 -584
rect 931 -586 946 -570
rect 995 -573 1025 -570
rect 995 -576 1031 -573
rect 961 -584 977 -582
rect 735 -596 750 -592
rect 653 -598 750 -596
rect 778 -598 946 -586
rect 962 -596 977 -592
rect 995 -595 1034 -576
rect 1053 -582 1060 -581
rect 1059 -589 1060 -582
rect 1043 -592 1044 -589
rect 1059 -592 1072 -589
rect 995 -596 1025 -595
rect 1034 -596 1040 -595
rect 1043 -596 1072 -592
rect 962 -597 1072 -596
rect 962 -598 1078 -597
rect 637 -606 688 -598
rect 637 -618 662 -606
rect 669 -618 688 -606
rect 719 -606 769 -598
rect 719 -614 735 -606
rect 742 -608 769 -606
rect 778 -608 999 -598
rect 742 -618 999 -608
rect 1028 -606 1078 -598
rect 1028 -615 1044 -606
rect 637 -626 688 -618
rect 735 -626 999 -618
rect 1025 -618 1044 -615
rect 1051 -618 1078 -606
rect 1025 -626 1078 -618
rect 653 -634 654 -626
rect 669 -634 682 -626
rect 653 -642 669 -634
rect 650 -649 669 -646
rect 650 -658 672 -649
rect 623 -668 672 -658
rect 623 -674 653 -668
rect 672 -673 677 -668
rect 595 -690 669 -674
rect 687 -682 717 -626
rect 752 -636 960 -626
rect 995 -630 1040 -626
rect 1043 -627 1044 -626
rect 1059 -627 1072 -626
rect 778 -666 967 -636
rect 793 -669 967 -666
rect 786 -672 967 -669
rect 595 -692 608 -690
rect 623 -692 657 -690
rect 595 -708 669 -692
rect 696 -696 709 -682
rect 724 -696 740 -680
rect 786 -685 797 -672
rect 579 -730 580 -714
rect 595 -730 608 -708
rect 623 -730 653 -708
rect 696 -712 758 -696
rect 786 -703 797 -687
rect 802 -692 812 -672
rect 822 -692 836 -672
rect 839 -685 848 -672
rect 864 -685 873 -672
rect 802 -703 836 -692
rect 839 -703 848 -687
rect 864 -703 873 -687
rect 880 -692 890 -672
rect 900 -692 914 -672
rect 915 -685 926 -672
rect 880 -703 914 -692
rect 915 -703 926 -687
rect 972 -696 988 -680
rect 995 -682 1025 -630
rect 1059 -634 1060 -627
rect 1044 -642 1060 -634
rect 1031 -674 1044 -655
rect 1059 -674 1089 -658
rect 1031 -690 1105 -674
rect 1031 -692 1044 -690
rect 1059 -692 1093 -690
rect 696 -714 709 -712
rect 724 -714 758 -712
rect 696 -730 758 -714
rect 802 -719 818 -716
rect 880 -719 910 -708
rect 958 -712 1004 -696
rect 1031 -708 1105 -692
rect 958 -714 992 -712
rect 957 -730 1004 -714
rect 1031 -730 1044 -708
rect 1059 -730 1089 -708
rect 1116 -730 1117 -714
rect 1132 -730 1145 -570
rect 1175 -674 1188 -570
rect 1233 -592 1234 -582
rect 1249 -592 1262 -582
rect 1233 -596 1262 -592
rect 1267 -596 1297 -570
rect 1315 -584 1331 -582
rect 1403 -584 1456 -570
rect 1404 -586 1468 -584
rect 1511 -586 1526 -570
rect 1575 -573 1605 -570
rect 1575 -576 1611 -573
rect 1541 -584 1557 -582
rect 1315 -596 1330 -592
rect 1233 -598 1330 -596
rect 1358 -598 1526 -586
rect 1542 -596 1557 -592
rect 1575 -595 1614 -576
rect 1633 -582 1640 -581
rect 1639 -589 1640 -582
rect 1623 -592 1624 -589
rect 1639 -592 1652 -589
rect 1575 -596 1605 -595
rect 1614 -596 1620 -595
rect 1623 -596 1652 -592
rect 1542 -597 1652 -596
rect 1542 -598 1658 -597
rect 1217 -606 1268 -598
rect 1217 -618 1242 -606
rect 1249 -618 1268 -606
rect 1299 -606 1349 -598
rect 1299 -614 1315 -606
rect 1322 -608 1349 -606
rect 1358 -608 1579 -598
rect 1322 -618 1579 -608
rect 1608 -606 1658 -598
rect 1608 -615 1624 -606
rect 1217 -626 1268 -618
rect 1315 -626 1579 -618
rect 1605 -618 1624 -615
rect 1631 -618 1658 -606
rect 1605 -626 1658 -618
rect 1233 -634 1234 -626
rect 1249 -634 1262 -626
rect 1233 -642 1249 -634
rect 1230 -649 1249 -646
rect 1230 -658 1252 -649
rect 1203 -668 1252 -658
rect 1203 -674 1233 -668
rect 1252 -673 1257 -668
rect 1175 -690 1249 -674
rect 1267 -682 1297 -626
rect 1332 -636 1540 -626
rect 1575 -630 1620 -626
rect 1623 -627 1624 -626
rect 1639 -627 1652 -626
rect 1358 -666 1547 -636
rect 1373 -669 1547 -666
rect 1366 -672 1547 -669
rect 1175 -692 1188 -690
rect 1203 -692 1237 -690
rect 1175 -708 1249 -692
rect 1276 -696 1289 -682
rect 1304 -696 1320 -680
rect 1366 -685 1377 -672
rect 1159 -730 1160 -714
rect 1175 -730 1188 -708
rect 1203 -730 1233 -708
rect 1276 -712 1338 -696
rect 1366 -703 1377 -687
rect 1382 -692 1392 -672
rect 1402 -692 1416 -672
rect 1419 -685 1428 -672
rect 1444 -685 1453 -672
rect 1382 -703 1416 -692
rect 1419 -703 1428 -687
rect 1444 -703 1453 -687
rect 1460 -692 1470 -672
rect 1480 -692 1494 -672
rect 1495 -685 1506 -672
rect 1460 -703 1494 -692
rect 1495 -703 1506 -687
rect 1552 -696 1568 -680
rect 1575 -682 1605 -630
rect 1639 -634 1640 -627
rect 1624 -642 1640 -634
rect 1611 -674 1624 -655
rect 1639 -674 1669 -658
rect 1611 -690 1685 -674
rect 1611 -692 1624 -690
rect 1639 -692 1673 -690
rect 1276 -714 1289 -712
rect 1304 -714 1338 -712
rect 1276 -730 1338 -714
rect 1382 -719 1398 -716
rect 1460 -719 1490 -708
rect 1538 -712 1584 -696
rect 1611 -708 1685 -692
rect 1538 -714 1572 -712
rect 1537 -730 1584 -714
rect 1611 -730 1624 -708
rect 1639 -730 1669 -708
rect 1696 -730 1697 -714
rect 1712 -730 1725 -570
rect 1755 -674 1768 -570
rect 1813 -592 1814 -582
rect 1829 -592 1842 -582
rect 1813 -596 1842 -592
rect 1847 -596 1877 -570
rect 1895 -584 1911 -582
rect 1983 -584 2036 -570
rect 1984 -586 2048 -584
rect 2091 -586 2106 -570
rect 2155 -573 2185 -570
rect 2155 -576 2191 -573
rect 2121 -584 2137 -582
rect 1895 -596 1910 -592
rect 1813 -598 1910 -596
rect 1938 -598 2106 -586
rect 2122 -596 2137 -592
rect 2155 -595 2194 -576
rect 2213 -582 2220 -581
rect 2219 -589 2220 -582
rect 2203 -592 2204 -589
rect 2219 -592 2232 -589
rect 2155 -596 2185 -595
rect 2194 -596 2200 -595
rect 2203 -596 2232 -592
rect 2122 -597 2232 -596
rect 2122 -598 2238 -597
rect 1797 -606 1848 -598
rect 1797 -618 1822 -606
rect 1829 -618 1848 -606
rect 1879 -606 1929 -598
rect 1879 -614 1895 -606
rect 1902 -608 1929 -606
rect 1938 -608 2159 -598
rect 1902 -618 2159 -608
rect 2188 -606 2238 -598
rect 2188 -615 2204 -606
rect 1797 -626 1848 -618
rect 1895 -626 2159 -618
rect 2185 -618 2204 -615
rect 2211 -618 2238 -606
rect 2185 -626 2238 -618
rect 1813 -634 1814 -626
rect 1829 -634 1842 -626
rect 1813 -642 1829 -634
rect 1810 -649 1829 -646
rect 1810 -658 1832 -649
rect 1783 -668 1832 -658
rect 1783 -674 1813 -668
rect 1832 -673 1837 -668
rect 1755 -690 1829 -674
rect 1847 -682 1877 -626
rect 1912 -636 2120 -626
rect 2155 -630 2200 -626
rect 2203 -627 2204 -626
rect 2219 -627 2232 -626
rect 1938 -666 2127 -636
rect 1953 -669 2127 -666
rect 1946 -672 2127 -669
rect 1755 -692 1768 -690
rect 1783 -692 1817 -690
rect 1755 -708 1829 -692
rect 1856 -696 1869 -682
rect 1884 -696 1900 -680
rect 1946 -685 1957 -672
rect 1739 -730 1740 -714
rect 1755 -730 1768 -708
rect 1783 -730 1813 -708
rect 1856 -712 1918 -696
rect 1946 -703 1957 -687
rect 1962 -692 1972 -672
rect 1982 -692 1996 -672
rect 1999 -685 2008 -672
rect 2024 -685 2033 -672
rect 1962 -703 1996 -692
rect 1999 -703 2008 -687
rect 2024 -703 2033 -687
rect 2040 -692 2050 -672
rect 2060 -692 2074 -672
rect 2075 -685 2086 -672
rect 2040 -703 2074 -692
rect 2075 -703 2086 -687
rect 2132 -696 2148 -680
rect 2155 -682 2185 -630
rect 2219 -634 2220 -627
rect 2204 -642 2220 -634
rect 2191 -674 2204 -655
rect 2219 -674 2249 -658
rect 2191 -690 2265 -674
rect 2191 -692 2204 -690
rect 2219 -692 2253 -690
rect 1856 -714 1869 -712
rect 1884 -714 1918 -712
rect 1856 -730 1918 -714
rect 1962 -719 1978 -716
rect 2040 -719 2070 -708
rect 2118 -712 2164 -696
rect 2191 -708 2265 -692
rect 2118 -714 2152 -712
rect 2117 -730 2164 -714
rect 2191 -730 2204 -708
rect 2219 -730 2249 -708
rect 2276 -730 2277 -714
rect 2292 -730 2305 -570
rect 2335 -674 2348 -570
rect 2393 -592 2394 -582
rect 2409 -592 2422 -582
rect 2393 -596 2422 -592
rect 2427 -596 2457 -570
rect 2475 -584 2491 -582
rect 2563 -584 2616 -570
rect 2564 -586 2628 -584
rect 2671 -586 2686 -570
rect 2735 -573 2765 -570
rect 2735 -576 2771 -573
rect 2701 -584 2717 -582
rect 2475 -596 2490 -592
rect 2393 -598 2490 -596
rect 2518 -598 2686 -586
rect 2702 -596 2717 -592
rect 2735 -595 2774 -576
rect 2793 -582 2800 -581
rect 2799 -589 2800 -582
rect 2783 -592 2784 -589
rect 2799 -592 2812 -589
rect 2735 -596 2765 -595
rect 2774 -596 2780 -595
rect 2783 -596 2812 -592
rect 2702 -597 2812 -596
rect 2702 -598 2818 -597
rect 2377 -606 2428 -598
rect 2377 -618 2402 -606
rect 2409 -618 2428 -606
rect 2459 -606 2509 -598
rect 2459 -614 2475 -606
rect 2482 -608 2509 -606
rect 2518 -608 2739 -598
rect 2482 -618 2739 -608
rect 2768 -606 2818 -598
rect 2768 -615 2784 -606
rect 2377 -626 2428 -618
rect 2475 -626 2739 -618
rect 2765 -618 2784 -615
rect 2791 -618 2818 -606
rect 2765 -626 2818 -618
rect 2393 -634 2394 -626
rect 2409 -634 2422 -626
rect 2393 -642 2409 -634
rect 2390 -649 2409 -646
rect 2390 -658 2412 -649
rect 2363 -668 2412 -658
rect 2363 -674 2393 -668
rect 2412 -673 2417 -668
rect 2335 -690 2409 -674
rect 2427 -682 2457 -626
rect 2492 -636 2700 -626
rect 2735 -630 2780 -626
rect 2783 -627 2784 -626
rect 2799 -627 2812 -626
rect 2518 -666 2707 -636
rect 2533 -669 2707 -666
rect 2526 -672 2707 -669
rect 2335 -692 2348 -690
rect 2363 -692 2397 -690
rect 2335 -708 2409 -692
rect 2436 -696 2449 -682
rect 2464 -696 2480 -680
rect 2526 -685 2537 -672
rect 2319 -730 2320 -714
rect 2335 -730 2348 -708
rect 2363 -730 2393 -708
rect 2436 -712 2498 -696
rect 2526 -703 2537 -687
rect 2542 -692 2552 -672
rect 2562 -692 2576 -672
rect 2579 -685 2588 -672
rect 2604 -685 2613 -672
rect 2542 -703 2576 -692
rect 2579 -703 2588 -687
rect 2604 -703 2613 -687
rect 2620 -692 2630 -672
rect 2640 -692 2654 -672
rect 2655 -685 2666 -672
rect 2620 -703 2654 -692
rect 2655 -703 2666 -687
rect 2712 -696 2728 -680
rect 2735 -682 2765 -630
rect 2799 -634 2800 -627
rect 2784 -642 2800 -634
rect 2771 -674 2784 -655
rect 2799 -674 2829 -658
rect 2771 -690 2845 -674
rect 2771 -692 2784 -690
rect 2799 -692 2833 -690
rect 2436 -714 2449 -712
rect 2464 -714 2498 -712
rect 2436 -730 2498 -714
rect 2542 -719 2558 -716
rect 2620 -719 2650 -708
rect 2698 -712 2744 -696
rect 2771 -708 2845 -692
rect 2698 -714 2732 -712
rect 2697 -730 2744 -714
rect 2771 -730 2784 -708
rect 2799 -730 2829 -708
rect 2856 -730 2857 -714
rect 2872 -730 2885 -570
rect 2915 -674 2928 -570
rect 2973 -592 2974 -582
rect 2989 -592 3002 -582
rect 2973 -596 3002 -592
rect 3007 -596 3037 -570
rect 3055 -584 3071 -582
rect 3143 -584 3196 -570
rect 3144 -586 3208 -584
rect 3251 -586 3266 -570
rect 3315 -573 3345 -570
rect 3315 -576 3351 -573
rect 3281 -584 3297 -582
rect 3055 -596 3070 -592
rect 2973 -598 3070 -596
rect 3098 -598 3266 -586
rect 3282 -596 3297 -592
rect 3315 -595 3354 -576
rect 3373 -582 3380 -581
rect 3379 -589 3380 -582
rect 3363 -592 3364 -589
rect 3379 -592 3392 -589
rect 3315 -596 3345 -595
rect 3354 -596 3360 -595
rect 3363 -596 3392 -592
rect 3282 -597 3392 -596
rect 3282 -598 3398 -597
rect 2957 -606 3008 -598
rect 2957 -618 2982 -606
rect 2989 -618 3008 -606
rect 3039 -606 3089 -598
rect 3039 -614 3055 -606
rect 3062 -608 3089 -606
rect 3098 -608 3319 -598
rect 3062 -618 3319 -608
rect 3348 -606 3398 -598
rect 3348 -615 3364 -606
rect 2957 -626 3008 -618
rect 3055 -626 3319 -618
rect 3345 -618 3364 -615
rect 3371 -618 3398 -606
rect 3345 -626 3398 -618
rect 2973 -634 2974 -626
rect 2989 -634 3002 -626
rect 2973 -642 2989 -634
rect 2970 -649 2989 -646
rect 2970 -658 2992 -649
rect 2943 -668 2992 -658
rect 2943 -674 2973 -668
rect 2992 -673 2997 -668
rect 2915 -690 2989 -674
rect 3007 -682 3037 -626
rect 3072 -636 3280 -626
rect 3315 -630 3360 -626
rect 3363 -627 3364 -626
rect 3379 -627 3392 -626
rect 3098 -666 3287 -636
rect 3113 -669 3287 -666
rect 3106 -672 3287 -669
rect 2915 -692 2928 -690
rect 2943 -692 2977 -690
rect 2915 -708 2989 -692
rect 3016 -696 3029 -682
rect 3044 -696 3060 -680
rect 3106 -685 3117 -672
rect 2899 -730 2900 -714
rect 2915 -730 2928 -708
rect 2943 -730 2973 -708
rect 3016 -712 3078 -696
rect 3106 -703 3117 -687
rect 3122 -692 3132 -672
rect 3142 -692 3156 -672
rect 3159 -685 3168 -672
rect 3184 -685 3193 -672
rect 3122 -703 3156 -692
rect 3159 -703 3168 -687
rect 3184 -703 3193 -687
rect 3200 -692 3210 -672
rect 3220 -692 3234 -672
rect 3235 -685 3246 -672
rect 3200 -703 3234 -692
rect 3235 -703 3246 -687
rect 3292 -696 3308 -680
rect 3315 -682 3345 -630
rect 3379 -634 3380 -627
rect 3364 -642 3380 -634
rect 3351 -674 3364 -655
rect 3379 -674 3409 -658
rect 3351 -690 3425 -674
rect 3351 -692 3364 -690
rect 3379 -692 3413 -690
rect 3016 -714 3029 -712
rect 3044 -714 3078 -712
rect 3016 -730 3078 -714
rect 3122 -719 3138 -716
rect 3200 -719 3230 -708
rect 3278 -712 3324 -696
rect 3351 -708 3425 -692
rect 3278 -714 3312 -712
rect 3277 -730 3324 -714
rect 3351 -730 3364 -708
rect 3379 -730 3409 -708
rect 3436 -730 3437 -714
rect 3452 -730 3465 -570
rect 3495 -674 3508 -570
rect 3553 -592 3554 -582
rect 3569 -592 3582 -582
rect 3553 -596 3582 -592
rect 3587 -596 3617 -570
rect 3635 -584 3651 -582
rect 3723 -584 3776 -570
rect 3724 -586 3788 -584
rect 3831 -586 3846 -570
rect 3895 -573 3925 -570
rect 3895 -576 3931 -573
rect 3861 -584 3877 -582
rect 3635 -596 3650 -592
rect 3553 -598 3650 -596
rect 3678 -598 3846 -586
rect 3862 -596 3877 -592
rect 3895 -595 3934 -576
rect 3953 -582 3960 -581
rect 3959 -589 3960 -582
rect 3943 -592 3944 -589
rect 3959 -592 3972 -589
rect 3895 -596 3925 -595
rect 3934 -596 3940 -595
rect 3943 -596 3972 -592
rect 3862 -597 3972 -596
rect 3862 -598 3978 -597
rect 3537 -606 3588 -598
rect 3537 -618 3562 -606
rect 3569 -618 3588 -606
rect 3619 -606 3669 -598
rect 3619 -614 3635 -606
rect 3642 -608 3669 -606
rect 3678 -608 3899 -598
rect 3642 -618 3899 -608
rect 3928 -606 3978 -598
rect 3928 -615 3944 -606
rect 3537 -626 3588 -618
rect 3635 -626 3899 -618
rect 3925 -618 3944 -615
rect 3951 -618 3978 -606
rect 3925 -626 3978 -618
rect 3553 -634 3554 -626
rect 3569 -634 3582 -626
rect 3553 -642 3569 -634
rect 3550 -649 3569 -646
rect 3550 -658 3572 -649
rect 3523 -668 3572 -658
rect 3523 -674 3553 -668
rect 3572 -673 3577 -668
rect 3495 -690 3569 -674
rect 3587 -682 3617 -626
rect 3652 -636 3860 -626
rect 3895 -630 3940 -626
rect 3943 -627 3944 -626
rect 3959 -627 3972 -626
rect 3678 -666 3867 -636
rect 3693 -669 3867 -666
rect 3686 -672 3867 -669
rect 3495 -692 3508 -690
rect 3523 -692 3557 -690
rect 3495 -708 3569 -692
rect 3596 -696 3609 -682
rect 3624 -696 3640 -680
rect 3686 -685 3697 -672
rect 3479 -730 3480 -714
rect 3495 -730 3508 -708
rect 3523 -730 3553 -708
rect 3596 -712 3658 -696
rect 3686 -703 3697 -687
rect 3702 -692 3712 -672
rect 3722 -692 3736 -672
rect 3739 -685 3748 -672
rect 3764 -685 3773 -672
rect 3702 -703 3736 -692
rect 3739 -703 3748 -687
rect 3764 -703 3773 -687
rect 3780 -692 3790 -672
rect 3800 -692 3814 -672
rect 3815 -685 3826 -672
rect 3780 -703 3814 -692
rect 3815 -703 3826 -687
rect 3872 -696 3888 -680
rect 3895 -682 3925 -630
rect 3959 -634 3960 -627
rect 3944 -642 3960 -634
rect 3931 -674 3944 -655
rect 3959 -674 3989 -658
rect 3931 -690 4005 -674
rect 3931 -692 3944 -690
rect 3959 -692 3993 -690
rect 3596 -714 3609 -712
rect 3624 -714 3658 -712
rect 3596 -730 3658 -714
rect 3702 -719 3718 -716
rect 3780 -719 3810 -708
rect 3858 -712 3904 -696
rect 3931 -708 4005 -692
rect 3858 -714 3892 -712
rect 3857 -730 3904 -714
rect 3931 -730 3944 -708
rect 3959 -730 3989 -708
rect 4016 -730 4017 -714
rect 4032 -730 4045 -570
rect 4075 -674 4088 -570
rect 4133 -592 4134 -582
rect 4149 -592 4162 -582
rect 4133 -596 4162 -592
rect 4167 -596 4197 -570
rect 4215 -584 4231 -582
rect 4303 -584 4356 -570
rect 4304 -586 4368 -584
rect 4411 -586 4426 -570
rect 4475 -573 4505 -570
rect 4475 -576 4511 -573
rect 4441 -584 4457 -582
rect 4215 -596 4230 -592
rect 4133 -598 4230 -596
rect 4258 -598 4426 -586
rect 4442 -596 4457 -592
rect 4475 -595 4514 -576
rect 4533 -582 4540 -581
rect 4539 -589 4540 -582
rect 4523 -592 4524 -589
rect 4539 -592 4552 -589
rect 4475 -596 4505 -595
rect 4514 -596 4520 -595
rect 4523 -596 4552 -592
rect 4442 -597 4552 -596
rect 4442 -598 4558 -597
rect 4117 -606 4168 -598
rect 4117 -618 4142 -606
rect 4149 -618 4168 -606
rect 4199 -606 4249 -598
rect 4199 -614 4215 -606
rect 4222 -608 4249 -606
rect 4258 -608 4479 -598
rect 4222 -618 4479 -608
rect 4508 -606 4558 -598
rect 4508 -615 4524 -606
rect 4117 -626 4168 -618
rect 4215 -626 4479 -618
rect 4505 -618 4524 -615
rect 4531 -618 4558 -606
rect 4505 -626 4558 -618
rect 4133 -634 4134 -626
rect 4149 -634 4162 -626
rect 4133 -642 4149 -634
rect 4130 -649 4149 -646
rect 4130 -658 4152 -649
rect 4103 -668 4152 -658
rect 4103 -674 4133 -668
rect 4152 -673 4157 -668
rect 4075 -690 4149 -674
rect 4167 -682 4197 -626
rect 4232 -636 4440 -626
rect 4475 -630 4520 -626
rect 4523 -627 4524 -626
rect 4539 -627 4552 -626
rect 4258 -666 4447 -636
rect 4273 -669 4447 -666
rect 4266 -672 4447 -669
rect 4075 -692 4088 -690
rect 4103 -692 4137 -690
rect 4075 -708 4149 -692
rect 4176 -696 4189 -682
rect 4204 -696 4220 -680
rect 4266 -685 4277 -672
rect 4059 -730 4060 -714
rect 4075 -730 4088 -708
rect 4103 -730 4133 -708
rect 4176 -712 4238 -696
rect 4266 -703 4277 -687
rect 4282 -692 4292 -672
rect 4302 -692 4316 -672
rect 4319 -685 4328 -672
rect 4344 -685 4353 -672
rect 4282 -703 4316 -692
rect 4319 -703 4328 -687
rect 4344 -703 4353 -687
rect 4360 -692 4370 -672
rect 4380 -692 4394 -672
rect 4395 -685 4406 -672
rect 4360 -703 4394 -692
rect 4395 -703 4406 -687
rect 4452 -696 4468 -680
rect 4475 -682 4505 -630
rect 4539 -634 4540 -627
rect 4524 -642 4540 -634
rect 4511 -674 4524 -655
rect 4539 -674 4569 -658
rect 4511 -690 4585 -674
rect 4511 -692 4524 -690
rect 4539 -692 4573 -690
rect 4176 -714 4189 -712
rect 4204 -714 4238 -712
rect 4176 -730 4238 -714
rect 4282 -719 4298 -716
rect 4360 -719 4390 -708
rect 4438 -712 4484 -696
rect 4511 -708 4585 -692
rect 4438 -714 4472 -712
rect 4437 -730 4484 -714
rect 4511 -730 4524 -708
rect 4539 -730 4569 -708
rect 4596 -730 4597 -714
rect 4612 -730 4625 -570
rect -7 -738 34 -730
rect -7 -764 8 -738
rect 15 -764 34 -738
rect 98 -742 160 -730
rect 172 -742 247 -730
rect 305 -742 380 -730
rect 392 -742 423 -730
rect 429 -742 464 -730
rect 98 -744 260 -742
rect -7 -772 34 -764
rect 116 -768 129 -744
rect 144 -746 159 -744
rect -1 -782 0 -772
rect 15 -782 28 -772
rect 43 -782 73 -768
rect 116 -782 159 -768
rect 183 -771 190 -764
rect 193 -768 260 -744
rect 292 -744 464 -742
rect 262 -766 290 -762
rect 292 -766 372 -744
rect 393 -746 408 -744
rect 262 -768 372 -766
rect 193 -772 372 -768
rect 166 -782 196 -772
rect 198 -782 351 -772
rect 359 -782 389 -772
rect 393 -782 423 -768
rect 451 -782 464 -744
rect 536 -738 571 -730
rect 536 -764 537 -738
rect 544 -764 571 -738
rect 479 -782 509 -768
rect 536 -772 571 -764
rect 573 -738 614 -730
rect 573 -764 588 -738
rect 595 -764 614 -738
rect 678 -742 740 -730
rect 752 -742 827 -730
rect 885 -742 960 -730
rect 972 -742 1003 -730
rect 1009 -742 1044 -730
rect 678 -744 840 -742
rect 573 -772 614 -764
rect 696 -768 709 -744
rect 724 -746 739 -744
rect 536 -782 537 -772
rect 552 -782 565 -772
rect 579 -782 580 -772
rect 595 -782 608 -772
rect 623 -782 653 -768
rect 696 -782 739 -768
rect 763 -771 770 -764
rect 773 -768 840 -744
rect 872 -744 1044 -742
rect 842 -766 870 -762
rect 872 -766 952 -744
rect 973 -746 988 -744
rect 842 -768 952 -766
rect 773 -772 952 -768
rect 746 -782 776 -772
rect 778 -782 931 -772
rect 939 -782 969 -772
rect 973 -782 1003 -768
rect 1031 -782 1044 -744
rect 1116 -738 1151 -730
rect 1116 -764 1117 -738
rect 1124 -764 1151 -738
rect 1059 -782 1089 -768
rect 1116 -772 1151 -764
rect 1153 -738 1194 -730
rect 1153 -764 1168 -738
rect 1175 -764 1194 -738
rect 1258 -742 1320 -730
rect 1332 -742 1407 -730
rect 1465 -742 1540 -730
rect 1552 -742 1583 -730
rect 1589 -742 1624 -730
rect 1258 -744 1420 -742
rect 1153 -772 1194 -764
rect 1276 -768 1289 -744
rect 1304 -746 1319 -744
rect 1116 -782 1117 -772
rect 1132 -782 1145 -772
rect 1159 -782 1160 -772
rect 1175 -782 1188 -772
rect 1203 -782 1233 -768
rect 1276 -782 1319 -768
rect 1343 -771 1350 -764
rect 1353 -768 1420 -744
rect 1452 -744 1624 -742
rect 1422 -766 1450 -762
rect 1452 -766 1532 -744
rect 1553 -746 1568 -744
rect 1422 -768 1532 -766
rect 1353 -772 1532 -768
rect 1326 -782 1356 -772
rect 1358 -782 1511 -772
rect 1519 -782 1549 -772
rect 1553 -782 1583 -768
rect 1611 -782 1624 -744
rect 1696 -738 1731 -730
rect 1696 -764 1697 -738
rect 1704 -764 1731 -738
rect 1639 -782 1669 -768
rect 1696 -772 1731 -764
rect 1733 -738 1774 -730
rect 1733 -764 1748 -738
rect 1755 -764 1774 -738
rect 1838 -742 1900 -730
rect 1912 -742 1987 -730
rect 2045 -742 2120 -730
rect 2132 -742 2163 -730
rect 2169 -742 2204 -730
rect 1838 -744 2000 -742
rect 1733 -772 1774 -764
rect 1856 -768 1869 -744
rect 1884 -746 1899 -744
rect 1696 -782 1697 -772
rect 1712 -782 1725 -772
rect 1739 -782 1740 -772
rect 1755 -782 1768 -772
rect 1783 -782 1813 -768
rect 1856 -782 1899 -768
rect 1923 -771 1930 -764
rect 1933 -768 2000 -744
rect 2032 -744 2204 -742
rect 2002 -766 2030 -762
rect 2032 -766 2112 -744
rect 2133 -746 2148 -744
rect 2002 -768 2112 -766
rect 1933 -772 2112 -768
rect 1906 -782 1936 -772
rect 1938 -782 2091 -772
rect 2099 -782 2129 -772
rect 2133 -782 2163 -768
rect 2191 -782 2204 -744
rect 2276 -738 2311 -730
rect 2276 -764 2277 -738
rect 2284 -764 2311 -738
rect 2219 -782 2249 -768
rect 2276 -772 2311 -764
rect 2313 -738 2354 -730
rect 2313 -764 2328 -738
rect 2335 -764 2354 -738
rect 2418 -742 2480 -730
rect 2492 -742 2567 -730
rect 2625 -742 2700 -730
rect 2712 -742 2743 -730
rect 2749 -742 2784 -730
rect 2418 -744 2580 -742
rect 2313 -772 2354 -764
rect 2436 -768 2449 -744
rect 2464 -746 2479 -744
rect 2276 -782 2277 -772
rect 2292 -782 2305 -772
rect 2319 -782 2320 -772
rect 2335 -782 2348 -772
rect 2363 -782 2393 -768
rect 2436 -782 2479 -768
rect 2503 -771 2510 -764
rect 2513 -768 2580 -744
rect 2612 -744 2784 -742
rect 2582 -766 2610 -762
rect 2612 -766 2692 -744
rect 2713 -746 2728 -744
rect 2582 -768 2692 -766
rect 2513 -772 2692 -768
rect 2486 -782 2516 -772
rect 2518 -782 2671 -772
rect 2679 -782 2709 -772
rect 2713 -782 2743 -768
rect 2771 -782 2784 -744
rect 2856 -738 2891 -730
rect 2856 -764 2857 -738
rect 2864 -764 2891 -738
rect 2799 -782 2829 -768
rect 2856 -772 2891 -764
rect 2893 -738 2934 -730
rect 2893 -764 2908 -738
rect 2915 -764 2934 -738
rect 2998 -742 3060 -730
rect 3072 -742 3147 -730
rect 3205 -742 3280 -730
rect 3292 -742 3323 -730
rect 3329 -742 3364 -730
rect 2998 -744 3160 -742
rect 2893 -772 2934 -764
rect 3016 -768 3029 -744
rect 3044 -746 3059 -744
rect 2856 -782 2857 -772
rect 2872 -782 2885 -772
rect 2899 -782 2900 -772
rect 2915 -782 2928 -772
rect 2943 -782 2973 -768
rect 3016 -782 3059 -768
rect 3083 -771 3090 -764
rect 3093 -768 3160 -744
rect 3192 -744 3364 -742
rect 3162 -766 3190 -762
rect 3192 -766 3272 -744
rect 3293 -746 3308 -744
rect 3162 -768 3272 -766
rect 3093 -772 3272 -768
rect 3066 -782 3096 -772
rect 3098 -782 3251 -772
rect 3259 -782 3289 -772
rect 3293 -782 3323 -768
rect 3351 -782 3364 -744
rect 3436 -738 3471 -730
rect 3436 -764 3437 -738
rect 3444 -764 3471 -738
rect 3379 -782 3409 -768
rect 3436 -772 3471 -764
rect 3473 -738 3514 -730
rect 3473 -764 3488 -738
rect 3495 -764 3514 -738
rect 3578 -742 3640 -730
rect 3652 -742 3727 -730
rect 3785 -742 3860 -730
rect 3872 -742 3903 -730
rect 3909 -742 3944 -730
rect 3578 -744 3740 -742
rect 3473 -772 3514 -764
rect 3596 -768 3609 -744
rect 3624 -746 3639 -744
rect 3436 -782 3437 -772
rect 3452 -782 3465 -772
rect 3479 -782 3480 -772
rect 3495 -782 3508 -772
rect 3523 -782 3553 -768
rect 3596 -782 3639 -768
rect 3663 -771 3670 -764
rect 3673 -768 3740 -744
rect 3772 -744 3944 -742
rect 3742 -766 3770 -762
rect 3772 -766 3852 -744
rect 3873 -746 3888 -744
rect 3742 -768 3852 -766
rect 3673 -772 3852 -768
rect 3646 -782 3676 -772
rect 3678 -782 3831 -772
rect 3839 -782 3869 -772
rect 3873 -782 3903 -768
rect 3931 -782 3944 -744
rect 4016 -738 4051 -730
rect 4016 -764 4017 -738
rect 4024 -764 4051 -738
rect 3959 -782 3989 -768
rect 4016 -772 4051 -764
rect 4053 -738 4094 -730
rect 4053 -764 4068 -738
rect 4075 -764 4094 -738
rect 4158 -742 4220 -730
rect 4232 -742 4307 -730
rect 4365 -742 4440 -730
rect 4452 -742 4483 -730
rect 4489 -742 4524 -730
rect 4158 -744 4320 -742
rect 4053 -772 4094 -764
rect 4176 -768 4189 -744
rect 4204 -746 4219 -744
rect 4016 -782 4017 -772
rect 4032 -782 4045 -772
rect 4059 -782 4060 -772
rect 4075 -782 4088 -772
rect 4103 -782 4133 -768
rect 4176 -782 4219 -768
rect 4243 -771 4250 -764
rect 4253 -768 4320 -744
rect 4352 -744 4524 -742
rect 4322 -766 4350 -762
rect 4352 -766 4432 -744
rect 4453 -746 4468 -744
rect 4322 -768 4432 -766
rect 4253 -772 4432 -768
rect 4226 -782 4256 -772
rect 4258 -782 4411 -772
rect 4419 -782 4449 -772
rect 4453 -782 4483 -768
rect 4511 -782 4524 -744
rect 4596 -738 4631 -730
rect 4596 -764 4597 -738
rect 4604 -764 4631 -738
rect 4539 -782 4569 -768
rect 4596 -772 4631 -764
rect 4596 -782 4597 -772
rect 4612 -782 4625 -772
rect -1 -788 4625 -782
rect 0 -796 4625 -788
rect 15 -826 28 -796
rect 43 -814 73 -796
rect 116 -810 130 -796
rect 166 -810 386 -796
rect 117 -812 130 -810
rect 83 -824 98 -812
rect 80 -826 102 -824
rect 107 -826 137 -812
rect 198 -814 351 -810
rect 180 -826 372 -814
rect 415 -826 445 -812
rect 451 -826 464 -796
rect 479 -814 509 -796
rect 552 -826 565 -796
rect 595 -826 608 -796
rect 623 -814 653 -796
rect 696 -810 710 -796
rect 746 -810 966 -796
rect 697 -812 710 -810
rect 663 -824 678 -812
rect 660 -826 682 -824
rect 687 -826 717 -812
rect 778 -814 931 -810
rect 760 -826 952 -814
rect 995 -826 1025 -812
rect 1031 -826 1044 -796
rect 1059 -814 1089 -796
rect 1132 -826 1145 -796
rect 1175 -826 1188 -796
rect 1203 -814 1233 -796
rect 1276 -810 1290 -796
rect 1326 -810 1546 -796
rect 1277 -812 1290 -810
rect 1243 -824 1258 -812
rect 1240 -826 1262 -824
rect 1267 -826 1297 -812
rect 1358 -814 1511 -810
rect 1340 -826 1532 -814
rect 1575 -826 1605 -812
rect 1611 -826 1624 -796
rect 1639 -814 1669 -796
rect 1712 -826 1725 -796
rect 1755 -826 1768 -796
rect 1783 -814 1813 -796
rect 1856 -810 1870 -796
rect 1906 -810 2126 -796
rect 1857 -812 1870 -810
rect 1823 -824 1838 -812
rect 1820 -826 1842 -824
rect 1847 -826 1877 -812
rect 1938 -814 2091 -810
rect 1920 -826 2112 -814
rect 2155 -826 2185 -812
rect 2191 -826 2204 -796
rect 2219 -814 2249 -796
rect 2292 -826 2305 -796
rect 2335 -826 2348 -796
rect 2363 -814 2393 -796
rect 2436 -810 2450 -796
rect 2486 -810 2706 -796
rect 2437 -812 2450 -810
rect 2403 -824 2418 -812
rect 2400 -826 2422 -824
rect 2427 -826 2457 -812
rect 2518 -814 2671 -810
rect 2500 -826 2692 -814
rect 2735 -826 2765 -812
rect 2771 -826 2784 -796
rect 2799 -814 2829 -796
rect 2872 -826 2885 -796
rect 2915 -826 2928 -796
rect 2943 -814 2973 -796
rect 3016 -810 3030 -796
rect 3066 -810 3286 -796
rect 3017 -812 3030 -810
rect 2983 -824 2998 -812
rect 2980 -826 3002 -824
rect 3007 -826 3037 -812
rect 3098 -814 3251 -810
rect 3080 -826 3272 -814
rect 3315 -826 3345 -812
rect 3351 -826 3364 -796
rect 3379 -814 3409 -796
rect 3452 -826 3465 -796
rect 3495 -826 3508 -796
rect 3523 -814 3553 -796
rect 3596 -810 3610 -796
rect 3646 -810 3866 -796
rect 3597 -812 3610 -810
rect 3563 -824 3578 -812
rect 3560 -826 3582 -824
rect 3587 -826 3617 -812
rect 3678 -814 3831 -810
rect 3660 -826 3852 -814
rect 3895 -826 3925 -812
rect 3931 -826 3944 -796
rect 3959 -814 3989 -796
rect 4032 -826 4045 -796
rect 4075 -826 4088 -796
rect 4103 -814 4133 -796
rect 4176 -810 4190 -796
rect 4226 -810 4446 -796
rect 4177 -812 4190 -810
rect 4143 -824 4158 -812
rect 4140 -826 4162 -824
rect 4167 -826 4197 -812
rect 4258 -814 4411 -810
rect 4240 -826 4432 -814
rect 4475 -826 4505 -812
rect 4511 -826 4524 -796
rect 4539 -814 4569 -796
rect 4612 -826 4625 -796
rect 0 -840 4625 -826
rect 15 -944 28 -840
rect 73 -862 74 -852
rect 89 -862 102 -852
rect 73 -866 102 -862
rect 107 -866 137 -840
rect 155 -854 171 -852
rect 243 -854 296 -840
rect 244 -856 308 -854
rect 155 -866 170 -862
rect 73 -868 170 -866
rect 57 -876 108 -868
rect 57 -888 82 -876
rect 89 -888 108 -876
rect 139 -876 189 -868
rect 139 -884 155 -876
rect 162 -878 189 -876
rect 198 -876 213 -872
rect 260 -876 292 -856
rect 351 -868 366 -840
rect 415 -843 445 -840
rect 415 -846 451 -843
rect 381 -854 397 -852
rect 382 -866 397 -862
rect 415 -865 454 -846
rect 473 -852 480 -851
rect 479 -859 480 -852
rect 463 -862 464 -859
rect 479 -862 492 -859
rect 415 -866 445 -865
rect 454 -866 460 -865
rect 463 -866 492 -862
rect 382 -867 492 -866
rect 382 -868 498 -867
rect 351 -876 419 -868
rect 198 -878 267 -876
rect 285 -878 419 -876
rect 162 -882 234 -878
rect 162 -884 287 -882
rect 162 -888 234 -884
rect 57 -896 108 -888
rect 155 -892 234 -888
rect 315 -892 419 -878
rect 448 -876 498 -868
rect 448 -885 464 -876
rect 155 -896 419 -892
rect 445 -888 464 -885
rect 471 -888 498 -876
rect 445 -896 498 -888
rect 73 -904 74 -896
rect 89 -904 102 -896
rect 73 -912 89 -904
rect 70 -919 89 -916
rect 70 -928 92 -919
rect 43 -938 92 -928
rect 43 -944 73 -938
rect 92 -943 97 -938
rect 15 -960 89 -944
rect 107 -952 137 -896
rect 172 -906 380 -896
rect 415 -900 460 -896
rect 463 -897 464 -896
rect 479 -897 492 -896
rect 339 -910 387 -906
rect 222 -932 252 -923
rect 315 -930 330 -923
rect 351 -932 387 -910
rect 198 -936 387 -932
rect 213 -939 387 -936
rect 206 -942 387 -939
rect 15 -962 28 -960
rect 43 -962 77 -960
rect 15 -978 89 -962
rect 116 -966 129 -952
rect 144 -966 160 -950
rect 206 -955 217 -942
rect -1 -1000 0 -984
rect 15 -1000 28 -978
rect 43 -1000 73 -978
rect 116 -982 178 -966
rect 206 -973 217 -957
rect 222 -962 232 -942
rect 242 -962 256 -942
rect 259 -955 268 -942
rect 284 -955 293 -942
rect 222 -973 256 -962
rect 259 -973 267 -957
rect 284 -973 293 -957
rect 300 -962 310 -942
rect 320 -962 334 -942
rect 335 -955 346 -942
rect 300 -973 334 -962
rect 335 -973 346 -957
rect 392 -966 408 -950
rect 415 -952 445 -900
rect 479 -904 480 -897
rect 464 -912 480 -904
rect 451 -944 464 -925
rect 479 -944 509 -928
rect 451 -960 525 -944
rect 451 -962 464 -960
rect 479 -962 513 -960
rect 116 -984 129 -982
rect 144 -984 178 -982
rect 116 -1000 178 -984
rect 222 -989 235 -986
rect 300 -989 330 -978
rect 378 -982 424 -966
rect 451 -978 525 -962
rect 378 -984 412 -982
rect 377 -1000 424 -984
rect 451 -1000 464 -978
rect 479 -1000 509 -978
rect 536 -1000 537 -984
rect 552 -1000 565 -840
rect 595 -944 608 -840
rect 653 -862 654 -852
rect 669 -862 682 -852
rect 653 -866 682 -862
rect 687 -866 717 -840
rect 735 -854 751 -852
rect 823 -854 876 -840
rect 824 -856 888 -854
rect 735 -866 750 -862
rect 653 -868 750 -866
rect 637 -876 688 -868
rect 637 -888 662 -876
rect 669 -888 688 -876
rect 719 -876 769 -868
rect 719 -884 735 -876
rect 742 -878 769 -876
rect 778 -876 793 -872
rect 840 -876 872 -856
rect 931 -868 946 -840
rect 995 -843 1025 -840
rect 995 -846 1031 -843
rect 961 -854 977 -852
rect 962 -866 977 -862
rect 995 -865 1034 -846
rect 1053 -852 1060 -851
rect 1059 -859 1060 -852
rect 1043 -862 1044 -859
rect 1059 -862 1072 -859
rect 995 -866 1025 -865
rect 1034 -866 1040 -865
rect 1043 -866 1072 -862
rect 962 -867 1072 -866
rect 962 -868 1078 -867
rect 931 -876 999 -868
rect 778 -878 847 -876
rect 865 -878 999 -876
rect 742 -882 814 -878
rect 742 -884 867 -882
rect 742 -888 814 -884
rect 637 -896 688 -888
rect 735 -892 814 -888
rect 895 -892 999 -878
rect 1028 -876 1078 -868
rect 1028 -885 1044 -876
rect 735 -896 999 -892
rect 1025 -888 1044 -885
rect 1051 -888 1078 -876
rect 1025 -896 1078 -888
rect 653 -904 654 -896
rect 669 -904 682 -896
rect 653 -912 669 -904
rect 650 -919 669 -916
rect 650 -928 672 -919
rect 623 -938 672 -928
rect 623 -944 653 -938
rect 672 -943 677 -938
rect 595 -960 669 -944
rect 687 -952 717 -896
rect 752 -906 960 -896
rect 995 -900 1040 -896
rect 1043 -897 1044 -896
rect 1059 -897 1072 -896
rect 919 -910 967 -906
rect 802 -932 832 -923
rect 895 -930 910 -923
rect 931 -932 967 -910
rect 778 -936 967 -932
rect 793 -939 967 -936
rect 786 -942 967 -939
rect 595 -962 608 -960
rect 623 -962 657 -960
rect 595 -978 669 -962
rect 696 -966 709 -952
rect 724 -966 740 -950
rect 786 -955 797 -942
rect 579 -1000 580 -984
rect 595 -1000 608 -978
rect 623 -1000 653 -978
rect 696 -982 758 -966
rect 786 -973 797 -957
rect 802 -962 812 -942
rect 822 -962 836 -942
rect 839 -955 848 -942
rect 864 -955 873 -942
rect 802 -973 836 -962
rect 839 -973 847 -957
rect 864 -973 873 -957
rect 880 -962 890 -942
rect 900 -962 914 -942
rect 915 -955 926 -942
rect 880 -973 914 -962
rect 915 -973 926 -957
rect 972 -966 988 -950
rect 995 -952 1025 -900
rect 1059 -904 1060 -897
rect 1044 -912 1060 -904
rect 1031 -944 1044 -925
rect 1059 -944 1089 -928
rect 1031 -960 1105 -944
rect 1031 -962 1044 -960
rect 1059 -962 1093 -960
rect 696 -984 709 -982
rect 724 -984 758 -982
rect 696 -1000 758 -984
rect 802 -989 815 -986
rect 880 -989 910 -978
rect 958 -982 1004 -966
rect 1031 -978 1105 -962
rect 958 -984 992 -982
rect 957 -1000 1004 -984
rect 1031 -1000 1044 -978
rect 1059 -1000 1089 -978
rect 1116 -1000 1117 -984
rect 1132 -1000 1145 -840
rect 1175 -944 1188 -840
rect 1233 -862 1234 -852
rect 1249 -862 1262 -852
rect 1233 -866 1262 -862
rect 1267 -866 1297 -840
rect 1315 -854 1331 -852
rect 1403 -854 1456 -840
rect 1404 -856 1468 -854
rect 1315 -866 1330 -862
rect 1233 -868 1330 -866
rect 1217 -876 1268 -868
rect 1217 -888 1242 -876
rect 1249 -888 1268 -876
rect 1299 -876 1349 -868
rect 1299 -884 1315 -876
rect 1322 -878 1349 -876
rect 1358 -876 1373 -872
rect 1420 -876 1452 -856
rect 1511 -868 1526 -840
rect 1575 -843 1605 -840
rect 1575 -846 1611 -843
rect 1541 -854 1557 -852
rect 1542 -866 1557 -862
rect 1575 -865 1614 -846
rect 1633 -852 1640 -851
rect 1639 -859 1640 -852
rect 1623 -862 1624 -859
rect 1639 -862 1652 -859
rect 1575 -866 1605 -865
rect 1614 -866 1620 -865
rect 1623 -866 1652 -862
rect 1542 -867 1652 -866
rect 1542 -868 1658 -867
rect 1511 -876 1579 -868
rect 1358 -878 1427 -876
rect 1445 -878 1579 -876
rect 1322 -882 1394 -878
rect 1322 -884 1447 -882
rect 1322 -888 1394 -884
rect 1217 -896 1268 -888
rect 1315 -892 1394 -888
rect 1475 -892 1579 -878
rect 1608 -876 1658 -868
rect 1608 -885 1624 -876
rect 1315 -896 1579 -892
rect 1605 -888 1624 -885
rect 1631 -888 1658 -876
rect 1605 -896 1658 -888
rect 1233 -904 1234 -896
rect 1249 -904 1262 -896
rect 1233 -912 1249 -904
rect 1230 -919 1249 -916
rect 1230 -928 1252 -919
rect 1203 -938 1252 -928
rect 1203 -944 1233 -938
rect 1252 -943 1257 -938
rect 1175 -960 1249 -944
rect 1267 -952 1297 -896
rect 1332 -906 1540 -896
rect 1575 -900 1620 -896
rect 1623 -897 1624 -896
rect 1639 -897 1652 -896
rect 1499 -910 1547 -906
rect 1382 -932 1412 -923
rect 1475 -930 1490 -923
rect 1511 -932 1547 -910
rect 1358 -936 1547 -932
rect 1373 -939 1547 -936
rect 1366 -942 1547 -939
rect 1175 -962 1188 -960
rect 1203 -962 1237 -960
rect 1175 -978 1249 -962
rect 1276 -966 1289 -952
rect 1304 -966 1320 -950
rect 1366 -955 1377 -942
rect 1159 -1000 1160 -984
rect 1175 -1000 1188 -978
rect 1203 -1000 1233 -978
rect 1276 -982 1338 -966
rect 1366 -973 1377 -957
rect 1382 -962 1392 -942
rect 1402 -962 1416 -942
rect 1419 -955 1428 -942
rect 1444 -955 1453 -942
rect 1382 -973 1416 -962
rect 1419 -973 1427 -957
rect 1444 -973 1453 -957
rect 1460 -962 1470 -942
rect 1480 -962 1494 -942
rect 1495 -955 1506 -942
rect 1460 -973 1494 -962
rect 1495 -973 1506 -957
rect 1552 -966 1568 -950
rect 1575 -952 1605 -900
rect 1639 -904 1640 -897
rect 1624 -912 1640 -904
rect 1611 -944 1624 -925
rect 1639 -944 1669 -928
rect 1611 -960 1685 -944
rect 1611 -962 1624 -960
rect 1639 -962 1673 -960
rect 1276 -984 1289 -982
rect 1304 -984 1338 -982
rect 1276 -1000 1338 -984
rect 1382 -989 1395 -986
rect 1460 -989 1490 -978
rect 1538 -982 1584 -966
rect 1611 -978 1685 -962
rect 1538 -984 1572 -982
rect 1537 -1000 1584 -984
rect 1611 -1000 1624 -978
rect 1639 -1000 1669 -978
rect 1696 -1000 1697 -984
rect 1712 -1000 1725 -840
rect 1755 -944 1768 -840
rect 1813 -862 1814 -852
rect 1829 -862 1842 -852
rect 1813 -866 1842 -862
rect 1847 -866 1877 -840
rect 1895 -854 1911 -852
rect 1983 -854 2036 -840
rect 1984 -856 2048 -854
rect 1895 -866 1910 -862
rect 1813 -868 1910 -866
rect 1797 -876 1848 -868
rect 1797 -888 1822 -876
rect 1829 -888 1848 -876
rect 1879 -876 1929 -868
rect 1879 -884 1895 -876
rect 1902 -878 1929 -876
rect 1938 -876 1953 -872
rect 2000 -876 2032 -856
rect 2091 -868 2106 -840
rect 2155 -843 2185 -840
rect 2155 -846 2191 -843
rect 2121 -854 2137 -852
rect 2122 -866 2137 -862
rect 2155 -865 2194 -846
rect 2213 -852 2220 -851
rect 2219 -859 2220 -852
rect 2203 -862 2204 -859
rect 2219 -862 2232 -859
rect 2155 -866 2185 -865
rect 2194 -866 2200 -865
rect 2203 -866 2232 -862
rect 2122 -867 2232 -866
rect 2122 -868 2238 -867
rect 2091 -876 2159 -868
rect 1938 -878 2007 -876
rect 2025 -878 2159 -876
rect 1902 -882 1974 -878
rect 1902 -884 2027 -882
rect 1902 -888 1974 -884
rect 1797 -896 1848 -888
rect 1895 -892 1974 -888
rect 2055 -892 2159 -878
rect 2188 -876 2238 -868
rect 2188 -885 2204 -876
rect 1895 -896 2159 -892
rect 2185 -888 2204 -885
rect 2211 -888 2238 -876
rect 2185 -896 2238 -888
rect 1813 -904 1814 -896
rect 1829 -904 1842 -896
rect 1813 -912 1829 -904
rect 1810 -919 1829 -916
rect 1810 -928 1832 -919
rect 1783 -938 1832 -928
rect 1783 -944 1813 -938
rect 1832 -943 1837 -938
rect 1755 -960 1829 -944
rect 1847 -952 1877 -896
rect 1912 -906 2120 -896
rect 2155 -900 2200 -896
rect 2203 -897 2204 -896
rect 2219 -897 2232 -896
rect 2079 -910 2127 -906
rect 1962 -932 1992 -923
rect 2055 -930 2070 -923
rect 2091 -932 2127 -910
rect 1938 -936 2127 -932
rect 1953 -939 2127 -936
rect 1946 -942 2127 -939
rect 1755 -962 1768 -960
rect 1783 -962 1817 -960
rect 1755 -978 1829 -962
rect 1856 -966 1869 -952
rect 1884 -966 1900 -950
rect 1946 -955 1957 -942
rect 1739 -1000 1740 -984
rect 1755 -1000 1768 -978
rect 1783 -1000 1813 -978
rect 1856 -982 1918 -966
rect 1946 -973 1957 -957
rect 1962 -962 1972 -942
rect 1982 -962 1996 -942
rect 1999 -955 2008 -942
rect 2024 -955 2033 -942
rect 1962 -973 1996 -962
rect 1999 -973 2007 -957
rect 2024 -973 2033 -957
rect 2040 -962 2050 -942
rect 2060 -962 2074 -942
rect 2075 -955 2086 -942
rect 2040 -973 2074 -962
rect 2075 -973 2086 -957
rect 2132 -966 2148 -950
rect 2155 -952 2185 -900
rect 2219 -904 2220 -897
rect 2204 -912 2220 -904
rect 2191 -944 2204 -925
rect 2219 -944 2249 -928
rect 2191 -960 2265 -944
rect 2191 -962 2204 -960
rect 2219 -962 2253 -960
rect 1856 -984 1869 -982
rect 1884 -984 1918 -982
rect 1856 -1000 1918 -984
rect 1962 -989 1975 -986
rect 2040 -989 2070 -978
rect 2118 -982 2164 -966
rect 2191 -978 2265 -962
rect 2118 -984 2152 -982
rect 2117 -1000 2164 -984
rect 2191 -1000 2204 -978
rect 2219 -1000 2249 -978
rect 2276 -1000 2277 -984
rect 2292 -1000 2305 -840
rect 2335 -944 2348 -840
rect 2393 -862 2394 -852
rect 2409 -862 2422 -852
rect 2393 -866 2422 -862
rect 2427 -866 2457 -840
rect 2475 -854 2491 -852
rect 2563 -854 2616 -840
rect 2564 -856 2628 -854
rect 2475 -866 2490 -862
rect 2393 -868 2490 -866
rect 2377 -876 2428 -868
rect 2377 -888 2402 -876
rect 2409 -888 2428 -876
rect 2459 -876 2509 -868
rect 2459 -884 2475 -876
rect 2482 -878 2509 -876
rect 2518 -876 2533 -872
rect 2580 -876 2612 -856
rect 2671 -868 2686 -840
rect 2735 -843 2765 -840
rect 2735 -846 2771 -843
rect 2701 -854 2717 -852
rect 2702 -866 2717 -862
rect 2735 -865 2774 -846
rect 2793 -852 2800 -851
rect 2799 -859 2800 -852
rect 2783 -862 2784 -859
rect 2799 -862 2812 -859
rect 2735 -866 2765 -865
rect 2774 -866 2780 -865
rect 2783 -866 2812 -862
rect 2702 -867 2812 -866
rect 2702 -868 2818 -867
rect 2671 -876 2739 -868
rect 2518 -878 2587 -876
rect 2605 -878 2739 -876
rect 2482 -882 2554 -878
rect 2482 -884 2607 -882
rect 2482 -888 2554 -884
rect 2377 -896 2428 -888
rect 2475 -892 2554 -888
rect 2635 -892 2739 -878
rect 2768 -876 2818 -868
rect 2768 -885 2784 -876
rect 2475 -896 2739 -892
rect 2765 -888 2784 -885
rect 2791 -888 2818 -876
rect 2765 -896 2818 -888
rect 2393 -904 2394 -896
rect 2409 -904 2422 -896
rect 2393 -912 2409 -904
rect 2390 -919 2409 -916
rect 2390 -928 2412 -919
rect 2363 -938 2412 -928
rect 2363 -944 2393 -938
rect 2412 -943 2417 -938
rect 2335 -960 2409 -944
rect 2427 -952 2457 -896
rect 2492 -906 2700 -896
rect 2735 -900 2780 -896
rect 2783 -897 2784 -896
rect 2799 -897 2812 -896
rect 2659 -910 2707 -906
rect 2542 -932 2572 -923
rect 2635 -930 2650 -923
rect 2671 -932 2707 -910
rect 2518 -936 2707 -932
rect 2533 -939 2707 -936
rect 2526 -942 2707 -939
rect 2335 -962 2348 -960
rect 2363 -962 2397 -960
rect 2335 -978 2409 -962
rect 2436 -966 2449 -952
rect 2464 -966 2480 -950
rect 2526 -955 2537 -942
rect 2319 -1000 2320 -984
rect 2335 -1000 2348 -978
rect 2363 -1000 2393 -978
rect 2436 -982 2498 -966
rect 2526 -973 2537 -957
rect 2542 -962 2552 -942
rect 2562 -962 2576 -942
rect 2579 -955 2588 -942
rect 2604 -955 2613 -942
rect 2542 -973 2576 -962
rect 2579 -973 2587 -957
rect 2604 -973 2613 -957
rect 2620 -962 2630 -942
rect 2640 -962 2654 -942
rect 2655 -955 2666 -942
rect 2620 -973 2654 -962
rect 2655 -973 2666 -957
rect 2712 -966 2728 -950
rect 2735 -952 2765 -900
rect 2799 -904 2800 -897
rect 2784 -912 2800 -904
rect 2771 -944 2784 -925
rect 2799 -944 2829 -928
rect 2771 -960 2845 -944
rect 2771 -962 2784 -960
rect 2799 -962 2833 -960
rect 2436 -984 2449 -982
rect 2464 -984 2498 -982
rect 2436 -1000 2498 -984
rect 2542 -989 2555 -986
rect 2620 -989 2650 -978
rect 2698 -982 2744 -966
rect 2771 -978 2845 -962
rect 2698 -984 2732 -982
rect 2697 -1000 2744 -984
rect 2771 -1000 2784 -978
rect 2799 -1000 2829 -978
rect 2856 -1000 2857 -984
rect 2872 -1000 2885 -840
rect 2915 -944 2928 -840
rect 2973 -862 2974 -852
rect 2989 -862 3002 -852
rect 2973 -866 3002 -862
rect 3007 -866 3037 -840
rect 3055 -854 3071 -852
rect 3143 -854 3196 -840
rect 3144 -856 3208 -854
rect 3055 -866 3070 -862
rect 2973 -868 3070 -866
rect 2957 -876 3008 -868
rect 2957 -888 2982 -876
rect 2989 -888 3008 -876
rect 3039 -876 3089 -868
rect 3039 -884 3055 -876
rect 3062 -878 3089 -876
rect 3098 -876 3113 -872
rect 3160 -876 3192 -856
rect 3251 -868 3266 -840
rect 3315 -843 3345 -840
rect 3315 -846 3351 -843
rect 3281 -854 3297 -852
rect 3282 -866 3297 -862
rect 3315 -865 3354 -846
rect 3373 -852 3380 -851
rect 3379 -859 3380 -852
rect 3363 -862 3364 -859
rect 3379 -862 3392 -859
rect 3315 -866 3345 -865
rect 3354 -866 3360 -865
rect 3363 -866 3392 -862
rect 3282 -867 3392 -866
rect 3282 -868 3398 -867
rect 3251 -876 3319 -868
rect 3098 -878 3167 -876
rect 3185 -878 3319 -876
rect 3062 -882 3134 -878
rect 3062 -884 3187 -882
rect 3062 -888 3134 -884
rect 2957 -896 3008 -888
rect 3055 -892 3134 -888
rect 3215 -892 3319 -878
rect 3348 -876 3398 -868
rect 3348 -885 3364 -876
rect 3055 -896 3319 -892
rect 3345 -888 3364 -885
rect 3371 -888 3398 -876
rect 3345 -896 3398 -888
rect 2973 -904 2974 -896
rect 2989 -904 3002 -896
rect 2973 -912 2989 -904
rect 2970 -919 2989 -916
rect 2970 -928 2992 -919
rect 2943 -938 2992 -928
rect 2943 -944 2973 -938
rect 2992 -943 2997 -938
rect 2915 -960 2989 -944
rect 3007 -952 3037 -896
rect 3072 -906 3280 -896
rect 3315 -900 3360 -896
rect 3363 -897 3364 -896
rect 3379 -897 3392 -896
rect 3239 -910 3287 -906
rect 3122 -932 3152 -923
rect 3215 -930 3230 -923
rect 3251 -932 3287 -910
rect 3098 -936 3287 -932
rect 3113 -939 3287 -936
rect 3106 -942 3287 -939
rect 2915 -962 2928 -960
rect 2943 -962 2977 -960
rect 2915 -978 2989 -962
rect 3016 -966 3029 -952
rect 3044 -966 3060 -950
rect 3106 -955 3117 -942
rect 2899 -1000 2900 -984
rect 2915 -1000 2928 -978
rect 2943 -1000 2973 -978
rect 3016 -982 3078 -966
rect 3106 -973 3117 -957
rect 3122 -962 3132 -942
rect 3142 -962 3156 -942
rect 3159 -955 3168 -942
rect 3184 -955 3193 -942
rect 3122 -973 3156 -962
rect 3159 -973 3167 -957
rect 3184 -973 3193 -957
rect 3200 -962 3210 -942
rect 3220 -962 3234 -942
rect 3235 -955 3246 -942
rect 3200 -973 3234 -962
rect 3235 -973 3246 -957
rect 3292 -966 3308 -950
rect 3315 -952 3345 -900
rect 3379 -904 3380 -897
rect 3364 -912 3380 -904
rect 3351 -944 3364 -925
rect 3379 -944 3409 -928
rect 3351 -960 3425 -944
rect 3351 -962 3364 -960
rect 3379 -962 3413 -960
rect 3016 -984 3029 -982
rect 3044 -984 3078 -982
rect 3016 -1000 3078 -984
rect 3122 -989 3135 -986
rect 3200 -989 3230 -978
rect 3278 -982 3324 -966
rect 3351 -978 3425 -962
rect 3278 -984 3312 -982
rect 3277 -1000 3324 -984
rect 3351 -1000 3364 -978
rect 3379 -1000 3409 -978
rect 3436 -1000 3437 -984
rect 3452 -1000 3465 -840
rect 3495 -944 3508 -840
rect 3553 -862 3554 -852
rect 3569 -862 3582 -852
rect 3553 -866 3582 -862
rect 3587 -866 3617 -840
rect 3635 -854 3651 -852
rect 3723 -854 3776 -840
rect 3724 -856 3788 -854
rect 3635 -866 3650 -862
rect 3553 -868 3650 -866
rect 3537 -876 3588 -868
rect 3537 -888 3562 -876
rect 3569 -888 3588 -876
rect 3619 -876 3669 -868
rect 3619 -884 3635 -876
rect 3642 -878 3669 -876
rect 3678 -876 3693 -872
rect 3740 -876 3772 -856
rect 3831 -868 3846 -840
rect 3895 -843 3925 -840
rect 3895 -846 3931 -843
rect 3861 -854 3877 -852
rect 3862 -866 3877 -862
rect 3895 -865 3934 -846
rect 3953 -852 3960 -851
rect 3959 -859 3960 -852
rect 3943 -862 3944 -859
rect 3959 -862 3972 -859
rect 3895 -866 3925 -865
rect 3934 -866 3940 -865
rect 3943 -866 3972 -862
rect 3862 -867 3972 -866
rect 3862 -868 3978 -867
rect 3831 -876 3899 -868
rect 3678 -878 3747 -876
rect 3765 -878 3899 -876
rect 3642 -882 3714 -878
rect 3642 -884 3767 -882
rect 3642 -888 3714 -884
rect 3537 -896 3588 -888
rect 3635 -892 3714 -888
rect 3795 -892 3899 -878
rect 3928 -876 3978 -868
rect 3928 -885 3944 -876
rect 3635 -896 3899 -892
rect 3925 -888 3944 -885
rect 3951 -888 3978 -876
rect 3925 -896 3978 -888
rect 3553 -904 3554 -896
rect 3569 -904 3582 -896
rect 3553 -912 3569 -904
rect 3550 -919 3569 -916
rect 3550 -928 3572 -919
rect 3523 -938 3572 -928
rect 3523 -944 3553 -938
rect 3572 -943 3577 -938
rect 3495 -960 3569 -944
rect 3587 -952 3617 -896
rect 3652 -906 3860 -896
rect 3895 -900 3940 -896
rect 3943 -897 3944 -896
rect 3959 -897 3972 -896
rect 3819 -910 3867 -906
rect 3702 -932 3732 -923
rect 3795 -930 3810 -923
rect 3831 -932 3867 -910
rect 3678 -936 3867 -932
rect 3693 -939 3867 -936
rect 3686 -942 3867 -939
rect 3495 -962 3508 -960
rect 3523 -962 3557 -960
rect 3495 -978 3569 -962
rect 3596 -966 3609 -952
rect 3624 -966 3640 -950
rect 3686 -955 3697 -942
rect 3479 -1000 3480 -984
rect 3495 -1000 3508 -978
rect 3523 -1000 3553 -978
rect 3596 -982 3658 -966
rect 3686 -973 3697 -957
rect 3702 -962 3712 -942
rect 3722 -962 3736 -942
rect 3739 -955 3748 -942
rect 3764 -955 3773 -942
rect 3702 -973 3736 -962
rect 3739 -973 3747 -957
rect 3764 -973 3773 -957
rect 3780 -962 3790 -942
rect 3800 -962 3814 -942
rect 3815 -955 3826 -942
rect 3780 -973 3814 -962
rect 3815 -973 3826 -957
rect 3872 -966 3888 -950
rect 3895 -952 3925 -900
rect 3959 -904 3960 -897
rect 3944 -912 3960 -904
rect 3931 -944 3944 -925
rect 3959 -944 3989 -928
rect 3931 -960 4005 -944
rect 3931 -962 3944 -960
rect 3959 -962 3993 -960
rect 3596 -984 3609 -982
rect 3624 -984 3658 -982
rect 3596 -1000 3658 -984
rect 3702 -989 3715 -986
rect 3780 -989 3810 -978
rect 3858 -982 3904 -966
rect 3931 -978 4005 -962
rect 3858 -984 3892 -982
rect 3857 -1000 3904 -984
rect 3931 -1000 3944 -978
rect 3959 -1000 3989 -978
rect 4016 -1000 4017 -984
rect 4032 -1000 4045 -840
rect 4075 -944 4088 -840
rect 4133 -862 4134 -852
rect 4149 -862 4162 -852
rect 4133 -866 4162 -862
rect 4167 -866 4197 -840
rect 4215 -854 4231 -852
rect 4303 -854 4356 -840
rect 4304 -856 4368 -854
rect 4215 -866 4230 -862
rect 4133 -868 4230 -866
rect 4117 -876 4168 -868
rect 4117 -888 4142 -876
rect 4149 -888 4168 -876
rect 4199 -876 4249 -868
rect 4199 -884 4215 -876
rect 4222 -878 4249 -876
rect 4258 -876 4273 -872
rect 4320 -876 4352 -856
rect 4411 -868 4426 -840
rect 4475 -843 4505 -840
rect 4475 -846 4511 -843
rect 4441 -854 4457 -852
rect 4442 -866 4457 -862
rect 4475 -865 4514 -846
rect 4533 -852 4540 -851
rect 4539 -859 4540 -852
rect 4523 -862 4524 -859
rect 4539 -862 4552 -859
rect 4475 -866 4505 -865
rect 4514 -866 4520 -865
rect 4523 -866 4552 -862
rect 4442 -867 4552 -866
rect 4442 -868 4558 -867
rect 4411 -876 4479 -868
rect 4258 -878 4327 -876
rect 4345 -878 4479 -876
rect 4222 -882 4294 -878
rect 4222 -884 4347 -882
rect 4222 -888 4294 -884
rect 4117 -896 4168 -888
rect 4215 -892 4294 -888
rect 4375 -892 4479 -878
rect 4508 -876 4558 -868
rect 4508 -885 4524 -876
rect 4215 -896 4479 -892
rect 4505 -888 4524 -885
rect 4531 -888 4558 -876
rect 4505 -896 4558 -888
rect 4133 -904 4134 -896
rect 4149 -904 4162 -896
rect 4133 -912 4149 -904
rect 4130 -919 4149 -916
rect 4130 -928 4152 -919
rect 4103 -938 4152 -928
rect 4103 -944 4133 -938
rect 4152 -943 4157 -938
rect 4075 -960 4149 -944
rect 4167 -952 4197 -896
rect 4232 -906 4440 -896
rect 4475 -900 4520 -896
rect 4523 -897 4524 -896
rect 4539 -897 4552 -896
rect 4399 -910 4447 -906
rect 4282 -932 4312 -923
rect 4375 -930 4390 -923
rect 4411 -932 4447 -910
rect 4258 -936 4447 -932
rect 4273 -939 4447 -936
rect 4266 -942 4447 -939
rect 4075 -962 4088 -960
rect 4103 -962 4137 -960
rect 4075 -978 4149 -962
rect 4176 -966 4189 -952
rect 4204 -966 4220 -950
rect 4266 -955 4277 -942
rect 4059 -1000 4060 -984
rect 4075 -1000 4088 -978
rect 4103 -1000 4133 -978
rect 4176 -982 4238 -966
rect 4266 -973 4277 -957
rect 4282 -962 4292 -942
rect 4302 -962 4316 -942
rect 4319 -955 4328 -942
rect 4344 -955 4353 -942
rect 4282 -973 4316 -962
rect 4319 -973 4327 -957
rect 4344 -973 4353 -957
rect 4360 -962 4370 -942
rect 4380 -962 4394 -942
rect 4395 -955 4406 -942
rect 4360 -973 4394 -962
rect 4395 -973 4406 -957
rect 4452 -966 4468 -950
rect 4475 -952 4505 -900
rect 4539 -904 4540 -897
rect 4524 -912 4540 -904
rect 4511 -944 4524 -925
rect 4539 -944 4569 -928
rect 4511 -960 4585 -944
rect 4511 -962 4524 -960
rect 4539 -962 4573 -960
rect 4176 -984 4189 -982
rect 4204 -984 4238 -982
rect 4176 -1000 4238 -984
rect 4282 -989 4295 -986
rect 4360 -989 4390 -978
rect 4438 -982 4484 -966
rect 4511 -978 4585 -962
rect 4438 -984 4472 -982
rect 4437 -1000 4484 -984
rect 4511 -1000 4524 -978
rect 4539 -1000 4569 -978
rect 4596 -1000 4597 -984
rect 4612 -1000 4625 -840
rect -7 -1008 34 -1000
rect -7 -1034 8 -1008
rect 15 -1034 34 -1008
rect 98 -1012 160 -1000
rect 172 -1012 247 -1000
rect 305 -1012 380 -1000
rect 392 -1012 423 -1000
rect 429 -1012 464 -1000
rect 98 -1014 260 -1012
rect -7 -1042 34 -1034
rect 116 -1042 129 -1014
rect 144 -1016 159 -1014
rect 183 -1041 190 -1034
rect 193 -1042 260 -1014
rect 292 -1014 464 -1012
rect 262 -1036 290 -1032
rect 292 -1036 372 -1014
rect 393 -1016 408 -1014
rect 262 -1038 372 -1036
rect 262 -1042 290 -1038
rect 292 -1042 372 -1038
rect -1 -1052 0 -1042
rect 15 -1052 28 -1042
rect 43 -1052 73 -1042
rect 116 -1052 159 -1042
rect 166 -1052 174 -1042
rect 193 -1050 196 -1042
rect 260 -1050 292 -1042
rect 193 -1052 359 -1050
rect 378 -1052 389 -1042
rect 393 -1052 423 -1042
rect 451 -1052 464 -1014
rect 536 -1008 571 -1000
rect 536 -1034 537 -1008
rect 544 -1034 571 -1008
rect 536 -1042 571 -1034
rect 573 -1008 614 -1000
rect 573 -1034 588 -1008
rect 595 -1034 614 -1008
rect 678 -1012 740 -1000
rect 752 -1012 827 -1000
rect 885 -1012 960 -1000
rect 972 -1012 1003 -1000
rect 1009 -1012 1044 -1000
rect 678 -1014 840 -1012
rect 573 -1042 614 -1034
rect 696 -1042 709 -1014
rect 724 -1016 739 -1014
rect 763 -1041 770 -1034
rect 773 -1042 840 -1014
rect 872 -1014 1044 -1012
rect 842 -1036 870 -1032
rect 872 -1036 952 -1014
rect 973 -1016 988 -1014
rect 842 -1038 952 -1036
rect 842 -1042 870 -1038
rect 872 -1042 952 -1038
rect 479 -1052 509 -1042
rect 536 -1052 537 -1042
rect 552 -1052 565 -1042
rect 579 -1052 580 -1042
rect 595 -1052 608 -1042
rect 623 -1052 653 -1042
rect 696 -1052 739 -1042
rect 746 -1052 754 -1042
rect 773 -1050 776 -1042
rect 840 -1050 872 -1042
rect 773 -1052 939 -1050
rect 958 -1052 969 -1042
rect 973 -1052 1003 -1042
rect 1031 -1052 1044 -1014
rect 1116 -1008 1151 -1000
rect 1116 -1034 1117 -1008
rect 1124 -1034 1151 -1008
rect 1116 -1042 1151 -1034
rect 1153 -1008 1194 -1000
rect 1153 -1034 1168 -1008
rect 1175 -1034 1194 -1008
rect 1258 -1012 1320 -1000
rect 1332 -1012 1407 -1000
rect 1465 -1012 1540 -1000
rect 1552 -1012 1583 -1000
rect 1589 -1012 1624 -1000
rect 1258 -1014 1420 -1012
rect 1153 -1042 1194 -1034
rect 1276 -1042 1289 -1014
rect 1304 -1016 1319 -1014
rect 1343 -1041 1350 -1034
rect 1353 -1042 1420 -1014
rect 1452 -1014 1624 -1012
rect 1422 -1036 1450 -1032
rect 1452 -1036 1532 -1014
rect 1553 -1016 1568 -1014
rect 1422 -1038 1532 -1036
rect 1422 -1042 1450 -1038
rect 1452 -1042 1532 -1038
rect 1059 -1052 1089 -1042
rect 1116 -1052 1117 -1042
rect 1132 -1052 1145 -1042
rect 1159 -1052 1160 -1042
rect 1175 -1052 1188 -1042
rect 1203 -1052 1233 -1042
rect 1276 -1052 1319 -1042
rect 1326 -1052 1334 -1042
rect 1353 -1050 1356 -1042
rect 1420 -1050 1452 -1042
rect 1353 -1052 1519 -1050
rect 1538 -1052 1549 -1042
rect 1553 -1052 1583 -1042
rect 1611 -1052 1624 -1014
rect 1696 -1008 1731 -1000
rect 1696 -1034 1697 -1008
rect 1704 -1034 1731 -1008
rect 1696 -1042 1731 -1034
rect 1733 -1008 1774 -1000
rect 1733 -1034 1748 -1008
rect 1755 -1034 1774 -1008
rect 1838 -1012 1900 -1000
rect 1912 -1012 1987 -1000
rect 2045 -1012 2120 -1000
rect 2132 -1012 2163 -1000
rect 2169 -1012 2204 -1000
rect 1838 -1014 2000 -1012
rect 1733 -1042 1774 -1034
rect 1856 -1042 1869 -1014
rect 1884 -1016 1899 -1014
rect 1923 -1041 1930 -1034
rect 1933 -1042 2000 -1014
rect 2032 -1014 2204 -1012
rect 2002 -1036 2030 -1032
rect 2032 -1036 2112 -1014
rect 2133 -1016 2148 -1014
rect 2002 -1038 2112 -1036
rect 2002 -1042 2030 -1038
rect 2032 -1042 2112 -1038
rect 1639 -1052 1669 -1042
rect 1696 -1052 1697 -1042
rect 1712 -1052 1725 -1042
rect 1739 -1052 1740 -1042
rect 1755 -1052 1768 -1042
rect 1783 -1052 1813 -1042
rect 1856 -1052 1899 -1042
rect 1906 -1052 1914 -1042
rect 1933 -1050 1936 -1042
rect 2000 -1050 2032 -1042
rect 1933 -1052 2099 -1050
rect 2118 -1052 2129 -1042
rect 2133 -1052 2163 -1042
rect 2191 -1052 2204 -1014
rect 2276 -1008 2311 -1000
rect 2276 -1034 2277 -1008
rect 2284 -1034 2311 -1008
rect 2276 -1042 2311 -1034
rect 2313 -1008 2354 -1000
rect 2313 -1034 2328 -1008
rect 2335 -1034 2354 -1008
rect 2418 -1012 2480 -1000
rect 2492 -1012 2567 -1000
rect 2625 -1012 2700 -1000
rect 2712 -1012 2743 -1000
rect 2749 -1012 2784 -1000
rect 2418 -1014 2580 -1012
rect 2313 -1042 2354 -1034
rect 2436 -1042 2449 -1014
rect 2464 -1016 2479 -1014
rect 2503 -1041 2510 -1034
rect 2513 -1042 2580 -1014
rect 2612 -1014 2784 -1012
rect 2582 -1036 2610 -1032
rect 2612 -1036 2692 -1014
rect 2713 -1016 2728 -1014
rect 2582 -1038 2692 -1036
rect 2582 -1042 2610 -1038
rect 2612 -1042 2692 -1038
rect 2219 -1052 2249 -1042
rect 2276 -1052 2277 -1042
rect 2292 -1052 2305 -1042
rect 2319 -1052 2320 -1042
rect 2335 -1052 2348 -1042
rect 2363 -1052 2393 -1042
rect 2436 -1052 2479 -1042
rect 2486 -1052 2494 -1042
rect 2513 -1050 2516 -1042
rect 2580 -1050 2612 -1042
rect 2513 -1052 2679 -1050
rect 2698 -1052 2709 -1042
rect 2713 -1052 2743 -1042
rect 2771 -1052 2784 -1014
rect 2856 -1008 2891 -1000
rect 2856 -1034 2857 -1008
rect 2864 -1034 2891 -1008
rect 2856 -1042 2891 -1034
rect 2893 -1008 2934 -1000
rect 2893 -1034 2908 -1008
rect 2915 -1034 2934 -1008
rect 2998 -1012 3060 -1000
rect 3072 -1012 3147 -1000
rect 3205 -1012 3280 -1000
rect 3292 -1012 3323 -1000
rect 3329 -1012 3364 -1000
rect 2998 -1014 3160 -1012
rect 2893 -1042 2934 -1034
rect 3016 -1042 3029 -1014
rect 3044 -1016 3059 -1014
rect 3083 -1041 3090 -1034
rect 3093 -1042 3160 -1014
rect 3192 -1014 3364 -1012
rect 3162 -1036 3190 -1032
rect 3192 -1036 3272 -1014
rect 3293 -1016 3308 -1014
rect 3162 -1038 3272 -1036
rect 3162 -1042 3190 -1038
rect 3192 -1042 3272 -1038
rect 2799 -1052 2829 -1042
rect 2856 -1052 2857 -1042
rect 2872 -1052 2885 -1042
rect 2899 -1052 2900 -1042
rect 2915 -1052 2928 -1042
rect 2943 -1052 2973 -1042
rect 3016 -1052 3059 -1042
rect 3066 -1052 3074 -1042
rect 3093 -1050 3096 -1042
rect 3160 -1050 3192 -1042
rect 3093 -1052 3259 -1050
rect 3278 -1052 3289 -1042
rect 3293 -1052 3323 -1042
rect 3351 -1052 3364 -1014
rect 3436 -1008 3471 -1000
rect 3436 -1034 3437 -1008
rect 3444 -1034 3471 -1008
rect 3436 -1042 3471 -1034
rect 3473 -1008 3514 -1000
rect 3473 -1034 3488 -1008
rect 3495 -1034 3514 -1008
rect 3578 -1012 3640 -1000
rect 3652 -1012 3727 -1000
rect 3785 -1012 3860 -1000
rect 3872 -1012 3903 -1000
rect 3909 -1012 3944 -1000
rect 3578 -1014 3740 -1012
rect 3473 -1042 3514 -1034
rect 3596 -1042 3609 -1014
rect 3624 -1016 3639 -1014
rect 3663 -1041 3670 -1034
rect 3673 -1042 3740 -1014
rect 3772 -1014 3944 -1012
rect 3742 -1036 3770 -1032
rect 3772 -1036 3852 -1014
rect 3873 -1016 3888 -1014
rect 3742 -1038 3852 -1036
rect 3742 -1042 3770 -1038
rect 3772 -1042 3852 -1038
rect 3379 -1052 3409 -1042
rect 3436 -1052 3437 -1042
rect 3452 -1052 3465 -1042
rect 3479 -1052 3480 -1042
rect 3495 -1052 3508 -1042
rect 3523 -1052 3553 -1042
rect 3596 -1052 3639 -1042
rect 3646 -1052 3654 -1042
rect 3673 -1050 3676 -1042
rect 3740 -1050 3772 -1042
rect 3673 -1052 3839 -1050
rect 3858 -1052 3869 -1042
rect 3873 -1052 3903 -1042
rect 3931 -1052 3944 -1014
rect 4016 -1008 4051 -1000
rect 4016 -1034 4017 -1008
rect 4024 -1034 4051 -1008
rect 4016 -1042 4051 -1034
rect 4053 -1008 4094 -1000
rect 4053 -1034 4068 -1008
rect 4075 -1034 4094 -1008
rect 4158 -1012 4220 -1000
rect 4232 -1012 4307 -1000
rect 4365 -1012 4440 -1000
rect 4452 -1012 4483 -1000
rect 4489 -1012 4524 -1000
rect 4158 -1014 4320 -1012
rect 4053 -1042 4094 -1034
rect 4176 -1042 4189 -1014
rect 4204 -1016 4219 -1014
rect 4243 -1041 4250 -1034
rect 4253 -1042 4320 -1014
rect 4352 -1014 4524 -1012
rect 4322 -1036 4350 -1032
rect 4352 -1036 4432 -1014
rect 4453 -1016 4468 -1014
rect 4322 -1038 4432 -1036
rect 4322 -1042 4350 -1038
rect 4352 -1042 4432 -1038
rect 3959 -1052 3989 -1042
rect 4016 -1052 4017 -1042
rect 4032 -1052 4045 -1042
rect 4059 -1052 4060 -1042
rect 4075 -1052 4088 -1042
rect 4103 -1052 4133 -1042
rect 4176 -1052 4219 -1042
rect 4226 -1052 4234 -1042
rect 4253 -1050 4256 -1042
rect 4320 -1050 4352 -1042
rect 4253 -1052 4419 -1050
rect 4438 -1052 4449 -1042
rect 4453 -1052 4483 -1042
rect 4511 -1052 4524 -1014
rect 4596 -1008 4631 -1000
rect 4596 -1034 4597 -1008
rect 4604 -1034 4631 -1008
rect 4596 -1042 4631 -1034
rect 4539 -1052 4569 -1042
rect 4596 -1052 4597 -1042
rect 4612 -1052 4625 -1042
rect -1 -1058 4625 -1052
rect 0 -1066 4625 -1058
rect 15 -1080 28 -1066
rect 43 -1084 73 -1066
rect 116 -1080 129 -1066
rect 166 -1079 174 -1066
rect 207 -1079 345 -1066
rect 378 -1079 386 -1066
rect 243 -1080 294 -1079
rect 451 -1080 464 -1066
rect 244 -1082 308 -1080
rect 479 -1084 509 -1066
rect 552 -1080 565 -1066
rect 595 -1080 608 -1066
rect 623 -1084 653 -1066
rect 696 -1080 709 -1066
rect 746 -1079 754 -1066
rect 787 -1079 925 -1066
rect 958 -1079 966 -1066
rect 823 -1080 874 -1079
rect 1031 -1080 1044 -1066
rect 824 -1082 888 -1080
rect 1059 -1084 1089 -1066
rect 1132 -1080 1145 -1066
rect 1175 -1080 1188 -1066
rect 1203 -1084 1233 -1066
rect 1276 -1080 1289 -1066
rect 1326 -1079 1334 -1066
rect 1367 -1079 1505 -1066
rect 1538 -1079 1546 -1066
rect 1403 -1080 1454 -1079
rect 1611 -1080 1624 -1066
rect 1404 -1082 1468 -1080
rect 1639 -1084 1669 -1066
rect 1712 -1080 1725 -1066
rect 1755 -1080 1768 -1066
rect 1783 -1084 1813 -1066
rect 1856 -1080 1869 -1066
rect 1906 -1079 1914 -1066
rect 1947 -1079 2085 -1066
rect 2118 -1079 2126 -1066
rect 1983 -1080 2034 -1079
rect 2191 -1080 2204 -1066
rect 1984 -1082 2048 -1080
rect 2219 -1084 2249 -1066
rect 2292 -1080 2305 -1066
rect 2335 -1080 2348 -1066
rect 2363 -1084 2393 -1066
rect 2436 -1080 2449 -1066
rect 2486 -1079 2494 -1066
rect 2527 -1079 2665 -1066
rect 2698 -1079 2706 -1066
rect 2563 -1080 2614 -1079
rect 2771 -1080 2784 -1066
rect 2564 -1082 2628 -1080
rect 2799 -1084 2829 -1066
rect 2872 -1080 2885 -1066
rect 2915 -1080 2928 -1066
rect 2943 -1084 2973 -1066
rect 3016 -1080 3029 -1066
rect 3066 -1079 3074 -1066
rect 3107 -1079 3245 -1066
rect 3278 -1079 3286 -1066
rect 3143 -1080 3194 -1079
rect 3351 -1080 3364 -1066
rect 3144 -1082 3208 -1080
rect 3379 -1084 3409 -1066
rect 3452 -1080 3465 -1066
rect 3495 -1080 3508 -1066
rect 3523 -1084 3553 -1066
rect 3596 -1080 3609 -1066
rect 3646 -1079 3654 -1066
rect 3687 -1079 3825 -1066
rect 3858 -1079 3866 -1066
rect 3723 -1080 3774 -1079
rect 3931 -1080 3944 -1066
rect 3724 -1082 3788 -1080
rect 3959 -1084 3989 -1066
rect 4032 -1080 4045 -1066
rect 4075 -1080 4088 -1066
rect 4103 -1084 4133 -1066
rect 4176 -1080 4189 -1066
rect 4226 -1079 4234 -1066
rect 4267 -1079 4405 -1066
rect 4438 -1079 4446 -1066
rect 4303 -1080 4354 -1079
rect 4511 -1080 4524 -1066
rect 4304 -1082 4368 -1080
rect 4539 -1084 4569 -1066
rect 4612 -1080 4625 -1066
<< pwell >>
rect 74 -896 89 -868
rect 464 -896 479 -867
rect 0 -1042 15 -1000
rect 537 -1042 552 -1000
rect 580 -1042 595 -1000
<< ndiffc >>
rect 74 -896 89 -868
rect 464 -896 479 -867
rect 654 -896 669 -868
rect 1044 -896 1059 -867
rect 1234 -896 1249 -868
rect 1624 -896 1639 -867
rect 1814 -896 1829 -868
rect 2204 -896 2219 -867
rect 2394 -896 2409 -868
rect 2784 -896 2799 -867
rect 2974 -896 2989 -868
rect 3364 -896 3379 -867
rect 3554 -896 3569 -868
rect 3944 -896 3959 -867
rect 4134 -896 4149 -868
rect 4524 -896 4539 -867
rect 0 -1042 15 -1000
rect 537 -1042 552 -1000
rect 580 -1042 595 -1000
rect 1117 -1042 1132 -1000
rect 1160 -1042 1175 -1000
rect 1697 -1042 1712 -1000
rect 1740 -1042 1755 -1000
rect 2277 -1042 2292 -1000
rect 2320 -1042 2335 -1000
rect 2857 -1042 2872 -1000
rect 2900 -1042 2915 -1000
rect 3437 -1042 3452 -1000
rect 3480 -1042 3495 -1000
rect 4017 -1042 4032 -1000
rect 4060 -1042 4075 -1000
rect 4597 -1042 4612 -1000
<< poly >>
rect 0 1050 30 1080
rect 0 780 30 810
rect 0 510 30 540
rect 0 240 30 270
rect 0 -30 30 0
rect 0 -300 30 -270
rect 0 -570 30 -540
rect 0 -840 30 -810
<< metal1 >>
rect 0 1036 15 1050
rect 0 912 15 946
rect 0 810 15 824
rect 0 766 15 780
rect 0 642 15 676
rect 0 540 15 554
rect 0 496 15 510
rect 0 372 15 406
rect 0 270 15 284
rect 0 226 15 240
rect 0 102 15 136
rect 0 0 15 14
rect 0 -44 15 -30
rect 0 -168 15 -134
rect 0 -270 15 -256
rect 0 -314 15 -300
rect 0 -438 15 -404
rect 0 -540 15 -526
rect 0 -584 15 -570
rect 0 -708 15 -674
rect 0 -810 15 -796
rect 0 -854 15 -840
rect 0 -978 15 -944
rect 0 -1080 15 -1066
use 10T_1x8_magic  10T_1x8_magic_0
timestamp 1667336911
transform 1 0 0 0 1 270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_1
timestamp 1667336911
transform 1 0 0 0 1 0
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_2
timestamp 1667336911
transform 1 0 0 0 1 810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_3
timestamp 1667336911
transform 1 0 0 0 1 540
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_4
timestamp 1667336911
transform 1 0 0 0 1 -1080
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_5
timestamp 1667336911
transform 1 0 0 0 1 -810
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_6
timestamp 1667336911
transform 1 0 0 0 1 -270
box -7 -4 4631 312
use 10T_1x8_magic  10T_1x8_magic_7
timestamp 1667336911
transform 1 0 0 0 1 -540
box -7 -4 4631 312
<< labels >>
rlabel locali 0 -1042 15 -1000 1 RBL1_0
port 1 ns signal output
rlabel locali 537 -1042 552 -1000 1 RBL0_0
port 2 ns signal output
rlabel locali 580 -1042 595 -1000 1 RBL1_1
port 3 ns signal output
rlabel locali 1117 -1042 1132 -1000 1 RBL0_1
port 4 ns signal output
rlabel locali 1160 -1042 1175 -1000 1 RBL1_2
port 5 ns signal output
rlabel locali 1697 -1042 1712 -1000 1 RBL0_2
port 6 ns signal output
rlabel locali 1740 -1042 1755 -1000 1 RBL1_3
port 7 ns signal output
rlabel locali 2277 -1042 2292 -1000 1 RBL0_3
port 8 ns signal output
rlabel locali 2320 -1042 2335 -1000 1 RBL1_4
port 9 ns signal output
rlabel locali 2857 -1042 2872 -1000 1 RBL0_4
port 10 ns signal output
rlabel locali 2900 -1042 2915 -1000 1 RBL1_5
port 11 ns signal output
rlabel locali 3437 -1042 3452 -1000 1 RBL0_5
port 12 ns signal output
rlabel locali 3480 -1042 3495 -1000 1 RBL1_6
port 13 ns signal output
rlabel locali 4017 -1042 4032 -1000 1 RBL0_6
port 14 ns signal output
rlabel locali 4060 -1042 4075 -1000 1 RBL1_7
port 15 ns signal output
rlabel locali 4597 -1042 4612 -1000 1 RBL0_7
port 16 ns signal output
rlabel locali 464 -896 479 -867 1 WBL_0
port 17 ns signal input
rlabel locali 74 -896 89 -868 1 WBLb_0
port 18 ns signal input
rlabel locali 1044 -896 1059 -867 1 WBL_1
port 19 ns signal input
rlabel locali 654 -896 669 -868 1 WBLb_1
port 20 ns signal input
rlabel locali 1624 -896 1639 -867 1 WBL_2
port 21 ns signal input
rlabel locali 1234 -896 1249 -868 1 WBLb_2
port 22 ns signal input
rlabel locali 2204 -896 2219 -867 1 WBL_3
port 23 ns signal input
rlabel locali 1814 -896 1829 -868 1 WBLb_3
port 24 ns signal input
rlabel locali 2784 -896 2799 -867 1 WBL_4
port 25 ns signal input
rlabel locali 2394 -896 2409 -868 1 WBLb_4
port 26 ns signal input
rlabel locali 3364 -896 3379 -867 1 WBL_5
port 27 ns signal input
rlabel locali 2974 -896 2989 -868 1 WBLb_5
port 28 ns signal input
rlabel locali 3944 -896 3959 -867 1 WBL_6
port 29 ns signal input
rlabel locali 3554 -896 3569 -868 1 WBLb_6
port 30 ns signal input
rlabel locali 4524 -896 4539 -867 1 WBL_7
port 31 ns signal input
rlabel locali 4134 -896 4149 -868 1 WBLb_7
port 32 ns signal input
rlabel poly 0 1050 30 1080 1 WWL_0
port 33 ew signal input
rlabel metal1 0 912 15 946 1 RWL_0
port 34 ew signal input
rlabel poly 0 780 30 810 1 WWL_1
port 35 ew signal input
rlabel metal1 0 642 15 676 1 RWL_1
port 36 ew signal input
rlabel poly 0 510 30 540 1 WWL_2
port 37 ew signal input
rlabel metal1 0 372 15 406 1 RWL_2
port 38 ew signal input
rlabel poly 0 240 30 270 1 WWL_3
port 39 ew signal input
rlabel metal1 0 102 15 136 1 RWL_3
port 40 ew signal input
rlabel poly 0 -30 30 0 1 WWL_4
port 41 ew signal input
rlabel metal1 0 -168 15 -134 1 RWL_4
port 42 ew signal input
rlabel poly 0 -300 30 -270 1 WWL_5
port 43 ew signal input
rlabel metal1 0 -438 15 -404 1 RWL_5
port 44 ew signal input
rlabel poly 0 -570 30 -540 1 WWL_6
port 45 ew signal input
rlabel metal1 0 -708 15 -674 1 RWL_6
port 46 ew signal input
rlabel poly 0 -840 30 -810 1 WWL_7
port 47 ew signal input
rlabel metal1 0 -978 15 -944 1 RWL_7
port 48 ew signal input
rlabel metal1 0 1036 15 1050 1 VDD
port 49 ew power bidirectional abutment
rlabel metal1 0 810 15 824 1 GND
port 50 ew ground bidirectional abutment
rlabel metal1 0 496 15 510 1 VDD
rlabel metal1 0 226 15 240 1 VDD
rlabel metal1 0 766 15 780 1 VDD
rlabel metal1 0 -44 15 -30 1 VDD
rlabel metal1 0 -584 15 -570 1 VDD
rlabel metal1 0 -854 15 -840 1 VDD
rlabel metal1 0 -314 15 -300 1 VDD
rlabel metal1 0 0 15 14 1 GND
rlabel metal1 0 270 15 284 1 GND
rlabel metal1 0 540 15 554 1 GND
rlabel metal1 0 -270 15 -256 1 GND
rlabel metal1 0 -1080 15 -1066 1 GND
rlabel metal1 0 -810 15 -796 1 GND
rlabel metal1 0 -540 15 -526 1 GND
<< end >>
