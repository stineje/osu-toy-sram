* SPICE3 file created from sky130_fd_bd_sram__sram_sp_cell.ext - technology: sky130A

** INV 0
Mpu_2 VPWR      right_net left_net   PWELL ppu   l=0.15  w=0.14
Mnp_1 VGND      right_net left_net   VSUBS npd   l=0.15  w=0.21
                                                               
** INV 1                                                       
Mpu_1 right_net left_net  VPWR       PWELL ppu   l=0.15  w=0.14
Mnp_0 right_net left_net  VGND       VSUBS npd   l=0.15  w=0.21

** Left side
Mpu_3 left_net  WL1       left_net   PWELL ppu   l=0.095 w=0.07
Mnp_1 left_net  WL1       bit_v      VSUBS npass l=0.15  w=0.14
                                                                
** Right side                                                   
Mpu_0 right_net WL2       right_net  PWELL ppu   l=0.095 w=0.07
Mnp_0 bit_b_v   WL2       right_net  VSUBS npass l=0.15  w=0.14

