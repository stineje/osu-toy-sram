* SPICE3 file created from sky130_fd_bd_sram__sram_sp_cell.ext - technology: sky130A

M1000 a_16_104# a_16_182# a_0_142# w_n26_116# npd w=0.21u l=0.15u
+  ad=0.0425p pd=0.92u as=0.0808p ps=1.28u
M1001 a_16_104# a_16_182# a_174_134# w_144_0# ppu w=0.14u l=0.15u
+  ad=0.035p pd=0.78u as=0.064p ps=1.14u
M1002 a_38_292# a_16_262# a_16_104# w_n26_116# npass w=0.14u l=0.15u
+  ad=0.0168p pd=0.52u as=0p ps=0u
M1003 a_174_134# a_16_104# a_16_182# w_144_0# ppu w=0.14u l=0.15u
+  ad=0p pd=0u as=0.0332p ps=0.72u
M1004 a_0_142# a_16_104# a_16_182# w_n26_116# npd w=0.21u l=0.15u
+  ad=0p pd=0u as=0.04375p ps=0.92u
M1005 a_16_104# a_16_262# a_16_104# w_144_0# ppu w=0.07u l=0.095u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_16_182# a_16_24# a_38_0# w_n26_116# npass w=0.14u l=0.15u
+  ad=0p pd=0u as=0.0168p ps=0.52u
M1007 a_16_182# a_16_24# a_16_182# w_144_0# ppu w=0.07u l=0.095u
+  ad=0p pd=0u as=0p ps=0u
