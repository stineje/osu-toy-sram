* FILE: 12T-OSU.sp

********************** begin header *****************************

* SPICE Header file for TSMC 3.3 0.35 process (scn4me_subm)

.OPTIONS post NOMOD probe measout captab 

**################################################
* Only Typical/Typical spice models included
.include '/programs/micromagic/mmi_local/ami05.mod'
**################################################

.param ln_min   =  0.4u
.param lp_min   =  0.4u

.PARAM vddp=3.30	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 25
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "12T-OSU" generated by MMI_SUE5.6.37 on Fri Nov 12 
*+ 13:58:25 CST 2021.

* start main CELL 12T-OSU
* .SUBCKT 12T-OSU BL BR SEL 
M_1 net_2 net_3 BR gnd n W='0.42*1u' L='0.15*1u' 
M_2 net_5 SEL net_2 gnd n W='0.42*1u' L='0.15*1u' 
M_3 net_6 SEL net_1 gnd n W='0.42*1u' L='0.15*1u' 
M_4 BL net_3 net_6 gnd n W='0.42*1u' L='0.15*1u' 
M_5 GND net_1 net_5 gnd n W='0.42*1u' L='0.15*1u' 
M_6 net_1 net_5 GND gnd n W='0.42*1u' L='0.15*1u' 
M_7 net_1 net_5 VDD vdd p W='0.42*1u' L='0.15*1u' 
M_8 VDD net_1 net_5 vdd p W='0.42*1u' L='0.15*1u' 
M_9 net_2 net_3 net_4 gnd n W='0.42*1u' L='0.15*1u' 
M_10 net_7 net_3 net_6 gnd n W='0.42*1u' L='0.15*1u' 
M_11 GND net_5 net_4 gnd n W='0.42*1u' L='0.15*1u' 
M_12 net_7 net_1 GND gnd n W='0.42*1u' L='0.15*1u' 
* .ENDS	$ 12T-OSU

.GLOBAL gnd vdd

.END

